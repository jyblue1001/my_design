* PEX produced on Fri Aug 22 11:19:30 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_19.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_19 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 VDDA.t219 bgr_11_0.1st_Vout_2.t7 bgr_11_0.PFET_GATE_10uA.t9 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1 two_stage_opamp_dummy_magic_26_0.VD1.t18 two_stage_opamp_dummy_magic_26_0.Vb1.t12 two_stage_opamp_dummy_magic_26_0.X.t16 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X2 VOUT-.t19 two_stage_opamp_dummy_magic_26_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 VOUT+.t19 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 two_stage_opamp_dummy_magic_26_0.V_source.t26 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t12 GNDA.t199 GNDA.t198 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X5 VDDA.t408 two_stage_opamp_dummy_magic_26_0.Y.t25 VOUT+.t17 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X6 VOUT-.t20 two_stage_opamp_dummy_magic_26_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X7 two_stage_opamp_dummy_magic_26_0.Y.t5 two_stage_opamp_dummy_magic_26_0.Vb2.t11 two_stage_opamp_dummy_magic_26_0.VD4.t19 two_stage_opamp_dummy_magic_26_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X8 GNDA.t140 GNDA.t138 two_stage_opamp_dummy_magic_26_0.Vb2.t4 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X9 two_stage_opamp_dummy_magic_26_0.X.t1 two_stage_opamp_dummy_magic_26_0.Vb2.t12 two_stage_opamp_dummy_magic_26_0.VD3.t19 two_stage_opamp_dummy_magic_26_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X10 VOUT-.t21 two_stage_opamp_dummy_magic_26_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X11 two_stage_opamp_dummy_magic_26_0.err_amp_mir.t0 GNDA.t136 GNDA.t137 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X12 two_stage_opamp_dummy_magic_26_0.X.t9 two_stage_opamp_dummy_magic_26_0.Vb1.t13 two_stage_opamp_dummy_magic_26_0.VD1.t17 GNDA.t255 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X13 VOUT-.t22 two_stage_opamp_dummy_magic_26_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t10 two_stage_opamp_dummy_magic_26_0.X.t25 GNDA.t189 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X15 VDDA.t52 bgr_11_0.V_TOP.t14 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t4 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X16 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t9 two_stage_opamp_dummy_magic_26_0.X.t26 GNDA.t188 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X17 bgr_11_0.1st_Vout_1.t7 bgr_11_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 VOUT+.t20 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 VOUT-.t23 two_stage_opamp_dummy_magic_26_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X20 two_stage_opamp_dummy_magic_26_0.Vb2.t8 bgr_11_0.NFET_GATE_10uA.t5 GNDA.t229 GNDA.t228 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X21 bgr_11_0.V_TOP.t15 VDDA.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 two_stage_opamp_dummy_magic_26_0.Vb1.t0 GNDA.t134 GNDA.t135 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X23 GNDA.t18 bgr_11_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_26_0.Vb2.t2 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X24 two_stage_opamp_dummy_magic_26_0.Y.t13 two_stage_opamp_dummy_magic_26_0.Vb1.t14 two_stage_opamp_dummy_magic_26_0.VD2.t19 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X25 VOUT-.t24 two_stage_opamp_dummy_magic_26_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X26 bgr_11_0.START_UP_NFET1.t0 bgr_11_0.START_UP_NFET1 GNDA.t8 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X27 bgr_11_0.1st_Vout_1.t1 bgr_11_0.V_mir1.t13 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X28 two_stage_opamp_dummy_magic_26_0.VD2.t3 VIN+.t0 two_stage_opamp_dummy_magic_26_0.V_source.t3 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X29 GNDA.t281 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_26_0.V_source.t25 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X30 two_stage_opamp_dummy_magic_26_0.V_err_mir_p.t3 two_stage_opamp_dummy_magic_26_0.V_err_gate.t6 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X31 VDDA.t374 VDDA.t372 two_stage_opamp_dummy_magic_26_0.VD4.t35 VDDA.t373 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X32 VDDA.t45 two_stage_opamp_dummy_magic_26_0.X.t27 VOUT-.t14 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X33 VOUT-.t25 two_stage_opamp_dummy_magic_26_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 bgr_11_0.V_TOP.t16 VDDA.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 VDDA.t206 two_stage_opamp_dummy_magic_26_0.X.t28 VOUT-.t13 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X36 VOUT+.t21 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t9 two_stage_opamp_dummy_magic_26_0.Y.t26 GNDA.t164 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X38 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t8 two_stage_opamp_dummy_magic_26_0.Y.t27 GNDA.t266 VDDA.t390 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X39 two_stage_opamp_dummy_magic_26_0.Vb2_2.t8 two_stage_opamp_dummy_magic_26_0.Vb2_2.t6 two_stage_opamp_dummy_magic_26_0.Vb2_2.t8 two_stage_opamp_dummy_magic_26_0.Vb2_2.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X40 two_stage_opamp_dummy_magic_26_0.VD3.t17 two_stage_opamp_dummy_magic_26_0.Vb2.t13 two_stage_opamp_dummy_magic_26_0.X.t22 two_stage_opamp_dummy_magic_26_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X41 two_stage_opamp_dummy_magic_26_0.VD3.t37 two_stage_opamp_dummy_magic_26_0.Vb3.t8 VDDA.t411 VDDA.t410 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X42 a_6350_30238.t0 bgr_11_0.Vin+.t1 GNDA.t152 sky130_fd_pr__res_xhigh_po_0p35 l=6
X43 bgr_11_0.V_TOP.t17 VDDA.t188 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 two_stage_opamp_dummy_magic_26_0.V_err_gate.t3 bgr_11_0.NFET_GATE_10uA.t7 GNDA.t233 GNDA.t232 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X45 VOUT+.t22 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X46 VOUT-.t26 two_stage_opamp_dummy_magic_26_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 VOUT-.t27 two_stage_opamp_dummy_magic_26_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 VDDA.t196 a_6540_22450.t11 a_6540_22450.t12 VDDA.t195 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X49 VOUT-.t28 two_stage_opamp_dummy_magic_26_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X50 VOUT-.t29 two_stage_opamp_dummy_magic_26_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 VOUT-.t30 two_stage_opamp_dummy_magic_26_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 VDDA.t204 bgr_11_0.V_mir1.t11 bgr_11_0.V_mir1.t12 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X53 two_stage_opamp_dummy_magic_26_0.Y.t1 two_stage_opamp_dummy_magic_26_0.Vb2.t14 two_stage_opamp_dummy_magic_26_0.VD4.t17 two_stage_opamp_dummy_magic_26_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X54 VOUT+.t23 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 VOUT+.t24 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t14 bgr_11_0.PFET_GATE_10uA.t10 VDDA.t257 VDDA.t256 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X57 VOUT+.t25 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 VDDA.t255 bgr_11_0.PFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t13 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X59 bgr_11_0.V_TOP.t18 VDDA.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 bgr_11_0.cap_res1.t20 bgr_11_0.V_TOP.t12 GNDA.t278 sky130_fd_pr__res_high_po_0p35 l=2.05
X61 VDDA.t39 two_stage_opamp_dummy_magic_26_0.Y.t28 VOUT+.t2 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X62 VDDA.t74 two_stage_opamp_dummy_magic_26_0.Y.t29 VOUT+.t4 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X63 VOUT+.t26 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 GNDA.t236 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t2 VOUT-.t15 GNDA.t235 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X65 VOUT-.t31 two_stage_opamp_dummy_magic_26_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 VOUT-.t32 two_stage_opamp_dummy_magic_26_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 bgr_11_0.V_TOP.t19 VDDA.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_26_0.X.t29 GNDA.t185 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X69 VOUT-.t33 two_stage_opamp_dummy_magic_26_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 VOUT-.t34 two_stage_opamp_dummy_magic_26_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 bgr_11_0.1st_Vout_2.t8 bgr_11_0.cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 VOUT+.t27 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 GNDA.t45 GNDA.t91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X74 VOUT+.t28 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 two_stage_opamp_dummy_magic_26_0.Y.t9 two_stage_opamp_dummy_magic_26_0.Vb2.t15 two_stage_opamp_dummy_magic_26_0.VD4.t15 two_stage_opamp_dummy_magic_26_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X76 two_stage_opamp_dummy_magic_26_0.Y.t11 two_stage_opamp_dummy_magic_26_0.Vb1.t15 two_stage_opamp_dummy_magic_26_0.VD2.t18 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X77 VOUT+.t29 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 VOUT+.t30 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 two_stage_opamp_dummy_magic_26_0.Y.t19 two_stage_opamp_dummy_magic_26_0.Vb1.t16 two_stage_opamp_dummy_magic_26_0.VD2.t17 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X80 VDDA.t138 two_stage_opamp_dummy_magic_26_0.Y.t30 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t9 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X81 VDDA.t217 bgr_11_0.1st_Vout_2.t9 bgr_11_0.PFET_GATE_10uA.t8 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X82 VOUT-.t35 two_stage_opamp_dummy_magic_26_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X83 two_stage_opamp_dummy_magic_26_0.VD2.t9 VIN+.t1 two_stage_opamp_dummy_magic_26_0.V_source.t34 GNDA.t234 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X84 bgr_11_0.1st_Vout_2.t10 bgr_11_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 GNDA.t273 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t14 two_stage_opamp_dummy_magic_26_0.V_source.t24 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X86 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t10 bgr_11_0.PFET_GATE_10uA.t12 VDDA.t253 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X87 two_stage_opamp_dummy_magic_26_0.VD3.t15 two_stage_opamp_dummy_magic_26_0.Vb2.t16 two_stage_opamp_dummy_magic_26_0.X.t8 two_stage_opamp_dummy_magic_26_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X88 VOUT+.t31 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 VOUT-.t36 two_stage_opamp_dummy_magic_26_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 bgr_11_0.Vin+.t0 GNDA.t6 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X91 VDDA.t176 two_stage_opamp_dummy_magic_26_0.X.t30 VOUT-.t12 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X92 VOUT-.t37 two_stage_opamp_dummy_magic_26_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X93 VOUT-.t38 two_stage_opamp_dummy_magic_26_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 VOUT+.t32 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 bgr_11_0.1st_Vout_1.t8 bgr_11_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X96 VOUT-.t39 two_stage_opamp_dummy_magic_26_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X97 VOUT-.t40 two_stage_opamp_dummy_magic_26_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 bgr_11_0.1st_Vout_2.t11 bgr_11_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X99 VOUT-.t41 two_stage_opamp_dummy_magic_26_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 bgr_11_0.V_TOP.t20 VDDA.t414 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t7 two_stage_opamp_dummy_magic_26_0.Y.t31 GNDA.t196 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X102 GNDA.t98 GNDA.t96 GNDA.t98 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X103 VDDA.t251 bgr_11_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t14 VDDA.t250 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X104 VOUT+.t33 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X105 VOUT+.t34 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t16 VDDA.t359 VDDA.t361 VDDA.t360 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X107 VDDA.t69 a_6540_22450.t13 bgr_11_0.1st_Vout_2.t1 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X108 VOUT+.t35 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 VOUT+.t36 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 VOUT-.t42 two_stage_opamp_dummy_magic_26_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 VDDA.t61 bgr_11_0.V_TOP.t21 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t3 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X112 VOUT+.t37 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 VOUT-.t43 two_stage_opamp_dummy_magic_26_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 VDDA.t83 two_stage_opamp_dummy_magic_26_0.X.t31 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t14 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X115 VOUT+.t38 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X116 two_stage_opamp_dummy_magic_26_0.VD3.t13 two_stage_opamp_dummy_magic_26_0.Vb2.t17 two_stage_opamp_dummy_magic_26_0.X.t6 two_stage_opamp_dummy_magic_26_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X117 VOUT-.t44 two_stage_opamp_dummy_magic_26_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 VOUT+.t39 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 VOUT+.t40 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 VDDA.t174 two_stage_opamp_dummy_magic_26_0.Y.t32 VOUT+.t12 VDDA.t173 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X121 VOUT-.t45 two_stage_opamp_dummy_magic_26_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 VOUT-.t46 two_stage_opamp_dummy_magic_26_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 bgr_11_0.1st_Vout_2.t12 bgr_11_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 bgr_11_0.V_TOP.t22 VDDA.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 two_stage_opamp_dummy_magic_26_0.Vb1.t5 two_stage_opamp_dummy_magic_26_0.Vb1.t4 two_stage_opamp_dummy_magic_26_0.Vb1_2.t4 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X126 VOUT+.t41 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 VOUT+.t42 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 VOUT-.t47 two_stage_opamp_dummy_magic_26_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 VOUT+.t43 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t6 VDDA.t369 VDDA.t371 VDDA.t370 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X131 two_stage_opamp_dummy_magic_26_0.VD4.t32 two_stage_opamp_dummy_magic_26_0.Vb3.t9 VDDA.t192 VDDA.t191 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X132 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_26_0.X.t32 GNDA.t186 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X133 two_stage_opamp_dummy_magic_26_0.VD1.t7 VIN-.t0 two_stage_opamp_dummy_magic_26_0.V_source.t29 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X134 two_stage_opamp_dummy_magic_26_0.Y.t18 two_stage_opamp_dummy_magic_26_0.Vb1.t17 two_stage_opamp_dummy_magic_26_0.VD2.t16 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X135 GNDA.t218 bgr_11_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_26_0.Vb3.t6 GNDA.t217 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X136 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t7 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X137 VOUT+.t44 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X138 VDDA.t158 a_6540_22450.t9 a_6540_22450.t10 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X139 VDDA.t147 two_stage_opamp_dummy_magic_26_0.Y.t33 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t8 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X140 bgr_11_0.START_UP.t5 bgr_11_0.V_TOP.t23 VDDA.t194 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X141 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_26_0.Y.t24 GNDA.t289 sky130_fd_pr__res_high_po_1p41 l=1.41
X142 VOUT-.t48 two_stage_opamp_dummy_magic_26_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 VOUT-.t49 two_stage_opamp_dummy_magic_26_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 GNDA.t151 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t15 two_stage_opamp_dummy_magic_26_0.V_p_mir.t2 GNDA.t150 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X145 VOUT-.t50 two_stage_opamp_dummy_magic_26_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 VOUT+.t45 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 two_stage_opamp_dummy_magic_26_0.VD2.t6 GNDA.t132 GNDA.t133 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X148 VOUT+.t46 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 a_11420_30238.t1 bgr_11_0.Vin-.t7 GNDA.t288 sky130_fd_pr__res_xhigh_po_0p35 l=6
X150 bgr_11_0.V_TOP.t10 VDDA.t366 VDDA.t368 VDDA.t367 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X151 GNDA.t272 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_26_0.V_source.t23 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X152 GNDA.t283 a_11950_28880.t0 GNDA.t282 sky130_fd_pr__res_xhigh_po_0p35 l=4
X153 GNDA.t100 GNDA.t99 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t1 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X154 two_stage_opamp_dummy_magic_26_0.VD1.t2 VIN-.t1 two_stage_opamp_dummy_magic_26_0.V_source.t6 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X155 VOUT+.t47 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 a_3810_3908.t0 two_stage_opamp_dummy_magic_26_0.V_tot.t3 GNDA.t200 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X157 VOUT+.t48 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X158 bgr_11_0.V_TOP.t24 VDDA.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 VDDA.t90 two_stage_opamp_dummy_magic_26_0.X.t33 VOUT-.t11 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X160 a_13840_3908.t1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t1 GNDA.t147 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X161 VOUT-.t51 two_stage_opamp_dummy_magic_26_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 VOUT+.t49 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 VDDA.t180 two_stage_opamp_dummy_magic_26_0.Vb3.t10 two_stage_opamp_dummy_magic_26_0.VD3.t34 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X164 VOUT+.t50 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VOUT+.t51 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 bgr_11_0.Vin+.t5 bgr_11_0.V_TOP.t25 VDDA.t150 VDDA.t149 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X167 VOUT+.t52 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 VOUT+.t53 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 VOUT+.t54 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 VDDA.t48 bgr_11_0.V_mir1.t14 bgr_11_0.1st_Vout_1.t2 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X171 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_26_0.Y.t34 GNDA.t11 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X172 two_stage_opamp_dummy_magic_26_0.V_source.t31 two_stage_opamp_dummy_magic_26_0.err_amp_out.t4 GNDA.t221 GNDA.t220 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X173 GNDA.t131 GNDA.t129 VOUT+.t6 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X174 VOUT-.t52 two_stage_opamp_dummy_magic_26_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X175 VOUT+.t55 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 VOUT-.t53 two_stage_opamp_dummy_magic_26_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 bgr_11_0.1st_Vout_2.t13 bgr_11_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 VDDA.t365 VDDA.t362 VDDA.t364 VDDA.t363 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.15
X179 VDDA.t358 VDDA.t355 VDDA.t357 VDDA.t356 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X180 VOUT-.t54 two_stage_opamp_dummy_magic_26_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 VOUT-.t55 two_stage_opamp_dummy_magic_26_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X182 VDDA.t249 bgr_11_0.PFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t9 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X183 VOUT-.t4 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t3 GNDA.t159 GNDA.t158 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X184 VOUT+.t56 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 VDDA.t382 two_stage_opamp_dummy_magic_26_0.X.t34 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t13 GNDA.t184 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X186 VOUT-.t56 two_stage_opamp_dummy_magic_26_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t14 bgr_11_0.NFET_GATE_10uA.t9 GNDA.t161 GNDA.t160 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X188 VDDA.t106 two_stage_opamp_dummy_magic_26_0.X.t35 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t12 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X189 VOUT+.t57 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 VOUT-.t57 two_stage_opamp_dummy_magic_26_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 VOUT+.t58 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X192 two_stage_opamp_dummy_magic_26_0.Vb2.t6 bgr_11_0.NFET_GATE_10uA.t10 GNDA.t213 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X193 VDDA.t8 bgr_11_0.V_TOP.t26 bgr_11_0.Vin-.t6 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X194 VDDA.t354 VDDA.t352 bgr_11_0.V_TOP.t9 VDDA.t353 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X195 VDDA.t146 two_stage_opamp_dummy_magic_26_0.Y.t35 VOUT+.t10 VDDA.t145 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X196 VOUT-.t58 two_stage_opamp_dummy_magic_26_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 GNDA.t45 GNDA.t44 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X198 VOUT+.t59 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 GNDA.t113 GNDA.t111 two_stage_opamp_dummy_magic_26_0.Vb1.t1 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X200 two_stage_opamp_dummy_magic_26_0.err_amp_out.t2 two_stage_opamp_dummy_magic_26_0.err_amp_mir.t5 GNDA.t216 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X201 GNDA.t270 two_stage_opamp_dummy_magic_26_0.Y.t36 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t5 VDDA.t401 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X202 two_stage_opamp_dummy_magic_26_0.VD4.t29 two_stage_opamp_dummy_magic_26_0.VD4.t27 two_stage_opamp_dummy_magic_26_0.Y.t6 two_stage_opamp_dummy_magic_26_0.VD4.t28 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X203 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t6 two_stage_opamp_dummy_magic_26_0.X.t36 GNDA.t182 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X204 bgr_11_0.1st_Vout_1.t9 bgr_11_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 GNDA.t45 GNDA.t128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X206 VDDA.t190 bgr_11_0.1st_Vout_1.t10 bgr_11_0.V_TOP.t5 VDDA.t189 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X207 VOUT-.t59 two_stage_opamp_dummy_magic_26_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 VOUT-.t60 two_stage_opamp_dummy_magic_26_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 VOUT-.t61 two_stage_opamp_dummy_magic_26_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 VOUT+.t0 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t4 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X211 bgr_11_0.START_UP.t1 bgr_11_0.START_UP.t0 bgr_11_0.START_UP_NFET1.t0 GNDA.t256 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X212 two_stage_opamp_dummy_magic_26_0.VD1.t8 VIN-.t2 two_stage_opamp_dummy_magic_26_0.V_source.t30 GNDA.t219 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X213 two_stage_opamp_dummy_magic_26_0.Y.t14 two_stage_opamp_dummy_magic_26_0.Vb1.t18 two_stage_opamp_dummy_magic_26_0.VD2.t15 GNDA.t234 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X214 VOUT-.t62 two_stage_opamp_dummy_magic_26_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X215 VOUT-.t63 two_stage_opamp_dummy_magic_26_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 two_stage_opamp_dummy_magic_26_0.X.t21 two_stage_opamp_dummy_magic_26_0.Vb2.t18 two_stage_opamp_dummy_magic_26_0.VD3.t11 two_stage_opamp_dummy_magic_26_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X217 VDDA.t125 GNDA.t125 GNDA.t127 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X218 VDDA.t417 two_stage_opamp_dummy_magic_26_0.Y.t37 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t7 GNDA.t279 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X219 VOUT+.t60 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 bgr_11_0.NFET_GATE_10uA.t2 bgr_11_0.NFET_GATE_10uA.t1 GNDA.t285 GNDA.t284 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X221 GNDA.t31 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t5 VOUT-.t0 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X222 VOUT-.t64 two_stage_opamp_dummy_magic_26_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 GNDA.t280 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t17 two_stage_opamp_dummy_magic_26_0.V_source.t22 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X224 GNDA.t124 GNDA.t121 GNDA.t123 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X225 VDDA.t183 bgr_11_0.V_TOP.t27 bgr_11_0.Vin+.t4 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X226 bgr_11_0.1st_Vout_1.t11 bgr_11_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 two_stage_opamp_dummy_magic_26_0.err_amp_out.t0 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_26_0.V_err_p.t0 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X228 VOUT+.t9 two_stage_opamp_dummy_magic_26_0.Y.t38 VDDA.t131 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X229 two_stage_opamp_dummy_magic_26_0.VD1.t1 VIN-.t3 two_stage_opamp_dummy_magic_26_0.V_source.t5 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X230 VOUT+.t61 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 VOUT-.t65 two_stage_opamp_dummy_magic_26_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 bgr_11_0.V_TOP.t28 VDDA.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X233 VDDA.t59 two_stage_opamp_dummy_magic_26_0.X.t37 VOUT-.t10 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X234 GNDA.t45 GNDA.t120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X235 a_3690_3908.t1 two_stage_opamp_dummy_magic_26_0.V_tot.t2 GNDA.t149 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X236 VDDA.t202 bgr_11_0.V_mir1.t9 bgr_11_0.V_mir1.t10 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X237 GNDA.t119 GNDA.t116 GNDA.t118 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X238 VDDA.t351 VDDA.t349 bgr_11_0.NFET_GATE_10uA.t4 VDDA.t350 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X239 bgr_11_0.1st_Vout_1.t12 bgr_11_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VOUT+.t62 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 GNDA.t115 GNDA.t114 two_stage_opamp_dummy_magic_26_0.VD1.t5 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X242 VDDA.t110 bgr_11_0.1st_Vout_1.t13 bgr_11_0.V_TOP.t1 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X243 VOUT-.t66 two_stage_opamp_dummy_magic_26_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X244 VOUT-.t67 two_stage_opamp_dummy_magic_26_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X245 VOUT-.t68 two_stage_opamp_dummy_magic_26_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 VOUT+.t63 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 VOUT+.t64 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 VOUT+.t65 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X249 VOUT+.t66 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 bgr_11_0.Vin+.t3 bgr_11_0.V_TOP.t29 VDDA.t119 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X251 two_stage_opamp_dummy_magic_26_0.X.t24 two_stage_opamp_dummy_magic_26_0.Vb2.t19 two_stage_opamp_dummy_magic_26_0.VD3.t9 two_stage_opamp_dummy_magic_26_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X252 GNDA.t110 GNDA.t109 two_stage_opamp_dummy_magic_26_0.VD2.t5 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X253 VDDA.t43 two_stage_opamp_dummy_magic_26_0.X.t38 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t11 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X254 VOUT+.t67 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X255 bgr_11_0.V_TOP.t30 VDDA.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 bgr_11_0.PFET_GATE_10uA.t7 bgr_11_0.1st_Vout_2.t14 VDDA.t215 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X257 two_stage_opamp_dummy_magic_26_0.Vb2.t10 bgr_11_0.NFET_GATE_10uA.t11 GNDA.t258 GNDA.t257 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X258 bgr_11_0.1st_Vout_1.t14 bgr_11_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 VDDA.t82 two_stage_opamp_dummy_magic_26_0.Vb3.t11 two_stage_opamp_dummy_magic_26_0.VD4.t23 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X260 VDDA.t185 bgr_11_0.V_mir1.t7 bgr_11_0.V_mir1.t8 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X261 VOUT-.t69 two_stage_opamp_dummy_magic_26_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 bgr_11_0.V_TOP.t31 VDDA.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 two_stage_opamp_dummy_magic_26_0.X.t14 two_stage_opamp_dummy_magic_26_0.Vb1.t19 two_stage_opamp_dummy_magic_26_0.VD1.t16 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X264 VOUT+.t68 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X265 VOUT-.t70 two_stage_opamp_dummy_magic_26_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X266 VOUT-.t71 two_stage_opamp_dummy_magic_26_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 VDDA.t213 bgr_11_0.1st_Vout_2.t15 bgr_11_0.PFET_GATE_10uA.t6 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X268 two_stage_opamp_dummy_magic_26_0.Vb3.t0 two_stage_opamp_dummy_magic_26_0.Vb2.t20 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X269 VOUT+.t69 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 VOUT+.t70 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X271 two_stage_opamp_dummy_magic_26_0.VD3.t36 VDDA.t346 VDDA.t348 VDDA.t347 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X272 GNDA.t264 a_11300_28630.t1 GNDA.t263 sky130_fd_pr__res_xhigh_po_0p35 l=6
X273 GNDA.t262 bgr_11_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t13 GNDA.t261 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X274 two_stage_opamp_dummy_magic_26_0.Vb2.t3 GNDA.t106 GNDA.t108 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X275 two_stage_opamp_dummy_magic_26_0.Y.t3 GNDA.t103 GNDA.t105 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X276 two_stage_opamp_dummy_magic_26_0.X.t17 two_stage_opamp_dummy_magic_26_0.Vb1.t20 two_stage_opamp_dummy_magic_26_0.VD1.t15 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X277 a_3810_3908.t1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t10 GNDA.t206 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X278 VDDA.t144 two_stage_opamp_dummy_magic_26_0.Y.t39 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t6 GNDA.t208 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X279 bgr_11_0.1st_Vout_2.t16 bgr_11_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X280 bgr_11_0.V_TOP.t32 VDDA.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 two_stage_opamp_dummy_magic_26_0.Vb1_2.t3 two_stage_opamp_dummy_magic_26_0.Vb1.t6 two_stage_opamp_dummy_magic_26_0.Vb1.t7 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X282 a_13960_3908.t1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t0 GNDA.t148 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X283 GNDA.t153 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_26_0.V_source.t21 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X284 two_stage_opamp_dummy_magic_26_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_26_0.V_err_gate.t0 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X285 VDDA.t1 two_stage_opamp_dummy_magic_26_0.V_err_gate.t7 two_stage_opamp_dummy_magic_26_0.V_err_p.t3 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X286 two_stage_opamp_dummy_magic_26_0.VD1.t6 GNDA.t101 GNDA.t102 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X287 VOUT-.t72 two_stage_opamp_dummy_magic_26_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 bgr_11_0.V_p_1.t1 bgr_11_0.Vin+.t6 bgr_11_0.1st_Vout_1.t3 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X289 VDDA.t376 a_6540_22450.t14 bgr_11_0.1st_Vout_2.t5 VDDA.t375 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X290 bgr_11_0.1st_Vout_1.t15 bgr_11_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 VOUT-.t73 two_stage_opamp_dummy_magic_26_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 VOUT+.t71 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 VOUT-.t74 two_stage_opamp_dummy_magic_26_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 VOUT+.t72 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X295 VOUT-.t75 two_stage_opamp_dummy_magic_26_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 VOUT+.t73 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X297 bgr_11_0.1st_Vout_2.t17 bgr_11_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 VOUT+.t74 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 VOUT+.t75 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 GNDA.t95 GNDA.t92 GNDA.t94 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X301 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t1 a_13940_106.t1 GNDA.t204 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X302 GNDA.t90 GNDA.t88 VDDA.t121 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X303 bgr_11_0.1st_Vout_1.t16 bgr_11_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 a_5700_30088.t1 a_5820_28824.t0 GNDA.t27 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X305 VOUT+.t76 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 bgr_11_0.1st_Vout_2.t18 bgr_11_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X307 VDDA.t247 bgr_11_0.PFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t12 VDDA.t246 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X308 VDDA.t200 two_stage_opamp_dummy_magic_26_0.Vb3.t12 two_stage_opamp_dummy_magic_26_0.VD4.t33 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X309 two_stage_opamp_dummy_magic_26_0.V_source.t20 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t19 GNDA.t277 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X310 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t16 VDDA.t343 VDDA.t345 VDDA.t344 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X311 VDDA.t388 two_stage_opamp_dummy_magic_26_0.X.t39 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t10 GNDA.t180 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X312 two_stage_opamp_dummy_magic_26_0.V_source.t19 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t20 GNDA.t271 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X313 two_stage_opamp_dummy_magic_26_0.V_source.t32 VIN+.t2 two_stage_opamp_dummy_magic_26_0.VD2.t7 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X314 VOUT+.t77 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X315 VOUT-.t76 two_stage_opamp_dummy_magic_26_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X316 a_6540_22450.t8 a_6540_22450.t7 VDDA.t163 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X317 bgr_11_0.1st_Vout_1.t17 bgr_11_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 VOUT-.t77 two_stage_opamp_dummy_magic_26_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 bgr_11_0.1st_Vout_2.t19 bgr_11_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 GNDA.t260 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t6 VOUT+.t15 GNDA.t259 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X321 GNDA.t45 GNDA.t47 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X322 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t10 VDDA.t340 VDDA.t342 VDDA.t341 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X323 GNDA.t269 two_stage_opamp_dummy_magic_26_0.Y.t40 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t4 VDDA.t400 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X324 VOUT+.t78 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 VOUT-.t78 two_stage_opamp_dummy_magic_26_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 two_stage_opamp_dummy_magic_26_0.X.t13 two_stage_opamp_dummy_magic_26_0.Vb1.t21 two_stage_opamp_dummy_magic_26_0.VD1.t14 GNDA.t219 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X327 VOUT+.t79 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 two_stage_opamp_dummy_magic_26_0.VD3.t7 two_stage_opamp_dummy_magic_26_0.Vb2.t21 two_stage_opamp_dummy_magic_26_0.X.t5 two_stage_opamp_dummy_magic_26_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X329 bgr_11_0.1st_Vout_2.t20 bgr_11_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 VOUT+.t80 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 VOUT-.t79 two_stage_opamp_dummy_magic_26_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 VOUT-.t80 two_stage_opamp_dummy_magic_26_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 two_stage_opamp_dummy_magic_26_0.X.t15 two_stage_opamp_dummy_magic_26_0.Vb1.t22 two_stage_opamp_dummy_magic_26_0.VD1.t13 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X334 VOUT-.t81 two_stage_opamp_dummy_magic_26_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X335 VOUT-.t82 two_stage_opamp_dummy_magic_26_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X336 VOUT+.t81 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 bgr_11_0.START_UP.t4 bgr_11_0.V_TOP.t33 VDDA.t29 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X338 VOUT+.t82 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 VDDA.t339 VDDA.t337 VDDA.t339 VDDA.t338 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0 ps=0 w=1 l=0.15
X340 VOUT-.t83 two_stage_opamp_dummy_magic_26_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 bgr_11_0.1st_Vout_1.t18 bgr_11_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X342 GNDA.t197 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t21 two_stage_opamp_dummy_magic_26_0.V_source.t18 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X343 VDDA.t378 bgr_11_0.V_mir1.t15 bgr_11_0.1st_Vout_1.t5 VDDA.t377 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X344 VDDA.t245 bgr_11_0.PFET_GATE_10uA.t16 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t8 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X345 VOUT+.t18 two_stage_opamp_dummy_magic_26_0.Y.t41 VDDA.t416 VDDA.t415 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X346 bgr_11_0.cap_res2.t0 bgr_11_0.PFET_GATE_10uA.t1 GNDA.t12 sky130_fd_pr__res_high_po_0p35 l=2.05
X347 two_stage_opamp_dummy_magic_26_0.VD4.t34 VDDA.t334 VDDA.t336 VDDA.t335 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X348 bgr_11_0.V_TOP.t34 VDDA.t379 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X349 VOUT-.t1 a_13940_106.t0 GNDA.t40 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X350 two_stage_opamp_dummy_magic_26_0.VD3.t30 two_stage_opamp_dummy_magic_26_0.Vb3.t13 VDDA.t154 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X351 two_stage_opamp_dummy_magic_26_0.err_amp_mir.t4 VDDA.t331 VDDA.t333 VDDA.t332 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X352 GNDA.t2 two_stage_opamp_dummy_magic_26_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_26_0.err_amp_mir.t2 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X353 VOUT-.t84 two_stage_opamp_dummy_magic_26_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 VOUT-.t85 two_stage_opamp_dummy_magic_26_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 VOUT+.t83 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 VOUT+.t84 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 VOUT+.t85 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X358 VOUT+.t86 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 VOUT+.t5 GNDA.t85 GNDA.t87 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X360 GNDA.t45 GNDA.t84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X361 GNDA.t83 GNDA.t81 two_stage_opamp_dummy_magic_26_0.X.t3 GNDA.t82 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X362 VOUT+.t87 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t0 a_3830_106.t1 GNDA.t142 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X364 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t13 bgr_11_0.PFET_GATE_10uA.t17 VDDA.t243 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X365 GNDA.t178 two_stage_opamp_dummy_magic_26_0.X.t40 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t5 VDDA.t391 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X366 two_stage_opamp_dummy_magic_26_0.VD3.t27 two_stage_opamp_dummy_magic_26_0.VD3.t25 two_stage_opamp_dummy_magic_26_0.X.t23 two_stage_opamp_dummy_magic_26_0.VD3.t26 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X367 VOUT+.t88 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X368 a_6350_30238.t1 a_6470_28630.t1 GNDA.t152 sky130_fd_pr__res_xhigh_po_0p35 l=6
X369 GNDA.t80 GNDA.t79 two_stage_opamp_dummy_magic_26_0.Y.t2 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X370 VOUT-.t86 two_stage_opamp_dummy_magic_26_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X371 VOUT-.t87 two_stage_opamp_dummy_magic_26_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 bgr_11_0.1st_Vout_2.t4 a_6540_22450.t15 VDDA.t198 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X373 VDDA.t165 bgr_11_0.1st_Vout_1.t19 bgr_11_0.V_TOP.t4 VDDA.t164 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X374 VOUT+.t89 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X375 two_stage_opamp_dummy_magic_26_0.V_source.t36 VIN+.t3 two_stage_opamp_dummy_magic_26_0.VD2.t20 GNDA.t253 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X376 VOUT-.t88 two_stage_opamp_dummy_magic_26_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 VDDA.t124 GNDA.t76 GNDA.t78 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X378 two_stage_opamp_dummy_magic_26_0.V_source.t17 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t22 GNDA.t154 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X379 two_stage_opamp_dummy_magic_26_0.V_err_gate.t1 two_stage_opamp_dummy_magic_26_0.V_tot.t4 two_stage_opamp_dummy_magic_26_0.V_err_mir_p.t1 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X380 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t0 GNDA.t74 GNDA.t75 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X381 VOUT+.t90 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 VDDA.t152 bgr_11_0.V_mir1.t16 bgr_11_0.1st_Vout_1.t4 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X383 two_stage_opamp_dummy_magic_26_0.VD4.t20 two_stage_opamp_dummy_magic_26_0.Vb3.t14 VDDA.t26 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X384 VOUT+.t91 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X385 VOUT-.t89 two_stage_opamp_dummy_magic_26_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X386 VOUT-.t90 two_stage_opamp_dummy_magic_26_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 VOUT+.t92 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 VOUT+.t93 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X389 VOUT-.t9 two_stage_opamp_dummy_magic_26_0.X.t41 VDDA.t384 VDDA.t383 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X390 bgr_11_0.V_TOP.t35 VDDA.t380 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_26_0.Vb3.t7 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t4 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X392 GNDA.t195 two_stage_opamp_dummy_magic_26_0.Y.t42 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t3 VDDA.t129 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X393 VOUT+.t94 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 VDDA.t161 two_stage_opamp_dummy_magic_26_0.Vb3.t15 two_stage_opamp_dummy_magic_26_0.VD3.t32 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X395 VOUT-.t91 two_stage_opamp_dummy_magic_26_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X396 GNDA.t73 GNDA.t72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X397 a_12070_30088.t1 a_11950_28880.t1 GNDA.t287 sky130_fd_pr__res_xhigh_po_0p35 l=4
X398 VOUT-.t92 two_stage_opamp_dummy_magic_26_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X399 VDDA.t63 bgr_11_0.V_TOP.t36 bgr_11_0.Vin+.t2 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X400 VOUT-.t93 two_stage_opamp_dummy_magic_26_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 VOUT-.t94 two_stage_opamp_dummy_magic_26_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 GNDA.t71 GNDA.t69 two_stage_opamp_dummy_magic_26_0.Vb3.t1 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X403 two_stage_opamp_dummy_magic_26_0.VD4.t37 two_stage_opamp_dummy_magic_26_0.Vb3.t16 VDDA.t419 VDDA.t418 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X404 VOUT+.t95 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 VOUT+.t96 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X406 two_stage_opamp_dummy_magic_26_0.X.t4 GNDA.t66 GNDA.t68 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X407 bgr_11_0.V_TOP.t0 bgr_11_0.START_UP.t6 bgr_11_0.Vin-.t1 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X408 a_6540_22450.t6 a_6540_22450.t5 VDDA.t108 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X409 bgr_11_0.1st_Vout_1.t20 bgr_11_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 VDDA.t287 VDDA.t285 bgr_11_0.V_TOP.t8 VDDA.t286 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X411 VOUT+.t16 two_stage_opamp_dummy_magic_26_0.Y.t43 VDDA.t399 VDDA.t398 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X412 VOUT+.t97 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 VOUT-.t95 two_stage_opamp_dummy_magic_26_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 VOUT+.t98 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t2 bgr_11_0.V_TOP.t37 VDDA.t65 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X416 VOUT+.t99 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 two_stage_opamp_dummy_magic_26_0.V_source.t35 two_stage_opamp_dummy_magic_26_0.Vb1.t23 two_stage_opamp_dummy_magic_26_0.Vb1_2.t0 GNDA.t254 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X418 GNDA.t176 two_stage_opamp_dummy_magic_26_0.X.t42 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t4 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X419 VOUT-.t96 two_stage_opamp_dummy_magic_26_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X420 VOUT-.t97 two_stage_opamp_dummy_magic_26_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 GNDA.t179 two_stage_opamp_dummy_magic_26_0.X.t43 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t3 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X422 VOUT-.t98 two_stage_opamp_dummy_magic_26_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 VOUT+.t100 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X424 VOUT-.t99 two_stage_opamp_dummy_magic_26_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X425 VOUT+.t101 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 VOUT-.t100 two_stage_opamp_dummy_magic_26_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 VDDA.t330 VDDA.t328 two_stage_opamp_dummy_magic_26_0.Vb1.t3 VDDA.t329 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X428 VDDA.t241 bgr_11_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t7 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X429 two_stage_opamp_dummy_magic_26_0.VD4.t22 two_stage_opamp_dummy_magic_26_0.Vb3.t17 VDDA.t41 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X430 two_stage_opamp_dummy_magic_26_0.VD4.t13 two_stage_opamp_dummy_magic_26_0.Vb2.t22 two_stage_opamp_dummy_magic_26_0.Y.t4 two_stage_opamp_dummy_magic_26_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X431 VOUT+.t102 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 two_stage_opamp_dummy_magic_26_0.VD2.t14 two_stage_opamp_dummy_magic_26_0.Vb1.t24 two_stage_opamp_dummy_magic_26_0.Y.t12 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X433 VOUT+.t103 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 VOUT+.t104 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 bgr_11_0.PFET_GATE_10uA.t5 bgr_11_0.1st_Vout_2.t21 VDDA.t211 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X436 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t6 bgr_11_0.PFET_GATE_10uA.t19 VDDA.t239 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X437 bgr_11_0.1st_Vout_1.t21 bgr_11_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 two_stage_opamp_dummy_magic_26_0.V_source.t39 VIN+.t4 two_stage_opamp_dummy_magic_26_0.VD2.t21 GNDA.t252 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X439 VOUT-.t101 two_stage_opamp_dummy_magic_26_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 VOUT+.t105 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 two_stage_opamp_dummy_magic_26_0.V_source.t16 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t23 GNDA.t155 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X442 VDDA.t86 two_stage_opamp_dummy_magic_26_0.Vb3.t18 two_stage_opamp_dummy_magic_26_0.VD3.t21 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X443 VDDA.t6 two_stage_opamp_dummy_magic_26_0.V_err_gate.t8 two_stage_opamp_dummy_magic_26_0.V_err_mir_p.t2 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X444 GNDA.t291 bgr_11_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t4 GNDA.t290 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X445 VDDA.t78 bgr_11_0.V_TOP.t38 bgr_11_0.START_UP.t3 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X446 VDDA.t413 two_stage_opamp_dummy_magic_26_0.Vb3.t19 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t2 VDDA.t412 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X447 VOUT+.t106 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X448 VOUT-.t8 two_stage_opamp_dummy_magic_26_0.X.t44 VDDA.t97 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X449 bgr_11_0.Vin-.t5 bgr_11_0.V_TOP.t39 VDDA.t80 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X450 VOUT+.t107 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X451 bgr_11_0.1st_Vout_1.t22 bgr_11_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 VOUT-.t7 two_stage_opamp_dummy_magic_26_0.X.t45 VDDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X453 GNDA.t250 VDDA.t325 VDDA.t327 VDDA.t326 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X454 GNDA.t276 two_stage_opamp_dummy_magic_26_0.Y.t44 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t2 VDDA.t406 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X455 two_stage_opamp_dummy_magic_26_0.X.t20 two_stage_opamp_dummy_magic_26_0.Vb2.t23 two_stage_opamp_dummy_magic_26_0.VD3.t5 two_stage_opamp_dummy_magic_26_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X456 VOUT-.t102 two_stage_opamp_dummy_magic_26_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 VOUT-.t103 two_stage_opamp_dummy_magic_26_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X458 VOUT+.t108 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 VOUT-.t104 two_stage_opamp_dummy_magic_26_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X460 VOUT+.t109 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 VOUT+.t110 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 GNDA.t249 VDDA.t421 bgr_11_0.V_TOP.t6 GNDA.t248 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X463 bgr_11_0.1st_Vout_1.t23 bgr_11_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 GNDA.t223 bgr_11_0.NFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_26_0.V_err_gate.t2 GNDA.t222 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X465 VOUT-.t105 two_stage_opamp_dummy_magic_26_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X466 VOUT+.t111 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 bgr_11_0.V_TOP.t40 VDDA.t170 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X468 GNDA.t157 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t24 two_stage_opamp_dummy_magic_26_0.V_source.t15 GNDA.t156 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X469 VDDA.t32 two_stage_opamp_dummy_magic_26_0.Vb3.t20 two_stage_opamp_dummy_magic_26_0.VD4.t21 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X470 GNDA.t65 GNDA.t63 VDDA.t95 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X471 bgr_11_0.1st_Vout_2.t2 a_6540_22450.t16 VDDA.t94 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X472 VDDA.t156 two_stage_opamp_dummy_magic_26_0.Vb3.t21 two_stage_opamp_dummy_magic_26_0.VD3.t31 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X473 VOUT+.t112 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 VOUT+.t113 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 VOUT+.t14 VDDA.t322 VDDA.t324 VDDA.t323 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X476 VOUT+.t8 two_stage_opamp_dummy_magic_26_0.Y.t45 VDDA.t112 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X477 bgr_11_0.V_p_1.t2 VDDA.t422 GNDA.t247 GNDA.t246 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X478 VOUT-.t106 two_stage_opamp_dummy_magic_26_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X479 VOUT-.t107 two_stage_opamp_dummy_magic_26_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 bgr_11_0.NFET_GATE_10uA.t3 bgr_11_0.PFET_GATE_10uA.t20 VDDA.t237 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X481 VOUT+.t114 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X482 VOUT-.t108 two_stage_opamp_dummy_magic_26_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X483 GNDA.t62 GNDA.t60 VOUT-.t3 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X484 two_stage_opamp_dummy_magic_26_0.Vb3.t5 bgr_11_0.NFET_GATE_10uA.t15 GNDA.t146 GNDA.t145 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X485 GNDA.t177 two_stage_opamp_dummy_magic_26_0.X.t46 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t2 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X486 VOUT-.t109 two_stage_opamp_dummy_magic_26_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X487 VOUT+.t115 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 bgr_11_0.1st_Vout_2.t22 bgr_11_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X489 bgr_11_0.V_mir1.t6 bgr_11_0.V_mir1.t5 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X490 VOUT+.t116 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X491 bgr_11_0.1st_Vout_2.t0 bgr_11_0.V_CUR_REF_REG.t3 bgr_11_0.V_p_2.t1 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X492 two_stage_opamp_dummy_magic_26_0.V_source.t27 VIN-.t4 two_stage_opamp_dummy_magic_26_0.VD1.t3 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X493 two_stage_opamp_dummy_magic_26_0.VD2.t13 two_stage_opamp_dummy_magic_26_0.Vb1.t25 two_stage_opamp_dummy_magic_26_0.Y.t15 GNDA.t253 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X494 bgr_11_0.1st_Vout_1.t24 bgr_11_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t5 two_stage_opamp_dummy_magic_26_0.Y.t46 VDDA.t115 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X496 two_stage_opamp_dummy_magic_26_0.V_source.t8 VIN+.t5 two_stage_opamp_dummy_magic_26_0.VD2.t4 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X497 bgr_11_0.1st_Vout_2.t23 bgr_11_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 two_stage_opamp_dummy_magic_26_0.V_source.t14 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t25 GNDA.t205 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X499 VOUT+.t7 a_3830_106.t0 GNDA.t141 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X500 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t3 bgr_11_0.NFET_GATE_10uA.t16 GNDA.t144 GNDA.t143 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X501 two_stage_opamp_dummy_magic_26_0.V_source.t37 VIN-.t5 two_stage_opamp_dummy_magic_26_0.VD1.t19 GNDA.t251 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X502 GNDA.t45 GNDA.t46 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X503 GNDA.t22 bgr_11_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t2 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X504 VOUT-.t6 two_stage_opamp_dummy_magic_26_0.X.t47 VDDA.t393 VDDA.t392 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X505 VOUT-.t110 two_stage_opamp_dummy_magic_26_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X506 two_stage_opamp_dummy_magic_26_0.VD3.t33 two_stage_opamp_dummy_magic_26_0.Vb3.t22 VDDA.t178 VDDA.t177 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X507 VOUT+.t117 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X508 VOUT+.t118 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 bgr_11_0.1st_Vout_2.t24 bgr_11_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 GNDA.t265 two_stage_opamp_dummy_magic_26_0.Y.t47 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t1 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X511 GNDA.t29 two_stage_opamp_dummy_magic_26_0.err_amp_out.t5 two_stage_opamp_dummy_magic_26_0.V_source.t7 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X512 two_stage_opamp_dummy_magic_26_0.Y.t22 two_stage_opamp_dummy_magic_26_0.VD4.t24 two_stage_opamp_dummy_magic_26_0.VD4.t26 two_stage_opamp_dummy_magic_26_0.VD4.t25 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X513 VDDA.t395 two_stage_opamp_dummy_magic_26_0.Vb3.t23 two_stage_opamp_dummy_magic_26_0.VD4.t36 VDDA.t394 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X514 VOUT-.t18 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t7 GNDA.t268 GNDA.t267 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X515 VOUT-.t111 two_stage_opamp_dummy_magic_26_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 bgr_11_0.1st_Vout_1.t25 bgr_11_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 GNDA.t238 bgr_11_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_26_0.Vb2.t9 GNDA.t237 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X518 VOUT+.t119 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 bgr_11_0.1st_Vout_2.t25 bgr_11_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X520 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t12 bgr_11_0.NFET_GATE_10uA.t19 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X521 bgr_11_0.PFET_GATE_10uA.t4 bgr_11_0.1st_Vout_2.t26 VDDA.t209 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X522 VDDA.t321 VDDA.t318 VDDA.t320 VDDA.t319 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X523 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t9 two_stage_opamp_dummy_magic_26_0.X.t48 VDDA.t381 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X524 VOUT-.t112 two_stage_opamp_dummy_magic_26_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 VOUT+.t120 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t8 two_stage_opamp_dummy_magic_26_0.X.t49 VDDA.t159 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X527 bgr_11_0.1st_Vout_1.t26 bgr_11_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 VOUT-.t113 two_stage_opamp_dummy_magic_26_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 VOUT-.t114 two_stage_opamp_dummy_magic_26_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 VOUT+.t1 two_stage_opamp_dummy_magic_26_0.Y.t48 VDDA.t36 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X531 VOUT-.t115 two_stage_opamp_dummy_magic_26_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 bgr_11_0.1st_Vout_2.t27 bgr_11_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 GNDA.t45 GNDA.t59 bgr_11_0.Vin-.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X534 VOUT-.t116 two_stage_opamp_dummy_magic_26_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 VOUT+.t121 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 GNDA.t58 GNDA.t57 two_stage_opamp_dummy_magic_26_0.err_amp_out.t1 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X537 VDDA.t317 VDDA.t315 GNDA.t245 VDDA.t316 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X538 VOUT+.t122 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X539 bgr_11_0.1st_Vout_2.t6 a_6540_22450.t17 VDDA.t403 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X540 VDDA.t140 two_stage_opamp_dummy_magic_26_0.Vb3.t24 two_stage_opamp_dummy_magic_26_0.VD4.t31 VDDA.t139 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X541 two_stage_opamp_dummy_magic_26_0.Y.t0 two_stage_opamp_dummy_magic_26_0.Vb2.t24 two_stage_opamp_dummy_magic_26_0.VD4.t11 two_stage_opamp_dummy_magic_26_0.VD4.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X542 bgr_11_0.1st_Vout_1.t27 bgr_11_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 bgr_11_0.V_TOP.t3 bgr_11_0.1st_Vout_1.t28 VDDA.t134 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X544 GNDA.t173 two_stage_opamp_dummy_magic_26_0.X.t50 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t1 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X545 VOUT-.t117 two_stage_opamp_dummy_magic_26_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 two_stage_opamp_dummy_magic_26_0.V_source.t4 VIN-.t6 two_stage_opamp_dummy_magic_26_0.VD1.t0 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X547 VOUT+.t123 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 two_stage_opamp_dummy_magic_26_0.Vb1_2.t2 two_stage_opamp_dummy_magic_26_0.Vb1.t8 two_stage_opamp_dummy_magic_26_0.Vb1.t9 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X549 VOUT-.t118 two_stage_opamp_dummy_magic_26_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 bgr_11_0.1st_Vout_1.t6 bgr_11_0.V_mir1.t17 VDDA.t397 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X551 two_stage_opamp_dummy_magic_26_0.VD2.t12 two_stage_opamp_dummy_magic_26_0.Vb1.t26 two_stage_opamp_dummy_magic_26_0.Y.t17 GNDA.t252 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X552 VOUT-.t119 two_stage_opamp_dummy_magic_26_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t4 two_stage_opamp_dummy_magic_26_0.Y.t49 VDDA.t72 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X554 VDDA.t314 VDDA.t312 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t15 VDDA.t313 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X555 two_stage_opamp_dummy_magic_26_0.Vb2.t5 two_stage_opamp_dummy_magic_26_0.Vb2_2.t3 two_stage_opamp_dummy_magic_26_0.Vb2_2.t5 two_stage_opamp_dummy_magic_26_0.Vb2_2.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X556 two_stage_opamp_dummy_magic_26_0.VD3.t29 two_stage_opamp_dummy_magic_26_0.Vb3.t25 VDDA.t142 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X557 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t3 two_stage_opamp_dummy_magic_26_0.Y.t50 VDDA.t137 GNDA.t202 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X558 VOUT-.t120 two_stage_opamp_dummy_magic_26_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X559 VOUT-.t121 two_stage_opamp_dummy_magic_26_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X560 bgr_11_0.PFET_GATE_10uA.t0 VDDA.t423 GNDA.t244 GNDA.t243 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X561 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t11 bgr_11_0.PFET_GATE_10uA.t21 VDDA.t235 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X562 VOUT-.t122 two_stage_opamp_dummy_magic_26_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 two_stage_opamp_dummy_magic_26_0.V_p_mir.t1 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t26 GNDA.t275 GNDA.t274 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X564 VDDA.t311 VDDA.t309 VDDA.t311 VDDA.t310 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X565 two_stage_opamp_dummy_magic_26_0.V_source.t13 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t27 GNDA.t169 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X566 two_stage_opamp_dummy_magic_26_0.V_source.t2 VIN+.t6 two_stage_opamp_dummy_magic_26_0.VD2.t2 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X567 VDDA.t308 VDDA.t306 VOUT+.t13 VDDA.t307 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X568 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t11 VIN-.t7 two_stage_opamp_dummy_magic_26_0.V_p_mir.t0 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X569 two_stage_opamp_dummy_magic_26_0.V_source.t40 VIN-.t8 two_stage_opamp_dummy_magic_26_0.VD1.t21 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X570 VDDA.t305 VDDA.t303 two_stage_opamp_dummy_magic_26_0.err_amp_out.t3 VDDA.t304 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X571 bgr_11_0.V_TOP.t41 VDDA.t171 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 VOUT-.t5 two_stage_opamp_dummy_magic_26_0.X.t51 VDDA.t386 VDDA.t385 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X573 VDDA.t302 VDDA.t300 bgr_11_0.PFET_GATE_10uA.t3 VDDA.t301 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X574 VDDA.t168 bgr_11_0.V_TOP.t42 bgr_11_0.START_UP.t2 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X575 VDDA.t299 VDDA.t297 two_stage_opamp_dummy_magic_26_0.Vb2_2.t9 VDDA.t298 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X576 VOUT+.t124 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X577 VOUT+.t125 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 VOUT-.t123 two_stage_opamp_dummy_magic_26_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X579 a_6540_22450.t4 a_6540_22450.t3 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X580 VOUT-.t124 two_stage_opamp_dummy_magic_26_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X581 bgr_11_0.V_TOP.t43 VDDA.t169 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X582 VOUT-.t125 two_stage_opamp_dummy_magic_26_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X583 a_13840_3908.t0 two_stage_opamp_dummy_magic_26_0.V_tot.t0 GNDA.t25 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X584 two_stage_opamp_dummy_magic_26_0.VD3.t28 two_stage_opamp_dummy_magic_26_0.Vb3.t26 VDDA.t92 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X585 a_11420_30238.t0 a_11300_28630.t0 GNDA.t210 sky130_fd_pr__res_xhigh_po_0p35 l=6
X586 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t7 two_stage_opamp_dummy_magic_26_0.X.t52 VDDA.t148 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X587 VOUT+.t126 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X588 VOUT-.t126 two_stage_opamp_dummy_magic_26_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X589 VDDA.t233 bgr_11_0.PFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t5 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X590 VOUT+.t127 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X591 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t4 bgr_11_0.PFET_GATE_10uA.t23 VDDA.t231 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X592 two_stage_opamp_dummy_magic_26_0.Y.t8 two_stage_opamp_dummy_magic_26_0.Vb2.t25 two_stage_opamp_dummy_magic_26_0.VD4.t9 two_stage_opamp_dummy_magic_26_0.VD4.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X593 bgr_11_0.V_TOP.t44 VDDA.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 VOUT+.t128 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X595 VOUT+.t129 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X596 VOUT-.t127 two_stage_opamp_dummy_magic_26_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X597 bgr_11_0.1st_Vout_1.t0 bgr_11_0.V_mir1.t18 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X598 VOUT+.t130 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X599 VOUT+.t131 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X600 bgr_11_0.V_mir1.t0 bgr_11_0.Vin-.t8 bgr_11_0.V_p_1.t0 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X601 two_stage_opamp_dummy_magic_26_0.VD1.t12 two_stage_opamp_dummy_magic_26_0.Vb1.t27 two_stage_opamp_dummy_magic_26_0.X.t12 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X602 VOUT-.t128 two_stage_opamp_dummy_magic_26_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X603 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t12 bgr_11_0.PFET_GATE_10uA.t24 VDDA.t229 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X604 VDDA.t227 bgr_11_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t11 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X605 GNDA.t242 VDDA.t294 VDDA.t296 VDDA.t295 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X606 VOUT-.t129 two_stage_opamp_dummy_magic_26_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 VOUT-.t130 two_stage_opamp_dummy_magic_26_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X608 VOUT-.t131 two_stage_opamp_dummy_magic_26_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 VDDA.t293 VDDA.t291 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t15 VDDA.t292 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X610 VOUT-.t132 two_stage_opamp_dummy_magic_26_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 two_stage_opamp_dummy_magic_26_0.Vb1.t11 two_stage_opamp_dummy_magic_26_0.Vb1.t10 two_stage_opamp_dummy_magic_26_0.Vb1_2.t1 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X612 VOUT+.t132 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 two_stage_opamp_dummy_magic_26_0.VD2.t11 two_stage_opamp_dummy_magic_26_0.Vb1.t28 two_stage_opamp_dummy_magic_26_0.Y.t20 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X614 VOUT+.t133 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X615 VOUT+.t3 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t8 GNDA.t16 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X616 two_stage_opamp_dummy_magic_26_0.VD1.t11 two_stage_opamp_dummy_magic_26_0.Vb1.t29 two_stage_opamp_dummy_magic_26_0.X.t11 GNDA.t251 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X617 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t2 two_stage_opamp_dummy_magic_26_0.Y.t51 VDDA.t128 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X618 VOUT+.t134 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X619 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t1 bgr_11_0.V_TOP.t45 VDDA.t105 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X620 bgr_11_0.V_TOP.t46 VDDA.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X621 GNDA.t168 a_5820_28824.t1 GNDA.t167 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X622 two_stage_opamp_dummy_magic_26_0.V_source.t12 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t28 GNDA.t34 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X623 bgr_11_0.V_TOP.t11 bgr_11_0.1st_Vout_1.t29 VDDA.t405 VDDA.t404 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X624 two_stage_opamp_dummy_magic_26_0.V_source.t28 VIN-.t9 two_stage_opamp_dummy_magic_26_0.VD1.t4 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X625 VOUT+.t135 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 two_stage_opamp_dummy_magic_26_0.V_err_p.t2 two_stage_opamp_dummy_magic_26_0.V_err_gate.t9 VDDA.t71 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X627 VOUT-.t17 VDDA.t288 VDDA.t290 VDDA.t289 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X628 VOUT+.t136 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 VOUT-.t133 two_stage_opamp_dummy_magic_26_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X630 two_stage_opamp_dummy_magic_26_0.VD4.t7 two_stage_opamp_dummy_magic_26_0.Vb2.t26 two_stage_opamp_dummy_magic_26_0.Y.t10 two_stage_opamp_dummy_magic_26_0.VD4.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X631 two_stage_opamp_dummy_magic_26_0.VD3.t3 two_stage_opamp_dummy_magic_26_0.Vb2.t27 two_stage_opamp_dummy_magic_26_0.X.t0 two_stage_opamp_dummy_magic_26_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X632 VOUT-.t134 two_stage_opamp_dummy_magic_26_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X633 VOUT-.t135 two_stage_opamp_dummy_magic_26_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X634 bgr_11_0.V_TOP.t2 bgr_11_0.1st_Vout_1.t30 VDDA.t127 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X635 VOUT-.t136 two_stage_opamp_dummy_magic_26_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X636 VOUT+.t137 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X637 VOUT-.t137 two_stage_opamp_dummy_magic_26_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 bgr_11_0.1st_Vout_2.t28 bgr_11_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 two_stage_opamp_dummy_magic_26_0.Vb2_2.t2 two_stage_opamp_dummy_magic_26_0.Vb2.t28 VDDA.t17 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X640 two_stage_opamp_dummy_magic_26_0.VD1.t20 VIN-.t10 two_stage_opamp_dummy_magic_26_0.V_source.t38 GNDA.t255 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X641 VOUT+.t138 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X642 VDDA.t284 VDDA.t282 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t5 VDDA.t283 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X643 VOUT+.t139 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X644 two_stage_opamp_dummy_magic_26_0.Vb3.t4 bgr_11_0.NFET_GATE_10uA.t20 GNDA.t193 GNDA.t192 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X645 VOUT-.t138 two_stage_opamp_dummy_magic_26_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X646 bgr_11_0.1st_Vout_1.t31 bgr_11_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X647 a_3690_3908.t0 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t10 GNDA.t24 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X648 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t6 two_stage_opamp_dummy_magic_26_0.X.t53 VDDA.t18 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X649 two_stage_opamp_dummy_magic_26_0.VD2.t8 VIN+.t7 two_stage_opamp_dummy_magic_26_0.V_source.t33 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X650 a_13960_3908.t0 two_stage_opamp_dummy_magic_26_0.V_tot.t1 GNDA.t32 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X651 VOUT+.t140 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X652 VOUT-.t139 two_stage_opamp_dummy_magic_26_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 GNDA.t215 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t9 VOUT+.t11 GNDA.t214 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X654 bgr_11_0.Vin-.t0 bgr_11_0.START_UP.t7 bgr_11_0.V_TOP.t13 VDDA.t420 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X655 VOUT-.t140 two_stage_opamp_dummy_magic_26_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 VOUT+.t141 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 VOUT+.t142 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X658 VOUT+.t143 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 VOUT-.t141 two_stage_opamp_dummy_magic_26_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X660 bgr_11_0.V_mir1.t4 bgr_11_0.V_mir1.t3 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X661 two_stage_opamp_dummy_magic_26_0.VD4.t5 two_stage_opamp_dummy_magic_26_0.Vb2.t29 two_stage_opamp_dummy_magic_26_0.Y.t21 two_stage_opamp_dummy_magic_26_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X662 VOUT+.t144 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 VOUT-.t2 GNDA.t54 GNDA.t56 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X664 bgr_11_0.V_p_2.t0 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t9 a_6540_22450.t0 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X665 two_stage_opamp_dummy_magic_26_0.VD4.t30 two_stage_opamp_dummy_magic_26_0.Vb3.t27 VDDA.t114 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X666 VOUT-.t142 two_stage_opamp_dummy_magic_26_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X667 VOUT-.t143 two_stage_opamp_dummy_magic_26_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X668 VOUT-.t144 two_stage_opamp_dummy_magic_26_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X669 bgr_11_0.V_TOP.t7 VDDA.t279 VDDA.t281 VDDA.t280 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X670 two_stage_opamp_dummy_magic_26_0.VD1.t10 two_stage_opamp_dummy_magic_26_0.Vb1.t30 two_stage_opamp_dummy_magic_26_0.X.t18 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X671 VOUT-.t145 two_stage_opamp_dummy_magic_26_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X672 VOUT+.t145 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X673 bgr_11_0.V_TOP.t47 VDDA.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X674 VDDA.t100 bgr_11_0.V_TOP.t48 bgr_11_0.Vin-.t4 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X675 VOUT+.t146 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X676 VOUT+.t147 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X677 VOUT-.t146 two_stage_opamp_dummy_magic_26_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X678 two_stage_opamp_dummy_magic_26_0.Vb2_2.t1 two_stage_opamp_dummy_magic_26_0.Vb2.t0 two_stage_opamp_dummy_magic_26_0.Vb2.t1 two_stage_opamp_dummy_magic_26_0.Vb2_2.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X679 two_stage_opamp_dummy_magic_26_0.X.t7 two_stage_opamp_dummy_magic_26_0.VD3.t22 two_stage_opamp_dummy_magic_26_0.VD3.t24 two_stage_opamp_dummy_magic_26_0.VD3.t23 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X680 two_stage_opamp_dummy_magic_26_0.Vb1.t2 bgr_11_0.PFET_GATE_10uA.t26 VDDA.t225 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X681 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t3 bgr_11_0.PFET_GATE_10uA.t27 VDDA.t223 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X682 VDDA.t67 two_stage_opamp_dummy_magic_26_0.Vb3.t28 two_stage_opamp_dummy_magic_26_0.VD3.t20 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X683 VOUT-.t147 two_stage_opamp_dummy_magic_26_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 two_stage_opamp_dummy_magic_26_0.VD2.t10 two_stage_opamp_dummy_magic_26_0.Vb1.t31 two_stage_opamp_dummy_magic_26_0.Y.t16 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X685 GNDA.t165 a_6470_28630.t0 GNDA.t152 sky130_fd_pr__res_xhigh_po_0p35 l=6
X686 two_stage_opamp_dummy_magic_26_0.VD1.t9 two_stage_opamp_dummy_magic_26_0.Vb1.t32 two_stage_opamp_dummy_magic_26_0.X.t10 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X687 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t1 two_stage_opamp_dummy_magic_26_0.Y.t52 VDDA.t172 GNDA.t225 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X688 VOUT+.t148 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 VOUT-.t148 two_stage_opamp_dummy_magic_26_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 GNDA.t53 GNDA.t51 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t11 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X691 two_stage_opamp_dummy_magic_26_0.VD4.t3 two_stage_opamp_dummy_magic_26_0.Vb2.t30 two_stage_opamp_dummy_magic_26_0.Y.t23 two_stage_opamp_dummy_magic_26_0.VD4.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X692 VDDA.t187 a_6540_22450.t18 bgr_11_0.1st_Vout_2.t3 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X693 bgr_11_0.1st_Vout_2.t29 bgr_11_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 two_stage_opamp_dummy_magic_26_0.V_source.t11 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t29 GNDA.t39 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X695 two_stage_opamp_dummy_magic_26_0.V_err_gate.t5 VDDA.t276 VDDA.t278 VDDA.t277 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X696 GNDA.t227 bgr_11_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_26_0.Vb2.t7 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X697 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t0 GNDA.t48 GNDA.t50 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X698 GNDA.t240 VDDA.t424 bgr_11_0.V_p_2.t2 GNDA.t239 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X699 bgr_11_0.V_mir1.t2 bgr_11_0.V_mir1.t1 VDDA.t88 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X700 two_stage_opamp_dummy_magic_26_0.V_err_p.t1 two_stage_opamp_dummy_magic_26_0.V_tot.t5 two_stage_opamp_dummy_magic_26_0.err_amp_mir.t3 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X701 VOUT+.t149 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 bgr_11_0.PFET_GATE_10uA.t2 VDDA.t273 VDDA.t275 VDDA.t274 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X703 VDDA.t272 VDDA.t270 GNDA.t241 VDDA.t271 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X704 VDDA.t269 VDDA.t267 two_stage_opamp_dummy_magic_26_0.VD3.t35 VDDA.t268 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X705 a_12070_30088.t0 bgr_11_0.V_CUR_REF_REG.t0 GNDA.t166 sky130_fd_pr__res_xhigh_po_0p35 l=4
X706 VDDA.t143 two_stage_opamp_dummy_magic_26_0.Y.t53 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t0 GNDA.t207 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X707 VOUT+.t150 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X708 bgr_11_0.1st_Vout_2.t30 bgr_11_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X709 GNDA.t43 GNDA.t41 bgr_11_0.NFET_GATE_10uA.t0 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X710 bgr_11_0.Vin-.t3 bgr_11_0.V_TOP.t49 VDDA.t102 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X711 two_stage_opamp_dummy_magic_26_0.VD4.t1 two_stage_opamp_dummy_magic_26_0.Vb2.t31 two_stage_opamp_dummy_magic_26_0.Y.t7 two_stage_opamp_dummy_magic_26_0.VD4.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X712 two_stage_opamp_dummy_magic_26_0.VD2.t1 VIN+.t8 two_stage_opamp_dummy_magic_26_0.V_source.t1 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X713 VOUT-.t149 two_stage_opamp_dummy_magic_26_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X714 VOUT+.t151 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 GNDA.t286 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_26_0.V_source.t10 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X716 GNDA.t224 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t31 two_stage_opamp_dummy_magic_26_0.V_source.t9 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X717 two_stage_opamp_dummy_magic_26_0.VD2.t0 VIN+.t9 two_stage_opamp_dummy_magic_26_0.V_source.t0 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X718 two_stage_opamp_dummy_magic_26_0.V_p_mir.t3 VIN+.t10 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t2 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X719 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t5 two_stage_opamp_dummy_magic_26_0.X.t54 VDDA.t409 GNDA.t170 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X720 VDDA.t266 VDDA.t264 two_stage_opamp_dummy_magic_26_0.V_err_gate.t4 VDDA.t265 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X721 VOUT-.t150 two_stage_opamp_dummy_magic_26_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X722 VOUT+.t152 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X723 VDDA.t136 a_6540_22450.t1 a_6540_22450.t2 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X724 VOUT-.t151 two_stage_opamp_dummy_magic_26_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 VOUT-.t152 two_stage_opamp_dummy_magic_26_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 VOUT+.t153 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 bgr_11_0.1st_Vout_2.t31 bgr_11_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 two_stage_opamp_dummy_magic_26_0.X.t19 two_stage_opamp_dummy_magic_26_0.Vb2.t32 two_stage_opamp_dummy_magic_26_0.VD3.t1 two_stage_opamp_dummy_magic_26_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X729 VDDA.t263 VDDA.t261 VOUT-.t16 VDDA.t262 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X730 VOUT+.t154 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X731 bgr_11_0.V_CUR_REF_REG.t2 VDDA.t258 VDDA.t260 VDDA.t259 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X732 VOUT+.t155 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X733 two_stage_opamp_dummy_magic_26_0.Vb3.t3 bgr_11_0.NFET_GATE_10uA.t22 GNDA.t231 GNDA.t230 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X734 two_stage_opamp_dummy_magic_26_0.cap_res_X.t0 two_stage_opamp_dummy_magic_26_0.X.t2 GNDA.t26 sky130_fd_pr__res_high_po_1p41 l=1.41
X735 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t0 two_stage_opamp_dummy_magic_26_0.Y.t54 GNDA.t10 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X736 VOUT+.t156 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 VDDA.t221 bgr_11_0.PFET_GATE_10uA.t28 bgr_11_0.V_CUR_REF_REG.t1 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X738 GNDA.t191 bgr_11_0.NFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_26_0.Vb3.t2 GNDA.t190 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X739 VOUT-.t153 two_stage_opamp_dummy_magic_26_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X740 bgr_11_0.1st_Vout_1.t32 bgr_11_0.cap_res1.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X741 a_5700_30088.t0 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t0 GNDA.t0 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X742 VOUT-.t154 two_stage_opamp_dummy_magic_26_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X743 bgr_11_0.1st_Vout_2.t32 bgr_11_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 VOUT-.t155 two_stage_opamp_dummy_magic_26_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 VOUT-.t156 two_stage_opamp_dummy_magic_26_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.t15 362.341
R1 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.t14 355.094
R2 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n10 302.183
R3 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.n6 302.183
R4 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n5 297.683
R5 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t26 194.809
R6 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t9 194.809
R7 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t21 194.809
R8 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t7 194.809
R9 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n11 166.03
R10 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n8 166.03
R11 bgr_11_0.1st_Vout_2.t0 bgr_11_0.1st_Vout_2.n12 49.5021
R12 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t5 39.4005
R13 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t2 39.4005
R14 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t3 39.4005
R15 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t4 39.4005
R16 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t1 39.4005
R17 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t6 39.4005
R18 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.n0 35.7185
R19 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t32 4.8295
R20 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t12 4.8295
R21 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t13 4.8295
R22 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t19 4.8295
R23 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t30 4.8295
R24 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t11 4.8295
R25 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t23 4.8295
R26 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t28 4.8295
R27 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t8 4.8295
R28 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t27 4.5005
R29 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t20 4.5005
R30 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t31 4.5005
R31 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t25 4.5005
R32 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t24 4.5005
R33 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t18 4.5005
R34 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t17 4.5005
R35 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t10 4.5005
R36 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t29 4.5005
R37 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t22 4.5005
R38 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t16 4.5005
R39 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n3 4.5005
R40 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n9 2.90725
R41 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.n2 2.2095
R42 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n4 1.1255
R43 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n7 1.1255
R44 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.n1 0.8935
R45 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.t26 758.64
R46 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.n0 510.991
R47 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n25 509.226
R48 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t22 369.534
R49 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t27 369.534
R50 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.t11 369.534
R51 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.t10 369.534
R52 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.t25 369.534
R53 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t24 369.534
R54 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.n11 301.933
R55 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n9 301.933
R56 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.n7 301.933
R57 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.n5 301.933
R58 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t20 249.034
R59 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t28 249.034
R60 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t12 192.8
R61 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.t16 192.8
R62 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.t23 192.8
R63 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.t14 192.8
R64 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.t19 192.8
R65 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t18 192.8
R66 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.t21 192.8
R67 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.t15 192.8
R68 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.t17 192.8
R69 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t13 192.8
R70 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.n20 176.733
R71 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.n19 176.733
R72 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.n22 176.733
R73 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.n23 176.733
R74 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.n17 166.541
R75 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.n3 166.343
R76 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.t1 119.118
R77 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.t0 104.474
R78 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n16 56.2338
R79 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n15 56.2338
R80 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.n2 56.2338
R81 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.n1 56.2338
R82 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n21 56.2338
R83 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n24 56.2338
R84 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t6 39.4005
R85 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t2 39.4005
R86 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t8 39.4005
R87 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t4 39.4005
R88 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.t9 39.4005
R89 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.t5 39.4005
R90 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.t3 39.4005
R91 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.t7 39.4005
R92 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.n14 10.5161
R93 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.n12 6.15675
R94 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n4 2.28175
R95 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n18 2.28175
R96 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.n13 1.40675
R97 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.n6 1.1255
R98 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n8 1.1255
R99 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.n10 1.1255
R100 VDDA.n2565 VDDA.t306 1231.74
R101 VDDA.n2568 VDDA.t322 1231.74
R102 VDDA.n2430 VDDA.t261 1231.74
R103 VDDA.n2433 VDDA.t288 1231.74
R104 VDDA.n2447 VDDA.t303 858.933
R105 VDDA.n2492 VDDA.t276 858.933
R106 VDDA.n2487 VDDA.t264 858.933
R107 VDDA.n543 VDDA.t331 858.933
R108 VDDA.t302 VDDA.n2121 708.125
R109 VDDA.n2144 VDDA.t302 708.125
R110 VDDA.n2141 VDDA.t275 708.125
R111 VDDA.t275 VDDA.n2122 708.125
R112 VDDA.t354 VDDA.n2101 708.125
R113 VDDA.n2154 VDDA.t354 708.125
R114 VDDA.n2151 VDDA.t281 708.125
R115 VDDA.t281 VDDA.n2102 708.125
R116 VDDA.t367 VDDA.n2231 676.966
R117 VDDA.n2458 VDDA.t309 661.375
R118 VDDA.n2461 VDDA.t340 661.375
R119 VDDA.n2509 VDDA.t372 661.375
R120 VDDA.n2506 VDDA.t334 661.375
R121 VDDA.n557 VDDA.t267 661.375
R122 VDDA.n560 VDDA.t346 661.375
R123 VDDA.n2143 VDDA.t301 657.76
R124 VDDA.n2153 VDDA.t353 657.76
R125 VDDA.n2232 VDDA.t286 643.038
R126 VDDA.t313 VDDA.n2265 643.037
R127 VDDA.n2266 VDDA.t344 643.037
R128 VDDA.t292 VDDA.n2250 643.037
R129 VDDA.n2251 VDDA.t360 643.037
R130 VDDA.n2260 VDDA.t356 642.992
R131 VDDA.t338 VDDA.n2259 642.992
R132 VDDA.n2245 VDDA.t259 642.992
R133 VDDA.t350 VDDA.n2244 642.992
R134 VDDA.n1916 VDDA.t362 605.143
R135 VDDA.n1937 VDDA.t328 589.076
R136 VDDA.n589 VDDA.t270 589.076
R137 VDDA.n592 VDDA.t294 589.076
R138 VDDA.n2545 VDDA.t315 589.076
R139 VDDA.n2542 VDDA.t325 589.076
R140 VDDA.n2183 VDDA.n2181 587.407
R141 VDDA.n2187 VDDA.n2184 587.407
R142 VDDA.n2213 VDDA.n2212 587.407
R143 VDDA.n2208 VDDA.n2174 587.407
R144 VDDA.n2212 VDDA.n2211 585
R145 VDDA.n2210 VDDA.n2208 585
R146 VDDA.n2194 VDDA.n2183 585
R147 VDDA.n2191 VDDA.n2184 585
R148 VDDA.t274 VDDA.n2142 540.818
R149 VDDA.t280 VDDA.n2152 540.818
R150 VDDA.n1927 VDDA.t330 464.281
R151 VDDA.t330 VDDA.n1543 464.281
R152 VDDA.n1922 VDDA.t365 464.281
R153 VDDA.t365 VDDA.n1921 464.281
R154 VDDA.n2474 VDDA.t297 456.526
R155 VDDA.n2471 VDDA.t318 456.526
R156 VDDA.n2253 VDDA.t337 441.2
R157 VDDA.n2261 VDDA.t355 441.2
R158 VDDA.n2242 VDDA.t349 441.2
R159 VDDA.n2246 VDDA.t258 441.2
R160 VDDA.n2233 VDDA.t285 413.084
R161 VDDA.n2230 VDDA.t366 413.084
R162 VDDA.n2262 VDDA.t312 409.067
R163 VDDA.n2267 VDDA.t343 409.067
R164 VDDA.t301 VDDA.t214 407.144
R165 VDDA.t214 VDDA.t186 407.144
R166 VDDA.t186 VDDA.t197 407.144
R167 VDDA.t197 VDDA.t195 407.144
R168 VDDA.t195 VDDA.t162 407.144
R169 VDDA.t162 VDDA.t218 407.144
R170 VDDA.t218 VDDA.t210 407.144
R171 VDDA.t210 VDDA.t68 407.144
R172 VDDA.t68 VDDA.t402 407.144
R173 VDDA.t402 VDDA.t135 407.144
R174 VDDA.t135 VDDA.t107 407.144
R175 VDDA.t107 VDDA.t216 407.144
R176 VDDA.t216 VDDA.t208 407.144
R177 VDDA.t208 VDDA.t375 407.144
R178 VDDA.t375 VDDA.t93 407.144
R179 VDDA.t93 VDDA.t157 407.144
R180 VDDA.t157 VDDA.t23 407.144
R181 VDDA.t23 VDDA.t212 407.144
R182 VDDA.t212 VDDA.t274 407.144
R183 VDDA.t353 VDDA.t404 407.144
R184 VDDA.t404 VDDA.t203 407.144
R185 VDDA.t203 VDDA.t9 407.144
R186 VDDA.t9 VDDA.t47 407.144
R187 VDDA.t47 VDDA.t11 407.144
R188 VDDA.t11 VDDA.t164 407.144
R189 VDDA.t164 VDDA.t133 407.144
R190 VDDA.t133 VDDA.t201 407.144
R191 VDDA.t201 VDDA.t122 407.144
R192 VDDA.t122 VDDA.t377 407.144
R193 VDDA.t377 VDDA.t13 407.144
R194 VDDA.t13 VDDA.t189 407.144
R195 VDDA.t189 VDDA.t126 407.144
R196 VDDA.t126 VDDA.t184 407.144
R197 VDDA.t184 VDDA.t87 407.144
R198 VDDA.t87 VDDA.t151 407.144
R199 VDDA.t151 VDDA.t396 407.144
R200 VDDA.t396 VDDA.t109 407.144
R201 VDDA.t109 VDDA.t280 407.144
R202 VDDA.n2473 VDDA.t298 397.784
R203 VDDA.t319 VDDA.n2472 397.784
R204 VDDA.n2247 VDDA.t291 390.322
R205 VDDA.n2252 VDDA.t359 390.322
R206 VDDA.t256 VDDA.t313 373.214
R207 VDDA.t246 VDDA.t256 373.214
R208 VDDA.t234 VDDA.t246 373.214
R209 VDDA.t254 VDDA.t234 373.214
R210 VDDA.t344 VDDA.t254 373.214
R211 VDDA.t232 VDDA.t338 373.214
R212 VDDA.t252 VDDA.t232 373.214
R213 VDDA.t244 VDDA.t252 373.214
R214 VDDA.t230 VDDA.t244 373.214
R215 VDDA.t248 VDDA.t230 373.214
R216 VDDA.t238 VDDA.t248 373.214
R217 VDDA.t240 VDDA.t238 373.214
R218 VDDA.t222 VDDA.t240 373.214
R219 VDDA.t356 VDDA.t222 373.214
R220 VDDA.t228 VDDA.t292 373.214
R221 VDDA.t250 VDDA.t228 373.214
R222 VDDA.t242 VDDA.t250 373.214
R223 VDDA.t226 VDDA.t242 373.214
R224 VDDA.t360 VDDA.t226 373.214
R225 VDDA.t236 VDDA.t350 373.214
R226 VDDA.t220 VDDA.t236 373.214
R227 VDDA.t259 VDDA.t220 373.214
R228 VDDA.t286 VDDA.t15 373.214
R229 VDDA.t15 VDDA.t420 373.214
R230 VDDA.t420 VDDA.t367 373.214
R231 VDDA.n2146 VDDA.t300 370.168
R232 VDDA.n2139 VDDA.t273 370.168
R233 VDDA.n2156 VDDA.t352 370.168
R234 VDDA.n2149 VDDA.t279 370.168
R235 VDDA.n2165 VDDA.t282 360.868
R236 VDDA.n2219 VDDA.t369 360.868
R237 VDDA.n2260 VDDA.t358 354.154
R238 VDDA.n2259 VDDA.t339 354.154
R239 VDDA.n2245 VDDA.t260 354.154
R240 VDDA.n2244 VDDA.t351 354.154
R241 VDDA.n2232 VDDA.t287 354.063
R242 VDDA.n2231 VDDA.t368 347.224
R243 VDDA.t271 VDDA.n590 343.882
R244 VDDA.n591 VDDA.t295 343.882
R245 VDDA.n2544 VDDA.t316 343.882
R246 VDDA.t326 VDDA.n2543 343.882
R247 VDDA.n2279 VDDA.n2249 342.197
R248 VDDA.n2280 VDDA.n2248 342.197
R249 VDDA.n2268 VDDA.n2264 341.769
R250 VDDA.n2269 VDDA.n2263 341.769
R251 VDDA.n2272 VDDA.n2258 336.341
R252 VDDA.n2273 VDDA.n2257 336.341
R253 VDDA.n2274 VDDA.n2256 336.341
R254 VDDA.n2275 VDDA.n2255 336.341
R255 VDDA.n2276 VDDA.n2254 336.341
R256 VDDA.n2283 VDDA.n2243 336.341
R257 VDDA.n2250 VDDA.t293 332.267
R258 VDDA.n2251 VDDA.t361 332.267
R259 VDDA.n2265 VDDA.t314 332.084
R260 VDDA.n2266 VDDA.t345 332.084
R261 VDDA.n2138 VDDA.n2137 299.231
R262 VDDA.n2136 VDDA.n2135 299.231
R263 VDDA.n2134 VDDA.n2133 299.231
R264 VDDA.n2132 VDDA.n2131 299.231
R265 VDDA.n2130 VDDA.n2129 299.231
R266 VDDA.n2128 VDDA.n2127 299.231
R267 VDDA.n2126 VDDA.n2125 299.231
R268 VDDA.n2124 VDDA.n2123 299.231
R269 VDDA.n2120 VDDA.n2119 299.231
R270 VDDA.n2118 VDDA.n2117 299.231
R271 VDDA.n2116 VDDA.n2115 299.231
R272 VDDA.n2114 VDDA.n2113 299.231
R273 VDDA.n2112 VDDA.n2111 299.231
R274 VDDA.n2110 VDDA.n2109 299.231
R275 VDDA.n2108 VDDA.n2107 299.231
R276 VDDA.n2106 VDDA.n2105 299.231
R277 VDDA.n2104 VDDA.n2103 299.231
R278 VDDA.n2100 VDDA.n2099 299.231
R279 VDDA.n2446 VDDA.t304 282.788
R280 VDDA.n2491 VDDA.t277 282.788
R281 VDDA.n1933 VDDA.t329 267.188
R282 VDDA.t363 VDDA.n1925 267.188
R283 VDDA.t298 VDDA.t16 259.091
R284 VDDA.t16 VDDA.t319 259.091
R285 VDDA.t64 VDDA.t283 251.471
R286 VDDA.t77 VDDA.t64 251.471
R287 VDDA.t193 VDDA.t77 251.471
R288 VDDA.t99 VDDA.t193 251.471
R289 VDDA.t79 VDDA.t99 251.471
R290 VDDA.t182 VDDA.t79 251.471
R291 VDDA.t118 VDDA.t182 251.471
R292 VDDA.t51 VDDA.t118 251.471
R293 VDDA.t104 VDDA.t51 251.471
R294 VDDA.t62 VDDA.t104 251.471
R295 VDDA.t149 VDDA.t62 251.471
R296 VDDA.t7 VDDA.t149 251.471
R297 VDDA.t101 VDDA.t7 251.471
R298 VDDA.t167 VDDA.t101 251.471
R299 VDDA.t28 VDDA.t167 251.471
R300 VDDA.t60 VDDA.t28 251.471
R301 VDDA.t370 VDDA.t60 251.471
R302 VDDA.n1924 VDDA.n1923 238.367
R303 VDDA.n1550 VDDA.n1546 238.367
R304 VDDA.n2215 VDDA.n2214 238.367
R305 VDDA.n2142 VDDA.n2141 238.367
R306 VDDA.n2142 VDDA.n2122 238.367
R307 VDDA.n2152 VDDA.n2151 238.367
R308 VDDA.n2152 VDDA.n2102 238.367
R309 VDDA.t283 VDDA.n2199 237.5
R310 VDDA.n2216 VDDA.t370 237.5
R311 VDDA.n542 VDDA.n541 222.524
R312 VDDA.n2450 VDDA.n2449 222.524
R313 VDDA.n2490 VDDA.t332 221.121
R314 VDDA.t265 VDDA.n2490 221.121
R315 VDDA.t329 VDDA.t224 217.708
R316 VDDA.t224 VDDA.t363 217.708
R317 VDDA.t391 VDDA.t271 217.708
R318 VDDA.t56 VDDA.t391 217.708
R319 VDDA.t19 VDDA.t56 217.708
R320 VDDA.t387 VDDA.t19 217.708
R321 VDDA.t84 VDDA.t387 217.708
R322 VDDA.t22 VDDA.t84 217.708
R323 VDDA.t54 VDDA.t22 217.708
R324 VDDA.t207 VDDA.t54 217.708
R325 VDDA.t4 VDDA.t207 217.708
R326 VDDA.t98 VDDA.t4 217.708
R327 VDDA.t295 VDDA.t98 217.708
R328 VDDA.t316 VDDA.t401 217.708
R329 VDDA.t401 VDDA.t390 217.708
R330 VDDA.t390 VDDA.t406 217.708
R331 VDDA.t406 VDDA.t132 217.708
R332 VDDA.t132 VDDA.t389 217.708
R333 VDDA.t389 VDDA.t37 217.708
R334 VDDA.t37 VDDA.t400 217.708
R335 VDDA.t400 VDDA.t34 217.708
R336 VDDA.t34 VDDA.t129 217.708
R337 VDDA.t129 VDDA.t116 217.708
R338 VDDA.t116 VDDA.t326 217.708
R339 VDDA.t310 VDDA.n2459 213.131
R340 VDDA.n2460 VDDA.t341 213.131
R341 VDDA.n2508 VDDA.t373 213.131
R342 VDDA.t335 VDDA.n2507 213.131
R343 VDDA.t268 VDDA.n558 213.131
R344 VDDA.n559 VDDA.t347 213.131
R345 VDDA.n1549 VDDA.n1547 185
R346 VDDA.n1920 VDDA.n1919 185
R347 VDDA.n1932 VDDA.n1931 185
R348 VDDA.n1933 VDDA.n1932 185
R349 VDDA.n1929 VDDA.n1926 185
R350 VDDA.n1928 VDDA.n1544 185
R351 VDDA.n1935 VDDA.n1934 185
R352 VDDA.n1934 VDDA.n1933 185
R353 VDDA.n2204 VDDA.n2202 185
R354 VDDA.n2211 VDDA.n2201 185
R355 VDDA.n2216 VDDA.n2201 185
R356 VDDA.n2210 VDDA.n2209 185
R357 VDDA.n2207 VDDA.n2176 185
R358 VDDA.n2218 VDDA.n2217 185
R359 VDDA.n2217 VDDA.n2216 185
R360 VDDA.n2198 VDDA.n2197 185
R361 VDDA.n2199 VDDA.n2198 185
R362 VDDA.n2195 VDDA.n2180 185
R363 VDDA.n2194 VDDA.n2193 185
R364 VDDA.n2192 VDDA.n2191 185
R365 VDDA.n2186 VDDA.n2185 185
R366 VDDA.n2188 VDDA.n2179 185
R367 VDDA.n2199 VDDA.n2179 185
R368 VDDA.t304 VDDA.t181 180.173
R369 VDDA.t181 VDDA.t70 180.173
R370 VDDA.t70 VDDA.t0 180.173
R371 VDDA.t0 VDDA.t166 180.173
R372 VDDA.t166 VDDA.t332 180.173
R373 VDDA.t33 VDDA.t265 180.173
R374 VDDA.t2 VDDA.t33 180.173
R375 VDDA.t5 VDDA.t2 180.173
R376 VDDA.t120 VDDA.t5 180.173
R377 VDDA.t277 VDDA.t120 180.173
R378 VDDA.n2473 VDDA.t299 168.139
R379 VDDA.n2472 VDDA.t321 168.139
R380 VDDA.n2470 VDDA.n2469 150.643
R381 VDDA.n1919 VDDA.n1547 150
R382 VDDA.n1932 VDDA.n1926 150
R383 VDDA.n1934 VDDA.n1544 150
R384 VDDA.n2202 VDDA.n2201 150
R385 VDDA.n2209 VDDA.n2201 150
R386 VDDA.n2217 VDDA.n2176 150
R387 VDDA.n2198 VDDA.n2180 150
R388 VDDA.n2193 VDDA.n2192 150
R389 VDDA.n2185 VDDA.n2179 150
R390 VDDA.n1552 VDDA.n1551 149.112
R391 VDDA.t412 VDDA.t310 146.155
R392 VDDA.t341 VDDA.t412 146.155
R393 VDDA.t373 VDDA.t113 146.155
R394 VDDA.t113 VDDA.t139 146.155
R395 VDDA.t139 VDDA.t40 146.155
R396 VDDA.t40 VDDA.t199 146.155
R397 VDDA.t199 VDDA.t25 146.155
R398 VDDA.t25 VDDA.t81 146.155
R399 VDDA.t81 VDDA.t191 146.155
R400 VDDA.t191 VDDA.t394 146.155
R401 VDDA.t394 VDDA.t418 146.155
R402 VDDA.t418 VDDA.t31 146.155
R403 VDDA.t31 VDDA.t335 146.155
R404 VDDA.t91 VDDA.t268 146.155
R405 VDDA.t155 VDDA.t91 146.155
R406 VDDA.t153 VDDA.t155 146.155
R407 VDDA.t179 VDDA.t153 146.155
R408 VDDA.t410 VDDA.t179 146.155
R409 VDDA.t66 VDDA.t410 146.155
R410 VDDA.t141 VDDA.t66 146.155
R411 VDDA.t85 VDDA.t141 146.155
R412 VDDA.t177 VDDA.t85 146.155
R413 VDDA.t160 VDDA.t177 146.155
R414 VDDA.t347 VDDA.t160 146.155
R415 VDDA.n2220 VDDA.n2173 141.712
R416 VDDA.n2221 VDDA.n2172 141.712
R417 VDDA.n2222 VDDA.n2171 141.712
R418 VDDA.n2223 VDDA.n2170 141.712
R419 VDDA.n2224 VDDA.n2169 141.712
R420 VDDA.n2225 VDDA.n2168 141.712
R421 VDDA.n2226 VDDA.n2167 141.712
R422 VDDA.n2227 VDDA.n2166 141.712
R423 VDDA.n590 VDDA.t272 136.701
R424 VDDA.n591 VDDA.t296 136.701
R425 VDDA.n2544 VDDA.t317 136.701
R426 VDDA.n2543 VDDA.t327 136.701
R427 VDDA.t284 VDDA.n2183 123.126
R428 VDDA.n2184 VDDA.t284 123.126
R429 VDDA.n2212 VDDA.t371 123.126
R430 VDDA.n2208 VDDA.t371 123.126
R431 VDDA.t307 VDDA.n2566 122.829
R432 VDDA.n2567 VDDA.t323 122.829
R433 VDDA.t262 VDDA.n2431 122.829
R434 VDDA.n2432 VDDA.t289 122.829
R435 VDDA.n2446 VDDA.t305 113.26
R436 VDDA.n2491 VDDA.t278 113.26
R437 VDDA.n2489 VDDA.t266 113.26
R438 VDDA.n2489 VDDA.t333 113.26
R439 VDDA.n2492 VDDA.n2491 82.7434
R440 VDDA.n2447 VDDA.n2446 82.7434
R441 VDDA.t130 VDDA.t307 81.6411
R442 VDDA.t73 VDDA.t130 81.6411
R443 VDDA.t111 VDDA.t73 81.6411
R444 VDDA.t173 VDDA.t111 81.6411
R445 VDDA.t35 VDDA.t173 81.6411
R446 VDDA.t145 VDDA.t35 81.6411
R447 VDDA.t415 VDDA.t145 81.6411
R448 VDDA.t407 VDDA.t415 81.6411
R449 VDDA.t398 VDDA.t407 81.6411
R450 VDDA.t38 VDDA.t398 81.6411
R451 VDDA.t323 VDDA.t38 81.6411
R452 VDDA.t383 VDDA.t262 81.6411
R453 VDDA.t205 VDDA.t383 81.6411
R454 VDDA.t20 VDDA.t205 81.6411
R455 VDDA.t44 VDDA.t20 81.6411
R456 VDDA.t96 VDDA.t44 81.6411
R457 VDDA.t175 VDDA.t96 81.6411
R458 VDDA.t392 VDDA.t175 81.6411
R459 VDDA.t89 VDDA.t392 81.6411
R460 VDDA.t385 VDDA.t89 81.6411
R461 VDDA.t58 VDDA.t385 81.6411
R462 VDDA.t289 VDDA.t58 81.6411
R463 VDDA.n2459 VDDA.t311 76.2576
R464 VDDA.n2460 VDDA.t342 76.2576
R465 VDDA.n2508 VDDA.t374 76.2576
R466 VDDA.n2507 VDDA.t336 76.2576
R467 VDDA.n558 VDDA.t269 76.2576
R468 VDDA.n559 VDDA.t348 76.2576
R469 VDDA.n2505 VDDA.n2504 71.388
R470 VDDA.n2503 VDDA.n2502 71.388
R471 VDDA.n2501 VDDA.n2500 71.388
R472 VDDA.n2499 VDDA.n2498 71.388
R473 VDDA.n2497 VDDA.n2496 71.388
R474 VDDA.n548 VDDA.n547 71.388
R475 VDDA.n550 VDDA.n549 71.388
R476 VDDA.n552 VDDA.n551 71.388
R477 VDDA.n554 VDDA.n553 71.388
R478 VDDA.n556 VDDA.n555 71.388
R479 VDDA.n2457 VDDA.n2456 68.4557
R480 VDDA.n1925 VDDA.n1924 65.8183
R481 VDDA.n1925 VDDA.n1546 65.8183
R482 VDDA.n1933 VDDA.n1545 65.8183
R483 VDDA.n2216 VDDA.n2215 65.8183
R484 VDDA.n2216 VDDA.n2200 65.8183
R485 VDDA.n2199 VDDA.n2177 65.8183
R486 VDDA.n2199 VDDA.n2178 65.8183
R487 VDDA.n2490 VDDA.n2489 61.6672
R488 VDDA.n2488 VDDA.n2487 60.8005
R489 VDDA.n2488 VDDA.n543 60.8005
R490 VDDA.n2090 VDDA.t421 58.8005
R491 VDDA.n2089 VDDA.t423 58.8005
R492 VDDA.n1924 VDDA.n1547 53.3664
R493 VDDA.n1919 VDDA.n1546 53.3664
R494 VDDA.n1926 VDDA.n1545 53.3664
R495 VDDA.n1545 VDDA.n1544 53.3664
R496 VDDA.n2209 VDDA.n2200 53.3664
R497 VDDA.n2215 VDDA.n2202 53.3664
R498 VDDA.n2200 VDDA.n2176 53.3664
R499 VDDA.n2180 VDDA.n2177 53.3664
R500 VDDA.n2192 VDDA.n2178 53.3664
R501 VDDA.n2193 VDDA.n2177 53.3664
R502 VDDA.n2185 VDDA.n2178 53.3664
R503 VDDA.n2089 VDDA.t424 49.1638
R504 VDDA.n2091 VDDA.t422 48.5162
R505 VDDA.n2566 VDDA.t308 40.9789
R506 VDDA.n2567 VDDA.t324 40.9789
R507 VDDA.n2431 VDDA.t263 40.9789
R508 VDDA.n2432 VDDA.t290 40.9789
R509 VDDA.n2264 VDDA.t235 39.4005
R510 VDDA.n2264 VDDA.t255 39.4005
R511 VDDA.n2263 VDDA.t257 39.4005
R512 VDDA.n2263 VDDA.t247 39.4005
R513 VDDA.n2258 VDDA.t223 39.4005
R514 VDDA.n2258 VDDA.t357 39.4005
R515 VDDA.n2257 VDDA.t239 39.4005
R516 VDDA.n2257 VDDA.t241 39.4005
R517 VDDA.n2256 VDDA.t231 39.4005
R518 VDDA.n2256 VDDA.t249 39.4005
R519 VDDA.n2255 VDDA.t253 39.4005
R520 VDDA.n2255 VDDA.t245 39.4005
R521 VDDA.t339 VDDA.n2254 39.4005
R522 VDDA.n2254 VDDA.t233 39.4005
R523 VDDA.n2249 VDDA.t243 39.4005
R524 VDDA.n2249 VDDA.t227 39.4005
R525 VDDA.n2248 VDDA.t229 39.4005
R526 VDDA.n2248 VDDA.t251 39.4005
R527 VDDA.n2243 VDDA.t237 39.4005
R528 VDDA.n2243 VDDA.t221 39.4005
R529 VDDA.n2137 VDDA.t24 39.4005
R530 VDDA.n2137 VDDA.t213 39.4005
R531 VDDA.n2135 VDDA.t94 39.4005
R532 VDDA.n2135 VDDA.t158 39.4005
R533 VDDA.n2133 VDDA.t209 39.4005
R534 VDDA.n2133 VDDA.t376 39.4005
R535 VDDA.n2131 VDDA.t108 39.4005
R536 VDDA.n2131 VDDA.t217 39.4005
R537 VDDA.n2129 VDDA.t403 39.4005
R538 VDDA.n2129 VDDA.t136 39.4005
R539 VDDA.n2127 VDDA.t211 39.4005
R540 VDDA.n2127 VDDA.t69 39.4005
R541 VDDA.n2125 VDDA.t163 39.4005
R542 VDDA.n2125 VDDA.t219 39.4005
R543 VDDA.n2123 VDDA.t198 39.4005
R544 VDDA.n2123 VDDA.t196 39.4005
R545 VDDA.n2119 VDDA.t215 39.4005
R546 VDDA.n2119 VDDA.t187 39.4005
R547 VDDA.n2117 VDDA.t397 39.4005
R548 VDDA.n2117 VDDA.t110 39.4005
R549 VDDA.n2115 VDDA.t88 39.4005
R550 VDDA.n2115 VDDA.t152 39.4005
R551 VDDA.n2113 VDDA.t127 39.4005
R552 VDDA.n2113 VDDA.t185 39.4005
R553 VDDA.n2111 VDDA.t14 39.4005
R554 VDDA.n2111 VDDA.t190 39.4005
R555 VDDA.n2109 VDDA.t123 39.4005
R556 VDDA.n2109 VDDA.t378 39.4005
R557 VDDA.n2107 VDDA.t134 39.4005
R558 VDDA.n2107 VDDA.t202 39.4005
R559 VDDA.n2105 VDDA.t12 39.4005
R560 VDDA.n2105 VDDA.t165 39.4005
R561 VDDA.n2103 VDDA.t10 39.4005
R562 VDDA.n2103 VDDA.t48 39.4005
R563 VDDA.n2099 VDDA.t405 39.4005
R564 VDDA.n2099 VDDA.t204 39.4005
R565 VDDA.n536 VDDA.n535 38.2695
R566 VDDA.n2557 VDDA.n2556 38.2695
R567 VDDA.n2559 VDDA.n2558 38.2695
R568 VDDA.n2561 VDDA.n2560 38.2695
R569 VDDA.n2563 VDDA.n2562 38.2695
R570 VDDA.n601 VDDA.n600 38.2695
R571 VDDA.n2422 VDDA.n2421 38.2695
R572 VDDA.n2424 VDDA.n2423 38.2695
R573 VDDA.n2426 VDDA.n2425 38.2695
R574 VDDA.n2428 VDDA.n2427 38.2695
R575 VDDA.n2267 VDDA.n2266 27.2462
R576 VDDA.n2265 VDDA.n2262 27.2462
R577 VDDA.n2252 VDDA.n2251 27.2462
R578 VDDA.n2250 VDDA.n2247 27.2462
R579 VDDA.n575 VDDA.n573 26.8887
R580 VDDA.n2527 VDDA.n2525 26.8887
R581 VDDA.n583 VDDA.n582 26.7741
R582 VDDA.n581 VDDA.n580 26.7741
R583 VDDA.n579 VDDA.n578 26.7741
R584 VDDA.n577 VDDA.n576 26.7741
R585 VDDA.n575 VDDA.n574 26.7741
R586 VDDA.n2527 VDDA.n2526 26.7741
R587 VDDA.n2529 VDDA.n2528 26.7741
R588 VDDA.n2531 VDDA.n2530 26.7741
R589 VDDA.n2533 VDDA.n2532 26.7741
R590 VDDA.n2535 VDDA.n2534 26.7741
R591 VDDA.n2261 VDDA.n2260 24.9931
R592 VDDA.n2259 VDDA.n2253 24.9931
R593 VDDA.n2246 VDDA.n2245 24.9931
R594 VDDA.n2244 VDDA.n2242 24.9931
R595 VDDA.n1611 VDDA.t46 24.1029
R596 VDDA.n2233 VDDA.n2232 22.9536
R597 VDDA.n2219 VDDA.n2218 22.8576
R598 VDDA.n2188 VDDA.n2165 22.8576
R599 VDDA.n2469 VDDA.t17 21.8894
R600 VDDA.n2469 VDDA.t320 21.8894
R601 VDDA.n2231 VDDA.n2230 20.4312
R602 VDDA.n1551 VDDA.t225 19.7005
R603 VDDA.n1551 VDDA.t364 19.7005
R604 VDDA.n541 VDDA.t3 15.7605
R605 VDDA.n541 VDDA.t6 15.7605
R606 VDDA.n2449 VDDA.t71 15.7605
R607 VDDA.n2449 VDDA.t1 15.7605
R608 VDDA.n2489 VDDA.n2488 13.9641
R609 VDDA.n2173 VDDA.t29 13.1338
R610 VDDA.n2173 VDDA.t61 13.1338
R611 VDDA.n2172 VDDA.t102 13.1338
R612 VDDA.n2172 VDDA.t168 13.1338
R613 VDDA.n2171 VDDA.t150 13.1338
R614 VDDA.n2171 VDDA.t8 13.1338
R615 VDDA.n2170 VDDA.t105 13.1338
R616 VDDA.n2170 VDDA.t63 13.1338
R617 VDDA.n2169 VDDA.t119 13.1338
R618 VDDA.n2169 VDDA.t52 13.1338
R619 VDDA.n2168 VDDA.t80 13.1338
R620 VDDA.n2168 VDDA.t183 13.1338
R621 VDDA.n2167 VDDA.t194 13.1338
R622 VDDA.n2167 VDDA.t100 13.1338
R623 VDDA.n2166 VDDA.t65 13.1338
R624 VDDA.n2166 VDDA.t78 13.1338
R625 VDDA.n2230 VDDA.n2229 11.37
R626 VDDA.n2234 VDDA.n2233 11.37
R627 VDDA.t311 VDDA.n2457 11.2576
R628 VDDA.n2457 VDDA.t413 11.2576
R629 VDDA.n2504 VDDA.t419 11.2576
R630 VDDA.n2504 VDDA.t32 11.2576
R631 VDDA.n2502 VDDA.t192 11.2576
R632 VDDA.n2502 VDDA.t395 11.2576
R633 VDDA.n2500 VDDA.t26 11.2576
R634 VDDA.n2500 VDDA.t82 11.2576
R635 VDDA.n2498 VDDA.t41 11.2576
R636 VDDA.n2498 VDDA.t200 11.2576
R637 VDDA.n2496 VDDA.t114 11.2576
R638 VDDA.n2496 VDDA.t140 11.2576
R639 VDDA.n547 VDDA.t178 11.2576
R640 VDDA.n547 VDDA.t161 11.2576
R641 VDDA.n549 VDDA.t142 11.2576
R642 VDDA.n549 VDDA.t86 11.2576
R643 VDDA.n551 VDDA.t411 11.2576
R644 VDDA.n551 VDDA.t67 11.2576
R645 VDDA.n553 VDDA.t154 11.2576
R646 VDDA.n553 VDDA.t180 11.2576
R647 VDDA.n555 VDDA.t92 11.2576
R648 VDDA.n555 VDDA.t156 11.2576
R649 VDDA.n2220 VDDA.n2219 11.0575
R650 VDDA.n2268 VDDA.n2267 10.9846
R651 VDDA.n2270 VDDA.n2262 10.87
R652 VDDA.n2277 VDDA.n2253 10.87
R653 VDDA.n2281 VDDA.n2247 10.87
R654 VDDA.n2284 VDDA.n2242 10.87
R655 VDDA.n2282 VDDA.n2246 10.87
R656 VDDA.n2278 VDDA.n2252 10.87
R657 VDDA.n2271 VDDA.n2261 10.87
R658 VDDA.n2228 VDDA.n2165 10.87
R659 VDDA.n2448 VDDA.n2447 10.8696
R660 VDDA.n2493 VDDA.n2492 10.869
R661 VDDA.n1923 VDDA.n1548 9.50883
R662 VDDA.n1931 VDDA.n1930 9.50883
R663 VDDA.n2197 VDDA.n2196 9.50883
R664 VDDA.n2189 VDDA.n2188 9.50883
R665 VDDA.n2214 VDDA.n2203 9.50883
R666 VDDA.n2218 VDDA.n2175 9.50883
R667 VDDA.n2145 VDDA.n2121 9.50883
R668 VDDA.n2155 VDDA.n2101 9.50883
R669 VDDA.n1920 VDDA.n1918 9.3005
R670 VDDA.n1549 VDDA.n1548 9.3005
R671 VDDA.n1917 VDDA.n1550 9.3005
R672 VDDA.n1928 VDDA.n1542 9.3005
R673 VDDA.n1930 VDDA.n1929 9.3005
R674 VDDA.n1936 VDDA.n1935 9.3005
R675 VDDA.n2207 VDDA.n2175 9.3005
R676 VDDA.n2210 VDDA.n2206 9.3005
R677 VDDA.n2211 VDDA.n2205 9.3005
R678 VDDA.n2204 VDDA.n2203 9.3005
R679 VDDA.n2189 VDDA.n2186 9.3005
R680 VDDA.n2191 VDDA.n2190 9.3005
R681 VDDA.n2194 VDDA.n2182 9.3005
R682 VDDA.n2196 VDDA.n2195 9.3005
R683 VDDA.n2145 VDDA.n2144 9.3005
R684 VDDA.n2155 VDDA.n2154 9.3005
R685 VDDA.n2487 VDDA.n2486 9.3005
R686 VDDA.n2486 VDDA.n543 9.3005
R687 VDDA.n1920 VDDA.n1549 9.14336
R688 VDDA.n1929 VDDA.n1928 9.14336
R689 VDDA.n2211 VDDA.n2204 9.14336
R690 VDDA.n2211 VDDA.n2210 9.14336
R691 VDDA.n2210 VDDA.n2207 9.14336
R692 VDDA.n2195 VDDA.n2194 9.14336
R693 VDDA.n2194 VDDA.n2191 9.14336
R694 VDDA.n2191 VDDA.n2186 9.14336
R695 VDDA.n582 VDDA.t409 8.0005
R696 VDDA.n582 VDDA.t124 8.0005
R697 VDDA.n580 VDDA.t18 8.0005
R698 VDDA.n580 VDDA.t388 8.0005
R699 VDDA.n578 VDDA.t148 8.0005
R700 VDDA.n578 VDDA.t43 8.0005
R701 VDDA.n576 VDDA.t381 8.0005
R702 VDDA.n576 VDDA.t382 8.0005
R703 VDDA.n574 VDDA.t159 8.0005
R704 VDDA.n574 VDDA.t106 8.0005
R705 VDDA.n573 VDDA.t95 8.0005
R706 VDDA.n573 VDDA.t83 8.0005
R707 VDDA.n2525 VDDA.t72 8.0005
R708 VDDA.n2525 VDDA.t125 8.0005
R709 VDDA.n2526 VDDA.t115 8.0005
R710 VDDA.n2526 VDDA.t147 8.0005
R711 VDDA.n2528 VDDA.t172 8.0005
R712 VDDA.n2528 VDDA.t138 8.0005
R713 VDDA.n2530 VDDA.t128 8.0005
R714 VDDA.n2530 VDDA.t144 8.0005
R715 VDDA.n2532 VDDA.t137 8.0005
R716 VDDA.n2532 VDDA.t417 8.0005
R717 VDDA.n2534 VDDA.t121 8.0005
R718 VDDA.n2534 VDDA.t143 8.0005
R719 VDDA.n535 VDDA.t399 6.56717
R720 VDDA.n535 VDDA.t39 6.56717
R721 VDDA.n2556 VDDA.t416 6.56717
R722 VDDA.n2556 VDDA.t408 6.56717
R723 VDDA.n2558 VDDA.t36 6.56717
R724 VDDA.n2558 VDDA.t146 6.56717
R725 VDDA.n2560 VDDA.t112 6.56717
R726 VDDA.n2560 VDDA.t174 6.56717
R727 VDDA.n2562 VDDA.t131 6.56717
R728 VDDA.n2562 VDDA.t74 6.56717
R729 VDDA.n600 VDDA.t386 6.56717
R730 VDDA.n600 VDDA.t59 6.56717
R731 VDDA.n2421 VDDA.t393 6.56717
R732 VDDA.n2421 VDDA.t90 6.56717
R733 VDDA.n2423 VDDA.t97 6.56717
R734 VDDA.n2423 VDDA.t176 6.56717
R735 VDDA.n2425 VDDA.t21 6.56717
R736 VDDA.n2425 VDDA.t45 6.56717
R737 VDDA.n2427 VDDA.t384 6.56717
R738 VDDA.n2427 VDDA.t206 6.56717
R739 VDDA.n1923 VDDA.n1922 5.33286
R740 VDDA.n1921 VDDA.n1550 5.33286
R741 VDDA.n1931 VDDA.n1927 5.33286
R742 VDDA.n1935 VDDA.n1543 5.33286
R743 VDDA.n2214 VDDA.n2213 5.33286
R744 VDDA.n2218 VDDA.n2174 5.33286
R745 VDDA.n2197 VDDA.n2181 5.33286
R746 VDDA.n2188 VDDA.n2187 5.33286
R747 VDDA.n2506 VDDA.n2505 4.8755
R748 VDDA.n557 VDDA.n556 4.8755
R749 VDDA.n1940 VDDA.n1939 4.5005
R750 VDDA.n1943 VDDA.n1942 4.5005
R751 VDDA.n1944 VDDA.n1540 4.5005
R752 VDDA.n1948 VDDA.n1945 4.5005
R753 VDDA.n1949 VDDA.n1539 4.5005
R754 VDDA.n1953 VDDA.n1952 4.5005
R755 VDDA.n1954 VDDA.n1538 4.5005
R756 VDDA.n1958 VDDA.n1955 4.5005
R757 VDDA.n1959 VDDA.n1537 4.5005
R758 VDDA.n1963 VDDA.n1962 4.5005
R759 VDDA.n1964 VDDA.n1536 4.5005
R760 VDDA.n1968 VDDA.n1965 4.5005
R761 VDDA.n1969 VDDA.n1535 4.5005
R762 VDDA.n1973 VDDA.n1972 4.5005
R763 VDDA.n1974 VDDA.n1534 4.5005
R764 VDDA.n1978 VDDA.n1975 4.5005
R765 VDDA.n1979 VDDA.n1533 4.5005
R766 VDDA.n1983 VDDA.n1982 4.5005
R767 VDDA.n1984 VDDA.n1532 4.5005
R768 VDDA.n1988 VDDA.n1985 4.5005
R769 VDDA.n1989 VDDA.n1531 4.5005
R770 VDDA.n1993 VDDA.n1992 4.5005
R771 VDDA.n1994 VDDA.n1530 4.5005
R772 VDDA.n1998 VDDA.n1995 4.5005
R773 VDDA.n1999 VDDA.n1529 4.5005
R774 VDDA.n2003 VDDA.n2002 4.5005
R775 VDDA.n2004 VDDA.n1528 4.5005
R776 VDDA.n2008 VDDA.n2005 4.5005
R777 VDDA.n2009 VDDA.n1527 4.5005
R778 VDDA.n2013 VDDA.n2012 4.5005
R779 VDDA.n2014 VDDA.n1526 4.5005
R780 VDDA.n2018 VDDA.n2015 4.5005
R781 VDDA.n2019 VDDA.n1525 4.5005
R782 VDDA.n2023 VDDA.n2022 4.5005
R783 VDDA.n2024 VDDA.n1524 4.5005
R784 VDDA.n2028 VDDA.n2025 4.5005
R785 VDDA.n2029 VDDA.n1523 4.5005
R786 VDDA.n2033 VDDA.n2032 4.5005
R787 VDDA.n2034 VDDA.n1522 4.5005
R788 VDDA.n2038 VDDA.n2035 4.5005
R789 VDDA.n2039 VDDA.n1521 4.5005
R790 VDDA.n2043 VDDA.n2042 4.5005
R791 VDDA.n2044 VDDA.n1520 4.5005
R792 VDDA.n2048 VDDA.n2045 4.5005
R793 VDDA.n2049 VDDA.n1519 4.5005
R794 VDDA.n2053 VDDA.n2052 4.5005
R795 VDDA.n1612 VDDA.n1611 4.5005
R796 VDDA.n1615 VDDA.n1614 4.5005
R797 VDDA.n1616 VDDA.n1605 4.5005
R798 VDDA.n1620 VDDA.n1617 4.5005
R799 VDDA.n1621 VDDA.n1604 4.5005
R800 VDDA.n1625 VDDA.n1624 4.5005
R801 VDDA.n1626 VDDA.n1603 4.5005
R802 VDDA.n1630 VDDA.n1627 4.5005
R803 VDDA.n1631 VDDA.n1602 4.5005
R804 VDDA.n1635 VDDA.n1634 4.5005
R805 VDDA.n1636 VDDA.n1601 4.5005
R806 VDDA.n1640 VDDA.n1637 4.5005
R807 VDDA.n1641 VDDA.n1600 4.5005
R808 VDDA.n1645 VDDA.n1644 4.5005
R809 VDDA.n1646 VDDA.n1599 4.5005
R810 VDDA.n1650 VDDA.n1647 4.5005
R811 VDDA.n1651 VDDA.n1598 4.5005
R812 VDDA.n1655 VDDA.n1654 4.5005
R813 VDDA.n1656 VDDA.n1597 4.5005
R814 VDDA.n1660 VDDA.n1657 4.5005
R815 VDDA.n1661 VDDA.n1596 4.5005
R816 VDDA.n1665 VDDA.n1664 4.5005
R817 VDDA.n1666 VDDA.n1595 4.5005
R818 VDDA.n1670 VDDA.n1667 4.5005
R819 VDDA.n1671 VDDA.n1594 4.5005
R820 VDDA.n1675 VDDA.n1674 4.5005
R821 VDDA.n1676 VDDA.n1593 4.5005
R822 VDDA.n1680 VDDA.n1677 4.5005
R823 VDDA.n1681 VDDA.n1592 4.5005
R824 VDDA.n1685 VDDA.n1684 4.5005
R825 VDDA.n1686 VDDA.n1591 4.5005
R826 VDDA.n1690 VDDA.n1687 4.5005
R827 VDDA.n1691 VDDA.n1590 4.5005
R828 VDDA.n1695 VDDA.n1694 4.5005
R829 VDDA.n1696 VDDA.n1589 4.5005
R830 VDDA.n1700 VDDA.n1697 4.5005
R831 VDDA.n1701 VDDA.n1588 4.5005
R832 VDDA.n1705 VDDA.n1704 4.5005
R833 VDDA.n1706 VDDA.n1587 4.5005
R834 VDDA.n1710 VDDA.n1707 4.5005
R835 VDDA.n1711 VDDA.n1586 4.5005
R836 VDDA.n1715 VDDA.n1714 4.5005
R837 VDDA.n1716 VDDA.n1585 4.5005
R838 VDDA.n1720 VDDA.n1717 4.5005
R839 VDDA.n1721 VDDA.n1584 4.5005
R840 VDDA.n1725 VDDA.n1724 4.5005
R841 VDDA.n2095 VDDA.n2094 4.5005
R842 VDDA.n2161 VDDA.n2160 4.5005
R843 VDDA.n2238 VDDA.n2237 4.5005
R844 VDDA.n2288 VDDA.n2287 4.5005
R845 VDDA.n2292 VDDA.n2291 4.5005
R846 VDDA.n2293 VDDA.n2080 4.5005
R847 VDDA.n2297 VDDA.n2294 4.5005
R848 VDDA.n2298 VDDA.n2079 4.5005
R849 VDDA.n2302 VDDA.n2301 4.5005
R850 VDDA.n2303 VDDA.n2078 4.5005
R851 VDDA.n2307 VDDA.n2304 4.5005
R852 VDDA.n2308 VDDA.n2077 4.5005
R853 VDDA.n2312 VDDA.n2311 4.5005
R854 VDDA.n2313 VDDA.n2076 4.5005
R855 VDDA.n2317 VDDA.n2314 4.5005
R856 VDDA.n2318 VDDA.n2075 4.5005
R857 VDDA.n2322 VDDA.n2321 4.5005
R858 VDDA.n2323 VDDA.n2074 4.5005
R859 VDDA.n2327 VDDA.n2324 4.5005
R860 VDDA.n2328 VDDA.n2073 4.5005
R861 VDDA.n2332 VDDA.n2331 4.5005
R862 VDDA.n2333 VDDA.n2072 4.5005
R863 VDDA.n2337 VDDA.n2334 4.5005
R864 VDDA.n2338 VDDA.n2071 4.5005
R865 VDDA.n2342 VDDA.n2341 4.5005
R866 VDDA.n2343 VDDA.n2070 4.5005
R867 VDDA.n2347 VDDA.n2344 4.5005
R868 VDDA.n2348 VDDA.n2069 4.5005
R869 VDDA.n2352 VDDA.n2351 4.5005
R870 VDDA.n2353 VDDA.n2068 4.5005
R871 VDDA.n2357 VDDA.n2354 4.5005
R872 VDDA.n2358 VDDA.n2067 4.5005
R873 VDDA.n2362 VDDA.n2361 4.5005
R874 VDDA.n2363 VDDA.n2066 4.5005
R875 VDDA.n2367 VDDA.n2364 4.5005
R876 VDDA.n2368 VDDA.n2065 4.5005
R877 VDDA.n2372 VDDA.n2371 4.5005
R878 VDDA.n2373 VDDA.n2064 4.5005
R879 VDDA.n2377 VDDA.n2374 4.5005
R880 VDDA.n2378 VDDA.n2063 4.5005
R881 VDDA.n2382 VDDA.n2381 4.5005
R882 VDDA.n2383 VDDA.n2062 4.5005
R883 VDDA.n2387 VDDA.n2384 4.5005
R884 VDDA.n2388 VDDA.n2061 4.5005
R885 VDDA.n2392 VDDA.n2391 4.5005
R886 VDDA.n2393 VDDA.n2060 4.5005
R887 VDDA.n2397 VDDA.n2394 4.5005
R888 VDDA.n2398 VDDA.n2059 4.5005
R889 VDDA.n2402 VDDA.n2401 4.5005
R890 VDDA.n2479 VDDA.n2453 4.5005
R891 VDDA.n2464 VDDA.n2455 4.5005
R892 VDDA.n93 VDDA.n87 4.5005
R893 VDDA.n95 VDDA.n94 4.5005
R894 VDDA.n96 VDDA.n86 4.5005
R895 VDDA.n100 VDDA.n99 4.5005
R896 VDDA.n101 VDDA.n83 4.5005
R897 VDDA.n103 VDDA.n102 4.5005
R898 VDDA.n104 VDDA.n82 4.5005
R899 VDDA.n108 VDDA.n107 4.5005
R900 VDDA.n109 VDDA.n79 4.5005
R901 VDDA.n111 VDDA.n110 4.5005
R902 VDDA.n112 VDDA.n78 4.5005
R903 VDDA.n116 VDDA.n115 4.5005
R904 VDDA.n117 VDDA.n75 4.5005
R905 VDDA.n119 VDDA.n118 4.5005
R906 VDDA.n120 VDDA.n74 4.5005
R907 VDDA.n124 VDDA.n123 4.5005
R908 VDDA.n125 VDDA.n71 4.5005
R909 VDDA.n127 VDDA.n126 4.5005
R910 VDDA.n128 VDDA.n70 4.5005
R911 VDDA.n132 VDDA.n131 4.5005
R912 VDDA.n133 VDDA.n67 4.5005
R913 VDDA.n135 VDDA.n134 4.5005
R914 VDDA.n136 VDDA.n66 4.5005
R915 VDDA.n140 VDDA.n139 4.5005
R916 VDDA.n141 VDDA.n63 4.5005
R917 VDDA.n143 VDDA.n142 4.5005
R918 VDDA.n144 VDDA.n62 4.5005
R919 VDDA.n148 VDDA.n147 4.5005
R920 VDDA.n149 VDDA.n59 4.5005
R921 VDDA.n151 VDDA.n150 4.5005
R922 VDDA.n152 VDDA.n58 4.5005
R923 VDDA.n156 VDDA.n155 4.5005
R924 VDDA.n157 VDDA.n55 4.5005
R925 VDDA.n159 VDDA.n158 4.5005
R926 VDDA.n160 VDDA.n54 4.5005
R927 VDDA.n164 VDDA.n163 4.5005
R928 VDDA.n165 VDDA.n51 4.5005
R929 VDDA.n167 VDDA.n166 4.5005
R930 VDDA.n168 VDDA.n50 4.5005
R931 VDDA.n172 VDDA.n171 4.5005
R932 VDDA.n173 VDDA.n47 4.5005
R933 VDDA.n175 VDDA.n174 4.5005
R934 VDDA.n176 VDDA.n46 4.5005
R935 VDDA.n180 VDDA.n179 4.5005
R936 VDDA.n181 VDDA.n45 4.5005
R937 VDDA.n2935 VDDA.n2934 4.5005
R938 VDDA.n2804 VDDA.n2803 4.5005
R939 VDDA.n2814 VDDA.n2813 4.5005
R940 VDDA.n2815 VDDA.n2802 4.5005
R941 VDDA.n2817 VDDA.n2816 4.5005
R942 VDDA.n2800 VDDA.n2799 4.5005
R943 VDDA.n2824 VDDA.n2823 4.5005
R944 VDDA.n2825 VDDA.n2798 4.5005
R945 VDDA.n2827 VDDA.n2826 4.5005
R946 VDDA.n2796 VDDA.n2795 4.5005
R947 VDDA.n2834 VDDA.n2833 4.5005
R948 VDDA.n2835 VDDA.n2794 4.5005
R949 VDDA.n2837 VDDA.n2836 4.5005
R950 VDDA.n2792 VDDA.n2791 4.5005
R951 VDDA.n2844 VDDA.n2843 4.5005
R952 VDDA.n2845 VDDA.n2790 4.5005
R953 VDDA.n2847 VDDA.n2846 4.5005
R954 VDDA.n2788 VDDA.n2787 4.5005
R955 VDDA.n2854 VDDA.n2853 4.5005
R956 VDDA.n2855 VDDA.n2786 4.5005
R957 VDDA.n2857 VDDA.n2856 4.5005
R958 VDDA.n2784 VDDA.n2783 4.5005
R959 VDDA.n2864 VDDA.n2863 4.5005
R960 VDDA.n2865 VDDA.n2782 4.5005
R961 VDDA.n2867 VDDA.n2866 4.5005
R962 VDDA.n2780 VDDA.n2779 4.5005
R963 VDDA.n2874 VDDA.n2873 4.5005
R964 VDDA.n2875 VDDA.n2778 4.5005
R965 VDDA.n2877 VDDA.n2876 4.5005
R966 VDDA.n2776 VDDA.n2775 4.5005
R967 VDDA.n2884 VDDA.n2883 4.5005
R968 VDDA.n2885 VDDA.n2774 4.5005
R969 VDDA.n2887 VDDA.n2886 4.5005
R970 VDDA.n2772 VDDA.n2771 4.5005
R971 VDDA.n2894 VDDA.n2893 4.5005
R972 VDDA.n2895 VDDA.n2770 4.5005
R973 VDDA.n2897 VDDA.n2896 4.5005
R974 VDDA.n2768 VDDA.n2767 4.5005
R975 VDDA.n2904 VDDA.n2903 4.5005
R976 VDDA.n2905 VDDA.n2766 4.5005
R977 VDDA.n2907 VDDA.n2906 4.5005
R978 VDDA.n2764 VDDA.n2763 4.5005
R979 VDDA.n2914 VDDA.n2913 4.5005
R980 VDDA.n2915 VDDA.n2762 4.5005
R981 VDDA.n2917 VDDA.n2916 4.5005
R982 VDDA.n2760 VDDA.n2759 4.5005
R983 VDDA.n2923 VDDA.n2922 4.5005
R984 VDDA.n2659 VDDA.n2655 4.5005
R985 VDDA.n2663 VDDA.n2662 4.5005
R986 VDDA.n2664 VDDA.n2652 4.5005
R987 VDDA.n2666 VDDA.n2665 4.5005
R988 VDDA.n2667 VDDA.n2651 4.5005
R989 VDDA.n2671 VDDA.n2670 4.5005
R990 VDDA.n2672 VDDA.n2648 4.5005
R991 VDDA.n2674 VDDA.n2673 4.5005
R992 VDDA.n2675 VDDA.n2647 4.5005
R993 VDDA.n2679 VDDA.n2678 4.5005
R994 VDDA.n2680 VDDA.n2644 4.5005
R995 VDDA.n2682 VDDA.n2681 4.5005
R996 VDDA.n2683 VDDA.n2643 4.5005
R997 VDDA.n2687 VDDA.n2686 4.5005
R998 VDDA.n2688 VDDA.n2640 4.5005
R999 VDDA.n2690 VDDA.n2689 4.5005
R1000 VDDA.n2691 VDDA.n2639 4.5005
R1001 VDDA.n2695 VDDA.n2694 4.5005
R1002 VDDA.n2696 VDDA.n2636 4.5005
R1003 VDDA.n2698 VDDA.n2697 4.5005
R1004 VDDA.n2699 VDDA.n2635 4.5005
R1005 VDDA.n2703 VDDA.n2702 4.5005
R1006 VDDA.n2704 VDDA.n2632 4.5005
R1007 VDDA.n2706 VDDA.n2705 4.5005
R1008 VDDA.n2707 VDDA.n2631 4.5005
R1009 VDDA.n2711 VDDA.n2710 4.5005
R1010 VDDA.n2712 VDDA.n2628 4.5005
R1011 VDDA.n2714 VDDA.n2713 4.5005
R1012 VDDA.n2715 VDDA.n2627 4.5005
R1013 VDDA.n2719 VDDA.n2718 4.5005
R1014 VDDA.n2720 VDDA.n2624 4.5005
R1015 VDDA.n2722 VDDA.n2721 4.5005
R1016 VDDA.n2723 VDDA.n2623 4.5005
R1017 VDDA.n2727 VDDA.n2726 4.5005
R1018 VDDA.n2728 VDDA.n2620 4.5005
R1019 VDDA.n2730 VDDA.n2729 4.5005
R1020 VDDA.n2731 VDDA.n2619 4.5005
R1021 VDDA.n2735 VDDA.n2734 4.5005
R1022 VDDA.n2736 VDDA.n2616 4.5005
R1023 VDDA.n2738 VDDA.n2737 4.5005
R1024 VDDA.n2739 VDDA.n2615 4.5005
R1025 VDDA.n2743 VDDA.n2742 4.5005
R1026 VDDA.n2744 VDDA.n2614 4.5005
R1027 VDDA.n2746 VDDA.n2745 4.5005
R1028 VDDA.n195 VDDA.n194 4.5005
R1029 VDDA.n2752 VDDA.n2751 4.5005
R1030 VDDA.n271 VDDA.n265 4.5005
R1031 VDDA.n273 VDDA.n272 4.5005
R1032 VDDA.n274 VDDA.n264 4.5005
R1033 VDDA.n278 VDDA.n277 4.5005
R1034 VDDA.n279 VDDA.n261 4.5005
R1035 VDDA.n281 VDDA.n280 4.5005
R1036 VDDA.n282 VDDA.n260 4.5005
R1037 VDDA.n286 VDDA.n285 4.5005
R1038 VDDA.n287 VDDA.n257 4.5005
R1039 VDDA.n289 VDDA.n288 4.5005
R1040 VDDA.n290 VDDA.n256 4.5005
R1041 VDDA.n294 VDDA.n293 4.5005
R1042 VDDA.n295 VDDA.n253 4.5005
R1043 VDDA.n297 VDDA.n296 4.5005
R1044 VDDA.n298 VDDA.n252 4.5005
R1045 VDDA.n302 VDDA.n301 4.5005
R1046 VDDA.n303 VDDA.n249 4.5005
R1047 VDDA.n305 VDDA.n304 4.5005
R1048 VDDA.n306 VDDA.n248 4.5005
R1049 VDDA.n310 VDDA.n309 4.5005
R1050 VDDA.n311 VDDA.n245 4.5005
R1051 VDDA.n313 VDDA.n312 4.5005
R1052 VDDA.n314 VDDA.n244 4.5005
R1053 VDDA.n318 VDDA.n317 4.5005
R1054 VDDA.n319 VDDA.n241 4.5005
R1055 VDDA.n321 VDDA.n320 4.5005
R1056 VDDA.n322 VDDA.n240 4.5005
R1057 VDDA.n326 VDDA.n325 4.5005
R1058 VDDA.n327 VDDA.n237 4.5005
R1059 VDDA.n329 VDDA.n328 4.5005
R1060 VDDA.n330 VDDA.n236 4.5005
R1061 VDDA.n334 VDDA.n333 4.5005
R1062 VDDA.n335 VDDA.n233 4.5005
R1063 VDDA.n337 VDDA.n336 4.5005
R1064 VDDA.n338 VDDA.n232 4.5005
R1065 VDDA.n342 VDDA.n341 4.5005
R1066 VDDA.n343 VDDA.n229 4.5005
R1067 VDDA.n345 VDDA.n344 4.5005
R1068 VDDA.n346 VDDA.n228 4.5005
R1069 VDDA.n350 VDDA.n349 4.5005
R1070 VDDA.n351 VDDA.n225 4.5005
R1071 VDDA.n353 VDDA.n352 4.5005
R1072 VDDA.n354 VDDA.n224 4.5005
R1073 VDDA.n358 VDDA.n357 4.5005
R1074 VDDA.n359 VDDA.n223 4.5005
R1075 VDDA.n2587 VDDA.n2586 4.5005
R1076 VDDA.n2583 VDDA.n2582 4.5005
R1077 VDDA.n2581 VDDA.n192 4.5005
R1078 VDDA.n2582 VDDA.n2581 4.5005
R1079 VDDA.n2755 VDDA.n193 4.5005
R1080 VDDA.n2757 VDDA.n2756 4.5005
R1081 VDDA.n2756 VDDA.n2755 4.5005
R1082 VDDA.n2926 VDDA.n2758 4.5005
R1083 VDDA.n2928 VDDA.n2927 4.5005
R1084 VDDA.n2927 VDDA.n2926 4.5005
R1085 VDDA.n2929 VDDA.n183 4.5005
R1086 VDDA.n2931 VDDA.n2930 4.5005
R1087 VDDA.n2930 VDDA.n2929 4.5005
R1088 VDDA.n410 VDDA.n409 4.5005
R1089 VDDA.n420 VDDA.n419 4.5005
R1090 VDDA.n421 VDDA.n408 4.5005
R1091 VDDA.n423 VDDA.n422 4.5005
R1092 VDDA.n406 VDDA.n405 4.5005
R1093 VDDA.n430 VDDA.n429 4.5005
R1094 VDDA.n431 VDDA.n404 4.5005
R1095 VDDA.n433 VDDA.n432 4.5005
R1096 VDDA.n402 VDDA.n401 4.5005
R1097 VDDA.n440 VDDA.n439 4.5005
R1098 VDDA.n441 VDDA.n400 4.5005
R1099 VDDA.n443 VDDA.n442 4.5005
R1100 VDDA.n398 VDDA.n397 4.5005
R1101 VDDA.n450 VDDA.n449 4.5005
R1102 VDDA.n451 VDDA.n396 4.5005
R1103 VDDA.n453 VDDA.n452 4.5005
R1104 VDDA.n394 VDDA.n393 4.5005
R1105 VDDA.n460 VDDA.n459 4.5005
R1106 VDDA.n461 VDDA.n392 4.5005
R1107 VDDA.n463 VDDA.n462 4.5005
R1108 VDDA.n390 VDDA.n389 4.5005
R1109 VDDA.n470 VDDA.n469 4.5005
R1110 VDDA.n471 VDDA.n388 4.5005
R1111 VDDA.n473 VDDA.n472 4.5005
R1112 VDDA.n386 VDDA.n385 4.5005
R1113 VDDA.n480 VDDA.n479 4.5005
R1114 VDDA.n481 VDDA.n384 4.5005
R1115 VDDA.n483 VDDA.n482 4.5005
R1116 VDDA.n382 VDDA.n381 4.5005
R1117 VDDA.n490 VDDA.n489 4.5005
R1118 VDDA.n491 VDDA.n380 4.5005
R1119 VDDA.n493 VDDA.n492 4.5005
R1120 VDDA.n378 VDDA.n377 4.5005
R1121 VDDA.n500 VDDA.n499 4.5005
R1122 VDDA.n501 VDDA.n376 4.5005
R1123 VDDA.n503 VDDA.n502 4.5005
R1124 VDDA.n374 VDDA.n373 4.5005
R1125 VDDA.n510 VDDA.n509 4.5005
R1126 VDDA.n511 VDDA.n372 4.5005
R1127 VDDA.n513 VDDA.n512 4.5005
R1128 VDDA.n370 VDDA.n369 4.5005
R1129 VDDA.n520 VDDA.n519 4.5005
R1130 VDDA.n521 VDDA.n368 4.5005
R1131 VDDA.n523 VDDA.n522 4.5005
R1132 VDDA.n366 VDDA.n365 4.5005
R1133 VDDA.n529 VDDA.n528 4.5005
R1134 VDDA.n530 VDDA.n364 4.5005
R1135 VDDA.n2570 VDDA.n532 4.5005
R1136 VDDA.n2572 VDDA.n2571 4.5005
R1137 VDDA.n2571 VDDA.n2570 4.5005
R1138 VDDA.n2510 VDDA.n2509 4.5005
R1139 VDDA.n2516 VDDA.n538 4.5005
R1140 VDDA.n2519 VDDA.n2518 4.5005
R1141 VDDA.n2522 VDDA.n2521 4.5005
R1142 VDDA.n2514 VDDA.n2494 4.5005
R1143 VDDA.n2515 VDDA.n540 4.5005
R1144 VDDA.n2515 VDDA.n2514 4.5005
R1145 VDDA.n2483 VDDA.n2451 4.5005
R1146 VDDA.n2486 VDDA.n2485 4.5005
R1147 VDDA.n561 VDDA.n560 4.5005
R1148 VDDA.n562 VDDA.n546 4.5005
R1149 VDDA.n569 VDDA.n568 4.5005
R1150 VDDA.n572 VDDA.n571 4.5005
R1151 VDDA.n2435 VDDA.n564 4.5005
R1152 VDDA.n2437 VDDA.n2436 4.5005
R1153 VDDA.n2436 VDDA.n2435 4.5005
R1154 VDDA.n1379 VDDA.n1375 4.5005
R1155 VDDA.n1383 VDDA.n1382 4.5005
R1156 VDDA.n1384 VDDA.n1372 4.5005
R1157 VDDA.n1386 VDDA.n1385 4.5005
R1158 VDDA.n1387 VDDA.n1371 4.5005
R1159 VDDA.n1391 VDDA.n1390 4.5005
R1160 VDDA.n1392 VDDA.n1368 4.5005
R1161 VDDA.n1394 VDDA.n1393 4.5005
R1162 VDDA.n1395 VDDA.n1367 4.5005
R1163 VDDA.n1399 VDDA.n1398 4.5005
R1164 VDDA.n1400 VDDA.n1364 4.5005
R1165 VDDA.n1402 VDDA.n1401 4.5005
R1166 VDDA.n1403 VDDA.n1363 4.5005
R1167 VDDA.n1407 VDDA.n1406 4.5005
R1168 VDDA.n1408 VDDA.n1360 4.5005
R1169 VDDA.n1410 VDDA.n1409 4.5005
R1170 VDDA.n1411 VDDA.n1359 4.5005
R1171 VDDA.n1415 VDDA.n1414 4.5005
R1172 VDDA.n1416 VDDA.n1356 4.5005
R1173 VDDA.n1418 VDDA.n1417 4.5005
R1174 VDDA.n1419 VDDA.n1355 4.5005
R1175 VDDA.n1423 VDDA.n1422 4.5005
R1176 VDDA.n1424 VDDA.n1352 4.5005
R1177 VDDA.n1426 VDDA.n1425 4.5005
R1178 VDDA.n1427 VDDA.n1351 4.5005
R1179 VDDA.n1431 VDDA.n1430 4.5005
R1180 VDDA.n1432 VDDA.n1348 4.5005
R1181 VDDA.n1434 VDDA.n1433 4.5005
R1182 VDDA.n1435 VDDA.n1347 4.5005
R1183 VDDA.n1439 VDDA.n1438 4.5005
R1184 VDDA.n1440 VDDA.n1344 4.5005
R1185 VDDA.n1442 VDDA.n1441 4.5005
R1186 VDDA.n1443 VDDA.n1343 4.5005
R1187 VDDA.n1447 VDDA.n1446 4.5005
R1188 VDDA.n1448 VDDA.n1340 4.5005
R1189 VDDA.n1450 VDDA.n1449 4.5005
R1190 VDDA.n1451 VDDA.n1339 4.5005
R1191 VDDA.n1455 VDDA.n1454 4.5005
R1192 VDDA.n1456 VDDA.n1336 4.5005
R1193 VDDA.n1458 VDDA.n1457 4.5005
R1194 VDDA.n1459 VDDA.n1335 4.5005
R1195 VDDA.n1463 VDDA.n1462 4.5005
R1196 VDDA.n1464 VDDA.n1334 4.5005
R1197 VDDA.n1466 VDDA.n1465 4.5005
R1198 VDDA.n610 VDDA.n609 4.5005
R1199 VDDA.n2409 VDDA.n2408 4.5005
R1200 VDDA.n2415 VDDA.n603 4.5005
R1201 VDDA.n686 VDDA.n680 4.5005
R1202 VDDA.n688 VDDA.n687 4.5005
R1203 VDDA.n689 VDDA.n679 4.5005
R1204 VDDA.n693 VDDA.n692 4.5005
R1205 VDDA.n694 VDDA.n676 4.5005
R1206 VDDA.n696 VDDA.n695 4.5005
R1207 VDDA.n697 VDDA.n675 4.5005
R1208 VDDA.n701 VDDA.n700 4.5005
R1209 VDDA.n702 VDDA.n672 4.5005
R1210 VDDA.n704 VDDA.n703 4.5005
R1211 VDDA.n705 VDDA.n671 4.5005
R1212 VDDA.n709 VDDA.n708 4.5005
R1213 VDDA.n710 VDDA.n668 4.5005
R1214 VDDA.n712 VDDA.n711 4.5005
R1215 VDDA.n713 VDDA.n667 4.5005
R1216 VDDA.n717 VDDA.n716 4.5005
R1217 VDDA.n718 VDDA.n664 4.5005
R1218 VDDA.n720 VDDA.n719 4.5005
R1219 VDDA.n721 VDDA.n663 4.5005
R1220 VDDA.n725 VDDA.n724 4.5005
R1221 VDDA.n726 VDDA.n660 4.5005
R1222 VDDA.n728 VDDA.n727 4.5005
R1223 VDDA.n729 VDDA.n659 4.5005
R1224 VDDA.n733 VDDA.n732 4.5005
R1225 VDDA.n734 VDDA.n656 4.5005
R1226 VDDA.n736 VDDA.n735 4.5005
R1227 VDDA.n737 VDDA.n655 4.5005
R1228 VDDA.n741 VDDA.n740 4.5005
R1229 VDDA.n742 VDDA.n652 4.5005
R1230 VDDA.n744 VDDA.n743 4.5005
R1231 VDDA.n745 VDDA.n651 4.5005
R1232 VDDA.n749 VDDA.n748 4.5005
R1233 VDDA.n750 VDDA.n648 4.5005
R1234 VDDA.n752 VDDA.n751 4.5005
R1235 VDDA.n753 VDDA.n647 4.5005
R1236 VDDA.n757 VDDA.n756 4.5005
R1237 VDDA.n758 VDDA.n644 4.5005
R1238 VDDA.n760 VDDA.n759 4.5005
R1239 VDDA.n761 VDDA.n643 4.5005
R1240 VDDA.n765 VDDA.n764 4.5005
R1241 VDDA.n766 VDDA.n640 4.5005
R1242 VDDA.n768 VDDA.n767 4.5005
R1243 VDDA.n769 VDDA.n639 4.5005
R1244 VDDA.n773 VDDA.n772 4.5005
R1245 VDDA.n774 VDDA.n638 4.5005
R1246 VDDA.n1307 VDDA.n1306 4.5005
R1247 VDDA.n1176 VDDA.n1175 4.5005
R1248 VDDA.n1186 VDDA.n1185 4.5005
R1249 VDDA.n1187 VDDA.n1174 4.5005
R1250 VDDA.n1189 VDDA.n1188 4.5005
R1251 VDDA.n1172 VDDA.n1171 4.5005
R1252 VDDA.n1196 VDDA.n1195 4.5005
R1253 VDDA.n1197 VDDA.n1170 4.5005
R1254 VDDA.n1199 VDDA.n1198 4.5005
R1255 VDDA.n1168 VDDA.n1167 4.5005
R1256 VDDA.n1206 VDDA.n1205 4.5005
R1257 VDDA.n1207 VDDA.n1166 4.5005
R1258 VDDA.n1209 VDDA.n1208 4.5005
R1259 VDDA.n1164 VDDA.n1163 4.5005
R1260 VDDA.n1216 VDDA.n1215 4.5005
R1261 VDDA.n1217 VDDA.n1162 4.5005
R1262 VDDA.n1219 VDDA.n1218 4.5005
R1263 VDDA.n1160 VDDA.n1159 4.5005
R1264 VDDA.n1226 VDDA.n1225 4.5005
R1265 VDDA.n1227 VDDA.n1158 4.5005
R1266 VDDA.n1229 VDDA.n1228 4.5005
R1267 VDDA.n1156 VDDA.n1155 4.5005
R1268 VDDA.n1236 VDDA.n1235 4.5005
R1269 VDDA.n1237 VDDA.n1154 4.5005
R1270 VDDA.n1239 VDDA.n1238 4.5005
R1271 VDDA.n1152 VDDA.n1151 4.5005
R1272 VDDA.n1246 VDDA.n1245 4.5005
R1273 VDDA.n1247 VDDA.n1150 4.5005
R1274 VDDA.n1249 VDDA.n1248 4.5005
R1275 VDDA.n1148 VDDA.n1147 4.5005
R1276 VDDA.n1256 VDDA.n1255 4.5005
R1277 VDDA.n1257 VDDA.n1146 4.5005
R1278 VDDA.n1259 VDDA.n1258 4.5005
R1279 VDDA.n1144 VDDA.n1143 4.5005
R1280 VDDA.n1266 VDDA.n1265 4.5005
R1281 VDDA.n1267 VDDA.n1142 4.5005
R1282 VDDA.n1269 VDDA.n1268 4.5005
R1283 VDDA.n1140 VDDA.n1139 4.5005
R1284 VDDA.n1276 VDDA.n1275 4.5005
R1285 VDDA.n1277 VDDA.n1138 4.5005
R1286 VDDA.n1279 VDDA.n1278 4.5005
R1287 VDDA.n1136 VDDA.n1135 4.5005
R1288 VDDA.n1286 VDDA.n1285 4.5005
R1289 VDDA.n1287 VDDA.n1134 4.5005
R1290 VDDA.n1289 VDDA.n1288 4.5005
R1291 VDDA.n1132 VDDA.n1131 4.5005
R1292 VDDA.n1295 VDDA.n1294 4.5005
R1293 VDDA.n1031 VDDA.n1027 4.5005
R1294 VDDA.n1035 VDDA.n1034 4.5005
R1295 VDDA.n1036 VDDA.n1024 4.5005
R1296 VDDA.n1038 VDDA.n1037 4.5005
R1297 VDDA.n1039 VDDA.n1023 4.5005
R1298 VDDA.n1043 VDDA.n1042 4.5005
R1299 VDDA.n1044 VDDA.n1020 4.5005
R1300 VDDA.n1046 VDDA.n1045 4.5005
R1301 VDDA.n1047 VDDA.n1019 4.5005
R1302 VDDA.n1051 VDDA.n1050 4.5005
R1303 VDDA.n1052 VDDA.n1016 4.5005
R1304 VDDA.n1054 VDDA.n1053 4.5005
R1305 VDDA.n1055 VDDA.n1015 4.5005
R1306 VDDA.n1059 VDDA.n1058 4.5005
R1307 VDDA.n1060 VDDA.n1012 4.5005
R1308 VDDA.n1062 VDDA.n1061 4.5005
R1309 VDDA.n1063 VDDA.n1011 4.5005
R1310 VDDA.n1067 VDDA.n1066 4.5005
R1311 VDDA.n1068 VDDA.n1008 4.5005
R1312 VDDA.n1070 VDDA.n1069 4.5005
R1313 VDDA.n1071 VDDA.n1007 4.5005
R1314 VDDA.n1075 VDDA.n1074 4.5005
R1315 VDDA.n1076 VDDA.n1004 4.5005
R1316 VDDA.n1078 VDDA.n1077 4.5005
R1317 VDDA.n1079 VDDA.n1003 4.5005
R1318 VDDA.n1083 VDDA.n1082 4.5005
R1319 VDDA.n1084 VDDA.n1000 4.5005
R1320 VDDA.n1086 VDDA.n1085 4.5005
R1321 VDDA.n1087 VDDA.n999 4.5005
R1322 VDDA.n1091 VDDA.n1090 4.5005
R1323 VDDA.n1092 VDDA.n996 4.5005
R1324 VDDA.n1094 VDDA.n1093 4.5005
R1325 VDDA.n1095 VDDA.n995 4.5005
R1326 VDDA.n1099 VDDA.n1098 4.5005
R1327 VDDA.n1100 VDDA.n992 4.5005
R1328 VDDA.n1102 VDDA.n1101 4.5005
R1329 VDDA.n1103 VDDA.n991 4.5005
R1330 VDDA.n1107 VDDA.n1106 4.5005
R1331 VDDA.n1108 VDDA.n988 4.5005
R1332 VDDA.n1110 VDDA.n1109 4.5005
R1333 VDDA.n1111 VDDA.n987 4.5005
R1334 VDDA.n1115 VDDA.n1114 4.5005
R1335 VDDA.n1116 VDDA.n986 4.5005
R1336 VDDA.n1118 VDDA.n1117 4.5005
R1337 VDDA.n787 VDDA.n786 4.5005
R1338 VDDA.n1124 VDDA.n1123 4.5005
R1339 VDDA.n1127 VDDA.n785 4.5005
R1340 VDDA.n1129 VDDA.n1128 4.5005
R1341 VDDA.n1128 VDDA.n1127 4.5005
R1342 VDDA.n1298 VDDA.n1130 4.5005
R1343 VDDA.n1300 VDDA.n1299 4.5005
R1344 VDDA.n1299 VDDA.n1298 4.5005
R1345 VDDA.n1303 VDDA.n1302 4.5005
R1346 VDDA.n1301 VDDA.n606 4.5005
R1347 VDDA.n1302 VDDA.n1301 4.5005
R1348 VDDA.n2413 VDDA.n607 4.5005
R1349 VDDA.n2414 VDDA.n605 4.5005
R1350 VDDA.n2414 VDDA.n2413 4.5005
R1351 VDDA.n955 VDDA.n952 4.5005
R1352 VDDA.n840 VDDA.n836 4.5005
R1353 VDDA.n844 VDDA.n841 4.5005
R1354 VDDA.n845 VDDA.n835 4.5005
R1355 VDDA.n849 VDDA.n848 4.5005
R1356 VDDA.n850 VDDA.n834 4.5005
R1357 VDDA.n854 VDDA.n851 4.5005
R1358 VDDA.n855 VDDA.n833 4.5005
R1359 VDDA.n859 VDDA.n858 4.5005
R1360 VDDA.n860 VDDA.n832 4.5005
R1361 VDDA.n864 VDDA.n861 4.5005
R1362 VDDA.n865 VDDA.n831 4.5005
R1363 VDDA.n869 VDDA.n868 4.5005
R1364 VDDA.n870 VDDA.n830 4.5005
R1365 VDDA.n874 VDDA.n871 4.5005
R1366 VDDA.n875 VDDA.n829 4.5005
R1367 VDDA.n879 VDDA.n878 4.5005
R1368 VDDA.n880 VDDA.n828 4.5005
R1369 VDDA.n884 VDDA.n881 4.5005
R1370 VDDA.n885 VDDA.n827 4.5005
R1371 VDDA.n889 VDDA.n888 4.5005
R1372 VDDA.n890 VDDA.n826 4.5005
R1373 VDDA.n894 VDDA.n891 4.5005
R1374 VDDA.n895 VDDA.n825 4.5005
R1375 VDDA.n899 VDDA.n898 4.5005
R1376 VDDA.n900 VDDA.n824 4.5005
R1377 VDDA.n904 VDDA.n901 4.5005
R1378 VDDA.n905 VDDA.n823 4.5005
R1379 VDDA.n909 VDDA.n908 4.5005
R1380 VDDA.n910 VDDA.n822 4.5005
R1381 VDDA.n914 VDDA.n911 4.5005
R1382 VDDA.n915 VDDA.n821 4.5005
R1383 VDDA.n919 VDDA.n918 4.5005
R1384 VDDA.n920 VDDA.n820 4.5005
R1385 VDDA.n924 VDDA.n921 4.5005
R1386 VDDA.n925 VDDA.n819 4.5005
R1387 VDDA.n929 VDDA.n928 4.5005
R1388 VDDA.n930 VDDA.n818 4.5005
R1389 VDDA.n934 VDDA.n931 4.5005
R1390 VDDA.n935 VDDA.n817 4.5005
R1391 VDDA.n939 VDDA.n938 4.5005
R1392 VDDA.n940 VDDA.n816 4.5005
R1393 VDDA.n944 VDDA.n941 4.5005
R1394 VDDA.n945 VDDA.n815 4.5005
R1395 VDDA.n949 VDDA.n948 4.5005
R1396 VDDA.n950 VDDA.n814 4.5005
R1397 VDDA.n959 VDDA.n958 4.5005
R1398 VDDA.n2144 VDDA.n2143 4.48641
R1399 VDDA.n2143 VDDA.n2121 4.48641
R1400 VDDA.n2154 VDDA.n2153 4.48641
R1401 VDDA.n2153 VDDA.n2101 4.48641
R1402 VDDA.n1922 VDDA.n1549 3.75335
R1403 VDDA.n1921 VDDA.n1920 3.75335
R1404 VDDA.n1929 VDDA.n1927 3.75335
R1405 VDDA.n1928 VDDA.n1543 3.75335
R1406 VDDA.n2213 VDDA.n2204 3.75335
R1407 VDDA.n2207 VDDA.n2174 3.75335
R1408 VDDA.n2195 VDDA.n2181 3.75335
R1409 VDDA.n2187 VDDA.n2186 3.75335
R1410 VDDA.n2055 VDDA.n2054 3.48486
R1411 VDDA.n1727 VDDA.n1726 3.47821
R1412 VDDA.n2404 VDDA.n2403 3.47821
R1413 VDDA.n92 VDDA.n20 3.47821
R1414 VDDA.n2806 VDDA.n2805 3.47821
R1415 VDDA.n2656 VDDA.n2590 3.47821
R1416 VDDA.n270 VDDA.n198 3.47821
R1417 VDDA.n412 VDDA.n411 3.47821
R1418 VDDA.n1376 VDDA.n1310 3.47821
R1419 VDDA.n685 VDDA.n613 3.47821
R1420 VDDA.n1178 VDDA.n1177 3.47821
R1421 VDDA.n1028 VDDA.n962 3.47821
R1422 VDDA.n839 VDDA.n789 3.47821
R1423 VDDA.n2140 VDDA.n2139 3.41464
R1424 VDDA.n2150 VDDA.n2149 3.41464
R1425 VDDA.n1518 VDDA.n1517 3.4105
R1426 VDDA.n2052 VDDA.n2051 3.4105
R1427 VDDA.n2050 VDDA.n2049 3.4105
R1428 VDDA.n2048 VDDA.n2047 3.4105
R1429 VDDA.n2046 VDDA.n1520 3.4105
R1430 VDDA.n2042 VDDA.n2041 3.4105
R1431 VDDA.n2040 VDDA.n2039 3.4105
R1432 VDDA.n2038 VDDA.n2037 3.4105
R1433 VDDA.n2036 VDDA.n1522 3.4105
R1434 VDDA.n2032 VDDA.n2031 3.4105
R1435 VDDA.n2030 VDDA.n2029 3.4105
R1436 VDDA.n2028 VDDA.n2027 3.4105
R1437 VDDA.n2026 VDDA.n1524 3.4105
R1438 VDDA.n2022 VDDA.n2021 3.4105
R1439 VDDA.n2020 VDDA.n2019 3.4105
R1440 VDDA.n2018 VDDA.n2017 3.4105
R1441 VDDA.n2016 VDDA.n1526 3.4105
R1442 VDDA.n2012 VDDA.n2011 3.4105
R1443 VDDA.n2010 VDDA.n2009 3.4105
R1444 VDDA.n2008 VDDA.n2007 3.4105
R1445 VDDA.n2006 VDDA.n1528 3.4105
R1446 VDDA.n2002 VDDA.n2001 3.4105
R1447 VDDA.n2000 VDDA.n1999 3.4105
R1448 VDDA.n1998 VDDA.n1997 3.4105
R1449 VDDA.n1996 VDDA.n1530 3.4105
R1450 VDDA.n1992 VDDA.n1991 3.4105
R1451 VDDA.n1990 VDDA.n1989 3.4105
R1452 VDDA.n1988 VDDA.n1987 3.4105
R1453 VDDA.n1986 VDDA.n1532 3.4105
R1454 VDDA.n1982 VDDA.n1981 3.4105
R1455 VDDA.n1980 VDDA.n1979 3.4105
R1456 VDDA.n1978 VDDA.n1977 3.4105
R1457 VDDA.n1976 VDDA.n1534 3.4105
R1458 VDDA.n1972 VDDA.n1971 3.4105
R1459 VDDA.n1970 VDDA.n1969 3.4105
R1460 VDDA.n1968 VDDA.n1967 3.4105
R1461 VDDA.n1966 VDDA.n1536 3.4105
R1462 VDDA.n1962 VDDA.n1961 3.4105
R1463 VDDA.n1960 VDDA.n1959 3.4105
R1464 VDDA.n1958 VDDA.n1957 3.4105
R1465 VDDA.n1956 VDDA.n1538 3.4105
R1466 VDDA.n1952 VDDA.n1951 3.4105
R1467 VDDA.n1950 VDDA.n1949 3.4105
R1468 VDDA.n1948 VDDA.n1947 3.4105
R1469 VDDA.n1946 VDDA.n1540 3.4105
R1470 VDDA.n1942 VDDA.n1941 3.4105
R1471 VDDA.n1940 VDDA.n1492 3.4105
R1472 VDDA.n1583 VDDA.n1582 3.4105
R1473 VDDA.n1724 VDDA.n1723 3.4105
R1474 VDDA.n1722 VDDA.n1721 3.4105
R1475 VDDA.n1720 VDDA.n1719 3.4105
R1476 VDDA.n1718 VDDA.n1585 3.4105
R1477 VDDA.n1714 VDDA.n1713 3.4105
R1478 VDDA.n1712 VDDA.n1711 3.4105
R1479 VDDA.n1710 VDDA.n1709 3.4105
R1480 VDDA.n1708 VDDA.n1587 3.4105
R1481 VDDA.n1704 VDDA.n1703 3.4105
R1482 VDDA.n1702 VDDA.n1701 3.4105
R1483 VDDA.n1700 VDDA.n1699 3.4105
R1484 VDDA.n1698 VDDA.n1589 3.4105
R1485 VDDA.n1694 VDDA.n1693 3.4105
R1486 VDDA.n1692 VDDA.n1691 3.4105
R1487 VDDA.n1690 VDDA.n1689 3.4105
R1488 VDDA.n1688 VDDA.n1591 3.4105
R1489 VDDA.n1684 VDDA.n1683 3.4105
R1490 VDDA.n1682 VDDA.n1681 3.4105
R1491 VDDA.n1680 VDDA.n1679 3.4105
R1492 VDDA.n1678 VDDA.n1593 3.4105
R1493 VDDA.n1674 VDDA.n1673 3.4105
R1494 VDDA.n1672 VDDA.n1671 3.4105
R1495 VDDA.n1670 VDDA.n1669 3.4105
R1496 VDDA.n1668 VDDA.n1595 3.4105
R1497 VDDA.n1664 VDDA.n1663 3.4105
R1498 VDDA.n1662 VDDA.n1661 3.4105
R1499 VDDA.n1660 VDDA.n1659 3.4105
R1500 VDDA.n1658 VDDA.n1597 3.4105
R1501 VDDA.n1654 VDDA.n1653 3.4105
R1502 VDDA.n1652 VDDA.n1651 3.4105
R1503 VDDA.n1650 VDDA.n1649 3.4105
R1504 VDDA.n1648 VDDA.n1599 3.4105
R1505 VDDA.n1644 VDDA.n1643 3.4105
R1506 VDDA.n1642 VDDA.n1641 3.4105
R1507 VDDA.n1640 VDDA.n1639 3.4105
R1508 VDDA.n1638 VDDA.n1601 3.4105
R1509 VDDA.n1634 VDDA.n1633 3.4105
R1510 VDDA.n1632 VDDA.n1631 3.4105
R1511 VDDA.n1630 VDDA.n1629 3.4105
R1512 VDDA.n1628 VDDA.n1603 3.4105
R1513 VDDA.n1624 VDDA.n1623 3.4105
R1514 VDDA.n1622 VDDA.n1621 3.4105
R1515 VDDA.n1620 VDDA.n1619 3.4105
R1516 VDDA.n1618 VDDA.n1605 3.4105
R1517 VDDA.n1614 VDDA.n1613 3.4105
R1518 VDDA.n1612 VDDA.n1558 3.4105
R1519 VDDA.n2058 VDDA.n2057 3.4105
R1520 VDDA.n2401 VDDA.n2400 3.4105
R1521 VDDA.n2399 VDDA.n2398 3.4105
R1522 VDDA.n2397 VDDA.n2396 3.4105
R1523 VDDA.n2395 VDDA.n2060 3.4105
R1524 VDDA.n2391 VDDA.n2390 3.4105
R1525 VDDA.n2389 VDDA.n2388 3.4105
R1526 VDDA.n2387 VDDA.n2386 3.4105
R1527 VDDA.n2385 VDDA.n2062 3.4105
R1528 VDDA.n2381 VDDA.n2380 3.4105
R1529 VDDA.n2379 VDDA.n2378 3.4105
R1530 VDDA.n2377 VDDA.n2376 3.4105
R1531 VDDA.n2375 VDDA.n2064 3.4105
R1532 VDDA.n2371 VDDA.n2370 3.4105
R1533 VDDA.n2369 VDDA.n2368 3.4105
R1534 VDDA.n2367 VDDA.n2366 3.4105
R1535 VDDA.n2365 VDDA.n2066 3.4105
R1536 VDDA.n2361 VDDA.n2360 3.4105
R1537 VDDA.n2359 VDDA.n2358 3.4105
R1538 VDDA.n2357 VDDA.n2356 3.4105
R1539 VDDA.n2355 VDDA.n2068 3.4105
R1540 VDDA.n2351 VDDA.n2350 3.4105
R1541 VDDA.n2349 VDDA.n2348 3.4105
R1542 VDDA.n2347 VDDA.n2346 3.4105
R1543 VDDA.n2345 VDDA.n2070 3.4105
R1544 VDDA.n2341 VDDA.n2340 3.4105
R1545 VDDA.n2339 VDDA.n2338 3.4105
R1546 VDDA.n2337 VDDA.n2336 3.4105
R1547 VDDA.n2335 VDDA.n2072 3.4105
R1548 VDDA.n2331 VDDA.n2330 3.4105
R1549 VDDA.n2329 VDDA.n2328 3.4105
R1550 VDDA.n2327 VDDA.n2326 3.4105
R1551 VDDA.n2325 VDDA.n2074 3.4105
R1552 VDDA.n2321 VDDA.n2320 3.4105
R1553 VDDA.n2319 VDDA.n2318 3.4105
R1554 VDDA.n2317 VDDA.n2316 3.4105
R1555 VDDA.n2315 VDDA.n2076 3.4105
R1556 VDDA.n2311 VDDA.n2310 3.4105
R1557 VDDA.n2309 VDDA.n2308 3.4105
R1558 VDDA.n2307 VDDA.n2306 3.4105
R1559 VDDA.n2305 VDDA.n2078 3.4105
R1560 VDDA.n2301 VDDA.n2300 3.4105
R1561 VDDA.n2299 VDDA.n2298 3.4105
R1562 VDDA.n2297 VDDA.n2296 3.4105
R1563 VDDA.n2295 VDDA.n2080 3.4105
R1564 VDDA.n45 VDDA.n44 3.4105
R1565 VDDA.n179 VDDA.n178 3.4105
R1566 VDDA.n177 VDDA.n176 3.4105
R1567 VDDA.n175 VDDA.n49 3.4105
R1568 VDDA.n48 VDDA.n47 3.4105
R1569 VDDA.n171 VDDA.n170 3.4105
R1570 VDDA.n169 VDDA.n168 3.4105
R1571 VDDA.n167 VDDA.n53 3.4105
R1572 VDDA.n52 VDDA.n51 3.4105
R1573 VDDA.n163 VDDA.n162 3.4105
R1574 VDDA.n161 VDDA.n160 3.4105
R1575 VDDA.n159 VDDA.n57 3.4105
R1576 VDDA.n56 VDDA.n55 3.4105
R1577 VDDA.n155 VDDA.n154 3.4105
R1578 VDDA.n153 VDDA.n152 3.4105
R1579 VDDA.n151 VDDA.n61 3.4105
R1580 VDDA.n60 VDDA.n59 3.4105
R1581 VDDA.n147 VDDA.n146 3.4105
R1582 VDDA.n145 VDDA.n144 3.4105
R1583 VDDA.n143 VDDA.n65 3.4105
R1584 VDDA.n64 VDDA.n63 3.4105
R1585 VDDA.n139 VDDA.n138 3.4105
R1586 VDDA.n137 VDDA.n136 3.4105
R1587 VDDA.n135 VDDA.n69 3.4105
R1588 VDDA.n68 VDDA.n67 3.4105
R1589 VDDA.n131 VDDA.n130 3.4105
R1590 VDDA.n129 VDDA.n128 3.4105
R1591 VDDA.n127 VDDA.n73 3.4105
R1592 VDDA.n72 VDDA.n71 3.4105
R1593 VDDA.n123 VDDA.n122 3.4105
R1594 VDDA.n121 VDDA.n120 3.4105
R1595 VDDA.n119 VDDA.n77 3.4105
R1596 VDDA.n76 VDDA.n75 3.4105
R1597 VDDA.n115 VDDA.n114 3.4105
R1598 VDDA.n113 VDDA.n112 3.4105
R1599 VDDA.n111 VDDA.n81 3.4105
R1600 VDDA.n80 VDDA.n79 3.4105
R1601 VDDA.n107 VDDA.n106 3.4105
R1602 VDDA.n105 VDDA.n104 3.4105
R1603 VDDA.n103 VDDA.n85 3.4105
R1604 VDDA.n84 VDDA.n83 3.4105
R1605 VDDA.n99 VDDA.n98 3.4105
R1606 VDDA.n97 VDDA.n96 3.4105
R1607 VDDA.n95 VDDA.n89 3.4105
R1608 VDDA.n88 VDDA.n87 3.4105
R1609 VDDA.n91 VDDA.n90 3.4105
R1610 VDDA.n2936 VDDA.n2935 3.4105
R1611 VDDA.n2920 VDDA.n2760 3.4105
R1612 VDDA.n2918 VDDA.n2917 3.4105
R1613 VDDA.n2762 VDDA.n2761 3.4105
R1614 VDDA.n2913 VDDA.n2912 3.4105
R1615 VDDA.n2910 VDDA.n2764 3.4105
R1616 VDDA.n2908 VDDA.n2907 3.4105
R1617 VDDA.n2766 VDDA.n2765 3.4105
R1618 VDDA.n2903 VDDA.n2902 3.4105
R1619 VDDA.n2900 VDDA.n2768 3.4105
R1620 VDDA.n2898 VDDA.n2897 3.4105
R1621 VDDA.n2770 VDDA.n2769 3.4105
R1622 VDDA.n2893 VDDA.n2892 3.4105
R1623 VDDA.n2890 VDDA.n2772 3.4105
R1624 VDDA.n2888 VDDA.n2887 3.4105
R1625 VDDA.n2774 VDDA.n2773 3.4105
R1626 VDDA.n2883 VDDA.n2882 3.4105
R1627 VDDA.n2880 VDDA.n2776 3.4105
R1628 VDDA.n2878 VDDA.n2877 3.4105
R1629 VDDA.n2778 VDDA.n2777 3.4105
R1630 VDDA.n2873 VDDA.n2872 3.4105
R1631 VDDA.n2870 VDDA.n2780 3.4105
R1632 VDDA.n2868 VDDA.n2867 3.4105
R1633 VDDA.n2782 VDDA.n2781 3.4105
R1634 VDDA.n2863 VDDA.n2862 3.4105
R1635 VDDA.n2860 VDDA.n2784 3.4105
R1636 VDDA.n2858 VDDA.n2857 3.4105
R1637 VDDA.n2786 VDDA.n2785 3.4105
R1638 VDDA.n2853 VDDA.n2852 3.4105
R1639 VDDA.n2850 VDDA.n2788 3.4105
R1640 VDDA.n2848 VDDA.n2847 3.4105
R1641 VDDA.n2790 VDDA.n2789 3.4105
R1642 VDDA.n2843 VDDA.n2842 3.4105
R1643 VDDA.n2840 VDDA.n2792 3.4105
R1644 VDDA.n2838 VDDA.n2837 3.4105
R1645 VDDA.n2794 VDDA.n2793 3.4105
R1646 VDDA.n2833 VDDA.n2832 3.4105
R1647 VDDA.n2830 VDDA.n2796 3.4105
R1648 VDDA.n2828 VDDA.n2827 3.4105
R1649 VDDA.n2798 VDDA.n2797 3.4105
R1650 VDDA.n2823 VDDA.n2822 3.4105
R1651 VDDA.n2820 VDDA.n2800 3.4105
R1652 VDDA.n2818 VDDA.n2817 3.4105
R1653 VDDA.n2802 VDDA.n2801 3.4105
R1654 VDDA.n2813 VDDA.n2812 3.4105
R1655 VDDA.n2810 VDDA.n2804 3.4105
R1656 VDDA.n2808 VDDA.n2807 3.4105
R1657 VDDA.n2922 VDDA.n2921 3.4105
R1658 VDDA.n196 VDDA.n195 3.4105
R1659 VDDA.n2747 VDDA.n2746 3.4105
R1660 VDDA.n2614 VDDA.n2613 3.4105
R1661 VDDA.n2742 VDDA.n2741 3.4105
R1662 VDDA.n2740 VDDA.n2739 3.4105
R1663 VDDA.n2738 VDDA.n2618 3.4105
R1664 VDDA.n2617 VDDA.n2616 3.4105
R1665 VDDA.n2734 VDDA.n2733 3.4105
R1666 VDDA.n2732 VDDA.n2731 3.4105
R1667 VDDA.n2730 VDDA.n2622 3.4105
R1668 VDDA.n2621 VDDA.n2620 3.4105
R1669 VDDA.n2726 VDDA.n2725 3.4105
R1670 VDDA.n2724 VDDA.n2723 3.4105
R1671 VDDA.n2722 VDDA.n2626 3.4105
R1672 VDDA.n2625 VDDA.n2624 3.4105
R1673 VDDA.n2718 VDDA.n2717 3.4105
R1674 VDDA.n2716 VDDA.n2715 3.4105
R1675 VDDA.n2714 VDDA.n2630 3.4105
R1676 VDDA.n2629 VDDA.n2628 3.4105
R1677 VDDA.n2710 VDDA.n2709 3.4105
R1678 VDDA.n2708 VDDA.n2707 3.4105
R1679 VDDA.n2706 VDDA.n2634 3.4105
R1680 VDDA.n2633 VDDA.n2632 3.4105
R1681 VDDA.n2702 VDDA.n2701 3.4105
R1682 VDDA.n2700 VDDA.n2699 3.4105
R1683 VDDA.n2698 VDDA.n2638 3.4105
R1684 VDDA.n2637 VDDA.n2636 3.4105
R1685 VDDA.n2694 VDDA.n2693 3.4105
R1686 VDDA.n2692 VDDA.n2691 3.4105
R1687 VDDA.n2690 VDDA.n2642 3.4105
R1688 VDDA.n2641 VDDA.n2640 3.4105
R1689 VDDA.n2686 VDDA.n2685 3.4105
R1690 VDDA.n2684 VDDA.n2683 3.4105
R1691 VDDA.n2682 VDDA.n2646 3.4105
R1692 VDDA.n2645 VDDA.n2644 3.4105
R1693 VDDA.n2678 VDDA.n2677 3.4105
R1694 VDDA.n2676 VDDA.n2675 3.4105
R1695 VDDA.n2674 VDDA.n2650 3.4105
R1696 VDDA.n2649 VDDA.n2648 3.4105
R1697 VDDA.n2670 VDDA.n2669 3.4105
R1698 VDDA.n2668 VDDA.n2667 3.4105
R1699 VDDA.n2666 VDDA.n2654 3.4105
R1700 VDDA.n2653 VDDA.n2652 3.4105
R1701 VDDA.n2662 VDDA.n2661 3.4105
R1702 VDDA.n2660 VDDA.n2659 3.4105
R1703 VDDA.n2658 VDDA.n2657 3.4105
R1704 VDDA.n2751 VDDA.n2750 3.4105
R1705 VDDA.n223 VDDA.n222 3.4105
R1706 VDDA.n357 VDDA.n356 3.4105
R1707 VDDA.n355 VDDA.n354 3.4105
R1708 VDDA.n353 VDDA.n227 3.4105
R1709 VDDA.n226 VDDA.n225 3.4105
R1710 VDDA.n349 VDDA.n348 3.4105
R1711 VDDA.n347 VDDA.n346 3.4105
R1712 VDDA.n345 VDDA.n231 3.4105
R1713 VDDA.n230 VDDA.n229 3.4105
R1714 VDDA.n341 VDDA.n340 3.4105
R1715 VDDA.n339 VDDA.n338 3.4105
R1716 VDDA.n337 VDDA.n235 3.4105
R1717 VDDA.n234 VDDA.n233 3.4105
R1718 VDDA.n333 VDDA.n332 3.4105
R1719 VDDA.n331 VDDA.n330 3.4105
R1720 VDDA.n329 VDDA.n239 3.4105
R1721 VDDA.n238 VDDA.n237 3.4105
R1722 VDDA.n325 VDDA.n324 3.4105
R1723 VDDA.n323 VDDA.n322 3.4105
R1724 VDDA.n321 VDDA.n243 3.4105
R1725 VDDA.n242 VDDA.n241 3.4105
R1726 VDDA.n317 VDDA.n316 3.4105
R1727 VDDA.n315 VDDA.n314 3.4105
R1728 VDDA.n313 VDDA.n247 3.4105
R1729 VDDA.n246 VDDA.n245 3.4105
R1730 VDDA.n309 VDDA.n308 3.4105
R1731 VDDA.n307 VDDA.n306 3.4105
R1732 VDDA.n305 VDDA.n251 3.4105
R1733 VDDA.n250 VDDA.n249 3.4105
R1734 VDDA.n301 VDDA.n300 3.4105
R1735 VDDA.n299 VDDA.n298 3.4105
R1736 VDDA.n297 VDDA.n255 3.4105
R1737 VDDA.n254 VDDA.n253 3.4105
R1738 VDDA.n293 VDDA.n292 3.4105
R1739 VDDA.n291 VDDA.n290 3.4105
R1740 VDDA.n289 VDDA.n259 3.4105
R1741 VDDA.n258 VDDA.n257 3.4105
R1742 VDDA.n285 VDDA.n284 3.4105
R1743 VDDA.n283 VDDA.n282 3.4105
R1744 VDDA.n281 VDDA.n263 3.4105
R1745 VDDA.n262 VDDA.n261 3.4105
R1746 VDDA.n277 VDDA.n276 3.4105
R1747 VDDA.n275 VDDA.n274 3.4105
R1748 VDDA.n273 VDDA.n267 3.4105
R1749 VDDA.n266 VDDA.n265 3.4105
R1750 VDDA.n269 VDDA.n268 3.4105
R1751 VDDA.n2588 VDDA.n2587 3.4105
R1752 VDDA.n526 VDDA.n366 3.4105
R1753 VDDA.n524 VDDA.n523 3.4105
R1754 VDDA.n368 VDDA.n367 3.4105
R1755 VDDA.n519 VDDA.n518 3.4105
R1756 VDDA.n516 VDDA.n370 3.4105
R1757 VDDA.n514 VDDA.n513 3.4105
R1758 VDDA.n372 VDDA.n371 3.4105
R1759 VDDA.n509 VDDA.n508 3.4105
R1760 VDDA.n506 VDDA.n374 3.4105
R1761 VDDA.n504 VDDA.n503 3.4105
R1762 VDDA.n376 VDDA.n375 3.4105
R1763 VDDA.n499 VDDA.n498 3.4105
R1764 VDDA.n496 VDDA.n378 3.4105
R1765 VDDA.n494 VDDA.n493 3.4105
R1766 VDDA.n380 VDDA.n379 3.4105
R1767 VDDA.n489 VDDA.n488 3.4105
R1768 VDDA.n486 VDDA.n382 3.4105
R1769 VDDA.n484 VDDA.n483 3.4105
R1770 VDDA.n384 VDDA.n383 3.4105
R1771 VDDA.n479 VDDA.n478 3.4105
R1772 VDDA.n476 VDDA.n386 3.4105
R1773 VDDA.n474 VDDA.n473 3.4105
R1774 VDDA.n388 VDDA.n387 3.4105
R1775 VDDA.n469 VDDA.n468 3.4105
R1776 VDDA.n466 VDDA.n390 3.4105
R1777 VDDA.n464 VDDA.n463 3.4105
R1778 VDDA.n392 VDDA.n391 3.4105
R1779 VDDA.n459 VDDA.n458 3.4105
R1780 VDDA.n456 VDDA.n394 3.4105
R1781 VDDA.n454 VDDA.n453 3.4105
R1782 VDDA.n396 VDDA.n395 3.4105
R1783 VDDA.n449 VDDA.n448 3.4105
R1784 VDDA.n446 VDDA.n398 3.4105
R1785 VDDA.n444 VDDA.n443 3.4105
R1786 VDDA.n400 VDDA.n399 3.4105
R1787 VDDA.n439 VDDA.n438 3.4105
R1788 VDDA.n436 VDDA.n402 3.4105
R1789 VDDA.n434 VDDA.n433 3.4105
R1790 VDDA.n404 VDDA.n403 3.4105
R1791 VDDA.n429 VDDA.n428 3.4105
R1792 VDDA.n426 VDDA.n406 3.4105
R1793 VDDA.n424 VDDA.n423 3.4105
R1794 VDDA.n408 VDDA.n407 3.4105
R1795 VDDA.n419 VDDA.n418 3.4105
R1796 VDDA.n416 VDDA.n410 3.4105
R1797 VDDA.n414 VDDA.n413 3.4105
R1798 VDDA.n528 VDDA.n527 3.4105
R1799 VDDA.n611 VDDA.n610 3.4105
R1800 VDDA.n1467 VDDA.n1466 3.4105
R1801 VDDA.n1334 VDDA.n1333 3.4105
R1802 VDDA.n1462 VDDA.n1461 3.4105
R1803 VDDA.n1460 VDDA.n1459 3.4105
R1804 VDDA.n1458 VDDA.n1338 3.4105
R1805 VDDA.n1337 VDDA.n1336 3.4105
R1806 VDDA.n1454 VDDA.n1453 3.4105
R1807 VDDA.n1452 VDDA.n1451 3.4105
R1808 VDDA.n1450 VDDA.n1342 3.4105
R1809 VDDA.n1341 VDDA.n1340 3.4105
R1810 VDDA.n1446 VDDA.n1445 3.4105
R1811 VDDA.n1444 VDDA.n1443 3.4105
R1812 VDDA.n1442 VDDA.n1346 3.4105
R1813 VDDA.n1345 VDDA.n1344 3.4105
R1814 VDDA.n1438 VDDA.n1437 3.4105
R1815 VDDA.n1436 VDDA.n1435 3.4105
R1816 VDDA.n1434 VDDA.n1350 3.4105
R1817 VDDA.n1349 VDDA.n1348 3.4105
R1818 VDDA.n1430 VDDA.n1429 3.4105
R1819 VDDA.n1428 VDDA.n1427 3.4105
R1820 VDDA.n1426 VDDA.n1354 3.4105
R1821 VDDA.n1353 VDDA.n1352 3.4105
R1822 VDDA.n1422 VDDA.n1421 3.4105
R1823 VDDA.n1420 VDDA.n1419 3.4105
R1824 VDDA.n1418 VDDA.n1358 3.4105
R1825 VDDA.n1357 VDDA.n1356 3.4105
R1826 VDDA.n1414 VDDA.n1413 3.4105
R1827 VDDA.n1412 VDDA.n1411 3.4105
R1828 VDDA.n1410 VDDA.n1362 3.4105
R1829 VDDA.n1361 VDDA.n1360 3.4105
R1830 VDDA.n1406 VDDA.n1405 3.4105
R1831 VDDA.n1404 VDDA.n1403 3.4105
R1832 VDDA.n1402 VDDA.n1366 3.4105
R1833 VDDA.n1365 VDDA.n1364 3.4105
R1834 VDDA.n1398 VDDA.n1397 3.4105
R1835 VDDA.n1396 VDDA.n1395 3.4105
R1836 VDDA.n1394 VDDA.n1370 3.4105
R1837 VDDA.n1369 VDDA.n1368 3.4105
R1838 VDDA.n1390 VDDA.n1389 3.4105
R1839 VDDA.n1388 VDDA.n1387 3.4105
R1840 VDDA.n1386 VDDA.n1374 3.4105
R1841 VDDA.n1373 VDDA.n1372 3.4105
R1842 VDDA.n1382 VDDA.n1381 3.4105
R1843 VDDA.n1380 VDDA.n1379 3.4105
R1844 VDDA.n1378 VDDA.n1377 3.4105
R1845 VDDA.n2408 VDDA.n2407 3.4105
R1846 VDDA.n638 VDDA.n637 3.4105
R1847 VDDA.n772 VDDA.n771 3.4105
R1848 VDDA.n770 VDDA.n769 3.4105
R1849 VDDA.n768 VDDA.n642 3.4105
R1850 VDDA.n641 VDDA.n640 3.4105
R1851 VDDA.n764 VDDA.n763 3.4105
R1852 VDDA.n762 VDDA.n761 3.4105
R1853 VDDA.n760 VDDA.n646 3.4105
R1854 VDDA.n645 VDDA.n644 3.4105
R1855 VDDA.n756 VDDA.n755 3.4105
R1856 VDDA.n754 VDDA.n753 3.4105
R1857 VDDA.n752 VDDA.n650 3.4105
R1858 VDDA.n649 VDDA.n648 3.4105
R1859 VDDA.n748 VDDA.n747 3.4105
R1860 VDDA.n746 VDDA.n745 3.4105
R1861 VDDA.n744 VDDA.n654 3.4105
R1862 VDDA.n653 VDDA.n652 3.4105
R1863 VDDA.n740 VDDA.n739 3.4105
R1864 VDDA.n738 VDDA.n737 3.4105
R1865 VDDA.n736 VDDA.n658 3.4105
R1866 VDDA.n657 VDDA.n656 3.4105
R1867 VDDA.n732 VDDA.n731 3.4105
R1868 VDDA.n730 VDDA.n729 3.4105
R1869 VDDA.n728 VDDA.n662 3.4105
R1870 VDDA.n661 VDDA.n660 3.4105
R1871 VDDA.n724 VDDA.n723 3.4105
R1872 VDDA.n722 VDDA.n721 3.4105
R1873 VDDA.n720 VDDA.n666 3.4105
R1874 VDDA.n665 VDDA.n664 3.4105
R1875 VDDA.n716 VDDA.n715 3.4105
R1876 VDDA.n714 VDDA.n713 3.4105
R1877 VDDA.n712 VDDA.n670 3.4105
R1878 VDDA.n669 VDDA.n668 3.4105
R1879 VDDA.n708 VDDA.n707 3.4105
R1880 VDDA.n706 VDDA.n705 3.4105
R1881 VDDA.n704 VDDA.n674 3.4105
R1882 VDDA.n673 VDDA.n672 3.4105
R1883 VDDA.n700 VDDA.n699 3.4105
R1884 VDDA.n698 VDDA.n697 3.4105
R1885 VDDA.n696 VDDA.n678 3.4105
R1886 VDDA.n677 VDDA.n676 3.4105
R1887 VDDA.n692 VDDA.n691 3.4105
R1888 VDDA.n690 VDDA.n689 3.4105
R1889 VDDA.n688 VDDA.n682 3.4105
R1890 VDDA.n681 VDDA.n680 3.4105
R1891 VDDA.n684 VDDA.n683 3.4105
R1892 VDDA.n1308 VDDA.n1307 3.4105
R1893 VDDA.n1292 VDDA.n1132 3.4105
R1894 VDDA.n1290 VDDA.n1289 3.4105
R1895 VDDA.n1134 VDDA.n1133 3.4105
R1896 VDDA.n1285 VDDA.n1284 3.4105
R1897 VDDA.n1282 VDDA.n1136 3.4105
R1898 VDDA.n1280 VDDA.n1279 3.4105
R1899 VDDA.n1138 VDDA.n1137 3.4105
R1900 VDDA.n1275 VDDA.n1274 3.4105
R1901 VDDA.n1272 VDDA.n1140 3.4105
R1902 VDDA.n1270 VDDA.n1269 3.4105
R1903 VDDA.n1142 VDDA.n1141 3.4105
R1904 VDDA.n1265 VDDA.n1264 3.4105
R1905 VDDA.n1262 VDDA.n1144 3.4105
R1906 VDDA.n1260 VDDA.n1259 3.4105
R1907 VDDA.n1146 VDDA.n1145 3.4105
R1908 VDDA.n1255 VDDA.n1254 3.4105
R1909 VDDA.n1252 VDDA.n1148 3.4105
R1910 VDDA.n1250 VDDA.n1249 3.4105
R1911 VDDA.n1150 VDDA.n1149 3.4105
R1912 VDDA.n1245 VDDA.n1244 3.4105
R1913 VDDA.n1242 VDDA.n1152 3.4105
R1914 VDDA.n1240 VDDA.n1239 3.4105
R1915 VDDA.n1154 VDDA.n1153 3.4105
R1916 VDDA.n1235 VDDA.n1234 3.4105
R1917 VDDA.n1232 VDDA.n1156 3.4105
R1918 VDDA.n1230 VDDA.n1229 3.4105
R1919 VDDA.n1158 VDDA.n1157 3.4105
R1920 VDDA.n1225 VDDA.n1224 3.4105
R1921 VDDA.n1222 VDDA.n1160 3.4105
R1922 VDDA.n1220 VDDA.n1219 3.4105
R1923 VDDA.n1162 VDDA.n1161 3.4105
R1924 VDDA.n1215 VDDA.n1214 3.4105
R1925 VDDA.n1212 VDDA.n1164 3.4105
R1926 VDDA.n1210 VDDA.n1209 3.4105
R1927 VDDA.n1166 VDDA.n1165 3.4105
R1928 VDDA.n1205 VDDA.n1204 3.4105
R1929 VDDA.n1202 VDDA.n1168 3.4105
R1930 VDDA.n1200 VDDA.n1199 3.4105
R1931 VDDA.n1170 VDDA.n1169 3.4105
R1932 VDDA.n1195 VDDA.n1194 3.4105
R1933 VDDA.n1192 VDDA.n1172 3.4105
R1934 VDDA.n1190 VDDA.n1189 3.4105
R1935 VDDA.n1174 VDDA.n1173 3.4105
R1936 VDDA.n1185 VDDA.n1184 3.4105
R1937 VDDA.n1182 VDDA.n1176 3.4105
R1938 VDDA.n1180 VDDA.n1179 3.4105
R1939 VDDA.n1294 VDDA.n1293 3.4105
R1940 VDDA.n788 VDDA.n787 3.4105
R1941 VDDA.n1119 VDDA.n1118 3.4105
R1942 VDDA.n986 VDDA.n985 3.4105
R1943 VDDA.n1114 VDDA.n1113 3.4105
R1944 VDDA.n1112 VDDA.n1111 3.4105
R1945 VDDA.n1110 VDDA.n990 3.4105
R1946 VDDA.n989 VDDA.n988 3.4105
R1947 VDDA.n1106 VDDA.n1105 3.4105
R1948 VDDA.n1104 VDDA.n1103 3.4105
R1949 VDDA.n1102 VDDA.n994 3.4105
R1950 VDDA.n993 VDDA.n992 3.4105
R1951 VDDA.n1098 VDDA.n1097 3.4105
R1952 VDDA.n1096 VDDA.n1095 3.4105
R1953 VDDA.n1094 VDDA.n998 3.4105
R1954 VDDA.n997 VDDA.n996 3.4105
R1955 VDDA.n1090 VDDA.n1089 3.4105
R1956 VDDA.n1088 VDDA.n1087 3.4105
R1957 VDDA.n1086 VDDA.n1002 3.4105
R1958 VDDA.n1001 VDDA.n1000 3.4105
R1959 VDDA.n1082 VDDA.n1081 3.4105
R1960 VDDA.n1080 VDDA.n1079 3.4105
R1961 VDDA.n1078 VDDA.n1006 3.4105
R1962 VDDA.n1005 VDDA.n1004 3.4105
R1963 VDDA.n1074 VDDA.n1073 3.4105
R1964 VDDA.n1072 VDDA.n1071 3.4105
R1965 VDDA.n1070 VDDA.n1010 3.4105
R1966 VDDA.n1009 VDDA.n1008 3.4105
R1967 VDDA.n1066 VDDA.n1065 3.4105
R1968 VDDA.n1064 VDDA.n1063 3.4105
R1969 VDDA.n1062 VDDA.n1014 3.4105
R1970 VDDA.n1013 VDDA.n1012 3.4105
R1971 VDDA.n1058 VDDA.n1057 3.4105
R1972 VDDA.n1056 VDDA.n1055 3.4105
R1973 VDDA.n1054 VDDA.n1018 3.4105
R1974 VDDA.n1017 VDDA.n1016 3.4105
R1975 VDDA.n1050 VDDA.n1049 3.4105
R1976 VDDA.n1048 VDDA.n1047 3.4105
R1977 VDDA.n1046 VDDA.n1022 3.4105
R1978 VDDA.n1021 VDDA.n1020 3.4105
R1979 VDDA.n1042 VDDA.n1041 3.4105
R1980 VDDA.n1040 VDDA.n1039 3.4105
R1981 VDDA.n1038 VDDA.n1026 3.4105
R1982 VDDA.n1025 VDDA.n1024 3.4105
R1983 VDDA.n1034 VDDA.n1033 3.4105
R1984 VDDA.n1032 VDDA.n1031 3.4105
R1985 VDDA.n1030 VDDA.n1029 3.4105
R1986 VDDA.n1123 VDDA.n1122 3.4105
R1987 VDDA.n814 VDDA.n813 3.4105
R1988 VDDA.n948 VDDA.n947 3.4105
R1989 VDDA.n946 VDDA.n945 3.4105
R1990 VDDA.n944 VDDA.n943 3.4105
R1991 VDDA.n942 VDDA.n816 3.4105
R1992 VDDA.n938 VDDA.n937 3.4105
R1993 VDDA.n936 VDDA.n935 3.4105
R1994 VDDA.n934 VDDA.n933 3.4105
R1995 VDDA.n932 VDDA.n818 3.4105
R1996 VDDA.n928 VDDA.n927 3.4105
R1997 VDDA.n926 VDDA.n925 3.4105
R1998 VDDA.n924 VDDA.n923 3.4105
R1999 VDDA.n922 VDDA.n820 3.4105
R2000 VDDA.n918 VDDA.n917 3.4105
R2001 VDDA.n916 VDDA.n915 3.4105
R2002 VDDA.n914 VDDA.n913 3.4105
R2003 VDDA.n912 VDDA.n822 3.4105
R2004 VDDA.n908 VDDA.n907 3.4105
R2005 VDDA.n906 VDDA.n905 3.4105
R2006 VDDA.n904 VDDA.n903 3.4105
R2007 VDDA.n902 VDDA.n824 3.4105
R2008 VDDA.n898 VDDA.n897 3.4105
R2009 VDDA.n896 VDDA.n895 3.4105
R2010 VDDA.n894 VDDA.n893 3.4105
R2011 VDDA.n892 VDDA.n826 3.4105
R2012 VDDA.n888 VDDA.n887 3.4105
R2013 VDDA.n886 VDDA.n885 3.4105
R2014 VDDA.n884 VDDA.n883 3.4105
R2015 VDDA.n882 VDDA.n828 3.4105
R2016 VDDA.n878 VDDA.n877 3.4105
R2017 VDDA.n876 VDDA.n875 3.4105
R2018 VDDA.n874 VDDA.n873 3.4105
R2019 VDDA.n872 VDDA.n830 3.4105
R2020 VDDA.n868 VDDA.n867 3.4105
R2021 VDDA.n866 VDDA.n865 3.4105
R2022 VDDA.n864 VDDA.n863 3.4105
R2023 VDDA.n862 VDDA.n832 3.4105
R2024 VDDA.n858 VDDA.n857 3.4105
R2025 VDDA.n856 VDDA.n855 3.4105
R2026 VDDA.n854 VDDA.n853 3.4105
R2027 VDDA.n852 VDDA.n834 3.4105
R2028 VDDA.n848 VDDA.n847 3.4105
R2029 VDDA.n846 VDDA.n845 3.4105
R2030 VDDA.n844 VDDA.n843 3.4105
R2031 VDDA.n842 VDDA.n836 3.4105
R2032 VDDA.n838 VDDA.n837 3.4105
R2033 VDDA.n960 VDDA.n959 3.4105
R2034 VDDA.n961 VDDA.n789 3.4105
R2035 VDDA.n961 VDDA.n960 3.4105
R2036 VDDA.n1121 VDDA.n962 3.4105
R2037 VDDA.n1122 VDDA.n1121 3.4105
R2038 VDDA.n1177 VDDA.n612 3.4105
R2039 VDDA.n1293 VDDA.n612 3.4105
R2040 VDDA.n1309 VDDA.n613 3.4105
R2041 VDDA.n1309 VDDA.n1308 3.4105
R2042 VDDA.n2406 VDDA.n1310 3.4105
R2043 VDDA.n2407 VDDA.n2406 3.4105
R2044 VDDA.n2405 VDDA.n2404 3.4105
R2045 VDDA.n411 VDDA.n197 3.4105
R2046 VDDA.n527 VDDA.n197 3.4105
R2047 VDDA.n2589 VDDA.n198 3.4105
R2048 VDDA.n2589 VDDA.n2588 3.4105
R2049 VDDA.n2749 VDDA.n2590 3.4105
R2050 VDDA.n2750 VDDA.n2749 3.4105
R2051 VDDA.n2805 VDDA.n19 3.4105
R2052 VDDA.n2921 VDDA.n19 3.4105
R2053 VDDA.n2937 VDDA.n20 3.4105
R2054 VDDA.n2937 VDDA.n2936 3.4105
R2055 VDDA.n1728 VDDA.n1558 3.4105
R2056 VDDA.n1728 VDDA.n1727 3.4105
R2057 VDDA.n2056 VDDA.n1492 3.4105
R2058 VDDA.n2056 VDDA.n2055 3.4105
R2059 VDDA.n1729 VDDA.n1557 3.4105
R2060 VDDA.n1794 VDDA.n1729 3.4105
R2061 VDDA.n3124 VDDA.n17 3.4105
R2062 VDDA.n3124 VDDA.n16 3.4105
R2063 VDDA.n3124 VDDA.n18 3.4105
R2064 VDDA.n3124 VDDA.n3123 3.4105
R2065 VDDA.n3123 VDDA.n2974 3.4105
R2066 VDDA.n2971 VDDA.n16 3.4105
R2067 VDDA.n3093 VDDA.n2971 3.4105
R2068 VDDA.n3090 VDDA.n2971 3.4105
R2069 VDDA.n3095 VDDA.n2971 3.4105
R2070 VDDA.n3089 VDDA.n2971 3.4105
R2071 VDDA.n3097 VDDA.n2971 3.4105
R2072 VDDA.n3088 VDDA.n2971 3.4105
R2073 VDDA.n3099 VDDA.n2971 3.4105
R2074 VDDA.n3087 VDDA.n2971 3.4105
R2075 VDDA.n3101 VDDA.n2971 3.4105
R2076 VDDA.n3086 VDDA.n2971 3.4105
R2077 VDDA.n3103 VDDA.n2971 3.4105
R2078 VDDA.n3085 VDDA.n2971 3.4105
R2079 VDDA.n3105 VDDA.n2971 3.4105
R2080 VDDA.n3084 VDDA.n2971 3.4105
R2081 VDDA.n3107 VDDA.n2971 3.4105
R2082 VDDA.n3083 VDDA.n2971 3.4105
R2083 VDDA.n3109 VDDA.n2971 3.4105
R2084 VDDA.n3082 VDDA.n2971 3.4105
R2085 VDDA.n3111 VDDA.n2971 3.4105
R2086 VDDA.n3081 VDDA.n2971 3.4105
R2087 VDDA.n3113 VDDA.n2971 3.4105
R2088 VDDA.n3080 VDDA.n2971 3.4105
R2089 VDDA.n3115 VDDA.n2971 3.4105
R2090 VDDA.n3079 VDDA.n2971 3.4105
R2091 VDDA.n3117 VDDA.n2971 3.4105
R2092 VDDA.n3078 VDDA.n2971 3.4105
R2093 VDDA.n3119 VDDA.n2971 3.4105
R2094 VDDA.n3077 VDDA.n2971 3.4105
R2095 VDDA.n3121 VDDA.n2971 3.4105
R2096 VDDA.n3076 VDDA.n2971 3.4105
R2097 VDDA.n2971 VDDA.n18 3.4105
R2098 VDDA.n3123 VDDA.n2971 3.4105
R2099 VDDA.n2977 VDDA.n16 3.4105
R2100 VDDA.n3093 VDDA.n2977 3.4105
R2101 VDDA.n3090 VDDA.n2977 3.4105
R2102 VDDA.n3095 VDDA.n2977 3.4105
R2103 VDDA.n3089 VDDA.n2977 3.4105
R2104 VDDA.n3097 VDDA.n2977 3.4105
R2105 VDDA.n3088 VDDA.n2977 3.4105
R2106 VDDA.n3099 VDDA.n2977 3.4105
R2107 VDDA.n3087 VDDA.n2977 3.4105
R2108 VDDA.n3101 VDDA.n2977 3.4105
R2109 VDDA.n3086 VDDA.n2977 3.4105
R2110 VDDA.n3103 VDDA.n2977 3.4105
R2111 VDDA.n3085 VDDA.n2977 3.4105
R2112 VDDA.n3105 VDDA.n2977 3.4105
R2113 VDDA.n3084 VDDA.n2977 3.4105
R2114 VDDA.n3107 VDDA.n2977 3.4105
R2115 VDDA.n3083 VDDA.n2977 3.4105
R2116 VDDA.n3109 VDDA.n2977 3.4105
R2117 VDDA.n3082 VDDA.n2977 3.4105
R2118 VDDA.n3111 VDDA.n2977 3.4105
R2119 VDDA.n3081 VDDA.n2977 3.4105
R2120 VDDA.n3113 VDDA.n2977 3.4105
R2121 VDDA.n3080 VDDA.n2977 3.4105
R2122 VDDA.n3115 VDDA.n2977 3.4105
R2123 VDDA.n3079 VDDA.n2977 3.4105
R2124 VDDA.n3117 VDDA.n2977 3.4105
R2125 VDDA.n3078 VDDA.n2977 3.4105
R2126 VDDA.n3119 VDDA.n2977 3.4105
R2127 VDDA.n3077 VDDA.n2977 3.4105
R2128 VDDA.n3121 VDDA.n2977 3.4105
R2129 VDDA.n3076 VDDA.n2977 3.4105
R2130 VDDA.n2977 VDDA.n18 3.4105
R2131 VDDA.n3123 VDDA.n2977 3.4105
R2132 VDDA.n2970 VDDA.n16 3.4105
R2133 VDDA.n3093 VDDA.n2970 3.4105
R2134 VDDA.n3090 VDDA.n2970 3.4105
R2135 VDDA.n3095 VDDA.n2970 3.4105
R2136 VDDA.n3089 VDDA.n2970 3.4105
R2137 VDDA.n3097 VDDA.n2970 3.4105
R2138 VDDA.n3088 VDDA.n2970 3.4105
R2139 VDDA.n3099 VDDA.n2970 3.4105
R2140 VDDA.n3087 VDDA.n2970 3.4105
R2141 VDDA.n3101 VDDA.n2970 3.4105
R2142 VDDA.n3086 VDDA.n2970 3.4105
R2143 VDDA.n3103 VDDA.n2970 3.4105
R2144 VDDA.n3085 VDDA.n2970 3.4105
R2145 VDDA.n3105 VDDA.n2970 3.4105
R2146 VDDA.n3084 VDDA.n2970 3.4105
R2147 VDDA.n3107 VDDA.n2970 3.4105
R2148 VDDA.n3083 VDDA.n2970 3.4105
R2149 VDDA.n3109 VDDA.n2970 3.4105
R2150 VDDA.n3082 VDDA.n2970 3.4105
R2151 VDDA.n3111 VDDA.n2970 3.4105
R2152 VDDA.n3081 VDDA.n2970 3.4105
R2153 VDDA.n3113 VDDA.n2970 3.4105
R2154 VDDA.n3080 VDDA.n2970 3.4105
R2155 VDDA.n3115 VDDA.n2970 3.4105
R2156 VDDA.n3079 VDDA.n2970 3.4105
R2157 VDDA.n3117 VDDA.n2970 3.4105
R2158 VDDA.n3078 VDDA.n2970 3.4105
R2159 VDDA.n3119 VDDA.n2970 3.4105
R2160 VDDA.n3077 VDDA.n2970 3.4105
R2161 VDDA.n3121 VDDA.n2970 3.4105
R2162 VDDA.n3076 VDDA.n2970 3.4105
R2163 VDDA.n2970 VDDA.n18 3.4105
R2164 VDDA.n3123 VDDA.n2970 3.4105
R2165 VDDA.n2980 VDDA.n16 3.4105
R2166 VDDA.n3093 VDDA.n2980 3.4105
R2167 VDDA.n3090 VDDA.n2980 3.4105
R2168 VDDA.n3095 VDDA.n2980 3.4105
R2169 VDDA.n3089 VDDA.n2980 3.4105
R2170 VDDA.n3097 VDDA.n2980 3.4105
R2171 VDDA.n3088 VDDA.n2980 3.4105
R2172 VDDA.n3099 VDDA.n2980 3.4105
R2173 VDDA.n3087 VDDA.n2980 3.4105
R2174 VDDA.n3101 VDDA.n2980 3.4105
R2175 VDDA.n3086 VDDA.n2980 3.4105
R2176 VDDA.n3103 VDDA.n2980 3.4105
R2177 VDDA.n3085 VDDA.n2980 3.4105
R2178 VDDA.n3105 VDDA.n2980 3.4105
R2179 VDDA.n3084 VDDA.n2980 3.4105
R2180 VDDA.n3107 VDDA.n2980 3.4105
R2181 VDDA.n3083 VDDA.n2980 3.4105
R2182 VDDA.n3109 VDDA.n2980 3.4105
R2183 VDDA.n3082 VDDA.n2980 3.4105
R2184 VDDA.n3111 VDDA.n2980 3.4105
R2185 VDDA.n3081 VDDA.n2980 3.4105
R2186 VDDA.n3113 VDDA.n2980 3.4105
R2187 VDDA.n3080 VDDA.n2980 3.4105
R2188 VDDA.n3115 VDDA.n2980 3.4105
R2189 VDDA.n3079 VDDA.n2980 3.4105
R2190 VDDA.n3117 VDDA.n2980 3.4105
R2191 VDDA.n3078 VDDA.n2980 3.4105
R2192 VDDA.n3119 VDDA.n2980 3.4105
R2193 VDDA.n3077 VDDA.n2980 3.4105
R2194 VDDA.n3121 VDDA.n2980 3.4105
R2195 VDDA.n3076 VDDA.n2980 3.4105
R2196 VDDA.n2980 VDDA.n18 3.4105
R2197 VDDA.n3123 VDDA.n2980 3.4105
R2198 VDDA.n2969 VDDA.n16 3.4105
R2199 VDDA.n3093 VDDA.n2969 3.4105
R2200 VDDA.n3090 VDDA.n2969 3.4105
R2201 VDDA.n3095 VDDA.n2969 3.4105
R2202 VDDA.n3089 VDDA.n2969 3.4105
R2203 VDDA.n3097 VDDA.n2969 3.4105
R2204 VDDA.n3088 VDDA.n2969 3.4105
R2205 VDDA.n3099 VDDA.n2969 3.4105
R2206 VDDA.n3087 VDDA.n2969 3.4105
R2207 VDDA.n3101 VDDA.n2969 3.4105
R2208 VDDA.n3086 VDDA.n2969 3.4105
R2209 VDDA.n3103 VDDA.n2969 3.4105
R2210 VDDA.n3085 VDDA.n2969 3.4105
R2211 VDDA.n3105 VDDA.n2969 3.4105
R2212 VDDA.n3084 VDDA.n2969 3.4105
R2213 VDDA.n3107 VDDA.n2969 3.4105
R2214 VDDA.n3083 VDDA.n2969 3.4105
R2215 VDDA.n3109 VDDA.n2969 3.4105
R2216 VDDA.n3082 VDDA.n2969 3.4105
R2217 VDDA.n3111 VDDA.n2969 3.4105
R2218 VDDA.n3081 VDDA.n2969 3.4105
R2219 VDDA.n3113 VDDA.n2969 3.4105
R2220 VDDA.n3080 VDDA.n2969 3.4105
R2221 VDDA.n3115 VDDA.n2969 3.4105
R2222 VDDA.n3079 VDDA.n2969 3.4105
R2223 VDDA.n3117 VDDA.n2969 3.4105
R2224 VDDA.n3078 VDDA.n2969 3.4105
R2225 VDDA.n3119 VDDA.n2969 3.4105
R2226 VDDA.n3077 VDDA.n2969 3.4105
R2227 VDDA.n3121 VDDA.n2969 3.4105
R2228 VDDA.n3076 VDDA.n2969 3.4105
R2229 VDDA.n2969 VDDA.n18 3.4105
R2230 VDDA.n3123 VDDA.n2969 3.4105
R2231 VDDA.n2983 VDDA.n16 3.4105
R2232 VDDA.n3093 VDDA.n2983 3.4105
R2233 VDDA.n3090 VDDA.n2983 3.4105
R2234 VDDA.n3095 VDDA.n2983 3.4105
R2235 VDDA.n3089 VDDA.n2983 3.4105
R2236 VDDA.n3097 VDDA.n2983 3.4105
R2237 VDDA.n3088 VDDA.n2983 3.4105
R2238 VDDA.n3099 VDDA.n2983 3.4105
R2239 VDDA.n3087 VDDA.n2983 3.4105
R2240 VDDA.n3101 VDDA.n2983 3.4105
R2241 VDDA.n3086 VDDA.n2983 3.4105
R2242 VDDA.n3103 VDDA.n2983 3.4105
R2243 VDDA.n3085 VDDA.n2983 3.4105
R2244 VDDA.n3105 VDDA.n2983 3.4105
R2245 VDDA.n3084 VDDA.n2983 3.4105
R2246 VDDA.n3107 VDDA.n2983 3.4105
R2247 VDDA.n3083 VDDA.n2983 3.4105
R2248 VDDA.n3109 VDDA.n2983 3.4105
R2249 VDDA.n3082 VDDA.n2983 3.4105
R2250 VDDA.n3111 VDDA.n2983 3.4105
R2251 VDDA.n3081 VDDA.n2983 3.4105
R2252 VDDA.n3113 VDDA.n2983 3.4105
R2253 VDDA.n3080 VDDA.n2983 3.4105
R2254 VDDA.n3115 VDDA.n2983 3.4105
R2255 VDDA.n3079 VDDA.n2983 3.4105
R2256 VDDA.n3117 VDDA.n2983 3.4105
R2257 VDDA.n3078 VDDA.n2983 3.4105
R2258 VDDA.n3119 VDDA.n2983 3.4105
R2259 VDDA.n3077 VDDA.n2983 3.4105
R2260 VDDA.n3121 VDDA.n2983 3.4105
R2261 VDDA.n3076 VDDA.n2983 3.4105
R2262 VDDA.n2983 VDDA.n18 3.4105
R2263 VDDA.n3123 VDDA.n2983 3.4105
R2264 VDDA.n2968 VDDA.n16 3.4105
R2265 VDDA.n3093 VDDA.n2968 3.4105
R2266 VDDA.n3090 VDDA.n2968 3.4105
R2267 VDDA.n3095 VDDA.n2968 3.4105
R2268 VDDA.n3089 VDDA.n2968 3.4105
R2269 VDDA.n3097 VDDA.n2968 3.4105
R2270 VDDA.n3088 VDDA.n2968 3.4105
R2271 VDDA.n3099 VDDA.n2968 3.4105
R2272 VDDA.n3087 VDDA.n2968 3.4105
R2273 VDDA.n3101 VDDA.n2968 3.4105
R2274 VDDA.n3086 VDDA.n2968 3.4105
R2275 VDDA.n3103 VDDA.n2968 3.4105
R2276 VDDA.n3085 VDDA.n2968 3.4105
R2277 VDDA.n3105 VDDA.n2968 3.4105
R2278 VDDA.n3084 VDDA.n2968 3.4105
R2279 VDDA.n3107 VDDA.n2968 3.4105
R2280 VDDA.n3083 VDDA.n2968 3.4105
R2281 VDDA.n3109 VDDA.n2968 3.4105
R2282 VDDA.n3082 VDDA.n2968 3.4105
R2283 VDDA.n3111 VDDA.n2968 3.4105
R2284 VDDA.n3081 VDDA.n2968 3.4105
R2285 VDDA.n3113 VDDA.n2968 3.4105
R2286 VDDA.n3080 VDDA.n2968 3.4105
R2287 VDDA.n3115 VDDA.n2968 3.4105
R2288 VDDA.n3079 VDDA.n2968 3.4105
R2289 VDDA.n3117 VDDA.n2968 3.4105
R2290 VDDA.n3078 VDDA.n2968 3.4105
R2291 VDDA.n3119 VDDA.n2968 3.4105
R2292 VDDA.n3077 VDDA.n2968 3.4105
R2293 VDDA.n3121 VDDA.n2968 3.4105
R2294 VDDA.n3076 VDDA.n2968 3.4105
R2295 VDDA.n2968 VDDA.n18 3.4105
R2296 VDDA.n3123 VDDA.n2968 3.4105
R2297 VDDA.n2986 VDDA.n16 3.4105
R2298 VDDA.n3093 VDDA.n2986 3.4105
R2299 VDDA.n3090 VDDA.n2986 3.4105
R2300 VDDA.n3095 VDDA.n2986 3.4105
R2301 VDDA.n3089 VDDA.n2986 3.4105
R2302 VDDA.n3097 VDDA.n2986 3.4105
R2303 VDDA.n3088 VDDA.n2986 3.4105
R2304 VDDA.n3099 VDDA.n2986 3.4105
R2305 VDDA.n3087 VDDA.n2986 3.4105
R2306 VDDA.n3101 VDDA.n2986 3.4105
R2307 VDDA.n3086 VDDA.n2986 3.4105
R2308 VDDA.n3103 VDDA.n2986 3.4105
R2309 VDDA.n3085 VDDA.n2986 3.4105
R2310 VDDA.n3105 VDDA.n2986 3.4105
R2311 VDDA.n3084 VDDA.n2986 3.4105
R2312 VDDA.n3107 VDDA.n2986 3.4105
R2313 VDDA.n3083 VDDA.n2986 3.4105
R2314 VDDA.n3109 VDDA.n2986 3.4105
R2315 VDDA.n3082 VDDA.n2986 3.4105
R2316 VDDA.n3111 VDDA.n2986 3.4105
R2317 VDDA.n3081 VDDA.n2986 3.4105
R2318 VDDA.n3113 VDDA.n2986 3.4105
R2319 VDDA.n3080 VDDA.n2986 3.4105
R2320 VDDA.n3115 VDDA.n2986 3.4105
R2321 VDDA.n3079 VDDA.n2986 3.4105
R2322 VDDA.n3117 VDDA.n2986 3.4105
R2323 VDDA.n3078 VDDA.n2986 3.4105
R2324 VDDA.n3119 VDDA.n2986 3.4105
R2325 VDDA.n3077 VDDA.n2986 3.4105
R2326 VDDA.n3121 VDDA.n2986 3.4105
R2327 VDDA.n3076 VDDA.n2986 3.4105
R2328 VDDA.n2986 VDDA.n18 3.4105
R2329 VDDA.n3123 VDDA.n2986 3.4105
R2330 VDDA.n2967 VDDA.n16 3.4105
R2331 VDDA.n3093 VDDA.n2967 3.4105
R2332 VDDA.n3090 VDDA.n2967 3.4105
R2333 VDDA.n3095 VDDA.n2967 3.4105
R2334 VDDA.n3089 VDDA.n2967 3.4105
R2335 VDDA.n3097 VDDA.n2967 3.4105
R2336 VDDA.n3088 VDDA.n2967 3.4105
R2337 VDDA.n3099 VDDA.n2967 3.4105
R2338 VDDA.n3087 VDDA.n2967 3.4105
R2339 VDDA.n3101 VDDA.n2967 3.4105
R2340 VDDA.n3086 VDDA.n2967 3.4105
R2341 VDDA.n3103 VDDA.n2967 3.4105
R2342 VDDA.n3085 VDDA.n2967 3.4105
R2343 VDDA.n3105 VDDA.n2967 3.4105
R2344 VDDA.n3084 VDDA.n2967 3.4105
R2345 VDDA.n3107 VDDA.n2967 3.4105
R2346 VDDA.n3083 VDDA.n2967 3.4105
R2347 VDDA.n3109 VDDA.n2967 3.4105
R2348 VDDA.n3082 VDDA.n2967 3.4105
R2349 VDDA.n3111 VDDA.n2967 3.4105
R2350 VDDA.n3081 VDDA.n2967 3.4105
R2351 VDDA.n3113 VDDA.n2967 3.4105
R2352 VDDA.n3080 VDDA.n2967 3.4105
R2353 VDDA.n3115 VDDA.n2967 3.4105
R2354 VDDA.n3079 VDDA.n2967 3.4105
R2355 VDDA.n3117 VDDA.n2967 3.4105
R2356 VDDA.n3078 VDDA.n2967 3.4105
R2357 VDDA.n3119 VDDA.n2967 3.4105
R2358 VDDA.n3077 VDDA.n2967 3.4105
R2359 VDDA.n3121 VDDA.n2967 3.4105
R2360 VDDA.n3076 VDDA.n2967 3.4105
R2361 VDDA.n2967 VDDA.n18 3.4105
R2362 VDDA.n3123 VDDA.n2967 3.4105
R2363 VDDA.n2989 VDDA.n16 3.4105
R2364 VDDA.n3093 VDDA.n2989 3.4105
R2365 VDDA.n3090 VDDA.n2989 3.4105
R2366 VDDA.n3095 VDDA.n2989 3.4105
R2367 VDDA.n3089 VDDA.n2989 3.4105
R2368 VDDA.n3097 VDDA.n2989 3.4105
R2369 VDDA.n3088 VDDA.n2989 3.4105
R2370 VDDA.n3099 VDDA.n2989 3.4105
R2371 VDDA.n3087 VDDA.n2989 3.4105
R2372 VDDA.n3101 VDDA.n2989 3.4105
R2373 VDDA.n3086 VDDA.n2989 3.4105
R2374 VDDA.n3103 VDDA.n2989 3.4105
R2375 VDDA.n3085 VDDA.n2989 3.4105
R2376 VDDA.n3105 VDDA.n2989 3.4105
R2377 VDDA.n3084 VDDA.n2989 3.4105
R2378 VDDA.n3107 VDDA.n2989 3.4105
R2379 VDDA.n3083 VDDA.n2989 3.4105
R2380 VDDA.n3109 VDDA.n2989 3.4105
R2381 VDDA.n3082 VDDA.n2989 3.4105
R2382 VDDA.n3111 VDDA.n2989 3.4105
R2383 VDDA.n3081 VDDA.n2989 3.4105
R2384 VDDA.n3113 VDDA.n2989 3.4105
R2385 VDDA.n3080 VDDA.n2989 3.4105
R2386 VDDA.n3115 VDDA.n2989 3.4105
R2387 VDDA.n3079 VDDA.n2989 3.4105
R2388 VDDA.n3117 VDDA.n2989 3.4105
R2389 VDDA.n3078 VDDA.n2989 3.4105
R2390 VDDA.n3119 VDDA.n2989 3.4105
R2391 VDDA.n3077 VDDA.n2989 3.4105
R2392 VDDA.n3121 VDDA.n2989 3.4105
R2393 VDDA.n3076 VDDA.n2989 3.4105
R2394 VDDA.n2989 VDDA.n18 3.4105
R2395 VDDA.n3123 VDDA.n2989 3.4105
R2396 VDDA.n2966 VDDA.n16 3.4105
R2397 VDDA.n3093 VDDA.n2966 3.4105
R2398 VDDA.n3090 VDDA.n2966 3.4105
R2399 VDDA.n3095 VDDA.n2966 3.4105
R2400 VDDA.n3089 VDDA.n2966 3.4105
R2401 VDDA.n3097 VDDA.n2966 3.4105
R2402 VDDA.n3088 VDDA.n2966 3.4105
R2403 VDDA.n3099 VDDA.n2966 3.4105
R2404 VDDA.n3087 VDDA.n2966 3.4105
R2405 VDDA.n3101 VDDA.n2966 3.4105
R2406 VDDA.n3086 VDDA.n2966 3.4105
R2407 VDDA.n3103 VDDA.n2966 3.4105
R2408 VDDA.n3085 VDDA.n2966 3.4105
R2409 VDDA.n3105 VDDA.n2966 3.4105
R2410 VDDA.n3084 VDDA.n2966 3.4105
R2411 VDDA.n3107 VDDA.n2966 3.4105
R2412 VDDA.n3083 VDDA.n2966 3.4105
R2413 VDDA.n3109 VDDA.n2966 3.4105
R2414 VDDA.n3082 VDDA.n2966 3.4105
R2415 VDDA.n3111 VDDA.n2966 3.4105
R2416 VDDA.n3081 VDDA.n2966 3.4105
R2417 VDDA.n3113 VDDA.n2966 3.4105
R2418 VDDA.n3080 VDDA.n2966 3.4105
R2419 VDDA.n3115 VDDA.n2966 3.4105
R2420 VDDA.n3079 VDDA.n2966 3.4105
R2421 VDDA.n3117 VDDA.n2966 3.4105
R2422 VDDA.n3078 VDDA.n2966 3.4105
R2423 VDDA.n3119 VDDA.n2966 3.4105
R2424 VDDA.n3077 VDDA.n2966 3.4105
R2425 VDDA.n3121 VDDA.n2966 3.4105
R2426 VDDA.n3076 VDDA.n2966 3.4105
R2427 VDDA.n2966 VDDA.n18 3.4105
R2428 VDDA.n3123 VDDA.n2966 3.4105
R2429 VDDA.n2992 VDDA.n16 3.4105
R2430 VDDA.n3093 VDDA.n2992 3.4105
R2431 VDDA.n3090 VDDA.n2992 3.4105
R2432 VDDA.n3095 VDDA.n2992 3.4105
R2433 VDDA.n3089 VDDA.n2992 3.4105
R2434 VDDA.n3097 VDDA.n2992 3.4105
R2435 VDDA.n3088 VDDA.n2992 3.4105
R2436 VDDA.n3099 VDDA.n2992 3.4105
R2437 VDDA.n3087 VDDA.n2992 3.4105
R2438 VDDA.n3101 VDDA.n2992 3.4105
R2439 VDDA.n3086 VDDA.n2992 3.4105
R2440 VDDA.n3103 VDDA.n2992 3.4105
R2441 VDDA.n3085 VDDA.n2992 3.4105
R2442 VDDA.n3105 VDDA.n2992 3.4105
R2443 VDDA.n3084 VDDA.n2992 3.4105
R2444 VDDA.n3107 VDDA.n2992 3.4105
R2445 VDDA.n3083 VDDA.n2992 3.4105
R2446 VDDA.n3109 VDDA.n2992 3.4105
R2447 VDDA.n3082 VDDA.n2992 3.4105
R2448 VDDA.n3111 VDDA.n2992 3.4105
R2449 VDDA.n3081 VDDA.n2992 3.4105
R2450 VDDA.n3113 VDDA.n2992 3.4105
R2451 VDDA.n3080 VDDA.n2992 3.4105
R2452 VDDA.n3115 VDDA.n2992 3.4105
R2453 VDDA.n3079 VDDA.n2992 3.4105
R2454 VDDA.n3117 VDDA.n2992 3.4105
R2455 VDDA.n3078 VDDA.n2992 3.4105
R2456 VDDA.n3119 VDDA.n2992 3.4105
R2457 VDDA.n3077 VDDA.n2992 3.4105
R2458 VDDA.n3121 VDDA.n2992 3.4105
R2459 VDDA.n3076 VDDA.n2992 3.4105
R2460 VDDA.n2992 VDDA.n18 3.4105
R2461 VDDA.n3123 VDDA.n2992 3.4105
R2462 VDDA.n2965 VDDA.n16 3.4105
R2463 VDDA.n3093 VDDA.n2965 3.4105
R2464 VDDA.n3090 VDDA.n2965 3.4105
R2465 VDDA.n3095 VDDA.n2965 3.4105
R2466 VDDA.n3089 VDDA.n2965 3.4105
R2467 VDDA.n3097 VDDA.n2965 3.4105
R2468 VDDA.n3088 VDDA.n2965 3.4105
R2469 VDDA.n3099 VDDA.n2965 3.4105
R2470 VDDA.n3087 VDDA.n2965 3.4105
R2471 VDDA.n3101 VDDA.n2965 3.4105
R2472 VDDA.n3086 VDDA.n2965 3.4105
R2473 VDDA.n3103 VDDA.n2965 3.4105
R2474 VDDA.n3085 VDDA.n2965 3.4105
R2475 VDDA.n3105 VDDA.n2965 3.4105
R2476 VDDA.n3084 VDDA.n2965 3.4105
R2477 VDDA.n3107 VDDA.n2965 3.4105
R2478 VDDA.n3083 VDDA.n2965 3.4105
R2479 VDDA.n3109 VDDA.n2965 3.4105
R2480 VDDA.n3082 VDDA.n2965 3.4105
R2481 VDDA.n3111 VDDA.n2965 3.4105
R2482 VDDA.n3081 VDDA.n2965 3.4105
R2483 VDDA.n3113 VDDA.n2965 3.4105
R2484 VDDA.n3080 VDDA.n2965 3.4105
R2485 VDDA.n3115 VDDA.n2965 3.4105
R2486 VDDA.n3079 VDDA.n2965 3.4105
R2487 VDDA.n3117 VDDA.n2965 3.4105
R2488 VDDA.n3078 VDDA.n2965 3.4105
R2489 VDDA.n3119 VDDA.n2965 3.4105
R2490 VDDA.n3077 VDDA.n2965 3.4105
R2491 VDDA.n3121 VDDA.n2965 3.4105
R2492 VDDA.n3076 VDDA.n2965 3.4105
R2493 VDDA.n2965 VDDA.n18 3.4105
R2494 VDDA.n3123 VDDA.n2965 3.4105
R2495 VDDA.n2995 VDDA.n16 3.4105
R2496 VDDA.n3093 VDDA.n2995 3.4105
R2497 VDDA.n3090 VDDA.n2995 3.4105
R2498 VDDA.n3095 VDDA.n2995 3.4105
R2499 VDDA.n3089 VDDA.n2995 3.4105
R2500 VDDA.n3097 VDDA.n2995 3.4105
R2501 VDDA.n3088 VDDA.n2995 3.4105
R2502 VDDA.n3099 VDDA.n2995 3.4105
R2503 VDDA.n3087 VDDA.n2995 3.4105
R2504 VDDA.n3101 VDDA.n2995 3.4105
R2505 VDDA.n3086 VDDA.n2995 3.4105
R2506 VDDA.n3103 VDDA.n2995 3.4105
R2507 VDDA.n3085 VDDA.n2995 3.4105
R2508 VDDA.n3105 VDDA.n2995 3.4105
R2509 VDDA.n3084 VDDA.n2995 3.4105
R2510 VDDA.n3107 VDDA.n2995 3.4105
R2511 VDDA.n3083 VDDA.n2995 3.4105
R2512 VDDA.n3109 VDDA.n2995 3.4105
R2513 VDDA.n3082 VDDA.n2995 3.4105
R2514 VDDA.n3111 VDDA.n2995 3.4105
R2515 VDDA.n3081 VDDA.n2995 3.4105
R2516 VDDA.n3113 VDDA.n2995 3.4105
R2517 VDDA.n3080 VDDA.n2995 3.4105
R2518 VDDA.n3115 VDDA.n2995 3.4105
R2519 VDDA.n3079 VDDA.n2995 3.4105
R2520 VDDA.n3117 VDDA.n2995 3.4105
R2521 VDDA.n3078 VDDA.n2995 3.4105
R2522 VDDA.n3119 VDDA.n2995 3.4105
R2523 VDDA.n3077 VDDA.n2995 3.4105
R2524 VDDA.n3121 VDDA.n2995 3.4105
R2525 VDDA.n3076 VDDA.n2995 3.4105
R2526 VDDA.n2995 VDDA.n18 3.4105
R2527 VDDA.n3123 VDDA.n2995 3.4105
R2528 VDDA.n2964 VDDA.n16 3.4105
R2529 VDDA.n3093 VDDA.n2964 3.4105
R2530 VDDA.n3090 VDDA.n2964 3.4105
R2531 VDDA.n3095 VDDA.n2964 3.4105
R2532 VDDA.n3089 VDDA.n2964 3.4105
R2533 VDDA.n3097 VDDA.n2964 3.4105
R2534 VDDA.n3088 VDDA.n2964 3.4105
R2535 VDDA.n3099 VDDA.n2964 3.4105
R2536 VDDA.n3087 VDDA.n2964 3.4105
R2537 VDDA.n3101 VDDA.n2964 3.4105
R2538 VDDA.n3086 VDDA.n2964 3.4105
R2539 VDDA.n3103 VDDA.n2964 3.4105
R2540 VDDA.n3085 VDDA.n2964 3.4105
R2541 VDDA.n3105 VDDA.n2964 3.4105
R2542 VDDA.n3084 VDDA.n2964 3.4105
R2543 VDDA.n3107 VDDA.n2964 3.4105
R2544 VDDA.n3083 VDDA.n2964 3.4105
R2545 VDDA.n3109 VDDA.n2964 3.4105
R2546 VDDA.n3082 VDDA.n2964 3.4105
R2547 VDDA.n3111 VDDA.n2964 3.4105
R2548 VDDA.n3081 VDDA.n2964 3.4105
R2549 VDDA.n3113 VDDA.n2964 3.4105
R2550 VDDA.n3080 VDDA.n2964 3.4105
R2551 VDDA.n3115 VDDA.n2964 3.4105
R2552 VDDA.n3079 VDDA.n2964 3.4105
R2553 VDDA.n3117 VDDA.n2964 3.4105
R2554 VDDA.n3078 VDDA.n2964 3.4105
R2555 VDDA.n3119 VDDA.n2964 3.4105
R2556 VDDA.n3077 VDDA.n2964 3.4105
R2557 VDDA.n3121 VDDA.n2964 3.4105
R2558 VDDA.n3076 VDDA.n2964 3.4105
R2559 VDDA.n2964 VDDA.n18 3.4105
R2560 VDDA.n3123 VDDA.n2964 3.4105
R2561 VDDA.n2998 VDDA.n16 3.4105
R2562 VDDA.n3093 VDDA.n2998 3.4105
R2563 VDDA.n3090 VDDA.n2998 3.4105
R2564 VDDA.n3095 VDDA.n2998 3.4105
R2565 VDDA.n3089 VDDA.n2998 3.4105
R2566 VDDA.n3097 VDDA.n2998 3.4105
R2567 VDDA.n3088 VDDA.n2998 3.4105
R2568 VDDA.n3099 VDDA.n2998 3.4105
R2569 VDDA.n3087 VDDA.n2998 3.4105
R2570 VDDA.n3101 VDDA.n2998 3.4105
R2571 VDDA.n3086 VDDA.n2998 3.4105
R2572 VDDA.n3103 VDDA.n2998 3.4105
R2573 VDDA.n3085 VDDA.n2998 3.4105
R2574 VDDA.n3105 VDDA.n2998 3.4105
R2575 VDDA.n3084 VDDA.n2998 3.4105
R2576 VDDA.n3107 VDDA.n2998 3.4105
R2577 VDDA.n3083 VDDA.n2998 3.4105
R2578 VDDA.n3109 VDDA.n2998 3.4105
R2579 VDDA.n3082 VDDA.n2998 3.4105
R2580 VDDA.n3111 VDDA.n2998 3.4105
R2581 VDDA.n3081 VDDA.n2998 3.4105
R2582 VDDA.n3113 VDDA.n2998 3.4105
R2583 VDDA.n3080 VDDA.n2998 3.4105
R2584 VDDA.n3115 VDDA.n2998 3.4105
R2585 VDDA.n3079 VDDA.n2998 3.4105
R2586 VDDA.n3117 VDDA.n2998 3.4105
R2587 VDDA.n3078 VDDA.n2998 3.4105
R2588 VDDA.n3119 VDDA.n2998 3.4105
R2589 VDDA.n3077 VDDA.n2998 3.4105
R2590 VDDA.n3121 VDDA.n2998 3.4105
R2591 VDDA.n3076 VDDA.n2998 3.4105
R2592 VDDA.n2998 VDDA.n18 3.4105
R2593 VDDA.n3123 VDDA.n2998 3.4105
R2594 VDDA.n2963 VDDA.n16 3.4105
R2595 VDDA.n3093 VDDA.n2963 3.4105
R2596 VDDA.n3090 VDDA.n2963 3.4105
R2597 VDDA.n3095 VDDA.n2963 3.4105
R2598 VDDA.n3089 VDDA.n2963 3.4105
R2599 VDDA.n3097 VDDA.n2963 3.4105
R2600 VDDA.n3088 VDDA.n2963 3.4105
R2601 VDDA.n3099 VDDA.n2963 3.4105
R2602 VDDA.n3087 VDDA.n2963 3.4105
R2603 VDDA.n3101 VDDA.n2963 3.4105
R2604 VDDA.n3086 VDDA.n2963 3.4105
R2605 VDDA.n3103 VDDA.n2963 3.4105
R2606 VDDA.n3085 VDDA.n2963 3.4105
R2607 VDDA.n3105 VDDA.n2963 3.4105
R2608 VDDA.n3084 VDDA.n2963 3.4105
R2609 VDDA.n3107 VDDA.n2963 3.4105
R2610 VDDA.n3083 VDDA.n2963 3.4105
R2611 VDDA.n3109 VDDA.n2963 3.4105
R2612 VDDA.n3082 VDDA.n2963 3.4105
R2613 VDDA.n3111 VDDA.n2963 3.4105
R2614 VDDA.n3081 VDDA.n2963 3.4105
R2615 VDDA.n3113 VDDA.n2963 3.4105
R2616 VDDA.n3080 VDDA.n2963 3.4105
R2617 VDDA.n3115 VDDA.n2963 3.4105
R2618 VDDA.n3079 VDDA.n2963 3.4105
R2619 VDDA.n3117 VDDA.n2963 3.4105
R2620 VDDA.n3078 VDDA.n2963 3.4105
R2621 VDDA.n3119 VDDA.n2963 3.4105
R2622 VDDA.n3077 VDDA.n2963 3.4105
R2623 VDDA.n3121 VDDA.n2963 3.4105
R2624 VDDA.n3076 VDDA.n2963 3.4105
R2625 VDDA.n2963 VDDA.n18 3.4105
R2626 VDDA.n3123 VDDA.n2963 3.4105
R2627 VDDA.n3001 VDDA.n16 3.4105
R2628 VDDA.n3093 VDDA.n3001 3.4105
R2629 VDDA.n3090 VDDA.n3001 3.4105
R2630 VDDA.n3095 VDDA.n3001 3.4105
R2631 VDDA.n3089 VDDA.n3001 3.4105
R2632 VDDA.n3097 VDDA.n3001 3.4105
R2633 VDDA.n3088 VDDA.n3001 3.4105
R2634 VDDA.n3099 VDDA.n3001 3.4105
R2635 VDDA.n3087 VDDA.n3001 3.4105
R2636 VDDA.n3101 VDDA.n3001 3.4105
R2637 VDDA.n3086 VDDA.n3001 3.4105
R2638 VDDA.n3103 VDDA.n3001 3.4105
R2639 VDDA.n3085 VDDA.n3001 3.4105
R2640 VDDA.n3105 VDDA.n3001 3.4105
R2641 VDDA.n3084 VDDA.n3001 3.4105
R2642 VDDA.n3107 VDDA.n3001 3.4105
R2643 VDDA.n3083 VDDA.n3001 3.4105
R2644 VDDA.n3109 VDDA.n3001 3.4105
R2645 VDDA.n3082 VDDA.n3001 3.4105
R2646 VDDA.n3111 VDDA.n3001 3.4105
R2647 VDDA.n3081 VDDA.n3001 3.4105
R2648 VDDA.n3113 VDDA.n3001 3.4105
R2649 VDDA.n3080 VDDA.n3001 3.4105
R2650 VDDA.n3115 VDDA.n3001 3.4105
R2651 VDDA.n3079 VDDA.n3001 3.4105
R2652 VDDA.n3117 VDDA.n3001 3.4105
R2653 VDDA.n3078 VDDA.n3001 3.4105
R2654 VDDA.n3119 VDDA.n3001 3.4105
R2655 VDDA.n3077 VDDA.n3001 3.4105
R2656 VDDA.n3121 VDDA.n3001 3.4105
R2657 VDDA.n3076 VDDA.n3001 3.4105
R2658 VDDA.n3001 VDDA.n18 3.4105
R2659 VDDA.n3123 VDDA.n3001 3.4105
R2660 VDDA.n2962 VDDA.n16 3.4105
R2661 VDDA.n3093 VDDA.n2962 3.4105
R2662 VDDA.n3090 VDDA.n2962 3.4105
R2663 VDDA.n3095 VDDA.n2962 3.4105
R2664 VDDA.n3089 VDDA.n2962 3.4105
R2665 VDDA.n3097 VDDA.n2962 3.4105
R2666 VDDA.n3088 VDDA.n2962 3.4105
R2667 VDDA.n3099 VDDA.n2962 3.4105
R2668 VDDA.n3087 VDDA.n2962 3.4105
R2669 VDDA.n3101 VDDA.n2962 3.4105
R2670 VDDA.n3086 VDDA.n2962 3.4105
R2671 VDDA.n3103 VDDA.n2962 3.4105
R2672 VDDA.n3085 VDDA.n2962 3.4105
R2673 VDDA.n3105 VDDA.n2962 3.4105
R2674 VDDA.n3084 VDDA.n2962 3.4105
R2675 VDDA.n3107 VDDA.n2962 3.4105
R2676 VDDA.n3083 VDDA.n2962 3.4105
R2677 VDDA.n3109 VDDA.n2962 3.4105
R2678 VDDA.n3082 VDDA.n2962 3.4105
R2679 VDDA.n3111 VDDA.n2962 3.4105
R2680 VDDA.n3081 VDDA.n2962 3.4105
R2681 VDDA.n3113 VDDA.n2962 3.4105
R2682 VDDA.n3080 VDDA.n2962 3.4105
R2683 VDDA.n3115 VDDA.n2962 3.4105
R2684 VDDA.n3079 VDDA.n2962 3.4105
R2685 VDDA.n3117 VDDA.n2962 3.4105
R2686 VDDA.n3078 VDDA.n2962 3.4105
R2687 VDDA.n3119 VDDA.n2962 3.4105
R2688 VDDA.n3077 VDDA.n2962 3.4105
R2689 VDDA.n3121 VDDA.n2962 3.4105
R2690 VDDA.n3076 VDDA.n2962 3.4105
R2691 VDDA.n2962 VDDA.n18 3.4105
R2692 VDDA.n3123 VDDA.n2962 3.4105
R2693 VDDA.n3004 VDDA.n16 3.4105
R2694 VDDA.n3093 VDDA.n3004 3.4105
R2695 VDDA.n3090 VDDA.n3004 3.4105
R2696 VDDA.n3095 VDDA.n3004 3.4105
R2697 VDDA.n3089 VDDA.n3004 3.4105
R2698 VDDA.n3097 VDDA.n3004 3.4105
R2699 VDDA.n3088 VDDA.n3004 3.4105
R2700 VDDA.n3099 VDDA.n3004 3.4105
R2701 VDDA.n3087 VDDA.n3004 3.4105
R2702 VDDA.n3101 VDDA.n3004 3.4105
R2703 VDDA.n3086 VDDA.n3004 3.4105
R2704 VDDA.n3103 VDDA.n3004 3.4105
R2705 VDDA.n3085 VDDA.n3004 3.4105
R2706 VDDA.n3105 VDDA.n3004 3.4105
R2707 VDDA.n3084 VDDA.n3004 3.4105
R2708 VDDA.n3107 VDDA.n3004 3.4105
R2709 VDDA.n3083 VDDA.n3004 3.4105
R2710 VDDA.n3109 VDDA.n3004 3.4105
R2711 VDDA.n3082 VDDA.n3004 3.4105
R2712 VDDA.n3111 VDDA.n3004 3.4105
R2713 VDDA.n3081 VDDA.n3004 3.4105
R2714 VDDA.n3113 VDDA.n3004 3.4105
R2715 VDDA.n3080 VDDA.n3004 3.4105
R2716 VDDA.n3115 VDDA.n3004 3.4105
R2717 VDDA.n3079 VDDA.n3004 3.4105
R2718 VDDA.n3117 VDDA.n3004 3.4105
R2719 VDDA.n3078 VDDA.n3004 3.4105
R2720 VDDA.n3119 VDDA.n3004 3.4105
R2721 VDDA.n3077 VDDA.n3004 3.4105
R2722 VDDA.n3121 VDDA.n3004 3.4105
R2723 VDDA.n3076 VDDA.n3004 3.4105
R2724 VDDA.n3004 VDDA.n18 3.4105
R2725 VDDA.n3123 VDDA.n3004 3.4105
R2726 VDDA.n2961 VDDA.n16 3.4105
R2727 VDDA.n3093 VDDA.n2961 3.4105
R2728 VDDA.n3090 VDDA.n2961 3.4105
R2729 VDDA.n3095 VDDA.n2961 3.4105
R2730 VDDA.n3089 VDDA.n2961 3.4105
R2731 VDDA.n3097 VDDA.n2961 3.4105
R2732 VDDA.n3088 VDDA.n2961 3.4105
R2733 VDDA.n3099 VDDA.n2961 3.4105
R2734 VDDA.n3087 VDDA.n2961 3.4105
R2735 VDDA.n3101 VDDA.n2961 3.4105
R2736 VDDA.n3086 VDDA.n2961 3.4105
R2737 VDDA.n3103 VDDA.n2961 3.4105
R2738 VDDA.n3085 VDDA.n2961 3.4105
R2739 VDDA.n3105 VDDA.n2961 3.4105
R2740 VDDA.n3084 VDDA.n2961 3.4105
R2741 VDDA.n3107 VDDA.n2961 3.4105
R2742 VDDA.n3083 VDDA.n2961 3.4105
R2743 VDDA.n3109 VDDA.n2961 3.4105
R2744 VDDA.n3082 VDDA.n2961 3.4105
R2745 VDDA.n3111 VDDA.n2961 3.4105
R2746 VDDA.n3081 VDDA.n2961 3.4105
R2747 VDDA.n3113 VDDA.n2961 3.4105
R2748 VDDA.n3080 VDDA.n2961 3.4105
R2749 VDDA.n3115 VDDA.n2961 3.4105
R2750 VDDA.n3079 VDDA.n2961 3.4105
R2751 VDDA.n3117 VDDA.n2961 3.4105
R2752 VDDA.n3078 VDDA.n2961 3.4105
R2753 VDDA.n3119 VDDA.n2961 3.4105
R2754 VDDA.n3077 VDDA.n2961 3.4105
R2755 VDDA.n3121 VDDA.n2961 3.4105
R2756 VDDA.n3076 VDDA.n2961 3.4105
R2757 VDDA.n2961 VDDA.n18 3.4105
R2758 VDDA.n3123 VDDA.n2961 3.4105
R2759 VDDA.n3007 VDDA.n16 3.4105
R2760 VDDA.n3093 VDDA.n3007 3.4105
R2761 VDDA.n3090 VDDA.n3007 3.4105
R2762 VDDA.n3095 VDDA.n3007 3.4105
R2763 VDDA.n3089 VDDA.n3007 3.4105
R2764 VDDA.n3097 VDDA.n3007 3.4105
R2765 VDDA.n3088 VDDA.n3007 3.4105
R2766 VDDA.n3099 VDDA.n3007 3.4105
R2767 VDDA.n3087 VDDA.n3007 3.4105
R2768 VDDA.n3101 VDDA.n3007 3.4105
R2769 VDDA.n3086 VDDA.n3007 3.4105
R2770 VDDA.n3103 VDDA.n3007 3.4105
R2771 VDDA.n3085 VDDA.n3007 3.4105
R2772 VDDA.n3105 VDDA.n3007 3.4105
R2773 VDDA.n3084 VDDA.n3007 3.4105
R2774 VDDA.n3107 VDDA.n3007 3.4105
R2775 VDDA.n3083 VDDA.n3007 3.4105
R2776 VDDA.n3109 VDDA.n3007 3.4105
R2777 VDDA.n3082 VDDA.n3007 3.4105
R2778 VDDA.n3111 VDDA.n3007 3.4105
R2779 VDDA.n3081 VDDA.n3007 3.4105
R2780 VDDA.n3113 VDDA.n3007 3.4105
R2781 VDDA.n3080 VDDA.n3007 3.4105
R2782 VDDA.n3115 VDDA.n3007 3.4105
R2783 VDDA.n3079 VDDA.n3007 3.4105
R2784 VDDA.n3117 VDDA.n3007 3.4105
R2785 VDDA.n3078 VDDA.n3007 3.4105
R2786 VDDA.n3119 VDDA.n3007 3.4105
R2787 VDDA.n3077 VDDA.n3007 3.4105
R2788 VDDA.n3121 VDDA.n3007 3.4105
R2789 VDDA.n3076 VDDA.n3007 3.4105
R2790 VDDA.n3007 VDDA.n18 3.4105
R2791 VDDA.n3123 VDDA.n3007 3.4105
R2792 VDDA.n2960 VDDA.n16 3.4105
R2793 VDDA.n3093 VDDA.n2960 3.4105
R2794 VDDA.n3090 VDDA.n2960 3.4105
R2795 VDDA.n3095 VDDA.n2960 3.4105
R2796 VDDA.n3089 VDDA.n2960 3.4105
R2797 VDDA.n3097 VDDA.n2960 3.4105
R2798 VDDA.n3088 VDDA.n2960 3.4105
R2799 VDDA.n3099 VDDA.n2960 3.4105
R2800 VDDA.n3087 VDDA.n2960 3.4105
R2801 VDDA.n3101 VDDA.n2960 3.4105
R2802 VDDA.n3086 VDDA.n2960 3.4105
R2803 VDDA.n3103 VDDA.n2960 3.4105
R2804 VDDA.n3085 VDDA.n2960 3.4105
R2805 VDDA.n3105 VDDA.n2960 3.4105
R2806 VDDA.n3084 VDDA.n2960 3.4105
R2807 VDDA.n3107 VDDA.n2960 3.4105
R2808 VDDA.n3083 VDDA.n2960 3.4105
R2809 VDDA.n3109 VDDA.n2960 3.4105
R2810 VDDA.n3082 VDDA.n2960 3.4105
R2811 VDDA.n3111 VDDA.n2960 3.4105
R2812 VDDA.n3081 VDDA.n2960 3.4105
R2813 VDDA.n3113 VDDA.n2960 3.4105
R2814 VDDA.n3080 VDDA.n2960 3.4105
R2815 VDDA.n3115 VDDA.n2960 3.4105
R2816 VDDA.n3079 VDDA.n2960 3.4105
R2817 VDDA.n3117 VDDA.n2960 3.4105
R2818 VDDA.n3078 VDDA.n2960 3.4105
R2819 VDDA.n3119 VDDA.n2960 3.4105
R2820 VDDA.n3077 VDDA.n2960 3.4105
R2821 VDDA.n3121 VDDA.n2960 3.4105
R2822 VDDA.n3076 VDDA.n2960 3.4105
R2823 VDDA.n2960 VDDA.n18 3.4105
R2824 VDDA.n3123 VDDA.n2960 3.4105
R2825 VDDA.n3010 VDDA.n16 3.4105
R2826 VDDA.n3093 VDDA.n3010 3.4105
R2827 VDDA.n3090 VDDA.n3010 3.4105
R2828 VDDA.n3095 VDDA.n3010 3.4105
R2829 VDDA.n3089 VDDA.n3010 3.4105
R2830 VDDA.n3097 VDDA.n3010 3.4105
R2831 VDDA.n3088 VDDA.n3010 3.4105
R2832 VDDA.n3099 VDDA.n3010 3.4105
R2833 VDDA.n3087 VDDA.n3010 3.4105
R2834 VDDA.n3101 VDDA.n3010 3.4105
R2835 VDDA.n3086 VDDA.n3010 3.4105
R2836 VDDA.n3103 VDDA.n3010 3.4105
R2837 VDDA.n3085 VDDA.n3010 3.4105
R2838 VDDA.n3105 VDDA.n3010 3.4105
R2839 VDDA.n3084 VDDA.n3010 3.4105
R2840 VDDA.n3107 VDDA.n3010 3.4105
R2841 VDDA.n3083 VDDA.n3010 3.4105
R2842 VDDA.n3109 VDDA.n3010 3.4105
R2843 VDDA.n3082 VDDA.n3010 3.4105
R2844 VDDA.n3111 VDDA.n3010 3.4105
R2845 VDDA.n3081 VDDA.n3010 3.4105
R2846 VDDA.n3113 VDDA.n3010 3.4105
R2847 VDDA.n3080 VDDA.n3010 3.4105
R2848 VDDA.n3115 VDDA.n3010 3.4105
R2849 VDDA.n3079 VDDA.n3010 3.4105
R2850 VDDA.n3117 VDDA.n3010 3.4105
R2851 VDDA.n3078 VDDA.n3010 3.4105
R2852 VDDA.n3119 VDDA.n3010 3.4105
R2853 VDDA.n3077 VDDA.n3010 3.4105
R2854 VDDA.n3121 VDDA.n3010 3.4105
R2855 VDDA.n3076 VDDA.n3010 3.4105
R2856 VDDA.n3010 VDDA.n18 3.4105
R2857 VDDA.n3123 VDDA.n3010 3.4105
R2858 VDDA.n2959 VDDA.n16 3.4105
R2859 VDDA.n3093 VDDA.n2959 3.4105
R2860 VDDA.n3090 VDDA.n2959 3.4105
R2861 VDDA.n3095 VDDA.n2959 3.4105
R2862 VDDA.n3089 VDDA.n2959 3.4105
R2863 VDDA.n3097 VDDA.n2959 3.4105
R2864 VDDA.n3088 VDDA.n2959 3.4105
R2865 VDDA.n3099 VDDA.n2959 3.4105
R2866 VDDA.n3087 VDDA.n2959 3.4105
R2867 VDDA.n3101 VDDA.n2959 3.4105
R2868 VDDA.n3086 VDDA.n2959 3.4105
R2869 VDDA.n3103 VDDA.n2959 3.4105
R2870 VDDA.n3085 VDDA.n2959 3.4105
R2871 VDDA.n3105 VDDA.n2959 3.4105
R2872 VDDA.n3084 VDDA.n2959 3.4105
R2873 VDDA.n3107 VDDA.n2959 3.4105
R2874 VDDA.n3083 VDDA.n2959 3.4105
R2875 VDDA.n3109 VDDA.n2959 3.4105
R2876 VDDA.n3082 VDDA.n2959 3.4105
R2877 VDDA.n3111 VDDA.n2959 3.4105
R2878 VDDA.n3081 VDDA.n2959 3.4105
R2879 VDDA.n3113 VDDA.n2959 3.4105
R2880 VDDA.n3080 VDDA.n2959 3.4105
R2881 VDDA.n3115 VDDA.n2959 3.4105
R2882 VDDA.n3079 VDDA.n2959 3.4105
R2883 VDDA.n3117 VDDA.n2959 3.4105
R2884 VDDA.n3078 VDDA.n2959 3.4105
R2885 VDDA.n3119 VDDA.n2959 3.4105
R2886 VDDA.n3077 VDDA.n2959 3.4105
R2887 VDDA.n3121 VDDA.n2959 3.4105
R2888 VDDA.n3076 VDDA.n2959 3.4105
R2889 VDDA.n2959 VDDA.n18 3.4105
R2890 VDDA.n3123 VDDA.n2959 3.4105
R2891 VDDA.n3013 VDDA.n16 3.4105
R2892 VDDA.n3093 VDDA.n3013 3.4105
R2893 VDDA.n3090 VDDA.n3013 3.4105
R2894 VDDA.n3095 VDDA.n3013 3.4105
R2895 VDDA.n3089 VDDA.n3013 3.4105
R2896 VDDA.n3097 VDDA.n3013 3.4105
R2897 VDDA.n3088 VDDA.n3013 3.4105
R2898 VDDA.n3099 VDDA.n3013 3.4105
R2899 VDDA.n3087 VDDA.n3013 3.4105
R2900 VDDA.n3101 VDDA.n3013 3.4105
R2901 VDDA.n3086 VDDA.n3013 3.4105
R2902 VDDA.n3103 VDDA.n3013 3.4105
R2903 VDDA.n3085 VDDA.n3013 3.4105
R2904 VDDA.n3105 VDDA.n3013 3.4105
R2905 VDDA.n3084 VDDA.n3013 3.4105
R2906 VDDA.n3107 VDDA.n3013 3.4105
R2907 VDDA.n3083 VDDA.n3013 3.4105
R2908 VDDA.n3109 VDDA.n3013 3.4105
R2909 VDDA.n3082 VDDA.n3013 3.4105
R2910 VDDA.n3111 VDDA.n3013 3.4105
R2911 VDDA.n3081 VDDA.n3013 3.4105
R2912 VDDA.n3113 VDDA.n3013 3.4105
R2913 VDDA.n3080 VDDA.n3013 3.4105
R2914 VDDA.n3115 VDDA.n3013 3.4105
R2915 VDDA.n3079 VDDA.n3013 3.4105
R2916 VDDA.n3117 VDDA.n3013 3.4105
R2917 VDDA.n3078 VDDA.n3013 3.4105
R2918 VDDA.n3119 VDDA.n3013 3.4105
R2919 VDDA.n3077 VDDA.n3013 3.4105
R2920 VDDA.n3121 VDDA.n3013 3.4105
R2921 VDDA.n3076 VDDA.n3013 3.4105
R2922 VDDA.n3013 VDDA.n18 3.4105
R2923 VDDA.n3123 VDDA.n3013 3.4105
R2924 VDDA.n2958 VDDA.n16 3.4105
R2925 VDDA.n3093 VDDA.n2958 3.4105
R2926 VDDA.n3090 VDDA.n2958 3.4105
R2927 VDDA.n3095 VDDA.n2958 3.4105
R2928 VDDA.n3089 VDDA.n2958 3.4105
R2929 VDDA.n3097 VDDA.n2958 3.4105
R2930 VDDA.n3088 VDDA.n2958 3.4105
R2931 VDDA.n3099 VDDA.n2958 3.4105
R2932 VDDA.n3087 VDDA.n2958 3.4105
R2933 VDDA.n3101 VDDA.n2958 3.4105
R2934 VDDA.n3086 VDDA.n2958 3.4105
R2935 VDDA.n3103 VDDA.n2958 3.4105
R2936 VDDA.n3085 VDDA.n2958 3.4105
R2937 VDDA.n3105 VDDA.n2958 3.4105
R2938 VDDA.n3084 VDDA.n2958 3.4105
R2939 VDDA.n3107 VDDA.n2958 3.4105
R2940 VDDA.n3083 VDDA.n2958 3.4105
R2941 VDDA.n3109 VDDA.n2958 3.4105
R2942 VDDA.n3082 VDDA.n2958 3.4105
R2943 VDDA.n3111 VDDA.n2958 3.4105
R2944 VDDA.n3081 VDDA.n2958 3.4105
R2945 VDDA.n3113 VDDA.n2958 3.4105
R2946 VDDA.n3080 VDDA.n2958 3.4105
R2947 VDDA.n3115 VDDA.n2958 3.4105
R2948 VDDA.n3079 VDDA.n2958 3.4105
R2949 VDDA.n3117 VDDA.n2958 3.4105
R2950 VDDA.n3078 VDDA.n2958 3.4105
R2951 VDDA.n3119 VDDA.n2958 3.4105
R2952 VDDA.n3077 VDDA.n2958 3.4105
R2953 VDDA.n3121 VDDA.n2958 3.4105
R2954 VDDA.n3076 VDDA.n2958 3.4105
R2955 VDDA.n2958 VDDA.n18 3.4105
R2956 VDDA.n3123 VDDA.n2958 3.4105
R2957 VDDA.n3016 VDDA.n16 3.4105
R2958 VDDA.n3093 VDDA.n3016 3.4105
R2959 VDDA.n3090 VDDA.n3016 3.4105
R2960 VDDA.n3095 VDDA.n3016 3.4105
R2961 VDDA.n3089 VDDA.n3016 3.4105
R2962 VDDA.n3097 VDDA.n3016 3.4105
R2963 VDDA.n3088 VDDA.n3016 3.4105
R2964 VDDA.n3099 VDDA.n3016 3.4105
R2965 VDDA.n3087 VDDA.n3016 3.4105
R2966 VDDA.n3101 VDDA.n3016 3.4105
R2967 VDDA.n3086 VDDA.n3016 3.4105
R2968 VDDA.n3103 VDDA.n3016 3.4105
R2969 VDDA.n3085 VDDA.n3016 3.4105
R2970 VDDA.n3105 VDDA.n3016 3.4105
R2971 VDDA.n3084 VDDA.n3016 3.4105
R2972 VDDA.n3107 VDDA.n3016 3.4105
R2973 VDDA.n3083 VDDA.n3016 3.4105
R2974 VDDA.n3109 VDDA.n3016 3.4105
R2975 VDDA.n3082 VDDA.n3016 3.4105
R2976 VDDA.n3111 VDDA.n3016 3.4105
R2977 VDDA.n3081 VDDA.n3016 3.4105
R2978 VDDA.n3113 VDDA.n3016 3.4105
R2979 VDDA.n3080 VDDA.n3016 3.4105
R2980 VDDA.n3115 VDDA.n3016 3.4105
R2981 VDDA.n3079 VDDA.n3016 3.4105
R2982 VDDA.n3117 VDDA.n3016 3.4105
R2983 VDDA.n3078 VDDA.n3016 3.4105
R2984 VDDA.n3119 VDDA.n3016 3.4105
R2985 VDDA.n3077 VDDA.n3016 3.4105
R2986 VDDA.n3121 VDDA.n3016 3.4105
R2987 VDDA.n3076 VDDA.n3016 3.4105
R2988 VDDA.n3016 VDDA.n18 3.4105
R2989 VDDA.n3123 VDDA.n3016 3.4105
R2990 VDDA.n2957 VDDA.n16 3.4105
R2991 VDDA.n3093 VDDA.n2957 3.4105
R2992 VDDA.n3090 VDDA.n2957 3.4105
R2993 VDDA.n3095 VDDA.n2957 3.4105
R2994 VDDA.n3089 VDDA.n2957 3.4105
R2995 VDDA.n3097 VDDA.n2957 3.4105
R2996 VDDA.n3088 VDDA.n2957 3.4105
R2997 VDDA.n3099 VDDA.n2957 3.4105
R2998 VDDA.n3087 VDDA.n2957 3.4105
R2999 VDDA.n3101 VDDA.n2957 3.4105
R3000 VDDA.n3086 VDDA.n2957 3.4105
R3001 VDDA.n3103 VDDA.n2957 3.4105
R3002 VDDA.n3085 VDDA.n2957 3.4105
R3003 VDDA.n3105 VDDA.n2957 3.4105
R3004 VDDA.n3084 VDDA.n2957 3.4105
R3005 VDDA.n3107 VDDA.n2957 3.4105
R3006 VDDA.n3083 VDDA.n2957 3.4105
R3007 VDDA.n3109 VDDA.n2957 3.4105
R3008 VDDA.n3082 VDDA.n2957 3.4105
R3009 VDDA.n3111 VDDA.n2957 3.4105
R3010 VDDA.n3081 VDDA.n2957 3.4105
R3011 VDDA.n3113 VDDA.n2957 3.4105
R3012 VDDA.n3080 VDDA.n2957 3.4105
R3013 VDDA.n3115 VDDA.n2957 3.4105
R3014 VDDA.n3079 VDDA.n2957 3.4105
R3015 VDDA.n3117 VDDA.n2957 3.4105
R3016 VDDA.n3078 VDDA.n2957 3.4105
R3017 VDDA.n3119 VDDA.n2957 3.4105
R3018 VDDA.n3077 VDDA.n2957 3.4105
R3019 VDDA.n3121 VDDA.n2957 3.4105
R3020 VDDA.n3076 VDDA.n2957 3.4105
R3021 VDDA.n2957 VDDA.n18 3.4105
R3022 VDDA.n3123 VDDA.n2957 3.4105
R3023 VDDA.n3019 VDDA.n16 3.4105
R3024 VDDA.n3093 VDDA.n3019 3.4105
R3025 VDDA.n3090 VDDA.n3019 3.4105
R3026 VDDA.n3095 VDDA.n3019 3.4105
R3027 VDDA.n3089 VDDA.n3019 3.4105
R3028 VDDA.n3097 VDDA.n3019 3.4105
R3029 VDDA.n3088 VDDA.n3019 3.4105
R3030 VDDA.n3099 VDDA.n3019 3.4105
R3031 VDDA.n3087 VDDA.n3019 3.4105
R3032 VDDA.n3101 VDDA.n3019 3.4105
R3033 VDDA.n3086 VDDA.n3019 3.4105
R3034 VDDA.n3103 VDDA.n3019 3.4105
R3035 VDDA.n3085 VDDA.n3019 3.4105
R3036 VDDA.n3105 VDDA.n3019 3.4105
R3037 VDDA.n3084 VDDA.n3019 3.4105
R3038 VDDA.n3107 VDDA.n3019 3.4105
R3039 VDDA.n3083 VDDA.n3019 3.4105
R3040 VDDA.n3109 VDDA.n3019 3.4105
R3041 VDDA.n3082 VDDA.n3019 3.4105
R3042 VDDA.n3111 VDDA.n3019 3.4105
R3043 VDDA.n3081 VDDA.n3019 3.4105
R3044 VDDA.n3113 VDDA.n3019 3.4105
R3045 VDDA.n3080 VDDA.n3019 3.4105
R3046 VDDA.n3115 VDDA.n3019 3.4105
R3047 VDDA.n3079 VDDA.n3019 3.4105
R3048 VDDA.n3117 VDDA.n3019 3.4105
R3049 VDDA.n3078 VDDA.n3019 3.4105
R3050 VDDA.n3119 VDDA.n3019 3.4105
R3051 VDDA.n3077 VDDA.n3019 3.4105
R3052 VDDA.n3121 VDDA.n3019 3.4105
R3053 VDDA.n3076 VDDA.n3019 3.4105
R3054 VDDA.n3019 VDDA.n18 3.4105
R3055 VDDA.n3123 VDDA.n3019 3.4105
R3056 VDDA.n2956 VDDA.n16 3.4105
R3057 VDDA.n3093 VDDA.n2956 3.4105
R3058 VDDA.n3090 VDDA.n2956 3.4105
R3059 VDDA.n3095 VDDA.n2956 3.4105
R3060 VDDA.n3089 VDDA.n2956 3.4105
R3061 VDDA.n3097 VDDA.n2956 3.4105
R3062 VDDA.n3088 VDDA.n2956 3.4105
R3063 VDDA.n3099 VDDA.n2956 3.4105
R3064 VDDA.n3087 VDDA.n2956 3.4105
R3065 VDDA.n3101 VDDA.n2956 3.4105
R3066 VDDA.n3086 VDDA.n2956 3.4105
R3067 VDDA.n3103 VDDA.n2956 3.4105
R3068 VDDA.n3085 VDDA.n2956 3.4105
R3069 VDDA.n3105 VDDA.n2956 3.4105
R3070 VDDA.n3084 VDDA.n2956 3.4105
R3071 VDDA.n3107 VDDA.n2956 3.4105
R3072 VDDA.n3083 VDDA.n2956 3.4105
R3073 VDDA.n3109 VDDA.n2956 3.4105
R3074 VDDA.n3082 VDDA.n2956 3.4105
R3075 VDDA.n3111 VDDA.n2956 3.4105
R3076 VDDA.n3081 VDDA.n2956 3.4105
R3077 VDDA.n3113 VDDA.n2956 3.4105
R3078 VDDA.n3080 VDDA.n2956 3.4105
R3079 VDDA.n3115 VDDA.n2956 3.4105
R3080 VDDA.n3079 VDDA.n2956 3.4105
R3081 VDDA.n3117 VDDA.n2956 3.4105
R3082 VDDA.n3078 VDDA.n2956 3.4105
R3083 VDDA.n3119 VDDA.n2956 3.4105
R3084 VDDA.n3077 VDDA.n2956 3.4105
R3085 VDDA.n3121 VDDA.n2956 3.4105
R3086 VDDA.n3076 VDDA.n2956 3.4105
R3087 VDDA.n2956 VDDA.n18 3.4105
R3088 VDDA.n3123 VDDA.n2956 3.4105
R3089 VDDA.n3022 VDDA.n16 3.4105
R3090 VDDA.n3093 VDDA.n3022 3.4105
R3091 VDDA.n3090 VDDA.n3022 3.4105
R3092 VDDA.n3095 VDDA.n3022 3.4105
R3093 VDDA.n3089 VDDA.n3022 3.4105
R3094 VDDA.n3097 VDDA.n3022 3.4105
R3095 VDDA.n3088 VDDA.n3022 3.4105
R3096 VDDA.n3099 VDDA.n3022 3.4105
R3097 VDDA.n3087 VDDA.n3022 3.4105
R3098 VDDA.n3101 VDDA.n3022 3.4105
R3099 VDDA.n3086 VDDA.n3022 3.4105
R3100 VDDA.n3103 VDDA.n3022 3.4105
R3101 VDDA.n3085 VDDA.n3022 3.4105
R3102 VDDA.n3105 VDDA.n3022 3.4105
R3103 VDDA.n3084 VDDA.n3022 3.4105
R3104 VDDA.n3107 VDDA.n3022 3.4105
R3105 VDDA.n3083 VDDA.n3022 3.4105
R3106 VDDA.n3109 VDDA.n3022 3.4105
R3107 VDDA.n3082 VDDA.n3022 3.4105
R3108 VDDA.n3111 VDDA.n3022 3.4105
R3109 VDDA.n3081 VDDA.n3022 3.4105
R3110 VDDA.n3113 VDDA.n3022 3.4105
R3111 VDDA.n3080 VDDA.n3022 3.4105
R3112 VDDA.n3115 VDDA.n3022 3.4105
R3113 VDDA.n3079 VDDA.n3022 3.4105
R3114 VDDA.n3117 VDDA.n3022 3.4105
R3115 VDDA.n3078 VDDA.n3022 3.4105
R3116 VDDA.n3119 VDDA.n3022 3.4105
R3117 VDDA.n3077 VDDA.n3022 3.4105
R3118 VDDA.n3121 VDDA.n3022 3.4105
R3119 VDDA.n3076 VDDA.n3022 3.4105
R3120 VDDA.n3022 VDDA.n18 3.4105
R3121 VDDA.n3123 VDDA.n3022 3.4105
R3122 VDDA.n2955 VDDA.n16 3.4105
R3123 VDDA.n3093 VDDA.n2955 3.4105
R3124 VDDA.n3090 VDDA.n2955 3.4105
R3125 VDDA.n3095 VDDA.n2955 3.4105
R3126 VDDA.n3089 VDDA.n2955 3.4105
R3127 VDDA.n3097 VDDA.n2955 3.4105
R3128 VDDA.n3088 VDDA.n2955 3.4105
R3129 VDDA.n3099 VDDA.n2955 3.4105
R3130 VDDA.n3087 VDDA.n2955 3.4105
R3131 VDDA.n3101 VDDA.n2955 3.4105
R3132 VDDA.n3086 VDDA.n2955 3.4105
R3133 VDDA.n3103 VDDA.n2955 3.4105
R3134 VDDA.n3085 VDDA.n2955 3.4105
R3135 VDDA.n3105 VDDA.n2955 3.4105
R3136 VDDA.n3084 VDDA.n2955 3.4105
R3137 VDDA.n3107 VDDA.n2955 3.4105
R3138 VDDA.n3083 VDDA.n2955 3.4105
R3139 VDDA.n3109 VDDA.n2955 3.4105
R3140 VDDA.n3082 VDDA.n2955 3.4105
R3141 VDDA.n3111 VDDA.n2955 3.4105
R3142 VDDA.n3081 VDDA.n2955 3.4105
R3143 VDDA.n3113 VDDA.n2955 3.4105
R3144 VDDA.n3080 VDDA.n2955 3.4105
R3145 VDDA.n3115 VDDA.n2955 3.4105
R3146 VDDA.n3079 VDDA.n2955 3.4105
R3147 VDDA.n3117 VDDA.n2955 3.4105
R3148 VDDA.n3078 VDDA.n2955 3.4105
R3149 VDDA.n3119 VDDA.n2955 3.4105
R3150 VDDA.n3077 VDDA.n2955 3.4105
R3151 VDDA.n3121 VDDA.n2955 3.4105
R3152 VDDA.n3076 VDDA.n2955 3.4105
R3153 VDDA.n2955 VDDA.n18 3.4105
R3154 VDDA.n3123 VDDA.n2955 3.4105
R3155 VDDA.n3025 VDDA.n16 3.4105
R3156 VDDA.n3093 VDDA.n3025 3.4105
R3157 VDDA.n3090 VDDA.n3025 3.4105
R3158 VDDA.n3095 VDDA.n3025 3.4105
R3159 VDDA.n3089 VDDA.n3025 3.4105
R3160 VDDA.n3097 VDDA.n3025 3.4105
R3161 VDDA.n3088 VDDA.n3025 3.4105
R3162 VDDA.n3099 VDDA.n3025 3.4105
R3163 VDDA.n3087 VDDA.n3025 3.4105
R3164 VDDA.n3101 VDDA.n3025 3.4105
R3165 VDDA.n3086 VDDA.n3025 3.4105
R3166 VDDA.n3103 VDDA.n3025 3.4105
R3167 VDDA.n3085 VDDA.n3025 3.4105
R3168 VDDA.n3105 VDDA.n3025 3.4105
R3169 VDDA.n3084 VDDA.n3025 3.4105
R3170 VDDA.n3107 VDDA.n3025 3.4105
R3171 VDDA.n3083 VDDA.n3025 3.4105
R3172 VDDA.n3109 VDDA.n3025 3.4105
R3173 VDDA.n3082 VDDA.n3025 3.4105
R3174 VDDA.n3111 VDDA.n3025 3.4105
R3175 VDDA.n3081 VDDA.n3025 3.4105
R3176 VDDA.n3113 VDDA.n3025 3.4105
R3177 VDDA.n3080 VDDA.n3025 3.4105
R3178 VDDA.n3115 VDDA.n3025 3.4105
R3179 VDDA.n3079 VDDA.n3025 3.4105
R3180 VDDA.n3117 VDDA.n3025 3.4105
R3181 VDDA.n3078 VDDA.n3025 3.4105
R3182 VDDA.n3119 VDDA.n3025 3.4105
R3183 VDDA.n3077 VDDA.n3025 3.4105
R3184 VDDA.n3121 VDDA.n3025 3.4105
R3185 VDDA.n3076 VDDA.n3025 3.4105
R3186 VDDA.n3025 VDDA.n18 3.4105
R3187 VDDA.n3123 VDDA.n3025 3.4105
R3188 VDDA.n2954 VDDA.n16 3.4105
R3189 VDDA.n3093 VDDA.n2954 3.4105
R3190 VDDA.n3090 VDDA.n2954 3.4105
R3191 VDDA.n3095 VDDA.n2954 3.4105
R3192 VDDA.n3089 VDDA.n2954 3.4105
R3193 VDDA.n3097 VDDA.n2954 3.4105
R3194 VDDA.n3088 VDDA.n2954 3.4105
R3195 VDDA.n3099 VDDA.n2954 3.4105
R3196 VDDA.n3087 VDDA.n2954 3.4105
R3197 VDDA.n3101 VDDA.n2954 3.4105
R3198 VDDA.n3086 VDDA.n2954 3.4105
R3199 VDDA.n3103 VDDA.n2954 3.4105
R3200 VDDA.n3085 VDDA.n2954 3.4105
R3201 VDDA.n3105 VDDA.n2954 3.4105
R3202 VDDA.n3084 VDDA.n2954 3.4105
R3203 VDDA.n3107 VDDA.n2954 3.4105
R3204 VDDA.n3083 VDDA.n2954 3.4105
R3205 VDDA.n3109 VDDA.n2954 3.4105
R3206 VDDA.n3082 VDDA.n2954 3.4105
R3207 VDDA.n3111 VDDA.n2954 3.4105
R3208 VDDA.n3081 VDDA.n2954 3.4105
R3209 VDDA.n3113 VDDA.n2954 3.4105
R3210 VDDA.n3080 VDDA.n2954 3.4105
R3211 VDDA.n3115 VDDA.n2954 3.4105
R3212 VDDA.n3079 VDDA.n2954 3.4105
R3213 VDDA.n3117 VDDA.n2954 3.4105
R3214 VDDA.n3078 VDDA.n2954 3.4105
R3215 VDDA.n3119 VDDA.n2954 3.4105
R3216 VDDA.n3077 VDDA.n2954 3.4105
R3217 VDDA.n3121 VDDA.n2954 3.4105
R3218 VDDA.n3076 VDDA.n2954 3.4105
R3219 VDDA.n2954 VDDA.n18 3.4105
R3220 VDDA.n3123 VDDA.n2954 3.4105
R3221 VDDA.n3028 VDDA.n16 3.4105
R3222 VDDA.n3093 VDDA.n3028 3.4105
R3223 VDDA.n3090 VDDA.n3028 3.4105
R3224 VDDA.n3095 VDDA.n3028 3.4105
R3225 VDDA.n3089 VDDA.n3028 3.4105
R3226 VDDA.n3097 VDDA.n3028 3.4105
R3227 VDDA.n3088 VDDA.n3028 3.4105
R3228 VDDA.n3099 VDDA.n3028 3.4105
R3229 VDDA.n3087 VDDA.n3028 3.4105
R3230 VDDA.n3101 VDDA.n3028 3.4105
R3231 VDDA.n3086 VDDA.n3028 3.4105
R3232 VDDA.n3103 VDDA.n3028 3.4105
R3233 VDDA.n3085 VDDA.n3028 3.4105
R3234 VDDA.n3105 VDDA.n3028 3.4105
R3235 VDDA.n3084 VDDA.n3028 3.4105
R3236 VDDA.n3107 VDDA.n3028 3.4105
R3237 VDDA.n3083 VDDA.n3028 3.4105
R3238 VDDA.n3109 VDDA.n3028 3.4105
R3239 VDDA.n3082 VDDA.n3028 3.4105
R3240 VDDA.n3111 VDDA.n3028 3.4105
R3241 VDDA.n3081 VDDA.n3028 3.4105
R3242 VDDA.n3113 VDDA.n3028 3.4105
R3243 VDDA.n3080 VDDA.n3028 3.4105
R3244 VDDA.n3115 VDDA.n3028 3.4105
R3245 VDDA.n3079 VDDA.n3028 3.4105
R3246 VDDA.n3117 VDDA.n3028 3.4105
R3247 VDDA.n3078 VDDA.n3028 3.4105
R3248 VDDA.n3119 VDDA.n3028 3.4105
R3249 VDDA.n3077 VDDA.n3028 3.4105
R3250 VDDA.n3121 VDDA.n3028 3.4105
R3251 VDDA.n3076 VDDA.n3028 3.4105
R3252 VDDA.n3028 VDDA.n18 3.4105
R3253 VDDA.n3123 VDDA.n3028 3.4105
R3254 VDDA.n2953 VDDA.n16 3.4105
R3255 VDDA.n3093 VDDA.n2953 3.4105
R3256 VDDA.n3090 VDDA.n2953 3.4105
R3257 VDDA.n3095 VDDA.n2953 3.4105
R3258 VDDA.n3089 VDDA.n2953 3.4105
R3259 VDDA.n3097 VDDA.n2953 3.4105
R3260 VDDA.n3088 VDDA.n2953 3.4105
R3261 VDDA.n3099 VDDA.n2953 3.4105
R3262 VDDA.n3087 VDDA.n2953 3.4105
R3263 VDDA.n3101 VDDA.n2953 3.4105
R3264 VDDA.n3086 VDDA.n2953 3.4105
R3265 VDDA.n3103 VDDA.n2953 3.4105
R3266 VDDA.n3085 VDDA.n2953 3.4105
R3267 VDDA.n3105 VDDA.n2953 3.4105
R3268 VDDA.n3084 VDDA.n2953 3.4105
R3269 VDDA.n3107 VDDA.n2953 3.4105
R3270 VDDA.n3083 VDDA.n2953 3.4105
R3271 VDDA.n3109 VDDA.n2953 3.4105
R3272 VDDA.n3082 VDDA.n2953 3.4105
R3273 VDDA.n3111 VDDA.n2953 3.4105
R3274 VDDA.n3081 VDDA.n2953 3.4105
R3275 VDDA.n3113 VDDA.n2953 3.4105
R3276 VDDA.n3080 VDDA.n2953 3.4105
R3277 VDDA.n3115 VDDA.n2953 3.4105
R3278 VDDA.n3079 VDDA.n2953 3.4105
R3279 VDDA.n3117 VDDA.n2953 3.4105
R3280 VDDA.n3078 VDDA.n2953 3.4105
R3281 VDDA.n3119 VDDA.n2953 3.4105
R3282 VDDA.n3077 VDDA.n2953 3.4105
R3283 VDDA.n3121 VDDA.n2953 3.4105
R3284 VDDA.n3076 VDDA.n2953 3.4105
R3285 VDDA.n2953 VDDA.n18 3.4105
R3286 VDDA.n3123 VDDA.n2953 3.4105
R3287 VDDA.n3031 VDDA.n16 3.4105
R3288 VDDA.n3093 VDDA.n3031 3.4105
R3289 VDDA.n3090 VDDA.n3031 3.4105
R3290 VDDA.n3095 VDDA.n3031 3.4105
R3291 VDDA.n3089 VDDA.n3031 3.4105
R3292 VDDA.n3097 VDDA.n3031 3.4105
R3293 VDDA.n3088 VDDA.n3031 3.4105
R3294 VDDA.n3099 VDDA.n3031 3.4105
R3295 VDDA.n3087 VDDA.n3031 3.4105
R3296 VDDA.n3101 VDDA.n3031 3.4105
R3297 VDDA.n3086 VDDA.n3031 3.4105
R3298 VDDA.n3103 VDDA.n3031 3.4105
R3299 VDDA.n3085 VDDA.n3031 3.4105
R3300 VDDA.n3105 VDDA.n3031 3.4105
R3301 VDDA.n3084 VDDA.n3031 3.4105
R3302 VDDA.n3107 VDDA.n3031 3.4105
R3303 VDDA.n3083 VDDA.n3031 3.4105
R3304 VDDA.n3109 VDDA.n3031 3.4105
R3305 VDDA.n3082 VDDA.n3031 3.4105
R3306 VDDA.n3111 VDDA.n3031 3.4105
R3307 VDDA.n3081 VDDA.n3031 3.4105
R3308 VDDA.n3113 VDDA.n3031 3.4105
R3309 VDDA.n3080 VDDA.n3031 3.4105
R3310 VDDA.n3115 VDDA.n3031 3.4105
R3311 VDDA.n3079 VDDA.n3031 3.4105
R3312 VDDA.n3117 VDDA.n3031 3.4105
R3313 VDDA.n3078 VDDA.n3031 3.4105
R3314 VDDA.n3119 VDDA.n3031 3.4105
R3315 VDDA.n3077 VDDA.n3031 3.4105
R3316 VDDA.n3121 VDDA.n3031 3.4105
R3317 VDDA.n3076 VDDA.n3031 3.4105
R3318 VDDA.n3031 VDDA.n18 3.4105
R3319 VDDA.n3123 VDDA.n3031 3.4105
R3320 VDDA.n2952 VDDA.n16 3.4105
R3321 VDDA.n3093 VDDA.n2952 3.4105
R3322 VDDA.n3090 VDDA.n2952 3.4105
R3323 VDDA.n3095 VDDA.n2952 3.4105
R3324 VDDA.n3089 VDDA.n2952 3.4105
R3325 VDDA.n3097 VDDA.n2952 3.4105
R3326 VDDA.n3088 VDDA.n2952 3.4105
R3327 VDDA.n3099 VDDA.n2952 3.4105
R3328 VDDA.n3087 VDDA.n2952 3.4105
R3329 VDDA.n3101 VDDA.n2952 3.4105
R3330 VDDA.n3086 VDDA.n2952 3.4105
R3331 VDDA.n3103 VDDA.n2952 3.4105
R3332 VDDA.n3085 VDDA.n2952 3.4105
R3333 VDDA.n3105 VDDA.n2952 3.4105
R3334 VDDA.n3084 VDDA.n2952 3.4105
R3335 VDDA.n3107 VDDA.n2952 3.4105
R3336 VDDA.n3083 VDDA.n2952 3.4105
R3337 VDDA.n3109 VDDA.n2952 3.4105
R3338 VDDA.n3082 VDDA.n2952 3.4105
R3339 VDDA.n3111 VDDA.n2952 3.4105
R3340 VDDA.n3081 VDDA.n2952 3.4105
R3341 VDDA.n3113 VDDA.n2952 3.4105
R3342 VDDA.n3080 VDDA.n2952 3.4105
R3343 VDDA.n3115 VDDA.n2952 3.4105
R3344 VDDA.n3079 VDDA.n2952 3.4105
R3345 VDDA.n3117 VDDA.n2952 3.4105
R3346 VDDA.n3078 VDDA.n2952 3.4105
R3347 VDDA.n3119 VDDA.n2952 3.4105
R3348 VDDA.n3077 VDDA.n2952 3.4105
R3349 VDDA.n3121 VDDA.n2952 3.4105
R3350 VDDA.n3076 VDDA.n2952 3.4105
R3351 VDDA.n2952 VDDA.n18 3.4105
R3352 VDDA.n3123 VDDA.n2952 3.4105
R3353 VDDA.n3034 VDDA.n16 3.4105
R3354 VDDA.n3093 VDDA.n3034 3.4105
R3355 VDDA.n3090 VDDA.n3034 3.4105
R3356 VDDA.n3095 VDDA.n3034 3.4105
R3357 VDDA.n3089 VDDA.n3034 3.4105
R3358 VDDA.n3097 VDDA.n3034 3.4105
R3359 VDDA.n3088 VDDA.n3034 3.4105
R3360 VDDA.n3099 VDDA.n3034 3.4105
R3361 VDDA.n3087 VDDA.n3034 3.4105
R3362 VDDA.n3101 VDDA.n3034 3.4105
R3363 VDDA.n3086 VDDA.n3034 3.4105
R3364 VDDA.n3103 VDDA.n3034 3.4105
R3365 VDDA.n3085 VDDA.n3034 3.4105
R3366 VDDA.n3105 VDDA.n3034 3.4105
R3367 VDDA.n3084 VDDA.n3034 3.4105
R3368 VDDA.n3107 VDDA.n3034 3.4105
R3369 VDDA.n3083 VDDA.n3034 3.4105
R3370 VDDA.n3109 VDDA.n3034 3.4105
R3371 VDDA.n3082 VDDA.n3034 3.4105
R3372 VDDA.n3111 VDDA.n3034 3.4105
R3373 VDDA.n3081 VDDA.n3034 3.4105
R3374 VDDA.n3113 VDDA.n3034 3.4105
R3375 VDDA.n3080 VDDA.n3034 3.4105
R3376 VDDA.n3115 VDDA.n3034 3.4105
R3377 VDDA.n3079 VDDA.n3034 3.4105
R3378 VDDA.n3117 VDDA.n3034 3.4105
R3379 VDDA.n3078 VDDA.n3034 3.4105
R3380 VDDA.n3119 VDDA.n3034 3.4105
R3381 VDDA.n3077 VDDA.n3034 3.4105
R3382 VDDA.n3121 VDDA.n3034 3.4105
R3383 VDDA.n3076 VDDA.n3034 3.4105
R3384 VDDA.n3034 VDDA.n18 3.4105
R3385 VDDA.n3123 VDDA.n3034 3.4105
R3386 VDDA.n2951 VDDA.n16 3.4105
R3387 VDDA.n3093 VDDA.n2951 3.4105
R3388 VDDA.n3090 VDDA.n2951 3.4105
R3389 VDDA.n3095 VDDA.n2951 3.4105
R3390 VDDA.n3089 VDDA.n2951 3.4105
R3391 VDDA.n3097 VDDA.n2951 3.4105
R3392 VDDA.n3088 VDDA.n2951 3.4105
R3393 VDDA.n3099 VDDA.n2951 3.4105
R3394 VDDA.n3087 VDDA.n2951 3.4105
R3395 VDDA.n3101 VDDA.n2951 3.4105
R3396 VDDA.n3086 VDDA.n2951 3.4105
R3397 VDDA.n3103 VDDA.n2951 3.4105
R3398 VDDA.n3085 VDDA.n2951 3.4105
R3399 VDDA.n3105 VDDA.n2951 3.4105
R3400 VDDA.n3084 VDDA.n2951 3.4105
R3401 VDDA.n3107 VDDA.n2951 3.4105
R3402 VDDA.n3083 VDDA.n2951 3.4105
R3403 VDDA.n3109 VDDA.n2951 3.4105
R3404 VDDA.n3082 VDDA.n2951 3.4105
R3405 VDDA.n3111 VDDA.n2951 3.4105
R3406 VDDA.n3081 VDDA.n2951 3.4105
R3407 VDDA.n3113 VDDA.n2951 3.4105
R3408 VDDA.n3080 VDDA.n2951 3.4105
R3409 VDDA.n3115 VDDA.n2951 3.4105
R3410 VDDA.n3079 VDDA.n2951 3.4105
R3411 VDDA.n3117 VDDA.n2951 3.4105
R3412 VDDA.n3078 VDDA.n2951 3.4105
R3413 VDDA.n3119 VDDA.n2951 3.4105
R3414 VDDA.n3077 VDDA.n2951 3.4105
R3415 VDDA.n3121 VDDA.n2951 3.4105
R3416 VDDA.n3076 VDDA.n2951 3.4105
R3417 VDDA.n2951 VDDA.n18 3.4105
R3418 VDDA.n3123 VDDA.n2951 3.4105
R3419 VDDA.n3037 VDDA.n16 3.4105
R3420 VDDA.n3093 VDDA.n3037 3.4105
R3421 VDDA.n3090 VDDA.n3037 3.4105
R3422 VDDA.n3095 VDDA.n3037 3.4105
R3423 VDDA.n3089 VDDA.n3037 3.4105
R3424 VDDA.n3097 VDDA.n3037 3.4105
R3425 VDDA.n3088 VDDA.n3037 3.4105
R3426 VDDA.n3099 VDDA.n3037 3.4105
R3427 VDDA.n3087 VDDA.n3037 3.4105
R3428 VDDA.n3101 VDDA.n3037 3.4105
R3429 VDDA.n3086 VDDA.n3037 3.4105
R3430 VDDA.n3103 VDDA.n3037 3.4105
R3431 VDDA.n3085 VDDA.n3037 3.4105
R3432 VDDA.n3105 VDDA.n3037 3.4105
R3433 VDDA.n3084 VDDA.n3037 3.4105
R3434 VDDA.n3107 VDDA.n3037 3.4105
R3435 VDDA.n3083 VDDA.n3037 3.4105
R3436 VDDA.n3109 VDDA.n3037 3.4105
R3437 VDDA.n3082 VDDA.n3037 3.4105
R3438 VDDA.n3111 VDDA.n3037 3.4105
R3439 VDDA.n3081 VDDA.n3037 3.4105
R3440 VDDA.n3113 VDDA.n3037 3.4105
R3441 VDDA.n3080 VDDA.n3037 3.4105
R3442 VDDA.n3115 VDDA.n3037 3.4105
R3443 VDDA.n3079 VDDA.n3037 3.4105
R3444 VDDA.n3117 VDDA.n3037 3.4105
R3445 VDDA.n3078 VDDA.n3037 3.4105
R3446 VDDA.n3119 VDDA.n3037 3.4105
R3447 VDDA.n3077 VDDA.n3037 3.4105
R3448 VDDA.n3121 VDDA.n3037 3.4105
R3449 VDDA.n3076 VDDA.n3037 3.4105
R3450 VDDA.n3037 VDDA.n18 3.4105
R3451 VDDA.n3123 VDDA.n3037 3.4105
R3452 VDDA.n2950 VDDA.n16 3.4105
R3453 VDDA.n3093 VDDA.n2950 3.4105
R3454 VDDA.n3090 VDDA.n2950 3.4105
R3455 VDDA.n3095 VDDA.n2950 3.4105
R3456 VDDA.n3089 VDDA.n2950 3.4105
R3457 VDDA.n3097 VDDA.n2950 3.4105
R3458 VDDA.n3088 VDDA.n2950 3.4105
R3459 VDDA.n3099 VDDA.n2950 3.4105
R3460 VDDA.n3087 VDDA.n2950 3.4105
R3461 VDDA.n3101 VDDA.n2950 3.4105
R3462 VDDA.n3086 VDDA.n2950 3.4105
R3463 VDDA.n3103 VDDA.n2950 3.4105
R3464 VDDA.n3085 VDDA.n2950 3.4105
R3465 VDDA.n3105 VDDA.n2950 3.4105
R3466 VDDA.n3084 VDDA.n2950 3.4105
R3467 VDDA.n3107 VDDA.n2950 3.4105
R3468 VDDA.n3083 VDDA.n2950 3.4105
R3469 VDDA.n3109 VDDA.n2950 3.4105
R3470 VDDA.n3082 VDDA.n2950 3.4105
R3471 VDDA.n3111 VDDA.n2950 3.4105
R3472 VDDA.n3081 VDDA.n2950 3.4105
R3473 VDDA.n3113 VDDA.n2950 3.4105
R3474 VDDA.n3080 VDDA.n2950 3.4105
R3475 VDDA.n3115 VDDA.n2950 3.4105
R3476 VDDA.n3079 VDDA.n2950 3.4105
R3477 VDDA.n3117 VDDA.n2950 3.4105
R3478 VDDA.n3078 VDDA.n2950 3.4105
R3479 VDDA.n3119 VDDA.n2950 3.4105
R3480 VDDA.n3077 VDDA.n2950 3.4105
R3481 VDDA.n3121 VDDA.n2950 3.4105
R3482 VDDA.n3076 VDDA.n2950 3.4105
R3483 VDDA.n2950 VDDA.n18 3.4105
R3484 VDDA.n3123 VDDA.n2950 3.4105
R3485 VDDA.n3040 VDDA.n16 3.4105
R3486 VDDA.n3093 VDDA.n3040 3.4105
R3487 VDDA.n3090 VDDA.n3040 3.4105
R3488 VDDA.n3095 VDDA.n3040 3.4105
R3489 VDDA.n3089 VDDA.n3040 3.4105
R3490 VDDA.n3097 VDDA.n3040 3.4105
R3491 VDDA.n3088 VDDA.n3040 3.4105
R3492 VDDA.n3099 VDDA.n3040 3.4105
R3493 VDDA.n3087 VDDA.n3040 3.4105
R3494 VDDA.n3101 VDDA.n3040 3.4105
R3495 VDDA.n3086 VDDA.n3040 3.4105
R3496 VDDA.n3103 VDDA.n3040 3.4105
R3497 VDDA.n3085 VDDA.n3040 3.4105
R3498 VDDA.n3105 VDDA.n3040 3.4105
R3499 VDDA.n3084 VDDA.n3040 3.4105
R3500 VDDA.n3107 VDDA.n3040 3.4105
R3501 VDDA.n3083 VDDA.n3040 3.4105
R3502 VDDA.n3109 VDDA.n3040 3.4105
R3503 VDDA.n3082 VDDA.n3040 3.4105
R3504 VDDA.n3111 VDDA.n3040 3.4105
R3505 VDDA.n3081 VDDA.n3040 3.4105
R3506 VDDA.n3113 VDDA.n3040 3.4105
R3507 VDDA.n3080 VDDA.n3040 3.4105
R3508 VDDA.n3115 VDDA.n3040 3.4105
R3509 VDDA.n3079 VDDA.n3040 3.4105
R3510 VDDA.n3117 VDDA.n3040 3.4105
R3511 VDDA.n3078 VDDA.n3040 3.4105
R3512 VDDA.n3119 VDDA.n3040 3.4105
R3513 VDDA.n3077 VDDA.n3040 3.4105
R3514 VDDA.n3121 VDDA.n3040 3.4105
R3515 VDDA.n3076 VDDA.n3040 3.4105
R3516 VDDA.n3040 VDDA.n18 3.4105
R3517 VDDA.n3123 VDDA.n3040 3.4105
R3518 VDDA.n2949 VDDA.n16 3.4105
R3519 VDDA.n3093 VDDA.n2949 3.4105
R3520 VDDA.n3090 VDDA.n2949 3.4105
R3521 VDDA.n3095 VDDA.n2949 3.4105
R3522 VDDA.n3089 VDDA.n2949 3.4105
R3523 VDDA.n3097 VDDA.n2949 3.4105
R3524 VDDA.n3088 VDDA.n2949 3.4105
R3525 VDDA.n3099 VDDA.n2949 3.4105
R3526 VDDA.n3087 VDDA.n2949 3.4105
R3527 VDDA.n3101 VDDA.n2949 3.4105
R3528 VDDA.n3086 VDDA.n2949 3.4105
R3529 VDDA.n3103 VDDA.n2949 3.4105
R3530 VDDA.n3085 VDDA.n2949 3.4105
R3531 VDDA.n3105 VDDA.n2949 3.4105
R3532 VDDA.n3084 VDDA.n2949 3.4105
R3533 VDDA.n3107 VDDA.n2949 3.4105
R3534 VDDA.n3083 VDDA.n2949 3.4105
R3535 VDDA.n3109 VDDA.n2949 3.4105
R3536 VDDA.n3082 VDDA.n2949 3.4105
R3537 VDDA.n3111 VDDA.n2949 3.4105
R3538 VDDA.n3081 VDDA.n2949 3.4105
R3539 VDDA.n3113 VDDA.n2949 3.4105
R3540 VDDA.n3080 VDDA.n2949 3.4105
R3541 VDDA.n3115 VDDA.n2949 3.4105
R3542 VDDA.n3079 VDDA.n2949 3.4105
R3543 VDDA.n3117 VDDA.n2949 3.4105
R3544 VDDA.n3078 VDDA.n2949 3.4105
R3545 VDDA.n3119 VDDA.n2949 3.4105
R3546 VDDA.n3077 VDDA.n2949 3.4105
R3547 VDDA.n3121 VDDA.n2949 3.4105
R3548 VDDA.n3076 VDDA.n2949 3.4105
R3549 VDDA.n2949 VDDA.n18 3.4105
R3550 VDDA.n3123 VDDA.n2949 3.4105
R3551 VDDA.n3043 VDDA.n16 3.4105
R3552 VDDA.n3093 VDDA.n3043 3.4105
R3553 VDDA.n3090 VDDA.n3043 3.4105
R3554 VDDA.n3095 VDDA.n3043 3.4105
R3555 VDDA.n3089 VDDA.n3043 3.4105
R3556 VDDA.n3097 VDDA.n3043 3.4105
R3557 VDDA.n3088 VDDA.n3043 3.4105
R3558 VDDA.n3099 VDDA.n3043 3.4105
R3559 VDDA.n3087 VDDA.n3043 3.4105
R3560 VDDA.n3101 VDDA.n3043 3.4105
R3561 VDDA.n3086 VDDA.n3043 3.4105
R3562 VDDA.n3103 VDDA.n3043 3.4105
R3563 VDDA.n3085 VDDA.n3043 3.4105
R3564 VDDA.n3105 VDDA.n3043 3.4105
R3565 VDDA.n3084 VDDA.n3043 3.4105
R3566 VDDA.n3107 VDDA.n3043 3.4105
R3567 VDDA.n3083 VDDA.n3043 3.4105
R3568 VDDA.n3109 VDDA.n3043 3.4105
R3569 VDDA.n3082 VDDA.n3043 3.4105
R3570 VDDA.n3111 VDDA.n3043 3.4105
R3571 VDDA.n3081 VDDA.n3043 3.4105
R3572 VDDA.n3113 VDDA.n3043 3.4105
R3573 VDDA.n3080 VDDA.n3043 3.4105
R3574 VDDA.n3115 VDDA.n3043 3.4105
R3575 VDDA.n3079 VDDA.n3043 3.4105
R3576 VDDA.n3117 VDDA.n3043 3.4105
R3577 VDDA.n3078 VDDA.n3043 3.4105
R3578 VDDA.n3119 VDDA.n3043 3.4105
R3579 VDDA.n3077 VDDA.n3043 3.4105
R3580 VDDA.n3121 VDDA.n3043 3.4105
R3581 VDDA.n3076 VDDA.n3043 3.4105
R3582 VDDA.n3043 VDDA.n18 3.4105
R3583 VDDA.n3123 VDDA.n3043 3.4105
R3584 VDDA.n2948 VDDA.n16 3.4105
R3585 VDDA.n3093 VDDA.n2948 3.4105
R3586 VDDA.n3090 VDDA.n2948 3.4105
R3587 VDDA.n3095 VDDA.n2948 3.4105
R3588 VDDA.n3089 VDDA.n2948 3.4105
R3589 VDDA.n3097 VDDA.n2948 3.4105
R3590 VDDA.n3088 VDDA.n2948 3.4105
R3591 VDDA.n3099 VDDA.n2948 3.4105
R3592 VDDA.n3087 VDDA.n2948 3.4105
R3593 VDDA.n3101 VDDA.n2948 3.4105
R3594 VDDA.n3086 VDDA.n2948 3.4105
R3595 VDDA.n3103 VDDA.n2948 3.4105
R3596 VDDA.n3085 VDDA.n2948 3.4105
R3597 VDDA.n3105 VDDA.n2948 3.4105
R3598 VDDA.n3084 VDDA.n2948 3.4105
R3599 VDDA.n3107 VDDA.n2948 3.4105
R3600 VDDA.n3083 VDDA.n2948 3.4105
R3601 VDDA.n3109 VDDA.n2948 3.4105
R3602 VDDA.n3082 VDDA.n2948 3.4105
R3603 VDDA.n3111 VDDA.n2948 3.4105
R3604 VDDA.n3081 VDDA.n2948 3.4105
R3605 VDDA.n3113 VDDA.n2948 3.4105
R3606 VDDA.n3080 VDDA.n2948 3.4105
R3607 VDDA.n3115 VDDA.n2948 3.4105
R3608 VDDA.n3079 VDDA.n2948 3.4105
R3609 VDDA.n3117 VDDA.n2948 3.4105
R3610 VDDA.n3078 VDDA.n2948 3.4105
R3611 VDDA.n3119 VDDA.n2948 3.4105
R3612 VDDA.n3077 VDDA.n2948 3.4105
R3613 VDDA.n3121 VDDA.n2948 3.4105
R3614 VDDA.n3076 VDDA.n2948 3.4105
R3615 VDDA.n2948 VDDA.n18 3.4105
R3616 VDDA.n3123 VDDA.n2948 3.4105
R3617 VDDA.n3046 VDDA.n16 3.4105
R3618 VDDA.n3093 VDDA.n3046 3.4105
R3619 VDDA.n3090 VDDA.n3046 3.4105
R3620 VDDA.n3095 VDDA.n3046 3.4105
R3621 VDDA.n3089 VDDA.n3046 3.4105
R3622 VDDA.n3097 VDDA.n3046 3.4105
R3623 VDDA.n3088 VDDA.n3046 3.4105
R3624 VDDA.n3099 VDDA.n3046 3.4105
R3625 VDDA.n3087 VDDA.n3046 3.4105
R3626 VDDA.n3101 VDDA.n3046 3.4105
R3627 VDDA.n3086 VDDA.n3046 3.4105
R3628 VDDA.n3103 VDDA.n3046 3.4105
R3629 VDDA.n3085 VDDA.n3046 3.4105
R3630 VDDA.n3105 VDDA.n3046 3.4105
R3631 VDDA.n3084 VDDA.n3046 3.4105
R3632 VDDA.n3107 VDDA.n3046 3.4105
R3633 VDDA.n3083 VDDA.n3046 3.4105
R3634 VDDA.n3109 VDDA.n3046 3.4105
R3635 VDDA.n3082 VDDA.n3046 3.4105
R3636 VDDA.n3111 VDDA.n3046 3.4105
R3637 VDDA.n3081 VDDA.n3046 3.4105
R3638 VDDA.n3113 VDDA.n3046 3.4105
R3639 VDDA.n3080 VDDA.n3046 3.4105
R3640 VDDA.n3115 VDDA.n3046 3.4105
R3641 VDDA.n3079 VDDA.n3046 3.4105
R3642 VDDA.n3117 VDDA.n3046 3.4105
R3643 VDDA.n3078 VDDA.n3046 3.4105
R3644 VDDA.n3119 VDDA.n3046 3.4105
R3645 VDDA.n3077 VDDA.n3046 3.4105
R3646 VDDA.n3121 VDDA.n3046 3.4105
R3647 VDDA.n3076 VDDA.n3046 3.4105
R3648 VDDA.n3046 VDDA.n18 3.4105
R3649 VDDA.n3123 VDDA.n3046 3.4105
R3650 VDDA.n2947 VDDA.n16 3.4105
R3651 VDDA.n3093 VDDA.n2947 3.4105
R3652 VDDA.n3090 VDDA.n2947 3.4105
R3653 VDDA.n3095 VDDA.n2947 3.4105
R3654 VDDA.n3089 VDDA.n2947 3.4105
R3655 VDDA.n3097 VDDA.n2947 3.4105
R3656 VDDA.n3088 VDDA.n2947 3.4105
R3657 VDDA.n3099 VDDA.n2947 3.4105
R3658 VDDA.n3087 VDDA.n2947 3.4105
R3659 VDDA.n3101 VDDA.n2947 3.4105
R3660 VDDA.n3086 VDDA.n2947 3.4105
R3661 VDDA.n3103 VDDA.n2947 3.4105
R3662 VDDA.n3085 VDDA.n2947 3.4105
R3663 VDDA.n3105 VDDA.n2947 3.4105
R3664 VDDA.n3084 VDDA.n2947 3.4105
R3665 VDDA.n3107 VDDA.n2947 3.4105
R3666 VDDA.n3083 VDDA.n2947 3.4105
R3667 VDDA.n3109 VDDA.n2947 3.4105
R3668 VDDA.n3082 VDDA.n2947 3.4105
R3669 VDDA.n3111 VDDA.n2947 3.4105
R3670 VDDA.n3081 VDDA.n2947 3.4105
R3671 VDDA.n3113 VDDA.n2947 3.4105
R3672 VDDA.n3080 VDDA.n2947 3.4105
R3673 VDDA.n3115 VDDA.n2947 3.4105
R3674 VDDA.n3079 VDDA.n2947 3.4105
R3675 VDDA.n3117 VDDA.n2947 3.4105
R3676 VDDA.n3078 VDDA.n2947 3.4105
R3677 VDDA.n3119 VDDA.n2947 3.4105
R3678 VDDA.n3077 VDDA.n2947 3.4105
R3679 VDDA.n3121 VDDA.n2947 3.4105
R3680 VDDA.n3076 VDDA.n2947 3.4105
R3681 VDDA.n2947 VDDA.n18 3.4105
R3682 VDDA.n3123 VDDA.n2947 3.4105
R3683 VDDA.n3049 VDDA.n16 3.4105
R3684 VDDA.n3093 VDDA.n3049 3.4105
R3685 VDDA.n3090 VDDA.n3049 3.4105
R3686 VDDA.n3095 VDDA.n3049 3.4105
R3687 VDDA.n3089 VDDA.n3049 3.4105
R3688 VDDA.n3097 VDDA.n3049 3.4105
R3689 VDDA.n3088 VDDA.n3049 3.4105
R3690 VDDA.n3099 VDDA.n3049 3.4105
R3691 VDDA.n3087 VDDA.n3049 3.4105
R3692 VDDA.n3101 VDDA.n3049 3.4105
R3693 VDDA.n3086 VDDA.n3049 3.4105
R3694 VDDA.n3103 VDDA.n3049 3.4105
R3695 VDDA.n3085 VDDA.n3049 3.4105
R3696 VDDA.n3105 VDDA.n3049 3.4105
R3697 VDDA.n3084 VDDA.n3049 3.4105
R3698 VDDA.n3107 VDDA.n3049 3.4105
R3699 VDDA.n3083 VDDA.n3049 3.4105
R3700 VDDA.n3109 VDDA.n3049 3.4105
R3701 VDDA.n3082 VDDA.n3049 3.4105
R3702 VDDA.n3111 VDDA.n3049 3.4105
R3703 VDDA.n3081 VDDA.n3049 3.4105
R3704 VDDA.n3113 VDDA.n3049 3.4105
R3705 VDDA.n3080 VDDA.n3049 3.4105
R3706 VDDA.n3115 VDDA.n3049 3.4105
R3707 VDDA.n3079 VDDA.n3049 3.4105
R3708 VDDA.n3117 VDDA.n3049 3.4105
R3709 VDDA.n3078 VDDA.n3049 3.4105
R3710 VDDA.n3119 VDDA.n3049 3.4105
R3711 VDDA.n3077 VDDA.n3049 3.4105
R3712 VDDA.n3121 VDDA.n3049 3.4105
R3713 VDDA.n3076 VDDA.n3049 3.4105
R3714 VDDA.n3049 VDDA.n18 3.4105
R3715 VDDA.n3123 VDDA.n3049 3.4105
R3716 VDDA.n2946 VDDA.n16 3.4105
R3717 VDDA.n3093 VDDA.n2946 3.4105
R3718 VDDA.n3090 VDDA.n2946 3.4105
R3719 VDDA.n3095 VDDA.n2946 3.4105
R3720 VDDA.n3089 VDDA.n2946 3.4105
R3721 VDDA.n3097 VDDA.n2946 3.4105
R3722 VDDA.n3088 VDDA.n2946 3.4105
R3723 VDDA.n3099 VDDA.n2946 3.4105
R3724 VDDA.n3087 VDDA.n2946 3.4105
R3725 VDDA.n3101 VDDA.n2946 3.4105
R3726 VDDA.n3086 VDDA.n2946 3.4105
R3727 VDDA.n3103 VDDA.n2946 3.4105
R3728 VDDA.n3085 VDDA.n2946 3.4105
R3729 VDDA.n3105 VDDA.n2946 3.4105
R3730 VDDA.n3084 VDDA.n2946 3.4105
R3731 VDDA.n3107 VDDA.n2946 3.4105
R3732 VDDA.n3083 VDDA.n2946 3.4105
R3733 VDDA.n3109 VDDA.n2946 3.4105
R3734 VDDA.n3082 VDDA.n2946 3.4105
R3735 VDDA.n3111 VDDA.n2946 3.4105
R3736 VDDA.n3081 VDDA.n2946 3.4105
R3737 VDDA.n3113 VDDA.n2946 3.4105
R3738 VDDA.n3080 VDDA.n2946 3.4105
R3739 VDDA.n3115 VDDA.n2946 3.4105
R3740 VDDA.n3079 VDDA.n2946 3.4105
R3741 VDDA.n3117 VDDA.n2946 3.4105
R3742 VDDA.n3078 VDDA.n2946 3.4105
R3743 VDDA.n3119 VDDA.n2946 3.4105
R3744 VDDA.n3077 VDDA.n2946 3.4105
R3745 VDDA.n3121 VDDA.n2946 3.4105
R3746 VDDA.n3076 VDDA.n2946 3.4105
R3747 VDDA.n2946 VDDA.n18 3.4105
R3748 VDDA.n3123 VDDA.n2946 3.4105
R3749 VDDA.n3052 VDDA.n16 3.4105
R3750 VDDA.n3093 VDDA.n3052 3.4105
R3751 VDDA.n3090 VDDA.n3052 3.4105
R3752 VDDA.n3095 VDDA.n3052 3.4105
R3753 VDDA.n3089 VDDA.n3052 3.4105
R3754 VDDA.n3097 VDDA.n3052 3.4105
R3755 VDDA.n3088 VDDA.n3052 3.4105
R3756 VDDA.n3099 VDDA.n3052 3.4105
R3757 VDDA.n3087 VDDA.n3052 3.4105
R3758 VDDA.n3101 VDDA.n3052 3.4105
R3759 VDDA.n3086 VDDA.n3052 3.4105
R3760 VDDA.n3103 VDDA.n3052 3.4105
R3761 VDDA.n3085 VDDA.n3052 3.4105
R3762 VDDA.n3105 VDDA.n3052 3.4105
R3763 VDDA.n3084 VDDA.n3052 3.4105
R3764 VDDA.n3107 VDDA.n3052 3.4105
R3765 VDDA.n3083 VDDA.n3052 3.4105
R3766 VDDA.n3109 VDDA.n3052 3.4105
R3767 VDDA.n3082 VDDA.n3052 3.4105
R3768 VDDA.n3111 VDDA.n3052 3.4105
R3769 VDDA.n3081 VDDA.n3052 3.4105
R3770 VDDA.n3113 VDDA.n3052 3.4105
R3771 VDDA.n3080 VDDA.n3052 3.4105
R3772 VDDA.n3115 VDDA.n3052 3.4105
R3773 VDDA.n3079 VDDA.n3052 3.4105
R3774 VDDA.n3117 VDDA.n3052 3.4105
R3775 VDDA.n3078 VDDA.n3052 3.4105
R3776 VDDA.n3119 VDDA.n3052 3.4105
R3777 VDDA.n3077 VDDA.n3052 3.4105
R3778 VDDA.n3121 VDDA.n3052 3.4105
R3779 VDDA.n3076 VDDA.n3052 3.4105
R3780 VDDA.n3052 VDDA.n18 3.4105
R3781 VDDA.n3123 VDDA.n3052 3.4105
R3782 VDDA.n2945 VDDA.n16 3.4105
R3783 VDDA.n3093 VDDA.n2945 3.4105
R3784 VDDA.n3090 VDDA.n2945 3.4105
R3785 VDDA.n3095 VDDA.n2945 3.4105
R3786 VDDA.n3089 VDDA.n2945 3.4105
R3787 VDDA.n3097 VDDA.n2945 3.4105
R3788 VDDA.n3088 VDDA.n2945 3.4105
R3789 VDDA.n3099 VDDA.n2945 3.4105
R3790 VDDA.n3087 VDDA.n2945 3.4105
R3791 VDDA.n3101 VDDA.n2945 3.4105
R3792 VDDA.n3086 VDDA.n2945 3.4105
R3793 VDDA.n3103 VDDA.n2945 3.4105
R3794 VDDA.n3085 VDDA.n2945 3.4105
R3795 VDDA.n3105 VDDA.n2945 3.4105
R3796 VDDA.n3084 VDDA.n2945 3.4105
R3797 VDDA.n3107 VDDA.n2945 3.4105
R3798 VDDA.n3083 VDDA.n2945 3.4105
R3799 VDDA.n3109 VDDA.n2945 3.4105
R3800 VDDA.n3082 VDDA.n2945 3.4105
R3801 VDDA.n3111 VDDA.n2945 3.4105
R3802 VDDA.n3081 VDDA.n2945 3.4105
R3803 VDDA.n3113 VDDA.n2945 3.4105
R3804 VDDA.n3080 VDDA.n2945 3.4105
R3805 VDDA.n3115 VDDA.n2945 3.4105
R3806 VDDA.n3079 VDDA.n2945 3.4105
R3807 VDDA.n3117 VDDA.n2945 3.4105
R3808 VDDA.n3078 VDDA.n2945 3.4105
R3809 VDDA.n3119 VDDA.n2945 3.4105
R3810 VDDA.n3077 VDDA.n2945 3.4105
R3811 VDDA.n3121 VDDA.n2945 3.4105
R3812 VDDA.n3076 VDDA.n2945 3.4105
R3813 VDDA.n2945 VDDA.n18 3.4105
R3814 VDDA.n3123 VDDA.n2945 3.4105
R3815 VDDA.n3055 VDDA.n16 3.4105
R3816 VDDA.n3093 VDDA.n3055 3.4105
R3817 VDDA.n3090 VDDA.n3055 3.4105
R3818 VDDA.n3095 VDDA.n3055 3.4105
R3819 VDDA.n3089 VDDA.n3055 3.4105
R3820 VDDA.n3097 VDDA.n3055 3.4105
R3821 VDDA.n3088 VDDA.n3055 3.4105
R3822 VDDA.n3099 VDDA.n3055 3.4105
R3823 VDDA.n3087 VDDA.n3055 3.4105
R3824 VDDA.n3101 VDDA.n3055 3.4105
R3825 VDDA.n3086 VDDA.n3055 3.4105
R3826 VDDA.n3103 VDDA.n3055 3.4105
R3827 VDDA.n3085 VDDA.n3055 3.4105
R3828 VDDA.n3105 VDDA.n3055 3.4105
R3829 VDDA.n3084 VDDA.n3055 3.4105
R3830 VDDA.n3107 VDDA.n3055 3.4105
R3831 VDDA.n3083 VDDA.n3055 3.4105
R3832 VDDA.n3109 VDDA.n3055 3.4105
R3833 VDDA.n3082 VDDA.n3055 3.4105
R3834 VDDA.n3111 VDDA.n3055 3.4105
R3835 VDDA.n3081 VDDA.n3055 3.4105
R3836 VDDA.n3113 VDDA.n3055 3.4105
R3837 VDDA.n3080 VDDA.n3055 3.4105
R3838 VDDA.n3115 VDDA.n3055 3.4105
R3839 VDDA.n3079 VDDA.n3055 3.4105
R3840 VDDA.n3117 VDDA.n3055 3.4105
R3841 VDDA.n3078 VDDA.n3055 3.4105
R3842 VDDA.n3119 VDDA.n3055 3.4105
R3843 VDDA.n3077 VDDA.n3055 3.4105
R3844 VDDA.n3121 VDDA.n3055 3.4105
R3845 VDDA.n3076 VDDA.n3055 3.4105
R3846 VDDA.n3055 VDDA.n18 3.4105
R3847 VDDA.n3123 VDDA.n3055 3.4105
R3848 VDDA.n2944 VDDA.n16 3.4105
R3849 VDDA.n3093 VDDA.n2944 3.4105
R3850 VDDA.n3090 VDDA.n2944 3.4105
R3851 VDDA.n3095 VDDA.n2944 3.4105
R3852 VDDA.n3089 VDDA.n2944 3.4105
R3853 VDDA.n3097 VDDA.n2944 3.4105
R3854 VDDA.n3088 VDDA.n2944 3.4105
R3855 VDDA.n3099 VDDA.n2944 3.4105
R3856 VDDA.n3087 VDDA.n2944 3.4105
R3857 VDDA.n3101 VDDA.n2944 3.4105
R3858 VDDA.n3086 VDDA.n2944 3.4105
R3859 VDDA.n3103 VDDA.n2944 3.4105
R3860 VDDA.n3085 VDDA.n2944 3.4105
R3861 VDDA.n3105 VDDA.n2944 3.4105
R3862 VDDA.n3084 VDDA.n2944 3.4105
R3863 VDDA.n3107 VDDA.n2944 3.4105
R3864 VDDA.n3083 VDDA.n2944 3.4105
R3865 VDDA.n3109 VDDA.n2944 3.4105
R3866 VDDA.n3082 VDDA.n2944 3.4105
R3867 VDDA.n3111 VDDA.n2944 3.4105
R3868 VDDA.n3081 VDDA.n2944 3.4105
R3869 VDDA.n3113 VDDA.n2944 3.4105
R3870 VDDA.n3080 VDDA.n2944 3.4105
R3871 VDDA.n3115 VDDA.n2944 3.4105
R3872 VDDA.n3079 VDDA.n2944 3.4105
R3873 VDDA.n3117 VDDA.n2944 3.4105
R3874 VDDA.n3078 VDDA.n2944 3.4105
R3875 VDDA.n3119 VDDA.n2944 3.4105
R3876 VDDA.n3077 VDDA.n2944 3.4105
R3877 VDDA.n3121 VDDA.n2944 3.4105
R3878 VDDA.n3076 VDDA.n2944 3.4105
R3879 VDDA.n2944 VDDA.n18 3.4105
R3880 VDDA.n3123 VDDA.n2944 3.4105
R3881 VDDA.n3058 VDDA.n16 3.4105
R3882 VDDA.n3093 VDDA.n3058 3.4105
R3883 VDDA.n3090 VDDA.n3058 3.4105
R3884 VDDA.n3095 VDDA.n3058 3.4105
R3885 VDDA.n3089 VDDA.n3058 3.4105
R3886 VDDA.n3097 VDDA.n3058 3.4105
R3887 VDDA.n3088 VDDA.n3058 3.4105
R3888 VDDA.n3099 VDDA.n3058 3.4105
R3889 VDDA.n3087 VDDA.n3058 3.4105
R3890 VDDA.n3101 VDDA.n3058 3.4105
R3891 VDDA.n3086 VDDA.n3058 3.4105
R3892 VDDA.n3103 VDDA.n3058 3.4105
R3893 VDDA.n3085 VDDA.n3058 3.4105
R3894 VDDA.n3105 VDDA.n3058 3.4105
R3895 VDDA.n3084 VDDA.n3058 3.4105
R3896 VDDA.n3107 VDDA.n3058 3.4105
R3897 VDDA.n3083 VDDA.n3058 3.4105
R3898 VDDA.n3109 VDDA.n3058 3.4105
R3899 VDDA.n3082 VDDA.n3058 3.4105
R3900 VDDA.n3111 VDDA.n3058 3.4105
R3901 VDDA.n3081 VDDA.n3058 3.4105
R3902 VDDA.n3113 VDDA.n3058 3.4105
R3903 VDDA.n3080 VDDA.n3058 3.4105
R3904 VDDA.n3115 VDDA.n3058 3.4105
R3905 VDDA.n3079 VDDA.n3058 3.4105
R3906 VDDA.n3117 VDDA.n3058 3.4105
R3907 VDDA.n3078 VDDA.n3058 3.4105
R3908 VDDA.n3119 VDDA.n3058 3.4105
R3909 VDDA.n3077 VDDA.n3058 3.4105
R3910 VDDA.n3121 VDDA.n3058 3.4105
R3911 VDDA.n3076 VDDA.n3058 3.4105
R3912 VDDA.n3058 VDDA.n18 3.4105
R3913 VDDA.n3123 VDDA.n3058 3.4105
R3914 VDDA.n2943 VDDA.n16 3.4105
R3915 VDDA.n3093 VDDA.n2943 3.4105
R3916 VDDA.n3090 VDDA.n2943 3.4105
R3917 VDDA.n3095 VDDA.n2943 3.4105
R3918 VDDA.n3089 VDDA.n2943 3.4105
R3919 VDDA.n3097 VDDA.n2943 3.4105
R3920 VDDA.n3088 VDDA.n2943 3.4105
R3921 VDDA.n3099 VDDA.n2943 3.4105
R3922 VDDA.n3087 VDDA.n2943 3.4105
R3923 VDDA.n3101 VDDA.n2943 3.4105
R3924 VDDA.n3086 VDDA.n2943 3.4105
R3925 VDDA.n3103 VDDA.n2943 3.4105
R3926 VDDA.n3085 VDDA.n2943 3.4105
R3927 VDDA.n3105 VDDA.n2943 3.4105
R3928 VDDA.n3084 VDDA.n2943 3.4105
R3929 VDDA.n3107 VDDA.n2943 3.4105
R3930 VDDA.n3083 VDDA.n2943 3.4105
R3931 VDDA.n3109 VDDA.n2943 3.4105
R3932 VDDA.n3082 VDDA.n2943 3.4105
R3933 VDDA.n3111 VDDA.n2943 3.4105
R3934 VDDA.n3081 VDDA.n2943 3.4105
R3935 VDDA.n3113 VDDA.n2943 3.4105
R3936 VDDA.n3080 VDDA.n2943 3.4105
R3937 VDDA.n3115 VDDA.n2943 3.4105
R3938 VDDA.n3079 VDDA.n2943 3.4105
R3939 VDDA.n3117 VDDA.n2943 3.4105
R3940 VDDA.n3078 VDDA.n2943 3.4105
R3941 VDDA.n3119 VDDA.n2943 3.4105
R3942 VDDA.n3077 VDDA.n2943 3.4105
R3943 VDDA.n3121 VDDA.n2943 3.4105
R3944 VDDA.n3076 VDDA.n2943 3.4105
R3945 VDDA.n2943 VDDA.n18 3.4105
R3946 VDDA.n3123 VDDA.n2943 3.4105
R3947 VDDA.n3061 VDDA.n16 3.4105
R3948 VDDA.n3093 VDDA.n3061 3.4105
R3949 VDDA.n3090 VDDA.n3061 3.4105
R3950 VDDA.n3095 VDDA.n3061 3.4105
R3951 VDDA.n3089 VDDA.n3061 3.4105
R3952 VDDA.n3097 VDDA.n3061 3.4105
R3953 VDDA.n3088 VDDA.n3061 3.4105
R3954 VDDA.n3099 VDDA.n3061 3.4105
R3955 VDDA.n3087 VDDA.n3061 3.4105
R3956 VDDA.n3101 VDDA.n3061 3.4105
R3957 VDDA.n3086 VDDA.n3061 3.4105
R3958 VDDA.n3103 VDDA.n3061 3.4105
R3959 VDDA.n3085 VDDA.n3061 3.4105
R3960 VDDA.n3105 VDDA.n3061 3.4105
R3961 VDDA.n3084 VDDA.n3061 3.4105
R3962 VDDA.n3107 VDDA.n3061 3.4105
R3963 VDDA.n3083 VDDA.n3061 3.4105
R3964 VDDA.n3109 VDDA.n3061 3.4105
R3965 VDDA.n3082 VDDA.n3061 3.4105
R3966 VDDA.n3111 VDDA.n3061 3.4105
R3967 VDDA.n3081 VDDA.n3061 3.4105
R3968 VDDA.n3113 VDDA.n3061 3.4105
R3969 VDDA.n3080 VDDA.n3061 3.4105
R3970 VDDA.n3115 VDDA.n3061 3.4105
R3971 VDDA.n3079 VDDA.n3061 3.4105
R3972 VDDA.n3117 VDDA.n3061 3.4105
R3973 VDDA.n3078 VDDA.n3061 3.4105
R3974 VDDA.n3119 VDDA.n3061 3.4105
R3975 VDDA.n3077 VDDA.n3061 3.4105
R3976 VDDA.n3121 VDDA.n3061 3.4105
R3977 VDDA.n3076 VDDA.n3061 3.4105
R3978 VDDA.n3061 VDDA.n18 3.4105
R3979 VDDA.n3123 VDDA.n3061 3.4105
R3980 VDDA.n2942 VDDA.n16 3.4105
R3981 VDDA.n3093 VDDA.n2942 3.4105
R3982 VDDA.n3090 VDDA.n2942 3.4105
R3983 VDDA.n3095 VDDA.n2942 3.4105
R3984 VDDA.n3089 VDDA.n2942 3.4105
R3985 VDDA.n3097 VDDA.n2942 3.4105
R3986 VDDA.n3088 VDDA.n2942 3.4105
R3987 VDDA.n3099 VDDA.n2942 3.4105
R3988 VDDA.n3087 VDDA.n2942 3.4105
R3989 VDDA.n3101 VDDA.n2942 3.4105
R3990 VDDA.n3086 VDDA.n2942 3.4105
R3991 VDDA.n3103 VDDA.n2942 3.4105
R3992 VDDA.n3085 VDDA.n2942 3.4105
R3993 VDDA.n3105 VDDA.n2942 3.4105
R3994 VDDA.n3084 VDDA.n2942 3.4105
R3995 VDDA.n3107 VDDA.n2942 3.4105
R3996 VDDA.n3083 VDDA.n2942 3.4105
R3997 VDDA.n3109 VDDA.n2942 3.4105
R3998 VDDA.n3082 VDDA.n2942 3.4105
R3999 VDDA.n3111 VDDA.n2942 3.4105
R4000 VDDA.n3081 VDDA.n2942 3.4105
R4001 VDDA.n3113 VDDA.n2942 3.4105
R4002 VDDA.n3080 VDDA.n2942 3.4105
R4003 VDDA.n3115 VDDA.n2942 3.4105
R4004 VDDA.n3079 VDDA.n2942 3.4105
R4005 VDDA.n3117 VDDA.n2942 3.4105
R4006 VDDA.n3078 VDDA.n2942 3.4105
R4007 VDDA.n3119 VDDA.n2942 3.4105
R4008 VDDA.n3077 VDDA.n2942 3.4105
R4009 VDDA.n3121 VDDA.n2942 3.4105
R4010 VDDA.n3076 VDDA.n2942 3.4105
R4011 VDDA.n2942 VDDA.n18 3.4105
R4012 VDDA.n3123 VDDA.n2942 3.4105
R4013 VDDA.n3064 VDDA.n16 3.4105
R4014 VDDA.n3093 VDDA.n3064 3.4105
R4015 VDDA.n3090 VDDA.n3064 3.4105
R4016 VDDA.n3095 VDDA.n3064 3.4105
R4017 VDDA.n3089 VDDA.n3064 3.4105
R4018 VDDA.n3097 VDDA.n3064 3.4105
R4019 VDDA.n3088 VDDA.n3064 3.4105
R4020 VDDA.n3099 VDDA.n3064 3.4105
R4021 VDDA.n3087 VDDA.n3064 3.4105
R4022 VDDA.n3101 VDDA.n3064 3.4105
R4023 VDDA.n3086 VDDA.n3064 3.4105
R4024 VDDA.n3103 VDDA.n3064 3.4105
R4025 VDDA.n3085 VDDA.n3064 3.4105
R4026 VDDA.n3105 VDDA.n3064 3.4105
R4027 VDDA.n3084 VDDA.n3064 3.4105
R4028 VDDA.n3107 VDDA.n3064 3.4105
R4029 VDDA.n3083 VDDA.n3064 3.4105
R4030 VDDA.n3109 VDDA.n3064 3.4105
R4031 VDDA.n3082 VDDA.n3064 3.4105
R4032 VDDA.n3111 VDDA.n3064 3.4105
R4033 VDDA.n3081 VDDA.n3064 3.4105
R4034 VDDA.n3113 VDDA.n3064 3.4105
R4035 VDDA.n3080 VDDA.n3064 3.4105
R4036 VDDA.n3115 VDDA.n3064 3.4105
R4037 VDDA.n3079 VDDA.n3064 3.4105
R4038 VDDA.n3117 VDDA.n3064 3.4105
R4039 VDDA.n3078 VDDA.n3064 3.4105
R4040 VDDA.n3119 VDDA.n3064 3.4105
R4041 VDDA.n3077 VDDA.n3064 3.4105
R4042 VDDA.n3121 VDDA.n3064 3.4105
R4043 VDDA.n3076 VDDA.n3064 3.4105
R4044 VDDA.n3064 VDDA.n18 3.4105
R4045 VDDA.n3123 VDDA.n3064 3.4105
R4046 VDDA.n2941 VDDA.n16 3.4105
R4047 VDDA.n3093 VDDA.n2941 3.4105
R4048 VDDA.n3090 VDDA.n2941 3.4105
R4049 VDDA.n3095 VDDA.n2941 3.4105
R4050 VDDA.n3089 VDDA.n2941 3.4105
R4051 VDDA.n3097 VDDA.n2941 3.4105
R4052 VDDA.n3088 VDDA.n2941 3.4105
R4053 VDDA.n3099 VDDA.n2941 3.4105
R4054 VDDA.n3087 VDDA.n2941 3.4105
R4055 VDDA.n3101 VDDA.n2941 3.4105
R4056 VDDA.n3086 VDDA.n2941 3.4105
R4057 VDDA.n3103 VDDA.n2941 3.4105
R4058 VDDA.n3085 VDDA.n2941 3.4105
R4059 VDDA.n3105 VDDA.n2941 3.4105
R4060 VDDA.n3084 VDDA.n2941 3.4105
R4061 VDDA.n3107 VDDA.n2941 3.4105
R4062 VDDA.n3083 VDDA.n2941 3.4105
R4063 VDDA.n3109 VDDA.n2941 3.4105
R4064 VDDA.n3082 VDDA.n2941 3.4105
R4065 VDDA.n3111 VDDA.n2941 3.4105
R4066 VDDA.n3081 VDDA.n2941 3.4105
R4067 VDDA.n3113 VDDA.n2941 3.4105
R4068 VDDA.n3080 VDDA.n2941 3.4105
R4069 VDDA.n3115 VDDA.n2941 3.4105
R4070 VDDA.n3079 VDDA.n2941 3.4105
R4071 VDDA.n3117 VDDA.n2941 3.4105
R4072 VDDA.n3078 VDDA.n2941 3.4105
R4073 VDDA.n3119 VDDA.n2941 3.4105
R4074 VDDA.n3077 VDDA.n2941 3.4105
R4075 VDDA.n3121 VDDA.n2941 3.4105
R4076 VDDA.n3076 VDDA.n2941 3.4105
R4077 VDDA.n2941 VDDA.n18 3.4105
R4078 VDDA.n3123 VDDA.n2941 3.4105
R4079 VDDA.n3067 VDDA.n16 3.4105
R4080 VDDA.n3093 VDDA.n3067 3.4105
R4081 VDDA.n3090 VDDA.n3067 3.4105
R4082 VDDA.n3095 VDDA.n3067 3.4105
R4083 VDDA.n3089 VDDA.n3067 3.4105
R4084 VDDA.n3097 VDDA.n3067 3.4105
R4085 VDDA.n3088 VDDA.n3067 3.4105
R4086 VDDA.n3099 VDDA.n3067 3.4105
R4087 VDDA.n3087 VDDA.n3067 3.4105
R4088 VDDA.n3101 VDDA.n3067 3.4105
R4089 VDDA.n3086 VDDA.n3067 3.4105
R4090 VDDA.n3103 VDDA.n3067 3.4105
R4091 VDDA.n3085 VDDA.n3067 3.4105
R4092 VDDA.n3105 VDDA.n3067 3.4105
R4093 VDDA.n3084 VDDA.n3067 3.4105
R4094 VDDA.n3107 VDDA.n3067 3.4105
R4095 VDDA.n3083 VDDA.n3067 3.4105
R4096 VDDA.n3109 VDDA.n3067 3.4105
R4097 VDDA.n3082 VDDA.n3067 3.4105
R4098 VDDA.n3111 VDDA.n3067 3.4105
R4099 VDDA.n3081 VDDA.n3067 3.4105
R4100 VDDA.n3113 VDDA.n3067 3.4105
R4101 VDDA.n3080 VDDA.n3067 3.4105
R4102 VDDA.n3115 VDDA.n3067 3.4105
R4103 VDDA.n3079 VDDA.n3067 3.4105
R4104 VDDA.n3117 VDDA.n3067 3.4105
R4105 VDDA.n3078 VDDA.n3067 3.4105
R4106 VDDA.n3119 VDDA.n3067 3.4105
R4107 VDDA.n3077 VDDA.n3067 3.4105
R4108 VDDA.n3121 VDDA.n3067 3.4105
R4109 VDDA.n3076 VDDA.n3067 3.4105
R4110 VDDA.n3067 VDDA.n18 3.4105
R4111 VDDA.n3123 VDDA.n3067 3.4105
R4112 VDDA.n2940 VDDA.n16 3.4105
R4113 VDDA.n3093 VDDA.n2940 3.4105
R4114 VDDA.n3090 VDDA.n2940 3.4105
R4115 VDDA.n3095 VDDA.n2940 3.4105
R4116 VDDA.n3089 VDDA.n2940 3.4105
R4117 VDDA.n3097 VDDA.n2940 3.4105
R4118 VDDA.n3088 VDDA.n2940 3.4105
R4119 VDDA.n3099 VDDA.n2940 3.4105
R4120 VDDA.n3087 VDDA.n2940 3.4105
R4121 VDDA.n3101 VDDA.n2940 3.4105
R4122 VDDA.n3086 VDDA.n2940 3.4105
R4123 VDDA.n3103 VDDA.n2940 3.4105
R4124 VDDA.n3085 VDDA.n2940 3.4105
R4125 VDDA.n3105 VDDA.n2940 3.4105
R4126 VDDA.n3084 VDDA.n2940 3.4105
R4127 VDDA.n3107 VDDA.n2940 3.4105
R4128 VDDA.n3083 VDDA.n2940 3.4105
R4129 VDDA.n3109 VDDA.n2940 3.4105
R4130 VDDA.n3082 VDDA.n2940 3.4105
R4131 VDDA.n3111 VDDA.n2940 3.4105
R4132 VDDA.n3081 VDDA.n2940 3.4105
R4133 VDDA.n3113 VDDA.n2940 3.4105
R4134 VDDA.n3080 VDDA.n2940 3.4105
R4135 VDDA.n3115 VDDA.n2940 3.4105
R4136 VDDA.n3079 VDDA.n2940 3.4105
R4137 VDDA.n3117 VDDA.n2940 3.4105
R4138 VDDA.n3078 VDDA.n2940 3.4105
R4139 VDDA.n3119 VDDA.n2940 3.4105
R4140 VDDA.n3077 VDDA.n2940 3.4105
R4141 VDDA.n3121 VDDA.n2940 3.4105
R4142 VDDA.n3076 VDDA.n2940 3.4105
R4143 VDDA.n2940 VDDA.n18 3.4105
R4144 VDDA.n3123 VDDA.n2940 3.4105
R4145 VDDA.n3070 VDDA.n16 3.4105
R4146 VDDA.n3093 VDDA.n3070 3.4105
R4147 VDDA.n3090 VDDA.n3070 3.4105
R4148 VDDA.n3095 VDDA.n3070 3.4105
R4149 VDDA.n3089 VDDA.n3070 3.4105
R4150 VDDA.n3097 VDDA.n3070 3.4105
R4151 VDDA.n3088 VDDA.n3070 3.4105
R4152 VDDA.n3099 VDDA.n3070 3.4105
R4153 VDDA.n3087 VDDA.n3070 3.4105
R4154 VDDA.n3101 VDDA.n3070 3.4105
R4155 VDDA.n3086 VDDA.n3070 3.4105
R4156 VDDA.n3103 VDDA.n3070 3.4105
R4157 VDDA.n3085 VDDA.n3070 3.4105
R4158 VDDA.n3105 VDDA.n3070 3.4105
R4159 VDDA.n3084 VDDA.n3070 3.4105
R4160 VDDA.n3107 VDDA.n3070 3.4105
R4161 VDDA.n3083 VDDA.n3070 3.4105
R4162 VDDA.n3109 VDDA.n3070 3.4105
R4163 VDDA.n3082 VDDA.n3070 3.4105
R4164 VDDA.n3111 VDDA.n3070 3.4105
R4165 VDDA.n3081 VDDA.n3070 3.4105
R4166 VDDA.n3113 VDDA.n3070 3.4105
R4167 VDDA.n3080 VDDA.n3070 3.4105
R4168 VDDA.n3115 VDDA.n3070 3.4105
R4169 VDDA.n3079 VDDA.n3070 3.4105
R4170 VDDA.n3117 VDDA.n3070 3.4105
R4171 VDDA.n3078 VDDA.n3070 3.4105
R4172 VDDA.n3119 VDDA.n3070 3.4105
R4173 VDDA.n3077 VDDA.n3070 3.4105
R4174 VDDA.n3121 VDDA.n3070 3.4105
R4175 VDDA.n3076 VDDA.n3070 3.4105
R4176 VDDA.n3070 VDDA.n18 3.4105
R4177 VDDA.n3123 VDDA.n3070 3.4105
R4178 VDDA.n2939 VDDA.n16 3.4105
R4179 VDDA.n3093 VDDA.n2939 3.4105
R4180 VDDA.n3090 VDDA.n2939 3.4105
R4181 VDDA.n3095 VDDA.n2939 3.4105
R4182 VDDA.n3089 VDDA.n2939 3.4105
R4183 VDDA.n3097 VDDA.n2939 3.4105
R4184 VDDA.n3088 VDDA.n2939 3.4105
R4185 VDDA.n3099 VDDA.n2939 3.4105
R4186 VDDA.n3087 VDDA.n2939 3.4105
R4187 VDDA.n3101 VDDA.n2939 3.4105
R4188 VDDA.n3086 VDDA.n2939 3.4105
R4189 VDDA.n3103 VDDA.n2939 3.4105
R4190 VDDA.n3085 VDDA.n2939 3.4105
R4191 VDDA.n3105 VDDA.n2939 3.4105
R4192 VDDA.n3084 VDDA.n2939 3.4105
R4193 VDDA.n3107 VDDA.n2939 3.4105
R4194 VDDA.n3083 VDDA.n2939 3.4105
R4195 VDDA.n3109 VDDA.n2939 3.4105
R4196 VDDA.n3082 VDDA.n2939 3.4105
R4197 VDDA.n3111 VDDA.n2939 3.4105
R4198 VDDA.n3081 VDDA.n2939 3.4105
R4199 VDDA.n3113 VDDA.n2939 3.4105
R4200 VDDA.n3080 VDDA.n2939 3.4105
R4201 VDDA.n3115 VDDA.n2939 3.4105
R4202 VDDA.n3079 VDDA.n2939 3.4105
R4203 VDDA.n3117 VDDA.n2939 3.4105
R4204 VDDA.n3078 VDDA.n2939 3.4105
R4205 VDDA.n3119 VDDA.n2939 3.4105
R4206 VDDA.n3077 VDDA.n2939 3.4105
R4207 VDDA.n3121 VDDA.n2939 3.4105
R4208 VDDA.n3076 VDDA.n2939 3.4105
R4209 VDDA.n2939 VDDA.n18 3.4105
R4210 VDDA.n3123 VDDA.n2939 3.4105
R4211 VDDA.n3073 VDDA.n16 3.4105
R4212 VDDA.n3093 VDDA.n3073 3.4105
R4213 VDDA.n3090 VDDA.n3073 3.4105
R4214 VDDA.n3095 VDDA.n3073 3.4105
R4215 VDDA.n3089 VDDA.n3073 3.4105
R4216 VDDA.n3097 VDDA.n3073 3.4105
R4217 VDDA.n3088 VDDA.n3073 3.4105
R4218 VDDA.n3099 VDDA.n3073 3.4105
R4219 VDDA.n3087 VDDA.n3073 3.4105
R4220 VDDA.n3101 VDDA.n3073 3.4105
R4221 VDDA.n3086 VDDA.n3073 3.4105
R4222 VDDA.n3103 VDDA.n3073 3.4105
R4223 VDDA.n3085 VDDA.n3073 3.4105
R4224 VDDA.n3105 VDDA.n3073 3.4105
R4225 VDDA.n3084 VDDA.n3073 3.4105
R4226 VDDA.n3107 VDDA.n3073 3.4105
R4227 VDDA.n3083 VDDA.n3073 3.4105
R4228 VDDA.n3109 VDDA.n3073 3.4105
R4229 VDDA.n3082 VDDA.n3073 3.4105
R4230 VDDA.n3111 VDDA.n3073 3.4105
R4231 VDDA.n3081 VDDA.n3073 3.4105
R4232 VDDA.n3113 VDDA.n3073 3.4105
R4233 VDDA.n3080 VDDA.n3073 3.4105
R4234 VDDA.n3115 VDDA.n3073 3.4105
R4235 VDDA.n3079 VDDA.n3073 3.4105
R4236 VDDA.n3117 VDDA.n3073 3.4105
R4237 VDDA.n3078 VDDA.n3073 3.4105
R4238 VDDA.n3119 VDDA.n3073 3.4105
R4239 VDDA.n3077 VDDA.n3073 3.4105
R4240 VDDA.n3121 VDDA.n3073 3.4105
R4241 VDDA.n3076 VDDA.n3073 3.4105
R4242 VDDA.n3073 VDDA.n18 3.4105
R4243 VDDA.n3123 VDDA.n3073 3.4105
R4244 VDDA.n2938 VDDA.n16 3.4105
R4245 VDDA.n3093 VDDA.n2938 3.4105
R4246 VDDA.n3090 VDDA.n2938 3.4105
R4247 VDDA.n3095 VDDA.n2938 3.4105
R4248 VDDA.n3089 VDDA.n2938 3.4105
R4249 VDDA.n3097 VDDA.n2938 3.4105
R4250 VDDA.n3088 VDDA.n2938 3.4105
R4251 VDDA.n3099 VDDA.n2938 3.4105
R4252 VDDA.n3087 VDDA.n2938 3.4105
R4253 VDDA.n3101 VDDA.n2938 3.4105
R4254 VDDA.n3086 VDDA.n2938 3.4105
R4255 VDDA.n3103 VDDA.n2938 3.4105
R4256 VDDA.n3085 VDDA.n2938 3.4105
R4257 VDDA.n3105 VDDA.n2938 3.4105
R4258 VDDA.n3084 VDDA.n2938 3.4105
R4259 VDDA.n3107 VDDA.n2938 3.4105
R4260 VDDA.n3083 VDDA.n2938 3.4105
R4261 VDDA.n3109 VDDA.n2938 3.4105
R4262 VDDA.n3082 VDDA.n2938 3.4105
R4263 VDDA.n3111 VDDA.n2938 3.4105
R4264 VDDA.n3081 VDDA.n2938 3.4105
R4265 VDDA.n3113 VDDA.n2938 3.4105
R4266 VDDA.n3080 VDDA.n2938 3.4105
R4267 VDDA.n3115 VDDA.n2938 3.4105
R4268 VDDA.n3079 VDDA.n2938 3.4105
R4269 VDDA.n3117 VDDA.n2938 3.4105
R4270 VDDA.n3078 VDDA.n2938 3.4105
R4271 VDDA.n3119 VDDA.n2938 3.4105
R4272 VDDA.n3077 VDDA.n2938 3.4105
R4273 VDDA.n3121 VDDA.n2938 3.4105
R4274 VDDA.n3076 VDDA.n2938 3.4105
R4275 VDDA.n2938 VDDA.n18 3.4105
R4276 VDDA.n3123 VDDA.n2938 3.4105
R4277 VDDA.n3122 VDDA.n3093 3.4105
R4278 VDDA.n3122 VDDA.n3090 3.4105
R4279 VDDA.n3122 VDDA.n3095 3.4105
R4280 VDDA.n3122 VDDA.n3089 3.4105
R4281 VDDA.n3122 VDDA.n3097 3.4105
R4282 VDDA.n3122 VDDA.n3088 3.4105
R4283 VDDA.n3122 VDDA.n3099 3.4105
R4284 VDDA.n3122 VDDA.n3087 3.4105
R4285 VDDA.n3122 VDDA.n3101 3.4105
R4286 VDDA.n3122 VDDA.n3086 3.4105
R4287 VDDA.n3122 VDDA.n3103 3.4105
R4288 VDDA.n3122 VDDA.n3085 3.4105
R4289 VDDA.n3122 VDDA.n3105 3.4105
R4290 VDDA.n3122 VDDA.n3084 3.4105
R4291 VDDA.n3122 VDDA.n3107 3.4105
R4292 VDDA.n3122 VDDA.n3083 3.4105
R4293 VDDA.n3122 VDDA.n3109 3.4105
R4294 VDDA.n3122 VDDA.n3082 3.4105
R4295 VDDA.n3122 VDDA.n3111 3.4105
R4296 VDDA.n3122 VDDA.n3081 3.4105
R4297 VDDA.n3122 VDDA.n3113 3.4105
R4298 VDDA.n3122 VDDA.n3080 3.4105
R4299 VDDA.n3122 VDDA.n3115 3.4105
R4300 VDDA.n3122 VDDA.n3079 3.4105
R4301 VDDA.n3122 VDDA.n3117 3.4105
R4302 VDDA.n3122 VDDA.n3078 3.4105
R4303 VDDA.n3122 VDDA.n3119 3.4105
R4304 VDDA.n3122 VDDA.n3077 3.4105
R4305 VDDA.n3122 VDDA.n3121 3.4105
R4306 VDDA.n3122 VDDA.n3076 3.4105
R4307 VDDA.n3122 VDDA.n18 3.4105
R4308 VDDA.n3123 VDDA.n3122 3.4105
R4309 VDDA.n2141 VDDA.n2140 3.11118
R4310 VDDA.n2151 VDDA.n2150 3.11118
R4311 VDDA.n2140 VDDA.n2122 3.04304
R4312 VDDA.n2150 VDDA.n2102 3.04304
R4313 VDDA.n593 VDDA.n589 2.96402
R4314 VDDA.n2546 VDDA.n2542 2.96402
R4315 VDDA.n2472 VDDA.n2471 2.8255
R4316 VDDA.n2474 VDDA.n2473 2.8255
R4317 VDDA.n592 VDDA.n591 2.423
R4318 VDDA.n590 VDDA.n589 2.423
R4319 VDDA.n2543 VDDA.n2542 2.423
R4320 VDDA.n2545 VDDA.n2544 2.423
R4321 VDDA.n2054 VDDA.n2053 2.41009
R4322 VDDA.n2512 VDDA.n2510 2.3971
R4323 VDDA.n2443 VDDA.n561 2.39632
R4324 VDDA.n1939 VDDA.n1938 2.36299
R4325 VDDA.n93 VDDA.n92 2.30736
R4326 VDDA.n2806 VDDA.n2803 2.30736
R4327 VDDA.n2656 VDDA.n2655 2.30736
R4328 VDDA.n271 VDDA.n270 2.30736
R4329 VDDA.n412 VDDA.n409 2.30736
R4330 VDDA.n1376 VDDA.n1375 2.30736
R4331 VDDA.n686 VDDA.n685 2.30736
R4332 VDDA.n1178 VDDA.n1175 2.30736
R4333 VDDA.n1028 VDDA.n1027 2.30736
R4334 VDDA.n1726 VDDA.n1725 2.30736
R4335 VDDA.n2403 VDDA.n2402 2.30736
R4336 VDDA.n840 VDDA.n839 2.30736
R4337 VDDA.n1914 VDDA.n1552 2.2948
R4338 VDDA.n1915 VDDA.n1914 2.2948
R4339 VDDA.n593 VDDA.n592 2.27652
R4340 VDDA.n2546 VDDA.n2545 2.27652
R4341 VDDA.n2096 VDDA.n2088 2.26187
R4342 VDDA.n2162 VDDA.n2086 2.26187
R4343 VDDA.n2239 VDDA.n2084 2.26187
R4344 VDDA.n2289 VDDA.n2082 2.26187
R4345 VDDA.n2463 VDDA.n2454 2.26187
R4346 VDDA.n2465 VDDA.n2463 2.26187
R4347 VDDA.n2577 VDDA.n2576 2.26187
R4348 VDDA.n2552 VDDA.n2551 2.26187
R4349 VDDA.n2539 VDDA.n2517 2.26187
R4350 VDDA.n2523 VDDA.n2520 2.26187
R4351 VDDA.n2524 VDDA.n2523 2.26187
R4352 VDDA.n2442 VDDA.n2441 2.26187
R4353 VDDA.n586 VDDA.n585 2.26187
R4354 VDDA.n2417 VDDA.n2416 2.26187
R4355 VDDA.n2416 VDDA.n602 2.26187
R4356 VDDA.n954 VDDA.n951 2.26187
R4357 VDDA.n954 VDDA.n953 2.26187
R4358 VDDA.n2093 VDDA.n2088 2.26187
R4359 VDDA.n587 VDDA.n586 2.26187
R4360 VDDA.n598 VDDA.n597 2.26187
R4361 VDDA.n2481 VDDA.n2480 2.26187
R4362 VDDA.n1913 VDDA.n1553 2.2505
R4363 VDDA.n1912 VDDA.n1911 2.2505
R4364 VDDA.n1555 VDDA.n1554 2.2505
R4365 VDDA.n1733 VDDA.n1730 2.2505
R4366 VDDA.n1903 VDDA.n1902 2.2505
R4367 VDDA.n1901 VDDA.n1732 2.2505
R4368 VDDA.n1900 VDDA.n1899 2.2505
R4369 VDDA.n1735 VDDA.n1734 2.2505
R4370 VDDA.n1893 VDDA.n1892 2.2505
R4371 VDDA.n1891 VDDA.n1739 2.2505
R4372 VDDA.n1890 VDDA.n1889 2.2505
R4373 VDDA.n1741 VDDA.n1740 2.2505
R4374 VDDA.n1883 VDDA.n1882 2.2505
R4375 VDDA.n1881 VDDA.n1745 2.2505
R4376 VDDA.n1880 VDDA.n1879 2.2505
R4377 VDDA.n1747 VDDA.n1746 2.2505
R4378 VDDA.n1873 VDDA.n1872 2.2505
R4379 VDDA.n1871 VDDA.n1751 2.2505
R4380 VDDA.n1870 VDDA.n1869 2.2505
R4381 VDDA.n1753 VDDA.n1752 2.2505
R4382 VDDA.n1863 VDDA.n1862 2.2505
R4383 VDDA.n1861 VDDA.n1757 2.2505
R4384 VDDA.n1860 VDDA.n1859 2.2505
R4385 VDDA.n1759 VDDA.n1758 2.2505
R4386 VDDA.n1853 VDDA.n1852 2.2505
R4387 VDDA.n1851 VDDA.n1763 2.2505
R4388 VDDA.n1850 VDDA.n1849 2.2505
R4389 VDDA.n1765 VDDA.n1764 2.2505
R4390 VDDA.n1843 VDDA.n1842 2.2505
R4391 VDDA.n1841 VDDA.n1769 2.2505
R4392 VDDA.n1840 VDDA.n1839 2.2505
R4393 VDDA.n1771 VDDA.n1770 2.2505
R4394 VDDA.n1833 VDDA.n1832 2.2505
R4395 VDDA.n1831 VDDA.n1775 2.2505
R4396 VDDA.n1830 VDDA.n1829 2.2505
R4397 VDDA.n1777 VDDA.n1776 2.2505
R4398 VDDA.n1823 VDDA.n1822 2.2505
R4399 VDDA.n1821 VDDA.n1781 2.2505
R4400 VDDA.n1820 VDDA.n1819 2.2505
R4401 VDDA.n1783 VDDA.n1782 2.2505
R4402 VDDA.n1813 VDDA.n1812 2.2505
R4403 VDDA.n1811 VDDA.n1787 2.2505
R4404 VDDA.n1810 VDDA.n1809 2.2505
R4405 VDDA.n1789 VDDA.n1788 2.2505
R4406 VDDA.n1803 VDDA.n1802 2.2505
R4407 VDDA.n1801 VDDA.n1793 2.2505
R4408 VDDA.n2097 VDDA.n2087 2.24063
R4409 VDDA.n2163 VDDA.n2085 2.24063
R4410 VDDA.n2240 VDDA.n2083 2.24063
R4411 VDDA.n2290 VDDA.n2081 2.24063
R4412 VDDA.n2482 VDDA.n2481 2.24063
R4413 VDDA.n2476 VDDA.n2452 2.24063
R4414 VDDA.n2478 VDDA.n2477 2.24063
R4415 VDDA.n2468 VDDA.n2467 2.24063
R4416 VDDA.n2584 VDDA.n192 2.24063
R4417 VDDA.n362 VDDA.n361 2.24063
R4418 VDDA.n2757 VDDA.n190 2.24063
R4419 VDDA.n191 VDDA.n189 2.24063
R4420 VDDA.n2928 VDDA.n187 2.24063
R4421 VDDA.n188 VDDA.n186 2.24063
R4422 VDDA.n2932 VDDA.n2931 2.24063
R4423 VDDA.n185 VDDA.n184 2.24063
R4424 VDDA.n2575 VDDA.n363 2.24063
R4425 VDDA.n2573 VDDA.n2572 2.24063
R4426 VDDA.n534 VDDA.n533 2.24063
R4427 VDDA.n2550 VDDA.n537 2.24063
R4428 VDDA.n2541 VDDA.n2540 2.24063
R4429 VDDA.n2511 VDDA.n540 2.24063
R4430 VDDA.n2495 VDDA.n539 2.24063
R4431 VDDA.n2485 VDDA.n2484 2.24063
R4432 VDDA.n2451 VDDA.n544 2.24063
R4433 VDDA.n2440 VDDA.n545 2.24063
R4434 VDDA.n595 VDDA.n594 2.24063
R4435 VDDA.n597 VDDA.n596 2.24063
R4436 VDDA.n585 VDDA.n584 2.24063
R4437 VDDA.n2438 VDDA.n2437 2.24063
R4438 VDDA.n566 VDDA.n565 2.24063
R4439 VDDA.n1129 VDDA.n782 2.24063
R4440 VDDA.n783 VDDA.n781 2.24063
R4441 VDDA.n1300 VDDA.n779 2.24063
R4442 VDDA.n780 VDDA.n778 2.24063
R4443 VDDA.n1304 VDDA.n606 2.24063
R4444 VDDA.n777 VDDA.n776 2.24063
R4445 VDDA.n2410 VDDA.n605 2.24063
R4446 VDDA.n608 VDDA.n604 2.24063
R4447 VDDA.n2093 VDDA.n2092 2.24063
R4448 VDDA.n2098 VDDA.n2086 2.24063
R4449 VDDA.n2159 VDDA.n2158 2.24063
R4450 VDDA.n2164 VDDA.n2084 2.24063
R4451 VDDA.n2236 VDDA.n2235 2.24063
R4452 VDDA.n2241 VDDA.n2082 2.24063
R4453 VDDA.n2286 VDDA.n2285 2.24063
R4454 VDDA.n2466 VDDA.n2465 2.24063
R4455 VDDA.n2585 VDDA.n360 2.24063
R4456 VDDA.n2754 VDDA.n2753 2.24063
R4457 VDDA.n2925 VDDA.n2924 2.24063
R4458 VDDA.n2933 VDDA.n182 2.24063
R4459 VDDA.n2578 VDDA.n2577 2.24063
R4460 VDDA.n2580 VDDA.n2579 2.24063
R4461 VDDA.n2574 VDDA.n531 2.24063
R4462 VDDA.n2553 VDDA.n2552 2.24063
R4463 VDDA.n2555 VDDA.n2554 2.24063
R4464 VDDA.n2549 VDDA.n2517 2.24063
R4465 VDDA.n2548 VDDA.n2547 2.24063
R4466 VDDA.n2538 VDDA.n2520 2.24063
R4467 VDDA.n2537 VDDA.n2536 2.24063
R4468 VDDA.n2513 VDDA.n2512 2.24063
R4469 VDDA.n2443 VDDA.n2442 2.24063
R4470 VDDA.n2445 VDDA.n2444 2.24063
R4471 VDDA.n599 VDDA.n567 2.24063
R4472 VDDA.n588 VDDA.n570 2.24063
R4473 VDDA.n2439 VDDA.n563 2.24063
R4474 VDDA.n2418 VDDA.n2417 2.24063
R4475 VDDA.n2420 VDDA.n2419 2.24063
R4476 VDDA.n1126 VDDA.n1125 2.24063
R4477 VDDA.n1297 VDDA.n1296 2.24063
R4478 VDDA.n1305 VDDA.n775 2.24063
R4479 VDDA.n2412 VDDA.n2411 2.24063
R4480 VDDA.n957 VDDA.n951 2.24063
R4481 VDDA.n956 VDDA.n784 2.24063
R4482 VDDA.n2568 VDDA.n2567 1.97758
R4483 VDDA.n2566 VDDA.n2565 1.97758
R4484 VDDA.n2433 VDDA.n2432 1.97758
R4485 VDDA.n2431 VDDA.n2430 1.97758
R4486 VDDA.n2139 VDDA.n2138 1.90331
R4487 VDDA.n2461 VDDA.n2460 1.888
R4488 VDDA.n2459 VDDA.n2458 1.888
R4489 VDDA.n2507 VDDA.n2506 1.888
R4490 VDDA.n2509 VDDA.n2508 1.888
R4491 VDDA.n560 VDDA.n559 1.888
R4492 VDDA.n558 VDDA.n557 1.888
R4493 VDDA.n2569 VDDA.n2568 1.88069
R4494 VDDA.n2565 VDDA.n2564 1.88069
R4495 VDDA.n2434 VDDA.n2433 1.88069
R4496 VDDA.n2430 VDDA.n2429 1.88069
R4497 VDDA.n2934 VDDA.n2933 1.79738
R4498 VDDA.n2924 VDDA.n2923 1.79738
R4499 VDDA.n2753 VDDA.n2752 1.79738
R4500 VDDA.n2586 VDDA.n2585 1.79738
R4501 VDDA.n2578 VDDA.n529 1.79738
R4502 VDDA.n2411 VDDA.n2409 1.79738
R4503 VDDA.n1306 VDDA.n1305 1.79738
R4504 VDDA.n1296 VDDA.n1295 1.79738
R4505 VDDA.n1125 VDDA.n1124 1.79738
R4506 VDDA.n958 VDDA.n957 1.79738
R4507 VDDA.n2147 VDDA.n2146 1.77831
R4508 VDDA.n2149 VDDA.n2148 1.77831
R4509 VDDA.n2157 VDDA.n2156 1.77831
R4510 VDDA.n2291 VDDA.n1469 1.7622
R4511 VDDA.n1800 VDDA.n1794 1.74133
R4512 VDDA.n3124 VDDA.n15 1.70583
R4513 VDDA.n3124 VDDA.n14 1.70583
R4514 VDDA.n3124 VDDA.n13 1.70583
R4515 VDDA.n3124 VDDA.n12 1.70583
R4516 VDDA.n3124 VDDA.n11 1.70583
R4517 VDDA.n3124 VDDA.n10 1.70583
R4518 VDDA.n3124 VDDA.n9 1.70583
R4519 VDDA.n3124 VDDA.n8 1.70583
R4520 VDDA.n3124 VDDA.n7 1.70583
R4521 VDDA.n3124 VDDA.n6 1.70583
R4522 VDDA.n3124 VDDA.n5 1.70583
R4523 VDDA.n3124 VDDA.n4 1.70583
R4524 VDDA.n3124 VDDA.n3 1.70583
R4525 VDDA.n3124 VDDA.n2 1.70583
R4526 VDDA.n3124 VDDA.n1 1.70583
R4527 VDDA.n3092 VDDA.n2974 1.70583
R4528 VDDA.n3094 VDDA.n2974 1.70583
R4529 VDDA.n3096 VDDA.n2974 1.70583
R4530 VDDA.n3098 VDDA.n2974 1.70583
R4531 VDDA.n3100 VDDA.n2974 1.70583
R4532 VDDA.n3102 VDDA.n2974 1.70583
R4533 VDDA.n3104 VDDA.n2974 1.70583
R4534 VDDA.n3106 VDDA.n2974 1.70583
R4535 VDDA.n3108 VDDA.n2974 1.70583
R4536 VDDA.n3110 VDDA.n2974 1.70583
R4537 VDDA.n3112 VDDA.n2974 1.70583
R4538 VDDA.n3114 VDDA.n2974 1.70583
R4539 VDDA.n3116 VDDA.n2974 1.70583
R4540 VDDA.n3118 VDDA.n2974 1.70583
R4541 VDDA.n3120 VDDA.n2974 1.70583
R4542 VDDA.n3075 VDDA.n2974 1.70583
R4543 VDDA.n3122 VDDA.n3091 1.70583
R4544 VDDA.n2972 VDDA.n0 1.70567
R4545 VDDA.n2973 VDDA.n17 1.70567
R4546 VDDA.n2975 VDDA.n2972 1.70567
R4547 VDDA.n2976 VDDA.n17 1.70567
R4548 VDDA.n2978 VDDA.n2972 1.70567
R4549 VDDA.n2979 VDDA.n17 1.70567
R4550 VDDA.n2981 VDDA.n2972 1.70567
R4551 VDDA.n2982 VDDA.n17 1.70567
R4552 VDDA.n2984 VDDA.n2972 1.70567
R4553 VDDA.n2985 VDDA.n17 1.70567
R4554 VDDA.n2987 VDDA.n2972 1.70567
R4555 VDDA.n2988 VDDA.n17 1.70567
R4556 VDDA.n2990 VDDA.n2972 1.70567
R4557 VDDA.n2991 VDDA.n17 1.70567
R4558 VDDA.n2993 VDDA.n2972 1.70567
R4559 VDDA.n2994 VDDA.n17 1.70567
R4560 VDDA.n2996 VDDA.n2972 1.70567
R4561 VDDA.n2997 VDDA.n17 1.70567
R4562 VDDA.n2999 VDDA.n2972 1.70567
R4563 VDDA.n3000 VDDA.n17 1.70567
R4564 VDDA.n3002 VDDA.n2972 1.70567
R4565 VDDA.n3003 VDDA.n17 1.70567
R4566 VDDA.n3005 VDDA.n2972 1.70567
R4567 VDDA.n3006 VDDA.n17 1.70567
R4568 VDDA.n3008 VDDA.n2972 1.70567
R4569 VDDA.n3009 VDDA.n17 1.70567
R4570 VDDA.n3011 VDDA.n2972 1.70567
R4571 VDDA.n3012 VDDA.n17 1.70567
R4572 VDDA.n3014 VDDA.n2972 1.70567
R4573 VDDA.n3015 VDDA.n17 1.70567
R4574 VDDA.n3017 VDDA.n2972 1.70567
R4575 VDDA.n3018 VDDA.n17 1.70567
R4576 VDDA.n3020 VDDA.n2972 1.70567
R4577 VDDA.n3021 VDDA.n17 1.70567
R4578 VDDA.n3024 VDDA.n17 1.70567
R4579 VDDA.n3026 VDDA.n2972 1.70567
R4580 VDDA.n3027 VDDA.n17 1.70567
R4581 VDDA.n3029 VDDA.n2972 1.70567
R4582 VDDA.n3030 VDDA.n17 1.70567
R4583 VDDA.n3032 VDDA.n2972 1.70567
R4584 VDDA.n3033 VDDA.n17 1.70567
R4585 VDDA.n3035 VDDA.n2972 1.70567
R4586 VDDA.n3036 VDDA.n17 1.70567
R4587 VDDA.n3038 VDDA.n2972 1.70567
R4588 VDDA.n3039 VDDA.n17 1.70567
R4589 VDDA.n3041 VDDA.n2972 1.70567
R4590 VDDA.n3042 VDDA.n17 1.70567
R4591 VDDA.n3044 VDDA.n2972 1.70567
R4592 VDDA.n3045 VDDA.n17 1.70567
R4593 VDDA.n3047 VDDA.n2972 1.70567
R4594 VDDA.n3048 VDDA.n17 1.70567
R4595 VDDA.n3050 VDDA.n2972 1.70567
R4596 VDDA.n3051 VDDA.n17 1.70567
R4597 VDDA.n3053 VDDA.n2972 1.70567
R4598 VDDA.n3054 VDDA.n17 1.70567
R4599 VDDA.n3056 VDDA.n2972 1.70567
R4600 VDDA.n3057 VDDA.n17 1.70567
R4601 VDDA.n3059 VDDA.n2972 1.70567
R4602 VDDA.n3060 VDDA.n17 1.70567
R4603 VDDA.n3062 VDDA.n2972 1.70567
R4604 VDDA.n3063 VDDA.n17 1.70567
R4605 VDDA.n3065 VDDA.n2972 1.70567
R4606 VDDA.n3066 VDDA.n17 1.70567
R4607 VDDA.n3068 VDDA.n2972 1.70567
R4608 VDDA.n3069 VDDA.n17 1.70567
R4609 VDDA.n3071 VDDA.n2972 1.70567
R4610 VDDA.n3072 VDDA.n17 1.70567
R4611 VDDA.n3074 VDDA.n2972 1.70567
R4612 VDDA.n1799 VDDA.n1798 1.7055
R4613 VDDA.n1795 VDDA.n1793 1.7055
R4614 VDDA.n1804 VDDA.n1803 1.7055
R4615 VDDA.n1806 VDDA.n1789 1.7055
R4616 VDDA.n1809 VDDA.n1808 1.7055
R4617 VDDA.n1790 VDDA.n1787 1.7055
R4618 VDDA.n1814 VDDA.n1813 1.7055
R4619 VDDA.n1816 VDDA.n1783 1.7055
R4620 VDDA.n1819 VDDA.n1818 1.7055
R4621 VDDA.n1784 VDDA.n1781 1.7055
R4622 VDDA.n1824 VDDA.n1823 1.7055
R4623 VDDA.n1826 VDDA.n1777 1.7055
R4624 VDDA.n1829 VDDA.n1828 1.7055
R4625 VDDA.n1778 VDDA.n1775 1.7055
R4626 VDDA.n1834 VDDA.n1833 1.7055
R4627 VDDA.n1836 VDDA.n1771 1.7055
R4628 VDDA.n1839 VDDA.n1838 1.7055
R4629 VDDA.n1772 VDDA.n1769 1.7055
R4630 VDDA.n1844 VDDA.n1843 1.7055
R4631 VDDA.n1846 VDDA.n1765 1.7055
R4632 VDDA.n1849 VDDA.n1848 1.7055
R4633 VDDA.n1766 VDDA.n1763 1.7055
R4634 VDDA.n1854 VDDA.n1853 1.7055
R4635 VDDA.n1856 VDDA.n1759 1.7055
R4636 VDDA.n1859 VDDA.n1858 1.7055
R4637 VDDA.n1760 VDDA.n1757 1.7055
R4638 VDDA.n1864 VDDA.n1863 1.7055
R4639 VDDA.n1866 VDDA.n1753 1.7055
R4640 VDDA.n1869 VDDA.n1868 1.7055
R4641 VDDA.n1754 VDDA.n1751 1.7055
R4642 VDDA.n1874 VDDA.n1873 1.7055
R4643 VDDA.n1876 VDDA.n1747 1.7055
R4644 VDDA.n1879 VDDA.n1878 1.7055
R4645 VDDA.n1748 VDDA.n1745 1.7055
R4646 VDDA.n1884 VDDA.n1883 1.7055
R4647 VDDA.n1886 VDDA.n1741 1.7055
R4648 VDDA.n1889 VDDA.n1888 1.7055
R4649 VDDA.n1742 VDDA.n1739 1.7055
R4650 VDDA.n1894 VDDA.n1893 1.7055
R4651 VDDA.n1896 VDDA.n1735 1.7055
R4652 VDDA.n1899 VDDA.n1898 1.7055
R4653 VDDA.n1736 VDDA.n1732 1.7055
R4654 VDDA.n1904 VDDA.n1903 1.7055
R4655 VDDA.n1906 VDDA.n1730 1.7055
R4656 VDDA.n1908 VDDA.n1555 1.7055
R4657 VDDA.n1911 VDDA.n1910 1.7055
R4658 VDDA.n1557 VDDA.n1553 1.7055
R4659 VDDA.n3023 VDDA.n2972 1.70549
R4660 VDDA.n1791 VDDA.n1729 1.69989
R4661 VDDA.n1825 VDDA.n1729 1.69989
R4662 VDDA.n1773 VDDA.n1729 1.69989
R4663 VDDA.n1855 VDDA.n1729 1.69989
R4664 VDDA.n1755 VDDA.n1729 1.69989
R4665 VDDA.n1885 VDDA.n1729 1.69989
R4666 VDDA.n1737 VDDA.n1729 1.69989
R4667 VDDA.n1807 VDDA.n1516 1.69938
R4668 VDDA.n1786 VDDA.n1516 1.69938
R4669 VDDA.n1780 VDDA.n1516 1.69938
R4670 VDDA.n1827 VDDA.n1516 1.69938
R4671 VDDA.n1837 VDDA.n1516 1.69938
R4672 VDDA.n1768 VDDA.n1516 1.69938
R4673 VDDA.n1762 VDDA.n1516 1.69938
R4674 VDDA.n1857 VDDA.n1516 1.69938
R4675 VDDA.n1867 VDDA.n1516 1.69938
R4676 VDDA.n1750 VDDA.n1516 1.69938
R4677 VDDA.n1744 VDDA.n1516 1.69938
R4678 VDDA.n1887 VDDA.n1516 1.69938
R4679 VDDA.n1897 VDDA.n1516 1.69938
R4680 VDDA.n1731 VDDA.n1516 1.69938
R4681 VDDA.n1556 VDDA.n1516 1.69938
R4682 VDDA.n1797 VDDA.n1516 1.69938
R4683 VDDA.n1796 VDDA.n1729 1.69888
R4684 VDDA.n1792 VDDA.n1516 1.69888
R4685 VDDA.n1805 VDDA.n1729 1.69888
R4686 VDDA.n1815 VDDA.n1729 1.69888
R4687 VDDA.n1817 VDDA.n1516 1.69888
R4688 VDDA.n1785 VDDA.n1729 1.69888
R4689 VDDA.n1779 VDDA.n1729 1.69888
R4690 VDDA.n1774 VDDA.n1516 1.69888
R4691 VDDA.n1835 VDDA.n1729 1.69888
R4692 VDDA.n1845 VDDA.n1729 1.69888
R4693 VDDA.n1847 VDDA.n1516 1.69888
R4694 VDDA.n1767 VDDA.n1729 1.69888
R4695 VDDA.n1761 VDDA.n1729 1.69888
R4696 VDDA.n1756 VDDA.n1516 1.69888
R4697 VDDA.n1865 VDDA.n1729 1.69888
R4698 VDDA.n1875 VDDA.n1729 1.69888
R4699 VDDA.n1877 VDDA.n1516 1.69888
R4700 VDDA.n1749 VDDA.n1729 1.69888
R4701 VDDA.n1743 VDDA.n1729 1.69888
R4702 VDDA.n1738 VDDA.n1516 1.69888
R4703 VDDA.n1895 VDDA.n1729 1.69888
R4704 VDDA.n1905 VDDA.n1729 1.69888
R4705 VDDA.n1907 VDDA.n1516 1.69888
R4706 VDDA.n1909 VDDA.n1729 1.69888
R4707 VDDA.n961 VDDA.n810 1.69433
R4708 VDDA.n961 VDDA.n807 1.69433
R4709 VDDA.n961 VDDA.n804 1.69433
R4710 VDDA.n961 VDDA.n801 1.69433
R4711 VDDA.n961 VDDA.n798 1.69433
R4712 VDDA.n961 VDDA.n795 1.69433
R4713 VDDA.n961 VDDA.n792 1.69433
R4714 VDDA.n1121 VDDA.n983 1.69433
R4715 VDDA.n1121 VDDA.n980 1.69433
R4716 VDDA.n1121 VDDA.n977 1.69433
R4717 VDDA.n1121 VDDA.n974 1.69433
R4718 VDDA.n1121 VDDA.n971 1.69433
R4719 VDDA.n1121 VDDA.n968 1.69433
R4720 VDDA.n1121 VDDA.n965 1.69433
R4721 VDDA.n1281 VDDA.n612 1.69433
R4722 VDDA.n1263 VDDA.n612 1.69433
R4723 VDDA.n1251 VDDA.n612 1.69433
R4724 VDDA.n1233 VDDA.n612 1.69433
R4725 VDDA.n1221 VDDA.n612 1.69433
R4726 VDDA.n1203 VDDA.n612 1.69433
R4727 VDDA.n1191 VDDA.n612 1.69433
R4728 VDDA.n1309 VDDA.n634 1.69433
R4729 VDDA.n1309 VDDA.n631 1.69433
R4730 VDDA.n1309 VDDA.n628 1.69433
R4731 VDDA.n1309 VDDA.n625 1.69433
R4732 VDDA.n1309 VDDA.n622 1.69433
R4733 VDDA.n1309 VDDA.n619 1.69433
R4734 VDDA.n1309 VDDA.n616 1.69433
R4735 VDDA.n2406 VDDA.n1331 1.69433
R4736 VDDA.n2406 VDDA.n1328 1.69433
R4737 VDDA.n2406 VDDA.n1325 1.69433
R4738 VDDA.n2406 VDDA.n1322 1.69433
R4739 VDDA.n2406 VDDA.n1319 1.69433
R4740 VDDA.n2406 VDDA.n1316 1.69433
R4741 VDDA.n2406 VDDA.n1313 1.69433
R4742 VDDA.n2405 VDDA.n1489 1.69433
R4743 VDDA.n2405 VDDA.n1486 1.69433
R4744 VDDA.n2405 VDDA.n1483 1.69433
R4745 VDDA.n2405 VDDA.n1480 1.69433
R4746 VDDA.n2405 VDDA.n1477 1.69433
R4747 VDDA.n2405 VDDA.n1474 1.69433
R4748 VDDA.n2405 VDDA.n1471 1.69433
R4749 VDDA.n515 VDDA.n197 1.69433
R4750 VDDA.n497 VDDA.n197 1.69433
R4751 VDDA.n485 VDDA.n197 1.69433
R4752 VDDA.n467 VDDA.n197 1.69433
R4753 VDDA.n455 VDDA.n197 1.69433
R4754 VDDA.n437 VDDA.n197 1.69433
R4755 VDDA.n425 VDDA.n197 1.69433
R4756 VDDA.n2589 VDDA.n219 1.69433
R4757 VDDA.n2589 VDDA.n216 1.69433
R4758 VDDA.n2589 VDDA.n213 1.69433
R4759 VDDA.n2589 VDDA.n210 1.69433
R4760 VDDA.n2589 VDDA.n207 1.69433
R4761 VDDA.n2589 VDDA.n204 1.69433
R4762 VDDA.n2589 VDDA.n201 1.69433
R4763 VDDA.n2749 VDDA.n2611 1.69433
R4764 VDDA.n2749 VDDA.n2608 1.69433
R4765 VDDA.n2749 VDDA.n2605 1.69433
R4766 VDDA.n2749 VDDA.n2602 1.69433
R4767 VDDA.n2749 VDDA.n2599 1.69433
R4768 VDDA.n2749 VDDA.n2596 1.69433
R4769 VDDA.n2749 VDDA.n2593 1.69433
R4770 VDDA.n2909 VDDA.n19 1.69433
R4771 VDDA.n2891 VDDA.n19 1.69433
R4772 VDDA.n2879 VDDA.n19 1.69433
R4773 VDDA.n2861 VDDA.n19 1.69433
R4774 VDDA.n2849 VDDA.n19 1.69433
R4775 VDDA.n2831 VDDA.n19 1.69433
R4776 VDDA.n2819 VDDA.n19 1.69433
R4777 VDDA.n2937 VDDA.n41 1.69433
R4778 VDDA.n2937 VDDA.n38 1.69433
R4779 VDDA.n2937 VDDA.n35 1.69433
R4780 VDDA.n2937 VDDA.n32 1.69433
R4781 VDDA.n2937 VDDA.n29 1.69433
R4782 VDDA.n2937 VDDA.n26 1.69433
R4783 VDDA.n2937 VDDA.n23 1.69433
R4784 VDDA.n1728 VDDA.n1579 1.69433
R4785 VDDA.n1728 VDDA.n1576 1.69433
R4786 VDDA.n1728 VDDA.n1573 1.69433
R4787 VDDA.n1728 VDDA.n1570 1.69433
R4788 VDDA.n1728 VDDA.n1567 1.69433
R4789 VDDA.n1728 VDDA.n1564 1.69433
R4790 VDDA.n1728 VDDA.n1561 1.69433
R4791 VDDA.n2056 VDDA.n1513 1.69328
R4792 VDDA.n2056 VDDA.n1510 1.69328
R4793 VDDA.n2056 VDDA.n1507 1.69328
R4794 VDDA.n2056 VDDA.n1504 1.69328
R4795 VDDA.n2056 VDDA.n1501 1.69328
R4796 VDDA.n2056 VDDA.n1498 1.69328
R4797 VDDA.n2056 VDDA.n1495 1.69328
R4798 VDDA.n961 VDDA.n812 1.6924
R4799 VDDA.n961 VDDA.n811 1.6924
R4800 VDDA.n961 VDDA.n809 1.6924
R4801 VDDA.n961 VDDA.n808 1.6924
R4802 VDDA.n961 VDDA.n806 1.6924
R4803 VDDA.n961 VDDA.n805 1.6924
R4804 VDDA.n961 VDDA.n803 1.6924
R4805 VDDA.n961 VDDA.n802 1.6924
R4806 VDDA.n961 VDDA.n800 1.6924
R4807 VDDA.n961 VDDA.n799 1.6924
R4808 VDDA.n961 VDDA.n797 1.6924
R4809 VDDA.n961 VDDA.n796 1.6924
R4810 VDDA.n961 VDDA.n794 1.6924
R4811 VDDA.n961 VDDA.n793 1.6924
R4812 VDDA.n961 VDDA.n791 1.6924
R4813 VDDA.n961 VDDA.n790 1.6924
R4814 VDDA.n1121 VDDA.n1120 1.6924
R4815 VDDA.n1121 VDDA.n984 1.6924
R4816 VDDA.n1121 VDDA.n982 1.6924
R4817 VDDA.n1121 VDDA.n981 1.6924
R4818 VDDA.n1121 VDDA.n979 1.6924
R4819 VDDA.n1121 VDDA.n978 1.6924
R4820 VDDA.n1121 VDDA.n976 1.6924
R4821 VDDA.n1121 VDDA.n975 1.6924
R4822 VDDA.n1121 VDDA.n973 1.6924
R4823 VDDA.n1121 VDDA.n972 1.6924
R4824 VDDA.n1121 VDDA.n970 1.6924
R4825 VDDA.n1121 VDDA.n969 1.6924
R4826 VDDA.n1121 VDDA.n967 1.6924
R4827 VDDA.n1121 VDDA.n966 1.6924
R4828 VDDA.n1121 VDDA.n964 1.6924
R4829 VDDA.n1121 VDDA.n963 1.6924
R4830 VDDA.n1291 VDDA.n612 1.6924
R4831 VDDA.n1283 VDDA.n612 1.6924
R4832 VDDA.n1273 VDDA.n612 1.6924
R4833 VDDA.n1271 VDDA.n612 1.6924
R4834 VDDA.n1261 VDDA.n612 1.6924
R4835 VDDA.n1253 VDDA.n612 1.6924
R4836 VDDA.n1243 VDDA.n612 1.6924
R4837 VDDA.n1241 VDDA.n612 1.6924
R4838 VDDA.n1231 VDDA.n612 1.6924
R4839 VDDA.n1223 VDDA.n612 1.6924
R4840 VDDA.n1213 VDDA.n612 1.6924
R4841 VDDA.n1211 VDDA.n612 1.6924
R4842 VDDA.n1201 VDDA.n612 1.6924
R4843 VDDA.n1193 VDDA.n612 1.6924
R4844 VDDA.n1183 VDDA.n612 1.6924
R4845 VDDA.n1181 VDDA.n612 1.6924
R4846 VDDA.n1309 VDDA.n636 1.6924
R4847 VDDA.n1309 VDDA.n635 1.6924
R4848 VDDA.n1309 VDDA.n633 1.6924
R4849 VDDA.n1309 VDDA.n632 1.6924
R4850 VDDA.n1309 VDDA.n630 1.6924
R4851 VDDA.n1309 VDDA.n629 1.6924
R4852 VDDA.n1309 VDDA.n627 1.6924
R4853 VDDA.n1309 VDDA.n626 1.6924
R4854 VDDA.n1309 VDDA.n624 1.6924
R4855 VDDA.n1309 VDDA.n623 1.6924
R4856 VDDA.n1309 VDDA.n621 1.6924
R4857 VDDA.n1309 VDDA.n620 1.6924
R4858 VDDA.n1309 VDDA.n618 1.6924
R4859 VDDA.n1309 VDDA.n617 1.6924
R4860 VDDA.n1309 VDDA.n615 1.6924
R4861 VDDA.n1309 VDDA.n614 1.6924
R4862 VDDA.n2406 VDDA.n1468 1.6924
R4863 VDDA.n2406 VDDA.n1332 1.6924
R4864 VDDA.n2406 VDDA.n1330 1.6924
R4865 VDDA.n2406 VDDA.n1329 1.6924
R4866 VDDA.n2406 VDDA.n1327 1.6924
R4867 VDDA.n2406 VDDA.n1326 1.6924
R4868 VDDA.n2406 VDDA.n1324 1.6924
R4869 VDDA.n2406 VDDA.n1323 1.6924
R4870 VDDA.n2406 VDDA.n1321 1.6924
R4871 VDDA.n2406 VDDA.n1320 1.6924
R4872 VDDA.n2406 VDDA.n1318 1.6924
R4873 VDDA.n2406 VDDA.n1317 1.6924
R4874 VDDA.n2406 VDDA.n1315 1.6924
R4875 VDDA.n2406 VDDA.n1314 1.6924
R4876 VDDA.n2406 VDDA.n1312 1.6924
R4877 VDDA.n2406 VDDA.n1311 1.6924
R4878 VDDA.n2405 VDDA.n1491 1.6924
R4879 VDDA.n2405 VDDA.n1490 1.6924
R4880 VDDA.n2405 VDDA.n1488 1.6924
R4881 VDDA.n2405 VDDA.n1487 1.6924
R4882 VDDA.n2405 VDDA.n1485 1.6924
R4883 VDDA.n2405 VDDA.n1484 1.6924
R4884 VDDA.n2405 VDDA.n1482 1.6924
R4885 VDDA.n2405 VDDA.n1481 1.6924
R4886 VDDA.n2405 VDDA.n1479 1.6924
R4887 VDDA.n2405 VDDA.n1478 1.6924
R4888 VDDA.n2405 VDDA.n1476 1.6924
R4889 VDDA.n2405 VDDA.n1475 1.6924
R4890 VDDA.n2405 VDDA.n1473 1.6924
R4891 VDDA.n2405 VDDA.n1472 1.6924
R4892 VDDA.n2405 VDDA.n1470 1.6924
R4893 VDDA.n525 VDDA.n197 1.6924
R4894 VDDA.n517 VDDA.n197 1.6924
R4895 VDDA.n507 VDDA.n197 1.6924
R4896 VDDA.n505 VDDA.n197 1.6924
R4897 VDDA.n495 VDDA.n197 1.6924
R4898 VDDA.n487 VDDA.n197 1.6924
R4899 VDDA.n477 VDDA.n197 1.6924
R4900 VDDA.n475 VDDA.n197 1.6924
R4901 VDDA.n465 VDDA.n197 1.6924
R4902 VDDA.n457 VDDA.n197 1.6924
R4903 VDDA.n447 VDDA.n197 1.6924
R4904 VDDA.n445 VDDA.n197 1.6924
R4905 VDDA.n435 VDDA.n197 1.6924
R4906 VDDA.n427 VDDA.n197 1.6924
R4907 VDDA.n417 VDDA.n197 1.6924
R4908 VDDA.n415 VDDA.n197 1.6924
R4909 VDDA.n2589 VDDA.n221 1.6924
R4910 VDDA.n2589 VDDA.n220 1.6924
R4911 VDDA.n2589 VDDA.n218 1.6924
R4912 VDDA.n2589 VDDA.n217 1.6924
R4913 VDDA.n2589 VDDA.n215 1.6924
R4914 VDDA.n2589 VDDA.n214 1.6924
R4915 VDDA.n2589 VDDA.n212 1.6924
R4916 VDDA.n2589 VDDA.n211 1.6924
R4917 VDDA.n2589 VDDA.n209 1.6924
R4918 VDDA.n2589 VDDA.n208 1.6924
R4919 VDDA.n2589 VDDA.n206 1.6924
R4920 VDDA.n2589 VDDA.n205 1.6924
R4921 VDDA.n2589 VDDA.n203 1.6924
R4922 VDDA.n2589 VDDA.n202 1.6924
R4923 VDDA.n2589 VDDA.n200 1.6924
R4924 VDDA.n2589 VDDA.n199 1.6924
R4925 VDDA.n2749 VDDA.n2748 1.6924
R4926 VDDA.n2749 VDDA.n2612 1.6924
R4927 VDDA.n2749 VDDA.n2610 1.6924
R4928 VDDA.n2749 VDDA.n2609 1.6924
R4929 VDDA.n2749 VDDA.n2607 1.6924
R4930 VDDA.n2749 VDDA.n2606 1.6924
R4931 VDDA.n2749 VDDA.n2604 1.6924
R4932 VDDA.n2749 VDDA.n2603 1.6924
R4933 VDDA.n2749 VDDA.n2601 1.6924
R4934 VDDA.n2749 VDDA.n2600 1.6924
R4935 VDDA.n2749 VDDA.n2598 1.6924
R4936 VDDA.n2749 VDDA.n2597 1.6924
R4937 VDDA.n2749 VDDA.n2595 1.6924
R4938 VDDA.n2749 VDDA.n2594 1.6924
R4939 VDDA.n2749 VDDA.n2592 1.6924
R4940 VDDA.n2749 VDDA.n2591 1.6924
R4941 VDDA.n2919 VDDA.n19 1.6924
R4942 VDDA.n2911 VDDA.n19 1.6924
R4943 VDDA.n2901 VDDA.n19 1.6924
R4944 VDDA.n2899 VDDA.n19 1.6924
R4945 VDDA.n2889 VDDA.n19 1.6924
R4946 VDDA.n2881 VDDA.n19 1.6924
R4947 VDDA.n2871 VDDA.n19 1.6924
R4948 VDDA.n2869 VDDA.n19 1.6924
R4949 VDDA.n2859 VDDA.n19 1.6924
R4950 VDDA.n2851 VDDA.n19 1.6924
R4951 VDDA.n2841 VDDA.n19 1.6924
R4952 VDDA.n2839 VDDA.n19 1.6924
R4953 VDDA.n2829 VDDA.n19 1.6924
R4954 VDDA.n2821 VDDA.n19 1.6924
R4955 VDDA.n2811 VDDA.n19 1.6924
R4956 VDDA.n2809 VDDA.n19 1.6924
R4957 VDDA.n2937 VDDA.n43 1.6924
R4958 VDDA.n2937 VDDA.n42 1.6924
R4959 VDDA.n2937 VDDA.n40 1.6924
R4960 VDDA.n2937 VDDA.n39 1.6924
R4961 VDDA.n2937 VDDA.n37 1.6924
R4962 VDDA.n2937 VDDA.n36 1.6924
R4963 VDDA.n2937 VDDA.n34 1.6924
R4964 VDDA.n2937 VDDA.n33 1.6924
R4965 VDDA.n2937 VDDA.n31 1.6924
R4966 VDDA.n2937 VDDA.n30 1.6924
R4967 VDDA.n2937 VDDA.n28 1.6924
R4968 VDDA.n2937 VDDA.n27 1.6924
R4969 VDDA.n2937 VDDA.n25 1.6924
R4970 VDDA.n2937 VDDA.n24 1.6924
R4971 VDDA.n2937 VDDA.n22 1.6924
R4972 VDDA.n2937 VDDA.n21 1.6924
R4973 VDDA.n1728 VDDA.n1581 1.6924
R4974 VDDA.n1728 VDDA.n1580 1.6924
R4975 VDDA.n1728 VDDA.n1578 1.6924
R4976 VDDA.n1728 VDDA.n1577 1.6924
R4977 VDDA.n1728 VDDA.n1575 1.6924
R4978 VDDA.n1728 VDDA.n1574 1.6924
R4979 VDDA.n1728 VDDA.n1572 1.6924
R4980 VDDA.n1728 VDDA.n1571 1.6924
R4981 VDDA.n1728 VDDA.n1569 1.6924
R4982 VDDA.n1728 VDDA.n1568 1.6924
R4983 VDDA.n1728 VDDA.n1566 1.6924
R4984 VDDA.n1728 VDDA.n1565 1.6924
R4985 VDDA.n1728 VDDA.n1563 1.6924
R4986 VDDA.n1728 VDDA.n1562 1.6924
R4987 VDDA.n1728 VDDA.n1560 1.6924
R4988 VDDA.n1728 VDDA.n1559 1.6924
R4989 VDDA.n2056 VDDA.n1515 1.69118
R4990 VDDA.n2056 VDDA.n1514 1.69118
R4991 VDDA.n2056 VDDA.n1512 1.69118
R4992 VDDA.n2056 VDDA.n1511 1.69118
R4993 VDDA.n2056 VDDA.n1509 1.69118
R4994 VDDA.n2056 VDDA.n1508 1.69118
R4995 VDDA.n2056 VDDA.n1506 1.69118
R4996 VDDA.n2056 VDDA.n1505 1.69118
R4997 VDDA.n2056 VDDA.n1503 1.69118
R4998 VDDA.n2056 VDDA.n1502 1.69118
R4999 VDDA.n2056 VDDA.n1500 1.69118
R5000 VDDA.n2056 VDDA.n1499 1.69118
R5001 VDDA.n2056 VDDA.n1497 1.69118
R5002 VDDA.n2056 VDDA.n1496 1.69118
R5003 VDDA.n2056 VDDA.n1494 1.69118
R5004 VDDA.n2056 VDDA.n1493 1.69118
R5005 VDDA.n2458 VDDA.n2456 1.63212
R5006 VDDA.n2471 VDDA.n2470 1.63212
R5007 VDDA.n2462 VDDA.n2461 1.56962
R5008 VDDA.n2475 VDDA.n2474 1.56962
R5009 VDDA.n1938 VDDA.n1541 1.56177
R5010 VDDA.n1915 VDDA.n1541 1.50969
R5011 VDDA.n1552 VDDA.n1541 1.44719
R5012 VDDA.n2092 VDDA.n2091 1.26222
R5013 VDDA.n1801 VDDA.n1800 1.20209
R5014 VDDA.n2550 VDDA.n2549 1.14633
R5015 VDDA.n2436 VDDA.n599 1.14633
R5016 VDDA.n2405 VDDA.n1469 1.12311
R5017 VDDA.n2540 VDDA.n2538 1.06821
R5018 VDDA.n596 VDDA.n588 1.06821
R5019 VDDA.n2575 VDDA.n2574 0.953625
R5020 VDDA.n2418 VDDA.n2414 0.953625
R5021 VDDA.n2098 VDDA.n2097 0.943208
R5022 VDDA.n2448 VDDA.n2445 0.932792
R5023 VDDA.n2514 VDDA.n2493 0.932792
R5024 VDDA.n2235 VDDA.n2234 0.880708
R5025 VDDA.n2158 VDDA.n2157 0.865083
R5026 VDDA.n2285 VDDA.n2284 0.807792
R5027 VDDA.n2090 VDDA.n2089 0.75233
R5028 VDDA.n2164 VDDA.n2163 0.672375
R5029 VDDA.n2091 VDDA.n2090 0.648711
R5030 VDDA.n2582 VDDA.n2580 0.646333
R5031 VDDA.n2413 VDDA.n606 0.646333
R5032 VDDA.n3123 VDDA.n2937 0.546104
R5033 VDDA.n2570 VDDA.n2569 0.521333
R5034 VDDA.n2429 VDDA.n2420 0.521333
R5035 VDDA.n2553 VDDA.n2515 0.495292
R5036 VDDA.n2440 VDDA.n2439 0.495292
R5037 VDDA.n2292 VDDA.n2290 0.448417
R5038 VDDA.n2483 VDDA.n2482 0.417167
R5039 VDDA.n2510 VDDA.n2497 0.3755
R5040 VDDA.n2499 VDDA.n2497 0.3755
R5041 VDDA.n2501 VDDA.n2499 0.3755
R5042 VDDA.n2503 VDDA.n2501 0.3755
R5043 VDDA.n2505 VDDA.n2503 0.3755
R5044 VDDA.n556 VDDA.n554 0.3755
R5045 VDDA.n554 VDDA.n552 0.3755
R5046 VDDA.n552 VDDA.n550 0.3755
R5047 VDDA.n550 VDDA.n548 0.3755
R5048 VDDA.n561 VDDA.n548 0.3755
R5049 VDDA.n2148 VDDA.n2147 0.333833
R5050 VDDA.n2229 VDDA.n2228 0.328625
R5051 VDDA.n584 VDDA.n583 0.323417
R5052 VDDA.n2536 VDDA.n2535 0.323417
R5053 VDDA.n2282 VDDA.n2281 0.292167
R5054 VDDA.n2278 VDDA.n2277 0.292167
R5055 VDDA.n2271 VDDA.n2270 0.292167
R5056 VDDA.n2241 VDDA.n2240 0.292167
R5057 VDDA.n2755 VDDA.n192 0.28175
R5058 VDDA.n2926 VDDA.n2757 0.28175
R5059 VDDA.n2929 VDDA.n2928 0.28175
R5060 VDDA.n1127 VDDA.n784 0.28175
R5061 VDDA.n1298 VDDA.n1129 0.28175
R5062 VDDA.n1302 VDDA.n1300 0.28175
R5063 VDDA.n594 VDDA.n593 0.266125
R5064 VDDA.n2547 VDDA.n2546 0.266125
R5065 VDDA.n2564 VDDA.n2555 0.266125
R5066 VDDA.n2435 VDDA.n2434 0.266125
R5067 VDDA.n2146 VDDA.n2145 0.2505
R5068 VDDA.n2156 VDDA.n2155 0.2505
R5069 VDDA.n1917 VDDA.n1916 0.229667
R5070 VDDA.n1937 VDDA.n1936 0.229667
R5071 VDDA.n2234 VDDA.n2229 0.229667
R5072 VDDA.n2466 VDDA.n2462 0.214042
R5073 VDDA.n2476 VDDA.n2475 0.214042
R5074 VDDA.n1918 VDDA.n1548 0.208833
R5075 VDDA.n1918 VDDA.n1917 0.208833
R5076 VDDA.n1930 VDDA.n1542 0.208833
R5077 VDDA.n1936 VDDA.n1542 0.208833
R5078 VDDA.n2196 VDDA.n2182 0.208833
R5079 VDDA.n2190 VDDA.n2182 0.208833
R5080 VDDA.n2190 VDDA.n2189 0.208833
R5081 VDDA.n2205 VDDA.n2203 0.208833
R5082 VDDA.n2206 VDDA.n2205 0.208833
R5083 VDDA.n2206 VDDA.n2175 0.208833
R5084 VDDA.n2228 VDDA.n2227 0.188
R5085 VDDA.n2227 VDDA.n2226 0.188
R5086 VDDA.n2226 VDDA.n2225 0.188
R5087 VDDA.n2225 VDDA.n2224 0.188
R5088 VDDA.n2224 VDDA.n2223 0.188
R5089 VDDA.n2223 VDDA.n2222 0.188
R5090 VDDA.n2222 VDDA.n2221 0.188
R5091 VDDA.n2221 VDDA.n2220 0.188
R5092 VDDA.n2450 VDDA.n2448 0.172375
R5093 VDDA.n2485 VDDA.n2450 0.172375
R5094 VDDA.n2451 VDDA.n542 0.172375
R5095 VDDA.n2493 VDDA.n542 0.172375
R5096 VDDA.t117 VDDA.t414 0.1603
R5097 VDDA.t30 VDDA.t76 0.1603
R5098 VDDA.t49 VDDA.t55 0.1603
R5099 VDDA.t170 VDDA.t379 0.1603
R5100 VDDA.t27 VDDA.t42 0.1603
R5101 VDDA.n1944 VDDA.n1943 0.159591
R5102 VDDA.n1945 VDDA.n1944 0.159591
R5103 VDDA.n1945 VDDA.n1539 0.159591
R5104 VDDA.n1955 VDDA.n1537 0.159591
R5105 VDDA.n1963 VDDA.n1537 0.159591
R5106 VDDA.n1964 VDDA.n1963 0.159591
R5107 VDDA.n1974 VDDA.n1973 0.159591
R5108 VDDA.n1975 VDDA.n1974 0.159591
R5109 VDDA.n1975 VDDA.n1533 0.159591
R5110 VDDA.n1985 VDDA.n1531 0.159591
R5111 VDDA.n1993 VDDA.n1531 0.159591
R5112 VDDA.n1994 VDDA.n1993 0.159591
R5113 VDDA.n2004 VDDA.n2003 0.159591
R5114 VDDA.n2005 VDDA.n2004 0.159591
R5115 VDDA.n2005 VDDA.n1527 0.159591
R5116 VDDA.n2015 VDDA.n1525 0.159591
R5117 VDDA.n2023 VDDA.n1525 0.159591
R5118 VDDA.n2024 VDDA.n2023 0.159591
R5119 VDDA.n2034 VDDA.n2033 0.159591
R5120 VDDA.n2035 VDDA.n2034 0.159591
R5121 VDDA.n2035 VDDA.n1521 0.159591
R5122 VDDA.n2045 VDDA.n1519 0.159591
R5123 VDDA.n2053 VDDA.n1519 0.159591
R5124 VDDA.n1942 VDDA.n1540 0.159591
R5125 VDDA.n1948 VDDA.n1540 0.159591
R5126 VDDA.n1949 VDDA.n1948 0.159591
R5127 VDDA.n1959 VDDA.n1958 0.159591
R5128 VDDA.n1962 VDDA.n1959 0.159591
R5129 VDDA.n1962 VDDA.n1536 0.159591
R5130 VDDA.n1972 VDDA.n1534 0.159591
R5131 VDDA.n1978 VDDA.n1534 0.159591
R5132 VDDA.n1979 VDDA.n1978 0.159591
R5133 VDDA.n1989 VDDA.n1988 0.159591
R5134 VDDA.n1992 VDDA.n1989 0.159591
R5135 VDDA.n1992 VDDA.n1530 0.159591
R5136 VDDA.n2002 VDDA.n1528 0.159591
R5137 VDDA.n2008 VDDA.n1528 0.159591
R5138 VDDA.n2009 VDDA.n2008 0.159591
R5139 VDDA.n2019 VDDA.n2018 0.159591
R5140 VDDA.n2022 VDDA.n2019 0.159591
R5141 VDDA.n2022 VDDA.n1524 0.159591
R5142 VDDA.n2032 VDDA.n1522 0.159591
R5143 VDDA.n2038 VDDA.n1522 0.159591
R5144 VDDA.n2039 VDDA.n2038 0.159591
R5145 VDDA.n2049 VDDA.n2048 0.159591
R5146 VDDA.n2052 VDDA.n2049 0.159591
R5147 VDDA.n2052 VDDA.n1518 0.159591
R5148 VDDA.n1607 VDDA.t53 0.159278
R5149 VDDA.n1608 VDDA.t50 0.159278
R5150 VDDA.n1609 VDDA.t188 0.159278
R5151 VDDA.n1610 VDDA.t169 0.159278
R5152 VDDA.n1943 VDDA.n1939 0.148227
R5153 VDDA.n1953 VDDA.n1539 0.148227
R5154 VDDA.n1955 VDDA.n1954 0.148227
R5155 VDDA.n1965 VDDA.n1964 0.148227
R5156 VDDA.n1973 VDDA.n1535 0.148227
R5157 VDDA.n1983 VDDA.n1533 0.148227
R5158 VDDA.n1985 VDDA.n1984 0.148227
R5159 VDDA.n1995 VDDA.n1994 0.148227
R5160 VDDA.n2003 VDDA.n1529 0.148227
R5161 VDDA.n2013 VDDA.n1527 0.148227
R5162 VDDA.n2015 VDDA.n2014 0.148227
R5163 VDDA.n2025 VDDA.n2024 0.148227
R5164 VDDA.n2033 VDDA.n1523 0.148227
R5165 VDDA.n2043 VDDA.n1521 0.148227
R5166 VDDA.n2045 VDDA.n2044 0.148227
R5167 VDDA.n1942 VDDA.n1940 0.148227
R5168 VDDA.n1952 VDDA.n1949 0.148227
R5169 VDDA.n1958 VDDA.n1538 0.148227
R5170 VDDA.n1968 VDDA.n1536 0.148227
R5171 VDDA.n1972 VDDA.n1969 0.148227
R5172 VDDA.n1982 VDDA.n1979 0.148227
R5173 VDDA.n1988 VDDA.n1532 0.148227
R5174 VDDA.n1998 VDDA.n1530 0.148227
R5175 VDDA.n2002 VDDA.n1999 0.148227
R5176 VDDA.n2012 VDDA.n2009 0.148227
R5177 VDDA.n2018 VDDA.n1526 0.148227
R5178 VDDA.n2028 VDDA.n1524 0.148227
R5179 VDDA.n2032 VDDA.n2029 0.148227
R5180 VDDA.n2042 VDDA.n2039 0.148227
R5181 VDDA.n2048 VDDA.n1520 0.148227
R5182 VDDA.n1614 VDDA.n1605 0.146333
R5183 VDDA.n1620 VDDA.n1605 0.146333
R5184 VDDA.n1621 VDDA.n1620 0.146333
R5185 VDDA.n1631 VDDA.n1630 0.146333
R5186 VDDA.n1634 VDDA.n1631 0.146333
R5187 VDDA.n1634 VDDA.n1601 0.146333
R5188 VDDA.n1644 VDDA.n1599 0.146333
R5189 VDDA.n1650 VDDA.n1599 0.146333
R5190 VDDA.n1651 VDDA.n1650 0.146333
R5191 VDDA.n1661 VDDA.n1660 0.146333
R5192 VDDA.n1664 VDDA.n1661 0.146333
R5193 VDDA.n1664 VDDA.n1595 0.146333
R5194 VDDA.n1674 VDDA.n1593 0.146333
R5195 VDDA.n1680 VDDA.n1593 0.146333
R5196 VDDA.n1681 VDDA.n1680 0.146333
R5197 VDDA.n1691 VDDA.n1690 0.146333
R5198 VDDA.n1694 VDDA.n1691 0.146333
R5199 VDDA.n1694 VDDA.n1589 0.146333
R5200 VDDA.n1704 VDDA.n1587 0.146333
R5201 VDDA.n1710 VDDA.n1587 0.146333
R5202 VDDA.n1711 VDDA.n1710 0.146333
R5203 VDDA.n1721 VDDA.n1720 0.146333
R5204 VDDA.n1724 VDDA.n1721 0.146333
R5205 VDDA.n1724 VDDA.n1583 0.146333
R5206 VDDA.n2291 VDDA.n2080 0.146333
R5207 VDDA.n2297 VDDA.n2080 0.146333
R5208 VDDA.n2298 VDDA.n2297 0.146333
R5209 VDDA.n2308 VDDA.n2307 0.146333
R5210 VDDA.n2311 VDDA.n2308 0.146333
R5211 VDDA.n2311 VDDA.n2076 0.146333
R5212 VDDA.n2321 VDDA.n2074 0.146333
R5213 VDDA.n2327 VDDA.n2074 0.146333
R5214 VDDA.n2328 VDDA.n2327 0.146333
R5215 VDDA.n2338 VDDA.n2337 0.146333
R5216 VDDA.n2341 VDDA.n2338 0.146333
R5217 VDDA.n2341 VDDA.n2070 0.146333
R5218 VDDA.n2351 VDDA.n2068 0.146333
R5219 VDDA.n2357 VDDA.n2068 0.146333
R5220 VDDA.n2358 VDDA.n2357 0.146333
R5221 VDDA.n2368 VDDA.n2367 0.146333
R5222 VDDA.n2371 VDDA.n2368 0.146333
R5223 VDDA.n2371 VDDA.n2064 0.146333
R5224 VDDA.n2381 VDDA.n2062 0.146333
R5225 VDDA.n2387 VDDA.n2062 0.146333
R5226 VDDA.n2388 VDDA.n2387 0.146333
R5227 VDDA.n2398 VDDA.n2397 0.146333
R5228 VDDA.n2401 VDDA.n2398 0.146333
R5229 VDDA.n2401 VDDA.n2058 0.146333
R5230 VDDA.n91 VDDA.n87 0.146333
R5231 VDDA.n95 VDDA.n87 0.146333
R5232 VDDA.n96 VDDA.n95 0.146333
R5233 VDDA.n104 VDDA.n103 0.146333
R5234 VDDA.n107 VDDA.n104 0.146333
R5235 VDDA.n107 VDDA.n79 0.146333
R5236 VDDA.n115 VDDA.n75 0.146333
R5237 VDDA.n119 VDDA.n75 0.146333
R5238 VDDA.n120 VDDA.n119 0.146333
R5239 VDDA.n128 VDDA.n127 0.146333
R5240 VDDA.n131 VDDA.n128 0.146333
R5241 VDDA.n131 VDDA.n67 0.146333
R5242 VDDA.n139 VDDA.n63 0.146333
R5243 VDDA.n143 VDDA.n63 0.146333
R5244 VDDA.n144 VDDA.n143 0.146333
R5245 VDDA.n152 VDDA.n151 0.146333
R5246 VDDA.n155 VDDA.n152 0.146333
R5247 VDDA.n155 VDDA.n55 0.146333
R5248 VDDA.n163 VDDA.n51 0.146333
R5249 VDDA.n167 VDDA.n51 0.146333
R5250 VDDA.n168 VDDA.n167 0.146333
R5251 VDDA.n176 VDDA.n175 0.146333
R5252 VDDA.n179 VDDA.n176 0.146333
R5253 VDDA.n179 VDDA.n45 0.146333
R5254 VDDA.n2807 VDDA.n2804 0.146333
R5255 VDDA.n2813 VDDA.n2804 0.146333
R5256 VDDA.n2813 VDDA.n2802 0.146333
R5257 VDDA.n2823 VDDA.n2798 0.146333
R5258 VDDA.n2827 VDDA.n2798 0.146333
R5259 VDDA.n2827 VDDA.n2796 0.146333
R5260 VDDA.n2837 VDDA.n2792 0.146333
R5261 VDDA.n2843 VDDA.n2792 0.146333
R5262 VDDA.n2843 VDDA.n2790 0.146333
R5263 VDDA.n2853 VDDA.n2786 0.146333
R5264 VDDA.n2857 VDDA.n2786 0.146333
R5265 VDDA.n2857 VDDA.n2784 0.146333
R5266 VDDA.n2867 VDDA.n2780 0.146333
R5267 VDDA.n2873 VDDA.n2780 0.146333
R5268 VDDA.n2873 VDDA.n2778 0.146333
R5269 VDDA.n2883 VDDA.n2774 0.146333
R5270 VDDA.n2887 VDDA.n2774 0.146333
R5271 VDDA.n2887 VDDA.n2772 0.146333
R5272 VDDA.n2897 VDDA.n2768 0.146333
R5273 VDDA.n2903 VDDA.n2768 0.146333
R5274 VDDA.n2903 VDDA.n2766 0.146333
R5275 VDDA.n2913 VDDA.n2762 0.146333
R5276 VDDA.n2917 VDDA.n2762 0.146333
R5277 VDDA.n2917 VDDA.n2760 0.146333
R5278 VDDA.n2659 VDDA.n2658 0.146333
R5279 VDDA.n2662 VDDA.n2659 0.146333
R5280 VDDA.n2662 VDDA.n2652 0.146333
R5281 VDDA.n2670 VDDA.n2648 0.146333
R5282 VDDA.n2674 VDDA.n2648 0.146333
R5283 VDDA.n2675 VDDA.n2674 0.146333
R5284 VDDA.n2683 VDDA.n2682 0.146333
R5285 VDDA.n2686 VDDA.n2683 0.146333
R5286 VDDA.n2686 VDDA.n2640 0.146333
R5287 VDDA.n2694 VDDA.n2636 0.146333
R5288 VDDA.n2698 VDDA.n2636 0.146333
R5289 VDDA.n2699 VDDA.n2698 0.146333
R5290 VDDA.n2707 VDDA.n2706 0.146333
R5291 VDDA.n2710 VDDA.n2707 0.146333
R5292 VDDA.n2710 VDDA.n2628 0.146333
R5293 VDDA.n2718 VDDA.n2624 0.146333
R5294 VDDA.n2722 VDDA.n2624 0.146333
R5295 VDDA.n2723 VDDA.n2722 0.146333
R5296 VDDA.n2731 VDDA.n2730 0.146333
R5297 VDDA.n2734 VDDA.n2731 0.146333
R5298 VDDA.n2734 VDDA.n2616 0.146333
R5299 VDDA.n2742 VDDA.n2614 0.146333
R5300 VDDA.n2746 VDDA.n2614 0.146333
R5301 VDDA.n2746 VDDA.n195 0.146333
R5302 VDDA.n269 VDDA.n265 0.146333
R5303 VDDA.n273 VDDA.n265 0.146333
R5304 VDDA.n274 VDDA.n273 0.146333
R5305 VDDA.n282 VDDA.n281 0.146333
R5306 VDDA.n285 VDDA.n282 0.146333
R5307 VDDA.n285 VDDA.n257 0.146333
R5308 VDDA.n293 VDDA.n253 0.146333
R5309 VDDA.n297 VDDA.n253 0.146333
R5310 VDDA.n298 VDDA.n297 0.146333
R5311 VDDA.n306 VDDA.n305 0.146333
R5312 VDDA.n309 VDDA.n306 0.146333
R5313 VDDA.n309 VDDA.n245 0.146333
R5314 VDDA.n317 VDDA.n241 0.146333
R5315 VDDA.n321 VDDA.n241 0.146333
R5316 VDDA.n322 VDDA.n321 0.146333
R5317 VDDA.n330 VDDA.n329 0.146333
R5318 VDDA.n333 VDDA.n330 0.146333
R5319 VDDA.n333 VDDA.n233 0.146333
R5320 VDDA.n341 VDDA.n229 0.146333
R5321 VDDA.n345 VDDA.n229 0.146333
R5322 VDDA.n346 VDDA.n345 0.146333
R5323 VDDA.n354 VDDA.n353 0.146333
R5324 VDDA.n357 VDDA.n354 0.146333
R5325 VDDA.n357 VDDA.n223 0.146333
R5326 VDDA.n413 VDDA.n410 0.146333
R5327 VDDA.n419 VDDA.n410 0.146333
R5328 VDDA.n419 VDDA.n408 0.146333
R5329 VDDA.n429 VDDA.n404 0.146333
R5330 VDDA.n433 VDDA.n404 0.146333
R5331 VDDA.n433 VDDA.n402 0.146333
R5332 VDDA.n443 VDDA.n398 0.146333
R5333 VDDA.n449 VDDA.n398 0.146333
R5334 VDDA.n449 VDDA.n396 0.146333
R5335 VDDA.n459 VDDA.n392 0.146333
R5336 VDDA.n463 VDDA.n392 0.146333
R5337 VDDA.n463 VDDA.n390 0.146333
R5338 VDDA.n473 VDDA.n386 0.146333
R5339 VDDA.n479 VDDA.n386 0.146333
R5340 VDDA.n479 VDDA.n384 0.146333
R5341 VDDA.n489 VDDA.n380 0.146333
R5342 VDDA.n493 VDDA.n380 0.146333
R5343 VDDA.n493 VDDA.n378 0.146333
R5344 VDDA.n503 VDDA.n374 0.146333
R5345 VDDA.n509 VDDA.n374 0.146333
R5346 VDDA.n509 VDDA.n372 0.146333
R5347 VDDA.n519 VDDA.n368 0.146333
R5348 VDDA.n523 VDDA.n368 0.146333
R5349 VDDA.n523 VDDA.n366 0.146333
R5350 VDDA.n1379 VDDA.n1378 0.146333
R5351 VDDA.n1382 VDDA.n1379 0.146333
R5352 VDDA.n1382 VDDA.n1372 0.146333
R5353 VDDA.n1390 VDDA.n1368 0.146333
R5354 VDDA.n1394 VDDA.n1368 0.146333
R5355 VDDA.n1395 VDDA.n1394 0.146333
R5356 VDDA.n1403 VDDA.n1402 0.146333
R5357 VDDA.n1406 VDDA.n1403 0.146333
R5358 VDDA.n1406 VDDA.n1360 0.146333
R5359 VDDA.n1414 VDDA.n1356 0.146333
R5360 VDDA.n1418 VDDA.n1356 0.146333
R5361 VDDA.n1419 VDDA.n1418 0.146333
R5362 VDDA.n1427 VDDA.n1426 0.146333
R5363 VDDA.n1430 VDDA.n1427 0.146333
R5364 VDDA.n1430 VDDA.n1348 0.146333
R5365 VDDA.n1438 VDDA.n1344 0.146333
R5366 VDDA.n1442 VDDA.n1344 0.146333
R5367 VDDA.n1443 VDDA.n1442 0.146333
R5368 VDDA.n1451 VDDA.n1450 0.146333
R5369 VDDA.n1454 VDDA.n1451 0.146333
R5370 VDDA.n1454 VDDA.n1336 0.146333
R5371 VDDA.n1462 VDDA.n1334 0.146333
R5372 VDDA.n1466 VDDA.n1334 0.146333
R5373 VDDA.n1466 VDDA.n610 0.146333
R5374 VDDA.n684 VDDA.n680 0.146333
R5375 VDDA.n688 VDDA.n680 0.146333
R5376 VDDA.n689 VDDA.n688 0.146333
R5377 VDDA.n697 VDDA.n696 0.146333
R5378 VDDA.n700 VDDA.n697 0.146333
R5379 VDDA.n700 VDDA.n672 0.146333
R5380 VDDA.n708 VDDA.n668 0.146333
R5381 VDDA.n712 VDDA.n668 0.146333
R5382 VDDA.n713 VDDA.n712 0.146333
R5383 VDDA.n721 VDDA.n720 0.146333
R5384 VDDA.n724 VDDA.n721 0.146333
R5385 VDDA.n724 VDDA.n660 0.146333
R5386 VDDA.n732 VDDA.n656 0.146333
R5387 VDDA.n736 VDDA.n656 0.146333
R5388 VDDA.n737 VDDA.n736 0.146333
R5389 VDDA.n745 VDDA.n744 0.146333
R5390 VDDA.n748 VDDA.n745 0.146333
R5391 VDDA.n748 VDDA.n648 0.146333
R5392 VDDA.n756 VDDA.n644 0.146333
R5393 VDDA.n760 VDDA.n644 0.146333
R5394 VDDA.n761 VDDA.n760 0.146333
R5395 VDDA.n769 VDDA.n768 0.146333
R5396 VDDA.n772 VDDA.n769 0.146333
R5397 VDDA.n772 VDDA.n638 0.146333
R5398 VDDA.n1179 VDDA.n1176 0.146333
R5399 VDDA.n1185 VDDA.n1176 0.146333
R5400 VDDA.n1185 VDDA.n1174 0.146333
R5401 VDDA.n1195 VDDA.n1170 0.146333
R5402 VDDA.n1199 VDDA.n1170 0.146333
R5403 VDDA.n1199 VDDA.n1168 0.146333
R5404 VDDA.n1209 VDDA.n1164 0.146333
R5405 VDDA.n1215 VDDA.n1164 0.146333
R5406 VDDA.n1215 VDDA.n1162 0.146333
R5407 VDDA.n1225 VDDA.n1158 0.146333
R5408 VDDA.n1229 VDDA.n1158 0.146333
R5409 VDDA.n1229 VDDA.n1156 0.146333
R5410 VDDA.n1239 VDDA.n1152 0.146333
R5411 VDDA.n1245 VDDA.n1152 0.146333
R5412 VDDA.n1245 VDDA.n1150 0.146333
R5413 VDDA.n1255 VDDA.n1146 0.146333
R5414 VDDA.n1259 VDDA.n1146 0.146333
R5415 VDDA.n1259 VDDA.n1144 0.146333
R5416 VDDA.n1269 VDDA.n1140 0.146333
R5417 VDDA.n1275 VDDA.n1140 0.146333
R5418 VDDA.n1275 VDDA.n1138 0.146333
R5419 VDDA.n1285 VDDA.n1134 0.146333
R5420 VDDA.n1289 VDDA.n1134 0.146333
R5421 VDDA.n1289 VDDA.n1132 0.146333
R5422 VDDA.n1031 VDDA.n1030 0.146333
R5423 VDDA.n1034 VDDA.n1031 0.146333
R5424 VDDA.n1034 VDDA.n1024 0.146333
R5425 VDDA.n1042 VDDA.n1020 0.146333
R5426 VDDA.n1046 VDDA.n1020 0.146333
R5427 VDDA.n1047 VDDA.n1046 0.146333
R5428 VDDA.n1055 VDDA.n1054 0.146333
R5429 VDDA.n1058 VDDA.n1055 0.146333
R5430 VDDA.n1058 VDDA.n1012 0.146333
R5431 VDDA.n1066 VDDA.n1008 0.146333
R5432 VDDA.n1070 VDDA.n1008 0.146333
R5433 VDDA.n1071 VDDA.n1070 0.146333
R5434 VDDA.n1079 VDDA.n1078 0.146333
R5435 VDDA.n1082 VDDA.n1079 0.146333
R5436 VDDA.n1082 VDDA.n1000 0.146333
R5437 VDDA.n1090 VDDA.n996 0.146333
R5438 VDDA.n1094 VDDA.n996 0.146333
R5439 VDDA.n1095 VDDA.n1094 0.146333
R5440 VDDA.n1103 VDDA.n1102 0.146333
R5441 VDDA.n1106 VDDA.n1103 0.146333
R5442 VDDA.n1106 VDDA.n988 0.146333
R5443 VDDA.n1114 VDDA.n986 0.146333
R5444 VDDA.n1118 VDDA.n986 0.146333
R5445 VDDA.n1118 VDDA.n787 0.146333
R5446 VDDA.n838 VDDA.n836 0.146333
R5447 VDDA.n844 VDDA.n836 0.146333
R5448 VDDA.n845 VDDA.n844 0.146333
R5449 VDDA.n855 VDDA.n854 0.146333
R5450 VDDA.n858 VDDA.n855 0.146333
R5451 VDDA.n858 VDDA.n832 0.146333
R5452 VDDA.n868 VDDA.n830 0.146333
R5453 VDDA.n874 VDDA.n830 0.146333
R5454 VDDA.n875 VDDA.n874 0.146333
R5455 VDDA.n885 VDDA.n884 0.146333
R5456 VDDA.n888 VDDA.n885 0.146333
R5457 VDDA.n888 VDDA.n826 0.146333
R5458 VDDA.n898 VDDA.n824 0.146333
R5459 VDDA.n904 VDDA.n824 0.146333
R5460 VDDA.n905 VDDA.n904 0.146333
R5461 VDDA.n915 VDDA.n914 0.146333
R5462 VDDA.n918 VDDA.n915 0.146333
R5463 VDDA.n918 VDDA.n820 0.146333
R5464 VDDA.n928 VDDA.n818 0.146333
R5465 VDDA.n934 VDDA.n818 0.146333
R5466 VDDA.n935 VDDA.n934 0.146333
R5467 VDDA.n945 VDDA.n944 0.146333
R5468 VDDA.n948 VDDA.n945 0.146333
R5469 VDDA.n948 VDDA.n814 0.146333
R5470 VDDA.n1954 VDDA.n1953 0.136864
R5471 VDDA.n1965 VDDA.n1535 0.136864
R5472 VDDA.n1984 VDDA.n1983 0.136864
R5473 VDDA.n1995 VDDA.n1529 0.136864
R5474 VDDA.n2014 VDDA.n2013 0.136864
R5475 VDDA.n2025 VDDA.n1523 0.136864
R5476 VDDA.n2044 VDDA.n2043 0.136864
R5477 VDDA.n1952 VDDA.n1538 0.136864
R5478 VDDA.n1969 VDDA.n1968 0.136864
R5479 VDDA.n1982 VDDA.n1532 0.136864
R5480 VDDA.n1999 VDDA.n1998 0.136864
R5481 VDDA.n2012 VDDA.n1526 0.136864
R5482 VDDA.n2029 VDDA.n2028 0.136864
R5483 VDDA.n2042 VDDA.n1520 0.136864
R5484 VDDA.n1610 VDDA.t171 0.1368
R5485 VDDA.n1610 VDDA.t117 0.1368
R5486 VDDA.n1609 VDDA.t380 0.1368
R5487 VDDA.n1609 VDDA.t30 0.1368
R5488 VDDA.n1608 VDDA.t103 0.1368
R5489 VDDA.n1608 VDDA.t49 0.1368
R5490 VDDA.n1607 VDDA.t57 0.1368
R5491 VDDA.n1607 VDDA.t170 0.1368
R5492 VDDA.n1606 VDDA.t75 0.1368
R5493 VDDA.n1606 VDDA.t27 0.1368
R5494 VDDA.n1614 VDDA.n1612 0.135917
R5495 VDDA.n1624 VDDA.n1621 0.135917
R5496 VDDA.n1630 VDDA.n1603 0.135917
R5497 VDDA.n1640 VDDA.n1601 0.135917
R5498 VDDA.n1644 VDDA.n1641 0.135917
R5499 VDDA.n1654 VDDA.n1651 0.135917
R5500 VDDA.n1660 VDDA.n1597 0.135917
R5501 VDDA.n1670 VDDA.n1595 0.135917
R5502 VDDA.n1674 VDDA.n1671 0.135917
R5503 VDDA.n1684 VDDA.n1681 0.135917
R5504 VDDA.n1690 VDDA.n1591 0.135917
R5505 VDDA.n1700 VDDA.n1589 0.135917
R5506 VDDA.n1704 VDDA.n1701 0.135917
R5507 VDDA.n1714 VDDA.n1711 0.135917
R5508 VDDA.n1720 VDDA.n1585 0.135917
R5509 VDDA.n2301 VDDA.n2298 0.135917
R5510 VDDA.n2307 VDDA.n2078 0.135917
R5511 VDDA.n2317 VDDA.n2076 0.135917
R5512 VDDA.n2321 VDDA.n2318 0.135917
R5513 VDDA.n2331 VDDA.n2328 0.135917
R5514 VDDA.n2337 VDDA.n2072 0.135917
R5515 VDDA.n2347 VDDA.n2070 0.135917
R5516 VDDA.n2351 VDDA.n2348 0.135917
R5517 VDDA.n2361 VDDA.n2358 0.135917
R5518 VDDA.n2367 VDDA.n2066 0.135917
R5519 VDDA.n2377 VDDA.n2064 0.135917
R5520 VDDA.n2381 VDDA.n2378 0.135917
R5521 VDDA.n2391 VDDA.n2388 0.135917
R5522 VDDA.n2397 VDDA.n2060 0.135917
R5523 VDDA.n99 VDDA.n96 0.135917
R5524 VDDA.n103 VDDA.n83 0.135917
R5525 VDDA.n111 VDDA.n79 0.135917
R5526 VDDA.n115 VDDA.n112 0.135917
R5527 VDDA.n123 VDDA.n120 0.135917
R5528 VDDA.n127 VDDA.n71 0.135917
R5529 VDDA.n135 VDDA.n67 0.135917
R5530 VDDA.n139 VDDA.n136 0.135917
R5531 VDDA.n147 VDDA.n144 0.135917
R5532 VDDA.n151 VDDA.n59 0.135917
R5533 VDDA.n159 VDDA.n55 0.135917
R5534 VDDA.n163 VDDA.n160 0.135917
R5535 VDDA.n171 VDDA.n168 0.135917
R5536 VDDA.n175 VDDA.n47 0.135917
R5537 VDDA.n2935 VDDA.n45 0.135917
R5538 VDDA.n2817 VDDA.n2802 0.135917
R5539 VDDA.n2823 VDDA.n2800 0.135917
R5540 VDDA.n2833 VDDA.n2796 0.135917
R5541 VDDA.n2837 VDDA.n2794 0.135917
R5542 VDDA.n2847 VDDA.n2790 0.135917
R5543 VDDA.n2853 VDDA.n2788 0.135917
R5544 VDDA.n2863 VDDA.n2784 0.135917
R5545 VDDA.n2867 VDDA.n2782 0.135917
R5546 VDDA.n2877 VDDA.n2778 0.135917
R5547 VDDA.n2883 VDDA.n2776 0.135917
R5548 VDDA.n2893 VDDA.n2772 0.135917
R5549 VDDA.n2897 VDDA.n2770 0.135917
R5550 VDDA.n2907 VDDA.n2766 0.135917
R5551 VDDA.n2913 VDDA.n2764 0.135917
R5552 VDDA.n2922 VDDA.n2760 0.135917
R5553 VDDA.n2666 VDDA.n2652 0.135917
R5554 VDDA.n2670 VDDA.n2667 0.135917
R5555 VDDA.n2678 VDDA.n2675 0.135917
R5556 VDDA.n2682 VDDA.n2644 0.135917
R5557 VDDA.n2690 VDDA.n2640 0.135917
R5558 VDDA.n2694 VDDA.n2691 0.135917
R5559 VDDA.n2702 VDDA.n2699 0.135917
R5560 VDDA.n2706 VDDA.n2632 0.135917
R5561 VDDA.n2714 VDDA.n2628 0.135917
R5562 VDDA.n2718 VDDA.n2715 0.135917
R5563 VDDA.n2726 VDDA.n2723 0.135917
R5564 VDDA.n2730 VDDA.n2620 0.135917
R5565 VDDA.n2738 VDDA.n2616 0.135917
R5566 VDDA.n2742 VDDA.n2739 0.135917
R5567 VDDA.n2751 VDDA.n195 0.135917
R5568 VDDA.n277 VDDA.n274 0.135917
R5569 VDDA.n281 VDDA.n261 0.135917
R5570 VDDA.n289 VDDA.n257 0.135917
R5571 VDDA.n293 VDDA.n290 0.135917
R5572 VDDA.n301 VDDA.n298 0.135917
R5573 VDDA.n305 VDDA.n249 0.135917
R5574 VDDA.n313 VDDA.n245 0.135917
R5575 VDDA.n317 VDDA.n314 0.135917
R5576 VDDA.n325 VDDA.n322 0.135917
R5577 VDDA.n329 VDDA.n237 0.135917
R5578 VDDA.n337 VDDA.n233 0.135917
R5579 VDDA.n341 VDDA.n338 0.135917
R5580 VDDA.n349 VDDA.n346 0.135917
R5581 VDDA.n353 VDDA.n225 0.135917
R5582 VDDA.n2587 VDDA.n223 0.135917
R5583 VDDA.n423 VDDA.n408 0.135917
R5584 VDDA.n429 VDDA.n406 0.135917
R5585 VDDA.n439 VDDA.n402 0.135917
R5586 VDDA.n443 VDDA.n400 0.135917
R5587 VDDA.n453 VDDA.n396 0.135917
R5588 VDDA.n459 VDDA.n394 0.135917
R5589 VDDA.n469 VDDA.n390 0.135917
R5590 VDDA.n473 VDDA.n388 0.135917
R5591 VDDA.n483 VDDA.n384 0.135917
R5592 VDDA.n489 VDDA.n382 0.135917
R5593 VDDA.n499 VDDA.n378 0.135917
R5594 VDDA.n503 VDDA.n376 0.135917
R5595 VDDA.n513 VDDA.n372 0.135917
R5596 VDDA.n519 VDDA.n370 0.135917
R5597 VDDA.n528 VDDA.n366 0.135917
R5598 VDDA.n1386 VDDA.n1372 0.135917
R5599 VDDA.n1390 VDDA.n1387 0.135917
R5600 VDDA.n1398 VDDA.n1395 0.135917
R5601 VDDA.n1402 VDDA.n1364 0.135917
R5602 VDDA.n1410 VDDA.n1360 0.135917
R5603 VDDA.n1414 VDDA.n1411 0.135917
R5604 VDDA.n1422 VDDA.n1419 0.135917
R5605 VDDA.n1426 VDDA.n1352 0.135917
R5606 VDDA.n1434 VDDA.n1348 0.135917
R5607 VDDA.n1438 VDDA.n1435 0.135917
R5608 VDDA.n1446 VDDA.n1443 0.135917
R5609 VDDA.n1450 VDDA.n1340 0.135917
R5610 VDDA.n1458 VDDA.n1336 0.135917
R5611 VDDA.n1462 VDDA.n1459 0.135917
R5612 VDDA.n2408 VDDA.n610 0.135917
R5613 VDDA.n692 VDDA.n689 0.135917
R5614 VDDA.n696 VDDA.n676 0.135917
R5615 VDDA.n704 VDDA.n672 0.135917
R5616 VDDA.n708 VDDA.n705 0.135917
R5617 VDDA.n716 VDDA.n713 0.135917
R5618 VDDA.n720 VDDA.n664 0.135917
R5619 VDDA.n728 VDDA.n660 0.135917
R5620 VDDA.n732 VDDA.n729 0.135917
R5621 VDDA.n740 VDDA.n737 0.135917
R5622 VDDA.n744 VDDA.n652 0.135917
R5623 VDDA.n752 VDDA.n648 0.135917
R5624 VDDA.n756 VDDA.n753 0.135917
R5625 VDDA.n764 VDDA.n761 0.135917
R5626 VDDA.n768 VDDA.n640 0.135917
R5627 VDDA.n1307 VDDA.n638 0.135917
R5628 VDDA.n1189 VDDA.n1174 0.135917
R5629 VDDA.n1195 VDDA.n1172 0.135917
R5630 VDDA.n1205 VDDA.n1168 0.135917
R5631 VDDA.n1209 VDDA.n1166 0.135917
R5632 VDDA.n1219 VDDA.n1162 0.135917
R5633 VDDA.n1225 VDDA.n1160 0.135917
R5634 VDDA.n1235 VDDA.n1156 0.135917
R5635 VDDA.n1239 VDDA.n1154 0.135917
R5636 VDDA.n1249 VDDA.n1150 0.135917
R5637 VDDA.n1255 VDDA.n1148 0.135917
R5638 VDDA.n1265 VDDA.n1144 0.135917
R5639 VDDA.n1269 VDDA.n1142 0.135917
R5640 VDDA.n1279 VDDA.n1138 0.135917
R5641 VDDA.n1285 VDDA.n1136 0.135917
R5642 VDDA.n1294 VDDA.n1132 0.135917
R5643 VDDA.n1038 VDDA.n1024 0.135917
R5644 VDDA.n1042 VDDA.n1039 0.135917
R5645 VDDA.n1050 VDDA.n1047 0.135917
R5646 VDDA.n1054 VDDA.n1016 0.135917
R5647 VDDA.n1062 VDDA.n1012 0.135917
R5648 VDDA.n1066 VDDA.n1063 0.135917
R5649 VDDA.n1074 VDDA.n1071 0.135917
R5650 VDDA.n1078 VDDA.n1004 0.135917
R5651 VDDA.n1086 VDDA.n1000 0.135917
R5652 VDDA.n1090 VDDA.n1087 0.135917
R5653 VDDA.n1098 VDDA.n1095 0.135917
R5654 VDDA.n1102 VDDA.n992 0.135917
R5655 VDDA.n1110 VDDA.n988 0.135917
R5656 VDDA.n1114 VDDA.n1111 0.135917
R5657 VDDA.n1123 VDDA.n787 0.135917
R5658 VDDA.n848 VDDA.n845 0.135917
R5659 VDDA.n854 VDDA.n834 0.135917
R5660 VDDA.n864 VDDA.n832 0.135917
R5661 VDDA.n868 VDDA.n865 0.135917
R5662 VDDA.n878 VDDA.n875 0.135917
R5663 VDDA.n884 VDDA.n828 0.135917
R5664 VDDA.n894 VDDA.n826 0.135917
R5665 VDDA.n898 VDDA.n895 0.135917
R5666 VDDA.n908 VDDA.n905 0.135917
R5667 VDDA.n914 VDDA.n822 0.135917
R5668 VDDA.n924 VDDA.n820 0.135917
R5669 VDDA.n928 VDDA.n925 0.135917
R5670 VDDA.n938 VDDA.n935 0.135917
R5671 VDDA.n944 VDDA.n816 0.135917
R5672 VDDA.n959 VDDA.n814 0.135917
R5673 VDDA.n1624 VDDA.n1603 0.1255
R5674 VDDA.n1641 VDDA.n1640 0.1255
R5675 VDDA.n1654 VDDA.n1597 0.1255
R5676 VDDA.n1671 VDDA.n1670 0.1255
R5677 VDDA.n1684 VDDA.n1591 0.1255
R5678 VDDA.n1701 VDDA.n1700 0.1255
R5679 VDDA.n1714 VDDA.n1585 0.1255
R5680 VDDA.n2284 VDDA.n2283 0.1255
R5681 VDDA.n2283 VDDA.n2282 0.1255
R5682 VDDA.n2157 VDDA.n2100 0.1255
R5683 VDDA.n2104 VDDA.n2100 0.1255
R5684 VDDA.n2106 VDDA.n2104 0.1255
R5685 VDDA.n2108 VDDA.n2106 0.1255
R5686 VDDA.n2110 VDDA.n2108 0.1255
R5687 VDDA.n2112 VDDA.n2110 0.1255
R5688 VDDA.n2114 VDDA.n2112 0.1255
R5689 VDDA.n2116 VDDA.n2114 0.1255
R5690 VDDA.n2118 VDDA.n2116 0.1255
R5691 VDDA.n2148 VDDA.n2118 0.1255
R5692 VDDA.n2147 VDDA.n2120 0.1255
R5693 VDDA.n2124 VDDA.n2120 0.1255
R5694 VDDA.n2126 VDDA.n2124 0.1255
R5695 VDDA.n2128 VDDA.n2126 0.1255
R5696 VDDA.n2130 VDDA.n2128 0.1255
R5697 VDDA.n2132 VDDA.n2130 0.1255
R5698 VDDA.n2134 VDDA.n2132 0.1255
R5699 VDDA.n2136 VDDA.n2134 0.1255
R5700 VDDA.n2138 VDDA.n2136 0.1255
R5701 VDDA.n2301 VDDA.n2078 0.1255
R5702 VDDA.n2318 VDDA.n2317 0.1255
R5703 VDDA.n2331 VDDA.n2072 0.1255
R5704 VDDA.n2348 VDDA.n2347 0.1255
R5705 VDDA.n2361 VDDA.n2066 0.1255
R5706 VDDA.n2378 VDDA.n2377 0.1255
R5707 VDDA.n2391 VDDA.n2060 0.1255
R5708 VDDA.n2462 VDDA.n2456 0.1255
R5709 VDDA.n2475 VDDA.n2470 0.1255
R5710 VDDA.n99 VDDA.n83 0.1255
R5711 VDDA.n112 VDDA.n111 0.1255
R5712 VDDA.n123 VDDA.n71 0.1255
R5713 VDDA.n136 VDDA.n135 0.1255
R5714 VDDA.n147 VDDA.n59 0.1255
R5715 VDDA.n160 VDDA.n159 0.1255
R5716 VDDA.n171 VDDA.n47 0.1255
R5717 VDDA.n2817 VDDA.n2800 0.1255
R5718 VDDA.n2833 VDDA.n2794 0.1255
R5719 VDDA.n2847 VDDA.n2788 0.1255
R5720 VDDA.n2863 VDDA.n2782 0.1255
R5721 VDDA.n2877 VDDA.n2776 0.1255
R5722 VDDA.n2893 VDDA.n2770 0.1255
R5723 VDDA.n2907 VDDA.n2764 0.1255
R5724 VDDA.n2667 VDDA.n2666 0.1255
R5725 VDDA.n2678 VDDA.n2644 0.1255
R5726 VDDA.n2691 VDDA.n2690 0.1255
R5727 VDDA.n2702 VDDA.n2632 0.1255
R5728 VDDA.n2715 VDDA.n2714 0.1255
R5729 VDDA.n2726 VDDA.n2620 0.1255
R5730 VDDA.n2739 VDDA.n2738 0.1255
R5731 VDDA.n277 VDDA.n261 0.1255
R5732 VDDA.n290 VDDA.n289 0.1255
R5733 VDDA.n301 VDDA.n249 0.1255
R5734 VDDA.n314 VDDA.n313 0.1255
R5735 VDDA.n325 VDDA.n237 0.1255
R5736 VDDA.n338 VDDA.n337 0.1255
R5737 VDDA.n349 VDDA.n225 0.1255
R5738 VDDA.n423 VDDA.n406 0.1255
R5739 VDDA.n439 VDDA.n400 0.1255
R5740 VDDA.n453 VDDA.n394 0.1255
R5741 VDDA.n469 VDDA.n388 0.1255
R5742 VDDA.n483 VDDA.n382 0.1255
R5743 VDDA.n499 VDDA.n376 0.1255
R5744 VDDA.n513 VDDA.n370 0.1255
R5745 VDDA.n1387 VDDA.n1386 0.1255
R5746 VDDA.n1398 VDDA.n1364 0.1255
R5747 VDDA.n1411 VDDA.n1410 0.1255
R5748 VDDA.n1422 VDDA.n1352 0.1255
R5749 VDDA.n1435 VDDA.n1434 0.1255
R5750 VDDA.n1446 VDDA.n1340 0.1255
R5751 VDDA.n1459 VDDA.n1458 0.1255
R5752 VDDA.n692 VDDA.n676 0.1255
R5753 VDDA.n705 VDDA.n704 0.1255
R5754 VDDA.n716 VDDA.n664 0.1255
R5755 VDDA.n729 VDDA.n728 0.1255
R5756 VDDA.n740 VDDA.n652 0.1255
R5757 VDDA.n753 VDDA.n752 0.1255
R5758 VDDA.n764 VDDA.n640 0.1255
R5759 VDDA.n1189 VDDA.n1172 0.1255
R5760 VDDA.n1205 VDDA.n1166 0.1255
R5761 VDDA.n1219 VDDA.n1160 0.1255
R5762 VDDA.n1235 VDDA.n1154 0.1255
R5763 VDDA.n1249 VDDA.n1148 0.1255
R5764 VDDA.n1265 VDDA.n1142 0.1255
R5765 VDDA.n1279 VDDA.n1136 0.1255
R5766 VDDA.n1039 VDDA.n1038 0.1255
R5767 VDDA.n1050 VDDA.n1016 0.1255
R5768 VDDA.n1063 VDDA.n1062 0.1255
R5769 VDDA.n1074 VDDA.n1004 0.1255
R5770 VDDA.n1087 VDDA.n1086 0.1255
R5771 VDDA.n1098 VDDA.n992 0.1255
R5772 VDDA.n1111 VDDA.n1110 0.1255
R5773 VDDA.n848 VDDA.n834 0.1255
R5774 VDDA.n865 VDDA.n864 0.1255
R5775 VDDA.n878 VDDA.n828 0.1255
R5776 VDDA.n895 VDDA.n894 0.1255
R5777 VDDA.n908 VDDA.n822 0.1255
R5778 VDDA.n925 VDDA.n924 0.1255
R5779 VDDA.n938 VDDA.n816 0.1255
R5780 VDDA.n1916 VDDA.n1915 0.123287
R5781 VDDA.n1938 VDDA.n1937 0.123287
R5782 VDDA.n2281 VDDA.n2280 0.115083
R5783 VDDA.n2280 VDDA.n2279 0.115083
R5784 VDDA.n2279 VDDA.n2278 0.115083
R5785 VDDA.n2276 VDDA.n2275 0.115083
R5786 VDDA.n2275 VDDA.n2274 0.115083
R5787 VDDA.n2274 VDDA.n2273 0.115083
R5788 VDDA.n2273 VDDA.n2272 0.115083
R5789 VDDA.n2270 VDDA.n2269 0.115083
R5790 VDDA.n2269 VDDA.n2268 0.115083
R5791 VDDA.n577 VDDA.n575 0.115083
R5792 VDDA.n579 VDDA.n577 0.115083
R5793 VDDA.n581 VDDA.n579 0.115083
R5794 VDDA.n583 VDDA.n581 0.115083
R5795 VDDA.n2535 VDDA.n2533 0.115083
R5796 VDDA.n2533 VDDA.n2531 0.115083
R5797 VDDA.n2531 VDDA.n2529 0.115083
R5798 VDDA.n2529 VDDA.n2527 0.115083
R5799 VDDA.n2564 VDDA.n2563 0.115083
R5800 VDDA.n2563 VDDA.n2561 0.115083
R5801 VDDA.n2561 VDDA.n2559 0.115083
R5802 VDDA.n2559 VDDA.n2557 0.115083
R5803 VDDA.n2557 VDDA.n536 0.115083
R5804 VDDA.n2569 VDDA.n536 0.115083
R5805 VDDA.n2429 VDDA.n2428 0.115083
R5806 VDDA.n2428 VDDA.n2426 0.115083
R5807 VDDA.n2426 VDDA.n2424 0.115083
R5808 VDDA.n2424 VDDA.n2422 0.115083
R5809 VDDA.n2422 VDDA.n601 0.115083
R5810 VDDA.n2434 VDDA.n601 0.115083
R5811 VDDA.n2478 VDDA.n2468 0.09425
R5812 VDDA.n2485 VDDA.n2451 0.0838333
R5813 VDDA.n1911 VDDA.n1555 0.076587
R5814 VDDA.n1730 VDDA.n1555 0.076587
R5815 VDDA.n1903 VDDA.n1730 0.076587
R5816 VDDA.n1893 VDDA.n1735 0.076587
R5817 VDDA.n1893 VDDA.n1739 0.076587
R5818 VDDA.n1889 VDDA.n1739 0.076587
R5819 VDDA.n1879 VDDA.n1745 0.076587
R5820 VDDA.n1879 VDDA.n1747 0.076587
R5821 VDDA.n1873 VDDA.n1747 0.076587
R5822 VDDA.n1863 VDDA.n1753 0.076587
R5823 VDDA.n1863 VDDA.n1757 0.076587
R5824 VDDA.n1859 VDDA.n1757 0.076587
R5825 VDDA.n1849 VDDA.n1763 0.076587
R5826 VDDA.n1849 VDDA.n1765 0.076587
R5827 VDDA.n1843 VDDA.n1765 0.076587
R5828 VDDA.n1833 VDDA.n1771 0.076587
R5829 VDDA.n1833 VDDA.n1775 0.076587
R5830 VDDA.n1829 VDDA.n1775 0.076587
R5831 VDDA.n1819 VDDA.n1781 0.076587
R5832 VDDA.n1819 VDDA.n1783 0.076587
R5833 VDDA.n1813 VDDA.n1783 0.076587
R5834 VDDA.n1803 VDDA.n1789 0.076587
R5835 VDDA.n1803 VDDA.n1793 0.076587
R5836 VDDA.n1799 VDDA.n1793 0.076587
R5837 VDDA.n1912 VDDA.n1554 0.076587
R5838 VDDA.n1733 VDDA.n1554 0.076587
R5839 VDDA.n1902 VDDA.n1733 0.076587
R5840 VDDA.n1892 VDDA.n1734 0.076587
R5841 VDDA.n1892 VDDA.n1891 0.076587
R5842 VDDA.n1891 VDDA.n1890 0.076587
R5843 VDDA.n1881 VDDA.n1880 0.076587
R5844 VDDA.n1880 VDDA.n1746 0.076587
R5845 VDDA.n1872 VDDA.n1746 0.076587
R5846 VDDA.n1862 VDDA.n1752 0.076587
R5847 VDDA.n1862 VDDA.n1861 0.076587
R5848 VDDA.n1861 VDDA.n1860 0.076587
R5849 VDDA.n1851 VDDA.n1850 0.076587
R5850 VDDA.n1850 VDDA.n1764 0.076587
R5851 VDDA.n1842 VDDA.n1764 0.076587
R5852 VDDA.n1832 VDDA.n1770 0.076587
R5853 VDDA.n1832 VDDA.n1831 0.076587
R5854 VDDA.n1831 VDDA.n1830 0.076587
R5855 VDDA.n1821 VDDA.n1820 0.076587
R5856 VDDA.n1820 VDDA.n1782 0.076587
R5857 VDDA.n1812 VDDA.n1782 0.076587
R5858 VDDA.n1802 VDDA.n1788 0.076587
R5859 VDDA.n1802 VDDA.n1801 0.076587
R5860 VDDA.n1616 VDDA.n1615 0.0734167
R5861 VDDA.n1617 VDDA.n1616 0.0734167
R5862 VDDA.n1617 VDDA.n1604 0.0734167
R5863 VDDA.n1627 VDDA.n1602 0.0734167
R5864 VDDA.n1635 VDDA.n1602 0.0734167
R5865 VDDA.n1636 VDDA.n1635 0.0734167
R5866 VDDA.n1646 VDDA.n1645 0.0734167
R5867 VDDA.n1647 VDDA.n1646 0.0734167
R5868 VDDA.n1647 VDDA.n1598 0.0734167
R5869 VDDA.n1657 VDDA.n1596 0.0734167
R5870 VDDA.n1665 VDDA.n1596 0.0734167
R5871 VDDA.n1666 VDDA.n1665 0.0734167
R5872 VDDA.n1676 VDDA.n1675 0.0734167
R5873 VDDA.n1677 VDDA.n1676 0.0734167
R5874 VDDA.n1677 VDDA.n1592 0.0734167
R5875 VDDA.n1687 VDDA.n1590 0.0734167
R5876 VDDA.n1695 VDDA.n1590 0.0734167
R5877 VDDA.n1696 VDDA.n1695 0.0734167
R5878 VDDA.n1706 VDDA.n1705 0.0734167
R5879 VDDA.n1707 VDDA.n1706 0.0734167
R5880 VDDA.n1707 VDDA.n1586 0.0734167
R5881 VDDA.n1717 VDDA.n1584 0.0734167
R5882 VDDA.n1725 VDDA.n1584 0.0734167
R5883 VDDA.n2293 VDDA.n2292 0.0734167
R5884 VDDA.n2294 VDDA.n2293 0.0734167
R5885 VDDA.n2294 VDDA.n2079 0.0734167
R5886 VDDA.n2304 VDDA.n2077 0.0734167
R5887 VDDA.n2312 VDDA.n2077 0.0734167
R5888 VDDA.n2313 VDDA.n2312 0.0734167
R5889 VDDA.n2323 VDDA.n2322 0.0734167
R5890 VDDA.n2324 VDDA.n2323 0.0734167
R5891 VDDA.n2324 VDDA.n2073 0.0734167
R5892 VDDA.n2334 VDDA.n2071 0.0734167
R5893 VDDA.n2342 VDDA.n2071 0.0734167
R5894 VDDA.n2343 VDDA.n2342 0.0734167
R5895 VDDA.n2353 VDDA.n2352 0.0734167
R5896 VDDA.n2354 VDDA.n2353 0.0734167
R5897 VDDA.n2354 VDDA.n2067 0.0734167
R5898 VDDA.n2364 VDDA.n2065 0.0734167
R5899 VDDA.n2372 VDDA.n2065 0.0734167
R5900 VDDA.n2373 VDDA.n2372 0.0734167
R5901 VDDA.n2383 VDDA.n2382 0.0734167
R5902 VDDA.n2384 VDDA.n2383 0.0734167
R5903 VDDA.n2384 VDDA.n2061 0.0734167
R5904 VDDA.n2394 VDDA.n2059 0.0734167
R5905 VDDA.n2402 VDDA.n2059 0.0734167
R5906 VDDA.n94 VDDA.n93 0.0734167
R5907 VDDA.n94 VDDA.n86 0.0734167
R5908 VDDA.n102 VDDA.n82 0.0734167
R5909 VDDA.n108 VDDA.n82 0.0734167
R5910 VDDA.n109 VDDA.n108 0.0734167
R5911 VDDA.n117 VDDA.n116 0.0734167
R5912 VDDA.n118 VDDA.n117 0.0734167
R5913 VDDA.n118 VDDA.n74 0.0734167
R5914 VDDA.n126 VDDA.n70 0.0734167
R5915 VDDA.n132 VDDA.n70 0.0734167
R5916 VDDA.n133 VDDA.n132 0.0734167
R5917 VDDA.n141 VDDA.n140 0.0734167
R5918 VDDA.n142 VDDA.n141 0.0734167
R5919 VDDA.n142 VDDA.n62 0.0734167
R5920 VDDA.n150 VDDA.n58 0.0734167
R5921 VDDA.n156 VDDA.n58 0.0734167
R5922 VDDA.n157 VDDA.n156 0.0734167
R5923 VDDA.n165 VDDA.n164 0.0734167
R5924 VDDA.n166 VDDA.n165 0.0734167
R5925 VDDA.n166 VDDA.n50 0.0734167
R5926 VDDA.n174 VDDA.n46 0.0734167
R5927 VDDA.n180 VDDA.n46 0.0734167
R5928 VDDA.n181 VDDA.n180 0.0734167
R5929 VDDA.n2814 VDDA.n2803 0.0734167
R5930 VDDA.n2815 VDDA.n2814 0.0734167
R5931 VDDA.n2825 VDDA.n2824 0.0734167
R5932 VDDA.n2826 VDDA.n2825 0.0734167
R5933 VDDA.n2826 VDDA.n2795 0.0734167
R5934 VDDA.n2836 VDDA.n2791 0.0734167
R5935 VDDA.n2844 VDDA.n2791 0.0734167
R5936 VDDA.n2845 VDDA.n2844 0.0734167
R5937 VDDA.n2855 VDDA.n2854 0.0734167
R5938 VDDA.n2856 VDDA.n2855 0.0734167
R5939 VDDA.n2856 VDDA.n2783 0.0734167
R5940 VDDA.n2866 VDDA.n2779 0.0734167
R5941 VDDA.n2874 VDDA.n2779 0.0734167
R5942 VDDA.n2875 VDDA.n2874 0.0734167
R5943 VDDA.n2885 VDDA.n2884 0.0734167
R5944 VDDA.n2886 VDDA.n2885 0.0734167
R5945 VDDA.n2886 VDDA.n2771 0.0734167
R5946 VDDA.n2896 VDDA.n2767 0.0734167
R5947 VDDA.n2904 VDDA.n2767 0.0734167
R5948 VDDA.n2905 VDDA.n2904 0.0734167
R5949 VDDA.n2915 VDDA.n2914 0.0734167
R5950 VDDA.n2916 VDDA.n2915 0.0734167
R5951 VDDA.n2916 VDDA.n2759 0.0734167
R5952 VDDA.n2663 VDDA.n2655 0.0734167
R5953 VDDA.n2664 VDDA.n2663 0.0734167
R5954 VDDA.n2672 VDDA.n2671 0.0734167
R5955 VDDA.n2673 VDDA.n2672 0.0734167
R5956 VDDA.n2673 VDDA.n2647 0.0734167
R5957 VDDA.n2681 VDDA.n2643 0.0734167
R5958 VDDA.n2687 VDDA.n2643 0.0734167
R5959 VDDA.n2688 VDDA.n2687 0.0734167
R5960 VDDA.n2696 VDDA.n2695 0.0734167
R5961 VDDA.n2697 VDDA.n2696 0.0734167
R5962 VDDA.n2697 VDDA.n2635 0.0734167
R5963 VDDA.n2705 VDDA.n2631 0.0734167
R5964 VDDA.n2711 VDDA.n2631 0.0734167
R5965 VDDA.n2712 VDDA.n2711 0.0734167
R5966 VDDA.n2720 VDDA.n2719 0.0734167
R5967 VDDA.n2721 VDDA.n2720 0.0734167
R5968 VDDA.n2721 VDDA.n2623 0.0734167
R5969 VDDA.n2729 VDDA.n2619 0.0734167
R5970 VDDA.n2735 VDDA.n2619 0.0734167
R5971 VDDA.n2736 VDDA.n2735 0.0734167
R5972 VDDA.n2744 VDDA.n2743 0.0734167
R5973 VDDA.n2745 VDDA.n2744 0.0734167
R5974 VDDA.n2745 VDDA.n194 0.0734167
R5975 VDDA.n272 VDDA.n271 0.0734167
R5976 VDDA.n272 VDDA.n264 0.0734167
R5977 VDDA.n280 VDDA.n260 0.0734167
R5978 VDDA.n286 VDDA.n260 0.0734167
R5979 VDDA.n287 VDDA.n286 0.0734167
R5980 VDDA.n295 VDDA.n294 0.0734167
R5981 VDDA.n296 VDDA.n295 0.0734167
R5982 VDDA.n296 VDDA.n252 0.0734167
R5983 VDDA.n304 VDDA.n248 0.0734167
R5984 VDDA.n310 VDDA.n248 0.0734167
R5985 VDDA.n311 VDDA.n310 0.0734167
R5986 VDDA.n319 VDDA.n318 0.0734167
R5987 VDDA.n320 VDDA.n319 0.0734167
R5988 VDDA.n320 VDDA.n240 0.0734167
R5989 VDDA.n328 VDDA.n236 0.0734167
R5990 VDDA.n334 VDDA.n236 0.0734167
R5991 VDDA.n335 VDDA.n334 0.0734167
R5992 VDDA.n343 VDDA.n342 0.0734167
R5993 VDDA.n344 VDDA.n343 0.0734167
R5994 VDDA.n344 VDDA.n228 0.0734167
R5995 VDDA.n352 VDDA.n224 0.0734167
R5996 VDDA.n358 VDDA.n224 0.0734167
R5997 VDDA.n359 VDDA.n358 0.0734167
R5998 VDDA.n420 VDDA.n409 0.0734167
R5999 VDDA.n421 VDDA.n420 0.0734167
R6000 VDDA.n431 VDDA.n430 0.0734167
R6001 VDDA.n432 VDDA.n431 0.0734167
R6002 VDDA.n432 VDDA.n401 0.0734167
R6003 VDDA.n442 VDDA.n397 0.0734167
R6004 VDDA.n450 VDDA.n397 0.0734167
R6005 VDDA.n451 VDDA.n450 0.0734167
R6006 VDDA.n461 VDDA.n460 0.0734167
R6007 VDDA.n462 VDDA.n461 0.0734167
R6008 VDDA.n462 VDDA.n389 0.0734167
R6009 VDDA.n472 VDDA.n385 0.0734167
R6010 VDDA.n480 VDDA.n385 0.0734167
R6011 VDDA.n481 VDDA.n480 0.0734167
R6012 VDDA.n491 VDDA.n490 0.0734167
R6013 VDDA.n492 VDDA.n491 0.0734167
R6014 VDDA.n492 VDDA.n377 0.0734167
R6015 VDDA.n502 VDDA.n373 0.0734167
R6016 VDDA.n510 VDDA.n373 0.0734167
R6017 VDDA.n511 VDDA.n510 0.0734167
R6018 VDDA.n521 VDDA.n520 0.0734167
R6019 VDDA.n522 VDDA.n521 0.0734167
R6020 VDDA.n522 VDDA.n365 0.0734167
R6021 VDDA.n1383 VDDA.n1375 0.0734167
R6022 VDDA.n1384 VDDA.n1383 0.0734167
R6023 VDDA.n1392 VDDA.n1391 0.0734167
R6024 VDDA.n1393 VDDA.n1392 0.0734167
R6025 VDDA.n1393 VDDA.n1367 0.0734167
R6026 VDDA.n1401 VDDA.n1363 0.0734167
R6027 VDDA.n1407 VDDA.n1363 0.0734167
R6028 VDDA.n1408 VDDA.n1407 0.0734167
R6029 VDDA.n1416 VDDA.n1415 0.0734167
R6030 VDDA.n1417 VDDA.n1416 0.0734167
R6031 VDDA.n1417 VDDA.n1355 0.0734167
R6032 VDDA.n1425 VDDA.n1351 0.0734167
R6033 VDDA.n1431 VDDA.n1351 0.0734167
R6034 VDDA.n1432 VDDA.n1431 0.0734167
R6035 VDDA.n1440 VDDA.n1439 0.0734167
R6036 VDDA.n1441 VDDA.n1440 0.0734167
R6037 VDDA.n1441 VDDA.n1343 0.0734167
R6038 VDDA.n1449 VDDA.n1339 0.0734167
R6039 VDDA.n1455 VDDA.n1339 0.0734167
R6040 VDDA.n1456 VDDA.n1455 0.0734167
R6041 VDDA.n1464 VDDA.n1463 0.0734167
R6042 VDDA.n1465 VDDA.n1464 0.0734167
R6043 VDDA.n1465 VDDA.n609 0.0734167
R6044 VDDA.n687 VDDA.n686 0.0734167
R6045 VDDA.n687 VDDA.n679 0.0734167
R6046 VDDA.n695 VDDA.n675 0.0734167
R6047 VDDA.n701 VDDA.n675 0.0734167
R6048 VDDA.n702 VDDA.n701 0.0734167
R6049 VDDA.n710 VDDA.n709 0.0734167
R6050 VDDA.n711 VDDA.n710 0.0734167
R6051 VDDA.n711 VDDA.n667 0.0734167
R6052 VDDA.n719 VDDA.n663 0.0734167
R6053 VDDA.n725 VDDA.n663 0.0734167
R6054 VDDA.n726 VDDA.n725 0.0734167
R6055 VDDA.n734 VDDA.n733 0.0734167
R6056 VDDA.n735 VDDA.n734 0.0734167
R6057 VDDA.n735 VDDA.n655 0.0734167
R6058 VDDA.n743 VDDA.n651 0.0734167
R6059 VDDA.n749 VDDA.n651 0.0734167
R6060 VDDA.n750 VDDA.n749 0.0734167
R6061 VDDA.n758 VDDA.n757 0.0734167
R6062 VDDA.n759 VDDA.n758 0.0734167
R6063 VDDA.n759 VDDA.n643 0.0734167
R6064 VDDA.n767 VDDA.n639 0.0734167
R6065 VDDA.n773 VDDA.n639 0.0734167
R6066 VDDA.n774 VDDA.n773 0.0734167
R6067 VDDA.n1186 VDDA.n1175 0.0734167
R6068 VDDA.n1187 VDDA.n1186 0.0734167
R6069 VDDA.n1197 VDDA.n1196 0.0734167
R6070 VDDA.n1198 VDDA.n1197 0.0734167
R6071 VDDA.n1198 VDDA.n1167 0.0734167
R6072 VDDA.n1208 VDDA.n1163 0.0734167
R6073 VDDA.n1216 VDDA.n1163 0.0734167
R6074 VDDA.n1217 VDDA.n1216 0.0734167
R6075 VDDA.n1227 VDDA.n1226 0.0734167
R6076 VDDA.n1228 VDDA.n1227 0.0734167
R6077 VDDA.n1228 VDDA.n1155 0.0734167
R6078 VDDA.n1238 VDDA.n1151 0.0734167
R6079 VDDA.n1246 VDDA.n1151 0.0734167
R6080 VDDA.n1247 VDDA.n1246 0.0734167
R6081 VDDA.n1257 VDDA.n1256 0.0734167
R6082 VDDA.n1258 VDDA.n1257 0.0734167
R6083 VDDA.n1258 VDDA.n1143 0.0734167
R6084 VDDA.n1268 VDDA.n1139 0.0734167
R6085 VDDA.n1276 VDDA.n1139 0.0734167
R6086 VDDA.n1277 VDDA.n1276 0.0734167
R6087 VDDA.n1287 VDDA.n1286 0.0734167
R6088 VDDA.n1288 VDDA.n1287 0.0734167
R6089 VDDA.n1288 VDDA.n1131 0.0734167
R6090 VDDA.n1035 VDDA.n1027 0.0734167
R6091 VDDA.n1036 VDDA.n1035 0.0734167
R6092 VDDA.n1044 VDDA.n1043 0.0734167
R6093 VDDA.n1045 VDDA.n1044 0.0734167
R6094 VDDA.n1045 VDDA.n1019 0.0734167
R6095 VDDA.n1053 VDDA.n1015 0.0734167
R6096 VDDA.n1059 VDDA.n1015 0.0734167
R6097 VDDA.n1060 VDDA.n1059 0.0734167
R6098 VDDA.n1068 VDDA.n1067 0.0734167
R6099 VDDA.n1069 VDDA.n1068 0.0734167
R6100 VDDA.n1069 VDDA.n1007 0.0734167
R6101 VDDA.n1077 VDDA.n1003 0.0734167
R6102 VDDA.n1083 VDDA.n1003 0.0734167
R6103 VDDA.n1084 VDDA.n1083 0.0734167
R6104 VDDA.n1092 VDDA.n1091 0.0734167
R6105 VDDA.n1093 VDDA.n1092 0.0734167
R6106 VDDA.n1093 VDDA.n995 0.0734167
R6107 VDDA.n1101 VDDA.n991 0.0734167
R6108 VDDA.n1107 VDDA.n991 0.0734167
R6109 VDDA.n1108 VDDA.n1107 0.0734167
R6110 VDDA.n1116 VDDA.n1115 0.0734167
R6111 VDDA.n1117 VDDA.n1116 0.0734167
R6112 VDDA.n1117 VDDA.n786 0.0734167
R6113 VDDA.n841 VDDA.n840 0.0734167
R6114 VDDA.n841 VDDA.n835 0.0734167
R6115 VDDA.n851 VDDA.n833 0.0734167
R6116 VDDA.n859 VDDA.n833 0.0734167
R6117 VDDA.n860 VDDA.n859 0.0734167
R6118 VDDA.n870 VDDA.n869 0.0734167
R6119 VDDA.n871 VDDA.n870 0.0734167
R6120 VDDA.n871 VDDA.n829 0.0734167
R6121 VDDA.n881 VDDA.n827 0.0734167
R6122 VDDA.n889 VDDA.n827 0.0734167
R6123 VDDA.n890 VDDA.n889 0.0734167
R6124 VDDA.n900 VDDA.n899 0.0734167
R6125 VDDA.n901 VDDA.n900 0.0734167
R6126 VDDA.n901 VDDA.n823 0.0734167
R6127 VDDA.n911 VDDA.n821 0.0734167
R6128 VDDA.n919 VDDA.n821 0.0734167
R6129 VDDA.n920 VDDA.n919 0.0734167
R6130 VDDA.n930 VDDA.n929 0.0734167
R6131 VDDA.n931 VDDA.n930 0.0734167
R6132 VDDA.n931 VDDA.n817 0.0734167
R6133 VDDA.n941 VDDA.n815 0.0734167
R6134 VDDA.n949 VDDA.n815 0.0734167
R6135 VDDA.n950 VDDA.n949 0.0734167
R6136 VDDA.n2054 VDDA.n1518 0.0725159
R6137 VDDA.n1911 VDDA.n1553 0.0711522
R6138 VDDA.n1903 VDDA.n1732 0.0711522
R6139 VDDA.n1899 VDDA.n1735 0.0711522
R6140 VDDA.n1889 VDDA.n1741 0.0711522
R6141 VDDA.n1883 VDDA.n1745 0.0711522
R6142 VDDA.n1873 VDDA.n1751 0.0711522
R6143 VDDA.n1869 VDDA.n1753 0.0711522
R6144 VDDA.n1859 VDDA.n1759 0.0711522
R6145 VDDA.n1853 VDDA.n1763 0.0711522
R6146 VDDA.n1843 VDDA.n1769 0.0711522
R6147 VDDA.n1839 VDDA.n1771 0.0711522
R6148 VDDA.n1829 VDDA.n1777 0.0711522
R6149 VDDA.n1823 VDDA.n1781 0.0711522
R6150 VDDA.n1813 VDDA.n1787 0.0711522
R6151 VDDA.n1809 VDDA.n1789 0.0711522
R6152 VDDA.n1913 VDDA.n1912 0.0711522
R6153 VDDA.n1902 VDDA.n1901 0.0711522
R6154 VDDA.n1900 VDDA.n1734 0.0711522
R6155 VDDA.n1890 VDDA.n1740 0.0711522
R6156 VDDA.n1882 VDDA.n1881 0.0711522
R6157 VDDA.n1872 VDDA.n1871 0.0711522
R6158 VDDA.n1870 VDDA.n1752 0.0711522
R6159 VDDA.n1860 VDDA.n1758 0.0711522
R6160 VDDA.n1852 VDDA.n1851 0.0711522
R6161 VDDA.n1842 VDDA.n1841 0.0711522
R6162 VDDA.n1840 VDDA.n1770 0.0711522
R6163 VDDA.n1830 VDDA.n1776 0.0711522
R6164 VDDA.n1822 VDDA.n1821 0.0711522
R6165 VDDA.n1812 VDDA.n1811 0.0711522
R6166 VDDA.n1810 VDDA.n1788 0.0711522
R6167 VDDA.n1615 VDDA.n1611 0.0682083
R6168 VDDA.n1625 VDDA.n1604 0.0682083
R6169 VDDA.n1627 VDDA.n1626 0.0682083
R6170 VDDA.n1637 VDDA.n1636 0.0682083
R6171 VDDA.n1645 VDDA.n1600 0.0682083
R6172 VDDA.n1655 VDDA.n1598 0.0682083
R6173 VDDA.n1657 VDDA.n1656 0.0682083
R6174 VDDA.n1667 VDDA.n1666 0.0682083
R6175 VDDA.n1675 VDDA.n1594 0.0682083
R6176 VDDA.n1685 VDDA.n1592 0.0682083
R6177 VDDA.n1687 VDDA.n1686 0.0682083
R6178 VDDA.n1697 VDDA.n1696 0.0682083
R6179 VDDA.n1705 VDDA.n1588 0.0682083
R6180 VDDA.n1715 VDDA.n1586 0.0682083
R6181 VDDA.n1717 VDDA.n1716 0.0682083
R6182 VDDA.n2277 VDDA.n2276 0.0682083
R6183 VDDA.n2272 VDDA.n2271 0.0682083
R6184 VDDA.n2302 VDDA.n2079 0.0682083
R6185 VDDA.n2304 VDDA.n2303 0.0682083
R6186 VDDA.n2314 VDDA.n2313 0.0682083
R6187 VDDA.n2322 VDDA.n2075 0.0682083
R6188 VDDA.n2332 VDDA.n2073 0.0682083
R6189 VDDA.n2334 VDDA.n2333 0.0682083
R6190 VDDA.n2344 VDDA.n2343 0.0682083
R6191 VDDA.n2352 VDDA.n2069 0.0682083
R6192 VDDA.n2362 VDDA.n2067 0.0682083
R6193 VDDA.n2364 VDDA.n2363 0.0682083
R6194 VDDA.n2374 VDDA.n2373 0.0682083
R6195 VDDA.n2382 VDDA.n2063 0.0682083
R6196 VDDA.n2392 VDDA.n2061 0.0682083
R6197 VDDA.n2394 VDDA.n2393 0.0682083
R6198 VDDA.n100 VDDA.n86 0.0682083
R6199 VDDA.n102 VDDA.n101 0.0682083
R6200 VDDA.n110 VDDA.n109 0.0682083
R6201 VDDA.n116 VDDA.n78 0.0682083
R6202 VDDA.n124 VDDA.n74 0.0682083
R6203 VDDA.n126 VDDA.n125 0.0682083
R6204 VDDA.n134 VDDA.n133 0.0682083
R6205 VDDA.n140 VDDA.n66 0.0682083
R6206 VDDA.n148 VDDA.n62 0.0682083
R6207 VDDA.n150 VDDA.n149 0.0682083
R6208 VDDA.n158 VDDA.n157 0.0682083
R6209 VDDA.n164 VDDA.n54 0.0682083
R6210 VDDA.n172 VDDA.n50 0.0682083
R6211 VDDA.n174 VDDA.n173 0.0682083
R6212 VDDA.n2934 VDDA.n181 0.0682083
R6213 VDDA.n2816 VDDA.n2815 0.0682083
R6214 VDDA.n2824 VDDA.n2799 0.0682083
R6215 VDDA.n2834 VDDA.n2795 0.0682083
R6216 VDDA.n2836 VDDA.n2835 0.0682083
R6217 VDDA.n2846 VDDA.n2845 0.0682083
R6218 VDDA.n2854 VDDA.n2787 0.0682083
R6219 VDDA.n2864 VDDA.n2783 0.0682083
R6220 VDDA.n2866 VDDA.n2865 0.0682083
R6221 VDDA.n2876 VDDA.n2875 0.0682083
R6222 VDDA.n2884 VDDA.n2775 0.0682083
R6223 VDDA.n2894 VDDA.n2771 0.0682083
R6224 VDDA.n2896 VDDA.n2895 0.0682083
R6225 VDDA.n2906 VDDA.n2905 0.0682083
R6226 VDDA.n2914 VDDA.n2763 0.0682083
R6227 VDDA.n2923 VDDA.n2759 0.0682083
R6228 VDDA.n2665 VDDA.n2664 0.0682083
R6229 VDDA.n2671 VDDA.n2651 0.0682083
R6230 VDDA.n2679 VDDA.n2647 0.0682083
R6231 VDDA.n2681 VDDA.n2680 0.0682083
R6232 VDDA.n2689 VDDA.n2688 0.0682083
R6233 VDDA.n2695 VDDA.n2639 0.0682083
R6234 VDDA.n2703 VDDA.n2635 0.0682083
R6235 VDDA.n2705 VDDA.n2704 0.0682083
R6236 VDDA.n2713 VDDA.n2712 0.0682083
R6237 VDDA.n2719 VDDA.n2627 0.0682083
R6238 VDDA.n2727 VDDA.n2623 0.0682083
R6239 VDDA.n2729 VDDA.n2728 0.0682083
R6240 VDDA.n2737 VDDA.n2736 0.0682083
R6241 VDDA.n2743 VDDA.n2615 0.0682083
R6242 VDDA.n2752 VDDA.n194 0.0682083
R6243 VDDA.n278 VDDA.n264 0.0682083
R6244 VDDA.n280 VDDA.n279 0.0682083
R6245 VDDA.n288 VDDA.n287 0.0682083
R6246 VDDA.n294 VDDA.n256 0.0682083
R6247 VDDA.n302 VDDA.n252 0.0682083
R6248 VDDA.n304 VDDA.n303 0.0682083
R6249 VDDA.n312 VDDA.n311 0.0682083
R6250 VDDA.n318 VDDA.n244 0.0682083
R6251 VDDA.n326 VDDA.n240 0.0682083
R6252 VDDA.n328 VDDA.n327 0.0682083
R6253 VDDA.n336 VDDA.n335 0.0682083
R6254 VDDA.n342 VDDA.n232 0.0682083
R6255 VDDA.n350 VDDA.n228 0.0682083
R6256 VDDA.n352 VDDA.n351 0.0682083
R6257 VDDA.n2586 VDDA.n359 0.0682083
R6258 VDDA.n422 VDDA.n421 0.0682083
R6259 VDDA.n430 VDDA.n405 0.0682083
R6260 VDDA.n440 VDDA.n401 0.0682083
R6261 VDDA.n442 VDDA.n441 0.0682083
R6262 VDDA.n452 VDDA.n451 0.0682083
R6263 VDDA.n460 VDDA.n393 0.0682083
R6264 VDDA.n470 VDDA.n389 0.0682083
R6265 VDDA.n472 VDDA.n471 0.0682083
R6266 VDDA.n482 VDDA.n481 0.0682083
R6267 VDDA.n490 VDDA.n381 0.0682083
R6268 VDDA.n500 VDDA.n377 0.0682083
R6269 VDDA.n502 VDDA.n501 0.0682083
R6270 VDDA.n512 VDDA.n511 0.0682083
R6271 VDDA.n520 VDDA.n369 0.0682083
R6272 VDDA.n529 VDDA.n365 0.0682083
R6273 VDDA.n1385 VDDA.n1384 0.0682083
R6274 VDDA.n1391 VDDA.n1371 0.0682083
R6275 VDDA.n1399 VDDA.n1367 0.0682083
R6276 VDDA.n1401 VDDA.n1400 0.0682083
R6277 VDDA.n1409 VDDA.n1408 0.0682083
R6278 VDDA.n1415 VDDA.n1359 0.0682083
R6279 VDDA.n1423 VDDA.n1355 0.0682083
R6280 VDDA.n1425 VDDA.n1424 0.0682083
R6281 VDDA.n1433 VDDA.n1432 0.0682083
R6282 VDDA.n1439 VDDA.n1347 0.0682083
R6283 VDDA.n1447 VDDA.n1343 0.0682083
R6284 VDDA.n1449 VDDA.n1448 0.0682083
R6285 VDDA.n1457 VDDA.n1456 0.0682083
R6286 VDDA.n1463 VDDA.n1335 0.0682083
R6287 VDDA.n2409 VDDA.n609 0.0682083
R6288 VDDA.n693 VDDA.n679 0.0682083
R6289 VDDA.n695 VDDA.n694 0.0682083
R6290 VDDA.n703 VDDA.n702 0.0682083
R6291 VDDA.n709 VDDA.n671 0.0682083
R6292 VDDA.n717 VDDA.n667 0.0682083
R6293 VDDA.n719 VDDA.n718 0.0682083
R6294 VDDA.n727 VDDA.n726 0.0682083
R6295 VDDA.n733 VDDA.n659 0.0682083
R6296 VDDA.n741 VDDA.n655 0.0682083
R6297 VDDA.n743 VDDA.n742 0.0682083
R6298 VDDA.n751 VDDA.n750 0.0682083
R6299 VDDA.n757 VDDA.n647 0.0682083
R6300 VDDA.n765 VDDA.n643 0.0682083
R6301 VDDA.n767 VDDA.n766 0.0682083
R6302 VDDA.n1306 VDDA.n774 0.0682083
R6303 VDDA.n1188 VDDA.n1187 0.0682083
R6304 VDDA.n1196 VDDA.n1171 0.0682083
R6305 VDDA.n1206 VDDA.n1167 0.0682083
R6306 VDDA.n1208 VDDA.n1207 0.0682083
R6307 VDDA.n1218 VDDA.n1217 0.0682083
R6308 VDDA.n1226 VDDA.n1159 0.0682083
R6309 VDDA.n1236 VDDA.n1155 0.0682083
R6310 VDDA.n1238 VDDA.n1237 0.0682083
R6311 VDDA.n1248 VDDA.n1247 0.0682083
R6312 VDDA.n1256 VDDA.n1147 0.0682083
R6313 VDDA.n1266 VDDA.n1143 0.0682083
R6314 VDDA.n1268 VDDA.n1267 0.0682083
R6315 VDDA.n1278 VDDA.n1277 0.0682083
R6316 VDDA.n1286 VDDA.n1135 0.0682083
R6317 VDDA.n1295 VDDA.n1131 0.0682083
R6318 VDDA.n1037 VDDA.n1036 0.0682083
R6319 VDDA.n1043 VDDA.n1023 0.0682083
R6320 VDDA.n1051 VDDA.n1019 0.0682083
R6321 VDDA.n1053 VDDA.n1052 0.0682083
R6322 VDDA.n1061 VDDA.n1060 0.0682083
R6323 VDDA.n1067 VDDA.n1011 0.0682083
R6324 VDDA.n1075 VDDA.n1007 0.0682083
R6325 VDDA.n1077 VDDA.n1076 0.0682083
R6326 VDDA.n1085 VDDA.n1084 0.0682083
R6327 VDDA.n1091 VDDA.n999 0.0682083
R6328 VDDA.n1099 VDDA.n995 0.0682083
R6329 VDDA.n1101 VDDA.n1100 0.0682083
R6330 VDDA.n1109 VDDA.n1108 0.0682083
R6331 VDDA.n1115 VDDA.n987 0.0682083
R6332 VDDA.n1124 VDDA.n786 0.0682083
R6333 VDDA.n849 VDDA.n835 0.0682083
R6334 VDDA.n851 VDDA.n850 0.0682083
R6335 VDDA.n861 VDDA.n860 0.0682083
R6336 VDDA.n869 VDDA.n831 0.0682083
R6337 VDDA.n879 VDDA.n829 0.0682083
R6338 VDDA.n881 VDDA.n880 0.0682083
R6339 VDDA.n891 VDDA.n890 0.0682083
R6340 VDDA.n899 VDDA.n825 0.0682083
R6341 VDDA.n909 VDDA.n823 0.0682083
R6342 VDDA.n911 VDDA.n910 0.0682083
R6343 VDDA.n921 VDDA.n920 0.0682083
R6344 VDDA.n929 VDDA.n819 0.0682083
R6345 VDDA.n939 VDDA.n817 0.0682083
R6346 VDDA.n941 VDDA.n940 0.0682083
R6347 VDDA.n958 VDDA.n950 0.0682083
R6348 VDDA.n92 VDDA.n91 0.0672139
R6349 VDDA.n2807 VDDA.n2806 0.0672139
R6350 VDDA.n2658 VDDA.n2656 0.0672139
R6351 VDDA.n270 VDDA.n269 0.0672139
R6352 VDDA.n413 VDDA.n412 0.0672139
R6353 VDDA.n1378 VDDA.n1376 0.0672139
R6354 VDDA.n685 VDDA.n684 0.0672139
R6355 VDDA.n1179 VDDA.n1178 0.0672139
R6356 VDDA.n1030 VDDA.n1028 0.0672139
R6357 VDDA.n1726 VDDA.n1583 0.0672139
R6358 VDDA.n2403 VDDA.n2058 0.0672139
R6359 VDDA.n839 VDDA.n838 0.0672139
R6360 VDDA.n1899 VDDA.n1732 0.0657174
R6361 VDDA.n1883 VDDA.n1741 0.0657174
R6362 VDDA.n1869 VDDA.n1751 0.0657174
R6363 VDDA.n1853 VDDA.n1759 0.0657174
R6364 VDDA.n1839 VDDA.n1769 0.0657174
R6365 VDDA.n1823 VDDA.n1777 0.0657174
R6366 VDDA.n1809 VDDA.n1787 0.0657174
R6367 VDDA.n1901 VDDA.n1900 0.0657174
R6368 VDDA.n1882 VDDA.n1740 0.0657174
R6369 VDDA.n1871 VDDA.n1870 0.0657174
R6370 VDDA.n1852 VDDA.n1758 0.0657174
R6371 VDDA.n1841 VDDA.n1840 0.0657174
R6372 VDDA.n1822 VDDA.n1776 0.0657174
R6373 VDDA.n1811 VDDA.n1810 0.0657174
R6374 VDDA.n1626 VDDA.n1625 0.063
R6375 VDDA.n1637 VDDA.n1600 0.063
R6376 VDDA.n1656 VDDA.n1655 0.063
R6377 VDDA.n1667 VDDA.n1594 0.063
R6378 VDDA.n1686 VDDA.n1685 0.063
R6379 VDDA.n1697 VDDA.n1588 0.063
R6380 VDDA.n1716 VDDA.n1715 0.063
R6381 VDDA.n2303 VDDA.n2302 0.063
R6382 VDDA.n2314 VDDA.n2075 0.063
R6383 VDDA.n2333 VDDA.n2332 0.063
R6384 VDDA.n2344 VDDA.n2069 0.063
R6385 VDDA.n2363 VDDA.n2362 0.063
R6386 VDDA.n2374 VDDA.n2063 0.063
R6387 VDDA.n2393 VDDA.n2392 0.063
R6388 VDDA.n101 VDDA.n100 0.063
R6389 VDDA.n110 VDDA.n78 0.063
R6390 VDDA.n125 VDDA.n124 0.063
R6391 VDDA.n134 VDDA.n66 0.063
R6392 VDDA.n149 VDDA.n148 0.063
R6393 VDDA.n158 VDDA.n54 0.063
R6394 VDDA.n173 VDDA.n172 0.063
R6395 VDDA.n2816 VDDA.n2799 0.063
R6396 VDDA.n2835 VDDA.n2834 0.063
R6397 VDDA.n2846 VDDA.n2787 0.063
R6398 VDDA.n2865 VDDA.n2864 0.063
R6399 VDDA.n2876 VDDA.n2775 0.063
R6400 VDDA.n2895 VDDA.n2894 0.063
R6401 VDDA.n2906 VDDA.n2763 0.063
R6402 VDDA.n2665 VDDA.n2651 0.063
R6403 VDDA.n2680 VDDA.n2679 0.063
R6404 VDDA.n2689 VDDA.n2639 0.063
R6405 VDDA.n2704 VDDA.n2703 0.063
R6406 VDDA.n2713 VDDA.n2627 0.063
R6407 VDDA.n2728 VDDA.n2727 0.063
R6408 VDDA.n2737 VDDA.n2615 0.063
R6409 VDDA.n279 VDDA.n278 0.063
R6410 VDDA.n288 VDDA.n256 0.063
R6411 VDDA.n303 VDDA.n302 0.063
R6412 VDDA.n312 VDDA.n244 0.063
R6413 VDDA.n327 VDDA.n326 0.063
R6414 VDDA.n336 VDDA.n232 0.063
R6415 VDDA.n351 VDDA.n350 0.063
R6416 VDDA.n422 VDDA.n405 0.063
R6417 VDDA.n441 VDDA.n440 0.063
R6418 VDDA.n452 VDDA.n393 0.063
R6419 VDDA.n471 VDDA.n470 0.063
R6420 VDDA.n482 VDDA.n381 0.063
R6421 VDDA.n501 VDDA.n500 0.063
R6422 VDDA.n512 VDDA.n369 0.063
R6423 VDDA.n1385 VDDA.n1371 0.063
R6424 VDDA.n1400 VDDA.n1399 0.063
R6425 VDDA.n1409 VDDA.n1359 0.063
R6426 VDDA.n1424 VDDA.n1423 0.063
R6427 VDDA.n1433 VDDA.n1347 0.063
R6428 VDDA.n1448 VDDA.n1447 0.063
R6429 VDDA.n1457 VDDA.n1335 0.063
R6430 VDDA.n694 VDDA.n693 0.063
R6431 VDDA.n703 VDDA.n671 0.063
R6432 VDDA.n718 VDDA.n717 0.063
R6433 VDDA.n727 VDDA.n659 0.063
R6434 VDDA.n742 VDDA.n741 0.063
R6435 VDDA.n751 VDDA.n647 0.063
R6436 VDDA.n766 VDDA.n765 0.063
R6437 VDDA.n1188 VDDA.n1171 0.063
R6438 VDDA.n1207 VDDA.n1206 0.063
R6439 VDDA.n1218 VDDA.n1159 0.063
R6440 VDDA.n1237 VDDA.n1236 0.063
R6441 VDDA.n1248 VDDA.n1147 0.063
R6442 VDDA.n1267 VDDA.n1266 0.063
R6443 VDDA.n1278 VDDA.n1135 0.063
R6444 VDDA.n1037 VDDA.n1023 0.063
R6445 VDDA.n1052 VDDA.n1051 0.063
R6446 VDDA.n1061 VDDA.n1011 0.063
R6447 VDDA.n1076 VDDA.n1075 0.063
R6448 VDDA.n1085 VDDA.n999 0.063
R6449 VDDA.n1100 VDDA.n1099 0.063
R6450 VDDA.n1109 VDDA.n987 0.063
R6451 VDDA.n850 VDDA.n849 0.063
R6452 VDDA.n861 VDDA.n831 0.063
R6453 VDDA.n880 VDDA.n879 0.063
R6454 VDDA.n891 VDDA.n825 0.063
R6455 VDDA.n910 VDDA.n909 0.063
R6456 VDDA.n921 VDDA.n819 0.063
R6457 VDDA.n940 VDDA.n939 0.063
R6458 VDDA.n1947 VDDA.n1946 0.0603182
R6459 VDDA.n1961 VDDA.n1960 0.0603182
R6460 VDDA.n1977 VDDA.n1976 0.0603182
R6461 VDDA.n1991 VDDA.n1990 0.0603182
R6462 VDDA.n2007 VDDA.n2006 0.0603182
R6463 VDDA.n2021 VDDA.n2020 0.0603182
R6464 VDDA.n2037 VDDA.n2036 0.0603182
R6465 VDDA.n2051 VDDA.n2050 0.0603182
R6466 VDDA.n1941 VDDA.n1492 0.0560455
R6467 VDDA.n1951 VDDA.n1950 0.0560455
R6468 VDDA.n1957 VDDA.n1956 0.0560455
R6469 VDDA.n1967 VDDA.n1966 0.0560455
R6470 VDDA.n1971 VDDA.n1970 0.0560455
R6471 VDDA.n1981 VDDA.n1980 0.0560455
R6472 VDDA.n1987 VDDA.n1986 0.0560455
R6473 VDDA.n1997 VDDA.n1996 0.0560455
R6474 VDDA.n2001 VDDA.n2000 0.0560455
R6475 VDDA.n2011 VDDA.n2010 0.0560455
R6476 VDDA.n2017 VDDA.n2016 0.0560455
R6477 VDDA.n2027 VDDA.n2026 0.0560455
R6478 VDDA.n2031 VDDA.n2030 0.0560455
R6479 VDDA.n2041 VDDA.n2040 0.0560455
R6480 VDDA.n2047 VDDA.n2046 0.0560455
R6481 VDDA.n2055 VDDA.n1517 0.0560455
R6482 VDDA.n1619 VDDA.n1618 0.0553333
R6483 VDDA.n1633 VDDA.n1632 0.0553333
R6484 VDDA.n1649 VDDA.n1648 0.0553333
R6485 VDDA.n1663 VDDA.n1662 0.0553333
R6486 VDDA.n1679 VDDA.n1678 0.0553333
R6487 VDDA.n1693 VDDA.n1692 0.0553333
R6488 VDDA.n1709 VDDA.n1708 0.0553333
R6489 VDDA.n1723 VDDA.n1722 0.0553333
R6490 VDDA.n2296 VDDA.n2295 0.0553333
R6491 VDDA.n2310 VDDA.n2309 0.0553333
R6492 VDDA.n2326 VDDA.n2325 0.0553333
R6493 VDDA.n2340 VDDA.n2339 0.0553333
R6494 VDDA.n2356 VDDA.n2355 0.0553333
R6495 VDDA.n2370 VDDA.n2369 0.0553333
R6496 VDDA.n2386 VDDA.n2385 0.0553333
R6497 VDDA.n2400 VDDA.n2399 0.0553333
R6498 VDDA.n89 VDDA.n88 0.0553333
R6499 VDDA.n106 VDDA.n105 0.0553333
R6500 VDDA.n77 VDDA.n76 0.0553333
R6501 VDDA.n130 VDDA.n129 0.0553333
R6502 VDDA.n65 VDDA.n64 0.0553333
R6503 VDDA.n154 VDDA.n153 0.0553333
R6504 VDDA.n53 VDDA.n52 0.0553333
R6505 VDDA.n178 VDDA.n177 0.0553333
R6506 VDDA.n2812 VDDA.n2810 0.0553333
R6507 VDDA.n2828 VDDA.n2797 0.0553333
R6508 VDDA.n2842 VDDA.n2840 0.0553333
R6509 VDDA.n2858 VDDA.n2785 0.0553333
R6510 VDDA.n2872 VDDA.n2870 0.0553333
R6511 VDDA.n2888 VDDA.n2773 0.0553333
R6512 VDDA.n2902 VDDA.n2900 0.0553333
R6513 VDDA.n2918 VDDA.n2761 0.0553333
R6514 VDDA.n2661 VDDA.n2660 0.0553333
R6515 VDDA.n2650 VDDA.n2649 0.0553333
R6516 VDDA.n2685 VDDA.n2684 0.0553333
R6517 VDDA.n2638 VDDA.n2637 0.0553333
R6518 VDDA.n2709 VDDA.n2708 0.0553333
R6519 VDDA.n2626 VDDA.n2625 0.0553333
R6520 VDDA.n2733 VDDA.n2732 0.0553333
R6521 VDDA.n2747 VDDA.n2613 0.0553333
R6522 VDDA.n267 VDDA.n266 0.0553333
R6523 VDDA.n284 VDDA.n283 0.0553333
R6524 VDDA.n255 VDDA.n254 0.0553333
R6525 VDDA.n308 VDDA.n307 0.0553333
R6526 VDDA.n243 VDDA.n242 0.0553333
R6527 VDDA.n332 VDDA.n331 0.0553333
R6528 VDDA.n231 VDDA.n230 0.0553333
R6529 VDDA.n356 VDDA.n355 0.0553333
R6530 VDDA.n418 VDDA.n416 0.0553333
R6531 VDDA.n434 VDDA.n403 0.0553333
R6532 VDDA.n448 VDDA.n446 0.0553333
R6533 VDDA.n464 VDDA.n391 0.0553333
R6534 VDDA.n478 VDDA.n476 0.0553333
R6535 VDDA.n494 VDDA.n379 0.0553333
R6536 VDDA.n508 VDDA.n506 0.0553333
R6537 VDDA.n524 VDDA.n367 0.0553333
R6538 VDDA.n1381 VDDA.n1380 0.0553333
R6539 VDDA.n1370 VDDA.n1369 0.0553333
R6540 VDDA.n1405 VDDA.n1404 0.0553333
R6541 VDDA.n1358 VDDA.n1357 0.0553333
R6542 VDDA.n1429 VDDA.n1428 0.0553333
R6543 VDDA.n1346 VDDA.n1345 0.0553333
R6544 VDDA.n1453 VDDA.n1452 0.0553333
R6545 VDDA.n1467 VDDA.n1333 0.0553333
R6546 VDDA.n682 VDDA.n681 0.0553333
R6547 VDDA.n699 VDDA.n698 0.0553333
R6548 VDDA.n670 VDDA.n669 0.0553333
R6549 VDDA.n723 VDDA.n722 0.0553333
R6550 VDDA.n658 VDDA.n657 0.0553333
R6551 VDDA.n747 VDDA.n746 0.0553333
R6552 VDDA.n646 VDDA.n645 0.0553333
R6553 VDDA.n771 VDDA.n770 0.0553333
R6554 VDDA.n1184 VDDA.n1182 0.0553333
R6555 VDDA.n1200 VDDA.n1169 0.0553333
R6556 VDDA.n1214 VDDA.n1212 0.0553333
R6557 VDDA.n1230 VDDA.n1157 0.0553333
R6558 VDDA.n1244 VDDA.n1242 0.0553333
R6559 VDDA.n1260 VDDA.n1145 0.0553333
R6560 VDDA.n1274 VDDA.n1272 0.0553333
R6561 VDDA.n1290 VDDA.n1133 0.0553333
R6562 VDDA.n1033 VDDA.n1032 0.0553333
R6563 VDDA.n1022 VDDA.n1021 0.0553333
R6564 VDDA.n1057 VDDA.n1056 0.0553333
R6565 VDDA.n1010 VDDA.n1009 0.0553333
R6566 VDDA.n1081 VDDA.n1080 0.0553333
R6567 VDDA.n998 VDDA.n997 0.0553333
R6568 VDDA.n1105 VDDA.n1104 0.0553333
R6569 VDDA.n1119 VDDA.n985 0.0553333
R6570 VDDA.n843 VDDA.n842 0.0553333
R6571 VDDA.n857 VDDA.n856 0.0553333
R6572 VDDA.n873 VDDA.n872 0.0553333
R6573 VDDA.n887 VDDA.n886 0.0553333
R6574 VDDA.n903 VDDA.n902 0.0553333
R6575 VDDA.n917 VDDA.n916 0.0553333
R6576 VDDA.n933 VDDA.n932 0.0553333
R6577 VDDA.n947 VDDA.n946 0.0553333
R6578 VDDA.n1613 VDDA.n1558 0.0514167
R6579 VDDA.n1623 VDDA.n1622 0.0514167
R6580 VDDA.n1629 VDDA.n1628 0.0514167
R6581 VDDA.n1639 VDDA.n1638 0.0514167
R6582 VDDA.n1643 VDDA.n1642 0.0514167
R6583 VDDA.n1653 VDDA.n1652 0.0514167
R6584 VDDA.n1659 VDDA.n1658 0.0514167
R6585 VDDA.n1669 VDDA.n1668 0.0514167
R6586 VDDA.n1673 VDDA.n1672 0.0514167
R6587 VDDA.n1683 VDDA.n1682 0.0514167
R6588 VDDA.n1689 VDDA.n1688 0.0514167
R6589 VDDA.n1699 VDDA.n1698 0.0514167
R6590 VDDA.n1703 VDDA.n1702 0.0514167
R6591 VDDA.n1713 VDDA.n1712 0.0514167
R6592 VDDA.n1719 VDDA.n1718 0.0514167
R6593 VDDA.n1727 VDDA.n1582 0.0514167
R6594 VDDA.n2300 VDDA.n2299 0.0514167
R6595 VDDA.n2306 VDDA.n2305 0.0514167
R6596 VDDA.n2316 VDDA.n2315 0.0514167
R6597 VDDA.n2320 VDDA.n2319 0.0514167
R6598 VDDA.n2330 VDDA.n2329 0.0514167
R6599 VDDA.n2336 VDDA.n2335 0.0514167
R6600 VDDA.n2346 VDDA.n2345 0.0514167
R6601 VDDA.n2350 VDDA.n2349 0.0514167
R6602 VDDA.n2360 VDDA.n2359 0.0514167
R6603 VDDA.n2366 VDDA.n2365 0.0514167
R6604 VDDA.n2376 VDDA.n2375 0.0514167
R6605 VDDA.n2380 VDDA.n2379 0.0514167
R6606 VDDA.n2390 VDDA.n2389 0.0514167
R6607 VDDA.n2396 VDDA.n2395 0.0514167
R6608 VDDA.n2404 VDDA.n2057 0.0514167
R6609 VDDA.n90 VDDA.n20 0.0514167
R6610 VDDA.n98 VDDA.n97 0.0514167
R6611 VDDA.n85 VDDA.n84 0.0514167
R6612 VDDA.n81 VDDA.n80 0.0514167
R6613 VDDA.n114 VDDA.n113 0.0514167
R6614 VDDA.n122 VDDA.n121 0.0514167
R6615 VDDA.n73 VDDA.n72 0.0514167
R6616 VDDA.n69 VDDA.n68 0.0514167
R6617 VDDA.n138 VDDA.n137 0.0514167
R6618 VDDA.n146 VDDA.n145 0.0514167
R6619 VDDA.n61 VDDA.n60 0.0514167
R6620 VDDA.n57 VDDA.n56 0.0514167
R6621 VDDA.n162 VDDA.n161 0.0514167
R6622 VDDA.n170 VDDA.n169 0.0514167
R6623 VDDA.n49 VDDA.n48 0.0514167
R6624 VDDA.n2936 VDDA.n44 0.0514167
R6625 VDDA.n2808 VDDA.n2805 0.0514167
R6626 VDDA.n2818 VDDA.n2801 0.0514167
R6627 VDDA.n2822 VDDA.n2820 0.0514167
R6628 VDDA.n2832 VDDA.n2830 0.0514167
R6629 VDDA.n2838 VDDA.n2793 0.0514167
R6630 VDDA.n2848 VDDA.n2789 0.0514167
R6631 VDDA.n2852 VDDA.n2850 0.0514167
R6632 VDDA.n2862 VDDA.n2860 0.0514167
R6633 VDDA.n2868 VDDA.n2781 0.0514167
R6634 VDDA.n2878 VDDA.n2777 0.0514167
R6635 VDDA.n2882 VDDA.n2880 0.0514167
R6636 VDDA.n2892 VDDA.n2890 0.0514167
R6637 VDDA.n2898 VDDA.n2769 0.0514167
R6638 VDDA.n2908 VDDA.n2765 0.0514167
R6639 VDDA.n2912 VDDA.n2910 0.0514167
R6640 VDDA.n2921 VDDA.n2920 0.0514167
R6641 VDDA.n2657 VDDA.n2590 0.0514167
R6642 VDDA.n2654 VDDA.n2653 0.0514167
R6643 VDDA.n2669 VDDA.n2668 0.0514167
R6644 VDDA.n2677 VDDA.n2676 0.0514167
R6645 VDDA.n2646 VDDA.n2645 0.0514167
R6646 VDDA.n2642 VDDA.n2641 0.0514167
R6647 VDDA.n2693 VDDA.n2692 0.0514167
R6648 VDDA.n2701 VDDA.n2700 0.0514167
R6649 VDDA.n2634 VDDA.n2633 0.0514167
R6650 VDDA.n2630 VDDA.n2629 0.0514167
R6651 VDDA.n2717 VDDA.n2716 0.0514167
R6652 VDDA.n2725 VDDA.n2724 0.0514167
R6653 VDDA.n2622 VDDA.n2621 0.0514167
R6654 VDDA.n2618 VDDA.n2617 0.0514167
R6655 VDDA.n2741 VDDA.n2740 0.0514167
R6656 VDDA.n2750 VDDA.n196 0.0514167
R6657 VDDA.n268 VDDA.n198 0.0514167
R6658 VDDA.n276 VDDA.n275 0.0514167
R6659 VDDA.n263 VDDA.n262 0.0514167
R6660 VDDA.n259 VDDA.n258 0.0514167
R6661 VDDA.n292 VDDA.n291 0.0514167
R6662 VDDA.n300 VDDA.n299 0.0514167
R6663 VDDA.n251 VDDA.n250 0.0514167
R6664 VDDA.n247 VDDA.n246 0.0514167
R6665 VDDA.n316 VDDA.n315 0.0514167
R6666 VDDA.n324 VDDA.n323 0.0514167
R6667 VDDA.n239 VDDA.n238 0.0514167
R6668 VDDA.n235 VDDA.n234 0.0514167
R6669 VDDA.n340 VDDA.n339 0.0514167
R6670 VDDA.n348 VDDA.n347 0.0514167
R6671 VDDA.n227 VDDA.n226 0.0514167
R6672 VDDA.n2588 VDDA.n222 0.0514167
R6673 VDDA.n414 VDDA.n411 0.0514167
R6674 VDDA.n424 VDDA.n407 0.0514167
R6675 VDDA.n428 VDDA.n426 0.0514167
R6676 VDDA.n438 VDDA.n436 0.0514167
R6677 VDDA.n444 VDDA.n399 0.0514167
R6678 VDDA.n454 VDDA.n395 0.0514167
R6679 VDDA.n458 VDDA.n456 0.0514167
R6680 VDDA.n468 VDDA.n466 0.0514167
R6681 VDDA.n474 VDDA.n387 0.0514167
R6682 VDDA.n484 VDDA.n383 0.0514167
R6683 VDDA.n488 VDDA.n486 0.0514167
R6684 VDDA.n498 VDDA.n496 0.0514167
R6685 VDDA.n504 VDDA.n375 0.0514167
R6686 VDDA.n514 VDDA.n371 0.0514167
R6687 VDDA.n518 VDDA.n516 0.0514167
R6688 VDDA.n527 VDDA.n526 0.0514167
R6689 VDDA.n1377 VDDA.n1310 0.0514167
R6690 VDDA.n1374 VDDA.n1373 0.0514167
R6691 VDDA.n1389 VDDA.n1388 0.0514167
R6692 VDDA.n1397 VDDA.n1396 0.0514167
R6693 VDDA.n1366 VDDA.n1365 0.0514167
R6694 VDDA.n1362 VDDA.n1361 0.0514167
R6695 VDDA.n1413 VDDA.n1412 0.0514167
R6696 VDDA.n1421 VDDA.n1420 0.0514167
R6697 VDDA.n1354 VDDA.n1353 0.0514167
R6698 VDDA.n1350 VDDA.n1349 0.0514167
R6699 VDDA.n1437 VDDA.n1436 0.0514167
R6700 VDDA.n1445 VDDA.n1444 0.0514167
R6701 VDDA.n1342 VDDA.n1341 0.0514167
R6702 VDDA.n1338 VDDA.n1337 0.0514167
R6703 VDDA.n1461 VDDA.n1460 0.0514167
R6704 VDDA.n2407 VDDA.n611 0.0514167
R6705 VDDA.n683 VDDA.n613 0.0514167
R6706 VDDA.n691 VDDA.n690 0.0514167
R6707 VDDA.n678 VDDA.n677 0.0514167
R6708 VDDA.n674 VDDA.n673 0.0514167
R6709 VDDA.n707 VDDA.n706 0.0514167
R6710 VDDA.n715 VDDA.n714 0.0514167
R6711 VDDA.n666 VDDA.n665 0.0514167
R6712 VDDA.n662 VDDA.n661 0.0514167
R6713 VDDA.n731 VDDA.n730 0.0514167
R6714 VDDA.n739 VDDA.n738 0.0514167
R6715 VDDA.n654 VDDA.n653 0.0514167
R6716 VDDA.n650 VDDA.n649 0.0514167
R6717 VDDA.n755 VDDA.n754 0.0514167
R6718 VDDA.n763 VDDA.n762 0.0514167
R6719 VDDA.n642 VDDA.n641 0.0514167
R6720 VDDA.n1308 VDDA.n637 0.0514167
R6721 VDDA.n1180 VDDA.n1177 0.0514167
R6722 VDDA.n1190 VDDA.n1173 0.0514167
R6723 VDDA.n1194 VDDA.n1192 0.0514167
R6724 VDDA.n1204 VDDA.n1202 0.0514167
R6725 VDDA.n1210 VDDA.n1165 0.0514167
R6726 VDDA.n1220 VDDA.n1161 0.0514167
R6727 VDDA.n1224 VDDA.n1222 0.0514167
R6728 VDDA.n1234 VDDA.n1232 0.0514167
R6729 VDDA.n1240 VDDA.n1153 0.0514167
R6730 VDDA.n1250 VDDA.n1149 0.0514167
R6731 VDDA.n1254 VDDA.n1252 0.0514167
R6732 VDDA.n1264 VDDA.n1262 0.0514167
R6733 VDDA.n1270 VDDA.n1141 0.0514167
R6734 VDDA.n1280 VDDA.n1137 0.0514167
R6735 VDDA.n1284 VDDA.n1282 0.0514167
R6736 VDDA.n1293 VDDA.n1292 0.0514167
R6737 VDDA.n1029 VDDA.n962 0.0514167
R6738 VDDA.n1026 VDDA.n1025 0.0514167
R6739 VDDA.n1041 VDDA.n1040 0.0514167
R6740 VDDA.n1049 VDDA.n1048 0.0514167
R6741 VDDA.n1018 VDDA.n1017 0.0514167
R6742 VDDA.n1014 VDDA.n1013 0.0514167
R6743 VDDA.n1065 VDDA.n1064 0.0514167
R6744 VDDA.n1073 VDDA.n1072 0.0514167
R6745 VDDA.n1006 VDDA.n1005 0.0514167
R6746 VDDA.n1002 VDDA.n1001 0.0514167
R6747 VDDA.n1089 VDDA.n1088 0.0514167
R6748 VDDA.n1097 VDDA.n1096 0.0514167
R6749 VDDA.n994 VDDA.n993 0.0514167
R6750 VDDA.n990 VDDA.n989 0.0514167
R6751 VDDA.n1113 VDDA.n1112 0.0514167
R6752 VDDA.n1122 VDDA.n788 0.0514167
R6753 VDDA.n837 VDDA.n789 0.0514167
R6754 VDDA.n847 VDDA.n846 0.0514167
R6755 VDDA.n853 VDDA.n852 0.0514167
R6756 VDDA.n863 VDDA.n862 0.0514167
R6757 VDDA.n867 VDDA.n866 0.0514167
R6758 VDDA.n877 VDDA.n876 0.0514167
R6759 VDDA.n883 VDDA.n882 0.0514167
R6760 VDDA.n893 VDDA.n892 0.0514167
R6761 VDDA.n897 VDDA.n896 0.0514167
R6762 VDDA.n907 VDDA.n906 0.0514167
R6763 VDDA.n913 VDDA.n912 0.0514167
R6764 VDDA.n923 VDDA.n922 0.0514167
R6765 VDDA.n927 VDDA.n926 0.0514167
R6766 VDDA.n937 VDDA.n936 0.0514167
R6767 VDDA.n943 VDDA.n942 0.0514167
R6768 VDDA.n960 VDDA.n813 0.0514167
R6769 VDDA.n2405 VDDA.n2056 0.0497766
R6770 VDDA.n2295 VDDA.n1469 0.0459984
R6771 VDDA.n2484 VDDA.n544 0.0429747
R6772 VDDA.n361 VDDA.n192 0.0421667
R6773 VDDA.n2757 VDDA.n189 0.0421667
R6774 VDDA.n2928 VDDA.n186 0.0421667
R6775 VDDA.n2931 VDDA.n184 0.0421667
R6776 VDDA.n2572 VDDA.n533 0.0421667
R6777 VDDA.n2495 VDDA.n540 0.0421667
R6778 VDDA.n2437 VDDA.n565 0.0421667
R6779 VDDA.n1129 VDDA.n781 0.0421667
R6780 VDDA.n1300 VDDA.n778 0.0421667
R6781 VDDA.n776 VDDA.n606 0.0421667
R6782 VDDA.n608 VDDA.n605 0.0421667
R6783 VDDA.n1800 VDDA.n1799 0.0352506
R6784 VDDA.n1914 VDDA.n1913 0.0331087
R6785 VDDA.n1946 VDDA.n1493 0.030649
R6786 VDDA.n1950 VDDA.n1494 0.030649
R6787 VDDA.n1960 VDDA.n1496 0.030649
R6788 VDDA.n1966 VDDA.n1497 0.030649
R6789 VDDA.n1976 VDDA.n1499 0.030649
R6790 VDDA.n1980 VDDA.n1500 0.030649
R6791 VDDA.n1990 VDDA.n1502 0.030649
R6792 VDDA.n1996 VDDA.n1503 0.030649
R6793 VDDA.n2006 VDDA.n1505 0.030649
R6794 VDDA.n2010 VDDA.n1506 0.030649
R6795 VDDA.n2020 VDDA.n1508 0.030649
R6796 VDDA.n2026 VDDA.n1509 0.030649
R6797 VDDA.n2036 VDDA.n1511 0.030649
R6798 VDDA.n2040 VDDA.n1512 0.030649
R6799 VDDA.n2050 VDDA.n1514 0.030649
R6800 VDDA.n1517 VDDA.n1515 0.030649
R6801 VDDA.n2051 VDDA.n1515 0.030649
R6802 VDDA.n2047 VDDA.n1514 0.030649
R6803 VDDA.n2037 VDDA.n1512 0.030649
R6804 VDDA.n2031 VDDA.n1511 0.030649
R6805 VDDA.n2021 VDDA.n1509 0.030649
R6806 VDDA.n2017 VDDA.n1508 0.030649
R6807 VDDA.n2007 VDDA.n1506 0.030649
R6808 VDDA.n2001 VDDA.n1505 0.030649
R6809 VDDA.n1991 VDDA.n1503 0.030649
R6810 VDDA.n1987 VDDA.n1502 0.030649
R6811 VDDA.n1977 VDDA.n1500 0.030649
R6812 VDDA.n1971 VDDA.n1499 0.030649
R6813 VDDA.n1961 VDDA.n1497 0.030649
R6814 VDDA.n1957 VDDA.n1496 0.030649
R6815 VDDA.n1947 VDDA.n1494 0.030649
R6816 VDDA.n1941 VDDA.n1493 0.030649
R6817 VDDA.n1618 VDDA.n1559 0.028198
R6818 VDDA.n1622 VDDA.n1560 0.028198
R6819 VDDA.n1632 VDDA.n1562 0.028198
R6820 VDDA.n1638 VDDA.n1563 0.028198
R6821 VDDA.n1648 VDDA.n1565 0.028198
R6822 VDDA.n1652 VDDA.n1566 0.028198
R6823 VDDA.n1662 VDDA.n1568 0.028198
R6824 VDDA.n1668 VDDA.n1569 0.028198
R6825 VDDA.n1678 VDDA.n1571 0.028198
R6826 VDDA.n1682 VDDA.n1572 0.028198
R6827 VDDA.n1692 VDDA.n1574 0.028198
R6828 VDDA.n1698 VDDA.n1575 0.028198
R6829 VDDA.n1708 VDDA.n1577 0.028198
R6830 VDDA.n1712 VDDA.n1578 0.028198
R6831 VDDA.n1722 VDDA.n1580 0.028198
R6832 VDDA.n1582 VDDA.n1581 0.028198
R6833 VDDA.n2299 VDDA.n1470 0.028198
R6834 VDDA.n2309 VDDA.n1472 0.028198
R6835 VDDA.n2315 VDDA.n1473 0.028198
R6836 VDDA.n2325 VDDA.n1475 0.028198
R6837 VDDA.n2329 VDDA.n1476 0.028198
R6838 VDDA.n2339 VDDA.n1478 0.028198
R6839 VDDA.n2345 VDDA.n1479 0.028198
R6840 VDDA.n2355 VDDA.n1481 0.028198
R6841 VDDA.n2359 VDDA.n1482 0.028198
R6842 VDDA.n2369 VDDA.n1484 0.028198
R6843 VDDA.n2375 VDDA.n1485 0.028198
R6844 VDDA.n2385 VDDA.n1487 0.028198
R6845 VDDA.n2389 VDDA.n1488 0.028198
R6846 VDDA.n2399 VDDA.n1490 0.028198
R6847 VDDA.n2057 VDDA.n1491 0.028198
R6848 VDDA.n88 VDDA.n21 0.028198
R6849 VDDA.n97 VDDA.n22 0.028198
R6850 VDDA.n105 VDDA.n24 0.028198
R6851 VDDA.n80 VDDA.n25 0.028198
R6852 VDDA.n76 VDDA.n27 0.028198
R6853 VDDA.n121 VDDA.n28 0.028198
R6854 VDDA.n129 VDDA.n30 0.028198
R6855 VDDA.n68 VDDA.n31 0.028198
R6856 VDDA.n64 VDDA.n33 0.028198
R6857 VDDA.n145 VDDA.n34 0.028198
R6858 VDDA.n153 VDDA.n36 0.028198
R6859 VDDA.n56 VDDA.n37 0.028198
R6860 VDDA.n52 VDDA.n39 0.028198
R6861 VDDA.n169 VDDA.n40 0.028198
R6862 VDDA.n177 VDDA.n42 0.028198
R6863 VDDA.n44 VDDA.n43 0.028198
R6864 VDDA.n2810 VDDA.n2809 0.028198
R6865 VDDA.n2811 VDDA.n2801 0.028198
R6866 VDDA.n2821 VDDA.n2797 0.028198
R6867 VDDA.n2830 VDDA.n2829 0.028198
R6868 VDDA.n2840 VDDA.n2839 0.028198
R6869 VDDA.n2841 VDDA.n2789 0.028198
R6870 VDDA.n2851 VDDA.n2785 0.028198
R6871 VDDA.n2860 VDDA.n2859 0.028198
R6872 VDDA.n2870 VDDA.n2869 0.028198
R6873 VDDA.n2871 VDDA.n2777 0.028198
R6874 VDDA.n2881 VDDA.n2773 0.028198
R6875 VDDA.n2890 VDDA.n2889 0.028198
R6876 VDDA.n2900 VDDA.n2899 0.028198
R6877 VDDA.n2901 VDDA.n2765 0.028198
R6878 VDDA.n2911 VDDA.n2761 0.028198
R6879 VDDA.n2920 VDDA.n2919 0.028198
R6880 VDDA.n2660 VDDA.n2591 0.028198
R6881 VDDA.n2653 VDDA.n2592 0.028198
R6882 VDDA.n2649 VDDA.n2594 0.028198
R6883 VDDA.n2676 VDDA.n2595 0.028198
R6884 VDDA.n2684 VDDA.n2597 0.028198
R6885 VDDA.n2641 VDDA.n2598 0.028198
R6886 VDDA.n2637 VDDA.n2600 0.028198
R6887 VDDA.n2700 VDDA.n2601 0.028198
R6888 VDDA.n2708 VDDA.n2603 0.028198
R6889 VDDA.n2629 VDDA.n2604 0.028198
R6890 VDDA.n2625 VDDA.n2606 0.028198
R6891 VDDA.n2724 VDDA.n2607 0.028198
R6892 VDDA.n2732 VDDA.n2609 0.028198
R6893 VDDA.n2617 VDDA.n2610 0.028198
R6894 VDDA.n2613 VDDA.n2612 0.028198
R6895 VDDA.n2748 VDDA.n196 0.028198
R6896 VDDA.n266 VDDA.n199 0.028198
R6897 VDDA.n275 VDDA.n200 0.028198
R6898 VDDA.n283 VDDA.n202 0.028198
R6899 VDDA.n258 VDDA.n203 0.028198
R6900 VDDA.n254 VDDA.n205 0.028198
R6901 VDDA.n299 VDDA.n206 0.028198
R6902 VDDA.n307 VDDA.n208 0.028198
R6903 VDDA.n246 VDDA.n209 0.028198
R6904 VDDA.n242 VDDA.n211 0.028198
R6905 VDDA.n323 VDDA.n212 0.028198
R6906 VDDA.n331 VDDA.n214 0.028198
R6907 VDDA.n234 VDDA.n215 0.028198
R6908 VDDA.n230 VDDA.n217 0.028198
R6909 VDDA.n347 VDDA.n218 0.028198
R6910 VDDA.n355 VDDA.n220 0.028198
R6911 VDDA.n222 VDDA.n221 0.028198
R6912 VDDA.n416 VDDA.n415 0.028198
R6913 VDDA.n417 VDDA.n407 0.028198
R6914 VDDA.n427 VDDA.n403 0.028198
R6915 VDDA.n436 VDDA.n435 0.028198
R6916 VDDA.n446 VDDA.n445 0.028198
R6917 VDDA.n447 VDDA.n395 0.028198
R6918 VDDA.n457 VDDA.n391 0.028198
R6919 VDDA.n466 VDDA.n465 0.028198
R6920 VDDA.n476 VDDA.n475 0.028198
R6921 VDDA.n477 VDDA.n383 0.028198
R6922 VDDA.n487 VDDA.n379 0.028198
R6923 VDDA.n496 VDDA.n495 0.028198
R6924 VDDA.n506 VDDA.n505 0.028198
R6925 VDDA.n507 VDDA.n371 0.028198
R6926 VDDA.n517 VDDA.n367 0.028198
R6927 VDDA.n526 VDDA.n525 0.028198
R6928 VDDA.n1380 VDDA.n1311 0.028198
R6929 VDDA.n1373 VDDA.n1312 0.028198
R6930 VDDA.n1369 VDDA.n1314 0.028198
R6931 VDDA.n1396 VDDA.n1315 0.028198
R6932 VDDA.n1404 VDDA.n1317 0.028198
R6933 VDDA.n1361 VDDA.n1318 0.028198
R6934 VDDA.n1357 VDDA.n1320 0.028198
R6935 VDDA.n1420 VDDA.n1321 0.028198
R6936 VDDA.n1428 VDDA.n1323 0.028198
R6937 VDDA.n1349 VDDA.n1324 0.028198
R6938 VDDA.n1345 VDDA.n1326 0.028198
R6939 VDDA.n1444 VDDA.n1327 0.028198
R6940 VDDA.n1452 VDDA.n1329 0.028198
R6941 VDDA.n1337 VDDA.n1330 0.028198
R6942 VDDA.n1333 VDDA.n1332 0.028198
R6943 VDDA.n1468 VDDA.n611 0.028198
R6944 VDDA.n681 VDDA.n614 0.028198
R6945 VDDA.n690 VDDA.n615 0.028198
R6946 VDDA.n698 VDDA.n617 0.028198
R6947 VDDA.n673 VDDA.n618 0.028198
R6948 VDDA.n669 VDDA.n620 0.028198
R6949 VDDA.n714 VDDA.n621 0.028198
R6950 VDDA.n722 VDDA.n623 0.028198
R6951 VDDA.n661 VDDA.n624 0.028198
R6952 VDDA.n657 VDDA.n626 0.028198
R6953 VDDA.n738 VDDA.n627 0.028198
R6954 VDDA.n746 VDDA.n629 0.028198
R6955 VDDA.n649 VDDA.n630 0.028198
R6956 VDDA.n645 VDDA.n632 0.028198
R6957 VDDA.n762 VDDA.n633 0.028198
R6958 VDDA.n770 VDDA.n635 0.028198
R6959 VDDA.n637 VDDA.n636 0.028198
R6960 VDDA.n1182 VDDA.n1181 0.028198
R6961 VDDA.n1183 VDDA.n1173 0.028198
R6962 VDDA.n1193 VDDA.n1169 0.028198
R6963 VDDA.n1202 VDDA.n1201 0.028198
R6964 VDDA.n1212 VDDA.n1211 0.028198
R6965 VDDA.n1213 VDDA.n1161 0.028198
R6966 VDDA.n1223 VDDA.n1157 0.028198
R6967 VDDA.n1232 VDDA.n1231 0.028198
R6968 VDDA.n1242 VDDA.n1241 0.028198
R6969 VDDA.n1243 VDDA.n1149 0.028198
R6970 VDDA.n1253 VDDA.n1145 0.028198
R6971 VDDA.n1262 VDDA.n1261 0.028198
R6972 VDDA.n1272 VDDA.n1271 0.028198
R6973 VDDA.n1273 VDDA.n1137 0.028198
R6974 VDDA.n1283 VDDA.n1133 0.028198
R6975 VDDA.n1292 VDDA.n1291 0.028198
R6976 VDDA.n1032 VDDA.n963 0.028198
R6977 VDDA.n1025 VDDA.n964 0.028198
R6978 VDDA.n1021 VDDA.n966 0.028198
R6979 VDDA.n1048 VDDA.n967 0.028198
R6980 VDDA.n1056 VDDA.n969 0.028198
R6981 VDDA.n1013 VDDA.n970 0.028198
R6982 VDDA.n1009 VDDA.n972 0.028198
R6983 VDDA.n1072 VDDA.n973 0.028198
R6984 VDDA.n1080 VDDA.n975 0.028198
R6985 VDDA.n1001 VDDA.n976 0.028198
R6986 VDDA.n997 VDDA.n978 0.028198
R6987 VDDA.n1096 VDDA.n979 0.028198
R6988 VDDA.n1104 VDDA.n981 0.028198
R6989 VDDA.n989 VDDA.n982 0.028198
R6990 VDDA.n985 VDDA.n984 0.028198
R6991 VDDA.n1120 VDDA.n788 0.028198
R6992 VDDA.n842 VDDA.n790 0.028198
R6993 VDDA.n846 VDDA.n791 0.028198
R6994 VDDA.n856 VDDA.n793 0.028198
R6995 VDDA.n862 VDDA.n794 0.028198
R6996 VDDA.n872 VDDA.n796 0.028198
R6997 VDDA.n876 VDDA.n797 0.028198
R6998 VDDA.n886 VDDA.n799 0.028198
R6999 VDDA.n892 VDDA.n800 0.028198
R7000 VDDA.n902 VDDA.n802 0.028198
R7001 VDDA.n906 VDDA.n803 0.028198
R7002 VDDA.n916 VDDA.n805 0.028198
R7003 VDDA.n922 VDDA.n806 0.028198
R7004 VDDA.n932 VDDA.n808 0.028198
R7005 VDDA.n936 VDDA.n809 0.028198
R7006 VDDA.n946 VDDA.n811 0.028198
R7007 VDDA.n813 VDDA.n812 0.028198
R7008 VDDA.n947 VDDA.n812 0.028198
R7009 VDDA.n943 VDDA.n811 0.028198
R7010 VDDA.n933 VDDA.n809 0.028198
R7011 VDDA.n927 VDDA.n808 0.028198
R7012 VDDA.n917 VDDA.n806 0.028198
R7013 VDDA.n913 VDDA.n805 0.028198
R7014 VDDA.n903 VDDA.n803 0.028198
R7015 VDDA.n897 VDDA.n802 0.028198
R7016 VDDA.n887 VDDA.n800 0.028198
R7017 VDDA.n883 VDDA.n799 0.028198
R7018 VDDA.n873 VDDA.n797 0.028198
R7019 VDDA.n867 VDDA.n796 0.028198
R7020 VDDA.n857 VDDA.n794 0.028198
R7021 VDDA.n853 VDDA.n793 0.028198
R7022 VDDA.n843 VDDA.n791 0.028198
R7023 VDDA.n837 VDDA.n790 0.028198
R7024 VDDA.n1120 VDDA.n1119 0.028198
R7025 VDDA.n1113 VDDA.n984 0.028198
R7026 VDDA.n1105 VDDA.n982 0.028198
R7027 VDDA.n994 VDDA.n981 0.028198
R7028 VDDA.n998 VDDA.n979 0.028198
R7029 VDDA.n1089 VDDA.n978 0.028198
R7030 VDDA.n1081 VDDA.n976 0.028198
R7031 VDDA.n1006 VDDA.n975 0.028198
R7032 VDDA.n1010 VDDA.n973 0.028198
R7033 VDDA.n1065 VDDA.n972 0.028198
R7034 VDDA.n1057 VDDA.n970 0.028198
R7035 VDDA.n1018 VDDA.n969 0.028198
R7036 VDDA.n1022 VDDA.n967 0.028198
R7037 VDDA.n1041 VDDA.n966 0.028198
R7038 VDDA.n1033 VDDA.n964 0.028198
R7039 VDDA.n1029 VDDA.n963 0.028198
R7040 VDDA.n1291 VDDA.n1290 0.028198
R7041 VDDA.n1284 VDDA.n1283 0.028198
R7042 VDDA.n1274 VDDA.n1273 0.028198
R7043 VDDA.n1271 VDDA.n1270 0.028198
R7044 VDDA.n1261 VDDA.n1260 0.028198
R7045 VDDA.n1254 VDDA.n1253 0.028198
R7046 VDDA.n1244 VDDA.n1243 0.028198
R7047 VDDA.n1241 VDDA.n1240 0.028198
R7048 VDDA.n1231 VDDA.n1230 0.028198
R7049 VDDA.n1224 VDDA.n1223 0.028198
R7050 VDDA.n1214 VDDA.n1213 0.028198
R7051 VDDA.n1211 VDDA.n1210 0.028198
R7052 VDDA.n1201 VDDA.n1200 0.028198
R7053 VDDA.n1194 VDDA.n1193 0.028198
R7054 VDDA.n1184 VDDA.n1183 0.028198
R7055 VDDA.n1181 VDDA.n1180 0.028198
R7056 VDDA.n771 VDDA.n636 0.028198
R7057 VDDA.n642 VDDA.n635 0.028198
R7058 VDDA.n646 VDDA.n633 0.028198
R7059 VDDA.n755 VDDA.n632 0.028198
R7060 VDDA.n747 VDDA.n630 0.028198
R7061 VDDA.n654 VDDA.n629 0.028198
R7062 VDDA.n658 VDDA.n627 0.028198
R7063 VDDA.n731 VDDA.n626 0.028198
R7064 VDDA.n723 VDDA.n624 0.028198
R7065 VDDA.n666 VDDA.n623 0.028198
R7066 VDDA.n670 VDDA.n621 0.028198
R7067 VDDA.n707 VDDA.n620 0.028198
R7068 VDDA.n699 VDDA.n618 0.028198
R7069 VDDA.n678 VDDA.n617 0.028198
R7070 VDDA.n682 VDDA.n615 0.028198
R7071 VDDA.n683 VDDA.n614 0.028198
R7072 VDDA.n1468 VDDA.n1467 0.028198
R7073 VDDA.n1461 VDDA.n1332 0.028198
R7074 VDDA.n1453 VDDA.n1330 0.028198
R7075 VDDA.n1342 VDDA.n1329 0.028198
R7076 VDDA.n1346 VDDA.n1327 0.028198
R7077 VDDA.n1437 VDDA.n1326 0.028198
R7078 VDDA.n1429 VDDA.n1324 0.028198
R7079 VDDA.n1354 VDDA.n1323 0.028198
R7080 VDDA.n1358 VDDA.n1321 0.028198
R7081 VDDA.n1413 VDDA.n1320 0.028198
R7082 VDDA.n1405 VDDA.n1318 0.028198
R7083 VDDA.n1366 VDDA.n1317 0.028198
R7084 VDDA.n1370 VDDA.n1315 0.028198
R7085 VDDA.n1389 VDDA.n1314 0.028198
R7086 VDDA.n1381 VDDA.n1312 0.028198
R7087 VDDA.n1377 VDDA.n1311 0.028198
R7088 VDDA.n2400 VDDA.n1491 0.028198
R7089 VDDA.n2396 VDDA.n1490 0.028198
R7090 VDDA.n2386 VDDA.n1488 0.028198
R7091 VDDA.n2380 VDDA.n1487 0.028198
R7092 VDDA.n2370 VDDA.n1485 0.028198
R7093 VDDA.n2366 VDDA.n1484 0.028198
R7094 VDDA.n2356 VDDA.n1482 0.028198
R7095 VDDA.n2350 VDDA.n1481 0.028198
R7096 VDDA.n2340 VDDA.n1479 0.028198
R7097 VDDA.n2336 VDDA.n1478 0.028198
R7098 VDDA.n2326 VDDA.n1476 0.028198
R7099 VDDA.n2320 VDDA.n1475 0.028198
R7100 VDDA.n2310 VDDA.n1473 0.028198
R7101 VDDA.n2306 VDDA.n1472 0.028198
R7102 VDDA.n2296 VDDA.n1470 0.028198
R7103 VDDA.n525 VDDA.n524 0.028198
R7104 VDDA.n518 VDDA.n517 0.028198
R7105 VDDA.n508 VDDA.n507 0.028198
R7106 VDDA.n505 VDDA.n504 0.028198
R7107 VDDA.n495 VDDA.n494 0.028198
R7108 VDDA.n488 VDDA.n487 0.028198
R7109 VDDA.n478 VDDA.n477 0.028198
R7110 VDDA.n475 VDDA.n474 0.028198
R7111 VDDA.n465 VDDA.n464 0.028198
R7112 VDDA.n458 VDDA.n457 0.028198
R7113 VDDA.n448 VDDA.n447 0.028198
R7114 VDDA.n445 VDDA.n444 0.028198
R7115 VDDA.n435 VDDA.n434 0.028198
R7116 VDDA.n428 VDDA.n427 0.028198
R7117 VDDA.n418 VDDA.n417 0.028198
R7118 VDDA.n415 VDDA.n414 0.028198
R7119 VDDA.n356 VDDA.n221 0.028198
R7120 VDDA.n227 VDDA.n220 0.028198
R7121 VDDA.n231 VDDA.n218 0.028198
R7122 VDDA.n340 VDDA.n217 0.028198
R7123 VDDA.n332 VDDA.n215 0.028198
R7124 VDDA.n239 VDDA.n214 0.028198
R7125 VDDA.n243 VDDA.n212 0.028198
R7126 VDDA.n316 VDDA.n211 0.028198
R7127 VDDA.n308 VDDA.n209 0.028198
R7128 VDDA.n251 VDDA.n208 0.028198
R7129 VDDA.n255 VDDA.n206 0.028198
R7130 VDDA.n292 VDDA.n205 0.028198
R7131 VDDA.n284 VDDA.n203 0.028198
R7132 VDDA.n263 VDDA.n202 0.028198
R7133 VDDA.n267 VDDA.n200 0.028198
R7134 VDDA.n268 VDDA.n199 0.028198
R7135 VDDA.n2748 VDDA.n2747 0.028198
R7136 VDDA.n2741 VDDA.n2612 0.028198
R7137 VDDA.n2733 VDDA.n2610 0.028198
R7138 VDDA.n2622 VDDA.n2609 0.028198
R7139 VDDA.n2626 VDDA.n2607 0.028198
R7140 VDDA.n2717 VDDA.n2606 0.028198
R7141 VDDA.n2709 VDDA.n2604 0.028198
R7142 VDDA.n2634 VDDA.n2603 0.028198
R7143 VDDA.n2638 VDDA.n2601 0.028198
R7144 VDDA.n2693 VDDA.n2600 0.028198
R7145 VDDA.n2685 VDDA.n2598 0.028198
R7146 VDDA.n2646 VDDA.n2597 0.028198
R7147 VDDA.n2650 VDDA.n2595 0.028198
R7148 VDDA.n2669 VDDA.n2594 0.028198
R7149 VDDA.n2661 VDDA.n2592 0.028198
R7150 VDDA.n2657 VDDA.n2591 0.028198
R7151 VDDA.n2919 VDDA.n2918 0.028198
R7152 VDDA.n2912 VDDA.n2911 0.028198
R7153 VDDA.n2902 VDDA.n2901 0.028198
R7154 VDDA.n2899 VDDA.n2898 0.028198
R7155 VDDA.n2889 VDDA.n2888 0.028198
R7156 VDDA.n2882 VDDA.n2881 0.028198
R7157 VDDA.n2872 VDDA.n2871 0.028198
R7158 VDDA.n2869 VDDA.n2868 0.028198
R7159 VDDA.n2859 VDDA.n2858 0.028198
R7160 VDDA.n2852 VDDA.n2851 0.028198
R7161 VDDA.n2842 VDDA.n2841 0.028198
R7162 VDDA.n2839 VDDA.n2838 0.028198
R7163 VDDA.n2829 VDDA.n2828 0.028198
R7164 VDDA.n2822 VDDA.n2821 0.028198
R7165 VDDA.n2812 VDDA.n2811 0.028198
R7166 VDDA.n2809 VDDA.n2808 0.028198
R7167 VDDA.n178 VDDA.n43 0.028198
R7168 VDDA.n49 VDDA.n42 0.028198
R7169 VDDA.n53 VDDA.n40 0.028198
R7170 VDDA.n162 VDDA.n39 0.028198
R7171 VDDA.n154 VDDA.n37 0.028198
R7172 VDDA.n61 VDDA.n36 0.028198
R7173 VDDA.n65 VDDA.n34 0.028198
R7174 VDDA.n138 VDDA.n33 0.028198
R7175 VDDA.n130 VDDA.n31 0.028198
R7176 VDDA.n73 VDDA.n30 0.028198
R7177 VDDA.n77 VDDA.n28 0.028198
R7178 VDDA.n114 VDDA.n27 0.028198
R7179 VDDA.n106 VDDA.n25 0.028198
R7180 VDDA.n85 VDDA.n24 0.028198
R7181 VDDA.n89 VDDA.n22 0.028198
R7182 VDDA.n90 VDDA.n21 0.028198
R7183 VDDA.n1723 VDDA.n1581 0.028198
R7184 VDDA.n1719 VDDA.n1580 0.028198
R7185 VDDA.n1709 VDDA.n1578 0.028198
R7186 VDDA.n1703 VDDA.n1577 0.028198
R7187 VDDA.n1693 VDDA.n1575 0.028198
R7188 VDDA.n1689 VDDA.n1574 0.028198
R7189 VDDA.n1679 VDDA.n1572 0.028198
R7190 VDDA.n1673 VDDA.n1571 0.028198
R7191 VDDA.n1663 VDDA.n1569 0.028198
R7192 VDDA.n1659 VDDA.n1568 0.028198
R7193 VDDA.n1649 VDDA.n1566 0.028198
R7194 VDDA.n1643 VDDA.n1565 0.028198
R7195 VDDA.n1633 VDDA.n1563 0.028198
R7196 VDDA.n1629 VDDA.n1562 0.028198
R7197 VDDA.n1619 VDDA.n1560 0.028198
R7198 VDDA.n1613 VDDA.n1559 0.028198
R7199 VDDA.n1956 VDDA.n1495 0.0264451
R7200 VDDA.n1970 VDDA.n1498 0.0264451
R7201 VDDA.n1986 VDDA.n1501 0.0264451
R7202 VDDA.n2000 VDDA.n1504 0.0264451
R7203 VDDA.n2016 VDDA.n1507 0.0264451
R7204 VDDA.n2030 VDDA.n1510 0.0264451
R7205 VDDA.n2046 VDDA.n1513 0.0264451
R7206 VDDA.n2041 VDDA.n1513 0.0264451
R7207 VDDA.n2027 VDDA.n1510 0.0264451
R7208 VDDA.n2011 VDDA.n1507 0.0264451
R7209 VDDA.n1997 VDDA.n1504 0.0264451
R7210 VDDA.n1981 VDDA.n1501 0.0264451
R7211 VDDA.n1967 VDDA.n1498 0.0264451
R7212 VDDA.n1951 VDDA.n1495 0.0264451
R7213 VDDA.n1628 VDDA.n1561 0.0243392
R7214 VDDA.n1642 VDDA.n1564 0.0243392
R7215 VDDA.n1658 VDDA.n1567 0.0243392
R7216 VDDA.n1672 VDDA.n1570 0.0243392
R7217 VDDA.n1688 VDDA.n1573 0.0243392
R7218 VDDA.n1702 VDDA.n1576 0.0243392
R7219 VDDA.n1718 VDDA.n1579 0.0243392
R7220 VDDA.n2305 VDDA.n1471 0.0243392
R7221 VDDA.n2319 VDDA.n1474 0.0243392
R7222 VDDA.n2335 VDDA.n1477 0.0243392
R7223 VDDA.n2349 VDDA.n1480 0.0243392
R7224 VDDA.n2365 VDDA.n1483 0.0243392
R7225 VDDA.n2379 VDDA.n1486 0.0243392
R7226 VDDA.n2395 VDDA.n1489 0.0243392
R7227 VDDA.n84 VDDA.n23 0.0243392
R7228 VDDA.n113 VDDA.n26 0.0243392
R7229 VDDA.n72 VDDA.n29 0.0243392
R7230 VDDA.n137 VDDA.n32 0.0243392
R7231 VDDA.n60 VDDA.n35 0.0243392
R7232 VDDA.n161 VDDA.n38 0.0243392
R7233 VDDA.n48 VDDA.n41 0.0243392
R7234 VDDA.n2820 VDDA.n2819 0.0243392
R7235 VDDA.n2831 VDDA.n2793 0.0243392
R7236 VDDA.n2850 VDDA.n2849 0.0243392
R7237 VDDA.n2861 VDDA.n2781 0.0243392
R7238 VDDA.n2880 VDDA.n2879 0.0243392
R7239 VDDA.n2891 VDDA.n2769 0.0243392
R7240 VDDA.n2910 VDDA.n2909 0.0243392
R7241 VDDA.n2668 VDDA.n2593 0.0243392
R7242 VDDA.n2645 VDDA.n2596 0.0243392
R7243 VDDA.n2692 VDDA.n2599 0.0243392
R7244 VDDA.n2633 VDDA.n2602 0.0243392
R7245 VDDA.n2716 VDDA.n2605 0.0243392
R7246 VDDA.n2621 VDDA.n2608 0.0243392
R7247 VDDA.n2740 VDDA.n2611 0.0243392
R7248 VDDA.n262 VDDA.n201 0.0243392
R7249 VDDA.n291 VDDA.n204 0.0243392
R7250 VDDA.n250 VDDA.n207 0.0243392
R7251 VDDA.n315 VDDA.n210 0.0243392
R7252 VDDA.n238 VDDA.n213 0.0243392
R7253 VDDA.n339 VDDA.n216 0.0243392
R7254 VDDA.n226 VDDA.n219 0.0243392
R7255 VDDA.n426 VDDA.n425 0.0243392
R7256 VDDA.n437 VDDA.n399 0.0243392
R7257 VDDA.n456 VDDA.n455 0.0243392
R7258 VDDA.n467 VDDA.n387 0.0243392
R7259 VDDA.n486 VDDA.n485 0.0243392
R7260 VDDA.n497 VDDA.n375 0.0243392
R7261 VDDA.n516 VDDA.n515 0.0243392
R7262 VDDA.n1388 VDDA.n1313 0.0243392
R7263 VDDA.n1365 VDDA.n1316 0.0243392
R7264 VDDA.n1412 VDDA.n1319 0.0243392
R7265 VDDA.n1353 VDDA.n1322 0.0243392
R7266 VDDA.n1436 VDDA.n1325 0.0243392
R7267 VDDA.n1341 VDDA.n1328 0.0243392
R7268 VDDA.n1460 VDDA.n1331 0.0243392
R7269 VDDA.n677 VDDA.n616 0.0243392
R7270 VDDA.n706 VDDA.n619 0.0243392
R7271 VDDA.n665 VDDA.n622 0.0243392
R7272 VDDA.n730 VDDA.n625 0.0243392
R7273 VDDA.n653 VDDA.n628 0.0243392
R7274 VDDA.n754 VDDA.n631 0.0243392
R7275 VDDA.n641 VDDA.n634 0.0243392
R7276 VDDA.n1192 VDDA.n1191 0.0243392
R7277 VDDA.n1203 VDDA.n1165 0.0243392
R7278 VDDA.n1222 VDDA.n1221 0.0243392
R7279 VDDA.n1233 VDDA.n1153 0.0243392
R7280 VDDA.n1252 VDDA.n1251 0.0243392
R7281 VDDA.n1263 VDDA.n1141 0.0243392
R7282 VDDA.n1282 VDDA.n1281 0.0243392
R7283 VDDA.n1040 VDDA.n965 0.0243392
R7284 VDDA.n1017 VDDA.n968 0.0243392
R7285 VDDA.n1064 VDDA.n971 0.0243392
R7286 VDDA.n1005 VDDA.n974 0.0243392
R7287 VDDA.n1088 VDDA.n977 0.0243392
R7288 VDDA.n993 VDDA.n980 0.0243392
R7289 VDDA.n1112 VDDA.n983 0.0243392
R7290 VDDA.n852 VDDA.n792 0.0243392
R7291 VDDA.n866 VDDA.n795 0.0243392
R7292 VDDA.n882 VDDA.n798 0.0243392
R7293 VDDA.n896 VDDA.n801 0.0243392
R7294 VDDA.n912 VDDA.n804 0.0243392
R7295 VDDA.n926 VDDA.n807 0.0243392
R7296 VDDA.n942 VDDA.n810 0.0243392
R7297 VDDA.n937 VDDA.n810 0.0243392
R7298 VDDA.n923 VDDA.n807 0.0243392
R7299 VDDA.n907 VDDA.n804 0.0243392
R7300 VDDA.n893 VDDA.n801 0.0243392
R7301 VDDA.n877 VDDA.n798 0.0243392
R7302 VDDA.n863 VDDA.n795 0.0243392
R7303 VDDA.n847 VDDA.n792 0.0243392
R7304 VDDA.n990 VDDA.n983 0.0243392
R7305 VDDA.n1097 VDDA.n980 0.0243392
R7306 VDDA.n1002 VDDA.n977 0.0243392
R7307 VDDA.n1073 VDDA.n974 0.0243392
R7308 VDDA.n1014 VDDA.n971 0.0243392
R7309 VDDA.n1049 VDDA.n968 0.0243392
R7310 VDDA.n1026 VDDA.n965 0.0243392
R7311 VDDA.n1281 VDDA.n1280 0.0243392
R7312 VDDA.n1264 VDDA.n1263 0.0243392
R7313 VDDA.n1251 VDDA.n1250 0.0243392
R7314 VDDA.n1234 VDDA.n1233 0.0243392
R7315 VDDA.n1221 VDDA.n1220 0.0243392
R7316 VDDA.n1204 VDDA.n1203 0.0243392
R7317 VDDA.n1191 VDDA.n1190 0.0243392
R7318 VDDA.n763 VDDA.n634 0.0243392
R7319 VDDA.n650 VDDA.n631 0.0243392
R7320 VDDA.n739 VDDA.n628 0.0243392
R7321 VDDA.n662 VDDA.n625 0.0243392
R7322 VDDA.n715 VDDA.n622 0.0243392
R7323 VDDA.n674 VDDA.n619 0.0243392
R7324 VDDA.n691 VDDA.n616 0.0243392
R7325 VDDA.n1338 VDDA.n1331 0.0243392
R7326 VDDA.n1445 VDDA.n1328 0.0243392
R7327 VDDA.n1350 VDDA.n1325 0.0243392
R7328 VDDA.n1421 VDDA.n1322 0.0243392
R7329 VDDA.n1362 VDDA.n1319 0.0243392
R7330 VDDA.n1397 VDDA.n1316 0.0243392
R7331 VDDA.n1374 VDDA.n1313 0.0243392
R7332 VDDA.n2390 VDDA.n1489 0.0243392
R7333 VDDA.n2376 VDDA.n1486 0.0243392
R7334 VDDA.n2360 VDDA.n1483 0.0243392
R7335 VDDA.n2346 VDDA.n1480 0.0243392
R7336 VDDA.n2330 VDDA.n1477 0.0243392
R7337 VDDA.n2316 VDDA.n1474 0.0243392
R7338 VDDA.n2300 VDDA.n1471 0.0243392
R7339 VDDA.n515 VDDA.n514 0.0243392
R7340 VDDA.n498 VDDA.n497 0.0243392
R7341 VDDA.n485 VDDA.n484 0.0243392
R7342 VDDA.n468 VDDA.n467 0.0243392
R7343 VDDA.n455 VDDA.n454 0.0243392
R7344 VDDA.n438 VDDA.n437 0.0243392
R7345 VDDA.n425 VDDA.n424 0.0243392
R7346 VDDA.n348 VDDA.n219 0.0243392
R7347 VDDA.n235 VDDA.n216 0.0243392
R7348 VDDA.n324 VDDA.n213 0.0243392
R7349 VDDA.n247 VDDA.n210 0.0243392
R7350 VDDA.n300 VDDA.n207 0.0243392
R7351 VDDA.n259 VDDA.n204 0.0243392
R7352 VDDA.n276 VDDA.n201 0.0243392
R7353 VDDA.n2618 VDDA.n2611 0.0243392
R7354 VDDA.n2725 VDDA.n2608 0.0243392
R7355 VDDA.n2630 VDDA.n2605 0.0243392
R7356 VDDA.n2701 VDDA.n2602 0.0243392
R7357 VDDA.n2642 VDDA.n2599 0.0243392
R7358 VDDA.n2677 VDDA.n2596 0.0243392
R7359 VDDA.n2654 VDDA.n2593 0.0243392
R7360 VDDA.n2909 VDDA.n2908 0.0243392
R7361 VDDA.n2892 VDDA.n2891 0.0243392
R7362 VDDA.n2879 VDDA.n2878 0.0243392
R7363 VDDA.n2862 VDDA.n2861 0.0243392
R7364 VDDA.n2849 VDDA.n2848 0.0243392
R7365 VDDA.n2832 VDDA.n2831 0.0243392
R7366 VDDA.n2819 VDDA.n2818 0.0243392
R7367 VDDA.n170 VDDA.n41 0.0243392
R7368 VDDA.n57 VDDA.n38 0.0243392
R7369 VDDA.n146 VDDA.n35 0.0243392
R7370 VDDA.n69 VDDA.n32 0.0243392
R7371 VDDA.n122 VDDA.n29 0.0243392
R7372 VDDA.n81 VDDA.n26 0.0243392
R7373 VDDA.n98 VDDA.n23 0.0243392
R7374 VDDA.n1713 VDDA.n1579 0.0243392
R7375 VDDA.n1699 VDDA.n1576 0.0243392
R7376 VDDA.n1683 VDDA.n1573 0.0243392
R7377 VDDA.n1669 VDDA.n1570 0.0243392
R7378 VDDA.n1653 VDDA.n1567 0.0243392
R7379 VDDA.n1639 VDDA.n1564 0.0243392
R7380 VDDA.n1623 VDDA.n1561 0.0243392
R7381 VDDA.n2285 VDDA.n2081 0.0217373
R7382 VDDA.n2235 VDDA.n2083 0.0217373
R7383 VDDA.n2158 VDDA.n2085 0.0217373
R7384 VDDA.n2092 VDDA.n2087 0.0217373
R7385 VDDA.n2096 VDDA.n2095 0.0217373
R7386 VDDA.n2162 VDDA.n2161 0.0217373
R7387 VDDA.n2239 VDDA.n2238 0.0217373
R7388 VDDA.n2289 VDDA.n2288 0.0217373
R7389 VDDA.n2094 VDDA.n2087 0.0217373
R7390 VDDA.n2097 VDDA.n2096 0.0217373
R7391 VDDA.n2160 VDDA.n2085 0.0217373
R7392 VDDA.n2163 VDDA.n2162 0.0217373
R7393 VDDA.n2237 VDDA.n2083 0.0217373
R7394 VDDA.n2240 VDDA.n2239 0.0217373
R7395 VDDA.n2287 VDDA.n2081 0.0217373
R7396 VDDA.n2290 VDDA.n2289 0.0217373
R7397 VDDA.n2467 VDDA.n2466 0.0217373
R7398 VDDA.n2463 VDDA.n2455 0.0217373
R7399 VDDA.n2477 VDDA.n2453 0.0217373
R7400 VDDA.n2468 VDDA.n2454 0.0217373
R7401 VDDA.n2482 VDDA.n2452 0.0217373
R7402 VDDA.n2486 VDDA.n544 0.0217373
R7403 VDDA.n2481 VDDA.n2453 0.0217373
R7404 VDDA.n2479 VDDA.n2452 0.0217373
R7405 VDDA.n2477 VDDA.n2476 0.0217373
R7406 VDDA.n2467 VDDA.n2455 0.0217373
R7407 VDDA.n2464 VDDA.n2454 0.0217373
R7408 VDDA.n2536 VDDA.n2524 0.0217373
R7409 VDDA.n2547 VDDA.n2541 0.0217373
R7410 VDDA.n2933 VDDA.n2932 0.0217373
R7411 VDDA.n2930 VDDA.n185 0.0217373
R7412 VDDA.n2924 VDDA.n187 0.0217373
R7413 VDDA.n2927 VDDA.n188 0.0217373
R7414 VDDA.n2753 VDDA.n190 0.0217373
R7415 VDDA.n2756 VDDA.n191 0.0217373
R7416 VDDA.n2585 VDDA.n2584 0.0217373
R7417 VDDA.n2581 VDDA.n362 0.0217373
R7418 VDDA.n2580 VDDA.n363 0.0217373
R7419 VDDA.n2584 VDDA.n2583 0.0217373
R7420 VDDA.n2583 VDDA.n362 0.0217373
R7421 VDDA.n193 VDDA.n190 0.0217373
R7422 VDDA.n193 VDDA.n191 0.0217373
R7423 VDDA.n2758 VDDA.n187 0.0217373
R7424 VDDA.n2758 VDDA.n188 0.0217373
R7425 VDDA.n2932 VDDA.n183 0.0217373
R7426 VDDA.n185 VDDA.n183 0.0217373
R7427 VDDA.n2576 VDDA.n364 0.0217373
R7428 VDDA.n2574 VDDA.n2573 0.0217373
R7429 VDDA.n2571 VDDA.n534 0.0217373
R7430 VDDA.n530 VDDA.n363 0.0217373
R7431 VDDA.n2576 VDDA.n2575 0.0217373
R7432 VDDA.n2555 VDDA.n537 0.0217373
R7433 VDDA.n2573 VDDA.n532 0.0217373
R7434 VDDA.n534 VDDA.n532 0.0217373
R7435 VDDA.n2512 VDDA.n2511 0.0217373
R7436 VDDA.n2515 VDDA.n539 0.0217373
R7437 VDDA.n2551 VDDA.n538 0.0217373
R7438 VDDA.n2539 VDDA.n2518 0.0217373
R7439 VDDA.n2523 VDDA.n2521 0.0217373
R7440 VDDA.n2516 VDDA.n537 0.0217373
R7441 VDDA.n2551 VDDA.n2550 0.0217373
R7442 VDDA.n2541 VDDA.n2519 0.0217373
R7443 VDDA.n2540 VDDA.n2539 0.0217373
R7444 VDDA.n2524 VDDA.n2522 0.0217373
R7445 VDDA.n2445 VDDA.n545 0.0217373
R7446 VDDA.n2511 VDDA.n2494 0.0217373
R7447 VDDA.n2494 VDDA.n539 0.0217373
R7448 VDDA.n2484 VDDA.n2483 0.0217373
R7449 VDDA.n2441 VDDA.n546 0.0217373
R7450 VDDA.n2439 VDDA.n2438 0.0217373
R7451 VDDA.n2436 VDDA.n566 0.0217373
R7452 VDDA.n595 VDDA.n568 0.0217373
R7453 VDDA.n585 VDDA.n571 0.0217373
R7454 VDDA.n562 VDDA.n545 0.0217373
R7455 VDDA.n2441 VDDA.n2440 0.0217373
R7456 VDDA.n597 VDDA.n569 0.0217373
R7457 VDDA.n596 VDDA.n595 0.0217373
R7458 VDDA.n586 VDDA.n572 0.0217373
R7459 VDDA.n2420 VDDA.n602 0.0217373
R7460 VDDA.n2438 VDDA.n564 0.0217373
R7461 VDDA.n566 VDDA.n564 0.0217373
R7462 VDDA.n2411 VDDA.n2410 0.0217373
R7463 VDDA.n2414 VDDA.n604 0.0217373
R7464 VDDA.n2416 VDDA.n603 0.0217373
R7465 VDDA.n2415 VDDA.n602 0.0217373
R7466 VDDA.n1305 VDDA.n1304 0.0217373
R7467 VDDA.n1301 VDDA.n777 0.0217373
R7468 VDDA.n1296 VDDA.n779 0.0217373
R7469 VDDA.n1299 VDDA.n780 0.0217373
R7470 VDDA.n1125 VDDA.n782 0.0217373
R7471 VDDA.n1128 VDDA.n783 0.0217373
R7472 VDDA.n953 VDDA.n784 0.0217373
R7473 VDDA.n785 VDDA.n782 0.0217373
R7474 VDDA.n785 VDDA.n783 0.0217373
R7475 VDDA.n1130 VDDA.n779 0.0217373
R7476 VDDA.n1130 VDDA.n780 0.0217373
R7477 VDDA.n1304 VDDA.n1303 0.0217373
R7478 VDDA.n1303 VDDA.n777 0.0217373
R7479 VDDA.n2410 VDDA.n607 0.0217373
R7480 VDDA.n607 VDDA.n604 0.0217373
R7481 VDDA.n955 VDDA.n954 0.0217373
R7482 VDDA.n953 VDDA.n952 0.0217373
R7483 VDDA.n2287 VDDA.n2082 0.0217373
R7484 VDDA.n2237 VDDA.n2084 0.0217373
R7485 VDDA.n2160 VDDA.n2086 0.0217373
R7486 VDDA.n2094 VDDA.n2088 0.0217373
R7487 VDDA.n2095 VDDA.n2093 0.0217373
R7488 VDDA.n2161 VDDA.n2159 0.0217373
R7489 VDDA.n2238 VDDA.n2236 0.0217373
R7490 VDDA.n2288 VDDA.n2286 0.0217373
R7491 VDDA.n2159 VDDA.n2098 0.0217373
R7492 VDDA.n2236 VDDA.n2164 0.0217373
R7493 VDDA.n2286 VDDA.n2241 0.0217373
R7494 VDDA.n572 VDDA.n570 0.0217373
R7495 VDDA.n569 VDDA.n567 0.0217373
R7496 VDDA.n2480 VDDA.n2478 0.0217373
R7497 VDDA.n2480 VDDA.n2479 0.0217373
R7498 VDDA.n2465 VDDA.n2464 0.0217373
R7499 VDDA.n2522 VDDA.n2520 0.0217373
R7500 VDDA.n2519 VDDA.n2517 0.0217373
R7501 VDDA.n2577 VDDA.n530 0.0217373
R7502 VDDA.n2582 VDDA.n360 0.0217373
R7503 VDDA.n2755 VDDA.n2754 0.0217373
R7504 VDDA.n2926 VDDA.n2925 0.0217373
R7505 VDDA.n2929 VDDA.n182 0.0217373
R7506 VDDA.n361 VDDA.n360 0.0217373
R7507 VDDA.n2754 VDDA.n189 0.0217373
R7508 VDDA.n2925 VDDA.n186 0.0217373
R7509 VDDA.n184 VDDA.n182 0.0217373
R7510 VDDA.n2579 VDDA.n364 0.0217373
R7511 VDDA.n2579 VDDA.n2578 0.0217373
R7512 VDDA.n2552 VDDA.n2516 0.0217373
R7513 VDDA.n2570 VDDA.n531 0.0217373
R7514 VDDA.n533 VDDA.n531 0.0217373
R7515 VDDA.n2554 VDDA.n538 0.0217373
R7516 VDDA.n2548 VDDA.n2518 0.0217373
R7517 VDDA.n2537 VDDA.n2521 0.0217373
R7518 VDDA.n2554 VDDA.n2553 0.0217373
R7519 VDDA.n2549 VDDA.n2548 0.0217373
R7520 VDDA.n2538 VDDA.n2537 0.0217373
R7521 VDDA.n2442 VDDA.n562 0.0217373
R7522 VDDA.n2514 VDDA.n2513 0.0217373
R7523 VDDA.n2513 VDDA.n2495 0.0217373
R7524 VDDA.n2444 VDDA.n546 0.0217373
R7525 VDDA.n598 VDDA.n568 0.0217373
R7526 VDDA.n587 VDDA.n571 0.0217373
R7527 VDDA.n2444 VDDA.n2443 0.0217373
R7528 VDDA.n599 VDDA.n598 0.0217373
R7529 VDDA.n594 VDDA.n567 0.0217373
R7530 VDDA.n588 VDDA.n587 0.0217373
R7531 VDDA.n584 VDDA.n570 0.0217373
R7532 VDDA.n2417 VDDA.n2415 0.0217373
R7533 VDDA.n2435 VDDA.n563 0.0217373
R7534 VDDA.n565 VDDA.n563 0.0217373
R7535 VDDA.n2419 VDDA.n603 0.0217373
R7536 VDDA.n2419 VDDA.n2418 0.0217373
R7537 VDDA.n952 VDDA.n951 0.0217373
R7538 VDDA.n1127 VDDA.n1126 0.0217373
R7539 VDDA.n1298 VDDA.n1297 0.0217373
R7540 VDDA.n1302 VDDA.n775 0.0217373
R7541 VDDA.n2413 VDDA.n2412 0.0217373
R7542 VDDA.n1126 VDDA.n781 0.0217373
R7543 VDDA.n1297 VDDA.n778 0.0217373
R7544 VDDA.n776 VDDA.n775 0.0217373
R7545 VDDA.n2412 VDDA.n608 0.0217373
R7546 VDDA.n956 VDDA.n955 0.0217373
R7547 VDDA.n957 VDDA.n956 0.0217373
R7548 VDDA VDDA.n3124 0.0164359
R7549 VDDA.n1909 VDDA.n1908 0.0152446
R7550 VDDA.n1907 VDDA.n1906 0.0152446
R7551 VDDA.n1905 VDDA.n1904 0.0152446
R7552 VDDA.n1895 VDDA.n1894 0.0152446
R7553 VDDA.n1742 VDDA.n1738 0.0152446
R7554 VDDA.n1888 VDDA.n1743 0.0152446
R7555 VDDA.n1878 VDDA.n1749 0.0152446
R7556 VDDA.n1877 VDDA.n1876 0.0152446
R7557 VDDA.n1875 VDDA.n1874 0.0152446
R7558 VDDA.n1865 VDDA.n1864 0.0152446
R7559 VDDA.n1760 VDDA.n1756 0.0152446
R7560 VDDA.n1858 VDDA.n1761 0.0152446
R7561 VDDA.n1848 VDDA.n1767 0.0152446
R7562 VDDA.n1847 VDDA.n1846 0.0152446
R7563 VDDA.n1845 VDDA.n1844 0.0152446
R7564 VDDA.n1835 VDDA.n1834 0.0152446
R7565 VDDA.n1778 VDDA.n1774 0.0152446
R7566 VDDA.n1828 VDDA.n1779 0.0152446
R7567 VDDA.n1818 VDDA.n1785 0.0152446
R7568 VDDA.n1817 VDDA.n1816 0.0152446
R7569 VDDA.n1815 VDDA.n1814 0.0152446
R7570 VDDA.n1805 VDDA.n1804 0.0152446
R7571 VDDA.n1795 VDDA.n1792 0.0152446
R7572 VDDA.n1798 VDDA.n1796 0.0152446
R7573 VDDA.n1796 VDDA.n1795 0.0152446
R7574 VDDA.n1804 VDDA.n1792 0.0152446
R7575 VDDA.n1806 VDDA.n1805 0.0152446
R7576 VDDA.n1816 VDDA.n1815 0.0152446
R7577 VDDA.n1818 VDDA.n1817 0.0152446
R7578 VDDA.n1785 VDDA.n1784 0.0152446
R7579 VDDA.n1779 VDDA.n1778 0.0152446
R7580 VDDA.n1834 VDDA.n1774 0.0152446
R7581 VDDA.n1836 VDDA.n1835 0.0152446
R7582 VDDA.n1846 VDDA.n1845 0.0152446
R7583 VDDA.n1848 VDDA.n1847 0.0152446
R7584 VDDA.n1767 VDDA.n1766 0.0152446
R7585 VDDA.n1761 VDDA.n1760 0.0152446
R7586 VDDA.n1864 VDDA.n1756 0.0152446
R7587 VDDA.n1866 VDDA.n1865 0.0152446
R7588 VDDA.n1876 VDDA.n1875 0.0152446
R7589 VDDA.n1878 VDDA.n1877 0.0152446
R7590 VDDA.n1749 VDDA.n1748 0.0152446
R7591 VDDA.n1743 VDDA.n1742 0.0152446
R7592 VDDA.n1894 VDDA.n1738 0.0152446
R7593 VDDA.n1896 VDDA.n1895 0.0152446
R7594 VDDA.n1906 VDDA.n1905 0.0152446
R7595 VDDA.n1908 VDDA.n1907 0.0152446
R7596 VDDA.n1910 VDDA.n1909 0.0152446
R7597 VDDA.n1910 VDDA.n1556 0.0142311
R7598 VDDA.n1736 VDDA.n1731 0.0142311
R7599 VDDA.n1897 VDDA.n1896 0.0142311
R7600 VDDA.n1887 VDDA.n1886 0.0142311
R7601 VDDA.n1748 VDDA.n1744 0.0142311
R7602 VDDA.n1754 VDDA.n1750 0.0142311
R7603 VDDA.n1867 VDDA.n1866 0.0142311
R7604 VDDA.n1857 VDDA.n1856 0.0142311
R7605 VDDA.n1766 VDDA.n1762 0.0142311
R7606 VDDA.n1772 VDDA.n1768 0.0142311
R7607 VDDA.n1837 VDDA.n1836 0.0142311
R7608 VDDA.n1827 VDDA.n1826 0.0142311
R7609 VDDA.n1784 VDDA.n1780 0.0142311
R7610 VDDA.n1790 VDDA.n1786 0.0142311
R7611 VDDA.n1807 VDDA.n1806 0.0142311
R7612 VDDA.n1797 VDDA.n1794 0.0142311
R7613 VDDA.n1798 VDDA.n1797 0.0142311
R7614 VDDA.n1808 VDDA.n1807 0.0142311
R7615 VDDA.n1814 VDDA.n1786 0.0142311
R7616 VDDA.n1824 VDDA.n1780 0.0142311
R7617 VDDA.n1828 VDDA.n1827 0.0142311
R7618 VDDA.n1838 VDDA.n1837 0.0142311
R7619 VDDA.n1844 VDDA.n1768 0.0142311
R7620 VDDA.n1854 VDDA.n1762 0.0142311
R7621 VDDA.n1858 VDDA.n1857 0.0142311
R7622 VDDA.n1868 VDDA.n1867 0.0142311
R7623 VDDA.n1874 VDDA.n1750 0.0142311
R7624 VDDA.n1884 VDDA.n1744 0.0142311
R7625 VDDA.n1888 VDDA.n1887 0.0142311
R7626 VDDA.n1898 VDDA.n1897 0.0142311
R7627 VDDA.n1904 VDDA.n1731 0.0142311
R7628 VDDA.n1557 VDDA.n1556 0.0142311
R7629 VDDA.n1729 VDDA.n1728 0.0141594
R7630 VDDA.n1898 VDDA.n1737 0.0132169
R7631 VDDA.n1885 VDDA.n1884 0.0132169
R7632 VDDA.n1868 VDDA.n1755 0.0132169
R7633 VDDA.n1855 VDDA.n1854 0.0132169
R7634 VDDA.n1838 VDDA.n1773 0.0132169
R7635 VDDA.n1825 VDDA.n1824 0.0132169
R7636 VDDA.n1808 VDDA.n1791 0.0132169
R7637 VDDA.n1791 VDDA.n1790 0.0132169
R7638 VDDA.n1826 VDDA.n1825 0.0132169
R7639 VDDA.n1773 VDDA.n1772 0.0132169
R7640 VDDA.n1856 VDDA.n1855 0.0132169
R7641 VDDA.n1755 VDDA.n1754 0.0132169
R7642 VDDA.n1886 VDDA.n1885 0.0132169
R7643 VDDA.n1737 VDDA.n1736 0.0132169
R7644 VDDA.n2406 VDDA.n1309 0.0107812
R7645 VDDA.n2589 VDDA.n197 0.0107812
R7646 VDDA.n1728 VDDA.n197 0.00894531
R7647 VDDA.n2406 VDDA.n2405 0.00887187
R7648 VDDA.n1121 VDDA.n961 0.00564062
R7649 VDDA.n1121 VDDA.n612 0.00564062
R7650 VDDA.n1309 VDDA.n612 0.00564062
R7651 VDDA.n2749 VDDA.n2589 0.00564062
R7652 VDDA.n2749 VDDA.n19 0.00564062
R7653 VDDA.n2937 VDDA.n19 0.00564062
R7654 VDDA.n2056 VDDA.n1516 0.00211562
R7655 VDDA.n3025 VDDA.n3023 0.00202782
R7656 VDDA.n3023 VDDA.n2955 0.00202782
R7657 VDDA.n2974 VDDA.n0 0.00166081
R7658 VDDA.n2973 VDDA.n2971 0.00166081
R7659 VDDA.n2977 VDDA.n2975 0.00166081
R7660 VDDA.n2976 VDDA.n2970 0.00166081
R7661 VDDA.n2980 VDDA.n2978 0.00166081
R7662 VDDA.n2979 VDDA.n2969 0.00166081
R7663 VDDA.n2983 VDDA.n2981 0.00166081
R7664 VDDA.n2982 VDDA.n2968 0.00166081
R7665 VDDA.n2986 VDDA.n2984 0.00166081
R7666 VDDA.n2985 VDDA.n2967 0.00166081
R7667 VDDA.n2989 VDDA.n2987 0.00166081
R7668 VDDA.n2988 VDDA.n2966 0.00166081
R7669 VDDA.n2992 VDDA.n2990 0.00166081
R7670 VDDA.n2991 VDDA.n2965 0.00166081
R7671 VDDA.n2995 VDDA.n2993 0.00166081
R7672 VDDA.n2994 VDDA.n2964 0.00166081
R7673 VDDA.n2998 VDDA.n2996 0.00166081
R7674 VDDA.n2997 VDDA.n2963 0.00166081
R7675 VDDA.n3001 VDDA.n2999 0.00166081
R7676 VDDA.n3000 VDDA.n2962 0.00166081
R7677 VDDA.n3004 VDDA.n3002 0.00166081
R7678 VDDA.n3003 VDDA.n2961 0.00166081
R7679 VDDA.n3007 VDDA.n3005 0.00166081
R7680 VDDA.n3006 VDDA.n2960 0.00166081
R7681 VDDA.n3010 VDDA.n3008 0.00166081
R7682 VDDA.n3009 VDDA.n2959 0.00166081
R7683 VDDA.n3013 VDDA.n3011 0.00166081
R7684 VDDA.n3012 VDDA.n2958 0.00166081
R7685 VDDA.n3016 VDDA.n3014 0.00166081
R7686 VDDA.n3015 VDDA.n2957 0.00166081
R7687 VDDA.n3019 VDDA.n3017 0.00166081
R7688 VDDA.n3018 VDDA.n2956 0.00166081
R7689 VDDA.n3022 VDDA.n3020 0.00166081
R7690 VDDA.n3021 VDDA.n2955 0.00166081
R7691 VDDA.n3024 VDDA.n2954 0.00166081
R7692 VDDA.n3028 VDDA.n3026 0.00166081
R7693 VDDA.n3027 VDDA.n2953 0.00166081
R7694 VDDA.n3031 VDDA.n3029 0.00166081
R7695 VDDA.n3030 VDDA.n2952 0.00166081
R7696 VDDA.n3034 VDDA.n3032 0.00166081
R7697 VDDA.n3033 VDDA.n2951 0.00166081
R7698 VDDA.n3037 VDDA.n3035 0.00166081
R7699 VDDA.n3036 VDDA.n2950 0.00166081
R7700 VDDA.n3040 VDDA.n3038 0.00166081
R7701 VDDA.n3039 VDDA.n2949 0.00166081
R7702 VDDA.n3043 VDDA.n3041 0.00166081
R7703 VDDA.n3042 VDDA.n2948 0.00166081
R7704 VDDA.n3046 VDDA.n3044 0.00166081
R7705 VDDA.n3045 VDDA.n2947 0.00166081
R7706 VDDA.n3049 VDDA.n3047 0.00166081
R7707 VDDA.n3048 VDDA.n2946 0.00166081
R7708 VDDA.n3052 VDDA.n3050 0.00166081
R7709 VDDA.n3051 VDDA.n2945 0.00166081
R7710 VDDA.n3055 VDDA.n3053 0.00166081
R7711 VDDA.n3054 VDDA.n2944 0.00166081
R7712 VDDA.n3058 VDDA.n3056 0.00166081
R7713 VDDA.n3057 VDDA.n2943 0.00166081
R7714 VDDA.n3061 VDDA.n3059 0.00166081
R7715 VDDA.n3060 VDDA.n2942 0.00166081
R7716 VDDA.n3064 VDDA.n3062 0.00166081
R7717 VDDA.n3063 VDDA.n2941 0.00166081
R7718 VDDA.n3067 VDDA.n3065 0.00166081
R7719 VDDA.n3066 VDDA.n2940 0.00166081
R7720 VDDA.n3070 VDDA.n3068 0.00166081
R7721 VDDA.n3069 VDDA.n2939 0.00166081
R7722 VDDA.n3073 VDDA.n3071 0.00166081
R7723 VDDA.n3072 VDDA.n2938 0.00166081
R7724 VDDA.n3122 VDDA.n3074 0.00166081
R7725 VDDA.n3124 VDDA.n0 0.00166081
R7726 VDDA.n2974 VDDA.n2973 0.00166081
R7727 VDDA.n2975 VDDA.n2971 0.00166081
R7728 VDDA.n2977 VDDA.n2976 0.00166081
R7729 VDDA.n2978 VDDA.n2970 0.00166081
R7730 VDDA.n2980 VDDA.n2979 0.00166081
R7731 VDDA.n2981 VDDA.n2969 0.00166081
R7732 VDDA.n2983 VDDA.n2982 0.00166081
R7733 VDDA.n2984 VDDA.n2968 0.00166081
R7734 VDDA.n2986 VDDA.n2985 0.00166081
R7735 VDDA.n2987 VDDA.n2967 0.00166081
R7736 VDDA.n2989 VDDA.n2988 0.00166081
R7737 VDDA.n2990 VDDA.n2966 0.00166081
R7738 VDDA.n2992 VDDA.n2991 0.00166081
R7739 VDDA.n2993 VDDA.n2965 0.00166081
R7740 VDDA.n2995 VDDA.n2994 0.00166081
R7741 VDDA.n2996 VDDA.n2964 0.00166081
R7742 VDDA.n2998 VDDA.n2997 0.00166081
R7743 VDDA.n2999 VDDA.n2963 0.00166081
R7744 VDDA.n3001 VDDA.n3000 0.00166081
R7745 VDDA.n3002 VDDA.n2962 0.00166081
R7746 VDDA.n3004 VDDA.n3003 0.00166081
R7747 VDDA.n3005 VDDA.n2961 0.00166081
R7748 VDDA.n3007 VDDA.n3006 0.00166081
R7749 VDDA.n3008 VDDA.n2960 0.00166081
R7750 VDDA.n3010 VDDA.n3009 0.00166081
R7751 VDDA.n3011 VDDA.n2959 0.00166081
R7752 VDDA.n3013 VDDA.n3012 0.00166081
R7753 VDDA.n3014 VDDA.n2958 0.00166081
R7754 VDDA.n3016 VDDA.n3015 0.00166081
R7755 VDDA.n3017 VDDA.n2957 0.00166081
R7756 VDDA.n3019 VDDA.n3018 0.00166081
R7757 VDDA.n3020 VDDA.n2956 0.00166081
R7758 VDDA.n3022 VDDA.n3021 0.00166081
R7759 VDDA.n3025 VDDA.n3024 0.00166081
R7760 VDDA.n3026 VDDA.n2954 0.00166081
R7761 VDDA.n3028 VDDA.n3027 0.00166081
R7762 VDDA.n3029 VDDA.n2953 0.00166081
R7763 VDDA.n3031 VDDA.n3030 0.00166081
R7764 VDDA.n3032 VDDA.n2952 0.00166081
R7765 VDDA.n3034 VDDA.n3033 0.00166081
R7766 VDDA.n3035 VDDA.n2951 0.00166081
R7767 VDDA.n3037 VDDA.n3036 0.00166081
R7768 VDDA.n3038 VDDA.n2950 0.00166081
R7769 VDDA.n3040 VDDA.n3039 0.00166081
R7770 VDDA.n3041 VDDA.n2949 0.00166081
R7771 VDDA.n3043 VDDA.n3042 0.00166081
R7772 VDDA.n3044 VDDA.n2948 0.00166081
R7773 VDDA.n3046 VDDA.n3045 0.00166081
R7774 VDDA.n3047 VDDA.n2947 0.00166081
R7775 VDDA.n3049 VDDA.n3048 0.00166081
R7776 VDDA.n3050 VDDA.n2946 0.00166081
R7777 VDDA.n3052 VDDA.n3051 0.00166081
R7778 VDDA.n3053 VDDA.n2945 0.00166081
R7779 VDDA.n3055 VDDA.n3054 0.00166081
R7780 VDDA.n3056 VDDA.n2944 0.00166081
R7781 VDDA.n3058 VDDA.n3057 0.00166081
R7782 VDDA.n3059 VDDA.n2943 0.00166081
R7783 VDDA.n3061 VDDA.n3060 0.00166081
R7784 VDDA.n3062 VDDA.n2942 0.00166081
R7785 VDDA.n3064 VDDA.n3063 0.00166081
R7786 VDDA.n3065 VDDA.n2941 0.00166081
R7787 VDDA.n3067 VDDA.n3066 0.00166081
R7788 VDDA.n3068 VDDA.n2940 0.00166081
R7789 VDDA.n3070 VDDA.n3069 0.00166081
R7790 VDDA.n3071 VDDA.n2939 0.00166081
R7791 VDDA.n3073 VDDA.n3072 0.00166081
R7792 VDDA.n3074 VDDA.n2938 0.00166081
R7793 VDDA.t53 VDDA.n1606 0.00152174
R7794 VDDA.t50 VDDA.n1607 0.00152174
R7795 VDDA.t188 VDDA.n1608 0.00152174
R7796 VDDA.t169 VDDA.n1609 0.00152174
R7797 VDDA.t46 VDDA.n1610 0.00152174
R7798 VDDA.n1729 VDDA.n1516 0.00138125
R7799 VDDA.n3076 VDDA.n3075 0.00133044
R7800 VDDA.n3076 VDDA.n1 0.00133044
R7801 VDDA.n3120 VDDA.n3077 0.00133044
R7802 VDDA.n3077 VDDA.n2 0.00133044
R7803 VDDA.n3118 VDDA.n3078 0.00133044
R7804 VDDA.n3078 VDDA.n3 0.00133044
R7805 VDDA.n3116 VDDA.n3079 0.00133044
R7806 VDDA.n3079 VDDA.n4 0.00133044
R7807 VDDA.n3114 VDDA.n3080 0.00133044
R7808 VDDA.n3080 VDDA.n5 0.00133044
R7809 VDDA.n3112 VDDA.n3081 0.00133044
R7810 VDDA.n3081 VDDA.n6 0.00133044
R7811 VDDA.n3110 VDDA.n3082 0.00133044
R7812 VDDA.n3082 VDDA.n7 0.00133044
R7813 VDDA.n3108 VDDA.n3083 0.00133044
R7814 VDDA.n3083 VDDA.n8 0.00133044
R7815 VDDA.n3106 VDDA.n3084 0.00133044
R7816 VDDA.n3084 VDDA.n9 0.00133044
R7817 VDDA.n3104 VDDA.n3085 0.00133044
R7818 VDDA.n3085 VDDA.n10 0.00133044
R7819 VDDA.n3102 VDDA.n3086 0.00133044
R7820 VDDA.n3086 VDDA.n11 0.00133044
R7821 VDDA.n3100 VDDA.n3087 0.00133044
R7822 VDDA.n3087 VDDA.n12 0.00133044
R7823 VDDA.n3098 VDDA.n3088 0.00133044
R7824 VDDA.n3088 VDDA.n13 0.00133044
R7825 VDDA.n3096 VDDA.n3089 0.00133044
R7826 VDDA.n3089 VDDA.n14 0.00133044
R7827 VDDA.n3094 VDDA.n3090 0.00133044
R7828 VDDA.n3090 VDDA.n15 0.00133044
R7829 VDDA.n3092 VDDA.n16 0.00133044
R7830 VDDA.n3091 VDDA.n17 0.00133044
R7831 VDDA.n3093 VDDA.n15 0.00133044
R7832 VDDA.n3095 VDDA.n14 0.00133044
R7833 VDDA.n3097 VDDA.n13 0.00133044
R7834 VDDA.n3099 VDDA.n12 0.00133044
R7835 VDDA.n3101 VDDA.n11 0.00133044
R7836 VDDA.n3103 VDDA.n10 0.00133044
R7837 VDDA.n3105 VDDA.n9 0.00133044
R7838 VDDA.n3107 VDDA.n8 0.00133044
R7839 VDDA.n3109 VDDA.n7 0.00133044
R7840 VDDA.n3111 VDDA.n6 0.00133044
R7841 VDDA.n3113 VDDA.n5 0.00133044
R7842 VDDA.n3115 VDDA.n4 0.00133044
R7843 VDDA.n3117 VDDA.n3 0.00133044
R7844 VDDA.n3119 VDDA.n2 0.00133044
R7845 VDDA.n3121 VDDA.n1 0.00133044
R7846 VDDA.n3093 VDDA.n3092 0.00133044
R7847 VDDA.n3095 VDDA.n3094 0.00133044
R7848 VDDA.n3097 VDDA.n3096 0.00133044
R7849 VDDA.n3099 VDDA.n3098 0.00133044
R7850 VDDA.n3101 VDDA.n3100 0.00133044
R7851 VDDA.n3103 VDDA.n3102 0.00133044
R7852 VDDA.n3105 VDDA.n3104 0.00133044
R7853 VDDA.n3107 VDDA.n3106 0.00133044
R7854 VDDA.n3109 VDDA.n3108 0.00133044
R7855 VDDA.n3111 VDDA.n3110 0.00133044
R7856 VDDA.n3113 VDDA.n3112 0.00133044
R7857 VDDA.n3115 VDDA.n3114 0.00133044
R7858 VDDA.n3117 VDDA.n3116 0.00133044
R7859 VDDA.n3119 VDDA.n3118 0.00133044
R7860 VDDA.n3121 VDDA.n3120 0.00133044
R7861 VDDA.n3075 VDDA.n18 0.00133044
R7862 VDDA.n3091 VDDA.n16 0.00133044
R7863 VDDA.n3123 VDDA.n2972 0.00116094
R7864 VDDA.n2972 VDDA.n18 0.00116094
R7865 two_stage_opamp_dummy_magic_26_0.Vb1.n1 two_stage_opamp_dummy_magic_26_0.Vb1.t28 484.212
R7866 two_stage_opamp_dummy_magic_26_0.Vb1.n1 two_stage_opamp_dummy_magic_26_0.Vb1.t18 484.212
R7867 two_stage_opamp_dummy_magic_26_0.Vb1.n1 two_stage_opamp_dummy_magic_26_0.Vb1.t26 484.212
R7868 two_stage_opamp_dummy_magic_26_0.Vb1.n1 two_stage_opamp_dummy_magic_26_0.Vb1.t17 484.212
R7869 two_stage_opamp_dummy_magic_26_0.Vb1.n2 two_stage_opamp_dummy_magic_26_0.Vb1.t25 484.212
R7870 two_stage_opamp_dummy_magic_26_0.Vb1.n2 two_stage_opamp_dummy_magic_26_0.Vb1.t15 484.212
R7871 two_stage_opamp_dummy_magic_26_0.Vb1.n2 two_stage_opamp_dummy_magic_26_0.Vb1.t31 484.212
R7872 two_stage_opamp_dummy_magic_26_0.Vb1.n2 two_stage_opamp_dummy_magic_26_0.Vb1.t16 484.212
R7873 two_stage_opamp_dummy_magic_26_0.Vb1.n2 two_stage_opamp_dummy_magic_26_0.Vb1.t24 484.212
R7874 two_stage_opamp_dummy_magic_26_0.Vb1.n2 two_stage_opamp_dummy_magic_26_0.Vb1.t14 484.212
R7875 two_stage_opamp_dummy_magic_26_0.Vb1.n3 two_stage_opamp_dummy_magic_26_0.Vb1.t12 484.212
R7876 two_stage_opamp_dummy_magic_26_0.Vb1.n3 two_stage_opamp_dummy_magic_26_0.Vb1.t22 484.212
R7877 two_stage_opamp_dummy_magic_26_0.Vb1.n3 two_stage_opamp_dummy_magic_26_0.Vb1.t32 484.212
R7878 two_stage_opamp_dummy_magic_26_0.Vb1.n3 two_stage_opamp_dummy_magic_26_0.Vb1.t20 484.212
R7879 two_stage_opamp_dummy_magic_26_0.Vb1.n4 two_stage_opamp_dummy_magic_26_0.Vb1.t29 484.212
R7880 two_stage_opamp_dummy_magic_26_0.Vb1.n4 two_stage_opamp_dummy_magic_26_0.Vb1.t21 484.212
R7881 two_stage_opamp_dummy_magic_26_0.Vb1.n4 two_stage_opamp_dummy_magic_26_0.Vb1.t30 484.212
R7882 two_stage_opamp_dummy_magic_26_0.Vb1.n4 two_stage_opamp_dummy_magic_26_0.Vb1.t19 484.212
R7883 two_stage_opamp_dummy_magic_26_0.Vb1.n4 two_stage_opamp_dummy_magic_26_0.Vb1.t27 484.212
R7884 two_stage_opamp_dummy_magic_26_0.Vb1.n4 two_stage_opamp_dummy_magic_26_0.Vb1.t13 484.212
R7885 two_stage_opamp_dummy_magic_26_0.Vb1.n8 two_stage_opamp_dummy_magic_26_0.Vb1.t8 449.868
R7886 two_stage_opamp_dummy_magic_26_0.Vb1.n7 two_stage_opamp_dummy_magic_26_0.Vb1.t10 449.868
R7887 two_stage_opamp_dummy_magic_26_0.Vb1.n8 two_stage_opamp_dummy_magic_26_0.Vb1.t4 273.134
R7888 two_stage_opamp_dummy_magic_26_0.Vb1.n7 two_stage_opamp_dummy_magic_26_0.Vb1.t6 273.134
R7889 two_stage_opamp_dummy_magic_26_0.Vb1.n11 two_stage_opamp_dummy_magic_26_0.Vb1.t23 161.363
R7890 two_stage_opamp_dummy_magic_26_0.Vb1.n5 two_stage_opamp_dummy_magic_26_0.Vb1.n9 161.3
R7891 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.Vb1.n6 151.863
R7892 two_stage_opamp_dummy_magic_26_0.Vb1.n13 two_stage_opamp_dummy_magic_26_0.Vb1.n12 49.3505
R7893 two_stage_opamp_dummy_magic_26_0.Vb1.n5 two_stage_opamp_dummy_magic_26_0.Vb1.n10 49.3505
R7894 two_stage_opamp_dummy_magic_26_0.Vb1.n16 two_stage_opamp_dummy_magic_26_0.Vb1.n15 49.3505
R7895 two_stage_opamp_dummy_magic_26_0.Vb1.n9 two_stage_opamp_dummy_magic_26_0.Vb1.n8 45.5227
R7896 two_stage_opamp_dummy_magic_26_0.Vb1.n9 two_stage_opamp_dummy_magic_26_0.Vb1.n7 45.5227
R7897 two_stage_opamp_dummy_magic_26_0.Vb1.n0 two_stage_opamp_dummy_magic_26_0.Vb1.n4 21.6489
R7898 two_stage_opamp_dummy_magic_26_0.Vb1.n1 two_stage_opamp_dummy_magic_26_0.Vb1.n0 21.3677
R7899 two_stage_opamp_dummy_magic_26_0.Vb1.n6 two_stage_opamp_dummy_magic_26_0.Vb1.t3 19.7005
R7900 two_stage_opamp_dummy_magic_26_0.Vb1.n6 two_stage_opamp_dummy_magic_26_0.Vb1.t2 19.7005
R7901 two_stage_opamp_dummy_magic_26_0.Vb1.n12 two_stage_opamp_dummy_magic_26_0.Vb1.t1 16.0005
R7902 two_stage_opamp_dummy_magic_26_0.Vb1.n12 two_stage_opamp_dummy_magic_26_0.Vb1.t11 16.0005
R7903 two_stage_opamp_dummy_magic_26_0.Vb1.n10 two_stage_opamp_dummy_magic_26_0.Vb1.t7 16.0005
R7904 two_stage_opamp_dummy_magic_26_0.Vb1.n10 two_stage_opamp_dummy_magic_26_0.Vb1.t5 16.0005
R7905 two_stage_opamp_dummy_magic_26_0.Vb1.n15 two_stage_opamp_dummy_magic_26_0.Vb1.t9 16.0005
R7906 two_stage_opamp_dummy_magic_26_0.Vb1.n15 two_stage_opamp_dummy_magic_26_0.Vb1.t0 16.0005
R7907 two_stage_opamp_dummy_magic_26_0.Vb1.n16 two_stage_opamp_dummy_magic_26_0.Vb1.n14 5.28175
R7908 two_stage_opamp_dummy_magic_26_0.Vb1.n14 two_stage_opamp_dummy_magic_26_0.Vb1.n13 5.28175
R7909 two_stage_opamp_dummy_magic_26_0.Vb1.n5 two_stage_opamp_dummy_magic_26_0.Vb1.n0 5.188
R7910 two_stage_opamp_dummy_magic_26_0.Vb1.n0 two_stage_opamp_dummy_magic_26_0.Vb1.n16 4.938
R7911 two_stage_opamp_dummy_magic_26_0.Vb1.n13 two_stage_opamp_dummy_magic_26_0.Vb1.n0 4.938
R7912 two_stage_opamp_dummy_magic_26_0.Vb1.n14 two_stage_opamp_dummy_magic_26_0.Vb1.n11 2.23569
R7913 two_stage_opamp_dummy_magic_26_0.Vb1.n4 two_stage_opamp_dummy_magic_26_0.Vb1.n3 1.54738
R7914 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.Vb1.n2 1.36769
R7915 two_stage_opamp_dummy_magic_26_0.Vb1.n2 two_stage_opamp_dummy_magic_26_0.Vb1.n1 1.03175
R7916 two_stage_opamp_dummy_magic_26_0.Vb1.n11 two_stage_opamp_dummy_magic_26_0.Vb1.n5 0.937224
R7917 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.Vb1.n3 0.852062
R7918 two_stage_opamp_dummy_magic_26_0.X.n76 two_stage_opamp_dummy_magic_26_0.X.t41 1172.87
R7919 two_stage_opamp_dummy_magic_26_0.X.n72 two_stage_opamp_dummy_magic_26_0.X.t37 1172.87
R7920 two_stage_opamp_dummy_magic_26_0.X.n76 two_stage_opamp_dummy_magic_26_0.X.t28 996.134
R7921 two_stage_opamp_dummy_magic_26_0.X.n77 two_stage_opamp_dummy_magic_26_0.X.t45 996.134
R7922 two_stage_opamp_dummy_magic_26_0.X.n78 two_stage_opamp_dummy_magic_26_0.X.t27 996.134
R7923 two_stage_opamp_dummy_magic_26_0.X.n79 two_stage_opamp_dummy_magic_26_0.X.t44 996.134
R7924 two_stage_opamp_dummy_magic_26_0.X.n75 two_stage_opamp_dummy_magic_26_0.X.t30 996.134
R7925 two_stage_opamp_dummy_magic_26_0.X.n74 two_stage_opamp_dummy_magic_26_0.X.t47 996.134
R7926 two_stage_opamp_dummy_magic_26_0.X.n73 two_stage_opamp_dummy_magic_26_0.X.t33 996.134
R7927 two_stage_opamp_dummy_magic_26_0.X.n72 two_stage_opamp_dummy_magic_26_0.X.t51 996.134
R7928 two_stage_opamp_dummy_magic_26_0.X.n35 two_stage_opamp_dummy_magic_26_0.X.t31 690.867
R7929 two_stage_opamp_dummy_magic_26_0.X.n34 two_stage_opamp_dummy_magic_26_0.X.t54 690.867
R7930 two_stage_opamp_dummy_magic_26_0.X.n44 two_stage_opamp_dummy_magic_26_0.X.t40 530.201
R7931 two_stage_opamp_dummy_magic_26_0.X.n43 two_stage_opamp_dummy_magic_26_0.X.t36 530.201
R7932 two_stage_opamp_dummy_magic_26_0.X.n41 two_stage_opamp_dummy_magic_26_0.X.t53 514.134
R7933 two_stage_opamp_dummy_magic_26_0.X.n40 two_stage_opamp_dummy_magic_26_0.X.t38 514.134
R7934 two_stage_opamp_dummy_magic_26_0.X.n39 two_stage_opamp_dummy_magic_26_0.X.t52 514.134
R7935 two_stage_opamp_dummy_magic_26_0.X.n38 two_stage_opamp_dummy_magic_26_0.X.t34 514.134
R7936 two_stage_opamp_dummy_magic_26_0.X.n37 two_stage_opamp_dummy_magic_26_0.X.t48 514.134
R7937 two_stage_opamp_dummy_magic_26_0.X.n36 two_stage_opamp_dummy_magic_26_0.X.t35 514.134
R7938 two_stage_opamp_dummy_magic_26_0.X.n35 two_stage_opamp_dummy_magic_26_0.X.t49 514.134
R7939 two_stage_opamp_dummy_magic_26_0.X.n34 two_stage_opamp_dummy_magic_26_0.X.t39 514.134
R7940 two_stage_opamp_dummy_magic_26_0.X.n44 two_stage_opamp_dummy_magic_26_0.X.t26 353.467
R7941 two_stage_opamp_dummy_magic_26_0.X.n45 two_stage_opamp_dummy_magic_26_0.X.t43 353.467
R7942 two_stage_opamp_dummy_magic_26_0.X.n46 two_stage_opamp_dummy_magic_26_0.X.t25 353.467
R7943 two_stage_opamp_dummy_magic_26_0.X.n47 two_stage_opamp_dummy_magic_26_0.X.t42 353.467
R7944 two_stage_opamp_dummy_magic_26_0.X.n48 two_stage_opamp_dummy_magic_26_0.X.t29 353.467
R7945 two_stage_opamp_dummy_magic_26_0.X.n49 two_stage_opamp_dummy_magic_26_0.X.t46 353.467
R7946 two_stage_opamp_dummy_magic_26_0.X.n50 two_stage_opamp_dummy_magic_26_0.X.t32 353.467
R7947 two_stage_opamp_dummy_magic_26_0.X.n43 two_stage_opamp_dummy_magic_26_0.X.t50 353.467
R7948 two_stage_opamp_dummy_magic_26_0.X.n75 two_stage_opamp_dummy_magic_26_0.X.n74 176.733
R7949 two_stage_opamp_dummy_magic_26_0.X.n74 two_stage_opamp_dummy_magic_26_0.X.n73 176.733
R7950 two_stage_opamp_dummy_magic_26_0.X.n73 two_stage_opamp_dummy_magic_26_0.X.n72 176.733
R7951 two_stage_opamp_dummy_magic_26_0.X.n77 two_stage_opamp_dummy_magic_26_0.X.n76 176.733
R7952 two_stage_opamp_dummy_magic_26_0.X.n78 two_stage_opamp_dummy_magic_26_0.X.n77 176.733
R7953 two_stage_opamp_dummy_magic_26_0.X.n79 two_stage_opamp_dummy_magic_26_0.X.n78 176.733
R7954 two_stage_opamp_dummy_magic_26_0.X.n45 two_stage_opamp_dummy_magic_26_0.X.n44 176.733
R7955 two_stage_opamp_dummy_magic_26_0.X.n46 two_stage_opamp_dummy_magic_26_0.X.n45 176.733
R7956 two_stage_opamp_dummy_magic_26_0.X.n47 two_stage_opamp_dummy_magic_26_0.X.n46 176.733
R7957 two_stage_opamp_dummy_magic_26_0.X.n48 two_stage_opamp_dummy_magic_26_0.X.n47 176.733
R7958 two_stage_opamp_dummy_magic_26_0.X.n49 two_stage_opamp_dummy_magic_26_0.X.n48 176.733
R7959 two_stage_opamp_dummy_magic_26_0.X.n50 two_stage_opamp_dummy_magic_26_0.X.n49 176.733
R7960 two_stage_opamp_dummy_magic_26_0.X.n36 two_stage_opamp_dummy_magic_26_0.X.n35 176.733
R7961 two_stage_opamp_dummy_magic_26_0.X.n37 two_stage_opamp_dummy_magic_26_0.X.n36 176.733
R7962 two_stage_opamp_dummy_magic_26_0.X.n38 two_stage_opamp_dummy_magic_26_0.X.n37 176.733
R7963 two_stage_opamp_dummy_magic_26_0.X.n39 two_stage_opamp_dummy_magic_26_0.X.n38 176.733
R7964 two_stage_opamp_dummy_magic_26_0.X.n40 two_stage_opamp_dummy_magic_26_0.X.n39 176.733
R7965 two_stage_opamp_dummy_magic_26_0.X.n41 two_stage_opamp_dummy_magic_26_0.X.n40 176.733
R7966 two_stage_opamp_dummy_magic_26_0.X.n52 two_stage_opamp_dummy_magic_26_0.X.n51 165.472
R7967 two_stage_opamp_dummy_magic_26_0.X.n52 two_stage_opamp_dummy_magic_26_0.X.n42 165.472
R7968 two_stage_opamp_dummy_magic_26_0.X.n82 two_stage_opamp_dummy_magic_26_0.X.n81 152
R7969 two_stage_opamp_dummy_magic_26_0.X.n83 two_stage_opamp_dummy_magic_26_0.X.n82 131.571
R7970 two_stage_opamp_dummy_magic_26_0.X.n82 two_stage_opamp_dummy_magic_26_0.X.n80 124.517
R7971 two_stage_opamp_dummy_magic_26_0.X.n60 two_stage_opamp_dummy_magic_26_0.X.n52 73.687
R7972 two_stage_opamp_dummy_magic_26_0.X.n11 two_stage_opamp_dummy_magic_26_0.X.n10 66.0338
R7973 two_stage_opamp_dummy_magic_26_0.X.n27 two_stage_opamp_dummy_magic_26_0.X.n26 66.0338
R7974 two_stage_opamp_dummy_magic_26_0.X.n24 two_stage_opamp_dummy_magic_26_0.X.n23 66.0338
R7975 two_stage_opamp_dummy_magic_26_0.X.n21 two_stage_opamp_dummy_magic_26_0.X.n20 66.0338
R7976 two_stage_opamp_dummy_magic_26_0.X.n17 two_stage_opamp_dummy_magic_26_0.X.n16 66.0338
R7977 two_stage_opamp_dummy_magic_26_0.X.n14 two_stage_opamp_dummy_magic_26_0.X.n13 66.0338
R7978 two_stage_opamp_dummy_magic_26_0.X.n109 two_stage_opamp_dummy_magic_26_0.X.n107 54.7984
R7979 two_stage_opamp_dummy_magic_26_0.X.n117 two_stage_opamp_dummy_magic_26_0.X.n116 54.4547
R7980 two_stage_opamp_dummy_magic_26_0.X.n115 two_stage_opamp_dummy_magic_26_0.X.n114 54.4547
R7981 two_stage_opamp_dummy_magic_26_0.X.n113 two_stage_opamp_dummy_magic_26_0.X.n112 54.4547
R7982 two_stage_opamp_dummy_magic_26_0.X.n111 two_stage_opamp_dummy_magic_26_0.X.n110 54.4547
R7983 two_stage_opamp_dummy_magic_26_0.X.n109 two_stage_opamp_dummy_magic_26_0.X.n108 54.4547
R7984 two_stage_opamp_dummy_magic_26_0.X.n66 two_stage_opamp_dummy_magic_26_0.X.t2 41.0384
R7985 two_stage_opamp_dummy_magic_26_0.X.n80 two_stage_opamp_dummy_magic_26_0.X.n75 40.1672
R7986 two_stage_opamp_dummy_magic_26_0.X.n80 two_stage_opamp_dummy_magic_26_0.X.n79 40.1672
R7987 two_stage_opamp_dummy_magic_26_0.X.n51 two_stage_opamp_dummy_magic_26_0.X.n43 40.1672
R7988 two_stage_opamp_dummy_magic_26_0.X.n51 two_stage_opamp_dummy_magic_26_0.X.n50 40.1672
R7989 two_stage_opamp_dummy_magic_26_0.X.n42 two_stage_opamp_dummy_magic_26_0.X.n34 40.1672
R7990 two_stage_opamp_dummy_magic_26_0.X.n42 two_stage_opamp_dummy_magic_26_0.X.n41 40.1672
R7991 two_stage_opamp_dummy_magic_26_0.X.n84 two_stage_opamp_dummy_magic_26_0.X.n83 16.3217
R7992 two_stage_opamp_dummy_magic_26_0.X.n116 two_stage_opamp_dummy_magic_26_0.X.t16 16.0005
R7993 two_stage_opamp_dummy_magic_26_0.X.n116 two_stage_opamp_dummy_magic_26_0.X.t4 16.0005
R7994 two_stage_opamp_dummy_magic_26_0.X.n114 two_stage_opamp_dummy_magic_26_0.X.t10 16.0005
R7995 two_stage_opamp_dummy_magic_26_0.X.n114 two_stage_opamp_dummy_magic_26_0.X.t15 16.0005
R7996 two_stage_opamp_dummy_magic_26_0.X.n112 two_stage_opamp_dummy_magic_26_0.X.t11 16.0005
R7997 two_stage_opamp_dummy_magic_26_0.X.n112 two_stage_opamp_dummy_magic_26_0.X.t17 16.0005
R7998 two_stage_opamp_dummy_magic_26_0.X.n110 two_stage_opamp_dummy_magic_26_0.X.t18 16.0005
R7999 two_stage_opamp_dummy_magic_26_0.X.n110 two_stage_opamp_dummy_magic_26_0.X.t13 16.0005
R8000 two_stage_opamp_dummy_magic_26_0.X.n108 two_stage_opamp_dummy_magic_26_0.X.t12 16.0005
R8001 two_stage_opamp_dummy_magic_26_0.X.n108 two_stage_opamp_dummy_magic_26_0.X.t14 16.0005
R8002 two_stage_opamp_dummy_magic_26_0.X.n107 two_stage_opamp_dummy_magic_26_0.X.t3 16.0005
R8003 two_stage_opamp_dummy_magic_26_0.X.n107 two_stage_opamp_dummy_magic_26_0.X.t9 16.0005
R8004 two_stage_opamp_dummy_magic_26_0.X.n81 two_stage_opamp_dummy_magic_26_0.X.n71 12.8005
R8005 two_stage_opamp_dummy_magic_26_0.X.n10 two_stage_opamp_dummy_magic_26_0.X.t23 11.2576
R8006 two_stage_opamp_dummy_magic_26_0.X.n10 two_stage_opamp_dummy_magic_26_0.X.t24 11.2576
R8007 two_stage_opamp_dummy_magic_26_0.X.n26 two_stage_opamp_dummy_magic_26_0.X.t22 11.2576
R8008 two_stage_opamp_dummy_magic_26_0.X.n26 two_stage_opamp_dummy_magic_26_0.X.t7 11.2576
R8009 two_stage_opamp_dummy_magic_26_0.X.n23 two_stage_opamp_dummy_magic_26_0.X.t8 11.2576
R8010 two_stage_opamp_dummy_magic_26_0.X.n23 two_stage_opamp_dummy_magic_26_0.X.t19 11.2576
R8011 two_stage_opamp_dummy_magic_26_0.X.n20 two_stage_opamp_dummy_magic_26_0.X.t5 11.2576
R8012 two_stage_opamp_dummy_magic_26_0.X.n20 two_stage_opamp_dummy_magic_26_0.X.t21 11.2576
R8013 two_stage_opamp_dummy_magic_26_0.X.n16 two_stage_opamp_dummy_magic_26_0.X.t0 11.2576
R8014 two_stage_opamp_dummy_magic_26_0.X.n16 two_stage_opamp_dummy_magic_26_0.X.t20 11.2576
R8015 two_stage_opamp_dummy_magic_26_0.X.n13 two_stage_opamp_dummy_magic_26_0.X.t6 11.2576
R8016 two_stage_opamp_dummy_magic_26_0.X.n13 two_stage_opamp_dummy_magic_26_0.X.t1 11.2576
R8017 two_stage_opamp_dummy_magic_26_0.X.n118 two_stage_opamp_dummy_magic_26_0.X.n117 10.9224
R8018 two_stage_opamp_dummy_magic_26_0.X.n81 two_stage_opamp_dummy_magic_26_0.X.n69 9.36264
R8019 two_stage_opamp_dummy_magic_26_0.X.n71 two_stage_opamp_dummy_magic_26_0.X.n70 9.3005
R8020 two_stage_opamp_dummy_magic_26_0.X.n102 two_stage_opamp_dummy_magic_26_0.X.n3 6.1255
R8021 two_stage_opamp_dummy_magic_26_0.X.n119 two_stage_opamp_dummy_magic_26_0.X.n118 5.84022
R8022 two_stage_opamp_dummy_magic_26_0.X.n102 two_stage_opamp_dummy_magic_26_0.X.n101 5.78175
R8023 two_stage_opamp_dummy_magic_26_0.X.n103 two_stage_opamp_dummy_magic_26_0.X.n2 5.78175
R8024 two_stage_opamp_dummy_magic_26_0.X.n122 two_stage_opamp_dummy_magic_26_0.X.n104 5.78175
R8025 two_stage_opamp_dummy_magic_26_0.X.n106 two_stage_opamp_dummy_magic_26_0.X.n105 5.78175
R8026 two_stage_opamp_dummy_magic_26_0.X.n27 two_stage_opamp_dummy_magic_26_0.X.n25 5.66717
R8027 two_stage_opamp_dummy_magic_26_0.X.n12 two_stage_opamp_dummy_magic_26_0.X.n11 5.66717
R8028 two_stage_opamp_dummy_magic_26_0.X.n15 two_stage_opamp_dummy_magic_26_0.X.n11 5.66717
R8029 two_stage_opamp_dummy_magic_26_0.X.n83 two_stage_opamp_dummy_magic_26_0.X.n71 5.33141
R8030 two_stage_opamp_dummy_magic_26_0.X.n28 two_stage_opamp_dummy_magic_26_0.X.n27 5.29217
R8031 two_stage_opamp_dummy_magic_26_0.X.n24 two_stage_opamp_dummy_magic_26_0.X.n8 5.29217
R8032 two_stage_opamp_dummy_magic_26_0.X.n25 two_stage_opamp_dummy_magic_26_0.X.n24 5.29217
R8033 two_stage_opamp_dummy_magic_26_0.X.n21 two_stage_opamp_dummy_magic_26_0.X.n19 5.29217
R8034 two_stage_opamp_dummy_magic_26_0.X.n22 two_stage_opamp_dummy_magic_26_0.X.n21 5.29217
R8035 two_stage_opamp_dummy_magic_26_0.X.n18 two_stage_opamp_dummy_magic_26_0.X.n17 5.29217
R8036 two_stage_opamp_dummy_magic_26_0.X.n17 two_stage_opamp_dummy_magic_26_0.X.n9 5.29217
R8037 two_stage_opamp_dummy_magic_26_0.X.n15 two_stage_opamp_dummy_magic_26_0.X.n14 5.29217
R8038 two_stage_opamp_dummy_magic_26_0.X.n14 two_stage_opamp_dummy_magic_26_0.X.n12 5.29217
R8039 two_stage_opamp_dummy_magic_26_0.X.n29 two_stage_opamp_dummy_magic_26_0.X.n7 4.5005
R8040 two_stage_opamp_dummy_magic_26_0.X.n55 two_stage_opamp_dummy_magic_26_0.X.n54 4.5005
R8041 two_stage_opamp_dummy_magic_26_0.X.n86 two_stage_opamp_dummy_magic_26_0.X.n31 4.5005
R8042 two_stage_opamp_dummy_magic_26_0.X.n88 two_stage_opamp_dummy_magic_26_0.X.n87 4.5005
R8043 two_stage_opamp_dummy_magic_26_0.X.n87 two_stage_opamp_dummy_magic_26_0.X.n86 4.5005
R8044 two_stage_opamp_dummy_magic_26_0.X.n85 two_stage_opamp_dummy_magic_26_0.X.n84 4.5005
R8045 two_stage_opamp_dummy_magic_26_0.X.n63 two_stage_opamp_dummy_magic_26_0.X.n62 4.5005
R8046 two_stage_opamp_dummy_magic_26_0.X.n94 two_stage_opamp_dummy_magic_26_0.X.n28 2.35465
R8047 two_stage_opamp_dummy_magic_26_0.X.n93 two_stage_opamp_dummy_magic_26_0.X.n92 2.26187
R8048 two_stage_opamp_dummy_magic_26_0.X.n56 two_stage_opamp_dummy_magic_26_0.X.n53 2.26187
R8049 two_stage_opamp_dummy_magic_26_0.X.n57 two_stage_opamp_dummy_magic_26_0.X.n56 2.26187
R8050 two_stage_opamp_dummy_magic_26_0.X.n65 two_stage_opamp_dummy_magic_26_0.X.n64 2.26187
R8051 two_stage_opamp_dummy_magic_26_0.X.n64 two_stage_opamp_dummy_magic_26_0.X.n61 2.26187
R8052 two_stage_opamp_dummy_magic_26_0.X.n58 two_stage_opamp_dummy_magic_26_0.X.n57 2.26187
R8053 two_stage_opamp_dummy_magic_26_0.X.n91 two_stage_opamp_dummy_magic_26_0.X.n6 2.24063
R8054 two_stage_opamp_dummy_magic_26_0.X.n89 two_stage_opamp_dummy_magic_26_0.X.n88 2.24063
R8055 two_stage_opamp_dummy_magic_26_0.X.n33 two_stage_opamp_dummy_magic_26_0.X.n32 2.24063
R8056 two_stage_opamp_dummy_magic_26_0.X.n94 two_stage_opamp_dummy_magic_26_0.X.n93 2.24063
R8057 two_stage_opamp_dummy_magic_26_0.X.n96 two_stage_opamp_dummy_magic_26_0.X.n95 2.24063
R8058 two_stage_opamp_dummy_magic_26_0.X.n59 two_stage_opamp_dummy_magic_26_0.X.n53 2.24063
R8059 two_stage_opamp_dummy_magic_26_0.X.n90 two_stage_opamp_dummy_magic_26_0.X.n30 2.24063
R8060 two_stage_opamp_dummy_magic_26_0.X.n66 two_stage_opamp_dummy_magic_26_0.X.n65 2.24063
R8061 two_stage_opamp_dummy_magic_26_0.X.n68 two_stage_opamp_dummy_magic_26_0.X.n67 2.24063
R8062 two_stage_opamp_dummy_magic_26_0.X.n85 two_stage_opamp_dummy_magic_26_0.X.n69 2.22018
R8063 two_stage_opamp_dummy_magic_26_0.X.n121 two_stage_opamp_dummy_magic_26_0.X.n120 1.5005
R8064 two_stage_opamp_dummy_magic_26_0.X.n122 two_stage_opamp_dummy_magic_26_0.X.n1 1.5005
R8065 two_stage_opamp_dummy_magic_26_0.X.n124 two_stage_opamp_dummy_magic_26_0.X.n123 1.5005
R8066 two_stage_opamp_dummy_magic_26_0.X.n2 two_stage_opamp_dummy_magic_26_0.X.n0 1.5005
R8067 two_stage_opamp_dummy_magic_26_0.X.n99 two_stage_opamp_dummy_magic_26_0.X.n5 1.5005
R8068 two_stage_opamp_dummy_magic_26_0.X.n101 two_stage_opamp_dummy_magic_26_0.X.n100 1.5005
R8069 two_stage_opamp_dummy_magic_26_0.X.n98 two_stage_opamp_dummy_magic_26_0.X.n4 1.5005
R8070 two_stage_opamp_dummy_magic_26_0.X.n97 two_stage_opamp_dummy_magic_26_0.X.n3 1.5005
R8071 two_stage_opamp_dummy_magic_26_0.X.n87 two_stage_opamp_dummy_magic_26_0.X.n60 0.850754
R8072 two_stage_opamp_dummy_magic_26_0.X.n85 two_stage_opamp_dummy_magic_26_0.X.n68 0.682792
R8073 two_stage_opamp_dummy_magic_26_0.X.n91 two_stage_opamp_dummy_magic_26_0.X.n90 0.646333
R8074 two_stage_opamp_dummy_magic_26_0.X.n97 two_stage_opamp_dummy_magic_26_0.X.n96 0.630708
R8075 two_stage_opamp_dummy_magic_26_0.X.n120 two_stage_opamp_dummy_magic_26_0.X.n119 0.564601
R8076 two_stage_opamp_dummy_magic_26_0.X.n86 two_stage_opamp_dummy_magic_26_0.X.n85 0.46925
R8077 two_stage_opamp_dummy_magic_26_0.X.n60 two_stage_opamp_dummy_magic_26_0.X.n59 0.37662
R8078 two_stage_opamp_dummy_magic_26_0.X.n12 two_stage_opamp_dummy_magic_26_0.X.n9 0.3755
R8079 two_stage_opamp_dummy_magic_26_0.X.n22 two_stage_opamp_dummy_magic_26_0.X.n9 0.3755
R8080 two_stage_opamp_dummy_magic_26_0.X.n25 two_stage_opamp_dummy_magic_26_0.X.n22 0.3755
R8081 two_stage_opamp_dummy_magic_26_0.X.n18 two_stage_opamp_dummy_magic_26_0.X.n15 0.3755
R8082 two_stage_opamp_dummy_magic_26_0.X.n19 two_stage_opamp_dummy_magic_26_0.X.n18 0.3755
R8083 two_stage_opamp_dummy_magic_26_0.X.n19 two_stage_opamp_dummy_magic_26_0.X.n8 0.3755
R8084 two_stage_opamp_dummy_magic_26_0.X.n28 two_stage_opamp_dummy_magic_26_0.X.n8 0.3755
R8085 two_stage_opamp_dummy_magic_26_0.X.n111 two_stage_opamp_dummy_magic_26_0.X.n109 0.34425
R8086 two_stage_opamp_dummy_magic_26_0.X.n113 two_stage_opamp_dummy_magic_26_0.X.n111 0.34425
R8087 two_stage_opamp_dummy_magic_26_0.X.n115 two_stage_opamp_dummy_magic_26_0.X.n113 0.34425
R8088 two_stage_opamp_dummy_magic_26_0.X.n117 two_stage_opamp_dummy_magic_26_0.X.n115 0.34425
R8089 two_stage_opamp_dummy_magic_26_0.X.n103 two_stage_opamp_dummy_magic_26_0.X.n102 0.34425
R8090 two_stage_opamp_dummy_magic_26_0.X.n104 two_stage_opamp_dummy_magic_26_0.X.n103 0.34425
R8091 two_stage_opamp_dummy_magic_26_0.X.n106 two_stage_opamp_dummy_magic_26_0.X.n104 0.34425
R8092 two_stage_opamp_dummy_magic_26_0.X.n118 two_stage_opamp_dummy_magic_26_0.X.n106 0.34425
R8093 two_stage_opamp_dummy_magic_26_0.X.n84 two_stage_opamp_dummy_magic_26_0.X.n70 0.1255
R8094 two_stage_opamp_dummy_magic_26_0.X.n70 two_stage_opamp_dummy_magic_26_0.X.n69 0.0626438
R8095 two_stage_opamp_dummy_magic_26_0.X.n4 two_stage_opamp_dummy_magic_26_0.X.n3 0.0577917
R8096 two_stage_opamp_dummy_magic_26_0.X.n101 two_stage_opamp_dummy_magic_26_0.X.n4 0.0577917
R8097 two_stage_opamp_dummy_magic_26_0.X.n101 two_stage_opamp_dummy_magic_26_0.X.n5 0.0577917
R8098 two_stage_opamp_dummy_magic_26_0.X.n5 two_stage_opamp_dummy_magic_26_0.X.n2 0.0577917
R8099 two_stage_opamp_dummy_magic_26_0.X.n123 two_stage_opamp_dummy_magic_26_0.X.n2 0.0577917
R8100 two_stage_opamp_dummy_magic_26_0.X.n123 two_stage_opamp_dummy_magic_26_0.X.n122 0.0577917
R8101 two_stage_opamp_dummy_magic_26_0.X.n122 two_stage_opamp_dummy_magic_26_0.X.n121 0.0577917
R8102 two_stage_opamp_dummy_magic_26_0.X.n121 two_stage_opamp_dummy_magic_26_0.X.n105 0.0577917
R8103 two_stage_opamp_dummy_magic_26_0.X.n98 two_stage_opamp_dummy_magic_26_0.X.n97 0.0577917
R8104 two_stage_opamp_dummy_magic_26_0.X.n100 two_stage_opamp_dummy_magic_26_0.X.n98 0.0577917
R8105 two_stage_opamp_dummy_magic_26_0.X.n100 two_stage_opamp_dummy_magic_26_0.X.n99 0.0577917
R8106 two_stage_opamp_dummy_magic_26_0.X.n99 two_stage_opamp_dummy_magic_26_0.X.n0 0.0577917
R8107 two_stage_opamp_dummy_magic_26_0.X.n124 two_stage_opamp_dummy_magic_26_0.X.n1 0.0577917
R8108 two_stage_opamp_dummy_magic_26_0.X.n120 two_stage_opamp_dummy_magic_26_0.X.n1 0.0577917
R8109 two_stage_opamp_dummy_magic_26_0.X.n119 two_stage_opamp_dummy_magic_26_0.X.n105 0.054517
R8110 two_stage_opamp_dummy_magic_26_0.X.n88 two_stage_opamp_dummy_magic_26_0.X.n32 0.0421667
R8111 two_stage_opamp_dummy_magic_26_0.X two_stage_opamp_dummy_magic_26_0.X.n124 0.0369583
R8112 two_stage_opamp_dummy_magic_26_0.X.n96 two_stage_opamp_dummy_magic_26_0.X.n6 0.0217373
R8113 two_stage_opamp_dummy_magic_26_0.X.n92 two_stage_opamp_dummy_magic_26_0.X.n7 0.0217373
R8114 two_stage_opamp_dummy_magic_26_0.X.n90 two_stage_opamp_dummy_magic_26_0.X.n89 0.0217373
R8115 two_stage_opamp_dummy_magic_26_0.X.n87 two_stage_opamp_dummy_magic_26_0.X.n33 0.0217373
R8116 two_stage_opamp_dummy_magic_26_0.X.n56 two_stage_opamp_dummy_magic_26_0.X.n54 0.0217373
R8117 two_stage_opamp_dummy_magic_26_0.X.n29 two_stage_opamp_dummy_magic_26_0.X.n6 0.0217373
R8118 two_stage_opamp_dummy_magic_26_0.X.n92 two_stage_opamp_dummy_magic_26_0.X.n91 0.0217373
R8119 two_stage_opamp_dummy_magic_26_0.X.n57 two_stage_opamp_dummy_magic_26_0.X.n55 0.0217373
R8120 two_stage_opamp_dummy_magic_26_0.X.n68 two_stage_opamp_dummy_magic_26_0.X.n61 0.0217373
R8121 two_stage_opamp_dummy_magic_26_0.X.n89 two_stage_opamp_dummy_magic_26_0.X.n31 0.0217373
R8122 two_stage_opamp_dummy_magic_26_0.X.n33 two_stage_opamp_dummy_magic_26_0.X.n31 0.0217373
R8123 two_stage_opamp_dummy_magic_26_0.X.n64 two_stage_opamp_dummy_magic_26_0.X.n62 0.0217373
R8124 two_stage_opamp_dummy_magic_26_0.X.n63 two_stage_opamp_dummy_magic_26_0.X.n61 0.0217373
R8125 two_stage_opamp_dummy_magic_26_0.X.n55 two_stage_opamp_dummy_magic_26_0.X.n53 0.0217373
R8126 two_stage_opamp_dummy_magic_26_0.X.n93 two_stage_opamp_dummy_magic_26_0.X.n29 0.0217373
R8127 two_stage_opamp_dummy_magic_26_0.X.n95 two_stage_opamp_dummy_magic_26_0.X.n7 0.0217373
R8128 two_stage_opamp_dummy_magic_26_0.X.n58 two_stage_opamp_dummy_magic_26_0.X.n54 0.0217373
R8129 two_stage_opamp_dummy_magic_26_0.X.n95 two_stage_opamp_dummy_magic_26_0.X.n94 0.0217373
R8130 two_stage_opamp_dummy_magic_26_0.X.n59 two_stage_opamp_dummy_magic_26_0.X.n58 0.0217373
R8131 two_stage_opamp_dummy_magic_26_0.X.n65 two_stage_opamp_dummy_magic_26_0.X.n63 0.0217373
R8132 two_stage_opamp_dummy_magic_26_0.X.n86 two_stage_opamp_dummy_magic_26_0.X.n30 0.0217373
R8133 two_stage_opamp_dummy_magic_26_0.X.n32 two_stage_opamp_dummy_magic_26_0.X.n30 0.0217373
R8134 two_stage_opamp_dummy_magic_26_0.X.n67 two_stage_opamp_dummy_magic_26_0.X.n62 0.0217373
R8135 two_stage_opamp_dummy_magic_26_0.X.n67 two_stage_opamp_dummy_magic_26_0.X.n66 0.0217373
R8136 two_stage_opamp_dummy_magic_26_0.X two_stage_opamp_dummy_magic_26_0.X.n0 0.0213333
R8137 two_stage_opamp_dummy_magic_26_0.VD1.n21 two_stage_opamp_dummy_magic_26_0.VD1.n12 49.7255
R8138 two_stage_opamp_dummy_magic_26_0.VD1.n1 two_stage_opamp_dummy_magic_26_0.VD1.n0 49.7255
R8139 two_stage_opamp_dummy_magic_26_0.VD1.n25 two_stage_opamp_dummy_magic_26_0.VD1.n24 49.7255
R8140 two_stage_opamp_dummy_magic_26_0.VD1.n11 two_stage_opamp_dummy_magic_26_0.VD1.n10 49.7255
R8141 two_stage_opamp_dummy_magic_26_0.VD1.n27 two_stage_opamp_dummy_magic_26_0.VD1.n9 49.7255
R8142 two_stage_opamp_dummy_magic_26_0.VD1.n15 two_stage_opamp_dummy_magic_26_0.VD1.n14 49.3505
R8143 two_stage_opamp_dummy_magic_26_0.VD1.n18 two_stage_opamp_dummy_magic_26_0.VD1.n17 49.3505
R8144 two_stage_opamp_dummy_magic_26_0.VD1.n5 two_stage_opamp_dummy_magic_26_0.VD1.n4 49.3505
R8145 two_stage_opamp_dummy_magic_26_0.VD1.n35 two_stage_opamp_dummy_magic_26_0.VD1.n34 49.3505
R8146 two_stage_opamp_dummy_magic_26_0.VD1.n31 two_stage_opamp_dummy_magic_26_0.VD1.n30 49.3505
R8147 two_stage_opamp_dummy_magic_26_0.VD1.n8 two_stage_opamp_dummy_magic_26_0.VD1.n7 49.3505
R8148 two_stage_opamp_dummy_magic_26_0.VD1.n12 two_stage_opamp_dummy_magic_26_0.VD1.t16 16.0005
R8149 two_stage_opamp_dummy_magic_26_0.VD1.n12 two_stage_opamp_dummy_magic_26_0.VD1.t10 16.0005
R8150 two_stage_opamp_dummy_magic_26_0.VD1.n0 two_stage_opamp_dummy_magic_26_0.VD1.t14 16.0005
R8151 two_stage_opamp_dummy_magic_26_0.VD1.n0 two_stage_opamp_dummy_magic_26_0.VD1.t11 16.0005
R8152 two_stage_opamp_dummy_magic_26_0.VD1.n24 two_stage_opamp_dummy_magic_26_0.VD1.t15 16.0005
R8153 two_stage_opamp_dummy_magic_26_0.VD1.n24 two_stage_opamp_dummy_magic_26_0.VD1.t9 16.0005
R8154 two_stage_opamp_dummy_magic_26_0.VD1.n10 two_stage_opamp_dummy_magic_26_0.VD1.t17 16.0005
R8155 two_stage_opamp_dummy_magic_26_0.VD1.n10 two_stage_opamp_dummy_magic_26_0.VD1.t12 16.0005
R8156 two_stage_opamp_dummy_magic_26_0.VD1.n14 two_stage_opamp_dummy_magic_26_0.VD1.t5 16.0005
R8157 two_stage_opamp_dummy_magic_26_0.VD1.n14 two_stage_opamp_dummy_magic_26_0.VD1.t20 16.0005
R8158 two_stage_opamp_dummy_magic_26_0.VD1.n17 two_stage_opamp_dummy_magic_26_0.VD1.t3 16.0005
R8159 two_stage_opamp_dummy_magic_26_0.VD1.n17 two_stage_opamp_dummy_magic_26_0.VD1.t7 16.0005
R8160 two_stage_opamp_dummy_magic_26_0.VD1.n4 two_stage_opamp_dummy_magic_26_0.VD1.t0 16.0005
R8161 two_stage_opamp_dummy_magic_26_0.VD1.n4 two_stage_opamp_dummy_magic_26_0.VD1.t8 16.0005
R8162 two_stage_opamp_dummy_magic_26_0.VD1.n34 two_stage_opamp_dummy_magic_26_0.VD1.t19 16.0005
R8163 two_stage_opamp_dummy_magic_26_0.VD1.n34 two_stage_opamp_dummy_magic_26_0.VD1.t2 16.0005
R8164 two_stage_opamp_dummy_magic_26_0.VD1.n30 two_stage_opamp_dummy_magic_26_0.VD1.t21 16.0005
R8165 two_stage_opamp_dummy_magic_26_0.VD1.n30 two_stage_opamp_dummy_magic_26_0.VD1.t1 16.0005
R8166 two_stage_opamp_dummy_magic_26_0.VD1.n7 two_stage_opamp_dummy_magic_26_0.VD1.t4 16.0005
R8167 two_stage_opamp_dummy_magic_26_0.VD1.n7 two_stage_opamp_dummy_magic_26_0.VD1.t6 16.0005
R8168 two_stage_opamp_dummy_magic_26_0.VD1.n9 two_stage_opamp_dummy_magic_26_0.VD1.t13 16.0005
R8169 two_stage_opamp_dummy_magic_26_0.VD1.n9 two_stage_opamp_dummy_magic_26_0.VD1.t18 16.0005
R8170 two_stage_opamp_dummy_magic_26_0.VD1.n21 two_stage_opamp_dummy_magic_26_0.VD1.n20 7.33383
R8171 two_stage_opamp_dummy_magic_26_0.VD1.n25 two_stage_opamp_dummy_magic_26_0.VD1.n3 7.33383
R8172 two_stage_opamp_dummy_magic_26_0.VD1.n13 two_stage_opamp_dummy_magic_26_0.VD1.n11 7.33383
R8173 two_stage_opamp_dummy_magic_26_0.VD1.n28 two_stage_opamp_dummy_magic_26_0.VD1.n27 7.33383
R8174 two_stage_opamp_dummy_magic_26_0.VD1.n32 two_stage_opamp_dummy_magic_26_0.VD1.n8 5.438
R8175 two_stage_opamp_dummy_magic_26_0.VD1.n16 two_stage_opamp_dummy_magic_26_0.VD1.n15 5.438
R8176 two_stage_opamp_dummy_magic_26_0.VD1.n28 two_stage_opamp_dummy_magic_26_0.VD1.n8 5.31821
R8177 two_stage_opamp_dummy_magic_26_0.VD1.n15 two_stage_opamp_dummy_magic_26_0.VD1.n13 5.31821
R8178 two_stage_opamp_dummy_magic_26_0.VD1.n19 two_stage_opamp_dummy_magic_26_0.VD1.n18 5.08383
R8179 two_stage_opamp_dummy_magic_26_0.VD1.n5 two_stage_opamp_dummy_magic_26_0.VD1.n2 5.08383
R8180 two_stage_opamp_dummy_magic_26_0.VD1.n36 two_stage_opamp_dummy_magic_26_0.VD1.n35 5.08383
R8181 two_stage_opamp_dummy_magic_26_0.VD1.n31 two_stage_opamp_dummy_magic_26_0.VD1.n29 5.08383
R8182 two_stage_opamp_dummy_magic_26_0.VD1.n27 two_stage_opamp_dummy_magic_26_0.VD1.n26 5.063
R8183 two_stage_opamp_dummy_magic_26_0.VD1.n22 two_stage_opamp_dummy_magic_26_0.VD1.n11 5.063
R8184 two_stage_opamp_dummy_magic_26_0.VD1.n18 two_stage_opamp_dummy_magic_26_0.VD1.n16 4.8755
R8185 two_stage_opamp_dummy_magic_26_0.VD1.n6 two_stage_opamp_dummy_magic_26_0.VD1.n5 4.8755
R8186 two_stage_opamp_dummy_magic_26_0.VD1.n35 two_stage_opamp_dummy_magic_26_0.VD1.n33 4.8755
R8187 two_stage_opamp_dummy_magic_26_0.VD1.n32 two_stage_opamp_dummy_magic_26_0.VD1.n31 4.8755
R8188 two_stage_opamp_dummy_magic_26_0.VD1 two_stage_opamp_dummy_magic_26_0.VD1.n37 4.60467
R8189 two_stage_opamp_dummy_magic_26_0.VD1.n26 two_stage_opamp_dummy_magic_26_0.VD1.n25 4.5005
R8190 two_stage_opamp_dummy_magic_26_0.VD1.n23 two_stage_opamp_dummy_magic_26_0.VD1.n1 4.5005
R8191 two_stage_opamp_dummy_magic_26_0.VD1.n22 two_stage_opamp_dummy_magic_26_0.VD1.n21 4.5005
R8192 two_stage_opamp_dummy_magic_26_0.VD1 two_stage_opamp_dummy_magic_26_0.VD1.n1 2.72967
R8193 two_stage_opamp_dummy_magic_26_0.VD1.n26 two_stage_opamp_dummy_magic_26_0.VD1.n23 0.563
R8194 two_stage_opamp_dummy_magic_26_0.VD1.n23 two_stage_opamp_dummy_magic_26_0.VD1.n22 0.563
R8195 two_stage_opamp_dummy_magic_26_0.VD1.n33 two_stage_opamp_dummy_magic_26_0.VD1.n32 0.563
R8196 two_stage_opamp_dummy_magic_26_0.VD1.n33 two_stage_opamp_dummy_magic_26_0.VD1.n6 0.563
R8197 two_stage_opamp_dummy_magic_26_0.VD1.n16 two_stage_opamp_dummy_magic_26_0.VD1.n6 0.563
R8198 two_stage_opamp_dummy_magic_26_0.VD1.n19 two_stage_opamp_dummy_magic_26_0.VD1.n13 0.234875
R8199 two_stage_opamp_dummy_magic_26_0.VD1.n20 two_stage_opamp_dummy_magic_26_0.VD1.n19 0.234875
R8200 two_stage_opamp_dummy_magic_26_0.VD1.n20 two_stage_opamp_dummy_magic_26_0.VD1.n2 0.234875
R8201 two_stage_opamp_dummy_magic_26_0.VD1.n37 two_stage_opamp_dummy_magic_26_0.VD1.n2 0.234875
R8202 two_stage_opamp_dummy_magic_26_0.VD1.n37 two_stage_opamp_dummy_magic_26_0.VD1.n36 0.234875
R8203 two_stage_opamp_dummy_magic_26_0.VD1.n36 two_stage_opamp_dummy_magic_26_0.VD1.n3 0.234875
R8204 two_stage_opamp_dummy_magic_26_0.VD1.n29 two_stage_opamp_dummy_magic_26_0.VD1.n3 0.234875
R8205 two_stage_opamp_dummy_magic_26_0.VD1.n29 two_stage_opamp_dummy_magic_26_0.VD1.n28 0.234875
R8206 GNDA.n3095 GNDA.n3094 396244
R8207 GNDA.n4633 GNDA.n430 254322
R8208 GNDA.n1743 GNDA.n642 203887
R8209 GNDA.n644 GNDA.n429 184643
R8210 GNDA.n4634 GNDA.n428 180896
R8211 GNDA.n4632 GNDA.t289 138700
R8212 GNDA.n1746 GNDA.n1743 132035
R8213 GNDA.n3094 GNDA.n3093 105027
R8214 GNDA.n4632 GNDA.n4631 100684
R8215 GNDA.n3094 GNDA.n3089 71214.8
R8216 GNDA.n3095 GNDA.t288 55812.1
R8217 GNDA.n3090 GNDA.n429 29432.8
R8218 GNDA.n3095 GNDA.n645 29017.7
R8219 GNDA.n1743 GNDA.t278 28013.5
R8220 GNDA.n4634 GNDA.n429 24514.3
R8221 GNDA.n3097 GNDA.n642 23898.2
R8222 GNDA.n645 GNDA.n640 21706.7
R8223 GNDA.n4632 GNDA.t149 17920.8
R8224 GNDA.n4648 GNDA.n4647 17109.1
R8225 GNDA.n3128 GNDA.n640 16116.7
R8226 GNDA.n3091 GNDA.n3090 13613.1
R8227 GNDA.n3096 GNDA.n640 13566.7
R8228 GNDA.n3092 GNDA.n3091 13460.8
R8229 GNDA.n3098 GNDA.n3097 13200
R8230 GNDA.n3129 GNDA.n640 13111.6
R8231 GNDA.n3088 GNDA.n428 11693.7
R8232 GNDA.n4631 GNDA.n430 10098.5
R8233 GNDA.n3097 GNDA.n3096 10046.7
R8234 GNDA.n3089 GNDA.n3088 9511.11
R8235 GNDA.n3090 GNDA.n428 8875.99
R8236 GNDA.n3152 GNDA.n625 7301.54
R8237 GNDA.n3037 GNDA.n3035 7286.54
R8238 GNDA.n4630 GNDA.n431 6490.78
R8239 GNDA.t12 GNDA.n4633 6488.11
R8240 GNDA.t3 GNDA.t33 6013.33
R8241 GNDA.n4631 GNDA.n4630 5937.42
R8242 GNDA.n3093 GNDA.n643 4738.46
R8243 GNDA.t67 GNDA.t3 4571.11
R8244 GNDA.n3095 GNDA.n643 4525.2
R8245 GNDA.n3096 GNDA.n3095 4525.2
R8246 GNDA.n3088 GNDA.t45 4106.67
R8247 GNDA.n3092 GNDA.n3089 4106.67
R8248 GNDA.n644 GNDA.n430 3428.05
R8249 GNDA.t67 GNDA.t1 2517.78
R8250 GNDA.n3129 GNDA.t112 2212.22
R8251 GNDA.n3095 GNDA.n429 2005.06
R8252 GNDA.n697 GNDA.n696 1684.55
R8253 GNDA.n4630 GNDA.n4629 1560.83
R8254 GNDA.n645 GNDA.n644 1336.71
R8255 GNDA.t112 GNDA.t254 1271.11
R8256 GNDA.t33 GNDA.n3129 1161.11
R8257 GNDA.n3093 GNDA.n3092 1031.25
R8258 GNDA.n642 GNDA.n625 857.37
R8259 GNDA.n3091 GNDA.n643 854.477
R8260 GNDA.n1744 GNDA.t63 749.742
R8261 GNDA.n4624 GNDA.t125 749.742
R8262 GNDA.n4627 GNDA.t88 749.742
R8263 GNDA.n3150 GNDA.t76 747.734
R8264 GNDA.t45 GNDA.n102 741.376
R8265 GNDA.n3023 GNDA.n3022 686.717
R8266 GNDA.n2408 GNDA.n2407 686.717
R8267 GNDA.n2400 GNDA.n2276 686.717
R8268 GNDA.n3014 GNDA.n708 686.717
R8269 GNDA.n2762 GNDA.t152 671.187
R8270 GNDA.n2386 GNDA.n2385 669.307
R8271 GNDA.n2291 GNDA.n2290 669.307
R8272 GNDA.n1274 GNDA.t136 659.367
R8273 GNDA.n1272 GNDA.t57 659.367
R8274 GNDA.n641 GNDA.t96 659.367
R8275 GNDA.n3125 GNDA.t121 659.367
R8276 GNDA.n4689 GNDA.n357 654.447
R8277 GNDA.n4633 GNDA.n4632 630.303
R8278 GNDA.n2241 GNDA.n2240 585.003
R8279 GNDA.n2513 GNDA.n2512 585.001
R8280 GNDA.n2501 GNDA.n2500 585.001
R8281 GNDA.n2320 GNDA.n2319 585.001
R8282 GNDA.n3062 GNDA.n3061 585.001
R8283 GNDA.n808 GNDA.n807 585.001
R8284 GNDA.n2976 GNDA.n2975 585.001
R8285 GNDA.n3049 GNDA.n3048 585.001
R8286 GNDA.n4704 GNDA.n4703 585
R8287 GNDA.n4705 GNDA.n4704 585
R8288 GNDA.n299 GNDA.n298 585
R8289 GNDA.n4706 GNDA.n299 585
R8290 GNDA.n4709 GNDA.n4708 585
R8291 GNDA.n4708 GNDA.n4707 585
R8292 GNDA.n4710 GNDA.n297 585
R8293 GNDA.n297 GNDA.n296 585
R8294 GNDA.n4712 GNDA.n4711 585
R8295 GNDA.n4713 GNDA.n4712 585
R8296 GNDA.n295 GNDA.n294 585
R8297 GNDA.n4714 GNDA.n295 585
R8298 GNDA.n4717 GNDA.n4716 585
R8299 GNDA.n4716 GNDA.n4715 585
R8300 GNDA.n4718 GNDA.n293 585
R8301 GNDA.n293 GNDA.n292 585
R8302 GNDA.n4720 GNDA.n4719 585
R8303 GNDA.n4721 GNDA.n4720 585
R8304 GNDA.n291 GNDA.n290 585
R8305 GNDA.n4722 GNDA.n291 585
R8306 GNDA.n4725 GNDA.n4724 585
R8307 GNDA.n4724 GNDA.n4723 585
R8308 GNDA.n4726 GNDA.n289 585
R8309 GNDA.n289 GNDA.n99 585
R8310 GNDA.n4688 GNDA.n4687 585
R8311 GNDA.n4686 GNDA.n355 585
R8312 GNDA.t45 GNDA.n355 585
R8313 GNDA.n5085 GNDA.n5084 585
R8314 GNDA.n131 GNDA.n129 585
R8315 GNDA.n242 GNDA.n241 585
R8316 GNDA.n244 GNDA.n243 585
R8317 GNDA.n246 GNDA.n245 585
R8318 GNDA.n248 GNDA.n247 585
R8319 GNDA.n250 GNDA.n249 585
R8320 GNDA.n252 GNDA.n251 585
R8321 GNDA.n254 GNDA.n253 585
R8322 GNDA.n256 GNDA.n255 585
R8323 GNDA.n258 GNDA.n257 585
R8324 GNDA.n260 GNDA.n259 585
R8325 GNDA.n2611 GNDA.n2610 585
R8326 GNDA.n2608 GNDA.n2607 585
R8327 GNDA.n2606 GNDA.n2605 585
R8328 GNDA.n2604 GNDA.n2603 585
R8329 GNDA.n2602 GNDA.n2601 585
R8330 GNDA.n2600 GNDA.n2599 585
R8331 GNDA.n2598 GNDA.n2597 585
R8332 GNDA.n2596 GNDA.n2595 585
R8333 GNDA.n2594 GNDA.n2593 585
R8334 GNDA.n2592 GNDA.n2591 585
R8335 GNDA.n2590 GNDA.n2589 585
R8336 GNDA.n135 GNDA.n132 585
R8337 GNDA.n2765 GNDA.n2764 585
R8338 GNDA.n2767 GNDA.n2766 585
R8339 GNDA.n2769 GNDA.n2768 585
R8340 GNDA.n2771 GNDA.n2770 585
R8341 GNDA.n2773 GNDA.n2772 585
R8342 GNDA.n2775 GNDA.n2774 585
R8343 GNDA.n2777 GNDA.n2776 585
R8344 GNDA.n2779 GNDA.n2778 585
R8345 GNDA.n2781 GNDA.n2780 585
R8346 GNDA.n2783 GNDA.n2782 585
R8347 GNDA.n2785 GNDA.n2784 585
R8348 GNDA.n2787 GNDA.n2786 585
R8349 GNDA.n5265 GNDA.n5264 585
R8350 GNDA.n5262 GNDA.n54 585
R8351 GNDA.n59 GNDA.n58 585
R8352 GNDA.n5257 GNDA.n5256 585
R8353 GNDA.n5255 GNDA.n5254 585
R8354 GNDA.n5181 GNDA.n63 585
R8355 GNDA.n5183 GNDA.n5182 585
R8356 GNDA.n5188 GNDA.n5187 585
R8357 GNDA.n5186 GNDA.n5179 585
R8358 GNDA.n5194 GNDA.n5193 585
R8359 GNDA.n5196 GNDA.n5195 585
R8360 GNDA.n5177 GNDA.n5176 585
R8361 GNDA.n4842 GNDA.n4841 585
R8362 GNDA.n4839 GNDA.n4838 585
R8363 GNDA.n4837 GNDA.n4836 585
R8364 GNDA.n4753 GNDA.n4729 585
R8365 GNDA.n4755 GNDA.n4754 585
R8366 GNDA.n4759 GNDA.n4758 585
R8367 GNDA.n4761 GNDA.n4760 585
R8368 GNDA.n4768 GNDA.n4767 585
R8369 GNDA.n4766 GNDA.n4751 585
R8370 GNDA.n4774 GNDA.n4773 585
R8371 GNDA.n4776 GNDA.n4775 585
R8372 GNDA.n4749 GNDA.n4748 585
R8373 GNDA.n328 GNDA.n325 585
R8374 GNDA.n329 GNDA.n323 585
R8375 GNDA.n330 GNDA.n322 585
R8376 GNDA.n320 GNDA.n318 585
R8377 GNDA.n336 GNDA.n317 585
R8378 GNDA.n337 GNDA.n315 585
R8379 GNDA.n338 GNDA.n314 585
R8380 GNDA.n312 GNDA.n310 585
R8381 GNDA.n344 GNDA.n309 585
R8382 GNDA.n345 GNDA.n307 585
R8383 GNDA.n346 GNDA.n306 585
R8384 GNDA.n302 GNDA.n301 585
R8385 GNDA.n133 GNDA.n85 585
R8386 GNDA.n5174 GNDA.n85 585
R8387 GNDA.n349 GNDA.n302 585
R8388 GNDA.n347 GNDA.n346 585
R8389 GNDA.n345 GNDA.n304 585
R8390 GNDA.n344 GNDA.n343 585
R8391 GNDA.n341 GNDA.n310 585
R8392 GNDA.n339 GNDA.n338 585
R8393 GNDA.n337 GNDA.n311 585
R8394 GNDA.n336 GNDA.n335 585
R8395 GNDA.n333 GNDA.n318 585
R8396 GNDA.n331 GNDA.n330 585
R8397 GNDA.n329 GNDA.n319 585
R8398 GNDA.n328 GNDA.n327 585
R8399 GNDA.n133 GNDA.n55 585
R8400 GNDA.n5174 GNDA.n55 585
R8401 GNDA.n5060 GNDA.n159 585
R8402 GNDA.n5061 GNDA.n150 585
R8403 GNDA.n5064 GNDA.n149 585
R8404 GNDA.n5065 GNDA.n148 585
R8405 GNDA.n5068 GNDA.n147 585
R8406 GNDA.n5069 GNDA.n146 585
R8407 GNDA.n5072 GNDA.n145 585
R8408 GNDA.n5074 GNDA.n144 585
R8409 GNDA.n5075 GNDA.n143 585
R8410 GNDA.n5076 GNDA.n142 585
R8411 GNDA.n151 GNDA.n134 585
R8412 GNDA.n5082 GNDA.n130 585
R8413 GNDA.n5082 GNDA.n5081 585
R8414 GNDA.n136 GNDA.n134 585
R8415 GNDA.n5077 GNDA.n5076 585
R8416 GNDA.n5075 GNDA.n141 585
R8417 GNDA.n5074 GNDA.n5073 585
R8418 GNDA.n5072 GNDA.n5071 585
R8419 GNDA.n5070 GNDA.n5069 585
R8420 GNDA.n5068 GNDA.n5067 585
R8421 GNDA.n5066 GNDA.n5065 585
R8422 GNDA.n5064 GNDA.n5063 585
R8423 GNDA.n5062 GNDA.n5061 585
R8424 GNDA.n5060 GNDA.n5059 585
R8425 GNDA.n2972 GNDA.n812 585
R8426 GNDA.n2970 GNDA.n2969 585
R8427 GNDA.n814 GNDA.n813 585
R8428 GNDA.n820 GNDA.n816 585
R8429 GNDA.n2962 GNDA.n2961 585
R8430 GNDA.n2959 GNDA.n818 585
R8431 GNDA.n2958 GNDA.n821 585
R8432 GNDA.n2956 GNDA.n2955 585
R8433 GNDA.n823 GNDA.n822 585
R8434 GNDA.n2950 GNDA.n2949 585
R8435 GNDA.n2947 GNDA.n827 585
R8436 GNDA.n2945 GNDA.n2944 585
R8437 GNDA.n2944 GNDA.n2943 585
R8438 GNDA.n827 GNDA.n826 585
R8439 GNDA.n2951 GNDA.n2950 585
R8440 GNDA.n2951 GNDA.n646 585
R8441 GNDA.n2952 GNDA.n823 585
R8442 GNDA.n2955 GNDA.n2954 585
R8443 GNDA.n825 GNDA.n821 585
R8444 GNDA.n818 GNDA.n817 585
R8445 GNDA.n2963 GNDA.n2962 585
R8446 GNDA.n2965 GNDA.n816 585
R8447 GNDA.n2966 GNDA.n814 585
R8448 GNDA.n2969 GNDA.n2968 585
R8449 GNDA.n815 GNDA.n812 585
R8450 GNDA.n815 GNDA.n646 585
R8451 GNDA.n2563 GNDA.n828 585
R8452 GNDA.n2562 GNDA.n2561 585
R8453 GNDA.n2559 GNDA.n829 585
R8454 GNDA.n2557 GNDA.n2556 585
R8455 GNDA.n2555 GNDA.n830 585
R8456 GNDA.n2554 GNDA.n2553 585
R8457 GNDA.n2551 GNDA.n831 585
R8458 GNDA.n2549 GNDA.n2548 585
R8459 GNDA.n2547 GNDA.n832 585
R8460 GNDA.n2546 GNDA.n2545 585
R8461 GNDA.n2543 GNDA.n833 585
R8462 GNDA.n2541 GNDA.n2540 585
R8463 GNDA.n2922 GNDA.n2921 585
R8464 GNDA.n2923 GNDA.n2572 585
R8465 GNDA.n2925 GNDA.n2924 585
R8466 GNDA.n2927 GNDA.n2570 585
R8467 GNDA.n2929 GNDA.n2928 585
R8468 GNDA.n2930 GNDA.n2569 585
R8469 GNDA.n2932 GNDA.n2931 585
R8470 GNDA.n2934 GNDA.n2567 585
R8471 GNDA.n2936 GNDA.n2935 585
R8472 GNDA.n2937 GNDA.n2566 585
R8473 GNDA.n2939 GNDA.n2938 585
R8474 GNDA.n2941 GNDA.n2565 585
R8475 GNDA.n2894 GNDA.n2893 585
R8476 GNDA.n2895 GNDA.n2867 585
R8477 GNDA.n2897 GNDA.n2896 585
R8478 GNDA.n2899 GNDA.n2865 585
R8479 GNDA.n2901 GNDA.n2900 585
R8480 GNDA.n2902 GNDA.n2864 585
R8481 GNDA.n2904 GNDA.n2903 585
R8482 GNDA.n2906 GNDA.n2862 585
R8483 GNDA.n2908 GNDA.n2907 585
R8484 GNDA.n2909 GNDA.n2861 585
R8485 GNDA.n2911 GNDA.n2910 585
R8486 GNDA.n2913 GNDA.n2860 585
R8487 GNDA.n4896 GNDA.n162 585
R8488 GNDA.n4896 GNDA.n161 585
R8489 GNDA.n4986 GNDA.n4985 585
R8490 GNDA.n4983 GNDA.n226 585
R8491 GNDA.n4873 GNDA.n4872 585
R8492 GNDA.n4978 GNDA.n4977 585
R8493 GNDA.n4976 GNDA.n4975 585
R8494 GNDA.n4902 GNDA.n4877 585
R8495 GNDA.n4904 GNDA.n4903 585
R8496 GNDA.n4909 GNDA.n4908 585
R8497 GNDA.n4907 GNDA.n4900 585
R8498 GNDA.n4915 GNDA.n4914 585
R8499 GNDA.n4917 GNDA.n4916 585
R8500 GNDA.n4898 GNDA.n4897 585
R8501 GNDA.n5058 GNDA.n162 585
R8502 GNDA.n5058 GNDA.n161 585
R8503 GNDA.n5057 GNDA.n5056 585
R8504 GNDA.n5054 GNDA.n5053 585
R8505 GNDA.n5052 GNDA.n5051 585
R8506 GNDA.n199 GNDA.n167 585
R8507 GNDA.n219 GNDA.n218 585
R8508 GNDA.n215 GNDA.n198 585
R8509 GNDA.n202 GNDA.n201 585
R8510 GNDA.n210 GNDA.n209 585
R8511 GNDA.n208 GNDA.n207 585
R8512 GNDA.n188 GNDA.n187 585
R8513 GNDA.n4991 GNDA.n4990 585
R8514 GNDA.n2573 GNDA.n189 585
R8515 GNDA.n2700 GNDA.n2576 585
R8516 GNDA.n2724 GNDA.n2702 585
R8517 GNDA.n2726 GNDA.n2725 585
R8518 GNDA.n2722 GNDA.n2721 585
R8519 GNDA.n2720 GNDA.n2719 585
R8520 GNDA.n2715 GNDA.n2714 585
R8521 GNDA.n2713 GNDA.n2712 585
R8522 GNDA.n2708 GNDA.n2707 585
R8523 GNDA.n2706 GNDA.n2627 585
R8524 GNDA.n2734 GNDA.n2733 585
R8525 GNDA.n2736 GNDA.n2735 585
R8526 GNDA.n2739 GNDA.n2738 585
R8527 GNDA.n3034 GNDA.n3033 585
R8528 GNDA.n3035 GNDA.n3034 585
R8529 GNDA.n3031 GNDA.n698 585
R8530 GNDA.n698 GNDA.n697 585
R8531 GNDA.n3038 GNDA.n694 585
R8532 GNDA.n3041 GNDA.n3040 585
R8533 GNDA.n3040 GNDA.n3039 585
R8534 GNDA.n693 GNDA.n692 585
R8535 GNDA.n695 GNDA.n693 585
R8536 GNDA.n2877 GNDA.n2876 585
R8537 GNDA.n2879 GNDA.n2876 585
R8538 GNDA.n2881 GNDA.n2878 585
R8539 GNDA.n2881 GNDA.n2880 585
R8540 GNDA.n2882 GNDA.n2875 585
R8541 GNDA.n2882 GNDA.n710 585
R8542 GNDA.n2884 GNDA.n2883 585
R8543 GNDA.n2883 GNDA.n709 585
R8544 GNDA.n2885 GNDA.n2873 585
R8545 GNDA.n2873 GNDA.n2872 585
R8546 GNDA.n2887 GNDA.n2886 585
R8547 GNDA.n2888 GNDA.n2887 585
R8548 GNDA.n2874 GNDA.n2870 585
R8549 GNDA.n2889 GNDA.n2870 585
R8550 GNDA.n2891 GNDA.n2871 585
R8551 GNDA.n2891 GNDA.n2890 585
R8552 GNDA.n2892 GNDA.n2868 585
R8553 GNDA.n2892 GNDA.n102 585
R8554 GNDA.n3037 GNDA.n3036 585
R8555 GNDA.n2624 GNDA.n2623 585
R8556 GNDA.n2744 GNDA.n2743 585
R8557 GNDA.n2745 GNDA.n2744 585
R8558 GNDA.n2621 GNDA.n2620 585
R8559 GNDA.n2746 GNDA.n2621 585
R8560 GNDA.n2749 GNDA.n2748 585
R8561 GNDA.n2748 GNDA.n2747 585
R8562 GNDA.n2750 GNDA.n2619 585
R8563 GNDA.n2622 GNDA.n2619 585
R8564 GNDA.n2752 GNDA.n2751 585
R8565 GNDA.n2752 GNDA.n108 585
R8566 GNDA.n2753 GNDA.n2618 585
R8567 GNDA.n2753 GNDA.n109 585
R8568 GNDA.n2756 GNDA.n2755 585
R8569 GNDA.n2755 GNDA.n2754 585
R8570 GNDA.n2757 GNDA.n2616 585
R8571 GNDA.n2616 GNDA.n2615 585
R8572 GNDA.n2759 GNDA.n2758 585
R8573 GNDA.n2760 GNDA.n2759 585
R8574 GNDA.n2617 GNDA.n2614 585
R8575 GNDA.n2761 GNDA.n2614 585
R8576 GNDA.n2763 GNDA.n2613 585
R8577 GNDA.n2763 GNDA.n2762 585
R8578 GNDA.n2740 GNDA.n103 585
R8579 GNDA.n5099 GNDA.n5098 585
R8580 GNDA.n5101 GNDA.n88 585
R8581 GNDA.n5172 GNDA.n5171 585
R8582 GNDA.n24 GNDA.n22 585
R8583 GNDA.n5270 GNDA.n5269 585
R8584 GNDA.n32 GNDA.n25 585
R8585 GNDA.n40 GNDA.n39 585
R8586 GNDA.n35 GNDA.n31 585
R8587 GNDA.n30 GNDA.n0 585
R8588 GNDA.n5106 GNDA.n1 585
R8589 GNDA.n5108 GNDA.n5107 585
R8590 GNDA.n5112 GNDA.n5111 585
R8591 GNDA.n5114 GNDA.n5113 585
R8592 GNDA.n5103 GNDA.n5102 585
R8593 GNDA.n5093 GNDA.n89 585
R8594 GNDA.n5097 GNDA.n89 585
R8595 GNDA.n5095 GNDA.n5094 585
R8596 GNDA.n5096 GNDA.n5095 585
R8597 GNDA.n5092 GNDA.n91 585
R8598 GNDA.n91 GNDA.n90 585
R8599 GNDA.n5091 GNDA.n5090 585
R8600 GNDA.n5090 GNDA.n5089 585
R8601 GNDA.n93 GNDA.n92 585
R8602 GNDA.n5088 GNDA.n93 585
R8603 GNDA.n4636 GNDA.n4635 585
R8604 GNDA.n4635 GNDA.n110 585
R8605 GNDA.n4638 GNDA.n4637 585
R8606 GNDA.n4639 GNDA.n4638 585
R8607 GNDA.n427 GNDA.n426 585
R8608 GNDA.n4640 GNDA.n427 585
R8609 GNDA.n4643 GNDA.n4642 585
R8610 GNDA.n4642 GNDA.n4641 585
R8611 GNDA.n4644 GNDA.n425 585
R8612 GNDA.n425 GNDA.n424 585
R8613 GNDA.n4646 GNDA.n4645 585
R8614 GNDA.n4647 GNDA.n4646 585
R8615 GNDA.n423 GNDA.n422 585
R8616 GNDA.n4648 GNDA.n423 585
R8617 GNDA.n4651 GNDA.n4650 585
R8618 GNDA.n4650 GNDA.n4649 585
R8619 GNDA.n4652 GNDA.n421 585
R8620 GNDA.n421 GNDA.n420 585
R8621 GNDA.n4654 GNDA.n4653 585
R8622 GNDA.n4655 GNDA.n4654 585
R8623 GNDA.n419 GNDA.n418 585
R8624 GNDA.n4656 GNDA.n419 585
R8625 GNDA.n4659 GNDA.n4658 585
R8626 GNDA.n4658 GNDA.n4657 585
R8627 GNDA.n4660 GNDA.n417 585
R8628 GNDA.n417 GNDA.n416 585
R8629 GNDA.n4662 GNDA.n4661 585
R8630 GNDA.n4663 GNDA.n4662 585
R8631 GNDA.n415 GNDA.n414 585
R8632 GNDA.n4664 GNDA.n415 585
R8633 GNDA.n4667 GNDA.n4666 585
R8634 GNDA.n4666 GNDA.n4665 585
R8635 GNDA.n4668 GNDA.n413 585
R8636 GNDA.n413 GNDA.n367 585
R8637 GNDA.n4670 GNDA.n4669 585
R8638 GNDA.n4671 GNDA.n4670 585
R8639 GNDA.n4675 GNDA.n4674 585
R8640 GNDA.n4674 GNDA.n4673 585
R8641 GNDA.n4676 GNDA.n363 585
R8642 GNDA.n363 GNDA.n362 585
R8643 GNDA.n4678 GNDA.n4677 585
R8644 GNDA.n4679 GNDA.n4678 585
R8645 GNDA.n364 GNDA.n361 585
R8646 GNDA.n4680 GNDA.n361 585
R8647 GNDA.n4682 GNDA.n360 585
R8648 GNDA.n4682 GNDA.n4681 585
R8649 GNDA.n4684 GNDA.n4683 585
R8650 GNDA.n4683 GNDA.n356 585
R8651 GNDA.n354 GNDA.n353 585
R8652 GNDA.n4690 GNDA.n354 585
R8653 GNDA.n4693 GNDA.n4692 585
R8654 GNDA.n4692 GNDA.n4691 585
R8655 GNDA.n4694 GNDA.n352 585
R8656 GNDA.n352 GNDA.n351 585
R8657 GNDA.n4696 GNDA.n4695 585
R8658 GNDA.n4697 GNDA.n4696 585
R8659 GNDA.n350 GNDA.n303 585
R8660 GNDA.n4698 GNDA.n350 585
R8661 GNDA.n4701 GNDA.n4700 585
R8662 GNDA.n4700 GNDA.n4699 585
R8663 GNDA.n389 GNDA.n83 585
R8664 GNDA.n390 GNDA.n388 585
R8665 GNDA.n395 GNDA.n386 585
R8666 GNDA.n396 GNDA.n384 585
R8667 GNDA.n397 GNDA.n383 585
R8668 GNDA.n381 GNDA.n379 585
R8669 GNDA.n403 GNDA.n378 585
R8670 GNDA.n404 GNDA.n376 585
R8671 GNDA.n405 GNDA.n375 585
R8672 GNDA.n373 GNDA.n371 585
R8673 GNDA.n410 GNDA.n370 585
R8674 GNDA.n411 GNDA.n366 585
R8675 GNDA.n5175 GNDA.n84 585
R8676 GNDA.n5175 GNDA.n5174 585
R8677 GNDA.n412 GNDA.n411 585
R8678 GNDA.n410 GNDA.n409 585
R8679 GNDA.n408 GNDA.n371 585
R8680 GNDA.n406 GNDA.n405 585
R8681 GNDA.n404 GNDA.n372 585
R8682 GNDA.n403 GNDA.n402 585
R8683 GNDA.n400 GNDA.n379 585
R8684 GNDA.n398 GNDA.n397 585
R8685 GNDA.n396 GNDA.n380 585
R8686 GNDA.n395 GNDA.n394 585
R8687 GNDA.n392 GNDA.n390 585
R8688 GNDA.n389 GNDA.n86 585
R8689 GNDA.n5173 GNDA.n84 585
R8690 GNDA.n5174 GNDA.n5173 585
R8691 GNDA.n2820 GNDA.n2819 585
R8692 GNDA.n2817 GNDA.n2578 585
R8693 GNDA.n2816 GNDA.n2815 585
R8694 GNDA.n2807 GNDA.n2580 585
R8695 GNDA.n2809 GNDA.n2808 585
R8696 GNDA.n2805 GNDA.n2582 585
R8697 GNDA.n2804 GNDA.n2803 585
R8698 GNDA.n2795 GNDA.n2584 585
R8699 GNDA.n2797 GNDA.n2796 585
R8700 GNDA.n2793 GNDA.n2586 585
R8701 GNDA.n2792 GNDA.n2791 585
R8702 GNDA.n2609 GNDA.n2588 585
R8703 GNDA.n2823 GNDA.n2575 585
R8704 GNDA.n2575 GNDA.n161 585
R8705 GNDA.n2788 GNDA.n2588 585
R8706 GNDA.n2791 GNDA.n2790 585
R8707 GNDA.n2586 GNDA.n2585 585
R8708 GNDA.n2585 GNDA.n111 585
R8709 GNDA.n2798 GNDA.n2797 585
R8710 GNDA.n2800 GNDA.n2584 585
R8711 GNDA.n2803 GNDA.n2802 585
R8712 GNDA.n2582 GNDA.n2581 585
R8713 GNDA.n2810 GNDA.n2809 585
R8714 GNDA.n2812 GNDA.n2580 585
R8715 GNDA.n2815 GNDA.n2814 585
R8716 GNDA.n2578 GNDA.n2577 585
R8717 GNDA.n2821 GNDA.n2820 585
R8718 GNDA.n2821 GNDA.n111 585
R8719 GNDA.n2823 GNDA.n2822 585
R8720 GNDA.n2822 GNDA.n161 585
R8721 GNDA.n2980 GNDA.n2979 585
R8722 GNDA.n2842 GNDA.n750 585
R8723 GNDA.n2844 GNDA.n2843 585
R8724 GNDA.n2849 GNDA.n2840 585
R8725 GNDA.n2850 GNDA.n2839 585
R8726 GNDA.n2851 GNDA.n2837 585
R8727 GNDA.n2836 GNDA.n2833 585
R8728 GNDA.n2856 GNDA.n2832 585
R8729 GNDA.n2857 GNDA.n2831 585
R8730 GNDA.n2828 GNDA.n2827 585
R8731 GNDA.n2918 GNDA.n2917 585
R8732 GNDA.n2920 GNDA.n2826 585
R8733 GNDA.n2914 GNDA.n2826 585
R8734 GNDA.n2917 GNDA.n2916 585
R8735 GNDA.n2859 GNDA.n2828 585
R8736 GNDA.n2859 GNDA.n711 585
R8737 GNDA.n2858 GNDA.n2857 585
R8738 GNDA.n2856 GNDA.n2855 585
R8739 GNDA.n2854 GNDA.n2833 585
R8740 GNDA.n2852 GNDA.n2851 585
R8741 GNDA.n2850 GNDA.n2834 585
R8742 GNDA.n2849 GNDA.n2848 585
R8743 GNDA.n2846 GNDA.n2844 585
R8744 GNDA.n750 GNDA.n749 585
R8745 GNDA.n2981 GNDA.n2980 585
R8746 GNDA.n2981 GNDA.n711 585
R8747 GNDA.n2292 GNDA.n2289 585
R8748 GNDA.n2294 GNDA.n2293 585
R8749 GNDA.n2293 GNDA.n675 585
R8750 GNDA.n2303 GNDA.n2302 585
R8751 GNDA.n2389 GNDA.n2388 585
R8752 GNDA.n2388 GNDA.n2387 585
R8753 GNDA.n2398 GNDA.n2278 585
R8754 GNDA.n2405 GNDA.n2277 585
R8755 GNDA.n2409 GNDA.n2277 585
R8756 GNDA.n2403 GNDA.n2402 585
R8757 GNDA.n3017 GNDA.n706 585
R8758 GNDA.n3020 GNDA.n3019 585
R8759 GNDA.n3021 GNDA.n3020 585
R8760 GNDA.n3012 GNDA.n3011 585
R8761 GNDA.n2973 GNDA.n811 585
R8762 GNDA.n2974 GNDA.n2973 585
R8763 GNDA.n2517 GNDA.n2516 585
R8764 GNDA.n2516 GNDA.n2515 585
R8765 GNDA.n2489 GNDA.n837 585
R8766 GNDA.n2514 GNDA.n837 585
R8767 GNDA.n2490 GNDA.n2248 585
R8768 GNDA.n2248 GNDA.n838 585
R8769 GNDA.n2498 GNDA.n2497 585
R8770 GNDA.n2499 GNDA.n2498 585
R8771 GNDA.n2252 GNDA.n2250 585
R8772 GNDA.n2250 GNDA.n2249 585
R8773 GNDA.n2414 GNDA.n2413 585
R8774 GNDA.n2413 GNDA.n106 585
R8775 GNDA.n2415 GNDA.n2411 585
R8776 GNDA.n2411 GNDA.n2410 585
R8777 GNDA.n2424 GNDA.n2423 585
R8778 GNDA.n2425 GNDA.n2424 585
R8779 GNDA.n2273 GNDA.n2272 585
R8780 GNDA.n2426 GNDA.n2273 585
R8781 GNDA.n2431 GNDA.n2430 585
R8782 GNDA.n2430 GNDA.n2429 585
R8783 GNDA.n2275 GNDA.n2274 585
R8784 GNDA.n2428 GNDA.n2275 585
R8785 GNDA.n2315 GNDA.n810 585
R8786 GNDA.n2427 GNDA.n810 585
R8787 GNDA.n2978 GNDA.n748 585
R8788 GNDA.n2978 GNDA.n2977 585
R8789 GNDA.n2317 GNDA.n811 585
R8790 GNDA.n2317 GNDA.n809 585
R8791 GNDA.n2323 GNDA.n2322 585
R8792 GNDA.n2322 GNDA.n2321 585
R8793 GNDA.n673 GNDA.n671 585
R8794 GNDA.n3063 GNDA.n673 585
R8795 GNDA.n3078 GNDA.n3077 585
R8796 GNDA.n3077 GNDA.n3076 585
R8797 GNDA.n3065 GNDA.n674 585
R8798 GNDA.n3075 GNDA.n674 585
R8799 GNDA.n3073 GNDA.n3072 585
R8800 GNDA.n3074 GNDA.n3073 585
R8801 GNDA.n3068 GNDA.n648 585
R8802 GNDA.n3064 GNDA.n648 585
R8803 GNDA.n3086 GNDA.n3085 585
R8804 GNDA.n3087 GNDA.n3086 585
R8805 GNDA.n650 GNDA.n649 585
R8806 GNDA.n2306 GNDA.n649 585
R8807 GNDA.n2310 GNDA.n2309 585
R8808 GNDA.n2309 GNDA.n2308 585
R8809 GNDA.n2313 GNDA.n2304 585
R8810 GNDA.n2307 GNDA.n2304 585
R8811 GNDA.n2382 GNDA.n2381 585
R8812 GNDA.n2383 GNDA.n2382 585
R8813 GNDA.n2379 GNDA.n806 585
R8814 GNDA.n2384 GNDA.n806 585
R8815 GNDA.n2982 GNDA.n748 585
R8816 GNDA.n2983 GNDA.n2982 585
R8817 GNDA.n803 GNDA.n747 585
R8818 GNDA.n2984 GNDA.n747 585
R8819 GNDA.n2986 GNDA.n745 585
R8820 GNDA.n2986 GNDA.n2985 585
R8821 GNDA.n3001 GNDA.n3000 585
R8822 GNDA.n3000 GNDA.n2999 585
R8823 GNDA.n2988 GNDA.n2987 585
R8824 GNDA.n2998 GNDA.n2987 585
R8825 GNDA.n2996 GNDA.n2995 585
R8826 GNDA.n2997 GNDA.n2996 585
R8827 GNDA.n2991 GNDA.n712 585
R8828 GNDA.n712 GNDA.n707 585
R8829 GNDA.n3009 GNDA.n3008 585
R8830 GNDA.n3010 GNDA.n3009 585
R8831 GNDA.n714 GNDA.n713 585
R8832 GNDA.n722 GNDA.n713 585
R8833 GNDA.n725 GNDA.n724 585
R8834 GNDA.n724 GNDA.n723 585
R8835 GNDA.n726 GNDA.n687 585
R8836 GNDA.n687 GNDA.n685 585
R8837 GNDA.n3046 GNDA.n3045 585
R8838 GNDA.n3047 GNDA.n3046 585
R8839 GNDA.n3043 GNDA.n688 585
R8840 GNDA.n688 GNDA.n686 585
R8841 GNDA.n2539 GNDA.n834 585
R8842 GNDA.n2538 GNDA.n2537 585
R8843 GNDA.n2536 GNDA.n2535 585
R8844 GNDA.n2534 GNDA.n2533 585
R8845 GNDA.n2532 GNDA.n2531 585
R8846 GNDA.n2530 GNDA.n2529 585
R8847 GNDA.n2528 GNDA.n2527 585
R8848 GNDA.n2526 GNDA.n2525 585
R8849 GNDA.n2524 GNDA.n2523 585
R8850 GNDA.n2522 GNDA.n2521 585
R8851 GNDA.n2520 GNDA.n2519 585
R8852 GNDA.n4867 GNDA.n280 585
R8853 GNDA.n262 GNDA.n261 585
R8854 GNDA.n264 GNDA.n263 585
R8855 GNDA.n266 GNDA.n265 585
R8856 GNDA.n268 GNDA.n267 585
R8857 GNDA.n270 GNDA.n269 585
R8858 GNDA.n272 GNDA.n271 585
R8859 GNDA.n274 GNDA.n273 585
R8860 GNDA.n275 GNDA.n240 585
R8861 GNDA.n278 GNDA.n277 585
R8862 GNDA.n276 GNDA.n239 585
R8863 GNDA.n229 GNDA.n228 585
R8864 GNDA.n4867 GNDA.n229 585
R8865 GNDA.n4870 GNDA.n4869 585
R8866 GNDA.n4870 GNDA.n227 585
R8867 GNDA.n4865 GNDA.n4864 585
R8868 GNDA.n4863 GNDA.n288 585
R8869 GNDA.n4862 GNDA.n287 585
R8870 GNDA.n4867 GNDA.n287 585
R8871 GNDA.n4861 GNDA.n4860 585
R8872 GNDA.n4859 GNDA.n4858 585
R8873 GNDA.n4857 GNDA.n4856 585
R8874 GNDA.n4855 GNDA.n4854 585
R8875 GNDA.n4853 GNDA.n4852 585
R8876 GNDA.n4851 GNDA.n4850 585
R8877 GNDA.n4849 GNDA.n4848 585
R8878 GNDA.n4847 GNDA.n4846 585
R8879 GNDA.n4845 GNDA.n4844 585
R8880 GNDA.n4844 GNDA.n4843 585
R8881 GNDA.n3860 GNDA.t129 524.808
R8882 GNDA.n4619 GNDA.t85 524.808
R8883 GNDA.n1749 GNDA.t60 524.808
R8884 GNDA.n3155 GNDA.t54 524.808
R8885 GNDA.n3137 GNDA.t79 508.743
R8886 GNDA.n3140 GNDA.t66 508.743
R8887 GNDA.n636 GNDA.t134 508.743
R8888 GNDA.n638 GNDA.t111 508.743
R8889 GNDA.n1321 GNDA.t103 499.442
R8890 GNDA.n3143 GNDA.t81 499.442
R8891 GNDA.n434 GNDA.t132 499.442
R8892 GNDA.n3147 GNDA.t114 499.442
R8893 GNDA.t45 GNDA.n88 486.94
R8894 GNDA.t45 GNDA.n103 486.94
R8895 GNDA.n3132 GNDA.t109 475.976
R8896 GNDA.n3132 GNDA.t74 475.976
R8897 GNDA.n631 GNDA.t99 475.976
R8898 GNDA.n631 GNDA.t101 475.976
R8899 GNDA.n680 GNDA.t116 425.134
R8900 GNDA.n2511 GNDA.t92 425.134
R8901 GNDA.n2242 GNDA.t41 409.067
R8902 GNDA.n3050 GNDA.t106 409.067
R8903 GNDA.n681 GNDA.t51 409.067
R8904 GNDA.n3060 GNDA.t69 409.067
R8905 GNDA.n2318 GNDA.t48 409.067
R8906 GNDA.n2502 GNDA.t138 409.067
R8907 GNDA.n4647 GNDA.n424 394.817
R8908 GNDA.n4641 GNDA.n4640 394.817
R8909 GNDA.n4640 GNDA.n4639 394.817
R8910 GNDA.n4639 GNDA.n110 394.817
R8911 GNDA.n5089 GNDA.n5088 394.817
R8912 GNDA.n5089 GNDA.n90 394.817
R8913 GNDA.n5096 GNDA.n90 394.817
R8914 GNDA.n5097 GNDA.n5096 394.817
R8915 GNDA.n5098 GNDA.n5097 394.817
R8916 GNDA.n5098 GNDA.n88 394.817
R8917 GNDA.n2762 GNDA.n2761 394.817
R8918 GNDA.n2761 GNDA.n2760 394.817
R8919 GNDA.n2760 GNDA.n2615 394.817
R8920 GNDA.n2754 GNDA.n2615 394.817
R8921 GNDA.n2754 GNDA.n109 394.817
R8922 GNDA.n2622 GNDA.n108 394.817
R8923 GNDA.n2747 GNDA.n2622 394.817
R8924 GNDA.n2747 GNDA.n2746 394.817
R8925 GNDA.n2746 GNDA.n2745 394.817
R8926 GNDA.n2745 GNDA.n2623 394.817
R8927 GNDA.n2623 GNDA.n103 394.817
R8928 GNDA.n2890 GNDA.n102 394.817
R8929 GNDA.n2890 GNDA.n2889 394.817
R8930 GNDA.n2889 GNDA.n2888 394.817
R8931 GNDA.n2888 GNDA.n2872 394.817
R8932 GNDA.n2872 GNDA.n709 394.817
R8933 GNDA.n2880 GNDA.n710 394.817
R8934 GNDA.n2880 GNDA.n2879 394.817
R8935 GNDA.n2879 GNDA.n695 394.817
R8936 GNDA.n3039 GNDA.n695 394.817
R8937 GNDA.n3039 GNDA.n3038 394.817
R8938 GNDA.n3038 GNDA.n3037 394.817
R8939 GNDA.n4634 GNDA.n424 377.269
R8940 GNDA.n300 GNDA.n96 370.214
R8941 GNDA.n4672 GNDA.n98 370.214
R8942 GNDA.n300 GNDA.n95 365.957
R8943 GNDA.n4672 GNDA.n97 365.957
R8944 GNDA.t45 GNDA.n94 172.876
R8945 GNDA.t45 GNDA.n95 327.661
R8946 GNDA.t45 GNDA.n97 327.661
R8947 GNDA.t45 GNDA.n647 172.876
R8948 GNDA.t45 GNDA.n646 172.615
R8949 GNDA.t45 GNDA.n96 323.404
R8950 GNDA.t45 GNDA.n98 323.404
R8951 GNDA.t45 GNDA.n711 172.615
R8952 GNDA.t67 GNDA.n3138 296.158
R8953 GNDA.n3139 GNDA.t67 296.158
R8954 GNDA.t112 GNDA.n637 296.158
R8955 GNDA.t112 GNDA.n639 296.158
R8956 GNDA.n433 GNDA.n431 292.5
R8957 GNDA.n1320 GNDA.n431 292.5
R8958 GNDA.t3 GNDA.n635 292.5
R8959 GNDA.t3 GNDA.n3136 292.5
R8960 GNDA.n3146 GNDA.n3145 292.5
R8961 GNDA.n3145 GNDA.n3144 292.5
R8962 GNDA.t45 GNDA.n110 267.598
R8963 GNDA.t45 GNDA.n109 267.598
R8964 GNDA.t45 GNDA.n709 267.598
R8965 GNDA.n3042 GNDA.n691 264.301
R8966 GNDA.n2742 GNDA.n2741 264.301
R8967 GNDA.n5100 GNDA.n87 264.301
R8968 GNDA.n2518 GNDA.n835 264.301
R8969 GNDA.n4868 GNDA.n4867 264.301
R8970 GNDA.n4867 GNDA.n234 264.301
R8971 GNDA.n3033 GNDA.t8 260
R8972 GNDA.n3031 GNDA.t8 260
R8973 GNDA.n2893 GNDA.n2892 259.416
R8974 GNDA.n2921 GNDA.n2920 259.416
R8975 GNDA.n2945 GNDA.n828 259.416
R8976 GNDA.n4674 GNDA.n366 259.416
R8977 GNDA.n2764 GNDA.n2763 259.416
R8978 GNDA.n2610 GNDA.n2609 259.416
R8979 GNDA.n5085 GNDA.n130 259.416
R8980 GNDA.n4704 GNDA.n301 259.416
R8981 GNDA.n4646 GNDA.n423 259.416
R8982 GNDA.n785 GNDA.n784 258.334
R8983 GNDA.n2342 GNDA.n2341 258.334
R8984 GNDA.n5030 GNDA.n5029 258.334
R8985 GNDA.n4815 GNDA.n4814 258.334
R8986 GNDA.n2683 GNDA.n2682 258.334
R8987 GNDA.n4954 GNDA.n4894 258.334
R8988 GNDA.n5233 GNDA.n80 258.334
R8989 GNDA.n2471 GNDA.n2258 258.334
R8990 GNDA.n5153 GNDA.n5152 258.334
R8991 GNDA.t45 GNDA.n4689 257.779
R8992 GNDA.n5087 GNDA.n5086 254.34
R8993 GNDA.n5087 GNDA.n128 254.34
R8994 GNDA.n5087 GNDA.n127 254.34
R8995 GNDA.n5087 GNDA.n126 254.34
R8996 GNDA.n5087 GNDA.n125 254.34
R8997 GNDA.n5087 GNDA.n124 254.34
R8998 GNDA.n5087 GNDA.n123 254.34
R8999 GNDA.n5087 GNDA.n122 254.34
R9000 GNDA.n5087 GNDA.n121 254.34
R9001 GNDA.n5087 GNDA.n120 254.34
R9002 GNDA.n5087 GNDA.n119 254.34
R9003 GNDA.n5087 GNDA.n118 254.34
R9004 GNDA.n5087 GNDA.n117 254.34
R9005 GNDA.n5087 GNDA.n116 254.34
R9006 GNDA.n5087 GNDA.n115 254.34
R9007 GNDA.n5087 GNDA.n114 254.34
R9008 GNDA.n5087 GNDA.n113 254.34
R9009 GNDA.n5087 GNDA.n112 254.34
R9010 GNDA.n5267 GNDA.n5266 254.34
R9011 GNDA.n5267 GNDA.n53 254.34
R9012 GNDA.n5267 GNDA.n52 254.34
R9013 GNDA.n5267 GNDA.n51 254.34
R9014 GNDA.n5267 GNDA.n50 254.34
R9015 GNDA.n5267 GNDA.n49 254.34
R9016 GNDA.n5267 GNDA.n48 254.34
R9017 GNDA.n5267 GNDA.n47 254.34
R9018 GNDA.n5267 GNDA.n46 254.34
R9019 GNDA.n5267 GNDA.n45 254.34
R9020 GNDA.n5267 GNDA.n44 254.34
R9021 GNDA.n5267 GNDA.n43 254.34
R9022 GNDA.n324 GNDA.n95 254.34
R9023 GNDA.n321 GNDA.n95 254.34
R9024 GNDA.n316 GNDA.n95 254.34
R9025 GNDA.n313 GNDA.n95 254.34
R9026 GNDA.n308 GNDA.n95 254.34
R9027 GNDA.n305 GNDA.n95 254.34
R9028 GNDA.n348 GNDA.n96 254.34
R9029 GNDA.n342 GNDA.n96 254.34
R9030 GNDA.n340 GNDA.n96 254.34
R9031 GNDA.n334 GNDA.n96 254.34
R9032 GNDA.n332 GNDA.n96 254.34
R9033 GNDA.n326 GNDA.n96 254.34
R9034 GNDA.n158 GNDA.n157 254.34
R9035 GNDA.n157 GNDA.n156 254.34
R9036 GNDA.n157 GNDA.n155 254.34
R9037 GNDA.n157 GNDA.n154 254.34
R9038 GNDA.n157 GNDA.n153 254.34
R9039 GNDA.n157 GNDA.n152 254.34
R9040 GNDA.n5080 GNDA.n5079 254.34
R9041 GNDA.n5079 GNDA.n5078 254.34
R9042 GNDA.n5079 GNDA.n140 254.34
R9043 GNDA.n5079 GNDA.n139 254.34
R9044 GNDA.n5079 GNDA.n138 254.34
R9045 GNDA.n5079 GNDA.n137 254.34
R9046 GNDA.n2971 GNDA.n94 254.34
R9047 GNDA.n819 GNDA.n94 254.34
R9048 GNDA.n2960 GNDA.n94 254.34
R9049 GNDA.n2957 GNDA.n94 254.34
R9050 GNDA.n2948 GNDA.n94 254.34
R9051 GNDA.n2946 GNDA.n94 254.34
R9052 GNDA.n2942 GNDA.n646 254.34
R9053 GNDA.n2953 GNDA.n646 254.34
R9054 GNDA.n824 GNDA.n646 254.34
R9055 GNDA.n2964 GNDA.n646 254.34
R9056 GNDA.n2967 GNDA.n646 254.34
R9057 GNDA.n2560 GNDA.n104 254.34
R9058 GNDA.n2558 GNDA.n104 254.34
R9059 GNDA.n2552 GNDA.n104 254.34
R9060 GNDA.n2550 GNDA.n104 254.34
R9061 GNDA.n2544 GNDA.n104 254.34
R9062 GNDA.n2542 GNDA.n104 254.34
R9063 GNDA.n2825 GNDA.n104 254.34
R9064 GNDA.n2926 GNDA.n104 254.34
R9065 GNDA.n2571 GNDA.n104 254.34
R9066 GNDA.n2933 GNDA.n104 254.34
R9067 GNDA.n2568 GNDA.n104 254.34
R9068 GNDA.n2940 GNDA.n104 254.34
R9069 GNDA.n2869 GNDA.n104 254.34
R9070 GNDA.n2898 GNDA.n104 254.34
R9071 GNDA.n2866 GNDA.n104 254.34
R9072 GNDA.n2905 GNDA.n104 254.34
R9073 GNDA.n2863 GNDA.n104 254.34
R9074 GNDA.n2912 GNDA.n104 254.34
R9075 GNDA.n4988 GNDA.n4987 254.34
R9076 GNDA.n4988 GNDA.n225 254.34
R9077 GNDA.n4988 GNDA.n224 254.34
R9078 GNDA.n4988 GNDA.n223 254.34
R9079 GNDA.n4988 GNDA.n222 254.34
R9080 GNDA.n4988 GNDA.n221 254.34
R9081 GNDA.n4988 GNDA.n163 254.34
R9082 GNDA.n4988 GNDA.n166 254.34
R9083 GNDA.n4988 GNDA.n220 254.34
R9084 GNDA.n4988 GNDA.n197 254.34
R9085 GNDA.n4988 GNDA.n196 254.34
R9086 GNDA.n4989 GNDA.n4988 254.34
R9087 GNDA.n4988 GNDA.n195 254.34
R9088 GNDA.n4988 GNDA.n194 254.34
R9089 GNDA.n4988 GNDA.n193 254.34
R9090 GNDA.n4988 GNDA.n192 254.34
R9091 GNDA.n4988 GNDA.n191 254.34
R9092 GNDA.n4988 GNDA.n190 254.34
R9093 GNDA.n5267 GNDA.n42 254.34
R9094 GNDA.n5268 GNDA.n5267 254.34
R9095 GNDA.n5267 GNDA.n41 254.34
R9096 GNDA.n5267 GNDA.n29 254.34
R9097 GNDA.n5267 GNDA.n28 254.34
R9098 GNDA.n5267 GNDA.n27 254.34
R9099 GNDA.n387 GNDA.n97 254.34
R9100 GNDA.n385 GNDA.n97 254.34
R9101 GNDA.n382 GNDA.n97 254.34
R9102 GNDA.n377 GNDA.n97 254.34
R9103 GNDA.n374 GNDA.n97 254.34
R9104 GNDA.n369 GNDA.n97 254.34
R9105 GNDA.n368 GNDA.n98 254.34
R9106 GNDA.n407 GNDA.n98 254.34
R9107 GNDA.n401 GNDA.n98 254.34
R9108 GNDA.n399 GNDA.n98 254.34
R9109 GNDA.n393 GNDA.n98 254.34
R9110 GNDA.n391 GNDA.n98 254.34
R9111 GNDA.n2818 GNDA.n101 254.34
R9112 GNDA.n2579 GNDA.n101 254.34
R9113 GNDA.n2806 GNDA.n101 254.34
R9114 GNDA.n2583 GNDA.n101 254.34
R9115 GNDA.n2794 GNDA.n101 254.34
R9116 GNDA.n2587 GNDA.n101 254.34
R9117 GNDA.n2789 GNDA.n111 254.34
R9118 GNDA.n2799 GNDA.n111 254.34
R9119 GNDA.n2801 GNDA.n111 254.34
R9120 GNDA.n2811 GNDA.n111 254.34
R9121 GNDA.n2813 GNDA.n111 254.34
R9122 GNDA.n805 GNDA.n647 254.34
R9123 GNDA.n2841 GNDA.n647 254.34
R9124 GNDA.n2838 GNDA.n647 254.34
R9125 GNDA.n2835 GNDA.n647 254.34
R9126 GNDA.n2830 GNDA.n647 254.34
R9127 GNDA.n2919 GNDA.n647 254.34
R9128 GNDA.n2915 GNDA.n711 254.34
R9129 GNDA.n2829 GNDA.n711 254.34
R9130 GNDA.n2853 GNDA.n711 254.34
R9131 GNDA.n2847 GNDA.n711 254.34
R9132 GNDA.n2845 GNDA.n711 254.34
R9133 GNDA.n4867 GNDA.n286 254.34
R9134 GNDA.n4867 GNDA.n285 254.34
R9135 GNDA.n4867 GNDA.n284 254.34
R9136 GNDA.n4867 GNDA.n283 254.34
R9137 GNDA.n4867 GNDA.n282 254.34
R9138 GNDA.n4867 GNDA.n281 254.34
R9139 GNDA.n4867 GNDA.n235 254.34
R9140 GNDA.n4867 GNDA.n236 254.34
R9141 GNDA.n4867 GNDA.n237 254.34
R9142 GNDA.n4867 GNDA.n238 254.34
R9143 GNDA.n4867 GNDA.n279 254.34
R9144 GNDA.n4867 GNDA.n4866 254.34
R9145 GNDA.n4867 GNDA.n230 254.34
R9146 GNDA.n4867 GNDA.n231 254.34
R9147 GNDA.n4867 GNDA.n232 254.34
R9148 GNDA.n4867 GNDA.n233 254.34
R9149 GNDA.n2291 GNDA.n675 250.349
R9150 GNDA.n2387 GNDA.n2386 250.349
R9151 GNDA.n2914 GNDA.n2913 249.663
R9152 GNDA.n2943 GNDA.n2941 249.663
R9153 GNDA.n2541 GNDA.n834 249.663
R9154 GNDA.n4700 GNDA.n349 249.663
R9155 GNDA.n2788 GNDA.n2787 249.663
R9156 GNDA.n5081 GNDA.n135 249.663
R9157 GNDA.n261 GNDA.n260 249.663
R9158 GNDA.n4865 GNDA.n289 249.663
R9159 GNDA.n4670 GNDA.n412 249.663
R9160 GNDA.n3020 GNDA.n706 246.25
R9161 GNDA.n3020 GNDA.n3011 246.25
R9162 GNDA.n2278 GNDA.n2277 246.25
R9163 GNDA.n2402 GNDA.n2277 246.25
R9164 GNDA.n3034 GNDA.n698 246.25
R9165 GNDA.n2409 GNDA.n2408 241.643
R9166 GNDA.n2409 GNDA.n2276 241.643
R9167 GNDA.n3022 GNDA.n3021 241.643
R9168 GNDA.n3021 GNDA.n708 241.643
R9169 GNDA.t256 GNDA.t93 227.873
R9170 GNDA.n3035 GNDA.t7 219.343
R9171 GNDA.n697 GNDA.t7 219.343
R9172 GNDA.n1273 GNDA.t1 197.133
R9173 GNDA.n1271 GNDA.t1 197.133
R9174 GNDA.n3127 GNDA.n3126 197.133
R9175 GNDA.n3100 GNDA.n3099 197.133
R9176 GNDA.n2388 GNDA.n2303 197
R9177 GNDA.n2293 GNDA.n2292 197
R9178 GNDA.n3036 GNDA.n688 197
R9179 GNDA.n2978 GNDA.n806 197
R9180 GNDA.n2973 GNDA.n810 197
R9181 GNDA.n2740 GNDA.n2739 197
R9182 GNDA.n2575 GNDA.n189 197
R9183 GNDA.n4897 GNDA.n4896 197
R9184 GNDA.n4748 GNDA.n85 197
R9185 GNDA.n5176 GNDA.n5175 197
R9186 GNDA.n5102 GNDA.n5101 197
R9187 GNDA.n2982 GNDA.n747 187.249
R9188 GNDA.n2322 GNDA.n2317 187.249
R9189 GNDA.n2516 GNDA.n280 187.249
R9190 GNDA.n2822 GNDA.n2576 187.249
R9191 GNDA.n5058 GNDA.n5057 187.249
R9192 GNDA.n4986 GNDA.n227 187.249
R9193 GNDA.n4843 GNDA.n4842 187.249
R9194 GNDA.n5265 GNDA.n55 187.249
R9195 GNDA.n5173 GNDA.n5172 187.249
R9196 GNDA.n786 GNDA.n785 185
R9197 GNDA.n788 GNDA.n787 185
R9198 GNDA.n790 GNDA.n789 185
R9199 GNDA.n792 GNDA.n791 185
R9200 GNDA.n794 GNDA.n793 185
R9201 GNDA.n796 GNDA.n795 185
R9202 GNDA.n798 GNDA.n797 185
R9203 GNDA.n800 GNDA.n799 185
R9204 GNDA.n801 GNDA.n743 185
R9205 GNDA.n768 GNDA.n767 185
R9206 GNDA.n770 GNDA.n769 185
R9207 GNDA.n772 GNDA.n771 185
R9208 GNDA.n774 GNDA.n773 185
R9209 GNDA.n776 GNDA.n775 185
R9210 GNDA.n778 GNDA.n777 185
R9211 GNDA.n780 GNDA.n779 185
R9212 GNDA.n782 GNDA.n781 185
R9213 GNDA.n784 GNDA.n783 185
R9214 GNDA.n735 GNDA.n690 185
R9215 GNDA.n752 GNDA.n751 185
R9216 GNDA.n754 GNDA.n753 185
R9217 GNDA.n756 GNDA.n755 185
R9218 GNDA.n758 GNDA.n757 185
R9219 GNDA.n760 GNDA.n759 185
R9220 GNDA.n762 GNDA.n761 185
R9221 GNDA.n764 GNDA.n763 185
R9222 GNDA.n766 GNDA.n765 185
R9223 GNDA.n734 GNDA.n689 185
R9224 GNDA.n728 GNDA.n727 185
R9225 GNDA.n721 GNDA.n716 185
R9226 GNDA.n3007 GNDA.n3006 185
R9227 GNDA.n2990 GNDA.n715 185
R9228 GNDA.n2994 GNDA.n2993 185
R9229 GNDA.n2992 GNDA.n2989 185
R9230 GNDA.n746 GNDA.n744 185
R9231 GNDA.n3003 GNDA.n3002 185
R9232 GNDA.n2341 GNDA.n2340 185
R9233 GNDA.n2339 GNDA.n2338 185
R9234 GNDA.n2337 GNDA.n2336 185
R9235 GNDA.n2335 GNDA.n2334 185
R9236 GNDA.n2333 GNDA.n2332 185
R9237 GNDA.n2331 GNDA.n2330 185
R9238 GNDA.n2329 GNDA.n2328 185
R9239 GNDA.n2327 GNDA.n2326 185
R9240 GNDA.n2325 GNDA.n669 185
R9241 GNDA.n2359 GNDA.n2358 185
R9242 GNDA.n2357 GNDA.n2356 185
R9243 GNDA.n2355 GNDA.n2354 185
R9244 GNDA.n2353 GNDA.n2352 185
R9245 GNDA.n2351 GNDA.n2350 185
R9246 GNDA.n2349 GNDA.n2348 185
R9247 GNDA.n2347 GNDA.n2346 185
R9248 GNDA.n2345 GNDA.n2344 185
R9249 GNDA.n2343 GNDA.n2342 185
R9250 GNDA.n2378 GNDA.n2377 185
R9251 GNDA.n2375 GNDA.n2374 185
R9252 GNDA.n2373 GNDA.n2372 185
R9253 GNDA.n2371 GNDA.n2370 185
R9254 GNDA.n2369 GNDA.n2368 185
R9255 GNDA.n2367 GNDA.n2366 185
R9256 GNDA.n2365 GNDA.n2364 185
R9257 GNDA.n2363 GNDA.n2362 185
R9258 GNDA.n2361 GNDA.n2360 185
R9259 GNDA.n2376 GNDA.n2314 185
R9260 GNDA.n2312 GNDA.n2311 185
R9261 GNDA.n2305 GNDA.n652 185
R9262 GNDA.n3084 GNDA.n3083 185
R9263 GNDA.n3067 GNDA.n651 185
R9264 GNDA.n3071 GNDA.n3070 185
R9265 GNDA.n3069 GNDA.n3066 185
R9266 GNDA.n672 GNDA.n670 185
R9267 GNDA.n3080 GNDA.n3079 185
R9268 GNDA.n5031 GNDA.n5030 185
R9269 GNDA.n5033 GNDA.n5032 185
R9270 GNDA.n5035 GNDA.n5034 185
R9271 GNDA.n5037 GNDA.n5036 185
R9272 GNDA.n5039 GNDA.n5038 185
R9273 GNDA.n5041 GNDA.n5040 185
R9274 GNDA.n5043 GNDA.n5042 185
R9275 GNDA.n5045 GNDA.n5044 185
R9276 GNDA.n5046 GNDA.n164 185
R9277 GNDA.n5013 GNDA.n5012 185
R9278 GNDA.n5015 GNDA.n5014 185
R9279 GNDA.n5017 GNDA.n5016 185
R9280 GNDA.n5019 GNDA.n5018 185
R9281 GNDA.n5021 GNDA.n5020 185
R9282 GNDA.n5023 GNDA.n5022 185
R9283 GNDA.n5025 GNDA.n5024 185
R9284 GNDA.n5027 GNDA.n5026 185
R9285 GNDA.n5029 GNDA.n5028 185
R9286 GNDA.n4995 GNDA.n4994 185
R9287 GNDA.n4997 GNDA.n4996 185
R9288 GNDA.n4999 GNDA.n4998 185
R9289 GNDA.n5001 GNDA.n5000 185
R9290 GNDA.n5003 GNDA.n5002 185
R9291 GNDA.n5005 GNDA.n5004 185
R9292 GNDA.n5007 GNDA.n5006 185
R9293 GNDA.n5009 GNDA.n5008 185
R9294 GNDA.n5011 GNDA.n5010 185
R9295 GNDA.n4993 GNDA.n4992 185
R9296 GNDA.n206 GNDA.n205 185
R9297 GNDA.n204 GNDA.n203 185
R9298 GNDA.n212 GNDA.n211 185
R9299 GNDA.n214 GNDA.n213 185
R9300 GNDA.n217 GNDA.n216 185
R9301 GNDA.n200 GNDA.n169 185
R9302 GNDA.n5050 GNDA.n5049 185
R9303 GNDA.n168 GNDA.n165 185
R9304 GNDA.n4816 GNDA.n4815 185
R9305 GNDA.n4818 GNDA.n4817 185
R9306 GNDA.n4820 GNDA.n4819 185
R9307 GNDA.n4822 GNDA.n4821 185
R9308 GNDA.n4824 GNDA.n4823 185
R9309 GNDA.n4826 GNDA.n4825 185
R9310 GNDA.n4828 GNDA.n4827 185
R9311 GNDA.n4830 GNDA.n4829 185
R9312 GNDA.n4831 GNDA.n4727 185
R9313 GNDA.n4798 GNDA.n4797 185
R9314 GNDA.n4800 GNDA.n4799 185
R9315 GNDA.n4802 GNDA.n4801 185
R9316 GNDA.n4804 GNDA.n4803 185
R9317 GNDA.n4806 GNDA.n4805 185
R9318 GNDA.n4808 GNDA.n4807 185
R9319 GNDA.n4810 GNDA.n4809 185
R9320 GNDA.n4812 GNDA.n4811 185
R9321 GNDA.n4814 GNDA.n4813 185
R9322 GNDA.n4780 GNDA.n4779 185
R9323 GNDA.n4782 GNDA.n4781 185
R9324 GNDA.n4784 GNDA.n4783 185
R9325 GNDA.n4786 GNDA.n4785 185
R9326 GNDA.n4788 GNDA.n4787 185
R9327 GNDA.n4790 GNDA.n4789 185
R9328 GNDA.n4792 GNDA.n4791 185
R9329 GNDA.n4794 GNDA.n4793 185
R9330 GNDA.n4796 GNDA.n4795 185
R9331 GNDA.n2684 GNDA.n2683 185
R9332 GNDA.n2686 GNDA.n2685 185
R9333 GNDA.n2688 GNDA.n2687 185
R9334 GNDA.n2690 GNDA.n2689 185
R9335 GNDA.n2692 GNDA.n2691 185
R9336 GNDA.n2694 GNDA.n2693 185
R9337 GNDA.n2696 GNDA.n2695 185
R9338 GNDA.n2698 GNDA.n2697 185
R9339 GNDA.n2699 GNDA.n2647 185
R9340 GNDA.n2666 GNDA.n2665 185
R9341 GNDA.n2668 GNDA.n2667 185
R9342 GNDA.n2670 GNDA.n2669 185
R9343 GNDA.n2672 GNDA.n2671 185
R9344 GNDA.n2674 GNDA.n2673 185
R9345 GNDA.n2676 GNDA.n2675 185
R9346 GNDA.n2678 GNDA.n2677 185
R9347 GNDA.n2680 GNDA.n2679 185
R9348 GNDA.n2682 GNDA.n2681 185
R9349 GNDA.n2639 GNDA.n2625 185
R9350 GNDA.n2650 GNDA.n2649 185
R9351 GNDA.n2652 GNDA.n2651 185
R9352 GNDA.n2654 GNDA.n2653 185
R9353 GNDA.n2656 GNDA.n2655 185
R9354 GNDA.n2658 GNDA.n2657 185
R9355 GNDA.n2660 GNDA.n2659 185
R9356 GNDA.n2662 GNDA.n2661 185
R9357 GNDA.n2664 GNDA.n2663 185
R9358 GNDA.n2629 GNDA.n2626 185
R9359 GNDA.n2732 GNDA.n2731 185
R9360 GNDA.n2705 GNDA.n2628 185
R9361 GNDA.n2711 GNDA.n2710 185
R9362 GNDA.n2709 GNDA.n2704 185
R9363 GNDA.n2718 GNDA.n2717 185
R9364 GNDA.n2716 GNDA.n2703 185
R9365 GNDA.n2723 GNDA.n2648 185
R9366 GNDA.n2728 GNDA.n2727 185
R9367 GNDA.n4956 GNDA.n4894 185
R9368 GNDA.n4970 GNDA.n4969 185
R9369 GNDA.n4968 GNDA.n4895 185
R9370 GNDA.n4967 GNDA.n4966 185
R9371 GNDA.n4965 GNDA.n4964 185
R9372 GNDA.n4963 GNDA.n4962 185
R9373 GNDA.n4961 GNDA.n4960 185
R9374 GNDA.n4959 GNDA.n4958 185
R9375 GNDA.n4957 GNDA.n4871 185
R9376 GNDA.n4939 GNDA.n4938 185
R9377 GNDA.n4941 GNDA.n4940 185
R9378 GNDA.n4943 GNDA.n4942 185
R9379 GNDA.n4945 GNDA.n4944 185
R9380 GNDA.n4947 GNDA.n4946 185
R9381 GNDA.n4949 GNDA.n4948 185
R9382 GNDA.n4951 GNDA.n4950 185
R9383 GNDA.n4953 GNDA.n4952 185
R9384 GNDA.n4955 GNDA.n4954 185
R9385 GNDA.n4921 GNDA.n4920 185
R9386 GNDA.n4923 GNDA.n4922 185
R9387 GNDA.n4925 GNDA.n4924 185
R9388 GNDA.n4927 GNDA.n4926 185
R9389 GNDA.n4929 GNDA.n4928 185
R9390 GNDA.n4931 GNDA.n4930 185
R9391 GNDA.n4933 GNDA.n4932 185
R9392 GNDA.n4935 GNDA.n4934 185
R9393 GNDA.n4937 GNDA.n4936 185
R9394 GNDA.n4919 GNDA.n4918 185
R9395 GNDA.n4913 GNDA.n4912 185
R9396 GNDA.n4911 GNDA.n4910 185
R9397 GNDA.n4906 GNDA.n4905 185
R9398 GNDA.n4901 GNDA.n4879 185
R9399 GNDA.n4974 GNDA.n4973 185
R9400 GNDA.n4878 GNDA.n4876 185
R9401 GNDA.n4980 GNDA.n4979 185
R9402 GNDA.n4982 GNDA.n4981 185
R9403 GNDA.n3023 GNDA.n705 185
R9404 GNDA.n3015 GNDA.n3014 185
R9405 GNDA.n2407 GNDA.n2406 185
R9406 GNDA.n2406 GNDA.n2405 185
R9407 GNDA.n2407 GNDA.n2397 185
R9408 GNDA.n2400 GNDA.n2397 185
R9409 GNDA.n5235 GNDA.n80 185
R9410 GNDA.n5249 GNDA.n5248 185
R9411 GNDA.n5247 GNDA.n81 185
R9412 GNDA.n5246 GNDA.n5245 185
R9413 GNDA.n5244 GNDA.n5243 185
R9414 GNDA.n5242 GNDA.n5241 185
R9415 GNDA.n5240 GNDA.n5239 185
R9416 GNDA.n5238 GNDA.n5237 185
R9417 GNDA.n5236 GNDA.n57 185
R9418 GNDA.n5218 GNDA.n5217 185
R9419 GNDA.n5220 GNDA.n5219 185
R9420 GNDA.n5222 GNDA.n5221 185
R9421 GNDA.n5224 GNDA.n5223 185
R9422 GNDA.n5226 GNDA.n5225 185
R9423 GNDA.n5228 GNDA.n5227 185
R9424 GNDA.n5230 GNDA.n5229 185
R9425 GNDA.n5232 GNDA.n5231 185
R9426 GNDA.n5234 GNDA.n5233 185
R9427 GNDA.n5200 GNDA.n5199 185
R9428 GNDA.n5202 GNDA.n5201 185
R9429 GNDA.n5204 GNDA.n5203 185
R9430 GNDA.n5206 GNDA.n5205 185
R9431 GNDA.n5208 GNDA.n5207 185
R9432 GNDA.n5210 GNDA.n5209 185
R9433 GNDA.n5212 GNDA.n5211 185
R9434 GNDA.n5214 GNDA.n5213 185
R9435 GNDA.n5216 GNDA.n5215 185
R9436 GNDA.n5198 GNDA.n5197 185
R9437 GNDA.n5192 GNDA.n5191 185
R9438 GNDA.n5190 GNDA.n5189 185
R9439 GNDA.n5185 GNDA.n5184 185
R9440 GNDA.n5180 GNDA.n65 185
R9441 GNDA.n5253 GNDA.n5252 185
R9442 GNDA.n64 GNDA.n62 185
R9443 GNDA.n5259 GNDA.n5258 185
R9444 GNDA.n5261 GNDA.n5260 185
R9445 GNDA.n4778 GNDA.n4777 185
R9446 GNDA.n4772 GNDA.n4771 185
R9447 GNDA.n4770 GNDA.n4769 185
R9448 GNDA.n4765 GNDA.n4764 185
R9449 GNDA.n4763 GNDA.n4762 185
R9450 GNDA.n4757 GNDA.n4756 185
R9451 GNDA.n4752 GNDA.n4731 185
R9452 GNDA.n4835 GNDA.n4834 185
R9453 GNDA.n4730 GNDA.n4728 185
R9454 GNDA.n2471 GNDA.n2470 185
R9455 GNDA.n2473 GNDA.n2257 185
R9456 GNDA.n2476 GNDA.n2475 185
R9457 GNDA.n2477 GNDA.n2256 185
R9458 GNDA.n2479 GNDA.n2478 185
R9459 GNDA.n2481 GNDA.n2255 185
R9460 GNDA.n2484 GNDA.n2483 185
R9461 GNDA.n2485 GNDA.n2254 185
R9462 GNDA.n2487 GNDA.n2486 185
R9463 GNDA.n2453 GNDA.n2262 185
R9464 GNDA.n2455 GNDA.n2454 185
R9465 GNDA.n2457 GNDA.n2261 185
R9466 GNDA.n2460 GNDA.n2459 185
R9467 GNDA.n2461 GNDA.n2260 185
R9468 GNDA.n2463 GNDA.n2462 185
R9469 GNDA.n2465 GNDA.n2259 185
R9470 GNDA.n2468 GNDA.n2467 185
R9471 GNDA.n2469 GNDA.n2258 185
R9472 GNDA.n2437 GNDA.n2436 185
R9473 GNDA.n2438 GNDA.n2267 185
R9474 GNDA.n2440 GNDA.n2439 185
R9475 GNDA.n2442 GNDA.n2265 185
R9476 GNDA.n2444 GNDA.n2443 185
R9477 GNDA.n2445 GNDA.n2264 185
R9478 GNDA.n2447 GNDA.n2446 185
R9479 GNDA.n2449 GNDA.n2263 185
R9480 GNDA.n2452 GNDA.n2451 185
R9481 GNDA.n2435 GNDA.n2270 185
R9482 GNDA.n2433 GNDA.n2432 185
R9483 GNDA.n2422 GNDA.n2271 185
R9484 GNDA.n2421 GNDA.n2420 185
R9485 GNDA.n2418 GNDA.n2416 185
R9486 GNDA.n2412 GNDA.n2253 185
R9487 GNDA.n2496 GNDA.n2495 185
R9488 GNDA.n2493 GNDA.n2251 185
R9489 GNDA.n2492 GNDA.n2491 185
R9490 GNDA.n5154 GNDA.n5153 185
R9491 GNDA.n5156 GNDA.n5155 185
R9492 GNDA.n5158 GNDA.n5157 185
R9493 GNDA.n5160 GNDA.n5159 185
R9494 GNDA.n5162 GNDA.n5161 185
R9495 GNDA.n5164 GNDA.n5163 185
R9496 GNDA.n5166 GNDA.n5165 185
R9497 GNDA.n5168 GNDA.n5167 185
R9498 GNDA.n5169 GNDA.n20 185
R9499 GNDA.n5136 GNDA.n5135 185
R9500 GNDA.n5138 GNDA.n5137 185
R9501 GNDA.n5140 GNDA.n5139 185
R9502 GNDA.n5142 GNDA.n5141 185
R9503 GNDA.n5144 GNDA.n5143 185
R9504 GNDA.n5146 GNDA.n5145 185
R9505 GNDA.n5148 GNDA.n5147 185
R9506 GNDA.n5150 GNDA.n5149 185
R9507 GNDA.n5152 GNDA.n5151 185
R9508 GNDA.n5118 GNDA.n5117 185
R9509 GNDA.n5120 GNDA.n5119 185
R9510 GNDA.n5122 GNDA.n5121 185
R9511 GNDA.n5124 GNDA.n5123 185
R9512 GNDA.n5126 GNDA.n5125 185
R9513 GNDA.n5128 GNDA.n5127 185
R9514 GNDA.n5130 GNDA.n5129 185
R9515 GNDA.n5132 GNDA.n5131 185
R9516 GNDA.n5134 GNDA.n5133 185
R9517 GNDA.n5116 GNDA.n5115 185
R9518 GNDA.n5110 GNDA.n5109 185
R9519 GNDA.n5105 GNDA.n3 185
R9520 GNDA.n5276 GNDA.n5275 185
R9521 GNDA.n34 GNDA.n2 185
R9522 GNDA.n38 GNDA.n37 185
R9523 GNDA.n36 GNDA.n33 185
R9524 GNDA.n23 GNDA.n21 185
R9525 GNDA.n5272 GNDA.n5271 185
R9526 GNDA.n2892 GNDA.n2891 175.546
R9527 GNDA.n2891 GNDA.n2870 175.546
R9528 GNDA.n2887 GNDA.n2870 175.546
R9529 GNDA.n2887 GNDA.n2873 175.546
R9530 GNDA.n2883 GNDA.n2873 175.546
R9531 GNDA.n2883 GNDA.n2882 175.546
R9532 GNDA.n2882 GNDA.n2881 175.546
R9533 GNDA.n2881 GNDA.n2876 175.546
R9534 GNDA.n2876 GNDA.n693 175.546
R9535 GNDA.n3040 GNDA.n693 175.546
R9536 GNDA.n3040 GNDA.n694 175.546
R9537 GNDA.n2986 GNDA.n747 175.546
R9538 GNDA.n3000 GNDA.n2986 175.546
R9539 GNDA.n3000 GNDA.n2987 175.546
R9540 GNDA.n2996 GNDA.n2987 175.546
R9541 GNDA.n2996 GNDA.n712 175.546
R9542 GNDA.n3009 GNDA.n712 175.546
R9543 GNDA.n3009 GNDA.n713 175.546
R9544 GNDA.n724 GNDA.n713 175.546
R9545 GNDA.n724 GNDA.n687 175.546
R9546 GNDA.n3046 GNDA.n687 175.546
R9547 GNDA.n3046 GNDA.n688 175.546
R9548 GNDA.n2916 GNDA.n2859 175.546
R9549 GNDA.n2859 GNDA.n2858 175.546
R9550 GNDA.n2855 GNDA.n2854 175.546
R9551 GNDA.n2852 GNDA.n2834 175.546
R9552 GNDA.n2848 GNDA.n2846 175.546
R9553 GNDA.n2981 GNDA.n749 175.546
R9554 GNDA.n2911 GNDA.n2861 175.546
R9555 GNDA.n2907 GNDA.n2906 175.546
R9556 GNDA.n2904 GNDA.n2864 175.546
R9557 GNDA.n2900 GNDA.n2899 175.546
R9558 GNDA.n2897 GNDA.n2867 175.546
R9559 GNDA.n2918 GNDA.n2827 175.546
R9560 GNDA.n2832 GNDA.n2831 175.546
R9561 GNDA.n2837 GNDA.n2836 175.546
R9562 GNDA.n2840 GNDA.n2839 175.546
R9563 GNDA.n2843 GNDA.n2842 175.546
R9564 GNDA.n2939 GNDA.n2566 175.546
R9565 GNDA.n2935 GNDA.n2934 175.546
R9566 GNDA.n2932 GNDA.n2569 175.546
R9567 GNDA.n2928 GNDA.n2927 175.546
R9568 GNDA.n2925 GNDA.n2572 175.546
R9569 GNDA.n2322 GNDA.n673 175.546
R9570 GNDA.n3077 GNDA.n673 175.546
R9571 GNDA.n3077 GNDA.n674 175.546
R9572 GNDA.n3073 GNDA.n674 175.546
R9573 GNDA.n3073 GNDA.n648 175.546
R9574 GNDA.n3086 GNDA.n648 175.546
R9575 GNDA.n3086 GNDA.n649 175.546
R9576 GNDA.n2309 GNDA.n649 175.546
R9577 GNDA.n2309 GNDA.n2304 175.546
R9578 GNDA.n2382 GNDA.n2304 175.546
R9579 GNDA.n2382 GNDA.n806 175.546
R9580 GNDA.n2951 GNDA.n826 175.546
R9581 GNDA.n2952 GNDA.n2951 175.546
R9582 GNDA.n2954 GNDA.n825 175.546
R9583 GNDA.n2963 GNDA.n817 175.546
R9584 GNDA.n2966 GNDA.n2965 175.546
R9585 GNDA.n2968 GNDA.n815 175.546
R9586 GNDA.n2537 GNDA.n2536 175.546
R9587 GNDA.n2533 GNDA.n2532 175.546
R9588 GNDA.n2529 GNDA.n2528 175.546
R9589 GNDA.n2525 GNDA.n2524 175.546
R9590 GNDA.n2521 GNDA.n2520 175.546
R9591 GNDA.n2545 GNDA.n2543 175.546
R9592 GNDA.n2549 GNDA.n832 175.546
R9593 GNDA.n2553 GNDA.n2551 175.546
R9594 GNDA.n2557 GNDA.n830 175.546
R9595 GNDA.n2561 GNDA.n2559 175.546
R9596 GNDA.n2516 GNDA.n837 175.546
R9597 GNDA.n2248 GNDA.n837 175.546
R9598 GNDA.n2498 GNDA.n2248 175.546
R9599 GNDA.n2498 GNDA.n2250 175.546
R9600 GNDA.n2413 GNDA.n2250 175.546
R9601 GNDA.n2413 GNDA.n2411 175.546
R9602 GNDA.n2424 GNDA.n2411 175.546
R9603 GNDA.n2424 GNDA.n2273 175.546
R9604 GNDA.n2430 GNDA.n2273 175.546
R9605 GNDA.n2430 GNDA.n2275 175.546
R9606 GNDA.n2275 GNDA.n810 175.546
R9607 GNDA.n2949 GNDA.n2947 175.546
R9608 GNDA.n2956 GNDA.n822 175.546
R9609 GNDA.n2959 GNDA.n2958 175.546
R9610 GNDA.n2961 GNDA.n820 175.546
R9611 GNDA.n2970 GNDA.n813 175.546
R9612 GNDA.n373 GNDA.n370 175.546
R9613 GNDA.n376 GNDA.n375 175.546
R9614 GNDA.n381 GNDA.n378 175.546
R9615 GNDA.n384 GNDA.n383 175.546
R9616 GNDA.n388 GNDA.n386 175.546
R9617 GNDA.n4700 GNDA.n350 175.546
R9618 GNDA.n4696 GNDA.n350 175.546
R9619 GNDA.n4696 GNDA.n352 175.546
R9620 GNDA.n4692 GNDA.n352 175.546
R9621 GNDA.n4692 GNDA.n354 175.546
R9622 GNDA.n4683 GNDA.n354 175.546
R9623 GNDA.n4683 GNDA.n4682 175.546
R9624 GNDA.n4682 GNDA.n361 175.546
R9625 GNDA.n4678 GNDA.n361 175.546
R9626 GNDA.n4678 GNDA.n363 175.546
R9627 GNDA.n4674 GNDA.n363 175.546
R9628 GNDA.n347 GNDA.n304 175.546
R9629 GNDA.n343 GNDA.n341 175.546
R9630 GNDA.n339 GNDA.n311 175.546
R9631 GNDA.n335 GNDA.n333 175.546
R9632 GNDA.n331 GNDA.n319 175.546
R9633 GNDA.n2763 GNDA.n2614 175.546
R9634 GNDA.n2759 GNDA.n2614 175.546
R9635 GNDA.n2759 GNDA.n2616 175.546
R9636 GNDA.n2755 GNDA.n2616 175.546
R9637 GNDA.n2755 GNDA.n2753 175.546
R9638 GNDA.n2753 GNDA.n2752 175.546
R9639 GNDA.n2752 GNDA.n2619 175.546
R9640 GNDA.n2748 GNDA.n2619 175.546
R9641 GNDA.n2748 GNDA.n2621 175.546
R9642 GNDA.n2744 GNDA.n2621 175.546
R9643 GNDA.n2744 GNDA.n2624 175.546
R9644 GNDA.n2725 GNDA.n2724 175.546
R9645 GNDA.n2721 GNDA.n2720 175.546
R9646 GNDA.n2714 GNDA.n2713 175.546
R9647 GNDA.n2707 GNDA.n2706 175.546
R9648 GNDA.n2735 GNDA.n2734 175.546
R9649 GNDA.n2790 GNDA.n2585 175.546
R9650 GNDA.n2798 GNDA.n2585 175.546
R9651 GNDA.n2802 GNDA.n2800 175.546
R9652 GNDA.n2810 GNDA.n2581 175.546
R9653 GNDA.n2814 GNDA.n2812 175.546
R9654 GNDA.n2821 GNDA.n2577 175.546
R9655 GNDA.n2784 GNDA.n2783 175.546
R9656 GNDA.n2780 GNDA.n2779 175.546
R9657 GNDA.n2776 GNDA.n2775 175.546
R9658 GNDA.n2772 GNDA.n2771 175.546
R9659 GNDA.n2768 GNDA.n2767 175.546
R9660 GNDA.n2793 GNDA.n2792 175.546
R9661 GNDA.n2796 GNDA.n2795 175.546
R9662 GNDA.n2805 GNDA.n2804 175.546
R9663 GNDA.n2808 GNDA.n2807 175.546
R9664 GNDA.n2817 GNDA.n2816 175.546
R9665 GNDA.n5053 GNDA.n5052 175.546
R9666 GNDA.n219 GNDA.n199 175.546
R9667 GNDA.n201 GNDA.n198 175.546
R9668 GNDA.n209 GNDA.n208 175.546
R9669 GNDA.n4990 GNDA.n188 175.546
R9670 GNDA.n5077 GNDA.n136 175.546
R9671 GNDA.n5073 GNDA.n141 175.546
R9672 GNDA.n5071 GNDA.n5070 175.546
R9673 GNDA.n5067 GNDA.n5066 175.546
R9674 GNDA.n5063 GNDA.n5062 175.546
R9675 GNDA.n2591 GNDA.n2590 175.546
R9676 GNDA.n2595 GNDA.n2594 175.546
R9677 GNDA.n2599 GNDA.n2598 175.546
R9678 GNDA.n2603 GNDA.n2602 175.546
R9679 GNDA.n2607 GNDA.n2606 175.546
R9680 GNDA.n151 GNDA.n142 175.546
R9681 GNDA.n144 GNDA.n143 175.546
R9682 GNDA.n146 GNDA.n145 175.546
R9683 GNDA.n148 GNDA.n147 175.546
R9684 GNDA.n150 GNDA.n149 175.546
R9685 GNDA.n4872 GNDA.n226 175.546
R9686 GNDA.n4977 GNDA.n4976 175.546
R9687 GNDA.n4903 GNDA.n4902 175.546
R9688 GNDA.n4908 GNDA.n4907 175.546
R9689 GNDA.n4916 GNDA.n4915 175.546
R9690 GNDA.n265 GNDA.n264 175.546
R9691 GNDA.n269 GNDA.n268 175.546
R9692 GNDA.n273 GNDA.n272 175.546
R9693 GNDA.n278 GNDA.n240 175.546
R9694 GNDA.n239 GNDA.n229 175.546
R9695 GNDA.n4869 GNDA.n229 175.546
R9696 GNDA.n257 GNDA.n256 175.546
R9697 GNDA.n253 GNDA.n252 175.546
R9698 GNDA.n249 GNDA.n248 175.546
R9699 GNDA.n245 GNDA.n244 175.546
R9700 GNDA.n241 GNDA.n129 175.546
R9701 GNDA.n307 GNDA.n306 175.546
R9702 GNDA.n312 GNDA.n309 175.546
R9703 GNDA.n315 GNDA.n314 175.546
R9704 GNDA.n320 GNDA.n317 175.546
R9705 GNDA.n323 GNDA.n322 175.546
R9706 GNDA.n4838 GNDA.n4837 175.546
R9707 GNDA.n4754 GNDA.n4753 175.546
R9708 GNDA.n4760 GNDA.n4759 175.546
R9709 GNDA.n4767 GNDA.n4766 175.546
R9710 GNDA.n4775 GNDA.n4774 175.546
R9711 GNDA.n288 GNDA.n287 175.546
R9712 GNDA.n4860 GNDA.n287 175.546
R9713 GNDA.n4858 GNDA.n4857 175.546
R9714 GNDA.n4854 GNDA.n4853 175.546
R9715 GNDA.n4850 GNDA.n4849 175.546
R9716 GNDA.n4846 GNDA.n4845 175.546
R9717 GNDA.n4724 GNDA.n289 175.546
R9718 GNDA.n4724 GNDA.n291 175.546
R9719 GNDA.n4720 GNDA.n291 175.546
R9720 GNDA.n4720 GNDA.n293 175.546
R9721 GNDA.n4716 GNDA.n293 175.546
R9722 GNDA.n4716 GNDA.n295 175.546
R9723 GNDA.n4712 GNDA.n295 175.546
R9724 GNDA.n4712 GNDA.n297 175.546
R9725 GNDA.n4708 GNDA.n297 175.546
R9726 GNDA.n4708 GNDA.n299 175.546
R9727 GNDA.n4704 GNDA.n299 175.546
R9728 GNDA.n58 GNDA.n54 175.546
R9729 GNDA.n5256 GNDA.n5255 175.546
R9730 GNDA.n5182 GNDA.n5181 175.546
R9731 GNDA.n5187 GNDA.n5186 175.546
R9732 GNDA.n5195 GNDA.n5194 175.546
R9733 GNDA.n409 GNDA.n408 175.546
R9734 GNDA.n406 GNDA.n372 175.546
R9735 GNDA.n402 GNDA.n400 175.546
R9736 GNDA.n398 GNDA.n380 175.546
R9737 GNDA.n394 GNDA.n392 175.546
R9738 GNDA.n4670 GNDA.n413 175.546
R9739 GNDA.n4666 GNDA.n413 175.546
R9740 GNDA.n4666 GNDA.n415 175.546
R9741 GNDA.n4662 GNDA.n415 175.546
R9742 GNDA.n4662 GNDA.n417 175.546
R9743 GNDA.n4658 GNDA.n417 175.546
R9744 GNDA.n4658 GNDA.n419 175.546
R9745 GNDA.n4654 GNDA.n419 175.546
R9746 GNDA.n4654 GNDA.n421 175.546
R9747 GNDA.n4650 GNDA.n421 175.546
R9748 GNDA.n4650 GNDA.n423 175.546
R9749 GNDA.n5269 GNDA.n24 175.546
R9750 GNDA.n40 GNDA.n25 175.546
R9751 GNDA.n31 GNDA.n30 175.546
R9752 GNDA.n5107 GNDA.n5106 175.546
R9753 GNDA.n5113 GNDA.n5112 175.546
R9754 GNDA.n4646 GNDA.n425 175.546
R9755 GNDA.n4642 GNDA.n425 175.546
R9756 GNDA.n4642 GNDA.n427 175.546
R9757 GNDA.n4638 GNDA.n427 175.546
R9758 GNDA.n4638 GNDA.n4635 175.546
R9759 GNDA.n4635 GNDA.n93 175.546
R9760 GNDA.n5090 GNDA.n93 175.546
R9761 GNDA.n5090 GNDA.n91 175.546
R9762 GNDA.n5095 GNDA.n91 175.546
R9763 GNDA.n5095 GNDA.n89 175.546
R9764 GNDA.n5099 GNDA.n89 175.546
R9765 GNDA.n157 GNDA.n100 173.881
R9766 GNDA.t45 GNDA.n101 172.876
R9767 GNDA.t45 GNDA.n111 172.615
R9768 GNDA.n5079 GNDA.n100 171.624
R9769 GNDA.n735 GNDA.n734 163.333
R9770 GNDA.n2377 GNDA.n2376 163.333
R9771 GNDA.n4994 GNDA.n4993 163.333
R9772 GNDA.n4779 GNDA.n4778 163.333
R9773 GNDA.n2639 GNDA.n2629 163.333
R9774 GNDA.n4920 GNDA.n4919 163.333
R9775 GNDA.n5199 GNDA.n5198 163.333
R9776 GNDA.n2436 GNDA.n2435 163.333
R9777 GNDA.n5117 GNDA.n5116 163.333
R9778 GNDA.n3133 GNDA.n3132 161.3
R9779 GNDA.n632 GNDA.n631 161.3
R9780 GNDA.n4688 GNDA.n355 157.601
R9781 GNDA.n781 GNDA.n780 150
R9782 GNDA.n777 GNDA.n776 150
R9783 GNDA.n773 GNDA.n772 150
R9784 GNDA.n769 GNDA.n768 150
R9785 GNDA.n765 GNDA.n764 150
R9786 GNDA.n761 GNDA.n760 150
R9787 GNDA.n757 GNDA.n756 150
R9788 GNDA.n753 GNDA.n752 150
R9789 GNDA.n3003 GNDA.n744 150
R9790 GNDA.n2993 GNDA.n2992 150
R9791 GNDA.n3006 GNDA.n715 150
R9792 GNDA.n728 GNDA.n716 150
R9793 GNDA.n789 GNDA.n788 150
R9794 GNDA.n793 GNDA.n792 150
R9795 GNDA.n797 GNDA.n796 150
R9796 GNDA.n799 GNDA.n743 150
R9797 GNDA.n2346 GNDA.n2345 150
R9798 GNDA.n2350 GNDA.n2349 150
R9799 GNDA.n2354 GNDA.n2353 150
R9800 GNDA.n2358 GNDA.n2357 150
R9801 GNDA.n2362 GNDA.n2361 150
R9802 GNDA.n2366 GNDA.n2365 150
R9803 GNDA.n2370 GNDA.n2369 150
R9804 GNDA.n2374 GNDA.n2373 150
R9805 GNDA.n3080 GNDA.n670 150
R9806 GNDA.n3070 GNDA.n3069 150
R9807 GNDA.n3083 GNDA.n651 150
R9808 GNDA.n2311 GNDA.n652 150
R9809 GNDA.n2338 GNDA.n2337 150
R9810 GNDA.n2334 GNDA.n2333 150
R9811 GNDA.n2330 GNDA.n2329 150
R9812 GNDA.n2326 GNDA.n669 150
R9813 GNDA.n5026 GNDA.n5025 150
R9814 GNDA.n5022 GNDA.n5021 150
R9815 GNDA.n5018 GNDA.n5017 150
R9816 GNDA.n5014 GNDA.n5013 150
R9817 GNDA.n5010 GNDA.n5009 150
R9818 GNDA.n5006 GNDA.n5005 150
R9819 GNDA.n5002 GNDA.n5001 150
R9820 GNDA.n4998 GNDA.n4997 150
R9821 GNDA.n5049 GNDA.n168 150
R9822 GNDA.n216 GNDA.n169 150
R9823 GNDA.n213 GNDA.n212 150
R9824 GNDA.n205 GNDA.n204 150
R9825 GNDA.n5034 GNDA.n5033 150
R9826 GNDA.n5038 GNDA.n5037 150
R9827 GNDA.n5042 GNDA.n5041 150
R9828 GNDA.n5046 GNDA.n5045 150
R9829 GNDA.n4811 GNDA.n4810 150
R9830 GNDA.n4807 GNDA.n4806 150
R9831 GNDA.n4803 GNDA.n4802 150
R9832 GNDA.n4799 GNDA.n4798 150
R9833 GNDA.n4795 GNDA.n4794 150
R9834 GNDA.n4791 GNDA.n4790 150
R9835 GNDA.n4787 GNDA.n4786 150
R9836 GNDA.n4783 GNDA.n4782 150
R9837 GNDA.n4834 GNDA.n4730 150
R9838 GNDA.n4756 GNDA.n4731 150
R9839 GNDA.n4764 GNDA.n4763 150
R9840 GNDA.n4771 GNDA.n4770 150
R9841 GNDA.n4819 GNDA.n4818 150
R9842 GNDA.n4823 GNDA.n4822 150
R9843 GNDA.n4827 GNDA.n4826 150
R9844 GNDA.n4831 GNDA.n4830 150
R9845 GNDA.n2679 GNDA.n2678 150
R9846 GNDA.n2675 GNDA.n2674 150
R9847 GNDA.n2671 GNDA.n2670 150
R9848 GNDA.n2667 GNDA.n2666 150
R9849 GNDA.n2663 GNDA.n2662 150
R9850 GNDA.n2659 GNDA.n2658 150
R9851 GNDA.n2655 GNDA.n2654 150
R9852 GNDA.n2651 GNDA.n2650 150
R9853 GNDA.n2728 GNDA.n2648 150
R9854 GNDA.n2717 GNDA.n2716 150
R9855 GNDA.n2710 GNDA.n2709 150
R9856 GNDA.n2731 GNDA.n2628 150
R9857 GNDA.n2687 GNDA.n2686 150
R9858 GNDA.n2691 GNDA.n2690 150
R9859 GNDA.n2695 GNDA.n2694 150
R9860 GNDA.n2697 GNDA.n2647 150
R9861 GNDA.n4952 GNDA.n4951 150
R9862 GNDA.n4948 GNDA.n4947 150
R9863 GNDA.n4944 GNDA.n4943 150
R9864 GNDA.n4940 GNDA.n4939 150
R9865 GNDA.n4936 GNDA.n4935 150
R9866 GNDA.n4932 GNDA.n4931 150
R9867 GNDA.n4928 GNDA.n4927 150
R9868 GNDA.n4924 GNDA.n4923 150
R9869 GNDA.n4981 GNDA.n4980 150
R9870 GNDA.n4973 GNDA.n4878 150
R9871 GNDA.n4905 GNDA.n4879 150
R9872 GNDA.n4912 GNDA.n4911 150
R9873 GNDA.n4970 GNDA.n4895 150
R9874 GNDA.n4966 GNDA.n4965 150
R9875 GNDA.n4962 GNDA.n4961 150
R9876 GNDA.n4958 GNDA.n4957 150
R9877 GNDA.n5231 GNDA.n5230 150
R9878 GNDA.n5227 GNDA.n5226 150
R9879 GNDA.n5223 GNDA.n5222 150
R9880 GNDA.n5219 GNDA.n5218 150
R9881 GNDA.n5215 GNDA.n5214 150
R9882 GNDA.n5211 GNDA.n5210 150
R9883 GNDA.n5207 GNDA.n5206 150
R9884 GNDA.n5203 GNDA.n5202 150
R9885 GNDA.n5260 GNDA.n5259 150
R9886 GNDA.n5252 GNDA.n64 150
R9887 GNDA.n5184 GNDA.n65 150
R9888 GNDA.n5191 GNDA.n5190 150
R9889 GNDA.n5249 GNDA.n81 150
R9890 GNDA.n5245 GNDA.n5244 150
R9891 GNDA.n5241 GNDA.n5240 150
R9892 GNDA.n5237 GNDA.n5236 150
R9893 GNDA.n2467 GNDA.n2465 150
R9894 GNDA.n2463 GNDA.n2260 150
R9895 GNDA.n2459 GNDA.n2457 150
R9896 GNDA.n2455 GNDA.n2262 150
R9897 GNDA.n2451 GNDA.n2449 150
R9898 GNDA.n2447 GNDA.n2264 150
R9899 GNDA.n2443 GNDA.n2442 150
R9900 GNDA.n2440 GNDA.n2267 150
R9901 GNDA.n2493 GNDA.n2492 150
R9902 GNDA.n2495 GNDA.n2253 150
R9903 GNDA.n2420 GNDA.n2418 150
R9904 GNDA.n2433 GNDA.n2271 150
R9905 GNDA.n2475 GNDA.n2473 150
R9906 GNDA.n2479 GNDA.n2256 150
R9907 GNDA.n2483 GNDA.n2481 150
R9908 GNDA.n2487 GNDA.n2254 150
R9909 GNDA.n5149 GNDA.n5148 150
R9910 GNDA.n5145 GNDA.n5144 150
R9911 GNDA.n5141 GNDA.n5140 150
R9912 GNDA.n5137 GNDA.n5136 150
R9913 GNDA.n5133 GNDA.n5132 150
R9914 GNDA.n5129 GNDA.n5128 150
R9915 GNDA.n5125 GNDA.n5124 150
R9916 GNDA.n5121 GNDA.n5120 150
R9917 GNDA.n5272 GNDA.n21 150
R9918 GNDA.n37 GNDA.n36 150
R9919 GNDA.n5275 GNDA.n2 150
R9920 GNDA.n5109 GNDA.n3 150
R9921 GNDA.n5157 GNDA.n5156 150
R9922 GNDA.n5161 GNDA.n5160 150
R9923 GNDA.n5165 GNDA.n5164 150
R9924 GNDA.n5167 GNDA.n20 150
R9925 GNDA.n4623 GNDA.n4622 148.017
R9926 GNDA.n4629 GNDA.n4628 148.017
R9927 GNDA.n3152 GNDA.n3151 148.017
R9928 GNDA.n1746 GNDA.n1745 148.017
R9929 GNDA.n3051 GNDA.n684 136.145
R9930 GNDA.n3052 GNDA.n683 136.145
R9931 GNDA.n3053 GNDA.n682 136.145
R9932 GNDA.n3056 GNDA.n679 136.145
R9933 GNDA.n3057 GNDA.n678 136.145
R9934 GNDA.n3058 GNDA.n677 136.145
R9935 GNDA.n2506 GNDA.n2505 136.145
R9936 GNDA.n2507 GNDA.n2504 136.145
R9937 GNDA.n2508 GNDA.n2503 136.145
R9938 GNDA.n2247 GNDA.n2246 136.145
R9939 GNDA.n2245 GNDA.n2244 136.145
R9940 GNDA.n2406 GNDA.n2399 134.268
R9941 GNDA.n2399 GNDA.n2397 134.268
R9942 GNDA.n835 GNDA.n281 132.721
R9943 GNDA.n4622 GNDA.t24 130.847
R9944 GNDA.n3049 GNDA.t108 130.001
R9945 GNDA.n2975 GNDA.t53 130.001
R9946 GNDA.n807 GNDA.t119 130.001
R9947 GNDA.n3061 GNDA.t71 130.001
R9948 GNDA.n2319 GNDA.t50 130.001
R9949 GNDA.n2501 GNDA.t140 130.001
R9950 GNDA.n2512 GNDA.t95 130.001
R9951 GNDA.n2241 GNDA.t43 130
R9952 GNDA.n5088 GNDA.t45 127.219
R9953 GNDA.t45 GNDA.n108 127.219
R9954 GNDA.t45 GNDA.n710 127.219
R9955 GNDA.n2982 GNDA.n2981 124.832
R9956 GNDA.n2979 GNDA.n2978 124.832
R9957 GNDA.n2317 GNDA.n815 124.832
R9958 GNDA.n2973 GNDA.n2972 124.832
R9959 GNDA.n5175 GNDA.n83 124.832
R9960 GNDA.n327 GNDA.n55 124.832
R9961 GNDA.n2822 GNDA.n2821 124.832
R9962 GNDA.n2819 GNDA.n2575 124.832
R9963 GNDA.n5059 GNDA.n5058 124.832
R9964 GNDA.n4896 GNDA.n159 124.832
R9965 GNDA.n325 GNDA.n85 124.832
R9966 GNDA.n5173 GNDA.n86 124.832
R9967 GNDA.n1306 GNDA.n1305 121.136
R9968 GNDA.n1308 GNDA.n1307 121.136
R9969 GNDA.n1310 GNDA.n1309 121.136
R9970 GNDA.n1312 GNDA.n1311 121.136
R9971 GNDA.n1314 GNDA.n1313 121.136
R9972 GNDA.n1316 GNDA.n1315 121.136
R9973 GNDA.n1366 GNDA.n1365 121.136
R9974 GNDA.n1368 GNDA.n1367 121.136
R9975 GNDA.n1370 GNDA.n1369 121.136
R9976 GNDA.n1372 GNDA.n1371 121.136
R9977 GNDA.n1374 GNDA.n1373 121.136
R9978 GNDA.n1376 GNDA.n1375 121.136
R9979 GNDA.n2210 GNDA.t168 111.799
R9980 GNDA.n2209 GNDA.t165 111.331
R9981 GNDA.n2227 GNDA.t283 111.206
R9982 GNDA.n2227 GNDA.t264 111.076
R9983 GNDA.n4705 GNDA.n300 105.719
R9984 GNDA.n4673 GNDA.n4672 105.719
R9985 GNDA.n4699 GNDA.n300 103.457
R9986 GNDA.n4672 GNDA.n4671 103.457
R9987 GNDA.n3011 GNDA.n708 101.718
R9988 GNDA.n2402 GNDA.n2276 101.718
R9989 GNDA.n2408 GNDA.n2278 101.718
R9990 GNDA.n3022 GNDA.n706 101.718
R9991 GNDA.t45 GNDA.n104 47.6748
R9992 GNDA.n3018 GNDA.n705 91.069
R9993 GNDA.n3013 GNDA.n705 91.069
R9994 GNDA.n3015 GNDA.n704 91.069
R9995 GNDA.n3016 GNDA.n3015 91.069
R9996 GNDA.n2406 GNDA.n2401 91.069
R9997 GNDA.n2404 GNDA.n2397 91.069
R9998 GNDA.n2515 GNDA.n2514 90.1439
R9999 GNDA.n2426 GNDA.n2425 90.1439
R10000 GNDA.n3076 GNDA.n3063 90.1439
R10001 GNDA.n2998 GNDA.n2997 90.1439
R10002 GNDA.n723 GNDA.n685 90.1439
R10003 GNDA.n3047 GNDA.n686 90.1439
R10004 GNDA.n2500 GNDA.n838 87.1391
R10005 GNDA.t45 GNDA.n809 87.1391
R10006 GNDA.n2292 GNDA.n2291 84.306
R10007 GNDA.n2386 GNDA.n2303 84.306
R10008 GNDA.n2249 GNDA.t13 83.1328
R10009 GNDA.n2410 GNDA.t21 82.1312
R10010 GNDA.n3074 GNDA.t217 82.1312
R10011 GNDA.n2999 GNDA.t228 82.1312
R10012 GNDA.n696 GNDA.t239 78.5658
R10013 GNDA.n2429 GNDA.t143 78.1248
R10014 GNDA.n2306 GNDA.t145 78.1248
R10015 GNDA.t261 GNDA.n707 78.1248
R10016 GNDA.t45 GNDA.n100 76.3879
R10017 GNDA.n2915 GNDA.n2914 76.3222
R10018 GNDA.n2858 GNDA.n2829 76.3222
R10019 GNDA.n2854 GNDA.n2853 76.3222
R10020 GNDA.n2847 GNDA.n2834 76.3222
R10021 GNDA.n2846 GNDA.n2845 76.3222
R10022 GNDA.n2912 GNDA.n2911 76.3222
R10023 GNDA.n2907 GNDA.n2863 76.3222
R10024 GNDA.n2905 GNDA.n2904 76.3222
R10025 GNDA.n2900 GNDA.n2866 76.3222
R10026 GNDA.n2898 GNDA.n2897 76.3222
R10027 GNDA.n2893 GNDA.n2869 76.3222
R10028 GNDA.n2919 GNDA.n2918 76.3222
R10029 GNDA.n2831 GNDA.n2830 76.3222
R10030 GNDA.n2836 GNDA.n2835 76.3222
R10031 GNDA.n2839 GNDA.n2838 76.3222
R10032 GNDA.n2843 GNDA.n2841 76.3222
R10033 GNDA.n2979 GNDA.n805 76.3222
R10034 GNDA.n2940 GNDA.n2939 76.3222
R10035 GNDA.n2935 GNDA.n2568 76.3222
R10036 GNDA.n2933 GNDA.n2932 76.3222
R10037 GNDA.n2928 GNDA.n2571 76.3222
R10038 GNDA.n2926 GNDA.n2925 76.3222
R10039 GNDA.n2921 GNDA.n2825 76.3222
R10040 GNDA.n2943 GNDA.n2942 76.3222
R10041 GNDA.n2953 GNDA.n2952 76.3222
R10042 GNDA.n825 GNDA.n824 76.3222
R10043 GNDA.n2964 GNDA.n2963 76.3222
R10044 GNDA.n2967 GNDA.n2966 76.3222
R10045 GNDA.n834 GNDA.n286 76.3222
R10046 GNDA.n2536 GNDA.n285 76.3222
R10047 GNDA.n2532 GNDA.n284 76.3222
R10048 GNDA.n2528 GNDA.n283 76.3222
R10049 GNDA.n2524 GNDA.n282 76.3222
R10050 GNDA.n2520 GNDA.n281 76.3222
R10051 GNDA.n2543 GNDA.n2542 76.3222
R10052 GNDA.n2544 GNDA.n832 76.3222
R10053 GNDA.n2551 GNDA.n2550 76.3222
R10054 GNDA.n2552 GNDA.n830 76.3222
R10055 GNDA.n2559 GNDA.n2558 76.3222
R10056 GNDA.n2560 GNDA.n828 76.3222
R10057 GNDA.n2946 GNDA.n2945 76.3222
R10058 GNDA.n2949 GNDA.n2948 76.3222
R10059 GNDA.n2957 GNDA.n2956 76.3222
R10060 GNDA.n2960 GNDA.n2959 76.3222
R10061 GNDA.n820 GNDA.n819 76.3222
R10062 GNDA.n2971 GNDA.n2970 76.3222
R10063 GNDA.n370 GNDA.n369 76.3222
R10064 GNDA.n375 GNDA.n374 76.3222
R10065 GNDA.n378 GNDA.n377 76.3222
R10066 GNDA.n383 GNDA.n382 76.3222
R10067 GNDA.n386 GNDA.n385 76.3222
R10068 GNDA.n387 GNDA.n83 76.3222
R10069 GNDA.n349 GNDA.n348 76.3222
R10070 GNDA.n342 GNDA.n304 76.3222
R10071 GNDA.n341 GNDA.n340 76.3222
R10072 GNDA.n334 GNDA.n311 76.3222
R10073 GNDA.n333 GNDA.n332 76.3222
R10074 GNDA.n326 GNDA.n319 76.3222
R10075 GNDA.n2576 GNDA.n195 76.3222
R10076 GNDA.n2725 GNDA.n194 76.3222
R10077 GNDA.n2720 GNDA.n193 76.3222
R10078 GNDA.n2713 GNDA.n192 76.3222
R10079 GNDA.n2706 GNDA.n191 76.3222
R10080 GNDA.n2735 GNDA.n190 76.3222
R10081 GNDA.n2789 GNDA.n2788 76.3222
R10082 GNDA.n2799 GNDA.n2798 76.3222
R10083 GNDA.n2802 GNDA.n2801 76.3222
R10084 GNDA.n2811 GNDA.n2810 76.3222
R10085 GNDA.n2814 GNDA.n2813 76.3222
R10086 GNDA.n2784 GNDA.n112 76.3222
R10087 GNDA.n2780 GNDA.n113 76.3222
R10088 GNDA.n2776 GNDA.n114 76.3222
R10089 GNDA.n2772 GNDA.n115 76.3222
R10090 GNDA.n2768 GNDA.n116 76.3222
R10091 GNDA.n2764 GNDA.n117 76.3222
R10092 GNDA.n2792 GNDA.n2587 76.3222
R10093 GNDA.n2796 GNDA.n2794 76.3222
R10094 GNDA.n2804 GNDA.n2583 76.3222
R10095 GNDA.n2808 GNDA.n2806 76.3222
R10096 GNDA.n2816 GNDA.n2579 76.3222
R10097 GNDA.n2819 GNDA.n2818 76.3222
R10098 GNDA.n5057 GNDA.n163 76.3222
R10099 GNDA.n5052 GNDA.n166 76.3222
R10100 GNDA.n220 GNDA.n219 76.3222
R10101 GNDA.n201 GNDA.n197 76.3222
R10102 GNDA.n208 GNDA.n196 76.3222
R10103 GNDA.n4990 GNDA.n4989 76.3222
R10104 GNDA.n5081 GNDA.n5080 76.3222
R10105 GNDA.n5078 GNDA.n5077 76.3222
R10106 GNDA.n5073 GNDA.n140 76.3222
R10107 GNDA.n5070 GNDA.n139 76.3222
R10108 GNDA.n5066 GNDA.n138 76.3222
R10109 GNDA.n5062 GNDA.n137 76.3222
R10110 GNDA.n2590 GNDA.n118 76.3222
R10111 GNDA.n2594 GNDA.n119 76.3222
R10112 GNDA.n2598 GNDA.n120 76.3222
R10113 GNDA.n2602 GNDA.n121 76.3222
R10114 GNDA.n2606 GNDA.n122 76.3222
R10115 GNDA.n2610 GNDA.n123 76.3222
R10116 GNDA.n152 GNDA.n151 76.3222
R10117 GNDA.n153 GNDA.n143 76.3222
R10118 GNDA.n154 GNDA.n145 76.3222
R10119 GNDA.n155 GNDA.n147 76.3222
R10120 GNDA.n156 GNDA.n149 76.3222
R10121 GNDA.n159 GNDA.n158 76.3222
R10122 GNDA.n4987 GNDA.n4986 76.3222
R10123 GNDA.n4872 GNDA.n225 76.3222
R10124 GNDA.n4976 GNDA.n224 76.3222
R10125 GNDA.n4903 GNDA.n223 76.3222
R10126 GNDA.n4907 GNDA.n222 76.3222
R10127 GNDA.n4916 GNDA.n221 76.3222
R10128 GNDA.n261 GNDA.n235 76.3222
R10129 GNDA.n265 GNDA.n236 76.3222
R10130 GNDA.n269 GNDA.n237 76.3222
R10131 GNDA.n273 GNDA.n238 76.3222
R10132 GNDA.n279 GNDA.n278 76.3222
R10133 GNDA.n257 GNDA.n124 76.3222
R10134 GNDA.n253 GNDA.n125 76.3222
R10135 GNDA.n249 GNDA.n126 76.3222
R10136 GNDA.n245 GNDA.n127 76.3222
R10137 GNDA.n241 GNDA.n128 76.3222
R10138 GNDA.n5086 GNDA.n5085 76.3222
R10139 GNDA.n306 GNDA.n305 76.3222
R10140 GNDA.n309 GNDA.n308 76.3222
R10141 GNDA.n314 GNDA.n313 76.3222
R10142 GNDA.n317 GNDA.n316 76.3222
R10143 GNDA.n322 GNDA.n321 76.3222
R10144 GNDA.n325 GNDA.n324 76.3222
R10145 GNDA.n4838 GNDA.n48 76.3222
R10146 GNDA.n4753 GNDA.n47 76.3222
R10147 GNDA.n4759 GNDA.n46 76.3222
R10148 GNDA.n4767 GNDA.n45 76.3222
R10149 GNDA.n4774 GNDA.n44 76.3222
R10150 GNDA.n4748 GNDA.n43 76.3222
R10151 GNDA.n4866 GNDA.n4865 76.3222
R10152 GNDA.n4860 GNDA.n230 76.3222
R10153 GNDA.n4857 GNDA.n231 76.3222
R10154 GNDA.n4853 GNDA.n232 76.3222
R10155 GNDA.n4849 GNDA.n233 76.3222
R10156 GNDA.n5086 GNDA.n129 76.3222
R10157 GNDA.n244 GNDA.n128 76.3222
R10158 GNDA.n248 GNDA.n127 76.3222
R10159 GNDA.n252 GNDA.n126 76.3222
R10160 GNDA.n256 GNDA.n125 76.3222
R10161 GNDA.n260 GNDA.n124 76.3222
R10162 GNDA.n2607 GNDA.n123 76.3222
R10163 GNDA.n2603 GNDA.n122 76.3222
R10164 GNDA.n2599 GNDA.n121 76.3222
R10165 GNDA.n2595 GNDA.n120 76.3222
R10166 GNDA.n2591 GNDA.n119 76.3222
R10167 GNDA.n135 GNDA.n118 76.3222
R10168 GNDA.n2767 GNDA.n117 76.3222
R10169 GNDA.n2771 GNDA.n116 76.3222
R10170 GNDA.n2775 GNDA.n115 76.3222
R10171 GNDA.n2779 GNDA.n114 76.3222
R10172 GNDA.n2783 GNDA.n113 76.3222
R10173 GNDA.n2787 GNDA.n112 76.3222
R10174 GNDA.n5266 GNDA.n54 76.3222
R10175 GNDA.n5256 GNDA.n53 76.3222
R10176 GNDA.n5181 GNDA.n52 76.3222
R10177 GNDA.n5187 GNDA.n51 76.3222
R10178 GNDA.n5194 GNDA.n50 76.3222
R10179 GNDA.n5176 GNDA.n49 76.3222
R10180 GNDA.n5266 GNDA.n5265 76.3222
R10181 GNDA.n58 GNDA.n53 76.3222
R10182 GNDA.n5255 GNDA.n52 76.3222
R10183 GNDA.n5182 GNDA.n51 76.3222
R10184 GNDA.n5186 GNDA.n50 76.3222
R10185 GNDA.n5195 GNDA.n49 76.3222
R10186 GNDA.n4842 GNDA.n48 76.3222
R10187 GNDA.n4837 GNDA.n47 76.3222
R10188 GNDA.n4754 GNDA.n46 76.3222
R10189 GNDA.n4760 GNDA.n45 76.3222
R10190 GNDA.n4766 GNDA.n44 76.3222
R10191 GNDA.n4775 GNDA.n43 76.3222
R10192 GNDA.n324 GNDA.n323 76.3222
R10193 GNDA.n321 GNDA.n320 76.3222
R10194 GNDA.n316 GNDA.n315 76.3222
R10195 GNDA.n313 GNDA.n312 76.3222
R10196 GNDA.n308 GNDA.n307 76.3222
R10197 GNDA.n305 GNDA.n301 76.3222
R10198 GNDA.n348 GNDA.n347 76.3222
R10199 GNDA.n343 GNDA.n342 76.3222
R10200 GNDA.n340 GNDA.n339 76.3222
R10201 GNDA.n335 GNDA.n334 76.3222
R10202 GNDA.n332 GNDA.n331 76.3222
R10203 GNDA.n327 GNDA.n326 76.3222
R10204 GNDA.n158 GNDA.n150 76.3222
R10205 GNDA.n156 GNDA.n148 76.3222
R10206 GNDA.n155 GNDA.n146 76.3222
R10207 GNDA.n154 GNDA.n144 76.3222
R10208 GNDA.n153 GNDA.n142 76.3222
R10209 GNDA.n152 GNDA.n130 76.3222
R10210 GNDA.n5080 GNDA.n136 76.3222
R10211 GNDA.n5078 GNDA.n141 76.3222
R10212 GNDA.n5071 GNDA.n140 76.3222
R10213 GNDA.n5067 GNDA.n139 76.3222
R10214 GNDA.n5063 GNDA.n138 76.3222
R10215 GNDA.n5059 GNDA.n137 76.3222
R10216 GNDA.n2972 GNDA.n2971 76.3222
R10217 GNDA.n819 GNDA.n813 76.3222
R10218 GNDA.n2961 GNDA.n2960 76.3222
R10219 GNDA.n2958 GNDA.n2957 76.3222
R10220 GNDA.n2948 GNDA.n822 76.3222
R10221 GNDA.n2947 GNDA.n2946 76.3222
R10222 GNDA.n2942 GNDA.n826 76.3222
R10223 GNDA.n2954 GNDA.n2953 76.3222
R10224 GNDA.n824 GNDA.n817 76.3222
R10225 GNDA.n2965 GNDA.n2964 76.3222
R10226 GNDA.n2968 GNDA.n2967 76.3222
R10227 GNDA.n2561 GNDA.n2560 76.3222
R10228 GNDA.n2558 GNDA.n2557 76.3222
R10229 GNDA.n2553 GNDA.n2552 76.3222
R10230 GNDA.n2550 GNDA.n2549 76.3222
R10231 GNDA.n2545 GNDA.n2544 76.3222
R10232 GNDA.n2542 GNDA.n2541 76.3222
R10233 GNDA.n2825 GNDA.n2572 76.3222
R10234 GNDA.n2927 GNDA.n2926 76.3222
R10235 GNDA.n2571 GNDA.n2569 76.3222
R10236 GNDA.n2934 GNDA.n2933 76.3222
R10237 GNDA.n2568 GNDA.n2566 76.3222
R10238 GNDA.n2941 GNDA.n2940 76.3222
R10239 GNDA.n2869 GNDA.n2867 76.3222
R10240 GNDA.n2899 GNDA.n2898 76.3222
R10241 GNDA.n2866 GNDA.n2864 76.3222
R10242 GNDA.n2906 GNDA.n2905 76.3222
R10243 GNDA.n2863 GNDA.n2861 76.3222
R10244 GNDA.n2913 GNDA.n2912 76.3222
R10245 GNDA.n4987 GNDA.n226 76.3222
R10246 GNDA.n4977 GNDA.n225 76.3222
R10247 GNDA.n4902 GNDA.n224 76.3222
R10248 GNDA.n4908 GNDA.n223 76.3222
R10249 GNDA.n4915 GNDA.n222 76.3222
R10250 GNDA.n4897 GNDA.n221 76.3222
R10251 GNDA.n5053 GNDA.n163 76.3222
R10252 GNDA.n199 GNDA.n166 76.3222
R10253 GNDA.n220 GNDA.n198 76.3222
R10254 GNDA.n209 GNDA.n197 76.3222
R10255 GNDA.n196 GNDA.n188 76.3222
R10256 GNDA.n4989 GNDA.n189 76.3222
R10257 GNDA.n2724 GNDA.n195 76.3222
R10258 GNDA.n2721 GNDA.n194 76.3222
R10259 GNDA.n2714 GNDA.n193 76.3222
R10260 GNDA.n2707 GNDA.n192 76.3222
R10261 GNDA.n2734 GNDA.n191 76.3222
R10262 GNDA.n2739 GNDA.n190 76.3222
R10263 GNDA.n412 GNDA.n368 76.3222
R10264 GNDA.n408 GNDA.n407 76.3222
R10265 GNDA.n401 GNDA.n372 76.3222
R10266 GNDA.n400 GNDA.n399 76.3222
R10267 GNDA.n393 GNDA.n380 76.3222
R10268 GNDA.n392 GNDA.n391 76.3222
R10269 GNDA.n42 GNDA.n24 76.3222
R10270 GNDA.n5268 GNDA.n25 76.3222
R10271 GNDA.n41 GNDA.n31 76.3222
R10272 GNDA.n5106 GNDA.n29 76.3222
R10273 GNDA.n5112 GNDA.n28 76.3222
R10274 GNDA.n5102 GNDA.n27 76.3222
R10275 GNDA.n5172 GNDA.n42 76.3222
R10276 GNDA.n5269 GNDA.n5268 76.3222
R10277 GNDA.n41 GNDA.n40 76.3222
R10278 GNDA.n30 GNDA.n29 76.3222
R10279 GNDA.n5107 GNDA.n28 76.3222
R10280 GNDA.n5113 GNDA.n27 76.3222
R10281 GNDA.n388 GNDA.n387 76.3222
R10282 GNDA.n385 GNDA.n384 76.3222
R10283 GNDA.n382 GNDA.n381 76.3222
R10284 GNDA.n377 GNDA.n376 76.3222
R10285 GNDA.n374 GNDA.n373 76.3222
R10286 GNDA.n369 GNDA.n366 76.3222
R10287 GNDA.n409 GNDA.n368 76.3222
R10288 GNDA.n407 GNDA.n406 76.3222
R10289 GNDA.n402 GNDA.n401 76.3222
R10290 GNDA.n399 GNDA.n398 76.3222
R10291 GNDA.n394 GNDA.n393 76.3222
R10292 GNDA.n391 GNDA.n86 76.3222
R10293 GNDA.n2818 GNDA.n2817 76.3222
R10294 GNDA.n2807 GNDA.n2579 76.3222
R10295 GNDA.n2806 GNDA.n2805 76.3222
R10296 GNDA.n2795 GNDA.n2583 76.3222
R10297 GNDA.n2794 GNDA.n2793 76.3222
R10298 GNDA.n2609 GNDA.n2587 76.3222
R10299 GNDA.n2790 GNDA.n2789 76.3222
R10300 GNDA.n2800 GNDA.n2799 76.3222
R10301 GNDA.n2801 GNDA.n2581 76.3222
R10302 GNDA.n2812 GNDA.n2811 76.3222
R10303 GNDA.n2813 GNDA.n2577 76.3222
R10304 GNDA.n2842 GNDA.n805 76.3222
R10305 GNDA.n2841 GNDA.n2840 76.3222
R10306 GNDA.n2838 GNDA.n2837 76.3222
R10307 GNDA.n2835 GNDA.n2832 76.3222
R10308 GNDA.n2830 GNDA.n2827 76.3222
R10309 GNDA.n2920 GNDA.n2919 76.3222
R10310 GNDA.n2916 GNDA.n2915 76.3222
R10311 GNDA.n2855 GNDA.n2829 76.3222
R10312 GNDA.n2853 GNDA.n2852 76.3222
R10313 GNDA.n2848 GNDA.n2847 76.3222
R10314 GNDA.n2845 GNDA.n749 76.3222
R10315 GNDA.n2537 GNDA.n286 76.3222
R10316 GNDA.n2533 GNDA.n285 76.3222
R10317 GNDA.n2529 GNDA.n284 76.3222
R10318 GNDA.n2525 GNDA.n283 76.3222
R10319 GNDA.n2521 GNDA.n282 76.3222
R10320 GNDA.n264 GNDA.n235 76.3222
R10321 GNDA.n268 GNDA.n236 76.3222
R10322 GNDA.n272 GNDA.n237 76.3222
R10323 GNDA.n240 GNDA.n238 76.3222
R10324 GNDA.n279 GNDA.n239 76.3222
R10325 GNDA.n4866 GNDA.n288 76.3222
R10326 GNDA.n4858 GNDA.n230 76.3222
R10327 GNDA.n4854 GNDA.n231 76.3222
R10328 GNDA.n4850 GNDA.n232 76.3222
R10329 GNDA.n4846 GNDA.n233 76.3222
R10330 GNDA.n768 GNDA.n730 74.5978
R10331 GNDA.n765 GNDA.n730 74.5978
R10332 GNDA.n2358 GNDA.n658 74.5978
R10333 GNDA.n2361 GNDA.n658 74.5978
R10334 GNDA.n5013 GNDA.n175 74.5978
R10335 GNDA.n5010 GNDA.n175 74.5978
R10336 GNDA.n4798 GNDA.n4737 74.5978
R10337 GNDA.n4795 GNDA.n4737 74.5978
R10338 GNDA.n2666 GNDA.n2635 74.5978
R10339 GNDA.n2663 GNDA.n2635 74.5978
R10340 GNDA.n4939 GNDA.n4884 74.5978
R10341 GNDA.n4936 GNDA.n4884 74.5978
R10342 GNDA.n5218 GNDA.n70 74.5978
R10343 GNDA.n5215 GNDA.n70 74.5978
R10344 GNDA.n2450 GNDA.n2262 74.5978
R10345 GNDA.n2451 GNDA.n2450 74.5978
R10346 GNDA.n5136 GNDA.n9 74.5978
R10347 GNDA.n5133 GNDA.n9 74.5978
R10348 GNDA.n2977 GNDA.n808 74.1184
R10349 GNDA.n2427 GNDA.t290 72.1152
R10350 GNDA.n2307 GNDA.t117 72.1152
R10351 GNDA.t107 GNDA.n722 72.1152
R10352 GNDA.t45 GNDA.t152 70.1899
R10353 GNDA.n4689 GNDA.n4688 69.4466
R10354 GNDA.n3004 GNDA.n3003 69.3109
R10355 GNDA.n3004 GNDA.n743 69.3109
R10356 GNDA.n3081 GNDA.n3080 69.3109
R10357 GNDA.n3081 GNDA.n669 69.3109
R10358 GNDA.n5047 GNDA.n168 69.3109
R10359 GNDA.n5047 GNDA.n5046 69.3109
R10360 GNDA.n4832 GNDA.n4730 69.3109
R10361 GNDA.n4832 GNDA.n4831 69.3109
R10362 GNDA.n2729 GNDA.n2728 69.3109
R10363 GNDA.n2729 GNDA.n2647 69.3109
R10364 GNDA.n4981 GNDA.n4874 69.3109
R10365 GNDA.n4957 GNDA.n4874 69.3109
R10366 GNDA.n5260 GNDA.n60 69.3109
R10367 GNDA.n5236 GNDA.n60 69.3109
R10368 GNDA.n2492 GNDA.n2488 69.3109
R10369 GNDA.n2488 GNDA.n2487 69.3109
R10370 GNDA.n5273 GNDA.n5272 69.3109
R10371 GNDA.n5273 GNDA.n20 69.3109
R10372 GNDA.n2984 GNDA.t52 68.1089
R10373 GNDA.n2977 GNDA.n2976 66.1057
R10374 GNDA.t128 GNDA.n742 65.8183
R10375 GNDA.t128 GNDA.n741 65.8183
R10376 GNDA.t128 GNDA.n740 65.8183
R10377 GNDA.t128 GNDA.n739 65.8183
R10378 GNDA.t128 GNDA.n720 65.8183
R10379 GNDA.t128 GNDA.n737 65.8183
R10380 GNDA.t128 GNDA.n718 65.8183
R10381 GNDA.t128 GNDA.n738 65.8183
R10382 GNDA.t128 GNDA.n736 65.8183
R10383 GNDA.t128 GNDA.n733 65.8183
R10384 GNDA.t128 GNDA.n732 65.8183
R10385 GNDA.t128 GNDA.n731 65.8183
R10386 GNDA.t128 GNDA.n729 65.8183
R10387 GNDA.n3005 GNDA.t128 65.8183
R10388 GNDA.t128 GNDA.n719 65.8183
R10389 GNDA.t128 GNDA.n717 65.8183
R10390 GNDA.t72 GNDA.n668 65.8183
R10391 GNDA.t72 GNDA.n667 65.8183
R10392 GNDA.t72 GNDA.n666 65.8183
R10393 GNDA.t72 GNDA.n665 65.8183
R10394 GNDA.t72 GNDA.n656 65.8183
R10395 GNDA.t72 GNDA.n663 65.8183
R10396 GNDA.t72 GNDA.n654 65.8183
R10397 GNDA.t72 GNDA.n664 65.8183
R10398 GNDA.t72 GNDA.n662 65.8183
R10399 GNDA.t72 GNDA.n661 65.8183
R10400 GNDA.t72 GNDA.n660 65.8183
R10401 GNDA.t72 GNDA.n659 65.8183
R10402 GNDA.t72 GNDA.n657 65.8183
R10403 GNDA.n3082 GNDA.t72 65.8183
R10404 GNDA.t72 GNDA.n655 65.8183
R10405 GNDA.t72 GNDA.n653 65.8183
R10406 GNDA.t59 GNDA.n185 65.8183
R10407 GNDA.t59 GNDA.n184 65.8183
R10408 GNDA.t59 GNDA.n183 65.8183
R10409 GNDA.t59 GNDA.n182 65.8183
R10410 GNDA.t59 GNDA.n173 65.8183
R10411 GNDA.t59 GNDA.n180 65.8183
R10412 GNDA.t59 GNDA.n170 65.8183
R10413 GNDA.t59 GNDA.n181 65.8183
R10414 GNDA.t59 GNDA.n179 65.8183
R10415 GNDA.t59 GNDA.n178 65.8183
R10416 GNDA.t59 GNDA.n177 65.8183
R10417 GNDA.t59 GNDA.n176 65.8183
R10418 GNDA.t59 GNDA.n174 65.8183
R10419 GNDA.t59 GNDA.n172 65.8183
R10420 GNDA.t59 GNDA.n171 65.8183
R10421 GNDA.n5048 GNDA.t59 65.8183
R10422 GNDA.t44 GNDA.n4747 65.8183
R10423 GNDA.t44 GNDA.n4746 65.8183
R10424 GNDA.t44 GNDA.n4745 65.8183
R10425 GNDA.t44 GNDA.n4744 65.8183
R10426 GNDA.t44 GNDA.n4735 65.8183
R10427 GNDA.t44 GNDA.n4742 65.8183
R10428 GNDA.t44 GNDA.n4732 65.8183
R10429 GNDA.t44 GNDA.n4743 65.8183
R10430 GNDA.t44 GNDA.n4741 65.8183
R10431 GNDA.t44 GNDA.n4740 65.8183
R10432 GNDA.t44 GNDA.n4739 65.8183
R10433 GNDA.t44 GNDA.n4738 65.8183
R10434 GNDA.t84 GNDA.n2646 65.8183
R10435 GNDA.t84 GNDA.n2645 65.8183
R10436 GNDA.t84 GNDA.n2644 65.8183
R10437 GNDA.t84 GNDA.n2643 65.8183
R10438 GNDA.t84 GNDA.n2634 65.8183
R10439 GNDA.t84 GNDA.n2641 65.8183
R10440 GNDA.t84 GNDA.n2631 65.8183
R10441 GNDA.t84 GNDA.n2642 65.8183
R10442 GNDA.t84 GNDA.n2640 65.8183
R10443 GNDA.t84 GNDA.n2638 65.8183
R10444 GNDA.t84 GNDA.n2637 65.8183
R10445 GNDA.t84 GNDA.n2636 65.8183
R10446 GNDA.n2730 GNDA.t84 65.8183
R10447 GNDA.t84 GNDA.n2633 65.8183
R10448 GNDA.t84 GNDA.n2632 65.8183
R10449 GNDA.t84 GNDA.n2630 65.8183
R10450 GNDA.t120 GNDA.n4971 65.8183
R10451 GNDA.t120 GNDA.n4893 65.8183
R10452 GNDA.t120 GNDA.n4892 65.8183
R10453 GNDA.t120 GNDA.n4891 65.8183
R10454 GNDA.t120 GNDA.n4882 65.8183
R10455 GNDA.t120 GNDA.n4889 65.8183
R10456 GNDA.t120 GNDA.n4880 65.8183
R10457 GNDA.t120 GNDA.n4890 65.8183
R10458 GNDA.t120 GNDA.n4888 65.8183
R10459 GNDA.t120 GNDA.n4887 65.8183
R10460 GNDA.t120 GNDA.n4886 65.8183
R10461 GNDA.t120 GNDA.n4885 65.8183
R10462 GNDA.t120 GNDA.n4883 65.8183
R10463 GNDA.t120 GNDA.n4881 65.8183
R10464 GNDA.n4972 GNDA.t120 65.8183
R10465 GNDA.t120 GNDA.n4875 65.8183
R10466 GNDA.t46 GNDA.n5250 65.8183
R10467 GNDA.t46 GNDA.n79 65.8183
R10468 GNDA.t46 GNDA.n78 65.8183
R10469 GNDA.t46 GNDA.n77 65.8183
R10470 GNDA.t46 GNDA.n68 65.8183
R10471 GNDA.t46 GNDA.n75 65.8183
R10472 GNDA.t46 GNDA.n66 65.8183
R10473 GNDA.t46 GNDA.n76 65.8183
R10474 GNDA.t46 GNDA.n74 65.8183
R10475 GNDA.t46 GNDA.n73 65.8183
R10476 GNDA.t46 GNDA.n72 65.8183
R10477 GNDA.t46 GNDA.n71 65.8183
R10478 GNDA.t46 GNDA.n69 65.8183
R10479 GNDA.t46 GNDA.n67 65.8183
R10480 GNDA.n5251 GNDA.t46 65.8183
R10481 GNDA.t46 GNDA.n61 65.8183
R10482 GNDA.t44 GNDA.n4736 65.8183
R10483 GNDA.t44 GNDA.n4734 65.8183
R10484 GNDA.t44 GNDA.n4733 65.8183
R10485 GNDA.n4833 GNDA.t44 65.8183
R10486 GNDA.n2472 GNDA.t91 65.8183
R10487 GNDA.n2474 GNDA.t91 65.8183
R10488 GNDA.n2480 GNDA.t91 65.8183
R10489 GNDA.n2482 GNDA.t91 65.8183
R10490 GNDA.n2456 GNDA.t91 65.8183
R10491 GNDA.n2458 GNDA.t91 65.8183
R10492 GNDA.n2464 GNDA.t91 65.8183
R10493 GNDA.n2466 GNDA.t91 65.8183
R10494 GNDA.n2269 GNDA.t91 65.8183
R10495 GNDA.n2441 GNDA.t91 65.8183
R10496 GNDA.n2266 GNDA.t91 65.8183
R10497 GNDA.n2448 GNDA.t91 65.8183
R10498 GNDA.n2434 GNDA.t91 65.8183
R10499 GNDA.n2419 GNDA.t91 65.8183
R10500 GNDA.n2417 GNDA.t91 65.8183
R10501 GNDA.n2494 GNDA.t91 65.8183
R10502 GNDA.t47 GNDA.n19 65.8183
R10503 GNDA.t47 GNDA.n18 65.8183
R10504 GNDA.t47 GNDA.n17 65.8183
R10505 GNDA.t47 GNDA.n16 65.8183
R10506 GNDA.t47 GNDA.n7 65.8183
R10507 GNDA.t47 GNDA.n14 65.8183
R10508 GNDA.t47 GNDA.n5 65.8183
R10509 GNDA.t47 GNDA.n15 65.8183
R10510 GNDA.t47 GNDA.n13 65.8183
R10511 GNDA.t47 GNDA.n12 65.8183
R10512 GNDA.t47 GNDA.n11 65.8183
R10513 GNDA.t47 GNDA.n10 65.8183
R10514 GNDA.t47 GNDA.n8 65.8183
R10515 GNDA.n5274 GNDA.t47 65.8183
R10516 GNDA.t47 GNDA.n6 65.8183
R10517 GNDA.t47 GNDA.n4 65.8183
R10518 GNDA.t278 GNDA.t166 64.5933
R10519 GNDA.n3048 GNDA.n3047 63.1009
R10520 GNDA.t0 GNDA.t12 63.0554
R10521 GNDA.n3138 GNDA.t80 62.2505
R10522 GNDA.n3139 GNDA.t68 62.2505
R10523 GNDA.n1320 GNDA.t105 62.2505
R10524 GNDA.n3144 GNDA.t83 62.2505
R10525 GNDA.n3135 GNDA.t110 62.2505
R10526 GNDA.n3130 GNDA.t75 62.2505
R10527 GNDA.n634 GNDA.t100 62.2505
R10528 GNDA.n630 GNDA.t102 62.2505
R10529 GNDA.n433 GNDA.t133 62.2505
R10530 GNDA.n3146 GNDA.t115 62.2505
R10531 GNDA.n637 GNDA.t135 62.2505
R10532 GNDA.n639 GNDA.t113 62.2505
R10533 GNDA.n3075 GNDA.t192 62.0993
R10534 GNDA.n2985 GNDA.t237 62.0993
R10535 GNDA.n4621 GNDA.n4620 59.2425
R10536 GNDA.n3154 GNDA.n3153 59.2425
R10537 GNDA.n1748 GNDA.n1747 59.2425
R10538 GNDA.n3859 GNDA.n432 59.2425
R10539 GNDA.t226 GNDA.n2428 58.0929
R10540 GNDA.n2308 GNDA.t190 58.0929
R10541 GNDA.t128 GNDA.n3004 57.8461
R10542 GNDA.t72 GNDA.n3081 57.8461
R10543 GNDA.t59 GNDA.n5047 57.8461
R10544 GNDA.t84 GNDA.n2729 57.8461
R10545 GNDA.t120 GNDA.n4874 57.8461
R10546 GNDA.t46 GNDA.n60 57.8461
R10547 GNDA.t44 GNDA.n4832 57.8461
R10548 GNDA.n2488 GNDA.t91 57.8461
R10549 GNDA.t47 GNDA.n5273 57.8461
R10550 GNDA.n2321 GNDA.n675 57.0913
R10551 GNDA.n694 GNDA.n691 56.3995
R10552 GNDA.n2741 GNDA.n2624 56.3995
R10553 GNDA.n4869 GNDA.n4868 56.3995
R10554 GNDA.n4845 GNDA.n234 56.3995
R10555 GNDA.n3036 GNDA.n691 56.3995
R10556 GNDA.n2741 GNDA.n2740 56.3995
R10557 GNDA.n5100 GNDA.n5099 56.3995
R10558 GNDA.n5101 GNDA.n5100 56.3995
R10559 GNDA.n835 GNDA.n280 56.3995
R10560 GNDA.n4868 GNDA.n227 56.3995
R10561 GNDA.n4843 GNDA.n234 56.3995
R10562 GNDA.t128 GNDA.n730 55.2026
R10563 GNDA.t72 GNDA.n658 55.2026
R10564 GNDA.t59 GNDA.n175 55.2026
R10565 GNDA.t44 GNDA.n4737 55.2026
R10566 GNDA.t84 GNDA.n2635 55.2026
R10567 GNDA.t120 GNDA.n4884 55.2026
R10568 GNDA.t46 GNDA.n70 55.2026
R10569 GNDA.n2450 GNDA.t91 55.2026
R10570 GNDA.t47 GNDA.n9 55.2026
R10571 GNDA.n784 GNDA.n738 53.3664
R10572 GNDA.n780 GNDA.n718 53.3664
R10573 GNDA.n776 GNDA.n737 53.3664
R10574 GNDA.n772 GNDA.n720 53.3664
R10575 GNDA.n761 GNDA.n731 53.3664
R10576 GNDA.n757 GNDA.n732 53.3664
R10577 GNDA.n753 GNDA.n733 53.3664
R10578 GNDA.n736 GNDA.n735 53.3664
R10579 GNDA.n744 GNDA.n717 53.3664
R10580 GNDA.n2993 GNDA.n719 53.3664
R10581 GNDA.n3006 GNDA.n3005 53.3664
R10582 GNDA.n729 GNDA.n728 53.3664
R10583 GNDA.n788 GNDA.n742 53.3664
R10584 GNDA.n789 GNDA.n741 53.3664
R10585 GNDA.n793 GNDA.n740 53.3664
R10586 GNDA.n797 GNDA.n739 53.3664
R10587 GNDA.n785 GNDA.n742 53.3664
R10588 GNDA.n792 GNDA.n741 53.3664
R10589 GNDA.n796 GNDA.n740 53.3664
R10590 GNDA.n799 GNDA.n739 53.3664
R10591 GNDA.n769 GNDA.n720 53.3664
R10592 GNDA.n773 GNDA.n737 53.3664
R10593 GNDA.n777 GNDA.n718 53.3664
R10594 GNDA.n781 GNDA.n738 53.3664
R10595 GNDA.n752 GNDA.n736 53.3664
R10596 GNDA.n756 GNDA.n733 53.3664
R10597 GNDA.n760 GNDA.n732 53.3664
R10598 GNDA.n764 GNDA.n731 53.3664
R10599 GNDA.n734 GNDA.n729 53.3664
R10600 GNDA.n3005 GNDA.n716 53.3664
R10601 GNDA.n719 GNDA.n715 53.3664
R10602 GNDA.n2992 GNDA.n717 53.3664
R10603 GNDA.n2342 GNDA.n664 53.3664
R10604 GNDA.n2346 GNDA.n654 53.3664
R10605 GNDA.n2350 GNDA.n663 53.3664
R10606 GNDA.n2354 GNDA.n656 53.3664
R10607 GNDA.n2365 GNDA.n659 53.3664
R10608 GNDA.n2369 GNDA.n660 53.3664
R10609 GNDA.n2373 GNDA.n661 53.3664
R10610 GNDA.n2377 GNDA.n662 53.3664
R10611 GNDA.n670 GNDA.n653 53.3664
R10612 GNDA.n3070 GNDA.n655 53.3664
R10613 GNDA.n3083 GNDA.n3082 53.3664
R10614 GNDA.n2311 GNDA.n657 53.3664
R10615 GNDA.n2338 GNDA.n668 53.3664
R10616 GNDA.n2337 GNDA.n667 53.3664
R10617 GNDA.n2333 GNDA.n666 53.3664
R10618 GNDA.n2329 GNDA.n665 53.3664
R10619 GNDA.n2341 GNDA.n668 53.3664
R10620 GNDA.n2334 GNDA.n667 53.3664
R10621 GNDA.n2330 GNDA.n666 53.3664
R10622 GNDA.n2326 GNDA.n665 53.3664
R10623 GNDA.n2357 GNDA.n656 53.3664
R10624 GNDA.n2353 GNDA.n663 53.3664
R10625 GNDA.n2349 GNDA.n654 53.3664
R10626 GNDA.n2345 GNDA.n664 53.3664
R10627 GNDA.n2374 GNDA.n662 53.3664
R10628 GNDA.n2370 GNDA.n661 53.3664
R10629 GNDA.n2366 GNDA.n660 53.3664
R10630 GNDA.n2362 GNDA.n659 53.3664
R10631 GNDA.n2376 GNDA.n657 53.3664
R10632 GNDA.n3082 GNDA.n652 53.3664
R10633 GNDA.n655 GNDA.n651 53.3664
R10634 GNDA.n3069 GNDA.n653 53.3664
R10635 GNDA.n5029 GNDA.n181 53.3664
R10636 GNDA.n5025 GNDA.n170 53.3664
R10637 GNDA.n5021 GNDA.n180 53.3664
R10638 GNDA.n5017 GNDA.n173 53.3664
R10639 GNDA.n5006 GNDA.n176 53.3664
R10640 GNDA.n5002 GNDA.n177 53.3664
R10641 GNDA.n4998 GNDA.n178 53.3664
R10642 GNDA.n4994 GNDA.n179 53.3664
R10643 GNDA.n5049 GNDA.n5048 53.3664
R10644 GNDA.n216 GNDA.n171 53.3664
R10645 GNDA.n212 GNDA.n172 53.3664
R10646 GNDA.n205 GNDA.n174 53.3664
R10647 GNDA.n5033 GNDA.n185 53.3664
R10648 GNDA.n5034 GNDA.n184 53.3664
R10649 GNDA.n5038 GNDA.n183 53.3664
R10650 GNDA.n5042 GNDA.n182 53.3664
R10651 GNDA.n5030 GNDA.n185 53.3664
R10652 GNDA.n5037 GNDA.n184 53.3664
R10653 GNDA.n5041 GNDA.n183 53.3664
R10654 GNDA.n5045 GNDA.n182 53.3664
R10655 GNDA.n5014 GNDA.n173 53.3664
R10656 GNDA.n5018 GNDA.n180 53.3664
R10657 GNDA.n5022 GNDA.n170 53.3664
R10658 GNDA.n5026 GNDA.n181 53.3664
R10659 GNDA.n4997 GNDA.n179 53.3664
R10660 GNDA.n5001 GNDA.n178 53.3664
R10661 GNDA.n5005 GNDA.n177 53.3664
R10662 GNDA.n5009 GNDA.n176 53.3664
R10663 GNDA.n4993 GNDA.n174 53.3664
R10664 GNDA.n204 GNDA.n172 53.3664
R10665 GNDA.n213 GNDA.n171 53.3664
R10666 GNDA.n5048 GNDA.n169 53.3664
R10667 GNDA.n4814 GNDA.n4743 53.3664
R10668 GNDA.n4810 GNDA.n4732 53.3664
R10669 GNDA.n4806 GNDA.n4742 53.3664
R10670 GNDA.n4802 GNDA.n4735 53.3664
R10671 GNDA.n4791 GNDA.n4738 53.3664
R10672 GNDA.n4787 GNDA.n4739 53.3664
R10673 GNDA.n4783 GNDA.n4740 53.3664
R10674 GNDA.n4779 GNDA.n4741 53.3664
R10675 GNDA.n4834 GNDA.n4833 53.3664
R10676 GNDA.n4756 GNDA.n4733 53.3664
R10677 GNDA.n4764 GNDA.n4734 53.3664
R10678 GNDA.n4771 GNDA.n4736 53.3664
R10679 GNDA.n4818 GNDA.n4747 53.3664
R10680 GNDA.n4819 GNDA.n4746 53.3664
R10681 GNDA.n4823 GNDA.n4745 53.3664
R10682 GNDA.n4827 GNDA.n4744 53.3664
R10683 GNDA.n4815 GNDA.n4747 53.3664
R10684 GNDA.n4822 GNDA.n4746 53.3664
R10685 GNDA.n4826 GNDA.n4745 53.3664
R10686 GNDA.n4830 GNDA.n4744 53.3664
R10687 GNDA.n4799 GNDA.n4735 53.3664
R10688 GNDA.n4803 GNDA.n4742 53.3664
R10689 GNDA.n4807 GNDA.n4732 53.3664
R10690 GNDA.n4811 GNDA.n4743 53.3664
R10691 GNDA.n4782 GNDA.n4741 53.3664
R10692 GNDA.n4786 GNDA.n4740 53.3664
R10693 GNDA.n4790 GNDA.n4739 53.3664
R10694 GNDA.n4794 GNDA.n4738 53.3664
R10695 GNDA.n2682 GNDA.n2642 53.3664
R10696 GNDA.n2678 GNDA.n2631 53.3664
R10697 GNDA.n2674 GNDA.n2641 53.3664
R10698 GNDA.n2670 GNDA.n2634 53.3664
R10699 GNDA.n2659 GNDA.n2636 53.3664
R10700 GNDA.n2655 GNDA.n2637 53.3664
R10701 GNDA.n2651 GNDA.n2638 53.3664
R10702 GNDA.n2640 GNDA.n2639 53.3664
R10703 GNDA.n2648 GNDA.n2630 53.3664
R10704 GNDA.n2717 GNDA.n2632 53.3664
R10705 GNDA.n2710 GNDA.n2633 53.3664
R10706 GNDA.n2731 GNDA.n2730 53.3664
R10707 GNDA.n2686 GNDA.n2646 53.3664
R10708 GNDA.n2687 GNDA.n2645 53.3664
R10709 GNDA.n2691 GNDA.n2644 53.3664
R10710 GNDA.n2695 GNDA.n2643 53.3664
R10711 GNDA.n2683 GNDA.n2646 53.3664
R10712 GNDA.n2690 GNDA.n2645 53.3664
R10713 GNDA.n2694 GNDA.n2644 53.3664
R10714 GNDA.n2697 GNDA.n2643 53.3664
R10715 GNDA.n2667 GNDA.n2634 53.3664
R10716 GNDA.n2671 GNDA.n2641 53.3664
R10717 GNDA.n2675 GNDA.n2631 53.3664
R10718 GNDA.n2679 GNDA.n2642 53.3664
R10719 GNDA.n2650 GNDA.n2640 53.3664
R10720 GNDA.n2654 GNDA.n2638 53.3664
R10721 GNDA.n2658 GNDA.n2637 53.3664
R10722 GNDA.n2662 GNDA.n2636 53.3664
R10723 GNDA.n2730 GNDA.n2629 53.3664
R10724 GNDA.n2633 GNDA.n2628 53.3664
R10725 GNDA.n2709 GNDA.n2632 53.3664
R10726 GNDA.n2716 GNDA.n2630 53.3664
R10727 GNDA.n4954 GNDA.n4890 53.3664
R10728 GNDA.n4951 GNDA.n4880 53.3664
R10729 GNDA.n4947 GNDA.n4889 53.3664
R10730 GNDA.n4943 GNDA.n4882 53.3664
R10731 GNDA.n4932 GNDA.n4885 53.3664
R10732 GNDA.n4928 GNDA.n4886 53.3664
R10733 GNDA.n4924 GNDA.n4887 53.3664
R10734 GNDA.n4920 GNDA.n4888 53.3664
R10735 GNDA.n4980 GNDA.n4875 53.3664
R10736 GNDA.n4973 GNDA.n4972 53.3664
R10737 GNDA.n4905 GNDA.n4881 53.3664
R10738 GNDA.n4912 GNDA.n4883 53.3664
R10739 GNDA.n4971 GNDA.n4970 53.3664
R10740 GNDA.n4895 GNDA.n4893 53.3664
R10741 GNDA.n4965 GNDA.n4892 53.3664
R10742 GNDA.n4961 GNDA.n4891 53.3664
R10743 GNDA.n4971 GNDA.n4894 53.3664
R10744 GNDA.n4966 GNDA.n4893 53.3664
R10745 GNDA.n4962 GNDA.n4892 53.3664
R10746 GNDA.n4958 GNDA.n4891 53.3664
R10747 GNDA.n4940 GNDA.n4882 53.3664
R10748 GNDA.n4944 GNDA.n4889 53.3664
R10749 GNDA.n4948 GNDA.n4880 53.3664
R10750 GNDA.n4952 GNDA.n4890 53.3664
R10751 GNDA.n4923 GNDA.n4888 53.3664
R10752 GNDA.n4927 GNDA.n4887 53.3664
R10753 GNDA.n4931 GNDA.n4886 53.3664
R10754 GNDA.n4935 GNDA.n4885 53.3664
R10755 GNDA.n4919 GNDA.n4883 53.3664
R10756 GNDA.n4911 GNDA.n4881 53.3664
R10757 GNDA.n4972 GNDA.n4879 53.3664
R10758 GNDA.n4878 GNDA.n4875 53.3664
R10759 GNDA.n5233 GNDA.n76 53.3664
R10760 GNDA.n5230 GNDA.n66 53.3664
R10761 GNDA.n5226 GNDA.n75 53.3664
R10762 GNDA.n5222 GNDA.n68 53.3664
R10763 GNDA.n5211 GNDA.n71 53.3664
R10764 GNDA.n5207 GNDA.n72 53.3664
R10765 GNDA.n5203 GNDA.n73 53.3664
R10766 GNDA.n5199 GNDA.n74 53.3664
R10767 GNDA.n5259 GNDA.n61 53.3664
R10768 GNDA.n5252 GNDA.n5251 53.3664
R10769 GNDA.n5184 GNDA.n67 53.3664
R10770 GNDA.n5191 GNDA.n69 53.3664
R10771 GNDA.n5250 GNDA.n5249 53.3664
R10772 GNDA.n81 GNDA.n79 53.3664
R10773 GNDA.n5244 GNDA.n78 53.3664
R10774 GNDA.n5240 GNDA.n77 53.3664
R10775 GNDA.n5250 GNDA.n80 53.3664
R10776 GNDA.n5245 GNDA.n79 53.3664
R10777 GNDA.n5241 GNDA.n78 53.3664
R10778 GNDA.n5237 GNDA.n77 53.3664
R10779 GNDA.n5219 GNDA.n68 53.3664
R10780 GNDA.n5223 GNDA.n75 53.3664
R10781 GNDA.n5227 GNDA.n66 53.3664
R10782 GNDA.n5231 GNDA.n76 53.3664
R10783 GNDA.n5202 GNDA.n74 53.3664
R10784 GNDA.n5206 GNDA.n73 53.3664
R10785 GNDA.n5210 GNDA.n72 53.3664
R10786 GNDA.n5214 GNDA.n71 53.3664
R10787 GNDA.n5198 GNDA.n69 53.3664
R10788 GNDA.n5190 GNDA.n67 53.3664
R10789 GNDA.n5251 GNDA.n65 53.3664
R10790 GNDA.n64 GNDA.n61 53.3664
R10791 GNDA.n4778 GNDA.n4736 53.3664
R10792 GNDA.n4770 GNDA.n4734 53.3664
R10793 GNDA.n4763 GNDA.n4733 53.3664
R10794 GNDA.n4833 GNDA.n4731 53.3664
R10795 GNDA.n2466 GNDA.n2258 53.3664
R10796 GNDA.n2465 GNDA.n2464 53.3664
R10797 GNDA.n2458 GNDA.n2260 53.3664
R10798 GNDA.n2457 GNDA.n2456 53.3664
R10799 GNDA.n2448 GNDA.n2447 53.3664
R10800 GNDA.n2443 GNDA.n2266 53.3664
R10801 GNDA.n2441 GNDA.n2440 53.3664
R10802 GNDA.n2436 GNDA.n2269 53.3664
R10803 GNDA.n2494 GNDA.n2493 53.3664
R10804 GNDA.n2417 GNDA.n2253 53.3664
R10805 GNDA.n2420 GNDA.n2419 53.3664
R10806 GNDA.n2434 GNDA.n2433 53.3664
R10807 GNDA.n2473 GNDA.n2472 53.3664
R10808 GNDA.n2475 GNDA.n2474 53.3664
R10809 GNDA.n2480 GNDA.n2479 53.3664
R10810 GNDA.n2483 GNDA.n2482 53.3664
R10811 GNDA.n2472 GNDA.n2471 53.3664
R10812 GNDA.n2474 GNDA.n2256 53.3664
R10813 GNDA.n2481 GNDA.n2480 53.3664
R10814 GNDA.n2482 GNDA.n2254 53.3664
R10815 GNDA.n2456 GNDA.n2455 53.3664
R10816 GNDA.n2459 GNDA.n2458 53.3664
R10817 GNDA.n2464 GNDA.n2463 53.3664
R10818 GNDA.n2467 GNDA.n2466 53.3664
R10819 GNDA.n2269 GNDA.n2267 53.3664
R10820 GNDA.n2442 GNDA.n2441 53.3664
R10821 GNDA.n2266 GNDA.n2264 53.3664
R10822 GNDA.n2449 GNDA.n2448 53.3664
R10823 GNDA.n2435 GNDA.n2434 53.3664
R10824 GNDA.n2419 GNDA.n2271 53.3664
R10825 GNDA.n2418 GNDA.n2417 53.3664
R10826 GNDA.n2495 GNDA.n2494 53.3664
R10827 GNDA.n5152 GNDA.n15 53.3664
R10828 GNDA.n5148 GNDA.n5 53.3664
R10829 GNDA.n5144 GNDA.n14 53.3664
R10830 GNDA.n5140 GNDA.n7 53.3664
R10831 GNDA.n5129 GNDA.n10 53.3664
R10832 GNDA.n5125 GNDA.n11 53.3664
R10833 GNDA.n5121 GNDA.n12 53.3664
R10834 GNDA.n5117 GNDA.n13 53.3664
R10835 GNDA.n21 GNDA.n4 53.3664
R10836 GNDA.n37 GNDA.n6 53.3664
R10837 GNDA.n5275 GNDA.n5274 53.3664
R10838 GNDA.n5109 GNDA.n8 53.3664
R10839 GNDA.n5156 GNDA.n19 53.3664
R10840 GNDA.n5157 GNDA.n18 53.3664
R10841 GNDA.n5161 GNDA.n17 53.3664
R10842 GNDA.n5165 GNDA.n16 53.3664
R10843 GNDA.n5153 GNDA.n19 53.3664
R10844 GNDA.n5160 GNDA.n18 53.3664
R10845 GNDA.n5164 GNDA.n17 53.3664
R10846 GNDA.n5167 GNDA.n16 53.3664
R10847 GNDA.n5137 GNDA.n7 53.3664
R10848 GNDA.n5141 GNDA.n14 53.3664
R10849 GNDA.n5145 GNDA.n5 53.3664
R10850 GNDA.n5149 GNDA.n15 53.3664
R10851 GNDA.n5120 GNDA.n13 53.3664
R10852 GNDA.n5124 GNDA.n12 53.3664
R10853 GNDA.n5128 GNDA.n11 53.3664
R10854 GNDA.n5132 GNDA.n10 53.3664
R10855 GNDA.n5116 GNDA.n8 53.3664
R10856 GNDA.n5274 GNDA.n3 53.3664
R10857 GNDA.n6 GNDA.n2 53.3664
R10858 GNDA.n36 GNDA.n4 53.3664
R10859 GNDA.t200 GNDA.t149 53.2263
R10860 GNDA.n2513 GNDA.n838 53.085
R10861 GNDA.n2321 GNDA.n2320 53.085
R10862 GNDA.n2387 GNDA.n2384 53.085
R10863 GNDA.n2428 GNDA.t212 52.0834
R10864 GNDA.n2308 GNDA.t230 52.0834
R10865 GNDA.n3010 GNDA.t17 52.0834
R10866 GNDA.n4723 GNDA.n99 50.8806
R10867 GNDA.n4723 GNDA.n4722 50.8806
R10868 GNDA.n4722 GNDA.n4721 50.8806
R10869 GNDA.n4721 GNDA.n292 50.8806
R10870 GNDA.n4715 GNDA.n292 50.8806
R10871 GNDA.n4714 GNDA.n4713 50.8806
R10872 GNDA.n4713 GNDA.n296 50.8806
R10873 GNDA.n4707 GNDA.n296 50.8806
R10874 GNDA.n4707 GNDA.n4706 50.8806
R10875 GNDA.n4706 GNDA.n4705 50.8806
R10876 GNDA.n4699 GNDA.n4698 50.8806
R10877 GNDA.n4698 GNDA.n4697 50.8806
R10878 GNDA.n4697 GNDA.n351 50.8806
R10879 GNDA.n4691 GNDA.n351 50.8806
R10880 GNDA.n4691 GNDA.n4690 50.8806
R10881 GNDA.n4681 GNDA.n356 50.8806
R10882 GNDA.n4681 GNDA.n4680 50.8806
R10883 GNDA.n4680 GNDA.n4679 50.8806
R10884 GNDA.n4679 GNDA.n362 50.8806
R10885 GNDA.n4673 GNDA.n362 50.8806
R10886 GNDA.n4671 GNDA.n367 50.8806
R10887 GNDA.n4665 GNDA.n367 50.8806
R10888 GNDA.n4665 GNDA.n4664 50.8806
R10889 GNDA.n4664 GNDA.n4663 50.8806
R10890 GNDA.n4663 GNDA.n416 50.8806
R10891 GNDA.n4657 GNDA.n4656 50.8806
R10892 GNDA.n4656 GNDA.n4655 50.8806
R10893 GNDA.n4655 GNDA.n420 50.8806
R10894 GNDA.n4649 GNDA.n420 50.8806
R10895 GNDA.n4649 GNDA.n4648 50.8806
R10896 GNDA.n3145 GNDA.n625 50.7468
R10897 GNDA.t187 GNDA.t174 48.7908
R10898 GNDA.t183 GNDA.t175 48.7908
R10899 GNDA.t184 GNDA.t172 48.7908
R10900 GNDA.t181 GNDA.t171 48.7908
R10901 GNDA.t180 GNDA.t170 48.7908
R10902 GNDA.t202 GNDA.t207 48.7908
R10903 GNDA.t194 GNDA.t279 48.7908
R10904 GNDA.t225 GNDA.t208 48.7908
R10905 GNDA.t163 GNDA.t203 48.7908
R10906 GNDA.t38 GNDA.t209 48.7908
R10907 GNDA.t139 GNDA.n106 48.077
R10908 GNDA.t70 GNDA.n3075 48.077
R10909 GNDA.n2985 GNDA.t160 48.077
R10910 GNDA.t45 GNDA.n5087 47.6748
R10911 GNDA.t45 GNDA.n106 47.0754
R10912 GNDA.n2983 GNDA.t243 47.0754
R10913 GNDA.t64 GNDA.t61 46.5731
R10914 GNDA.t55 GNDA.t77 46.5731
R10915 GNDA.t130 GNDA.t89 46.5731
R10916 GNDA.t126 GNDA.t86 46.5731
R10917 GNDA.t248 GNDA.n2974 46.0738
R10918 GNDA.t24 GNDA.t141 44.3553
R10919 GNDA.t206 GNDA.t142 44.3553
R10920 GNDA.n2320 GNDA.n809 43.069
R10921 GNDA.t45 GNDA.n3087 43.069
R10922 GNDA.t45 GNDA.n3010 43.069
R10923 GNDA.n3076 GNDA.t70 42.0674
R10924 GNDA.t160 GNDA.n2984 42.0674
R10925 GNDA.n3064 GNDA.t6 41.0658
R10926 GNDA.n1273 GNDA.t137 40.4338
R10927 GNDA.n1271 GNDA.t58 40.4338
R10928 GNDA.n3126 GNDA.t124 40.4338
R10929 GNDA.t98 GNDA.n3100 40.4338
R10930 GNDA.t104 GNDA.n431 40.299
R10931 GNDA.n3145 GNDA.t82 40.299
R10932 GNDA.t45 GNDA.t243 40.0642
R10933 GNDA.t212 GNDA.n2427 38.0611
R10934 GNDA.t230 GNDA.n2307 38.0611
R10935 GNDA.t174 GNDA.t158 37.7021
R10936 GNDA.t30 GNDA.t180 37.7021
R10937 GNDA.t15 GNDA.t202 37.7021
R10938 GNDA.t209 GNDA.t214 37.7021
R10939 GNDA.n3124 GNDA.n3123 37.5297
R10940 GNDA.n3122 GNDA.n3121 37.5297
R10941 GNDA.n3120 GNDA.n3119 37.5297
R10942 GNDA.n3118 GNDA.n3117 37.5297
R10943 GNDA.n3116 GNDA.n3115 37.5297
R10944 GNDA.n3114 GNDA.n3113 37.5297
R10945 GNDA.n3112 GNDA.n3111 37.5297
R10946 GNDA.n3110 GNDA.n3109 37.5297
R10947 GNDA.n3108 GNDA.n3107 37.5297
R10948 GNDA.n3106 GNDA.n3105 37.5297
R10949 GNDA.n3104 GNDA.n3103 37.5297
R10950 GNDA.n3102 GNDA.n3101 37.5297
R10951 GNDA.n2514 GNDA.n2513 37.0595
R10952 GNDA.n2249 GNDA.t201 37.0595
R10953 GNDA.n2387 GNDA.n2383 37.0595
R10954 GNDA.t49 GNDA.t248 35.0563
R10955 GNDA.n1341 GNDA.n1340 34.5991
R10956 GNDA.n1747 GNDA.t64 33.2666
R10957 GNDA.n3153 GNDA.t77 33.2666
R10958 GNDA.t89 GNDA.n432 33.2666
R10959 GNDA.n4621 GNDA.t126 33.2666
R10960 GNDA.t210 GNDA.t288 33.1455
R10961 GNDA.n2407 GNDA.n2396 33.0531
R10962 GNDA.n722 GNDA.t9 33.0531
R10963 GNDA.t45 GNDA.n26 32.9056
R10964 GNDA.t45 GNDA.n107 32.9056
R10965 GNDA.t234 GNDA.t37 32.8363
R10966 GNDA.t37 GNDA.t104 32.8363
R10967 GNDA.t255 GNDA.t82 32.8363
R10968 GNDA.t162 GNDA.t255 32.8363
R10969 GNDA.n3024 GNDA.n3023 32.3969
R10970 GNDA.t190 GNDA.n2306 32.0515
R10971 GNDA.n434 GNDA.n433 31.5738
R10972 GNDA.n4686 GNDA.n4685 31.3605
R10973 GNDA.n1745 GNDA.t65 31.1255
R10974 GNDA.n4623 GNDA.t127 31.1255
R10975 GNDA.n4628 GNDA.t90 31.1255
R10976 GNDA.n3151 GNDA.t78 31.1255
R10977 GNDA.t42 GNDA.t284 30.3834
R10978 GNDA.t284 GNDA.t222 30.3834
R10979 GNDA.t222 GNDA.t232 30.3834
R10980 GNDA.n3062 GNDA.n675 30.0483
R10981 GNDA.n1321 GNDA.n1320 29.8672
R10982 GNDA.n3144 GNDA.n3143 29.8672
R10983 GNDA.n3147 GNDA.n3146 29.8672
R10984 GNDA.n2974 GNDA.t290 29.0467
R10985 GNDA.t175 GNDA.t235 28.8311
R10986 GNDA.t267 GNDA.t181 28.8311
R10987 GNDA.t259 GNDA.t194 28.8311
R10988 GNDA.t203 GNDA.t4 28.8311
R10989 GNDA.t192 GNDA.n3074 28.0451
R10990 GNDA.t52 GNDA.n2983 28.0451
R10991 GNDA.n786 GNDA.n783 27.5561
R10992 GNDA.n2343 GNDA.n2340 27.5561
R10993 GNDA.n5031 GNDA.n5028 27.5561
R10994 GNDA.n4816 GNDA.n4813 27.5561
R10995 GNDA.n2684 GNDA.n2681 27.5561
R10996 GNDA.n4956 GNDA.n4955 27.5561
R10997 GNDA.n5235 GNDA.n5234 27.5561
R10998 GNDA.n2470 GNDA.n2469 27.5561
R10999 GNDA.n5154 GNDA.n5151 27.5561
R11000 GNDA.n2384 GNDA.n808 27.0435
R11001 GNDA.n3021 GNDA.n707 27.0435
R11002 GNDA.n3048 GNDA.n685 27.0435
R11003 GNDA.n767 GNDA.n766 26.6672
R11004 GNDA.n2360 GNDA.n2359 26.6672
R11005 GNDA.n5012 GNDA.n5011 26.6672
R11006 GNDA.n4797 GNDA.n4796 26.6672
R11007 GNDA.n2665 GNDA.n2664 26.6672
R11008 GNDA.n4938 GNDA.n4937 26.6672
R11009 GNDA.n5217 GNDA.n5216 26.6672
R11010 GNDA.n2453 GNDA.n2452 26.6672
R11011 GNDA.n5135 GNDA.n5134 26.6672
R11012 GNDA.n1747 GNDA.n1746 26.6134
R11013 GNDA.n3153 GNDA.n3152 26.6134
R11014 GNDA.n4629 GNDA.n432 26.6134
R11015 GNDA.n4622 GNDA.n4621 26.6134
R11016 GNDA.n4715 GNDA.t45 26.5712
R11017 GNDA.n4690 GNDA.t45 26.5712
R11018 GNDA.t45 GNDA.n416 26.5712
R11019 GNDA.t252 GNDA.n3127 25.3736
R11020 GNDA.n3099 GNDA.t211 25.3736
R11021 GNDA.n2399 GNDA.n2398 25.3679
R11022 GNDA.t256 GNDA.t226 25.0403
R11023 GNDA.t237 GNDA.t7 25.0403
R11024 GNDA.t45 GNDA.n4714 24.3099
R11025 GNDA.t45 GNDA.n356 24.3099
R11026 GNDA.n4657 GNDA.t45 24.3099
R11027 GNDA.n696 GNDA.n686 24.0387
R11028 GNDA.n684 GNDA.t36 24.0005
R11029 GNDA.n684 GNDA.t18 24.0005
R11030 GNDA.n683 GNDA.t229 24.0005
R11031 GNDA.n683 GNDA.t262 24.0005
R11032 GNDA.n682 GNDA.t161 24.0005
R11033 GNDA.n682 GNDA.t238 24.0005
R11034 GNDA.n679 GNDA.t231 24.0005
R11035 GNDA.n679 GNDA.t118 24.0005
R11036 GNDA.n678 GNDA.t146 24.0005
R11037 GNDA.n678 GNDA.t191 24.0005
R11038 GNDA.n677 GNDA.t193 24.0005
R11039 GNDA.n677 GNDA.t218 24.0005
R11040 GNDA.n2505 GNDA.t213 24.0005
R11041 GNDA.n2505 GNDA.t291 24.0005
R11042 GNDA.n2504 GNDA.t144 24.0005
R11043 GNDA.n2504 GNDA.t227 24.0005
R11044 GNDA.n2503 GNDA.t258 24.0005
R11045 GNDA.n2503 GNDA.t22 24.0005
R11046 GNDA.n2246 GNDA.t233 24.0005
R11047 GNDA.n2246 GNDA.t94 24.0005
R11048 GNDA.n2244 GNDA.t285 24.0005
R11049 GNDA.n2244 GNDA.t223 24.0005
R11050 GNDA.n2240 GNDA.t263 23.4782
R11051 GNDA.n2410 GNDA.n2409 23.0371
R11052 GNDA.n807 GNDA.n680 22.53
R11053 GNDA.n3050 GNDA.n3049 20.8233
R11054 GNDA.n2975 GNDA.n681 20.8233
R11055 GNDA.n3061 GNDA.n3060 20.8233
R11056 GNDA.n2319 GNDA.n2318 20.8233
R11057 GNDA.n2502 GNDA.n2501 20.8233
R11058 GNDA.n2512 GNDA.n2511 20.8233
R11059 GNDA.n2242 GNDA.n2241 20.8233
R11060 GNDA.n2976 GNDA.t45 20.0324
R11061 GNDA.t235 GNDA.t184 19.9602
R11062 GNDA.t172 GNDA.t267 19.9602
R11063 GNDA.t208 GNDA.t259 19.9602
R11064 GNDA.t4 GNDA.t225 19.9602
R11065 GNDA.n1305 GNDA.t164 19.7005
R11066 GNDA.n1305 GNDA.t250 19.7005
R11067 GNDA.n1307 GNDA.t10 19.7005
R11068 GNDA.n1307 GNDA.t195 19.7005
R11069 GNDA.n1309 GNDA.t11 19.7005
R11070 GNDA.n1309 GNDA.t269 19.7005
R11071 GNDA.n1311 GNDA.t196 19.7005
R11072 GNDA.n1311 GNDA.t265 19.7005
R11073 GNDA.n1313 GNDA.t266 19.7005
R11074 GNDA.n1313 GNDA.t276 19.7005
R11075 GNDA.n1315 GNDA.t245 19.7005
R11076 GNDA.n1315 GNDA.t270 19.7005
R11077 GNDA.n1365 GNDA.t182 19.7005
R11078 GNDA.n1365 GNDA.t242 19.7005
R11079 GNDA.n1367 GNDA.t186 19.7005
R11080 GNDA.n1367 GNDA.t173 19.7005
R11081 GNDA.n1369 GNDA.t185 19.7005
R11082 GNDA.n1369 GNDA.t177 19.7005
R11083 GNDA.n1371 GNDA.t189 19.7005
R11084 GNDA.n1371 GNDA.t176 19.7005
R11085 GNDA.n1373 GNDA.t188 19.7005
R11086 GNDA.n1373 GNDA.t179 19.7005
R11087 GNDA.n1375 GNDA.t241 19.7005
R11088 GNDA.n1375 GNDA.t178 19.7005
R11089 GNDA.n4634 GNDA.t167 19.2245
R11090 GNDA.t167 GNDA.t27 18.4556
R11091 GNDA.t27 GNDA.t0 18.4556
R11092 GNDA.t166 GNDA.t287 18.4556
R11093 GNDA.t287 GNDA.t282 18.4556
R11094 GNDA.n2383 GNDA.t117 18.0292
R11095 GNDA.t14 GNDA.t150 17.9109
R11096 GNDA.t20 GNDA.t122 17.9109
R11097 GNDA.t97 GNDA.t23 17.9109
R11098 GNDA.t220 GNDA.t251 17.9109
R11099 GNDA.n2894 GNDA.n2868 17.5843
R11100 GNDA.n2765 GNDA.n2613 17.5843
R11101 GNDA.n4645 GNDA.n422 17.5843
R11102 GNDA.n4641 GNDA.n4634 17.5479
R11103 GNDA.n262 GNDA.n259 16.9379
R11104 GNDA.n4864 GNDA.n4726 16.9379
R11105 GNDA.n2540 GNDA.n2539 16.9379
R11106 GNDA.n5083 GNDA.n133 16.7709
R11107 GNDA.n2564 GNDA.n162 16.7709
R11108 GNDA.n2612 GNDA.n84 16.7709
R11109 GNDA.n2824 GNDA.n2823 16.7709
R11110 GNDA.t45 GNDA.n105 16.4553
R11111 GNDA.n787 GNDA.n786 16.0005
R11112 GNDA.n790 GNDA.n787 16.0005
R11113 GNDA.n791 GNDA.n790 16.0005
R11114 GNDA.n794 GNDA.n791 16.0005
R11115 GNDA.n795 GNDA.n794 16.0005
R11116 GNDA.n798 GNDA.n795 16.0005
R11117 GNDA.n800 GNDA.n798 16.0005
R11118 GNDA.n801 GNDA.n800 16.0005
R11119 GNDA.n783 GNDA.n782 16.0005
R11120 GNDA.n782 GNDA.n779 16.0005
R11121 GNDA.n779 GNDA.n778 16.0005
R11122 GNDA.n778 GNDA.n775 16.0005
R11123 GNDA.n775 GNDA.n774 16.0005
R11124 GNDA.n774 GNDA.n771 16.0005
R11125 GNDA.n771 GNDA.n770 16.0005
R11126 GNDA.n770 GNDA.n767 16.0005
R11127 GNDA.n766 GNDA.n763 16.0005
R11128 GNDA.n763 GNDA.n762 16.0005
R11129 GNDA.n762 GNDA.n759 16.0005
R11130 GNDA.n759 GNDA.n758 16.0005
R11131 GNDA.n758 GNDA.n755 16.0005
R11132 GNDA.n755 GNDA.n754 16.0005
R11133 GNDA.n754 GNDA.n751 16.0005
R11134 GNDA.n751 GNDA.n690 16.0005
R11135 GNDA.n2340 GNDA.n2339 16.0005
R11136 GNDA.n2339 GNDA.n2336 16.0005
R11137 GNDA.n2336 GNDA.n2335 16.0005
R11138 GNDA.n2335 GNDA.n2332 16.0005
R11139 GNDA.n2332 GNDA.n2331 16.0005
R11140 GNDA.n2331 GNDA.n2328 16.0005
R11141 GNDA.n2328 GNDA.n2327 16.0005
R11142 GNDA.n2327 GNDA.n2325 16.0005
R11143 GNDA.n2344 GNDA.n2343 16.0005
R11144 GNDA.n2347 GNDA.n2344 16.0005
R11145 GNDA.n2348 GNDA.n2347 16.0005
R11146 GNDA.n2351 GNDA.n2348 16.0005
R11147 GNDA.n2352 GNDA.n2351 16.0005
R11148 GNDA.n2355 GNDA.n2352 16.0005
R11149 GNDA.n2356 GNDA.n2355 16.0005
R11150 GNDA.n2359 GNDA.n2356 16.0005
R11151 GNDA.n2363 GNDA.n2360 16.0005
R11152 GNDA.n2364 GNDA.n2363 16.0005
R11153 GNDA.n2367 GNDA.n2364 16.0005
R11154 GNDA.n2368 GNDA.n2367 16.0005
R11155 GNDA.n2371 GNDA.n2368 16.0005
R11156 GNDA.n2372 GNDA.n2371 16.0005
R11157 GNDA.n2375 GNDA.n2372 16.0005
R11158 GNDA.n2378 GNDA.n2375 16.0005
R11159 GNDA.n5032 GNDA.n5031 16.0005
R11160 GNDA.n5035 GNDA.n5032 16.0005
R11161 GNDA.n5036 GNDA.n5035 16.0005
R11162 GNDA.n5039 GNDA.n5036 16.0005
R11163 GNDA.n5040 GNDA.n5039 16.0005
R11164 GNDA.n5043 GNDA.n5040 16.0005
R11165 GNDA.n5044 GNDA.n5043 16.0005
R11166 GNDA.n5044 GNDA.n164 16.0005
R11167 GNDA.n5028 GNDA.n5027 16.0005
R11168 GNDA.n5027 GNDA.n5024 16.0005
R11169 GNDA.n5024 GNDA.n5023 16.0005
R11170 GNDA.n5023 GNDA.n5020 16.0005
R11171 GNDA.n5020 GNDA.n5019 16.0005
R11172 GNDA.n5019 GNDA.n5016 16.0005
R11173 GNDA.n5016 GNDA.n5015 16.0005
R11174 GNDA.n5015 GNDA.n5012 16.0005
R11175 GNDA.n5011 GNDA.n5008 16.0005
R11176 GNDA.n5008 GNDA.n5007 16.0005
R11177 GNDA.n5007 GNDA.n5004 16.0005
R11178 GNDA.n5004 GNDA.n5003 16.0005
R11179 GNDA.n5003 GNDA.n5000 16.0005
R11180 GNDA.n5000 GNDA.n4999 16.0005
R11181 GNDA.n4999 GNDA.n4996 16.0005
R11182 GNDA.n4996 GNDA.n4995 16.0005
R11183 GNDA.n4817 GNDA.n4816 16.0005
R11184 GNDA.n4820 GNDA.n4817 16.0005
R11185 GNDA.n4821 GNDA.n4820 16.0005
R11186 GNDA.n4824 GNDA.n4821 16.0005
R11187 GNDA.n4825 GNDA.n4824 16.0005
R11188 GNDA.n4828 GNDA.n4825 16.0005
R11189 GNDA.n4829 GNDA.n4828 16.0005
R11190 GNDA.n4829 GNDA.n4727 16.0005
R11191 GNDA.n4813 GNDA.n4812 16.0005
R11192 GNDA.n4812 GNDA.n4809 16.0005
R11193 GNDA.n4809 GNDA.n4808 16.0005
R11194 GNDA.n4808 GNDA.n4805 16.0005
R11195 GNDA.n4805 GNDA.n4804 16.0005
R11196 GNDA.n4804 GNDA.n4801 16.0005
R11197 GNDA.n4801 GNDA.n4800 16.0005
R11198 GNDA.n4800 GNDA.n4797 16.0005
R11199 GNDA.n4796 GNDA.n4793 16.0005
R11200 GNDA.n4793 GNDA.n4792 16.0005
R11201 GNDA.n4792 GNDA.n4789 16.0005
R11202 GNDA.n4789 GNDA.n4788 16.0005
R11203 GNDA.n4788 GNDA.n4785 16.0005
R11204 GNDA.n4785 GNDA.n4784 16.0005
R11205 GNDA.n4784 GNDA.n4781 16.0005
R11206 GNDA.n4781 GNDA.n4780 16.0005
R11207 GNDA.n2685 GNDA.n2684 16.0005
R11208 GNDA.n2688 GNDA.n2685 16.0005
R11209 GNDA.n2689 GNDA.n2688 16.0005
R11210 GNDA.n2692 GNDA.n2689 16.0005
R11211 GNDA.n2693 GNDA.n2692 16.0005
R11212 GNDA.n2696 GNDA.n2693 16.0005
R11213 GNDA.n2698 GNDA.n2696 16.0005
R11214 GNDA.n2699 GNDA.n2698 16.0005
R11215 GNDA.n2681 GNDA.n2680 16.0005
R11216 GNDA.n2680 GNDA.n2677 16.0005
R11217 GNDA.n2677 GNDA.n2676 16.0005
R11218 GNDA.n2676 GNDA.n2673 16.0005
R11219 GNDA.n2673 GNDA.n2672 16.0005
R11220 GNDA.n2672 GNDA.n2669 16.0005
R11221 GNDA.n2669 GNDA.n2668 16.0005
R11222 GNDA.n2668 GNDA.n2665 16.0005
R11223 GNDA.n2664 GNDA.n2661 16.0005
R11224 GNDA.n2661 GNDA.n2660 16.0005
R11225 GNDA.n2660 GNDA.n2657 16.0005
R11226 GNDA.n2657 GNDA.n2656 16.0005
R11227 GNDA.n2656 GNDA.n2653 16.0005
R11228 GNDA.n2653 GNDA.n2652 16.0005
R11229 GNDA.n2652 GNDA.n2649 16.0005
R11230 GNDA.n2649 GNDA.n2625 16.0005
R11231 GNDA.n4969 GNDA.n4956 16.0005
R11232 GNDA.n4969 GNDA.n4968 16.0005
R11233 GNDA.n4968 GNDA.n4967 16.0005
R11234 GNDA.n4967 GNDA.n4964 16.0005
R11235 GNDA.n4964 GNDA.n4963 16.0005
R11236 GNDA.n4963 GNDA.n4960 16.0005
R11237 GNDA.n4960 GNDA.n4959 16.0005
R11238 GNDA.n4959 GNDA.n4871 16.0005
R11239 GNDA.n4955 GNDA.n4953 16.0005
R11240 GNDA.n4953 GNDA.n4950 16.0005
R11241 GNDA.n4950 GNDA.n4949 16.0005
R11242 GNDA.n4949 GNDA.n4946 16.0005
R11243 GNDA.n4946 GNDA.n4945 16.0005
R11244 GNDA.n4945 GNDA.n4942 16.0005
R11245 GNDA.n4942 GNDA.n4941 16.0005
R11246 GNDA.n4941 GNDA.n4938 16.0005
R11247 GNDA.n4937 GNDA.n4934 16.0005
R11248 GNDA.n4934 GNDA.n4933 16.0005
R11249 GNDA.n4933 GNDA.n4930 16.0005
R11250 GNDA.n4930 GNDA.n4929 16.0005
R11251 GNDA.n4929 GNDA.n4926 16.0005
R11252 GNDA.n4926 GNDA.n4925 16.0005
R11253 GNDA.n4925 GNDA.n4922 16.0005
R11254 GNDA.n4922 GNDA.n4921 16.0005
R11255 GNDA.n5248 GNDA.n5235 16.0005
R11256 GNDA.n5248 GNDA.n5247 16.0005
R11257 GNDA.n5247 GNDA.n5246 16.0005
R11258 GNDA.n5246 GNDA.n5243 16.0005
R11259 GNDA.n5243 GNDA.n5242 16.0005
R11260 GNDA.n5242 GNDA.n5239 16.0005
R11261 GNDA.n5239 GNDA.n5238 16.0005
R11262 GNDA.n5238 GNDA.n57 16.0005
R11263 GNDA.n5234 GNDA.n5232 16.0005
R11264 GNDA.n5232 GNDA.n5229 16.0005
R11265 GNDA.n5229 GNDA.n5228 16.0005
R11266 GNDA.n5228 GNDA.n5225 16.0005
R11267 GNDA.n5225 GNDA.n5224 16.0005
R11268 GNDA.n5224 GNDA.n5221 16.0005
R11269 GNDA.n5221 GNDA.n5220 16.0005
R11270 GNDA.n5220 GNDA.n5217 16.0005
R11271 GNDA.n5216 GNDA.n5213 16.0005
R11272 GNDA.n5213 GNDA.n5212 16.0005
R11273 GNDA.n5212 GNDA.n5209 16.0005
R11274 GNDA.n5209 GNDA.n5208 16.0005
R11275 GNDA.n5208 GNDA.n5205 16.0005
R11276 GNDA.n5205 GNDA.n5204 16.0005
R11277 GNDA.n5204 GNDA.n5201 16.0005
R11278 GNDA.n5201 GNDA.n5200 16.0005
R11279 GNDA.n2470 GNDA.n2257 16.0005
R11280 GNDA.n2476 GNDA.n2257 16.0005
R11281 GNDA.n2477 GNDA.n2476 16.0005
R11282 GNDA.n2478 GNDA.n2477 16.0005
R11283 GNDA.n2478 GNDA.n2255 16.0005
R11284 GNDA.n2484 GNDA.n2255 16.0005
R11285 GNDA.n2485 GNDA.n2484 16.0005
R11286 GNDA.n2486 GNDA.n2485 16.0005
R11287 GNDA.n2469 GNDA.n2468 16.0005
R11288 GNDA.n2468 GNDA.n2259 16.0005
R11289 GNDA.n2462 GNDA.n2259 16.0005
R11290 GNDA.n2462 GNDA.n2461 16.0005
R11291 GNDA.n2461 GNDA.n2460 16.0005
R11292 GNDA.n2460 GNDA.n2261 16.0005
R11293 GNDA.n2454 GNDA.n2261 16.0005
R11294 GNDA.n2454 GNDA.n2453 16.0005
R11295 GNDA.n2452 GNDA.n2263 16.0005
R11296 GNDA.n2446 GNDA.n2263 16.0005
R11297 GNDA.n2446 GNDA.n2445 16.0005
R11298 GNDA.n2445 GNDA.n2444 16.0005
R11299 GNDA.n2444 GNDA.n2265 16.0005
R11300 GNDA.n2439 GNDA.n2265 16.0005
R11301 GNDA.n2439 GNDA.n2438 16.0005
R11302 GNDA.n2438 GNDA.n2437 16.0005
R11303 GNDA.n5155 GNDA.n5154 16.0005
R11304 GNDA.n5158 GNDA.n5155 16.0005
R11305 GNDA.n5159 GNDA.n5158 16.0005
R11306 GNDA.n5162 GNDA.n5159 16.0005
R11307 GNDA.n5163 GNDA.n5162 16.0005
R11308 GNDA.n5166 GNDA.n5163 16.0005
R11309 GNDA.n5168 GNDA.n5166 16.0005
R11310 GNDA.n5169 GNDA.n5168 16.0005
R11311 GNDA.n5151 GNDA.n5150 16.0005
R11312 GNDA.n5150 GNDA.n5147 16.0005
R11313 GNDA.n5147 GNDA.n5146 16.0005
R11314 GNDA.n5146 GNDA.n5143 16.0005
R11315 GNDA.n5143 GNDA.n5142 16.0005
R11316 GNDA.n5142 GNDA.n5139 16.0005
R11317 GNDA.n5139 GNDA.n5138 16.0005
R11318 GNDA.n5138 GNDA.n5135 16.0005
R11319 GNDA.n5134 GNDA.n5131 16.0005
R11320 GNDA.n5131 GNDA.n5130 16.0005
R11321 GNDA.n5130 GNDA.n5127 16.0005
R11322 GNDA.n5127 GNDA.n5126 16.0005
R11323 GNDA.n5126 GNDA.n5123 16.0005
R11324 GNDA.n5123 GNDA.n5122 16.0005
R11325 GNDA.n5122 GNDA.n5119 16.0005
R11326 GNDA.n5119 GNDA.n5118 16.0005
R11327 GNDA.n1743 GNDA.t147 15.3505
R11328 GNDA.t45 GNDA.t257 15.0244
R11329 GNDA.t35 GNDA.t45 15.0244
R11330 GNDA.t19 GNDA.t107 15.0244
R11331 GNDA.t198 GNDA.t14 14.9259
R11332 GNDA.t150 GNDA.t253 14.9259
R11333 GNDA.t274 GNDA.t20 14.9259
R11334 GNDA.t122 GNDA.t252 14.9259
R11335 GNDA.t211 GNDA.t97 14.9259
R11336 GNDA.t23 GNDA.t28 14.9259
R11337 GNDA.t219 GNDA.t220 14.9259
R11338 GNDA.t251 GNDA.t156 14.9259
R11339 GNDA.n5267 GNDA.n26 14.555
R11340 GNDA.n4988 GNDA.n107 14.555
R11341 GNDA.n435 GNDA.n434 13.9533
R11342 GNDA.n3148 GNDA.n3147 13.9533
R11343 GNDA.t263 GNDA.t42 13.8109
R11344 GNDA.n3946 GNDA.n3945 13.5941
R11345 GNDA.n1737 GNDA.n1407 13.5941
R11346 GNDA.n3949 GNDA.n3948 13.5697
R11347 GNDA.n1403 GNDA.n1402 13.5697
R11348 GNDA.t253 GNDA.n3128 13.4333
R11349 GNDA.n3098 GNDA.t219 13.4333
R11350 GNDA.n2385 GNDA.n2302 12.8005
R11351 GNDA.n2389 GNDA.n2302 12.8005
R11352 GNDA.n2290 GNDA.n2289 12.8005
R11353 GNDA.n2294 GNDA.n2289 12.8005
R11354 GNDA.n4687 GNDA.n357 12.8005
R11355 GNDA.n4687 GNDA.n4686 12.8005
R11356 GNDA.n3859 GNDA.t131 12.6791
R11357 GNDA.n4620 GNDA.t87 12.6791
R11358 GNDA.n1748 GNDA.t62 12.6791
R11359 GNDA.n3154 GNDA.t56 12.6791
R11360 GNDA.t143 GNDA.n2426 12.0196
R11361 GNDA.n3087 GNDA.t145 12.0196
R11362 GNDA.n2997 GNDA.t261 12.0196
R11363 GNDA.n2871 GNDA.n2868 11.6369
R11364 GNDA.n2874 GNDA.n2871 11.6369
R11365 GNDA.n2886 GNDA.n2874 11.6369
R11366 GNDA.n2886 GNDA.n2885 11.6369
R11367 GNDA.n2885 GNDA.n2884 11.6369
R11368 GNDA.n2884 GNDA.n2875 11.6369
R11369 GNDA.n2878 GNDA.n2875 11.6369
R11370 GNDA.n2878 GNDA.n2877 11.6369
R11371 GNDA.n2877 GNDA.n692 11.6369
R11372 GNDA.n3041 GNDA.n692 11.6369
R11373 GNDA.n2910 GNDA.n2860 11.6369
R11374 GNDA.n2910 GNDA.n2909 11.6369
R11375 GNDA.n2909 GNDA.n2908 11.6369
R11376 GNDA.n2908 GNDA.n2862 11.6369
R11377 GNDA.n2903 GNDA.n2862 11.6369
R11378 GNDA.n2903 GNDA.n2902 11.6369
R11379 GNDA.n2902 GNDA.n2901 11.6369
R11380 GNDA.n2901 GNDA.n2865 11.6369
R11381 GNDA.n2896 GNDA.n2865 11.6369
R11382 GNDA.n2896 GNDA.n2895 11.6369
R11383 GNDA.n2895 GNDA.n2894 11.6369
R11384 GNDA.n2938 GNDA.n2565 11.6369
R11385 GNDA.n2938 GNDA.n2937 11.6369
R11386 GNDA.n2937 GNDA.n2936 11.6369
R11387 GNDA.n2936 GNDA.n2567 11.6369
R11388 GNDA.n2931 GNDA.n2567 11.6369
R11389 GNDA.n2931 GNDA.n2930 11.6369
R11390 GNDA.n2930 GNDA.n2929 11.6369
R11391 GNDA.n2929 GNDA.n2570 11.6369
R11392 GNDA.n2924 GNDA.n2570 11.6369
R11393 GNDA.n2924 GNDA.n2923 11.6369
R11394 GNDA.n2923 GNDA.n2922 11.6369
R11395 GNDA.n2617 GNDA.n2613 11.6369
R11396 GNDA.n2758 GNDA.n2617 11.6369
R11397 GNDA.n2758 GNDA.n2757 11.6369
R11398 GNDA.n2757 GNDA.n2756 11.6369
R11399 GNDA.n2756 GNDA.n2618 11.6369
R11400 GNDA.n2751 GNDA.n2618 11.6369
R11401 GNDA.n2751 GNDA.n2750 11.6369
R11402 GNDA.n2750 GNDA.n2749 11.6369
R11403 GNDA.n2749 GNDA.n2620 11.6369
R11404 GNDA.n2743 GNDA.n2620 11.6369
R11405 GNDA.n2786 GNDA.n2785 11.6369
R11406 GNDA.n2785 GNDA.n2782 11.6369
R11407 GNDA.n2782 GNDA.n2781 11.6369
R11408 GNDA.n2781 GNDA.n2778 11.6369
R11409 GNDA.n2778 GNDA.n2777 11.6369
R11410 GNDA.n2777 GNDA.n2774 11.6369
R11411 GNDA.n2774 GNDA.n2773 11.6369
R11412 GNDA.n2773 GNDA.n2770 11.6369
R11413 GNDA.n2770 GNDA.n2769 11.6369
R11414 GNDA.n2769 GNDA.n2766 11.6369
R11415 GNDA.n2766 GNDA.n2765 11.6369
R11416 GNDA.n2589 GNDA.n132 11.6369
R11417 GNDA.n2592 GNDA.n2589 11.6369
R11418 GNDA.n2593 GNDA.n2592 11.6369
R11419 GNDA.n2596 GNDA.n2593 11.6369
R11420 GNDA.n2597 GNDA.n2596 11.6369
R11421 GNDA.n2600 GNDA.n2597 11.6369
R11422 GNDA.n2601 GNDA.n2600 11.6369
R11423 GNDA.n2604 GNDA.n2601 11.6369
R11424 GNDA.n2605 GNDA.n2604 11.6369
R11425 GNDA.n2608 GNDA.n2605 11.6369
R11426 GNDA.n2611 GNDA.n2608 11.6369
R11427 GNDA.n263 GNDA.n262 11.6369
R11428 GNDA.n266 GNDA.n263 11.6369
R11429 GNDA.n267 GNDA.n266 11.6369
R11430 GNDA.n270 GNDA.n267 11.6369
R11431 GNDA.n271 GNDA.n270 11.6369
R11432 GNDA.n274 GNDA.n271 11.6369
R11433 GNDA.n275 GNDA.n274 11.6369
R11434 GNDA.n277 GNDA.n275 11.6369
R11435 GNDA.n277 GNDA.n276 11.6369
R11436 GNDA.n276 GNDA.n228 11.6369
R11437 GNDA.n259 GNDA.n258 11.6369
R11438 GNDA.n258 GNDA.n255 11.6369
R11439 GNDA.n255 GNDA.n254 11.6369
R11440 GNDA.n254 GNDA.n251 11.6369
R11441 GNDA.n251 GNDA.n250 11.6369
R11442 GNDA.n250 GNDA.n247 11.6369
R11443 GNDA.n247 GNDA.n246 11.6369
R11444 GNDA.n246 GNDA.n243 11.6369
R11445 GNDA.n243 GNDA.n242 11.6369
R11446 GNDA.n242 GNDA.n131 11.6369
R11447 GNDA.n5084 GNDA.n131 11.6369
R11448 GNDA.n4864 GNDA.n4863 11.6369
R11449 GNDA.n4863 GNDA.n4862 11.6369
R11450 GNDA.n4862 GNDA.n4861 11.6369
R11451 GNDA.n4861 GNDA.n4859 11.6369
R11452 GNDA.n4859 GNDA.n4856 11.6369
R11453 GNDA.n4856 GNDA.n4855 11.6369
R11454 GNDA.n4855 GNDA.n4852 11.6369
R11455 GNDA.n4852 GNDA.n4851 11.6369
R11456 GNDA.n4851 GNDA.n4848 11.6369
R11457 GNDA.n4848 GNDA.n4847 11.6369
R11458 GNDA.n4726 GNDA.n4725 11.6369
R11459 GNDA.n4725 GNDA.n290 11.6369
R11460 GNDA.n4719 GNDA.n290 11.6369
R11461 GNDA.n4719 GNDA.n4718 11.6369
R11462 GNDA.n4718 GNDA.n4717 11.6369
R11463 GNDA.n4717 GNDA.n294 11.6369
R11464 GNDA.n4711 GNDA.n294 11.6369
R11465 GNDA.n4711 GNDA.n4710 11.6369
R11466 GNDA.n4710 GNDA.n4709 11.6369
R11467 GNDA.n4709 GNDA.n298 11.6369
R11468 GNDA.n4703 GNDA.n298 11.6369
R11469 GNDA.n2539 GNDA.n2538 11.6369
R11470 GNDA.n2538 GNDA.n2535 11.6369
R11471 GNDA.n2535 GNDA.n2534 11.6369
R11472 GNDA.n2534 GNDA.n2531 11.6369
R11473 GNDA.n2531 GNDA.n2530 11.6369
R11474 GNDA.n2530 GNDA.n2527 11.6369
R11475 GNDA.n2527 GNDA.n2526 11.6369
R11476 GNDA.n2526 GNDA.n2523 11.6369
R11477 GNDA.n2523 GNDA.n2522 11.6369
R11478 GNDA.n2522 GNDA.n2519 11.6369
R11479 GNDA.n2540 GNDA.n833 11.6369
R11480 GNDA.n2546 GNDA.n833 11.6369
R11481 GNDA.n2547 GNDA.n2546 11.6369
R11482 GNDA.n2548 GNDA.n2547 11.6369
R11483 GNDA.n2548 GNDA.n831 11.6369
R11484 GNDA.n2554 GNDA.n831 11.6369
R11485 GNDA.n2555 GNDA.n2554 11.6369
R11486 GNDA.n2556 GNDA.n2555 11.6369
R11487 GNDA.n2556 GNDA.n829 11.6369
R11488 GNDA.n2562 GNDA.n829 11.6369
R11489 GNDA.n2563 GNDA.n2562 11.6369
R11490 GNDA.n4645 GNDA.n4644 11.6369
R11491 GNDA.n4644 GNDA.n4643 11.6369
R11492 GNDA.n4643 GNDA.n426 11.6369
R11493 GNDA.n4637 GNDA.n426 11.6369
R11494 GNDA.n4637 GNDA.n4636 11.6369
R11495 GNDA.n4636 GNDA.n92 11.6369
R11496 GNDA.n5091 GNDA.n92 11.6369
R11497 GNDA.n5092 GNDA.n5091 11.6369
R11498 GNDA.n5094 GNDA.n5092 11.6369
R11499 GNDA.n5094 GNDA.n5093 11.6369
R11500 GNDA.n4669 GNDA.n4668 11.6369
R11501 GNDA.n4668 GNDA.n4667 11.6369
R11502 GNDA.n4667 GNDA.n414 11.6369
R11503 GNDA.n4661 GNDA.n414 11.6369
R11504 GNDA.n4661 GNDA.n4660 11.6369
R11505 GNDA.n4660 GNDA.n4659 11.6369
R11506 GNDA.n4659 GNDA.n418 11.6369
R11507 GNDA.n4653 GNDA.n418 11.6369
R11508 GNDA.n4653 GNDA.n4652 11.6369
R11509 GNDA.n4652 GNDA.n4651 11.6369
R11510 GNDA.n4651 GNDA.n422 11.6369
R11511 GNDA.n4701 GNDA.n303 11.6369
R11512 GNDA.n4695 GNDA.n303 11.6369
R11513 GNDA.n4695 GNDA.n4694 11.6369
R11514 GNDA.n4694 GNDA.n4693 11.6369
R11515 GNDA.n4693 GNDA.n353 11.6369
R11516 GNDA.n4684 GNDA.n360 11.6369
R11517 GNDA.n364 GNDA.n360 11.6369
R11518 GNDA.n4677 GNDA.n364 11.6369
R11519 GNDA.n4677 GNDA.n4676 11.6369
R11520 GNDA.n4676 GNDA.n4675 11.6369
R11521 GNDA.t32 GNDA.t26 11.4882
R11522 GNDA.t45 GNDA.n99 11.3072
R11523 GNDA.n1322 GNDA.n1321 11.245
R11524 GNDA.n3143 GNDA.n3142 11.245
R11525 GNDA.t158 GNDA.t183 11.0892
R11526 GNDA.t171 GNDA.t30 11.0892
R11527 GNDA.t279 GNDA.t15 11.0892
R11528 GNDA.t214 GNDA.t163 11.0892
R11529 GNDA.n3051 GNDA.n3050 10.9846
R11530 GNDA.n2243 GNDA.n2242 10.87
R11531 GNDA.n2511 GNDA.n2510 10.87
R11532 GNDA.n2509 GNDA.n2502 10.87
R11533 GNDA.n2318 GNDA.n676 10.87
R11534 GNDA.n3060 GNDA.n3059 10.87
R11535 GNDA.n3055 GNDA.n680 10.87
R11536 GNDA.n3054 GNDA.n681 10.87
R11537 GNDA.n636 GNDA.n543 10.5474
R11538 GNDA.n638 GNDA.n586 10.5474
R11539 GNDA.n3129 GNDA.t198 10.4483
R11540 GNDA.n3129 GNDA.t156 10.4483
R11541 GNDA.t148 GNDA.t204 9.90372
R11542 GNDA.t147 GNDA.t40 9.90372
R11543 GNDA.n2240 GNDA.t210 9.66779
R11544 GNDA.n1340 GNDA.t216 9.6005
R11545 GNDA.n1340 GNDA.t2 9.6005
R11546 GNDA.n3123 GNDA.t275 9.6005
R11547 GNDA.n3123 GNDA.t123 9.6005
R11548 GNDA.n3121 GNDA.t199 9.6005
R11549 GNDA.n3121 GNDA.t151 9.6005
R11550 GNDA.n3119 GNDA.t39 9.6005
R11551 GNDA.n3119 GNDA.t197 9.6005
R11552 GNDA.n3117 GNDA.t34 9.6005
R11553 GNDA.n3117 GNDA.t153 9.6005
R11554 GNDA.n3115 GNDA.t169 9.6005
R11555 GNDA.n3115 GNDA.t280 9.6005
R11556 GNDA.n3113 GNDA.t277 9.6005
R11557 GNDA.n3113 GNDA.t224 9.6005
R11558 GNDA.n3111 GNDA.t205 9.6005
R11559 GNDA.n3111 GNDA.t272 9.6005
R11560 GNDA.n3109 GNDA.t155 9.6005
R11561 GNDA.n3109 GNDA.t273 9.6005
R11562 GNDA.n3107 GNDA.t154 9.6005
R11563 GNDA.n3107 GNDA.t281 9.6005
R11564 GNDA.n3105 GNDA.t271 9.6005
R11565 GNDA.n3105 GNDA.t286 9.6005
R11566 GNDA.n3103 GNDA.t221 9.6005
R11567 GNDA.n3103 GNDA.t157 9.6005
R11568 GNDA.n3101 GNDA.t98 9.6005
R11569 GNDA.n3101 GNDA.t29 9.6005
R11570 GNDA.n3015 GNDA.t240 9.6005
R11571 GNDA.n705 GNDA.t244 9.6005
R11572 GNDA.n2397 GNDA.t247 9.6005
R11573 GNDA.n2406 GNDA.t249 9.6005
R11574 GNDA.n2385 GNDA.n2300 9.36264
R11575 GNDA.n2290 GNDA.n2287 9.36264
R11576 GNDA.n2207 GNDA.n357 9.36264
R11577 GNDA.n2302 GNDA.n2301 9.3005
R11578 GNDA.n2390 GNDA.n2389 9.3005
R11579 GNDA.n2289 GNDA.n2288 9.3005
R11580 GNDA.n2295 GNDA.n2294 9.3005
R11581 GNDA.n4687 GNDA.n358 9.3005
R11582 GNDA.n4686 GNDA.n359 9.3005
R11583 GNDA.t141 GNDA.t206 8.87147
R11584 GNDA.t142 GNDA.t200 8.87147
R11585 GNDA.n3032 GNDA.n3030 8.62751
R11586 GNDA.n5174 GNDA.n26 8.60107
R11587 GNDA.n161 GNDA.n107 8.60107
R11588 GNDA.n2515 GNDA.t93 8.01325
R11589 GNDA.n2425 GNDA.t21 8.01325
R11590 GNDA.t217 GNDA.n3064 8.01325
R11591 GNDA.t228 GNDA.n2998 8.01325
R11592 GNDA.n3127 GNDA.t234 7.46319
R11593 GNDA.n3099 GNDA.t162 7.46319
R11594 GNDA.n2499 GNDA.t13 7.01165
R11595 GNDA.n2429 GNDA.t256 7.01165
R11596 GNDA.n2922 GNDA.n2824 6.72373
R11597 GNDA.n2612 GNDA.n2611 6.72373
R11598 GNDA.n5084 GNDA.n5083 6.72373
R11599 GNDA.n4703 GNDA.n4702 6.72373
R11600 GNDA.n2564 GNDA.n2563 6.72373
R11601 GNDA.n4675 GNDA.n365 6.72373
R11602 GNDA.n2860 GNDA.n2824 6.20656
R11603 GNDA.n2565 GNDA.n2564 6.20656
R11604 GNDA.n2786 GNDA.n2612 6.20656
R11605 GNDA.n5083 GNDA.n132 6.20656
R11606 GNDA.n4669 GNDA.n365 6.20656
R11607 GNDA.n4702 GNDA.n4701 6.20656
R11608 GNDA.n4685 GNDA.n353 6.07727
R11609 GNDA.t45 GNDA.t6 6.01006
R11610 GNDA.n2407 GNDA.n2398 5.81868
R11611 GNDA.n2405 GNDA.n2398 5.81868
R11612 GNDA.n4685 GNDA.n4684 5.5601
R11613 GNDA.n3044 GNDA.n690 5.51161
R11614 GNDA.n2380 GNDA.n2378 5.51161
R11615 GNDA.n4995 GNDA.n186 5.51161
R11616 GNDA.n4780 GNDA.n4750 5.51161
R11617 GNDA.n2737 GNDA.n2625 5.51161
R11618 GNDA.n4921 GNDA.n4899 5.51161
R11619 GNDA.n5200 GNDA.n5178 5.51161
R11620 GNDA.n2437 GNDA.n2268 5.51161
R11621 GNDA.n5118 GNDA.n5104 5.51161
R11622 GNDA.n3095 GNDA.t282 5.38323
R11623 GNDA.n3043 GNDA.n3042 5.1717
R11624 GNDA.n2742 GNDA.n2738 5.1717
R11625 GNDA.n5103 GNDA.n87 5.1717
R11626 GNDA.t201 GNDA.t139 5.00847
R11627 GNDA.n2409 GNDA.t257 5.00847
R11628 GNDA.t45 GNDA.t49 5.00847
R11629 GNDA.n3021 GNDA.t35 5.00847
R11630 GNDA.t9 GNDA.t17 5.00847
R11631 GNDA.n4985 GNDA.n4870 4.9157
R11632 GNDA.n4844 GNDA.n4841 4.9157
R11633 GNDA.n2518 GNDA.n2517 4.9157
R11634 GNDA.n3102 GNDA.n641 4.67238
R11635 GNDA.n3125 GNDA.n3124 4.67238
R11636 GNDA.n3133 GNDA.n3131 4.65331
R11637 GNDA.n632 GNDA.n627 4.65331
R11638 GNDA.n1304 GNDA.n1289 4.5005
R11639 GNDA.n1303 GNDA.n1302 4.5005
R11640 GNDA.n1304 GNDA.n1303 4.5005
R11641 GNDA.n1280 GNDA.n1279 4.5005
R11642 GNDA.n1283 GNDA.n1282 4.5005
R11643 GNDA.n1286 GNDA.n1285 4.5005
R11644 GNDA.n1338 GNDA.n1275 4.5005
R11645 GNDA.n1337 GNDA.n1336 4.5005
R11646 GNDA.n1338 GNDA.n1337 4.5005
R11647 GNDA.n1346 GNDA.n1345 4.5005
R11648 GNDA.n1352 GNDA.n1351 4.5005
R11649 GNDA.n1355 GNDA.n628 4.5005
R11650 GNDA.n1356 GNDA.n1355 4.5005
R11651 GNDA.n1357 GNDA.n1356 4.5005
R11652 GNDA.n1364 GNDA.n1260 4.5005
R11653 GNDA.n1363 GNDA.n1362 4.5005
R11654 GNDA.n1364 GNDA.n1363 4.5005
R11655 GNDA.n1380 GNDA.n1379 4.5005
R11656 GNDA.n1386 GNDA.n1256 4.5005
R11657 GNDA.n1387 GNDA.n1255 4.5005
R11658 GNDA.n1387 GNDA.n1386 4.5005
R11659 GNDA.n1299 GNDA.n1298 4.5005
R11660 GNDA.n1299 GNDA.n436 4.5005
R11661 GNDA.n1296 GNDA.n436 4.5005
R11662 GNDA.n3706 GNDA.n3705 4.5005
R11663 GNDA.n3704 GNDA.n3626 4.5005
R11664 GNDA.n3703 GNDA.n3702 4.5005
R11665 GNDA.n3701 GNDA.n3631 4.5005
R11666 GNDA.n3700 GNDA.n3699 4.5005
R11667 GNDA.n3698 GNDA.n3632 4.5005
R11668 GNDA.n3697 GNDA.n3696 4.5005
R11669 GNDA.n3695 GNDA.n3639 4.5005
R11670 GNDA.n3694 GNDA.n3693 4.5005
R11671 GNDA.n3692 GNDA.n3640 4.5005
R11672 GNDA.n3691 GNDA.n3690 4.5005
R11673 GNDA.n3689 GNDA.n3647 4.5005
R11674 GNDA.n3688 GNDA.n3687 4.5005
R11675 GNDA.n3686 GNDA.n3648 4.5005
R11676 GNDA.n3685 GNDA.n3684 4.5005
R11677 GNDA.n3683 GNDA.n3655 4.5005
R11678 GNDA.n3682 GNDA.n3681 4.5005
R11679 GNDA.n3680 GNDA.n3656 4.5005
R11680 GNDA.n3679 GNDA.n3678 4.5005
R11681 GNDA.n3677 GNDA.n3663 4.5005
R11682 GNDA.n3676 GNDA.n3675 4.5005
R11683 GNDA.n3674 GNDA.n3664 4.5005
R11684 GNDA.n3385 GNDA.n3384 4.5005
R11685 GNDA.n591 GNDA.n590 4.5005
R11686 GNDA.n3330 GNDA.n3329 4.5005
R11687 GNDA.n3334 GNDA.n3331 4.5005
R11688 GNDA.n3335 GNDA.n3328 4.5005
R11689 GNDA.n3339 GNDA.n3338 4.5005
R11690 GNDA.n3340 GNDA.n3327 4.5005
R11691 GNDA.n3344 GNDA.n3341 4.5005
R11692 GNDA.n3345 GNDA.n3326 4.5005
R11693 GNDA.n3349 GNDA.n3348 4.5005
R11694 GNDA.n3350 GNDA.n3325 4.5005
R11695 GNDA.n3354 GNDA.n3351 4.5005
R11696 GNDA.n3355 GNDA.n3324 4.5005
R11697 GNDA.n3359 GNDA.n3358 4.5005
R11698 GNDA.n3360 GNDA.n3323 4.5005
R11699 GNDA.n3364 GNDA.n3361 4.5005
R11700 GNDA.n3365 GNDA.n3322 4.5005
R11701 GNDA.n3369 GNDA.n3368 4.5005
R11702 GNDA.n3370 GNDA.n3321 4.5005
R11703 GNDA.n3374 GNDA.n3371 4.5005
R11704 GNDA.n3375 GNDA.n3320 4.5005
R11705 GNDA.n3379 GNDA.n3378 4.5005
R11706 GNDA.n4582 GNDA.n4581 4.5005
R11707 GNDA.n475 GNDA.n474 4.5005
R11708 GNDA.n4527 GNDA.n4526 4.5005
R11709 GNDA.n4531 GNDA.n4528 4.5005
R11710 GNDA.n4532 GNDA.n4525 4.5005
R11711 GNDA.n4536 GNDA.n4535 4.5005
R11712 GNDA.n4537 GNDA.n4524 4.5005
R11713 GNDA.n4541 GNDA.n4538 4.5005
R11714 GNDA.n4542 GNDA.n4523 4.5005
R11715 GNDA.n4546 GNDA.n4545 4.5005
R11716 GNDA.n4547 GNDA.n4522 4.5005
R11717 GNDA.n4551 GNDA.n4548 4.5005
R11718 GNDA.n4552 GNDA.n4521 4.5005
R11719 GNDA.n4556 GNDA.n4555 4.5005
R11720 GNDA.n4557 GNDA.n4520 4.5005
R11721 GNDA.n4561 GNDA.n4558 4.5005
R11722 GNDA.n4562 GNDA.n4519 4.5005
R11723 GNDA.n4566 GNDA.n4565 4.5005
R11724 GNDA.n4567 GNDA.n4518 4.5005
R11725 GNDA.n4571 GNDA.n4568 4.5005
R11726 GNDA.n4572 GNDA.n4517 4.5005
R11727 GNDA.n4576 GNDA.n4575 4.5005
R11728 GNDA.n4447 GNDA.n4446 4.5005
R11729 GNDA.n4450 GNDA.n4449 4.5005
R11730 GNDA.n4451 GNDA.n4445 4.5005
R11731 GNDA.n4455 GNDA.n4452 4.5005
R11732 GNDA.n4456 GNDA.n4444 4.5005
R11733 GNDA.n4460 GNDA.n4459 4.5005
R11734 GNDA.n4461 GNDA.n4443 4.5005
R11735 GNDA.n4465 GNDA.n4462 4.5005
R11736 GNDA.n4466 GNDA.n4442 4.5005
R11737 GNDA.n4470 GNDA.n4469 4.5005
R11738 GNDA.n4471 GNDA.n4441 4.5005
R11739 GNDA.n4475 GNDA.n4472 4.5005
R11740 GNDA.n4476 GNDA.n4440 4.5005
R11741 GNDA.n4480 GNDA.n4479 4.5005
R11742 GNDA.n4481 GNDA.n4439 4.5005
R11743 GNDA.n4485 GNDA.n4482 4.5005
R11744 GNDA.n4486 GNDA.n4438 4.5005
R11745 GNDA.n4490 GNDA.n4489 4.5005
R11746 GNDA.n4491 GNDA.n4437 4.5005
R11747 GNDA.n4495 GNDA.n4492 4.5005
R11748 GNDA.n4496 GNDA.n4436 4.5005
R11749 GNDA.n4500 GNDA.n4499 4.5005
R11750 GNDA.n4365 GNDA.n4364 4.5005
R11751 GNDA.n4368 GNDA.n4367 4.5005
R11752 GNDA.n4369 GNDA.n4363 4.5005
R11753 GNDA.n4373 GNDA.n4370 4.5005
R11754 GNDA.n4374 GNDA.n4362 4.5005
R11755 GNDA.n4378 GNDA.n4377 4.5005
R11756 GNDA.n4379 GNDA.n4361 4.5005
R11757 GNDA.n4383 GNDA.n4380 4.5005
R11758 GNDA.n4384 GNDA.n4360 4.5005
R11759 GNDA.n4388 GNDA.n4387 4.5005
R11760 GNDA.n4389 GNDA.n4359 4.5005
R11761 GNDA.n4393 GNDA.n4390 4.5005
R11762 GNDA.n4394 GNDA.n4358 4.5005
R11763 GNDA.n4398 GNDA.n4397 4.5005
R11764 GNDA.n4399 GNDA.n4357 4.5005
R11765 GNDA.n4403 GNDA.n4400 4.5005
R11766 GNDA.n4404 GNDA.n4356 4.5005
R11767 GNDA.n4408 GNDA.n4407 4.5005
R11768 GNDA.n4409 GNDA.n4355 4.5005
R11769 GNDA.n4413 GNDA.n4410 4.5005
R11770 GNDA.n4414 GNDA.n4354 4.5005
R11771 GNDA.n4418 GNDA.n4417 4.5005
R11772 GNDA.n4283 GNDA.n4282 4.5005
R11773 GNDA.n4286 GNDA.n4285 4.5005
R11774 GNDA.n4287 GNDA.n4281 4.5005
R11775 GNDA.n4291 GNDA.n4288 4.5005
R11776 GNDA.n4292 GNDA.n4280 4.5005
R11777 GNDA.n4296 GNDA.n4295 4.5005
R11778 GNDA.n4297 GNDA.n4279 4.5005
R11779 GNDA.n4301 GNDA.n4298 4.5005
R11780 GNDA.n4302 GNDA.n4278 4.5005
R11781 GNDA.n4306 GNDA.n4305 4.5005
R11782 GNDA.n4307 GNDA.n4277 4.5005
R11783 GNDA.n4311 GNDA.n4308 4.5005
R11784 GNDA.n4312 GNDA.n4276 4.5005
R11785 GNDA.n4316 GNDA.n4315 4.5005
R11786 GNDA.n4317 GNDA.n4275 4.5005
R11787 GNDA.n4321 GNDA.n4318 4.5005
R11788 GNDA.n4322 GNDA.n4274 4.5005
R11789 GNDA.n4326 GNDA.n4325 4.5005
R11790 GNDA.n4327 GNDA.n4273 4.5005
R11791 GNDA.n4331 GNDA.n4328 4.5005
R11792 GNDA.n4332 GNDA.n4272 4.5005
R11793 GNDA.n4336 GNDA.n4335 4.5005
R11794 GNDA.n4201 GNDA.n4200 4.5005
R11795 GNDA.n4204 GNDA.n4203 4.5005
R11796 GNDA.n4205 GNDA.n4199 4.5005
R11797 GNDA.n4209 GNDA.n4206 4.5005
R11798 GNDA.n4210 GNDA.n4198 4.5005
R11799 GNDA.n4214 GNDA.n4213 4.5005
R11800 GNDA.n4215 GNDA.n4197 4.5005
R11801 GNDA.n4219 GNDA.n4216 4.5005
R11802 GNDA.n4220 GNDA.n4196 4.5005
R11803 GNDA.n4224 GNDA.n4223 4.5005
R11804 GNDA.n4225 GNDA.n4195 4.5005
R11805 GNDA.n4229 GNDA.n4226 4.5005
R11806 GNDA.n4230 GNDA.n4194 4.5005
R11807 GNDA.n4234 GNDA.n4233 4.5005
R11808 GNDA.n4235 GNDA.n4193 4.5005
R11809 GNDA.n4239 GNDA.n4236 4.5005
R11810 GNDA.n4240 GNDA.n4192 4.5005
R11811 GNDA.n4244 GNDA.n4243 4.5005
R11812 GNDA.n4245 GNDA.n4191 4.5005
R11813 GNDA.n4249 GNDA.n4246 4.5005
R11814 GNDA.n4250 GNDA.n4190 4.5005
R11815 GNDA.n4254 GNDA.n4253 4.5005
R11816 GNDA.n3955 GNDA.n3954 4.5005
R11817 GNDA.n3958 GNDA.n3957 4.5005
R11818 GNDA.n3959 GNDA.n501 4.5005
R11819 GNDA.n3963 GNDA.n3960 4.5005
R11820 GNDA.n3964 GNDA.n500 4.5005
R11821 GNDA.n3968 GNDA.n3967 4.5005
R11822 GNDA.n3969 GNDA.n499 4.5005
R11823 GNDA.n3973 GNDA.n3970 4.5005
R11824 GNDA.n3974 GNDA.n498 4.5005
R11825 GNDA.n3978 GNDA.n3977 4.5005
R11826 GNDA.n3979 GNDA.n497 4.5005
R11827 GNDA.n3983 GNDA.n3980 4.5005
R11828 GNDA.n3984 GNDA.n496 4.5005
R11829 GNDA.n3988 GNDA.n3987 4.5005
R11830 GNDA.n3989 GNDA.n495 4.5005
R11831 GNDA.n3993 GNDA.n3990 4.5005
R11832 GNDA.n3994 GNDA.n494 4.5005
R11833 GNDA.n3998 GNDA.n3997 4.5005
R11834 GNDA.n3999 GNDA.n493 4.5005
R11835 GNDA.n4003 GNDA.n4000 4.5005
R11836 GNDA.n4004 GNDA.n492 4.5005
R11837 GNDA.n4008 GNDA.n4007 4.5005
R11838 GNDA.n4119 GNDA.n4118 4.5005
R11839 GNDA.n4122 GNDA.n4121 4.5005
R11840 GNDA.n4123 GNDA.n4117 4.5005
R11841 GNDA.n4127 GNDA.n4124 4.5005
R11842 GNDA.n4128 GNDA.n4116 4.5005
R11843 GNDA.n4132 GNDA.n4131 4.5005
R11844 GNDA.n4133 GNDA.n4115 4.5005
R11845 GNDA.n4137 GNDA.n4134 4.5005
R11846 GNDA.n4138 GNDA.n4114 4.5005
R11847 GNDA.n4142 GNDA.n4141 4.5005
R11848 GNDA.n4143 GNDA.n4113 4.5005
R11849 GNDA.n4147 GNDA.n4144 4.5005
R11850 GNDA.n4148 GNDA.n4112 4.5005
R11851 GNDA.n4152 GNDA.n4151 4.5005
R11852 GNDA.n4153 GNDA.n4111 4.5005
R11853 GNDA.n4157 GNDA.n4154 4.5005
R11854 GNDA.n4158 GNDA.n4110 4.5005
R11855 GNDA.n4162 GNDA.n4161 4.5005
R11856 GNDA.n4163 GNDA.n4109 4.5005
R11857 GNDA.n4167 GNDA.n4164 4.5005
R11858 GNDA.n4168 GNDA.n4108 4.5005
R11859 GNDA.n4172 GNDA.n4171 4.5005
R11860 GNDA.n4037 GNDA.n4036 4.5005
R11861 GNDA.n4040 GNDA.n4039 4.5005
R11862 GNDA.n4041 GNDA.n4035 4.5005
R11863 GNDA.n4045 GNDA.n4042 4.5005
R11864 GNDA.n4046 GNDA.n4034 4.5005
R11865 GNDA.n4050 GNDA.n4049 4.5005
R11866 GNDA.n4051 GNDA.n4033 4.5005
R11867 GNDA.n4055 GNDA.n4052 4.5005
R11868 GNDA.n4056 GNDA.n4032 4.5005
R11869 GNDA.n4060 GNDA.n4059 4.5005
R11870 GNDA.n4061 GNDA.n4031 4.5005
R11871 GNDA.n4065 GNDA.n4062 4.5005
R11872 GNDA.n4066 GNDA.n4030 4.5005
R11873 GNDA.n4070 GNDA.n4069 4.5005
R11874 GNDA.n4071 GNDA.n4029 4.5005
R11875 GNDA.n4075 GNDA.n4072 4.5005
R11876 GNDA.n4076 GNDA.n4028 4.5005
R11877 GNDA.n4080 GNDA.n4079 4.5005
R11878 GNDA.n4081 GNDA.n4027 4.5005
R11879 GNDA.n4085 GNDA.n4082 4.5005
R11880 GNDA.n4086 GNDA.n4026 4.5005
R11881 GNDA.n4090 GNDA.n4089 4.5005
R11882 GNDA.n3943 GNDA.n3942 4.5005
R11883 GNDA.n3864 GNDA.n3863 4.5005
R11884 GNDA.n3886 GNDA.n3865 4.5005
R11885 GNDA.n3887 GNDA.n3866 4.5005
R11886 GNDA.n3888 GNDA.n3867 4.5005
R11887 GNDA.n3889 GNDA.n3868 4.5005
R11888 GNDA.n3890 GNDA.n3869 4.5005
R11889 GNDA.n3891 GNDA.n3870 4.5005
R11890 GNDA.n3892 GNDA.n3871 4.5005
R11891 GNDA.n3893 GNDA.n3872 4.5005
R11892 GNDA.n3894 GNDA.n3873 4.5005
R11893 GNDA.n3895 GNDA.n3874 4.5005
R11894 GNDA.n3896 GNDA.n3875 4.5005
R11895 GNDA.n3897 GNDA.n3876 4.5005
R11896 GNDA.n3898 GNDA.n3877 4.5005
R11897 GNDA.n3899 GNDA.n3878 4.5005
R11898 GNDA.n3900 GNDA.n3879 4.5005
R11899 GNDA.n3901 GNDA.n3880 4.5005
R11900 GNDA.n3902 GNDA.n3881 4.5005
R11901 GNDA.n3903 GNDA.n3882 4.5005
R11902 GNDA.n3904 GNDA.n3883 4.5005
R11903 GNDA.n3905 GNDA.n3884 4.5005
R11904 GNDA.n1735 GNDA.n1734 4.5005
R11905 GNDA.n1409 GNDA.n1408 4.5005
R11906 GNDA.n1680 GNDA.n1679 4.5005
R11907 GNDA.n1684 GNDA.n1681 4.5005
R11908 GNDA.n1685 GNDA.n1678 4.5005
R11909 GNDA.n1689 GNDA.n1688 4.5005
R11910 GNDA.n1690 GNDA.n1677 4.5005
R11911 GNDA.n1694 GNDA.n1691 4.5005
R11912 GNDA.n1695 GNDA.n1676 4.5005
R11913 GNDA.n1699 GNDA.n1698 4.5005
R11914 GNDA.n1700 GNDA.n1675 4.5005
R11915 GNDA.n1704 GNDA.n1701 4.5005
R11916 GNDA.n1705 GNDA.n1674 4.5005
R11917 GNDA.n1709 GNDA.n1708 4.5005
R11918 GNDA.n1710 GNDA.n1673 4.5005
R11919 GNDA.n1714 GNDA.n1711 4.5005
R11920 GNDA.n1715 GNDA.n1672 4.5005
R11921 GNDA.n1719 GNDA.n1718 4.5005
R11922 GNDA.n1720 GNDA.n1671 4.5005
R11923 GNDA.n1724 GNDA.n1721 4.5005
R11924 GNDA.n1725 GNDA.n1670 4.5005
R11925 GNDA.n1729 GNDA.n1728 4.5005
R11926 GNDA.n3853 GNDA.n3852 4.5005
R11927 GNDA.n511 GNDA.n510 4.5005
R11928 GNDA.n3798 GNDA.n3797 4.5005
R11929 GNDA.n3802 GNDA.n3799 4.5005
R11930 GNDA.n3803 GNDA.n3796 4.5005
R11931 GNDA.n3807 GNDA.n3806 4.5005
R11932 GNDA.n3808 GNDA.n3795 4.5005
R11933 GNDA.n3812 GNDA.n3809 4.5005
R11934 GNDA.n3813 GNDA.n3794 4.5005
R11935 GNDA.n3817 GNDA.n3816 4.5005
R11936 GNDA.n3818 GNDA.n3793 4.5005
R11937 GNDA.n3822 GNDA.n3819 4.5005
R11938 GNDA.n3823 GNDA.n3792 4.5005
R11939 GNDA.n3827 GNDA.n3826 4.5005
R11940 GNDA.n3828 GNDA.n3791 4.5005
R11941 GNDA.n3832 GNDA.n3829 4.5005
R11942 GNDA.n3833 GNDA.n3790 4.5005
R11943 GNDA.n3837 GNDA.n3836 4.5005
R11944 GNDA.n3838 GNDA.n3789 4.5005
R11945 GNDA.n3842 GNDA.n3839 4.5005
R11946 GNDA.n3843 GNDA.n3788 4.5005
R11947 GNDA.n3847 GNDA.n3846 4.5005
R11948 GNDA.n3718 GNDA.n3717 4.5005
R11949 GNDA.n3721 GNDA.n3720 4.5005
R11950 GNDA.n3722 GNDA.n537 4.5005
R11951 GNDA.n3726 GNDA.n3723 4.5005
R11952 GNDA.n3727 GNDA.n536 4.5005
R11953 GNDA.n3731 GNDA.n3730 4.5005
R11954 GNDA.n3732 GNDA.n535 4.5005
R11955 GNDA.n3736 GNDA.n3733 4.5005
R11956 GNDA.n3737 GNDA.n534 4.5005
R11957 GNDA.n3741 GNDA.n3740 4.5005
R11958 GNDA.n3742 GNDA.n533 4.5005
R11959 GNDA.n3746 GNDA.n3743 4.5005
R11960 GNDA.n3747 GNDA.n532 4.5005
R11961 GNDA.n3751 GNDA.n3750 4.5005
R11962 GNDA.n3752 GNDA.n531 4.5005
R11963 GNDA.n3756 GNDA.n3753 4.5005
R11964 GNDA.n3757 GNDA.n530 4.5005
R11965 GNDA.n3761 GNDA.n3760 4.5005
R11966 GNDA.n3762 GNDA.n529 4.5005
R11967 GNDA.n3766 GNDA.n3763 4.5005
R11968 GNDA.n3767 GNDA.n528 4.5005
R11969 GNDA.n3771 GNDA.n3770 4.5005
R11970 GNDA.n3619 GNDA.n3618 4.5005
R11971 GNDA.n551 GNDA.n550 4.5005
R11972 GNDA.n3564 GNDA.n3563 4.5005
R11973 GNDA.n3568 GNDA.n3565 4.5005
R11974 GNDA.n3569 GNDA.n3562 4.5005
R11975 GNDA.n3573 GNDA.n3572 4.5005
R11976 GNDA.n3574 GNDA.n3561 4.5005
R11977 GNDA.n3578 GNDA.n3575 4.5005
R11978 GNDA.n3579 GNDA.n3560 4.5005
R11979 GNDA.n3583 GNDA.n3582 4.5005
R11980 GNDA.n3584 GNDA.n3559 4.5005
R11981 GNDA.n3588 GNDA.n3585 4.5005
R11982 GNDA.n3589 GNDA.n3558 4.5005
R11983 GNDA.n3593 GNDA.n3592 4.5005
R11984 GNDA.n3594 GNDA.n3557 4.5005
R11985 GNDA.n3598 GNDA.n3595 4.5005
R11986 GNDA.n3599 GNDA.n3556 4.5005
R11987 GNDA.n3603 GNDA.n3602 4.5005
R11988 GNDA.n3604 GNDA.n3555 4.5005
R11989 GNDA.n3608 GNDA.n3605 4.5005
R11990 GNDA.n3609 GNDA.n3554 4.5005
R11991 GNDA.n3613 GNDA.n3612 4.5005
R11992 GNDA.n3484 GNDA.n3483 4.5005
R11993 GNDA.n3487 GNDA.n3486 4.5005
R11994 GNDA.n3488 GNDA.n577 4.5005
R11995 GNDA.n3492 GNDA.n3489 4.5005
R11996 GNDA.n3493 GNDA.n576 4.5005
R11997 GNDA.n3497 GNDA.n3496 4.5005
R11998 GNDA.n3498 GNDA.n575 4.5005
R11999 GNDA.n3502 GNDA.n3499 4.5005
R12000 GNDA.n3503 GNDA.n574 4.5005
R12001 GNDA.n3507 GNDA.n3506 4.5005
R12002 GNDA.n3508 GNDA.n573 4.5005
R12003 GNDA.n3512 GNDA.n3509 4.5005
R12004 GNDA.n3513 GNDA.n572 4.5005
R12005 GNDA.n3517 GNDA.n3516 4.5005
R12006 GNDA.n3518 GNDA.n571 4.5005
R12007 GNDA.n3522 GNDA.n3519 4.5005
R12008 GNDA.n3523 GNDA.n570 4.5005
R12009 GNDA.n3527 GNDA.n3526 4.5005
R12010 GNDA.n3528 GNDA.n569 4.5005
R12011 GNDA.n3532 GNDA.n3529 4.5005
R12012 GNDA.n3533 GNDA.n568 4.5005
R12013 GNDA.n3537 GNDA.n3536 4.5005
R12014 GNDA.n3472 GNDA.n3471 4.5005
R12015 GNDA.n3393 GNDA.n3392 4.5005
R12016 GNDA.n3415 GNDA.n3394 4.5005
R12017 GNDA.n3416 GNDA.n3395 4.5005
R12018 GNDA.n3417 GNDA.n3396 4.5005
R12019 GNDA.n3418 GNDA.n3397 4.5005
R12020 GNDA.n3419 GNDA.n3398 4.5005
R12021 GNDA.n3420 GNDA.n3399 4.5005
R12022 GNDA.n3421 GNDA.n3400 4.5005
R12023 GNDA.n3422 GNDA.n3401 4.5005
R12024 GNDA.n3423 GNDA.n3402 4.5005
R12025 GNDA.n3424 GNDA.n3403 4.5005
R12026 GNDA.n3425 GNDA.n3404 4.5005
R12027 GNDA.n3426 GNDA.n3405 4.5005
R12028 GNDA.n3427 GNDA.n3406 4.5005
R12029 GNDA.n3428 GNDA.n3407 4.5005
R12030 GNDA.n3429 GNDA.n3408 4.5005
R12031 GNDA.n3430 GNDA.n3409 4.5005
R12032 GNDA.n3431 GNDA.n3410 4.5005
R12033 GNDA.n3432 GNDA.n3411 4.5005
R12034 GNDA.n3433 GNDA.n3412 4.5005
R12035 GNDA.n3434 GNDA.n3413 4.5005
R12036 GNDA.n3250 GNDA.n3249 4.5005
R12037 GNDA.n3253 GNDA.n3252 4.5005
R12038 GNDA.n3254 GNDA.n617 4.5005
R12039 GNDA.n3258 GNDA.n3255 4.5005
R12040 GNDA.n3259 GNDA.n616 4.5005
R12041 GNDA.n3263 GNDA.n3262 4.5005
R12042 GNDA.n3264 GNDA.n615 4.5005
R12043 GNDA.n3268 GNDA.n3265 4.5005
R12044 GNDA.n3269 GNDA.n614 4.5005
R12045 GNDA.n3273 GNDA.n3272 4.5005
R12046 GNDA.n3274 GNDA.n613 4.5005
R12047 GNDA.n3278 GNDA.n3275 4.5005
R12048 GNDA.n3279 GNDA.n612 4.5005
R12049 GNDA.n3283 GNDA.n3282 4.5005
R12050 GNDA.n3284 GNDA.n611 4.5005
R12051 GNDA.n3288 GNDA.n3285 4.5005
R12052 GNDA.n3289 GNDA.n610 4.5005
R12053 GNDA.n3293 GNDA.n3292 4.5005
R12054 GNDA.n3294 GNDA.n609 4.5005
R12055 GNDA.n3298 GNDA.n3295 4.5005
R12056 GNDA.n3299 GNDA.n608 4.5005
R12057 GNDA.n3303 GNDA.n3302 4.5005
R12058 GNDA.n3238 GNDA.n3237 4.5005
R12059 GNDA.n3159 GNDA.n3158 4.5005
R12060 GNDA.n3181 GNDA.n3160 4.5005
R12061 GNDA.n3182 GNDA.n3161 4.5005
R12062 GNDA.n3183 GNDA.n3162 4.5005
R12063 GNDA.n3184 GNDA.n3163 4.5005
R12064 GNDA.n3185 GNDA.n3164 4.5005
R12065 GNDA.n3186 GNDA.n3165 4.5005
R12066 GNDA.n3187 GNDA.n3166 4.5005
R12067 GNDA.n3188 GNDA.n3167 4.5005
R12068 GNDA.n3189 GNDA.n3168 4.5005
R12069 GNDA.n3190 GNDA.n3169 4.5005
R12070 GNDA.n3191 GNDA.n3170 4.5005
R12071 GNDA.n3192 GNDA.n3171 4.5005
R12072 GNDA.n3193 GNDA.n3172 4.5005
R12073 GNDA.n3194 GNDA.n3173 4.5005
R12074 GNDA.n3195 GNDA.n3174 4.5005
R12075 GNDA.n3196 GNDA.n3175 4.5005
R12076 GNDA.n3197 GNDA.n3176 4.5005
R12077 GNDA.n3198 GNDA.n3177 4.5005
R12078 GNDA.n3199 GNDA.n3178 4.5005
R12079 GNDA.n3200 GNDA.n3179 4.5005
R12080 GNDA.n1600 GNDA.n1599 4.5005
R12081 GNDA.n1603 GNDA.n1602 4.5005
R12082 GNDA.n1604 GNDA.n1598 4.5005
R12083 GNDA.n1608 GNDA.n1605 4.5005
R12084 GNDA.n1609 GNDA.n1597 4.5005
R12085 GNDA.n1613 GNDA.n1612 4.5005
R12086 GNDA.n1614 GNDA.n1596 4.5005
R12087 GNDA.n1618 GNDA.n1615 4.5005
R12088 GNDA.n1619 GNDA.n1595 4.5005
R12089 GNDA.n1623 GNDA.n1622 4.5005
R12090 GNDA.n1624 GNDA.n1594 4.5005
R12091 GNDA.n1628 GNDA.n1625 4.5005
R12092 GNDA.n1629 GNDA.n1593 4.5005
R12093 GNDA.n1633 GNDA.n1632 4.5005
R12094 GNDA.n1634 GNDA.n1592 4.5005
R12095 GNDA.n1638 GNDA.n1635 4.5005
R12096 GNDA.n1639 GNDA.n1591 4.5005
R12097 GNDA.n1643 GNDA.n1642 4.5005
R12098 GNDA.n1644 GNDA.n1590 4.5005
R12099 GNDA.n1648 GNDA.n1645 4.5005
R12100 GNDA.n1649 GNDA.n1589 4.5005
R12101 GNDA.n1653 GNDA.n1652 4.5005
R12102 GNDA.n1518 GNDA.n1517 4.5005
R12103 GNDA.n1521 GNDA.n1520 4.5005
R12104 GNDA.n1522 GNDA.n1516 4.5005
R12105 GNDA.n1526 GNDA.n1523 4.5005
R12106 GNDA.n1527 GNDA.n1515 4.5005
R12107 GNDA.n1531 GNDA.n1530 4.5005
R12108 GNDA.n1532 GNDA.n1514 4.5005
R12109 GNDA.n1536 GNDA.n1533 4.5005
R12110 GNDA.n1537 GNDA.n1513 4.5005
R12111 GNDA.n1541 GNDA.n1540 4.5005
R12112 GNDA.n1542 GNDA.n1512 4.5005
R12113 GNDA.n1546 GNDA.n1543 4.5005
R12114 GNDA.n1547 GNDA.n1511 4.5005
R12115 GNDA.n1551 GNDA.n1550 4.5005
R12116 GNDA.n1552 GNDA.n1510 4.5005
R12117 GNDA.n1556 GNDA.n1553 4.5005
R12118 GNDA.n1557 GNDA.n1509 4.5005
R12119 GNDA.n1561 GNDA.n1560 4.5005
R12120 GNDA.n1562 GNDA.n1508 4.5005
R12121 GNDA.n1566 GNDA.n1563 4.5005
R12122 GNDA.n1567 GNDA.n1507 4.5005
R12123 GNDA.n1571 GNDA.n1570 4.5005
R12124 GNDA.n1436 GNDA.n1435 4.5005
R12125 GNDA.n1439 GNDA.n1438 4.5005
R12126 GNDA.n1440 GNDA.n1434 4.5005
R12127 GNDA.n1444 GNDA.n1441 4.5005
R12128 GNDA.n1445 GNDA.n1433 4.5005
R12129 GNDA.n1449 GNDA.n1448 4.5005
R12130 GNDA.n1450 GNDA.n1432 4.5005
R12131 GNDA.n1454 GNDA.n1451 4.5005
R12132 GNDA.n1455 GNDA.n1431 4.5005
R12133 GNDA.n1459 GNDA.n1458 4.5005
R12134 GNDA.n1460 GNDA.n1430 4.5005
R12135 GNDA.n1464 GNDA.n1461 4.5005
R12136 GNDA.n1465 GNDA.n1429 4.5005
R12137 GNDA.n1469 GNDA.n1468 4.5005
R12138 GNDA.n1470 GNDA.n1428 4.5005
R12139 GNDA.n1474 GNDA.n1471 4.5005
R12140 GNDA.n1475 GNDA.n1427 4.5005
R12141 GNDA.n1479 GNDA.n1478 4.5005
R12142 GNDA.n1480 GNDA.n1426 4.5005
R12143 GNDA.n1484 GNDA.n1481 4.5005
R12144 GNDA.n1485 GNDA.n1425 4.5005
R12145 GNDA.n1489 GNDA.n1488 4.5005
R12146 GNDA.n1249 GNDA.n1248 4.5005
R12147 GNDA.n1170 GNDA.n1169 4.5005
R12148 GNDA.n1192 GNDA.n1171 4.5005
R12149 GNDA.n1193 GNDA.n1172 4.5005
R12150 GNDA.n1194 GNDA.n1173 4.5005
R12151 GNDA.n1195 GNDA.n1174 4.5005
R12152 GNDA.n1196 GNDA.n1175 4.5005
R12153 GNDA.n1197 GNDA.n1176 4.5005
R12154 GNDA.n1198 GNDA.n1177 4.5005
R12155 GNDA.n1199 GNDA.n1178 4.5005
R12156 GNDA.n1200 GNDA.n1179 4.5005
R12157 GNDA.n1201 GNDA.n1180 4.5005
R12158 GNDA.n1202 GNDA.n1181 4.5005
R12159 GNDA.n1203 GNDA.n1182 4.5005
R12160 GNDA.n1204 GNDA.n1183 4.5005
R12161 GNDA.n1205 GNDA.n1184 4.5005
R12162 GNDA.n1206 GNDA.n1185 4.5005
R12163 GNDA.n1207 GNDA.n1186 4.5005
R12164 GNDA.n1208 GNDA.n1187 4.5005
R12165 GNDA.n1209 GNDA.n1188 4.5005
R12166 GNDA.n1210 GNDA.n1189 4.5005
R12167 GNDA.n1211 GNDA.n1190 4.5005
R12168 GNDA.n1868 GNDA.n1867 4.5005
R12169 GNDA.n1871 GNDA.n1870 4.5005
R12170 GNDA.n1872 GNDA.n1165 4.5005
R12171 GNDA.n1876 GNDA.n1873 4.5005
R12172 GNDA.n1877 GNDA.n1164 4.5005
R12173 GNDA.n1881 GNDA.n1880 4.5005
R12174 GNDA.n1882 GNDA.n1163 4.5005
R12175 GNDA.n1886 GNDA.n1883 4.5005
R12176 GNDA.n1887 GNDA.n1162 4.5005
R12177 GNDA.n1891 GNDA.n1890 4.5005
R12178 GNDA.n1892 GNDA.n1161 4.5005
R12179 GNDA.n1896 GNDA.n1893 4.5005
R12180 GNDA.n1897 GNDA.n1160 4.5005
R12181 GNDA.n1901 GNDA.n1900 4.5005
R12182 GNDA.n1902 GNDA.n1159 4.5005
R12183 GNDA.n1906 GNDA.n1903 4.5005
R12184 GNDA.n1907 GNDA.n1158 4.5005
R12185 GNDA.n1911 GNDA.n1910 4.5005
R12186 GNDA.n1912 GNDA.n1157 4.5005
R12187 GNDA.n1916 GNDA.n1913 4.5005
R12188 GNDA.n1917 GNDA.n1156 4.5005
R12189 GNDA.n1921 GNDA.n1920 4.5005
R12190 GNDA.n1840 GNDA.n1839 4.5005
R12191 GNDA.n1838 GNDA.n1773 4.5005
R12192 GNDA.n1837 GNDA.n1836 4.5005
R12193 GNDA.n1835 GNDA.n1776 4.5005
R12194 GNDA.n1834 GNDA.n1833 4.5005
R12195 GNDA.n1832 GNDA.n1777 4.5005
R12196 GNDA.n1831 GNDA.n1830 4.5005
R12197 GNDA.n1829 GNDA.n1782 4.5005
R12198 GNDA.n1828 GNDA.n1827 4.5005
R12199 GNDA.n1826 GNDA.n1783 4.5005
R12200 GNDA.n1825 GNDA.n1824 4.5005
R12201 GNDA.n1823 GNDA.n1788 4.5005
R12202 GNDA.n1822 GNDA.n1821 4.5005
R12203 GNDA.n1820 GNDA.n1789 4.5005
R12204 GNDA.n1819 GNDA.n1818 4.5005
R12205 GNDA.n1817 GNDA.n1794 4.5005
R12206 GNDA.n1816 GNDA.n1815 4.5005
R12207 GNDA.n1814 GNDA.n1795 4.5005
R12208 GNDA.n1813 GNDA.n1812 4.5005
R12209 GNDA.n1811 GNDA.n1800 4.5005
R12210 GNDA.n1810 GNDA.n1809 4.5005
R12211 GNDA.n1808 GNDA.n1801 4.5005
R12212 GNDA.n1849 GNDA.n1847 4.5005
R12213 GNDA.n1851 GNDA.n1850 4.5005
R12214 GNDA.n1850 GNDA.n1849 4.5005
R12215 GNDA.n1854 GNDA.n1852 4.5005
R12216 GNDA.n1856 GNDA.n1855 4.5005
R12217 GNDA.n1855 GNDA.n1854 4.5005
R12218 GNDA.n1859 GNDA.n1857 4.5005
R12219 GNDA.n1861 GNDA.n1860 4.5005
R12220 GNDA.n1860 GNDA.n1859 4.5005
R12221 GNDA.n1862 GNDA.n1767 4.5005
R12222 GNDA.n1863 GNDA.n1862 4.5005
R12223 GNDA.n1864 GNDA.n1863 4.5005
R12224 GNDA.n1763 GNDA.n1168 4.5005
R12225 GNDA.n1766 GNDA.n1168 4.5005
R12226 GNDA.n1766 GNDA.n1167 4.5005
R12227 GNDA.n1755 GNDA.n1392 4.5005
R12228 GNDA.n1758 GNDA.n1392 4.5005
R12229 GNDA.n1758 GNDA.n1391 4.5005
R12230 GNDA.n1751 GNDA.n1397 4.5005
R12231 GNDA.n1754 GNDA.n1397 4.5005
R12232 GNDA.n1754 GNDA.n1396 4.5005
R12233 GNDA.n1739 GNDA.n1403 4.5005
R12234 GNDA.n1742 GNDA.n1403 4.5005
R12235 GNDA.n1742 GNDA.n1401 4.5005
R12236 GNDA.n3243 GNDA.n3242 4.5005
R12237 GNDA.n3242 GNDA.n3241 4.5005
R12238 GNDA.n3241 GNDA.n3157 4.5005
R12239 GNDA.n3244 GNDA.n588 4.5005
R12240 GNDA.n3245 GNDA.n3244 4.5005
R12241 GNDA.n3246 GNDA.n3245 4.5005
R12242 GNDA.n3477 GNDA.n3476 4.5005
R12243 GNDA.n3476 GNDA.n3475 4.5005
R12244 GNDA.n3475 GNDA.n3391 4.5005
R12245 GNDA.n3478 GNDA.n548 4.5005
R12246 GNDA.n3479 GNDA.n3478 4.5005
R12247 GNDA.n3480 GNDA.n3479 4.5005
R12248 GNDA.n3624 GNDA.n3623 4.5005
R12249 GNDA.n3623 GNDA.n3622 4.5005
R12250 GNDA.n3622 GNDA.n549 4.5005
R12251 GNDA.n3712 GNDA.n508 4.5005
R12252 GNDA.n3713 GNDA.n3712 4.5005
R12253 GNDA.n3714 GNDA.n3713 4.5005
R12254 GNDA.n3858 GNDA.n3857 4.5005
R12255 GNDA.n3857 GNDA.n3856 4.5005
R12256 GNDA.n3856 GNDA.n509 4.5005
R12257 GNDA.n4614 GNDA.n439 4.5005
R12258 GNDA.n4617 GNDA.n439 4.5005
R12259 GNDA.n4617 GNDA.n438 4.5005
R12260 GNDA.n4610 GNDA.n444 4.5005
R12261 GNDA.n4613 GNDA.n444 4.5005
R12262 GNDA.n4613 GNDA.n443 4.5005
R12263 GNDA.n3949 GNDA.n437 4.5005
R12264 GNDA.n3950 GNDA.n3949 4.5005
R12265 GNDA.n3951 GNDA.n3950 4.5005
R12266 GNDA.n4602 GNDA.n453 4.5005
R12267 GNDA.n4605 GNDA.n453 4.5005
R12268 GNDA.n4605 GNDA.n452 4.5005
R12269 GNDA.n4598 GNDA.n458 4.5005
R12270 GNDA.n4601 GNDA.n458 4.5005
R12271 GNDA.n4601 GNDA.n457 4.5005
R12272 GNDA.n4594 GNDA.n463 4.5005
R12273 GNDA.n4597 GNDA.n463 4.5005
R12274 GNDA.n4597 GNDA.n462 4.5005
R12275 GNDA.n4590 GNDA.n468 4.5005
R12276 GNDA.n4593 GNDA.n468 4.5005
R12277 GNDA.n4593 GNDA.n467 4.5005
R12278 GNDA.n4586 GNDA.n473 4.5005
R12279 GNDA.n4589 GNDA.n473 4.5005
R12280 GNDA.n4589 GNDA.n472 4.5005
R12281 GNDA.n1759 GNDA.n1388 4.5005
R12282 GNDA.n1762 GNDA.n1388 4.5005
R12283 GNDA.n1762 GNDA.n1253 4.5005
R12284 GNDA.n4606 GNDA.n449 4.5005
R12285 GNDA.n4609 GNDA.n449 4.5005
R12286 GNDA.n4609 GNDA.n448 4.5005
R12287 GNDA.n3390 GNDA.n3389 4.5005
R12288 GNDA.n3389 GNDA.n3388 4.5005
R12289 GNDA.n3388 GNDA.n589 4.5005
R12290 GNDA.n3711 GNDA.n3710 4.5005
R12291 GNDA.n3710 GNDA.n3709 4.5005
R12292 GNDA.n3709 GNDA.n3625 4.5005
R12293 GNDA.n2296 GNDA.n2295 4.5005
R12294 GNDA.n2391 GNDA.n2390 4.5005
R12295 GNDA.n2286 GNDA.n2285 4.5005
R12296 GNDA.n2396 GNDA.n2279 4.5005
R12297 GNDA.n2395 GNDA.n703 4.5005
R12298 GNDA.n2396 GNDA.n2395 4.5005
R12299 GNDA.n2165 GNDA.n2159 4.5005
R12300 GNDA.n2167 GNDA.n2166 4.5005
R12301 GNDA.n2168 GNDA.n2158 4.5005
R12302 GNDA.n2172 GNDA.n2171 4.5005
R12303 GNDA.n2173 GNDA.n2155 4.5005
R12304 GNDA.n2175 GNDA.n2174 4.5005
R12305 GNDA.n2176 GNDA.n2154 4.5005
R12306 GNDA.n2180 GNDA.n2179 4.5005
R12307 GNDA.n2181 GNDA.n2151 4.5005
R12308 GNDA.n2183 GNDA.n2182 4.5005
R12309 GNDA.n2184 GNDA.n2150 4.5005
R12310 GNDA.n2188 GNDA.n2187 4.5005
R12311 GNDA.n2189 GNDA.n2147 4.5005
R12312 GNDA.n2191 GNDA.n2190 4.5005
R12313 GNDA.n2192 GNDA.n2146 4.5005
R12314 GNDA.n2196 GNDA.n2195 4.5005
R12315 GNDA.n2197 GNDA.n2143 4.5005
R12316 GNDA.n2199 GNDA.n2198 4.5005
R12317 GNDA.n2200 GNDA.n2142 4.5005
R12318 GNDA.n2204 GNDA.n2203 4.5005
R12319 GNDA.n2205 GNDA.n2141 4.5005
R12320 GNDA.n2219 GNDA.n2218 4.5005
R12321 GNDA.n702 GNDA.n701 4.5005
R12322 GNDA.n2212 GNDA.n2211 4.5005
R12323 GNDA.n2215 GNDA.n699 4.5005
R12324 GNDA.n2211 GNDA.n699 4.5005
R12325 GNDA.n2208 GNDA.n359 4.5005
R12326 GNDA.n2231 GNDA.n2230 4.5005
R12327 GNDA.n2234 GNDA.n840 4.5005
R12328 GNDA.n2078 GNDA.n2074 4.5005
R12329 GNDA.n2082 GNDA.n2081 4.5005
R12330 GNDA.n2083 GNDA.n2073 4.5005
R12331 GNDA.n2087 GNDA.n2084 4.5005
R12332 GNDA.n2088 GNDA.n2072 4.5005
R12333 GNDA.n2092 GNDA.n2091 4.5005
R12334 GNDA.n2093 GNDA.n2071 4.5005
R12335 GNDA.n2097 GNDA.n2094 4.5005
R12336 GNDA.n2098 GNDA.n2070 4.5005
R12337 GNDA.n2102 GNDA.n2101 4.5005
R12338 GNDA.n2103 GNDA.n2069 4.5005
R12339 GNDA.n2107 GNDA.n2104 4.5005
R12340 GNDA.n2108 GNDA.n2068 4.5005
R12341 GNDA.n2112 GNDA.n2111 4.5005
R12342 GNDA.n2113 GNDA.n2067 4.5005
R12343 GNDA.n2117 GNDA.n2114 4.5005
R12344 GNDA.n2118 GNDA.n2066 4.5005
R12345 GNDA.n2122 GNDA.n2121 4.5005
R12346 GNDA.n2123 GNDA.n2065 4.5005
R12347 GNDA.n2125 GNDA.n2124 4.5005
R12348 GNDA.n844 GNDA.n843 4.5005
R12349 GNDA.n2225 GNDA.n2224 4.5005
R12350 GNDA.n3128 GNDA.t274 4.47811
R12351 GNDA.t28 GNDA.n3098 4.47811
R12352 GNDA.n346 GNDA.n302 4.26717
R12353 GNDA.n346 GNDA.n345 4.26717
R12354 GNDA.n345 GNDA.n344 4.26717
R12355 GNDA.n344 GNDA.n310 4.26717
R12356 GNDA.n338 GNDA.n310 4.26717
R12357 GNDA.n338 GNDA.n337 4.26717
R12358 GNDA.n337 GNDA.n336 4.26717
R12359 GNDA.n336 GNDA.n318 4.26717
R12360 GNDA.n330 GNDA.n318 4.26717
R12361 GNDA.n330 GNDA.n329 4.26717
R12362 GNDA.n329 GNDA.n328 4.26717
R12363 GNDA.n5082 GNDA.n134 4.26717
R12364 GNDA.n5076 GNDA.n134 4.26717
R12365 GNDA.n5076 GNDA.n5075 4.26717
R12366 GNDA.n5075 GNDA.n5074 4.26717
R12367 GNDA.n5074 GNDA.n5072 4.26717
R12368 GNDA.n5072 GNDA.n5069 4.26717
R12369 GNDA.n5069 GNDA.n5068 4.26717
R12370 GNDA.n5068 GNDA.n5065 4.26717
R12371 GNDA.n5065 GNDA.n5064 4.26717
R12372 GNDA.n5064 GNDA.n5061 4.26717
R12373 GNDA.n5061 GNDA.n5060 4.26717
R12374 GNDA.n2944 GNDA.n827 4.26717
R12375 GNDA.n2950 GNDA.n827 4.26717
R12376 GNDA.n2950 GNDA.n823 4.26717
R12377 GNDA.n2955 GNDA.n823 4.26717
R12378 GNDA.n2955 GNDA.n821 4.26717
R12379 GNDA.n821 GNDA.n818 4.26717
R12380 GNDA.n2962 GNDA.n818 4.26717
R12381 GNDA.n2962 GNDA.n816 4.26717
R12382 GNDA.n816 GNDA.n814 4.26717
R12383 GNDA.n2969 GNDA.n814 4.26717
R12384 GNDA.n2969 GNDA.n812 4.26717
R12385 GNDA.n411 GNDA.n410 4.26717
R12386 GNDA.n410 GNDA.n371 4.26717
R12387 GNDA.n405 GNDA.n371 4.26717
R12388 GNDA.n405 GNDA.n404 4.26717
R12389 GNDA.n404 GNDA.n403 4.26717
R12390 GNDA.n403 GNDA.n379 4.26717
R12391 GNDA.n397 GNDA.n379 4.26717
R12392 GNDA.n397 GNDA.n396 4.26717
R12393 GNDA.n396 GNDA.n395 4.26717
R12394 GNDA.n395 GNDA.n390 4.26717
R12395 GNDA.n390 GNDA.n389 4.26717
R12396 GNDA.n2791 GNDA.n2588 4.26717
R12397 GNDA.n2791 GNDA.n2586 4.26717
R12398 GNDA.n2797 GNDA.n2586 4.26717
R12399 GNDA.n2797 GNDA.n2584 4.26717
R12400 GNDA.n2803 GNDA.n2584 4.26717
R12401 GNDA.n2803 GNDA.n2582 4.26717
R12402 GNDA.n2809 GNDA.n2582 4.26717
R12403 GNDA.n2809 GNDA.n2580 4.26717
R12404 GNDA.n2815 GNDA.n2580 4.26717
R12405 GNDA.n2815 GNDA.n2578 4.26717
R12406 GNDA.n2820 GNDA.n2578 4.26717
R12407 GNDA.n2917 GNDA.n2826 4.26717
R12408 GNDA.n2917 GNDA.n2828 4.26717
R12409 GNDA.n2857 GNDA.n2828 4.26717
R12410 GNDA.n2857 GNDA.n2856 4.26717
R12411 GNDA.n2856 GNDA.n2833 4.26717
R12412 GNDA.n2851 GNDA.n2833 4.26717
R12413 GNDA.n2851 GNDA.n2850 4.26717
R12414 GNDA.n2850 GNDA.n2849 4.26717
R12415 GNDA.n2849 GNDA.n2844 4.26717
R12416 GNDA.n2844 GNDA.n750 4.26717
R12417 GNDA.n2980 GNDA.n750 4.26717
R12418 GNDA.t232 GNDA.t246 4.14363
R12419 GNDA.n4702 GNDA.n302 3.93531
R12420 GNDA.n5083 GNDA.n5082 3.93531
R12421 GNDA.n2944 GNDA.n2564 3.93531
R12422 GNDA.n411 GNDA.n365 3.93531
R12423 GNDA.n2612 GNDA.n2588 3.93531
R12424 GNDA.n2826 GNDA.n2824 3.93531
R12425 GNDA.n4619 GNDA.n4618 3.84081
R12426 GNDA.n3156 GNDA.n3155 3.84081
R12427 GNDA.n1750 GNDA.n1749 3.84081
R12428 GNDA.n3861 GNDA.n3860 3.84045
R12429 GNDA.n3002 GNDA.n745 3.7893
R12430 GNDA.n3001 GNDA.n746 3.7893
R12431 GNDA.n2989 GNDA.n2988 3.7893
R12432 GNDA.n2995 GNDA.n2994 3.7893
R12433 GNDA.n2991 GNDA.n2990 3.7893
R12434 GNDA.n721 GNDA.n714 3.7893
R12435 GNDA.n727 GNDA.n725 3.7893
R12436 GNDA.n726 GNDA.n689 3.7893
R12437 GNDA.n3079 GNDA.n671 3.7893
R12438 GNDA.n3078 GNDA.n672 3.7893
R12439 GNDA.n3066 GNDA.n3065 3.7893
R12440 GNDA.n3072 GNDA.n3071 3.7893
R12441 GNDA.n3068 GNDA.n3067 3.7893
R12442 GNDA.n2305 GNDA.n650 3.7893
R12443 GNDA.n2312 GNDA.n2310 3.7893
R12444 GNDA.n2314 GNDA.n2313 3.7893
R12445 GNDA.n5054 GNDA.n165 3.7893
R12446 GNDA.n5051 GNDA.n5050 3.7893
R12447 GNDA.n200 GNDA.n167 3.7893
R12448 GNDA.n218 GNDA.n217 3.7893
R12449 GNDA.n215 GNDA.n214 3.7893
R12450 GNDA.n210 GNDA.n203 3.7893
R12451 GNDA.n207 GNDA.n206 3.7893
R12452 GNDA.n4992 GNDA.n187 3.7893
R12453 GNDA.n2727 GNDA.n2702 3.7893
R12454 GNDA.n2726 GNDA.n2723 3.7893
R12455 GNDA.n2722 GNDA.n2703 3.7893
R12456 GNDA.n2719 GNDA.n2718 3.7893
R12457 GNDA.n2715 GNDA.n2704 3.7893
R12458 GNDA.n2708 GNDA.n2705 3.7893
R12459 GNDA.n2732 GNDA.n2627 3.7893
R12460 GNDA.n2733 GNDA.n2626 3.7893
R12461 GNDA.n4983 GNDA.n4982 3.7893
R12462 GNDA.n4979 GNDA.n4873 3.7893
R12463 GNDA.n4978 GNDA.n4876 3.7893
R12464 GNDA.n4975 GNDA.n4974 3.7893
R12465 GNDA.n4901 GNDA.n4877 3.7893
R12466 GNDA.n4910 GNDA.n4909 3.7893
R12467 GNDA.n4913 GNDA.n4900 3.7893
R12468 GNDA.n4918 GNDA.n4914 3.7893
R12469 GNDA.n5262 GNDA.n5261 3.7893
R12470 GNDA.n5258 GNDA.n59 3.7893
R12471 GNDA.n5257 GNDA.n62 3.7893
R12472 GNDA.n5254 GNDA.n5253 3.7893
R12473 GNDA.n5180 GNDA.n63 3.7893
R12474 GNDA.n5189 GNDA.n5188 3.7893
R12475 GNDA.n5192 GNDA.n5179 3.7893
R12476 GNDA.n5197 GNDA.n5193 3.7893
R12477 GNDA.n4839 GNDA.n4728 3.7893
R12478 GNDA.n4836 GNDA.n4835 3.7893
R12479 GNDA.n4752 GNDA.n4729 3.7893
R12480 GNDA.n4757 GNDA.n4755 3.7893
R12481 GNDA.n4762 GNDA.n4758 3.7893
R12482 GNDA.n4769 GNDA.n4768 3.7893
R12483 GNDA.n4772 GNDA.n4751 3.7893
R12484 GNDA.n4777 GNDA.n4773 3.7893
R12485 GNDA.n2491 GNDA.n2489 3.7893
R12486 GNDA.n2490 GNDA.n2251 3.7893
R12487 GNDA.n2497 GNDA.n2496 3.7893
R12488 GNDA.n2412 GNDA.n2252 3.7893
R12489 GNDA.n2416 GNDA.n2414 3.7893
R12490 GNDA.n2423 GNDA.n2422 3.7893
R12491 GNDA.n2432 GNDA.n2272 3.7893
R12492 GNDA.n2431 GNDA.n2270 3.7893
R12493 GNDA.n5271 GNDA.n22 3.7893
R12494 GNDA.n5270 GNDA.n23 3.7893
R12495 GNDA.n33 GNDA.n32 3.7893
R12496 GNDA.n39 GNDA.n38 3.7893
R12497 GNDA.n35 GNDA.n34 3.7893
R12498 GNDA.n5105 GNDA.n1 3.7893
R12499 GNDA.n5110 GNDA.n5108 3.7893
R12500 GNDA.n5115 GNDA.n5111 3.7893
R12501 GNDA GNDA.n3007 3.7381
R12502 GNDA GNDA.n3084 3.7381
R12503 GNDA.n211 GNDA 3.7381
R12504 GNDA GNDA.n2711 3.7381
R12505 GNDA.n4906 GNDA 3.7381
R12506 GNDA.n5185 GNDA 3.7381
R12507 GNDA.n4765 GNDA 3.7381
R12508 GNDA.n2421 GNDA 3.7381
R12509 GNDA GNDA.n5276 3.7381
R12510 GNDA.n3136 GNDA.n3130 3.65764
R12511 GNDA.n3136 GNDA.n3135 3.65764
R12512 GNDA.n635 GNDA.n630 3.65764
R12513 GNDA.n635 GNDA.n634 3.65764
R12514 GNDA.n1806 GNDA.n1129 3.50398
R12515 GNDA.n2075 GNDA.n2053 3.47871
R12516 GNDA.n3672 GNDA.n3671 3.47821
R12517 GNDA.n3381 GNDA.n3380 3.47821
R12518 GNDA.n4578 GNDA.n4577 3.47821
R12519 GNDA.n4502 GNDA.n4501 3.47821
R12520 GNDA.n4420 GNDA.n4419 3.47821
R12521 GNDA.n4338 GNDA.n4337 3.47821
R12522 GNDA.n4256 GNDA.n4255 3.47821
R12523 GNDA.n4010 GNDA.n4009 3.47821
R12524 GNDA.n4174 GNDA.n4173 3.47821
R12525 GNDA.n4092 GNDA.n4091 3.47821
R12526 GNDA.n3907 GNDA.n3906 3.47821
R12527 GNDA.n1731 GNDA.n1730 3.47821
R12528 GNDA.n3849 GNDA.n3848 3.47821
R12529 GNDA.n3773 GNDA.n3772 3.47821
R12530 GNDA.n3615 GNDA.n3614 3.47821
R12531 GNDA.n3539 GNDA.n3538 3.47821
R12532 GNDA.n3436 GNDA.n3435 3.47821
R12533 GNDA.n3305 GNDA.n3304 3.47821
R12534 GNDA.n3202 GNDA.n3201 3.47821
R12535 GNDA.n1655 GNDA.n1654 3.47821
R12536 GNDA.n1573 GNDA.n1572 3.47821
R12537 GNDA.n1491 GNDA.n1490 3.47821
R12538 GNDA.n1213 GNDA.n1212 3.47821
R12539 GNDA.n1923 GNDA.n1922 3.47821
R12540 GNDA.n2164 GNDA.n2128 3.47821
R12541 GNDA.n1839 GNDA.n1130 3.43627
R12542 GNDA.n3948 GNDA.t5 3.42907
R12543 GNDA.n3948 GNDA.t215 3.42907
R12544 GNDA.n3945 GNDA.t16 3.42907
R12545 GNDA.n3945 GNDA.t260 3.42907
R12546 GNDA.n1407 GNDA.t268 3.42907
R12547 GNDA.n1407 GNDA.t31 3.42907
R12548 GNDA.n1402 GNDA.t159 3.42907
R12549 GNDA.n1402 GNDA.t236 3.42907
R12550 GNDA.n3673 GNDA.n3670 3.4105
R12551 GNDA.n3674 GNDA.n3668 3.4105
R12552 GNDA.n3675 GNDA.n3667 3.4105
R12553 GNDA.n3665 GNDA.n3663 3.4105
R12554 GNDA.n3679 GNDA.n3662 3.4105
R12555 GNDA.n3680 GNDA.n3660 3.4105
R12556 GNDA.n3681 GNDA.n3659 3.4105
R12557 GNDA.n3657 GNDA.n3655 3.4105
R12558 GNDA.n3685 GNDA.n3654 3.4105
R12559 GNDA.n3686 GNDA.n3652 3.4105
R12560 GNDA.n3687 GNDA.n3651 3.4105
R12561 GNDA.n3649 GNDA.n3647 3.4105
R12562 GNDA.n3691 GNDA.n3646 3.4105
R12563 GNDA.n3692 GNDA.n3644 3.4105
R12564 GNDA.n3693 GNDA.n3643 3.4105
R12565 GNDA.n3641 GNDA.n3639 3.4105
R12566 GNDA.n3697 GNDA.n3638 3.4105
R12567 GNDA.n3698 GNDA.n3636 3.4105
R12568 GNDA.n3699 GNDA.n3635 3.4105
R12569 GNDA.n3633 GNDA.n3631 3.4105
R12570 GNDA.n3703 GNDA.n3630 3.4105
R12571 GNDA.n3704 GNDA.n3628 3.4105
R12572 GNDA.n3705 GNDA.n3627 3.4105
R12573 GNDA.n3319 GNDA.n3318 3.4105
R12574 GNDA.n3378 GNDA.n3377 3.4105
R12575 GNDA.n3376 GNDA.n3375 3.4105
R12576 GNDA.n3374 GNDA.n3373 3.4105
R12577 GNDA.n3372 GNDA.n3321 3.4105
R12578 GNDA.n3368 GNDA.n3367 3.4105
R12579 GNDA.n3366 GNDA.n3365 3.4105
R12580 GNDA.n3364 GNDA.n3363 3.4105
R12581 GNDA.n3362 GNDA.n3323 3.4105
R12582 GNDA.n3358 GNDA.n3357 3.4105
R12583 GNDA.n3356 GNDA.n3355 3.4105
R12584 GNDA.n3354 GNDA.n3353 3.4105
R12585 GNDA.n3352 GNDA.n3325 3.4105
R12586 GNDA.n3348 GNDA.n3347 3.4105
R12587 GNDA.n3346 GNDA.n3345 3.4105
R12588 GNDA.n3344 GNDA.n3343 3.4105
R12589 GNDA.n3342 GNDA.n3327 3.4105
R12590 GNDA.n3338 GNDA.n3337 3.4105
R12591 GNDA.n3336 GNDA.n3335 3.4105
R12592 GNDA.n3334 GNDA.n3333 3.4105
R12593 GNDA.n3332 GNDA.n3329 3.4105
R12594 GNDA.n592 GNDA.n591 3.4105
R12595 GNDA.n3384 GNDA.n3383 3.4105
R12596 GNDA.n4516 GNDA.n4515 3.4105
R12597 GNDA.n4575 GNDA.n4574 3.4105
R12598 GNDA.n4573 GNDA.n4572 3.4105
R12599 GNDA.n4571 GNDA.n4570 3.4105
R12600 GNDA.n4569 GNDA.n4518 3.4105
R12601 GNDA.n4565 GNDA.n4564 3.4105
R12602 GNDA.n4563 GNDA.n4562 3.4105
R12603 GNDA.n4561 GNDA.n4560 3.4105
R12604 GNDA.n4559 GNDA.n4520 3.4105
R12605 GNDA.n4555 GNDA.n4554 3.4105
R12606 GNDA.n4553 GNDA.n4552 3.4105
R12607 GNDA.n4551 GNDA.n4550 3.4105
R12608 GNDA.n4549 GNDA.n4522 3.4105
R12609 GNDA.n4545 GNDA.n4544 3.4105
R12610 GNDA.n4543 GNDA.n4542 3.4105
R12611 GNDA.n4541 GNDA.n4540 3.4105
R12612 GNDA.n4539 GNDA.n4524 3.4105
R12613 GNDA.n4535 GNDA.n4534 3.4105
R12614 GNDA.n4533 GNDA.n4532 3.4105
R12615 GNDA.n4531 GNDA.n4530 3.4105
R12616 GNDA.n4529 GNDA.n4526 3.4105
R12617 GNDA.n476 GNDA.n475 3.4105
R12618 GNDA.n4581 GNDA.n4580 3.4105
R12619 GNDA.n4435 GNDA.n4434 3.4105
R12620 GNDA.n4499 GNDA.n4498 3.4105
R12621 GNDA.n4497 GNDA.n4496 3.4105
R12622 GNDA.n4495 GNDA.n4494 3.4105
R12623 GNDA.n4493 GNDA.n4437 3.4105
R12624 GNDA.n4489 GNDA.n4488 3.4105
R12625 GNDA.n4487 GNDA.n4486 3.4105
R12626 GNDA.n4485 GNDA.n4484 3.4105
R12627 GNDA.n4483 GNDA.n4439 3.4105
R12628 GNDA.n4479 GNDA.n4478 3.4105
R12629 GNDA.n4477 GNDA.n4476 3.4105
R12630 GNDA.n4475 GNDA.n4474 3.4105
R12631 GNDA.n4473 GNDA.n4441 3.4105
R12632 GNDA.n4469 GNDA.n4468 3.4105
R12633 GNDA.n4467 GNDA.n4466 3.4105
R12634 GNDA.n4465 GNDA.n4464 3.4105
R12635 GNDA.n4463 GNDA.n4443 3.4105
R12636 GNDA.n4459 GNDA.n4458 3.4105
R12637 GNDA.n4457 GNDA.n4456 3.4105
R12638 GNDA.n4455 GNDA.n4454 3.4105
R12639 GNDA.n4453 GNDA.n4445 3.4105
R12640 GNDA.n4449 GNDA.n4448 3.4105
R12641 GNDA.n4447 GNDA.n4422 3.4105
R12642 GNDA.n4353 GNDA.n4352 3.4105
R12643 GNDA.n4417 GNDA.n4416 3.4105
R12644 GNDA.n4415 GNDA.n4414 3.4105
R12645 GNDA.n4413 GNDA.n4412 3.4105
R12646 GNDA.n4411 GNDA.n4355 3.4105
R12647 GNDA.n4407 GNDA.n4406 3.4105
R12648 GNDA.n4405 GNDA.n4404 3.4105
R12649 GNDA.n4403 GNDA.n4402 3.4105
R12650 GNDA.n4401 GNDA.n4357 3.4105
R12651 GNDA.n4397 GNDA.n4396 3.4105
R12652 GNDA.n4395 GNDA.n4394 3.4105
R12653 GNDA.n4393 GNDA.n4392 3.4105
R12654 GNDA.n4391 GNDA.n4359 3.4105
R12655 GNDA.n4387 GNDA.n4386 3.4105
R12656 GNDA.n4385 GNDA.n4384 3.4105
R12657 GNDA.n4383 GNDA.n4382 3.4105
R12658 GNDA.n4381 GNDA.n4361 3.4105
R12659 GNDA.n4377 GNDA.n4376 3.4105
R12660 GNDA.n4375 GNDA.n4374 3.4105
R12661 GNDA.n4373 GNDA.n4372 3.4105
R12662 GNDA.n4371 GNDA.n4363 3.4105
R12663 GNDA.n4367 GNDA.n4366 3.4105
R12664 GNDA.n4365 GNDA.n4340 3.4105
R12665 GNDA.n4271 GNDA.n4270 3.4105
R12666 GNDA.n4335 GNDA.n4334 3.4105
R12667 GNDA.n4333 GNDA.n4332 3.4105
R12668 GNDA.n4331 GNDA.n4330 3.4105
R12669 GNDA.n4329 GNDA.n4273 3.4105
R12670 GNDA.n4325 GNDA.n4324 3.4105
R12671 GNDA.n4323 GNDA.n4322 3.4105
R12672 GNDA.n4321 GNDA.n4320 3.4105
R12673 GNDA.n4319 GNDA.n4275 3.4105
R12674 GNDA.n4315 GNDA.n4314 3.4105
R12675 GNDA.n4313 GNDA.n4312 3.4105
R12676 GNDA.n4311 GNDA.n4310 3.4105
R12677 GNDA.n4309 GNDA.n4277 3.4105
R12678 GNDA.n4305 GNDA.n4304 3.4105
R12679 GNDA.n4303 GNDA.n4302 3.4105
R12680 GNDA.n4301 GNDA.n4300 3.4105
R12681 GNDA.n4299 GNDA.n4279 3.4105
R12682 GNDA.n4295 GNDA.n4294 3.4105
R12683 GNDA.n4293 GNDA.n4292 3.4105
R12684 GNDA.n4291 GNDA.n4290 3.4105
R12685 GNDA.n4289 GNDA.n4281 3.4105
R12686 GNDA.n4285 GNDA.n4284 3.4105
R12687 GNDA.n4283 GNDA.n4258 3.4105
R12688 GNDA.n4189 GNDA.n4188 3.4105
R12689 GNDA.n4253 GNDA.n4252 3.4105
R12690 GNDA.n4251 GNDA.n4250 3.4105
R12691 GNDA.n4249 GNDA.n4248 3.4105
R12692 GNDA.n4247 GNDA.n4191 3.4105
R12693 GNDA.n4243 GNDA.n4242 3.4105
R12694 GNDA.n4241 GNDA.n4240 3.4105
R12695 GNDA.n4239 GNDA.n4238 3.4105
R12696 GNDA.n4237 GNDA.n4193 3.4105
R12697 GNDA.n4233 GNDA.n4232 3.4105
R12698 GNDA.n4231 GNDA.n4230 3.4105
R12699 GNDA.n4229 GNDA.n4228 3.4105
R12700 GNDA.n4227 GNDA.n4195 3.4105
R12701 GNDA.n4223 GNDA.n4222 3.4105
R12702 GNDA.n4221 GNDA.n4220 3.4105
R12703 GNDA.n4219 GNDA.n4218 3.4105
R12704 GNDA.n4217 GNDA.n4197 3.4105
R12705 GNDA.n4213 GNDA.n4212 3.4105
R12706 GNDA.n4211 GNDA.n4210 3.4105
R12707 GNDA.n4209 GNDA.n4208 3.4105
R12708 GNDA.n4207 GNDA.n4199 3.4105
R12709 GNDA.n4203 GNDA.n4202 3.4105
R12710 GNDA.n4201 GNDA.n4176 3.4105
R12711 GNDA.n491 GNDA.n490 3.4105
R12712 GNDA.n4007 GNDA.n4006 3.4105
R12713 GNDA.n4005 GNDA.n4004 3.4105
R12714 GNDA.n4003 GNDA.n4002 3.4105
R12715 GNDA.n4001 GNDA.n493 3.4105
R12716 GNDA.n3997 GNDA.n3996 3.4105
R12717 GNDA.n3995 GNDA.n3994 3.4105
R12718 GNDA.n3993 GNDA.n3992 3.4105
R12719 GNDA.n3991 GNDA.n495 3.4105
R12720 GNDA.n3987 GNDA.n3986 3.4105
R12721 GNDA.n3985 GNDA.n3984 3.4105
R12722 GNDA.n3983 GNDA.n3982 3.4105
R12723 GNDA.n3981 GNDA.n497 3.4105
R12724 GNDA.n3977 GNDA.n3976 3.4105
R12725 GNDA.n3975 GNDA.n3974 3.4105
R12726 GNDA.n3973 GNDA.n3972 3.4105
R12727 GNDA.n3971 GNDA.n499 3.4105
R12728 GNDA.n3967 GNDA.n3966 3.4105
R12729 GNDA.n3965 GNDA.n3964 3.4105
R12730 GNDA.n3963 GNDA.n3962 3.4105
R12731 GNDA.n3961 GNDA.n501 3.4105
R12732 GNDA.n3957 GNDA.n3956 3.4105
R12733 GNDA.n3955 GNDA.n478 3.4105
R12734 GNDA.n4107 GNDA.n4106 3.4105
R12735 GNDA.n4171 GNDA.n4170 3.4105
R12736 GNDA.n4169 GNDA.n4168 3.4105
R12737 GNDA.n4167 GNDA.n4166 3.4105
R12738 GNDA.n4165 GNDA.n4109 3.4105
R12739 GNDA.n4161 GNDA.n4160 3.4105
R12740 GNDA.n4159 GNDA.n4158 3.4105
R12741 GNDA.n4157 GNDA.n4156 3.4105
R12742 GNDA.n4155 GNDA.n4111 3.4105
R12743 GNDA.n4151 GNDA.n4150 3.4105
R12744 GNDA.n4149 GNDA.n4148 3.4105
R12745 GNDA.n4147 GNDA.n4146 3.4105
R12746 GNDA.n4145 GNDA.n4113 3.4105
R12747 GNDA.n4141 GNDA.n4140 3.4105
R12748 GNDA.n4139 GNDA.n4138 3.4105
R12749 GNDA.n4137 GNDA.n4136 3.4105
R12750 GNDA.n4135 GNDA.n4115 3.4105
R12751 GNDA.n4131 GNDA.n4130 3.4105
R12752 GNDA.n4129 GNDA.n4128 3.4105
R12753 GNDA.n4127 GNDA.n4126 3.4105
R12754 GNDA.n4125 GNDA.n4117 3.4105
R12755 GNDA.n4121 GNDA.n4120 3.4105
R12756 GNDA.n4119 GNDA.n4094 3.4105
R12757 GNDA.n4025 GNDA.n4024 3.4105
R12758 GNDA.n4089 GNDA.n4088 3.4105
R12759 GNDA.n4087 GNDA.n4086 3.4105
R12760 GNDA.n4085 GNDA.n4084 3.4105
R12761 GNDA.n4083 GNDA.n4027 3.4105
R12762 GNDA.n4079 GNDA.n4078 3.4105
R12763 GNDA.n4077 GNDA.n4076 3.4105
R12764 GNDA.n4075 GNDA.n4074 3.4105
R12765 GNDA.n4073 GNDA.n4029 3.4105
R12766 GNDA.n4069 GNDA.n4068 3.4105
R12767 GNDA.n4067 GNDA.n4066 3.4105
R12768 GNDA.n4065 GNDA.n4064 3.4105
R12769 GNDA.n4063 GNDA.n4031 3.4105
R12770 GNDA.n4059 GNDA.n4058 3.4105
R12771 GNDA.n4057 GNDA.n4056 3.4105
R12772 GNDA.n4055 GNDA.n4054 3.4105
R12773 GNDA.n4053 GNDA.n4033 3.4105
R12774 GNDA.n4049 GNDA.n4048 3.4105
R12775 GNDA.n4047 GNDA.n4046 3.4105
R12776 GNDA.n4045 GNDA.n4044 3.4105
R12777 GNDA.n4043 GNDA.n4035 3.4105
R12778 GNDA.n4039 GNDA.n4038 3.4105
R12779 GNDA.n4037 GNDA.n4012 3.4105
R12780 GNDA.n3908 GNDA.n3885 3.4105
R12781 GNDA.n3910 GNDA.n3884 3.4105
R12782 GNDA.n3911 GNDA.n3883 3.4105
R12783 GNDA.n3913 GNDA.n3882 3.4105
R12784 GNDA.n3914 GNDA.n3881 3.4105
R12785 GNDA.n3916 GNDA.n3880 3.4105
R12786 GNDA.n3917 GNDA.n3879 3.4105
R12787 GNDA.n3919 GNDA.n3878 3.4105
R12788 GNDA.n3920 GNDA.n3877 3.4105
R12789 GNDA.n3922 GNDA.n3876 3.4105
R12790 GNDA.n3923 GNDA.n3875 3.4105
R12791 GNDA.n3925 GNDA.n3874 3.4105
R12792 GNDA.n3926 GNDA.n3873 3.4105
R12793 GNDA.n3928 GNDA.n3872 3.4105
R12794 GNDA.n3929 GNDA.n3871 3.4105
R12795 GNDA.n3931 GNDA.n3870 3.4105
R12796 GNDA.n3932 GNDA.n3869 3.4105
R12797 GNDA.n3934 GNDA.n3868 3.4105
R12798 GNDA.n3935 GNDA.n3867 3.4105
R12799 GNDA.n3937 GNDA.n3866 3.4105
R12800 GNDA.n3938 GNDA.n3865 3.4105
R12801 GNDA.n3940 GNDA.n3864 3.4105
R12802 GNDA.n3942 GNDA.n3941 3.4105
R12803 GNDA.n1669 GNDA.n1668 3.4105
R12804 GNDA.n1728 GNDA.n1727 3.4105
R12805 GNDA.n1726 GNDA.n1725 3.4105
R12806 GNDA.n1724 GNDA.n1723 3.4105
R12807 GNDA.n1722 GNDA.n1671 3.4105
R12808 GNDA.n1718 GNDA.n1717 3.4105
R12809 GNDA.n1716 GNDA.n1715 3.4105
R12810 GNDA.n1714 GNDA.n1713 3.4105
R12811 GNDA.n1712 GNDA.n1673 3.4105
R12812 GNDA.n1708 GNDA.n1707 3.4105
R12813 GNDA.n1706 GNDA.n1705 3.4105
R12814 GNDA.n1704 GNDA.n1703 3.4105
R12815 GNDA.n1702 GNDA.n1675 3.4105
R12816 GNDA.n1698 GNDA.n1697 3.4105
R12817 GNDA.n1696 GNDA.n1695 3.4105
R12818 GNDA.n1694 GNDA.n1693 3.4105
R12819 GNDA.n1692 GNDA.n1677 3.4105
R12820 GNDA.n1688 GNDA.n1687 3.4105
R12821 GNDA.n1686 GNDA.n1685 3.4105
R12822 GNDA.n1684 GNDA.n1683 3.4105
R12823 GNDA.n1682 GNDA.n1679 3.4105
R12824 GNDA.n1410 GNDA.n1409 3.4105
R12825 GNDA.n1734 GNDA.n1733 3.4105
R12826 GNDA.n3787 GNDA.n3786 3.4105
R12827 GNDA.n3846 GNDA.n3845 3.4105
R12828 GNDA.n3844 GNDA.n3843 3.4105
R12829 GNDA.n3842 GNDA.n3841 3.4105
R12830 GNDA.n3840 GNDA.n3789 3.4105
R12831 GNDA.n3836 GNDA.n3835 3.4105
R12832 GNDA.n3834 GNDA.n3833 3.4105
R12833 GNDA.n3832 GNDA.n3831 3.4105
R12834 GNDA.n3830 GNDA.n3791 3.4105
R12835 GNDA.n3826 GNDA.n3825 3.4105
R12836 GNDA.n3824 GNDA.n3823 3.4105
R12837 GNDA.n3822 GNDA.n3821 3.4105
R12838 GNDA.n3820 GNDA.n3793 3.4105
R12839 GNDA.n3816 GNDA.n3815 3.4105
R12840 GNDA.n3814 GNDA.n3813 3.4105
R12841 GNDA.n3812 GNDA.n3811 3.4105
R12842 GNDA.n3810 GNDA.n3795 3.4105
R12843 GNDA.n3806 GNDA.n3805 3.4105
R12844 GNDA.n3804 GNDA.n3803 3.4105
R12845 GNDA.n3802 GNDA.n3801 3.4105
R12846 GNDA.n3800 GNDA.n3797 3.4105
R12847 GNDA.n512 GNDA.n511 3.4105
R12848 GNDA.n3852 GNDA.n3851 3.4105
R12849 GNDA.n527 GNDA.n526 3.4105
R12850 GNDA.n3770 GNDA.n3769 3.4105
R12851 GNDA.n3768 GNDA.n3767 3.4105
R12852 GNDA.n3766 GNDA.n3765 3.4105
R12853 GNDA.n3764 GNDA.n529 3.4105
R12854 GNDA.n3760 GNDA.n3759 3.4105
R12855 GNDA.n3758 GNDA.n3757 3.4105
R12856 GNDA.n3756 GNDA.n3755 3.4105
R12857 GNDA.n3754 GNDA.n531 3.4105
R12858 GNDA.n3750 GNDA.n3749 3.4105
R12859 GNDA.n3748 GNDA.n3747 3.4105
R12860 GNDA.n3746 GNDA.n3745 3.4105
R12861 GNDA.n3744 GNDA.n533 3.4105
R12862 GNDA.n3740 GNDA.n3739 3.4105
R12863 GNDA.n3738 GNDA.n3737 3.4105
R12864 GNDA.n3736 GNDA.n3735 3.4105
R12865 GNDA.n3734 GNDA.n535 3.4105
R12866 GNDA.n3730 GNDA.n3729 3.4105
R12867 GNDA.n3728 GNDA.n3727 3.4105
R12868 GNDA.n3726 GNDA.n3725 3.4105
R12869 GNDA.n3724 GNDA.n537 3.4105
R12870 GNDA.n3720 GNDA.n3719 3.4105
R12871 GNDA.n3718 GNDA.n514 3.4105
R12872 GNDA.n3553 GNDA.n3552 3.4105
R12873 GNDA.n3612 GNDA.n3611 3.4105
R12874 GNDA.n3610 GNDA.n3609 3.4105
R12875 GNDA.n3608 GNDA.n3607 3.4105
R12876 GNDA.n3606 GNDA.n3555 3.4105
R12877 GNDA.n3602 GNDA.n3601 3.4105
R12878 GNDA.n3600 GNDA.n3599 3.4105
R12879 GNDA.n3598 GNDA.n3597 3.4105
R12880 GNDA.n3596 GNDA.n3557 3.4105
R12881 GNDA.n3592 GNDA.n3591 3.4105
R12882 GNDA.n3590 GNDA.n3589 3.4105
R12883 GNDA.n3588 GNDA.n3587 3.4105
R12884 GNDA.n3586 GNDA.n3559 3.4105
R12885 GNDA.n3582 GNDA.n3581 3.4105
R12886 GNDA.n3580 GNDA.n3579 3.4105
R12887 GNDA.n3578 GNDA.n3577 3.4105
R12888 GNDA.n3576 GNDA.n3561 3.4105
R12889 GNDA.n3572 GNDA.n3571 3.4105
R12890 GNDA.n3570 GNDA.n3569 3.4105
R12891 GNDA.n3568 GNDA.n3567 3.4105
R12892 GNDA.n3566 GNDA.n3563 3.4105
R12893 GNDA.n552 GNDA.n551 3.4105
R12894 GNDA.n3618 GNDA.n3617 3.4105
R12895 GNDA.n567 GNDA.n566 3.4105
R12896 GNDA.n3536 GNDA.n3535 3.4105
R12897 GNDA.n3534 GNDA.n3533 3.4105
R12898 GNDA.n3532 GNDA.n3531 3.4105
R12899 GNDA.n3530 GNDA.n569 3.4105
R12900 GNDA.n3526 GNDA.n3525 3.4105
R12901 GNDA.n3524 GNDA.n3523 3.4105
R12902 GNDA.n3522 GNDA.n3521 3.4105
R12903 GNDA.n3520 GNDA.n571 3.4105
R12904 GNDA.n3516 GNDA.n3515 3.4105
R12905 GNDA.n3514 GNDA.n3513 3.4105
R12906 GNDA.n3512 GNDA.n3511 3.4105
R12907 GNDA.n3510 GNDA.n573 3.4105
R12908 GNDA.n3506 GNDA.n3505 3.4105
R12909 GNDA.n3504 GNDA.n3503 3.4105
R12910 GNDA.n3502 GNDA.n3501 3.4105
R12911 GNDA.n3500 GNDA.n575 3.4105
R12912 GNDA.n3496 GNDA.n3495 3.4105
R12913 GNDA.n3494 GNDA.n3493 3.4105
R12914 GNDA.n3492 GNDA.n3491 3.4105
R12915 GNDA.n3490 GNDA.n577 3.4105
R12916 GNDA.n3486 GNDA.n3485 3.4105
R12917 GNDA.n3484 GNDA.n554 3.4105
R12918 GNDA.n3437 GNDA.n3414 3.4105
R12919 GNDA.n3439 GNDA.n3413 3.4105
R12920 GNDA.n3440 GNDA.n3412 3.4105
R12921 GNDA.n3442 GNDA.n3411 3.4105
R12922 GNDA.n3443 GNDA.n3410 3.4105
R12923 GNDA.n3445 GNDA.n3409 3.4105
R12924 GNDA.n3446 GNDA.n3408 3.4105
R12925 GNDA.n3448 GNDA.n3407 3.4105
R12926 GNDA.n3449 GNDA.n3406 3.4105
R12927 GNDA.n3451 GNDA.n3405 3.4105
R12928 GNDA.n3452 GNDA.n3404 3.4105
R12929 GNDA.n3454 GNDA.n3403 3.4105
R12930 GNDA.n3455 GNDA.n3402 3.4105
R12931 GNDA.n3457 GNDA.n3401 3.4105
R12932 GNDA.n3458 GNDA.n3400 3.4105
R12933 GNDA.n3460 GNDA.n3399 3.4105
R12934 GNDA.n3461 GNDA.n3398 3.4105
R12935 GNDA.n3463 GNDA.n3397 3.4105
R12936 GNDA.n3464 GNDA.n3396 3.4105
R12937 GNDA.n3466 GNDA.n3395 3.4105
R12938 GNDA.n3467 GNDA.n3394 3.4105
R12939 GNDA.n3469 GNDA.n3393 3.4105
R12940 GNDA.n3471 GNDA.n3470 3.4105
R12941 GNDA.n607 GNDA.n606 3.4105
R12942 GNDA.n3302 GNDA.n3301 3.4105
R12943 GNDA.n3300 GNDA.n3299 3.4105
R12944 GNDA.n3298 GNDA.n3297 3.4105
R12945 GNDA.n3296 GNDA.n609 3.4105
R12946 GNDA.n3292 GNDA.n3291 3.4105
R12947 GNDA.n3290 GNDA.n3289 3.4105
R12948 GNDA.n3288 GNDA.n3287 3.4105
R12949 GNDA.n3286 GNDA.n611 3.4105
R12950 GNDA.n3282 GNDA.n3281 3.4105
R12951 GNDA.n3280 GNDA.n3279 3.4105
R12952 GNDA.n3278 GNDA.n3277 3.4105
R12953 GNDA.n3276 GNDA.n613 3.4105
R12954 GNDA.n3272 GNDA.n3271 3.4105
R12955 GNDA.n3270 GNDA.n3269 3.4105
R12956 GNDA.n3268 GNDA.n3267 3.4105
R12957 GNDA.n3266 GNDA.n615 3.4105
R12958 GNDA.n3262 GNDA.n3261 3.4105
R12959 GNDA.n3260 GNDA.n3259 3.4105
R12960 GNDA.n3258 GNDA.n3257 3.4105
R12961 GNDA.n3256 GNDA.n617 3.4105
R12962 GNDA.n3252 GNDA.n3251 3.4105
R12963 GNDA.n3250 GNDA.n594 3.4105
R12964 GNDA.n3203 GNDA.n3180 3.4105
R12965 GNDA.n3205 GNDA.n3179 3.4105
R12966 GNDA.n3206 GNDA.n3178 3.4105
R12967 GNDA.n3208 GNDA.n3177 3.4105
R12968 GNDA.n3209 GNDA.n3176 3.4105
R12969 GNDA.n3211 GNDA.n3175 3.4105
R12970 GNDA.n3212 GNDA.n3174 3.4105
R12971 GNDA.n3214 GNDA.n3173 3.4105
R12972 GNDA.n3215 GNDA.n3172 3.4105
R12973 GNDA.n3217 GNDA.n3171 3.4105
R12974 GNDA.n3218 GNDA.n3170 3.4105
R12975 GNDA.n3220 GNDA.n3169 3.4105
R12976 GNDA.n3221 GNDA.n3168 3.4105
R12977 GNDA.n3223 GNDA.n3167 3.4105
R12978 GNDA.n3224 GNDA.n3166 3.4105
R12979 GNDA.n3226 GNDA.n3165 3.4105
R12980 GNDA.n3227 GNDA.n3164 3.4105
R12981 GNDA.n3229 GNDA.n3163 3.4105
R12982 GNDA.n3230 GNDA.n3162 3.4105
R12983 GNDA.n3232 GNDA.n3161 3.4105
R12984 GNDA.n3233 GNDA.n3160 3.4105
R12985 GNDA.n3235 GNDA.n3159 3.4105
R12986 GNDA.n3237 GNDA.n3236 3.4105
R12987 GNDA.n1588 GNDA.n1587 3.4105
R12988 GNDA.n1652 GNDA.n1651 3.4105
R12989 GNDA.n1650 GNDA.n1649 3.4105
R12990 GNDA.n1648 GNDA.n1647 3.4105
R12991 GNDA.n1646 GNDA.n1590 3.4105
R12992 GNDA.n1642 GNDA.n1641 3.4105
R12993 GNDA.n1640 GNDA.n1639 3.4105
R12994 GNDA.n1638 GNDA.n1637 3.4105
R12995 GNDA.n1636 GNDA.n1592 3.4105
R12996 GNDA.n1632 GNDA.n1631 3.4105
R12997 GNDA.n1630 GNDA.n1629 3.4105
R12998 GNDA.n1628 GNDA.n1627 3.4105
R12999 GNDA.n1626 GNDA.n1594 3.4105
R13000 GNDA.n1622 GNDA.n1621 3.4105
R13001 GNDA.n1620 GNDA.n1619 3.4105
R13002 GNDA.n1618 GNDA.n1617 3.4105
R13003 GNDA.n1616 GNDA.n1596 3.4105
R13004 GNDA.n1612 GNDA.n1611 3.4105
R13005 GNDA.n1610 GNDA.n1609 3.4105
R13006 GNDA.n1608 GNDA.n1607 3.4105
R13007 GNDA.n1606 GNDA.n1598 3.4105
R13008 GNDA.n1602 GNDA.n1601 3.4105
R13009 GNDA.n1600 GNDA.n1575 3.4105
R13010 GNDA.n1506 GNDA.n1505 3.4105
R13011 GNDA.n1570 GNDA.n1569 3.4105
R13012 GNDA.n1568 GNDA.n1567 3.4105
R13013 GNDA.n1566 GNDA.n1565 3.4105
R13014 GNDA.n1564 GNDA.n1508 3.4105
R13015 GNDA.n1560 GNDA.n1559 3.4105
R13016 GNDA.n1558 GNDA.n1557 3.4105
R13017 GNDA.n1556 GNDA.n1555 3.4105
R13018 GNDA.n1554 GNDA.n1510 3.4105
R13019 GNDA.n1550 GNDA.n1549 3.4105
R13020 GNDA.n1548 GNDA.n1547 3.4105
R13021 GNDA.n1546 GNDA.n1545 3.4105
R13022 GNDA.n1544 GNDA.n1512 3.4105
R13023 GNDA.n1540 GNDA.n1539 3.4105
R13024 GNDA.n1538 GNDA.n1537 3.4105
R13025 GNDA.n1536 GNDA.n1535 3.4105
R13026 GNDA.n1534 GNDA.n1514 3.4105
R13027 GNDA.n1530 GNDA.n1529 3.4105
R13028 GNDA.n1528 GNDA.n1527 3.4105
R13029 GNDA.n1526 GNDA.n1525 3.4105
R13030 GNDA.n1524 GNDA.n1516 3.4105
R13031 GNDA.n1520 GNDA.n1519 3.4105
R13032 GNDA.n1518 GNDA.n1493 3.4105
R13033 GNDA.n1424 GNDA.n1423 3.4105
R13034 GNDA.n1488 GNDA.n1487 3.4105
R13035 GNDA.n1486 GNDA.n1485 3.4105
R13036 GNDA.n1484 GNDA.n1483 3.4105
R13037 GNDA.n1482 GNDA.n1426 3.4105
R13038 GNDA.n1478 GNDA.n1477 3.4105
R13039 GNDA.n1476 GNDA.n1475 3.4105
R13040 GNDA.n1474 GNDA.n1473 3.4105
R13041 GNDA.n1472 GNDA.n1428 3.4105
R13042 GNDA.n1468 GNDA.n1467 3.4105
R13043 GNDA.n1466 GNDA.n1465 3.4105
R13044 GNDA.n1464 GNDA.n1463 3.4105
R13045 GNDA.n1462 GNDA.n1430 3.4105
R13046 GNDA.n1458 GNDA.n1457 3.4105
R13047 GNDA.n1456 GNDA.n1455 3.4105
R13048 GNDA.n1454 GNDA.n1453 3.4105
R13049 GNDA.n1452 GNDA.n1432 3.4105
R13050 GNDA.n1448 GNDA.n1447 3.4105
R13051 GNDA.n1446 GNDA.n1445 3.4105
R13052 GNDA.n1444 GNDA.n1443 3.4105
R13053 GNDA.n1442 GNDA.n1434 3.4105
R13054 GNDA.n1438 GNDA.n1437 3.4105
R13055 GNDA.n1436 GNDA.n1411 3.4105
R13056 GNDA.n1214 GNDA.n1191 3.4105
R13057 GNDA.n1216 GNDA.n1190 3.4105
R13058 GNDA.n1217 GNDA.n1189 3.4105
R13059 GNDA.n1219 GNDA.n1188 3.4105
R13060 GNDA.n1220 GNDA.n1187 3.4105
R13061 GNDA.n1222 GNDA.n1186 3.4105
R13062 GNDA.n1223 GNDA.n1185 3.4105
R13063 GNDA.n1225 GNDA.n1184 3.4105
R13064 GNDA.n1226 GNDA.n1183 3.4105
R13065 GNDA.n1228 GNDA.n1182 3.4105
R13066 GNDA.n1229 GNDA.n1181 3.4105
R13067 GNDA.n1231 GNDA.n1180 3.4105
R13068 GNDA.n1232 GNDA.n1179 3.4105
R13069 GNDA.n1234 GNDA.n1178 3.4105
R13070 GNDA.n1235 GNDA.n1177 3.4105
R13071 GNDA.n1237 GNDA.n1176 3.4105
R13072 GNDA.n1238 GNDA.n1175 3.4105
R13073 GNDA.n1240 GNDA.n1174 3.4105
R13074 GNDA.n1241 GNDA.n1173 3.4105
R13075 GNDA.n1243 GNDA.n1172 3.4105
R13076 GNDA.n1244 GNDA.n1171 3.4105
R13077 GNDA.n1246 GNDA.n1170 3.4105
R13078 GNDA.n1248 GNDA.n1247 3.4105
R13079 GNDA.n1155 GNDA.n1154 3.4105
R13080 GNDA.n1920 GNDA.n1919 3.4105
R13081 GNDA.n1918 GNDA.n1917 3.4105
R13082 GNDA.n1916 GNDA.n1915 3.4105
R13083 GNDA.n1914 GNDA.n1157 3.4105
R13084 GNDA.n1910 GNDA.n1909 3.4105
R13085 GNDA.n1908 GNDA.n1907 3.4105
R13086 GNDA.n1906 GNDA.n1905 3.4105
R13087 GNDA.n1904 GNDA.n1159 3.4105
R13088 GNDA.n1900 GNDA.n1899 3.4105
R13089 GNDA.n1898 GNDA.n1897 3.4105
R13090 GNDA.n1896 GNDA.n1895 3.4105
R13091 GNDA.n1894 GNDA.n1161 3.4105
R13092 GNDA.n1890 GNDA.n1889 3.4105
R13093 GNDA.n1888 GNDA.n1887 3.4105
R13094 GNDA.n1886 GNDA.n1885 3.4105
R13095 GNDA.n1884 GNDA.n1163 3.4105
R13096 GNDA.n1880 GNDA.n1879 3.4105
R13097 GNDA.n1878 GNDA.n1877 3.4105
R13098 GNDA.n1876 GNDA.n1875 3.4105
R13099 GNDA.n1874 GNDA.n1165 3.4105
R13100 GNDA.n1870 GNDA.n1869 3.4105
R13101 GNDA.n1868 GNDA.n1141 3.4105
R13102 GNDA.n1924 GNDA.n1141 3.4105
R13103 GNDA.n1924 GNDA.n1923 3.4105
R13104 GNDA.n1247 GNDA.n1153 3.4105
R13105 GNDA.n1213 GNDA.n1153 3.4105
R13106 GNDA.n1492 GNDA.n1411 3.4105
R13107 GNDA.n1492 GNDA.n1491 3.4105
R13108 GNDA.n1574 GNDA.n1493 3.4105
R13109 GNDA.n1574 GNDA.n1573 3.4105
R13110 GNDA.n1656 GNDA.n1575 3.4105
R13111 GNDA.n1656 GNDA.n1655 3.4105
R13112 GNDA.n3236 GNDA.n593 3.4105
R13113 GNDA.n3202 GNDA.n593 3.4105
R13114 GNDA.n3306 GNDA.n594 3.4105
R13115 GNDA.n3306 GNDA.n3305 3.4105
R13116 GNDA.n3470 GNDA.n553 3.4105
R13117 GNDA.n3436 GNDA.n553 3.4105
R13118 GNDA.n3540 GNDA.n554 3.4105
R13119 GNDA.n3540 GNDA.n3539 3.4105
R13120 GNDA.n3617 GNDA.n3616 3.4105
R13121 GNDA.n3616 GNDA.n3615 3.4105
R13122 GNDA.n3774 GNDA.n514 3.4105
R13123 GNDA.n3774 GNDA.n3773 3.4105
R13124 GNDA.n3851 GNDA.n3850 3.4105
R13125 GNDA.n3850 GNDA.n3849 3.4105
R13126 GNDA.n1733 GNDA.n1732 3.4105
R13127 GNDA.n1732 GNDA.n1731 3.4105
R13128 GNDA.n3941 GNDA.n477 3.4105
R13129 GNDA.n3907 GNDA.n477 3.4105
R13130 GNDA.n4093 GNDA.n4012 3.4105
R13131 GNDA.n4093 GNDA.n4092 3.4105
R13132 GNDA.n4175 GNDA.n4094 3.4105
R13133 GNDA.n4175 GNDA.n4174 3.4105
R13134 GNDA.n4011 GNDA.n478 3.4105
R13135 GNDA.n4011 GNDA.n4010 3.4105
R13136 GNDA.n4257 GNDA.n4176 3.4105
R13137 GNDA.n4257 GNDA.n4256 3.4105
R13138 GNDA.n4339 GNDA.n4258 3.4105
R13139 GNDA.n4339 GNDA.n4338 3.4105
R13140 GNDA.n4421 GNDA.n4340 3.4105
R13141 GNDA.n4421 GNDA.n4420 3.4105
R13142 GNDA.n4503 GNDA.n4422 3.4105
R13143 GNDA.n4503 GNDA.n4502 3.4105
R13144 GNDA.n4580 GNDA.n4579 3.4105
R13145 GNDA.n4579 GNDA.n4578 3.4105
R13146 GNDA.n3383 GNDA.n3382 3.4105
R13147 GNDA.n3382 GNDA.n3381 3.4105
R13148 GNDA.n3627 GNDA.n513 3.4105
R13149 GNDA.n3671 GNDA.n513 3.4105
R13150 GNDA.n1807 GNDA.n1805 3.4105
R13151 GNDA.n1808 GNDA.n1804 3.4105
R13152 GNDA.n1809 GNDA.n1803 3.4105
R13153 GNDA.n1802 GNDA.n1800 3.4105
R13154 GNDA.n1813 GNDA.n1799 3.4105
R13155 GNDA.n1814 GNDA.n1798 3.4105
R13156 GNDA.n1815 GNDA.n1797 3.4105
R13157 GNDA.n1796 GNDA.n1794 3.4105
R13158 GNDA.n1819 GNDA.n1793 3.4105
R13159 GNDA.n1820 GNDA.n1792 3.4105
R13160 GNDA.n1821 GNDA.n1791 3.4105
R13161 GNDA.n1790 GNDA.n1788 3.4105
R13162 GNDA.n1825 GNDA.n1787 3.4105
R13163 GNDA.n1826 GNDA.n1786 3.4105
R13164 GNDA.n1827 GNDA.n1785 3.4105
R13165 GNDA.n1784 GNDA.n1782 3.4105
R13166 GNDA.n1831 GNDA.n1781 3.4105
R13167 GNDA.n1832 GNDA.n1780 3.4105
R13168 GNDA.n1833 GNDA.n1779 3.4105
R13169 GNDA.n1778 GNDA.n1776 3.4105
R13170 GNDA.n1837 GNDA.n1775 3.4105
R13171 GNDA.n1838 GNDA.n1774 3.4105
R13172 GNDA.n2141 GNDA.n2140 3.4105
R13173 GNDA.n2203 GNDA.n2202 3.4105
R13174 GNDA.n2201 GNDA.n2200 3.4105
R13175 GNDA.n2199 GNDA.n2145 3.4105
R13176 GNDA.n2144 GNDA.n2143 3.4105
R13177 GNDA.n2195 GNDA.n2194 3.4105
R13178 GNDA.n2193 GNDA.n2192 3.4105
R13179 GNDA.n2191 GNDA.n2149 3.4105
R13180 GNDA.n2148 GNDA.n2147 3.4105
R13181 GNDA.n2187 GNDA.n2186 3.4105
R13182 GNDA.n2185 GNDA.n2184 3.4105
R13183 GNDA.n2183 GNDA.n2153 3.4105
R13184 GNDA.n2152 GNDA.n2151 3.4105
R13185 GNDA.n2179 GNDA.n2178 3.4105
R13186 GNDA.n2177 GNDA.n2176 3.4105
R13187 GNDA.n2175 GNDA.n2157 3.4105
R13188 GNDA.n2156 GNDA.n2155 3.4105
R13189 GNDA.n2171 GNDA.n2170 3.4105
R13190 GNDA.n2169 GNDA.n2168 3.4105
R13191 GNDA.n2167 GNDA.n2161 3.4105
R13192 GNDA.n2160 GNDA.n2159 3.4105
R13193 GNDA.n2163 GNDA.n2162 3.4105
R13194 GNDA.n2220 GNDA.n2219 3.4105
R13195 GNDA.n845 GNDA.n844 3.4105
R13196 GNDA.n2126 GNDA.n2125 3.4105
R13197 GNDA.n2065 GNDA.n2064 3.4105
R13198 GNDA.n2121 GNDA.n2120 3.4105
R13199 GNDA.n2119 GNDA.n2118 3.4105
R13200 GNDA.n2117 GNDA.n2116 3.4105
R13201 GNDA.n2115 GNDA.n2067 3.4105
R13202 GNDA.n2111 GNDA.n2110 3.4105
R13203 GNDA.n2109 GNDA.n2108 3.4105
R13204 GNDA.n2107 GNDA.n2106 3.4105
R13205 GNDA.n2105 GNDA.n2069 3.4105
R13206 GNDA.n2101 GNDA.n2100 3.4105
R13207 GNDA.n2099 GNDA.n2098 3.4105
R13208 GNDA.n2097 GNDA.n2096 3.4105
R13209 GNDA.n2095 GNDA.n2071 3.4105
R13210 GNDA.n2091 GNDA.n2090 3.4105
R13211 GNDA.n2089 GNDA.n2088 3.4105
R13212 GNDA.n2087 GNDA.n2086 3.4105
R13213 GNDA.n2085 GNDA.n2073 3.4105
R13214 GNDA.n2081 GNDA.n2080 3.4105
R13215 GNDA.n2079 GNDA.n2078 3.4105
R13216 GNDA.n2077 GNDA.n2076 3.4105
R13217 GNDA.n2224 GNDA.n2223 3.4105
R13218 GNDA.n2222 GNDA.n2053 3.4105
R13219 GNDA.n2223 GNDA.n2222 3.4105
R13220 GNDA.n2221 GNDA.n2128 3.4105
R13221 GNDA.n2221 GNDA.n2220 3.4105
R13222 GNDA.n2050 GNDA.n880 3.4105
R13223 GNDA.n2050 GNDA.n2049 3.4105
R13224 GNDA.n2049 GNDA.n863 3.4105
R13225 GNDA.n899 GNDA.n880 3.4105
R13226 GNDA.n2017 GNDA.n899 3.4105
R13227 GNDA.n945 GNDA.n899 3.4105
R13228 GNDA.n2019 GNDA.n899 3.4105
R13229 GNDA.n944 GNDA.n899 3.4105
R13230 GNDA.n2021 GNDA.n899 3.4105
R13231 GNDA.n943 GNDA.n899 3.4105
R13232 GNDA.n2023 GNDA.n899 3.4105
R13233 GNDA.n942 GNDA.n899 3.4105
R13234 GNDA.n2025 GNDA.n899 3.4105
R13235 GNDA.n941 GNDA.n899 3.4105
R13236 GNDA.n2027 GNDA.n899 3.4105
R13237 GNDA.n940 GNDA.n899 3.4105
R13238 GNDA.n2029 GNDA.n899 3.4105
R13239 GNDA.n939 GNDA.n899 3.4105
R13240 GNDA.n2031 GNDA.n899 3.4105
R13241 GNDA.n938 GNDA.n899 3.4105
R13242 GNDA.n2033 GNDA.n899 3.4105
R13243 GNDA.n937 GNDA.n899 3.4105
R13244 GNDA.n2035 GNDA.n899 3.4105
R13245 GNDA.n936 GNDA.n899 3.4105
R13246 GNDA.n2037 GNDA.n899 3.4105
R13247 GNDA.n935 GNDA.n899 3.4105
R13248 GNDA.n2039 GNDA.n899 3.4105
R13249 GNDA.n934 GNDA.n899 3.4105
R13250 GNDA.n2041 GNDA.n899 3.4105
R13251 GNDA.n933 GNDA.n899 3.4105
R13252 GNDA.n2043 GNDA.n899 3.4105
R13253 GNDA.n932 GNDA.n899 3.4105
R13254 GNDA.n2045 GNDA.n899 3.4105
R13255 GNDA.n931 GNDA.n899 3.4105
R13256 GNDA.n2047 GNDA.n899 3.4105
R13257 GNDA.n2049 GNDA.n899 3.4105
R13258 GNDA.n896 GNDA.n880 3.4105
R13259 GNDA.n2017 GNDA.n896 3.4105
R13260 GNDA.n945 GNDA.n896 3.4105
R13261 GNDA.n2019 GNDA.n896 3.4105
R13262 GNDA.n944 GNDA.n896 3.4105
R13263 GNDA.n2021 GNDA.n896 3.4105
R13264 GNDA.n943 GNDA.n896 3.4105
R13265 GNDA.n2023 GNDA.n896 3.4105
R13266 GNDA.n942 GNDA.n896 3.4105
R13267 GNDA.n2025 GNDA.n896 3.4105
R13268 GNDA.n941 GNDA.n896 3.4105
R13269 GNDA.n2027 GNDA.n896 3.4105
R13270 GNDA.n940 GNDA.n896 3.4105
R13271 GNDA.n2029 GNDA.n896 3.4105
R13272 GNDA.n939 GNDA.n896 3.4105
R13273 GNDA.n2031 GNDA.n896 3.4105
R13274 GNDA.n938 GNDA.n896 3.4105
R13275 GNDA.n2033 GNDA.n896 3.4105
R13276 GNDA.n937 GNDA.n896 3.4105
R13277 GNDA.n2035 GNDA.n896 3.4105
R13278 GNDA.n936 GNDA.n896 3.4105
R13279 GNDA.n2037 GNDA.n896 3.4105
R13280 GNDA.n935 GNDA.n896 3.4105
R13281 GNDA.n2039 GNDA.n896 3.4105
R13282 GNDA.n934 GNDA.n896 3.4105
R13283 GNDA.n2041 GNDA.n896 3.4105
R13284 GNDA.n933 GNDA.n896 3.4105
R13285 GNDA.n2043 GNDA.n896 3.4105
R13286 GNDA.n932 GNDA.n896 3.4105
R13287 GNDA.n2045 GNDA.n896 3.4105
R13288 GNDA.n931 GNDA.n896 3.4105
R13289 GNDA.n2047 GNDA.n896 3.4105
R13290 GNDA.n2049 GNDA.n896 3.4105
R13291 GNDA.n901 GNDA.n880 3.4105
R13292 GNDA.n2017 GNDA.n901 3.4105
R13293 GNDA.n945 GNDA.n901 3.4105
R13294 GNDA.n2019 GNDA.n901 3.4105
R13295 GNDA.n944 GNDA.n901 3.4105
R13296 GNDA.n2021 GNDA.n901 3.4105
R13297 GNDA.n943 GNDA.n901 3.4105
R13298 GNDA.n2023 GNDA.n901 3.4105
R13299 GNDA.n942 GNDA.n901 3.4105
R13300 GNDA.n2025 GNDA.n901 3.4105
R13301 GNDA.n941 GNDA.n901 3.4105
R13302 GNDA.n2027 GNDA.n901 3.4105
R13303 GNDA.n940 GNDA.n901 3.4105
R13304 GNDA.n2029 GNDA.n901 3.4105
R13305 GNDA.n939 GNDA.n901 3.4105
R13306 GNDA.n2031 GNDA.n901 3.4105
R13307 GNDA.n938 GNDA.n901 3.4105
R13308 GNDA.n2033 GNDA.n901 3.4105
R13309 GNDA.n937 GNDA.n901 3.4105
R13310 GNDA.n2035 GNDA.n901 3.4105
R13311 GNDA.n936 GNDA.n901 3.4105
R13312 GNDA.n2037 GNDA.n901 3.4105
R13313 GNDA.n935 GNDA.n901 3.4105
R13314 GNDA.n2039 GNDA.n901 3.4105
R13315 GNDA.n934 GNDA.n901 3.4105
R13316 GNDA.n2041 GNDA.n901 3.4105
R13317 GNDA.n933 GNDA.n901 3.4105
R13318 GNDA.n2043 GNDA.n901 3.4105
R13319 GNDA.n932 GNDA.n901 3.4105
R13320 GNDA.n2045 GNDA.n901 3.4105
R13321 GNDA.n931 GNDA.n901 3.4105
R13322 GNDA.n2047 GNDA.n901 3.4105
R13323 GNDA.n2049 GNDA.n901 3.4105
R13324 GNDA.n895 GNDA.n880 3.4105
R13325 GNDA.n2017 GNDA.n895 3.4105
R13326 GNDA.n945 GNDA.n895 3.4105
R13327 GNDA.n2019 GNDA.n895 3.4105
R13328 GNDA.n944 GNDA.n895 3.4105
R13329 GNDA.n2021 GNDA.n895 3.4105
R13330 GNDA.n943 GNDA.n895 3.4105
R13331 GNDA.n2023 GNDA.n895 3.4105
R13332 GNDA.n942 GNDA.n895 3.4105
R13333 GNDA.n2025 GNDA.n895 3.4105
R13334 GNDA.n941 GNDA.n895 3.4105
R13335 GNDA.n2027 GNDA.n895 3.4105
R13336 GNDA.n940 GNDA.n895 3.4105
R13337 GNDA.n2029 GNDA.n895 3.4105
R13338 GNDA.n939 GNDA.n895 3.4105
R13339 GNDA.n2031 GNDA.n895 3.4105
R13340 GNDA.n938 GNDA.n895 3.4105
R13341 GNDA.n2033 GNDA.n895 3.4105
R13342 GNDA.n937 GNDA.n895 3.4105
R13343 GNDA.n2035 GNDA.n895 3.4105
R13344 GNDA.n936 GNDA.n895 3.4105
R13345 GNDA.n2037 GNDA.n895 3.4105
R13346 GNDA.n935 GNDA.n895 3.4105
R13347 GNDA.n2039 GNDA.n895 3.4105
R13348 GNDA.n934 GNDA.n895 3.4105
R13349 GNDA.n2041 GNDA.n895 3.4105
R13350 GNDA.n933 GNDA.n895 3.4105
R13351 GNDA.n2043 GNDA.n895 3.4105
R13352 GNDA.n932 GNDA.n895 3.4105
R13353 GNDA.n2045 GNDA.n895 3.4105
R13354 GNDA.n931 GNDA.n895 3.4105
R13355 GNDA.n2047 GNDA.n895 3.4105
R13356 GNDA.n2049 GNDA.n895 3.4105
R13357 GNDA.n903 GNDA.n880 3.4105
R13358 GNDA.n2017 GNDA.n903 3.4105
R13359 GNDA.n945 GNDA.n903 3.4105
R13360 GNDA.n2019 GNDA.n903 3.4105
R13361 GNDA.n944 GNDA.n903 3.4105
R13362 GNDA.n2021 GNDA.n903 3.4105
R13363 GNDA.n943 GNDA.n903 3.4105
R13364 GNDA.n2023 GNDA.n903 3.4105
R13365 GNDA.n942 GNDA.n903 3.4105
R13366 GNDA.n2025 GNDA.n903 3.4105
R13367 GNDA.n941 GNDA.n903 3.4105
R13368 GNDA.n2027 GNDA.n903 3.4105
R13369 GNDA.n940 GNDA.n903 3.4105
R13370 GNDA.n2029 GNDA.n903 3.4105
R13371 GNDA.n939 GNDA.n903 3.4105
R13372 GNDA.n2031 GNDA.n903 3.4105
R13373 GNDA.n938 GNDA.n903 3.4105
R13374 GNDA.n2033 GNDA.n903 3.4105
R13375 GNDA.n937 GNDA.n903 3.4105
R13376 GNDA.n2035 GNDA.n903 3.4105
R13377 GNDA.n936 GNDA.n903 3.4105
R13378 GNDA.n2037 GNDA.n903 3.4105
R13379 GNDA.n935 GNDA.n903 3.4105
R13380 GNDA.n2039 GNDA.n903 3.4105
R13381 GNDA.n934 GNDA.n903 3.4105
R13382 GNDA.n2041 GNDA.n903 3.4105
R13383 GNDA.n933 GNDA.n903 3.4105
R13384 GNDA.n2043 GNDA.n903 3.4105
R13385 GNDA.n932 GNDA.n903 3.4105
R13386 GNDA.n2045 GNDA.n903 3.4105
R13387 GNDA.n931 GNDA.n903 3.4105
R13388 GNDA.n2047 GNDA.n903 3.4105
R13389 GNDA.n2049 GNDA.n903 3.4105
R13390 GNDA.n894 GNDA.n880 3.4105
R13391 GNDA.n2017 GNDA.n894 3.4105
R13392 GNDA.n945 GNDA.n894 3.4105
R13393 GNDA.n2019 GNDA.n894 3.4105
R13394 GNDA.n944 GNDA.n894 3.4105
R13395 GNDA.n2021 GNDA.n894 3.4105
R13396 GNDA.n943 GNDA.n894 3.4105
R13397 GNDA.n2023 GNDA.n894 3.4105
R13398 GNDA.n942 GNDA.n894 3.4105
R13399 GNDA.n2025 GNDA.n894 3.4105
R13400 GNDA.n941 GNDA.n894 3.4105
R13401 GNDA.n2027 GNDA.n894 3.4105
R13402 GNDA.n940 GNDA.n894 3.4105
R13403 GNDA.n2029 GNDA.n894 3.4105
R13404 GNDA.n939 GNDA.n894 3.4105
R13405 GNDA.n2031 GNDA.n894 3.4105
R13406 GNDA.n938 GNDA.n894 3.4105
R13407 GNDA.n2033 GNDA.n894 3.4105
R13408 GNDA.n937 GNDA.n894 3.4105
R13409 GNDA.n2035 GNDA.n894 3.4105
R13410 GNDA.n936 GNDA.n894 3.4105
R13411 GNDA.n2037 GNDA.n894 3.4105
R13412 GNDA.n935 GNDA.n894 3.4105
R13413 GNDA.n2039 GNDA.n894 3.4105
R13414 GNDA.n934 GNDA.n894 3.4105
R13415 GNDA.n2041 GNDA.n894 3.4105
R13416 GNDA.n933 GNDA.n894 3.4105
R13417 GNDA.n2043 GNDA.n894 3.4105
R13418 GNDA.n932 GNDA.n894 3.4105
R13419 GNDA.n2045 GNDA.n894 3.4105
R13420 GNDA.n931 GNDA.n894 3.4105
R13421 GNDA.n2047 GNDA.n894 3.4105
R13422 GNDA.n2049 GNDA.n894 3.4105
R13423 GNDA.n905 GNDA.n880 3.4105
R13424 GNDA.n2017 GNDA.n905 3.4105
R13425 GNDA.n945 GNDA.n905 3.4105
R13426 GNDA.n2019 GNDA.n905 3.4105
R13427 GNDA.n944 GNDA.n905 3.4105
R13428 GNDA.n2021 GNDA.n905 3.4105
R13429 GNDA.n943 GNDA.n905 3.4105
R13430 GNDA.n2023 GNDA.n905 3.4105
R13431 GNDA.n942 GNDA.n905 3.4105
R13432 GNDA.n2025 GNDA.n905 3.4105
R13433 GNDA.n941 GNDA.n905 3.4105
R13434 GNDA.n2027 GNDA.n905 3.4105
R13435 GNDA.n940 GNDA.n905 3.4105
R13436 GNDA.n2029 GNDA.n905 3.4105
R13437 GNDA.n939 GNDA.n905 3.4105
R13438 GNDA.n2031 GNDA.n905 3.4105
R13439 GNDA.n938 GNDA.n905 3.4105
R13440 GNDA.n2033 GNDA.n905 3.4105
R13441 GNDA.n937 GNDA.n905 3.4105
R13442 GNDA.n2035 GNDA.n905 3.4105
R13443 GNDA.n936 GNDA.n905 3.4105
R13444 GNDA.n2037 GNDA.n905 3.4105
R13445 GNDA.n935 GNDA.n905 3.4105
R13446 GNDA.n2039 GNDA.n905 3.4105
R13447 GNDA.n934 GNDA.n905 3.4105
R13448 GNDA.n2041 GNDA.n905 3.4105
R13449 GNDA.n933 GNDA.n905 3.4105
R13450 GNDA.n2043 GNDA.n905 3.4105
R13451 GNDA.n932 GNDA.n905 3.4105
R13452 GNDA.n2045 GNDA.n905 3.4105
R13453 GNDA.n931 GNDA.n905 3.4105
R13454 GNDA.n2047 GNDA.n905 3.4105
R13455 GNDA.n2049 GNDA.n905 3.4105
R13456 GNDA.n893 GNDA.n880 3.4105
R13457 GNDA.n2017 GNDA.n893 3.4105
R13458 GNDA.n945 GNDA.n893 3.4105
R13459 GNDA.n2019 GNDA.n893 3.4105
R13460 GNDA.n944 GNDA.n893 3.4105
R13461 GNDA.n2021 GNDA.n893 3.4105
R13462 GNDA.n943 GNDA.n893 3.4105
R13463 GNDA.n2023 GNDA.n893 3.4105
R13464 GNDA.n942 GNDA.n893 3.4105
R13465 GNDA.n2025 GNDA.n893 3.4105
R13466 GNDA.n941 GNDA.n893 3.4105
R13467 GNDA.n2027 GNDA.n893 3.4105
R13468 GNDA.n940 GNDA.n893 3.4105
R13469 GNDA.n2029 GNDA.n893 3.4105
R13470 GNDA.n939 GNDA.n893 3.4105
R13471 GNDA.n2031 GNDA.n893 3.4105
R13472 GNDA.n938 GNDA.n893 3.4105
R13473 GNDA.n2033 GNDA.n893 3.4105
R13474 GNDA.n937 GNDA.n893 3.4105
R13475 GNDA.n2035 GNDA.n893 3.4105
R13476 GNDA.n936 GNDA.n893 3.4105
R13477 GNDA.n2037 GNDA.n893 3.4105
R13478 GNDA.n935 GNDA.n893 3.4105
R13479 GNDA.n2039 GNDA.n893 3.4105
R13480 GNDA.n934 GNDA.n893 3.4105
R13481 GNDA.n2041 GNDA.n893 3.4105
R13482 GNDA.n933 GNDA.n893 3.4105
R13483 GNDA.n2043 GNDA.n893 3.4105
R13484 GNDA.n932 GNDA.n893 3.4105
R13485 GNDA.n2045 GNDA.n893 3.4105
R13486 GNDA.n931 GNDA.n893 3.4105
R13487 GNDA.n2047 GNDA.n893 3.4105
R13488 GNDA.n2049 GNDA.n893 3.4105
R13489 GNDA.n907 GNDA.n880 3.4105
R13490 GNDA.n2017 GNDA.n907 3.4105
R13491 GNDA.n945 GNDA.n907 3.4105
R13492 GNDA.n2019 GNDA.n907 3.4105
R13493 GNDA.n944 GNDA.n907 3.4105
R13494 GNDA.n2021 GNDA.n907 3.4105
R13495 GNDA.n943 GNDA.n907 3.4105
R13496 GNDA.n2023 GNDA.n907 3.4105
R13497 GNDA.n942 GNDA.n907 3.4105
R13498 GNDA.n2025 GNDA.n907 3.4105
R13499 GNDA.n941 GNDA.n907 3.4105
R13500 GNDA.n2027 GNDA.n907 3.4105
R13501 GNDA.n940 GNDA.n907 3.4105
R13502 GNDA.n2029 GNDA.n907 3.4105
R13503 GNDA.n939 GNDA.n907 3.4105
R13504 GNDA.n2031 GNDA.n907 3.4105
R13505 GNDA.n938 GNDA.n907 3.4105
R13506 GNDA.n2033 GNDA.n907 3.4105
R13507 GNDA.n937 GNDA.n907 3.4105
R13508 GNDA.n2035 GNDA.n907 3.4105
R13509 GNDA.n936 GNDA.n907 3.4105
R13510 GNDA.n2037 GNDA.n907 3.4105
R13511 GNDA.n935 GNDA.n907 3.4105
R13512 GNDA.n2039 GNDA.n907 3.4105
R13513 GNDA.n934 GNDA.n907 3.4105
R13514 GNDA.n2041 GNDA.n907 3.4105
R13515 GNDA.n933 GNDA.n907 3.4105
R13516 GNDA.n2043 GNDA.n907 3.4105
R13517 GNDA.n932 GNDA.n907 3.4105
R13518 GNDA.n2045 GNDA.n907 3.4105
R13519 GNDA.n931 GNDA.n907 3.4105
R13520 GNDA.n2047 GNDA.n907 3.4105
R13521 GNDA.n2049 GNDA.n907 3.4105
R13522 GNDA.n892 GNDA.n880 3.4105
R13523 GNDA.n2017 GNDA.n892 3.4105
R13524 GNDA.n945 GNDA.n892 3.4105
R13525 GNDA.n2019 GNDA.n892 3.4105
R13526 GNDA.n944 GNDA.n892 3.4105
R13527 GNDA.n2021 GNDA.n892 3.4105
R13528 GNDA.n943 GNDA.n892 3.4105
R13529 GNDA.n2023 GNDA.n892 3.4105
R13530 GNDA.n942 GNDA.n892 3.4105
R13531 GNDA.n2025 GNDA.n892 3.4105
R13532 GNDA.n941 GNDA.n892 3.4105
R13533 GNDA.n2027 GNDA.n892 3.4105
R13534 GNDA.n940 GNDA.n892 3.4105
R13535 GNDA.n2029 GNDA.n892 3.4105
R13536 GNDA.n939 GNDA.n892 3.4105
R13537 GNDA.n2031 GNDA.n892 3.4105
R13538 GNDA.n938 GNDA.n892 3.4105
R13539 GNDA.n2033 GNDA.n892 3.4105
R13540 GNDA.n937 GNDA.n892 3.4105
R13541 GNDA.n2035 GNDA.n892 3.4105
R13542 GNDA.n936 GNDA.n892 3.4105
R13543 GNDA.n2037 GNDA.n892 3.4105
R13544 GNDA.n935 GNDA.n892 3.4105
R13545 GNDA.n2039 GNDA.n892 3.4105
R13546 GNDA.n934 GNDA.n892 3.4105
R13547 GNDA.n2041 GNDA.n892 3.4105
R13548 GNDA.n933 GNDA.n892 3.4105
R13549 GNDA.n2043 GNDA.n892 3.4105
R13550 GNDA.n932 GNDA.n892 3.4105
R13551 GNDA.n2045 GNDA.n892 3.4105
R13552 GNDA.n931 GNDA.n892 3.4105
R13553 GNDA.n2047 GNDA.n892 3.4105
R13554 GNDA.n2049 GNDA.n892 3.4105
R13555 GNDA.n909 GNDA.n880 3.4105
R13556 GNDA.n2017 GNDA.n909 3.4105
R13557 GNDA.n945 GNDA.n909 3.4105
R13558 GNDA.n2019 GNDA.n909 3.4105
R13559 GNDA.n944 GNDA.n909 3.4105
R13560 GNDA.n2021 GNDA.n909 3.4105
R13561 GNDA.n943 GNDA.n909 3.4105
R13562 GNDA.n2023 GNDA.n909 3.4105
R13563 GNDA.n942 GNDA.n909 3.4105
R13564 GNDA.n2025 GNDA.n909 3.4105
R13565 GNDA.n941 GNDA.n909 3.4105
R13566 GNDA.n2027 GNDA.n909 3.4105
R13567 GNDA.n940 GNDA.n909 3.4105
R13568 GNDA.n2029 GNDA.n909 3.4105
R13569 GNDA.n939 GNDA.n909 3.4105
R13570 GNDA.n2031 GNDA.n909 3.4105
R13571 GNDA.n938 GNDA.n909 3.4105
R13572 GNDA.n2033 GNDA.n909 3.4105
R13573 GNDA.n937 GNDA.n909 3.4105
R13574 GNDA.n2035 GNDA.n909 3.4105
R13575 GNDA.n936 GNDA.n909 3.4105
R13576 GNDA.n2037 GNDA.n909 3.4105
R13577 GNDA.n935 GNDA.n909 3.4105
R13578 GNDA.n2039 GNDA.n909 3.4105
R13579 GNDA.n934 GNDA.n909 3.4105
R13580 GNDA.n2041 GNDA.n909 3.4105
R13581 GNDA.n933 GNDA.n909 3.4105
R13582 GNDA.n2043 GNDA.n909 3.4105
R13583 GNDA.n932 GNDA.n909 3.4105
R13584 GNDA.n2045 GNDA.n909 3.4105
R13585 GNDA.n931 GNDA.n909 3.4105
R13586 GNDA.n2047 GNDA.n909 3.4105
R13587 GNDA.n2049 GNDA.n909 3.4105
R13588 GNDA.n891 GNDA.n880 3.4105
R13589 GNDA.n2017 GNDA.n891 3.4105
R13590 GNDA.n945 GNDA.n891 3.4105
R13591 GNDA.n2019 GNDA.n891 3.4105
R13592 GNDA.n944 GNDA.n891 3.4105
R13593 GNDA.n2021 GNDA.n891 3.4105
R13594 GNDA.n943 GNDA.n891 3.4105
R13595 GNDA.n2023 GNDA.n891 3.4105
R13596 GNDA.n942 GNDA.n891 3.4105
R13597 GNDA.n2025 GNDA.n891 3.4105
R13598 GNDA.n941 GNDA.n891 3.4105
R13599 GNDA.n2027 GNDA.n891 3.4105
R13600 GNDA.n940 GNDA.n891 3.4105
R13601 GNDA.n2029 GNDA.n891 3.4105
R13602 GNDA.n939 GNDA.n891 3.4105
R13603 GNDA.n2031 GNDA.n891 3.4105
R13604 GNDA.n938 GNDA.n891 3.4105
R13605 GNDA.n2033 GNDA.n891 3.4105
R13606 GNDA.n937 GNDA.n891 3.4105
R13607 GNDA.n2035 GNDA.n891 3.4105
R13608 GNDA.n936 GNDA.n891 3.4105
R13609 GNDA.n2037 GNDA.n891 3.4105
R13610 GNDA.n935 GNDA.n891 3.4105
R13611 GNDA.n2039 GNDA.n891 3.4105
R13612 GNDA.n934 GNDA.n891 3.4105
R13613 GNDA.n2041 GNDA.n891 3.4105
R13614 GNDA.n933 GNDA.n891 3.4105
R13615 GNDA.n2043 GNDA.n891 3.4105
R13616 GNDA.n932 GNDA.n891 3.4105
R13617 GNDA.n2045 GNDA.n891 3.4105
R13618 GNDA.n931 GNDA.n891 3.4105
R13619 GNDA.n2047 GNDA.n891 3.4105
R13620 GNDA.n2049 GNDA.n891 3.4105
R13621 GNDA.n911 GNDA.n880 3.4105
R13622 GNDA.n2017 GNDA.n911 3.4105
R13623 GNDA.n945 GNDA.n911 3.4105
R13624 GNDA.n2019 GNDA.n911 3.4105
R13625 GNDA.n944 GNDA.n911 3.4105
R13626 GNDA.n2021 GNDA.n911 3.4105
R13627 GNDA.n943 GNDA.n911 3.4105
R13628 GNDA.n2023 GNDA.n911 3.4105
R13629 GNDA.n942 GNDA.n911 3.4105
R13630 GNDA.n2025 GNDA.n911 3.4105
R13631 GNDA.n941 GNDA.n911 3.4105
R13632 GNDA.n2027 GNDA.n911 3.4105
R13633 GNDA.n940 GNDA.n911 3.4105
R13634 GNDA.n2029 GNDA.n911 3.4105
R13635 GNDA.n939 GNDA.n911 3.4105
R13636 GNDA.n2031 GNDA.n911 3.4105
R13637 GNDA.n938 GNDA.n911 3.4105
R13638 GNDA.n2033 GNDA.n911 3.4105
R13639 GNDA.n937 GNDA.n911 3.4105
R13640 GNDA.n2035 GNDA.n911 3.4105
R13641 GNDA.n936 GNDA.n911 3.4105
R13642 GNDA.n2037 GNDA.n911 3.4105
R13643 GNDA.n935 GNDA.n911 3.4105
R13644 GNDA.n2039 GNDA.n911 3.4105
R13645 GNDA.n934 GNDA.n911 3.4105
R13646 GNDA.n2041 GNDA.n911 3.4105
R13647 GNDA.n933 GNDA.n911 3.4105
R13648 GNDA.n2043 GNDA.n911 3.4105
R13649 GNDA.n932 GNDA.n911 3.4105
R13650 GNDA.n2045 GNDA.n911 3.4105
R13651 GNDA.n931 GNDA.n911 3.4105
R13652 GNDA.n2047 GNDA.n911 3.4105
R13653 GNDA.n2049 GNDA.n911 3.4105
R13654 GNDA.n890 GNDA.n880 3.4105
R13655 GNDA.n2017 GNDA.n890 3.4105
R13656 GNDA.n945 GNDA.n890 3.4105
R13657 GNDA.n2019 GNDA.n890 3.4105
R13658 GNDA.n944 GNDA.n890 3.4105
R13659 GNDA.n2021 GNDA.n890 3.4105
R13660 GNDA.n943 GNDA.n890 3.4105
R13661 GNDA.n2023 GNDA.n890 3.4105
R13662 GNDA.n942 GNDA.n890 3.4105
R13663 GNDA.n2025 GNDA.n890 3.4105
R13664 GNDA.n941 GNDA.n890 3.4105
R13665 GNDA.n2027 GNDA.n890 3.4105
R13666 GNDA.n940 GNDA.n890 3.4105
R13667 GNDA.n2029 GNDA.n890 3.4105
R13668 GNDA.n939 GNDA.n890 3.4105
R13669 GNDA.n2031 GNDA.n890 3.4105
R13670 GNDA.n938 GNDA.n890 3.4105
R13671 GNDA.n2033 GNDA.n890 3.4105
R13672 GNDA.n937 GNDA.n890 3.4105
R13673 GNDA.n2035 GNDA.n890 3.4105
R13674 GNDA.n936 GNDA.n890 3.4105
R13675 GNDA.n2037 GNDA.n890 3.4105
R13676 GNDA.n935 GNDA.n890 3.4105
R13677 GNDA.n2039 GNDA.n890 3.4105
R13678 GNDA.n934 GNDA.n890 3.4105
R13679 GNDA.n2041 GNDA.n890 3.4105
R13680 GNDA.n933 GNDA.n890 3.4105
R13681 GNDA.n2043 GNDA.n890 3.4105
R13682 GNDA.n932 GNDA.n890 3.4105
R13683 GNDA.n2045 GNDA.n890 3.4105
R13684 GNDA.n931 GNDA.n890 3.4105
R13685 GNDA.n2047 GNDA.n890 3.4105
R13686 GNDA.n2049 GNDA.n890 3.4105
R13687 GNDA.n913 GNDA.n880 3.4105
R13688 GNDA.n2017 GNDA.n913 3.4105
R13689 GNDA.n945 GNDA.n913 3.4105
R13690 GNDA.n2019 GNDA.n913 3.4105
R13691 GNDA.n944 GNDA.n913 3.4105
R13692 GNDA.n2021 GNDA.n913 3.4105
R13693 GNDA.n943 GNDA.n913 3.4105
R13694 GNDA.n2023 GNDA.n913 3.4105
R13695 GNDA.n942 GNDA.n913 3.4105
R13696 GNDA.n2025 GNDA.n913 3.4105
R13697 GNDA.n941 GNDA.n913 3.4105
R13698 GNDA.n2027 GNDA.n913 3.4105
R13699 GNDA.n940 GNDA.n913 3.4105
R13700 GNDA.n2029 GNDA.n913 3.4105
R13701 GNDA.n939 GNDA.n913 3.4105
R13702 GNDA.n2031 GNDA.n913 3.4105
R13703 GNDA.n938 GNDA.n913 3.4105
R13704 GNDA.n2033 GNDA.n913 3.4105
R13705 GNDA.n937 GNDA.n913 3.4105
R13706 GNDA.n2035 GNDA.n913 3.4105
R13707 GNDA.n936 GNDA.n913 3.4105
R13708 GNDA.n2037 GNDA.n913 3.4105
R13709 GNDA.n935 GNDA.n913 3.4105
R13710 GNDA.n2039 GNDA.n913 3.4105
R13711 GNDA.n934 GNDA.n913 3.4105
R13712 GNDA.n2041 GNDA.n913 3.4105
R13713 GNDA.n933 GNDA.n913 3.4105
R13714 GNDA.n2043 GNDA.n913 3.4105
R13715 GNDA.n932 GNDA.n913 3.4105
R13716 GNDA.n2045 GNDA.n913 3.4105
R13717 GNDA.n931 GNDA.n913 3.4105
R13718 GNDA.n2047 GNDA.n913 3.4105
R13719 GNDA.n2049 GNDA.n913 3.4105
R13720 GNDA.n889 GNDA.n880 3.4105
R13721 GNDA.n2017 GNDA.n889 3.4105
R13722 GNDA.n945 GNDA.n889 3.4105
R13723 GNDA.n2019 GNDA.n889 3.4105
R13724 GNDA.n944 GNDA.n889 3.4105
R13725 GNDA.n2021 GNDA.n889 3.4105
R13726 GNDA.n943 GNDA.n889 3.4105
R13727 GNDA.n2023 GNDA.n889 3.4105
R13728 GNDA.n942 GNDA.n889 3.4105
R13729 GNDA.n2025 GNDA.n889 3.4105
R13730 GNDA.n941 GNDA.n889 3.4105
R13731 GNDA.n2027 GNDA.n889 3.4105
R13732 GNDA.n940 GNDA.n889 3.4105
R13733 GNDA.n2029 GNDA.n889 3.4105
R13734 GNDA.n939 GNDA.n889 3.4105
R13735 GNDA.n2031 GNDA.n889 3.4105
R13736 GNDA.n938 GNDA.n889 3.4105
R13737 GNDA.n2033 GNDA.n889 3.4105
R13738 GNDA.n937 GNDA.n889 3.4105
R13739 GNDA.n2035 GNDA.n889 3.4105
R13740 GNDA.n936 GNDA.n889 3.4105
R13741 GNDA.n2037 GNDA.n889 3.4105
R13742 GNDA.n935 GNDA.n889 3.4105
R13743 GNDA.n2039 GNDA.n889 3.4105
R13744 GNDA.n934 GNDA.n889 3.4105
R13745 GNDA.n2041 GNDA.n889 3.4105
R13746 GNDA.n933 GNDA.n889 3.4105
R13747 GNDA.n2043 GNDA.n889 3.4105
R13748 GNDA.n932 GNDA.n889 3.4105
R13749 GNDA.n2045 GNDA.n889 3.4105
R13750 GNDA.n931 GNDA.n889 3.4105
R13751 GNDA.n2047 GNDA.n889 3.4105
R13752 GNDA.n2049 GNDA.n889 3.4105
R13753 GNDA.n915 GNDA.n880 3.4105
R13754 GNDA.n2017 GNDA.n915 3.4105
R13755 GNDA.n945 GNDA.n915 3.4105
R13756 GNDA.n2019 GNDA.n915 3.4105
R13757 GNDA.n944 GNDA.n915 3.4105
R13758 GNDA.n2021 GNDA.n915 3.4105
R13759 GNDA.n943 GNDA.n915 3.4105
R13760 GNDA.n2023 GNDA.n915 3.4105
R13761 GNDA.n942 GNDA.n915 3.4105
R13762 GNDA.n2025 GNDA.n915 3.4105
R13763 GNDA.n941 GNDA.n915 3.4105
R13764 GNDA.n2027 GNDA.n915 3.4105
R13765 GNDA.n940 GNDA.n915 3.4105
R13766 GNDA.n2029 GNDA.n915 3.4105
R13767 GNDA.n939 GNDA.n915 3.4105
R13768 GNDA.n2031 GNDA.n915 3.4105
R13769 GNDA.n938 GNDA.n915 3.4105
R13770 GNDA.n2033 GNDA.n915 3.4105
R13771 GNDA.n937 GNDA.n915 3.4105
R13772 GNDA.n2035 GNDA.n915 3.4105
R13773 GNDA.n936 GNDA.n915 3.4105
R13774 GNDA.n2037 GNDA.n915 3.4105
R13775 GNDA.n935 GNDA.n915 3.4105
R13776 GNDA.n2039 GNDA.n915 3.4105
R13777 GNDA.n934 GNDA.n915 3.4105
R13778 GNDA.n2041 GNDA.n915 3.4105
R13779 GNDA.n933 GNDA.n915 3.4105
R13780 GNDA.n2043 GNDA.n915 3.4105
R13781 GNDA.n932 GNDA.n915 3.4105
R13782 GNDA.n2045 GNDA.n915 3.4105
R13783 GNDA.n931 GNDA.n915 3.4105
R13784 GNDA.n2047 GNDA.n915 3.4105
R13785 GNDA.n2049 GNDA.n915 3.4105
R13786 GNDA.n888 GNDA.n880 3.4105
R13787 GNDA.n2017 GNDA.n888 3.4105
R13788 GNDA.n945 GNDA.n888 3.4105
R13789 GNDA.n2019 GNDA.n888 3.4105
R13790 GNDA.n944 GNDA.n888 3.4105
R13791 GNDA.n2021 GNDA.n888 3.4105
R13792 GNDA.n943 GNDA.n888 3.4105
R13793 GNDA.n2023 GNDA.n888 3.4105
R13794 GNDA.n942 GNDA.n888 3.4105
R13795 GNDA.n2025 GNDA.n888 3.4105
R13796 GNDA.n941 GNDA.n888 3.4105
R13797 GNDA.n2027 GNDA.n888 3.4105
R13798 GNDA.n940 GNDA.n888 3.4105
R13799 GNDA.n2029 GNDA.n888 3.4105
R13800 GNDA.n939 GNDA.n888 3.4105
R13801 GNDA.n2031 GNDA.n888 3.4105
R13802 GNDA.n938 GNDA.n888 3.4105
R13803 GNDA.n2033 GNDA.n888 3.4105
R13804 GNDA.n937 GNDA.n888 3.4105
R13805 GNDA.n2035 GNDA.n888 3.4105
R13806 GNDA.n936 GNDA.n888 3.4105
R13807 GNDA.n2037 GNDA.n888 3.4105
R13808 GNDA.n935 GNDA.n888 3.4105
R13809 GNDA.n2039 GNDA.n888 3.4105
R13810 GNDA.n934 GNDA.n888 3.4105
R13811 GNDA.n2041 GNDA.n888 3.4105
R13812 GNDA.n933 GNDA.n888 3.4105
R13813 GNDA.n2043 GNDA.n888 3.4105
R13814 GNDA.n932 GNDA.n888 3.4105
R13815 GNDA.n2045 GNDA.n888 3.4105
R13816 GNDA.n931 GNDA.n888 3.4105
R13817 GNDA.n2047 GNDA.n888 3.4105
R13818 GNDA.n2049 GNDA.n888 3.4105
R13819 GNDA.n917 GNDA.n880 3.4105
R13820 GNDA.n2017 GNDA.n917 3.4105
R13821 GNDA.n945 GNDA.n917 3.4105
R13822 GNDA.n2019 GNDA.n917 3.4105
R13823 GNDA.n944 GNDA.n917 3.4105
R13824 GNDA.n2021 GNDA.n917 3.4105
R13825 GNDA.n943 GNDA.n917 3.4105
R13826 GNDA.n2023 GNDA.n917 3.4105
R13827 GNDA.n942 GNDA.n917 3.4105
R13828 GNDA.n2025 GNDA.n917 3.4105
R13829 GNDA.n941 GNDA.n917 3.4105
R13830 GNDA.n2027 GNDA.n917 3.4105
R13831 GNDA.n940 GNDA.n917 3.4105
R13832 GNDA.n2029 GNDA.n917 3.4105
R13833 GNDA.n939 GNDA.n917 3.4105
R13834 GNDA.n2031 GNDA.n917 3.4105
R13835 GNDA.n938 GNDA.n917 3.4105
R13836 GNDA.n2033 GNDA.n917 3.4105
R13837 GNDA.n937 GNDA.n917 3.4105
R13838 GNDA.n2035 GNDA.n917 3.4105
R13839 GNDA.n936 GNDA.n917 3.4105
R13840 GNDA.n2037 GNDA.n917 3.4105
R13841 GNDA.n935 GNDA.n917 3.4105
R13842 GNDA.n2039 GNDA.n917 3.4105
R13843 GNDA.n934 GNDA.n917 3.4105
R13844 GNDA.n2041 GNDA.n917 3.4105
R13845 GNDA.n933 GNDA.n917 3.4105
R13846 GNDA.n2043 GNDA.n917 3.4105
R13847 GNDA.n932 GNDA.n917 3.4105
R13848 GNDA.n2045 GNDA.n917 3.4105
R13849 GNDA.n931 GNDA.n917 3.4105
R13850 GNDA.n2047 GNDA.n917 3.4105
R13851 GNDA.n2049 GNDA.n917 3.4105
R13852 GNDA.n887 GNDA.n880 3.4105
R13853 GNDA.n2017 GNDA.n887 3.4105
R13854 GNDA.n945 GNDA.n887 3.4105
R13855 GNDA.n2019 GNDA.n887 3.4105
R13856 GNDA.n944 GNDA.n887 3.4105
R13857 GNDA.n2021 GNDA.n887 3.4105
R13858 GNDA.n943 GNDA.n887 3.4105
R13859 GNDA.n2023 GNDA.n887 3.4105
R13860 GNDA.n942 GNDA.n887 3.4105
R13861 GNDA.n2025 GNDA.n887 3.4105
R13862 GNDA.n941 GNDA.n887 3.4105
R13863 GNDA.n2027 GNDA.n887 3.4105
R13864 GNDA.n940 GNDA.n887 3.4105
R13865 GNDA.n2029 GNDA.n887 3.4105
R13866 GNDA.n939 GNDA.n887 3.4105
R13867 GNDA.n2031 GNDA.n887 3.4105
R13868 GNDA.n938 GNDA.n887 3.4105
R13869 GNDA.n2033 GNDA.n887 3.4105
R13870 GNDA.n937 GNDA.n887 3.4105
R13871 GNDA.n2035 GNDA.n887 3.4105
R13872 GNDA.n936 GNDA.n887 3.4105
R13873 GNDA.n2037 GNDA.n887 3.4105
R13874 GNDA.n935 GNDA.n887 3.4105
R13875 GNDA.n2039 GNDA.n887 3.4105
R13876 GNDA.n934 GNDA.n887 3.4105
R13877 GNDA.n2041 GNDA.n887 3.4105
R13878 GNDA.n933 GNDA.n887 3.4105
R13879 GNDA.n2043 GNDA.n887 3.4105
R13880 GNDA.n932 GNDA.n887 3.4105
R13881 GNDA.n2045 GNDA.n887 3.4105
R13882 GNDA.n931 GNDA.n887 3.4105
R13883 GNDA.n2047 GNDA.n887 3.4105
R13884 GNDA.n2049 GNDA.n887 3.4105
R13885 GNDA.n919 GNDA.n880 3.4105
R13886 GNDA.n2017 GNDA.n919 3.4105
R13887 GNDA.n945 GNDA.n919 3.4105
R13888 GNDA.n2019 GNDA.n919 3.4105
R13889 GNDA.n944 GNDA.n919 3.4105
R13890 GNDA.n2021 GNDA.n919 3.4105
R13891 GNDA.n943 GNDA.n919 3.4105
R13892 GNDA.n2023 GNDA.n919 3.4105
R13893 GNDA.n942 GNDA.n919 3.4105
R13894 GNDA.n2025 GNDA.n919 3.4105
R13895 GNDA.n941 GNDA.n919 3.4105
R13896 GNDA.n2027 GNDA.n919 3.4105
R13897 GNDA.n940 GNDA.n919 3.4105
R13898 GNDA.n2029 GNDA.n919 3.4105
R13899 GNDA.n939 GNDA.n919 3.4105
R13900 GNDA.n2031 GNDA.n919 3.4105
R13901 GNDA.n938 GNDA.n919 3.4105
R13902 GNDA.n2033 GNDA.n919 3.4105
R13903 GNDA.n937 GNDA.n919 3.4105
R13904 GNDA.n2035 GNDA.n919 3.4105
R13905 GNDA.n936 GNDA.n919 3.4105
R13906 GNDA.n2037 GNDA.n919 3.4105
R13907 GNDA.n935 GNDA.n919 3.4105
R13908 GNDA.n2039 GNDA.n919 3.4105
R13909 GNDA.n934 GNDA.n919 3.4105
R13910 GNDA.n2041 GNDA.n919 3.4105
R13911 GNDA.n933 GNDA.n919 3.4105
R13912 GNDA.n2043 GNDA.n919 3.4105
R13913 GNDA.n932 GNDA.n919 3.4105
R13914 GNDA.n2045 GNDA.n919 3.4105
R13915 GNDA.n931 GNDA.n919 3.4105
R13916 GNDA.n2047 GNDA.n919 3.4105
R13917 GNDA.n2049 GNDA.n919 3.4105
R13918 GNDA.n886 GNDA.n880 3.4105
R13919 GNDA.n2017 GNDA.n886 3.4105
R13920 GNDA.n945 GNDA.n886 3.4105
R13921 GNDA.n2019 GNDA.n886 3.4105
R13922 GNDA.n944 GNDA.n886 3.4105
R13923 GNDA.n2021 GNDA.n886 3.4105
R13924 GNDA.n943 GNDA.n886 3.4105
R13925 GNDA.n2023 GNDA.n886 3.4105
R13926 GNDA.n942 GNDA.n886 3.4105
R13927 GNDA.n2025 GNDA.n886 3.4105
R13928 GNDA.n941 GNDA.n886 3.4105
R13929 GNDA.n2027 GNDA.n886 3.4105
R13930 GNDA.n940 GNDA.n886 3.4105
R13931 GNDA.n2029 GNDA.n886 3.4105
R13932 GNDA.n939 GNDA.n886 3.4105
R13933 GNDA.n2031 GNDA.n886 3.4105
R13934 GNDA.n938 GNDA.n886 3.4105
R13935 GNDA.n2033 GNDA.n886 3.4105
R13936 GNDA.n937 GNDA.n886 3.4105
R13937 GNDA.n2035 GNDA.n886 3.4105
R13938 GNDA.n936 GNDA.n886 3.4105
R13939 GNDA.n2037 GNDA.n886 3.4105
R13940 GNDA.n935 GNDA.n886 3.4105
R13941 GNDA.n2039 GNDA.n886 3.4105
R13942 GNDA.n934 GNDA.n886 3.4105
R13943 GNDA.n2041 GNDA.n886 3.4105
R13944 GNDA.n933 GNDA.n886 3.4105
R13945 GNDA.n2043 GNDA.n886 3.4105
R13946 GNDA.n932 GNDA.n886 3.4105
R13947 GNDA.n2045 GNDA.n886 3.4105
R13948 GNDA.n931 GNDA.n886 3.4105
R13949 GNDA.n2047 GNDA.n886 3.4105
R13950 GNDA.n2049 GNDA.n886 3.4105
R13951 GNDA.n921 GNDA.n880 3.4105
R13952 GNDA.n2017 GNDA.n921 3.4105
R13953 GNDA.n945 GNDA.n921 3.4105
R13954 GNDA.n2019 GNDA.n921 3.4105
R13955 GNDA.n944 GNDA.n921 3.4105
R13956 GNDA.n2021 GNDA.n921 3.4105
R13957 GNDA.n943 GNDA.n921 3.4105
R13958 GNDA.n2023 GNDA.n921 3.4105
R13959 GNDA.n942 GNDA.n921 3.4105
R13960 GNDA.n2025 GNDA.n921 3.4105
R13961 GNDA.n941 GNDA.n921 3.4105
R13962 GNDA.n2027 GNDA.n921 3.4105
R13963 GNDA.n940 GNDA.n921 3.4105
R13964 GNDA.n2029 GNDA.n921 3.4105
R13965 GNDA.n939 GNDA.n921 3.4105
R13966 GNDA.n2031 GNDA.n921 3.4105
R13967 GNDA.n938 GNDA.n921 3.4105
R13968 GNDA.n2033 GNDA.n921 3.4105
R13969 GNDA.n937 GNDA.n921 3.4105
R13970 GNDA.n2035 GNDA.n921 3.4105
R13971 GNDA.n936 GNDA.n921 3.4105
R13972 GNDA.n2037 GNDA.n921 3.4105
R13973 GNDA.n935 GNDA.n921 3.4105
R13974 GNDA.n2039 GNDA.n921 3.4105
R13975 GNDA.n934 GNDA.n921 3.4105
R13976 GNDA.n2041 GNDA.n921 3.4105
R13977 GNDA.n933 GNDA.n921 3.4105
R13978 GNDA.n2043 GNDA.n921 3.4105
R13979 GNDA.n932 GNDA.n921 3.4105
R13980 GNDA.n2045 GNDA.n921 3.4105
R13981 GNDA.n931 GNDA.n921 3.4105
R13982 GNDA.n2047 GNDA.n921 3.4105
R13983 GNDA.n2049 GNDA.n921 3.4105
R13984 GNDA.n885 GNDA.n880 3.4105
R13985 GNDA.n2017 GNDA.n885 3.4105
R13986 GNDA.n945 GNDA.n885 3.4105
R13987 GNDA.n2019 GNDA.n885 3.4105
R13988 GNDA.n944 GNDA.n885 3.4105
R13989 GNDA.n2021 GNDA.n885 3.4105
R13990 GNDA.n943 GNDA.n885 3.4105
R13991 GNDA.n2023 GNDA.n885 3.4105
R13992 GNDA.n942 GNDA.n885 3.4105
R13993 GNDA.n2025 GNDA.n885 3.4105
R13994 GNDA.n941 GNDA.n885 3.4105
R13995 GNDA.n2027 GNDA.n885 3.4105
R13996 GNDA.n940 GNDA.n885 3.4105
R13997 GNDA.n2029 GNDA.n885 3.4105
R13998 GNDA.n939 GNDA.n885 3.4105
R13999 GNDA.n2031 GNDA.n885 3.4105
R14000 GNDA.n938 GNDA.n885 3.4105
R14001 GNDA.n2033 GNDA.n885 3.4105
R14002 GNDA.n937 GNDA.n885 3.4105
R14003 GNDA.n2035 GNDA.n885 3.4105
R14004 GNDA.n936 GNDA.n885 3.4105
R14005 GNDA.n2037 GNDA.n885 3.4105
R14006 GNDA.n935 GNDA.n885 3.4105
R14007 GNDA.n2039 GNDA.n885 3.4105
R14008 GNDA.n934 GNDA.n885 3.4105
R14009 GNDA.n2041 GNDA.n885 3.4105
R14010 GNDA.n933 GNDA.n885 3.4105
R14011 GNDA.n2043 GNDA.n885 3.4105
R14012 GNDA.n932 GNDA.n885 3.4105
R14013 GNDA.n2045 GNDA.n885 3.4105
R14014 GNDA.n931 GNDA.n885 3.4105
R14015 GNDA.n2047 GNDA.n885 3.4105
R14016 GNDA.n2049 GNDA.n885 3.4105
R14017 GNDA.n923 GNDA.n880 3.4105
R14018 GNDA.n2017 GNDA.n923 3.4105
R14019 GNDA.n945 GNDA.n923 3.4105
R14020 GNDA.n2019 GNDA.n923 3.4105
R14021 GNDA.n944 GNDA.n923 3.4105
R14022 GNDA.n2021 GNDA.n923 3.4105
R14023 GNDA.n943 GNDA.n923 3.4105
R14024 GNDA.n2023 GNDA.n923 3.4105
R14025 GNDA.n942 GNDA.n923 3.4105
R14026 GNDA.n2025 GNDA.n923 3.4105
R14027 GNDA.n941 GNDA.n923 3.4105
R14028 GNDA.n2027 GNDA.n923 3.4105
R14029 GNDA.n940 GNDA.n923 3.4105
R14030 GNDA.n2029 GNDA.n923 3.4105
R14031 GNDA.n939 GNDA.n923 3.4105
R14032 GNDA.n2031 GNDA.n923 3.4105
R14033 GNDA.n938 GNDA.n923 3.4105
R14034 GNDA.n2033 GNDA.n923 3.4105
R14035 GNDA.n937 GNDA.n923 3.4105
R14036 GNDA.n2035 GNDA.n923 3.4105
R14037 GNDA.n936 GNDA.n923 3.4105
R14038 GNDA.n2037 GNDA.n923 3.4105
R14039 GNDA.n935 GNDA.n923 3.4105
R14040 GNDA.n2039 GNDA.n923 3.4105
R14041 GNDA.n934 GNDA.n923 3.4105
R14042 GNDA.n2041 GNDA.n923 3.4105
R14043 GNDA.n933 GNDA.n923 3.4105
R14044 GNDA.n2043 GNDA.n923 3.4105
R14045 GNDA.n932 GNDA.n923 3.4105
R14046 GNDA.n2045 GNDA.n923 3.4105
R14047 GNDA.n931 GNDA.n923 3.4105
R14048 GNDA.n2047 GNDA.n923 3.4105
R14049 GNDA.n2049 GNDA.n923 3.4105
R14050 GNDA.n884 GNDA.n880 3.4105
R14051 GNDA.n2017 GNDA.n884 3.4105
R14052 GNDA.n945 GNDA.n884 3.4105
R14053 GNDA.n2019 GNDA.n884 3.4105
R14054 GNDA.n944 GNDA.n884 3.4105
R14055 GNDA.n2021 GNDA.n884 3.4105
R14056 GNDA.n943 GNDA.n884 3.4105
R14057 GNDA.n2023 GNDA.n884 3.4105
R14058 GNDA.n942 GNDA.n884 3.4105
R14059 GNDA.n2025 GNDA.n884 3.4105
R14060 GNDA.n941 GNDA.n884 3.4105
R14061 GNDA.n2027 GNDA.n884 3.4105
R14062 GNDA.n940 GNDA.n884 3.4105
R14063 GNDA.n2029 GNDA.n884 3.4105
R14064 GNDA.n939 GNDA.n884 3.4105
R14065 GNDA.n2031 GNDA.n884 3.4105
R14066 GNDA.n938 GNDA.n884 3.4105
R14067 GNDA.n2033 GNDA.n884 3.4105
R14068 GNDA.n937 GNDA.n884 3.4105
R14069 GNDA.n2035 GNDA.n884 3.4105
R14070 GNDA.n936 GNDA.n884 3.4105
R14071 GNDA.n2037 GNDA.n884 3.4105
R14072 GNDA.n935 GNDA.n884 3.4105
R14073 GNDA.n2039 GNDA.n884 3.4105
R14074 GNDA.n934 GNDA.n884 3.4105
R14075 GNDA.n2041 GNDA.n884 3.4105
R14076 GNDA.n933 GNDA.n884 3.4105
R14077 GNDA.n2043 GNDA.n884 3.4105
R14078 GNDA.n932 GNDA.n884 3.4105
R14079 GNDA.n2045 GNDA.n884 3.4105
R14080 GNDA.n931 GNDA.n884 3.4105
R14081 GNDA.n2047 GNDA.n884 3.4105
R14082 GNDA.n2049 GNDA.n884 3.4105
R14083 GNDA.n925 GNDA.n880 3.4105
R14084 GNDA.n2017 GNDA.n925 3.4105
R14085 GNDA.n945 GNDA.n925 3.4105
R14086 GNDA.n2019 GNDA.n925 3.4105
R14087 GNDA.n944 GNDA.n925 3.4105
R14088 GNDA.n2021 GNDA.n925 3.4105
R14089 GNDA.n943 GNDA.n925 3.4105
R14090 GNDA.n2023 GNDA.n925 3.4105
R14091 GNDA.n942 GNDA.n925 3.4105
R14092 GNDA.n2025 GNDA.n925 3.4105
R14093 GNDA.n941 GNDA.n925 3.4105
R14094 GNDA.n2027 GNDA.n925 3.4105
R14095 GNDA.n940 GNDA.n925 3.4105
R14096 GNDA.n2029 GNDA.n925 3.4105
R14097 GNDA.n939 GNDA.n925 3.4105
R14098 GNDA.n2031 GNDA.n925 3.4105
R14099 GNDA.n938 GNDA.n925 3.4105
R14100 GNDA.n2033 GNDA.n925 3.4105
R14101 GNDA.n937 GNDA.n925 3.4105
R14102 GNDA.n2035 GNDA.n925 3.4105
R14103 GNDA.n936 GNDA.n925 3.4105
R14104 GNDA.n2037 GNDA.n925 3.4105
R14105 GNDA.n935 GNDA.n925 3.4105
R14106 GNDA.n2039 GNDA.n925 3.4105
R14107 GNDA.n934 GNDA.n925 3.4105
R14108 GNDA.n2041 GNDA.n925 3.4105
R14109 GNDA.n933 GNDA.n925 3.4105
R14110 GNDA.n2043 GNDA.n925 3.4105
R14111 GNDA.n932 GNDA.n925 3.4105
R14112 GNDA.n2045 GNDA.n925 3.4105
R14113 GNDA.n931 GNDA.n925 3.4105
R14114 GNDA.n2047 GNDA.n925 3.4105
R14115 GNDA.n2049 GNDA.n925 3.4105
R14116 GNDA.n883 GNDA.n880 3.4105
R14117 GNDA.n2017 GNDA.n883 3.4105
R14118 GNDA.n945 GNDA.n883 3.4105
R14119 GNDA.n2019 GNDA.n883 3.4105
R14120 GNDA.n944 GNDA.n883 3.4105
R14121 GNDA.n2021 GNDA.n883 3.4105
R14122 GNDA.n943 GNDA.n883 3.4105
R14123 GNDA.n2023 GNDA.n883 3.4105
R14124 GNDA.n942 GNDA.n883 3.4105
R14125 GNDA.n2025 GNDA.n883 3.4105
R14126 GNDA.n941 GNDA.n883 3.4105
R14127 GNDA.n2027 GNDA.n883 3.4105
R14128 GNDA.n940 GNDA.n883 3.4105
R14129 GNDA.n2029 GNDA.n883 3.4105
R14130 GNDA.n939 GNDA.n883 3.4105
R14131 GNDA.n2031 GNDA.n883 3.4105
R14132 GNDA.n938 GNDA.n883 3.4105
R14133 GNDA.n2033 GNDA.n883 3.4105
R14134 GNDA.n937 GNDA.n883 3.4105
R14135 GNDA.n2035 GNDA.n883 3.4105
R14136 GNDA.n936 GNDA.n883 3.4105
R14137 GNDA.n2037 GNDA.n883 3.4105
R14138 GNDA.n935 GNDA.n883 3.4105
R14139 GNDA.n2039 GNDA.n883 3.4105
R14140 GNDA.n934 GNDA.n883 3.4105
R14141 GNDA.n2041 GNDA.n883 3.4105
R14142 GNDA.n933 GNDA.n883 3.4105
R14143 GNDA.n2043 GNDA.n883 3.4105
R14144 GNDA.n932 GNDA.n883 3.4105
R14145 GNDA.n2045 GNDA.n883 3.4105
R14146 GNDA.n931 GNDA.n883 3.4105
R14147 GNDA.n2047 GNDA.n883 3.4105
R14148 GNDA.n2049 GNDA.n883 3.4105
R14149 GNDA.n927 GNDA.n880 3.4105
R14150 GNDA.n2017 GNDA.n927 3.4105
R14151 GNDA.n945 GNDA.n927 3.4105
R14152 GNDA.n2019 GNDA.n927 3.4105
R14153 GNDA.n944 GNDA.n927 3.4105
R14154 GNDA.n2021 GNDA.n927 3.4105
R14155 GNDA.n943 GNDA.n927 3.4105
R14156 GNDA.n2023 GNDA.n927 3.4105
R14157 GNDA.n942 GNDA.n927 3.4105
R14158 GNDA.n2025 GNDA.n927 3.4105
R14159 GNDA.n941 GNDA.n927 3.4105
R14160 GNDA.n2027 GNDA.n927 3.4105
R14161 GNDA.n940 GNDA.n927 3.4105
R14162 GNDA.n2029 GNDA.n927 3.4105
R14163 GNDA.n939 GNDA.n927 3.4105
R14164 GNDA.n2031 GNDA.n927 3.4105
R14165 GNDA.n938 GNDA.n927 3.4105
R14166 GNDA.n2033 GNDA.n927 3.4105
R14167 GNDA.n937 GNDA.n927 3.4105
R14168 GNDA.n2035 GNDA.n927 3.4105
R14169 GNDA.n936 GNDA.n927 3.4105
R14170 GNDA.n2037 GNDA.n927 3.4105
R14171 GNDA.n935 GNDA.n927 3.4105
R14172 GNDA.n2039 GNDA.n927 3.4105
R14173 GNDA.n934 GNDA.n927 3.4105
R14174 GNDA.n2041 GNDA.n927 3.4105
R14175 GNDA.n933 GNDA.n927 3.4105
R14176 GNDA.n2043 GNDA.n927 3.4105
R14177 GNDA.n932 GNDA.n927 3.4105
R14178 GNDA.n2045 GNDA.n927 3.4105
R14179 GNDA.n931 GNDA.n927 3.4105
R14180 GNDA.n2047 GNDA.n927 3.4105
R14181 GNDA.n2049 GNDA.n927 3.4105
R14182 GNDA.n882 GNDA.n880 3.4105
R14183 GNDA.n2017 GNDA.n882 3.4105
R14184 GNDA.n945 GNDA.n882 3.4105
R14185 GNDA.n2019 GNDA.n882 3.4105
R14186 GNDA.n944 GNDA.n882 3.4105
R14187 GNDA.n2021 GNDA.n882 3.4105
R14188 GNDA.n943 GNDA.n882 3.4105
R14189 GNDA.n2023 GNDA.n882 3.4105
R14190 GNDA.n942 GNDA.n882 3.4105
R14191 GNDA.n2025 GNDA.n882 3.4105
R14192 GNDA.n941 GNDA.n882 3.4105
R14193 GNDA.n2027 GNDA.n882 3.4105
R14194 GNDA.n940 GNDA.n882 3.4105
R14195 GNDA.n2029 GNDA.n882 3.4105
R14196 GNDA.n939 GNDA.n882 3.4105
R14197 GNDA.n2031 GNDA.n882 3.4105
R14198 GNDA.n938 GNDA.n882 3.4105
R14199 GNDA.n2033 GNDA.n882 3.4105
R14200 GNDA.n937 GNDA.n882 3.4105
R14201 GNDA.n2035 GNDA.n882 3.4105
R14202 GNDA.n936 GNDA.n882 3.4105
R14203 GNDA.n2037 GNDA.n882 3.4105
R14204 GNDA.n935 GNDA.n882 3.4105
R14205 GNDA.n2039 GNDA.n882 3.4105
R14206 GNDA.n934 GNDA.n882 3.4105
R14207 GNDA.n2041 GNDA.n882 3.4105
R14208 GNDA.n933 GNDA.n882 3.4105
R14209 GNDA.n2043 GNDA.n882 3.4105
R14210 GNDA.n932 GNDA.n882 3.4105
R14211 GNDA.n2045 GNDA.n882 3.4105
R14212 GNDA.n931 GNDA.n882 3.4105
R14213 GNDA.n2047 GNDA.n882 3.4105
R14214 GNDA.n2049 GNDA.n882 3.4105
R14215 GNDA.n929 GNDA.n880 3.4105
R14216 GNDA.n2017 GNDA.n929 3.4105
R14217 GNDA.n945 GNDA.n929 3.4105
R14218 GNDA.n2019 GNDA.n929 3.4105
R14219 GNDA.n944 GNDA.n929 3.4105
R14220 GNDA.n2021 GNDA.n929 3.4105
R14221 GNDA.n943 GNDA.n929 3.4105
R14222 GNDA.n2023 GNDA.n929 3.4105
R14223 GNDA.n942 GNDA.n929 3.4105
R14224 GNDA.n2025 GNDA.n929 3.4105
R14225 GNDA.n941 GNDA.n929 3.4105
R14226 GNDA.n2027 GNDA.n929 3.4105
R14227 GNDA.n940 GNDA.n929 3.4105
R14228 GNDA.n2029 GNDA.n929 3.4105
R14229 GNDA.n939 GNDA.n929 3.4105
R14230 GNDA.n2031 GNDA.n929 3.4105
R14231 GNDA.n938 GNDA.n929 3.4105
R14232 GNDA.n2033 GNDA.n929 3.4105
R14233 GNDA.n937 GNDA.n929 3.4105
R14234 GNDA.n2035 GNDA.n929 3.4105
R14235 GNDA.n936 GNDA.n929 3.4105
R14236 GNDA.n2037 GNDA.n929 3.4105
R14237 GNDA.n935 GNDA.n929 3.4105
R14238 GNDA.n2039 GNDA.n929 3.4105
R14239 GNDA.n934 GNDA.n929 3.4105
R14240 GNDA.n2041 GNDA.n929 3.4105
R14241 GNDA.n933 GNDA.n929 3.4105
R14242 GNDA.n2043 GNDA.n929 3.4105
R14243 GNDA.n932 GNDA.n929 3.4105
R14244 GNDA.n2045 GNDA.n929 3.4105
R14245 GNDA.n931 GNDA.n929 3.4105
R14246 GNDA.n2047 GNDA.n929 3.4105
R14247 GNDA.n2049 GNDA.n929 3.4105
R14248 GNDA.n881 GNDA.n880 3.4105
R14249 GNDA.n2017 GNDA.n881 3.4105
R14250 GNDA.n945 GNDA.n881 3.4105
R14251 GNDA.n2019 GNDA.n881 3.4105
R14252 GNDA.n944 GNDA.n881 3.4105
R14253 GNDA.n2021 GNDA.n881 3.4105
R14254 GNDA.n943 GNDA.n881 3.4105
R14255 GNDA.n2023 GNDA.n881 3.4105
R14256 GNDA.n942 GNDA.n881 3.4105
R14257 GNDA.n2025 GNDA.n881 3.4105
R14258 GNDA.n941 GNDA.n881 3.4105
R14259 GNDA.n2027 GNDA.n881 3.4105
R14260 GNDA.n940 GNDA.n881 3.4105
R14261 GNDA.n2029 GNDA.n881 3.4105
R14262 GNDA.n939 GNDA.n881 3.4105
R14263 GNDA.n2031 GNDA.n881 3.4105
R14264 GNDA.n938 GNDA.n881 3.4105
R14265 GNDA.n2033 GNDA.n881 3.4105
R14266 GNDA.n937 GNDA.n881 3.4105
R14267 GNDA.n2035 GNDA.n881 3.4105
R14268 GNDA.n936 GNDA.n881 3.4105
R14269 GNDA.n2037 GNDA.n881 3.4105
R14270 GNDA.n935 GNDA.n881 3.4105
R14271 GNDA.n2039 GNDA.n881 3.4105
R14272 GNDA.n934 GNDA.n881 3.4105
R14273 GNDA.n2041 GNDA.n881 3.4105
R14274 GNDA.n933 GNDA.n881 3.4105
R14275 GNDA.n2043 GNDA.n881 3.4105
R14276 GNDA.n932 GNDA.n881 3.4105
R14277 GNDA.n2045 GNDA.n881 3.4105
R14278 GNDA.n931 GNDA.n881 3.4105
R14279 GNDA.n2047 GNDA.n881 3.4105
R14280 GNDA.n2049 GNDA.n881 3.4105
R14281 GNDA.n2048 GNDA.n2017 3.4105
R14282 GNDA.n2048 GNDA.n945 3.4105
R14283 GNDA.n2048 GNDA.n2019 3.4105
R14284 GNDA.n2048 GNDA.n944 3.4105
R14285 GNDA.n2048 GNDA.n2021 3.4105
R14286 GNDA.n2048 GNDA.n943 3.4105
R14287 GNDA.n2048 GNDA.n2023 3.4105
R14288 GNDA.n2048 GNDA.n942 3.4105
R14289 GNDA.n2048 GNDA.n2025 3.4105
R14290 GNDA.n2048 GNDA.n941 3.4105
R14291 GNDA.n2048 GNDA.n2027 3.4105
R14292 GNDA.n2048 GNDA.n940 3.4105
R14293 GNDA.n2048 GNDA.n2029 3.4105
R14294 GNDA.n2048 GNDA.n939 3.4105
R14295 GNDA.n2048 GNDA.n2031 3.4105
R14296 GNDA.n2048 GNDA.n938 3.4105
R14297 GNDA.n2048 GNDA.n2033 3.4105
R14298 GNDA.n2048 GNDA.n937 3.4105
R14299 GNDA.n2048 GNDA.n2035 3.4105
R14300 GNDA.n2048 GNDA.n936 3.4105
R14301 GNDA.n2048 GNDA.n2037 3.4105
R14302 GNDA.n2048 GNDA.n935 3.4105
R14303 GNDA.n2048 GNDA.n2039 3.4105
R14304 GNDA.n2048 GNDA.n934 3.4105
R14305 GNDA.n2048 GNDA.n2041 3.4105
R14306 GNDA.n2048 GNDA.n933 3.4105
R14307 GNDA.n2048 GNDA.n2043 3.4105
R14308 GNDA.n2048 GNDA.n932 3.4105
R14309 GNDA.n2048 GNDA.n2045 3.4105
R14310 GNDA.n2048 GNDA.n931 3.4105
R14311 GNDA.n2048 GNDA.n2047 3.4105
R14312 GNDA.n2049 GNDA.n2048 3.4105
R14313 GNDA.n1960 GNDA.n1045 3.4105
R14314 GNDA.n1960 GNDA.n1959 3.4105
R14315 GNDA.n1926 GNDA.n1062 3.4105
R14316 GNDA.n1062 GNDA.n1045 3.4105
R14317 GNDA.n1959 GNDA.n1062 3.4105
R14318 GNDA.n1926 GNDA.n1065 3.4105
R14319 GNDA.n1128 GNDA.n1065 3.4105
R14320 GNDA.n1928 GNDA.n1065 3.4105
R14321 GNDA.n1127 GNDA.n1065 3.4105
R14322 GNDA.n1930 GNDA.n1065 3.4105
R14323 GNDA.n1126 GNDA.n1065 3.4105
R14324 GNDA.n1932 GNDA.n1065 3.4105
R14325 GNDA.n1125 GNDA.n1065 3.4105
R14326 GNDA.n1934 GNDA.n1065 3.4105
R14327 GNDA.n1124 GNDA.n1065 3.4105
R14328 GNDA.n1936 GNDA.n1065 3.4105
R14329 GNDA.n1123 GNDA.n1065 3.4105
R14330 GNDA.n1938 GNDA.n1065 3.4105
R14331 GNDA.n1122 GNDA.n1065 3.4105
R14332 GNDA.n1940 GNDA.n1065 3.4105
R14333 GNDA.n1121 GNDA.n1065 3.4105
R14334 GNDA.n1942 GNDA.n1065 3.4105
R14335 GNDA.n1120 GNDA.n1065 3.4105
R14336 GNDA.n1944 GNDA.n1065 3.4105
R14337 GNDA.n1119 GNDA.n1065 3.4105
R14338 GNDA.n1946 GNDA.n1065 3.4105
R14339 GNDA.n1118 GNDA.n1065 3.4105
R14340 GNDA.n1948 GNDA.n1065 3.4105
R14341 GNDA.n1117 GNDA.n1065 3.4105
R14342 GNDA.n1950 GNDA.n1065 3.4105
R14343 GNDA.n1116 GNDA.n1065 3.4105
R14344 GNDA.n1952 GNDA.n1065 3.4105
R14345 GNDA.n1115 GNDA.n1065 3.4105
R14346 GNDA.n1954 GNDA.n1065 3.4105
R14347 GNDA.n1114 GNDA.n1065 3.4105
R14348 GNDA.n1956 GNDA.n1065 3.4105
R14349 GNDA.n1065 GNDA.n1045 3.4105
R14350 GNDA.n1959 GNDA.n1065 3.4105
R14351 GNDA.n1926 GNDA.n1061 3.4105
R14352 GNDA.n1128 GNDA.n1061 3.4105
R14353 GNDA.n1928 GNDA.n1061 3.4105
R14354 GNDA.n1127 GNDA.n1061 3.4105
R14355 GNDA.n1930 GNDA.n1061 3.4105
R14356 GNDA.n1126 GNDA.n1061 3.4105
R14357 GNDA.n1932 GNDA.n1061 3.4105
R14358 GNDA.n1125 GNDA.n1061 3.4105
R14359 GNDA.n1934 GNDA.n1061 3.4105
R14360 GNDA.n1124 GNDA.n1061 3.4105
R14361 GNDA.n1936 GNDA.n1061 3.4105
R14362 GNDA.n1123 GNDA.n1061 3.4105
R14363 GNDA.n1938 GNDA.n1061 3.4105
R14364 GNDA.n1122 GNDA.n1061 3.4105
R14365 GNDA.n1940 GNDA.n1061 3.4105
R14366 GNDA.n1121 GNDA.n1061 3.4105
R14367 GNDA.n1942 GNDA.n1061 3.4105
R14368 GNDA.n1120 GNDA.n1061 3.4105
R14369 GNDA.n1944 GNDA.n1061 3.4105
R14370 GNDA.n1119 GNDA.n1061 3.4105
R14371 GNDA.n1946 GNDA.n1061 3.4105
R14372 GNDA.n1118 GNDA.n1061 3.4105
R14373 GNDA.n1948 GNDA.n1061 3.4105
R14374 GNDA.n1117 GNDA.n1061 3.4105
R14375 GNDA.n1950 GNDA.n1061 3.4105
R14376 GNDA.n1116 GNDA.n1061 3.4105
R14377 GNDA.n1952 GNDA.n1061 3.4105
R14378 GNDA.n1115 GNDA.n1061 3.4105
R14379 GNDA.n1954 GNDA.n1061 3.4105
R14380 GNDA.n1114 GNDA.n1061 3.4105
R14381 GNDA.n1956 GNDA.n1061 3.4105
R14382 GNDA.n1061 GNDA.n1045 3.4105
R14383 GNDA.n1959 GNDA.n1061 3.4105
R14384 GNDA.n1926 GNDA.n1067 3.4105
R14385 GNDA.n1128 GNDA.n1067 3.4105
R14386 GNDA.n1928 GNDA.n1067 3.4105
R14387 GNDA.n1127 GNDA.n1067 3.4105
R14388 GNDA.n1930 GNDA.n1067 3.4105
R14389 GNDA.n1126 GNDA.n1067 3.4105
R14390 GNDA.n1932 GNDA.n1067 3.4105
R14391 GNDA.n1125 GNDA.n1067 3.4105
R14392 GNDA.n1934 GNDA.n1067 3.4105
R14393 GNDA.n1124 GNDA.n1067 3.4105
R14394 GNDA.n1936 GNDA.n1067 3.4105
R14395 GNDA.n1123 GNDA.n1067 3.4105
R14396 GNDA.n1938 GNDA.n1067 3.4105
R14397 GNDA.n1122 GNDA.n1067 3.4105
R14398 GNDA.n1940 GNDA.n1067 3.4105
R14399 GNDA.n1121 GNDA.n1067 3.4105
R14400 GNDA.n1942 GNDA.n1067 3.4105
R14401 GNDA.n1120 GNDA.n1067 3.4105
R14402 GNDA.n1944 GNDA.n1067 3.4105
R14403 GNDA.n1119 GNDA.n1067 3.4105
R14404 GNDA.n1946 GNDA.n1067 3.4105
R14405 GNDA.n1118 GNDA.n1067 3.4105
R14406 GNDA.n1948 GNDA.n1067 3.4105
R14407 GNDA.n1117 GNDA.n1067 3.4105
R14408 GNDA.n1950 GNDA.n1067 3.4105
R14409 GNDA.n1116 GNDA.n1067 3.4105
R14410 GNDA.n1952 GNDA.n1067 3.4105
R14411 GNDA.n1115 GNDA.n1067 3.4105
R14412 GNDA.n1954 GNDA.n1067 3.4105
R14413 GNDA.n1114 GNDA.n1067 3.4105
R14414 GNDA.n1956 GNDA.n1067 3.4105
R14415 GNDA.n1067 GNDA.n1045 3.4105
R14416 GNDA.n1959 GNDA.n1067 3.4105
R14417 GNDA.n1926 GNDA.n1060 3.4105
R14418 GNDA.n1128 GNDA.n1060 3.4105
R14419 GNDA.n1928 GNDA.n1060 3.4105
R14420 GNDA.n1127 GNDA.n1060 3.4105
R14421 GNDA.n1930 GNDA.n1060 3.4105
R14422 GNDA.n1126 GNDA.n1060 3.4105
R14423 GNDA.n1932 GNDA.n1060 3.4105
R14424 GNDA.n1125 GNDA.n1060 3.4105
R14425 GNDA.n1934 GNDA.n1060 3.4105
R14426 GNDA.n1124 GNDA.n1060 3.4105
R14427 GNDA.n1936 GNDA.n1060 3.4105
R14428 GNDA.n1123 GNDA.n1060 3.4105
R14429 GNDA.n1938 GNDA.n1060 3.4105
R14430 GNDA.n1122 GNDA.n1060 3.4105
R14431 GNDA.n1940 GNDA.n1060 3.4105
R14432 GNDA.n1121 GNDA.n1060 3.4105
R14433 GNDA.n1942 GNDA.n1060 3.4105
R14434 GNDA.n1120 GNDA.n1060 3.4105
R14435 GNDA.n1944 GNDA.n1060 3.4105
R14436 GNDA.n1119 GNDA.n1060 3.4105
R14437 GNDA.n1946 GNDA.n1060 3.4105
R14438 GNDA.n1118 GNDA.n1060 3.4105
R14439 GNDA.n1948 GNDA.n1060 3.4105
R14440 GNDA.n1117 GNDA.n1060 3.4105
R14441 GNDA.n1950 GNDA.n1060 3.4105
R14442 GNDA.n1116 GNDA.n1060 3.4105
R14443 GNDA.n1952 GNDA.n1060 3.4105
R14444 GNDA.n1115 GNDA.n1060 3.4105
R14445 GNDA.n1954 GNDA.n1060 3.4105
R14446 GNDA.n1114 GNDA.n1060 3.4105
R14447 GNDA.n1956 GNDA.n1060 3.4105
R14448 GNDA.n1060 GNDA.n1045 3.4105
R14449 GNDA.n1959 GNDA.n1060 3.4105
R14450 GNDA.n1926 GNDA.n1069 3.4105
R14451 GNDA.n1128 GNDA.n1069 3.4105
R14452 GNDA.n1928 GNDA.n1069 3.4105
R14453 GNDA.n1127 GNDA.n1069 3.4105
R14454 GNDA.n1930 GNDA.n1069 3.4105
R14455 GNDA.n1126 GNDA.n1069 3.4105
R14456 GNDA.n1932 GNDA.n1069 3.4105
R14457 GNDA.n1125 GNDA.n1069 3.4105
R14458 GNDA.n1934 GNDA.n1069 3.4105
R14459 GNDA.n1124 GNDA.n1069 3.4105
R14460 GNDA.n1936 GNDA.n1069 3.4105
R14461 GNDA.n1123 GNDA.n1069 3.4105
R14462 GNDA.n1938 GNDA.n1069 3.4105
R14463 GNDA.n1122 GNDA.n1069 3.4105
R14464 GNDA.n1940 GNDA.n1069 3.4105
R14465 GNDA.n1121 GNDA.n1069 3.4105
R14466 GNDA.n1942 GNDA.n1069 3.4105
R14467 GNDA.n1120 GNDA.n1069 3.4105
R14468 GNDA.n1944 GNDA.n1069 3.4105
R14469 GNDA.n1119 GNDA.n1069 3.4105
R14470 GNDA.n1946 GNDA.n1069 3.4105
R14471 GNDA.n1118 GNDA.n1069 3.4105
R14472 GNDA.n1948 GNDA.n1069 3.4105
R14473 GNDA.n1117 GNDA.n1069 3.4105
R14474 GNDA.n1950 GNDA.n1069 3.4105
R14475 GNDA.n1116 GNDA.n1069 3.4105
R14476 GNDA.n1952 GNDA.n1069 3.4105
R14477 GNDA.n1115 GNDA.n1069 3.4105
R14478 GNDA.n1954 GNDA.n1069 3.4105
R14479 GNDA.n1114 GNDA.n1069 3.4105
R14480 GNDA.n1956 GNDA.n1069 3.4105
R14481 GNDA.n1069 GNDA.n1045 3.4105
R14482 GNDA.n1959 GNDA.n1069 3.4105
R14483 GNDA.n1926 GNDA.n1059 3.4105
R14484 GNDA.n1128 GNDA.n1059 3.4105
R14485 GNDA.n1928 GNDA.n1059 3.4105
R14486 GNDA.n1127 GNDA.n1059 3.4105
R14487 GNDA.n1930 GNDA.n1059 3.4105
R14488 GNDA.n1126 GNDA.n1059 3.4105
R14489 GNDA.n1932 GNDA.n1059 3.4105
R14490 GNDA.n1125 GNDA.n1059 3.4105
R14491 GNDA.n1934 GNDA.n1059 3.4105
R14492 GNDA.n1124 GNDA.n1059 3.4105
R14493 GNDA.n1936 GNDA.n1059 3.4105
R14494 GNDA.n1123 GNDA.n1059 3.4105
R14495 GNDA.n1938 GNDA.n1059 3.4105
R14496 GNDA.n1122 GNDA.n1059 3.4105
R14497 GNDA.n1940 GNDA.n1059 3.4105
R14498 GNDA.n1121 GNDA.n1059 3.4105
R14499 GNDA.n1942 GNDA.n1059 3.4105
R14500 GNDA.n1120 GNDA.n1059 3.4105
R14501 GNDA.n1944 GNDA.n1059 3.4105
R14502 GNDA.n1119 GNDA.n1059 3.4105
R14503 GNDA.n1946 GNDA.n1059 3.4105
R14504 GNDA.n1118 GNDA.n1059 3.4105
R14505 GNDA.n1948 GNDA.n1059 3.4105
R14506 GNDA.n1117 GNDA.n1059 3.4105
R14507 GNDA.n1950 GNDA.n1059 3.4105
R14508 GNDA.n1116 GNDA.n1059 3.4105
R14509 GNDA.n1952 GNDA.n1059 3.4105
R14510 GNDA.n1115 GNDA.n1059 3.4105
R14511 GNDA.n1954 GNDA.n1059 3.4105
R14512 GNDA.n1114 GNDA.n1059 3.4105
R14513 GNDA.n1956 GNDA.n1059 3.4105
R14514 GNDA.n1059 GNDA.n1045 3.4105
R14515 GNDA.n1959 GNDA.n1059 3.4105
R14516 GNDA.n1926 GNDA.n1071 3.4105
R14517 GNDA.n1128 GNDA.n1071 3.4105
R14518 GNDA.n1928 GNDA.n1071 3.4105
R14519 GNDA.n1127 GNDA.n1071 3.4105
R14520 GNDA.n1930 GNDA.n1071 3.4105
R14521 GNDA.n1126 GNDA.n1071 3.4105
R14522 GNDA.n1932 GNDA.n1071 3.4105
R14523 GNDA.n1125 GNDA.n1071 3.4105
R14524 GNDA.n1934 GNDA.n1071 3.4105
R14525 GNDA.n1124 GNDA.n1071 3.4105
R14526 GNDA.n1936 GNDA.n1071 3.4105
R14527 GNDA.n1123 GNDA.n1071 3.4105
R14528 GNDA.n1938 GNDA.n1071 3.4105
R14529 GNDA.n1122 GNDA.n1071 3.4105
R14530 GNDA.n1940 GNDA.n1071 3.4105
R14531 GNDA.n1121 GNDA.n1071 3.4105
R14532 GNDA.n1942 GNDA.n1071 3.4105
R14533 GNDA.n1120 GNDA.n1071 3.4105
R14534 GNDA.n1944 GNDA.n1071 3.4105
R14535 GNDA.n1119 GNDA.n1071 3.4105
R14536 GNDA.n1946 GNDA.n1071 3.4105
R14537 GNDA.n1118 GNDA.n1071 3.4105
R14538 GNDA.n1948 GNDA.n1071 3.4105
R14539 GNDA.n1117 GNDA.n1071 3.4105
R14540 GNDA.n1950 GNDA.n1071 3.4105
R14541 GNDA.n1116 GNDA.n1071 3.4105
R14542 GNDA.n1952 GNDA.n1071 3.4105
R14543 GNDA.n1115 GNDA.n1071 3.4105
R14544 GNDA.n1954 GNDA.n1071 3.4105
R14545 GNDA.n1114 GNDA.n1071 3.4105
R14546 GNDA.n1956 GNDA.n1071 3.4105
R14547 GNDA.n1071 GNDA.n1045 3.4105
R14548 GNDA.n1959 GNDA.n1071 3.4105
R14549 GNDA.n1926 GNDA.n1058 3.4105
R14550 GNDA.n1128 GNDA.n1058 3.4105
R14551 GNDA.n1928 GNDA.n1058 3.4105
R14552 GNDA.n1127 GNDA.n1058 3.4105
R14553 GNDA.n1930 GNDA.n1058 3.4105
R14554 GNDA.n1126 GNDA.n1058 3.4105
R14555 GNDA.n1932 GNDA.n1058 3.4105
R14556 GNDA.n1125 GNDA.n1058 3.4105
R14557 GNDA.n1934 GNDA.n1058 3.4105
R14558 GNDA.n1124 GNDA.n1058 3.4105
R14559 GNDA.n1936 GNDA.n1058 3.4105
R14560 GNDA.n1123 GNDA.n1058 3.4105
R14561 GNDA.n1938 GNDA.n1058 3.4105
R14562 GNDA.n1122 GNDA.n1058 3.4105
R14563 GNDA.n1940 GNDA.n1058 3.4105
R14564 GNDA.n1121 GNDA.n1058 3.4105
R14565 GNDA.n1942 GNDA.n1058 3.4105
R14566 GNDA.n1120 GNDA.n1058 3.4105
R14567 GNDA.n1944 GNDA.n1058 3.4105
R14568 GNDA.n1119 GNDA.n1058 3.4105
R14569 GNDA.n1946 GNDA.n1058 3.4105
R14570 GNDA.n1118 GNDA.n1058 3.4105
R14571 GNDA.n1948 GNDA.n1058 3.4105
R14572 GNDA.n1117 GNDA.n1058 3.4105
R14573 GNDA.n1950 GNDA.n1058 3.4105
R14574 GNDA.n1116 GNDA.n1058 3.4105
R14575 GNDA.n1952 GNDA.n1058 3.4105
R14576 GNDA.n1115 GNDA.n1058 3.4105
R14577 GNDA.n1954 GNDA.n1058 3.4105
R14578 GNDA.n1114 GNDA.n1058 3.4105
R14579 GNDA.n1956 GNDA.n1058 3.4105
R14580 GNDA.n1058 GNDA.n1045 3.4105
R14581 GNDA.n1959 GNDA.n1058 3.4105
R14582 GNDA.n1926 GNDA.n1073 3.4105
R14583 GNDA.n1128 GNDA.n1073 3.4105
R14584 GNDA.n1928 GNDA.n1073 3.4105
R14585 GNDA.n1127 GNDA.n1073 3.4105
R14586 GNDA.n1930 GNDA.n1073 3.4105
R14587 GNDA.n1126 GNDA.n1073 3.4105
R14588 GNDA.n1932 GNDA.n1073 3.4105
R14589 GNDA.n1125 GNDA.n1073 3.4105
R14590 GNDA.n1934 GNDA.n1073 3.4105
R14591 GNDA.n1124 GNDA.n1073 3.4105
R14592 GNDA.n1936 GNDA.n1073 3.4105
R14593 GNDA.n1123 GNDA.n1073 3.4105
R14594 GNDA.n1938 GNDA.n1073 3.4105
R14595 GNDA.n1122 GNDA.n1073 3.4105
R14596 GNDA.n1940 GNDA.n1073 3.4105
R14597 GNDA.n1121 GNDA.n1073 3.4105
R14598 GNDA.n1942 GNDA.n1073 3.4105
R14599 GNDA.n1120 GNDA.n1073 3.4105
R14600 GNDA.n1944 GNDA.n1073 3.4105
R14601 GNDA.n1119 GNDA.n1073 3.4105
R14602 GNDA.n1946 GNDA.n1073 3.4105
R14603 GNDA.n1118 GNDA.n1073 3.4105
R14604 GNDA.n1948 GNDA.n1073 3.4105
R14605 GNDA.n1117 GNDA.n1073 3.4105
R14606 GNDA.n1950 GNDA.n1073 3.4105
R14607 GNDA.n1116 GNDA.n1073 3.4105
R14608 GNDA.n1952 GNDA.n1073 3.4105
R14609 GNDA.n1115 GNDA.n1073 3.4105
R14610 GNDA.n1954 GNDA.n1073 3.4105
R14611 GNDA.n1114 GNDA.n1073 3.4105
R14612 GNDA.n1956 GNDA.n1073 3.4105
R14613 GNDA.n1073 GNDA.n1045 3.4105
R14614 GNDA.n1959 GNDA.n1073 3.4105
R14615 GNDA.n1926 GNDA.n1057 3.4105
R14616 GNDA.n1128 GNDA.n1057 3.4105
R14617 GNDA.n1928 GNDA.n1057 3.4105
R14618 GNDA.n1127 GNDA.n1057 3.4105
R14619 GNDA.n1930 GNDA.n1057 3.4105
R14620 GNDA.n1126 GNDA.n1057 3.4105
R14621 GNDA.n1932 GNDA.n1057 3.4105
R14622 GNDA.n1125 GNDA.n1057 3.4105
R14623 GNDA.n1934 GNDA.n1057 3.4105
R14624 GNDA.n1124 GNDA.n1057 3.4105
R14625 GNDA.n1936 GNDA.n1057 3.4105
R14626 GNDA.n1123 GNDA.n1057 3.4105
R14627 GNDA.n1938 GNDA.n1057 3.4105
R14628 GNDA.n1122 GNDA.n1057 3.4105
R14629 GNDA.n1940 GNDA.n1057 3.4105
R14630 GNDA.n1121 GNDA.n1057 3.4105
R14631 GNDA.n1942 GNDA.n1057 3.4105
R14632 GNDA.n1120 GNDA.n1057 3.4105
R14633 GNDA.n1944 GNDA.n1057 3.4105
R14634 GNDA.n1119 GNDA.n1057 3.4105
R14635 GNDA.n1946 GNDA.n1057 3.4105
R14636 GNDA.n1118 GNDA.n1057 3.4105
R14637 GNDA.n1948 GNDA.n1057 3.4105
R14638 GNDA.n1117 GNDA.n1057 3.4105
R14639 GNDA.n1950 GNDA.n1057 3.4105
R14640 GNDA.n1116 GNDA.n1057 3.4105
R14641 GNDA.n1952 GNDA.n1057 3.4105
R14642 GNDA.n1115 GNDA.n1057 3.4105
R14643 GNDA.n1954 GNDA.n1057 3.4105
R14644 GNDA.n1114 GNDA.n1057 3.4105
R14645 GNDA.n1956 GNDA.n1057 3.4105
R14646 GNDA.n1057 GNDA.n1045 3.4105
R14647 GNDA.n1959 GNDA.n1057 3.4105
R14648 GNDA.n1926 GNDA.n1075 3.4105
R14649 GNDA.n1128 GNDA.n1075 3.4105
R14650 GNDA.n1928 GNDA.n1075 3.4105
R14651 GNDA.n1127 GNDA.n1075 3.4105
R14652 GNDA.n1930 GNDA.n1075 3.4105
R14653 GNDA.n1126 GNDA.n1075 3.4105
R14654 GNDA.n1932 GNDA.n1075 3.4105
R14655 GNDA.n1125 GNDA.n1075 3.4105
R14656 GNDA.n1934 GNDA.n1075 3.4105
R14657 GNDA.n1124 GNDA.n1075 3.4105
R14658 GNDA.n1936 GNDA.n1075 3.4105
R14659 GNDA.n1123 GNDA.n1075 3.4105
R14660 GNDA.n1938 GNDA.n1075 3.4105
R14661 GNDA.n1122 GNDA.n1075 3.4105
R14662 GNDA.n1940 GNDA.n1075 3.4105
R14663 GNDA.n1121 GNDA.n1075 3.4105
R14664 GNDA.n1942 GNDA.n1075 3.4105
R14665 GNDA.n1120 GNDA.n1075 3.4105
R14666 GNDA.n1944 GNDA.n1075 3.4105
R14667 GNDA.n1119 GNDA.n1075 3.4105
R14668 GNDA.n1946 GNDA.n1075 3.4105
R14669 GNDA.n1118 GNDA.n1075 3.4105
R14670 GNDA.n1948 GNDA.n1075 3.4105
R14671 GNDA.n1117 GNDA.n1075 3.4105
R14672 GNDA.n1950 GNDA.n1075 3.4105
R14673 GNDA.n1116 GNDA.n1075 3.4105
R14674 GNDA.n1952 GNDA.n1075 3.4105
R14675 GNDA.n1115 GNDA.n1075 3.4105
R14676 GNDA.n1954 GNDA.n1075 3.4105
R14677 GNDA.n1114 GNDA.n1075 3.4105
R14678 GNDA.n1956 GNDA.n1075 3.4105
R14679 GNDA.n1075 GNDA.n1045 3.4105
R14680 GNDA.n1959 GNDA.n1075 3.4105
R14681 GNDA.n1926 GNDA.n1056 3.4105
R14682 GNDA.n1128 GNDA.n1056 3.4105
R14683 GNDA.n1928 GNDA.n1056 3.4105
R14684 GNDA.n1127 GNDA.n1056 3.4105
R14685 GNDA.n1930 GNDA.n1056 3.4105
R14686 GNDA.n1126 GNDA.n1056 3.4105
R14687 GNDA.n1932 GNDA.n1056 3.4105
R14688 GNDA.n1125 GNDA.n1056 3.4105
R14689 GNDA.n1934 GNDA.n1056 3.4105
R14690 GNDA.n1124 GNDA.n1056 3.4105
R14691 GNDA.n1936 GNDA.n1056 3.4105
R14692 GNDA.n1123 GNDA.n1056 3.4105
R14693 GNDA.n1938 GNDA.n1056 3.4105
R14694 GNDA.n1122 GNDA.n1056 3.4105
R14695 GNDA.n1940 GNDA.n1056 3.4105
R14696 GNDA.n1121 GNDA.n1056 3.4105
R14697 GNDA.n1942 GNDA.n1056 3.4105
R14698 GNDA.n1120 GNDA.n1056 3.4105
R14699 GNDA.n1944 GNDA.n1056 3.4105
R14700 GNDA.n1119 GNDA.n1056 3.4105
R14701 GNDA.n1946 GNDA.n1056 3.4105
R14702 GNDA.n1118 GNDA.n1056 3.4105
R14703 GNDA.n1948 GNDA.n1056 3.4105
R14704 GNDA.n1117 GNDA.n1056 3.4105
R14705 GNDA.n1950 GNDA.n1056 3.4105
R14706 GNDA.n1116 GNDA.n1056 3.4105
R14707 GNDA.n1952 GNDA.n1056 3.4105
R14708 GNDA.n1115 GNDA.n1056 3.4105
R14709 GNDA.n1954 GNDA.n1056 3.4105
R14710 GNDA.n1114 GNDA.n1056 3.4105
R14711 GNDA.n1956 GNDA.n1056 3.4105
R14712 GNDA.n1056 GNDA.n1045 3.4105
R14713 GNDA.n1959 GNDA.n1056 3.4105
R14714 GNDA.n1926 GNDA.n1077 3.4105
R14715 GNDA.n1128 GNDA.n1077 3.4105
R14716 GNDA.n1928 GNDA.n1077 3.4105
R14717 GNDA.n1127 GNDA.n1077 3.4105
R14718 GNDA.n1930 GNDA.n1077 3.4105
R14719 GNDA.n1126 GNDA.n1077 3.4105
R14720 GNDA.n1932 GNDA.n1077 3.4105
R14721 GNDA.n1125 GNDA.n1077 3.4105
R14722 GNDA.n1934 GNDA.n1077 3.4105
R14723 GNDA.n1124 GNDA.n1077 3.4105
R14724 GNDA.n1936 GNDA.n1077 3.4105
R14725 GNDA.n1123 GNDA.n1077 3.4105
R14726 GNDA.n1938 GNDA.n1077 3.4105
R14727 GNDA.n1122 GNDA.n1077 3.4105
R14728 GNDA.n1940 GNDA.n1077 3.4105
R14729 GNDA.n1121 GNDA.n1077 3.4105
R14730 GNDA.n1942 GNDA.n1077 3.4105
R14731 GNDA.n1120 GNDA.n1077 3.4105
R14732 GNDA.n1944 GNDA.n1077 3.4105
R14733 GNDA.n1119 GNDA.n1077 3.4105
R14734 GNDA.n1946 GNDA.n1077 3.4105
R14735 GNDA.n1118 GNDA.n1077 3.4105
R14736 GNDA.n1948 GNDA.n1077 3.4105
R14737 GNDA.n1117 GNDA.n1077 3.4105
R14738 GNDA.n1950 GNDA.n1077 3.4105
R14739 GNDA.n1116 GNDA.n1077 3.4105
R14740 GNDA.n1952 GNDA.n1077 3.4105
R14741 GNDA.n1115 GNDA.n1077 3.4105
R14742 GNDA.n1954 GNDA.n1077 3.4105
R14743 GNDA.n1114 GNDA.n1077 3.4105
R14744 GNDA.n1956 GNDA.n1077 3.4105
R14745 GNDA.n1077 GNDA.n1045 3.4105
R14746 GNDA.n1959 GNDA.n1077 3.4105
R14747 GNDA.n1926 GNDA.n1055 3.4105
R14748 GNDA.n1128 GNDA.n1055 3.4105
R14749 GNDA.n1928 GNDA.n1055 3.4105
R14750 GNDA.n1127 GNDA.n1055 3.4105
R14751 GNDA.n1930 GNDA.n1055 3.4105
R14752 GNDA.n1126 GNDA.n1055 3.4105
R14753 GNDA.n1932 GNDA.n1055 3.4105
R14754 GNDA.n1125 GNDA.n1055 3.4105
R14755 GNDA.n1934 GNDA.n1055 3.4105
R14756 GNDA.n1124 GNDA.n1055 3.4105
R14757 GNDA.n1936 GNDA.n1055 3.4105
R14758 GNDA.n1123 GNDA.n1055 3.4105
R14759 GNDA.n1938 GNDA.n1055 3.4105
R14760 GNDA.n1122 GNDA.n1055 3.4105
R14761 GNDA.n1940 GNDA.n1055 3.4105
R14762 GNDA.n1121 GNDA.n1055 3.4105
R14763 GNDA.n1942 GNDA.n1055 3.4105
R14764 GNDA.n1120 GNDA.n1055 3.4105
R14765 GNDA.n1944 GNDA.n1055 3.4105
R14766 GNDA.n1119 GNDA.n1055 3.4105
R14767 GNDA.n1946 GNDA.n1055 3.4105
R14768 GNDA.n1118 GNDA.n1055 3.4105
R14769 GNDA.n1948 GNDA.n1055 3.4105
R14770 GNDA.n1117 GNDA.n1055 3.4105
R14771 GNDA.n1950 GNDA.n1055 3.4105
R14772 GNDA.n1116 GNDA.n1055 3.4105
R14773 GNDA.n1952 GNDA.n1055 3.4105
R14774 GNDA.n1115 GNDA.n1055 3.4105
R14775 GNDA.n1954 GNDA.n1055 3.4105
R14776 GNDA.n1114 GNDA.n1055 3.4105
R14777 GNDA.n1956 GNDA.n1055 3.4105
R14778 GNDA.n1055 GNDA.n1045 3.4105
R14779 GNDA.n1959 GNDA.n1055 3.4105
R14780 GNDA.n1926 GNDA.n1079 3.4105
R14781 GNDA.n1128 GNDA.n1079 3.4105
R14782 GNDA.n1928 GNDA.n1079 3.4105
R14783 GNDA.n1127 GNDA.n1079 3.4105
R14784 GNDA.n1930 GNDA.n1079 3.4105
R14785 GNDA.n1126 GNDA.n1079 3.4105
R14786 GNDA.n1932 GNDA.n1079 3.4105
R14787 GNDA.n1125 GNDA.n1079 3.4105
R14788 GNDA.n1934 GNDA.n1079 3.4105
R14789 GNDA.n1124 GNDA.n1079 3.4105
R14790 GNDA.n1936 GNDA.n1079 3.4105
R14791 GNDA.n1123 GNDA.n1079 3.4105
R14792 GNDA.n1938 GNDA.n1079 3.4105
R14793 GNDA.n1122 GNDA.n1079 3.4105
R14794 GNDA.n1940 GNDA.n1079 3.4105
R14795 GNDA.n1121 GNDA.n1079 3.4105
R14796 GNDA.n1942 GNDA.n1079 3.4105
R14797 GNDA.n1120 GNDA.n1079 3.4105
R14798 GNDA.n1944 GNDA.n1079 3.4105
R14799 GNDA.n1119 GNDA.n1079 3.4105
R14800 GNDA.n1946 GNDA.n1079 3.4105
R14801 GNDA.n1118 GNDA.n1079 3.4105
R14802 GNDA.n1948 GNDA.n1079 3.4105
R14803 GNDA.n1117 GNDA.n1079 3.4105
R14804 GNDA.n1950 GNDA.n1079 3.4105
R14805 GNDA.n1116 GNDA.n1079 3.4105
R14806 GNDA.n1952 GNDA.n1079 3.4105
R14807 GNDA.n1115 GNDA.n1079 3.4105
R14808 GNDA.n1954 GNDA.n1079 3.4105
R14809 GNDA.n1114 GNDA.n1079 3.4105
R14810 GNDA.n1956 GNDA.n1079 3.4105
R14811 GNDA.n1079 GNDA.n1045 3.4105
R14812 GNDA.n1959 GNDA.n1079 3.4105
R14813 GNDA.n1926 GNDA.n1054 3.4105
R14814 GNDA.n1128 GNDA.n1054 3.4105
R14815 GNDA.n1928 GNDA.n1054 3.4105
R14816 GNDA.n1127 GNDA.n1054 3.4105
R14817 GNDA.n1930 GNDA.n1054 3.4105
R14818 GNDA.n1126 GNDA.n1054 3.4105
R14819 GNDA.n1932 GNDA.n1054 3.4105
R14820 GNDA.n1125 GNDA.n1054 3.4105
R14821 GNDA.n1934 GNDA.n1054 3.4105
R14822 GNDA.n1124 GNDA.n1054 3.4105
R14823 GNDA.n1936 GNDA.n1054 3.4105
R14824 GNDA.n1123 GNDA.n1054 3.4105
R14825 GNDA.n1938 GNDA.n1054 3.4105
R14826 GNDA.n1122 GNDA.n1054 3.4105
R14827 GNDA.n1940 GNDA.n1054 3.4105
R14828 GNDA.n1121 GNDA.n1054 3.4105
R14829 GNDA.n1942 GNDA.n1054 3.4105
R14830 GNDA.n1120 GNDA.n1054 3.4105
R14831 GNDA.n1944 GNDA.n1054 3.4105
R14832 GNDA.n1119 GNDA.n1054 3.4105
R14833 GNDA.n1946 GNDA.n1054 3.4105
R14834 GNDA.n1118 GNDA.n1054 3.4105
R14835 GNDA.n1948 GNDA.n1054 3.4105
R14836 GNDA.n1117 GNDA.n1054 3.4105
R14837 GNDA.n1950 GNDA.n1054 3.4105
R14838 GNDA.n1116 GNDA.n1054 3.4105
R14839 GNDA.n1952 GNDA.n1054 3.4105
R14840 GNDA.n1115 GNDA.n1054 3.4105
R14841 GNDA.n1954 GNDA.n1054 3.4105
R14842 GNDA.n1114 GNDA.n1054 3.4105
R14843 GNDA.n1956 GNDA.n1054 3.4105
R14844 GNDA.n1054 GNDA.n1045 3.4105
R14845 GNDA.n1959 GNDA.n1054 3.4105
R14846 GNDA.n1926 GNDA.n1081 3.4105
R14847 GNDA.n1128 GNDA.n1081 3.4105
R14848 GNDA.n1928 GNDA.n1081 3.4105
R14849 GNDA.n1127 GNDA.n1081 3.4105
R14850 GNDA.n1930 GNDA.n1081 3.4105
R14851 GNDA.n1126 GNDA.n1081 3.4105
R14852 GNDA.n1932 GNDA.n1081 3.4105
R14853 GNDA.n1125 GNDA.n1081 3.4105
R14854 GNDA.n1934 GNDA.n1081 3.4105
R14855 GNDA.n1124 GNDA.n1081 3.4105
R14856 GNDA.n1936 GNDA.n1081 3.4105
R14857 GNDA.n1123 GNDA.n1081 3.4105
R14858 GNDA.n1938 GNDA.n1081 3.4105
R14859 GNDA.n1122 GNDA.n1081 3.4105
R14860 GNDA.n1940 GNDA.n1081 3.4105
R14861 GNDA.n1121 GNDA.n1081 3.4105
R14862 GNDA.n1942 GNDA.n1081 3.4105
R14863 GNDA.n1120 GNDA.n1081 3.4105
R14864 GNDA.n1944 GNDA.n1081 3.4105
R14865 GNDA.n1119 GNDA.n1081 3.4105
R14866 GNDA.n1946 GNDA.n1081 3.4105
R14867 GNDA.n1118 GNDA.n1081 3.4105
R14868 GNDA.n1948 GNDA.n1081 3.4105
R14869 GNDA.n1117 GNDA.n1081 3.4105
R14870 GNDA.n1950 GNDA.n1081 3.4105
R14871 GNDA.n1116 GNDA.n1081 3.4105
R14872 GNDA.n1952 GNDA.n1081 3.4105
R14873 GNDA.n1115 GNDA.n1081 3.4105
R14874 GNDA.n1954 GNDA.n1081 3.4105
R14875 GNDA.n1114 GNDA.n1081 3.4105
R14876 GNDA.n1956 GNDA.n1081 3.4105
R14877 GNDA.n1081 GNDA.n1045 3.4105
R14878 GNDA.n1959 GNDA.n1081 3.4105
R14879 GNDA.n1926 GNDA.n1053 3.4105
R14880 GNDA.n1128 GNDA.n1053 3.4105
R14881 GNDA.n1928 GNDA.n1053 3.4105
R14882 GNDA.n1127 GNDA.n1053 3.4105
R14883 GNDA.n1930 GNDA.n1053 3.4105
R14884 GNDA.n1126 GNDA.n1053 3.4105
R14885 GNDA.n1932 GNDA.n1053 3.4105
R14886 GNDA.n1125 GNDA.n1053 3.4105
R14887 GNDA.n1934 GNDA.n1053 3.4105
R14888 GNDA.n1124 GNDA.n1053 3.4105
R14889 GNDA.n1936 GNDA.n1053 3.4105
R14890 GNDA.n1123 GNDA.n1053 3.4105
R14891 GNDA.n1938 GNDA.n1053 3.4105
R14892 GNDA.n1122 GNDA.n1053 3.4105
R14893 GNDA.n1940 GNDA.n1053 3.4105
R14894 GNDA.n1121 GNDA.n1053 3.4105
R14895 GNDA.n1942 GNDA.n1053 3.4105
R14896 GNDA.n1120 GNDA.n1053 3.4105
R14897 GNDA.n1944 GNDA.n1053 3.4105
R14898 GNDA.n1119 GNDA.n1053 3.4105
R14899 GNDA.n1946 GNDA.n1053 3.4105
R14900 GNDA.n1118 GNDA.n1053 3.4105
R14901 GNDA.n1948 GNDA.n1053 3.4105
R14902 GNDA.n1117 GNDA.n1053 3.4105
R14903 GNDA.n1950 GNDA.n1053 3.4105
R14904 GNDA.n1116 GNDA.n1053 3.4105
R14905 GNDA.n1952 GNDA.n1053 3.4105
R14906 GNDA.n1115 GNDA.n1053 3.4105
R14907 GNDA.n1954 GNDA.n1053 3.4105
R14908 GNDA.n1114 GNDA.n1053 3.4105
R14909 GNDA.n1956 GNDA.n1053 3.4105
R14910 GNDA.n1053 GNDA.n1045 3.4105
R14911 GNDA.n1959 GNDA.n1053 3.4105
R14912 GNDA.n1926 GNDA.n1083 3.4105
R14913 GNDA.n1128 GNDA.n1083 3.4105
R14914 GNDA.n1928 GNDA.n1083 3.4105
R14915 GNDA.n1127 GNDA.n1083 3.4105
R14916 GNDA.n1930 GNDA.n1083 3.4105
R14917 GNDA.n1126 GNDA.n1083 3.4105
R14918 GNDA.n1932 GNDA.n1083 3.4105
R14919 GNDA.n1125 GNDA.n1083 3.4105
R14920 GNDA.n1934 GNDA.n1083 3.4105
R14921 GNDA.n1124 GNDA.n1083 3.4105
R14922 GNDA.n1936 GNDA.n1083 3.4105
R14923 GNDA.n1123 GNDA.n1083 3.4105
R14924 GNDA.n1938 GNDA.n1083 3.4105
R14925 GNDA.n1122 GNDA.n1083 3.4105
R14926 GNDA.n1940 GNDA.n1083 3.4105
R14927 GNDA.n1121 GNDA.n1083 3.4105
R14928 GNDA.n1942 GNDA.n1083 3.4105
R14929 GNDA.n1120 GNDA.n1083 3.4105
R14930 GNDA.n1944 GNDA.n1083 3.4105
R14931 GNDA.n1119 GNDA.n1083 3.4105
R14932 GNDA.n1946 GNDA.n1083 3.4105
R14933 GNDA.n1118 GNDA.n1083 3.4105
R14934 GNDA.n1948 GNDA.n1083 3.4105
R14935 GNDA.n1117 GNDA.n1083 3.4105
R14936 GNDA.n1950 GNDA.n1083 3.4105
R14937 GNDA.n1116 GNDA.n1083 3.4105
R14938 GNDA.n1952 GNDA.n1083 3.4105
R14939 GNDA.n1115 GNDA.n1083 3.4105
R14940 GNDA.n1954 GNDA.n1083 3.4105
R14941 GNDA.n1114 GNDA.n1083 3.4105
R14942 GNDA.n1956 GNDA.n1083 3.4105
R14943 GNDA.n1083 GNDA.n1045 3.4105
R14944 GNDA.n1959 GNDA.n1083 3.4105
R14945 GNDA.n1926 GNDA.n1052 3.4105
R14946 GNDA.n1128 GNDA.n1052 3.4105
R14947 GNDA.n1928 GNDA.n1052 3.4105
R14948 GNDA.n1127 GNDA.n1052 3.4105
R14949 GNDA.n1930 GNDA.n1052 3.4105
R14950 GNDA.n1126 GNDA.n1052 3.4105
R14951 GNDA.n1932 GNDA.n1052 3.4105
R14952 GNDA.n1125 GNDA.n1052 3.4105
R14953 GNDA.n1934 GNDA.n1052 3.4105
R14954 GNDA.n1124 GNDA.n1052 3.4105
R14955 GNDA.n1936 GNDA.n1052 3.4105
R14956 GNDA.n1123 GNDA.n1052 3.4105
R14957 GNDA.n1938 GNDA.n1052 3.4105
R14958 GNDA.n1122 GNDA.n1052 3.4105
R14959 GNDA.n1940 GNDA.n1052 3.4105
R14960 GNDA.n1121 GNDA.n1052 3.4105
R14961 GNDA.n1942 GNDA.n1052 3.4105
R14962 GNDA.n1120 GNDA.n1052 3.4105
R14963 GNDA.n1944 GNDA.n1052 3.4105
R14964 GNDA.n1119 GNDA.n1052 3.4105
R14965 GNDA.n1946 GNDA.n1052 3.4105
R14966 GNDA.n1118 GNDA.n1052 3.4105
R14967 GNDA.n1948 GNDA.n1052 3.4105
R14968 GNDA.n1117 GNDA.n1052 3.4105
R14969 GNDA.n1950 GNDA.n1052 3.4105
R14970 GNDA.n1116 GNDA.n1052 3.4105
R14971 GNDA.n1952 GNDA.n1052 3.4105
R14972 GNDA.n1115 GNDA.n1052 3.4105
R14973 GNDA.n1954 GNDA.n1052 3.4105
R14974 GNDA.n1114 GNDA.n1052 3.4105
R14975 GNDA.n1956 GNDA.n1052 3.4105
R14976 GNDA.n1052 GNDA.n1045 3.4105
R14977 GNDA.n1959 GNDA.n1052 3.4105
R14978 GNDA.n1926 GNDA.n1085 3.4105
R14979 GNDA.n1128 GNDA.n1085 3.4105
R14980 GNDA.n1928 GNDA.n1085 3.4105
R14981 GNDA.n1127 GNDA.n1085 3.4105
R14982 GNDA.n1930 GNDA.n1085 3.4105
R14983 GNDA.n1126 GNDA.n1085 3.4105
R14984 GNDA.n1932 GNDA.n1085 3.4105
R14985 GNDA.n1125 GNDA.n1085 3.4105
R14986 GNDA.n1934 GNDA.n1085 3.4105
R14987 GNDA.n1124 GNDA.n1085 3.4105
R14988 GNDA.n1936 GNDA.n1085 3.4105
R14989 GNDA.n1123 GNDA.n1085 3.4105
R14990 GNDA.n1938 GNDA.n1085 3.4105
R14991 GNDA.n1122 GNDA.n1085 3.4105
R14992 GNDA.n1940 GNDA.n1085 3.4105
R14993 GNDA.n1121 GNDA.n1085 3.4105
R14994 GNDA.n1942 GNDA.n1085 3.4105
R14995 GNDA.n1120 GNDA.n1085 3.4105
R14996 GNDA.n1944 GNDA.n1085 3.4105
R14997 GNDA.n1119 GNDA.n1085 3.4105
R14998 GNDA.n1946 GNDA.n1085 3.4105
R14999 GNDA.n1118 GNDA.n1085 3.4105
R15000 GNDA.n1948 GNDA.n1085 3.4105
R15001 GNDA.n1117 GNDA.n1085 3.4105
R15002 GNDA.n1950 GNDA.n1085 3.4105
R15003 GNDA.n1116 GNDA.n1085 3.4105
R15004 GNDA.n1952 GNDA.n1085 3.4105
R15005 GNDA.n1115 GNDA.n1085 3.4105
R15006 GNDA.n1954 GNDA.n1085 3.4105
R15007 GNDA.n1114 GNDA.n1085 3.4105
R15008 GNDA.n1956 GNDA.n1085 3.4105
R15009 GNDA.n1085 GNDA.n1045 3.4105
R15010 GNDA.n1959 GNDA.n1085 3.4105
R15011 GNDA.n1926 GNDA.n1051 3.4105
R15012 GNDA.n1128 GNDA.n1051 3.4105
R15013 GNDA.n1928 GNDA.n1051 3.4105
R15014 GNDA.n1127 GNDA.n1051 3.4105
R15015 GNDA.n1930 GNDA.n1051 3.4105
R15016 GNDA.n1126 GNDA.n1051 3.4105
R15017 GNDA.n1932 GNDA.n1051 3.4105
R15018 GNDA.n1125 GNDA.n1051 3.4105
R15019 GNDA.n1934 GNDA.n1051 3.4105
R15020 GNDA.n1124 GNDA.n1051 3.4105
R15021 GNDA.n1936 GNDA.n1051 3.4105
R15022 GNDA.n1123 GNDA.n1051 3.4105
R15023 GNDA.n1938 GNDA.n1051 3.4105
R15024 GNDA.n1122 GNDA.n1051 3.4105
R15025 GNDA.n1940 GNDA.n1051 3.4105
R15026 GNDA.n1121 GNDA.n1051 3.4105
R15027 GNDA.n1942 GNDA.n1051 3.4105
R15028 GNDA.n1120 GNDA.n1051 3.4105
R15029 GNDA.n1944 GNDA.n1051 3.4105
R15030 GNDA.n1119 GNDA.n1051 3.4105
R15031 GNDA.n1946 GNDA.n1051 3.4105
R15032 GNDA.n1118 GNDA.n1051 3.4105
R15033 GNDA.n1948 GNDA.n1051 3.4105
R15034 GNDA.n1117 GNDA.n1051 3.4105
R15035 GNDA.n1950 GNDA.n1051 3.4105
R15036 GNDA.n1116 GNDA.n1051 3.4105
R15037 GNDA.n1952 GNDA.n1051 3.4105
R15038 GNDA.n1115 GNDA.n1051 3.4105
R15039 GNDA.n1954 GNDA.n1051 3.4105
R15040 GNDA.n1114 GNDA.n1051 3.4105
R15041 GNDA.n1956 GNDA.n1051 3.4105
R15042 GNDA.n1051 GNDA.n1045 3.4105
R15043 GNDA.n1959 GNDA.n1051 3.4105
R15044 GNDA.n1926 GNDA.n1087 3.4105
R15045 GNDA.n1128 GNDA.n1087 3.4105
R15046 GNDA.n1928 GNDA.n1087 3.4105
R15047 GNDA.n1127 GNDA.n1087 3.4105
R15048 GNDA.n1930 GNDA.n1087 3.4105
R15049 GNDA.n1126 GNDA.n1087 3.4105
R15050 GNDA.n1932 GNDA.n1087 3.4105
R15051 GNDA.n1125 GNDA.n1087 3.4105
R15052 GNDA.n1934 GNDA.n1087 3.4105
R15053 GNDA.n1124 GNDA.n1087 3.4105
R15054 GNDA.n1936 GNDA.n1087 3.4105
R15055 GNDA.n1123 GNDA.n1087 3.4105
R15056 GNDA.n1938 GNDA.n1087 3.4105
R15057 GNDA.n1122 GNDA.n1087 3.4105
R15058 GNDA.n1940 GNDA.n1087 3.4105
R15059 GNDA.n1121 GNDA.n1087 3.4105
R15060 GNDA.n1942 GNDA.n1087 3.4105
R15061 GNDA.n1120 GNDA.n1087 3.4105
R15062 GNDA.n1944 GNDA.n1087 3.4105
R15063 GNDA.n1119 GNDA.n1087 3.4105
R15064 GNDA.n1946 GNDA.n1087 3.4105
R15065 GNDA.n1118 GNDA.n1087 3.4105
R15066 GNDA.n1948 GNDA.n1087 3.4105
R15067 GNDA.n1117 GNDA.n1087 3.4105
R15068 GNDA.n1950 GNDA.n1087 3.4105
R15069 GNDA.n1116 GNDA.n1087 3.4105
R15070 GNDA.n1952 GNDA.n1087 3.4105
R15071 GNDA.n1115 GNDA.n1087 3.4105
R15072 GNDA.n1954 GNDA.n1087 3.4105
R15073 GNDA.n1114 GNDA.n1087 3.4105
R15074 GNDA.n1956 GNDA.n1087 3.4105
R15075 GNDA.n1087 GNDA.n1045 3.4105
R15076 GNDA.n1959 GNDA.n1087 3.4105
R15077 GNDA.n1926 GNDA.n1050 3.4105
R15078 GNDA.n1128 GNDA.n1050 3.4105
R15079 GNDA.n1928 GNDA.n1050 3.4105
R15080 GNDA.n1127 GNDA.n1050 3.4105
R15081 GNDA.n1930 GNDA.n1050 3.4105
R15082 GNDA.n1126 GNDA.n1050 3.4105
R15083 GNDA.n1932 GNDA.n1050 3.4105
R15084 GNDA.n1125 GNDA.n1050 3.4105
R15085 GNDA.n1934 GNDA.n1050 3.4105
R15086 GNDA.n1124 GNDA.n1050 3.4105
R15087 GNDA.n1936 GNDA.n1050 3.4105
R15088 GNDA.n1123 GNDA.n1050 3.4105
R15089 GNDA.n1938 GNDA.n1050 3.4105
R15090 GNDA.n1122 GNDA.n1050 3.4105
R15091 GNDA.n1940 GNDA.n1050 3.4105
R15092 GNDA.n1121 GNDA.n1050 3.4105
R15093 GNDA.n1942 GNDA.n1050 3.4105
R15094 GNDA.n1120 GNDA.n1050 3.4105
R15095 GNDA.n1944 GNDA.n1050 3.4105
R15096 GNDA.n1119 GNDA.n1050 3.4105
R15097 GNDA.n1946 GNDA.n1050 3.4105
R15098 GNDA.n1118 GNDA.n1050 3.4105
R15099 GNDA.n1948 GNDA.n1050 3.4105
R15100 GNDA.n1117 GNDA.n1050 3.4105
R15101 GNDA.n1950 GNDA.n1050 3.4105
R15102 GNDA.n1116 GNDA.n1050 3.4105
R15103 GNDA.n1952 GNDA.n1050 3.4105
R15104 GNDA.n1115 GNDA.n1050 3.4105
R15105 GNDA.n1954 GNDA.n1050 3.4105
R15106 GNDA.n1114 GNDA.n1050 3.4105
R15107 GNDA.n1956 GNDA.n1050 3.4105
R15108 GNDA.n1050 GNDA.n1045 3.4105
R15109 GNDA.n1959 GNDA.n1050 3.4105
R15110 GNDA.n1926 GNDA.n1089 3.4105
R15111 GNDA.n1128 GNDA.n1089 3.4105
R15112 GNDA.n1928 GNDA.n1089 3.4105
R15113 GNDA.n1127 GNDA.n1089 3.4105
R15114 GNDA.n1930 GNDA.n1089 3.4105
R15115 GNDA.n1126 GNDA.n1089 3.4105
R15116 GNDA.n1932 GNDA.n1089 3.4105
R15117 GNDA.n1125 GNDA.n1089 3.4105
R15118 GNDA.n1934 GNDA.n1089 3.4105
R15119 GNDA.n1124 GNDA.n1089 3.4105
R15120 GNDA.n1936 GNDA.n1089 3.4105
R15121 GNDA.n1123 GNDA.n1089 3.4105
R15122 GNDA.n1938 GNDA.n1089 3.4105
R15123 GNDA.n1122 GNDA.n1089 3.4105
R15124 GNDA.n1940 GNDA.n1089 3.4105
R15125 GNDA.n1121 GNDA.n1089 3.4105
R15126 GNDA.n1942 GNDA.n1089 3.4105
R15127 GNDA.n1120 GNDA.n1089 3.4105
R15128 GNDA.n1944 GNDA.n1089 3.4105
R15129 GNDA.n1119 GNDA.n1089 3.4105
R15130 GNDA.n1946 GNDA.n1089 3.4105
R15131 GNDA.n1118 GNDA.n1089 3.4105
R15132 GNDA.n1948 GNDA.n1089 3.4105
R15133 GNDA.n1117 GNDA.n1089 3.4105
R15134 GNDA.n1950 GNDA.n1089 3.4105
R15135 GNDA.n1116 GNDA.n1089 3.4105
R15136 GNDA.n1952 GNDA.n1089 3.4105
R15137 GNDA.n1115 GNDA.n1089 3.4105
R15138 GNDA.n1954 GNDA.n1089 3.4105
R15139 GNDA.n1114 GNDA.n1089 3.4105
R15140 GNDA.n1956 GNDA.n1089 3.4105
R15141 GNDA.n1089 GNDA.n1045 3.4105
R15142 GNDA.n1959 GNDA.n1089 3.4105
R15143 GNDA.n1926 GNDA.n1049 3.4105
R15144 GNDA.n1128 GNDA.n1049 3.4105
R15145 GNDA.n1928 GNDA.n1049 3.4105
R15146 GNDA.n1127 GNDA.n1049 3.4105
R15147 GNDA.n1930 GNDA.n1049 3.4105
R15148 GNDA.n1126 GNDA.n1049 3.4105
R15149 GNDA.n1932 GNDA.n1049 3.4105
R15150 GNDA.n1125 GNDA.n1049 3.4105
R15151 GNDA.n1934 GNDA.n1049 3.4105
R15152 GNDA.n1124 GNDA.n1049 3.4105
R15153 GNDA.n1936 GNDA.n1049 3.4105
R15154 GNDA.n1123 GNDA.n1049 3.4105
R15155 GNDA.n1938 GNDA.n1049 3.4105
R15156 GNDA.n1122 GNDA.n1049 3.4105
R15157 GNDA.n1940 GNDA.n1049 3.4105
R15158 GNDA.n1121 GNDA.n1049 3.4105
R15159 GNDA.n1942 GNDA.n1049 3.4105
R15160 GNDA.n1120 GNDA.n1049 3.4105
R15161 GNDA.n1944 GNDA.n1049 3.4105
R15162 GNDA.n1119 GNDA.n1049 3.4105
R15163 GNDA.n1946 GNDA.n1049 3.4105
R15164 GNDA.n1118 GNDA.n1049 3.4105
R15165 GNDA.n1948 GNDA.n1049 3.4105
R15166 GNDA.n1117 GNDA.n1049 3.4105
R15167 GNDA.n1950 GNDA.n1049 3.4105
R15168 GNDA.n1116 GNDA.n1049 3.4105
R15169 GNDA.n1952 GNDA.n1049 3.4105
R15170 GNDA.n1115 GNDA.n1049 3.4105
R15171 GNDA.n1954 GNDA.n1049 3.4105
R15172 GNDA.n1114 GNDA.n1049 3.4105
R15173 GNDA.n1956 GNDA.n1049 3.4105
R15174 GNDA.n1049 GNDA.n1045 3.4105
R15175 GNDA.n1959 GNDA.n1049 3.4105
R15176 GNDA.n1926 GNDA.n1091 3.4105
R15177 GNDA.n1128 GNDA.n1091 3.4105
R15178 GNDA.n1928 GNDA.n1091 3.4105
R15179 GNDA.n1127 GNDA.n1091 3.4105
R15180 GNDA.n1930 GNDA.n1091 3.4105
R15181 GNDA.n1126 GNDA.n1091 3.4105
R15182 GNDA.n1932 GNDA.n1091 3.4105
R15183 GNDA.n1125 GNDA.n1091 3.4105
R15184 GNDA.n1934 GNDA.n1091 3.4105
R15185 GNDA.n1124 GNDA.n1091 3.4105
R15186 GNDA.n1936 GNDA.n1091 3.4105
R15187 GNDA.n1123 GNDA.n1091 3.4105
R15188 GNDA.n1938 GNDA.n1091 3.4105
R15189 GNDA.n1122 GNDA.n1091 3.4105
R15190 GNDA.n1940 GNDA.n1091 3.4105
R15191 GNDA.n1121 GNDA.n1091 3.4105
R15192 GNDA.n1942 GNDA.n1091 3.4105
R15193 GNDA.n1120 GNDA.n1091 3.4105
R15194 GNDA.n1944 GNDA.n1091 3.4105
R15195 GNDA.n1119 GNDA.n1091 3.4105
R15196 GNDA.n1946 GNDA.n1091 3.4105
R15197 GNDA.n1118 GNDA.n1091 3.4105
R15198 GNDA.n1948 GNDA.n1091 3.4105
R15199 GNDA.n1117 GNDA.n1091 3.4105
R15200 GNDA.n1950 GNDA.n1091 3.4105
R15201 GNDA.n1116 GNDA.n1091 3.4105
R15202 GNDA.n1952 GNDA.n1091 3.4105
R15203 GNDA.n1115 GNDA.n1091 3.4105
R15204 GNDA.n1954 GNDA.n1091 3.4105
R15205 GNDA.n1114 GNDA.n1091 3.4105
R15206 GNDA.n1956 GNDA.n1091 3.4105
R15207 GNDA.n1091 GNDA.n1045 3.4105
R15208 GNDA.n1959 GNDA.n1091 3.4105
R15209 GNDA.n1926 GNDA.n1048 3.4105
R15210 GNDA.n1128 GNDA.n1048 3.4105
R15211 GNDA.n1928 GNDA.n1048 3.4105
R15212 GNDA.n1127 GNDA.n1048 3.4105
R15213 GNDA.n1930 GNDA.n1048 3.4105
R15214 GNDA.n1126 GNDA.n1048 3.4105
R15215 GNDA.n1932 GNDA.n1048 3.4105
R15216 GNDA.n1125 GNDA.n1048 3.4105
R15217 GNDA.n1934 GNDA.n1048 3.4105
R15218 GNDA.n1124 GNDA.n1048 3.4105
R15219 GNDA.n1936 GNDA.n1048 3.4105
R15220 GNDA.n1123 GNDA.n1048 3.4105
R15221 GNDA.n1938 GNDA.n1048 3.4105
R15222 GNDA.n1122 GNDA.n1048 3.4105
R15223 GNDA.n1940 GNDA.n1048 3.4105
R15224 GNDA.n1121 GNDA.n1048 3.4105
R15225 GNDA.n1942 GNDA.n1048 3.4105
R15226 GNDA.n1120 GNDA.n1048 3.4105
R15227 GNDA.n1944 GNDA.n1048 3.4105
R15228 GNDA.n1119 GNDA.n1048 3.4105
R15229 GNDA.n1946 GNDA.n1048 3.4105
R15230 GNDA.n1118 GNDA.n1048 3.4105
R15231 GNDA.n1948 GNDA.n1048 3.4105
R15232 GNDA.n1117 GNDA.n1048 3.4105
R15233 GNDA.n1950 GNDA.n1048 3.4105
R15234 GNDA.n1116 GNDA.n1048 3.4105
R15235 GNDA.n1952 GNDA.n1048 3.4105
R15236 GNDA.n1115 GNDA.n1048 3.4105
R15237 GNDA.n1954 GNDA.n1048 3.4105
R15238 GNDA.n1114 GNDA.n1048 3.4105
R15239 GNDA.n1956 GNDA.n1048 3.4105
R15240 GNDA.n1048 GNDA.n1045 3.4105
R15241 GNDA.n1959 GNDA.n1048 3.4105
R15242 GNDA.n1926 GNDA.n1093 3.4105
R15243 GNDA.n1128 GNDA.n1093 3.4105
R15244 GNDA.n1928 GNDA.n1093 3.4105
R15245 GNDA.n1127 GNDA.n1093 3.4105
R15246 GNDA.n1930 GNDA.n1093 3.4105
R15247 GNDA.n1126 GNDA.n1093 3.4105
R15248 GNDA.n1932 GNDA.n1093 3.4105
R15249 GNDA.n1125 GNDA.n1093 3.4105
R15250 GNDA.n1934 GNDA.n1093 3.4105
R15251 GNDA.n1124 GNDA.n1093 3.4105
R15252 GNDA.n1936 GNDA.n1093 3.4105
R15253 GNDA.n1123 GNDA.n1093 3.4105
R15254 GNDA.n1938 GNDA.n1093 3.4105
R15255 GNDA.n1122 GNDA.n1093 3.4105
R15256 GNDA.n1940 GNDA.n1093 3.4105
R15257 GNDA.n1121 GNDA.n1093 3.4105
R15258 GNDA.n1942 GNDA.n1093 3.4105
R15259 GNDA.n1120 GNDA.n1093 3.4105
R15260 GNDA.n1944 GNDA.n1093 3.4105
R15261 GNDA.n1119 GNDA.n1093 3.4105
R15262 GNDA.n1946 GNDA.n1093 3.4105
R15263 GNDA.n1118 GNDA.n1093 3.4105
R15264 GNDA.n1948 GNDA.n1093 3.4105
R15265 GNDA.n1117 GNDA.n1093 3.4105
R15266 GNDA.n1950 GNDA.n1093 3.4105
R15267 GNDA.n1116 GNDA.n1093 3.4105
R15268 GNDA.n1952 GNDA.n1093 3.4105
R15269 GNDA.n1115 GNDA.n1093 3.4105
R15270 GNDA.n1954 GNDA.n1093 3.4105
R15271 GNDA.n1114 GNDA.n1093 3.4105
R15272 GNDA.n1956 GNDA.n1093 3.4105
R15273 GNDA.n1093 GNDA.n1045 3.4105
R15274 GNDA.n1959 GNDA.n1093 3.4105
R15275 GNDA.n1926 GNDA.n1047 3.4105
R15276 GNDA.n1128 GNDA.n1047 3.4105
R15277 GNDA.n1928 GNDA.n1047 3.4105
R15278 GNDA.n1127 GNDA.n1047 3.4105
R15279 GNDA.n1930 GNDA.n1047 3.4105
R15280 GNDA.n1126 GNDA.n1047 3.4105
R15281 GNDA.n1932 GNDA.n1047 3.4105
R15282 GNDA.n1125 GNDA.n1047 3.4105
R15283 GNDA.n1934 GNDA.n1047 3.4105
R15284 GNDA.n1124 GNDA.n1047 3.4105
R15285 GNDA.n1936 GNDA.n1047 3.4105
R15286 GNDA.n1123 GNDA.n1047 3.4105
R15287 GNDA.n1938 GNDA.n1047 3.4105
R15288 GNDA.n1122 GNDA.n1047 3.4105
R15289 GNDA.n1940 GNDA.n1047 3.4105
R15290 GNDA.n1121 GNDA.n1047 3.4105
R15291 GNDA.n1942 GNDA.n1047 3.4105
R15292 GNDA.n1120 GNDA.n1047 3.4105
R15293 GNDA.n1944 GNDA.n1047 3.4105
R15294 GNDA.n1119 GNDA.n1047 3.4105
R15295 GNDA.n1946 GNDA.n1047 3.4105
R15296 GNDA.n1118 GNDA.n1047 3.4105
R15297 GNDA.n1948 GNDA.n1047 3.4105
R15298 GNDA.n1117 GNDA.n1047 3.4105
R15299 GNDA.n1950 GNDA.n1047 3.4105
R15300 GNDA.n1116 GNDA.n1047 3.4105
R15301 GNDA.n1952 GNDA.n1047 3.4105
R15302 GNDA.n1115 GNDA.n1047 3.4105
R15303 GNDA.n1954 GNDA.n1047 3.4105
R15304 GNDA.n1114 GNDA.n1047 3.4105
R15305 GNDA.n1956 GNDA.n1047 3.4105
R15306 GNDA.n1047 GNDA.n1045 3.4105
R15307 GNDA.n1959 GNDA.n1047 3.4105
R15308 GNDA.n1926 GNDA.n1095 3.4105
R15309 GNDA.n1128 GNDA.n1095 3.4105
R15310 GNDA.n1928 GNDA.n1095 3.4105
R15311 GNDA.n1127 GNDA.n1095 3.4105
R15312 GNDA.n1930 GNDA.n1095 3.4105
R15313 GNDA.n1126 GNDA.n1095 3.4105
R15314 GNDA.n1932 GNDA.n1095 3.4105
R15315 GNDA.n1125 GNDA.n1095 3.4105
R15316 GNDA.n1934 GNDA.n1095 3.4105
R15317 GNDA.n1124 GNDA.n1095 3.4105
R15318 GNDA.n1936 GNDA.n1095 3.4105
R15319 GNDA.n1123 GNDA.n1095 3.4105
R15320 GNDA.n1938 GNDA.n1095 3.4105
R15321 GNDA.n1122 GNDA.n1095 3.4105
R15322 GNDA.n1940 GNDA.n1095 3.4105
R15323 GNDA.n1121 GNDA.n1095 3.4105
R15324 GNDA.n1942 GNDA.n1095 3.4105
R15325 GNDA.n1120 GNDA.n1095 3.4105
R15326 GNDA.n1944 GNDA.n1095 3.4105
R15327 GNDA.n1119 GNDA.n1095 3.4105
R15328 GNDA.n1946 GNDA.n1095 3.4105
R15329 GNDA.n1118 GNDA.n1095 3.4105
R15330 GNDA.n1948 GNDA.n1095 3.4105
R15331 GNDA.n1117 GNDA.n1095 3.4105
R15332 GNDA.n1950 GNDA.n1095 3.4105
R15333 GNDA.n1116 GNDA.n1095 3.4105
R15334 GNDA.n1952 GNDA.n1095 3.4105
R15335 GNDA.n1115 GNDA.n1095 3.4105
R15336 GNDA.n1954 GNDA.n1095 3.4105
R15337 GNDA.n1114 GNDA.n1095 3.4105
R15338 GNDA.n1956 GNDA.n1095 3.4105
R15339 GNDA.n1095 GNDA.n1045 3.4105
R15340 GNDA.n1959 GNDA.n1095 3.4105
R15341 GNDA.n1926 GNDA.n1046 3.4105
R15342 GNDA.n1128 GNDA.n1046 3.4105
R15343 GNDA.n1928 GNDA.n1046 3.4105
R15344 GNDA.n1127 GNDA.n1046 3.4105
R15345 GNDA.n1930 GNDA.n1046 3.4105
R15346 GNDA.n1126 GNDA.n1046 3.4105
R15347 GNDA.n1932 GNDA.n1046 3.4105
R15348 GNDA.n1125 GNDA.n1046 3.4105
R15349 GNDA.n1934 GNDA.n1046 3.4105
R15350 GNDA.n1124 GNDA.n1046 3.4105
R15351 GNDA.n1936 GNDA.n1046 3.4105
R15352 GNDA.n1123 GNDA.n1046 3.4105
R15353 GNDA.n1938 GNDA.n1046 3.4105
R15354 GNDA.n1122 GNDA.n1046 3.4105
R15355 GNDA.n1940 GNDA.n1046 3.4105
R15356 GNDA.n1121 GNDA.n1046 3.4105
R15357 GNDA.n1942 GNDA.n1046 3.4105
R15358 GNDA.n1120 GNDA.n1046 3.4105
R15359 GNDA.n1944 GNDA.n1046 3.4105
R15360 GNDA.n1119 GNDA.n1046 3.4105
R15361 GNDA.n1946 GNDA.n1046 3.4105
R15362 GNDA.n1118 GNDA.n1046 3.4105
R15363 GNDA.n1948 GNDA.n1046 3.4105
R15364 GNDA.n1117 GNDA.n1046 3.4105
R15365 GNDA.n1950 GNDA.n1046 3.4105
R15366 GNDA.n1116 GNDA.n1046 3.4105
R15367 GNDA.n1952 GNDA.n1046 3.4105
R15368 GNDA.n1115 GNDA.n1046 3.4105
R15369 GNDA.n1954 GNDA.n1046 3.4105
R15370 GNDA.n1114 GNDA.n1046 3.4105
R15371 GNDA.n1956 GNDA.n1046 3.4105
R15372 GNDA.n1046 GNDA.n1045 3.4105
R15373 GNDA.n1959 GNDA.n1046 3.4105
R15374 GNDA.n1958 GNDA.n1926 3.4105
R15375 GNDA.n1958 GNDA.n1128 3.4105
R15376 GNDA.n1958 GNDA.n1928 3.4105
R15377 GNDA.n1958 GNDA.n1127 3.4105
R15378 GNDA.n1958 GNDA.n1930 3.4105
R15379 GNDA.n1958 GNDA.n1126 3.4105
R15380 GNDA.n1958 GNDA.n1932 3.4105
R15381 GNDA.n1958 GNDA.n1125 3.4105
R15382 GNDA.n1958 GNDA.n1934 3.4105
R15383 GNDA.n1958 GNDA.n1124 3.4105
R15384 GNDA.n1958 GNDA.n1936 3.4105
R15385 GNDA.n1958 GNDA.n1123 3.4105
R15386 GNDA.n1958 GNDA.n1938 3.4105
R15387 GNDA.n1958 GNDA.n1122 3.4105
R15388 GNDA.n1958 GNDA.n1940 3.4105
R15389 GNDA.n1958 GNDA.n1121 3.4105
R15390 GNDA.n1958 GNDA.n1942 3.4105
R15391 GNDA.n1958 GNDA.n1120 3.4105
R15392 GNDA.n1958 GNDA.n1944 3.4105
R15393 GNDA.n1958 GNDA.n1119 3.4105
R15394 GNDA.n1958 GNDA.n1946 3.4105
R15395 GNDA.n1958 GNDA.n1118 3.4105
R15396 GNDA.n1958 GNDA.n1948 3.4105
R15397 GNDA.n1958 GNDA.n1117 3.4105
R15398 GNDA.n1958 GNDA.n1950 3.4105
R15399 GNDA.n1958 GNDA.n1116 3.4105
R15400 GNDA.n1958 GNDA.n1952 3.4105
R15401 GNDA.n1958 GNDA.n1115 3.4105
R15402 GNDA.n1958 GNDA.n1954 3.4105
R15403 GNDA.n1958 GNDA.n1114 3.4105
R15404 GNDA.n1958 GNDA.n1956 3.4105
R15405 GNDA.n1959 GNDA.n1958 3.4105
R15406 GNDA.n1027 GNDA.n963 3.4105
R15407 GNDA.n1991 GNDA.n963 3.4105
R15408 GNDA.n2011 GNDA.n963 3.4105
R15409 GNDA.n2010 GNDA.n1962 3.4105
R15410 GNDA.n2010 GNDA.n1026 3.4105
R15411 GNDA.n2010 GNDA.n1964 3.4105
R15412 GNDA.n2010 GNDA.n1025 3.4105
R15413 GNDA.n2010 GNDA.n1966 3.4105
R15414 GNDA.n2010 GNDA.n1024 3.4105
R15415 GNDA.n2010 GNDA.n1968 3.4105
R15416 GNDA.n2010 GNDA.n1023 3.4105
R15417 GNDA.n2010 GNDA.n1970 3.4105
R15418 GNDA.n2010 GNDA.n1022 3.4105
R15419 GNDA.n2010 GNDA.n1972 3.4105
R15420 GNDA.n2010 GNDA.n1021 3.4105
R15421 GNDA.n2010 GNDA.n1974 3.4105
R15422 GNDA.n2010 GNDA.n1020 3.4105
R15423 GNDA.n2010 GNDA.n1976 3.4105
R15424 GNDA.n2010 GNDA.n1019 3.4105
R15425 GNDA.n2010 GNDA.n1978 3.4105
R15426 GNDA.n2010 GNDA.n1018 3.4105
R15427 GNDA.n2010 GNDA.n1980 3.4105
R15428 GNDA.n2010 GNDA.n1017 3.4105
R15429 GNDA.n2010 GNDA.n1982 3.4105
R15430 GNDA.n2010 GNDA.n1016 3.4105
R15431 GNDA.n2010 GNDA.n1984 3.4105
R15432 GNDA.n2010 GNDA.n1015 3.4105
R15433 GNDA.n2010 GNDA.n1986 3.4105
R15434 GNDA.n2010 GNDA.n1014 3.4105
R15435 GNDA.n2010 GNDA.n1988 3.4105
R15436 GNDA.n2010 GNDA.n1013 3.4105
R15437 GNDA.n2010 GNDA.n1990 3.4105
R15438 GNDA.n2010 GNDA.n1991 3.4105
R15439 GNDA.n2011 GNDA.n2010 3.4105
R15440 GNDA.n2013 GNDA.n979 3.4105
R15441 GNDA.n1027 GNDA.n979 3.4105
R15442 GNDA.n1962 GNDA.n979 3.4105
R15443 GNDA.n1026 GNDA.n979 3.4105
R15444 GNDA.n1964 GNDA.n979 3.4105
R15445 GNDA.n1025 GNDA.n979 3.4105
R15446 GNDA.n1966 GNDA.n979 3.4105
R15447 GNDA.n1024 GNDA.n979 3.4105
R15448 GNDA.n1968 GNDA.n979 3.4105
R15449 GNDA.n1023 GNDA.n979 3.4105
R15450 GNDA.n1970 GNDA.n979 3.4105
R15451 GNDA.n1022 GNDA.n979 3.4105
R15452 GNDA.n1972 GNDA.n979 3.4105
R15453 GNDA.n1021 GNDA.n979 3.4105
R15454 GNDA.n1974 GNDA.n979 3.4105
R15455 GNDA.n1020 GNDA.n979 3.4105
R15456 GNDA.n1976 GNDA.n979 3.4105
R15457 GNDA.n1019 GNDA.n979 3.4105
R15458 GNDA.n1978 GNDA.n979 3.4105
R15459 GNDA.n1018 GNDA.n979 3.4105
R15460 GNDA.n1980 GNDA.n979 3.4105
R15461 GNDA.n1017 GNDA.n979 3.4105
R15462 GNDA.n1982 GNDA.n979 3.4105
R15463 GNDA.n1016 GNDA.n979 3.4105
R15464 GNDA.n1984 GNDA.n979 3.4105
R15465 GNDA.n1015 GNDA.n979 3.4105
R15466 GNDA.n1986 GNDA.n979 3.4105
R15467 GNDA.n1014 GNDA.n979 3.4105
R15468 GNDA.n1988 GNDA.n979 3.4105
R15469 GNDA.n1013 GNDA.n979 3.4105
R15470 GNDA.n1990 GNDA.n979 3.4105
R15471 GNDA.n1991 GNDA.n979 3.4105
R15472 GNDA.n2011 GNDA.n979 3.4105
R15473 GNDA.n2013 GNDA.n981 3.4105
R15474 GNDA.n1027 GNDA.n981 3.4105
R15475 GNDA.n1962 GNDA.n981 3.4105
R15476 GNDA.n1026 GNDA.n981 3.4105
R15477 GNDA.n1964 GNDA.n981 3.4105
R15478 GNDA.n1025 GNDA.n981 3.4105
R15479 GNDA.n1966 GNDA.n981 3.4105
R15480 GNDA.n1024 GNDA.n981 3.4105
R15481 GNDA.n1968 GNDA.n981 3.4105
R15482 GNDA.n1023 GNDA.n981 3.4105
R15483 GNDA.n1970 GNDA.n981 3.4105
R15484 GNDA.n1022 GNDA.n981 3.4105
R15485 GNDA.n1972 GNDA.n981 3.4105
R15486 GNDA.n1021 GNDA.n981 3.4105
R15487 GNDA.n1974 GNDA.n981 3.4105
R15488 GNDA.n1020 GNDA.n981 3.4105
R15489 GNDA.n1976 GNDA.n981 3.4105
R15490 GNDA.n1019 GNDA.n981 3.4105
R15491 GNDA.n1978 GNDA.n981 3.4105
R15492 GNDA.n1018 GNDA.n981 3.4105
R15493 GNDA.n1980 GNDA.n981 3.4105
R15494 GNDA.n1017 GNDA.n981 3.4105
R15495 GNDA.n1982 GNDA.n981 3.4105
R15496 GNDA.n1016 GNDA.n981 3.4105
R15497 GNDA.n1984 GNDA.n981 3.4105
R15498 GNDA.n1015 GNDA.n981 3.4105
R15499 GNDA.n1986 GNDA.n981 3.4105
R15500 GNDA.n1014 GNDA.n981 3.4105
R15501 GNDA.n1988 GNDA.n981 3.4105
R15502 GNDA.n1013 GNDA.n981 3.4105
R15503 GNDA.n1990 GNDA.n981 3.4105
R15504 GNDA.n1991 GNDA.n981 3.4105
R15505 GNDA.n2011 GNDA.n981 3.4105
R15506 GNDA.n2013 GNDA.n978 3.4105
R15507 GNDA.n1027 GNDA.n978 3.4105
R15508 GNDA.n1962 GNDA.n978 3.4105
R15509 GNDA.n1026 GNDA.n978 3.4105
R15510 GNDA.n1964 GNDA.n978 3.4105
R15511 GNDA.n1025 GNDA.n978 3.4105
R15512 GNDA.n1966 GNDA.n978 3.4105
R15513 GNDA.n1024 GNDA.n978 3.4105
R15514 GNDA.n1968 GNDA.n978 3.4105
R15515 GNDA.n1023 GNDA.n978 3.4105
R15516 GNDA.n1970 GNDA.n978 3.4105
R15517 GNDA.n1022 GNDA.n978 3.4105
R15518 GNDA.n1972 GNDA.n978 3.4105
R15519 GNDA.n1021 GNDA.n978 3.4105
R15520 GNDA.n1974 GNDA.n978 3.4105
R15521 GNDA.n1020 GNDA.n978 3.4105
R15522 GNDA.n1976 GNDA.n978 3.4105
R15523 GNDA.n1019 GNDA.n978 3.4105
R15524 GNDA.n1978 GNDA.n978 3.4105
R15525 GNDA.n1018 GNDA.n978 3.4105
R15526 GNDA.n1980 GNDA.n978 3.4105
R15527 GNDA.n1017 GNDA.n978 3.4105
R15528 GNDA.n1982 GNDA.n978 3.4105
R15529 GNDA.n1016 GNDA.n978 3.4105
R15530 GNDA.n1984 GNDA.n978 3.4105
R15531 GNDA.n1015 GNDA.n978 3.4105
R15532 GNDA.n1986 GNDA.n978 3.4105
R15533 GNDA.n1014 GNDA.n978 3.4105
R15534 GNDA.n1988 GNDA.n978 3.4105
R15535 GNDA.n1013 GNDA.n978 3.4105
R15536 GNDA.n1990 GNDA.n978 3.4105
R15537 GNDA.n1991 GNDA.n978 3.4105
R15538 GNDA.n2011 GNDA.n978 3.4105
R15539 GNDA.n2013 GNDA.n982 3.4105
R15540 GNDA.n1027 GNDA.n982 3.4105
R15541 GNDA.n1962 GNDA.n982 3.4105
R15542 GNDA.n1026 GNDA.n982 3.4105
R15543 GNDA.n1964 GNDA.n982 3.4105
R15544 GNDA.n1025 GNDA.n982 3.4105
R15545 GNDA.n1966 GNDA.n982 3.4105
R15546 GNDA.n1024 GNDA.n982 3.4105
R15547 GNDA.n1968 GNDA.n982 3.4105
R15548 GNDA.n1023 GNDA.n982 3.4105
R15549 GNDA.n1970 GNDA.n982 3.4105
R15550 GNDA.n1022 GNDA.n982 3.4105
R15551 GNDA.n1972 GNDA.n982 3.4105
R15552 GNDA.n1021 GNDA.n982 3.4105
R15553 GNDA.n1974 GNDA.n982 3.4105
R15554 GNDA.n1020 GNDA.n982 3.4105
R15555 GNDA.n1976 GNDA.n982 3.4105
R15556 GNDA.n1019 GNDA.n982 3.4105
R15557 GNDA.n1978 GNDA.n982 3.4105
R15558 GNDA.n1018 GNDA.n982 3.4105
R15559 GNDA.n1980 GNDA.n982 3.4105
R15560 GNDA.n1017 GNDA.n982 3.4105
R15561 GNDA.n1982 GNDA.n982 3.4105
R15562 GNDA.n1016 GNDA.n982 3.4105
R15563 GNDA.n1984 GNDA.n982 3.4105
R15564 GNDA.n1015 GNDA.n982 3.4105
R15565 GNDA.n1986 GNDA.n982 3.4105
R15566 GNDA.n1014 GNDA.n982 3.4105
R15567 GNDA.n1988 GNDA.n982 3.4105
R15568 GNDA.n1013 GNDA.n982 3.4105
R15569 GNDA.n1990 GNDA.n982 3.4105
R15570 GNDA.n1991 GNDA.n982 3.4105
R15571 GNDA.n2011 GNDA.n982 3.4105
R15572 GNDA.n2013 GNDA.n977 3.4105
R15573 GNDA.n1027 GNDA.n977 3.4105
R15574 GNDA.n1962 GNDA.n977 3.4105
R15575 GNDA.n1026 GNDA.n977 3.4105
R15576 GNDA.n1964 GNDA.n977 3.4105
R15577 GNDA.n1025 GNDA.n977 3.4105
R15578 GNDA.n1966 GNDA.n977 3.4105
R15579 GNDA.n1024 GNDA.n977 3.4105
R15580 GNDA.n1968 GNDA.n977 3.4105
R15581 GNDA.n1023 GNDA.n977 3.4105
R15582 GNDA.n1970 GNDA.n977 3.4105
R15583 GNDA.n1022 GNDA.n977 3.4105
R15584 GNDA.n1972 GNDA.n977 3.4105
R15585 GNDA.n1021 GNDA.n977 3.4105
R15586 GNDA.n1974 GNDA.n977 3.4105
R15587 GNDA.n1020 GNDA.n977 3.4105
R15588 GNDA.n1976 GNDA.n977 3.4105
R15589 GNDA.n1019 GNDA.n977 3.4105
R15590 GNDA.n1978 GNDA.n977 3.4105
R15591 GNDA.n1018 GNDA.n977 3.4105
R15592 GNDA.n1980 GNDA.n977 3.4105
R15593 GNDA.n1017 GNDA.n977 3.4105
R15594 GNDA.n1982 GNDA.n977 3.4105
R15595 GNDA.n1016 GNDA.n977 3.4105
R15596 GNDA.n1984 GNDA.n977 3.4105
R15597 GNDA.n1015 GNDA.n977 3.4105
R15598 GNDA.n1986 GNDA.n977 3.4105
R15599 GNDA.n1014 GNDA.n977 3.4105
R15600 GNDA.n1988 GNDA.n977 3.4105
R15601 GNDA.n1013 GNDA.n977 3.4105
R15602 GNDA.n1990 GNDA.n977 3.4105
R15603 GNDA.n1991 GNDA.n977 3.4105
R15604 GNDA.n2011 GNDA.n977 3.4105
R15605 GNDA.n2013 GNDA.n983 3.4105
R15606 GNDA.n1027 GNDA.n983 3.4105
R15607 GNDA.n1962 GNDA.n983 3.4105
R15608 GNDA.n1026 GNDA.n983 3.4105
R15609 GNDA.n1964 GNDA.n983 3.4105
R15610 GNDA.n1025 GNDA.n983 3.4105
R15611 GNDA.n1966 GNDA.n983 3.4105
R15612 GNDA.n1024 GNDA.n983 3.4105
R15613 GNDA.n1968 GNDA.n983 3.4105
R15614 GNDA.n1023 GNDA.n983 3.4105
R15615 GNDA.n1970 GNDA.n983 3.4105
R15616 GNDA.n1022 GNDA.n983 3.4105
R15617 GNDA.n1972 GNDA.n983 3.4105
R15618 GNDA.n1021 GNDA.n983 3.4105
R15619 GNDA.n1974 GNDA.n983 3.4105
R15620 GNDA.n1020 GNDA.n983 3.4105
R15621 GNDA.n1976 GNDA.n983 3.4105
R15622 GNDA.n1019 GNDA.n983 3.4105
R15623 GNDA.n1978 GNDA.n983 3.4105
R15624 GNDA.n1018 GNDA.n983 3.4105
R15625 GNDA.n1980 GNDA.n983 3.4105
R15626 GNDA.n1017 GNDA.n983 3.4105
R15627 GNDA.n1982 GNDA.n983 3.4105
R15628 GNDA.n1016 GNDA.n983 3.4105
R15629 GNDA.n1984 GNDA.n983 3.4105
R15630 GNDA.n1015 GNDA.n983 3.4105
R15631 GNDA.n1986 GNDA.n983 3.4105
R15632 GNDA.n1014 GNDA.n983 3.4105
R15633 GNDA.n1988 GNDA.n983 3.4105
R15634 GNDA.n1013 GNDA.n983 3.4105
R15635 GNDA.n1990 GNDA.n983 3.4105
R15636 GNDA.n1991 GNDA.n983 3.4105
R15637 GNDA.n2011 GNDA.n983 3.4105
R15638 GNDA.n2013 GNDA.n976 3.4105
R15639 GNDA.n1027 GNDA.n976 3.4105
R15640 GNDA.n1962 GNDA.n976 3.4105
R15641 GNDA.n1026 GNDA.n976 3.4105
R15642 GNDA.n1964 GNDA.n976 3.4105
R15643 GNDA.n1025 GNDA.n976 3.4105
R15644 GNDA.n1966 GNDA.n976 3.4105
R15645 GNDA.n1024 GNDA.n976 3.4105
R15646 GNDA.n1968 GNDA.n976 3.4105
R15647 GNDA.n1023 GNDA.n976 3.4105
R15648 GNDA.n1970 GNDA.n976 3.4105
R15649 GNDA.n1022 GNDA.n976 3.4105
R15650 GNDA.n1972 GNDA.n976 3.4105
R15651 GNDA.n1021 GNDA.n976 3.4105
R15652 GNDA.n1974 GNDA.n976 3.4105
R15653 GNDA.n1020 GNDA.n976 3.4105
R15654 GNDA.n1976 GNDA.n976 3.4105
R15655 GNDA.n1019 GNDA.n976 3.4105
R15656 GNDA.n1978 GNDA.n976 3.4105
R15657 GNDA.n1018 GNDA.n976 3.4105
R15658 GNDA.n1980 GNDA.n976 3.4105
R15659 GNDA.n1017 GNDA.n976 3.4105
R15660 GNDA.n1982 GNDA.n976 3.4105
R15661 GNDA.n1016 GNDA.n976 3.4105
R15662 GNDA.n1984 GNDA.n976 3.4105
R15663 GNDA.n1015 GNDA.n976 3.4105
R15664 GNDA.n1986 GNDA.n976 3.4105
R15665 GNDA.n1014 GNDA.n976 3.4105
R15666 GNDA.n1988 GNDA.n976 3.4105
R15667 GNDA.n1013 GNDA.n976 3.4105
R15668 GNDA.n1990 GNDA.n976 3.4105
R15669 GNDA.n1991 GNDA.n976 3.4105
R15670 GNDA.n2011 GNDA.n976 3.4105
R15671 GNDA.n2013 GNDA.n984 3.4105
R15672 GNDA.n1027 GNDA.n984 3.4105
R15673 GNDA.n1962 GNDA.n984 3.4105
R15674 GNDA.n1026 GNDA.n984 3.4105
R15675 GNDA.n1964 GNDA.n984 3.4105
R15676 GNDA.n1025 GNDA.n984 3.4105
R15677 GNDA.n1966 GNDA.n984 3.4105
R15678 GNDA.n1024 GNDA.n984 3.4105
R15679 GNDA.n1968 GNDA.n984 3.4105
R15680 GNDA.n1023 GNDA.n984 3.4105
R15681 GNDA.n1970 GNDA.n984 3.4105
R15682 GNDA.n1022 GNDA.n984 3.4105
R15683 GNDA.n1972 GNDA.n984 3.4105
R15684 GNDA.n1021 GNDA.n984 3.4105
R15685 GNDA.n1974 GNDA.n984 3.4105
R15686 GNDA.n1020 GNDA.n984 3.4105
R15687 GNDA.n1976 GNDA.n984 3.4105
R15688 GNDA.n1019 GNDA.n984 3.4105
R15689 GNDA.n1978 GNDA.n984 3.4105
R15690 GNDA.n1018 GNDA.n984 3.4105
R15691 GNDA.n1980 GNDA.n984 3.4105
R15692 GNDA.n1017 GNDA.n984 3.4105
R15693 GNDA.n1982 GNDA.n984 3.4105
R15694 GNDA.n1016 GNDA.n984 3.4105
R15695 GNDA.n1984 GNDA.n984 3.4105
R15696 GNDA.n1015 GNDA.n984 3.4105
R15697 GNDA.n1986 GNDA.n984 3.4105
R15698 GNDA.n1014 GNDA.n984 3.4105
R15699 GNDA.n1988 GNDA.n984 3.4105
R15700 GNDA.n1013 GNDA.n984 3.4105
R15701 GNDA.n1990 GNDA.n984 3.4105
R15702 GNDA.n1991 GNDA.n984 3.4105
R15703 GNDA.n2011 GNDA.n984 3.4105
R15704 GNDA.n2013 GNDA.n975 3.4105
R15705 GNDA.n1027 GNDA.n975 3.4105
R15706 GNDA.n1962 GNDA.n975 3.4105
R15707 GNDA.n1026 GNDA.n975 3.4105
R15708 GNDA.n1964 GNDA.n975 3.4105
R15709 GNDA.n1025 GNDA.n975 3.4105
R15710 GNDA.n1966 GNDA.n975 3.4105
R15711 GNDA.n1024 GNDA.n975 3.4105
R15712 GNDA.n1968 GNDA.n975 3.4105
R15713 GNDA.n1023 GNDA.n975 3.4105
R15714 GNDA.n1970 GNDA.n975 3.4105
R15715 GNDA.n1022 GNDA.n975 3.4105
R15716 GNDA.n1972 GNDA.n975 3.4105
R15717 GNDA.n1021 GNDA.n975 3.4105
R15718 GNDA.n1974 GNDA.n975 3.4105
R15719 GNDA.n1020 GNDA.n975 3.4105
R15720 GNDA.n1976 GNDA.n975 3.4105
R15721 GNDA.n1019 GNDA.n975 3.4105
R15722 GNDA.n1978 GNDA.n975 3.4105
R15723 GNDA.n1018 GNDA.n975 3.4105
R15724 GNDA.n1980 GNDA.n975 3.4105
R15725 GNDA.n1017 GNDA.n975 3.4105
R15726 GNDA.n1982 GNDA.n975 3.4105
R15727 GNDA.n1016 GNDA.n975 3.4105
R15728 GNDA.n1984 GNDA.n975 3.4105
R15729 GNDA.n1015 GNDA.n975 3.4105
R15730 GNDA.n1986 GNDA.n975 3.4105
R15731 GNDA.n1014 GNDA.n975 3.4105
R15732 GNDA.n1988 GNDA.n975 3.4105
R15733 GNDA.n1013 GNDA.n975 3.4105
R15734 GNDA.n1990 GNDA.n975 3.4105
R15735 GNDA.n1991 GNDA.n975 3.4105
R15736 GNDA.n2011 GNDA.n975 3.4105
R15737 GNDA.n2013 GNDA.n985 3.4105
R15738 GNDA.n1027 GNDA.n985 3.4105
R15739 GNDA.n1962 GNDA.n985 3.4105
R15740 GNDA.n1026 GNDA.n985 3.4105
R15741 GNDA.n1964 GNDA.n985 3.4105
R15742 GNDA.n1025 GNDA.n985 3.4105
R15743 GNDA.n1966 GNDA.n985 3.4105
R15744 GNDA.n1024 GNDA.n985 3.4105
R15745 GNDA.n1968 GNDA.n985 3.4105
R15746 GNDA.n1023 GNDA.n985 3.4105
R15747 GNDA.n1970 GNDA.n985 3.4105
R15748 GNDA.n1022 GNDA.n985 3.4105
R15749 GNDA.n1972 GNDA.n985 3.4105
R15750 GNDA.n1021 GNDA.n985 3.4105
R15751 GNDA.n1974 GNDA.n985 3.4105
R15752 GNDA.n1020 GNDA.n985 3.4105
R15753 GNDA.n1976 GNDA.n985 3.4105
R15754 GNDA.n1019 GNDA.n985 3.4105
R15755 GNDA.n1978 GNDA.n985 3.4105
R15756 GNDA.n1018 GNDA.n985 3.4105
R15757 GNDA.n1980 GNDA.n985 3.4105
R15758 GNDA.n1017 GNDA.n985 3.4105
R15759 GNDA.n1982 GNDA.n985 3.4105
R15760 GNDA.n1016 GNDA.n985 3.4105
R15761 GNDA.n1984 GNDA.n985 3.4105
R15762 GNDA.n1015 GNDA.n985 3.4105
R15763 GNDA.n1986 GNDA.n985 3.4105
R15764 GNDA.n1014 GNDA.n985 3.4105
R15765 GNDA.n1988 GNDA.n985 3.4105
R15766 GNDA.n1013 GNDA.n985 3.4105
R15767 GNDA.n1990 GNDA.n985 3.4105
R15768 GNDA.n1991 GNDA.n985 3.4105
R15769 GNDA.n2011 GNDA.n985 3.4105
R15770 GNDA.n2013 GNDA.n974 3.4105
R15771 GNDA.n1027 GNDA.n974 3.4105
R15772 GNDA.n1962 GNDA.n974 3.4105
R15773 GNDA.n1026 GNDA.n974 3.4105
R15774 GNDA.n1964 GNDA.n974 3.4105
R15775 GNDA.n1025 GNDA.n974 3.4105
R15776 GNDA.n1966 GNDA.n974 3.4105
R15777 GNDA.n1024 GNDA.n974 3.4105
R15778 GNDA.n1968 GNDA.n974 3.4105
R15779 GNDA.n1023 GNDA.n974 3.4105
R15780 GNDA.n1970 GNDA.n974 3.4105
R15781 GNDA.n1022 GNDA.n974 3.4105
R15782 GNDA.n1972 GNDA.n974 3.4105
R15783 GNDA.n1021 GNDA.n974 3.4105
R15784 GNDA.n1974 GNDA.n974 3.4105
R15785 GNDA.n1020 GNDA.n974 3.4105
R15786 GNDA.n1976 GNDA.n974 3.4105
R15787 GNDA.n1019 GNDA.n974 3.4105
R15788 GNDA.n1978 GNDA.n974 3.4105
R15789 GNDA.n1018 GNDA.n974 3.4105
R15790 GNDA.n1980 GNDA.n974 3.4105
R15791 GNDA.n1017 GNDA.n974 3.4105
R15792 GNDA.n1982 GNDA.n974 3.4105
R15793 GNDA.n1016 GNDA.n974 3.4105
R15794 GNDA.n1984 GNDA.n974 3.4105
R15795 GNDA.n1015 GNDA.n974 3.4105
R15796 GNDA.n1986 GNDA.n974 3.4105
R15797 GNDA.n1014 GNDA.n974 3.4105
R15798 GNDA.n1988 GNDA.n974 3.4105
R15799 GNDA.n1013 GNDA.n974 3.4105
R15800 GNDA.n1990 GNDA.n974 3.4105
R15801 GNDA.n1991 GNDA.n974 3.4105
R15802 GNDA.n2011 GNDA.n974 3.4105
R15803 GNDA.n2013 GNDA.n986 3.4105
R15804 GNDA.n1027 GNDA.n986 3.4105
R15805 GNDA.n1962 GNDA.n986 3.4105
R15806 GNDA.n1026 GNDA.n986 3.4105
R15807 GNDA.n1964 GNDA.n986 3.4105
R15808 GNDA.n1025 GNDA.n986 3.4105
R15809 GNDA.n1966 GNDA.n986 3.4105
R15810 GNDA.n1024 GNDA.n986 3.4105
R15811 GNDA.n1968 GNDA.n986 3.4105
R15812 GNDA.n1023 GNDA.n986 3.4105
R15813 GNDA.n1970 GNDA.n986 3.4105
R15814 GNDA.n1022 GNDA.n986 3.4105
R15815 GNDA.n1972 GNDA.n986 3.4105
R15816 GNDA.n1021 GNDA.n986 3.4105
R15817 GNDA.n1974 GNDA.n986 3.4105
R15818 GNDA.n1020 GNDA.n986 3.4105
R15819 GNDA.n1976 GNDA.n986 3.4105
R15820 GNDA.n1019 GNDA.n986 3.4105
R15821 GNDA.n1978 GNDA.n986 3.4105
R15822 GNDA.n1018 GNDA.n986 3.4105
R15823 GNDA.n1980 GNDA.n986 3.4105
R15824 GNDA.n1017 GNDA.n986 3.4105
R15825 GNDA.n1982 GNDA.n986 3.4105
R15826 GNDA.n1016 GNDA.n986 3.4105
R15827 GNDA.n1984 GNDA.n986 3.4105
R15828 GNDA.n1015 GNDA.n986 3.4105
R15829 GNDA.n1986 GNDA.n986 3.4105
R15830 GNDA.n1014 GNDA.n986 3.4105
R15831 GNDA.n1988 GNDA.n986 3.4105
R15832 GNDA.n1013 GNDA.n986 3.4105
R15833 GNDA.n1990 GNDA.n986 3.4105
R15834 GNDA.n1991 GNDA.n986 3.4105
R15835 GNDA.n2011 GNDA.n986 3.4105
R15836 GNDA.n2013 GNDA.n973 3.4105
R15837 GNDA.n1027 GNDA.n973 3.4105
R15838 GNDA.n1962 GNDA.n973 3.4105
R15839 GNDA.n1026 GNDA.n973 3.4105
R15840 GNDA.n1964 GNDA.n973 3.4105
R15841 GNDA.n1025 GNDA.n973 3.4105
R15842 GNDA.n1966 GNDA.n973 3.4105
R15843 GNDA.n1024 GNDA.n973 3.4105
R15844 GNDA.n1968 GNDA.n973 3.4105
R15845 GNDA.n1023 GNDA.n973 3.4105
R15846 GNDA.n1970 GNDA.n973 3.4105
R15847 GNDA.n1022 GNDA.n973 3.4105
R15848 GNDA.n1972 GNDA.n973 3.4105
R15849 GNDA.n1021 GNDA.n973 3.4105
R15850 GNDA.n1974 GNDA.n973 3.4105
R15851 GNDA.n1020 GNDA.n973 3.4105
R15852 GNDA.n1976 GNDA.n973 3.4105
R15853 GNDA.n1019 GNDA.n973 3.4105
R15854 GNDA.n1978 GNDA.n973 3.4105
R15855 GNDA.n1018 GNDA.n973 3.4105
R15856 GNDA.n1980 GNDA.n973 3.4105
R15857 GNDA.n1017 GNDA.n973 3.4105
R15858 GNDA.n1982 GNDA.n973 3.4105
R15859 GNDA.n1016 GNDA.n973 3.4105
R15860 GNDA.n1984 GNDA.n973 3.4105
R15861 GNDA.n1015 GNDA.n973 3.4105
R15862 GNDA.n1986 GNDA.n973 3.4105
R15863 GNDA.n1014 GNDA.n973 3.4105
R15864 GNDA.n1988 GNDA.n973 3.4105
R15865 GNDA.n1013 GNDA.n973 3.4105
R15866 GNDA.n1990 GNDA.n973 3.4105
R15867 GNDA.n1991 GNDA.n973 3.4105
R15868 GNDA.n2011 GNDA.n973 3.4105
R15869 GNDA.n2013 GNDA.n987 3.4105
R15870 GNDA.n1027 GNDA.n987 3.4105
R15871 GNDA.n1962 GNDA.n987 3.4105
R15872 GNDA.n1026 GNDA.n987 3.4105
R15873 GNDA.n1964 GNDA.n987 3.4105
R15874 GNDA.n1025 GNDA.n987 3.4105
R15875 GNDA.n1966 GNDA.n987 3.4105
R15876 GNDA.n1024 GNDA.n987 3.4105
R15877 GNDA.n1968 GNDA.n987 3.4105
R15878 GNDA.n1023 GNDA.n987 3.4105
R15879 GNDA.n1970 GNDA.n987 3.4105
R15880 GNDA.n1022 GNDA.n987 3.4105
R15881 GNDA.n1972 GNDA.n987 3.4105
R15882 GNDA.n1021 GNDA.n987 3.4105
R15883 GNDA.n1974 GNDA.n987 3.4105
R15884 GNDA.n1020 GNDA.n987 3.4105
R15885 GNDA.n1976 GNDA.n987 3.4105
R15886 GNDA.n1019 GNDA.n987 3.4105
R15887 GNDA.n1978 GNDA.n987 3.4105
R15888 GNDA.n1018 GNDA.n987 3.4105
R15889 GNDA.n1980 GNDA.n987 3.4105
R15890 GNDA.n1017 GNDA.n987 3.4105
R15891 GNDA.n1982 GNDA.n987 3.4105
R15892 GNDA.n1016 GNDA.n987 3.4105
R15893 GNDA.n1984 GNDA.n987 3.4105
R15894 GNDA.n1015 GNDA.n987 3.4105
R15895 GNDA.n1986 GNDA.n987 3.4105
R15896 GNDA.n1014 GNDA.n987 3.4105
R15897 GNDA.n1988 GNDA.n987 3.4105
R15898 GNDA.n1013 GNDA.n987 3.4105
R15899 GNDA.n1990 GNDA.n987 3.4105
R15900 GNDA.n1991 GNDA.n987 3.4105
R15901 GNDA.n2011 GNDA.n987 3.4105
R15902 GNDA.n2013 GNDA.n972 3.4105
R15903 GNDA.n1027 GNDA.n972 3.4105
R15904 GNDA.n1962 GNDA.n972 3.4105
R15905 GNDA.n1026 GNDA.n972 3.4105
R15906 GNDA.n1964 GNDA.n972 3.4105
R15907 GNDA.n1025 GNDA.n972 3.4105
R15908 GNDA.n1966 GNDA.n972 3.4105
R15909 GNDA.n1024 GNDA.n972 3.4105
R15910 GNDA.n1968 GNDA.n972 3.4105
R15911 GNDA.n1023 GNDA.n972 3.4105
R15912 GNDA.n1970 GNDA.n972 3.4105
R15913 GNDA.n1022 GNDA.n972 3.4105
R15914 GNDA.n1972 GNDA.n972 3.4105
R15915 GNDA.n1021 GNDA.n972 3.4105
R15916 GNDA.n1974 GNDA.n972 3.4105
R15917 GNDA.n1020 GNDA.n972 3.4105
R15918 GNDA.n1976 GNDA.n972 3.4105
R15919 GNDA.n1019 GNDA.n972 3.4105
R15920 GNDA.n1978 GNDA.n972 3.4105
R15921 GNDA.n1018 GNDA.n972 3.4105
R15922 GNDA.n1980 GNDA.n972 3.4105
R15923 GNDA.n1017 GNDA.n972 3.4105
R15924 GNDA.n1982 GNDA.n972 3.4105
R15925 GNDA.n1016 GNDA.n972 3.4105
R15926 GNDA.n1984 GNDA.n972 3.4105
R15927 GNDA.n1015 GNDA.n972 3.4105
R15928 GNDA.n1986 GNDA.n972 3.4105
R15929 GNDA.n1014 GNDA.n972 3.4105
R15930 GNDA.n1988 GNDA.n972 3.4105
R15931 GNDA.n1013 GNDA.n972 3.4105
R15932 GNDA.n1990 GNDA.n972 3.4105
R15933 GNDA.n1991 GNDA.n972 3.4105
R15934 GNDA.n2011 GNDA.n972 3.4105
R15935 GNDA.n2013 GNDA.n988 3.4105
R15936 GNDA.n1027 GNDA.n988 3.4105
R15937 GNDA.n1962 GNDA.n988 3.4105
R15938 GNDA.n1026 GNDA.n988 3.4105
R15939 GNDA.n1964 GNDA.n988 3.4105
R15940 GNDA.n1025 GNDA.n988 3.4105
R15941 GNDA.n1966 GNDA.n988 3.4105
R15942 GNDA.n1024 GNDA.n988 3.4105
R15943 GNDA.n1968 GNDA.n988 3.4105
R15944 GNDA.n1023 GNDA.n988 3.4105
R15945 GNDA.n1970 GNDA.n988 3.4105
R15946 GNDA.n1022 GNDA.n988 3.4105
R15947 GNDA.n1972 GNDA.n988 3.4105
R15948 GNDA.n1021 GNDA.n988 3.4105
R15949 GNDA.n1974 GNDA.n988 3.4105
R15950 GNDA.n1020 GNDA.n988 3.4105
R15951 GNDA.n1976 GNDA.n988 3.4105
R15952 GNDA.n1019 GNDA.n988 3.4105
R15953 GNDA.n1978 GNDA.n988 3.4105
R15954 GNDA.n1018 GNDA.n988 3.4105
R15955 GNDA.n1980 GNDA.n988 3.4105
R15956 GNDA.n1017 GNDA.n988 3.4105
R15957 GNDA.n1982 GNDA.n988 3.4105
R15958 GNDA.n1016 GNDA.n988 3.4105
R15959 GNDA.n1984 GNDA.n988 3.4105
R15960 GNDA.n1015 GNDA.n988 3.4105
R15961 GNDA.n1986 GNDA.n988 3.4105
R15962 GNDA.n1014 GNDA.n988 3.4105
R15963 GNDA.n1988 GNDA.n988 3.4105
R15964 GNDA.n1013 GNDA.n988 3.4105
R15965 GNDA.n1990 GNDA.n988 3.4105
R15966 GNDA.n1991 GNDA.n988 3.4105
R15967 GNDA.n2011 GNDA.n988 3.4105
R15968 GNDA.n2013 GNDA.n971 3.4105
R15969 GNDA.n1027 GNDA.n971 3.4105
R15970 GNDA.n1962 GNDA.n971 3.4105
R15971 GNDA.n1026 GNDA.n971 3.4105
R15972 GNDA.n1964 GNDA.n971 3.4105
R15973 GNDA.n1025 GNDA.n971 3.4105
R15974 GNDA.n1966 GNDA.n971 3.4105
R15975 GNDA.n1024 GNDA.n971 3.4105
R15976 GNDA.n1968 GNDA.n971 3.4105
R15977 GNDA.n1023 GNDA.n971 3.4105
R15978 GNDA.n1970 GNDA.n971 3.4105
R15979 GNDA.n1022 GNDA.n971 3.4105
R15980 GNDA.n1972 GNDA.n971 3.4105
R15981 GNDA.n1021 GNDA.n971 3.4105
R15982 GNDA.n1974 GNDA.n971 3.4105
R15983 GNDA.n1020 GNDA.n971 3.4105
R15984 GNDA.n1976 GNDA.n971 3.4105
R15985 GNDA.n1019 GNDA.n971 3.4105
R15986 GNDA.n1978 GNDA.n971 3.4105
R15987 GNDA.n1018 GNDA.n971 3.4105
R15988 GNDA.n1980 GNDA.n971 3.4105
R15989 GNDA.n1017 GNDA.n971 3.4105
R15990 GNDA.n1982 GNDA.n971 3.4105
R15991 GNDA.n1016 GNDA.n971 3.4105
R15992 GNDA.n1984 GNDA.n971 3.4105
R15993 GNDA.n1015 GNDA.n971 3.4105
R15994 GNDA.n1986 GNDA.n971 3.4105
R15995 GNDA.n1014 GNDA.n971 3.4105
R15996 GNDA.n1988 GNDA.n971 3.4105
R15997 GNDA.n1013 GNDA.n971 3.4105
R15998 GNDA.n1990 GNDA.n971 3.4105
R15999 GNDA.n1991 GNDA.n971 3.4105
R16000 GNDA.n2011 GNDA.n971 3.4105
R16001 GNDA.n2013 GNDA.n989 3.4105
R16002 GNDA.n1027 GNDA.n989 3.4105
R16003 GNDA.n1962 GNDA.n989 3.4105
R16004 GNDA.n1026 GNDA.n989 3.4105
R16005 GNDA.n1964 GNDA.n989 3.4105
R16006 GNDA.n1025 GNDA.n989 3.4105
R16007 GNDA.n1966 GNDA.n989 3.4105
R16008 GNDA.n1024 GNDA.n989 3.4105
R16009 GNDA.n1968 GNDA.n989 3.4105
R16010 GNDA.n1023 GNDA.n989 3.4105
R16011 GNDA.n1970 GNDA.n989 3.4105
R16012 GNDA.n1022 GNDA.n989 3.4105
R16013 GNDA.n1972 GNDA.n989 3.4105
R16014 GNDA.n1021 GNDA.n989 3.4105
R16015 GNDA.n1974 GNDA.n989 3.4105
R16016 GNDA.n1020 GNDA.n989 3.4105
R16017 GNDA.n1976 GNDA.n989 3.4105
R16018 GNDA.n1019 GNDA.n989 3.4105
R16019 GNDA.n1978 GNDA.n989 3.4105
R16020 GNDA.n1018 GNDA.n989 3.4105
R16021 GNDA.n1980 GNDA.n989 3.4105
R16022 GNDA.n1017 GNDA.n989 3.4105
R16023 GNDA.n1982 GNDA.n989 3.4105
R16024 GNDA.n1016 GNDA.n989 3.4105
R16025 GNDA.n1984 GNDA.n989 3.4105
R16026 GNDA.n1015 GNDA.n989 3.4105
R16027 GNDA.n1986 GNDA.n989 3.4105
R16028 GNDA.n1014 GNDA.n989 3.4105
R16029 GNDA.n1988 GNDA.n989 3.4105
R16030 GNDA.n1013 GNDA.n989 3.4105
R16031 GNDA.n1990 GNDA.n989 3.4105
R16032 GNDA.n1991 GNDA.n989 3.4105
R16033 GNDA.n2011 GNDA.n989 3.4105
R16034 GNDA.n2013 GNDA.n970 3.4105
R16035 GNDA.n1027 GNDA.n970 3.4105
R16036 GNDA.n1962 GNDA.n970 3.4105
R16037 GNDA.n1026 GNDA.n970 3.4105
R16038 GNDA.n1964 GNDA.n970 3.4105
R16039 GNDA.n1025 GNDA.n970 3.4105
R16040 GNDA.n1966 GNDA.n970 3.4105
R16041 GNDA.n1024 GNDA.n970 3.4105
R16042 GNDA.n1968 GNDA.n970 3.4105
R16043 GNDA.n1023 GNDA.n970 3.4105
R16044 GNDA.n1970 GNDA.n970 3.4105
R16045 GNDA.n1022 GNDA.n970 3.4105
R16046 GNDA.n1972 GNDA.n970 3.4105
R16047 GNDA.n1021 GNDA.n970 3.4105
R16048 GNDA.n1974 GNDA.n970 3.4105
R16049 GNDA.n1020 GNDA.n970 3.4105
R16050 GNDA.n1976 GNDA.n970 3.4105
R16051 GNDA.n1019 GNDA.n970 3.4105
R16052 GNDA.n1978 GNDA.n970 3.4105
R16053 GNDA.n1018 GNDA.n970 3.4105
R16054 GNDA.n1980 GNDA.n970 3.4105
R16055 GNDA.n1017 GNDA.n970 3.4105
R16056 GNDA.n1982 GNDA.n970 3.4105
R16057 GNDA.n1016 GNDA.n970 3.4105
R16058 GNDA.n1984 GNDA.n970 3.4105
R16059 GNDA.n1015 GNDA.n970 3.4105
R16060 GNDA.n1986 GNDA.n970 3.4105
R16061 GNDA.n1014 GNDA.n970 3.4105
R16062 GNDA.n1988 GNDA.n970 3.4105
R16063 GNDA.n1013 GNDA.n970 3.4105
R16064 GNDA.n1990 GNDA.n970 3.4105
R16065 GNDA.n1991 GNDA.n970 3.4105
R16066 GNDA.n2011 GNDA.n970 3.4105
R16067 GNDA.n2013 GNDA.n990 3.4105
R16068 GNDA.n1027 GNDA.n990 3.4105
R16069 GNDA.n1962 GNDA.n990 3.4105
R16070 GNDA.n1026 GNDA.n990 3.4105
R16071 GNDA.n1964 GNDA.n990 3.4105
R16072 GNDA.n1025 GNDA.n990 3.4105
R16073 GNDA.n1966 GNDA.n990 3.4105
R16074 GNDA.n1024 GNDA.n990 3.4105
R16075 GNDA.n1968 GNDA.n990 3.4105
R16076 GNDA.n1023 GNDA.n990 3.4105
R16077 GNDA.n1970 GNDA.n990 3.4105
R16078 GNDA.n1022 GNDA.n990 3.4105
R16079 GNDA.n1972 GNDA.n990 3.4105
R16080 GNDA.n1021 GNDA.n990 3.4105
R16081 GNDA.n1974 GNDA.n990 3.4105
R16082 GNDA.n1020 GNDA.n990 3.4105
R16083 GNDA.n1976 GNDA.n990 3.4105
R16084 GNDA.n1019 GNDA.n990 3.4105
R16085 GNDA.n1978 GNDA.n990 3.4105
R16086 GNDA.n1018 GNDA.n990 3.4105
R16087 GNDA.n1980 GNDA.n990 3.4105
R16088 GNDA.n1017 GNDA.n990 3.4105
R16089 GNDA.n1982 GNDA.n990 3.4105
R16090 GNDA.n1016 GNDA.n990 3.4105
R16091 GNDA.n1984 GNDA.n990 3.4105
R16092 GNDA.n1015 GNDA.n990 3.4105
R16093 GNDA.n1986 GNDA.n990 3.4105
R16094 GNDA.n1014 GNDA.n990 3.4105
R16095 GNDA.n1988 GNDA.n990 3.4105
R16096 GNDA.n1013 GNDA.n990 3.4105
R16097 GNDA.n1990 GNDA.n990 3.4105
R16098 GNDA.n1991 GNDA.n990 3.4105
R16099 GNDA.n2011 GNDA.n990 3.4105
R16100 GNDA.n2013 GNDA.n969 3.4105
R16101 GNDA.n1027 GNDA.n969 3.4105
R16102 GNDA.n1962 GNDA.n969 3.4105
R16103 GNDA.n1026 GNDA.n969 3.4105
R16104 GNDA.n1964 GNDA.n969 3.4105
R16105 GNDA.n1025 GNDA.n969 3.4105
R16106 GNDA.n1966 GNDA.n969 3.4105
R16107 GNDA.n1024 GNDA.n969 3.4105
R16108 GNDA.n1968 GNDA.n969 3.4105
R16109 GNDA.n1023 GNDA.n969 3.4105
R16110 GNDA.n1970 GNDA.n969 3.4105
R16111 GNDA.n1022 GNDA.n969 3.4105
R16112 GNDA.n1972 GNDA.n969 3.4105
R16113 GNDA.n1021 GNDA.n969 3.4105
R16114 GNDA.n1974 GNDA.n969 3.4105
R16115 GNDA.n1020 GNDA.n969 3.4105
R16116 GNDA.n1976 GNDA.n969 3.4105
R16117 GNDA.n1019 GNDA.n969 3.4105
R16118 GNDA.n1978 GNDA.n969 3.4105
R16119 GNDA.n1018 GNDA.n969 3.4105
R16120 GNDA.n1980 GNDA.n969 3.4105
R16121 GNDA.n1017 GNDA.n969 3.4105
R16122 GNDA.n1982 GNDA.n969 3.4105
R16123 GNDA.n1016 GNDA.n969 3.4105
R16124 GNDA.n1984 GNDA.n969 3.4105
R16125 GNDA.n1015 GNDA.n969 3.4105
R16126 GNDA.n1986 GNDA.n969 3.4105
R16127 GNDA.n1014 GNDA.n969 3.4105
R16128 GNDA.n1988 GNDA.n969 3.4105
R16129 GNDA.n1013 GNDA.n969 3.4105
R16130 GNDA.n1990 GNDA.n969 3.4105
R16131 GNDA.n1991 GNDA.n969 3.4105
R16132 GNDA.n2011 GNDA.n969 3.4105
R16133 GNDA.n2013 GNDA.n991 3.4105
R16134 GNDA.n1027 GNDA.n991 3.4105
R16135 GNDA.n1962 GNDA.n991 3.4105
R16136 GNDA.n1026 GNDA.n991 3.4105
R16137 GNDA.n1964 GNDA.n991 3.4105
R16138 GNDA.n1025 GNDA.n991 3.4105
R16139 GNDA.n1966 GNDA.n991 3.4105
R16140 GNDA.n1024 GNDA.n991 3.4105
R16141 GNDA.n1968 GNDA.n991 3.4105
R16142 GNDA.n1023 GNDA.n991 3.4105
R16143 GNDA.n1970 GNDA.n991 3.4105
R16144 GNDA.n1022 GNDA.n991 3.4105
R16145 GNDA.n1972 GNDA.n991 3.4105
R16146 GNDA.n1021 GNDA.n991 3.4105
R16147 GNDA.n1974 GNDA.n991 3.4105
R16148 GNDA.n1020 GNDA.n991 3.4105
R16149 GNDA.n1976 GNDA.n991 3.4105
R16150 GNDA.n1019 GNDA.n991 3.4105
R16151 GNDA.n1978 GNDA.n991 3.4105
R16152 GNDA.n1018 GNDA.n991 3.4105
R16153 GNDA.n1980 GNDA.n991 3.4105
R16154 GNDA.n1017 GNDA.n991 3.4105
R16155 GNDA.n1982 GNDA.n991 3.4105
R16156 GNDA.n1016 GNDA.n991 3.4105
R16157 GNDA.n1984 GNDA.n991 3.4105
R16158 GNDA.n1015 GNDA.n991 3.4105
R16159 GNDA.n1986 GNDA.n991 3.4105
R16160 GNDA.n1014 GNDA.n991 3.4105
R16161 GNDA.n1988 GNDA.n991 3.4105
R16162 GNDA.n1013 GNDA.n991 3.4105
R16163 GNDA.n1990 GNDA.n991 3.4105
R16164 GNDA.n1991 GNDA.n991 3.4105
R16165 GNDA.n2011 GNDA.n991 3.4105
R16166 GNDA.n2013 GNDA.n968 3.4105
R16167 GNDA.n1027 GNDA.n968 3.4105
R16168 GNDA.n1962 GNDA.n968 3.4105
R16169 GNDA.n1026 GNDA.n968 3.4105
R16170 GNDA.n1964 GNDA.n968 3.4105
R16171 GNDA.n1025 GNDA.n968 3.4105
R16172 GNDA.n1966 GNDA.n968 3.4105
R16173 GNDA.n1024 GNDA.n968 3.4105
R16174 GNDA.n1968 GNDA.n968 3.4105
R16175 GNDA.n1023 GNDA.n968 3.4105
R16176 GNDA.n1970 GNDA.n968 3.4105
R16177 GNDA.n1022 GNDA.n968 3.4105
R16178 GNDA.n1972 GNDA.n968 3.4105
R16179 GNDA.n1021 GNDA.n968 3.4105
R16180 GNDA.n1974 GNDA.n968 3.4105
R16181 GNDA.n1020 GNDA.n968 3.4105
R16182 GNDA.n1976 GNDA.n968 3.4105
R16183 GNDA.n1019 GNDA.n968 3.4105
R16184 GNDA.n1978 GNDA.n968 3.4105
R16185 GNDA.n1018 GNDA.n968 3.4105
R16186 GNDA.n1980 GNDA.n968 3.4105
R16187 GNDA.n1017 GNDA.n968 3.4105
R16188 GNDA.n1982 GNDA.n968 3.4105
R16189 GNDA.n1016 GNDA.n968 3.4105
R16190 GNDA.n1984 GNDA.n968 3.4105
R16191 GNDA.n1015 GNDA.n968 3.4105
R16192 GNDA.n1986 GNDA.n968 3.4105
R16193 GNDA.n1014 GNDA.n968 3.4105
R16194 GNDA.n1988 GNDA.n968 3.4105
R16195 GNDA.n1013 GNDA.n968 3.4105
R16196 GNDA.n1990 GNDA.n968 3.4105
R16197 GNDA.n1991 GNDA.n968 3.4105
R16198 GNDA.n2011 GNDA.n968 3.4105
R16199 GNDA.n2013 GNDA.n992 3.4105
R16200 GNDA.n1027 GNDA.n992 3.4105
R16201 GNDA.n1962 GNDA.n992 3.4105
R16202 GNDA.n1026 GNDA.n992 3.4105
R16203 GNDA.n1964 GNDA.n992 3.4105
R16204 GNDA.n1025 GNDA.n992 3.4105
R16205 GNDA.n1966 GNDA.n992 3.4105
R16206 GNDA.n1024 GNDA.n992 3.4105
R16207 GNDA.n1968 GNDA.n992 3.4105
R16208 GNDA.n1023 GNDA.n992 3.4105
R16209 GNDA.n1970 GNDA.n992 3.4105
R16210 GNDA.n1022 GNDA.n992 3.4105
R16211 GNDA.n1972 GNDA.n992 3.4105
R16212 GNDA.n1021 GNDA.n992 3.4105
R16213 GNDA.n1974 GNDA.n992 3.4105
R16214 GNDA.n1020 GNDA.n992 3.4105
R16215 GNDA.n1976 GNDA.n992 3.4105
R16216 GNDA.n1019 GNDA.n992 3.4105
R16217 GNDA.n1978 GNDA.n992 3.4105
R16218 GNDA.n1018 GNDA.n992 3.4105
R16219 GNDA.n1980 GNDA.n992 3.4105
R16220 GNDA.n1017 GNDA.n992 3.4105
R16221 GNDA.n1982 GNDA.n992 3.4105
R16222 GNDA.n1016 GNDA.n992 3.4105
R16223 GNDA.n1984 GNDA.n992 3.4105
R16224 GNDA.n1015 GNDA.n992 3.4105
R16225 GNDA.n1986 GNDA.n992 3.4105
R16226 GNDA.n1014 GNDA.n992 3.4105
R16227 GNDA.n1988 GNDA.n992 3.4105
R16228 GNDA.n1013 GNDA.n992 3.4105
R16229 GNDA.n1990 GNDA.n992 3.4105
R16230 GNDA.n1991 GNDA.n992 3.4105
R16231 GNDA.n2011 GNDA.n992 3.4105
R16232 GNDA.n2013 GNDA.n967 3.4105
R16233 GNDA.n1027 GNDA.n967 3.4105
R16234 GNDA.n1962 GNDA.n967 3.4105
R16235 GNDA.n1026 GNDA.n967 3.4105
R16236 GNDA.n1964 GNDA.n967 3.4105
R16237 GNDA.n1025 GNDA.n967 3.4105
R16238 GNDA.n1966 GNDA.n967 3.4105
R16239 GNDA.n1024 GNDA.n967 3.4105
R16240 GNDA.n1968 GNDA.n967 3.4105
R16241 GNDA.n1023 GNDA.n967 3.4105
R16242 GNDA.n1970 GNDA.n967 3.4105
R16243 GNDA.n1022 GNDA.n967 3.4105
R16244 GNDA.n1972 GNDA.n967 3.4105
R16245 GNDA.n1021 GNDA.n967 3.4105
R16246 GNDA.n1974 GNDA.n967 3.4105
R16247 GNDA.n1020 GNDA.n967 3.4105
R16248 GNDA.n1976 GNDA.n967 3.4105
R16249 GNDA.n1019 GNDA.n967 3.4105
R16250 GNDA.n1978 GNDA.n967 3.4105
R16251 GNDA.n1018 GNDA.n967 3.4105
R16252 GNDA.n1980 GNDA.n967 3.4105
R16253 GNDA.n1017 GNDA.n967 3.4105
R16254 GNDA.n1982 GNDA.n967 3.4105
R16255 GNDA.n1016 GNDA.n967 3.4105
R16256 GNDA.n1984 GNDA.n967 3.4105
R16257 GNDA.n1015 GNDA.n967 3.4105
R16258 GNDA.n1986 GNDA.n967 3.4105
R16259 GNDA.n1014 GNDA.n967 3.4105
R16260 GNDA.n1988 GNDA.n967 3.4105
R16261 GNDA.n1013 GNDA.n967 3.4105
R16262 GNDA.n1990 GNDA.n967 3.4105
R16263 GNDA.n1991 GNDA.n967 3.4105
R16264 GNDA.n2011 GNDA.n967 3.4105
R16265 GNDA.n2013 GNDA.n993 3.4105
R16266 GNDA.n1027 GNDA.n993 3.4105
R16267 GNDA.n1962 GNDA.n993 3.4105
R16268 GNDA.n1026 GNDA.n993 3.4105
R16269 GNDA.n1964 GNDA.n993 3.4105
R16270 GNDA.n1025 GNDA.n993 3.4105
R16271 GNDA.n1966 GNDA.n993 3.4105
R16272 GNDA.n1024 GNDA.n993 3.4105
R16273 GNDA.n1968 GNDA.n993 3.4105
R16274 GNDA.n1023 GNDA.n993 3.4105
R16275 GNDA.n1970 GNDA.n993 3.4105
R16276 GNDA.n1022 GNDA.n993 3.4105
R16277 GNDA.n1972 GNDA.n993 3.4105
R16278 GNDA.n1021 GNDA.n993 3.4105
R16279 GNDA.n1974 GNDA.n993 3.4105
R16280 GNDA.n1020 GNDA.n993 3.4105
R16281 GNDA.n1976 GNDA.n993 3.4105
R16282 GNDA.n1019 GNDA.n993 3.4105
R16283 GNDA.n1978 GNDA.n993 3.4105
R16284 GNDA.n1018 GNDA.n993 3.4105
R16285 GNDA.n1980 GNDA.n993 3.4105
R16286 GNDA.n1017 GNDA.n993 3.4105
R16287 GNDA.n1982 GNDA.n993 3.4105
R16288 GNDA.n1016 GNDA.n993 3.4105
R16289 GNDA.n1984 GNDA.n993 3.4105
R16290 GNDA.n1015 GNDA.n993 3.4105
R16291 GNDA.n1986 GNDA.n993 3.4105
R16292 GNDA.n1014 GNDA.n993 3.4105
R16293 GNDA.n1988 GNDA.n993 3.4105
R16294 GNDA.n1013 GNDA.n993 3.4105
R16295 GNDA.n1990 GNDA.n993 3.4105
R16296 GNDA.n1991 GNDA.n993 3.4105
R16297 GNDA.n2011 GNDA.n993 3.4105
R16298 GNDA.n2013 GNDA.n966 3.4105
R16299 GNDA.n1027 GNDA.n966 3.4105
R16300 GNDA.n1962 GNDA.n966 3.4105
R16301 GNDA.n1026 GNDA.n966 3.4105
R16302 GNDA.n1964 GNDA.n966 3.4105
R16303 GNDA.n1025 GNDA.n966 3.4105
R16304 GNDA.n1966 GNDA.n966 3.4105
R16305 GNDA.n1024 GNDA.n966 3.4105
R16306 GNDA.n1968 GNDA.n966 3.4105
R16307 GNDA.n1023 GNDA.n966 3.4105
R16308 GNDA.n1970 GNDA.n966 3.4105
R16309 GNDA.n1022 GNDA.n966 3.4105
R16310 GNDA.n1972 GNDA.n966 3.4105
R16311 GNDA.n1021 GNDA.n966 3.4105
R16312 GNDA.n1974 GNDA.n966 3.4105
R16313 GNDA.n1020 GNDA.n966 3.4105
R16314 GNDA.n1976 GNDA.n966 3.4105
R16315 GNDA.n1019 GNDA.n966 3.4105
R16316 GNDA.n1978 GNDA.n966 3.4105
R16317 GNDA.n1018 GNDA.n966 3.4105
R16318 GNDA.n1980 GNDA.n966 3.4105
R16319 GNDA.n1017 GNDA.n966 3.4105
R16320 GNDA.n1982 GNDA.n966 3.4105
R16321 GNDA.n1016 GNDA.n966 3.4105
R16322 GNDA.n1984 GNDA.n966 3.4105
R16323 GNDA.n1015 GNDA.n966 3.4105
R16324 GNDA.n1986 GNDA.n966 3.4105
R16325 GNDA.n1014 GNDA.n966 3.4105
R16326 GNDA.n1988 GNDA.n966 3.4105
R16327 GNDA.n1013 GNDA.n966 3.4105
R16328 GNDA.n1990 GNDA.n966 3.4105
R16329 GNDA.n1991 GNDA.n966 3.4105
R16330 GNDA.n2011 GNDA.n966 3.4105
R16331 GNDA.n2013 GNDA.n994 3.4105
R16332 GNDA.n1027 GNDA.n994 3.4105
R16333 GNDA.n1962 GNDA.n994 3.4105
R16334 GNDA.n1026 GNDA.n994 3.4105
R16335 GNDA.n1964 GNDA.n994 3.4105
R16336 GNDA.n1025 GNDA.n994 3.4105
R16337 GNDA.n1966 GNDA.n994 3.4105
R16338 GNDA.n1024 GNDA.n994 3.4105
R16339 GNDA.n1968 GNDA.n994 3.4105
R16340 GNDA.n1023 GNDA.n994 3.4105
R16341 GNDA.n1970 GNDA.n994 3.4105
R16342 GNDA.n1022 GNDA.n994 3.4105
R16343 GNDA.n1972 GNDA.n994 3.4105
R16344 GNDA.n1021 GNDA.n994 3.4105
R16345 GNDA.n1974 GNDA.n994 3.4105
R16346 GNDA.n1020 GNDA.n994 3.4105
R16347 GNDA.n1976 GNDA.n994 3.4105
R16348 GNDA.n1019 GNDA.n994 3.4105
R16349 GNDA.n1978 GNDA.n994 3.4105
R16350 GNDA.n1018 GNDA.n994 3.4105
R16351 GNDA.n1980 GNDA.n994 3.4105
R16352 GNDA.n1017 GNDA.n994 3.4105
R16353 GNDA.n1982 GNDA.n994 3.4105
R16354 GNDA.n1016 GNDA.n994 3.4105
R16355 GNDA.n1984 GNDA.n994 3.4105
R16356 GNDA.n1015 GNDA.n994 3.4105
R16357 GNDA.n1986 GNDA.n994 3.4105
R16358 GNDA.n1014 GNDA.n994 3.4105
R16359 GNDA.n1988 GNDA.n994 3.4105
R16360 GNDA.n1013 GNDA.n994 3.4105
R16361 GNDA.n1990 GNDA.n994 3.4105
R16362 GNDA.n1991 GNDA.n994 3.4105
R16363 GNDA.n2011 GNDA.n994 3.4105
R16364 GNDA.n2013 GNDA.n965 3.4105
R16365 GNDA.n1027 GNDA.n965 3.4105
R16366 GNDA.n1962 GNDA.n965 3.4105
R16367 GNDA.n1026 GNDA.n965 3.4105
R16368 GNDA.n1964 GNDA.n965 3.4105
R16369 GNDA.n1025 GNDA.n965 3.4105
R16370 GNDA.n1966 GNDA.n965 3.4105
R16371 GNDA.n1024 GNDA.n965 3.4105
R16372 GNDA.n1968 GNDA.n965 3.4105
R16373 GNDA.n1023 GNDA.n965 3.4105
R16374 GNDA.n1970 GNDA.n965 3.4105
R16375 GNDA.n1022 GNDA.n965 3.4105
R16376 GNDA.n1972 GNDA.n965 3.4105
R16377 GNDA.n1021 GNDA.n965 3.4105
R16378 GNDA.n1974 GNDA.n965 3.4105
R16379 GNDA.n1020 GNDA.n965 3.4105
R16380 GNDA.n1976 GNDA.n965 3.4105
R16381 GNDA.n1019 GNDA.n965 3.4105
R16382 GNDA.n1978 GNDA.n965 3.4105
R16383 GNDA.n1018 GNDA.n965 3.4105
R16384 GNDA.n1980 GNDA.n965 3.4105
R16385 GNDA.n1017 GNDA.n965 3.4105
R16386 GNDA.n1982 GNDA.n965 3.4105
R16387 GNDA.n1016 GNDA.n965 3.4105
R16388 GNDA.n1984 GNDA.n965 3.4105
R16389 GNDA.n1015 GNDA.n965 3.4105
R16390 GNDA.n1986 GNDA.n965 3.4105
R16391 GNDA.n1014 GNDA.n965 3.4105
R16392 GNDA.n1988 GNDA.n965 3.4105
R16393 GNDA.n1013 GNDA.n965 3.4105
R16394 GNDA.n1990 GNDA.n965 3.4105
R16395 GNDA.n1991 GNDA.n965 3.4105
R16396 GNDA.n2011 GNDA.n965 3.4105
R16397 GNDA.n2013 GNDA.n995 3.4105
R16398 GNDA.n1027 GNDA.n995 3.4105
R16399 GNDA.n1962 GNDA.n995 3.4105
R16400 GNDA.n1026 GNDA.n995 3.4105
R16401 GNDA.n1964 GNDA.n995 3.4105
R16402 GNDA.n1025 GNDA.n995 3.4105
R16403 GNDA.n1966 GNDA.n995 3.4105
R16404 GNDA.n1024 GNDA.n995 3.4105
R16405 GNDA.n1968 GNDA.n995 3.4105
R16406 GNDA.n1023 GNDA.n995 3.4105
R16407 GNDA.n1970 GNDA.n995 3.4105
R16408 GNDA.n1022 GNDA.n995 3.4105
R16409 GNDA.n1972 GNDA.n995 3.4105
R16410 GNDA.n1021 GNDA.n995 3.4105
R16411 GNDA.n1974 GNDA.n995 3.4105
R16412 GNDA.n1020 GNDA.n995 3.4105
R16413 GNDA.n1976 GNDA.n995 3.4105
R16414 GNDA.n1019 GNDA.n995 3.4105
R16415 GNDA.n1978 GNDA.n995 3.4105
R16416 GNDA.n1018 GNDA.n995 3.4105
R16417 GNDA.n1980 GNDA.n995 3.4105
R16418 GNDA.n1017 GNDA.n995 3.4105
R16419 GNDA.n1982 GNDA.n995 3.4105
R16420 GNDA.n1016 GNDA.n995 3.4105
R16421 GNDA.n1984 GNDA.n995 3.4105
R16422 GNDA.n1015 GNDA.n995 3.4105
R16423 GNDA.n1986 GNDA.n995 3.4105
R16424 GNDA.n1014 GNDA.n995 3.4105
R16425 GNDA.n1988 GNDA.n995 3.4105
R16426 GNDA.n1013 GNDA.n995 3.4105
R16427 GNDA.n1990 GNDA.n995 3.4105
R16428 GNDA.n1991 GNDA.n995 3.4105
R16429 GNDA.n2011 GNDA.n995 3.4105
R16430 GNDA.n2013 GNDA.n964 3.4105
R16431 GNDA.n1027 GNDA.n964 3.4105
R16432 GNDA.n1962 GNDA.n964 3.4105
R16433 GNDA.n1026 GNDA.n964 3.4105
R16434 GNDA.n1964 GNDA.n964 3.4105
R16435 GNDA.n1025 GNDA.n964 3.4105
R16436 GNDA.n1966 GNDA.n964 3.4105
R16437 GNDA.n1024 GNDA.n964 3.4105
R16438 GNDA.n1968 GNDA.n964 3.4105
R16439 GNDA.n1023 GNDA.n964 3.4105
R16440 GNDA.n1970 GNDA.n964 3.4105
R16441 GNDA.n1022 GNDA.n964 3.4105
R16442 GNDA.n1972 GNDA.n964 3.4105
R16443 GNDA.n1021 GNDA.n964 3.4105
R16444 GNDA.n1974 GNDA.n964 3.4105
R16445 GNDA.n1020 GNDA.n964 3.4105
R16446 GNDA.n1976 GNDA.n964 3.4105
R16447 GNDA.n1019 GNDA.n964 3.4105
R16448 GNDA.n1978 GNDA.n964 3.4105
R16449 GNDA.n1018 GNDA.n964 3.4105
R16450 GNDA.n1980 GNDA.n964 3.4105
R16451 GNDA.n1017 GNDA.n964 3.4105
R16452 GNDA.n1982 GNDA.n964 3.4105
R16453 GNDA.n1016 GNDA.n964 3.4105
R16454 GNDA.n1984 GNDA.n964 3.4105
R16455 GNDA.n1015 GNDA.n964 3.4105
R16456 GNDA.n1986 GNDA.n964 3.4105
R16457 GNDA.n1014 GNDA.n964 3.4105
R16458 GNDA.n1988 GNDA.n964 3.4105
R16459 GNDA.n1013 GNDA.n964 3.4105
R16460 GNDA.n1990 GNDA.n964 3.4105
R16461 GNDA.n1991 GNDA.n964 3.4105
R16462 GNDA.n2011 GNDA.n964 3.4105
R16463 GNDA.n2013 GNDA.n2012 3.4105
R16464 GNDA.n2012 GNDA.n1027 3.4105
R16465 GNDA.n2012 GNDA.n1962 3.4105
R16466 GNDA.n2012 GNDA.n1026 3.4105
R16467 GNDA.n2012 GNDA.n1964 3.4105
R16468 GNDA.n2012 GNDA.n1025 3.4105
R16469 GNDA.n2012 GNDA.n1966 3.4105
R16470 GNDA.n2012 GNDA.n1024 3.4105
R16471 GNDA.n2012 GNDA.n1968 3.4105
R16472 GNDA.n2012 GNDA.n1023 3.4105
R16473 GNDA.n2012 GNDA.n1970 3.4105
R16474 GNDA.n2012 GNDA.n1022 3.4105
R16475 GNDA.n2012 GNDA.n1972 3.4105
R16476 GNDA.n2012 GNDA.n1021 3.4105
R16477 GNDA.n2012 GNDA.n1974 3.4105
R16478 GNDA.n2012 GNDA.n1020 3.4105
R16479 GNDA.n2012 GNDA.n1976 3.4105
R16480 GNDA.n2012 GNDA.n1019 3.4105
R16481 GNDA.n2012 GNDA.n1978 3.4105
R16482 GNDA.n2012 GNDA.n1018 3.4105
R16483 GNDA.n2012 GNDA.n1980 3.4105
R16484 GNDA.n2012 GNDA.n1017 3.4105
R16485 GNDA.n2012 GNDA.n1982 3.4105
R16486 GNDA.n2012 GNDA.n1016 3.4105
R16487 GNDA.n2012 GNDA.n1984 3.4105
R16488 GNDA.n2012 GNDA.n1015 3.4105
R16489 GNDA.n2012 GNDA.n1986 3.4105
R16490 GNDA.n2012 GNDA.n1014 3.4105
R16491 GNDA.n2012 GNDA.n1988 3.4105
R16492 GNDA.n2012 GNDA.n1013 3.4105
R16493 GNDA.n2012 GNDA.n1990 3.4105
R16494 GNDA.n2012 GNDA.n1012 3.4105
R16495 GNDA.n2012 GNDA.n1991 3.4105
R16496 GNDA.n2012 GNDA.n2011 3.4105
R16497 GNDA.n3138 GNDA.n3137 3.39217
R16498 GNDA.n3140 GNDA.n3139 3.39217
R16499 GNDA.n637 GNDA.n636 3.39217
R16500 GNDA.n639 GNDA.n638 3.39217
R16501 GNDA.n3134 GNDA.n3130 3.13621
R16502 GNDA.n3135 GNDA.n3134 3.13621
R16503 GNDA.n633 GNDA.n630 3.13621
R16504 GNDA.n634 GNDA.n633 3.13621
R16505 GNDA.n3030 GNDA.n699 3.04346
R16506 GNDA.n2500 GNDA.n2499 3.00528
R16507 GNDA.n3063 GNDA.n3062 3.00528
R16508 GNDA.n2999 GNDA.t7 3.00528
R16509 GNDA.n723 GNDA.t19 3.00528
R16510 GNDA.n3017 GNDA.n704 2.86505
R16511 GNDA.n3018 GNDA.n3017 2.86505
R16512 GNDA.n3016 GNDA.n3012 2.86505
R16513 GNDA.n3013 GNDA.n3012 2.86505
R16514 GNDA.n3019 GNDA.n3018 2.86505
R16515 GNDA.n3014 GNDA.n3013 2.86505
R16516 GNDA.n3023 GNDA.n704 2.86505
R16517 GNDA.n3019 GNDA.n3016 2.86505
R16518 GNDA.n2404 GNDA.n2403 2.86505
R16519 GNDA.n2403 GNDA.n2401 2.86505
R16520 GNDA.n2401 GNDA.n2400 2.86505
R16521 GNDA.n2405 GNDA.n2404 2.86505
R16522 GNDA.n2237 GNDA.n2233 2.69842
R16523 GNDA.n803 GNDA.n802 2.6629
R16524 GNDA.n2324 GNDA.n2323 2.6629
R16525 GNDA.n2379 GNDA.n804 2.6629
R16526 GNDA.n5056 GNDA.n5055 2.6629
R16527 GNDA.n2574 GNDA.n2573 2.6629
R16528 GNDA.n2701 GNDA.n2700 2.6629
R16529 GNDA.n4985 GNDA.n4984 2.6629
R16530 GNDA.n4898 GNDA.n160 2.6629
R16531 GNDA.n5264 GNDA.n5263 2.6629
R16532 GNDA.n5177 GNDA.n82 2.6629
R16533 GNDA.n4841 GNDA.n4840 2.6629
R16534 GNDA.n4749 GNDA.n56 2.6629
R16535 GNDA.n2517 GNDA.n836 2.6629
R16536 GNDA.n2316 GNDA.n2315 2.6629
R16537 GNDA.n5171 GNDA.n5170 2.6629
R16538 GNDA.t45 GNDA.t93 2.59854
R16539 GNDA.n804 GNDA.n803 2.4581
R16540 GNDA.n3044 GNDA.n3043 2.4581
R16541 GNDA.n2323 GNDA.n2316 2.4581
R16542 GNDA.n2380 GNDA.n2379 2.4581
R16543 GNDA.n5056 GNDA.n160 2.4581
R16544 GNDA.n2573 GNDA.n186 2.4581
R16545 GNDA.n2700 GNDA.n2574 2.4581
R16546 GNDA.n2738 GNDA.n2737 2.4581
R16547 GNDA.n4899 GNDA.n4898 2.4581
R16548 GNDA.n5264 GNDA.n56 2.4581
R16549 GNDA.n5178 GNDA.n5177 2.4581
R16550 GNDA.n4750 GNDA.n4749 2.4581
R16551 GNDA.n2315 GNDA.n2268 2.4581
R16552 GNDA.n5171 GNDA.n82 2.4581
R16553 GNDA.n5104 GNDA.n5103 2.4581
R16554 GNDA.n3033 GNDA.n3032 2.44675
R16555 GNDA.n3032 GNDA.n3031 2.44675
R16556 GNDA.n2075 GNDA.n2074 2.39683
R16557 GNDA.n2165 GNDA.n2164 2.30736
R16558 GNDA.n3672 GNDA.n3664 2.30736
R16559 GNDA.n3380 GNDA.n3379 2.30736
R16560 GNDA.n4577 GNDA.n4576 2.30736
R16561 GNDA.n4501 GNDA.n4500 2.30736
R16562 GNDA.n4419 GNDA.n4418 2.30736
R16563 GNDA.n4337 GNDA.n4336 2.30736
R16564 GNDA.n4255 GNDA.n4254 2.30736
R16565 GNDA.n4009 GNDA.n4008 2.30736
R16566 GNDA.n4173 GNDA.n4172 2.30736
R16567 GNDA.n4091 GNDA.n4090 2.30736
R16568 GNDA.n3906 GNDA.n3905 2.30736
R16569 GNDA.n1730 GNDA.n1729 2.30736
R16570 GNDA.n3848 GNDA.n3847 2.30736
R16571 GNDA.n3772 GNDA.n3771 2.30736
R16572 GNDA.n3614 GNDA.n3613 2.30736
R16573 GNDA.n3538 GNDA.n3537 2.30736
R16574 GNDA.n3435 GNDA.n3434 2.30736
R16575 GNDA.n3304 GNDA.n3303 2.30736
R16576 GNDA.n3201 GNDA.n3200 2.30736
R16577 GNDA.n1654 GNDA.n1653 2.30736
R16578 GNDA.n1572 GNDA.n1571 2.30736
R16579 GNDA.n1490 GNDA.n1489 2.30736
R16580 GNDA.n1212 GNDA.n1211 2.30736
R16581 GNDA.n1922 GNDA.n1921 2.30736
R16582 GNDA.n1806 GNDA.n1801 2.30736
R16583 GNDA.n4625 GNDA.n4624 2.29914
R16584 GNDA.n4627 GNDA.n4626 2.29914
R16585 GNDA.n3150 GNDA.n3149 2.29914
R16586 GNDA.n1744 GNDA.n626 2.29878
R16587 GNDA.n2226 GNDA.n2225 2.29738
R16588 GNDA.n1329 GNDA.n1278 2.26187
R16589 GNDA.n1287 GNDA.n1284 2.26187
R16590 GNDA.n1288 GNDA.n1287 2.26187
R16591 GNDA.n1347 GNDA.n1270 2.26187
R16592 GNDA.n1353 GNDA.n1268 2.26187
R16593 GNDA.n1381 GNDA.n1259 2.26187
R16594 GNDA.n1761 GNDA.n1389 2.26187
R16595 GNDA.n4608 GNDA.n450 2.26187
R16596 GNDA.n2299 GNDA.n2298 2.26187
R16597 GNDA.n3027 GNDA.n3026 2.26187
R16598 GNDA.n2232 GNDA.n842 2.26187
R16599 GNDA.n2236 GNDA.n2235 2.26187
R16600 GNDA.n2235 GNDA.n839 2.26187
R16601 GNDA.n1350 GNDA.n1267 2.26187
R16602 GNDA.n1301 GNDA.n1290 2.26187
R16603 GNDA.n1327 GNDA.n1326 2.26187
R16604 GNDA.n1332 GNDA.n1331 2.26187
R16605 GNDA.n1335 GNDA.n1276 2.26187
R16606 GNDA.n1344 GNDA.n1270 2.26187
R16607 GNDA.n1378 GNDA.n1259 2.26187
R16608 GNDA.n1848 GNDA.n1845 2.26187
R16609 GNDA.n1853 GNDA.n1842 2.26187
R16610 GNDA.n1858 GNDA.n1771 2.26187
R16611 GNDA.n3028 GNDA.n3027 2.26187
R16612 GNDA.n2281 GNDA.n2280 2.26187
R16613 GNDA.n1739 GNDA.n1406 2.24241
R16614 GNDA.n1740 GNDA.n1405 2.24241
R16615 GNDA.n3952 GNDA.n437 2.24241
R16616 GNDA.n504 GNDA.n503 2.24241
R16617 GNDA.n1302 GNDA.n1301 2.24063
R16618 GNDA.n1300 GNDA.n1291 2.24063
R16619 GNDA.n1331 GNDA.n1330 2.24063
R16620 GNDA.n1324 GNDA.n1323 2.24063
R16621 GNDA.n1326 GNDA.n1325 2.24063
R16622 GNDA.n1336 GNDA.n1335 2.24063
R16623 GNDA.n1334 GNDA.n1277 2.24063
R16624 GNDA.n1348 GNDA.n1269 2.24063
R16625 GNDA.n1354 GNDA.n1267 2.24063
R16626 GNDA.n1358 GNDA.n628 2.24063
R16627 GNDA.n1266 GNDA.n1265 2.24063
R16628 GNDA.n1359 GNDA.n1264 2.24063
R16629 GNDA.n1362 GNDA.n1361 2.24063
R16630 GNDA.n1263 GNDA.n1262 2.24063
R16631 GNDA.n1382 GNDA.n1258 2.24063
R16632 GNDA.n1383 GNDA.n1255 2.24063
R16633 GNDA.n1257 GNDA.n1254 2.24063
R16634 GNDA.n1298 GNDA.n1297 2.24063
R16635 GNDA.n1293 GNDA.n1292 2.24063
R16636 GNDA.n1295 GNDA.n1294 2.24063
R16637 GNDA.n1851 GNDA.n1845 2.24063
R16638 GNDA.n1846 GNDA.n1844 2.24063
R16639 GNDA.n1856 GNDA.n1842 2.24063
R16640 GNDA.n1843 GNDA.n1841 2.24063
R16641 GNDA.n1861 GNDA.n1771 2.24063
R16642 GNDA.n1772 GNDA.n1770 2.24063
R16643 GNDA.n1865 GNDA.n1767 2.24063
R16644 GNDA.n1769 GNDA.n1768 2.24063
R16645 GNDA.n1866 GNDA.n1166 2.24063
R16646 GNDA.n1763 GNDA.n1252 2.24063
R16647 GNDA.n1764 GNDA.n1251 2.24063
R16648 GNDA.n1765 GNDA.n1250 2.24063
R16649 GNDA.n1755 GNDA.n1395 2.24063
R16650 GNDA.n1756 GNDA.n1394 2.24063
R16651 GNDA.n1757 GNDA.n1393 2.24063
R16652 GNDA.n1751 GNDA.n1400 2.24063
R16653 GNDA.n1752 GNDA.n1399 2.24063
R16654 GNDA.n1753 GNDA.n1398 2.24063
R16655 GNDA.n1741 GNDA.n1404 2.24063
R16656 GNDA.n3243 GNDA.n622 2.24063
R16657 GNDA.n623 GNDA.n621 2.24063
R16658 GNDA.n3240 GNDA.n3239 2.24063
R16659 GNDA.n3247 GNDA.n588 2.24063
R16660 GNDA.n620 GNDA.n619 2.24063
R16661 GNDA.n3248 GNDA.n618 2.24063
R16662 GNDA.n3477 GNDA.n582 2.24063
R16663 GNDA.n583 GNDA.n581 2.24063
R16664 GNDA.n3474 GNDA.n3473 2.24063
R16665 GNDA.n3481 GNDA.n548 2.24063
R16666 GNDA.n580 GNDA.n579 2.24063
R16667 GNDA.n3482 GNDA.n578 2.24063
R16668 GNDA.n3624 GNDA.n546 2.24063
R16669 GNDA.n547 GNDA.n545 2.24063
R16670 GNDA.n3621 GNDA.n3620 2.24063
R16671 GNDA.n3715 GNDA.n508 2.24063
R16672 GNDA.n540 GNDA.n539 2.24063
R16673 GNDA.n3716 GNDA.n538 2.24063
R16674 GNDA.n3858 GNDA.n506 2.24063
R16675 GNDA.n507 GNDA.n505 2.24063
R16676 GNDA.n3855 GNDA.n3854 2.24063
R16677 GNDA.n4614 GNDA.n442 2.24063
R16678 GNDA.n4615 GNDA.n441 2.24063
R16679 GNDA.n4616 GNDA.n440 2.24063
R16680 GNDA.n4610 GNDA.n447 2.24063
R16681 GNDA.n4611 GNDA.n446 2.24063
R16682 GNDA.n4612 GNDA.n445 2.24063
R16683 GNDA.n3953 GNDA.n502 2.24063
R16684 GNDA.n4602 GNDA.n456 2.24063
R16685 GNDA.n4603 GNDA.n455 2.24063
R16686 GNDA.n4604 GNDA.n454 2.24063
R16687 GNDA.n4598 GNDA.n461 2.24063
R16688 GNDA.n4599 GNDA.n460 2.24063
R16689 GNDA.n4600 GNDA.n459 2.24063
R16690 GNDA.n4594 GNDA.n466 2.24063
R16691 GNDA.n4595 GNDA.n465 2.24063
R16692 GNDA.n4596 GNDA.n464 2.24063
R16693 GNDA.n4590 GNDA.n471 2.24063
R16694 GNDA.n4591 GNDA.n470 2.24063
R16695 GNDA.n4592 GNDA.n469 2.24063
R16696 GNDA.n4586 GNDA.n4585 2.24063
R16697 GNDA.n4587 GNDA.n4584 2.24063
R16698 GNDA.n4588 GNDA.n4583 2.24063
R16699 GNDA.n1759 GNDA.n1389 2.24063
R16700 GNDA.n1760 GNDA.n1390 2.24063
R16701 GNDA.n4606 GNDA.n450 2.24063
R16702 GNDA.n4607 GNDA.n451 2.24063
R16703 GNDA.n3390 GNDA.n585 2.24063
R16704 GNDA.n587 GNDA.n584 2.24063
R16705 GNDA.n3387 GNDA.n3386 2.24063
R16706 GNDA.n3711 GNDA.n542 2.24063
R16707 GNDA.n544 GNDA.n541 2.24063
R16708 GNDA.n3708 GNDA.n3707 2.24063
R16709 GNDA.n2298 GNDA.n2297 2.24063
R16710 GNDA.n2280 GNDA.n703 2.24063
R16711 GNDA.n2283 GNDA.n2282 2.24063
R16712 GNDA.n3026 GNDA.n3025 2.24063
R16713 GNDA.n2216 GNDA.n2215 2.24063
R16714 GNDA.n2214 GNDA.n2213 2.24063
R16715 GNDA.n2233 GNDA.n841 2.24063
R16716 GNDA.n1333 GNDA.n1278 2.24063
R16717 GNDA.n1328 GNDA.n1281 2.24063
R16718 GNDA.n1319 GNDA.n1284 2.24063
R16719 GNDA.n1318 GNDA.n1317 2.24063
R16720 GNDA.n1344 GNDA.n1343 2.24063
R16721 GNDA.n1349 GNDA.n1268 2.24063
R16722 GNDA.n1360 GNDA.n1261 2.24063
R16723 GNDA.n1378 GNDA.n1377 2.24063
R16724 GNDA.n1385 GNDA.n1384 2.24063
R16725 GNDA.n2394 GNDA.n2284 2.24063
R16726 GNDA.n2393 GNDA.n2392 2.24063
R16727 GNDA.n3029 GNDA.n700 2.24063
R16728 GNDA.n2217 GNDA.n2206 2.24063
R16729 GNDA.n2226 GNDA.n842 2.24063
R16730 GNDA.n2229 GNDA.n2228 2.24063
R16731 GNDA.n2237 GNDA.n2236 2.24063
R16732 GNDA.n2239 GNDA.n2238 2.24063
R16733 GNDA.n2296 GNDA.n2287 2.22018
R16734 GNDA.n2391 GNDA.n2300 2.22018
R16735 GNDA.n2208 GNDA.n2207 2.22018
R16736 GNDA.t61 GNDA.t187 2.21824
R16737 GNDA.t170 GNDA.t55 2.21824
R16738 GNDA.t207 GNDA.t130 2.21824
R16739 GNDA.t86 GNDA.t38 2.21824
R16740 GNDA.n1274 GNDA.n1273 2.19633
R16741 GNDA.n1272 GNDA.n1271 2.19633
R16742 GNDA.n3100 GNDA.n641 2.19633
R16743 GNDA.n328 GNDA.n56 2.18124
R16744 GNDA.n5060 GNDA.n160 2.18124
R16745 GNDA.n2316 GNDA.n812 2.18124
R16746 GNDA.n389 GNDA.n82 2.18124
R16747 GNDA.n2820 GNDA.n2574 2.18124
R16748 GNDA.n2980 GNDA.n804 2.18124
R16749 GNDA.n2218 GNDA.n2217 2.16717
R16750 GNDA.n3045 GNDA.n3044 2.1509
R16751 GNDA.n2381 GNDA.n2380 2.1509
R16752 GNDA.n4991 GNDA.n186 2.1509
R16753 GNDA.n2737 GNDA.n2736 2.1509
R16754 GNDA.n4917 GNDA.n4899 2.1509
R16755 GNDA.n5196 GNDA.n5178 2.1509
R16756 GNDA.n4776 GNDA.n4750 2.1509
R16757 GNDA.n2274 GNDA.n2268 2.1509
R16758 GNDA.n5114 GNDA.n5104 2.1509
R16759 GNDA.n802 GNDA.n801 2.13383
R16760 GNDA.n2325 GNDA.n2324 2.13383
R16761 GNDA.n5055 GNDA.n164 2.13383
R16762 GNDA.n4840 GNDA.n4727 2.13383
R16763 GNDA.n2701 GNDA.n2699 2.13383
R16764 GNDA.n4984 GNDA.n4871 2.13383
R16765 GNDA.n5263 GNDA.n57 2.13383
R16766 GNDA.n2486 GNDA.n836 2.13383
R16767 GNDA.n5170 GNDA.n5169 2.13383
R16768 GNDA.n4620 GNDA.n4619 2.09414
R16769 GNDA.n3155 GNDA.n3154 2.09414
R16770 GNDA.n1749 GNDA.n1748 2.09414
R16771 GNDA.n3860 GNDA.n3859 2.09414
R16772 GNDA.n133 GNDA.n56 2.08643
R16773 GNDA.n162 GNDA.n160 2.08643
R16774 GNDA.n2316 GNDA.n811 2.08643
R16775 GNDA.n84 GNDA.n82 2.08643
R16776 GNDA.n2823 GNDA.n2574 2.08643
R16777 GNDA.n804 GNDA.n748 2.08643
R16778 GNDA.n3125 GNDA.n543 2.0005
R16779 GNDA.n641 GNDA.n586 2.0005
R16780 GNDA.t204 GNDA.t32 1.98114
R16781 GNDA.t40 GNDA.t148 1.98114
R16782 GNDA.n802 GNDA.n745 1.9461
R16783 GNDA.n2324 GNDA.n671 1.9461
R16784 GNDA.n5055 GNDA.n5054 1.9461
R16785 GNDA.n2702 GNDA.n2701 1.9461
R16786 GNDA.n4984 GNDA.n4983 1.9461
R16787 GNDA.n5263 GNDA.n5262 1.9461
R16788 GNDA.n4840 GNDA.n4839 1.9461
R16789 GNDA.n2489 GNDA.n836 1.9461
R16790 GNDA.n5170 GNDA.n22 1.9461
R16791 GNDA.n3137 GNDA.n629 1.94497
R16792 GNDA.n3141 GNDA.n3140 1.94497
R16793 GNDA.n4624 GNDA.n4623 1.93383
R16794 GNDA.n4628 GNDA.n4627 1.93383
R16795 GNDA.n3151 GNDA.n3150 1.93383
R16796 GNDA.n1745 GNDA.n1744 1.93383
R16797 GNDA.n3126 GNDA.n3125 1.91062
R16798 GNDA.n1295 GNDA.n449 1.82342
R16799 GNDA.n1388 GNDA.n1387 1.82342
R16800 GNDA.n3025 GNDA.n3024 1.71925
R16801 GNDA.n2050 GNDA.n879 1.70567
R16802 GNDA.n2050 GNDA.n878 1.70567
R16803 GNDA.n2050 GNDA.n877 1.70567
R16804 GNDA.n2050 GNDA.n876 1.70567
R16805 GNDA.n2050 GNDA.n875 1.70567
R16806 GNDA.n2050 GNDA.n874 1.70567
R16807 GNDA.n2050 GNDA.n873 1.70567
R16808 GNDA.n2050 GNDA.n872 1.70567
R16809 GNDA.n2050 GNDA.n871 1.70567
R16810 GNDA.n2050 GNDA.n870 1.70567
R16811 GNDA.n2050 GNDA.n869 1.70567
R16812 GNDA.n2050 GNDA.n868 1.70567
R16813 GNDA.n2050 GNDA.n867 1.70567
R16814 GNDA.n2050 GNDA.n866 1.70567
R16815 GNDA.n2050 GNDA.n865 1.70567
R16816 GNDA.n2050 GNDA.n864 1.70567
R16817 GNDA.n2052 GNDA.n2051 1.70567
R16818 GNDA.n2016 GNDA.n863 1.70567
R16819 GNDA.n2018 GNDA.n863 1.70567
R16820 GNDA.n2020 GNDA.n863 1.70567
R16821 GNDA.n2022 GNDA.n863 1.70567
R16822 GNDA.n2024 GNDA.n863 1.70567
R16823 GNDA.n2026 GNDA.n863 1.70567
R16824 GNDA.n2028 GNDA.n863 1.70567
R16825 GNDA.n2030 GNDA.n863 1.70567
R16826 GNDA.n2032 GNDA.n863 1.70567
R16827 GNDA.n2034 GNDA.n863 1.70567
R16828 GNDA.n2036 GNDA.n863 1.70567
R16829 GNDA.n2038 GNDA.n863 1.70567
R16830 GNDA.n2040 GNDA.n863 1.70567
R16831 GNDA.n2042 GNDA.n863 1.70567
R16832 GNDA.n2044 GNDA.n863 1.70567
R16833 GNDA.n2046 GNDA.n863 1.70567
R16834 GNDA.n898 GNDA.n897 1.70567
R16835 GNDA.n2052 GNDA.n862 1.70567
R16836 GNDA.n900 GNDA.n897 1.70567
R16837 GNDA.n2052 GNDA.n861 1.70567
R16838 GNDA.n902 GNDA.n897 1.70567
R16839 GNDA.n2052 GNDA.n860 1.70567
R16840 GNDA.n904 GNDA.n897 1.70567
R16841 GNDA.n2052 GNDA.n859 1.70567
R16842 GNDA.n906 GNDA.n897 1.70567
R16843 GNDA.n2052 GNDA.n858 1.70567
R16844 GNDA.n908 GNDA.n897 1.70567
R16845 GNDA.n2052 GNDA.n857 1.70567
R16846 GNDA.n910 GNDA.n897 1.70567
R16847 GNDA.n2052 GNDA.n856 1.70567
R16848 GNDA.n912 GNDA.n897 1.70567
R16849 GNDA.n2052 GNDA.n855 1.70567
R16850 GNDA.n914 GNDA.n897 1.70567
R16851 GNDA.n2052 GNDA.n854 1.70567
R16852 GNDA.n916 GNDA.n897 1.70567
R16853 GNDA.n2052 GNDA.n853 1.70567
R16854 GNDA.n918 GNDA.n897 1.70567
R16855 GNDA.n2052 GNDA.n852 1.70567
R16856 GNDA.n920 GNDA.n897 1.70567
R16857 GNDA.n2052 GNDA.n851 1.70567
R16858 GNDA.n922 GNDA.n897 1.70567
R16859 GNDA.n2052 GNDA.n850 1.70567
R16860 GNDA.n924 GNDA.n897 1.70567
R16861 GNDA.n2052 GNDA.n849 1.70567
R16862 GNDA.n926 GNDA.n897 1.70567
R16863 GNDA.n2052 GNDA.n848 1.70567
R16864 GNDA.n928 GNDA.n897 1.70567
R16865 GNDA.n2052 GNDA.n847 1.70567
R16866 GNDA.n2048 GNDA.n846 1.70567
R16867 GNDA.n930 GNDA.n897 1.70567
R16868 GNDA.n1960 GNDA.n1044 1.70567
R16869 GNDA.n1960 GNDA.n1043 1.70567
R16870 GNDA.n1960 GNDA.n1042 1.70567
R16871 GNDA.n1960 GNDA.n1041 1.70567
R16872 GNDA.n1960 GNDA.n1040 1.70567
R16873 GNDA.n1960 GNDA.n1039 1.70567
R16874 GNDA.n1960 GNDA.n1038 1.70567
R16875 GNDA.n1960 GNDA.n1037 1.70567
R16876 GNDA.n1960 GNDA.n1036 1.70567
R16877 GNDA.n1960 GNDA.n1035 1.70567
R16878 GNDA.n1960 GNDA.n1034 1.70567
R16879 GNDA.n1960 GNDA.n1033 1.70567
R16880 GNDA.n1960 GNDA.n1032 1.70567
R16881 GNDA.n1960 GNDA.n1031 1.70567
R16882 GNDA.n1960 GNDA.n1030 1.70567
R16883 GNDA.n1960 GNDA.n1029 1.70567
R16884 GNDA.n1927 GNDA.n1062 1.70567
R16885 GNDA.n1929 GNDA.n1062 1.70567
R16886 GNDA.n1931 GNDA.n1062 1.70567
R16887 GNDA.n1933 GNDA.n1062 1.70567
R16888 GNDA.n1935 GNDA.n1062 1.70567
R16889 GNDA.n1937 GNDA.n1062 1.70567
R16890 GNDA.n1939 GNDA.n1062 1.70567
R16891 GNDA.n1941 GNDA.n1062 1.70567
R16892 GNDA.n1943 GNDA.n1062 1.70567
R16893 GNDA.n1945 GNDA.n1062 1.70567
R16894 GNDA.n1947 GNDA.n1062 1.70567
R16895 GNDA.n1949 GNDA.n1062 1.70567
R16896 GNDA.n1951 GNDA.n1062 1.70567
R16897 GNDA.n1953 GNDA.n1062 1.70567
R16898 GNDA.n1955 GNDA.n1062 1.70567
R16899 GNDA.n1063 GNDA.n1028 1.70567
R16900 GNDA.n1112 GNDA.n1096 1.70567
R16901 GNDA.n1064 GNDA.n1063 1.70567
R16902 GNDA.n1112 GNDA.n1097 1.70567
R16903 GNDA.n1066 GNDA.n1063 1.70567
R16904 GNDA.n1112 GNDA.n1098 1.70567
R16905 GNDA.n1068 GNDA.n1063 1.70567
R16906 GNDA.n1112 GNDA.n1099 1.70567
R16907 GNDA.n1070 GNDA.n1063 1.70567
R16908 GNDA.n1112 GNDA.n1100 1.70567
R16909 GNDA.n1072 GNDA.n1063 1.70567
R16910 GNDA.n1112 GNDA.n1101 1.70567
R16911 GNDA.n1074 GNDA.n1063 1.70567
R16912 GNDA.n1112 GNDA.n1102 1.70567
R16913 GNDA.n1076 GNDA.n1063 1.70567
R16914 GNDA.n1112 GNDA.n1103 1.70567
R16915 GNDA.n1078 GNDA.n1063 1.70567
R16916 GNDA.n1112 GNDA.n1104 1.70567
R16917 GNDA.n1080 GNDA.n1063 1.70567
R16918 GNDA.n1112 GNDA.n1105 1.70567
R16919 GNDA.n1082 GNDA.n1063 1.70567
R16920 GNDA.n1112 GNDA.n1106 1.70567
R16921 GNDA.n1084 GNDA.n1063 1.70567
R16922 GNDA.n1112 GNDA.n1107 1.70567
R16923 GNDA.n1086 GNDA.n1063 1.70567
R16924 GNDA.n1112 GNDA.n1108 1.70567
R16925 GNDA.n1088 GNDA.n1063 1.70567
R16926 GNDA.n1112 GNDA.n1109 1.70567
R16927 GNDA.n1090 GNDA.n1063 1.70567
R16928 GNDA.n1112 GNDA.n1110 1.70567
R16929 GNDA.n1092 GNDA.n1063 1.70567
R16930 GNDA.n1112 GNDA.n1111 1.70567
R16931 GNDA.n1094 GNDA.n1063 1.70567
R16932 GNDA.n1113 GNDA.n1112 1.70567
R16933 GNDA.n1958 GNDA.n1957 1.70567
R16934 GNDA.n2014 GNDA.n2013 1.70567
R16935 GNDA.n2015 GNDA.n962 1.70567
R16936 GNDA.n2015 GNDA.n961 1.70567
R16937 GNDA.n2015 GNDA.n960 1.70567
R16938 GNDA.n2015 GNDA.n959 1.70567
R16939 GNDA.n2015 GNDA.n958 1.70567
R16940 GNDA.n2015 GNDA.n957 1.70567
R16941 GNDA.n2015 GNDA.n956 1.70567
R16942 GNDA.n2015 GNDA.n955 1.70567
R16943 GNDA.n2015 GNDA.n954 1.70567
R16944 GNDA.n2015 GNDA.n953 1.70567
R16945 GNDA.n2015 GNDA.n952 1.70567
R16946 GNDA.n2015 GNDA.n951 1.70567
R16947 GNDA.n2015 GNDA.n950 1.70567
R16948 GNDA.n2015 GNDA.n949 1.70567
R16949 GNDA.n2015 GNDA.n948 1.70567
R16950 GNDA.n2015 GNDA.n947 1.70567
R16951 GNDA.n2015 GNDA.n946 1.70567
R16952 GNDA.n1961 GNDA.n963 1.70567
R16953 GNDA.n1963 GNDA.n963 1.70567
R16954 GNDA.n1965 GNDA.n963 1.70567
R16955 GNDA.n1967 GNDA.n963 1.70567
R16956 GNDA.n1969 GNDA.n963 1.70567
R16957 GNDA.n1971 GNDA.n963 1.70567
R16958 GNDA.n1973 GNDA.n963 1.70567
R16959 GNDA.n1975 GNDA.n963 1.70567
R16960 GNDA.n1977 GNDA.n963 1.70567
R16961 GNDA.n1979 GNDA.n963 1.70567
R16962 GNDA.n1981 GNDA.n963 1.70567
R16963 GNDA.n1983 GNDA.n963 1.70567
R16964 GNDA.n1985 GNDA.n963 1.70567
R16965 GNDA.n1987 GNDA.n963 1.70567
R16966 GNDA.n1989 GNDA.n963 1.70567
R16967 GNDA.n2010 GNDA.n980 1.70567
R16968 GNDA.n2008 GNDA.n2007 1.70567
R16969 GNDA.n2009 GNDA.n1012 1.70567
R16970 GNDA.n2007 GNDA.n1992 1.70567
R16971 GNDA.n1012 GNDA.n1011 1.70567
R16972 GNDA.n2007 GNDA.n1993 1.70567
R16973 GNDA.n1012 GNDA.n1010 1.70567
R16974 GNDA.n2007 GNDA.n1994 1.70567
R16975 GNDA.n1012 GNDA.n1009 1.70567
R16976 GNDA.n2007 GNDA.n1995 1.70567
R16977 GNDA.n1012 GNDA.n1008 1.70567
R16978 GNDA.n2007 GNDA.n1996 1.70567
R16979 GNDA.n1012 GNDA.n1007 1.70567
R16980 GNDA.n2007 GNDA.n1997 1.70567
R16981 GNDA.n1012 GNDA.n1006 1.70567
R16982 GNDA.n2007 GNDA.n1998 1.70567
R16983 GNDA.n1012 GNDA.n1005 1.70567
R16984 GNDA.n2007 GNDA.n1999 1.70567
R16985 GNDA.n1012 GNDA.n1004 1.70567
R16986 GNDA.n2007 GNDA.n2000 1.70567
R16987 GNDA.n1012 GNDA.n1003 1.70567
R16988 GNDA.n2007 GNDA.n2001 1.70567
R16989 GNDA.n1012 GNDA.n1002 1.70567
R16990 GNDA.n2007 GNDA.n2002 1.70567
R16991 GNDA.n1012 GNDA.n1001 1.70567
R16992 GNDA.n2007 GNDA.n2003 1.70567
R16993 GNDA.n1012 GNDA.n1000 1.70567
R16994 GNDA.n2007 GNDA.n2004 1.70567
R16995 GNDA.n1012 GNDA.n999 1.70567
R16996 GNDA.n2007 GNDA.n2005 1.70567
R16997 GNDA.n1012 GNDA.n998 1.70567
R16998 GNDA.n2007 GNDA.n2006 1.70567
R16999 GNDA.n1012 GNDA.n997 1.70567
R17000 GNDA.n2007 GNDA.n996 1.70567
R17001 GNDA.n1924 GNDA.n1150 1.69433
R17002 GNDA.n1924 GNDA.n1147 1.69433
R17003 GNDA.n1924 GNDA.n1144 1.69433
R17004 GNDA.n1221 GNDA.n1153 1.69433
R17005 GNDA.n1230 GNDA.n1153 1.69433
R17006 GNDA.n1239 GNDA.n1153 1.69433
R17007 GNDA.n1492 GNDA.n1420 1.69433
R17008 GNDA.n1492 GNDA.n1417 1.69433
R17009 GNDA.n1492 GNDA.n1414 1.69433
R17010 GNDA.n1574 GNDA.n1502 1.69433
R17011 GNDA.n1574 GNDA.n1499 1.69433
R17012 GNDA.n1574 GNDA.n1496 1.69433
R17013 GNDA.n1656 GNDA.n1584 1.69433
R17014 GNDA.n1656 GNDA.n1581 1.69433
R17015 GNDA.n1656 GNDA.n1578 1.69433
R17016 GNDA.n3210 GNDA.n593 1.69433
R17017 GNDA.n3219 GNDA.n593 1.69433
R17018 GNDA.n3228 GNDA.n593 1.69433
R17019 GNDA.n3306 GNDA.n603 1.69433
R17020 GNDA.n3306 GNDA.n600 1.69433
R17021 GNDA.n3306 GNDA.n597 1.69433
R17022 GNDA.n3444 GNDA.n553 1.69433
R17023 GNDA.n3453 GNDA.n553 1.69433
R17024 GNDA.n3462 GNDA.n553 1.69433
R17025 GNDA.n3540 GNDA.n563 1.69433
R17026 GNDA.n3540 GNDA.n560 1.69433
R17027 GNDA.n3540 GNDA.n557 1.69433
R17028 GNDA.n3616 GNDA.n3549 1.69433
R17029 GNDA.n3616 GNDA.n3546 1.69433
R17030 GNDA.n3616 GNDA.n3543 1.69433
R17031 GNDA.n3774 GNDA.n523 1.69433
R17032 GNDA.n3774 GNDA.n520 1.69433
R17033 GNDA.n3774 GNDA.n517 1.69433
R17034 GNDA.n3850 GNDA.n3783 1.69433
R17035 GNDA.n3850 GNDA.n3780 1.69433
R17036 GNDA.n3850 GNDA.n3777 1.69433
R17037 GNDA.n1732 GNDA.n1665 1.69433
R17038 GNDA.n1732 GNDA.n1662 1.69433
R17039 GNDA.n1732 GNDA.n1659 1.69433
R17040 GNDA.n3915 GNDA.n477 1.69433
R17041 GNDA.n3924 GNDA.n477 1.69433
R17042 GNDA.n3933 GNDA.n477 1.69433
R17043 GNDA.n4093 GNDA.n4021 1.69433
R17044 GNDA.n4093 GNDA.n4018 1.69433
R17045 GNDA.n4093 GNDA.n4015 1.69433
R17046 GNDA.n4175 GNDA.n4103 1.69433
R17047 GNDA.n4175 GNDA.n4100 1.69433
R17048 GNDA.n4175 GNDA.n4097 1.69433
R17049 GNDA.n4011 GNDA.n487 1.69433
R17050 GNDA.n4011 GNDA.n484 1.69433
R17051 GNDA.n4011 GNDA.n481 1.69433
R17052 GNDA.n4257 GNDA.n4185 1.69433
R17053 GNDA.n4257 GNDA.n4182 1.69433
R17054 GNDA.n4257 GNDA.n4179 1.69433
R17055 GNDA.n4339 GNDA.n4267 1.69433
R17056 GNDA.n4339 GNDA.n4264 1.69433
R17057 GNDA.n4339 GNDA.n4261 1.69433
R17058 GNDA.n4421 GNDA.n4349 1.69433
R17059 GNDA.n4421 GNDA.n4346 1.69433
R17060 GNDA.n4421 GNDA.n4343 1.69433
R17061 GNDA.n4503 GNDA.n4431 1.69433
R17062 GNDA.n4503 GNDA.n4428 1.69433
R17063 GNDA.n4503 GNDA.n4425 1.69433
R17064 GNDA.n4579 GNDA.n4512 1.69433
R17065 GNDA.n4579 GNDA.n4509 1.69433
R17066 GNDA.n4579 GNDA.n4506 1.69433
R17067 GNDA.n3382 GNDA.n3315 1.69433
R17068 GNDA.n3382 GNDA.n3312 1.69433
R17069 GNDA.n3382 GNDA.n3309 1.69433
R17070 GNDA.n3661 GNDA.n513 1.69433
R17071 GNDA.n3650 GNDA.n513 1.69433
R17072 GNDA.n3637 GNDA.n513 1.69433
R17073 GNDA.n2222 GNDA.n2062 1.69433
R17074 GNDA.n2222 GNDA.n2059 1.69433
R17075 GNDA.n2222 GNDA.n2056 1.69433
R17076 GNDA.n2221 GNDA.n2137 1.69433
R17077 GNDA.n2221 GNDA.n2134 1.69433
R17078 GNDA.n2221 GNDA.n2131 1.69433
R17079 GNDA.n1925 GNDA.n1139 1.69337
R17080 GNDA.n1925 GNDA.n1138 1.69337
R17081 GNDA.n1925 GNDA.n1136 1.69337
R17082 GNDA.n1925 GNDA.n1135 1.69337
R17083 GNDA.n1925 GNDA.n1133 1.69337
R17084 GNDA.n1925 GNDA.n1132 1.69337
R17085 GNDA.n1925 GNDA.n1130 1.69337
R17086 GNDA.n1925 GNDA.n1129 1.69337
R17087 GNDA.n1924 GNDA.n1152 1.6924
R17088 GNDA.n1924 GNDA.n1151 1.6924
R17089 GNDA.n1924 GNDA.n1149 1.6924
R17090 GNDA.n1924 GNDA.n1148 1.6924
R17091 GNDA.n1924 GNDA.n1146 1.6924
R17092 GNDA.n1924 GNDA.n1145 1.6924
R17093 GNDA.n1924 GNDA.n1143 1.6924
R17094 GNDA.n1924 GNDA.n1142 1.6924
R17095 GNDA.n1215 GNDA.n1153 1.6924
R17096 GNDA.n1218 GNDA.n1153 1.6924
R17097 GNDA.n1224 GNDA.n1153 1.6924
R17098 GNDA.n1227 GNDA.n1153 1.6924
R17099 GNDA.n1233 GNDA.n1153 1.6924
R17100 GNDA.n1236 GNDA.n1153 1.6924
R17101 GNDA.n1242 GNDA.n1153 1.6924
R17102 GNDA.n1245 GNDA.n1153 1.6924
R17103 GNDA.n1492 GNDA.n1422 1.6924
R17104 GNDA.n1492 GNDA.n1421 1.6924
R17105 GNDA.n1492 GNDA.n1419 1.6924
R17106 GNDA.n1492 GNDA.n1418 1.6924
R17107 GNDA.n1492 GNDA.n1416 1.6924
R17108 GNDA.n1492 GNDA.n1415 1.6924
R17109 GNDA.n1492 GNDA.n1413 1.6924
R17110 GNDA.n1492 GNDA.n1412 1.6924
R17111 GNDA.n1574 GNDA.n1504 1.6924
R17112 GNDA.n1574 GNDA.n1503 1.6924
R17113 GNDA.n1574 GNDA.n1501 1.6924
R17114 GNDA.n1574 GNDA.n1500 1.6924
R17115 GNDA.n1574 GNDA.n1498 1.6924
R17116 GNDA.n1574 GNDA.n1497 1.6924
R17117 GNDA.n1574 GNDA.n1495 1.6924
R17118 GNDA.n1574 GNDA.n1494 1.6924
R17119 GNDA.n1656 GNDA.n1586 1.6924
R17120 GNDA.n1656 GNDA.n1585 1.6924
R17121 GNDA.n1656 GNDA.n1583 1.6924
R17122 GNDA.n1656 GNDA.n1582 1.6924
R17123 GNDA.n1656 GNDA.n1580 1.6924
R17124 GNDA.n1656 GNDA.n1579 1.6924
R17125 GNDA.n1656 GNDA.n1577 1.6924
R17126 GNDA.n1656 GNDA.n1576 1.6924
R17127 GNDA.n3204 GNDA.n593 1.6924
R17128 GNDA.n3207 GNDA.n593 1.6924
R17129 GNDA.n3213 GNDA.n593 1.6924
R17130 GNDA.n3216 GNDA.n593 1.6924
R17131 GNDA.n3222 GNDA.n593 1.6924
R17132 GNDA.n3225 GNDA.n593 1.6924
R17133 GNDA.n3231 GNDA.n593 1.6924
R17134 GNDA.n3234 GNDA.n593 1.6924
R17135 GNDA.n3306 GNDA.n605 1.6924
R17136 GNDA.n3306 GNDA.n604 1.6924
R17137 GNDA.n3306 GNDA.n602 1.6924
R17138 GNDA.n3306 GNDA.n601 1.6924
R17139 GNDA.n3306 GNDA.n599 1.6924
R17140 GNDA.n3306 GNDA.n598 1.6924
R17141 GNDA.n3306 GNDA.n596 1.6924
R17142 GNDA.n3306 GNDA.n595 1.6924
R17143 GNDA.n3438 GNDA.n553 1.6924
R17144 GNDA.n3441 GNDA.n553 1.6924
R17145 GNDA.n3447 GNDA.n553 1.6924
R17146 GNDA.n3450 GNDA.n553 1.6924
R17147 GNDA.n3456 GNDA.n553 1.6924
R17148 GNDA.n3459 GNDA.n553 1.6924
R17149 GNDA.n3465 GNDA.n553 1.6924
R17150 GNDA.n3468 GNDA.n553 1.6924
R17151 GNDA.n3540 GNDA.n565 1.6924
R17152 GNDA.n3540 GNDA.n564 1.6924
R17153 GNDA.n3540 GNDA.n562 1.6924
R17154 GNDA.n3540 GNDA.n561 1.6924
R17155 GNDA.n3540 GNDA.n559 1.6924
R17156 GNDA.n3540 GNDA.n558 1.6924
R17157 GNDA.n3540 GNDA.n556 1.6924
R17158 GNDA.n3540 GNDA.n555 1.6924
R17159 GNDA.n3616 GNDA.n3551 1.6924
R17160 GNDA.n3616 GNDA.n3550 1.6924
R17161 GNDA.n3616 GNDA.n3548 1.6924
R17162 GNDA.n3616 GNDA.n3547 1.6924
R17163 GNDA.n3616 GNDA.n3545 1.6924
R17164 GNDA.n3616 GNDA.n3544 1.6924
R17165 GNDA.n3616 GNDA.n3542 1.6924
R17166 GNDA.n3616 GNDA.n3541 1.6924
R17167 GNDA.n3774 GNDA.n525 1.6924
R17168 GNDA.n3774 GNDA.n524 1.6924
R17169 GNDA.n3774 GNDA.n522 1.6924
R17170 GNDA.n3774 GNDA.n521 1.6924
R17171 GNDA.n3774 GNDA.n519 1.6924
R17172 GNDA.n3774 GNDA.n518 1.6924
R17173 GNDA.n3774 GNDA.n516 1.6924
R17174 GNDA.n3774 GNDA.n515 1.6924
R17175 GNDA.n3850 GNDA.n3785 1.6924
R17176 GNDA.n3850 GNDA.n3784 1.6924
R17177 GNDA.n3850 GNDA.n3782 1.6924
R17178 GNDA.n3850 GNDA.n3781 1.6924
R17179 GNDA.n3850 GNDA.n3779 1.6924
R17180 GNDA.n3850 GNDA.n3778 1.6924
R17181 GNDA.n3850 GNDA.n3776 1.6924
R17182 GNDA.n3850 GNDA.n3775 1.6924
R17183 GNDA.n1732 GNDA.n1667 1.6924
R17184 GNDA.n1732 GNDA.n1666 1.6924
R17185 GNDA.n1732 GNDA.n1664 1.6924
R17186 GNDA.n1732 GNDA.n1663 1.6924
R17187 GNDA.n1732 GNDA.n1661 1.6924
R17188 GNDA.n1732 GNDA.n1660 1.6924
R17189 GNDA.n1732 GNDA.n1658 1.6924
R17190 GNDA.n1732 GNDA.n1657 1.6924
R17191 GNDA.n3909 GNDA.n477 1.6924
R17192 GNDA.n3912 GNDA.n477 1.6924
R17193 GNDA.n3918 GNDA.n477 1.6924
R17194 GNDA.n3921 GNDA.n477 1.6924
R17195 GNDA.n3927 GNDA.n477 1.6924
R17196 GNDA.n3930 GNDA.n477 1.6924
R17197 GNDA.n3936 GNDA.n477 1.6924
R17198 GNDA.n3939 GNDA.n477 1.6924
R17199 GNDA.n4093 GNDA.n4023 1.6924
R17200 GNDA.n4093 GNDA.n4022 1.6924
R17201 GNDA.n4093 GNDA.n4020 1.6924
R17202 GNDA.n4093 GNDA.n4019 1.6924
R17203 GNDA.n4093 GNDA.n4017 1.6924
R17204 GNDA.n4093 GNDA.n4016 1.6924
R17205 GNDA.n4093 GNDA.n4014 1.6924
R17206 GNDA.n4093 GNDA.n4013 1.6924
R17207 GNDA.n4175 GNDA.n4105 1.6924
R17208 GNDA.n4175 GNDA.n4104 1.6924
R17209 GNDA.n4175 GNDA.n4102 1.6924
R17210 GNDA.n4175 GNDA.n4101 1.6924
R17211 GNDA.n4175 GNDA.n4099 1.6924
R17212 GNDA.n4175 GNDA.n4098 1.6924
R17213 GNDA.n4175 GNDA.n4096 1.6924
R17214 GNDA.n4175 GNDA.n4095 1.6924
R17215 GNDA.n4011 GNDA.n489 1.6924
R17216 GNDA.n4011 GNDA.n488 1.6924
R17217 GNDA.n4011 GNDA.n486 1.6924
R17218 GNDA.n4011 GNDA.n485 1.6924
R17219 GNDA.n4011 GNDA.n483 1.6924
R17220 GNDA.n4011 GNDA.n482 1.6924
R17221 GNDA.n4011 GNDA.n480 1.6924
R17222 GNDA.n4011 GNDA.n479 1.6924
R17223 GNDA.n4257 GNDA.n4187 1.6924
R17224 GNDA.n4257 GNDA.n4186 1.6924
R17225 GNDA.n4257 GNDA.n4184 1.6924
R17226 GNDA.n4257 GNDA.n4183 1.6924
R17227 GNDA.n4257 GNDA.n4181 1.6924
R17228 GNDA.n4257 GNDA.n4180 1.6924
R17229 GNDA.n4257 GNDA.n4178 1.6924
R17230 GNDA.n4257 GNDA.n4177 1.6924
R17231 GNDA.n4339 GNDA.n4269 1.6924
R17232 GNDA.n4339 GNDA.n4268 1.6924
R17233 GNDA.n4339 GNDA.n4266 1.6924
R17234 GNDA.n4339 GNDA.n4265 1.6924
R17235 GNDA.n4339 GNDA.n4263 1.6924
R17236 GNDA.n4339 GNDA.n4262 1.6924
R17237 GNDA.n4339 GNDA.n4260 1.6924
R17238 GNDA.n4339 GNDA.n4259 1.6924
R17239 GNDA.n4421 GNDA.n4351 1.6924
R17240 GNDA.n4421 GNDA.n4350 1.6924
R17241 GNDA.n4421 GNDA.n4348 1.6924
R17242 GNDA.n4421 GNDA.n4347 1.6924
R17243 GNDA.n4421 GNDA.n4345 1.6924
R17244 GNDA.n4421 GNDA.n4344 1.6924
R17245 GNDA.n4421 GNDA.n4342 1.6924
R17246 GNDA.n4421 GNDA.n4341 1.6924
R17247 GNDA.n4503 GNDA.n4433 1.6924
R17248 GNDA.n4503 GNDA.n4432 1.6924
R17249 GNDA.n4503 GNDA.n4430 1.6924
R17250 GNDA.n4503 GNDA.n4429 1.6924
R17251 GNDA.n4503 GNDA.n4427 1.6924
R17252 GNDA.n4503 GNDA.n4426 1.6924
R17253 GNDA.n4503 GNDA.n4424 1.6924
R17254 GNDA.n4503 GNDA.n4423 1.6924
R17255 GNDA.n4579 GNDA.n4514 1.6924
R17256 GNDA.n4579 GNDA.n4513 1.6924
R17257 GNDA.n4579 GNDA.n4511 1.6924
R17258 GNDA.n4579 GNDA.n4510 1.6924
R17259 GNDA.n4579 GNDA.n4508 1.6924
R17260 GNDA.n4579 GNDA.n4507 1.6924
R17261 GNDA.n4579 GNDA.n4505 1.6924
R17262 GNDA.n4579 GNDA.n4504 1.6924
R17263 GNDA.n3382 GNDA.n3317 1.6924
R17264 GNDA.n3382 GNDA.n3316 1.6924
R17265 GNDA.n3382 GNDA.n3314 1.6924
R17266 GNDA.n3382 GNDA.n3313 1.6924
R17267 GNDA.n3382 GNDA.n3311 1.6924
R17268 GNDA.n3382 GNDA.n3310 1.6924
R17269 GNDA.n3382 GNDA.n3308 1.6924
R17270 GNDA.n3382 GNDA.n3307 1.6924
R17271 GNDA.n3669 GNDA.n513 1.6924
R17272 GNDA.n3666 GNDA.n513 1.6924
R17273 GNDA.n3658 GNDA.n513 1.6924
R17274 GNDA.n3653 GNDA.n513 1.6924
R17275 GNDA.n3645 GNDA.n513 1.6924
R17276 GNDA.n3642 GNDA.n513 1.6924
R17277 GNDA.n3634 GNDA.n513 1.6924
R17278 GNDA.n3629 GNDA.n513 1.6924
R17279 GNDA.n2222 GNDA.n2127 1.6924
R17280 GNDA.n2222 GNDA.n2063 1.6924
R17281 GNDA.n2222 GNDA.n2061 1.6924
R17282 GNDA.n2222 GNDA.n2060 1.6924
R17283 GNDA.n2222 GNDA.n2058 1.6924
R17284 GNDA.n2222 GNDA.n2057 1.6924
R17285 GNDA.n2222 GNDA.n2055 1.6924
R17286 GNDA.n2222 GNDA.n2054 1.6924
R17287 GNDA.n2221 GNDA.n2139 1.6924
R17288 GNDA.n2221 GNDA.n2138 1.6924
R17289 GNDA.n2221 GNDA.n2136 1.6924
R17290 GNDA.n2221 GNDA.n2135 1.6924
R17291 GNDA.n2221 GNDA.n2133 1.6924
R17292 GNDA.n2221 GNDA.n2132 1.6924
R17293 GNDA.n2221 GNDA.n2130 1.6924
R17294 GNDA.n2221 GNDA.n2129 1.6924
R17295 GNDA.n1925 GNDA.n1140 1.6924
R17296 GNDA.n1925 GNDA.n1137 1.6924
R17297 GNDA.n1925 GNDA.n1134 1.6924
R17298 GNDA.n1925 GNDA.n1131 1.6924
R17299 GNDA.n1342 GNDA.n1272 1.56997
R17300 GNDA.n1339 GNDA.n1274 1.56997
R17301 GNDA.t246 GNDA.n105 1.51652
R17302 GNDA.n1738 GNDA.n1737 1.5005
R17303 GNDA.n3947 GNDA.n3946 1.5005
R17304 GNDA.n3042 GNDA.n3041 1.47392
R17305 GNDA.n2743 GNDA.n2742 1.47392
R17306 GNDA.n4870 GNDA.n228 1.47392
R17307 GNDA.n4847 GNDA.n4844 1.47392
R17308 GNDA.n2519 GNDA.n2518 1.47392
R17309 GNDA.n5093 GNDA.n87 1.47392
R17310 GNDA.n3710 GNDA.n543 1.27133
R17311 GNDA.n3389 GNDA.n586 1.27133
R17312 GNDA.n2209 GNDA.n2208 1.22446
R17313 GNDA.n1303 GNDA.n1299 1.07342
R17314 GNDA.n1384 GNDA.n1382 1.06821
R17315 GNDA.n1343 GNDA.n1342 1.063
R17316 GNDA.n1339 GNDA.n1338 1.063
R17317 GNDA.n2243 GNDA.n2239 1.05258
R17318 GNDA.n2211 GNDA.n2210 0.854667
R17319 GNDA.n3002 GNDA.n3001 0.8197
R17320 GNDA.n2988 GNDA.n746 0.8197
R17321 GNDA.n2995 GNDA.n2989 0.8197
R17322 GNDA.n2994 GNDA.n2991 0.8197
R17323 GNDA.n3007 GNDA.n714 0.8197
R17324 GNDA.n725 GNDA.n721 0.8197
R17325 GNDA.n727 GNDA.n726 0.8197
R17326 GNDA.n3045 GNDA.n689 0.8197
R17327 GNDA.n3079 GNDA.n3078 0.8197
R17328 GNDA.n3065 GNDA.n672 0.8197
R17329 GNDA.n3072 GNDA.n3066 0.8197
R17330 GNDA.n3071 GNDA.n3068 0.8197
R17331 GNDA.n3084 GNDA.n650 0.8197
R17332 GNDA.n2310 GNDA.n2305 0.8197
R17333 GNDA.n2313 GNDA.n2312 0.8197
R17334 GNDA.n2381 GNDA.n2314 0.8197
R17335 GNDA.n5051 GNDA.n165 0.8197
R17336 GNDA.n5050 GNDA.n167 0.8197
R17337 GNDA.n218 GNDA.n200 0.8197
R17338 GNDA.n217 GNDA.n215 0.8197
R17339 GNDA.n211 GNDA.n210 0.8197
R17340 GNDA.n207 GNDA.n203 0.8197
R17341 GNDA.n206 GNDA.n187 0.8197
R17342 GNDA.n4992 GNDA.n4991 0.8197
R17343 GNDA.n2727 GNDA.n2726 0.8197
R17344 GNDA.n2723 GNDA.n2722 0.8197
R17345 GNDA.n2719 GNDA.n2703 0.8197
R17346 GNDA.n2718 GNDA.n2715 0.8197
R17347 GNDA.n2711 GNDA.n2708 0.8197
R17348 GNDA.n2705 GNDA.n2627 0.8197
R17349 GNDA.n2733 GNDA.n2732 0.8197
R17350 GNDA.n2736 GNDA.n2626 0.8197
R17351 GNDA.n4982 GNDA.n4873 0.8197
R17352 GNDA.n4979 GNDA.n4978 0.8197
R17353 GNDA.n4975 GNDA.n4876 0.8197
R17354 GNDA.n4974 GNDA.n4877 0.8197
R17355 GNDA.n4909 GNDA.n4906 0.8197
R17356 GNDA.n4910 GNDA.n4900 0.8197
R17357 GNDA.n4914 GNDA.n4913 0.8197
R17358 GNDA.n4918 GNDA.n4917 0.8197
R17359 GNDA.n5261 GNDA.n59 0.8197
R17360 GNDA.n5258 GNDA.n5257 0.8197
R17361 GNDA.n5254 GNDA.n62 0.8197
R17362 GNDA.n5253 GNDA.n63 0.8197
R17363 GNDA.n5188 GNDA.n5185 0.8197
R17364 GNDA.n5189 GNDA.n5179 0.8197
R17365 GNDA.n5193 GNDA.n5192 0.8197
R17366 GNDA.n5197 GNDA.n5196 0.8197
R17367 GNDA.n4836 GNDA.n4728 0.8197
R17368 GNDA.n4835 GNDA.n4729 0.8197
R17369 GNDA.n4755 GNDA.n4752 0.8197
R17370 GNDA.n4758 GNDA.n4757 0.8197
R17371 GNDA.n4768 GNDA.n4765 0.8197
R17372 GNDA.n4769 GNDA.n4751 0.8197
R17373 GNDA.n4773 GNDA.n4772 0.8197
R17374 GNDA.n4777 GNDA.n4776 0.8197
R17375 GNDA.n2491 GNDA.n2490 0.8197
R17376 GNDA.n2497 GNDA.n2251 0.8197
R17377 GNDA.n2496 GNDA.n2252 0.8197
R17378 GNDA.n2414 GNDA.n2412 0.8197
R17379 GNDA.n2423 GNDA.n2421 0.8197
R17380 GNDA.n2422 GNDA.n2272 0.8197
R17381 GNDA.n2432 GNDA.n2431 0.8197
R17382 GNDA.n2274 GNDA.n2270 0.8197
R17383 GNDA.n5271 GNDA.n5270 0.8197
R17384 GNDA.n32 GNDA.n23 0.8197
R17385 GNDA.n39 GNDA.n33 0.8197
R17386 GNDA.n38 GNDA.n35 0.8197
R17387 GNDA.n5276 GNDA.n1 0.8197
R17388 GNDA.n5108 GNDA.n5105 0.8197
R17389 GNDA.n5111 GNDA.n5110 0.8197
R17390 GNDA.n5115 GNDA.n5114 0.8197
R17391 GNDA.n1306 GNDA.n1304 0.786958
R17392 GNDA.n1377 GNDA.n1376 0.786958
R17393 GNDA.n3149 GNDA.n3148 0.78175
R17394 GNDA.n4626 GNDA.n435 0.78175
R17395 GNDA.n3707 GNDA.n3706 0.776542
R17396 GNDA.n3386 GNDA.n3385 0.776542
R17397 GNDA.n4583 GNDA.n4582 0.776542
R17398 GNDA.n4446 GNDA.n469 0.776542
R17399 GNDA.n4364 GNDA.n464 0.776542
R17400 GNDA.n4282 GNDA.n459 0.776542
R17401 GNDA.n4200 GNDA.n454 0.776542
R17402 GNDA.n4118 GNDA.n445 0.776542
R17403 GNDA.n4036 GNDA.n440 0.776542
R17404 GNDA.n3854 GNDA.n3853 0.776542
R17405 GNDA.n3717 GNDA.n3716 0.776542
R17406 GNDA.n3620 GNDA.n3619 0.776542
R17407 GNDA.n3483 GNDA.n3482 0.776542
R17408 GNDA.n3473 GNDA.n3472 0.776542
R17409 GNDA.n3249 GNDA.n3248 0.776542
R17410 GNDA.n3239 GNDA.n3238 0.776542
R17411 GNDA.n1435 GNDA.n1393 0.776542
R17412 GNDA.n1250 GNDA.n1249 0.776542
R17413 GNDA.n1867 GNDA.n1866 0.776542
R17414 GNDA.n1860 GNDA.n1840 0.776542
R17415 GNDA.n2395 GNDA.n2394 0.776542
R17416 GNDA.n1517 GNDA.n1398 0.776542
R17417 GNDA.n3954 GNDA.n3953 0.77295
R17418 GNDA.n1599 GNDA.n1404 0.77295
R17419 GNDA.n3944 GNDA.n3943 0.755708
R17420 GNDA.n1736 GNDA.n1735 0.755708
R17421 GNDA.n3944 GNDA.n3862 0.751
R17422 GNDA.n1736 GNDA.n624 0.751
R17423 GNDA.n1255 GNDA.n626 0.729667
R17424 GNDA.n3148 GNDA.n627 0.729667
R17425 GNDA.n3131 GNDA.n435 0.729667
R17426 GNDA.n4625 GNDA.n436 0.729667
R17427 GNDA.n2222 GNDA.n2052 0.723198
R17428 GNDA.n2228 GNDA.n2227 0.71925
R17429 GNDA.n3142 GNDA.n3141 0.688
R17430 GNDA.n1322 GNDA.n629 0.688
R17431 GNDA.n3149 GNDA.n626 0.688
R17432 GNDA.n4626 GNDA.n4625 0.688
R17433 GNDA.n1926 GNDA.n1925 0.675611
R17434 GNDA.n3024 GNDA.n703 0.65675
R17435 GNDA.n2990 GNDA 0.5637
R17436 GNDA.n3067 GNDA 0.5637
R17437 GNDA.n214 GNDA 0.5637
R17438 GNDA GNDA.n2704 0.5637
R17439 GNDA GNDA.n4901 0.5637
R17440 GNDA GNDA.n5180 0.5637
R17441 GNDA.n4762 GNDA 0.5637
R17442 GNDA.n2416 GNDA 0.5637
R17443 GNDA.n34 GNDA 0.5637
R17444 GNDA.n1317 GNDA.n1316 0.464042
R17445 GNDA.n1366 GNDA.n1364 0.464042
R17446 GNDA.t26 GNDA.t25 0.396629
R17447 GNDA.n3141 GNDA.n629 0.396333
R17448 GNDA.n4867 GNDA.n105 0.383687
R17449 GNDA.n1330 GNDA.n1328 0.34425
R17450 GNDA.n1355 GNDA.n1354 0.34425
R17451 GNDA.n3104 GNDA.n3102 0.34425
R17452 GNDA.n3106 GNDA.n3104 0.34425
R17453 GNDA.n3108 GNDA.n3106 0.34425
R17454 GNDA.n3110 GNDA.n3108 0.34425
R17455 GNDA.n3112 GNDA.n3110 0.34425
R17456 GNDA.n3114 GNDA.n3112 0.34425
R17457 GNDA.n3116 GNDA.n3114 0.34425
R17458 GNDA.n3118 GNDA.n3116 0.34425
R17459 GNDA.n3120 GNDA.n3118 0.34425
R17460 GNDA.n3122 GNDA.n3120 0.34425
R17461 GNDA.n3124 GNDA.n3122 0.34425
R17462 GNDA.n2210 GNDA.n2209 0.339042
R17463 GNDA.n3131 GNDA.n627 0.313
R17464 GNDA.n3142 GNDA.n628 0.292167
R17465 GNDA.n1323 GNDA.n1322 0.292167
R17466 GNDA.n2048 GNDA.n2015 0.286759
R17467 GNDA.n1854 GNDA.n1851 0.28175
R17468 GNDA.n1859 GNDA.n1856 0.28175
R17469 GNDA.n1863 GNDA.n1861 0.28175
R17470 GNDA.n1767 GNDA.n1766 0.28175
R17471 GNDA.n1739 GNDA.n1738 0.28175
R17472 GNDA.n3245 GNDA.n3243 0.28175
R17473 GNDA.n3388 GNDA.n588 0.28175
R17474 GNDA.n3475 GNDA.n3390 0.28175
R17475 GNDA.n3479 GNDA.n3477 0.28175
R17476 GNDA.n3622 GNDA.n548 0.28175
R17477 GNDA.n3709 GNDA.n3624 0.28175
R17478 GNDA.n3713 GNDA.n3711 0.28175
R17479 GNDA.n3856 GNDA.n508 0.28175
R17480 GNDA.n3950 GNDA.n3947 0.28175
R17481 GNDA.n4614 GNDA.n4613 0.28175
R17482 GNDA.n4602 GNDA.n4601 0.28175
R17483 GNDA.n4598 GNDA.n4597 0.28175
R17484 GNDA.n4594 GNDA.n4593 0.28175
R17485 GNDA.n4590 GNDA.n4589 0.28175
R17486 GNDA.n1751 GNDA.n1750 0.271333
R17487 GNDA.n3008 GNDA 0.2565
R17488 GNDA.n3085 GNDA 0.2565
R17489 GNDA.n202 GNDA 0.2565
R17490 GNDA.n2712 GNDA 0.2565
R17491 GNDA.n4904 GNDA 0.2565
R17492 GNDA.n5183 GNDA 0.2565
R17493 GNDA GNDA.n4761 0.2565
R17494 GNDA GNDA.n2415 0.2565
R17495 GNDA GNDA.n0 0.2565
R17496 GNDA.n2012 GNDA.n1960 0.229919
R17497 GNDA.n3134 GNDA.n3133 0.208833
R17498 GNDA.n633 GNDA.n632 0.208833
R17499 GNDA.n1755 GNDA.n1754 0.198417
R17500 GNDA.n3241 GNDA.n3156 0.198417
R17501 GNDA.n3861 GNDA.n3858 0.198417
R17502 GNDA.n4618 GNDA.n4617 0.188
R17503 GNDA.n2297 GNDA.n2296 0.188
R17504 GNDA.n2392 GNDA.n2391 0.188
R17505 GNDA.n1325 GNDA.n1319 0.167167
R17506 GNDA.n1360 GNDA.n1359 0.167167
R17507 GNDA.n3059 GNDA.n676 0.15675
R17508 GNDA.n2510 GNDA.n2509 0.151542
R17509 GNDA.n3055 GNDA.n3054 0.151542
R17510 GNDA.n3030 GNDA.n3029 0.147453
R17511 GNDA.n3704 GNDA.n3703 0.146333
R17512 GNDA.n3703 GNDA.n3631 0.146333
R17513 GNDA.n3699 GNDA.n3631 0.146333
R17514 GNDA.n3693 GNDA.n3639 0.146333
R17515 GNDA.n3693 GNDA.n3692 0.146333
R17516 GNDA.n3692 GNDA.n3691 0.146333
R17517 GNDA.n3686 GNDA.n3685 0.146333
R17518 GNDA.n3685 GNDA.n3655 0.146333
R17519 GNDA.n3681 GNDA.n3655 0.146333
R17520 GNDA.n3675 GNDA.n3663 0.146333
R17521 GNDA.n3675 GNDA.n3674 0.146333
R17522 GNDA.n3674 GNDA.n3673 0.146333
R17523 GNDA.n3329 GNDA.n591 0.146333
R17524 GNDA.n3334 GNDA.n3329 0.146333
R17525 GNDA.n3335 GNDA.n3334 0.146333
R17526 GNDA.n3345 GNDA.n3344 0.146333
R17527 GNDA.n3348 GNDA.n3345 0.146333
R17528 GNDA.n3348 GNDA.n3325 0.146333
R17529 GNDA.n3358 GNDA.n3323 0.146333
R17530 GNDA.n3364 GNDA.n3323 0.146333
R17531 GNDA.n3365 GNDA.n3364 0.146333
R17532 GNDA.n3375 GNDA.n3374 0.146333
R17533 GNDA.n3378 GNDA.n3375 0.146333
R17534 GNDA.n3378 GNDA.n3319 0.146333
R17535 GNDA.n4526 GNDA.n475 0.146333
R17536 GNDA.n4531 GNDA.n4526 0.146333
R17537 GNDA.n4532 GNDA.n4531 0.146333
R17538 GNDA.n4542 GNDA.n4541 0.146333
R17539 GNDA.n4545 GNDA.n4542 0.146333
R17540 GNDA.n4545 GNDA.n4522 0.146333
R17541 GNDA.n4555 GNDA.n4520 0.146333
R17542 GNDA.n4561 GNDA.n4520 0.146333
R17543 GNDA.n4562 GNDA.n4561 0.146333
R17544 GNDA.n4572 GNDA.n4571 0.146333
R17545 GNDA.n4575 GNDA.n4572 0.146333
R17546 GNDA.n4575 GNDA.n4516 0.146333
R17547 GNDA.n4449 GNDA.n4445 0.146333
R17548 GNDA.n4455 GNDA.n4445 0.146333
R17549 GNDA.n4456 GNDA.n4455 0.146333
R17550 GNDA.n4466 GNDA.n4465 0.146333
R17551 GNDA.n4469 GNDA.n4466 0.146333
R17552 GNDA.n4469 GNDA.n4441 0.146333
R17553 GNDA.n4479 GNDA.n4439 0.146333
R17554 GNDA.n4485 GNDA.n4439 0.146333
R17555 GNDA.n4486 GNDA.n4485 0.146333
R17556 GNDA.n4496 GNDA.n4495 0.146333
R17557 GNDA.n4499 GNDA.n4496 0.146333
R17558 GNDA.n4499 GNDA.n4435 0.146333
R17559 GNDA.n4367 GNDA.n4363 0.146333
R17560 GNDA.n4373 GNDA.n4363 0.146333
R17561 GNDA.n4374 GNDA.n4373 0.146333
R17562 GNDA.n4384 GNDA.n4383 0.146333
R17563 GNDA.n4387 GNDA.n4384 0.146333
R17564 GNDA.n4387 GNDA.n4359 0.146333
R17565 GNDA.n4397 GNDA.n4357 0.146333
R17566 GNDA.n4403 GNDA.n4357 0.146333
R17567 GNDA.n4404 GNDA.n4403 0.146333
R17568 GNDA.n4414 GNDA.n4413 0.146333
R17569 GNDA.n4417 GNDA.n4414 0.146333
R17570 GNDA.n4417 GNDA.n4353 0.146333
R17571 GNDA.n4285 GNDA.n4281 0.146333
R17572 GNDA.n4291 GNDA.n4281 0.146333
R17573 GNDA.n4292 GNDA.n4291 0.146333
R17574 GNDA.n4302 GNDA.n4301 0.146333
R17575 GNDA.n4305 GNDA.n4302 0.146333
R17576 GNDA.n4305 GNDA.n4277 0.146333
R17577 GNDA.n4315 GNDA.n4275 0.146333
R17578 GNDA.n4321 GNDA.n4275 0.146333
R17579 GNDA.n4322 GNDA.n4321 0.146333
R17580 GNDA.n4332 GNDA.n4331 0.146333
R17581 GNDA.n4335 GNDA.n4332 0.146333
R17582 GNDA.n4335 GNDA.n4271 0.146333
R17583 GNDA.n4203 GNDA.n4199 0.146333
R17584 GNDA.n4209 GNDA.n4199 0.146333
R17585 GNDA.n4210 GNDA.n4209 0.146333
R17586 GNDA.n4220 GNDA.n4219 0.146333
R17587 GNDA.n4223 GNDA.n4220 0.146333
R17588 GNDA.n4223 GNDA.n4195 0.146333
R17589 GNDA.n4233 GNDA.n4193 0.146333
R17590 GNDA.n4239 GNDA.n4193 0.146333
R17591 GNDA.n4240 GNDA.n4239 0.146333
R17592 GNDA.n4250 GNDA.n4249 0.146333
R17593 GNDA.n4253 GNDA.n4250 0.146333
R17594 GNDA.n4253 GNDA.n4189 0.146333
R17595 GNDA.n3957 GNDA.n501 0.146333
R17596 GNDA.n3963 GNDA.n501 0.146333
R17597 GNDA.n3964 GNDA.n3963 0.146333
R17598 GNDA.n3974 GNDA.n3973 0.146333
R17599 GNDA.n3977 GNDA.n3974 0.146333
R17600 GNDA.n3977 GNDA.n497 0.146333
R17601 GNDA.n3987 GNDA.n495 0.146333
R17602 GNDA.n3993 GNDA.n495 0.146333
R17603 GNDA.n3994 GNDA.n3993 0.146333
R17604 GNDA.n4004 GNDA.n4003 0.146333
R17605 GNDA.n4007 GNDA.n4004 0.146333
R17606 GNDA.n4007 GNDA.n491 0.146333
R17607 GNDA.n4121 GNDA.n4117 0.146333
R17608 GNDA.n4127 GNDA.n4117 0.146333
R17609 GNDA.n4128 GNDA.n4127 0.146333
R17610 GNDA.n4138 GNDA.n4137 0.146333
R17611 GNDA.n4141 GNDA.n4138 0.146333
R17612 GNDA.n4141 GNDA.n4113 0.146333
R17613 GNDA.n4151 GNDA.n4111 0.146333
R17614 GNDA.n4157 GNDA.n4111 0.146333
R17615 GNDA.n4158 GNDA.n4157 0.146333
R17616 GNDA.n4168 GNDA.n4167 0.146333
R17617 GNDA.n4171 GNDA.n4168 0.146333
R17618 GNDA.n4171 GNDA.n4107 0.146333
R17619 GNDA.n4039 GNDA.n4035 0.146333
R17620 GNDA.n4045 GNDA.n4035 0.146333
R17621 GNDA.n4046 GNDA.n4045 0.146333
R17622 GNDA.n4056 GNDA.n4055 0.146333
R17623 GNDA.n4059 GNDA.n4056 0.146333
R17624 GNDA.n4059 GNDA.n4031 0.146333
R17625 GNDA.n4069 GNDA.n4029 0.146333
R17626 GNDA.n4075 GNDA.n4029 0.146333
R17627 GNDA.n4076 GNDA.n4075 0.146333
R17628 GNDA.n4086 GNDA.n4085 0.146333
R17629 GNDA.n4089 GNDA.n4086 0.146333
R17630 GNDA.n4089 GNDA.n4025 0.146333
R17631 GNDA.n3865 GNDA.n3864 0.146333
R17632 GNDA.n3866 GNDA.n3865 0.146333
R17633 GNDA.n3867 GNDA.n3866 0.146333
R17634 GNDA.n3871 GNDA.n3870 0.146333
R17635 GNDA.n3872 GNDA.n3871 0.146333
R17636 GNDA.n3873 GNDA.n3872 0.146333
R17637 GNDA.n3877 GNDA.n3876 0.146333
R17638 GNDA.n3878 GNDA.n3877 0.146333
R17639 GNDA.n3879 GNDA.n3878 0.146333
R17640 GNDA.n3883 GNDA.n3882 0.146333
R17641 GNDA.n3884 GNDA.n3883 0.146333
R17642 GNDA.n3885 GNDA.n3884 0.146333
R17643 GNDA.n1679 GNDA.n1409 0.146333
R17644 GNDA.n1684 GNDA.n1679 0.146333
R17645 GNDA.n1685 GNDA.n1684 0.146333
R17646 GNDA.n1695 GNDA.n1694 0.146333
R17647 GNDA.n1698 GNDA.n1695 0.146333
R17648 GNDA.n1698 GNDA.n1675 0.146333
R17649 GNDA.n1708 GNDA.n1673 0.146333
R17650 GNDA.n1714 GNDA.n1673 0.146333
R17651 GNDA.n1715 GNDA.n1714 0.146333
R17652 GNDA.n1725 GNDA.n1724 0.146333
R17653 GNDA.n1728 GNDA.n1725 0.146333
R17654 GNDA.n1728 GNDA.n1669 0.146333
R17655 GNDA.n3797 GNDA.n511 0.146333
R17656 GNDA.n3802 GNDA.n3797 0.146333
R17657 GNDA.n3803 GNDA.n3802 0.146333
R17658 GNDA.n3813 GNDA.n3812 0.146333
R17659 GNDA.n3816 GNDA.n3813 0.146333
R17660 GNDA.n3816 GNDA.n3793 0.146333
R17661 GNDA.n3826 GNDA.n3791 0.146333
R17662 GNDA.n3832 GNDA.n3791 0.146333
R17663 GNDA.n3833 GNDA.n3832 0.146333
R17664 GNDA.n3843 GNDA.n3842 0.146333
R17665 GNDA.n3846 GNDA.n3843 0.146333
R17666 GNDA.n3846 GNDA.n3787 0.146333
R17667 GNDA.n3720 GNDA.n537 0.146333
R17668 GNDA.n3726 GNDA.n537 0.146333
R17669 GNDA.n3727 GNDA.n3726 0.146333
R17670 GNDA.n3737 GNDA.n3736 0.146333
R17671 GNDA.n3740 GNDA.n3737 0.146333
R17672 GNDA.n3740 GNDA.n533 0.146333
R17673 GNDA.n3750 GNDA.n531 0.146333
R17674 GNDA.n3756 GNDA.n531 0.146333
R17675 GNDA.n3757 GNDA.n3756 0.146333
R17676 GNDA.n3767 GNDA.n3766 0.146333
R17677 GNDA.n3770 GNDA.n3767 0.146333
R17678 GNDA.n3770 GNDA.n527 0.146333
R17679 GNDA.n3563 GNDA.n551 0.146333
R17680 GNDA.n3568 GNDA.n3563 0.146333
R17681 GNDA.n3569 GNDA.n3568 0.146333
R17682 GNDA.n3579 GNDA.n3578 0.146333
R17683 GNDA.n3582 GNDA.n3579 0.146333
R17684 GNDA.n3582 GNDA.n3559 0.146333
R17685 GNDA.n3592 GNDA.n3557 0.146333
R17686 GNDA.n3598 GNDA.n3557 0.146333
R17687 GNDA.n3599 GNDA.n3598 0.146333
R17688 GNDA.n3609 GNDA.n3608 0.146333
R17689 GNDA.n3612 GNDA.n3609 0.146333
R17690 GNDA.n3612 GNDA.n3553 0.146333
R17691 GNDA.n3486 GNDA.n577 0.146333
R17692 GNDA.n3492 GNDA.n577 0.146333
R17693 GNDA.n3493 GNDA.n3492 0.146333
R17694 GNDA.n3503 GNDA.n3502 0.146333
R17695 GNDA.n3506 GNDA.n3503 0.146333
R17696 GNDA.n3506 GNDA.n573 0.146333
R17697 GNDA.n3516 GNDA.n571 0.146333
R17698 GNDA.n3522 GNDA.n571 0.146333
R17699 GNDA.n3523 GNDA.n3522 0.146333
R17700 GNDA.n3533 GNDA.n3532 0.146333
R17701 GNDA.n3536 GNDA.n3533 0.146333
R17702 GNDA.n3536 GNDA.n567 0.146333
R17703 GNDA.n3394 GNDA.n3393 0.146333
R17704 GNDA.n3395 GNDA.n3394 0.146333
R17705 GNDA.n3396 GNDA.n3395 0.146333
R17706 GNDA.n3400 GNDA.n3399 0.146333
R17707 GNDA.n3401 GNDA.n3400 0.146333
R17708 GNDA.n3402 GNDA.n3401 0.146333
R17709 GNDA.n3406 GNDA.n3405 0.146333
R17710 GNDA.n3407 GNDA.n3406 0.146333
R17711 GNDA.n3408 GNDA.n3407 0.146333
R17712 GNDA.n3412 GNDA.n3411 0.146333
R17713 GNDA.n3413 GNDA.n3412 0.146333
R17714 GNDA.n3414 GNDA.n3413 0.146333
R17715 GNDA.n3252 GNDA.n617 0.146333
R17716 GNDA.n3258 GNDA.n617 0.146333
R17717 GNDA.n3259 GNDA.n3258 0.146333
R17718 GNDA.n3269 GNDA.n3268 0.146333
R17719 GNDA.n3272 GNDA.n3269 0.146333
R17720 GNDA.n3272 GNDA.n613 0.146333
R17721 GNDA.n3282 GNDA.n611 0.146333
R17722 GNDA.n3288 GNDA.n611 0.146333
R17723 GNDA.n3289 GNDA.n3288 0.146333
R17724 GNDA.n3299 GNDA.n3298 0.146333
R17725 GNDA.n3302 GNDA.n3299 0.146333
R17726 GNDA.n3302 GNDA.n607 0.146333
R17727 GNDA.n3160 GNDA.n3159 0.146333
R17728 GNDA.n3161 GNDA.n3160 0.146333
R17729 GNDA.n3162 GNDA.n3161 0.146333
R17730 GNDA.n3166 GNDA.n3165 0.146333
R17731 GNDA.n3167 GNDA.n3166 0.146333
R17732 GNDA.n3168 GNDA.n3167 0.146333
R17733 GNDA.n3172 GNDA.n3171 0.146333
R17734 GNDA.n3173 GNDA.n3172 0.146333
R17735 GNDA.n3174 GNDA.n3173 0.146333
R17736 GNDA.n3178 GNDA.n3177 0.146333
R17737 GNDA.n3179 GNDA.n3178 0.146333
R17738 GNDA.n3180 GNDA.n3179 0.146333
R17739 GNDA.n1602 GNDA.n1598 0.146333
R17740 GNDA.n1608 GNDA.n1598 0.146333
R17741 GNDA.n1609 GNDA.n1608 0.146333
R17742 GNDA.n1619 GNDA.n1618 0.146333
R17743 GNDA.n1622 GNDA.n1619 0.146333
R17744 GNDA.n1622 GNDA.n1594 0.146333
R17745 GNDA.n1632 GNDA.n1592 0.146333
R17746 GNDA.n1638 GNDA.n1592 0.146333
R17747 GNDA.n1639 GNDA.n1638 0.146333
R17748 GNDA.n1649 GNDA.n1648 0.146333
R17749 GNDA.n1652 GNDA.n1649 0.146333
R17750 GNDA.n1652 GNDA.n1588 0.146333
R17751 GNDA.n1520 GNDA.n1516 0.146333
R17752 GNDA.n1526 GNDA.n1516 0.146333
R17753 GNDA.n1527 GNDA.n1526 0.146333
R17754 GNDA.n1537 GNDA.n1536 0.146333
R17755 GNDA.n1540 GNDA.n1537 0.146333
R17756 GNDA.n1540 GNDA.n1512 0.146333
R17757 GNDA.n1550 GNDA.n1510 0.146333
R17758 GNDA.n1556 GNDA.n1510 0.146333
R17759 GNDA.n1557 GNDA.n1556 0.146333
R17760 GNDA.n1567 GNDA.n1566 0.146333
R17761 GNDA.n1570 GNDA.n1567 0.146333
R17762 GNDA.n1570 GNDA.n1506 0.146333
R17763 GNDA.n1438 GNDA.n1434 0.146333
R17764 GNDA.n1444 GNDA.n1434 0.146333
R17765 GNDA.n1445 GNDA.n1444 0.146333
R17766 GNDA.n1455 GNDA.n1454 0.146333
R17767 GNDA.n1458 GNDA.n1455 0.146333
R17768 GNDA.n1458 GNDA.n1430 0.146333
R17769 GNDA.n1468 GNDA.n1428 0.146333
R17770 GNDA.n1474 GNDA.n1428 0.146333
R17771 GNDA.n1475 GNDA.n1474 0.146333
R17772 GNDA.n1485 GNDA.n1484 0.146333
R17773 GNDA.n1488 GNDA.n1485 0.146333
R17774 GNDA.n1488 GNDA.n1424 0.146333
R17775 GNDA.n1171 GNDA.n1170 0.146333
R17776 GNDA.n1172 GNDA.n1171 0.146333
R17777 GNDA.n1173 GNDA.n1172 0.146333
R17778 GNDA.n1177 GNDA.n1176 0.146333
R17779 GNDA.n1178 GNDA.n1177 0.146333
R17780 GNDA.n1179 GNDA.n1178 0.146333
R17781 GNDA.n1183 GNDA.n1182 0.146333
R17782 GNDA.n1184 GNDA.n1183 0.146333
R17783 GNDA.n1185 GNDA.n1184 0.146333
R17784 GNDA.n1189 GNDA.n1188 0.146333
R17785 GNDA.n1190 GNDA.n1189 0.146333
R17786 GNDA.n1191 GNDA.n1190 0.146333
R17787 GNDA.n1870 GNDA.n1165 0.146333
R17788 GNDA.n1876 GNDA.n1165 0.146333
R17789 GNDA.n1877 GNDA.n1876 0.146333
R17790 GNDA.n1887 GNDA.n1886 0.146333
R17791 GNDA.n1890 GNDA.n1887 0.146333
R17792 GNDA.n1890 GNDA.n1161 0.146333
R17793 GNDA.n1900 GNDA.n1159 0.146333
R17794 GNDA.n1906 GNDA.n1159 0.146333
R17795 GNDA.n1907 GNDA.n1906 0.146333
R17796 GNDA.n1917 GNDA.n1916 0.146333
R17797 GNDA.n1920 GNDA.n1917 0.146333
R17798 GNDA.n1920 GNDA.n1155 0.146333
R17799 GNDA.n1838 GNDA.n1837 0.146333
R17800 GNDA.n1837 GNDA.n1776 0.146333
R17801 GNDA.n1833 GNDA.n1776 0.146333
R17802 GNDA.n1827 GNDA.n1782 0.146333
R17803 GNDA.n1827 GNDA.n1826 0.146333
R17804 GNDA.n1826 GNDA.n1825 0.146333
R17805 GNDA.n1820 GNDA.n1819 0.146333
R17806 GNDA.n1819 GNDA.n1794 0.146333
R17807 GNDA.n1815 GNDA.n1794 0.146333
R17808 GNDA.n1809 GNDA.n1800 0.146333
R17809 GNDA.n1809 GNDA.n1808 0.146333
R17810 GNDA.n1808 GNDA.n1807 0.146333
R17811 GNDA.n2163 GNDA.n2159 0.146333
R17812 GNDA.n2167 GNDA.n2159 0.146333
R17813 GNDA.n2168 GNDA.n2167 0.146333
R17814 GNDA.n2176 GNDA.n2175 0.146333
R17815 GNDA.n2179 GNDA.n2176 0.146333
R17816 GNDA.n2179 GNDA.n2151 0.146333
R17817 GNDA.n2187 GNDA.n2147 0.146333
R17818 GNDA.n2191 GNDA.n2147 0.146333
R17819 GNDA.n2192 GNDA.n2191 0.146333
R17820 GNDA.n2200 GNDA.n2199 0.146333
R17821 GNDA.n2203 GNDA.n2200 0.146333
R17822 GNDA.n2203 GNDA.n2141 0.146333
R17823 GNDA.n2082 GNDA.n2074 0.146333
R17824 GNDA.n2083 GNDA.n2082 0.146333
R17825 GNDA.n2093 GNDA.n2092 0.146333
R17826 GNDA.n2094 GNDA.n2093 0.146333
R17827 GNDA.n2094 GNDA.n2070 0.146333
R17828 GNDA.n2104 GNDA.n2068 0.146333
R17829 GNDA.n2112 GNDA.n2068 0.146333
R17830 GNDA.n2113 GNDA.n2112 0.146333
R17831 GNDA.n2123 GNDA.n2122 0.146333
R17832 GNDA.n2124 GNDA.n2123 0.146333
R17833 GNDA.n2124 GNDA.n843 0.146333
R17834 GNDA.n2078 GNDA.n2077 0.146333
R17835 GNDA.n2081 GNDA.n2078 0.146333
R17836 GNDA.n2081 GNDA.n2073 0.146333
R17837 GNDA.n2091 GNDA.n2071 0.146333
R17838 GNDA.n2097 GNDA.n2071 0.146333
R17839 GNDA.n2098 GNDA.n2097 0.146333
R17840 GNDA.n2108 GNDA.n2107 0.146333
R17841 GNDA.n2111 GNDA.n2108 0.146333
R17842 GNDA.n2111 GNDA.n2067 0.146333
R17843 GNDA.n2121 GNDA.n2065 0.146333
R17844 GNDA.n2125 GNDA.n2065 0.146333
R17845 GNDA.n2125 GNDA.n844 0.146333
R17846 GNDA.n3705 GNDA.n3704 0.135917
R17847 GNDA.n3699 GNDA.n3698 0.135917
R17848 GNDA.n3697 GNDA.n3639 0.135917
R17849 GNDA.n3691 GNDA.n3647 0.135917
R17850 GNDA.n3687 GNDA.n3686 0.135917
R17851 GNDA.n3681 GNDA.n3680 0.135917
R17852 GNDA.n3679 GNDA.n3663 0.135917
R17853 GNDA.n3384 GNDA.n591 0.135917
R17854 GNDA.n3338 GNDA.n3335 0.135917
R17855 GNDA.n3344 GNDA.n3327 0.135917
R17856 GNDA.n3354 GNDA.n3325 0.135917
R17857 GNDA.n3358 GNDA.n3355 0.135917
R17858 GNDA.n3368 GNDA.n3365 0.135917
R17859 GNDA.n3374 GNDA.n3321 0.135917
R17860 GNDA.n4581 GNDA.n475 0.135917
R17861 GNDA.n4535 GNDA.n4532 0.135917
R17862 GNDA.n4541 GNDA.n4524 0.135917
R17863 GNDA.n4551 GNDA.n4522 0.135917
R17864 GNDA.n4555 GNDA.n4552 0.135917
R17865 GNDA.n4565 GNDA.n4562 0.135917
R17866 GNDA.n4571 GNDA.n4518 0.135917
R17867 GNDA.n4449 GNDA.n4447 0.135917
R17868 GNDA.n4459 GNDA.n4456 0.135917
R17869 GNDA.n4465 GNDA.n4443 0.135917
R17870 GNDA.n4475 GNDA.n4441 0.135917
R17871 GNDA.n4479 GNDA.n4476 0.135917
R17872 GNDA.n4489 GNDA.n4486 0.135917
R17873 GNDA.n4495 GNDA.n4437 0.135917
R17874 GNDA.n4367 GNDA.n4365 0.135917
R17875 GNDA.n4377 GNDA.n4374 0.135917
R17876 GNDA.n4383 GNDA.n4361 0.135917
R17877 GNDA.n4393 GNDA.n4359 0.135917
R17878 GNDA.n4397 GNDA.n4394 0.135917
R17879 GNDA.n4407 GNDA.n4404 0.135917
R17880 GNDA.n4413 GNDA.n4355 0.135917
R17881 GNDA.n4285 GNDA.n4283 0.135917
R17882 GNDA.n4295 GNDA.n4292 0.135917
R17883 GNDA.n4301 GNDA.n4279 0.135917
R17884 GNDA.n4311 GNDA.n4277 0.135917
R17885 GNDA.n4315 GNDA.n4312 0.135917
R17886 GNDA.n4325 GNDA.n4322 0.135917
R17887 GNDA.n4331 GNDA.n4273 0.135917
R17888 GNDA.n4203 GNDA.n4201 0.135917
R17889 GNDA.n4213 GNDA.n4210 0.135917
R17890 GNDA.n4219 GNDA.n4197 0.135917
R17891 GNDA.n4229 GNDA.n4195 0.135917
R17892 GNDA.n4233 GNDA.n4230 0.135917
R17893 GNDA.n4243 GNDA.n4240 0.135917
R17894 GNDA.n4249 GNDA.n4191 0.135917
R17895 GNDA.n3957 GNDA.n3955 0.135917
R17896 GNDA.n3967 GNDA.n3964 0.135917
R17897 GNDA.n3973 GNDA.n499 0.135917
R17898 GNDA.n3983 GNDA.n497 0.135917
R17899 GNDA.n3987 GNDA.n3984 0.135917
R17900 GNDA.n3997 GNDA.n3994 0.135917
R17901 GNDA.n4003 GNDA.n493 0.135917
R17902 GNDA.n4121 GNDA.n4119 0.135917
R17903 GNDA.n4131 GNDA.n4128 0.135917
R17904 GNDA.n4137 GNDA.n4115 0.135917
R17905 GNDA.n4147 GNDA.n4113 0.135917
R17906 GNDA.n4151 GNDA.n4148 0.135917
R17907 GNDA.n4161 GNDA.n4158 0.135917
R17908 GNDA.n4167 GNDA.n4109 0.135917
R17909 GNDA.n4039 GNDA.n4037 0.135917
R17910 GNDA.n4049 GNDA.n4046 0.135917
R17911 GNDA.n4055 GNDA.n4033 0.135917
R17912 GNDA.n4065 GNDA.n4031 0.135917
R17913 GNDA.n4069 GNDA.n4066 0.135917
R17914 GNDA.n4079 GNDA.n4076 0.135917
R17915 GNDA.n4085 GNDA.n4027 0.135917
R17916 GNDA.n3942 GNDA.n3864 0.135917
R17917 GNDA.n3868 GNDA.n3867 0.135917
R17918 GNDA.n3870 GNDA.n3869 0.135917
R17919 GNDA.n3874 GNDA.n3873 0.135917
R17920 GNDA.n3876 GNDA.n3875 0.135917
R17921 GNDA.n3880 GNDA.n3879 0.135917
R17922 GNDA.n3882 GNDA.n3881 0.135917
R17923 GNDA.n1734 GNDA.n1409 0.135917
R17924 GNDA.n1688 GNDA.n1685 0.135917
R17925 GNDA.n1694 GNDA.n1677 0.135917
R17926 GNDA.n1704 GNDA.n1675 0.135917
R17927 GNDA.n1708 GNDA.n1705 0.135917
R17928 GNDA.n1718 GNDA.n1715 0.135917
R17929 GNDA.n1724 GNDA.n1671 0.135917
R17930 GNDA.n3852 GNDA.n511 0.135917
R17931 GNDA.n3806 GNDA.n3803 0.135917
R17932 GNDA.n3812 GNDA.n3795 0.135917
R17933 GNDA.n3822 GNDA.n3793 0.135917
R17934 GNDA.n3826 GNDA.n3823 0.135917
R17935 GNDA.n3836 GNDA.n3833 0.135917
R17936 GNDA.n3842 GNDA.n3789 0.135917
R17937 GNDA.n3720 GNDA.n3718 0.135917
R17938 GNDA.n3730 GNDA.n3727 0.135917
R17939 GNDA.n3736 GNDA.n535 0.135917
R17940 GNDA.n3746 GNDA.n533 0.135917
R17941 GNDA.n3750 GNDA.n3747 0.135917
R17942 GNDA.n3760 GNDA.n3757 0.135917
R17943 GNDA.n3766 GNDA.n529 0.135917
R17944 GNDA.n3618 GNDA.n551 0.135917
R17945 GNDA.n3572 GNDA.n3569 0.135917
R17946 GNDA.n3578 GNDA.n3561 0.135917
R17947 GNDA.n3588 GNDA.n3559 0.135917
R17948 GNDA.n3592 GNDA.n3589 0.135917
R17949 GNDA.n3602 GNDA.n3599 0.135917
R17950 GNDA.n3608 GNDA.n3555 0.135917
R17951 GNDA.n3486 GNDA.n3484 0.135917
R17952 GNDA.n3496 GNDA.n3493 0.135917
R17953 GNDA.n3502 GNDA.n575 0.135917
R17954 GNDA.n3512 GNDA.n573 0.135917
R17955 GNDA.n3516 GNDA.n3513 0.135917
R17956 GNDA.n3526 GNDA.n3523 0.135917
R17957 GNDA.n3532 GNDA.n569 0.135917
R17958 GNDA.n3471 GNDA.n3393 0.135917
R17959 GNDA.n3397 GNDA.n3396 0.135917
R17960 GNDA.n3399 GNDA.n3398 0.135917
R17961 GNDA.n3403 GNDA.n3402 0.135917
R17962 GNDA.n3405 GNDA.n3404 0.135917
R17963 GNDA.n3409 GNDA.n3408 0.135917
R17964 GNDA.n3411 GNDA.n3410 0.135917
R17965 GNDA.n3252 GNDA.n3250 0.135917
R17966 GNDA.n3262 GNDA.n3259 0.135917
R17967 GNDA.n3268 GNDA.n615 0.135917
R17968 GNDA.n3278 GNDA.n613 0.135917
R17969 GNDA.n3282 GNDA.n3279 0.135917
R17970 GNDA.n3292 GNDA.n3289 0.135917
R17971 GNDA.n3298 GNDA.n609 0.135917
R17972 GNDA.n3237 GNDA.n3159 0.135917
R17973 GNDA.n3163 GNDA.n3162 0.135917
R17974 GNDA.n3165 GNDA.n3164 0.135917
R17975 GNDA.n3169 GNDA.n3168 0.135917
R17976 GNDA.n3171 GNDA.n3170 0.135917
R17977 GNDA.n3175 GNDA.n3174 0.135917
R17978 GNDA.n3177 GNDA.n3176 0.135917
R17979 GNDA.n1602 GNDA.n1600 0.135917
R17980 GNDA.n1612 GNDA.n1609 0.135917
R17981 GNDA.n1618 GNDA.n1596 0.135917
R17982 GNDA.n1628 GNDA.n1594 0.135917
R17983 GNDA.n1632 GNDA.n1629 0.135917
R17984 GNDA.n1642 GNDA.n1639 0.135917
R17985 GNDA.n1648 GNDA.n1590 0.135917
R17986 GNDA.n1520 GNDA.n1518 0.135917
R17987 GNDA.n1530 GNDA.n1527 0.135917
R17988 GNDA.n1536 GNDA.n1514 0.135917
R17989 GNDA.n1546 GNDA.n1512 0.135917
R17990 GNDA.n1550 GNDA.n1547 0.135917
R17991 GNDA.n1560 GNDA.n1557 0.135917
R17992 GNDA.n1566 GNDA.n1508 0.135917
R17993 GNDA.n1438 GNDA.n1436 0.135917
R17994 GNDA.n1448 GNDA.n1445 0.135917
R17995 GNDA.n1454 GNDA.n1432 0.135917
R17996 GNDA.n1464 GNDA.n1430 0.135917
R17997 GNDA.n1468 GNDA.n1465 0.135917
R17998 GNDA.n1478 GNDA.n1475 0.135917
R17999 GNDA.n1484 GNDA.n1426 0.135917
R18000 GNDA.n1248 GNDA.n1170 0.135917
R18001 GNDA.n1174 GNDA.n1173 0.135917
R18002 GNDA.n1176 GNDA.n1175 0.135917
R18003 GNDA.n1180 GNDA.n1179 0.135917
R18004 GNDA.n1182 GNDA.n1181 0.135917
R18005 GNDA.n1186 GNDA.n1185 0.135917
R18006 GNDA.n1188 GNDA.n1187 0.135917
R18007 GNDA.n1870 GNDA.n1868 0.135917
R18008 GNDA.n1880 GNDA.n1877 0.135917
R18009 GNDA.n1886 GNDA.n1163 0.135917
R18010 GNDA.n1896 GNDA.n1161 0.135917
R18011 GNDA.n1900 GNDA.n1897 0.135917
R18012 GNDA.n1910 GNDA.n1907 0.135917
R18013 GNDA.n1916 GNDA.n1157 0.135917
R18014 GNDA.n1839 GNDA.n1838 0.135917
R18015 GNDA.n1833 GNDA.n1832 0.135917
R18016 GNDA.n1831 GNDA.n1782 0.135917
R18017 GNDA.n1825 GNDA.n1788 0.135917
R18018 GNDA.n1821 GNDA.n1820 0.135917
R18019 GNDA.n1815 GNDA.n1814 0.135917
R18020 GNDA.n1813 GNDA.n1800 0.135917
R18021 GNDA.n2171 GNDA.n2168 0.135917
R18022 GNDA.n2175 GNDA.n2155 0.135917
R18023 GNDA.n2183 GNDA.n2151 0.135917
R18024 GNDA.n2187 GNDA.n2184 0.135917
R18025 GNDA.n2195 GNDA.n2192 0.135917
R18026 GNDA.n2199 GNDA.n2143 0.135917
R18027 GNDA.n2219 GNDA.n2141 0.135917
R18028 GNDA.n2084 GNDA.n2083 0.135917
R18029 GNDA.n2092 GNDA.n2072 0.135917
R18030 GNDA.n2102 GNDA.n2070 0.135917
R18031 GNDA.n2104 GNDA.n2103 0.135917
R18032 GNDA.n2114 GNDA.n2113 0.135917
R18033 GNDA.n2122 GNDA.n2066 0.135917
R18034 GNDA.n2225 GNDA.n843 0.135917
R18035 GNDA.n2087 GNDA.n2073 0.135917
R18036 GNDA.n2091 GNDA.n2088 0.135917
R18037 GNDA.n2101 GNDA.n2098 0.135917
R18038 GNDA.n2107 GNDA.n2069 0.135917
R18039 GNDA.n2117 GNDA.n2067 0.135917
R18040 GNDA.n2121 GNDA.n2118 0.135917
R18041 GNDA.n2224 GNDA.n844 0.135917
R18042 GNDA.n2222 GNDA.n2221 0.135331
R18043 GNDA.n3698 GNDA.n3697 0.1255
R18044 GNDA.n3687 GNDA.n3647 0.1255
R18045 GNDA.n3680 GNDA.n3679 0.1255
R18046 GNDA.n3338 GNDA.n3327 0.1255
R18047 GNDA.n3355 GNDA.n3354 0.1255
R18048 GNDA.n3368 GNDA.n3321 0.1255
R18049 GNDA.n4535 GNDA.n4524 0.1255
R18050 GNDA.n4552 GNDA.n4551 0.1255
R18051 GNDA.n4565 GNDA.n4518 0.1255
R18052 GNDA.n4459 GNDA.n4443 0.1255
R18053 GNDA.n4476 GNDA.n4475 0.1255
R18054 GNDA.n4489 GNDA.n4437 0.1255
R18055 GNDA.n4377 GNDA.n4361 0.1255
R18056 GNDA.n4394 GNDA.n4393 0.1255
R18057 GNDA.n4407 GNDA.n4355 0.1255
R18058 GNDA.n4295 GNDA.n4279 0.1255
R18059 GNDA.n4312 GNDA.n4311 0.1255
R18060 GNDA.n4325 GNDA.n4273 0.1255
R18061 GNDA.n4213 GNDA.n4197 0.1255
R18062 GNDA.n4230 GNDA.n4229 0.1255
R18063 GNDA.n4243 GNDA.n4191 0.1255
R18064 GNDA.n3967 GNDA.n499 0.1255
R18065 GNDA.n3984 GNDA.n3983 0.1255
R18066 GNDA.n3997 GNDA.n493 0.1255
R18067 GNDA.n4131 GNDA.n4115 0.1255
R18068 GNDA.n4148 GNDA.n4147 0.1255
R18069 GNDA.n4161 GNDA.n4109 0.1255
R18070 GNDA.n4049 GNDA.n4033 0.1255
R18071 GNDA.n4066 GNDA.n4065 0.1255
R18072 GNDA.n4079 GNDA.n4027 0.1255
R18073 GNDA.n3869 GNDA.n3868 0.1255
R18074 GNDA.n3875 GNDA.n3874 0.1255
R18075 GNDA.n3881 GNDA.n3880 0.1255
R18076 GNDA.n1688 GNDA.n1677 0.1255
R18077 GNDA.n1705 GNDA.n1704 0.1255
R18078 GNDA.n1718 GNDA.n1671 0.1255
R18079 GNDA.n3806 GNDA.n3795 0.1255
R18080 GNDA.n3823 GNDA.n3822 0.1255
R18081 GNDA.n3836 GNDA.n3789 0.1255
R18082 GNDA.n3730 GNDA.n535 0.1255
R18083 GNDA.n3747 GNDA.n3746 0.1255
R18084 GNDA.n3760 GNDA.n529 0.1255
R18085 GNDA.n3572 GNDA.n3561 0.1255
R18086 GNDA.n3589 GNDA.n3588 0.1255
R18087 GNDA.n3602 GNDA.n3555 0.1255
R18088 GNDA.n3496 GNDA.n575 0.1255
R18089 GNDA.n3513 GNDA.n3512 0.1255
R18090 GNDA.n3526 GNDA.n569 0.1255
R18091 GNDA.n3398 GNDA.n3397 0.1255
R18092 GNDA.n3404 GNDA.n3403 0.1255
R18093 GNDA.n3410 GNDA.n3409 0.1255
R18094 GNDA.n3262 GNDA.n615 0.1255
R18095 GNDA.n3279 GNDA.n3278 0.1255
R18096 GNDA.n3292 GNDA.n609 0.1255
R18097 GNDA.n3164 GNDA.n3163 0.1255
R18098 GNDA.n3170 GNDA.n3169 0.1255
R18099 GNDA.n3176 GNDA.n3175 0.1255
R18100 GNDA.n1612 GNDA.n1596 0.1255
R18101 GNDA.n1629 GNDA.n1628 0.1255
R18102 GNDA.n1642 GNDA.n1590 0.1255
R18103 GNDA.n1530 GNDA.n1514 0.1255
R18104 GNDA.n1547 GNDA.n1546 0.1255
R18105 GNDA.n1560 GNDA.n1508 0.1255
R18106 GNDA.n1448 GNDA.n1432 0.1255
R18107 GNDA.n1465 GNDA.n1464 0.1255
R18108 GNDA.n1478 GNDA.n1426 0.1255
R18109 GNDA.n1175 GNDA.n1174 0.1255
R18110 GNDA.n1181 GNDA.n1180 0.1255
R18111 GNDA.n1187 GNDA.n1186 0.1255
R18112 GNDA.n1880 GNDA.n1163 0.1255
R18113 GNDA.n1897 GNDA.n1896 0.1255
R18114 GNDA.n1910 GNDA.n1157 0.1255
R18115 GNDA.n1832 GNDA.n1831 0.1255
R18116 GNDA.n1821 GNDA.n1788 0.1255
R18117 GNDA.n1814 GNDA.n1813 0.1255
R18118 GNDA.n1759 GNDA.n1758 0.1255
R18119 GNDA.n4610 GNDA.n4609 0.1255
R18120 GNDA.n2390 GNDA.n2301 0.1255
R18121 GNDA.n2295 GNDA.n2288 0.1255
R18122 GNDA.n2171 GNDA.n2155 0.1255
R18123 GNDA.n2184 GNDA.n2183 0.1255
R18124 GNDA.n2195 GNDA.n2143 0.1255
R18125 GNDA.n359 GNDA.n358 0.1255
R18126 GNDA.n2084 GNDA.n2072 0.1255
R18127 GNDA.n2103 GNDA.n2102 0.1255
R18128 GNDA.n2114 GNDA.n2066 0.1255
R18129 GNDA.n2088 GNDA.n2087 0.1255
R18130 GNDA.n2101 GNDA.n2069 0.1255
R18131 GNDA.n2118 GNDA.n2117 0.1255
R18132 GNDA.n1316 GNDA.n1314 0.115083
R18133 GNDA.n1314 GNDA.n1312 0.115083
R18134 GNDA.n1312 GNDA.n1310 0.115083
R18135 GNDA.n1310 GNDA.n1308 0.115083
R18136 GNDA.n1308 GNDA.n1306 0.115083
R18137 GNDA.n1342 GNDA.n1341 0.115083
R18138 GNDA.n1341 GNDA.n1339 0.115083
R18139 GNDA.n1376 GNDA.n1374 0.115083
R18140 GNDA.n1374 GNDA.n1372 0.115083
R18141 GNDA.n1372 GNDA.n1370 0.115083
R18142 GNDA.n1370 GNDA.n1368 0.115083
R18143 GNDA.n1368 GNDA.n1366 0.115083
R18144 GNDA.n2245 GNDA.n2243 0.115083
R18145 GNDA.n2247 GNDA.n2245 0.115083
R18146 GNDA.n2509 GNDA.n2508 0.115083
R18147 GNDA.n2508 GNDA.n2507 0.115083
R18148 GNDA.n2507 GNDA.n2506 0.115083
R18149 GNDA.n2506 GNDA.n676 0.115083
R18150 GNDA.n3059 GNDA.n3058 0.115083
R18151 GNDA.n3058 GNDA.n3057 0.115083
R18152 GNDA.n3057 GNDA.n3056 0.115083
R18153 GNDA.n3054 GNDA.n3053 0.115083
R18154 GNDA.n3053 GNDA.n3052 0.115083
R18155 GNDA.n3052 GNDA.n3051 0.115083
R18156 GNDA.n3156 GNDA.n624 0.105167
R18157 GNDA.n3862 GNDA.n3861 0.105167
R18158 GNDA.n1750 GNDA.n1742 0.09425
R18159 GNDA.n4618 GNDA.n437 0.09425
R18160 GNDA.n2011 GNDA 0.0817953
R18161 GNDA.n1337 GNDA.n1333 0.0734167
R18162 GNDA.n1349 GNDA.n1348 0.0734167
R18163 GNDA.n3702 GNDA.n3626 0.0734167
R18164 GNDA.n3702 GNDA.n3701 0.0734167
R18165 GNDA.n3701 GNDA.n3700 0.0734167
R18166 GNDA.n3695 GNDA.n3694 0.0734167
R18167 GNDA.n3694 GNDA.n3640 0.0734167
R18168 GNDA.n3690 GNDA.n3640 0.0734167
R18169 GNDA.n3684 GNDA.n3648 0.0734167
R18170 GNDA.n3684 GNDA.n3683 0.0734167
R18171 GNDA.n3683 GNDA.n3682 0.0734167
R18172 GNDA.n3677 GNDA.n3676 0.0734167
R18173 GNDA.n3676 GNDA.n3664 0.0734167
R18174 GNDA.n3330 GNDA.n590 0.0734167
R18175 GNDA.n3331 GNDA.n3330 0.0734167
R18176 GNDA.n3331 GNDA.n3328 0.0734167
R18177 GNDA.n3341 GNDA.n3326 0.0734167
R18178 GNDA.n3349 GNDA.n3326 0.0734167
R18179 GNDA.n3350 GNDA.n3349 0.0734167
R18180 GNDA.n3360 GNDA.n3359 0.0734167
R18181 GNDA.n3361 GNDA.n3360 0.0734167
R18182 GNDA.n3361 GNDA.n3322 0.0734167
R18183 GNDA.n3371 GNDA.n3320 0.0734167
R18184 GNDA.n3379 GNDA.n3320 0.0734167
R18185 GNDA.n4527 GNDA.n474 0.0734167
R18186 GNDA.n4528 GNDA.n4527 0.0734167
R18187 GNDA.n4528 GNDA.n4525 0.0734167
R18188 GNDA.n4538 GNDA.n4523 0.0734167
R18189 GNDA.n4546 GNDA.n4523 0.0734167
R18190 GNDA.n4547 GNDA.n4546 0.0734167
R18191 GNDA.n4557 GNDA.n4556 0.0734167
R18192 GNDA.n4558 GNDA.n4557 0.0734167
R18193 GNDA.n4558 GNDA.n4519 0.0734167
R18194 GNDA.n4568 GNDA.n4517 0.0734167
R18195 GNDA.n4576 GNDA.n4517 0.0734167
R18196 GNDA.n4451 GNDA.n4450 0.0734167
R18197 GNDA.n4452 GNDA.n4451 0.0734167
R18198 GNDA.n4452 GNDA.n4444 0.0734167
R18199 GNDA.n4462 GNDA.n4442 0.0734167
R18200 GNDA.n4470 GNDA.n4442 0.0734167
R18201 GNDA.n4471 GNDA.n4470 0.0734167
R18202 GNDA.n4481 GNDA.n4480 0.0734167
R18203 GNDA.n4482 GNDA.n4481 0.0734167
R18204 GNDA.n4482 GNDA.n4438 0.0734167
R18205 GNDA.n4492 GNDA.n4436 0.0734167
R18206 GNDA.n4500 GNDA.n4436 0.0734167
R18207 GNDA.n4369 GNDA.n4368 0.0734167
R18208 GNDA.n4370 GNDA.n4369 0.0734167
R18209 GNDA.n4370 GNDA.n4362 0.0734167
R18210 GNDA.n4380 GNDA.n4360 0.0734167
R18211 GNDA.n4388 GNDA.n4360 0.0734167
R18212 GNDA.n4389 GNDA.n4388 0.0734167
R18213 GNDA.n4399 GNDA.n4398 0.0734167
R18214 GNDA.n4400 GNDA.n4399 0.0734167
R18215 GNDA.n4400 GNDA.n4356 0.0734167
R18216 GNDA.n4410 GNDA.n4354 0.0734167
R18217 GNDA.n4418 GNDA.n4354 0.0734167
R18218 GNDA.n4287 GNDA.n4286 0.0734167
R18219 GNDA.n4288 GNDA.n4287 0.0734167
R18220 GNDA.n4288 GNDA.n4280 0.0734167
R18221 GNDA.n4298 GNDA.n4278 0.0734167
R18222 GNDA.n4306 GNDA.n4278 0.0734167
R18223 GNDA.n4307 GNDA.n4306 0.0734167
R18224 GNDA.n4317 GNDA.n4316 0.0734167
R18225 GNDA.n4318 GNDA.n4317 0.0734167
R18226 GNDA.n4318 GNDA.n4274 0.0734167
R18227 GNDA.n4328 GNDA.n4272 0.0734167
R18228 GNDA.n4336 GNDA.n4272 0.0734167
R18229 GNDA.n4205 GNDA.n4204 0.0734167
R18230 GNDA.n4206 GNDA.n4205 0.0734167
R18231 GNDA.n4206 GNDA.n4198 0.0734167
R18232 GNDA.n4216 GNDA.n4196 0.0734167
R18233 GNDA.n4224 GNDA.n4196 0.0734167
R18234 GNDA.n4225 GNDA.n4224 0.0734167
R18235 GNDA.n4235 GNDA.n4234 0.0734167
R18236 GNDA.n4236 GNDA.n4235 0.0734167
R18237 GNDA.n4236 GNDA.n4192 0.0734167
R18238 GNDA.n4246 GNDA.n4190 0.0734167
R18239 GNDA.n4254 GNDA.n4190 0.0734167
R18240 GNDA.n3959 GNDA.n3958 0.0734167
R18241 GNDA.n3960 GNDA.n3959 0.0734167
R18242 GNDA.n3960 GNDA.n500 0.0734167
R18243 GNDA.n3970 GNDA.n498 0.0734167
R18244 GNDA.n3978 GNDA.n498 0.0734167
R18245 GNDA.n3979 GNDA.n3978 0.0734167
R18246 GNDA.n3989 GNDA.n3988 0.0734167
R18247 GNDA.n3990 GNDA.n3989 0.0734167
R18248 GNDA.n3990 GNDA.n494 0.0734167
R18249 GNDA.n4000 GNDA.n492 0.0734167
R18250 GNDA.n4008 GNDA.n492 0.0734167
R18251 GNDA.n4123 GNDA.n4122 0.0734167
R18252 GNDA.n4124 GNDA.n4123 0.0734167
R18253 GNDA.n4124 GNDA.n4116 0.0734167
R18254 GNDA.n4134 GNDA.n4114 0.0734167
R18255 GNDA.n4142 GNDA.n4114 0.0734167
R18256 GNDA.n4143 GNDA.n4142 0.0734167
R18257 GNDA.n4153 GNDA.n4152 0.0734167
R18258 GNDA.n4154 GNDA.n4153 0.0734167
R18259 GNDA.n4154 GNDA.n4110 0.0734167
R18260 GNDA.n4164 GNDA.n4108 0.0734167
R18261 GNDA.n4172 GNDA.n4108 0.0734167
R18262 GNDA.n4041 GNDA.n4040 0.0734167
R18263 GNDA.n4042 GNDA.n4041 0.0734167
R18264 GNDA.n4042 GNDA.n4034 0.0734167
R18265 GNDA.n4052 GNDA.n4032 0.0734167
R18266 GNDA.n4060 GNDA.n4032 0.0734167
R18267 GNDA.n4061 GNDA.n4060 0.0734167
R18268 GNDA.n4071 GNDA.n4070 0.0734167
R18269 GNDA.n4072 GNDA.n4071 0.0734167
R18270 GNDA.n4072 GNDA.n4028 0.0734167
R18271 GNDA.n4082 GNDA.n4026 0.0734167
R18272 GNDA.n4090 GNDA.n4026 0.0734167
R18273 GNDA.n3886 GNDA.n3863 0.0734167
R18274 GNDA.n3887 GNDA.n3886 0.0734167
R18275 GNDA.n3888 GNDA.n3887 0.0734167
R18276 GNDA.n3892 GNDA.n3891 0.0734167
R18277 GNDA.n3893 GNDA.n3892 0.0734167
R18278 GNDA.n3894 GNDA.n3893 0.0734167
R18279 GNDA.n3898 GNDA.n3897 0.0734167
R18280 GNDA.n3899 GNDA.n3898 0.0734167
R18281 GNDA.n3900 GNDA.n3899 0.0734167
R18282 GNDA.n3904 GNDA.n3903 0.0734167
R18283 GNDA.n3905 GNDA.n3904 0.0734167
R18284 GNDA.n1680 GNDA.n1408 0.0734167
R18285 GNDA.n1681 GNDA.n1680 0.0734167
R18286 GNDA.n1681 GNDA.n1678 0.0734167
R18287 GNDA.n1691 GNDA.n1676 0.0734167
R18288 GNDA.n1699 GNDA.n1676 0.0734167
R18289 GNDA.n1700 GNDA.n1699 0.0734167
R18290 GNDA.n1710 GNDA.n1709 0.0734167
R18291 GNDA.n1711 GNDA.n1710 0.0734167
R18292 GNDA.n1711 GNDA.n1672 0.0734167
R18293 GNDA.n1721 GNDA.n1670 0.0734167
R18294 GNDA.n1729 GNDA.n1670 0.0734167
R18295 GNDA.n3798 GNDA.n510 0.0734167
R18296 GNDA.n3799 GNDA.n3798 0.0734167
R18297 GNDA.n3799 GNDA.n3796 0.0734167
R18298 GNDA.n3809 GNDA.n3794 0.0734167
R18299 GNDA.n3817 GNDA.n3794 0.0734167
R18300 GNDA.n3818 GNDA.n3817 0.0734167
R18301 GNDA.n3828 GNDA.n3827 0.0734167
R18302 GNDA.n3829 GNDA.n3828 0.0734167
R18303 GNDA.n3829 GNDA.n3790 0.0734167
R18304 GNDA.n3839 GNDA.n3788 0.0734167
R18305 GNDA.n3847 GNDA.n3788 0.0734167
R18306 GNDA.n3722 GNDA.n3721 0.0734167
R18307 GNDA.n3723 GNDA.n3722 0.0734167
R18308 GNDA.n3723 GNDA.n536 0.0734167
R18309 GNDA.n3733 GNDA.n534 0.0734167
R18310 GNDA.n3741 GNDA.n534 0.0734167
R18311 GNDA.n3742 GNDA.n3741 0.0734167
R18312 GNDA.n3752 GNDA.n3751 0.0734167
R18313 GNDA.n3753 GNDA.n3752 0.0734167
R18314 GNDA.n3753 GNDA.n530 0.0734167
R18315 GNDA.n3763 GNDA.n528 0.0734167
R18316 GNDA.n3771 GNDA.n528 0.0734167
R18317 GNDA.n3564 GNDA.n550 0.0734167
R18318 GNDA.n3565 GNDA.n3564 0.0734167
R18319 GNDA.n3565 GNDA.n3562 0.0734167
R18320 GNDA.n3575 GNDA.n3560 0.0734167
R18321 GNDA.n3583 GNDA.n3560 0.0734167
R18322 GNDA.n3584 GNDA.n3583 0.0734167
R18323 GNDA.n3594 GNDA.n3593 0.0734167
R18324 GNDA.n3595 GNDA.n3594 0.0734167
R18325 GNDA.n3595 GNDA.n3556 0.0734167
R18326 GNDA.n3605 GNDA.n3554 0.0734167
R18327 GNDA.n3613 GNDA.n3554 0.0734167
R18328 GNDA.n3488 GNDA.n3487 0.0734167
R18329 GNDA.n3489 GNDA.n3488 0.0734167
R18330 GNDA.n3489 GNDA.n576 0.0734167
R18331 GNDA.n3499 GNDA.n574 0.0734167
R18332 GNDA.n3507 GNDA.n574 0.0734167
R18333 GNDA.n3508 GNDA.n3507 0.0734167
R18334 GNDA.n3518 GNDA.n3517 0.0734167
R18335 GNDA.n3519 GNDA.n3518 0.0734167
R18336 GNDA.n3519 GNDA.n570 0.0734167
R18337 GNDA.n3529 GNDA.n568 0.0734167
R18338 GNDA.n3537 GNDA.n568 0.0734167
R18339 GNDA.n3415 GNDA.n3392 0.0734167
R18340 GNDA.n3416 GNDA.n3415 0.0734167
R18341 GNDA.n3417 GNDA.n3416 0.0734167
R18342 GNDA.n3421 GNDA.n3420 0.0734167
R18343 GNDA.n3422 GNDA.n3421 0.0734167
R18344 GNDA.n3423 GNDA.n3422 0.0734167
R18345 GNDA.n3427 GNDA.n3426 0.0734167
R18346 GNDA.n3428 GNDA.n3427 0.0734167
R18347 GNDA.n3429 GNDA.n3428 0.0734167
R18348 GNDA.n3433 GNDA.n3432 0.0734167
R18349 GNDA.n3434 GNDA.n3433 0.0734167
R18350 GNDA.n3254 GNDA.n3253 0.0734167
R18351 GNDA.n3255 GNDA.n3254 0.0734167
R18352 GNDA.n3255 GNDA.n616 0.0734167
R18353 GNDA.n3265 GNDA.n614 0.0734167
R18354 GNDA.n3273 GNDA.n614 0.0734167
R18355 GNDA.n3274 GNDA.n3273 0.0734167
R18356 GNDA.n3284 GNDA.n3283 0.0734167
R18357 GNDA.n3285 GNDA.n3284 0.0734167
R18358 GNDA.n3285 GNDA.n610 0.0734167
R18359 GNDA.n3295 GNDA.n608 0.0734167
R18360 GNDA.n3303 GNDA.n608 0.0734167
R18361 GNDA.n3181 GNDA.n3158 0.0734167
R18362 GNDA.n3182 GNDA.n3181 0.0734167
R18363 GNDA.n3183 GNDA.n3182 0.0734167
R18364 GNDA.n3187 GNDA.n3186 0.0734167
R18365 GNDA.n3188 GNDA.n3187 0.0734167
R18366 GNDA.n3189 GNDA.n3188 0.0734167
R18367 GNDA.n3193 GNDA.n3192 0.0734167
R18368 GNDA.n3194 GNDA.n3193 0.0734167
R18369 GNDA.n3195 GNDA.n3194 0.0734167
R18370 GNDA.n3199 GNDA.n3198 0.0734167
R18371 GNDA.n3200 GNDA.n3199 0.0734167
R18372 GNDA.n1604 GNDA.n1603 0.0734167
R18373 GNDA.n1605 GNDA.n1604 0.0734167
R18374 GNDA.n1605 GNDA.n1597 0.0734167
R18375 GNDA.n1615 GNDA.n1595 0.0734167
R18376 GNDA.n1623 GNDA.n1595 0.0734167
R18377 GNDA.n1624 GNDA.n1623 0.0734167
R18378 GNDA.n1634 GNDA.n1633 0.0734167
R18379 GNDA.n1635 GNDA.n1634 0.0734167
R18380 GNDA.n1635 GNDA.n1591 0.0734167
R18381 GNDA.n1645 GNDA.n1589 0.0734167
R18382 GNDA.n1653 GNDA.n1589 0.0734167
R18383 GNDA.n1522 GNDA.n1521 0.0734167
R18384 GNDA.n1523 GNDA.n1522 0.0734167
R18385 GNDA.n1523 GNDA.n1515 0.0734167
R18386 GNDA.n1533 GNDA.n1513 0.0734167
R18387 GNDA.n1541 GNDA.n1513 0.0734167
R18388 GNDA.n1542 GNDA.n1541 0.0734167
R18389 GNDA.n1552 GNDA.n1551 0.0734167
R18390 GNDA.n1553 GNDA.n1552 0.0734167
R18391 GNDA.n1553 GNDA.n1509 0.0734167
R18392 GNDA.n1563 GNDA.n1507 0.0734167
R18393 GNDA.n1571 GNDA.n1507 0.0734167
R18394 GNDA.n1440 GNDA.n1439 0.0734167
R18395 GNDA.n1441 GNDA.n1440 0.0734167
R18396 GNDA.n1441 GNDA.n1433 0.0734167
R18397 GNDA.n1451 GNDA.n1431 0.0734167
R18398 GNDA.n1459 GNDA.n1431 0.0734167
R18399 GNDA.n1460 GNDA.n1459 0.0734167
R18400 GNDA.n1470 GNDA.n1469 0.0734167
R18401 GNDA.n1471 GNDA.n1470 0.0734167
R18402 GNDA.n1471 GNDA.n1427 0.0734167
R18403 GNDA.n1481 GNDA.n1425 0.0734167
R18404 GNDA.n1489 GNDA.n1425 0.0734167
R18405 GNDA.n1192 GNDA.n1169 0.0734167
R18406 GNDA.n1193 GNDA.n1192 0.0734167
R18407 GNDA.n1194 GNDA.n1193 0.0734167
R18408 GNDA.n1198 GNDA.n1197 0.0734167
R18409 GNDA.n1199 GNDA.n1198 0.0734167
R18410 GNDA.n1200 GNDA.n1199 0.0734167
R18411 GNDA.n1204 GNDA.n1203 0.0734167
R18412 GNDA.n1205 GNDA.n1204 0.0734167
R18413 GNDA.n1206 GNDA.n1205 0.0734167
R18414 GNDA.n1210 GNDA.n1209 0.0734167
R18415 GNDA.n1211 GNDA.n1210 0.0734167
R18416 GNDA.n1872 GNDA.n1871 0.0734167
R18417 GNDA.n1873 GNDA.n1872 0.0734167
R18418 GNDA.n1873 GNDA.n1164 0.0734167
R18419 GNDA.n1883 GNDA.n1162 0.0734167
R18420 GNDA.n1891 GNDA.n1162 0.0734167
R18421 GNDA.n1892 GNDA.n1891 0.0734167
R18422 GNDA.n1902 GNDA.n1901 0.0734167
R18423 GNDA.n1903 GNDA.n1902 0.0734167
R18424 GNDA.n1903 GNDA.n1158 0.0734167
R18425 GNDA.n1913 GNDA.n1156 0.0734167
R18426 GNDA.n1921 GNDA.n1156 0.0734167
R18427 GNDA.n1836 GNDA.n1773 0.0734167
R18428 GNDA.n1836 GNDA.n1835 0.0734167
R18429 GNDA.n1835 GNDA.n1834 0.0734167
R18430 GNDA.n1829 GNDA.n1828 0.0734167
R18431 GNDA.n1828 GNDA.n1783 0.0734167
R18432 GNDA.n1824 GNDA.n1783 0.0734167
R18433 GNDA.n1818 GNDA.n1789 0.0734167
R18434 GNDA.n1818 GNDA.n1817 0.0734167
R18435 GNDA.n1817 GNDA.n1816 0.0734167
R18436 GNDA.n1811 GNDA.n1810 0.0734167
R18437 GNDA.n1810 GNDA.n1801 0.0734167
R18438 GNDA.n1763 GNDA.n1762 0.0734167
R18439 GNDA.n4606 GNDA.n4605 0.0734167
R18440 GNDA.n2166 GNDA.n2165 0.0734167
R18441 GNDA.n2166 GNDA.n2158 0.0734167
R18442 GNDA.n2174 GNDA.n2154 0.0734167
R18443 GNDA.n2180 GNDA.n2154 0.0734167
R18444 GNDA.n2181 GNDA.n2180 0.0734167
R18445 GNDA.n2189 GNDA.n2188 0.0734167
R18446 GNDA.n2190 GNDA.n2189 0.0734167
R18447 GNDA.n2190 GNDA.n2146 0.0734167
R18448 GNDA.n2198 GNDA.n2142 0.0734167
R18449 GNDA.n2204 GNDA.n2142 0.0734167
R18450 GNDA.n2205 GNDA.n2204 0.0734167
R18451 GNDA.n3706 GNDA.n3626 0.0682083
R18452 GNDA.n3700 GNDA.n3632 0.0682083
R18453 GNDA.n3696 GNDA.n3695 0.0682083
R18454 GNDA.n3690 GNDA.n3689 0.0682083
R18455 GNDA.n3688 GNDA.n3648 0.0682083
R18456 GNDA.n3682 GNDA.n3656 0.0682083
R18457 GNDA.n3678 GNDA.n3677 0.0682083
R18458 GNDA.n3385 GNDA.n590 0.0682083
R18459 GNDA.n3339 GNDA.n3328 0.0682083
R18460 GNDA.n3341 GNDA.n3340 0.0682083
R18461 GNDA.n3351 GNDA.n3350 0.0682083
R18462 GNDA.n3359 GNDA.n3324 0.0682083
R18463 GNDA.n3369 GNDA.n3322 0.0682083
R18464 GNDA.n3371 GNDA.n3370 0.0682083
R18465 GNDA.n4582 GNDA.n474 0.0682083
R18466 GNDA.n4536 GNDA.n4525 0.0682083
R18467 GNDA.n4538 GNDA.n4537 0.0682083
R18468 GNDA.n4548 GNDA.n4547 0.0682083
R18469 GNDA.n4556 GNDA.n4521 0.0682083
R18470 GNDA.n4566 GNDA.n4519 0.0682083
R18471 GNDA.n4568 GNDA.n4567 0.0682083
R18472 GNDA.n4450 GNDA.n4446 0.0682083
R18473 GNDA.n4460 GNDA.n4444 0.0682083
R18474 GNDA.n4462 GNDA.n4461 0.0682083
R18475 GNDA.n4472 GNDA.n4471 0.0682083
R18476 GNDA.n4480 GNDA.n4440 0.0682083
R18477 GNDA.n4490 GNDA.n4438 0.0682083
R18478 GNDA.n4492 GNDA.n4491 0.0682083
R18479 GNDA.n4368 GNDA.n4364 0.0682083
R18480 GNDA.n4378 GNDA.n4362 0.0682083
R18481 GNDA.n4380 GNDA.n4379 0.0682083
R18482 GNDA.n4390 GNDA.n4389 0.0682083
R18483 GNDA.n4398 GNDA.n4358 0.0682083
R18484 GNDA.n4408 GNDA.n4356 0.0682083
R18485 GNDA.n4410 GNDA.n4409 0.0682083
R18486 GNDA.n4286 GNDA.n4282 0.0682083
R18487 GNDA.n4296 GNDA.n4280 0.0682083
R18488 GNDA.n4298 GNDA.n4297 0.0682083
R18489 GNDA.n4308 GNDA.n4307 0.0682083
R18490 GNDA.n4316 GNDA.n4276 0.0682083
R18491 GNDA.n4326 GNDA.n4274 0.0682083
R18492 GNDA.n4328 GNDA.n4327 0.0682083
R18493 GNDA.n4204 GNDA.n4200 0.0682083
R18494 GNDA.n4214 GNDA.n4198 0.0682083
R18495 GNDA.n4216 GNDA.n4215 0.0682083
R18496 GNDA.n4226 GNDA.n4225 0.0682083
R18497 GNDA.n4234 GNDA.n4194 0.0682083
R18498 GNDA.n4244 GNDA.n4192 0.0682083
R18499 GNDA.n4246 GNDA.n4245 0.0682083
R18500 GNDA.n3958 GNDA.n3954 0.0682083
R18501 GNDA.n3968 GNDA.n500 0.0682083
R18502 GNDA.n3970 GNDA.n3969 0.0682083
R18503 GNDA.n3980 GNDA.n3979 0.0682083
R18504 GNDA.n3988 GNDA.n496 0.0682083
R18505 GNDA.n3998 GNDA.n494 0.0682083
R18506 GNDA.n4000 GNDA.n3999 0.0682083
R18507 GNDA.n4122 GNDA.n4118 0.0682083
R18508 GNDA.n4132 GNDA.n4116 0.0682083
R18509 GNDA.n4134 GNDA.n4133 0.0682083
R18510 GNDA.n4144 GNDA.n4143 0.0682083
R18511 GNDA.n4152 GNDA.n4112 0.0682083
R18512 GNDA.n4162 GNDA.n4110 0.0682083
R18513 GNDA.n4164 GNDA.n4163 0.0682083
R18514 GNDA.n4040 GNDA.n4036 0.0682083
R18515 GNDA.n4050 GNDA.n4034 0.0682083
R18516 GNDA.n4052 GNDA.n4051 0.0682083
R18517 GNDA.n4062 GNDA.n4061 0.0682083
R18518 GNDA.n4070 GNDA.n4030 0.0682083
R18519 GNDA.n4080 GNDA.n4028 0.0682083
R18520 GNDA.n4082 GNDA.n4081 0.0682083
R18521 GNDA.n3943 GNDA.n3863 0.0682083
R18522 GNDA.n3889 GNDA.n3888 0.0682083
R18523 GNDA.n3891 GNDA.n3890 0.0682083
R18524 GNDA.n3895 GNDA.n3894 0.0682083
R18525 GNDA.n3897 GNDA.n3896 0.0682083
R18526 GNDA.n3901 GNDA.n3900 0.0682083
R18527 GNDA.n3903 GNDA.n3902 0.0682083
R18528 GNDA.n1735 GNDA.n1408 0.0682083
R18529 GNDA.n1689 GNDA.n1678 0.0682083
R18530 GNDA.n1691 GNDA.n1690 0.0682083
R18531 GNDA.n1701 GNDA.n1700 0.0682083
R18532 GNDA.n1709 GNDA.n1674 0.0682083
R18533 GNDA.n1719 GNDA.n1672 0.0682083
R18534 GNDA.n1721 GNDA.n1720 0.0682083
R18535 GNDA.n3853 GNDA.n510 0.0682083
R18536 GNDA.n3807 GNDA.n3796 0.0682083
R18537 GNDA.n3809 GNDA.n3808 0.0682083
R18538 GNDA.n3819 GNDA.n3818 0.0682083
R18539 GNDA.n3827 GNDA.n3792 0.0682083
R18540 GNDA.n3837 GNDA.n3790 0.0682083
R18541 GNDA.n3839 GNDA.n3838 0.0682083
R18542 GNDA.n3721 GNDA.n3717 0.0682083
R18543 GNDA.n3731 GNDA.n536 0.0682083
R18544 GNDA.n3733 GNDA.n3732 0.0682083
R18545 GNDA.n3743 GNDA.n3742 0.0682083
R18546 GNDA.n3751 GNDA.n532 0.0682083
R18547 GNDA.n3761 GNDA.n530 0.0682083
R18548 GNDA.n3763 GNDA.n3762 0.0682083
R18549 GNDA.n3619 GNDA.n550 0.0682083
R18550 GNDA.n3573 GNDA.n3562 0.0682083
R18551 GNDA.n3575 GNDA.n3574 0.0682083
R18552 GNDA.n3585 GNDA.n3584 0.0682083
R18553 GNDA.n3593 GNDA.n3558 0.0682083
R18554 GNDA.n3603 GNDA.n3556 0.0682083
R18555 GNDA.n3605 GNDA.n3604 0.0682083
R18556 GNDA.n3487 GNDA.n3483 0.0682083
R18557 GNDA.n3497 GNDA.n576 0.0682083
R18558 GNDA.n3499 GNDA.n3498 0.0682083
R18559 GNDA.n3509 GNDA.n3508 0.0682083
R18560 GNDA.n3517 GNDA.n572 0.0682083
R18561 GNDA.n3527 GNDA.n570 0.0682083
R18562 GNDA.n3529 GNDA.n3528 0.0682083
R18563 GNDA.n3472 GNDA.n3392 0.0682083
R18564 GNDA.n3418 GNDA.n3417 0.0682083
R18565 GNDA.n3420 GNDA.n3419 0.0682083
R18566 GNDA.n3424 GNDA.n3423 0.0682083
R18567 GNDA.n3426 GNDA.n3425 0.0682083
R18568 GNDA.n3430 GNDA.n3429 0.0682083
R18569 GNDA.n3432 GNDA.n3431 0.0682083
R18570 GNDA.n3253 GNDA.n3249 0.0682083
R18571 GNDA.n3263 GNDA.n616 0.0682083
R18572 GNDA.n3265 GNDA.n3264 0.0682083
R18573 GNDA.n3275 GNDA.n3274 0.0682083
R18574 GNDA.n3283 GNDA.n612 0.0682083
R18575 GNDA.n3293 GNDA.n610 0.0682083
R18576 GNDA.n3295 GNDA.n3294 0.0682083
R18577 GNDA.n3238 GNDA.n3158 0.0682083
R18578 GNDA.n3184 GNDA.n3183 0.0682083
R18579 GNDA.n3186 GNDA.n3185 0.0682083
R18580 GNDA.n3190 GNDA.n3189 0.0682083
R18581 GNDA.n3192 GNDA.n3191 0.0682083
R18582 GNDA.n3196 GNDA.n3195 0.0682083
R18583 GNDA.n3198 GNDA.n3197 0.0682083
R18584 GNDA.n1603 GNDA.n1599 0.0682083
R18585 GNDA.n1613 GNDA.n1597 0.0682083
R18586 GNDA.n1615 GNDA.n1614 0.0682083
R18587 GNDA.n1625 GNDA.n1624 0.0682083
R18588 GNDA.n1633 GNDA.n1593 0.0682083
R18589 GNDA.n1643 GNDA.n1591 0.0682083
R18590 GNDA.n1645 GNDA.n1644 0.0682083
R18591 GNDA.n1521 GNDA.n1517 0.0682083
R18592 GNDA.n1531 GNDA.n1515 0.0682083
R18593 GNDA.n1533 GNDA.n1532 0.0682083
R18594 GNDA.n1543 GNDA.n1542 0.0682083
R18595 GNDA.n1551 GNDA.n1511 0.0682083
R18596 GNDA.n1561 GNDA.n1509 0.0682083
R18597 GNDA.n1563 GNDA.n1562 0.0682083
R18598 GNDA.n1439 GNDA.n1435 0.0682083
R18599 GNDA.n1449 GNDA.n1433 0.0682083
R18600 GNDA.n1451 GNDA.n1450 0.0682083
R18601 GNDA.n1461 GNDA.n1460 0.0682083
R18602 GNDA.n1469 GNDA.n1429 0.0682083
R18603 GNDA.n1479 GNDA.n1427 0.0682083
R18604 GNDA.n1481 GNDA.n1480 0.0682083
R18605 GNDA.n1249 GNDA.n1169 0.0682083
R18606 GNDA.n1195 GNDA.n1194 0.0682083
R18607 GNDA.n1197 GNDA.n1196 0.0682083
R18608 GNDA.n1201 GNDA.n1200 0.0682083
R18609 GNDA.n1203 GNDA.n1202 0.0682083
R18610 GNDA.n1207 GNDA.n1206 0.0682083
R18611 GNDA.n1209 GNDA.n1208 0.0682083
R18612 GNDA.n1871 GNDA.n1867 0.0682083
R18613 GNDA.n1881 GNDA.n1164 0.0682083
R18614 GNDA.n1883 GNDA.n1882 0.0682083
R18615 GNDA.n1893 GNDA.n1892 0.0682083
R18616 GNDA.n1901 GNDA.n1160 0.0682083
R18617 GNDA.n1911 GNDA.n1158 0.0682083
R18618 GNDA.n1913 GNDA.n1912 0.0682083
R18619 GNDA.n1840 GNDA.n1773 0.0682083
R18620 GNDA.n1834 GNDA.n1777 0.0682083
R18621 GNDA.n1830 GNDA.n1829 0.0682083
R18622 GNDA.n1824 GNDA.n1823 0.0682083
R18623 GNDA.n1822 GNDA.n1789 0.0682083
R18624 GNDA.n1816 GNDA.n1795 0.0682083
R18625 GNDA.n1812 GNDA.n1811 0.0682083
R18626 GNDA.n2172 GNDA.n2158 0.0682083
R18627 GNDA.n2174 GNDA.n2173 0.0682083
R18628 GNDA.n2182 GNDA.n2181 0.0682083
R18629 GNDA.n2188 GNDA.n2150 0.0682083
R18630 GNDA.n2196 GNDA.n2146 0.0682083
R18631 GNDA.n2198 GNDA.n2197 0.0682083
R18632 GNDA.n2218 GNDA.n2205 0.0682083
R18633 GNDA.n2164 GNDA.n2163 0.0672139
R18634 GNDA.n3673 GNDA.n3672 0.0672139
R18635 GNDA.n3380 GNDA.n3319 0.0672139
R18636 GNDA.n4577 GNDA.n4516 0.0672139
R18637 GNDA.n4501 GNDA.n4435 0.0672139
R18638 GNDA.n4419 GNDA.n4353 0.0672139
R18639 GNDA.n4337 GNDA.n4271 0.0672139
R18640 GNDA.n4255 GNDA.n4189 0.0672139
R18641 GNDA.n4009 GNDA.n491 0.0672139
R18642 GNDA.n4173 GNDA.n4107 0.0672139
R18643 GNDA.n4091 GNDA.n4025 0.0672139
R18644 GNDA.n3906 GNDA.n3885 0.0672139
R18645 GNDA.n1730 GNDA.n1669 0.0672139
R18646 GNDA.n3848 GNDA.n3787 0.0672139
R18647 GNDA.n3772 GNDA.n527 0.0672139
R18648 GNDA.n3614 GNDA.n3553 0.0672139
R18649 GNDA.n3538 GNDA.n567 0.0672139
R18650 GNDA.n3435 GNDA.n3414 0.0672139
R18651 GNDA.n3304 GNDA.n607 0.0672139
R18652 GNDA.n3201 GNDA.n3180 0.0672139
R18653 GNDA.n1654 GNDA.n1588 0.0672139
R18654 GNDA.n1572 GNDA.n1506 0.0672139
R18655 GNDA.n1490 GNDA.n1424 0.0672139
R18656 GNDA.n1212 GNDA.n1191 0.0672139
R18657 GNDA.n1922 GNDA.n1155 0.0672139
R18658 GNDA.n1807 GNDA.n1806 0.0672139
R18659 GNDA.n2077 GNDA.n2075 0.0667303
R18660 GNDA.n3696 GNDA.n3632 0.063
R18661 GNDA.n3689 GNDA.n3688 0.063
R18662 GNDA.n3678 GNDA.n3656 0.063
R18663 GNDA.n3340 GNDA.n3339 0.063
R18664 GNDA.n3351 GNDA.n3324 0.063
R18665 GNDA.n3370 GNDA.n3369 0.063
R18666 GNDA.n4537 GNDA.n4536 0.063
R18667 GNDA.n4548 GNDA.n4521 0.063
R18668 GNDA.n4567 GNDA.n4566 0.063
R18669 GNDA.n4461 GNDA.n4460 0.063
R18670 GNDA.n4472 GNDA.n4440 0.063
R18671 GNDA.n4491 GNDA.n4490 0.063
R18672 GNDA.n4379 GNDA.n4378 0.063
R18673 GNDA.n4390 GNDA.n4358 0.063
R18674 GNDA.n4409 GNDA.n4408 0.063
R18675 GNDA.n4297 GNDA.n4296 0.063
R18676 GNDA.n4308 GNDA.n4276 0.063
R18677 GNDA.n4327 GNDA.n4326 0.063
R18678 GNDA.n4215 GNDA.n4214 0.063
R18679 GNDA.n4226 GNDA.n4194 0.063
R18680 GNDA.n4245 GNDA.n4244 0.063
R18681 GNDA.n3969 GNDA.n3968 0.063
R18682 GNDA.n3980 GNDA.n496 0.063
R18683 GNDA.n3999 GNDA.n3998 0.063
R18684 GNDA.n4133 GNDA.n4132 0.063
R18685 GNDA.n4144 GNDA.n4112 0.063
R18686 GNDA.n4163 GNDA.n4162 0.063
R18687 GNDA.n4051 GNDA.n4050 0.063
R18688 GNDA.n4062 GNDA.n4030 0.063
R18689 GNDA.n4081 GNDA.n4080 0.063
R18690 GNDA.n3890 GNDA.n3889 0.063
R18691 GNDA.n3896 GNDA.n3895 0.063
R18692 GNDA.n3902 GNDA.n3901 0.063
R18693 GNDA.n1690 GNDA.n1689 0.063
R18694 GNDA.n1701 GNDA.n1674 0.063
R18695 GNDA.n1720 GNDA.n1719 0.063
R18696 GNDA.n3808 GNDA.n3807 0.063
R18697 GNDA.n3819 GNDA.n3792 0.063
R18698 GNDA.n3838 GNDA.n3837 0.063
R18699 GNDA.n3732 GNDA.n3731 0.063
R18700 GNDA.n3743 GNDA.n532 0.063
R18701 GNDA.n3762 GNDA.n3761 0.063
R18702 GNDA.n3574 GNDA.n3573 0.063
R18703 GNDA.n3585 GNDA.n3558 0.063
R18704 GNDA.n3604 GNDA.n3603 0.063
R18705 GNDA.n3498 GNDA.n3497 0.063
R18706 GNDA.n3509 GNDA.n572 0.063
R18707 GNDA.n3528 GNDA.n3527 0.063
R18708 GNDA.n3419 GNDA.n3418 0.063
R18709 GNDA.n3425 GNDA.n3424 0.063
R18710 GNDA.n3431 GNDA.n3430 0.063
R18711 GNDA.n3264 GNDA.n3263 0.063
R18712 GNDA.n3275 GNDA.n612 0.063
R18713 GNDA.n3294 GNDA.n3293 0.063
R18714 GNDA.n3185 GNDA.n3184 0.063
R18715 GNDA.n3191 GNDA.n3190 0.063
R18716 GNDA.n3197 GNDA.n3196 0.063
R18717 GNDA.n1614 GNDA.n1613 0.063
R18718 GNDA.n1625 GNDA.n1593 0.063
R18719 GNDA.n1644 GNDA.n1643 0.063
R18720 GNDA.n1532 GNDA.n1531 0.063
R18721 GNDA.n1543 GNDA.n1511 0.063
R18722 GNDA.n1562 GNDA.n1561 0.063
R18723 GNDA.n1450 GNDA.n1449 0.063
R18724 GNDA.n1461 GNDA.n1429 0.063
R18725 GNDA.n1480 GNDA.n1479 0.063
R18726 GNDA.n1196 GNDA.n1195 0.063
R18727 GNDA.n1202 GNDA.n1201 0.063
R18728 GNDA.n1208 GNDA.n1207 0.063
R18729 GNDA.n1882 GNDA.n1881 0.063
R18730 GNDA.n1893 GNDA.n1160 0.063
R18731 GNDA.n1912 GNDA.n1911 0.063
R18732 GNDA.n1830 GNDA.n1777 0.063
R18733 GNDA.n1823 GNDA.n1822 0.063
R18734 GNDA.n1812 GNDA.n1795 0.063
R18735 GNDA.n2173 GNDA.n2172 0.063
R18736 GNDA.n2182 GNDA.n2150 0.063
R18737 GNDA.n2197 GNDA.n2196 0.063
R18738 GNDA.n2510 GNDA.n2247 0.063
R18739 GNDA.n3056 GNDA.n3055 0.063
R18740 GNDA.n1738 GNDA.n624 0.0629369
R18741 GNDA.n3947 GNDA.n3862 0.0629369
R18742 GNDA.n2301 GNDA.n2300 0.0626438
R18743 GNDA.n2288 GNDA.n2287 0.0626438
R18744 GNDA.n2207 GNDA.n358 0.0626438
R18745 GNDA.n3633 GNDA.n3630 0.0553333
R18746 GNDA.n3644 GNDA.n3643 0.0553333
R18747 GNDA.n3657 GNDA.n3654 0.0553333
R18748 GNDA.n3668 GNDA.n3667 0.0553333
R18749 GNDA.n3333 GNDA.n3332 0.0553333
R18750 GNDA.n3347 GNDA.n3346 0.0553333
R18751 GNDA.n3363 GNDA.n3362 0.0553333
R18752 GNDA.n3377 GNDA.n3376 0.0553333
R18753 GNDA.n4530 GNDA.n4529 0.0553333
R18754 GNDA.n4544 GNDA.n4543 0.0553333
R18755 GNDA.n4560 GNDA.n4559 0.0553333
R18756 GNDA.n4574 GNDA.n4573 0.0553333
R18757 GNDA.n4454 GNDA.n4453 0.0553333
R18758 GNDA.n4468 GNDA.n4467 0.0553333
R18759 GNDA.n4484 GNDA.n4483 0.0553333
R18760 GNDA.n4498 GNDA.n4497 0.0553333
R18761 GNDA.n4372 GNDA.n4371 0.0553333
R18762 GNDA.n4386 GNDA.n4385 0.0553333
R18763 GNDA.n4402 GNDA.n4401 0.0553333
R18764 GNDA.n4416 GNDA.n4415 0.0553333
R18765 GNDA.n4290 GNDA.n4289 0.0553333
R18766 GNDA.n4304 GNDA.n4303 0.0553333
R18767 GNDA.n4320 GNDA.n4319 0.0553333
R18768 GNDA.n4334 GNDA.n4333 0.0553333
R18769 GNDA.n4208 GNDA.n4207 0.0553333
R18770 GNDA.n4222 GNDA.n4221 0.0553333
R18771 GNDA.n4238 GNDA.n4237 0.0553333
R18772 GNDA.n4252 GNDA.n4251 0.0553333
R18773 GNDA.n3962 GNDA.n3961 0.0553333
R18774 GNDA.n3976 GNDA.n3975 0.0553333
R18775 GNDA.n3992 GNDA.n3991 0.0553333
R18776 GNDA.n4006 GNDA.n4005 0.0553333
R18777 GNDA.n4126 GNDA.n4125 0.0553333
R18778 GNDA.n4140 GNDA.n4139 0.0553333
R18779 GNDA.n4156 GNDA.n4155 0.0553333
R18780 GNDA.n4170 GNDA.n4169 0.0553333
R18781 GNDA.n4044 GNDA.n4043 0.0553333
R18782 GNDA.n4058 GNDA.n4057 0.0553333
R18783 GNDA.n4074 GNDA.n4073 0.0553333
R18784 GNDA.n4088 GNDA.n4087 0.0553333
R18785 GNDA.n3938 GNDA.n3937 0.0553333
R18786 GNDA.n3929 GNDA.n3928 0.0553333
R18787 GNDA.n3920 GNDA.n3919 0.0553333
R18788 GNDA.n3911 GNDA.n3910 0.0553333
R18789 GNDA.n1683 GNDA.n1682 0.0553333
R18790 GNDA.n1697 GNDA.n1696 0.0553333
R18791 GNDA.n1713 GNDA.n1712 0.0553333
R18792 GNDA.n1727 GNDA.n1726 0.0553333
R18793 GNDA.n3801 GNDA.n3800 0.0553333
R18794 GNDA.n3815 GNDA.n3814 0.0553333
R18795 GNDA.n3831 GNDA.n3830 0.0553333
R18796 GNDA.n3845 GNDA.n3844 0.0553333
R18797 GNDA.n3725 GNDA.n3724 0.0553333
R18798 GNDA.n3739 GNDA.n3738 0.0553333
R18799 GNDA.n3755 GNDA.n3754 0.0553333
R18800 GNDA.n3769 GNDA.n3768 0.0553333
R18801 GNDA.n3567 GNDA.n3566 0.0553333
R18802 GNDA.n3581 GNDA.n3580 0.0553333
R18803 GNDA.n3597 GNDA.n3596 0.0553333
R18804 GNDA.n3611 GNDA.n3610 0.0553333
R18805 GNDA.n3491 GNDA.n3490 0.0553333
R18806 GNDA.n3505 GNDA.n3504 0.0553333
R18807 GNDA.n3521 GNDA.n3520 0.0553333
R18808 GNDA.n3535 GNDA.n3534 0.0553333
R18809 GNDA.n3467 GNDA.n3466 0.0553333
R18810 GNDA.n3458 GNDA.n3457 0.0553333
R18811 GNDA.n3449 GNDA.n3448 0.0553333
R18812 GNDA.n3440 GNDA.n3439 0.0553333
R18813 GNDA.n3257 GNDA.n3256 0.0553333
R18814 GNDA.n3271 GNDA.n3270 0.0553333
R18815 GNDA.n3287 GNDA.n3286 0.0553333
R18816 GNDA.n3301 GNDA.n3300 0.0553333
R18817 GNDA.n3233 GNDA.n3232 0.0553333
R18818 GNDA.n3224 GNDA.n3223 0.0553333
R18819 GNDA.n3215 GNDA.n3214 0.0553333
R18820 GNDA.n3206 GNDA.n3205 0.0553333
R18821 GNDA.n1607 GNDA.n1606 0.0553333
R18822 GNDA.n1621 GNDA.n1620 0.0553333
R18823 GNDA.n1637 GNDA.n1636 0.0553333
R18824 GNDA.n1651 GNDA.n1650 0.0553333
R18825 GNDA.n1525 GNDA.n1524 0.0553333
R18826 GNDA.n1539 GNDA.n1538 0.0553333
R18827 GNDA.n1555 GNDA.n1554 0.0553333
R18828 GNDA.n1569 GNDA.n1568 0.0553333
R18829 GNDA.n1443 GNDA.n1442 0.0553333
R18830 GNDA.n1457 GNDA.n1456 0.0553333
R18831 GNDA.n1473 GNDA.n1472 0.0553333
R18832 GNDA.n1487 GNDA.n1486 0.0553333
R18833 GNDA.n1244 GNDA.n1243 0.0553333
R18834 GNDA.n1235 GNDA.n1234 0.0553333
R18835 GNDA.n1226 GNDA.n1225 0.0553333
R18836 GNDA.n1217 GNDA.n1216 0.0553333
R18837 GNDA.n1875 GNDA.n1874 0.0553333
R18838 GNDA.n1889 GNDA.n1888 0.0553333
R18839 GNDA.n1905 GNDA.n1904 0.0553333
R18840 GNDA.n1919 GNDA.n1918 0.0553333
R18841 GNDA.n1775 GNDA.n1774 0.0553333
R18842 GNDA.n1779 GNDA.n1778 0.0553333
R18843 GNDA.n1785 GNDA.n1784 0.0553333
R18844 GNDA.n1787 GNDA.n1786 0.0553333
R18845 GNDA.n1793 GNDA.n1792 0.0553333
R18846 GNDA.n1797 GNDA.n1796 0.0553333
R18847 GNDA.n1803 GNDA.n1802 0.0553333
R18848 GNDA.n1805 GNDA.n1804 0.0553333
R18849 GNDA.n2161 GNDA.n2160 0.0553333
R18850 GNDA.n2178 GNDA.n2177 0.0553333
R18851 GNDA.n2149 GNDA.n2148 0.0553333
R18852 GNDA.n2202 GNDA.n2201 0.0553333
R18853 GNDA.n2080 GNDA.n2079 0.0553333
R18854 GNDA.n2096 GNDA.n2095 0.0553333
R18855 GNDA.n2110 GNDA.n2109 0.0553333
R18856 GNDA.n2126 GNDA.n2064 0.0553333
R18857 GNDA.n3008 GNDA 0.0517
R18858 GNDA.n3085 GNDA 0.0517
R18859 GNDA GNDA.n202 0.0517
R18860 GNDA.n2712 GNDA 0.0517
R18861 GNDA GNDA.n4904 0.0517
R18862 GNDA GNDA.n5183 0.0517
R18863 GNDA.n4761 GNDA 0.0517
R18864 GNDA.n2415 GNDA 0.0517
R18865 GNDA GNDA.n0 0.0517
R18866 GNDA.n3628 GNDA.n3627 0.0514167
R18867 GNDA.n3636 GNDA.n3635 0.0514167
R18868 GNDA.n3641 GNDA.n3638 0.0514167
R18869 GNDA.n3649 GNDA.n3646 0.0514167
R18870 GNDA.n3652 GNDA.n3651 0.0514167
R18871 GNDA.n3660 GNDA.n3659 0.0514167
R18872 GNDA.n3665 GNDA.n3662 0.0514167
R18873 GNDA.n3671 GNDA.n3670 0.0514167
R18874 GNDA.n3383 GNDA.n592 0.0514167
R18875 GNDA.n3337 GNDA.n3336 0.0514167
R18876 GNDA.n3343 GNDA.n3342 0.0514167
R18877 GNDA.n3353 GNDA.n3352 0.0514167
R18878 GNDA.n3357 GNDA.n3356 0.0514167
R18879 GNDA.n3367 GNDA.n3366 0.0514167
R18880 GNDA.n3373 GNDA.n3372 0.0514167
R18881 GNDA.n3381 GNDA.n3318 0.0514167
R18882 GNDA.n4580 GNDA.n476 0.0514167
R18883 GNDA.n4534 GNDA.n4533 0.0514167
R18884 GNDA.n4540 GNDA.n4539 0.0514167
R18885 GNDA.n4550 GNDA.n4549 0.0514167
R18886 GNDA.n4554 GNDA.n4553 0.0514167
R18887 GNDA.n4564 GNDA.n4563 0.0514167
R18888 GNDA.n4570 GNDA.n4569 0.0514167
R18889 GNDA.n4578 GNDA.n4515 0.0514167
R18890 GNDA.n4448 GNDA.n4422 0.0514167
R18891 GNDA.n4458 GNDA.n4457 0.0514167
R18892 GNDA.n4464 GNDA.n4463 0.0514167
R18893 GNDA.n4474 GNDA.n4473 0.0514167
R18894 GNDA.n4478 GNDA.n4477 0.0514167
R18895 GNDA.n4488 GNDA.n4487 0.0514167
R18896 GNDA.n4494 GNDA.n4493 0.0514167
R18897 GNDA.n4502 GNDA.n4434 0.0514167
R18898 GNDA.n4366 GNDA.n4340 0.0514167
R18899 GNDA.n4376 GNDA.n4375 0.0514167
R18900 GNDA.n4382 GNDA.n4381 0.0514167
R18901 GNDA.n4392 GNDA.n4391 0.0514167
R18902 GNDA.n4396 GNDA.n4395 0.0514167
R18903 GNDA.n4406 GNDA.n4405 0.0514167
R18904 GNDA.n4412 GNDA.n4411 0.0514167
R18905 GNDA.n4420 GNDA.n4352 0.0514167
R18906 GNDA.n4284 GNDA.n4258 0.0514167
R18907 GNDA.n4294 GNDA.n4293 0.0514167
R18908 GNDA.n4300 GNDA.n4299 0.0514167
R18909 GNDA.n4310 GNDA.n4309 0.0514167
R18910 GNDA.n4314 GNDA.n4313 0.0514167
R18911 GNDA.n4324 GNDA.n4323 0.0514167
R18912 GNDA.n4330 GNDA.n4329 0.0514167
R18913 GNDA.n4338 GNDA.n4270 0.0514167
R18914 GNDA.n4202 GNDA.n4176 0.0514167
R18915 GNDA.n4212 GNDA.n4211 0.0514167
R18916 GNDA.n4218 GNDA.n4217 0.0514167
R18917 GNDA.n4228 GNDA.n4227 0.0514167
R18918 GNDA.n4232 GNDA.n4231 0.0514167
R18919 GNDA.n4242 GNDA.n4241 0.0514167
R18920 GNDA.n4248 GNDA.n4247 0.0514167
R18921 GNDA.n4256 GNDA.n4188 0.0514167
R18922 GNDA.n3956 GNDA.n478 0.0514167
R18923 GNDA.n3966 GNDA.n3965 0.0514167
R18924 GNDA.n3972 GNDA.n3971 0.0514167
R18925 GNDA.n3982 GNDA.n3981 0.0514167
R18926 GNDA.n3986 GNDA.n3985 0.0514167
R18927 GNDA.n3996 GNDA.n3995 0.0514167
R18928 GNDA.n4002 GNDA.n4001 0.0514167
R18929 GNDA.n4010 GNDA.n490 0.0514167
R18930 GNDA.n4120 GNDA.n4094 0.0514167
R18931 GNDA.n4130 GNDA.n4129 0.0514167
R18932 GNDA.n4136 GNDA.n4135 0.0514167
R18933 GNDA.n4146 GNDA.n4145 0.0514167
R18934 GNDA.n4150 GNDA.n4149 0.0514167
R18935 GNDA.n4160 GNDA.n4159 0.0514167
R18936 GNDA.n4166 GNDA.n4165 0.0514167
R18937 GNDA.n4174 GNDA.n4106 0.0514167
R18938 GNDA.n4038 GNDA.n4012 0.0514167
R18939 GNDA.n4048 GNDA.n4047 0.0514167
R18940 GNDA.n4054 GNDA.n4053 0.0514167
R18941 GNDA.n4064 GNDA.n4063 0.0514167
R18942 GNDA.n4068 GNDA.n4067 0.0514167
R18943 GNDA.n4078 GNDA.n4077 0.0514167
R18944 GNDA.n4084 GNDA.n4083 0.0514167
R18945 GNDA.n4092 GNDA.n4024 0.0514167
R18946 GNDA.n3941 GNDA.n3940 0.0514167
R18947 GNDA.n3935 GNDA.n3934 0.0514167
R18948 GNDA.n3932 GNDA.n3931 0.0514167
R18949 GNDA.n3926 GNDA.n3925 0.0514167
R18950 GNDA.n3923 GNDA.n3922 0.0514167
R18951 GNDA.n3917 GNDA.n3916 0.0514167
R18952 GNDA.n3914 GNDA.n3913 0.0514167
R18953 GNDA.n3908 GNDA.n3907 0.0514167
R18954 GNDA.n1733 GNDA.n1410 0.0514167
R18955 GNDA.n1687 GNDA.n1686 0.0514167
R18956 GNDA.n1693 GNDA.n1692 0.0514167
R18957 GNDA.n1703 GNDA.n1702 0.0514167
R18958 GNDA.n1707 GNDA.n1706 0.0514167
R18959 GNDA.n1717 GNDA.n1716 0.0514167
R18960 GNDA.n1723 GNDA.n1722 0.0514167
R18961 GNDA.n1731 GNDA.n1668 0.0514167
R18962 GNDA.n3851 GNDA.n512 0.0514167
R18963 GNDA.n3805 GNDA.n3804 0.0514167
R18964 GNDA.n3811 GNDA.n3810 0.0514167
R18965 GNDA.n3821 GNDA.n3820 0.0514167
R18966 GNDA.n3825 GNDA.n3824 0.0514167
R18967 GNDA.n3835 GNDA.n3834 0.0514167
R18968 GNDA.n3841 GNDA.n3840 0.0514167
R18969 GNDA.n3849 GNDA.n3786 0.0514167
R18970 GNDA.n3719 GNDA.n514 0.0514167
R18971 GNDA.n3729 GNDA.n3728 0.0514167
R18972 GNDA.n3735 GNDA.n3734 0.0514167
R18973 GNDA.n3745 GNDA.n3744 0.0514167
R18974 GNDA.n3749 GNDA.n3748 0.0514167
R18975 GNDA.n3759 GNDA.n3758 0.0514167
R18976 GNDA.n3765 GNDA.n3764 0.0514167
R18977 GNDA.n3773 GNDA.n526 0.0514167
R18978 GNDA.n3617 GNDA.n552 0.0514167
R18979 GNDA.n3571 GNDA.n3570 0.0514167
R18980 GNDA.n3577 GNDA.n3576 0.0514167
R18981 GNDA.n3587 GNDA.n3586 0.0514167
R18982 GNDA.n3591 GNDA.n3590 0.0514167
R18983 GNDA.n3601 GNDA.n3600 0.0514167
R18984 GNDA.n3607 GNDA.n3606 0.0514167
R18985 GNDA.n3615 GNDA.n3552 0.0514167
R18986 GNDA.n3485 GNDA.n554 0.0514167
R18987 GNDA.n3495 GNDA.n3494 0.0514167
R18988 GNDA.n3501 GNDA.n3500 0.0514167
R18989 GNDA.n3511 GNDA.n3510 0.0514167
R18990 GNDA.n3515 GNDA.n3514 0.0514167
R18991 GNDA.n3525 GNDA.n3524 0.0514167
R18992 GNDA.n3531 GNDA.n3530 0.0514167
R18993 GNDA.n3539 GNDA.n566 0.0514167
R18994 GNDA.n3470 GNDA.n3469 0.0514167
R18995 GNDA.n3464 GNDA.n3463 0.0514167
R18996 GNDA.n3461 GNDA.n3460 0.0514167
R18997 GNDA.n3455 GNDA.n3454 0.0514167
R18998 GNDA.n3452 GNDA.n3451 0.0514167
R18999 GNDA.n3446 GNDA.n3445 0.0514167
R19000 GNDA.n3443 GNDA.n3442 0.0514167
R19001 GNDA.n3437 GNDA.n3436 0.0514167
R19002 GNDA.n3251 GNDA.n594 0.0514167
R19003 GNDA.n3261 GNDA.n3260 0.0514167
R19004 GNDA.n3267 GNDA.n3266 0.0514167
R19005 GNDA.n3277 GNDA.n3276 0.0514167
R19006 GNDA.n3281 GNDA.n3280 0.0514167
R19007 GNDA.n3291 GNDA.n3290 0.0514167
R19008 GNDA.n3297 GNDA.n3296 0.0514167
R19009 GNDA.n3305 GNDA.n606 0.0514167
R19010 GNDA.n3236 GNDA.n3235 0.0514167
R19011 GNDA.n3230 GNDA.n3229 0.0514167
R19012 GNDA.n3227 GNDA.n3226 0.0514167
R19013 GNDA.n3221 GNDA.n3220 0.0514167
R19014 GNDA.n3218 GNDA.n3217 0.0514167
R19015 GNDA.n3212 GNDA.n3211 0.0514167
R19016 GNDA.n3209 GNDA.n3208 0.0514167
R19017 GNDA.n3203 GNDA.n3202 0.0514167
R19018 GNDA.n1601 GNDA.n1575 0.0514167
R19019 GNDA.n1611 GNDA.n1610 0.0514167
R19020 GNDA.n1617 GNDA.n1616 0.0514167
R19021 GNDA.n1627 GNDA.n1626 0.0514167
R19022 GNDA.n1631 GNDA.n1630 0.0514167
R19023 GNDA.n1641 GNDA.n1640 0.0514167
R19024 GNDA.n1647 GNDA.n1646 0.0514167
R19025 GNDA.n1655 GNDA.n1587 0.0514167
R19026 GNDA.n1519 GNDA.n1493 0.0514167
R19027 GNDA.n1529 GNDA.n1528 0.0514167
R19028 GNDA.n1535 GNDA.n1534 0.0514167
R19029 GNDA.n1545 GNDA.n1544 0.0514167
R19030 GNDA.n1549 GNDA.n1548 0.0514167
R19031 GNDA.n1559 GNDA.n1558 0.0514167
R19032 GNDA.n1565 GNDA.n1564 0.0514167
R19033 GNDA.n1573 GNDA.n1505 0.0514167
R19034 GNDA.n1437 GNDA.n1411 0.0514167
R19035 GNDA.n1447 GNDA.n1446 0.0514167
R19036 GNDA.n1453 GNDA.n1452 0.0514167
R19037 GNDA.n1463 GNDA.n1462 0.0514167
R19038 GNDA.n1467 GNDA.n1466 0.0514167
R19039 GNDA.n1477 GNDA.n1476 0.0514167
R19040 GNDA.n1483 GNDA.n1482 0.0514167
R19041 GNDA.n1491 GNDA.n1423 0.0514167
R19042 GNDA.n1247 GNDA.n1246 0.0514167
R19043 GNDA.n1241 GNDA.n1240 0.0514167
R19044 GNDA.n1238 GNDA.n1237 0.0514167
R19045 GNDA.n1232 GNDA.n1231 0.0514167
R19046 GNDA.n1229 GNDA.n1228 0.0514167
R19047 GNDA.n1223 GNDA.n1222 0.0514167
R19048 GNDA.n1220 GNDA.n1219 0.0514167
R19049 GNDA.n1214 GNDA.n1213 0.0514167
R19050 GNDA.n1869 GNDA.n1141 0.0514167
R19051 GNDA.n1879 GNDA.n1878 0.0514167
R19052 GNDA.n1885 GNDA.n1884 0.0514167
R19053 GNDA.n1895 GNDA.n1894 0.0514167
R19054 GNDA.n1899 GNDA.n1898 0.0514167
R19055 GNDA.n1909 GNDA.n1908 0.0514167
R19056 GNDA.n1915 GNDA.n1914 0.0514167
R19057 GNDA.n1923 GNDA.n1154 0.0514167
R19058 GNDA.n2162 GNDA.n2128 0.0514167
R19059 GNDA.n2170 GNDA.n2169 0.0514167
R19060 GNDA.n2157 GNDA.n2156 0.0514167
R19061 GNDA.n2153 GNDA.n2152 0.0514167
R19062 GNDA.n2186 GNDA.n2185 0.0514167
R19063 GNDA.n2194 GNDA.n2193 0.0514167
R19064 GNDA.n2145 GNDA.n2144 0.0514167
R19065 GNDA.n2220 GNDA.n2140 0.0514167
R19066 GNDA.n2076 GNDA.n2053 0.0514167
R19067 GNDA.n2086 GNDA.n2085 0.0514167
R19068 GNDA.n2090 GNDA.n2089 0.0514167
R19069 GNDA.n2100 GNDA.n2099 0.0514167
R19070 GNDA.n2106 GNDA.n2105 0.0514167
R19071 GNDA.n2116 GNDA.n2115 0.0514167
R19072 GNDA.n2120 GNDA.n2119 0.0514167
R19073 GNDA.n2223 GNDA.n845 0.0514167
R19074 GNDA.n1781 GNDA.n1780 0.0475
R19075 GNDA.n1791 GNDA.n1790 0.0475
R19076 GNDA.n1799 GNDA.n1798 0.0475
R19077 GNDA.n1302 GNDA.n1300 0.0421667
R19078 GNDA.n1265 GNDA.n628 0.0421667
R19079 GNDA.n1336 GNDA.n1334 0.0421667
R19080 GNDA.n1362 GNDA.n1263 0.0421667
R19081 GNDA.n1257 GNDA.n1255 0.0421667
R19082 GNDA.n1298 GNDA.n1293 0.0421667
R19083 GNDA.n3946 GNDA.n3944 0.0421667
R19084 GNDA.n1737 GNDA.n1736 0.0421667
R19085 GNDA.n1851 GNDA.n1844 0.0421667
R19086 GNDA.n1856 GNDA.n1841 0.0421667
R19087 GNDA.n1861 GNDA.n1770 0.0421667
R19088 GNDA.n1768 GNDA.n1767 0.0421667
R19089 GNDA.n1764 GNDA.n1763 0.0421667
R19090 GNDA.n1760 GNDA.n1759 0.0421667
R19091 GNDA.n1756 GNDA.n1755 0.0421667
R19092 GNDA.n1752 GNDA.n1751 0.0421667
R19093 GNDA.n1740 GNDA.n1739 0.0421667
R19094 GNDA.n3243 GNDA.n621 0.0421667
R19095 GNDA.n619 GNDA.n588 0.0421667
R19096 GNDA.n3390 GNDA.n584 0.0421667
R19097 GNDA.n3477 GNDA.n581 0.0421667
R19098 GNDA.n579 GNDA.n548 0.0421667
R19099 GNDA.n3624 GNDA.n545 0.0421667
R19100 GNDA.n3711 GNDA.n541 0.0421667
R19101 GNDA.n539 GNDA.n508 0.0421667
R19102 GNDA.n3858 GNDA.n505 0.0421667
R19103 GNDA.n503 GNDA.n437 0.0421667
R19104 GNDA.n4615 GNDA.n4614 0.0421667
R19105 GNDA.n4611 GNDA.n4610 0.0421667
R19106 GNDA.n4607 GNDA.n4606 0.0421667
R19107 GNDA.n4603 GNDA.n4602 0.0421667
R19108 GNDA.n4599 GNDA.n4598 0.0421667
R19109 GNDA.n4595 GNDA.n4594 0.0421667
R19110 GNDA.n4591 GNDA.n4590 0.0421667
R19111 GNDA.n4587 GNDA.n4586 0.0421667
R19112 GNDA.n2282 GNDA.n703 0.0421667
R19113 GNDA.n2215 GNDA.n2214 0.0421667
R19114 GNDA.n3630 GNDA.n3629 0.028198
R19115 GNDA.n3635 GNDA.n3634 0.028198
R19116 GNDA.n3643 GNDA.n3642 0.028198
R19117 GNDA.n3646 GNDA.n3645 0.028198
R19118 GNDA.n3654 GNDA.n3653 0.028198
R19119 GNDA.n3659 GNDA.n3658 0.028198
R19120 GNDA.n3667 GNDA.n3666 0.028198
R19121 GNDA.n3670 GNDA.n3669 0.028198
R19122 GNDA.n3332 GNDA.n3307 0.028198
R19123 GNDA.n3336 GNDA.n3308 0.028198
R19124 GNDA.n3346 GNDA.n3310 0.028198
R19125 GNDA.n3352 GNDA.n3311 0.028198
R19126 GNDA.n3362 GNDA.n3313 0.028198
R19127 GNDA.n3366 GNDA.n3314 0.028198
R19128 GNDA.n3376 GNDA.n3316 0.028198
R19129 GNDA.n3318 GNDA.n3317 0.028198
R19130 GNDA.n4529 GNDA.n4504 0.028198
R19131 GNDA.n4533 GNDA.n4505 0.028198
R19132 GNDA.n4543 GNDA.n4507 0.028198
R19133 GNDA.n4549 GNDA.n4508 0.028198
R19134 GNDA.n4559 GNDA.n4510 0.028198
R19135 GNDA.n4563 GNDA.n4511 0.028198
R19136 GNDA.n4573 GNDA.n4513 0.028198
R19137 GNDA.n4515 GNDA.n4514 0.028198
R19138 GNDA.n4453 GNDA.n4423 0.028198
R19139 GNDA.n4457 GNDA.n4424 0.028198
R19140 GNDA.n4467 GNDA.n4426 0.028198
R19141 GNDA.n4473 GNDA.n4427 0.028198
R19142 GNDA.n4483 GNDA.n4429 0.028198
R19143 GNDA.n4487 GNDA.n4430 0.028198
R19144 GNDA.n4497 GNDA.n4432 0.028198
R19145 GNDA.n4434 GNDA.n4433 0.028198
R19146 GNDA.n4371 GNDA.n4341 0.028198
R19147 GNDA.n4375 GNDA.n4342 0.028198
R19148 GNDA.n4385 GNDA.n4344 0.028198
R19149 GNDA.n4391 GNDA.n4345 0.028198
R19150 GNDA.n4401 GNDA.n4347 0.028198
R19151 GNDA.n4405 GNDA.n4348 0.028198
R19152 GNDA.n4415 GNDA.n4350 0.028198
R19153 GNDA.n4352 GNDA.n4351 0.028198
R19154 GNDA.n4289 GNDA.n4259 0.028198
R19155 GNDA.n4293 GNDA.n4260 0.028198
R19156 GNDA.n4303 GNDA.n4262 0.028198
R19157 GNDA.n4309 GNDA.n4263 0.028198
R19158 GNDA.n4319 GNDA.n4265 0.028198
R19159 GNDA.n4323 GNDA.n4266 0.028198
R19160 GNDA.n4333 GNDA.n4268 0.028198
R19161 GNDA.n4270 GNDA.n4269 0.028198
R19162 GNDA.n4207 GNDA.n4177 0.028198
R19163 GNDA.n4211 GNDA.n4178 0.028198
R19164 GNDA.n4221 GNDA.n4180 0.028198
R19165 GNDA.n4227 GNDA.n4181 0.028198
R19166 GNDA.n4237 GNDA.n4183 0.028198
R19167 GNDA.n4241 GNDA.n4184 0.028198
R19168 GNDA.n4251 GNDA.n4186 0.028198
R19169 GNDA.n4188 GNDA.n4187 0.028198
R19170 GNDA.n3961 GNDA.n479 0.028198
R19171 GNDA.n3965 GNDA.n480 0.028198
R19172 GNDA.n3975 GNDA.n482 0.028198
R19173 GNDA.n3981 GNDA.n483 0.028198
R19174 GNDA.n3991 GNDA.n485 0.028198
R19175 GNDA.n3995 GNDA.n486 0.028198
R19176 GNDA.n4005 GNDA.n488 0.028198
R19177 GNDA.n490 GNDA.n489 0.028198
R19178 GNDA.n4125 GNDA.n4095 0.028198
R19179 GNDA.n4129 GNDA.n4096 0.028198
R19180 GNDA.n4139 GNDA.n4098 0.028198
R19181 GNDA.n4145 GNDA.n4099 0.028198
R19182 GNDA.n4155 GNDA.n4101 0.028198
R19183 GNDA.n4159 GNDA.n4102 0.028198
R19184 GNDA.n4169 GNDA.n4104 0.028198
R19185 GNDA.n4106 GNDA.n4105 0.028198
R19186 GNDA.n4043 GNDA.n4013 0.028198
R19187 GNDA.n4047 GNDA.n4014 0.028198
R19188 GNDA.n4057 GNDA.n4016 0.028198
R19189 GNDA.n4063 GNDA.n4017 0.028198
R19190 GNDA.n4073 GNDA.n4019 0.028198
R19191 GNDA.n4077 GNDA.n4020 0.028198
R19192 GNDA.n4087 GNDA.n4022 0.028198
R19193 GNDA.n4024 GNDA.n4023 0.028198
R19194 GNDA.n3939 GNDA.n3938 0.028198
R19195 GNDA.n3936 GNDA.n3935 0.028198
R19196 GNDA.n3930 GNDA.n3929 0.028198
R19197 GNDA.n3927 GNDA.n3926 0.028198
R19198 GNDA.n3921 GNDA.n3920 0.028198
R19199 GNDA.n3918 GNDA.n3917 0.028198
R19200 GNDA.n3912 GNDA.n3911 0.028198
R19201 GNDA.n3909 GNDA.n3908 0.028198
R19202 GNDA.n1682 GNDA.n1657 0.028198
R19203 GNDA.n1686 GNDA.n1658 0.028198
R19204 GNDA.n1696 GNDA.n1660 0.028198
R19205 GNDA.n1702 GNDA.n1661 0.028198
R19206 GNDA.n1712 GNDA.n1663 0.028198
R19207 GNDA.n1716 GNDA.n1664 0.028198
R19208 GNDA.n1726 GNDA.n1666 0.028198
R19209 GNDA.n1668 GNDA.n1667 0.028198
R19210 GNDA.n3800 GNDA.n3775 0.028198
R19211 GNDA.n3804 GNDA.n3776 0.028198
R19212 GNDA.n3814 GNDA.n3778 0.028198
R19213 GNDA.n3820 GNDA.n3779 0.028198
R19214 GNDA.n3830 GNDA.n3781 0.028198
R19215 GNDA.n3834 GNDA.n3782 0.028198
R19216 GNDA.n3844 GNDA.n3784 0.028198
R19217 GNDA.n3786 GNDA.n3785 0.028198
R19218 GNDA.n3724 GNDA.n515 0.028198
R19219 GNDA.n3728 GNDA.n516 0.028198
R19220 GNDA.n3738 GNDA.n518 0.028198
R19221 GNDA.n3744 GNDA.n519 0.028198
R19222 GNDA.n3754 GNDA.n521 0.028198
R19223 GNDA.n3758 GNDA.n522 0.028198
R19224 GNDA.n3768 GNDA.n524 0.028198
R19225 GNDA.n526 GNDA.n525 0.028198
R19226 GNDA.n3566 GNDA.n3541 0.028198
R19227 GNDA.n3570 GNDA.n3542 0.028198
R19228 GNDA.n3580 GNDA.n3544 0.028198
R19229 GNDA.n3586 GNDA.n3545 0.028198
R19230 GNDA.n3596 GNDA.n3547 0.028198
R19231 GNDA.n3600 GNDA.n3548 0.028198
R19232 GNDA.n3610 GNDA.n3550 0.028198
R19233 GNDA.n3552 GNDA.n3551 0.028198
R19234 GNDA.n3490 GNDA.n555 0.028198
R19235 GNDA.n3494 GNDA.n556 0.028198
R19236 GNDA.n3504 GNDA.n558 0.028198
R19237 GNDA.n3510 GNDA.n559 0.028198
R19238 GNDA.n3520 GNDA.n561 0.028198
R19239 GNDA.n3524 GNDA.n562 0.028198
R19240 GNDA.n3534 GNDA.n564 0.028198
R19241 GNDA.n566 GNDA.n565 0.028198
R19242 GNDA.n3468 GNDA.n3467 0.028198
R19243 GNDA.n3465 GNDA.n3464 0.028198
R19244 GNDA.n3459 GNDA.n3458 0.028198
R19245 GNDA.n3456 GNDA.n3455 0.028198
R19246 GNDA.n3450 GNDA.n3449 0.028198
R19247 GNDA.n3447 GNDA.n3446 0.028198
R19248 GNDA.n3441 GNDA.n3440 0.028198
R19249 GNDA.n3438 GNDA.n3437 0.028198
R19250 GNDA.n3256 GNDA.n595 0.028198
R19251 GNDA.n3260 GNDA.n596 0.028198
R19252 GNDA.n3270 GNDA.n598 0.028198
R19253 GNDA.n3276 GNDA.n599 0.028198
R19254 GNDA.n3286 GNDA.n601 0.028198
R19255 GNDA.n3290 GNDA.n602 0.028198
R19256 GNDA.n3300 GNDA.n604 0.028198
R19257 GNDA.n606 GNDA.n605 0.028198
R19258 GNDA.n3234 GNDA.n3233 0.028198
R19259 GNDA.n3231 GNDA.n3230 0.028198
R19260 GNDA.n3225 GNDA.n3224 0.028198
R19261 GNDA.n3222 GNDA.n3221 0.028198
R19262 GNDA.n3216 GNDA.n3215 0.028198
R19263 GNDA.n3213 GNDA.n3212 0.028198
R19264 GNDA.n3207 GNDA.n3206 0.028198
R19265 GNDA.n3204 GNDA.n3203 0.028198
R19266 GNDA.n1606 GNDA.n1576 0.028198
R19267 GNDA.n1610 GNDA.n1577 0.028198
R19268 GNDA.n1620 GNDA.n1579 0.028198
R19269 GNDA.n1626 GNDA.n1580 0.028198
R19270 GNDA.n1636 GNDA.n1582 0.028198
R19271 GNDA.n1640 GNDA.n1583 0.028198
R19272 GNDA.n1650 GNDA.n1585 0.028198
R19273 GNDA.n1587 GNDA.n1586 0.028198
R19274 GNDA.n1524 GNDA.n1494 0.028198
R19275 GNDA.n1528 GNDA.n1495 0.028198
R19276 GNDA.n1538 GNDA.n1497 0.028198
R19277 GNDA.n1544 GNDA.n1498 0.028198
R19278 GNDA.n1554 GNDA.n1500 0.028198
R19279 GNDA.n1558 GNDA.n1501 0.028198
R19280 GNDA.n1568 GNDA.n1503 0.028198
R19281 GNDA.n1505 GNDA.n1504 0.028198
R19282 GNDA.n1442 GNDA.n1412 0.028198
R19283 GNDA.n1446 GNDA.n1413 0.028198
R19284 GNDA.n1456 GNDA.n1415 0.028198
R19285 GNDA.n1462 GNDA.n1416 0.028198
R19286 GNDA.n1472 GNDA.n1418 0.028198
R19287 GNDA.n1476 GNDA.n1419 0.028198
R19288 GNDA.n1486 GNDA.n1421 0.028198
R19289 GNDA.n1423 GNDA.n1422 0.028198
R19290 GNDA.n1245 GNDA.n1244 0.028198
R19291 GNDA.n1242 GNDA.n1241 0.028198
R19292 GNDA.n1236 GNDA.n1235 0.028198
R19293 GNDA.n1233 GNDA.n1232 0.028198
R19294 GNDA.n1227 GNDA.n1226 0.028198
R19295 GNDA.n1224 GNDA.n1223 0.028198
R19296 GNDA.n1218 GNDA.n1217 0.028198
R19297 GNDA.n1215 GNDA.n1214 0.028198
R19298 GNDA.n1874 GNDA.n1142 0.028198
R19299 GNDA.n1878 GNDA.n1143 0.028198
R19300 GNDA.n1888 GNDA.n1145 0.028198
R19301 GNDA.n1894 GNDA.n1146 0.028198
R19302 GNDA.n1904 GNDA.n1148 0.028198
R19303 GNDA.n1908 GNDA.n1149 0.028198
R19304 GNDA.n1918 GNDA.n1151 0.028198
R19305 GNDA.n1154 GNDA.n1152 0.028198
R19306 GNDA.n1919 GNDA.n1152 0.028198
R19307 GNDA.n1915 GNDA.n1151 0.028198
R19308 GNDA.n1905 GNDA.n1149 0.028198
R19309 GNDA.n1899 GNDA.n1148 0.028198
R19310 GNDA.n1889 GNDA.n1146 0.028198
R19311 GNDA.n1885 GNDA.n1145 0.028198
R19312 GNDA.n1875 GNDA.n1143 0.028198
R19313 GNDA.n1869 GNDA.n1142 0.028198
R19314 GNDA.n1216 GNDA.n1215 0.028198
R19315 GNDA.n1219 GNDA.n1218 0.028198
R19316 GNDA.n1225 GNDA.n1224 0.028198
R19317 GNDA.n1228 GNDA.n1227 0.028198
R19318 GNDA.n1234 GNDA.n1233 0.028198
R19319 GNDA.n1237 GNDA.n1236 0.028198
R19320 GNDA.n1243 GNDA.n1242 0.028198
R19321 GNDA.n1246 GNDA.n1245 0.028198
R19322 GNDA.n1487 GNDA.n1422 0.028198
R19323 GNDA.n1483 GNDA.n1421 0.028198
R19324 GNDA.n1473 GNDA.n1419 0.028198
R19325 GNDA.n1467 GNDA.n1418 0.028198
R19326 GNDA.n1457 GNDA.n1416 0.028198
R19327 GNDA.n1453 GNDA.n1415 0.028198
R19328 GNDA.n1443 GNDA.n1413 0.028198
R19329 GNDA.n1437 GNDA.n1412 0.028198
R19330 GNDA.n1569 GNDA.n1504 0.028198
R19331 GNDA.n1565 GNDA.n1503 0.028198
R19332 GNDA.n1555 GNDA.n1501 0.028198
R19333 GNDA.n1549 GNDA.n1500 0.028198
R19334 GNDA.n1539 GNDA.n1498 0.028198
R19335 GNDA.n1535 GNDA.n1497 0.028198
R19336 GNDA.n1525 GNDA.n1495 0.028198
R19337 GNDA.n1519 GNDA.n1494 0.028198
R19338 GNDA.n1651 GNDA.n1586 0.028198
R19339 GNDA.n1647 GNDA.n1585 0.028198
R19340 GNDA.n1637 GNDA.n1583 0.028198
R19341 GNDA.n1631 GNDA.n1582 0.028198
R19342 GNDA.n1621 GNDA.n1580 0.028198
R19343 GNDA.n1617 GNDA.n1579 0.028198
R19344 GNDA.n1607 GNDA.n1577 0.028198
R19345 GNDA.n1601 GNDA.n1576 0.028198
R19346 GNDA.n3205 GNDA.n3204 0.028198
R19347 GNDA.n3208 GNDA.n3207 0.028198
R19348 GNDA.n3214 GNDA.n3213 0.028198
R19349 GNDA.n3217 GNDA.n3216 0.028198
R19350 GNDA.n3223 GNDA.n3222 0.028198
R19351 GNDA.n3226 GNDA.n3225 0.028198
R19352 GNDA.n3232 GNDA.n3231 0.028198
R19353 GNDA.n3235 GNDA.n3234 0.028198
R19354 GNDA.n3301 GNDA.n605 0.028198
R19355 GNDA.n3297 GNDA.n604 0.028198
R19356 GNDA.n3287 GNDA.n602 0.028198
R19357 GNDA.n3281 GNDA.n601 0.028198
R19358 GNDA.n3271 GNDA.n599 0.028198
R19359 GNDA.n3267 GNDA.n598 0.028198
R19360 GNDA.n3257 GNDA.n596 0.028198
R19361 GNDA.n3251 GNDA.n595 0.028198
R19362 GNDA.n3439 GNDA.n3438 0.028198
R19363 GNDA.n3442 GNDA.n3441 0.028198
R19364 GNDA.n3448 GNDA.n3447 0.028198
R19365 GNDA.n3451 GNDA.n3450 0.028198
R19366 GNDA.n3457 GNDA.n3456 0.028198
R19367 GNDA.n3460 GNDA.n3459 0.028198
R19368 GNDA.n3466 GNDA.n3465 0.028198
R19369 GNDA.n3469 GNDA.n3468 0.028198
R19370 GNDA.n3535 GNDA.n565 0.028198
R19371 GNDA.n3531 GNDA.n564 0.028198
R19372 GNDA.n3521 GNDA.n562 0.028198
R19373 GNDA.n3515 GNDA.n561 0.028198
R19374 GNDA.n3505 GNDA.n559 0.028198
R19375 GNDA.n3501 GNDA.n558 0.028198
R19376 GNDA.n3491 GNDA.n556 0.028198
R19377 GNDA.n3485 GNDA.n555 0.028198
R19378 GNDA.n3611 GNDA.n3551 0.028198
R19379 GNDA.n3607 GNDA.n3550 0.028198
R19380 GNDA.n3597 GNDA.n3548 0.028198
R19381 GNDA.n3591 GNDA.n3547 0.028198
R19382 GNDA.n3581 GNDA.n3545 0.028198
R19383 GNDA.n3577 GNDA.n3544 0.028198
R19384 GNDA.n3567 GNDA.n3542 0.028198
R19385 GNDA.n3541 GNDA.n552 0.028198
R19386 GNDA.n3769 GNDA.n525 0.028198
R19387 GNDA.n3765 GNDA.n524 0.028198
R19388 GNDA.n3755 GNDA.n522 0.028198
R19389 GNDA.n3749 GNDA.n521 0.028198
R19390 GNDA.n3739 GNDA.n519 0.028198
R19391 GNDA.n3735 GNDA.n518 0.028198
R19392 GNDA.n3725 GNDA.n516 0.028198
R19393 GNDA.n3719 GNDA.n515 0.028198
R19394 GNDA.n3845 GNDA.n3785 0.028198
R19395 GNDA.n3841 GNDA.n3784 0.028198
R19396 GNDA.n3831 GNDA.n3782 0.028198
R19397 GNDA.n3825 GNDA.n3781 0.028198
R19398 GNDA.n3815 GNDA.n3779 0.028198
R19399 GNDA.n3811 GNDA.n3778 0.028198
R19400 GNDA.n3801 GNDA.n3776 0.028198
R19401 GNDA.n3775 GNDA.n512 0.028198
R19402 GNDA.n1727 GNDA.n1667 0.028198
R19403 GNDA.n1723 GNDA.n1666 0.028198
R19404 GNDA.n1713 GNDA.n1664 0.028198
R19405 GNDA.n1707 GNDA.n1663 0.028198
R19406 GNDA.n1697 GNDA.n1661 0.028198
R19407 GNDA.n1693 GNDA.n1660 0.028198
R19408 GNDA.n1683 GNDA.n1658 0.028198
R19409 GNDA.n1657 GNDA.n1410 0.028198
R19410 GNDA.n3910 GNDA.n3909 0.028198
R19411 GNDA.n3913 GNDA.n3912 0.028198
R19412 GNDA.n3919 GNDA.n3918 0.028198
R19413 GNDA.n3922 GNDA.n3921 0.028198
R19414 GNDA.n3928 GNDA.n3927 0.028198
R19415 GNDA.n3931 GNDA.n3930 0.028198
R19416 GNDA.n3937 GNDA.n3936 0.028198
R19417 GNDA.n3940 GNDA.n3939 0.028198
R19418 GNDA.n4088 GNDA.n4023 0.028198
R19419 GNDA.n4084 GNDA.n4022 0.028198
R19420 GNDA.n4074 GNDA.n4020 0.028198
R19421 GNDA.n4068 GNDA.n4019 0.028198
R19422 GNDA.n4058 GNDA.n4017 0.028198
R19423 GNDA.n4054 GNDA.n4016 0.028198
R19424 GNDA.n4044 GNDA.n4014 0.028198
R19425 GNDA.n4038 GNDA.n4013 0.028198
R19426 GNDA.n4170 GNDA.n4105 0.028198
R19427 GNDA.n4166 GNDA.n4104 0.028198
R19428 GNDA.n4156 GNDA.n4102 0.028198
R19429 GNDA.n4150 GNDA.n4101 0.028198
R19430 GNDA.n4140 GNDA.n4099 0.028198
R19431 GNDA.n4136 GNDA.n4098 0.028198
R19432 GNDA.n4126 GNDA.n4096 0.028198
R19433 GNDA.n4120 GNDA.n4095 0.028198
R19434 GNDA.n4006 GNDA.n489 0.028198
R19435 GNDA.n4002 GNDA.n488 0.028198
R19436 GNDA.n3992 GNDA.n486 0.028198
R19437 GNDA.n3986 GNDA.n485 0.028198
R19438 GNDA.n3976 GNDA.n483 0.028198
R19439 GNDA.n3972 GNDA.n482 0.028198
R19440 GNDA.n3962 GNDA.n480 0.028198
R19441 GNDA.n3956 GNDA.n479 0.028198
R19442 GNDA.n4252 GNDA.n4187 0.028198
R19443 GNDA.n4248 GNDA.n4186 0.028198
R19444 GNDA.n4238 GNDA.n4184 0.028198
R19445 GNDA.n4232 GNDA.n4183 0.028198
R19446 GNDA.n4222 GNDA.n4181 0.028198
R19447 GNDA.n4218 GNDA.n4180 0.028198
R19448 GNDA.n4208 GNDA.n4178 0.028198
R19449 GNDA.n4202 GNDA.n4177 0.028198
R19450 GNDA.n4334 GNDA.n4269 0.028198
R19451 GNDA.n4330 GNDA.n4268 0.028198
R19452 GNDA.n4320 GNDA.n4266 0.028198
R19453 GNDA.n4314 GNDA.n4265 0.028198
R19454 GNDA.n4304 GNDA.n4263 0.028198
R19455 GNDA.n4300 GNDA.n4262 0.028198
R19456 GNDA.n4290 GNDA.n4260 0.028198
R19457 GNDA.n4284 GNDA.n4259 0.028198
R19458 GNDA.n4416 GNDA.n4351 0.028198
R19459 GNDA.n4412 GNDA.n4350 0.028198
R19460 GNDA.n4402 GNDA.n4348 0.028198
R19461 GNDA.n4396 GNDA.n4347 0.028198
R19462 GNDA.n4386 GNDA.n4345 0.028198
R19463 GNDA.n4382 GNDA.n4344 0.028198
R19464 GNDA.n4372 GNDA.n4342 0.028198
R19465 GNDA.n4366 GNDA.n4341 0.028198
R19466 GNDA.n4498 GNDA.n4433 0.028198
R19467 GNDA.n4494 GNDA.n4432 0.028198
R19468 GNDA.n4484 GNDA.n4430 0.028198
R19469 GNDA.n4478 GNDA.n4429 0.028198
R19470 GNDA.n4468 GNDA.n4427 0.028198
R19471 GNDA.n4464 GNDA.n4426 0.028198
R19472 GNDA.n4454 GNDA.n4424 0.028198
R19473 GNDA.n4448 GNDA.n4423 0.028198
R19474 GNDA.n4574 GNDA.n4514 0.028198
R19475 GNDA.n4570 GNDA.n4513 0.028198
R19476 GNDA.n4560 GNDA.n4511 0.028198
R19477 GNDA.n4554 GNDA.n4510 0.028198
R19478 GNDA.n4544 GNDA.n4508 0.028198
R19479 GNDA.n4540 GNDA.n4507 0.028198
R19480 GNDA.n4530 GNDA.n4505 0.028198
R19481 GNDA.n4504 GNDA.n476 0.028198
R19482 GNDA.n3377 GNDA.n3317 0.028198
R19483 GNDA.n3373 GNDA.n3316 0.028198
R19484 GNDA.n3363 GNDA.n3314 0.028198
R19485 GNDA.n3357 GNDA.n3313 0.028198
R19486 GNDA.n3347 GNDA.n3311 0.028198
R19487 GNDA.n3343 GNDA.n3310 0.028198
R19488 GNDA.n3333 GNDA.n3308 0.028198
R19489 GNDA.n3307 GNDA.n592 0.028198
R19490 GNDA.n3669 GNDA.n3668 0.028198
R19491 GNDA.n3666 GNDA.n3665 0.028198
R19492 GNDA.n3658 GNDA.n3657 0.028198
R19493 GNDA.n3653 GNDA.n3652 0.028198
R19494 GNDA.n3645 GNDA.n3644 0.028198
R19495 GNDA.n3642 GNDA.n3641 0.028198
R19496 GNDA.n3634 GNDA.n3633 0.028198
R19497 GNDA.n3629 GNDA.n3628 0.028198
R19498 GNDA.n2160 GNDA.n2129 0.028198
R19499 GNDA.n2169 GNDA.n2130 0.028198
R19500 GNDA.n2177 GNDA.n2132 0.028198
R19501 GNDA.n2152 GNDA.n2133 0.028198
R19502 GNDA.n2148 GNDA.n2135 0.028198
R19503 GNDA.n2193 GNDA.n2136 0.028198
R19504 GNDA.n2201 GNDA.n2138 0.028198
R19505 GNDA.n2140 GNDA.n2139 0.028198
R19506 GNDA.n2079 GNDA.n2054 0.028198
R19507 GNDA.n2085 GNDA.n2055 0.028198
R19508 GNDA.n2095 GNDA.n2057 0.028198
R19509 GNDA.n2099 GNDA.n2058 0.028198
R19510 GNDA.n2109 GNDA.n2060 0.028198
R19511 GNDA.n2115 GNDA.n2061 0.028198
R19512 GNDA.n2064 GNDA.n2063 0.028198
R19513 GNDA.n2127 GNDA.n845 0.028198
R19514 GNDA.n2127 GNDA.n2126 0.028198
R19515 GNDA.n2120 GNDA.n2063 0.028198
R19516 GNDA.n2110 GNDA.n2061 0.028198
R19517 GNDA.n2106 GNDA.n2060 0.028198
R19518 GNDA.n2096 GNDA.n2058 0.028198
R19519 GNDA.n2090 GNDA.n2057 0.028198
R19520 GNDA.n2080 GNDA.n2055 0.028198
R19521 GNDA.n2076 GNDA.n2054 0.028198
R19522 GNDA.n2202 GNDA.n2139 0.028198
R19523 GNDA.n2145 GNDA.n2138 0.028198
R19524 GNDA.n2149 GNDA.n2136 0.028198
R19525 GNDA.n2186 GNDA.n2135 0.028198
R19526 GNDA.n2178 GNDA.n2133 0.028198
R19527 GNDA.n2157 GNDA.n2132 0.028198
R19528 GNDA.n2161 GNDA.n2130 0.028198
R19529 GNDA.n2162 GNDA.n2129 0.028198
R19530 GNDA.n1775 GNDA.n1131 0.028198
R19531 GNDA.n1785 GNDA.n1134 0.028198
R19532 GNDA.n1793 GNDA.n1137 0.028198
R19533 GNDA.n1803 GNDA.n1140 0.028198
R19534 GNDA.n1804 GNDA.n1140 0.028198
R19535 GNDA.n1796 GNDA.n1137 0.028198
R19536 GNDA.n1786 GNDA.n1134 0.028198
R19537 GNDA.n1778 GNDA.n1131 0.028198
R19538 GNDA.n1779 GNDA.n1132 0.0262697
R19539 GNDA.n1781 GNDA.n1133 0.0262697
R19540 GNDA.n1787 GNDA.n1135 0.0262697
R19541 GNDA.n1791 GNDA.n1136 0.0262697
R19542 GNDA.n1797 GNDA.n1138 0.0262697
R19543 GNDA.n1799 GNDA.n1139 0.0262697
R19544 GNDA.n1805 GNDA.n1129 0.0262697
R19545 GNDA.n1802 GNDA.n1139 0.0262697
R19546 GNDA.n1798 GNDA.n1138 0.0262697
R19547 GNDA.n1792 GNDA.n1136 0.0262697
R19548 GNDA.n1790 GNDA.n1135 0.0262697
R19549 GNDA.n1784 GNDA.n1133 0.0262697
R19550 GNDA.n1780 GNDA.n1132 0.0262697
R19551 GNDA.n1774 GNDA.n1130 0.0262697
R19552 GNDA.n3638 GNDA.n3637 0.0243392
R19553 GNDA.n3651 GNDA.n3650 0.0243392
R19554 GNDA.n3662 GNDA.n3661 0.0243392
R19555 GNDA.n3342 GNDA.n3309 0.0243392
R19556 GNDA.n3356 GNDA.n3312 0.0243392
R19557 GNDA.n3372 GNDA.n3315 0.0243392
R19558 GNDA.n4539 GNDA.n4506 0.0243392
R19559 GNDA.n4553 GNDA.n4509 0.0243392
R19560 GNDA.n4569 GNDA.n4512 0.0243392
R19561 GNDA.n4463 GNDA.n4425 0.0243392
R19562 GNDA.n4477 GNDA.n4428 0.0243392
R19563 GNDA.n4493 GNDA.n4431 0.0243392
R19564 GNDA.n4381 GNDA.n4343 0.0243392
R19565 GNDA.n4395 GNDA.n4346 0.0243392
R19566 GNDA.n4411 GNDA.n4349 0.0243392
R19567 GNDA.n4299 GNDA.n4261 0.0243392
R19568 GNDA.n4313 GNDA.n4264 0.0243392
R19569 GNDA.n4329 GNDA.n4267 0.0243392
R19570 GNDA.n4217 GNDA.n4179 0.0243392
R19571 GNDA.n4231 GNDA.n4182 0.0243392
R19572 GNDA.n4247 GNDA.n4185 0.0243392
R19573 GNDA.n3971 GNDA.n481 0.0243392
R19574 GNDA.n3985 GNDA.n484 0.0243392
R19575 GNDA.n4001 GNDA.n487 0.0243392
R19576 GNDA.n4135 GNDA.n4097 0.0243392
R19577 GNDA.n4149 GNDA.n4100 0.0243392
R19578 GNDA.n4165 GNDA.n4103 0.0243392
R19579 GNDA.n4053 GNDA.n4015 0.0243392
R19580 GNDA.n4067 GNDA.n4018 0.0243392
R19581 GNDA.n4083 GNDA.n4021 0.0243392
R19582 GNDA.n3933 GNDA.n3932 0.0243392
R19583 GNDA.n3924 GNDA.n3923 0.0243392
R19584 GNDA.n3915 GNDA.n3914 0.0243392
R19585 GNDA.n1692 GNDA.n1659 0.0243392
R19586 GNDA.n1706 GNDA.n1662 0.0243392
R19587 GNDA.n1722 GNDA.n1665 0.0243392
R19588 GNDA.n3810 GNDA.n3777 0.0243392
R19589 GNDA.n3824 GNDA.n3780 0.0243392
R19590 GNDA.n3840 GNDA.n3783 0.0243392
R19591 GNDA.n3734 GNDA.n517 0.0243392
R19592 GNDA.n3748 GNDA.n520 0.0243392
R19593 GNDA.n3764 GNDA.n523 0.0243392
R19594 GNDA.n3576 GNDA.n3543 0.0243392
R19595 GNDA.n3590 GNDA.n3546 0.0243392
R19596 GNDA.n3606 GNDA.n3549 0.0243392
R19597 GNDA.n3500 GNDA.n557 0.0243392
R19598 GNDA.n3514 GNDA.n560 0.0243392
R19599 GNDA.n3530 GNDA.n563 0.0243392
R19600 GNDA.n3462 GNDA.n3461 0.0243392
R19601 GNDA.n3453 GNDA.n3452 0.0243392
R19602 GNDA.n3444 GNDA.n3443 0.0243392
R19603 GNDA.n3266 GNDA.n597 0.0243392
R19604 GNDA.n3280 GNDA.n600 0.0243392
R19605 GNDA.n3296 GNDA.n603 0.0243392
R19606 GNDA.n3228 GNDA.n3227 0.0243392
R19607 GNDA.n3219 GNDA.n3218 0.0243392
R19608 GNDA.n3210 GNDA.n3209 0.0243392
R19609 GNDA.n1616 GNDA.n1578 0.0243392
R19610 GNDA.n1630 GNDA.n1581 0.0243392
R19611 GNDA.n1646 GNDA.n1584 0.0243392
R19612 GNDA.n1534 GNDA.n1496 0.0243392
R19613 GNDA.n1548 GNDA.n1499 0.0243392
R19614 GNDA.n1564 GNDA.n1502 0.0243392
R19615 GNDA.n1452 GNDA.n1414 0.0243392
R19616 GNDA.n1466 GNDA.n1417 0.0243392
R19617 GNDA.n1482 GNDA.n1420 0.0243392
R19618 GNDA.n1239 GNDA.n1238 0.0243392
R19619 GNDA.n1230 GNDA.n1229 0.0243392
R19620 GNDA.n1221 GNDA.n1220 0.0243392
R19621 GNDA.n1884 GNDA.n1144 0.0243392
R19622 GNDA.n1898 GNDA.n1147 0.0243392
R19623 GNDA.n1914 GNDA.n1150 0.0243392
R19624 GNDA.n1909 GNDA.n1150 0.0243392
R19625 GNDA.n1895 GNDA.n1147 0.0243392
R19626 GNDA.n1879 GNDA.n1144 0.0243392
R19627 GNDA.n1222 GNDA.n1221 0.0243392
R19628 GNDA.n1231 GNDA.n1230 0.0243392
R19629 GNDA.n1240 GNDA.n1239 0.0243392
R19630 GNDA.n1477 GNDA.n1420 0.0243392
R19631 GNDA.n1463 GNDA.n1417 0.0243392
R19632 GNDA.n1447 GNDA.n1414 0.0243392
R19633 GNDA.n1559 GNDA.n1502 0.0243392
R19634 GNDA.n1545 GNDA.n1499 0.0243392
R19635 GNDA.n1529 GNDA.n1496 0.0243392
R19636 GNDA.n1641 GNDA.n1584 0.0243392
R19637 GNDA.n1627 GNDA.n1581 0.0243392
R19638 GNDA.n1611 GNDA.n1578 0.0243392
R19639 GNDA.n3211 GNDA.n3210 0.0243392
R19640 GNDA.n3220 GNDA.n3219 0.0243392
R19641 GNDA.n3229 GNDA.n3228 0.0243392
R19642 GNDA.n3291 GNDA.n603 0.0243392
R19643 GNDA.n3277 GNDA.n600 0.0243392
R19644 GNDA.n3261 GNDA.n597 0.0243392
R19645 GNDA.n3445 GNDA.n3444 0.0243392
R19646 GNDA.n3454 GNDA.n3453 0.0243392
R19647 GNDA.n3463 GNDA.n3462 0.0243392
R19648 GNDA.n3525 GNDA.n563 0.0243392
R19649 GNDA.n3511 GNDA.n560 0.0243392
R19650 GNDA.n3495 GNDA.n557 0.0243392
R19651 GNDA.n3601 GNDA.n3549 0.0243392
R19652 GNDA.n3587 GNDA.n3546 0.0243392
R19653 GNDA.n3571 GNDA.n3543 0.0243392
R19654 GNDA.n3759 GNDA.n523 0.0243392
R19655 GNDA.n3745 GNDA.n520 0.0243392
R19656 GNDA.n3729 GNDA.n517 0.0243392
R19657 GNDA.n3835 GNDA.n3783 0.0243392
R19658 GNDA.n3821 GNDA.n3780 0.0243392
R19659 GNDA.n3805 GNDA.n3777 0.0243392
R19660 GNDA.n1717 GNDA.n1665 0.0243392
R19661 GNDA.n1703 GNDA.n1662 0.0243392
R19662 GNDA.n1687 GNDA.n1659 0.0243392
R19663 GNDA.n3916 GNDA.n3915 0.0243392
R19664 GNDA.n3925 GNDA.n3924 0.0243392
R19665 GNDA.n3934 GNDA.n3933 0.0243392
R19666 GNDA.n4078 GNDA.n4021 0.0243392
R19667 GNDA.n4064 GNDA.n4018 0.0243392
R19668 GNDA.n4048 GNDA.n4015 0.0243392
R19669 GNDA.n4160 GNDA.n4103 0.0243392
R19670 GNDA.n4146 GNDA.n4100 0.0243392
R19671 GNDA.n4130 GNDA.n4097 0.0243392
R19672 GNDA.n3996 GNDA.n487 0.0243392
R19673 GNDA.n3982 GNDA.n484 0.0243392
R19674 GNDA.n3966 GNDA.n481 0.0243392
R19675 GNDA.n4242 GNDA.n4185 0.0243392
R19676 GNDA.n4228 GNDA.n4182 0.0243392
R19677 GNDA.n4212 GNDA.n4179 0.0243392
R19678 GNDA.n4324 GNDA.n4267 0.0243392
R19679 GNDA.n4310 GNDA.n4264 0.0243392
R19680 GNDA.n4294 GNDA.n4261 0.0243392
R19681 GNDA.n4406 GNDA.n4349 0.0243392
R19682 GNDA.n4392 GNDA.n4346 0.0243392
R19683 GNDA.n4376 GNDA.n4343 0.0243392
R19684 GNDA.n4488 GNDA.n4431 0.0243392
R19685 GNDA.n4474 GNDA.n4428 0.0243392
R19686 GNDA.n4458 GNDA.n4425 0.0243392
R19687 GNDA.n4564 GNDA.n4512 0.0243392
R19688 GNDA.n4550 GNDA.n4509 0.0243392
R19689 GNDA.n4534 GNDA.n4506 0.0243392
R19690 GNDA.n3367 GNDA.n3315 0.0243392
R19691 GNDA.n3353 GNDA.n3312 0.0243392
R19692 GNDA.n3337 GNDA.n3309 0.0243392
R19693 GNDA.n3661 GNDA.n3660 0.0243392
R19694 GNDA.n3650 GNDA.n3649 0.0243392
R19695 GNDA.n3637 GNDA.n3636 0.0243392
R19696 GNDA.n2156 GNDA.n2131 0.0243392
R19697 GNDA.n2185 GNDA.n2134 0.0243392
R19698 GNDA.n2144 GNDA.n2137 0.0243392
R19699 GNDA.n2089 GNDA.n2056 0.0243392
R19700 GNDA.n2105 GNDA.n2059 0.0243392
R19701 GNDA.n2119 GNDA.n2062 0.0243392
R19702 GNDA.n2116 GNDA.n2062 0.0243392
R19703 GNDA.n2100 GNDA.n2059 0.0243392
R19704 GNDA.n2086 GNDA.n2056 0.0243392
R19705 GNDA.n2194 GNDA.n2137 0.0243392
R19706 GNDA.n2153 GNDA.n2134 0.0243392
R19707 GNDA.n2170 GNDA.n2131 0.0243392
R19708 GNDA.n1303 GNDA.n1291 0.0217373
R19709 GNDA.n1296 GNDA.n1292 0.0217373
R19710 GNDA.n1297 GNDA.n1296 0.0217373
R19711 GNDA.n451 GNDA.n448 0.0217373
R19712 GNDA.n450 GNDA.n448 0.0217373
R19713 GNDA.n1317 GNDA.n1288 0.0217373
R19714 GNDA.n1301 GNDA.n1289 0.0217373
R19715 GNDA.n1291 GNDA.n1289 0.0217373
R19716 GNDA.n1265 GNDA.n1264 0.0217373
R19717 GNDA.n1337 GNDA.n1277 0.0217373
R19718 GNDA.n1329 GNDA.n1279 0.0217373
R19719 GNDA.n1324 GNDA.n1282 0.0217373
R19720 GNDA.n1287 GNDA.n1285 0.0217373
R19721 GNDA.n1331 GNDA.n1280 0.0217373
R19722 GNDA.n1330 GNDA.n1329 0.0217373
R19723 GNDA.n1326 GNDA.n1283 0.0217373
R19724 GNDA.n1325 GNDA.n1324 0.0217373
R19725 GNDA.n1288 GNDA.n1286 0.0217373
R19726 GNDA.n1343 GNDA.n1269 0.0217373
R19727 GNDA.n1335 GNDA.n1275 0.0217373
R19728 GNDA.n1277 GNDA.n1275 0.0217373
R19729 GNDA.n1347 GNDA.n1346 0.0217373
R19730 GNDA.n1353 GNDA.n1352 0.0217373
R19731 GNDA.n1357 GNDA.n1266 0.0217373
R19732 GNDA.n1358 GNDA.n1357 0.0217373
R19733 GNDA.n1361 GNDA.n1360 0.0217373
R19734 GNDA.n1363 GNDA.n1262 0.0217373
R19735 GNDA.n1345 GNDA.n1269 0.0217373
R19736 GNDA.n1348 GNDA.n1347 0.0217373
R19737 GNDA.n1351 GNDA.n1267 0.0217373
R19738 GNDA.n1354 GNDA.n1353 0.0217373
R19739 GNDA.n1355 GNDA.n1266 0.0217373
R19740 GNDA.n1359 GNDA.n1358 0.0217373
R19741 GNDA.n1356 GNDA.n1264 0.0217373
R19742 GNDA.n1361 GNDA.n1260 0.0217373
R19743 GNDA.n1262 GNDA.n1260 0.0217373
R19744 GNDA.n1377 GNDA.n1258 0.0217373
R19745 GNDA.n1381 GNDA.n1380 0.0217373
R19746 GNDA.n1384 GNDA.n1383 0.0217373
R19747 GNDA.n1387 GNDA.n1254 0.0217373
R19748 GNDA.n1390 GNDA.n1253 0.0217373
R19749 GNDA.n1389 GNDA.n1253 0.0217373
R19750 GNDA.n1379 GNDA.n1258 0.0217373
R19751 GNDA.n1382 GNDA.n1381 0.0217373
R19752 GNDA.n1294 GNDA.n1293 0.0217373
R19753 GNDA.n1383 GNDA.n1256 0.0217373
R19754 GNDA.n1256 GNDA.n1254 0.0217373
R19755 GNDA.n1299 GNDA.n1292 0.0217373
R19756 GNDA.n1297 GNDA.n1295 0.0217373
R19757 GNDA.n1294 GNDA.n436 0.0217373
R19758 GNDA.n3625 GNDA.n544 0.0217373
R19759 GNDA.n3625 GNDA.n542 0.0217373
R19760 GNDA.n589 GNDA.n587 0.0217373
R19761 GNDA.n589 GNDA.n585 0.0217373
R19762 GNDA.n4584 GNDA.n472 0.0217373
R19763 GNDA.n4585 GNDA.n472 0.0217373
R19764 GNDA.n470 GNDA.n467 0.0217373
R19765 GNDA.n471 GNDA.n467 0.0217373
R19766 GNDA.n465 GNDA.n462 0.0217373
R19767 GNDA.n466 GNDA.n462 0.0217373
R19768 GNDA.n460 GNDA.n457 0.0217373
R19769 GNDA.n461 GNDA.n457 0.0217373
R19770 GNDA.n455 GNDA.n452 0.0217373
R19771 GNDA.n456 GNDA.n452 0.0217373
R19772 GNDA.n446 GNDA.n443 0.0217373
R19773 GNDA.n447 GNDA.n443 0.0217373
R19774 GNDA.n441 GNDA.n438 0.0217373
R19775 GNDA.n442 GNDA.n438 0.0217373
R19776 GNDA.n509 GNDA.n507 0.0217373
R19777 GNDA.n509 GNDA.n506 0.0217373
R19778 GNDA.n3714 GNDA.n540 0.0217373
R19779 GNDA.n3715 GNDA.n3714 0.0217373
R19780 GNDA.n549 GNDA.n547 0.0217373
R19781 GNDA.n549 GNDA.n546 0.0217373
R19782 GNDA.n3480 GNDA.n580 0.0217373
R19783 GNDA.n3481 GNDA.n3480 0.0217373
R19784 GNDA.n3391 GNDA.n583 0.0217373
R19785 GNDA.n3391 GNDA.n582 0.0217373
R19786 GNDA.n3246 GNDA.n620 0.0217373
R19787 GNDA.n3247 GNDA.n3246 0.0217373
R19788 GNDA.n3157 GNDA.n623 0.0217373
R19789 GNDA.n3157 GNDA.n622 0.0217373
R19790 GNDA.n1399 GNDA.n1396 0.0217373
R19791 GNDA.n1400 GNDA.n1396 0.0217373
R19792 GNDA.n1394 GNDA.n1391 0.0217373
R19793 GNDA.n1395 GNDA.n1391 0.0217373
R19794 GNDA.n1251 GNDA.n1167 0.0217373
R19795 GNDA.n1252 GNDA.n1167 0.0217373
R19796 GNDA.n1864 GNDA.n1769 0.0217373
R19797 GNDA.n1865 GNDA.n1864 0.0217373
R19798 GNDA.n1860 GNDA.n1772 0.0217373
R19799 GNDA.n1855 GNDA.n1843 0.0217373
R19800 GNDA.n1850 GNDA.n1846 0.0217373
R19801 GNDA.n1768 GNDA.n1166 0.0217373
R19802 GNDA.n1765 GNDA.n1764 0.0217373
R19803 GNDA.n1761 GNDA.n1760 0.0217373
R19804 GNDA.n1757 GNDA.n1756 0.0217373
R19805 GNDA.n1753 GNDA.n1752 0.0217373
R19806 GNDA.n1741 GNDA.n1740 0.0217373
R19807 GNDA.n3240 GNDA.n621 0.0217373
R19808 GNDA.n619 GNDA.n618 0.0217373
R19809 GNDA.n3387 GNDA.n584 0.0217373
R19810 GNDA.n3474 GNDA.n581 0.0217373
R19811 GNDA.n579 GNDA.n578 0.0217373
R19812 GNDA.n3621 GNDA.n545 0.0217373
R19813 GNDA.n3708 GNDA.n541 0.0217373
R19814 GNDA.n539 GNDA.n538 0.0217373
R19815 GNDA.n3855 GNDA.n505 0.0217373
R19816 GNDA.n503 GNDA.n502 0.0217373
R19817 GNDA.n4616 GNDA.n4615 0.0217373
R19818 GNDA.n4612 GNDA.n4611 0.0217373
R19819 GNDA.n4608 GNDA.n4607 0.0217373
R19820 GNDA.n4604 GNDA.n4603 0.0217373
R19821 GNDA.n4600 GNDA.n4599 0.0217373
R19822 GNDA.n4596 GNDA.n4595 0.0217373
R19823 GNDA.n4592 GNDA.n4591 0.0217373
R19824 GNDA.n4588 GNDA.n4587 0.0217373
R19825 GNDA.n1847 GNDA.n1845 0.0217373
R19826 GNDA.n1847 GNDA.n1846 0.0217373
R19827 GNDA.n1852 GNDA.n1842 0.0217373
R19828 GNDA.n1852 GNDA.n1843 0.0217373
R19829 GNDA.n1857 GNDA.n1771 0.0217373
R19830 GNDA.n1857 GNDA.n1772 0.0217373
R19831 GNDA.n1862 GNDA.n1769 0.0217373
R19832 GNDA.n1866 GNDA.n1865 0.0217373
R19833 GNDA.n1863 GNDA.n1166 0.0217373
R19834 GNDA.n1251 GNDA.n1168 0.0217373
R19835 GNDA.n1252 GNDA.n1250 0.0217373
R19836 GNDA.n1766 GNDA.n1765 0.0217373
R19837 GNDA.n1394 GNDA.n1392 0.0217373
R19838 GNDA.n1395 GNDA.n1393 0.0217373
R19839 GNDA.n1758 GNDA.n1757 0.0217373
R19840 GNDA.n1399 GNDA.n1397 0.0217373
R19841 GNDA.n1400 GNDA.n1398 0.0217373
R19842 GNDA.n1754 GNDA.n1753 0.0217373
R19843 GNDA.n1742 GNDA.n1741 0.0217373
R19844 GNDA.n3242 GNDA.n623 0.0217373
R19845 GNDA.n3239 GNDA.n622 0.0217373
R19846 GNDA.n3241 GNDA.n3240 0.0217373
R19847 GNDA.n3244 GNDA.n620 0.0217373
R19848 GNDA.n3248 GNDA.n3247 0.0217373
R19849 GNDA.n3245 GNDA.n618 0.0217373
R19850 GNDA.n3476 GNDA.n583 0.0217373
R19851 GNDA.n3473 GNDA.n582 0.0217373
R19852 GNDA.n3475 GNDA.n3474 0.0217373
R19853 GNDA.n3478 GNDA.n580 0.0217373
R19854 GNDA.n3482 GNDA.n3481 0.0217373
R19855 GNDA.n3479 GNDA.n578 0.0217373
R19856 GNDA.n3623 GNDA.n547 0.0217373
R19857 GNDA.n3620 GNDA.n546 0.0217373
R19858 GNDA.n3622 GNDA.n3621 0.0217373
R19859 GNDA.n3712 GNDA.n540 0.0217373
R19860 GNDA.n3716 GNDA.n3715 0.0217373
R19861 GNDA.n3713 GNDA.n538 0.0217373
R19862 GNDA.n3857 GNDA.n507 0.0217373
R19863 GNDA.n3854 GNDA.n506 0.0217373
R19864 GNDA.n3856 GNDA.n3855 0.0217373
R19865 GNDA.n441 GNDA.n439 0.0217373
R19866 GNDA.n442 GNDA.n440 0.0217373
R19867 GNDA.n4617 GNDA.n4616 0.0217373
R19868 GNDA.n446 GNDA.n444 0.0217373
R19869 GNDA.n447 GNDA.n445 0.0217373
R19870 GNDA.n4613 GNDA.n4612 0.0217373
R19871 GNDA.n3950 GNDA.n502 0.0217373
R19872 GNDA.n455 GNDA.n453 0.0217373
R19873 GNDA.n456 GNDA.n454 0.0217373
R19874 GNDA.n4605 GNDA.n4604 0.0217373
R19875 GNDA.n460 GNDA.n458 0.0217373
R19876 GNDA.n461 GNDA.n459 0.0217373
R19877 GNDA.n4601 GNDA.n4600 0.0217373
R19878 GNDA.n465 GNDA.n463 0.0217373
R19879 GNDA.n466 GNDA.n464 0.0217373
R19880 GNDA.n4597 GNDA.n4596 0.0217373
R19881 GNDA.n470 GNDA.n468 0.0217373
R19882 GNDA.n471 GNDA.n469 0.0217373
R19883 GNDA.n4593 GNDA.n4592 0.0217373
R19884 GNDA.n4584 GNDA.n473 0.0217373
R19885 GNDA.n4585 GNDA.n4583 0.0217373
R19886 GNDA.n4589 GNDA.n4588 0.0217373
R19887 GNDA.n1390 GNDA.n1388 0.0217373
R19888 GNDA.n1762 GNDA.n1761 0.0217373
R19889 GNDA.n451 GNDA.n449 0.0217373
R19890 GNDA.n4609 GNDA.n4608 0.0217373
R19891 GNDA.n3389 GNDA.n587 0.0217373
R19892 GNDA.n3386 GNDA.n585 0.0217373
R19893 GNDA.n3388 GNDA.n3387 0.0217373
R19894 GNDA.n3710 GNDA.n544 0.0217373
R19895 GNDA.n3707 GNDA.n542 0.0217373
R19896 GNDA.n3709 GNDA.n3708 0.0217373
R19897 GNDA.n2392 GNDA.n2299 0.0217373
R19898 GNDA.n2395 GNDA.n2283 0.0217373
R19899 GNDA.n2298 GNDA.n2285 0.0217373
R19900 GNDA.n2299 GNDA.n2286 0.0217373
R19901 GNDA.n2280 GNDA.n2279 0.0217373
R19902 GNDA.n2283 GNDA.n2279 0.0217373
R19903 GNDA.n2217 GNDA.n2216 0.0217373
R19904 GNDA.n2213 GNDA.n699 0.0217373
R19905 GNDA.n3026 GNDA.n701 0.0217373
R19906 GNDA.n3027 GNDA.n702 0.0217373
R19907 GNDA.n2216 GNDA.n2212 0.0217373
R19908 GNDA.n2213 GNDA.n2212 0.0217373
R19909 GNDA.n2239 GNDA.n839 0.0217373
R19910 GNDA.n2228 GNDA.n841 0.0217373
R19911 GNDA.n2232 GNDA.n2231 0.0217373
R19912 GNDA.n2235 GNDA.n840 0.0217373
R19913 GNDA.n2230 GNDA.n841 0.0217373
R19914 GNDA.n2233 GNDA.n2232 0.0217373
R19915 GNDA.n2234 GNDA.n839 0.0217373
R19916 GNDA.n1351 GNDA.n1268 0.0217373
R19917 GNDA.n1286 GNDA.n1284 0.0217373
R19918 GNDA.n1304 GNDA.n1290 0.0217373
R19919 GNDA.n1300 GNDA.n1290 0.0217373
R19920 GNDA.n1283 GNDA.n1281 0.0217373
R19921 GNDA.n1280 GNDA.n1278 0.0217373
R19922 GNDA.n1332 GNDA.n1279 0.0217373
R19923 GNDA.n1327 GNDA.n1282 0.0217373
R19924 GNDA.n1318 GNDA.n1285 0.0217373
R19925 GNDA.n1333 GNDA.n1332 0.0217373
R19926 GNDA.n1328 GNDA.n1327 0.0217373
R19927 GNDA.n1323 GNDA.n1281 0.0217373
R19928 GNDA.n1319 GNDA.n1318 0.0217373
R19929 GNDA.n1345 GNDA.n1270 0.0217373
R19930 GNDA.n1338 GNDA.n1276 0.0217373
R19931 GNDA.n1334 GNDA.n1276 0.0217373
R19932 GNDA.n1346 GNDA.n1344 0.0217373
R19933 GNDA.n1352 GNDA.n1350 0.0217373
R19934 GNDA.n1350 GNDA.n1349 0.0217373
R19935 GNDA.n1364 GNDA.n1261 0.0217373
R19936 GNDA.n1263 GNDA.n1261 0.0217373
R19937 GNDA.n1379 GNDA.n1259 0.0217373
R19938 GNDA.n1380 GNDA.n1378 0.0217373
R19939 GNDA.n1386 GNDA.n1385 0.0217373
R19940 GNDA.n1385 GNDA.n1257 0.0217373
R19941 GNDA.n1849 GNDA.n1848 0.0217373
R19942 GNDA.n1854 GNDA.n1853 0.0217373
R19943 GNDA.n1859 GNDA.n1858 0.0217373
R19944 GNDA.n1848 GNDA.n1844 0.0217373
R19945 GNDA.n1853 GNDA.n1841 0.0217373
R19946 GNDA.n1858 GNDA.n1770 0.0217373
R19947 GNDA.n2286 GNDA.n2284 0.0217373
R19948 GNDA.n2393 GNDA.n2285 0.0217373
R19949 GNDA.n2394 GNDA.n2393 0.0217373
R19950 GNDA.n2297 GNDA.n2284 0.0217373
R19951 GNDA.n2396 GNDA.n2281 0.0217373
R19952 GNDA.n702 GNDA.n700 0.0217373
R19953 GNDA.n2282 GNDA.n2281 0.0217373
R19954 GNDA.n3028 GNDA.n701 0.0217373
R19955 GNDA.n3029 GNDA.n3028 0.0217373
R19956 GNDA.n3025 GNDA.n700 0.0217373
R19957 GNDA.n2211 GNDA.n2206 0.0217373
R19958 GNDA.n2214 GNDA.n2206 0.0217373
R19959 GNDA.n2236 GNDA.n2234 0.0217373
R19960 GNDA.n2230 GNDA.n842 0.0217373
R19961 GNDA.n2231 GNDA.n2229 0.0217373
R19962 GNDA.n2238 GNDA.n840 0.0217373
R19963 GNDA.n2229 GNDA.n2226 0.0217373
R19964 GNDA.n2238 GNDA.n2237 0.0217373
R19965 GNDA.n3951 GNDA.n504 0.0181756
R19966 GNDA.n3952 GNDA.n3951 0.0181756
R19967 GNDA.n1405 GNDA.n1401 0.0181756
R19968 GNDA.n1406 GNDA.n1401 0.0181756
R19969 GNDA.n1405 GNDA.n1403 0.0181756
R19970 GNDA.n1406 GNDA.n1404 0.0181756
R19971 GNDA.n3949 GNDA.n504 0.0181756
R19972 GNDA.n3953 GNDA.n3952 0.0181756
R19973 GNDA.n1925 GNDA.n1924 0.0107812
R19974 GNDA.n1924 GNDA.n1153 0.0107812
R19975 GNDA.n1492 GNDA.n1153 0.0107812
R19976 GNDA.n1574 GNDA.n1492 0.0107812
R19977 GNDA.n1656 GNDA.n1574 0.0107812
R19978 GNDA.n1732 GNDA.n1656 0.0107812
R19979 GNDA.n1732 GNDA.n593 0.0107812
R19980 GNDA.n3306 GNDA.n593 0.0107812
R19981 GNDA.n3382 GNDA.n3306 0.0107812
R19982 GNDA.n3382 GNDA.n553 0.0107812
R19983 GNDA.n3540 GNDA.n553 0.0107812
R19984 GNDA.n3616 GNDA.n3540 0.0107812
R19985 GNDA.n3616 GNDA.n513 0.0107812
R19986 GNDA.n3774 GNDA.n513 0.0107812
R19987 GNDA.n3850 GNDA.n3774 0.0107812
R19988 GNDA.n3850 GNDA.n477 0.0107812
R19989 GNDA.n4011 GNDA.n477 0.0107812
R19990 GNDA.n4093 GNDA.n4011 0.0107812
R19991 GNDA.n4175 GNDA.n4093 0.0107812
R19992 GNDA.n4257 GNDA.n4175 0.0107812
R19993 GNDA.n4339 GNDA.n4257 0.0107812
R19994 GNDA.n4421 GNDA.n4339 0.0107812
R19995 GNDA.n4503 GNDA.n4421 0.0107812
R19996 GNDA.n4579 GNDA.n4503 0.0107812
R19997 GNDA.n1959 GNDA.n1063 0.00182188
R19998 GNDA.n1112 GNDA.n1045 0.00182188
R19999 GNDA.n2049 GNDA.n897 0.00182188
R20000 GNDA.n2007 GNDA.n1991 0.00182188
R20001 GNDA.n1957 GNDA.n1045 0.00166081
R20002 GNDA.n1112 GNDA.n1029 0.00166081
R20003 GNDA.n1955 GNDA.n1114 0.00166081
R20004 GNDA.n1114 GNDA.n1030 0.00166081
R20005 GNDA.n1953 GNDA.n1115 0.00166081
R20006 GNDA.n1115 GNDA.n1031 0.00166081
R20007 GNDA.n1951 GNDA.n1116 0.00166081
R20008 GNDA.n1116 GNDA.n1032 0.00166081
R20009 GNDA.n1949 GNDA.n1117 0.00166081
R20010 GNDA.n1117 GNDA.n1033 0.00166081
R20011 GNDA.n1947 GNDA.n1118 0.00166081
R20012 GNDA.n1118 GNDA.n1034 0.00166081
R20013 GNDA.n1945 GNDA.n1119 0.00166081
R20014 GNDA.n1119 GNDA.n1035 0.00166081
R20015 GNDA.n1943 GNDA.n1120 0.00166081
R20016 GNDA.n1120 GNDA.n1036 0.00166081
R20017 GNDA.n1941 GNDA.n1121 0.00166081
R20018 GNDA.n1121 GNDA.n1037 0.00166081
R20019 GNDA.n1939 GNDA.n1122 0.00166081
R20020 GNDA.n1122 GNDA.n1038 0.00166081
R20021 GNDA.n1937 GNDA.n1123 0.00166081
R20022 GNDA.n1123 GNDA.n1039 0.00166081
R20023 GNDA.n1935 GNDA.n1124 0.00166081
R20024 GNDA.n1124 GNDA.n1040 0.00166081
R20025 GNDA.n1933 GNDA.n1125 0.00166081
R20026 GNDA.n1125 GNDA.n1041 0.00166081
R20027 GNDA.n1931 GNDA.n1126 0.00166081
R20028 GNDA.n1126 GNDA.n1042 0.00166081
R20029 GNDA.n1929 GNDA.n1127 0.00166081
R20030 GNDA.n1127 GNDA.n1043 0.00166081
R20031 GNDA.n1927 GNDA.n1128 0.00166081
R20032 GNDA.n1128 GNDA.n1044 0.00166081
R20033 GNDA.n897 GNDA.n864 0.00166081
R20034 GNDA.n2046 GNDA.n931 0.00166081
R20035 GNDA.n931 GNDA.n865 0.00166081
R20036 GNDA.n2044 GNDA.n932 0.00166081
R20037 GNDA.n932 GNDA.n866 0.00166081
R20038 GNDA.n2042 GNDA.n933 0.00166081
R20039 GNDA.n933 GNDA.n867 0.00166081
R20040 GNDA.n2040 GNDA.n934 0.00166081
R20041 GNDA.n934 GNDA.n868 0.00166081
R20042 GNDA.n2038 GNDA.n935 0.00166081
R20043 GNDA.n935 GNDA.n869 0.00166081
R20044 GNDA.n2036 GNDA.n936 0.00166081
R20045 GNDA.n936 GNDA.n870 0.00166081
R20046 GNDA.n2034 GNDA.n937 0.00166081
R20047 GNDA.n937 GNDA.n871 0.00166081
R20048 GNDA.n2032 GNDA.n938 0.00166081
R20049 GNDA.n938 GNDA.n872 0.00166081
R20050 GNDA.n2030 GNDA.n939 0.00166081
R20051 GNDA.n939 GNDA.n873 0.00166081
R20052 GNDA.n2028 GNDA.n940 0.00166081
R20053 GNDA.n940 GNDA.n874 0.00166081
R20054 GNDA.n2026 GNDA.n941 0.00166081
R20055 GNDA.n941 GNDA.n875 0.00166081
R20056 GNDA.n2024 GNDA.n942 0.00166081
R20057 GNDA.n942 GNDA.n876 0.00166081
R20058 GNDA.n2022 GNDA.n943 0.00166081
R20059 GNDA.n943 GNDA.n877 0.00166081
R20060 GNDA.n2020 GNDA.n944 0.00166081
R20061 GNDA.n944 GNDA.n878 0.00166081
R20062 GNDA.n2018 GNDA.n945 0.00166081
R20063 GNDA.n945 GNDA.n879 0.00166081
R20064 GNDA.n2016 GNDA.n880 0.00166081
R20065 GNDA.n2052 GNDA.n846 0.00166081
R20066 GNDA.n2051 GNDA.n863 0.00166081
R20067 GNDA.n899 GNDA.n898 0.00166081
R20068 GNDA.n896 GNDA.n862 0.00166081
R20069 GNDA.n901 GNDA.n900 0.00166081
R20070 GNDA.n895 GNDA.n861 0.00166081
R20071 GNDA.n903 GNDA.n902 0.00166081
R20072 GNDA.n894 GNDA.n860 0.00166081
R20073 GNDA.n905 GNDA.n904 0.00166081
R20074 GNDA.n893 GNDA.n859 0.00166081
R20075 GNDA.n907 GNDA.n906 0.00166081
R20076 GNDA.n892 GNDA.n858 0.00166081
R20077 GNDA.n909 GNDA.n908 0.00166081
R20078 GNDA.n891 GNDA.n857 0.00166081
R20079 GNDA.n911 GNDA.n910 0.00166081
R20080 GNDA.n890 GNDA.n856 0.00166081
R20081 GNDA.n913 GNDA.n912 0.00166081
R20082 GNDA.n889 GNDA.n855 0.00166081
R20083 GNDA.n915 GNDA.n914 0.00166081
R20084 GNDA.n888 GNDA.n854 0.00166081
R20085 GNDA.n917 GNDA.n916 0.00166081
R20086 GNDA.n887 GNDA.n853 0.00166081
R20087 GNDA.n919 GNDA.n918 0.00166081
R20088 GNDA.n886 GNDA.n852 0.00166081
R20089 GNDA.n921 GNDA.n920 0.00166081
R20090 GNDA.n885 GNDA.n851 0.00166081
R20091 GNDA.n923 GNDA.n922 0.00166081
R20092 GNDA.n884 GNDA.n850 0.00166081
R20093 GNDA.n925 GNDA.n924 0.00166081
R20094 GNDA.n883 GNDA.n849 0.00166081
R20095 GNDA.n927 GNDA.n926 0.00166081
R20096 GNDA.n882 GNDA.n848 0.00166081
R20097 GNDA.n929 GNDA.n928 0.00166081
R20098 GNDA.n881 GNDA.n847 0.00166081
R20099 GNDA.n2048 GNDA.n930 0.00166081
R20100 GNDA.n2015 GNDA.n2014 0.00166081
R20101 GNDA.n2010 GNDA.n2008 0.00166081
R20102 GNDA.n2009 GNDA.n979 0.00166081
R20103 GNDA.n1992 GNDA.n981 0.00166081
R20104 GNDA.n1011 GNDA.n978 0.00166081
R20105 GNDA.n1993 GNDA.n982 0.00166081
R20106 GNDA.n1010 GNDA.n977 0.00166081
R20107 GNDA.n1994 GNDA.n983 0.00166081
R20108 GNDA.n1009 GNDA.n976 0.00166081
R20109 GNDA.n1995 GNDA.n984 0.00166081
R20110 GNDA.n1008 GNDA.n975 0.00166081
R20111 GNDA.n1996 GNDA.n985 0.00166081
R20112 GNDA.n1007 GNDA.n974 0.00166081
R20113 GNDA.n1997 GNDA.n986 0.00166081
R20114 GNDA.n1006 GNDA.n973 0.00166081
R20115 GNDA.n1998 GNDA.n987 0.00166081
R20116 GNDA.n1005 GNDA.n972 0.00166081
R20117 GNDA.n1999 GNDA.n988 0.00166081
R20118 GNDA.n1004 GNDA.n971 0.00166081
R20119 GNDA.n2000 GNDA.n989 0.00166081
R20120 GNDA.n1003 GNDA.n970 0.00166081
R20121 GNDA.n2001 GNDA.n990 0.00166081
R20122 GNDA.n1002 GNDA.n969 0.00166081
R20123 GNDA.n2002 GNDA.n991 0.00166081
R20124 GNDA.n1001 GNDA.n968 0.00166081
R20125 GNDA.n2003 GNDA.n992 0.00166081
R20126 GNDA.n1000 GNDA.n967 0.00166081
R20127 GNDA.n2004 GNDA.n993 0.00166081
R20128 GNDA.n999 GNDA.n966 0.00166081
R20129 GNDA.n2005 GNDA.n994 0.00166081
R20130 GNDA.n998 GNDA.n965 0.00166081
R20131 GNDA.n2006 GNDA.n995 0.00166081
R20132 GNDA.n997 GNDA.n964 0.00166081
R20133 GNDA.n2012 GNDA.n996 0.00166081
R20134 GNDA.n1062 GNDA.n1028 0.00166081
R20135 GNDA.n1096 GNDA.n1065 0.00166081
R20136 GNDA.n1064 GNDA.n1061 0.00166081
R20137 GNDA.n1097 GNDA.n1067 0.00166081
R20138 GNDA.n1066 GNDA.n1060 0.00166081
R20139 GNDA.n1098 GNDA.n1069 0.00166081
R20140 GNDA.n1068 GNDA.n1059 0.00166081
R20141 GNDA.n1099 GNDA.n1071 0.00166081
R20142 GNDA.n1070 GNDA.n1058 0.00166081
R20143 GNDA.n1100 GNDA.n1073 0.00166081
R20144 GNDA.n1072 GNDA.n1057 0.00166081
R20145 GNDA.n1101 GNDA.n1075 0.00166081
R20146 GNDA.n1074 GNDA.n1056 0.00166081
R20147 GNDA.n1102 GNDA.n1077 0.00166081
R20148 GNDA.n1076 GNDA.n1055 0.00166081
R20149 GNDA.n1103 GNDA.n1079 0.00166081
R20150 GNDA.n1078 GNDA.n1054 0.00166081
R20151 GNDA.n1104 GNDA.n1081 0.00166081
R20152 GNDA.n1080 GNDA.n1053 0.00166081
R20153 GNDA.n1105 GNDA.n1083 0.00166081
R20154 GNDA.n1082 GNDA.n1052 0.00166081
R20155 GNDA.n1106 GNDA.n1085 0.00166081
R20156 GNDA.n1084 GNDA.n1051 0.00166081
R20157 GNDA.n1107 GNDA.n1087 0.00166081
R20158 GNDA.n1086 GNDA.n1050 0.00166081
R20159 GNDA.n1108 GNDA.n1089 0.00166081
R20160 GNDA.n1088 GNDA.n1049 0.00166081
R20161 GNDA.n1109 GNDA.n1091 0.00166081
R20162 GNDA.n1090 GNDA.n1048 0.00166081
R20163 GNDA.n1110 GNDA.n1093 0.00166081
R20164 GNDA.n1092 GNDA.n1047 0.00166081
R20165 GNDA.n1111 GNDA.n1095 0.00166081
R20166 GNDA.n1094 GNDA.n1046 0.00166081
R20167 GNDA.n1958 GNDA.n1113 0.00166081
R20168 GNDA.n2051 GNDA.n2050 0.00166081
R20169 GNDA.n2017 GNDA.n879 0.00166081
R20170 GNDA.n2019 GNDA.n878 0.00166081
R20171 GNDA.n2021 GNDA.n877 0.00166081
R20172 GNDA.n2023 GNDA.n876 0.00166081
R20173 GNDA.n2025 GNDA.n875 0.00166081
R20174 GNDA.n2027 GNDA.n874 0.00166081
R20175 GNDA.n2029 GNDA.n873 0.00166081
R20176 GNDA.n2031 GNDA.n872 0.00166081
R20177 GNDA.n2033 GNDA.n871 0.00166081
R20178 GNDA.n2035 GNDA.n870 0.00166081
R20179 GNDA.n2037 GNDA.n869 0.00166081
R20180 GNDA.n2039 GNDA.n868 0.00166081
R20181 GNDA.n2041 GNDA.n867 0.00166081
R20182 GNDA.n2043 GNDA.n866 0.00166081
R20183 GNDA.n2045 GNDA.n865 0.00166081
R20184 GNDA.n2047 GNDA.n864 0.00166081
R20185 GNDA.n2017 GNDA.n2016 0.00166081
R20186 GNDA.n2019 GNDA.n2018 0.00166081
R20187 GNDA.n2021 GNDA.n2020 0.00166081
R20188 GNDA.n2023 GNDA.n2022 0.00166081
R20189 GNDA.n2025 GNDA.n2024 0.00166081
R20190 GNDA.n2027 GNDA.n2026 0.00166081
R20191 GNDA.n2029 GNDA.n2028 0.00166081
R20192 GNDA.n2031 GNDA.n2030 0.00166081
R20193 GNDA.n2033 GNDA.n2032 0.00166081
R20194 GNDA.n2035 GNDA.n2034 0.00166081
R20195 GNDA.n2037 GNDA.n2036 0.00166081
R20196 GNDA.n2039 GNDA.n2038 0.00166081
R20197 GNDA.n2041 GNDA.n2040 0.00166081
R20198 GNDA.n2043 GNDA.n2042 0.00166081
R20199 GNDA.n2045 GNDA.n2044 0.00166081
R20200 GNDA.n2047 GNDA.n2046 0.00166081
R20201 GNDA.n898 GNDA.n863 0.00166081
R20202 GNDA.n899 GNDA.n862 0.00166081
R20203 GNDA.n900 GNDA.n896 0.00166081
R20204 GNDA.n901 GNDA.n861 0.00166081
R20205 GNDA.n902 GNDA.n895 0.00166081
R20206 GNDA.n903 GNDA.n860 0.00166081
R20207 GNDA.n904 GNDA.n894 0.00166081
R20208 GNDA.n905 GNDA.n859 0.00166081
R20209 GNDA.n906 GNDA.n893 0.00166081
R20210 GNDA.n907 GNDA.n858 0.00166081
R20211 GNDA.n908 GNDA.n892 0.00166081
R20212 GNDA.n909 GNDA.n857 0.00166081
R20213 GNDA.n910 GNDA.n891 0.00166081
R20214 GNDA.n911 GNDA.n856 0.00166081
R20215 GNDA.n912 GNDA.n890 0.00166081
R20216 GNDA.n913 GNDA.n855 0.00166081
R20217 GNDA.n914 GNDA.n889 0.00166081
R20218 GNDA.n915 GNDA.n854 0.00166081
R20219 GNDA.n916 GNDA.n888 0.00166081
R20220 GNDA.n917 GNDA.n853 0.00166081
R20221 GNDA.n918 GNDA.n887 0.00166081
R20222 GNDA.n919 GNDA.n852 0.00166081
R20223 GNDA.n920 GNDA.n886 0.00166081
R20224 GNDA.n921 GNDA.n851 0.00166081
R20225 GNDA.n922 GNDA.n885 0.00166081
R20226 GNDA.n923 GNDA.n850 0.00166081
R20227 GNDA.n924 GNDA.n884 0.00166081
R20228 GNDA.n925 GNDA.n849 0.00166081
R20229 GNDA.n926 GNDA.n883 0.00166081
R20230 GNDA.n927 GNDA.n848 0.00166081
R20231 GNDA.n928 GNDA.n882 0.00166081
R20232 GNDA.n929 GNDA.n847 0.00166081
R20233 GNDA.n930 GNDA.n881 0.00166081
R20234 GNDA.n880 GNDA.n846 0.00166081
R20235 GNDA.n1926 GNDA.n1044 0.00166081
R20236 GNDA.n1928 GNDA.n1043 0.00166081
R20237 GNDA.n1930 GNDA.n1042 0.00166081
R20238 GNDA.n1932 GNDA.n1041 0.00166081
R20239 GNDA.n1934 GNDA.n1040 0.00166081
R20240 GNDA.n1936 GNDA.n1039 0.00166081
R20241 GNDA.n1938 GNDA.n1038 0.00166081
R20242 GNDA.n1940 GNDA.n1037 0.00166081
R20243 GNDA.n1942 GNDA.n1036 0.00166081
R20244 GNDA.n1944 GNDA.n1035 0.00166081
R20245 GNDA.n1946 GNDA.n1034 0.00166081
R20246 GNDA.n1948 GNDA.n1033 0.00166081
R20247 GNDA.n1950 GNDA.n1032 0.00166081
R20248 GNDA.n1952 GNDA.n1031 0.00166081
R20249 GNDA.n1954 GNDA.n1030 0.00166081
R20250 GNDA.n1956 GNDA.n1029 0.00166081
R20251 GNDA.n1960 GNDA.n1028 0.00166081
R20252 GNDA.n1928 GNDA.n1927 0.00166081
R20253 GNDA.n1930 GNDA.n1929 0.00166081
R20254 GNDA.n1932 GNDA.n1931 0.00166081
R20255 GNDA.n1934 GNDA.n1933 0.00166081
R20256 GNDA.n1936 GNDA.n1935 0.00166081
R20257 GNDA.n1938 GNDA.n1937 0.00166081
R20258 GNDA.n1940 GNDA.n1939 0.00166081
R20259 GNDA.n1942 GNDA.n1941 0.00166081
R20260 GNDA.n1944 GNDA.n1943 0.00166081
R20261 GNDA.n1946 GNDA.n1945 0.00166081
R20262 GNDA.n1948 GNDA.n1947 0.00166081
R20263 GNDA.n1950 GNDA.n1949 0.00166081
R20264 GNDA.n1952 GNDA.n1951 0.00166081
R20265 GNDA.n1954 GNDA.n1953 0.00166081
R20266 GNDA.n1956 GNDA.n1955 0.00166081
R20267 GNDA.n1096 GNDA.n1062 0.00166081
R20268 GNDA.n1065 GNDA.n1064 0.00166081
R20269 GNDA.n1097 GNDA.n1061 0.00166081
R20270 GNDA.n1067 GNDA.n1066 0.00166081
R20271 GNDA.n1098 GNDA.n1060 0.00166081
R20272 GNDA.n1069 GNDA.n1068 0.00166081
R20273 GNDA.n1099 GNDA.n1059 0.00166081
R20274 GNDA.n1071 GNDA.n1070 0.00166081
R20275 GNDA.n1100 GNDA.n1058 0.00166081
R20276 GNDA.n1073 GNDA.n1072 0.00166081
R20277 GNDA.n1101 GNDA.n1057 0.00166081
R20278 GNDA.n1075 GNDA.n1074 0.00166081
R20279 GNDA.n1102 GNDA.n1056 0.00166081
R20280 GNDA.n1077 GNDA.n1076 0.00166081
R20281 GNDA.n1103 GNDA.n1055 0.00166081
R20282 GNDA.n1079 GNDA.n1078 0.00166081
R20283 GNDA.n1104 GNDA.n1054 0.00166081
R20284 GNDA.n1081 GNDA.n1080 0.00166081
R20285 GNDA.n1105 GNDA.n1053 0.00166081
R20286 GNDA.n1083 GNDA.n1082 0.00166081
R20287 GNDA.n1106 GNDA.n1052 0.00166081
R20288 GNDA.n1085 GNDA.n1084 0.00166081
R20289 GNDA.n1107 GNDA.n1051 0.00166081
R20290 GNDA.n1087 GNDA.n1086 0.00166081
R20291 GNDA.n1108 GNDA.n1050 0.00166081
R20292 GNDA.n1089 GNDA.n1088 0.00166081
R20293 GNDA.n1109 GNDA.n1049 0.00166081
R20294 GNDA.n1091 GNDA.n1090 0.00166081
R20295 GNDA.n1110 GNDA.n1048 0.00166081
R20296 GNDA.n1093 GNDA.n1092 0.00166081
R20297 GNDA.n1111 GNDA.n1047 0.00166081
R20298 GNDA.n1095 GNDA.n1094 0.00166081
R20299 GNDA.n1113 GNDA.n1046 0.00166081
R20300 GNDA.n1957 GNDA.n1063 0.00166081
R20301 GNDA.n2011 GNDA.n946 0.00166081
R20302 GNDA.n1991 GNDA.n947 0.00166081
R20303 GNDA.n1989 GNDA.n1012 0.00166081
R20304 GNDA.n1990 GNDA.n948 0.00166081
R20305 GNDA.n1987 GNDA.n1013 0.00166081
R20306 GNDA.n1988 GNDA.n949 0.00166081
R20307 GNDA.n1985 GNDA.n1014 0.00166081
R20308 GNDA.n1986 GNDA.n950 0.00166081
R20309 GNDA.n1983 GNDA.n1015 0.00166081
R20310 GNDA.n1984 GNDA.n951 0.00166081
R20311 GNDA.n1981 GNDA.n1016 0.00166081
R20312 GNDA.n1982 GNDA.n952 0.00166081
R20313 GNDA.n1979 GNDA.n1017 0.00166081
R20314 GNDA.n1980 GNDA.n953 0.00166081
R20315 GNDA.n1977 GNDA.n1018 0.00166081
R20316 GNDA.n1978 GNDA.n954 0.00166081
R20317 GNDA.n1975 GNDA.n1019 0.00166081
R20318 GNDA.n1976 GNDA.n955 0.00166081
R20319 GNDA.n1973 GNDA.n1020 0.00166081
R20320 GNDA.n1974 GNDA.n956 0.00166081
R20321 GNDA.n1971 GNDA.n1021 0.00166081
R20322 GNDA.n1972 GNDA.n957 0.00166081
R20323 GNDA.n1969 GNDA.n1022 0.00166081
R20324 GNDA.n1970 GNDA.n958 0.00166081
R20325 GNDA.n1967 GNDA.n1023 0.00166081
R20326 GNDA.n1968 GNDA.n959 0.00166081
R20327 GNDA.n1965 GNDA.n1024 0.00166081
R20328 GNDA.n1966 GNDA.n960 0.00166081
R20329 GNDA.n1963 GNDA.n1025 0.00166081
R20330 GNDA.n1964 GNDA.n961 0.00166081
R20331 GNDA.n1961 GNDA.n1026 0.00166081
R20332 GNDA.n1962 GNDA.n962 0.00166081
R20333 GNDA.n1027 GNDA.n980 0.00166081
R20334 GNDA.n1027 GNDA.n962 0.00166081
R20335 GNDA.n1026 GNDA.n961 0.00166081
R20336 GNDA.n1025 GNDA.n960 0.00166081
R20337 GNDA.n1024 GNDA.n959 0.00166081
R20338 GNDA.n1023 GNDA.n958 0.00166081
R20339 GNDA.n1022 GNDA.n957 0.00166081
R20340 GNDA.n1021 GNDA.n956 0.00166081
R20341 GNDA.n1020 GNDA.n955 0.00166081
R20342 GNDA.n1019 GNDA.n954 0.00166081
R20343 GNDA.n1018 GNDA.n953 0.00166081
R20344 GNDA.n1017 GNDA.n952 0.00166081
R20345 GNDA.n1016 GNDA.n951 0.00166081
R20346 GNDA.n1015 GNDA.n950 0.00166081
R20347 GNDA.n1014 GNDA.n949 0.00166081
R20348 GNDA.n1013 GNDA.n948 0.00166081
R20349 GNDA.n1012 GNDA.n947 0.00166081
R20350 GNDA.n2007 GNDA.n946 0.00166081
R20351 GNDA.n2014 GNDA.n963 0.00166081
R20352 GNDA.n1962 GNDA.n1961 0.00166081
R20353 GNDA.n1964 GNDA.n1963 0.00166081
R20354 GNDA.n1966 GNDA.n1965 0.00166081
R20355 GNDA.n1968 GNDA.n1967 0.00166081
R20356 GNDA.n1970 GNDA.n1969 0.00166081
R20357 GNDA.n1972 GNDA.n1971 0.00166081
R20358 GNDA.n1974 GNDA.n1973 0.00166081
R20359 GNDA.n1976 GNDA.n1975 0.00166081
R20360 GNDA.n1978 GNDA.n1977 0.00166081
R20361 GNDA.n1980 GNDA.n1979 0.00166081
R20362 GNDA.n1982 GNDA.n1981 0.00166081
R20363 GNDA.n1984 GNDA.n1983 0.00166081
R20364 GNDA.n1986 GNDA.n1985 0.00166081
R20365 GNDA.n1988 GNDA.n1987 0.00166081
R20366 GNDA.n1990 GNDA.n1989 0.00166081
R20367 GNDA.n2008 GNDA.n963 0.00166081
R20368 GNDA.n2013 GNDA.n980 0.00166081
R20369 GNDA.n2010 GNDA.n2009 0.00166081
R20370 GNDA.n1992 GNDA.n979 0.00166081
R20371 GNDA.n1011 GNDA.n981 0.00166081
R20372 GNDA.n1993 GNDA.n978 0.00166081
R20373 GNDA.n1010 GNDA.n982 0.00166081
R20374 GNDA.n1994 GNDA.n977 0.00166081
R20375 GNDA.n1009 GNDA.n983 0.00166081
R20376 GNDA.n1995 GNDA.n976 0.00166081
R20377 GNDA.n1008 GNDA.n984 0.00166081
R20378 GNDA.n1996 GNDA.n975 0.00166081
R20379 GNDA.n1007 GNDA.n985 0.00166081
R20380 GNDA.n1997 GNDA.n974 0.00166081
R20381 GNDA.n1006 GNDA.n986 0.00166081
R20382 GNDA.n1998 GNDA.n973 0.00166081
R20383 GNDA.n1005 GNDA.n987 0.00166081
R20384 GNDA.n1999 GNDA.n972 0.00166081
R20385 GNDA.n1004 GNDA.n988 0.00166081
R20386 GNDA.n2000 GNDA.n971 0.00166081
R20387 GNDA.n1003 GNDA.n989 0.00166081
R20388 GNDA.n2001 GNDA.n970 0.00166081
R20389 GNDA.n1002 GNDA.n990 0.00166081
R20390 GNDA.n2002 GNDA.n969 0.00166081
R20391 GNDA.n1001 GNDA.n991 0.00166081
R20392 GNDA.n2003 GNDA.n968 0.00166081
R20393 GNDA.n1000 GNDA.n992 0.00166081
R20394 GNDA.n2004 GNDA.n967 0.00166081
R20395 GNDA.n999 GNDA.n993 0.00166081
R20396 GNDA.n2005 GNDA.n966 0.00166081
R20397 GNDA.n998 GNDA.n994 0.00166081
R20398 GNDA.n2006 GNDA.n965 0.00166081
R20399 GNDA.n997 GNDA.n995 0.00166081
R20400 GNDA.n996 GNDA.n964 0.00166081
R20401 VOUT-.n176 VOUT-.t1 110.386
R20402 VOUT-.n39 VOUT-.n38 34.9935
R20403 VOUT-.n28 VOUT-.n27 34.9935
R20404 VOUT-.n30 VOUT-.n29 34.9935
R20405 VOUT-.n33 VOUT-.n32 34.9935
R20406 VOUT-.n36 VOUT-.n35 34.9935
R20407 VOUT-.n42 VOUT-.n41 34.9935
R20408 VOUT-.n183 VOUT-.n182 9.73997
R20409 VOUT-.n179 VOUT-.n178 9.73997
R20410 VOUT-.n186 VOUT-.n185 9.73997
R20411 VOUT-.n184 VOUT-.n179 6.64633
R20412 VOUT-.n184 VOUT-.n183 6.64633
R20413 VOUT-.n38 VOUT-.t10 6.56717
R20414 VOUT-.n38 VOUT-.t17 6.56717
R20415 VOUT-.n27 VOUT-.t16 6.56717
R20416 VOUT-.n27 VOUT-.t9 6.56717
R20417 VOUT-.n29 VOUT-.t13 6.56717
R20418 VOUT-.n29 VOUT-.t7 6.56717
R20419 VOUT-.n32 VOUT-.t14 6.56717
R20420 VOUT-.n32 VOUT-.t8 6.56717
R20421 VOUT-.n35 VOUT-.t12 6.56717
R20422 VOUT-.n35 VOUT-.t6 6.56717
R20423 VOUT-.n41 VOUT-.t11 6.56717
R20424 VOUT-.n41 VOUT-.t5 6.56717
R20425 VOUT-.n31 VOUT-.n28 6.3755
R20426 VOUT-.n40 VOUT-.n39 6.3755
R20427 VOUT-.n186 VOUT-.n184 6.02133
R20428 VOUT-.n31 VOUT-.n30 5.813
R20429 VOUT-.n34 VOUT-.n33 5.813
R20430 VOUT-.n37 VOUT-.n36 5.813
R20431 VOUT-.n42 VOUT-.n40 5.813
R20432 VOUT-.n46 VOUT-.n26 5.063
R20433 VOUT-.n43 VOUT-.n19 5.063
R20434 VOUT-.n109 VOUT-.t140 4.8295
R20435 VOUT-.n108 VOUT-.t55 4.8295
R20436 VOUT-.n107 VOUT-.t100 4.8295
R20437 VOUT-.n122 VOUT-.t131 4.8295
R20438 VOUT-.n123 VOUT-.t43 4.8295
R20439 VOUT-.n125 VOUT-.t103 4.8295
R20440 VOUT-.n126 VOUT-.t86 4.8295
R20441 VOUT-.n128 VOUT-.t68 4.8295
R20442 VOUT-.n129 VOUT-.t49 4.8295
R20443 VOUT-.n131 VOUT-.t98 4.8295
R20444 VOUT-.n132 VOUT-.t80 4.8295
R20445 VOUT-.n134 VOUT-.t62 4.8295
R20446 VOUT-.n135 VOUT-.t44 4.8295
R20447 VOUT-.n137 VOUT-.t19 4.8295
R20448 VOUT-.n138 VOUT-.t141 4.8295
R20449 VOUT-.n140 VOUT-.t56 4.8295
R20450 VOUT-.n141 VOUT-.t36 4.8295
R20451 VOUT-.n143 VOUT-.t150 4.8295
R20452 VOUT-.n144 VOUT-.t133 4.8295
R20453 VOUT-.n146 VOUT-.t110 4.8295
R20454 VOUT-.n147 VOUT-.t97 4.8295
R20455 VOUT-.n71 VOUT-.t96 4.8295
R20456 VOUT-.n73 VOUT-.t59 4.8295
R20457 VOUT-.n86 VOUT-.t116 4.8295
R20458 VOUT-.n87 VOUT-.t102 4.8295
R20459 VOUT-.n89 VOUT-.t152 4.8295
R20460 VOUT-.n90 VOUT-.t135 4.8295
R20461 VOUT-.n92 VOUT-.t63 4.8295
R20462 VOUT-.n93 VOUT-.t30 4.8295
R20463 VOUT-.n95 VOUT-.t67 4.8295
R20464 VOUT-.n96 VOUT-.t48 4.8295
R20465 VOUT-.n98 VOUT-.t29 4.8295
R20466 VOUT-.n99 VOUT-.t149 4.8295
R20467 VOUT-.n101 VOUT-.t71 4.8295
R20468 VOUT-.n102 VOUT-.t54 4.8295
R20469 VOUT-.n104 VOUT-.t107 4.8295
R20470 VOUT-.n105 VOUT-.t92 4.8295
R20471 VOUT-.n149 VOUT-.t74 4.8295
R20472 VOUT-.n110 VOUT-.t42 4.8154
R20473 VOUT-.n113 VOUT-.t75 4.8154
R20474 VOUT-.n111 VOUT-.t155 4.81305
R20475 VOUT-.n114 VOUT-.t53 4.81305
R20476 VOUT-.n112 VOUT-.t35 4.806
R20477 VOUT-.n115 VOUT-.t90 4.806
R20478 VOUT-.n116 VOUT-.t124 4.806
R20479 VOUT-.n74 VOUT-.t145 4.806
R20480 VOUT-.n75 VOUT-.t118 4.806
R20481 VOUT-.n76 VOUT-.t138 4.806
R20482 VOUT-.n77 VOUT-.t38 4.806
R20483 VOUT-.n78 VOUT-.t153 4.806
R20484 VOUT-.n79 VOUT-.t57 4.806
R20485 VOUT-.n80 VOUT-.t91 4.806
R20486 VOUT-.n81 VOUT-.t126 4.806
R20487 VOUT-.n82 VOUT-.t106 4.806
R20488 VOUT-.n83 VOUT-.t147 4.806
R20489 VOUT-.n84 VOUT-.t46 4.806
R20490 VOUT-.n109 VOUT-.t25 4.5005
R20491 VOUT-.n108 VOUT-.t144 4.5005
R20492 VOUT-.n107 VOUT-.t65 4.5005
R20493 VOUT-.n121 VOUT-.t23 4.5005
R20494 VOUT-.n120 VOUT-.t47 4.5005
R20495 VOUT-.n119 VOUT-.t148 4.5005
R20496 VOUT-.n118 VOUT-.t108 4.5005
R20497 VOUT-.n117 VOUT-.t127 4.5005
R20498 VOUT-.n116 VOUT-.t94 4.5005
R20499 VOUT-.n115 VOUT-.t58 4.5005
R20500 VOUT-.n114 VOUT-.t154 4.5005
R20501 VOUT-.n113 VOUT-.t41 4.5005
R20502 VOUT-.n112 VOUT-.t139 4.5005
R20503 VOUT-.n111 VOUT-.t121 4.5005
R20504 VOUT-.n110 VOUT-.t146 4.5005
R20505 VOUT-.n122 VOUT-.t95 4.5005
R20506 VOUT-.n124 VOUT-.t61 4.5005
R20507 VOUT-.n123 VOUT-.t78 4.5005
R20508 VOUT-.n125 VOUT-.t70 4.5005
R20509 VOUT-.n127 VOUT-.t32 4.5005
R20510 VOUT-.n126 VOUT-.t119 4.5005
R20511 VOUT-.n128 VOUT-.t27 4.5005
R20512 VOUT-.n130 VOUT-.t130 4.5005
R20513 VOUT-.n129 VOUT-.t82 4.5005
R20514 VOUT-.n131 VOUT-.t66 4.5005
R20515 VOUT-.n133 VOUT-.t26 4.5005
R20516 VOUT-.n132 VOUT-.t112 4.5005
R20517 VOUT-.n134 VOUT-.t24 4.5005
R20518 VOUT-.n136 VOUT-.t125 4.5005
R20519 VOUT-.n135 VOUT-.t76 4.5005
R20520 VOUT-.n137 VOUT-.t122 4.5005
R20521 VOUT-.n139 VOUT-.t88 4.5005
R20522 VOUT-.n138 VOUT-.t37 4.5005
R20523 VOUT-.n140 VOUT-.t156 4.5005
R20524 VOUT-.n142 VOUT-.t120 4.5005
R20525 VOUT-.n141 VOUT-.t72 4.5005
R20526 VOUT-.n143 VOUT-.t114 4.5005
R20527 VOUT-.n145 VOUT-.t83 4.5005
R20528 VOUT-.n144 VOUT-.t31 4.5005
R20529 VOUT-.n146 VOUT-.t77 4.5005
R20530 VOUT-.n148 VOUT-.t45 4.5005
R20531 VOUT-.n147 VOUT-.t128 4.5005
R20532 VOUT-.n71 VOUT-.t64 4.5005
R20533 VOUT-.n72 VOUT-.t22 4.5005
R20534 VOUT-.n73 VOUT-.t20 4.5005
R20535 VOUT-.n85 VOUT-.t117 4.5005
R20536 VOUT-.n84 VOUT-.t143 4.5005
R20537 VOUT-.n83 VOUT-.t105 4.5005
R20538 VOUT-.n82 VOUT-.t69 4.5005
R20539 VOUT-.n81 VOUT-.t89 4.5005
R20540 VOUT-.n80 VOUT-.t52 4.5005
R20541 VOUT-.n79 VOUT-.t151 4.5005
R20542 VOUT-.n78 VOUT-.t111 4.5005
R20543 VOUT-.n77 VOUT-.t134 4.5005
R20544 VOUT-.n76 VOUT-.t101 4.5005
R20545 VOUT-.n75 VOUT-.t79 4.5005
R20546 VOUT-.n74 VOUT-.t104 4.5005
R20547 VOUT-.n86 VOUT-.t85 4.5005
R20548 VOUT-.n88 VOUT-.t51 4.5005
R20549 VOUT-.n87 VOUT-.t136 4.5005
R20550 VOUT-.n89 VOUT-.t115 4.5005
R20551 VOUT-.n91 VOUT-.t84 4.5005
R20552 VOUT-.n90 VOUT-.t33 4.5005
R20553 VOUT-.n92 VOUT-.t109 4.5005
R20554 VOUT-.n94 VOUT-.t21 4.5005
R20555 VOUT-.n93 VOUT-.t113 4.5005
R20556 VOUT-.n95 VOUT-.t28 4.5005
R20557 VOUT-.n97 VOUT-.t129 4.5005
R20558 VOUT-.n96 VOUT-.t81 4.5005
R20559 VOUT-.n98 VOUT-.t132 4.5005
R20560 VOUT-.n100 VOUT-.t99 4.5005
R20561 VOUT-.n99 VOUT-.t50 4.5005
R20562 VOUT-.n101 VOUT-.t34 4.5005
R20563 VOUT-.n103 VOUT-.t137 4.5005
R20564 VOUT-.n102 VOUT-.t87 4.5005
R20565 VOUT-.n104 VOUT-.t73 4.5005
R20566 VOUT-.n106 VOUT-.t39 4.5005
R20567 VOUT-.n105 VOUT-.t123 4.5005
R20568 VOUT-.n149 VOUT-.t40 4.5005
R20569 VOUT-.n150 VOUT-.t142 4.5005
R20570 VOUT-.n151 VOUT-.t93 4.5005
R20571 VOUT-.n152 VOUT-.t60 4.5005
R20572 VOUT-.n47 VOUT-.n46 4.5005
R20573 VOUT-.n45 VOUT-.n24 4.5005
R20574 VOUT-.n44 VOUT-.n23 4.5005
R20575 VOUT-.n43 VOUT-.n20 4.5005
R20576 VOUT-.n65 VOUT-.n64 4.5005
R20577 VOUT-.n16 VOUT-.n13 4.5005
R20578 VOUT-.n65 VOUT-.n13 4.5005
R20579 VOUT-.n66 VOUT-.n9 4.5005
R20580 VOUT-.n66 VOUT-.n11 4.5005
R20581 VOUT-.n66 VOUT-.n65 4.5005
R20582 VOUT-.n161 VOUT-.n69 4.5005
R20583 VOUT-.n162 VOUT-.n161 4.5005
R20584 VOUT-.n162 VOUT-.n5 4.5005
R20585 VOUT-.n163 VOUT-.n4 4.5005
R20586 VOUT-.n163 VOUT-.n162 4.5005
R20587 VOUT-.n175 VOUT-.n174 4.5005
R20588 VOUT-.n175 VOUT-.n1 4.5005
R20589 VOUT-.n171 VOUT-.n1 4.5005
R20590 VOUT-.n168 VOUT-.n1 4.5005
R20591 VOUT-.n169 VOUT-.n1 4.5005
R20592 VOUT-.n171 VOUT-.n170 4.5005
R20593 VOUT-.n170 VOUT-.n168 4.5005
R20594 VOUT-.n170 VOUT-.n169 4.5005
R20595 VOUT-.n182 VOUT-.t0 3.42907
R20596 VOUT-.n182 VOUT-.t2 3.42907
R20597 VOUT-.n178 VOUT-.t3 3.42907
R20598 VOUT-.n178 VOUT-.t4 3.42907
R20599 VOUT-.n185 VOUT-.t15 3.42907
R20600 VOUT-.n185 VOUT-.t18 3.42907
R20601 VOUT-.n63 VOUT-.n62 2.24601
R20602 VOUT-.n14 VOUT-.n8 2.24601
R20603 VOUT-.n173 VOUT-.n172 2.24601
R20604 VOUT-.n167 VOUT-.n166 2.24601
R20605 VOUT-.n160 VOUT-.n159 2.24477
R20606 VOUT-.n7 VOUT-.n2 2.24477
R20607 VOUT-.n66 VOUT-.n10 2.24063
R20608 VOUT-.n163 VOUT-.n3 2.24063
R20609 VOUT-.n170 VOUT-.n0 2.24063
R20610 VOUT-.n13 VOUT-.n12 2.24063
R20611 VOUT-.n161 VOUT-.n67 2.24063
R20612 VOUT-.n68 VOUT-.n5 2.24063
R20613 VOUT-.n174 VOUT-.n165 2.24063
R20614 VOUT-.n174 VOUT-.n164 2.24063
R20615 VOUT-.n64 VOUT-.n17 2.23934
R20616 VOUT-.n64 VOUT-.n15 2.23934
R20617 VOUT-.n183 VOUT-.n181 1.83719
R20618 VOUT-.n194 VOUT-.n179 1.72967
R20619 VOUT-.n187 VOUT-.n186 1.72967
R20620 VOUT-.n50 VOUT-.n25 1.5005
R20621 VOUT-.n52 VOUT-.n51 1.5005
R20622 VOUT-.n53 VOUT-.n22 1.5005
R20623 VOUT-.n55 VOUT-.n54 1.5005
R20624 VOUT-.n56 VOUT-.n21 1.5005
R20625 VOUT-.n58 VOUT-.n57 1.5005
R20626 VOUT-.n59 VOUT-.n18 1.5005
R20627 VOUT-.n61 VOUT-.n60 1.5005
R20628 VOUT-.n189 VOUT-.n188 1.5005
R20629 VOUT-.n190 VOUT-.n180 1.5005
R20630 VOUT-.n192 VOUT-.n191 1.5005
R20631 VOUT-.n193 VOUT-.n177 1.5005
R20632 VOUT-.n195 VOUT-.n194 1.5005
R20633 VOUT-.n30 VOUT-.n20 1.313
R20634 VOUT-.n33 VOUT-.n23 1.313
R20635 VOUT-.n36 VOUT-.n24 1.313
R20636 VOUT-.n47 VOUT-.n42 1.313
R20637 VOUT-.n28 VOUT-.n19 1.313
R20638 VOUT-.n39 VOUT-.n26 1.313
R20639 VOUT-.n159 VOUT-.n158 1.1455
R20640 VOUT-.n153 VOUT-.n6 1.13717
R20641 VOUT-.n155 VOUT-.n154 1.13717
R20642 VOUT-.n157 VOUT-.n156 1.13717
R20643 VOUT-.n162 VOUT-.n6 1.13717
R20644 VOUT-.n155 VOUT-.n7 1.13717
R20645 VOUT-.n156 VOUT-.n4 1.13717
R20646 VOUT-.n70 VOUT-.n69 1.13717
R20647 VOUT-.n49 VOUT-.n26 0.715216
R20648 VOUT-.n58 VOUT-.n20 0.65675
R20649 VOUT-.n54 VOUT-.n23 0.65675
R20650 VOUT-.n52 VOUT-.n24 0.65675
R20651 VOUT-.n48 VOUT-.n47 0.65675
R20652 VOUT-.n60 VOUT-.n19 0.65675
R20653 VOUT-.n158 VOUT-.n157 0.585
R20654 VOUT-.n50 VOUT-.n49 0.564601
R20655 VOUT-.n46 VOUT-.n45 0.563
R20656 VOUT-.n45 VOUT-.n44 0.563
R20657 VOUT-.n44 VOUT-.n43 0.563
R20658 VOUT-.n34 VOUT-.n31 0.563
R20659 VOUT-.n37 VOUT-.n34 0.563
R20660 VOUT-.n40 VOUT-.n37 0.563
R20661 VOUT-.n174 VOUT-.n163 0.5455
R20662 VOUT-.n62 VOUT-.n61 0.495292
R20663 VOUT-.n121 VOUT-.n107 0.3295
R20664 VOUT-.n121 VOUT-.n120 0.3295
R20665 VOUT-.n120 VOUT-.n119 0.3295
R20666 VOUT-.n119 VOUT-.n118 0.3295
R20667 VOUT-.n118 VOUT-.n117 0.3295
R20668 VOUT-.n117 VOUT-.n116 0.3295
R20669 VOUT-.n116 VOUT-.n115 0.3295
R20670 VOUT-.n115 VOUT-.n114 0.3295
R20671 VOUT-.n114 VOUT-.n113 0.3295
R20672 VOUT-.n113 VOUT-.n112 0.3295
R20673 VOUT-.n112 VOUT-.n111 0.3295
R20674 VOUT-.n111 VOUT-.n110 0.3295
R20675 VOUT-.n124 VOUT-.n122 0.3295
R20676 VOUT-.n124 VOUT-.n123 0.3295
R20677 VOUT-.n127 VOUT-.n125 0.3295
R20678 VOUT-.n127 VOUT-.n126 0.3295
R20679 VOUT-.n130 VOUT-.n128 0.3295
R20680 VOUT-.n130 VOUT-.n129 0.3295
R20681 VOUT-.n133 VOUT-.n131 0.3295
R20682 VOUT-.n133 VOUT-.n132 0.3295
R20683 VOUT-.n136 VOUT-.n134 0.3295
R20684 VOUT-.n136 VOUT-.n135 0.3295
R20685 VOUT-.n139 VOUT-.n137 0.3295
R20686 VOUT-.n139 VOUT-.n138 0.3295
R20687 VOUT-.n142 VOUT-.n140 0.3295
R20688 VOUT-.n142 VOUT-.n141 0.3295
R20689 VOUT-.n145 VOUT-.n143 0.3295
R20690 VOUT-.n145 VOUT-.n144 0.3295
R20691 VOUT-.n148 VOUT-.n146 0.3295
R20692 VOUT-.n148 VOUT-.n147 0.3295
R20693 VOUT-.n72 VOUT-.n71 0.3295
R20694 VOUT-.n85 VOUT-.n73 0.3295
R20695 VOUT-.n85 VOUT-.n84 0.3295
R20696 VOUT-.n84 VOUT-.n83 0.3295
R20697 VOUT-.n83 VOUT-.n82 0.3295
R20698 VOUT-.n82 VOUT-.n81 0.3295
R20699 VOUT-.n81 VOUT-.n80 0.3295
R20700 VOUT-.n80 VOUT-.n79 0.3295
R20701 VOUT-.n79 VOUT-.n78 0.3295
R20702 VOUT-.n78 VOUT-.n77 0.3295
R20703 VOUT-.n77 VOUT-.n76 0.3295
R20704 VOUT-.n76 VOUT-.n75 0.3295
R20705 VOUT-.n75 VOUT-.n74 0.3295
R20706 VOUT-.n88 VOUT-.n86 0.3295
R20707 VOUT-.n88 VOUT-.n87 0.3295
R20708 VOUT-.n91 VOUT-.n89 0.3295
R20709 VOUT-.n91 VOUT-.n90 0.3295
R20710 VOUT-.n94 VOUT-.n92 0.3295
R20711 VOUT-.n94 VOUT-.n93 0.3295
R20712 VOUT-.n97 VOUT-.n95 0.3295
R20713 VOUT-.n97 VOUT-.n96 0.3295
R20714 VOUT-.n100 VOUT-.n98 0.3295
R20715 VOUT-.n100 VOUT-.n99 0.3295
R20716 VOUT-.n103 VOUT-.n101 0.3295
R20717 VOUT-.n103 VOUT-.n102 0.3295
R20718 VOUT-.n106 VOUT-.n104 0.3295
R20719 VOUT-.n106 VOUT-.n105 0.3295
R20720 VOUT-.n150 VOUT-.n149 0.3295
R20721 VOUT-.n151 VOUT-.n150 0.3295
R20722 VOUT-.n189 VOUT-.n181 0.314966
R20723 VOUT-.n152 VOUT-.n151 0.3107
R20724 VOUT-.n117 VOUT-.n109 0.306
R20725 VOUT-.n118 VOUT-.n108 0.306
R20726 VOUT-.n124 VOUT-.n121 0.2825
R20727 VOUT-.n127 VOUT-.n124 0.2825
R20728 VOUT-.n130 VOUT-.n127 0.2825
R20729 VOUT-.n133 VOUT-.n130 0.2825
R20730 VOUT-.n136 VOUT-.n133 0.2825
R20731 VOUT-.n139 VOUT-.n136 0.2825
R20732 VOUT-.n142 VOUT-.n139 0.2825
R20733 VOUT-.n145 VOUT-.n142 0.2825
R20734 VOUT-.n148 VOUT-.n145 0.2825
R20735 VOUT-.n85 VOUT-.n72 0.2825
R20736 VOUT-.n88 VOUT-.n85 0.2825
R20737 VOUT-.n91 VOUT-.n88 0.2825
R20738 VOUT-.n94 VOUT-.n91 0.2825
R20739 VOUT-.n97 VOUT-.n94 0.2825
R20740 VOUT-.n100 VOUT-.n97 0.2825
R20741 VOUT-.n103 VOUT-.n100 0.2825
R20742 VOUT-.n106 VOUT-.n103 0.2825
R20743 VOUT-.n150 VOUT-.n106 0.2825
R20744 VOUT-.n150 VOUT-.n148 0.2825
R20745 VOUT-.n161 VOUT-.n66 0.2455
R20746 VOUT- VOUT-.n176 0.198417
R20747 VOUT-.n176 VOUT-.n175 0.193208
R20748 VOUT- VOUT-.n195 0.182792
R20749 VOUT-.n153 VOUT-.n152 0.138367
R20750 VOUT-.n187 VOUT-.n181 0.0891864
R20751 VOUT-.n60 VOUT-.n59 0.0577917
R20752 VOUT-.n59 VOUT-.n58 0.0577917
R20753 VOUT-.n58 VOUT-.n21 0.0577917
R20754 VOUT-.n54 VOUT-.n21 0.0577917
R20755 VOUT-.n54 VOUT-.n53 0.0577917
R20756 VOUT-.n53 VOUT-.n52 0.0577917
R20757 VOUT-.n52 VOUT-.n25 0.0577917
R20758 VOUT-.n48 VOUT-.n25 0.0577917
R20759 VOUT-.n61 VOUT-.n18 0.0577917
R20760 VOUT-.n57 VOUT-.n18 0.0577917
R20761 VOUT-.n57 VOUT-.n56 0.0577917
R20762 VOUT-.n56 VOUT-.n55 0.0577917
R20763 VOUT-.n55 VOUT-.n22 0.0577917
R20764 VOUT-.n51 VOUT-.n22 0.0577917
R20765 VOUT-.n51 VOUT-.n50 0.0577917
R20766 VOUT-.n49 VOUT-.n48 0.054517
R20767 VOUT-.n168 VOUT-.n167 0.047375
R20768 VOUT-.n172 VOUT-.n171 0.047375
R20769 VOUT-.n162 VOUT-.n7 0.0421667
R20770 VOUT-.n65 VOUT-.n14 0.0421667
R20771 VOUT-.n194 VOUT-.n193 0.0421667
R20772 VOUT-.n193 VOUT-.n192 0.0421667
R20773 VOUT-.n192 VOUT-.n180 0.0421667
R20774 VOUT-.n188 VOUT-.n180 0.0421667
R20775 VOUT-.n188 VOUT-.n187 0.0421667
R20776 VOUT-.n195 VOUT-.n177 0.0421667
R20777 VOUT-.n191 VOUT-.n177 0.0421667
R20778 VOUT-.n191 VOUT-.n190 0.0421667
R20779 VOUT-.n190 VOUT-.n189 0.0421667
R20780 VOUT-.n15 VOUT-.n14 0.0243161
R20781 VOUT-.n17 VOUT-.n9 0.0243161
R20782 VOUT-.n17 VOUT-.n16 0.0243161
R20783 VOUT-.n15 VOUT-.n11 0.0243161
R20784 VOUT-.n159 VOUT-.n3 0.0217373
R20785 VOUT-.n62 VOUT-.n10 0.0217373
R20786 VOUT-.n16 VOUT-.n10 0.0217373
R20787 VOUT-.n69 VOUT-.n3 0.0217373
R20788 VOUT-.n175 VOUT-.n0 0.0217373
R20789 VOUT-.n172 VOUT-.n0 0.0217373
R20790 VOUT-.n67 VOUT-.n7 0.0217373
R20791 VOUT-.n69 VOUT-.n68 0.0217373
R20792 VOUT-.n12 VOUT-.n9 0.0217373
R20793 VOUT-.n12 VOUT-.n11 0.0217373
R20794 VOUT-.n67 VOUT-.n4 0.0217373
R20795 VOUT-.n68 VOUT-.n4 0.0217373
R20796 VOUT-.n169 VOUT-.n164 0.0217373
R20797 VOUT-.n168 VOUT-.n165 0.0217373
R20798 VOUT-.n171 VOUT-.n165 0.0217373
R20799 VOUT-.n167 VOUT-.n164 0.0217373
R20800 VOUT-.n154 VOUT-.n153 0.0161667
R20801 VOUT-.n157 VOUT-.n154 0.0161667
R20802 VOUT-.n155 VOUT-.n6 0.0161667
R20803 VOUT-.n156 VOUT-.n155 0.0161667
R20804 VOUT-.n156 VOUT-.n70 0.0161667
R20805 VOUT-.n160 VOUT-.n5 0.0134654
R20806 VOUT-.n163 VOUT-.n2 0.0134654
R20807 VOUT-.n161 VOUT-.n160 0.0134654
R20808 VOUT-.n5 VOUT-.n2 0.0134654
R20809 VOUT-.n63 VOUT-.n13 0.0109778
R20810 VOUT-.n66 VOUT-.n8 0.0109778
R20811 VOUT-.n173 VOUT-.n1 0.0109778
R20812 VOUT-.n170 VOUT-.n166 0.0109778
R20813 VOUT-.n64 VOUT-.n63 0.0109778
R20814 VOUT-.n13 VOUT-.n8 0.0109778
R20815 VOUT-.n174 VOUT-.n173 0.0109778
R20816 VOUT-.n166 VOUT-.n1 0.0109778
R20817 VOUT-.n158 VOUT-.n70 0.00872683
R20818 two_stage_opamp_dummy_magic_26_0.cap_res_X two_stage_opamp_dummy_magic_26_0.cap_res_X.t0 49.8942
R20819 two_stage_opamp_dummy_magic_26_0.cap_res_X two_stage_opamp_dummy_magic_26_0.cap_res_X.t17 0.9405
R20820 two_stage_opamp_dummy_magic_26_0.cap_res_X.t11 two_stage_opamp_dummy_magic_26_0.cap_res_X.t115 0.1603
R20821 two_stage_opamp_dummy_magic_26_0.cap_res_X.t36 two_stage_opamp_dummy_magic_26_0.cap_res_X.t2 0.1603
R20822 two_stage_opamp_dummy_magic_26_0.cap_res_X.t18 two_stage_opamp_dummy_magic_26_0.cap_res_X.t122 0.1603
R20823 two_stage_opamp_dummy_magic_26_0.cap_res_X.t116 two_stage_opamp_dummy_magic_26_0.cap_res_X.t82 0.1603
R20824 two_stage_opamp_dummy_magic_26_0.cap_res_X.t3 two_stage_opamp_dummy_magic_26_0.cap_res_X.t104 0.1603
R20825 two_stage_opamp_dummy_magic_26_0.cap_res_X.t99 two_stage_opamp_dummy_magic_26_0.cap_res_X.t67 0.1603
R20826 two_stage_opamp_dummy_magic_26_0.cap_res_X.t63 two_stage_opamp_dummy_magic_26_0.cap_res_X.t33 0.1603
R20827 two_stage_opamp_dummy_magic_26_0.cap_res_X.t92 two_stage_opamp_dummy_magic_26_0.cap_res_X.t57 0.1603
R20828 two_stage_opamp_dummy_magic_26_0.cap_res_X.t79 two_stage_opamp_dummy_magic_26_0.cap_res_X.t114 0.1603
R20829 two_stage_opamp_dummy_magic_26_0.cap_res_X.t62 two_stage_opamp_dummy_magic_26_0.cap_res_X.t26 0.1603
R20830 two_stage_opamp_dummy_magic_26_0.cap_res_X.t38 two_stage_opamp_dummy_magic_26_0.cap_res_X.t71 0.1603
R20831 two_stage_opamp_dummy_magic_26_0.cap_res_X.t87 two_stage_opamp_dummy_magic_26_0.cap_res_X.t54 0.1603
R20832 two_stage_opamp_dummy_magic_26_0.cap_res_X.t75 two_stage_opamp_dummy_magic_26_0.cap_res_X.t108 0.1603
R20833 two_stage_opamp_dummy_magic_26_0.cap_res_X.t130 two_stage_opamp_dummy_magic_26_0.cap_res_X.t89 0.1603
R20834 two_stage_opamp_dummy_magic_26_0.cap_res_X.t45 two_stage_opamp_dummy_magic_26_0.cap_res_X.t77 0.1603
R20835 two_stage_opamp_dummy_magic_26_0.cap_res_X.t91 two_stage_opamp_dummy_magic_26_0.cap_res_X.t59 0.1603
R20836 two_stage_opamp_dummy_magic_26_0.cap_res_X.t81 two_stage_opamp_dummy_magic_26_0.cap_res_X.t113 0.1603
R20837 two_stage_opamp_dummy_magic_26_0.cap_res_X.t133 two_stage_opamp_dummy_magic_26_0.cap_res_X.t95 0.1603
R20838 two_stage_opamp_dummy_magic_26_0.cap_res_X.t120 two_stage_opamp_dummy_magic_26_0.cap_res_X.t16 0.1603
R20839 two_stage_opamp_dummy_magic_26_0.cap_res_X.t35 two_stage_opamp_dummy_magic_26_0.cap_res_X.t138 0.1603
R20840 two_stage_opamp_dummy_magic_26_0.cap_res_X.t85 two_stage_opamp_dummy_magic_26_0.cap_res_X.t121 0.1603
R20841 two_stage_opamp_dummy_magic_26_0.cap_res_X.t1 two_stage_opamp_dummy_magic_26_0.cap_res_X.t101 0.1603
R20842 two_stage_opamp_dummy_magic_26_0.cap_res_X.t126 two_stage_opamp_dummy_magic_26_0.cap_res_X.t24 0.1603
R20843 two_stage_opamp_dummy_magic_26_0.cap_res_X.t43 two_stage_opamp_dummy_magic_26_0.cap_res_X.t7 0.1603
R20844 two_stage_opamp_dummy_magic_26_0.cap_res_X.t29 two_stage_opamp_dummy_magic_26_0.cap_res_X.t60 0.1603
R20845 two_stage_opamp_dummy_magic_26_0.cap_res_X.t80 two_stage_opamp_dummy_magic_26_0.cap_res_X.t47 0.1603
R20846 two_stage_opamp_dummy_magic_26_0.cap_res_X.t64 two_stage_opamp_dummy_magic_26_0.cap_res_X.t97 0.1603
R20847 two_stage_opamp_dummy_magic_26_0.cap_res_X.t117 two_stage_opamp_dummy_magic_26_0.cap_res_X.t83 0.1603
R20848 two_stage_opamp_dummy_magic_26_0.cap_res_X.t34 two_stage_opamp_dummy_magic_26_0.cap_res_X.t65 0.1603
R20849 two_stage_opamp_dummy_magic_26_0.cap_res_X.t84 two_stage_opamp_dummy_magic_26_0.cap_res_X.t50 0.1603
R20850 two_stage_opamp_dummy_magic_26_0.cap_res_X.t70 two_stage_opamp_dummy_magic_26_0.cap_res_X.t103 0.1603
R20851 two_stage_opamp_dummy_magic_26_0.cap_res_X.t123 two_stage_opamp_dummy_magic_26_0.cap_res_X.t86 0.1603
R20852 two_stage_opamp_dummy_magic_26_0.cap_res_X.t107 two_stage_opamp_dummy_magic_26_0.cap_res_X.t8 0.1603
R20853 two_stage_opamp_dummy_magic_26_0.cap_res_X.t25 two_stage_opamp_dummy_magic_26_0.cap_res_X.t128 0.1603
R20854 two_stage_opamp_dummy_magic_26_0.cap_res_X.t76 two_stage_opamp_dummy_magic_26_0.cap_res_X.t109 0.1603
R20855 two_stage_opamp_dummy_magic_26_0.cap_res_X.t129 two_stage_opamp_dummy_magic_26_0.cap_res_X.t90 0.1603
R20856 two_stage_opamp_dummy_magic_26_0.cap_res_X.t44 two_stage_opamp_dummy_magic_26_0.cap_res_X.t127 0.1603
R20857 two_stage_opamp_dummy_magic_26_0.cap_res_X.t48 two_stage_opamp_dummy_magic_26_0.cap_res_X.t94 0.1603
R20858 two_stage_opamp_dummy_magic_26_0.cap_res_X.t124 two_stage_opamp_dummy_magic_26_0.cap_res_X.t22 0.1603
R20859 two_stage_opamp_dummy_magic_26_0.cap_res_X.t42 two_stage_opamp_dummy_magic_26_0.cap_res_X.t5 0.1603
R20860 two_stage_opamp_dummy_magic_26_0.cap_res_X.t21 two_stage_opamp_dummy_magic_26_0.cap_res_X.t55 0.1603
R20861 two_stage_opamp_dummy_magic_26_0.cap_res_X.t72 two_stage_opamp_dummy_magic_26_0.cap_res_X.t41 0.1603
R20862 two_stage_opamp_dummy_magic_26_0.cap_res_X.t53 two_stage_opamp_dummy_magic_26_0.cap_res_X.t12 0.1603
R20863 two_stage_opamp_dummy_magic_26_0.cap_res_X.t78 two_stage_opamp_dummy_magic_26_0.cap_res_X.t39 0.1603
R20864 two_stage_opamp_dummy_magic_26_0.cap_res_X.t56 two_stage_opamp_dummy_magic_26_0.cap_res_X.t19 0.1603
R20865 two_stage_opamp_dummy_magic_26_0.cap_res_X.t23 two_stage_opamp_dummy_magic_26_0.cap_res_X.t119 0.1603
R20866 two_stage_opamp_dummy_magic_26_0.cap_res_X.t46 two_stage_opamp_dummy_magic_26_0.cap_res_X.t4 0.1603
R20867 two_stage_opamp_dummy_magic_26_0.cap_res_X.t6 two_stage_opamp_dummy_magic_26_0.cap_res_X.t100 0.1603
R20868 two_stage_opamp_dummy_magic_26_0.cap_res_X.t105 two_stage_opamp_dummy_magic_26_0.cap_res_X.t66 0.1603
R20869 two_stage_opamp_dummy_magic_26_0.cap_res_X.t68 two_stage_opamp_dummy_magic_26_0.cap_res_X.t31 0.1603
R20870 two_stage_opamp_dummy_magic_26_0.cap_res_X.t88 two_stage_opamp_dummy_magic_26_0.cap_res_X.t51 0.1603
R20871 two_stage_opamp_dummy_magic_26_0.cap_res_X.t52 two_stage_opamp_dummy_magic_26_0.cap_res_X.t10 0.1603
R20872 two_stage_opamp_dummy_magic_26_0.cap_res_X.t14 two_stage_opamp_dummy_magic_26_0.cap_res_X.t111 0.1603
R20873 two_stage_opamp_dummy_magic_26_0.cap_res_X.t137 two_stage_opamp_dummy_magic_26_0.cap_res_X.t98 0.1603
R20874 two_stage_opamp_dummy_magic_26_0.cap_res_X.t93 two_stage_opamp_dummy_magic_26_0.cap_res_X.t61 0.1603
R20875 two_stage_opamp_dummy_magic_26_0.cap_res_X.t9 two_stage_opamp_dummy_magic_26_0.cap_res_X.t110 0.1603
R20876 two_stage_opamp_dummy_magic_26_0.cap_res_X.t13 two_stage_opamp_dummy_magic_26_0.cap_res_X.t102 0.1603
R20877 two_stage_opamp_dummy_magic_26_0.cap_res_X.t49 two_stage_opamp_dummy_magic_26_0.cap_res_X.t13 0.1603
R20878 two_stage_opamp_dummy_magic_26_0.cap_res_X.t132 two_stage_opamp_dummy_magic_26_0.cap_res_X.t30 0.1603
R20879 two_stage_opamp_dummy_magic_26_0.cap_res_X.t17 two_stage_opamp_dummy_magic_26_0.cap_res_X.t132 0.1603
R20880 two_stage_opamp_dummy_magic_26_0.cap_res_X.t40 two_stage_opamp_dummy_magic_26_0.cap_res_X.n10 0.159278
R20881 two_stage_opamp_dummy_magic_26_0.cap_res_X.t106 two_stage_opamp_dummy_magic_26_0.cap_res_X.n11 0.159278
R20882 two_stage_opamp_dummy_magic_26_0.cap_res_X.t73 two_stage_opamp_dummy_magic_26_0.cap_res_X.n12 0.159278
R20883 two_stage_opamp_dummy_magic_26_0.cap_res_X.t136 two_stage_opamp_dummy_magic_26_0.cap_res_X.n13 0.159278
R20884 two_stage_opamp_dummy_magic_26_0.cap_res_X.t28 two_stage_opamp_dummy_magic_26_0.cap_res_X.n14 0.159278
R20885 two_stage_opamp_dummy_magic_26_0.cap_res_X.t58 two_stage_opamp_dummy_magic_26_0.cap_res_X.n15 0.159278
R20886 two_stage_opamp_dummy_magic_26_0.cap_res_X.t20 two_stage_opamp_dummy_magic_26_0.cap_res_X.n16 0.159278
R20887 two_stage_opamp_dummy_magic_26_0.cap_res_X.t118 two_stage_opamp_dummy_magic_26_0.cap_res_X.n17 0.159278
R20888 two_stage_opamp_dummy_magic_26_0.cap_res_X.t15 two_stage_opamp_dummy_magic_26_0.cap_res_X.n18 0.159278
R20889 two_stage_opamp_dummy_magic_26_0.cap_res_X.t112 two_stage_opamp_dummy_magic_26_0.cap_res_X.n19 0.159278
R20890 two_stage_opamp_dummy_magic_26_0.cap_res_X.t74 two_stage_opamp_dummy_magic_26_0.cap_res_X.n20 0.159278
R20891 two_stage_opamp_dummy_magic_26_0.cap_res_X.t37 two_stage_opamp_dummy_magic_26_0.cap_res_X.n21 0.159278
R20892 two_stage_opamp_dummy_magic_26_0.cap_res_X.t69 two_stage_opamp_dummy_magic_26_0.cap_res_X.n22 0.159278
R20893 two_stage_opamp_dummy_magic_26_0.cap_res_X.t32 two_stage_opamp_dummy_magic_26_0.cap_res_X.n23 0.159278
R20894 two_stage_opamp_dummy_magic_26_0.cap_res_X.t131 two_stage_opamp_dummy_magic_26_0.cap_res_X.n24 0.159278
R20895 two_stage_opamp_dummy_magic_26_0.cap_res_X.t27 two_stage_opamp_dummy_magic_26_0.cap_res_X.n25 0.159278
R20896 two_stage_opamp_dummy_magic_26_0.cap_res_X.t125 two_stage_opamp_dummy_magic_26_0.cap_res_X.n26 0.159278
R20897 two_stage_opamp_dummy_magic_26_0.cap_res_X.t96 two_stage_opamp_dummy_magic_26_0.cap_res_X.n27 0.159278
R20898 two_stage_opamp_dummy_magic_26_0.cap_res_X.t134 two_stage_opamp_dummy_magic_26_0.cap_res_X.n28 0.159278
R20899 two_stage_opamp_dummy_magic_26_0.cap_res_X.n29 two_stage_opamp_dummy_magic_26_0.cap_res_X.t92 0.1368
R20900 two_stage_opamp_dummy_magic_26_0.cap_res_X.n28 two_stage_opamp_dummy_magic_26_0.cap_res_X.t79 0.1368
R20901 two_stage_opamp_dummy_magic_26_0.cap_res_X.n28 two_stage_opamp_dummy_magic_26_0.cap_res_X.t62 0.1368
R20902 two_stage_opamp_dummy_magic_26_0.cap_res_X.n27 two_stage_opamp_dummy_magic_26_0.cap_res_X.t38 0.1368
R20903 two_stage_opamp_dummy_magic_26_0.cap_res_X.n27 two_stage_opamp_dummy_magic_26_0.cap_res_X.t87 0.1368
R20904 two_stage_opamp_dummy_magic_26_0.cap_res_X.n26 two_stage_opamp_dummy_magic_26_0.cap_res_X.t75 0.1368
R20905 two_stage_opamp_dummy_magic_26_0.cap_res_X.n26 two_stage_opamp_dummy_magic_26_0.cap_res_X.t130 0.1368
R20906 two_stage_opamp_dummy_magic_26_0.cap_res_X.n25 two_stage_opamp_dummy_magic_26_0.cap_res_X.t45 0.1368
R20907 two_stage_opamp_dummy_magic_26_0.cap_res_X.n25 two_stage_opamp_dummy_magic_26_0.cap_res_X.t91 0.1368
R20908 two_stage_opamp_dummy_magic_26_0.cap_res_X.n24 two_stage_opamp_dummy_magic_26_0.cap_res_X.t81 0.1368
R20909 two_stage_opamp_dummy_magic_26_0.cap_res_X.n24 two_stage_opamp_dummy_magic_26_0.cap_res_X.t133 0.1368
R20910 two_stage_opamp_dummy_magic_26_0.cap_res_X.n23 two_stage_opamp_dummy_magic_26_0.cap_res_X.t120 0.1368
R20911 two_stage_opamp_dummy_magic_26_0.cap_res_X.n23 two_stage_opamp_dummy_magic_26_0.cap_res_X.t35 0.1368
R20912 two_stage_opamp_dummy_magic_26_0.cap_res_X.n22 two_stage_opamp_dummy_magic_26_0.cap_res_X.t85 0.1368
R20913 two_stage_opamp_dummy_magic_26_0.cap_res_X.n22 two_stage_opamp_dummy_magic_26_0.cap_res_X.t1 0.1368
R20914 two_stage_opamp_dummy_magic_26_0.cap_res_X.n21 two_stage_opamp_dummy_magic_26_0.cap_res_X.t126 0.1368
R20915 two_stage_opamp_dummy_magic_26_0.cap_res_X.n21 two_stage_opamp_dummy_magic_26_0.cap_res_X.t43 0.1368
R20916 two_stage_opamp_dummy_magic_26_0.cap_res_X.n20 two_stage_opamp_dummy_magic_26_0.cap_res_X.t29 0.1368
R20917 two_stage_opamp_dummy_magic_26_0.cap_res_X.n20 two_stage_opamp_dummy_magic_26_0.cap_res_X.t80 0.1368
R20918 two_stage_opamp_dummy_magic_26_0.cap_res_X.n19 two_stage_opamp_dummy_magic_26_0.cap_res_X.t64 0.1368
R20919 two_stage_opamp_dummy_magic_26_0.cap_res_X.n19 two_stage_opamp_dummy_magic_26_0.cap_res_X.t117 0.1368
R20920 two_stage_opamp_dummy_magic_26_0.cap_res_X.n18 two_stage_opamp_dummy_magic_26_0.cap_res_X.t34 0.1368
R20921 two_stage_opamp_dummy_magic_26_0.cap_res_X.n18 two_stage_opamp_dummy_magic_26_0.cap_res_X.t84 0.1368
R20922 two_stage_opamp_dummy_magic_26_0.cap_res_X.n17 two_stage_opamp_dummy_magic_26_0.cap_res_X.t70 0.1368
R20923 two_stage_opamp_dummy_magic_26_0.cap_res_X.n17 two_stage_opamp_dummy_magic_26_0.cap_res_X.t123 0.1368
R20924 two_stage_opamp_dummy_magic_26_0.cap_res_X.n16 two_stage_opamp_dummy_magic_26_0.cap_res_X.t107 0.1368
R20925 two_stage_opamp_dummy_magic_26_0.cap_res_X.n16 two_stage_opamp_dummy_magic_26_0.cap_res_X.t25 0.1368
R20926 two_stage_opamp_dummy_magic_26_0.cap_res_X.n15 two_stage_opamp_dummy_magic_26_0.cap_res_X.t76 0.1368
R20927 two_stage_opamp_dummy_magic_26_0.cap_res_X.n15 two_stage_opamp_dummy_magic_26_0.cap_res_X.t129 0.1368
R20928 two_stage_opamp_dummy_magic_26_0.cap_res_X.n14 two_stage_opamp_dummy_magic_26_0.cap_res_X.t44 0.1368
R20929 two_stage_opamp_dummy_magic_26_0.cap_res_X.n14 two_stage_opamp_dummy_magic_26_0.cap_res_X.t48 0.1368
R20930 two_stage_opamp_dummy_magic_26_0.cap_res_X.n13 two_stage_opamp_dummy_magic_26_0.cap_res_X.t124 0.1368
R20931 two_stage_opamp_dummy_magic_26_0.cap_res_X.n13 two_stage_opamp_dummy_magic_26_0.cap_res_X.t42 0.1368
R20932 two_stage_opamp_dummy_magic_26_0.cap_res_X.n12 two_stage_opamp_dummy_magic_26_0.cap_res_X.t21 0.1368
R20933 two_stage_opamp_dummy_magic_26_0.cap_res_X.n12 two_stage_opamp_dummy_magic_26_0.cap_res_X.t72 0.1368
R20934 two_stage_opamp_dummy_magic_26_0.cap_res_X.n11 two_stage_opamp_dummy_magic_26_0.cap_res_X.t137 0.1368
R20935 two_stage_opamp_dummy_magic_26_0.cap_res_X.n10 two_stage_opamp_dummy_magic_26_0.cap_res_X.t93 0.1368
R20936 two_stage_opamp_dummy_magic_26_0.cap_res_X.t110 two_stage_opamp_dummy_magic_26_0.cap_res_X.n29 0.1368
R20937 two_stage_opamp_dummy_magic_26_0.cap_res_X.n30 two_stage_opamp_dummy_magic_26_0.cap_res_X.t9 0.1368
R20938 two_stage_opamp_dummy_magic_26_0.cap_res_X.n31 two_stage_opamp_dummy_magic_26_0.cap_res_X.t11 0.114322
R20939 two_stage_opamp_dummy_magic_26_0.cap_res_X.n0 two_stage_opamp_dummy_magic_26_0.cap_res_X.t53 0.114322
R20940 two_stage_opamp_dummy_magic_26_0.cap_res_X.n32 two_stage_opamp_dummy_magic_26_0.cap_res_X.n31 0.1133
R20941 two_stage_opamp_dummy_magic_26_0.cap_res_X.n33 two_stage_opamp_dummy_magic_26_0.cap_res_X.n32 0.1133
R20942 two_stage_opamp_dummy_magic_26_0.cap_res_X.n34 two_stage_opamp_dummy_magic_26_0.cap_res_X.n33 0.1133
R20943 two_stage_opamp_dummy_magic_26_0.cap_res_X.n35 two_stage_opamp_dummy_magic_26_0.cap_res_X.n34 0.1133
R20944 two_stage_opamp_dummy_magic_26_0.cap_res_X.n36 two_stage_opamp_dummy_magic_26_0.cap_res_X.n35 0.1133
R20945 two_stage_opamp_dummy_magic_26_0.cap_res_X.n1 two_stage_opamp_dummy_magic_26_0.cap_res_X.n0 0.1133
R20946 two_stage_opamp_dummy_magic_26_0.cap_res_X.n2 two_stage_opamp_dummy_magic_26_0.cap_res_X.n1 0.1133
R20947 two_stage_opamp_dummy_magic_26_0.cap_res_X.n3 two_stage_opamp_dummy_magic_26_0.cap_res_X.n2 0.1133
R20948 two_stage_opamp_dummy_magic_26_0.cap_res_X.n4 two_stage_opamp_dummy_magic_26_0.cap_res_X.n3 0.1133
R20949 two_stage_opamp_dummy_magic_26_0.cap_res_X.n5 two_stage_opamp_dummy_magic_26_0.cap_res_X.n4 0.1133
R20950 two_stage_opamp_dummy_magic_26_0.cap_res_X.n6 two_stage_opamp_dummy_magic_26_0.cap_res_X.n5 0.1133
R20951 two_stage_opamp_dummy_magic_26_0.cap_res_X.n7 two_stage_opamp_dummy_magic_26_0.cap_res_X.n6 0.1133
R20952 two_stage_opamp_dummy_magic_26_0.cap_res_X.n8 two_stage_opamp_dummy_magic_26_0.cap_res_X.n7 0.1133
R20953 two_stage_opamp_dummy_magic_26_0.cap_res_X.n9 two_stage_opamp_dummy_magic_26_0.cap_res_X.n8 0.1133
R20954 two_stage_opamp_dummy_magic_26_0.cap_res_X.n11 two_stage_opamp_dummy_magic_26_0.cap_res_X.n9 0.1133
R20955 two_stage_opamp_dummy_magic_26_0.cap_res_X.n37 two_stage_opamp_dummy_magic_26_0.cap_res_X.n30 0.1133
R20956 two_stage_opamp_dummy_magic_26_0.cap_res_X.n37 two_stage_opamp_dummy_magic_26_0.cap_res_X.n36 0.1133
R20957 two_stage_opamp_dummy_magic_26_0.cap_res_X.n31 two_stage_opamp_dummy_magic_26_0.cap_res_X.t36 0.00152174
R20958 two_stage_opamp_dummy_magic_26_0.cap_res_X.n32 two_stage_opamp_dummy_magic_26_0.cap_res_X.t18 0.00152174
R20959 two_stage_opamp_dummy_magic_26_0.cap_res_X.n33 two_stage_opamp_dummy_magic_26_0.cap_res_X.t116 0.00152174
R20960 two_stage_opamp_dummy_magic_26_0.cap_res_X.n34 two_stage_opamp_dummy_magic_26_0.cap_res_X.t3 0.00152174
R20961 two_stage_opamp_dummy_magic_26_0.cap_res_X.n35 two_stage_opamp_dummy_magic_26_0.cap_res_X.t99 0.00152174
R20962 two_stage_opamp_dummy_magic_26_0.cap_res_X.n36 two_stage_opamp_dummy_magic_26_0.cap_res_X.t63 0.00152174
R20963 two_stage_opamp_dummy_magic_26_0.cap_res_X.n0 two_stage_opamp_dummy_magic_26_0.cap_res_X.t78 0.00152174
R20964 two_stage_opamp_dummy_magic_26_0.cap_res_X.n1 two_stage_opamp_dummy_magic_26_0.cap_res_X.t56 0.00152174
R20965 two_stage_opamp_dummy_magic_26_0.cap_res_X.n2 two_stage_opamp_dummy_magic_26_0.cap_res_X.t23 0.00152174
R20966 two_stage_opamp_dummy_magic_26_0.cap_res_X.n3 two_stage_opamp_dummy_magic_26_0.cap_res_X.t46 0.00152174
R20967 two_stage_opamp_dummy_magic_26_0.cap_res_X.n4 two_stage_opamp_dummy_magic_26_0.cap_res_X.t6 0.00152174
R20968 two_stage_opamp_dummy_magic_26_0.cap_res_X.n5 two_stage_opamp_dummy_magic_26_0.cap_res_X.t105 0.00152174
R20969 two_stage_opamp_dummy_magic_26_0.cap_res_X.n6 two_stage_opamp_dummy_magic_26_0.cap_res_X.t68 0.00152174
R20970 two_stage_opamp_dummy_magic_26_0.cap_res_X.n7 two_stage_opamp_dummy_magic_26_0.cap_res_X.t88 0.00152174
R20971 two_stage_opamp_dummy_magic_26_0.cap_res_X.n8 two_stage_opamp_dummy_magic_26_0.cap_res_X.t52 0.00152174
R20972 two_stage_opamp_dummy_magic_26_0.cap_res_X.n9 two_stage_opamp_dummy_magic_26_0.cap_res_X.t14 0.00152174
R20973 two_stage_opamp_dummy_magic_26_0.cap_res_X.n10 two_stage_opamp_dummy_magic_26_0.cap_res_X.t135 0.00152174
R20974 two_stage_opamp_dummy_magic_26_0.cap_res_X.n11 two_stage_opamp_dummy_magic_26_0.cap_res_X.t40 0.00152174
R20975 two_stage_opamp_dummy_magic_26_0.cap_res_X.n12 two_stage_opamp_dummy_magic_26_0.cap_res_X.t106 0.00152174
R20976 two_stage_opamp_dummy_magic_26_0.cap_res_X.n13 two_stage_opamp_dummy_magic_26_0.cap_res_X.t73 0.00152174
R20977 two_stage_opamp_dummy_magic_26_0.cap_res_X.n14 two_stage_opamp_dummy_magic_26_0.cap_res_X.t136 0.00152174
R20978 two_stage_opamp_dummy_magic_26_0.cap_res_X.n15 two_stage_opamp_dummy_magic_26_0.cap_res_X.t28 0.00152174
R20979 two_stage_opamp_dummy_magic_26_0.cap_res_X.n16 two_stage_opamp_dummy_magic_26_0.cap_res_X.t58 0.00152174
R20980 two_stage_opamp_dummy_magic_26_0.cap_res_X.n17 two_stage_opamp_dummy_magic_26_0.cap_res_X.t20 0.00152174
R20981 two_stage_opamp_dummy_magic_26_0.cap_res_X.n18 two_stage_opamp_dummy_magic_26_0.cap_res_X.t118 0.00152174
R20982 two_stage_opamp_dummy_magic_26_0.cap_res_X.n19 two_stage_opamp_dummy_magic_26_0.cap_res_X.t15 0.00152174
R20983 two_stage_opamp_dummy_magic_26_0.cap_res_X.n20 two_stage_opamp_dummy_magic_26_0.cap_res_X.t112 0.00152174
R20984 two_stage_opamp_dummy_magic_26_0.cap_res_X.n21 two_stage_opamp_dummy_magic_26_0.cap_res_X.t74 0.00152174
R20985 two_stage_opamp_dummy_magic_26_0.cap_res_X.n22 two_stage_opamp_dummy_magic_26_0.cap_res_X.t37 0.00152174
R20986 two_stage_opamp_dummy_magic_26_0.cap_res_X.n23 two_stage_opamp_dummy_magic_26_0.cap_res_X.t69 0.00152174
R20987 two_stage_opamp_dummy_magic_26_0.cap_res_X.n24 two_stage_opamp_dummy_magic_26_0.cap_res_X.t32 0.00152174
R20988 two_stage_opamp_dummy_magic_26_0.cap_res_X.n25 two_stage_opamp_dummy_magic_26_0.cap_res_X.t131 0.00152174
R20989 two_stage_opamp_dummy_magic_26_0.cap_res_X.n26 two_stage_opamp_dummy_magic_26_0.cap_res_X.t27 0.00152174
R20990 two_stage_opamp_dummy_magic_26_0.cap_res_X.n27 two_stage_opamp_dummy_magic_26_0.cap_res_X.t125 0.00152174
R20991 two_stage_opamp_dummy_magic_26_0.cap_res_X.n28 two_stage_opamp_dummy_magic_26_0.cap_res_X.t96 0.00152174
R20992 two_stage_opamp_dummy_magic_26_0.cap_res_X.n29 two_stage_opamp_dummy_magic_26_0.cap_res_X.t134 0.00152174
R20993 two_stage_opamp_dummy_magic_26_0.cap_res_X.n30 two_stage_opamp_dummy_magic_26_0.cap_res_X.t49 0.00152174
R20994 two_stage_opamp_dummy_magic_26_0.cap_res_X.t30 two_stage_opamp_dummy_magic_26_0.cap_res_X.n37 0.00152174
R20995 VOUT+.n194 VOUT+.t7 110.386
R20996 VOUT+.n47 VOUT+.n46 34.9935
R20997 VOUT+.n45 VOUT+.n44 34.9935
R20998 VOUT+.n59 VOUT+.n58 34.9935
R20999 VOUT+.n55 VOUT+.n54 34.9935
R21000 VOUT+.n52 VOUT+.n51 34.9935
R21001 VOUT+.n49 VOUT+.n48 34.9935
R21002 VOUT+.n2 VOUT+.n1 9.73997
R21003 VOUT+.n6 VOUT+.n5 9.73997
R21004 VOUT+.n9 VOUT+.n8 9.73997
R21005 VOUT+.n7 VOUT+.n6 6.64633
R21006 VOUT+.n7 VOUT+.n2 6.64633
R21007 VOUT+.n46 VOUT+.t2 6.56717
R21008 VOUT+.n46 VOUT+.t14 6.56717
R21009 VOUT+.n44 VOUT+.t13 6.56717
R21010 VOUT+.n44 VOUT+.t9 6.56717
R21011 VOUT+.n58 VOUT+.t4 6.56717
R21012 VOUT+.n58 VOUT+.t8 6.56717
R21013 VOUT+.n54 VOUT+.t12 6.56717
R21014 VOUT+.n54 VOUT+.t1 6.56717
R21015 VOUT+.n51 VOUT+.t10 6.56717
R21016 VOUT+.n51 VOUT+.t18 6.56717
R21017 VOUT+.n48 VOUT+.t17 6.56717
R21018 VOUT+.n48 VOUT+.t16 6.56717
R21019 VOUT+.n57 VOUT+.n45 6.3755
R21020 VOUT+.n50 VOUT+.n47 6.3755
R21021 VOUT+.n9 VOUT+.n7 6.02133
R21022 VOUT+.n59 VOUT+.n57 5.813
R21023 VOUT+.n56 VOUT+.n55 5.813
R21024 VOUT+.n53 VOUT+.n52 5.813
R21025 VOUT+.n50 VOUT+.n49 5.813
R21026 VOUT+.n60 VOUT+.n36 5.063
R21027 VOUT+.n63 VOUT+.n43 5.063
R21028 VOUT+.n133 VOUT+.t51 4.8295
R21029 VOUT+.n134 VOUT+.t86 4.8295
R21030 VOUT+.n146 VOUT+.t144 4.8295
R21031 VOUT+.n148 VOUT+.t122 4.8295
R21032 VOUT+.n149 VOUT+.t32 4.8295
R21033 VOUT+.n151 VOUT+.t138 4.8295
R21034 VOUT+.n152 VOUT+.t26 4.8295
R21035 VOUT+.n154 VOUT+.t104 4.8295
R21036 VOUT+.n155 VOUT+.t131 4.8295
R21037 VOUT+.n157 VOUT+.t132 4.8295
R21038 VOUT+.n158 VOUT+.t21 4.8295
R21039 VOUT+.n160 VOUT+.t96 4.8295
R21040 VOUT+.n161 VOUT+.t125 4.8295
R21041 VOUT+.n163 VOUT+.t58 4.8295
R21042 VOUT+.n164 VOUT+.t88 4.8295
R21043 VOUT+.n166 VOUT+.t90 4.8295
R21044 VOUT+.n167 VOUT+.t123 4.8295
R21045 VOUT+.n169 VOUT+.t48 4.8295
R21046 VOUT+.n170 VOUT+.t80 4.8295
R21047 VOUT+.n172 VOUT+.t149 4.8295
R21048 VOUT+.n173 VOUT+.t38 4.8295
R21049 VOUT+.n97 VOUT+.t141 4.8295
R21050 VOUT+.n110 VOUT+.t107 4.8295
R21051 VOUT+.n112 VOUT+.t155 4.8295
R21052 VOUT+.n113 VOUT+.t46 4.8295
R21053 VOUT+.n115 VOUT+.t50 4.8295
R21054 VOUT+.n116 VOUT+.t82 4.8295
R21055 VOUT+.n118 VOUT+.t40 4.8295
R21056 VOUT+.n119 VOUT+.t47 4.8295
R21057 VOUT+.n121 VOUT+.t103 4.8295
R21058 VOUT+.n122 VOUT+.t130 4.8295
R21059 VOUT+.n124 VOUT+.t66 4.8295
R21060 VOUT+.n125 VOUT+.t99 4.8295
R21061 VOUT+.n127 VOUT+.t109 4.8295
R21062 VOUT+.n128 VOUT+.t136 4.8295
R21063 VOUT+.n130 VOUT+.t145 4.8295
R21064 VOUT+.n131 VOUT+.t31 4.8295
R21065 VOUT+.n175 VOUT+.t142 4.8295
R21066 VOUT+.n139 VOUT+.t54 4.8154
R21067 VOUT+.n138 VOUT+.t89 4.8154
R21068 VOUT+.n136 VOUT+.t110 4.8154
R21069 VOUT+.n135 VOUT+.t143 4.8154
R21070 VOUT+.n141 VOUT+.t28 4.806
R21071 VOUT+.n140 VOUT+.t151 4.806
R21072 VOUT+.n137 VOUT+.t124 4.806
R21073 VOUT+.n109 VOUT+.t44 4.806
R21074 VOUT+.n108 VOUT+.t83 4.806
R21075 VOUT+.n107 VOUT+.t62 4.806
R21076 VOUT+.n106 VOUT+.t105 4.806
R21077 VOUT+.n105 VOUT+.t137 4.806
R21078 VOUT+.n104 VOUT+.t119 4.806
R21079 VOUT+.n103 VOUT+.t153 4.806
R21080 VOUT+.n102 VOUT+.t55 4.806
R21081 VOUT+.n101 VOUT+.t92 4.806
R21082 VOUT+.n100 VOUT+.t68 4.806
R21083 VOUT+.n99 VOUT+.t111 4.806
R21084 VOUT+.n133 VOUT+.t101 4.5005
R21085 VOUT+.n134 VOUT+.t135 4.5005
R21086 VOUT+.n135 VOUT+.t113 4.5005
R21087 VOUT+.n136 VOUT+.t70 4.5005
R21088 VOUT+.n137 VOUT+.t94 4.5005
R21089 VOUT+.n138 VOUT+.t56 4.5005
R21090 VOUT+.n139 VOUT+.t156 4.5005
R21091 VOUT+.n140 VOUT+.t120 4.5005
R21092 VOUT+.n141 VOUT+.t139 4.5005
R21093 VOUT+.n142 VOUT+.t106 4.5005
R21094 VOUT+.n143 VOUT+.t63 4.5005
R21095 VOUT+.n144 VOUT+.t87 4.5005
R21096 VOUT+.n145 VOUT+.t45 4.5005
R21097 VOUT+.n147 VOUT+.t39 4.5005
R21098 VOUT+.n146 VOUT+.t75 4.5005
R21099 VOUT+.n148 VOUT+.t81 4.5005
R21100 VOUT+.n150 VOUT+.t77 4.5005
R21101 VOUT+.n149 VOUT+.t116 4.5005
R21102 VOUT+.n151 VOUT+.t108 4.5005
R21103 VOUT+.n153 VOUT+.t78 4.5005
R21104 VOUT+.n152 VOUT+.t79 4.5005
R21105 VOUT+.n154 VOUT+.t65 4.5005
R21106 VOUT+.n156 VOUT+.t34 4.5005
R21107 VOUT+.n155 VOUT+.t36 4.5005
R21108 VOUT+.n157 VOUT+.t102 4.5005
R21109 VOUT+.n159 VOUT+.t73 4.5005
R21110 VOUT+.n158 VOUT+.t74 4.5005
R21111 VOUT+.n160 VOUT+.t60 4.5005
R21112 VOUT+.n162 VOUT+.t29 4.5005
R21113 VOUT+.n161 VOUT+.t30 4.5005
R21114 VOUT+.n163 VOUT+.t19 4.5005
R21115 VOUT+.n165 VOUT+.t133 4.5005
R21116 VOUT+.n164 VOUT+.t134 4.5005
R21117 VOUT+.n166 VOUT+.t57 4.5005
R21118 VOUT+.n168 VOUT+.t24 4.5005
R21119 VOUT+.n167 VOUT+.t25 4.5005
R21120 VOUT+.n169 VOUT+.t152 4.5005
R21121 VOUT+.n171 VOUT+.t126 4.5005
R21122 VOUT+.n170 VOUT+.t127 4.5005
R21123 VOUT+.n172 VOUT+.t117 4.5005
R21124 VOUT+.n174 VOUT+.t91 4.5005
R21125 VOUT+.n173 VOUT+.t93 4.5005
R21126 VOUT+.n98 VOUT+.t37 4.5005
R21127 VOUT+.n97 VOUT+.t71 4.5005
R21128 VOUT+.n99 VOUT+.t67 4.5005
R21129 VOUT+.n100 VOUT+.t22 4.5005
R21130 VOUT+.n101 VOUT+.t52 4.5005
R21131 VOUT+.n102 VOUT+.t150 4.5005
R21132 VOUT+.n103 VOUT+.t118 4.5005
R21133 VOUT+.n104 VOUT+.t76 4.5005
R21134 VOUT+.n105 VOUT+.t100 4.5005
R21135 VOUT+.n106 VOUT+.t61 4.5005
R21136 VOUT+.n107 VOUT+.t20 4.5005
R21137 VOUT+.n108 VOUT+.t41 4.5005
R21138 VOUT+.n109 VOUT+.t148 4.5005
R21139 VOUT+.n111 VOUT+.t140 4.5005
R21140 VOUT+.n110 VOUT+.t27 4.5005
R21141 VOUT+.n112 VOUT+.t121 4.5005
R21142 VOUT+.n114 VOUT+.t97 4.5005
R21143 VOUT+.n113 VOUT+.t98 4.5005
R21144 VOUT+.n115 VOUT+.t154 4.5005
R21145 VOUT+.n117 VOUT+.t128 4.5005
R21146 VOUT+.n116 VOUT+.t129 4.5005
R21147 VOUT+.n118 VOUT+.t95 4.5005
R21148 VOUT+.n120 VOUT+.t59 4.5005
R21149 VOUT+.n119 VOUT+.t112 4.5005
R21150 VOUT+.n121 VOUT+.t64 4.5005
R21151 VOUT+.n123 VOUT+.t33 4.5005
R21152 VOUT+.n122 VOUT+.t35 4.5005
R21153 VOUT+.n124 VOUT+.t23 4.5005
R21154 VOUT+.n126 VOUT+.t146 4.5005
R21155 VOUT+.n125 VOUT+.t147 4.5005
R21156 VOUT+.n127 VOUT+.t69 4.5005
R21157 VOUT+.n129 VOUT+.t42 4.5005
R21158 VOUT+.n128 VOUT+.t43 4.5005
R21159 VOUT+.n130 VOUT+.t114 4.5005
R21160 VOUT+.n132 VOUT+.t84 4.5005
R21161 VOUT+.n131 VOUT+.t85 4.5005
R21162 VOUT+.n177 VOUT+.t72 4.5005
R21163 VOUT+.n176 VOUT+.t49 4.5005
R21164 VOUT+.n175 VOUT+.t53 4.5005
R21165 VOUT+.n178 VOUT+.t115 4.5005
R21166 VOUT+.n60 VOUT+.n37 4.5005
R21167 VOUT+.n61 VOUT+.n40 4.5005
R21168 VOUT+.n62 VOUT+.n41 4.5005
R21169 VOUT+.n64 VOUT+.n63 4.5005
R21170 VOUT+.n87 VOUT+.n86 4.5005
R21171 VOUT+.n83 VOUT+.n80 4.5005
R21172 VOUT+.n87 VOUT+.n80 4.5005
R21173 VOUT+.n88 VOUT+.n32 4.5005
R21174 VOUT+.n88 VOUT+.n34 4.5005
R21175 VOUT+.n88 VOUT+.n87 4.5005
R21176 VOUT+.n183 VOUT+.n91 4.5005
R21177 VOUT+.n184 VOUT+.n183 4.5005
R21178 VOUT+.n184 VOUT+.n28 4.5005
R21179 VOUT+.n185 VOUT+.n27 4.5005
R21180 VOUT+.n185 VOUT+.n184 4.5005
R21181 VOUT+.n189 VOUT+.n188 4.5005
R21182 VOUT+.n188 VOUT+.n19 4.5005
R21183 VOUT+.n22 VOUT+.n19 4.5005
R21184 VOUT+.n191 VOUT+.n19 4.5005
R21185 VOUT+.n193 VOUT+.n19 4.5005
R21186 VOUT+.n192 VOUT+.n22 4.5005
R21187 VOUT+.n192 VOUT+.n191 4.5005
R21188 VOUT+.n193 VOUT+.n192 4.5005
R21189 VOUT+.n1 VOUT+.t11 3.42907
R21190 VOUT+.n1 VOUT+.t5 3.42907
R21191 VOUT+.n5 VOUT+.t6 3.42907
R21192 VOUT+.n5 VOUT+.t3 3.42907
R21193 VOUT+.n8 VOUT+.t15 3.42907
R21194 VOUT+.n8 VOUT+.t0 3.42907
R21195 VOUT+.n85 VOUT+.n33 2.26725
R21196 VOUT+.n81 VOUT+.n31 2.24601
R21197 VOUT+.n187 VOUT+.n186 2.24601
R21198 VOUT+.n24 VOUT+.n21 2.24601
R21199 VOUT+.n182 VOUT+.n181 2.24477
R21200 VOUT+.n30 VOUT+.n25 2.24477
R21201 VOUT+.n88 VOUT+.n33 2.24063
R21202 VOUT+.n185 VOUT+.n26 2.24063
R21203 VOUT+.n192 VOUT+.n23 2.24063
R21204 VOUT+.n80 VOUT+.n79 2.24063
R21205 VOUT+.n183 VOUT+.n89 2.24063
R21206 VOUT+.n90 VOUT+.n28 2.24063
R21207 VOUT+.n190 VOUT+.n189 2.24063
R21208 VOUT+.n189 VOUT+.n20 2.24063
R21209 VOUT+.n86 VOUT+.n84 2.23934
R21210 VOUT+.n86 VOUT+.n82 2.23934
R21211 VOUT+.n6 VOUT+.n4 1.83719
R21212 VOUT+.n10 VOUT+.n9 1.72967
R21213 VOUT+.n17 VOUT+.n2 1.72967
R21214 VOUT+.n78 VOUT+.n77 1.5005
R21215 VOUT+.n76 VOUT+.n35 1.5005
R21216 VOUT+.n75 VOUT+.n74 1.5005
R21217 VOUT+.n73 VOUT+.n38 1.5005
R21218 VOUT+.n72 VOUT+.n71 1.5005
R21219 VOUT+.n70 VOUT+.n39 1.5005
R21220 VOUT+.n69 VOUT+.n68 1.5005
R21221 VOUT+.n67 VOUT+.n42 1.5005
R21222 VOUT+.n18 VOUT+.n17 1.5005
R21223 VOUT+.n16 VOUT+.n0 1.5005
R21224 VOUT+.n15 VOUT+.n14 1.5005
R21225 VOUT+.n13 VOUT+.n3 1.5005
R21226 VOUT+.n12 VOUT+.n11 1.5005
R21227 VOUT+.n64 VOUT+.n59 1.313
R21228 VOUT+.n55 VOUT+.n41 1.313
R21229 VOUT+.n52 VOUT+.n40 1.313
R21230 VOUT+.n49 VOUT+.n37 1.313
R21231 VOUT+.n45 VOUT+.n43 1.313
R21232 VOUT+.n47 VOUT+.n36 1.313
R21233 VOUT+.n184 VOUT+.n29 1.1455
R21234 VOUT+.n95 VOUT+.n94 1.13717
R21235 VOUT+.n96 VOUT+.n92 1.13717
R21236 VOUT+.n180 VOUT+.n179 1.13717
R21237 VOUT+.n93 VOUT+.n30 1.13717
R21238 VOUT+.n94 VOUT+.n27 1.13717
R21239 VOUT+.n92 VOUT+.n91 1.13717
R21240 VOUT+.n181 VOUT+.n180 1.13717
R21241 VOUT+.n66 VOUT+.n43 0.715216
R21242 VOUT+.n65 VOUT+.n64 0.65675
R21243 VOUT+.n69 VOUT+.n41 0.65675
R21244 VOUT+.n71 VOUT+.n40 0.65675
R21245 VOUT+.n75 VOUT+.n37 0.65675
R21246 VOUT+.n77 VOUT+.n36 0.65675
R21247 VOUT+.n95 VOUT+.n29 0.585
R21248 VOUT+.n67 VOUT+.n66 0.564601
R21249 VOUT+.n61 VOUT+.n60 0.563
R21250 VOUT+.n62 VOUT+.n61 0.563
R21251 VOUT+.n63 VOUT+.n62 0.563
R21252 VOUT+.n57 VOUT+.n56 0.563
R21253 VOUT+.n56 VOUT+.n53 0.563
R21254 VOUT+.n53 VOUT+.n50 0.563
R21255 VOUT+.n189 VOUT+.n185 0.5455
R21256 VOUT+.n87 VOUT+.n78 0.495292
R21257 VOUT+.n136 VOUT+.n135 0.3295
R21258 VOUT+.n137 VOUT+.n136 0.3295
R21259 VOUT+.n138 VOUT+.n137 0.3295
R21260 VOUT+.n139 VOUT+.n138 0.3295
R21261 VOUT+.n140 VOUT+.n139 0.3295
R21262 VOUT+.n141 VOUT+.n140 0.3295
R21263 VOUT+.n142 VOUT+.n141 0.3295
R21264 VOUT+.n143 VOUT+.n142 0.3295
R21265 VOUT+.n144 VOUT+.n143 0.3295
R21266 VOUT+.n145 VOUT+.n144 0.3295
R21267 VOUT+.n147 VOUT+.n145 0.3295
R21268 VOUT+.n147 VOUT+.n146 0.3295
R21269 VOUT+.n150 VOUT+.n148 0.3295
R21270 VOUT+.n150 VOUT+.n149 0.3295
R21271 VOUT+.n153 VOUT+.n151 0.3295
R21272 VOUT+.n153 VOUT+.n152 0.3295
R21273 VOUT+.n156 VOUT+.n154 0.3295
R21274 VOUT+.n156 VOUT+.n155 0.3295
R21275 VOUT+.n159 VOUT+.n157 0.3295
R21276 VOUT+.n159 VOUT+.n158 0.3295
R21277 VOUT+.n162 VOUT+.n160 0.3295
R21278 VOUT+.n162 VOUT+.n161 0.3295
R21279 VOUT+.n165 VOUT+.n163 0.3295
R21280 VOUT+.n165 VOUT+.n164 0.3295
R21281 VOUT+.n168 VOUT+.n166 0.3295
R21282 VOUT+.n168 VOUT+.n167 0.3295
R21283 VOUT+.n171 VOUT+.n169 0.3295
R21284 VOUT+.n171 VOUT+.n170 0.3295
R21285 VOUT+.n174 VOUT+.n172 0.3295
R21286 VOUT+.n174 VOUT+.n173 0.3295
R21287 VOUT+.n98 VOUT+.n97 0.3295
R21288 VOUT+.n100 VOUT+.n99 0.3295
R21289 VOUT+.n101 VOUT+.n100 0.3295
R21290 VOUT+.n102 VOUT+.n101 0.3295
R21291 VOUT+.n103 VOUT+.n102 0.3295
R21292 VOUT+.n104 VOUT+.n103 0.3295
R21293 VOUT+.n105 VOUT+.n104 0.3295
R21294 VOUT+.n106 VOUT+.n105 0.3295
R21295 VOUT+.n107 VOUT+.n106 0.3295
R21296 VOUT+.n108 VOUT+.n107 0.3295
R21297 VOUT+.n109 VOUT+.n108 0.3295
R21298 VOUT+.n111 VOUT+.n109 0.3295
R21299 VOUT+.n111 VOUT+.n110 0.3295
R21300 VOUT+.n114 VOUT+.n112 0.3295
R21301 VOUT+.n114 VOUT+.n113 0.3295
R21302 VOUT+.n117 VOUT+.n115 0.3295
R21303 VOUT+.n117 VOUT+.n116 0.3295
R21304 VOUT+.n120 VOUT+.n118 0.3295
R21305 VOUT+.n120 VOUT+.n119 0.3295
R21306 VOUT+.n123 VOUT+.n121 0.3295
R21307 VOUT+.n123 VOUT+.n122 0.3295
R21308 VOUT+.n126 VOUT+.n124 0.3295
R21309 VOUT+.n126 VOUT+.n125 0.3295
R21310 VOUT+.n129 VOUT+.n127 0.3295
R21311 VOUT+.n129 VOUT+.n128 0.3295
R21312 VOUT+.n132 VOUT+.n130 0.3295
R21313 VOUT+.n132 VOUT+.n131 0.3295
R21314 VOUT+.n177 VOUT+.n176 0.3295
R21315 VOUT+.n176 VOUT+.n175 0.3295
R21316 VOUT+.n12 VOUT+.n4 0.314966
R21317 VOUT+.n178 VOUT+.n177 0.313833
R21318 VOUT+.n143 VOUT+.n133 0.306
R21319 VOUT+.n142 VOUT+.n134 0.306
R21320 VOUT+.n150 VOUT+.n147 0.2825
R21321 VOUT+.n153 VOUT+.n150 0.2825
R21322 VOUT+.n156 VOUT+.n153 0.2825
R21323 VOUT+.n159 VOUT+.n156 0.2825
R21324 VOUT+.n162 VOUT+.n159 0.2825
R21325 VOUT+.n165 VOUT+.n162 0.2825
R21326 VOUT+.n168 VOUT+.n165 0.2825
R21327 VOUT+.n171 VOUT+.n168 0.2825
R21328 VOUT+.n174 VOUT+.n171 0.2825
R21329 VOUT+.n111 VOUT+.n98 0.2825
R21330 VOUT+.n114 VOUT+.n111 0.2825
R21331 VOUT+.n117 VOUT+.n114 0.2825
R21332 VOUT+.n120 VOUT+.n117 0.2825
R21333 VOUT+.n123 VOUT+.n120 0.2825
R21334 VOUT+.n126 VOUT+.n123 0.2825
R21335 VOUT+.n129 VOUT+.n126 0.2825
R21336 VOUT+.n132 VOUT+.n129 0.2825
R21337 VOUT+.n176 VOUT+.n132 0.2825
R21338 VOUT+.n176 VOUT+.n174 0.2825
R21339 VOUT+.n183 VOUT+.n88 0.2455
R21340 VOUT+ VOUT+.n194 0.198417
R21341 VOUT+.n194 VOUT+.n193 0.193208
R21342 VOUT+ VOUT+.n18 0.182792
R21343 VOUT+.n179 VOUT+.n178 0.138367
R21344 VOUT+.n10 VOUT+.n4 0.0891864
R21345 VOUT+.n65 VOUT+.n42 0.0577917
R21346 VOUT+.n69 VOUT+.n42 0.0577917
R21347 VOUT+.n70 VOUT+.n69 0.0577917
R21348 VOUT+.n71 VOUT+.n70 0.0577917
R21349 VOUT+.n71 VOUT+.n38 0.0577917
R21350 VOUT+.n75 VOUT+.n38 0.0577917
R21351 VOUT+.n76 VOUT+.n75 0.0577917
R21352 VOUT+.n77 VOUT+.n76 0.0577917
R21353 VOUT+.n68 VOUT+.n67 0.0577917
R21354 VOUT+.n68 VOUT+.n39 0.0577917
R21355 VOUT+.n72 VOUT+.n39 0.0577917
R21356 VOUT+.n73 VOUT+.n72 0.0577917
R21357 VOUT+.n74 VOUT+.n73 0.0577917
R21358 VOUT+.n74 VOUT+.n35 0.0577917
R21359 VOUT+.n78 VOUT+.n35 0.0577917
R21360 VOUT+.n66 VOUT+.n65 0.054517
R21361 VOUT+.n191 VOUT+.n24 0.047375
R21362 VOUT+.n186 VOUT+.n22 0.047375
R21363 VOUT+.n184 VOUT+.n30 0.0421667
R21364 VOUT+.n87 VOUT+.n81 0.0421667
R21365 VOUT+.n11 VOUT+.n10 0.0421667
R21366 VOUT+.n11 VOUT+.n3 0.0421667
R21367 VOUT+.n15 VOUT+.n3 0.0421667
R21368 VOUT+.n16 VOUT+.n15 0.0421667
R21369 VOUT+.n17 VOUT+.n16 0.0421667
R21370 VOUT+.n13 VOUT+.n12 0.0421667
R21371 VOUT+.n14 VOUT+.n13 0.0421667
R21372 VOUT+.n14 VOUT+.n0 0.0421667
R21373 VOUT+.n18 VOUT+.n0 0.0421667
R21374 VOUT+.n82 VOUT+.n81 0.0243161
R21375 VOUT+.n84 VOUT+.n32 0.0243161
R21376 VOUT+.n84 VOUT+.n83 0.0243161
R21377 VOUT+.n82 VOUT+.n34 0.0243161
R21378 VOUT+.n181 VOUT+.n26 0.0217373
R21379 VOUT+.n83 VOUT+.n33 0.0217373
R21380 VOUT+.n91 VOUT+.n26 0.0217373
R21381 VOUT+.n188 VOUT+.n23 0.0217373
R21382 VOUT+.n186 VOUT+.n23 0.0217373
R21383 VOUT+.n89 VOUT+.n30 0.0217373
R21384 VOUT+.n91 VOUT+.n90 0.0217373
R21385 VOUT+.n79 VOUT+.n32 0.0217373
R21386 VOUT+.n79 VOUT+.n34 0.0217373
R21387 VOUT+.n89 VOUT+.n27 0.0217373
R21388 VOUT+.n90 VOUT+.n27 0.0217373
R21389 VOUT+.n193 VOUT+.n20 0.0217373
R21390 VOUT+.n191 VOUT+.n190 0.0217373
R21391 VOUT+.n190 VOUT+.n22 0.0217373
R21392 VOUT+.n24 VOUT+.n20 0.0217373
R21393 VOUT+.n96 VOUT+.n95 0.0161667
R21394 VOUT+.n179 VOUT+.n96 0.0161667
R21395 VOUT+.n94 VOUT+.n93 0.0161667
R21396 VOUT+.n94 VOUT+.n92 0.0161667
R21397 VOUT+.n180 VOUT+.n92 0.0161667
R21398 VOUT+.n182 VOUT+.n28 0.0134654
R21399 VOUT+.n185 VOUT+.n25 0.0134654
R21400 VOUT+.n183 VOUT+.n182 0.0134654
R21401 VOUT+.n28 VOUT+.n25 0.0134654
R21402 VOUT+.n85 VOUT+.n80 0.0109778
R21403 VOUT+.n88 VOUT+.n31 0.0109778
R21404 VOUT+.n187 VOUT+.n19 0.0109778
R21405 VOUT+.n192 VOUT+.n21 0.0109778
R21406 VOUT+.n86 VOUT+.n85 0.0109778
R21407 VOUT+.n80 VOUT+.n31 0.0109778
R21408 VOUT+.n189 VOUT+.n187 0.0109778
R21409 VOUT+.n21 VOUT+.n19 0.0109778
R21410 VOUT+.n93 VOUT+.n29 0.00872683
R21411 two_stage_opamp_dummy_magic_26_0.cap_res_Y two_stage_opamp_dummy_magic_26_0.cap_res_Y.t138 49.895
R21412 two_stage_opamp_dummy_magic_26_0.cap_res_Y two_stage_opamp_dummy_magic_26_0.cap_res_Y.t70 0.9405
R21413 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t81 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t12 0.1603
R21414 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t40 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t124 0.1603
R21415 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t34 0.1603
R21416 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t130 0.1603
R21417 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t48 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t18 0.1603
R21418 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t120 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t25 0.1603
R21419 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t91 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t52 0.1603
R21420 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t82 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t135 0.1603
R21421 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t24 0.1603
R21422 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t31 0.1603
R21423 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t60 0.1603
R21424 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t22 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t68 0.1603
R21425 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t137 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t98 0.1603
R21426 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t33 0.1603
R21427 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t99 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t66 0.1603
R21428 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t76 0.1603
R21429 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t108 0.1603
R21430 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t118 0.1603
R21431 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t7 0.1603
R21432 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t14 0.1603
R21433 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t41 0.1603
R21434 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t125 0.1603
R21435 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t42 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t11 0.1603
R21436 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t113 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t20 0.1603
R21437 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t87 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t47 0.1603
R21438 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t57 0.1603
R21439 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t133 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t90 0.1603
R21440 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t121 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t26 0.1603
R21441 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t92 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t53 0.1603
R21442 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t109 0.1603
R21443 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t116 0.1603
R21444 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t74 0.1603
R21445 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t2 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t106 0.1603
R21446 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t110 0.1603
R21447 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t1 0.1603
R21448 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t129 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t49 0.1603
R21449 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t89 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t45 0.1603
R21450 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t88 0.1603
R21451 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t64 0.1603
R21452 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t6 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t101 0.1603
R21453 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t3 0.1603
R21454 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t80 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t37 0.1603
R21455 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t19 0.1603
R21456 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t95 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t51 0.1603
R21457 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t94 0.1603
R21458 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t73 0.1603
R21459 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t112 0.1603
R21460 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t85 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t15 0.1603
R21461 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t111 0.1603
R21462 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t105 0.1603
R21463 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t93 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t55 0.1603
R21464 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t43 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t13 0.1603
R21465 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t86 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t46 0.1603
R21466 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t32 0.1603
R21467 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t100 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t67 0.1603
R21468 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t102 0.1603
R21469 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t36 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t5 0.1603
R21470 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t128 0.1603
R21471 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t21 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t50 0.1603
R21472 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t70 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t21 0.1603
R21473 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n16 0.159278
R21474 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n17 0.159278
R21475 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t28 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n18 0.159278
R21476 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t97 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n19 0.159278
R21477 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t123 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n20 0.159278
R21478 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t10 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n21 0.159278
R21479 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n22 0.159278
R21480 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n23 0.159278
R21481 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n24 0.159278
R21482 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t65 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n25 0.159278
R21483 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n26 0.159278
R21484 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n27 0.159278
R21485 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t23 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n28 0.159278
R21486 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n29 0.159278
R21487 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t83 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n30 0.159278
R21488 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t122 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n31 0.159278
R21489 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n32 0.159278
R21490 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n33 0.159278
R21491 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n34 0.159278
R21492 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t81 0.1368
R21493 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t40 0.1368
R21494 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t75 0.1368
R21495 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t77 0.1368
R21496 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t48 0.1368
R21497 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t120 0.1368
R21498 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t91 0.1368
R21499 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t82 0.1368
R21500 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t54 0.1368
R21501 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t126 0.1368
R21502 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t96 0.1368
R21503 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t22 0.1368
R21504 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t137 0.1368
R21505 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t131 0.1368
R21506 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t99 0.1368
R21507 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t29 0.1368
R21508 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t4 0.1368
R21509 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t63 0.1368
R21510 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t39 0.1368
R21511 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t103 0.1368
R21512 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t84 0.1368
R21513 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t71 0.1368
R21514 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t42 0.1368
R21515 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t113 0.1368
R21516 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t87 0.1368
R21517 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t9 0.1368
R21518 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t133 0.1368
R21519 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t121 0.1368
R21520 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t92 0.1368
R21521 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t44 0.1368
R21522 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t61 0.1368
R21523 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t27 0.1368
R21524 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t2 0.1368
R21525 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t58 0.1368
R21526 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t35 0.1368
R21527 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t129 0.1368
R21528 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t85 0.1368
R21529 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n35 0.1368
R21530 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n36 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t69 0.1368
R21531 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t89 0.114322
R21532 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t43 0.114322
R21533 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n6 0.1133
R21534 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n7 0.1133
R21535 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n8 0.1133
R21536 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n9 0.1133
R21537 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n10 0.1133
R21538 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n11 0.1133
R21539 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n12 0.1133
R21540 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n13 0.1133
R21541 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n14 0.1133
R21542 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n15 0.1133
R21543 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n0 0.1133
R21544 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n1 0.1133
R21545 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n2 0.1133
R21546 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n3 0.1133
R21547 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n4 0.1133
R21548 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n37 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n5 0.1133
R21549 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n37 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n36 0.1133
R21550 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t134 0.00152174
R21551 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t104 0.00152174
R21552 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t6 0.00152174
R21553 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t38 0.00152174
R21554 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t80 0.00152174
R21555 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t56 0.00152174
R21556 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t95 0.00152174
R21557 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t136 0.00152174
R21558 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t115 0.00152174
R21559 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t8 0.00152174
R21560 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t119 0.00152174
R21561 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t16 0.00152174
R21562 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t59 0.00152174
R21563 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t28 0.00152174
R21564 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t97 0.00152174
R21565 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t123 0.00152174
R21566 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t10 0.00152174
R21567 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t114 0.00152174
R21568 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t72 0.00152174
R21569 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t107 0.00152174
R21570 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t65 0.00152174
R21571 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t30 0.00152174
R21572 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t132 0.00152174
R21573 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t23 0.00152174
R21574 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t127 0.00152174
R21575 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t83 0.00152174
R21576 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t122 0.00152174
R21577 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t78 0.00152174
R21578 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t79 0.00152174
R21579 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t117 0.00152174
R21580 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n36 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t93 0.00152174
R21581 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t86 0.00152174
R21582 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t62 0.00152174
R21583 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t100 0.00152174
R21584 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t0 0.00152174
R21585 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t36 0.00152174
R21586 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t17 0.00152174
R21587 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n37 0.00152174
R21588 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t26 610.534
R21589 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t24 610.534
R21590 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t15 433.8
R21591 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t12 433.8
R21592 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t21 433.8
R21593 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t29 433.8
R21594 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t18 433.8
R21595 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t28 433.8
R21596 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t17 433.8
R21597 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n34 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t27 433.8
R21598 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n35 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t31 433.8
R21599 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t25 433.8
R21600 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t14 433.8
R21601 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t23 433.8
R21602 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t13 433.8
R21603 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t22 433.8
R21604 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t30 433.8
R21605 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t20 433.8
R21606 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t19 433.8
R21607 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t16 433.8
R21608 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n14 287.264
R21609 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n18 287.264
R21610 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n15 287.264
R21611 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n21 287.264
R21612 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n35 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n34 176.733
R21613 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n34 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n33 176.733
R21614 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n32 176.733
R21615 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n31 176.733
R21616 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n30 176.733
R21617 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n29 176.733
R21618 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n28 176.733
R21619 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n27 176.733
R21620 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n6 176.733
R21621 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n7 176.733
R21622 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n8 176.733
R21623 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n9 176.733
R21624 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n10 176.733
R21625 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n11 176.733
R21626 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n25 176.733
R21627 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n37 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n36 161.986
R21628 two_stage_opamp_dummy_magic_26_0.V_tail_gate two_stage_opamp_dummy_magic_26_0.V_tail_gate.n13 161.986
R21629 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n22 63.1128
R21630 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n0 63.112
R21631 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n2 63.112
R21632 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n2 52.5725
R21633 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n20 52.5725
R21634 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n19 52.01
R21635 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n16 52.01
R21636 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n23 49.7255
R21637 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n4 49.7255
R21638 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_26_0.V_tail_gate 46.7517
R21639 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n36 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n35 45.5227
R21640 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n12 45.5227
R21641 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n13 45.5227
R21642 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n36 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n26 45.5227
R21643 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t7 39.4005
R21644 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t3 39.4005
R21645 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t9 39.4005
R21646 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t6 39.4005
R21647 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t8 39.4005
R21648 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t4 39.4005
R21649 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t5 39.4005
R21650 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t10 39.4005
R21651 two_stage_opamp_dummy_magic_26_0.V_tail_gate two_stage_opamp_dummy_magic_26_0.V_tail_gate.n3 16.3608
R21652 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t2 16.0005
R21653 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t0 16.0005
R21654 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t1 16.0005
R21655 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t11 16.0005
R21656 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n5 9.563
R21657 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n0 6.16966
R21658 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n37 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n24 2.35766
R21659 two_stage_opamp_dummy_magic_26_0.V_tail_gate two_stage_opamp_dummy_magic_26_0.V_tail_gate.n5 2.188
R21660 two_stage_opamp_dummy_magic_26_0.V_tail_gate two_stage_opamp_dummy_magic_26_0.V_tail_gate.n1 1.73143
R21661 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n37 1.44719
R21662 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n17 0.563
R21663 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n0 0.34059
R21664 two_stage_opamp_dummy_magic_26_0.V_source.n60 two_stage_opamp_dummy_magic_26_0.V_source.t35 67.42
R21665 two_stage_opamp_dummy_magic_26_0.V_source.n28 two_stage_opamp_dummy_magic_26_0.V_source.n27 49.3505
R21666 two_stage_opamp_dummy_magic_26_0.V_source.n26 two_stage_opamp_dummy_magic_26_0.V_source.n25 49.3505
R21667 two_stage_opamp_dummy_magic_26_0.V_source.n16 two_stage_opamp_dummy_magic_26_0.V_source.n15 49.3505
R21668 two_stage_opamp_dummy_magic_26_0.V_source.n34 two_stage_opamp_dummy_magic_26_0.V_source.n33 49.3505
R21669 two_stage_opamp_dummy_magic_26_0.V_source.n31 two_stage_opamp_dummy_magic_26_0.V_source.n30 49.3505
R21670 two_stage_opamp_dummy_magic_26_0.V_source.n43 two_stage_opamp_dummy_magic_26_0.V_source.n42 49.3505
R21671 two_stage_opamp_dummy_magic_26_0.V_source.n39 two_stage_opamp_dummy_magic_26_0.V_source.n38 49.3505
R21672 two_stage_opamp_dummy_magic_26_0.V_source.n37 two_stage_opamp_dummy_magic_26_0.V_source.n36 49.3505
R21673 two_stage_opamp_dummy_magic_26_0.V_source.n22 two_stage_opamp_dummy_magic_26_0.V_source.n21 49.3505
R21674 two_stage_opamp_dummy_magic_26_0.V_source.n18 two_stage_opamp_dummy_magic_26_0.V_source.n17 49.3505
R21675 two_stage_opamp_dummy_magic_26_0.V_source.n47 two_stage_opamp_dummy_magic_26_0.V_source.n46 32.3838
R21676 two_stage_opamp_dummy_magic_26_0.V_source.n49 two_stage_opamp_dummy_magic_26_0.V_source.n48 32.3838
R21677 two_stage_opamp_dummy_magic_26_0.V_source.n6 two_stage_opamp_dummy_magic_26_0.V_source.n5 32.3838
R21678 two_stage_opamp_dummy_magic_26_0.V_source.n54 two_stage_opamp_dummy_magic_26_0.V_source.n53 32.3838
R21679 two_stage_opamp_dummy_magic_26_0.V_source.n57 two_stage_opamp_dummy_magic_26_0.V_source.n56 32.3838
R21680 two_stage_opamp_dummy_magic_26_0.V_source.n9 two_stage_opamp_dummy_magic_26_0.V_source.n8 32.3838
R21681 two_stage_opamp_dummy_magic_26_0.V_source.n71 two_stage_opamp_dummy_magic_26_0.V_source.n70 32.3838
R21682 two_stage_opamp_dummy_magic_26_0.V_source.n74 two_stage_opamp_dummy_magic_26_0.V_source.n73 32.3838
R21683 two_stage_opamp_dummy_magic_26_0.V_source.n78 two_stage_opamp_dummy_magic_26_0.V_source.n77 32.3838
R21684 two_stage_opamp_dummy_magic_26_0.V_source.n68 two_stage_opamp_dummy_magic_26_0.V_source.n67 32.3838
R21685 two_stage_opamp_dummy_magic_26_0.V_source.n27 two_stage_opamp_dummy_magic_26_0.V_source.t5 16.0005
R21686 two_stage_opamp_dummy_magic_26_0.V_source.n27 two_stage_opamp_dummy_magic_26_0.V_source.t28 16.0005
R21687 two_stage_opamp_dummy_magic_26_0.V_source.n25 two_stage_opamp_dummy_magic_26_0.V_source.t6 16.0005
R21688 two_stage_opamp_dummy_magic_26_0.V_source.n25 two_stage_opamp_dummy_magic_26_0.V_source.t40 16.0005
R21689 two_stage_opamp_dummy_magic_26_0.V_source.n15 two_stage_opamp_dummy_magic_26_0.V_source.t38 16.0005
R21690 two_stage_opamp_dummy_magic_26_0.V_source.n15 two_stage_opamp_dummy_magic_26_0.V_source.t27 16.0005
R21691 two_stage_opamp_dummy_magic_26_0.V_source.n33 two_stage_opamp_dummy_magic_26_0.V_source.t0 16.0005
R21692 two_stage_opamp_dummy_magic_26_0.V_source.n33 two_stage_opamp_dummy_magic_26_0.V_source.t2 16.0005
R21693 two_stage_opamp_dummy_magic_26_0.V_source.n30 two_stage_opamp_dummy_magic_26_0.V_source.t33 16.0005
R21694 two_stage_opamp_dummy_magic_26_0.V_source.n30 two_stage_opamp_dummy_magic_26_0.V_source.t32 16.0005
R21695 two_stage_opamp_dummy_magic_26_0.V_source.n42 two_stage_opamp_dummy_magic_26_0.V_source.t1 16.0005
R21696 two_stage_opamp_dummy_magic_26_0.V_source.n42 two_stage_opamp_dummy_magic_26_0.V_source.t36 16.0005
R21697 two_stage_opamp_dummy_magic_26_0.V_source.n38 two_stage_opamp_dummy_magic_26_0.V_source.t3 16.0005
R21698 two_stage_opamp_dummy_magic_26_0.V_source.n38 two_stage_opamp_dummy_magic_26_0.V_source.t39 16.0005
R21699 two_stage_opamp_dummy_magic_26_0.V_source.n36 two_stage_opamp_dummy_magic_26_0.V_source.t34 16.0005
R21700 two_stage_opamp_dummy_magic_26_0.V_source.n36 two_stage_opamp_dummy_magic_26_0.V_source.t8 16.0005
R21701 two_stage_opamp_dummy_magic_26_0.V_source.n21 two_stage_opamp_dummy_magic_26_0.V_source.t30 16.0005
R21702 two_stage_opamp_dummy_magic_26_0.V_source.n21 two_stage_opamp_dummy_magic_26_0.V_source.t37 16.0005
R21703 two_stage_opamp_dummy_magic_26_0.V_source.n17 two_stage_opamp_dummy_magic_26_0.V_source.t29 16.0005
R21704 two_stage_opamp_dummy_magic_26_0.V_source.n17 two_stage_opamp_dummy_magic_26_0.V_source.t4 16.0005
R21705 two_stage_opamp_dummy_magic_26_0.V_source.n46 two_stage_opamp_dummy_magic_26_0.V_source.t22 9.6005
R21706 two_stage_opamp_dummy_magic_26_0.V_source.n46 two_stage_opamp_dummy_magic_26_0.V_source.t12 9.6005
R21707 two_stage_opamp_dummy_magic_26_0.V_source.n48 two_stage_opamp_dummy_magic_26_0.V_source.t21 9.6005
R21708 two_stage_opamp_dummy_magic_26_0.V_source.n48 two_stage_opamp_dummy_magic_26_0.V_source.t11 9.6005
R21709 two_stage_opamp_dummy_magic_26_0.V_source.n5 two_stage_opamp_dummy_magic_26_0.V_source.t7 9.6005
R21710 two_stage_opamp_dummy_magic_26_0.V_source.n5 two_stage_opamp_dummy_magic_26_0.V_source.t31 9.6005
R21711 two_stage_opamp_dummy_magic_26_0.V_source.n53 two_stage_opamp_dummy_magic_26_0.V_source.t10 9.6005
R21712 two_stage_opamp_dummy_magic_26_0.V_source.n53 two_stage_opamp_dummy_magic_26_0.V_source.t17 9.6005
R21713 two_stage_opamp_dummy_magic_26_0.V_source.n56 two_stage_opamp_dummy_magic_26_0.V_source.t15 9.6005
R21714 two_stage_opamp_dummy_magic_26_0.V_source.n56 two_stage_opamp_dummy_magic_26_0.V_source.t19 9.6005
R21715 two_stage_opamp_dummy_magic_26_0.V_source.n8 two_stage_opamp_dummy_magic_26_0.V_source.t25 9.6005
R21716 two_stage_opamp_dummy_magic_26_0.V_source.n8 two_stage_opamp_dummy_magic_26_0.V_source.t16 9.6005
R21717 two_stage_opamp_dummy_magic_26_0.V_source.n70 two_stage_opamp_dummy_magic_26_0.V_source.t9 9.6005
R21718 two_stage_opamp_dummy_magic_26_0.V_source.n70 two_stage_opamp_dummy_magic_26_0.V_source.t13 9.6005
R21719 two_stage_opamp_dummy_magic_26_0.V_source.n73 two_stage_opamp_dummy_magic_26_0.V_source.t23 9.6005
R21720 two_stage_opamp_dummy_magic_26_0.V_source.n73 two_stage_opamp_dummy_magic_26_0.V_source.t20 9.6005
R21721 two_stage_opamp_dummy_magic_26_0.V_source.n77 two_stage_opamp_dummy_magic_26_0.V_source.t24 9.6005
R21722 two_stage_opamp_dummy_magic_26_0.V_source.n77 two_stage_opamp_dummy_magic_26_0.V_source.t14 9.6005
R21723 two_stage_opamp_dummy_magic_26_0.V_source.n67 two_stage_opamp_dummy_magic_26_0.V_source.t18 9.6005
R21724 two_stage_opamp_dummy_magic_26_0.V_source.n67 two_stage_opamp_dummy_magic_26_0.V_source.t26 9.6005
R21725 two_stage_opamp_dummy_magic_26_0.V_source.n80 two_stage_opamp_dummy_magic_26_0.V_source.n6 5.85227
R21726 two_stage_opamp_dummy_magic_26_0.V_source.n37 two_stage_opamp_dummy_magic_26_0.V_source.n13 5.51092
R21727 two_stage_opamp_dummy_magic_26_0.V_source.n19 two_stage_opamp_dummy_magic_26_0.V_source.n16 5.51092
R21728 two_stage_opamp_dummy_magic_26_0.V_source.n40 two_stage_opamp_dummy_magic_26_0.V_source.n37 5.45883
R21729 two_stage_opamp_dummy_magic_26_0.V_source.n16 two_stage_opamp_dummy_magic_26_0.V_source.n14 5.45883
R21730 two_stage_opamp_dummy_magic_26_0.V_source.n71 two_stage_opamp_dummy_magic_26_0.V_source.n69 5.188
R21731 two_stage_opamp_dummy_magic_26_0.V_source.n74 two_stage_opamp_dummy_magic_26_0.V_source.n7 5.188
R21732 two_stage_opamp_dummy_magic_26_0.V_source.n79 two_stage_opamp_dummy_magic_26_0.V_source.n78 5.188
R21733 two_stage_opamp_dummy_magic_26_0.V_source.n44 two_stage_opamp_dummy_magic_26_0.V_source.n43 5.16717
R21734 two_stage_opamp_dummy_magic_26_0.V_source.n39 two_stage_opamp_dummy_magic_26_0.V_source.n13 5.16717
R21735 two_stage_opamp_dummy_magic_26_0.V_source.n22 two_stage_opamp_dummy_magic_26_0.V_source.n20 5.16717
R21736 two_stage_opamp_dummy_magic_26_0.V_source.n19 two_stage_opamp_dummy_magic_26_0.V_source.n18 5.16717
R21737 two_stage_opamp_dummy_magic_26_0.V_source.n35 two_stage_opamp_dummy_magic_26_0.V_source.n34 4.89633
R21738 two_stage_opamp_dummy_magic_26_0.V_source.n43 two_stage_opamp_dummy_magic_26_0.V_source.n41 4.89633
R21739 two_stage_opamp_dummy_magic_26_0.V_source.n40 two_stage_opamp_dummy_magic_26_0.V_source.n39 4.89633
R21740 two_stage_opamp_dummy_magic_26_0.V_source.n29 two_stage_opamp_dummy_magic_26_0.V_source.n28 4.89633
R21741 two_stage_opamp_dummy_magic_26_0.V_source.n32 two_stage_opamp_dummy_magic_26_0.V_source.n31 4.89633
R21742 two_stage_opamp_dummy_magic_26_0.V_source.n23 two_stage_opamp_dummy_magic_26_0.V_source.n22 4.89633
R21743 two_stage_opamp_dummy_magic_26_0.V_source.n18 two_stage_opamp_dummy_magic_26_0.V_source.n14 4.89633
R21744 two_stage_opamp_dummy_magic_26_0.V_source.n26 two_stage_opamp_dummy_magic_26_0.V_source.n24 4.89633
R21745 two_stage_opamp_dummy_magic_26_0.V_source.n61 two_stage_opamp_dummy_magic_26_0.V_source.n51 4.5005
R21746 two_stage_opamp_dummy_magic_26_0.V_source.n63 two_stage_opamp_dummy_magic_26_0.V_source.n62 4.5005
R21747 two_stage_opamp_dummy_magic_26_0.V_source.n62 two_stage_opamp_dummy_magic_26_0.V_source.n61 4.5005
R21748 two_stage_opamp_dummy_magic_26_0.V_source.n32 two_stage_opamp_dummy_magic_26_0.V_source.n29 3.6255
R21749 two_stage_opamp_dummy_magic_26_0.V_source.n47 two_stage_opamp_dummy_magic_26_0.V_source.n11 2.44497
R21750 two_stage_opamp_dummy_magic_26_0.V_source.n50 two_stage_opamp_dummy_magic_26_0.V_source.n49 2.44497
R21751 two_stage_opamp_dummy_magic_26_0.V_source.n55 two_stage_opamp_dummy_magic_26_0.V_source.n54 2.44497
R21752 two_stage_opamp_dummy_magic_26_0.V_source.n58 two_stage_opamp_dummy_magic_26_0.V_source.n57 2.44497
R21753 two_stage_opamp_dummy_magic_26_0.V_source.n10 two_stage_opamp_dummy_magic_26_0.V_source.n9 2.44497
R21754 two_stage_opamp_dummy_magic_26_0.V_source.n72 two_stage_opamp_dummy_magic_26_0.V_source.n71 2.44497
R21755 two_stage_opamp_dummy_magic_26_0.V_source.n75 two_stage_opamp_dummy_magic_26_0.V_source.n74 2.44497
R21756 two_stage_opamp_dummy_magic_26_0.V_source.n78 two_stage_opamp_dummy_magic_26_0.V_source.n76 2.44497
R21757 two_stage_opamp_dummy_magic_26_0.V_source.n59 two_stage_opamp_dummy_magic_26_0.V_source.n6 2.44497
R21758 two_stage_opamp_dummy_magic_26_0.V_source.n68 two_stage_opamp_dummy_magic_26_0.V_source.n66 2.44462
R21759 two_stage_opamp_dummy_magic_26_0.V_source.n64 two_stage_opamp_dummy_magic_26_0.V_source.n63 2.24063
R21760 two_stage_opamp_dummy_magic_26_0.V_source.n52 two_stage_opamp_dummy_magic_26_0.V_source.n0 2.24063
R21761 two_stage_opamp_dummy_magic_26_0.V_source.n65 two_stage_opamp_dummy_magic_26_0.V_source.n0 2.24063
R21762 two_stage_opamp_dummy_magic_26_0.V_source.n45 two_stage_opamp_dummy_magic_26_0.V_source.n12 2.2076
R21763 two_stage_opamp_dummy_magic_26_0.V_source.n1 two_stage_opamp_dummy_magic_26_0.V_source.n45 2.16822
R21764 two_stage_opamp_dummy_magic_26_0.V_source.n12 two_stage_opamp_dummy_magic_26_0.V_source.n3 2.16822
R21765 two_stage_opamp_dummy_magic_26_0.V_source.n69 two_stage_opamp_dummy_magic_26_0.V_source.n2 2.02255
R21766 two_stage_opamp_dummy_magic_26_0.V_source.n4 two_stage_opamp_dummy_magic_26_0.V_source.n80 1.36007
R21767 two_stage_opamp_dummy_magic_26_0.V_source.n61 two_stage_opamp_dummy_magic_26_0.V_source.n60 0.922375
R21768 two_stage_opamp_dummy_magic_26_0.V_source.n60 two_stage_opamp_dummy_magic_26_0.V_source.n59 2.64916
R21769 two_stage_opamp_dummy_magic_26_0.V_source.n80 two_stage_opamp_dummy_magic_26_0.V_source.n79 0.664374
R21770 two_stage_opamp_dummy_magic_26_0.V_source.n2 two_stage_opamp_dummy_magic_26_0.V_source.n47 0.6255
R21771 two_stage_opamp_dummy_magic_26_0.V_source.n2 two_stage_opamp_dummy_magic_26_0.V_source.n49 0.6255
R21772 two_stage_opamp_dummy_magic_26_0.V_source.n9 two_stage_opamp_dummy_magic_26_0.V_source.n4 0.6255
R21773 two_stage_opamp_dummy_magic_26_0.V_source.n57 two_stage_opamp_dummy_magic_26_0.V_source.n4 0.6255
R21774 two_stage_opamp_dummy_magic_26_0.V_source.n54 two_stage_opamp_dummy_magic_26_0.V_source.n4 0.6255
R21775 two_stage_opamp_dummy_magic_26_0.V_source.n2 two_stage_opamp_dummy_magic_26_0.V_source.n68 0.6255
R21776 two_stage_opamp_dummy_magic_26_0.V_source.n31 two_stage_opamp_dummy_magic_26_0.V_source.n1 0.604667
R21777 two_stage_opamp_dummy_magic_26_0.V_source.n34 two_stage_opamp_dummy_magic_26_0.V_source.n1 0.604667
R21778 two_stage_opamp_dummy_magic_26_0.V_source.n3 two_stage_opamp_dummy_magic_26_0.V_source.n26 0.604667
R21779 two_stage_opamp_dummy_magic_26_0.V_source.n28 two_stage_opamp_dummy_magic_26_0.V_source.n3 0.604667
R21780 two_stage_opamp_dummy_magic_26_0.V_source.n41 two_stage_opamp_dummy_magic_26_0.V_source.n40 0.563
R21781 two_stage_opamp_dummy_magic_26_0.V_source.n41 two_stage_opamp_dummy_magic_26_0.V_source.n35 0.563
R21782 two_stage_opamp_dummy_magic_26_0.V_source.n35 two_stage_opamp_dummy_magic_26_0.V_source.n32 0.563
R21783 two_stage_opamp_dummy_magic_26_0.V_source.n29 two_stage_opamp_dummy_magic_26_0.V_source.n24 0.563
R21784 two_stage_opamp_dummy_magic_26_0.V_source.n23 two_stage_opamp_dummy_magic_26_0.V_source.n14 0.563
R21785 two_stage_opamp_dummy_magic_26_0.V_source.n24 two_stage_opamp_dummy_magic_26_0.V_source.n23 0.563
R21786 two_stage_opamp_dummy_magic_26_0.V_source.n20 two_stage_opamp_dummy_magic_26_0.V_source.n12 0.510302
R21787 two_stage_opamp_dummy_magic_26_0.V_source.n45 two_stage_opamp_dummy_magic_26_0.V_source.n44 0.510302
R21788 two_stage_opamp_dummy_magic_26_0.V_source.n2 two_stage_opamp_dummy_magic_26_0.V_source.n1 0.450019
R21789 two_stage_opamp_dummy_magic_26_0.V_source two_stage_opamp_dummy_magic_26_0.V_source.n3 0.353865
R21790 two_stage_opamp_dummy_magic_26_0.V_source.n20 two_stage_opamp_dummy_magic_26_0.V_source.n19 0.34425
R21791 two_stage_opamp_dummy_magic_26_0.V_source.n44 two_stage_opamp_dummy_magic_26_0.V_source.n13 0.34425
R21792 two_stage_opamp_dummy_magic_26_0.V_source.n79 two_stage_opamp_dummy_magic_26_0.V_source.n7 0.34425
R21793 two_stage_opamp_dummy_magic_26_0.V_source.n69 two_stage_opamp_dummy_magic_26_0.V_source.n7 0.34425
R21794 two_stage_opamp_dummy_magic_26_0.V_source.n66 two_stage_opamp_dummy_magic_26_0.V_source.n65 1.63868
R21795 two_stage_opamp_dummy_magic_26_0.V_source.n59 two_stage_opamp_dummy_magic_26_0.V_source.n58 0.115083
R21796 two_stage_opamp_dummy_magic_26_0.V_source.n58 two_stage_opamp_dummy_magic_26_0.V_source.n55 0.115083
R21797 two_stage_opamp_dummy_magic_26_0.V_source.n55 two_stage_opamp_dummy_magic_26_0.V_source.n10 0.115083
R21798 two_stage_opamp_dummy_magic_26_0.V_source.n76 two_stage_opamp_dummy_magic_26_0.V_source.n10 0.115083
R21799 two_stage_opamp_dummy_magic_26_0.V_source.n76 two_stage_opamp_dummy_magic_26_0.V_source.n75 0.115083
R21800 two_stage_opamp_dummy_magic_26_0.V_source.n75 two_stage_opamp_dummy_magic_26_0.V_source.n72 0.115083
R21801 two_stage_opamp_dummy_magic_26_0.V_source.n72 two_stage_opamp_dummy_magic_26_0.V_source.n11 0.115083
R21802 two_stage_opamp_dummy_magic_26_0.V_source.n50 two_stage_opamp_dummy_magic_26_0.V_source.n11 0.115083
R21803 two_stage_opamp_dummy_magic_26_0.V_source.n66 two_stage_opamp_dummy_magic_26_0.V_source.n50 0.115083
R21804 two_stage_opamp_dummy_magic_26_0.V_source two_stage_opamp_dummy_magic_26_0.V_source.n4 0.0966538
R21805 two_stage_opamp_dummy_magic_26_0.V_source.n63 two_stage_opamp_dummy_magic_26_0.V_source.n0 0.0421667
R21806 two_stage_opamp_dummy_magic_26_0.V_source.n65 two_stage_opamp_dummy_magic_26_0.V_source.n64 0.0217373
R21807 two_stage_opamp_dummy_magic_26_0.V_source.n62 two_stage_opamp_dummy_magic_26_0.V_source.n52 0.0217373
R21808 two_stage_opamp_dummy_magic_26_0.V_source.n64 two_stage_opamp_dummy_magic_26_0.V_source.n51 0.0217373
R21809 two_stage_opamp_dummy_magic_26_0.V_source.n52 two_stage_opamp_dummy_magic_26_0.V_source.n51 0.0217373
R21810 two_stage_opamp_dummy_magic_26_0.V_source.n61 two_stage_opamp_dummy_magic_26_0.V_source.n0 0.0429746
R21811 two_stage_opamp_dummy_magic_26_0.Y.n68 two_stage_opamp_dummy_magic_26_0.Y.t38 1172.87
R21812 two_stage_opamp_dummy_magic_26_0.Y.n64 two_stage_opamp_dummy_magic_26_0.Y.t28 1172.87
R21813 two_stage_opamp_dummy_magic_26_0.Y.n68 two_stage_opamp_dummy_magic_26_0.Y.t29 996.134
R21814 two_stage_opamp_dummy_magic_26_0.Y.n69 two_stage_opamp_dummy_magic_26_0.Y.t45 996.134
R21815 two_stage_opamp_dummy_magic_26_0.Y.n70 two_stage_opamp_dummy_magic_26_0.Y.t32 996.134
R21816 two_stage_opamp_dummy_magic_26_0.Y.n71 two_stage_opamp_dummy_magic_26_0.Y.t48 996.134
R21817 two_stage_opamp_dummy_magic_26_0.Y.n67 two_stage_opamp_dummy_magic_26_0.Y.t35 996.134
R21818 two_stage_opamp_dummy_magic_26_0.Y.n66 two_stage_opamp_dummy_magic_26_0.Y.t41 996.134
R21819 two_stage_opamp_dummy_magic_26_0.Y.n65 two_stage_opamp_dummy_magic_26_0.Y.t25 996.134
R21820 two_stage_opamp_dummy_magic_26_0.Y.n64 two_stage_opamp_dummy_magic_26_0.Y.t43 996.134
R21821 two_stage_opamp_dummy_magic_26_0.Y.n86 two_stage_opamp_dummy_magic_26_0.Y.t53 690.867
R21822 two_stage_opamp_dummy_magic_26_0.Y.n79 two_stage_opamp_dummy_magic_26_0.Y.t49 690.867
R21823 two_stage_opamp_dummy_magic_26_0.Y.n95 two_stage_opamp_dummy_magic_26_0.Y.t36 530.201
R21824 two_stage_opamp_dummy_magic_26_0.Y.n88 two_stage_opamp_dummy_magic_26_0.Y.t26 530.201
R21825 two_stage_opamp_dummy_magic_26_0.Y.n86 two_stage_opamp_dummy_magic_26_0.Y.t50 514.134
R21826 two_stage_opamp_dummy_magic_26_0.Y.n79 two_stage_opamp_dummy_magic_26_0.Y.t33 514.134
R21827 two_stage_opamp_dummy_magic_26_0.Y.n80 two_stage_opamp_dummy_magic_26_0.Y.t46 514.134
R21828 two_stage_opamp_dummy_magic_26_0.Y.n81 two_stage_opamp_dummy_magic_26_0.Y.t30 514.134
R21829 two_stage_opamp_dummy_magic_26_0.Y.n82 two_stage_opamp_dummy_magic_26_0.Y.t52 514.134
R21830 two_stage_opamp_dummy_magic_26_0.Y.n83 two_stage_opamp_dummy_magic_26_0.Y.t39 514.134
R21831 two_stage_opamp_dummy_magic_26_0.Y.n84 two_stage_opamp_dummy_magic_26_0.Y.t51 514.134
R21832 two_stage_opamp_dummy_magic_26_0.Y.n85 two_stage_opamp_dummy_magic_26_0.Y.t37 514.134
R21833 two_stage_opamp_dummy_magic_26_0.Y.n95 two_stage_opamp_dummy_magic_26_0.Y.t27 353.467
R21834 two_stage_opamp_dummy_magic_26_0.Y.n94 two_stage_opamp_dummy_magic_26_0.Y.t44 353.467
R21835 two_stage_opamp_dummy_magic_26_0.Y.n93 two_stage_opamp_dummy_magic_26_0.Y.t31 353.467
R21836 two_stage_opamp_dummy_magic_26_0.Y.n92 two_stage_opamp_dummy_magic_26_0.Y.t47 353.467
R21837 two_stage_opamp_dummy_magic_26_0.Y.n91 two_stage_opamp_dummy_magic_26_0.Y.t34 353.467
R21838 two_stage_opamp_dummy_magic_26_0.Y.n90 two_stage_opamp_dummy_magic_26_0.Y.t40 353.467
R21839 two_stage_opamp_dummy_magic_26_0.Y.n89 two_stage_opamp_dummy_magic_26_0.Y.t54 353.467
R21840 two_stage_opamp_dummy_magic_26_0.Y.n88 two_stage_opamp_dummy_magic_26_0.Y.t42 353.467
R21841 two_stage_opamp_dummy_magic_26_0.Y.n67 two_stage_opamp_dummy_magic_26_0.Y.n66 176.733
R21842 two_stage_opamp_dummy_magic_26_0.Y.n66 two_stage_opamp_dummy_magic_26_0.Y.n65 176.733
R21843 two_stage_opamp_dummy_magic_26_0.Y.n65 two_stage_opamp_dummy_magic_26_0.Y.n64 176.733
R21844 two_stage_opamp_dummy_magic_26_0.Y.n69 two_stage_opamp_dummy_magic_26_0.Y.n68 176.733
R21845 two_stage_opamp_dummy_magic_26_0.Y.n70 two_stage_opamp_dummy_magic_26_0.Y.n69 176.733
R21846 two_stage_opamp_dummy_magic_26_0.Y.n71 two_stage_opamp_dummy_magic_26_0.Y.n70 176.733
R21847 two_stage_opamp_dummy_magic_26_0.Y.n94 two_stage_opamp_dummy_magic_26_0.Y.n93 176.733
R21848 two_stage_opamp_dummy_magic_26_0.Y.n93 two_stage_opamp_dummy_magic_26_0.Y.n92 176.733
R21849 two_stage_opamp_dummy_magic_26_0.Y.n92 two_stage_opamp_dummy_magic_26_0.Y.n91 176.733
R21850 two_stage_opamp_dummy_magic_26_0.Y.n91 two_stage_opamp_dummy_magic_26_0.Y.n90 176.733
R21851 two_stage_opamp_dummy_magic_26_0.Y.n90 two_stage_opamp_dummy_magic_26_0.Y.n89 176.733
R21852 two_stage_opamp_dummy_magic_26_0.Y.n89 two_stage_opamp_dummy_magic_26_0.Y.n88 176.733
R21853 two_stage_opamp_dummy_magic_26_0.Y.n85 two_stage_opamp_dummy_magic_26_0.Y.n84 176.733
R21854 two_stage_opamp_dummy_magic_26_0.Y.n84 two_stage_opamp_dummy_magic_26_0.Y.n83 176.733
R21855 two_stage_opamp_dummy_magic_26_0.Y.n83 two_stage_opamp_dummy_magic_26_0.Y.n82 176.733
R21856 two_stage_opamp_dummy_magic_26_0.Y.n82 two_stage_opamp_dummy_magic_26_0.Y.n81 176.733
R21857 two_stage_opamp_dummy_magic_26_0.Y.n81 two_stage_opamp_dummy_magic_26_0.Y.n80 176.733
R21858 two_stage_opamp_dummy_magic_26_0.Y.n80 two_stage_opamp_dummy_magic_26_0.Y.n79 176.733
R21859 two_stage_opamp_dummy_magic_26_0.Y.n97 two_stage_opamp_dummy_magic_26_0.Y.n96 165.472
R21860 two_stage_opamp_dummy_magic_26_0.Y.n97 two_stage_opamp_dummy_magic_26_0.Y.n87 165.472
R21861 two_stage_opamp_dummy_magic_26_0.Y.n74 two_stage_opamp_dummy_magic_26_0.Y.n73 152
R21862 two_stage_opamp_dummy_magic_26_0.Y.n75 two_stage_opamp_dummy_magic_26_0.Y.n74 131.571
R21863 two_stage_opamp_dummy_magic_26_0.Y.n74 two_stage_opamp_dummy_magic_26_0.Y.n72 124.517
R21864 two_stage_opamp_dummy_magic_26_0.Y.n105 two_stage_opamp_dummy_magic_26_0.Y.n97 73.6876
R21865 two_stage_opamp_dummy_magic_26_0.Y.n47 two_stage_opamp_dummy_magic_26_0.Y.n46 66.0338
R21866 two_stage_opamp_dummy_magic_26_0.Y.n31 two_stage_opamp_dummy_magic_26_0.Y.n30 66.0338
R21867 two_stage_opamp_dummy_magic_26_0.Y.n34 two_stage_opamp_dummy_magic_26_0.Y.n33 66.0338
R21868 two_stage_opamp_dummy_magic_26_0.Y.n37 two_stage_opamp_dummy_magic_26_0.Y.n36 66.0338
R21869 two_stage_opamp_dummy_magic_26_0.Y.n41 two_stage_opamp_dummy_magic_26_0.Y.n40 66.0338
R21870 two_stage_opamp_dummy_magic_26_0.Y.n44 two_stage_opamp_dummy_magic_26_0.Y.n43 66.0338
R21871 two_stage_opamp_dummy_magic_26_0.Y.n8 two_stage_opamp_dummy_magic_26_0.Y.n6 54.7984
R21872 two_stage_opamp_dummy_magic_26_0.Y.n8 two_stage_opamp_dummy_magic_26_0.Y.n7 54.4547
R21873 two_stage_opamp_dummy_magic_26_0.Y.n10 two_stage_opamp_dummy_magic_26_0.Y.n9 54.4547
R21874 two_stage_opamp_dummy_magic_26_0.Y.n12 two_stage_opamp_dummy_magic_26_0.Y.n11 54.4547
R21875 two_stage_opamp_dummy_magic_26_0.Y.n14 two_stage_opamp_dummy_magic_26_0.Y.n13 54.4547
R21876 two_stage_opamp_dummy_magic_26_0.Y.n16 two_stage_opamp_dummy_magic_26_0.Y.n15 54.4547
R21877 two_stage_opamp_dummy_magic_26_0.Y.n58 two_stage_opamp_dummy_magic_26_0.Y.t24 41.0384
R21878 two_stage_opamp_dummy_magic_26_0.Y.n72 two_stage_opamp_dummy_magic_26_0.Y.n67 40.1672
R21879 two_stage_opamp_dummy_magic_26_0.Y.n72 two_stage_opamp_dummy_magic_26_0.Y.n71 40.1672
R21880 two_stage_opamp_dummy_magic_26_0.Y.n96 two_stage_opamp_dummy_magic_26_0.Y.n94 40.1672
R21881 two_stage_opamp_dummy_magic_26_0.Y.n96 two_stage_opamp_dummy_magic_26_0.Y.n95 40.1672
R21882 two_stage_opamp_dummy_magic_26_0.Y.n87 two_stage_opamp_dummy_magic_26_0.Y.n85 40.1672
R21883 two_stage_opamp_dummy_magic_26_0.Y.n87 two_stage_opamp_dummy_magic_26_0.Y.n86 40.1672
R21884 two_stage_opamp_dummy_magic_26_0.Y.n76 two_stage_opamp_dummy_magic_26_0.Y.n75 16.3217
R21885 two_stage_opamp_dummy_magic_26_0.Y.n6 two_stage_opamp_dummy_magic_26_0.Y.t20 16.0005
R21886 two_stage_opamp_dummy_magic_26_0.Y.n6 two_stage_opamp_dummy_magic_26_0.Y.t3 16.0005
R21887 two_stage_opamp_dummy_magic_26_0.Y.n7 two_stage_opamp_dummy_magic_26_0.Y.t17 16.0005
R21888 two_stage_opamp_dummy_magic_26_0.Y.n7 two_stage_opamp_dummy_magic_26_0.Y.t14 16.0005
R21889 two_stage_opamp_dummy_magic_26_0.Y.n9 two_stage_opamp_dummy_magic_26_0.Y.t15 16.0005
R21890 two_stage_opamp_dummy_magic_26_0.Y.n9 two_stage_opamp_dummy_magic_26_0.Y.t18 16.0005
R21891 two_stage_opamp_dummy_magic_26_0.Y.n11 two_stage_opamp_dummy_magic_26_0.Y.t16 16.0005
R21892 two_stage_opamp_dummy_magic_26_0.Y.n11 two_stage_opamp_dummy_magic_26_0.Y.t11 16.0005
R21893 two_stage_opamp_dummy_magic_26_0.Y.n13 two_stage_opamp_dummy_magic_26_0.Y.t12 16.0005
R21894 two_stage_opamp_dummy_magic_26_0.Y.n13 two_stage_opamp_dummy_magic_26_0.Y.t19 16.0005
R21895 two_stage_opamp_dummy_magic_26_0.Y.n15 two_stage_opamp_dummy_magic_26_0.Y.t2 16.0005
R21896 two_stage_opamp_dummy_magic_26_0.Y.n15 two_stage_opamp_dummy_magic_26_0.Y.t13 16.0005
R21897 two_stage_opamp_dummy_magic_26_0.Y.n73 two_stage_opamp_dummy_magic_26_0.Y.n63 12.8005
R21898 two_stage_opamp_dummy_magic_26_0.Y.n46 two_stage_opamp_dummy_magic_26_0.Y.t6 11.2576
R21899 two_stage_opamp_dummy_magic_26_0.Y.n46 two_stage_opamp_dummy_magic_26_0.Y.t9 11.2576
R21900 two_stage_opamp_dummy_magic_26_0.Y.n30 two_stage_opamp_dummy_magic_26_0.Y.t10 11.2576
R21901 two_stage_opamp_dummy_magic_26_0.Y.n30 two_stage_opamp_dummy_magic_26_0.Y.t22 11.2576
R21902 two_stage_opamp_dummy_magic_26_0.Y.n33 two_stage_opamp_dummy_magic_26_0.Y.t23 11.2576
R21903 two_stage_opamp_dummy_magic_26_0.Y.n33 two_stage_opamp_dummy_magic_26_0.Y.t5 11.2576
R21904 two_stage_opamp_dummy_magic_26_0.Y.n36 two_stage_opamp_dummy_magic_26_0.Y.t4 11.2576
R21905 two_stage_opamp_dummy_magic_26_0.Y.n36 two_stage_opamp_dummy_magic_26_0.Y.t1 11.2576
R21906 two_stage_opamp_dummy_magic_26_0.Y.n40 two_stage_opamp_dummy_magic_26_0.Y.t21 11.2576
R21907 two_stage_opamp_dummy_magic_26_0.Y.n40 two_stage_opamp_dummy_magic_26_0.Y.t0 11.2576
R21908 two_stage_opamp_dummy_magic_26_0.Y.n43 two_stage_opamp_dummy_magic_26_0.Y.t7 11.2576
R21909 two_stage_opamp_dummy_magic_26_0.Y.n43 two_stage_opamp_dummy_magic_26_0.Y.t8 11.2576
R21910 two_stage_opamp_dummy_magic_26_0.Y.n17 two_stage_opamp_dummy_magic_26_0.Y.n16 10.9224
R21911 two_stage_opamp_dummy_magic_26_0.Y.n73 two_stage_opamp_dummy_magic_26_0.Y.n61 9.36264
R21912 two_stage_opamp_dummy_magic_26_0.Y.n63 two_stage_opamp_dummy_magic_26_0.Y.n62 9.3005
R21913 two_stage_opamp_dummy_magic_26_0.Y.n118 two_stage_opamp_dummy_magic_26_0.Y.n25 6.1255
R21914 two_stage_opamp_dummy_magic_26_0.Y.n18 two_stage_opamp_dummy_magic_26_0.Y.n17 5.84022
R21915 two_stage_opamp_dummy_magic_26_0.Y.n19 two_stage_opamp_dummy_magic_26_0.Y.n5 5.78175
R21916 two_stage_opamp_dummy_magic_26_0.Y.n21 two_stage_opamp_dummy_magic_26_0.Y.n4 5.78175
R21917 two_stage_opamp_dummy_magic_26_0.Y.n124 two_stage_opamp_dummy_magic_26_0.Y.n1 5.78175
R21918 two_stage_opamp_dummy_magic_26_0.Y.n120 two_stage_opamp_dummy_magic_26_0.Y.n25 5.78175
R21919 two_stage_opamp_dummy_magic_26_0.Y.n35 two_stage_opamp_dummy_magic_26_0.Y.n31 5.66717
R21920 two_stage_opamp_dummy_magic_26_0.Y.n32 two_stage_opamp_dummy_magic_26_0.Y.n31 5.66717
R21921 two_stage_opamp_dummy_magic_26_0.Y.n47 two_stage_opamp_dummy_magic_26_0.Y.n45 5.66717
R21922 two_stage_opamp_dummy_magic_26_0.Y.n75 two_stage_opamp_dummy_magic_26_0.Y.n63 5.33141
R21923 two_stage_opamp_dummy_magic_26_0.Y.n35 two_stage_opamp_dummy_magic_26_0.Y.n34 5.29217
R21924 two_stage_opamp_dummy_magic_26_0.Y.n34 two_stage_opamp_dummy_magic_26_0.Y.n32 5.29217
R21925 two_stage_opamp_dummy_magic_26_0.Y.n38 two_stage_opamp_dummy_magic_26_0.Y.n37 5.29217
R21926 two_stage_opamp_dummy_magic_26_0.Y.n37 two_stage_opamp_dummy_magic_26_0.Y.n29 5.29217
R21927 two_stage_opamp_dummy_magic_26_0.Y.n41 two_stage_opamp_dummy_magic_26_0.Y.n39 5.29217
R21928 two_stage_opamp_dummy_magic_26_0.Y.n42 two_stage_opamp_dummy_magic_26_0.Y.n41 5.29217
R21929 two_stage_opamp_dummy_magic_26_0.Y.n44 two_stage_opamp_dummy_magic_26_0.Y.n28 5.29217
R21930 two_stage_opamp_dummy_magic_26_0.Y.n45 two_stage_opamp_dummy_magic_26_0.Y.n44 5.29217
R21931 two_stage_opamp_dummy_magic_26_0.Y.n48 two_stage_opamp_dummy_magic_26_0.Y.n47 5.29217
R21932 two_stage_opamp_dummy_magic_26_0.Y.n49 two_stage_opamp_dummy_magic_26_0.Y.n27 4.5005
R21933 two_stage_opamp_dummy_magic_26_0.Y.n100 two_stage_opamp_dummy_magic_26_0.Y.n99 4.5005
R21934 two_stage_opamp_dummy_magic_26_0.Y.n106 two_stage_opamp_dummy_magic_26_0.Y.n51 4.5005
R21935 two_stage_opamp_dummy_magic_26_0.Y.n108 two_stage_opamp_dummy_magic_26_0.Y.n107 4.5005
R21936 two_stage_opamp_dummy_magic_26_0.Y.n107 two_stage_opamp_dummy_magic_26_0.Y.n106 4.5005
R21937 two_stage_opamp_dummy_magic_26_0.Y.n77 two_stage_opamp_dummy_magic_26_0.Y.n76 4.5005
R21938 two_stage_opamp_dummy_magic_26_0.Y.n55 two_stage_opamp_dummy_magic_26_0.Y.n54 4.5005
R21939 two_stage_opamp_dummy_magic_26_0.Y.n114 two_stage_opamp_dummy_magic_26_0.Y.n48 2.35543
R21940 two_stage_opamp_dummy_magic_26_0.Y.n101 two_stage_opamp_dummy_magic_26_0.Y.n98 2.26187
R21941 two_stage_opamp_dummy_magic_26_0.Y.n102 two_stage_opamp_dummy_magic_26_0.Y.n101 2.26187
R21942 two_stage_opamp_dummy_magic_26_0.Y.n56 two_stage_opamp_dummy_magic_26_0.Y.n53 2.26187
R21943 two_stage_opamp_dummy_magic_26_0.Y.n103 two_stage_opamp_dummy_magic_26_0.Y.n102 2.26187
R21944 two_stage_opamp_dummy_magic_26_0.Y.n113 two_stage_opamp_dummy_magic_26_0.Y.n112 2.26187
R21945 two_stage_opamp_dummy_magic_26_0.Y.n57 two_stage_opamp_dummy_magic_26_0.Y.n56 2.26187
R21946 two_stage_opamp_dummy_magic_26_0.Y.n116 two_stage_opamp_dummy_magic_26_0.Y.n26 2.24063
R21947 two_stage_opamp_dummy_magic_26_0.Y.n112 two_stage_opamp_dummy_magic_26_0.Y.n111 2.24063
R21948 two_stage_opamp_dummy_magic_26_0.Y.n109 two_stage_opamp_dummy_magic_26_0.Y.n108 2.24063
R21949 two_stage_opamp_dummy_magic_26_0.Y.n78 two_stage_opamp_dummy_magic_26_0.Y.n52 2.24063
R21950 two_stage_opamp_dummy_magic_26_0.Y.n60 two_stage_opamp_dummy_magic_26_0.Y.n53 2.24063
R21951 two_stage_opamp_dummy_magic_26_0.Y.n115 two_stage_opamp_dummy_magic_26_0.Y.n114 2.24063
R21952 two_stage_opamp_dummy_magic_26_0.Y.n104 two_stage_opamp_dummy_magic_26_0.Y.n98 2.24063
R21953 two_stage_opamp_dummy_magic_26_0.Y.n110 two_stage_opamp_dummy_magic_26_0.Y.n50 2.24063
R21954 two_stage_opamp_dummy_magic_26_0.Y.n59 two_stage_opamp_dummy_magic_26_0.Y.n58 2.24063
R21955 two_stage_opamp_dummy_magic_26_0.Y.n77 two_stage_opamp_dummy_magic_26_0.Y.n61 2.22018
R21956 two_stage_opamp_dummy_magic_26_0.Y.n118 two_stage_opamp_dummy_magic_26_0.Y.n117 1.5005
R21957 two_stage_opamp_dummy_magic_26_0.Y.n119 two_stage_opamp_dummy_magic_26_0.Y.n24 1.5005
R21958 two_stage_opamp_dummy_magic_26_0.Y.n121 two_stage_opamp_dummy_magic_26_0.Y.n120 1.5005
R21959 two_stage_opamp_dummy_magic_26_0.Y.n122 two_stage_opamp_dummy_magic_26_0.Y.n2 1.5005
R21960 two_stage_opamp_dummy_magic_26_0.Y.n124 two_stage_opamp_dummy_magic_26_0.Y.n123 1.5005
R21961 two_stage_opamp_dummy_magic_26_0.Y.n23 two_stage_opamp_dummy_magic_26_0.Y.n0 1.5005
R21962 two_stage_opamp_dummy_magic_26_0.Y.n22 two_stage_opamp_dummy_magic_26_0.Y.n21 1.5005
R21963 two_stage_opamp_dummy_magic_26_0.Y.n20 two_stage_opamp_dummy_magic_26_0.Y.n3 1.5005
R21964 two_stage_opamp_dummy_magic_26_0.Y.n107 two_stage_opamp_dummy_magic_26_0.Y.n105 0.850077
R21965 two_stage_opamp_dummy_magic_26_0.Y.n77 two_stage_opamp_dummy_magic_26_0.Y.n60 0.682792
R21966 two_stage_opamp_dummy_magic_26_0.Y.n111 two_stage_opamp_dummy_magic_26_0.Y.n110 0.646333
R21967 two_stage_opamp_dummy_magic_26_0.Y.n117 two_stage_opamp_dummy_magic_26_0.Y.n116 0.630708
R21968 two_stage_opamp_dummy_magic_26_0.Y.n18 two_stage_opamp_dummy_magic_26_0.Y.n3 0.564601
R21969 two_stage_opamp_dummy_magic_26_0.Y.n108 two_stage_opamp_dummy_magic_26_0.Y.n77 0.46925
R21970 two_stage_opamp_dummy_magic_26_0.Y.n105 two_stage_opamp_dummy_magic_26_0.Y.n104 0.376306
R21971 two_stage_opamp_dummy_magic_26_0.Y.n45 two_stage_opamp_dummy_magic_26_0.Y.n42 0.3755
R21972 two_stage_opamp_dummy_magic_26_0.Y.n42 two_stage_opamp_dummy_magic_26_0.Y.n29 0.3755
R21973 two_stage_opamp_dummy_magic_26_0.Y.n32 two_stage_opamp_dummy_magic_26_0.Y.n29 0.3755
R21974 two_stage_opamp_dummy_magic_26_0.Y.n48 two_stage_opamp_dummy_magic_26_0.Y.n28 0.3755
R21975 two_stage_opamp_dummy_magic_26_0.Y.n39 two_stage_opamp_dummy_magic_26_0.Y.n28 0.3755
R21976 two_stage_opamp_dummy_magic_26_0.Y.n39 two_stage_opamp_dummy_magic_26_0.Y.n38 0.3755
R21977 two_stage_opamp_dummy_magic_26_0.Y.n38 two_stage_opamp_dummy_magic_26_0.Y.n35 0.3755
R21978 two_stage_opamp_dummy_magic_26_0.Y.n16 two_stage_opamp_dummy_magic_26_0.Y.n14 0.34425
R21979 two_stage_opamp_dummy_magic_26_0.Y.n14 two_stage_opamp_dummy_magic_26_0.Y.n12 0.34425
R21980 two_stage_opamp_dummy_magic_26_0.Y.n12 two_stage_opamp_dummy_magic_26_0.Y.n10 0.34425
R21981 two_stage_opamp_dummy_magic_26_0.Y.n10 two_stage_opamp_dummy_magic_26_0.Y.n8 0.34425
R21982 two_stage_opamp_dummy_magic_26_0.Y.n17 two_stage_opamp_dummy_magic_26_0.Y.n5 0.34425
R21983 two_stage_opamp_dummy_magic_26_0.Y.n5 two_stage_opamp_dummy_magic_26_0.Y.n4 0.34425
R21984 two_stage_opamp_dummy_magic_26_0.Y.n4 two_stage_opamp_dummy_magic_26_0.Y.n1 0.34425
R21985 two_stage_opamp_dummy_magic_26_0.Y.n25 two_stage_opamp_dummy_magic_26_0.Y.n1 0.34425
R21986 two_stage_opamp_dummy_magic_26_0.Y.n76 two_stage_opamp_dummy_magic_26_0.Y.n62 0.1255
R21987 two_stage_opamp_dummy_magic_26_0.Y.n62 two_stage_opamp_dummy_magic_26_0.Y.n61 0.0626438
R21988 two_stage_opamp_dummy_magic_26_0.Y.n20 two_stage_opamp_dummy_magic_26_0.Y.n19 0.0577917
R21989 two_stage_opamp_dummy_magic_26_0.Y.n21 two_stage_opamp_dummy_magic_26_0.Y.n20 0.0577917
R21990 two_stage_opamp_dummy_magic_26_0.Y.n21 two_stage_opamp_dummy_magic_26_0.Y.n0 0.0577917
R21991 two_stage_opamp_dummy_magic_26_0.Y.n124 two_stage_opamp_dummy_magic_26_0.Y.n2 0.0577917
R21992 two_stage_opamp_dummy_magic_26_0.Y.n120 two_stage_opamp_dummy_magic_26_0.Y.n2 0.0577917
R21993 two_stage_opamp_dummy_magic_26_0.Y.n120 two_stage_opamp_dummy_magic_26_0.Y.n119 0.0577917
R21994 two_stage_opamp_dummy_magic_26_0.Y.n119 two_stage_opamp_dummy_magic_26_0.Y.n118 0.0577917
R21995 two_stage_opamp_dummy_magic_26_0.Y.n22 two_stage_opamp_dummy_magic_26_0.Y.n3 0.0577917
R21996 two_stage_opamp_dummy_magic_26_0.Y.n23 two_stage_opamp_dummy_magic_26_0.Y.n22 0.0577917
R21997 two_stage_opamp_dummy_magic_26_0.Y.n123 two_stage_opamp_dummy_magic_26_0.Y.n23 0.0577917
R21998 two_stage_opamp_dummy_magic_26_0.Y.n123 two_stage_opamp_dummy_magic_26_0.Y.n122 0.0577917
R21999 two_stage_opamp_dummy_magic_26_0.Y.n122 two_stage_opamp_dummy_magic_26_0.Y.n121 0.0577917
R22000 two_stage_opamp_dummy_magic_26_0.Y.n121 two_stage_opamp_dummy_magic_26_0.Y.n24 0.0577917
R22001 two_stage_opamp_dummy_magic_26_0.Y.n117 two_stage_opamp_dummy_magic_26_0.Y.n24 0.0577917
R22002 two_stage_opamp_dummy_magic_26_0.Y.n19 two_stage_opamp_dummy_magic_26_0.Y.n18 0.054517
R22003 two_stage_opamp_dummy_magic_26_0.Y.n108 two_stage_opamp_dummy_magic_26_0.Y.n52 0.0421667
R22004 two_stage_opamp_dummy_magic_26_0.Y two_stage_opamp_dummy_magic_26_0.Y.n0 0.0369583
R22005 two_stage_opamp_dummy_magic_26_0.Y.n49 two_stage_opamp_dummy_magic_26_0.Y.n26 0.0217373
R22006 two_stage_opamp_dummy_magic_26_0.Y.n110 two_stage_opamp_dummy_magic_26_0.Y.n109 0.0217373
R22007 two_stage_opamp_dummy_magic_26_0.Y.n107 two_stage_opamp_dummy_magic_26_0.Y.n78 0.0217373
R22008 two_stage_opamp_dummy_magic_26_0.Y.n101 two_stage_opamp_dummy_magic_26_0.Y.n99 0.0217373
R22009 two_stage_opamp_dummy_magic_26_0.Y.n112 two_stage_opamp_dummy_magic_26_0.Y.n27 0.0217373
R22010 two_stage_opamp_dummy_magic_26_0.Y.n111 two_stage_opamp_dummy_magic_26_0.Y.n26 0.0217373
R22011 two_stage_opamp_dummy_magic_26_0.Y.n102 two_stage_opamp_dummy_magic_26_0.Y.n100 0.0217373
R22012 two_stage_opamp_dummy_magic_26_0.Y.n109 two_stage_opamp_dummy_magic_26_0.Y.n51 0.0217373
R22013 two_stage_opamp_dummy_magic_26_0.Y.n78 two_stage_opamp_dummy_magic_26_0.Y.n51 0.0217373
R22014 two_stage_opamp_dummy_magic_26_0.Y.n55 two_stage_opamp_dummy_magic_26_0.Y.n53 0.0217373
R22015 two_stage_opamp_dummy_magic_26_0.Y.n56 two_stage_opamp_dummy_magic_26_0.Y.n54 0.0217373
R22016 two_stage_opamp_dummy_magic_26_0.Y.n100 two_stage_opamp_dummy_magic_26_0.Y.n98 0.0217373
R22017 two_stage_opamp_dummy_magic_26_0.Y.n115 two_stage_opamp_dummy_magic_26_0.Y.n27 0.0217373
R22018 two_stage_opamp_dummy_magic_26_0.Y.n113 two_stage_opamp_dummy_magic_26_0.Y.n49 0.0217373
R22019 two_stage_opamp_dummy_magic_26_0.Y.n103 two_stage_opamp_dummy_magic_26_0.Y.n99 0.0217373
R22020 two_stage_opamp_dummy_magic_26_0.Y.n114 two_stage_opamp_dummy_magic_26_0.Y.n113 0.0217373
R22021 two_stage_opamp_dummy_magic_26_0.Y.n116 two_stage_opamp_dummy_magic_26_0.Y.n115 0.0217373
R22022 two_stage_opamp_dummy_magic_26_0.Y.n104 two_stage_opamp_dummy_magic_26_0.Y.n103 0.0217373
R22023 two_stage_opamp_dummy_magic_26_0.Y.n106 two_stage_opamp_dummy_magic_26_0.Y.n50 0.0217373
R22024 two_stage_opamp_dummy_magic_26_0.Y.n59 two_stage_opamp_dummy_magic_26_0.Y.n54 0.0217373
R22025 two_stage_opamp_dummy_magic_26_0.Y.n52 two_stage_opamp_dummy_magic_26_0.Y.n50 0.0217373
R22026 two_stage_opamp_dummy_magic_26_0.Y.n57 two_stage_opamp_dummy_magic_26_0.Y.n55 0.0217373
R22027 two_stage_opamp_dummy_magic_26_0.Y.n58 two_stage_opamp_dummy_magic_26_0.Y.n57 0.0217373
R22028 two_stage_opamp_dummy_magic_26_0.Y.n60 two_stage_opamp_dummy_magic_26_0.Y.n59 0.0217373
R22029 two_stage_opamp_dummy_magic_26_0.Y two_stage_opamp_dummy_magic_26_0.Y.n124 0.0213333
R22030 two_stage_opamp_dummy_magic_26_0.Vb2.n2 two_stage_opamp_dummy_magic_26_0.Vb2.t26 752.515
R22031 two_stage_opamp_dummy_magic_26_0.Vb2.n0 two_stage_opamp_dummy_magic_26_0.Vb2.t19 752.515
R22032 two_stage_opamp_dummy_magic_26_0.Vb2.n4 two_stage_opamp_dummy_magic_26_0.Vb2.t15 752.234
R22033 two_stage_opamp_dummy_magic_26_0.Vb2.n4 two_stage_opamp_dummy_magic_26_0.Vb2.t31 752.234
R22034 two_stage_opamp_dummy_magic_26_0.Vb2.n3 two_stage_opamp_dummy_magic_26_0.Vb2.t25 752.234
R22035 two_stage_opamp_dummy_magic_26_0.Vb2.n3 two_stage_opamp_dummy_magic_26_0.Vb2.t29 752.234
R22036 two_stage_opamp_dummy_magic_26_0.Vb2.n3 two_stage_opamp_dummy_magic_26_0.Vb2.t24 752.234
R22037 two_stage_opamp_dummy_magic_26_0.Vb2.n3 two_stage_opamp_dummy_magic_26_0.Vb2.t22 752.234
R22038 two_stage_opamp_dummy_magic_26_0.Vb2.n2 two_stage_opamp_dummy_magic_26_0.Vb2.t14 752.234
R22039 two_stage_opamp_dummy_magic_26_0.Vb2.n2 two_stage_opamp_dummy_magic_26_0.Vb2.t30 752.234
R22040 two_stage_opamp_dummy_magic_26_0.Vb2.n2 two_stage_opamp_dummy_magic_26_0.Vb2.t11 752.234
R22041 two_stage_opamp_dummy_magic_26_0.Vb2.n5 two_stage_opamp_dummy_magic_26_0.Vb2.t13 752.234
R22042 two_stage_opamp_dummy_magic_26_0.Vb2.n5 two_stage_opamp_dummy_magic_26_0.Vb2.t32 752.234
R22043 two_stage_opamp_dummy_magic_26_0.Vb2.n1 two_stage_opamp_dummy_magic_26_0.Vb2.t16 752.234
R22044 two_stage_opamp_dummy_magic_26_0.Vb2.n1 two_stage_opamp_dummy_magic_26_0.Vb2.t18 752.234
R22045 two_stage_opamp_dummy_magic_26_0.Vb2.n1 two_stage_opamp_dummy_magic_26_0.Vb2.t21 752.234
R22046 two_stage_opamp_dummy_magic_26_0.Vb2.n1 two_stage_opamp_dummy_magic_26_0.Vb2.t23 752.234
R22047 two_stage_opamp_dummy_magic_26_0.Vb2.n0 two_stage_opamp_dummy_magic_26_0.Vb2.t27 752.234
R22048 two_stage_opamp_dummy_magic_26_0.Vb2.n0 two_stage_opamp_dummy_magic_26_0.Vb2.t12 752.234
R22049 two_stage_opamp_dummy_magic_26_0.Vb2.n0 two_stage_opamp_dummy_magic_26_0.Vb2.t17 752.234
R22050 two_stage_opamp_dummy_magic_26_0.Vb2.n14 two_stage_opamp_dummy_magic_26_0.Vb2.t20 746.673
R22051 two_stage_opamp_dummy_magic_26_0.Vb2.n17 two_stage_opamp_dummy_magic_26_0.Vb2.t0 745.726
R22052 two_stage_opamp_dummy_magic_26_0.Vb2.n15 two_stage_opamp_dummy_magic_26_0.Vb2.t28 587.551
R22053 two_stage_opamp_dummy_magic_26_0.Vb2.n8 two_stage_opamp_dummy_magic_26_0.Vb2.n6 140.546
R22054 two_stage_opamp_dummy_magic_26_0.Vb2.n12 two_stage_opamp_dummy_magic_26_0.Vb2.n11 139.297
R22055 two_stage_opamp_dummy_magic_26_0.Vb2.n10 two_stage_opamp_dummy_magic_26_0.Vb2.n9 139.297
R22056 two_stage_opamp_dummy_magic_26_0.Vb2.n8 two_stage_opamp_dummy_magic_26_0.Vb2.n7 139.297
R22057 two_stage_opamp_dummy_magic_26_0.Vb2.n13 two_stage_opamp_dummy_magic_26_0.Vb2.n12 82.6203
R22058 two_stage_opamp_dummy_magic_26_0.Vb2.n18 two_stage_opamp_dummy_magic_26_0.Vb2.n17 67.0547
R22059 two_stage_opamp_dummy_magic_26_0.Vb2.n11 two_stage_opamp_dummy_magic_26_0.Vb2.t4 24.0005
R22060 two_stage_opamp_dummy_magic_26_0.Vb2.n11 two_stage_opamp_dummy_magic_26_0.Vb2.t10 24.0005
R22061 two_stage_opamp_dummy_magic_26_0.Vb2.n9 two_stage_opamp_dummy_magic_26_0.Vb2.t7 24.0005
R22062 two_stage_opamp_dummy_magic_26_0.Vb2.n9 two_stage_opamp_dummy_magic_26_0.Vb2.t6 24.0005
R22063 two_stage_opamp_dummy_magic_26_0.Vb2.n7 two_stage_opamp_dummy_magic_26_0.Vb2.t9 24.0005
R22064 two_stage_opamp_dummy_magic_26_0.Vb2.n7 two_stage_opamp_dummy_magic_26_0.Vb2.t8 24.0005
R22065 two_stage_opamp_dummy_magic_26_0.Vb2.n6 two_stage_opamp_dummy_magic_26_0.Vb2.t2 24.0005
R22066 two_stage_opamp_dummy_magic_26_0.Vb2.n6 two_stage_opamp_dummy_magic_26_0.Vb2.t3 24.0005
R22067 two_stage_opamp_dummy_magic_26_0.Vb2.n16 two_stage_opamp_dummy_magic_26_0.Vb2.n4 17.6411
R22068 two_stage_opamp_dummy_magic_26_0.Vb2.n13 two_stage_opamp_dummy_magic_26_0.Vb2.n5 15.9693
R22069 two_stage_opamp_dummy_magic_26_0.Vb2.t1 two_stage_opamp_dummy_magic_26_0.Vb2.n18 11.2576
R22070 two_stage_opamp_dummy_magic_26_0.Vb2.n18 two_stage_opamp_dummy_magic_26_0.Vb2.t5 11.2576
R22071 two_stage_opamp_dummy_magic_26_0.Vb2.n15 two_stage_opamp_dummy_magic_26_0.Vb2.n14 7.06925
R22072 two_stage_opamp_dummy_magic_26_0.Vb2.n10 two_stage_opamp_dummy_magic_26_0.Vb2.n8 6.21925
R22073 two_stage_opamp_dummy_magic_26_0.Vb2.n17 two_stage_opamp_dummy_magic_26_0.Vb2.n16 4.5005
R22074 two_stage_opamp_dummy_magic_26_0.Vb2.n16 two_stage_opamp_dummy_magic_26_0.Vb2.n15 2.85988
R22075 two_stage_opamp_dummy_magic_26_0.Vb2.n14 two_stage_opamp_dummy_magic_26_0.Vb2.n13 1.838
R22076 two_stage_opamp_dummy_magic_26_0.Vb2.n12 two_stage_opamp_dummy_magic_26_0.Vb2.n10 1.2505
R22077 two_stage_opamp_dummy_magic_26_0.Vb2.n3 two_stage_opamp_dummy_magic_26_0.Vb2.n2 1.1255
R22078 two_stage_opamp_dummy_magic_26_0.Vb2.n4 two_stage_opamp_dummy_magic_26_0.Vb2.n3 1.1255
R22079 two_stage_opamp_dummy_magic_26_0.Vb2.n1 two_stage_opamp_dummy_magic_26_0.Vb2.n0 1.1255
R22080 two_stage_opamp_dummy_magic_26_0.Vb2.n5 two_stage_opamp_dummy_magic_26_0.Vb2.n1 1.1255
R22081 two_stage_opamp_dummy_magic_26_0.VD4.n18 two_stage_opamp_dummy_magic_26_0.VD4.t24 671.418
R22082 two_stage_opamp_dummy_magic_26_0.VD4.n15 two_stage_opamp_dummy_magic_26_0.VD4.t27 671.418
R22083 two_stage_opamp_dummy_magic_26_0.VD4.t28 two_stage_opamp_dummy_magic_26_0.VD4.n16 213.131
R22084 two_stage_opamp_dummy_magic_26_0.VD4.n17 two_stage_opamp_dummy_magic_26_0.VD4.t25 213.131
R22085 two_stage_opamp_dummy_magic_26_0.VD4.t14 two_stage_opamp_dummy_magic_26_0.VD4.t28 146.155
R22086 two_stage_opamp_dummy_magic_26_0.VD4.t0 two_stage_opamp_dummy_magic_26_0.VD4.t14 146.155
R22087 two_stage_opamp_dummy_magic_26_0.VD4.t8 two_stage_opamp_dummy_magic_26_0.VD4.t0 146.155
R22088 two_stage_opamp_dummy_magic_26_0.VD4.t4 two_stage_opamp_dummy_magic_26_0.VD4.t8 146.155
R22089 two_stage_opamp_dummy_magic_26_0.VD4.t10 two_stage_opamp_dummy_magic_26_0.VD4.t4 146.155
R22090 two_stage_opamp_dummy_magic_26_0.VD4.t12 two_stage_opamp_dummy_magic_26_0.VD4.t10 146.155
R22091 two_stage_opamp_dummy_magic_26_0.VD4.t16 two_stage_opamp_dummy_magic_26_0.VD4.t12 146.155
R22092 two_stage_opamp_dummy_magic_26_0.VD4.t2 two_stage_opamp_dummy_magic_26_0.VD4.t16 146.155
R22093 two_stage_opamp_dummy_magic_26_0.VD4.t18 two_stage_opamp_dummy_magic_26_0.VD4.t2 146.155
R22094 two_stage_opamp_dummy_magic_26_0.VD4.t6 two_stage_opamp_dummy_magic_26_0.VD4.t18 146.155
R22095 two_stage_opamp_dummy_magic_26_0.VD4.t25 two_stage_opamp_dummy_magic_26_0.VD4.t6 146.155
R22096 two_stage_opamp_dummy_magic_26_0.VD4.n16 two_stage_opamp_dummy_magic_26_0.VD4.t29 76.2576
R22097 two_stage_opamp_dummy_magic_26_0.VD4.n17 two_stage_opamp_dummy_magic_26_0.VD4.t26 76.2576
R22098 two_stage_opamp_dummy_magic_26_0.VD4.n33 two_stage_opamp_dummy_magic_26_0.VD4.n4 67.013
R22099 two_stage_opamp_dummy_magic_26_0.VD4.n32 two_stage_opamp_dummy_magic_26_0.VD4.n7 67.013
R22100 two_stage_opamp_dummy_magic_26_0.VD4.n31 two_stage_opamp_dummy_magic_26_0.VD4.n10 67.013
R22101 two_stage_opamp_dummy_magic_26_0.VD4.n14 two_stage_opamp_dummy_magic_26_0.VD4.n13 67.013
R22102 two_stage_opamp_dummy_magic_26_0.VD4.n0 two_stage_opamp_dummy_magic_26_0.VD4.n29 67.013
R22103 two_stage_opamp_dummy_magic_26_0.VD4.n25 two_stage_opamp_dummy_magic_26_0.VD4.n24 66.0338
R22104 two_stage_opamp_dummy_magic_26_0.VD4.n12 two_stage_opamp_dummy_magic_26_0.VD4.n11 66.0338
R22105 two_stage_opamp_dummy_magic_26_0.VD4.n9 two_stage_opamp_dummy_magic_26_0.VD4.n8 66.0338
R22106 two_stage_opamp_dummy_magic_26_0.VD4.n6 two_stage_opamp_dummy_magic_26_0.VD4.n5 66.0338
R22107 two_stage_opamp_dummy_magic_26_0.VD4.n20 two_stage_opamp_dummy_magic_26_0.VD4.n19 66.0338
R22108 two_stage_opamp_dummy_magic_26_0.VD4.n28 two_stage_opamp_dummy_magic_26_0.VD4.n27 66.0338
R22109 two_stage_opamp_dummy_magic_26_0.VD4.n4 two_stage_opamp_dummy_magic_26_0.VD4.t15 11.2576
R22110 two_stage_opamp_dummy_magic_26_0.VD4.n4 two_stage_opamp_dummy_magic_26_0.VD4.t1 11.2576
R22111 two_stage_opamp_dummy_magic_26_0.VD4.n7 two_stage_opamp_dummy_magic_26_0.VD4.t9 11.2576
R22112 two_stage_opamp_dummy_magic_26_0.VD4.n7 two_stage_opamp_dummy_magic_26_0.VD4.t5 11.2576
R22113 two_stage_opamp_dummy_magic_26_0.VD4.n10 two_stage_opamp_dummy_magic_26_0.VD4.t11 11.2576
R22114 two_stage_opamp_dummy_magic_26_0.VD4.n10 two_stage_opamp_dummy_magic_26_0.VD4.t13 11.2576
R22115 two_stage_opamp_dummy_magic_26_0.VD4.n24 two_stage_opamp_dummy_magic_26_0.VD4.t36 11.2576
R22116 two_stage_opamp_dummy_magic_26_0.VD4.n24 two_stage_opamp_dummy_magic_26_0.VD4.t37 11.2576
R22117 two_stage_opamp_dummy_magic_26_0.VD4.n11 two_stage_opamp_dummy_magic_26_0.VD4.t23 11.2576
R22118 two_stage_opamp_dummy_magic_26_0.VD4.n11 two_stage_opamp_dummy_magic_26_0.VD4.t32 11.2576
R22119 two_stage_opamp_dummy_magic_26_0.VD4.n8 two_stage_opamp_dummy_magic_26_0.VD4.t33 11.2576
R22120 two_stage_opamp_dummy_magic_26_0.VD4.n8 two_stage_opamp_dummy_magic_26_0.VD4.t20 11.2576
R22121 two_stage_opamp_dummy_magic_26_0.VD4.n5 two_stage_opamp_dummy_magic_26_0.VD4.t31 11.2576
R22122 two_stage_opamp_dummy_magic_26_0.VD4.n5 two_stage_opamp_dummy_magic_26_0.VD4.t22 11.2576
R22123 two_stage_opamp_dummy_magic_26_0.VD4.n19 two_stage_opamp_dummy_magic_26_0.VD4.t35 11.2576
R22124 two_stage_opamp_dummy_magic_26_0.VD4.n19 two_stage_opamp_dummy_magic_26_0.VD4.t30 11.2576
R22125 two_stage_opamp_dummy_magic_26_0.VD4.n27 two_stage_opamp_dummy_magic_26_0.VD4.t21 11.2576
R22126 two_stage_opamp_dummy_magic_26_0.VD4.n27 two_stage_opamp_dummy_magic_26_0.VD4.t34 11.2576
R22127 two_stage_opamp_dummy_magic_26_0.VD4.n13 two_stage_opamp_dummy_magic_26_0.VD4.t17 11.2576
R22128 two_stage_opamp_dummy_magic_26_0.VD4.n13 two_stage_opamp_dummy_magic_26_0.VD4.t3 11.2576
R22129 two_stage_opamp_dummy_magic_26_0.VD4.n29 two_stage_opamp_dummy_magic_26_0.VD4.t19 11.2576
R22130 two_stage_opamp_dummy_magic_26_0.VD4.n29 two_stage_opamp_dummy_magic_26_0.VD4.t7 11.2576
R22131 two_stage_opamp_dummy_magic_26_0.VD4.n21 two_stage_opamp_dummy_magic_26_0.VD4.n20 5.66717
R22132 two_stage_opamp_dummy_magic_26_0.VD4.n28 two_stage_opamp_dummy_magic_26_0.VD4.n26 5.66717
R22133 two_stage_opamp_dummy_magic_26_0.VD4.n23 two_stage_opamp_dummy_magic_26_0.VD4.n12 5.29217
R22134 two_stage_opamp_dummy_magic_26_0.VD4.n22 two_stage_opamp_dummy_magic_26_0.VD4.n9 5.29217
R22135 two_stage_opamp_dummy_magic_26_0.VD4.n21 two_stage_opamp_dummy_magic_26_0.VD4.n6 5.29217
R22136 two_stage_opamp_dummy_magic_26_0.VD4.n26 two_stage_opamp_dummy_magic_26_0.VD4.n25 5.29217
R22137 two_stage_opamp_dummy_magic_26_0.VD4.n16 two_stage_opamp_dummy_magic_26_0.VD4.n15 1.90883
R22138 two_stage_opamp_dummy_magic_26_0.VD4.n18 two_stage_opamp_dummy_magic_26_0.VD4.n17 1.90883
R22139 two_stage_opamp_dummy_magic_26_0.VD4.n31 two_stage_opamp_dummy_magic_26_0.VD4.n12 1.02133
R22140 two_stage_opamp_dummy_magic_26_0.VD4.n32 two_stage_opamp_dummy_magic_26_0.VD4.n9 1.02133
R22141 two_stage_opamp_dummy_magic_26_0.VD4.n33 two_stage_opamp_dummy_magic_26_0.VD4.n6 1.02133
R22142 two_stage_opamp_dummy_magic_26_0.VD4.n20 two_stage_opamp_dummy_magic_26_0.VD4.n2 1.02133
R22143 two_stage_opamp_dummy_magic_26_0.VD4.n0 two_stage_opamp_dummy_magic_26_0.VD4.n28 1.02133
R22144 two_stage_opamp_dummy_magic_26_0.VD4.n25 two_stage_opamp_dummy_magic_26_0.VD4.n14 1.02133
R22145 two_stage_opamp_dummy_magic_26_0.VD4 two_stage_opamp_dummy_magic_26_0.VD4.n2 0.65675
R22146 two_stage_opamp_dummy_magic_26_0.VD4.n31 two_stage_opamp_dummy_magic_26_0.VD4.n30 0.643357
R22147 two_stage_opamp_dummy_magic_26_0.VD4.n32 two_stage_opamp_dummy_magic_26_0.VD4.n3 0.643357
R22148 two_stage_opamp_dummy_magic_26_0.VD4.n34 two_stage_opamp_dummy_magic_26_0.VD4.n33 0.643357
R22149 two_stage_opamp_dummy_magic_26_0.VD4.n1 two_stage_opamp_dummy_magic_26_0.VD4.n0 0.0280497
R22150 two_stage_opamp_dummy_magic_26_0.VD4.n22 two_stage_opamp_dummy_magic_26_0.VD4.n21 0.3755
R22151 two_stage_opamp_dummy_magic_26_0.VD4.n23 two_stage_opamp_dummy_magic_26_0.VD4.n22 0.3755
R22152 two_stage_opamp_dummy_magic_26_0.VD4.n26 two_stage_opamp_dummy_magic_26_0.VD4.n23 0.3755
R22153 two_stage_opamp_dummy_magic_26_0.VD4.n0 two_stage_opamp_dummy_magic_26_0.VD4.n18 0.132669
R22154 two_stage_opamp_dummy_magic_26_0.VD4.n15 two_stage_opamp_dummy_magic_26_0.VD4.n2 0.104667
R22155 two_stage_opamp_dummy_magic_26_0.VD4.n1 two_stage_opamp_dummy_magic_26_0.VD4.n14 0.0473045
R22156 two_stage_opamp_dummy_magic_26_0.VD4.n34 two_stage_opamp_dummy_magic_26_0.VD4.n3 0.0540714
R22157 two_stage_opamp_dummy_magic_26_0.VD4.n30 two_stage_opamp_dummy_magic_26_0.VD4.n3 0.0540714
R22158 two_stage_opamp_dummy_magic_26_0.VD4.n30 two_stage_opamp_dummy_magic_26_0.VD4.n1 0.274553
R22159 two_stage_opamp_dummy_magic_26_0.VD4.n33 two_stage_opamp_dummy_magic_26_0.VD4.n2 0.0540714
R22160 two_stage_opamp_dummy_magic_26_0.VD4.n33 two_stage_opamp_dummy_magic_26_0.VD4.n32 0.0540714
R22161 two_stage_opamp_dummy_magic_26_0.VD4.n32 two_stage_opamp_dummy_magic_26_0.VD4.n31 0.0540714
R22162 two_stage_opamp_dummy_magic_26_0.VD4.n31 two_stage_opamp_dummy_magic_26_0.VD4.n14 0.0540714
R22163 two_stage_opamp_dummy_magic_26_0.VD4 two_stage_opamp_dummy_magic_26_0.VD4.n34 0.0406786
R22164 two_stage_opamp_dummy_magic_26_0.VD3.n3 two_stage_opamp_dummy_magic_26_0.VD3.t22 671.418
R22165 two_stage_opamp_dummy_magic_26_0.VD3.n16 two_stage_opamp_dummy_magic_26_0.VD3.t25 671.418
R22166 two_stage_opamp_dummy_magic_26_0.VD3.n15 two_stage_opamp_dummy_magic_26_0.VD3.t26 213.131
R22167 two_stage_opamp_dummy_magic_26_0.VD3.t23 two_stage_opamp_dummy_magic_26_0.VD3.n14 213.131
R22168 two_stage_opamp_dummy_magic_26_0.VD3.t26 two_stage_opamp_dummy_magic_26_0.VD3.t8 146.155
R22169 two_stage_opamp_dummy_magic_26_0.VD3.t8 two_stage_opamp_dummy_magic_26_0.VD3.t12 146.155
R22170 two_stage_opamp_dummy_magic_26_0.VD3.t12 two_stage_opamp_dummy_magic_26_0.VD3.t18 146.155
R22171 two_stage_opamp_dummy_magic_26_0.VD3.t18 two_stage_opamp_dummy_magic_26_0.VD3.t2 146.155
R22172 two_stage_opamp_dummy_magic_26_0.VD3.t2 two_stage_opamp_dummy_magic_26_0.VD3.t4 146.155
R22173 two_stage_opamp_dummy_magic_26_0.VD3.t4 two_stage_opamp_dummy_magic_26_0.VD3.t6 146.155
R22174 two_stage_opamp_dummy_magic_26_0.VD3.t6 two_stage_opamp_dummy_magic_26_0.VD3.t10 146.155
R22175 two_stage_opamp_dummy_magic_26_0.VD3.t10 two_stage_opamp_dummy_magic_26_0.VD3.t14 146.155
R22176 two_stage_opamp_dummy_magic_26_0.VD3.t14 two_stage_opamp_dummy_magic_26_0.VD3.t0 146.155
R22177 two_stage_opamp_dummy_magic_26_0.VD3.t0 two_stage_opamp_dummy_magic_26_0.VD3.t16 146.155
R22178 two_stage_opamp_dummy_magic_26_0.VD3.t16 two_stage_opamp_dummy_magic_26_0.VD3.t23 146.155
R22179 two_stage_opamp_dummy_magic_26_0.VD3.n15 two_stage_opamp_dummy_magic_26_0.VD3.t27 76.2576
R22180 two_stage_opamp_dummy_magic_26_0.VD3.n14 two_stage_opamp_dummy_magic_26_0.VD3.t24 76.2576
R22181 two_stage_opamp_dummy_magic_26_0.VD3.n0 two_stage_opamp_dummy_magic_26_0.VD3.n19 67.013
R22182 two_stage_opamp_dummy_magic_26_0.VD3.n13 two_stage_opamp_dummy_magic_26_0.VD3.n12 67.013
R22183 two_stage_opamp_dummy_magic_26_0.VD3.n32 two_stage_opamp_dummy_magic_26_0.VD3.n9 67.013
R22184 two_stage_opamp_dummy_magic_26_0.VD3.n33 two_stage_opamp_dummy_magic_26_0.VD3.n6 67.013
R22185 two_stage_opamp_dummy_magic_26_0.VD3.n29 two_stage_opamp_dummy_magic_26_0.VD3.n28 67.013
R22186 two_stage_opamp_dummy_magic_26_0.VD3.n5 two_stage_opamp_dummy_magic_26_0.VD3.n4 66.0338
R22187 two_stage_opamp_dummy_magic_26_0.VD3.n8 two_stage_opamp_dummy_magic_26_0.VD3.n7 66.0338
R22188 two_stage_opamp_dummy_magic_26_0.VD3.n11 two_stage_opamp_dummy_magic_26_0.VD3.n10 66.0338
R22189 two_stage_opamp_dummy_magic_26_0.VD3.n23 two_stage_opamp_dummy_magic_26_0.VD3.n22 66.0338
R22190 two_stage_opamp_dummy_magic_26_0.VD3.n18 two_stage_opamp_dummy_magic_26_0.VD3.n17 66.0338
R22191 two_stage_opamp_dummy_magic_26_0.VD3.n27 two_stage_opamp_dummy_magic_26_0.VD3.n26 66.0338
R22192 two_stage_opamp_dummy_magic_26_0.VD3.n19 two_stage_opamp_dummy_magic_26_0.VD3.t9 11.2576
R22193 two_stage_opamp_dummy_magic_26_0.VD3.n19 two_stage_opamp_dummy_magic_26_0.VD3.t13 11.2576
R22194 two_stage_opamp_dummy_magic_26_0.VD3.n12 two_stage_opamp_dummy_magic_26_0.VD3.t5 11.2576
R22195 two_stage_opamp_dummy_magic_26_0.VD3.n12 two_stage_opamp_dummy_magic_26_0.VD3.t7 11.2576
R22196 two_stage_opamp_dummy_magic_26_0.VD3.n9 two_stage_opamp_dummy_magic_26_0.VD3.t11 11.2576
R22197 two_stage_opamp_dummy_magic_26_0.VD3.n9 two_stage_opamp_dummy_magic_26_0.VD3.t15 11.2576
R22198 two_stage_opamp_dummy_magic_26_0.VD3.n6 two_stage_opamp_dummy_magic_26_0.VD3.t1 11.2576
R22199 two_stage_opamp_dummy_magic_26_0.VD3.n6 two_stage_opamp_dummy_magic_26_0.VD3.t17 11.2576
R22200 two_stage_opamp_dummy_magic_26_0.VD3.n4 two_stage_opamp_dummy_magic_26_0.VD3.t32 11.2576
R22201 two_stage_opamp_dummy_magic_26_0.VD3.n4 two_stage_opamp_dummy_magic_26_0.VD3.t36 11.2576
R22202 two_stage_opamp_dummy_magic_26_0.VD3.n7 two_stage_opamp_dummy_magic_26_0.VD3.t21 11.2576
R22203 two_stage_opamp_dummy_magic_26_0.VD3.n7 two_stage_opamp_dummy_magic_26_0.VD3.t33 11.2576
R22204 two_stage_opamp_dummy_magic_26_0.VD3.n10 two_stage_opamp_dummy_magic_26_0.VD3.t20 11.2576
R22205 two_stage_opamp_dummy_magic_26_0.VD3.n10 two_stage_opamp_dummy_magic_26_0.VD3.t29 11.2576
R22206 two_stage_opamp_dummy_magic_26_0.VD3.n22 two_stage_opamp_dummy_magic_26_0.VD3.t34 11.2576
R22207 two_stage_opamp_dummy_magic_26_0.VD3.n22 two_stage_opamp_dummy_magic_26_0.VD3.t37 11.2576
R22208 two_stage_opamp_dummy_magic_26_0.VD3.n17 two_stage_opamp_dummy_magic_26_0.VD3.t31 11.2576
R22209 two_stage_opamp_dummy_magic_26_0.VD3.n17 two_stage_opamp_dummy_magic_26_0.VD3.t30 11.2576
R22210 two_stage_opamp_dummy_magic_26_0.VD3.n26 two_stage_opamp_dummy_magic_26_0.VD3.t35 11.2576
R22211 two_stage_opamp_dummy_magic_26_0.VD3.n26 two_stage_opamp_dummy_magic_26_0.VD3.t28 11.2576
R22212 two_stage_opamp_dummy_magic_26_0.VD3.n28 two_stage_opamp_dummy_magic_26_0.VD3.t19 11.2576
R22213 two_stage_opamp_dummy_magic_26_0.VD3.n28 two_stage_opamp_dummy_magic_26_0.VD3.t3 11.2576
R22214 two_stage_opamp_dummy_magic_26_0.VD3.n27 two_stage_opamp_dummy_magic_26_0.VD3.n25 5.66717
R22215 two_stage_opamp_dummy_magic_26_0.VD3.n20 two_stage_opamp_dummy_magic_26_0.VD3.n5 5.66717
R22216 two_stage_opamp_dummy_magic_26_0.VD3.n20 two_stage_opamp_dummy_magic_26_0.VD3.n8 5.29217
R22217 two_stage_opamp_dummy_magic_26_0.VD3.n21 two_stage_opamp_dummy_magic_26_0.VD3.n11 5.29217
R22218 two_stage_opamp_dummy_magic_26_0.VD3.n24 two_stage_opamp_dummy_magic_26_0.VD3.n23 5.29217
R22219 two_stage_opamp_dummy_magic_26_0.VD3.n25 two_stage_opamp_dummy_magic_26_0.VD3.n18 5.29217
R22220 two_stage_opamp_dummy_magic_26_0.VD3.n16 two_stage_opamp_dummy_magic_26_0.VD3.n15 1.90883
R22221 two_stage_opamp_dummy_magic_26_0.VD3.n14 two_stage_opamp_dummy_magic_26_0.VD3.n3 1.90883
R22222 two_stage_opamp_dummy_magic_26_0.VD3.n33 two_stage_opamp_dummy_magic_26_0.VD3.n8 1.02133
R22223 two_stage_opamp_dummy_magic_26_0.VD3.n32 two_stage_opamp_dummy_magic_26_0.VD3.n11 1.02133
R22224 two_stage_opamp_dummy_magic_26_0.VD3.n23 two_stage_opamp_dummy_magic_26_0.VD3.n13 1.02133
R22225 two_stage_opamp_dummy_magic_26_0.VD3.n29 two_stage_opamp_dummy_magic_26_0.VD3.n18 1.02133
R22226 two_stage_opamp_dummy_magic_26_0.VD3.n0 two_stage_opamp_dummy_magic_26_0.VD3.n27 1.02133
R22227 two_stage_opamp_dummy_magic_26_0.VD3.n34 two_stage_opamp_dummy_magic_26_0.VD3.n5 1.02133
R22228 two_stage_opamp_dummy_magic_26_0.VD3 two_stage_opamp_dummy_magic_26_0.VD3.n34 0.65675
R22229 two_stage_opamp_dummy_magic_26_0.VD3.n33 two_stage_opamp_dummy_magic_26_0.VD3.n2 0.643357
R22230 two_stage_opamp_dummy_magic_26_0.VD3.n32 two_stage_opamp_dummy_magic_26_0.VD3.n31 0.643357
R22231 two_stage_opamp_dummy_magic_26_0.VD3.n30 two_stage_opamp_dummy_magic_26_0.VD3.n13 0.643357
R22232 two_stage_opamp_dummy_magic_26_0.VD3.n1 two_stage_opamp_dummy_magic_26_0.VD3.n0 0.0279681
R22233 two_stage_opamp_dummy_magic_26_0.VD3.n25 two_stage_opamp_dummy_magic_26_0.VD3.n24 0.3755
R22234 two_stage_opamp_dummy_magic_26_0.VD3.n24 two_stage_opamp_dummy_magic_26_0.VD3.n21 0.3755
R22235 two_stage_opamp_dummy_magic_26_0.VD3.n21 two_stage_opamp_dummy_magic_26_0.VD3.n20 0.3755
R22236 two_stage_opamp_dummy_magic_26_0.VD3.n0 two_stage_opamp_dummy_magic_26_0.VD3.n16 0.131952
R22237 two_stage_opamp_dummy_magic_26_0.VD3.n34 two_stage_opamp_dummy_magic_26_0.VD3.n3 0.104667
R22238 two_stage_opamp_dummy_magic_26_0.VD3.n29 two_stage_opamp_dummy_magic_26_0.VD3.n1 0.0471695
R22239 two_stage_opamp_dummy_magic_26_0.VD3.n30 two_stage_opamp_dummy_magic_26_0.VD3.n1 0.274589
R22240 two_stage_opamp_dummy_magic_26_0.VD3.n31 two_stage_opamp_dummy_magic_26_0.VD3.n30 0.0540714
R22241 two_stage_opamp_dummy_magic_26_0.VD3.n31 two_stage_opamp_dummy_magic_26_0.VD3.n2 0.0540714
R22242 two_stage_opamp_dummy_magic_26_0.VD3.n29 two_stage_opamp_dummy_magic_26_0.VD3.n13 0.0540714
R22243 two_stage_opamp_dummy_magic_26_0.VD3.n32 two_stage_opamp_dummy_magic_26_0.VD3.n13 0.0540714
R22244 two_stage_opamp_dummy_magic_26_0.VD3.n33 two_stage_opamp_dummy_magic_26_0.VD3.n32 0.0540714
R22245 two_stage_opamp_dummy_magic_26_0.VD3.n34 two_stage_opamp_dummy_magic_26_0.VD3.n33 0.0540714
R22246 two_stage_opamp_dummy_magic_26_0.VD3 two_stage_opamp_dummy_magic_26_0.VD3.n2 0.0406786
R22247 two_stage_opamp_dummy_magic_26_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_26_0.err_amp_mir.t5 573.044
R22248 two_stage_opamp_dummy_magic_26_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_26_0.err_amp_mir.t1 433.8
R22249 two_stage_opamp_dummy_magic_26_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_26_0.err_amp_mir.n0 184.09
R22250 two_stage_opamp_dummy_magic_26_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_26_0.err_amp_mir.n1 163.978
R22251 two_stage_opamp_dummy_magic_26_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_26_0.err_amp_mir.n2 33.0088
R22252 two_stage_opamp_dummy_magic_26_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_26_0.err_amp_mir.t3 15.7605
R22253 two_stage_opamp_dummy_magic_26_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_26_0.err_amp_mir.t4 15.7605
R22254 two_stage_opamp_dummy_magic_26_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_26_0.err_amp_mir.t2 9.6005
R22255 two_stage_opamp_dummy_magic_26_0.err_amp_mir.t0 two_stage_opamp_dummy_magic_26_0.err_amp_mir.n3 9.6005
R22256 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n0 344.837
R22257 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n1 344.274
R22258 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n3 292.5
R22259 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t0 121.785
R22260 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n7 118.861
R22261 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n9 118.861
R22262 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n13 118.861
R22263 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n16 118.861
R22264 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n19 118.861
R22265 bgr_11_0.V_CMFB_S1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n22 76.0943
R22266 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n2 52.3363
R22267 bgr_11_0.V_CMFB_S1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n4 52.2813
R22268 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t15 39.4005
R22269 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t12 39.4005
R22270 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t14 39.4005
R22271 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t13 39.4005
R22272 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t11 39.4005
R22273 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t16 39.4005
R22274 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t1 19.7005
R22275 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t6 19.7005
R22276 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t2 19.7005
R22277 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t7 19.7005
R22278 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t4 19.7005
R22279 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t8 19.7005
R22280 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t3 19.7005
R22281 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t10 19.7005
R22282 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t5 19.7005
R22283 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t9 19.7005
R22284 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n21 5.90675
R22285 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n8 5.60467
R22286 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n18 5.54217
R22287 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n6 5.54217
R22288 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n10 5.04217
R22289 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n12 5.04217
R22290 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n5 5.04217
R22291 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n20 5.04217
R22292 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n6 4.97967
R22293 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n14 4.97967
R22294 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n17 4.97967
R22295 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n15 0.563
R22296 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n6 0.563
R22297 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n11 0.563
R22298 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n5 0.563
R22299 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n5 0.563
R22300 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n21 344.178
R22301 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n22 334.772
R22302 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.t37 312.798
R22303 bgr_11_0.V_TOP bgr_11_0.V_TOP.t21 312.639
R22304 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.t45 312.5
R22305 bgr_11_0.V_TOP.n42 bgr_11_0.V_TOP.t33 310.401
R22306 bgr_11_0.V_TOP.n41 bgr_11_0.V_TOP.t42 310.401
R22307 bgr_11_0.V_TOP.n40 bgr_11_0.V_TOP.t49 310.401
R22308 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.t26 310.401
R22309 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.t25 310.401
R22310 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.t36 310.401
R22311 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.t27 310.401
R22312 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.t39 310.401
R22313 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.t48 310.401
R22314 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.t23 310.401
R22315 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.t38 310.401
R22316 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.t14 308
R22317 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.t29 305.901
R22318 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n30 301.933
R22319 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n28 301.933
R22320 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n26 301.933
R22321 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n20 297.433
R22322 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.t12 108.424
R22323 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.t6 99.5675
R22324 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t8 39.4005
R22325 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t0 39.4005
R22326 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t13 39.4005
R22327 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t10 39.4005
R22328 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t9 39.4005
R22329 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t11 39.4005
R22330 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.t1 39.4005
R22331 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.t7 39.4005
R22332 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t5 39.4005
R22333 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t2 39.4005
R22334 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t4 39.4005
R22335 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t3 39.4005
R22336 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.n18 29.1779
R22337 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n19 16.5063
R22338 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.n31 4.90675
R22339 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t24 4.8295
R22340 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t46 4.8295
R22341 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t34 4.8295
R22342 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t18 4.8295
R22343 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t22 4.8295
R22344 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t44 4.8295
R22345 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t47 4.8295
R22346 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.t35 4.8295
R22347 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.t41 4.8295
R22348 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t32 4.5005
R22349 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t19 4.5005
R22350 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t40 4.5005
R22351 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t31 4.5005
R22352 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t30 4.5005
R22353 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t17 4.5005
R22354 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t16 4.5005
R22355 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.t43 4.5005
R22356 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.t20 4.5005
R22357 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.t28 4.5005
R22358 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.t15 4.5005
R22359 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.n6 4.5005
R22360 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n0 4.5005
R22361 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.n34 4.5005
R22362 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n24 4.5005
R22363 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n23 1.59425
R22364 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n32 1.21925
R22365 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n25 1.1255
R22366 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n27 1.1255
R22367 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n29 1.1255
R22368 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.n8 0.3295
R22369 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n10 0.3295
R22370 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n12 0.3295
R22371 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.n14 0.3295
R22372 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.n17 0.3295
R22373 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.n16 0.3295
R22374 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n9 0.2825
R22375 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n11 0.2825
R22376 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.n13 0.2825
R22377 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.n15 0.2825
R22378 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.n1 0.28175
R22379 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.n2 0.28175
R22380 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.n3 0.28175
R22381 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.n4 0.28175
R22382 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.n5 0.28175
R22383 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.n35 0.28175
R22384 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.n36 0.28175
R22385 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.n37 0.28175
R22386 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.n38 0.28175
R22387 bgr_11_0.V_TOP.n40 bgr_11_0.V_TOP.n39 0.28175
R22388 bgr_11_0.V_TOP.n41 bgr_11_0.V_TOP.n40 0.28175
R22389 bgr_11_0.V_TOP.n42 bgr_11_0.V_TOP.n41 0.28175
R22390 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.n0 0.141125
R22391 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.n0 0.141125
R22392 bgr_11_0.V_TOP bgr_11_0.V_TOP.n42 0.141125
R22393 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n7 0.141125
R22394 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.n33 0.141125
R22395 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t7 651.343
R22396 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t8 647.968
R22397 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t9 537.922
R22398 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t0 117.243
R22399 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n1 107.266
R22400 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n4 105.016
R22401 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n2 105.016
R22402 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t3 13.1338
R22403 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t6 13.1338
R22404 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t4 13.1338
R22405 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t1 13.1338
R22406 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t5 13.1338
R22407 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t2 13.1338
R22408 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n5 7.32862
R22409 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n6 3.98488
R22410 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n3 2.2505
R22411 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n0 1.73488
R22412 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n7 1.53175
R22413 bgr_11_0.1st_Vout_1.n12 bgr_11_0.1st_Vout_1.t29 363.909
R22414 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.t13 351.88
R22415 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n22 299.25
R22416 bgr_11_0.1st_Vout_1.n14 bgr_11_0.1st_Vout_1.n13 299.25
R22417 bgr_11_0.1st_Vout_1.n18 bgr_11_0.1st_Vout_1.n17 297.807
R22418 bgr_11_0.1st_Vout_1.n20 bgr_11_0.1st_Vout_1.t30 194.809
R22419 bgr_11_0.1st_Vout_1.n20 bgr_11_0.1st_Vout_1.t10 194.809
R22420 bgr_11_0.1st_Vout_1.n15 bgr_11_0.1st_Vout_1.t28 194.809
R22421 bgr_11_0.1st_Vout_1.n15 bgr_11_0.1st_Vout_1.t19 194.809
R22422 bgr_11_0.1st_Vout_1.n21 bgr_11_0.1st_Vout_1.n20 163.097
R22423 bgr_11_0.1st_Vout_1.n16 bgr_11_0.1st_Vout_1.n15 163.097
R22424 bgr_11_0.1st_Vout_1.n18 bgr_11_0.1st_Vout_1.t3 49.4474
R22425 bgr_11_0.1st_Vout_1.n22 bgr_11_0.1st_Vout_1.t4 39.4005
R22426 bgr_11_0.1st_Vout_1.n22 bgr_11_0.1st_Vout_1.t6 39.4005
R22427 bgr_11_0.1st_Vout_1.n13 bgr_11_0.1st_Vout_1.t2 39.4005
R22428 bgr_11_0.1st_Vout_1.n13 bgr_11_0.1st_Vout_1.t0 39.4005
R22429 bgr_11_0.1st_Vout_1.n17 bgr_11_0.1st_Vout_1.t5 39.4005
R22430 bgr_11_0.1st_Vout_1.n17 bgr_11_0.1st_Vout_1.t1 39.4005
R22431 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t27 4.8295
R22432 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t14 4.8295
R22433 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.t32 4.8295
R22434 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t22 4.8295
R22435 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t25 4.8295
R22436 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t12 4.8295
R22437 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t16 4.8295
R22438 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t7 4.8295
R22439 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.t24 4.8295
R22440 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t18 4.5005
R22441 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t23 4.5005
R22442 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.t26 4.5005
R22443 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t31 4.5005
R22444 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t17 4.5005
R22445 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t21 4.5005
R22446 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t8 4.5005
R22447 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t11 4.5005
R22448 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.t15 4.5005
R22449 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.t20 4.5005
R22450 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.t9 4.5005
R22451 bgr_11_0.1st_Vout_1.n19 bgr_11_0.1st_Vout_1.n18 1.44719
R22452 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.n1 0.3295
R22453 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n3 0.3295
R22454 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.n5 0.3295
R22455 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.n7 0.3295
R22456 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.n9 0.3295
R22457 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.n10 0.3295
R22458 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n2 0.2825
R22459 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.n4 0.2825
R22460 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.n6 0.2825
R22461 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.n8 0.2825
R22462 bgr_11_0.1st_Vout_1.n19 bgr_11_0.1st_Vout_1.n16 0.2505
R22463 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n21 0.2505
R22464 bgr_11_0.1st_Vout_1.n14 bgr_11_0.1st_Vout_1.n12 0.21925
R22465 bgr_11_0.1st_Vout_1.n16 bgr_11_0.1st_Vout_1.n14 0.1255
R22466 bgr_11_0.1st_Vout_1.n21 bgr_11_0.1st_Vout_1.n19 0.1255
R22467 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n0 0.09425
R22468 bgr_11_0.1st_Vout_1.n12 bgr_11_0.1st_Vout_1.n11 10.102
R22469 bgr_11_0.cap_res1.t20 bgr_11_0.cap_res1.t13 121.983
R22470 bgr_11_0.cap_res1.t9 bgr_11_0.cap_res1.t17 0.1603
R22471 bgr_11_0.cap_res1.t16 bgr_11_0.cap_res1.t19 0.1603
R22472 bgr_11_0.cap_res1.t8 bgr_11_0.cap_res1.t15 0.1603
R22473 bgr_11_0.cap_res1.t1 bgr_11_0.cap_res1.t7 0.1603
R22474 bgr_11_0.cap_res1.t6 bgr_11_0.cap_res1.t14 0.1603
R22475 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t10 0.159278
R22476 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t3 0.159278
R22477 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t11 0.159278
R22478 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t18 0.159278
R22479 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t9 0.1368
R22480 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t5 0.1368
R22481 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t16 0.1368
R22482 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t12 0.1368
R22483 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t8 0.1368
R22484 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t4 0.1368
R22485 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t1 0.1368
R22486 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t0 0.1368
R22487 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t6 0.1368
R22488 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t2 0.1368
R22489 bgr_11_0.cap_res1.t10 bgr_11_0.cap_res1.n0 0.00152174
R22490 bgr_11_0.cap_res1.t3 bgr_11_0.cap_res1.n1 0.00152174
R22491 bgr_11_0.cap_res1.t11 bgr_11_0.cap_res1.n2 0.00152174
R22492 bgr_11_0.cap_res1.t18 bgr_11_0.cap_res1.n3 0.00152174
R22493 bgr_11_0.cap_res1.t13 bgr_11_0.cap_res1.n4 0.00152174
R22494 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t6 369.534
R22495 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t9 369.534
R22496 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.t22 369.534
R22497 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t20 369.534
R22498 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.t13 369.534
R22499 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.t11 369.534
R22500 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.t1 369.534
R22501 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n1 360.288
R22502 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.t7 249.034
R22503 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.t5 192.8
R22504 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.t12 192.8
R22505 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t19 192.8
R22506 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t18 192.8
R22507 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.t15 192.8
R22508 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.t23 192.8
R22509 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t8 192.8
R22510 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.t10 192.8
R22511 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.t17 192.8
R22512 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.t16 192.8
R22513 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.t21 192.8
R22514 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.t14 192.8
R22515 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.n4 176.733
R22516 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.n3 176.733
R22517 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.n8 176.733
R22518 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.n12 176.733
R22519 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.n13 176.733
R22520 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.n6 168.014
R22521 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.n10 166.343
R22522 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.n16 166.343
R22523 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n19 166.343
R22524 bgr_11_0.NFET_GATE_10uA.n20 bgr_11_0.NFET_GATE_10uA.n0 141.752
R22525 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n5 56.2338
R22526 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n2 56.2338
R22527 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.n9 56.2338
R22528 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.n7 56.2338
R22529 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n15 56.2338
R22530 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n14 56.2338
R22531 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.n18 56.2338
R22532 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t4 39.4005
R22533 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t3 39.4005
R22534 bgr_11_0.NFET_GATE_10uA.t0 bgr_11_0.NFET_GATE_10uA.n20 24.0005
R22535 bgr_11_0.NFET_GATE_10uA.n20 bgr_11_0.NFET_GATE_10uA.t2 24.0005
R22536 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n17 2.01612
R22537 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.n11 1.5005
R22538 two_stage_opamp_dummy_magic_26_0.VD2.n1 two_stage_opamp_dummy_magic_26_0.VD2.n0 49.7255
R22539 two_stage_opamp_dummy_magic_26_0.VD2.n25 two_stage_opamp_dummy_magic_26_0.VD2.n24 49.7255
R22540 two_stage_opamp_dummy_magic_26_0.VD2.n27 two_stage_opamp_dummy_magic_26_0.VD2.n9 49.7255
R22541 two_stage_opamp_dummy_magic_26_0.VD2.n21 two_stage_opamp_dummy_magic_26_0.VD2.n12 49.7255
R22542 two_stage_opamp_dummy_magic_26_0.VD2.n11 two_stage_opamp_dummy_magic_26_0.VD2.n10 49.7255
R22543 two_stage_opamp_dummy_magic_26_0.VD2.n15 two_stage_opamp_dummy_magic_26_0.VD2.n14 49.3505
R22544 two_stage_opamp_dummy_magic_26_0.VD2.n8 two_stage_opamp_dummy_magic_26_0.VD2.n7 49.3505
R22545 two_stage_opamp_dummy_magic_26_0.VD2.n31 two_stage_opamp_dummy_magic_26_0.VD2.n30 49.3505
R22546 two_stage_opamp_dummy_magic_26_0.VD2.n35 two_stage_opamp_dummy_magic_26_0.VD2.n34 49.3505
R22547 two_stage_opamp_dummy_magic_26_0.VD2.n5 two_stage_opamp_dummy_magic_26_0.VD2.n4 49.3505
R22548 two_stage_opamp_dummy_magic_26_0.VD2.n18 two_stage_opamp_dummy_magic_26_0.VD2.n17 49.3505
R22549 two_stage_opamp_dummy_magic_26_0.VD2.n14 two_stage_opamp_dummy_magic_26_0.VD2.t5 16.0005
R22550 two_stage_opamp_dummy_magic_26_0.VD2.n14 two_stage_opamp_dummy_magic_26_0.VD2.t8 16.0005
R22551 two_stage_opamp_dummy_magic_26_0.VD2.n7 two_stage_opamp_dummy_magic_26_0.VD2.t4 16.0005
R22552 two_stage_opamp_dummy_magic_26_0.VD2.n7 two_stage_opamp_dummy_magic_26_0.VD2.t6 16.0005
R22553 two_stage_opamp_dummy_magic_26_0.VD2.n30 two_stage_opamp_dummy_magic_26_0.VD2.t21 16.0005
R22554 two_stage_opamp_dummy_magic_26_0.VD2.n30 two_stage_opamp_dummy_magic_26_0.VD2.t9 16.0005
R22555 two_stage_opamp_dummy_magic_26_0.VD2.n34 two_stage_opamp_dummy_magic_26_0.VD2.t20 16.0005
R22556 two_stage_opamp_dummy_magic_26_0.VD2.n34 two_stage_opamp_dummy_magic_26_0.VD2.t3 16.0005
R22557 two_stage_opamp_dummy_magic_26_0.VD2.n4 two_stage_opamp_dummy_magic_26_0.VD2.t2 16.0005
R22558 two_stage_opamp_dummy_magic_26_0.VD2.n4 two_stage_opamp_dummy_magic_26_0.VD2.t1 16.0005
R22559 two_stage_opamp_dummy_magic_26_0.VD2.n0 two_stage_opamp_dummy_magic_26_0.VD2.t18 16.0005
R22560 two_stage_opamp_dummy_magic_26_0.VD2.n0 two_stage_opamp_dummy_magic_26_0.VD2.t13 16.0005
R22561 two_stage_opamp_dummy_magic_26_0.VD2.n24 two_stage_opamp_dummy_magic_26_0.VD2.t16 16.0005
R22562 two_stage_opamp_dummy_magic_26_0.VD2.n24 two_stage_opamp_dummy_magic_26_0.VD2.t12 16.0005
R22563 two_stage_opamp_dummy_magic_26_0.VD2.n9 two_stage_opamp_dummy_magic_26_0.VD2.t15 16.0005
R22564 two_stage_opamp_dummy_magic_26_0.VD2.n9 two_stage_opamp_dummy_magic_26_0.VD2.t11 16.0005
R22565 two_stage_opamp_dummy_magic_26_0.VD2.n12 two_stage_opamp_dummy_magic_26_0.VD2.t17 16.0005
R22566 two_stage_opamp_dummy_magic_26_0.VD2.n12 two_stage_opamp_dummy_magic_26_0.VD2.t10 16.0005
R22567 two_stage_opamp_dummy_magic_26_0.VD2.n17 two_stage_opamp_dummy_magic_26_0.VD2.t7 16.0005
R22568 two_stage_opamp_dummy_magic_26_0.VD2.n17 two_stage_opamp_dummy_magic_26_0.VD2.t0 16.0005
R22569 two_stage_opamp_dummy_magic_26_0.VD2.n10 two_stage_opamp_dummy_magic_26_0.VD2.t19 16.0005
R22570 two_stage_opamp_dummy_magic_26_0.VD2.n10 two_stage_opamp_dummy_magic_26_0.VD2.t14 16.0005
R22571 two_stage_opamp_dummy_magic_26_0.VD2.n25 two_stage_opamp_dummy_magic_26_0.VD2.n3 7.33383
R22572 two_stage_opamp_dummy_magic_26_0.VD2.n28 two_stage_opamp_dummy_magic_26_0.VD2.n27 7.33383
R22573 two_stage_opamp_dummy_magic_26_0.VD2.n21 two_stage_opamp_dummy_magic_26_0.VD2.n20 7.33383
R22574 two_stage_opamp_dummy_magic_26_0.VD2.n13 two_stage_opamp_dummy_magic_26_0.VD2.n11 7.33383
R22575 two_stage_opamp_dummy_magic_26_0.VD2.n32 two_stage_opamp_dummy_magic_26_0.VD2.n8 5.438
R22576 two_stage_opamp_dummy_magic_26_0.VD2.n16 two_stage_opamp_dummy_magic_26_0.VD2.n15 5.438
R22577 two_stage_opamp_dummy_magic_26_0.VD2.n28 two_stage_opamp_dummy_magic_26_0.VD2.n8 5.31821
R22578 two_stage_opamp_dummy_magic_26_0.VD2.n15 two_stage_opamp_dummy_magic_26_0.VD2.n13 5.31821
R22579 two_stage_opamp_dummy_magic_26_0.VD2.n31 two_stage_opamp_dummy_magic_26_0.VD2.n29 5.08383
R22580 two_stage_opamp_dummy_magic_26_0.VD2.n36 two_stage_opamp_dummy_magic_26_0.VD2.n35 5.08383
R22581 two_stage_opamp_dummy_magic_26_0.VD2.n5 two_stage_opamp_dummy_magic_26_0.VD2.n2 5.08383
R22582 two_stage_opamp_dummy_magic_26_0.VD2.n19 two_stage_opamp_dummy_magic_26_0.VD2.n18 5.08383
R22583 two_stage_opamp_dummy_magic_26_0.VD2.n27 two_stage_opamp_dummy_magic_26_0.VD2.n26 5.063
R22584 two_stage_opamp_dummy_magic_26_0.VD2.n22 two_stage_opamp_dummy_magic_26_0.VD2.n11 5.063
R22585 two_stage_opamp_dummy_magic_26_0.VD2.n32 two_stage_opamp_dummy_magic_26_0.VD2.n31 4.8755
R22586 two_stage_opamp_dummy_magic_26_0.VD2.n35 two_stage_opamp_dummy_magic_26_0.VD2.n33 4.8755
R22587 two_stage_opamp_dummy_magic_26_0.VD2.n6 two_stage_opamp_dummy_magic_26_0.VD2.n5 4.8755
R22588 two_stage_opamp_dummy_magic_26_0.VD2.n18 two_stage_opamp_dummy_magic_26_0.VD2.n16 4.8755
R22589 two_stage_opamp_dummy_magic_26_0.VD2 two_stage_opamp_dummy_magic_26_0.VD2.n37 4.60467
R22590 two_stage_opamp_dummy_magic_26_0.VD2.n26 two_stage_opamp_dummy_magic_26_0.VD2.n25 4.5005
R22591 two_stage_opamp_dummy_magic_26_0.VD2.n23 two_stage_opamp_dummy_magic_26_0.VD2.n1 4.5005
R22592 two_stage_opamp_dummy_magic_26_0.VD2.n22 two_stage_opamp_dummy_magic_26_0.VD2.n21 4.5005
R22593 two_stage_opamp_dummy_magic_26_0.VD2 two_stage_opamp_dummy_magic_26_0.VD2.n1 2.72967
R22594 two_stage_opamp_dummy_magic_26_0.VD2.n26 two_stage_opamp_dummy_magic_26_0.VD2.n23 0.563
R22595 two_stage_opamp_dummy_magic_26_0.VD2.n23 two_stage_opamp_dummy_magic_26_0.VD2.n22 0.563
R22596 two_stage_opamp_dummy_magic_26_0.VD2.n33 two_stage_opamp_dummy_magic_26_0.VD2.n32 0.563
R22597 two_stage_opamp_dummy_magic_26_0.VD2.n33 two_stage_opamp_dummy_magic_26_0.VD2.n6 0.563
R22598 two_stage_opamp_dummy_magic_26_0.VD2.n16 two_stage_opamp_dummy_magic_26_0.VD2.n6 0.563
R22599 two_stage_opamp_dummy_magic_26_0.VD2.n19 two_stage_opamp_dummy_magic_26_0.VD2.n13 0.234875
R22600 two_stage_opamp_dummy_magic_26_0.VD2.n20 two_stage_opamp_dummy_magic_26_0.VD2.n19 0.234875
R22601 two_stage_opamp_dummy_magic_26_0.VD2.n20 two_stage_opamp_dummy_magic_26_0.VD2.n2 0.234875
R22602 two_stage_opamp_dummy_magic_26_0.VD2.n37 two_stage_opamp_dummy_magic_26_0.VD2.n2 0.234875
R22603 two_stage_opamp_dummy_magic_26_0.VD2.n37 two_stage_opamp_dummy_magic_26_0.VD2.n36 0.234875
R22604 two_stage_opamp_dummy_magic_26_0.VD2.n36 two_stage_opamp_dummy_magic_26_0.VD2.n3 0.234875
R22605 two_stage_opamp_dummy_magic_26_0.VD2.n29 two_stage_opamp_dummy_magic_26_0.VD2.n3 0.234875
R22606 two_stage_opamp_dummy_magic_26_0.VD2.n29 two_stage_opamp_dummy_magic_26_0.VD2.n28 0.234875
R22607 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP_NFET1.t0 141.653
R22608 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.t18 310.488
R22609 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t13 310.488
R22610 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t17 310.488
R22611 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n8 297.433
R22612 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n3 297.433
R22613 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.n14 297.433
R22614 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.t11 184.097
R22615 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.t9 184.097
R22616 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.t7 184.097
R22617 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.n11 167.094
R22618 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.n5 167.094
R22619 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.n0 167.094
R22620 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.n13 161.3
R22621 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n7 161.3
R22622 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n2 161.3
R22623 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.t14 120.501
R22624 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.t5 120.501
R22625 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t15 120.501
R22626 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.t3 120.501
R22627 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t16 120.501
R22628 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.t1 120.501
R22629 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.t0 50.2004
R22630 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.n12 40.7027
R22631 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.n6 40.7027
R22632 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.n1 40.7027
R22633 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t10 39.4005
R22634 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t4 39.4005
R22635 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t8 39.4005
R22636 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t2 39.4005
R22637 bgr_11_0.V_mir1.t12 bgr_11_0.V_mir1.n15 39.4005
R22638 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.t6 39.4005
R22639 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n4 6.6255
R22640 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.n10 6.6255
R22641 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n9 4.5005
R22642 VIN+.n0 VIN+.t10 1097.62
R22643 VIN+ VIN+.n9 433.019
R22644 VIN+.n9 VIN+.t5 273.134
R22645 VIN+.n0 VIN+.t7 273.134
R22646 VIN+.n8 VIN+.t1 273.134
R22647 VIN+.n7 VIN+.t4 273.134
R22648 VIN+.n6 VIN+.t0 273.134
R22649 VIN+.n5 VIN+.t3 273.134
R22650 VIN+.n4 VIN+.t8 273.134
R22651 VIN+.n3 VIN+.t6 273.134
R22652 VIN+.n2 VIN+.t9 273.134
R22653 VIN+.n1 VIN+.t2 273.134
R22654 VIN+.n1 VIN+.n0 176.733
R22655 VIN+.n2 VIN+.n1 176.733
R22656 VIN+.n3 VIN+.n2 176.733
R22657 VIN+.n4 VIN+.n3 176.733
R22658 VIN+.n5 VIN+.n4 176.733
R22659 VIN+.n6 VIN+.n5 176.733
R22660 VIN+.n7 VIN+.n6 176.733
R22661 VIN+.n8 VIN+.n7 176.733
R22662 VIN+.n9 VIN+.n8 176.733
R22663 two_stage_opamp_dummy_magic_26_0.V_err_gate.n2 two_stage_opamp_dummy_magic_26_0.V_err_gate.t8 479.322
R22664 two_stage_opamp_dummy_magic_26_0.V_err_gate.n2 two_stage_opamp_dummy_magic_26_0.V_err_gate.t6 479.322
R22665 two_stage_opamp_dummy_magic_26_0.V_err_gate.n6 two_stage_opamp_dummy_magic_26_0.V_err_gate.t7 479.322
R22666 two_stage_opamp_dummy_magic_26_0.V_err_gate.n6 two_stage_opamp_dummy_magic_26_0.V_err_gate.t9 479.322
R22667 two_stage_opamp_dummy_magic_26_0.V_err_gate.n3 two_stage_opamp_dummy_magic_26_0.V_err_gate.n1 178.075
R22668 two_stage_opamp_dummy_magic_26_0.V_err_gate.n5 two_stage_opamp_dummy_magic_26_0.V_err_gate.n4 177.434
R22669 two_stage_opamp_dummy_magic_26_0.V_err_gate two_stage_opamp_dummy_magic_26_0.V_err_gate.n0 170.357
R22670 two_stage_opamp_dummy_magic_26_0.V_err_gate.n3 two_stage_opamp_dummy_magic_26_0.V_err_gate.n2 165.8
R22671 two_stage_opamp_dummy_magic_26_0.V_err_gate two_stage_opamp_dummy_magic_26_0.V_err_gate.n6 165.8
R22672 two_stage_opamp_dummy_magic_26_0.V_err_gate.n0 two_stage_opamp_dummy_magic_26_0.V_err_gate.t2 24.0005
R22673 two_stage_opamp_dummy_magic_26_0.V_err_gate.n0 two_stage_opamp_dummy_magic_26_0.V_err_gate.t3 24.0005
R22674 two_stage_opamp_dummy_magic_26_0.V_err_gate.n4 two_stage_opamp_dummy_magic_26_0.V_err_gate.t4 15.7605
R22675 two_stage_opamp_dummy_magic_26_0.V_err_gate.n4 two_stage_opamp_dummy_magic_26_0.V_err_gate.t1 15.7605
R22676 two_stage_opamp_dummy_magic_26_0.V_err_gate.n1 two_stage_opamp_dummy_magic_26_0.V_err_gate.t0 15.7605
R22677 two_stage_opamp_dummy_magic_26_0.V_err_gate.n1 two_stage_opamp_dummy_magic_26_0.V_err_gate.t5 15.7605
R22678 two_stage_opamp_dummy_magic_26_0.V_err_gate two_stage_opamp_dummy_magic_26_0.V_err_gate.n5 1.76612
R22679 two_stage_opamp_dummy_magic_26_0.V_err_gate.n5 two_stage_opamp_dummy_magic_26_0.V_err_gate.n3 0.641125
R22680 two_stage_opamp_dummy_magic_26_0.V_err_mir_p two_stage_opamp_dummy_magic_26_0.V_err_mir_p.n0 186.762
R22681 two_stage_opamp_dummy_magic_26_0.V_err_mir_p two_stage_opamp_dummy_magic_26_0.V_err_mir_p.n1 177.201
R22682 two_stage_opamp_dummy_magic_26_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_26_0.V_err_mir_p.t1 15.7605
R22683 two_stage_opamp_dummy_magic_26_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_26_0.V_err_mir_p.t3 15.7605
R22684 two_stage_opamp_dummy_magic_26_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_26_0.V_err_mir_p.t2 15.7605
R22685 two_stage_opamp_dummy_magic_26_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_26_0.V_err_mir_p.t0 15.7605
R22686 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n0 345.264
R22687 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n1 344.7
R22688 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n3 292.5
R22689 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t10 121.931
R22690 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n7 118.861
R22691 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n9 118.861
R22692 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n13 118.861
R22693 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n16 118.861
R22694 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n19 118.861
R22695 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n22 74.1255
R22696 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n2 52.763
R22697 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n4 51.8547
R22698 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t13 39.4005
R22699 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t16 39.4005
R22700 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t12 39.4005
R22701 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t11 39.4005
R22702 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t15 39.4005
R22703 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t14 39.4005
R22704 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t5 19.7005
R22705 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t8 19.7005
R22706 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t2 19.7005
R22707 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t7 19.7005
R22708 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t1 19.7005
R22709 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t6 19.7005
R22710 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t4 19.7005
R22711 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t0 19.7005
R22712 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t3 19.7005
R22713 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t9 19.7005
R22714 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n21 5.90675
R22715 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n8 5.60467
R22716 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n18 5.54217
R22717 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n6 5.54217
R22718 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n10 5.04217
R22719 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n12 5.04217
R22720 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n5 5.04217
R22721 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n20 5.04217
R22722 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n6 4.97967
R22723 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n14 4.97967
R22724 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n17 4.97967
R22725 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n15 0.563
R22726 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n6 0.563
R22727 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n11 0.563
R22728 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n5 0.563
R22729 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n5 0.563
R22730 two_stage_opamp_dummy_magic_26_0.Vb2_2.n2 two_stage_opamp_dummy_magic_26_0.Vb2_2.t6 661.375
R22731 two_stage_opamp_dummy_magic_26_0.Vb2_2.n4 two_stage_opamp_dummy_magic_26_0.Vb2_2.t3 661.375
R22732 two_stage_opamp_dummy_magic_26_0.Vb2_2.t7 two_stage_opamp_dummy_magic_26_0.Vb2_2.n0 213.131
R22733 two_stage_opamp_dummy_magic_26_0.Vb2_2.n3 two_stage_opamp_dummy_magic_26_0.Vb2_2.t4 213.131
R22734 two_stage_opamp_dummy_magic_26_0.Vb2_2.n6 two_stage_opamp_dummy_magic_26_0.Vb2_2.n1 154.994
R22735 two_stage_opamp_dummy_magic_26_0.Vb2_2.t0 two_stage_opamp_dummy_magic_26_0.Vb2_2.t7 146.155
R22736 two_stage_opamp_dummy_magic_26_0.Vb2_2.t4 two_stage_opamp_dummy_magic_26_0.Vb2_2.t0 146.155
R22737 two_stage_opamp_dummy_magic_26_0.Vb2_2.t8 two_stage_opamp_dummy_magic_26_0.Vb2_2.n0 76.2576
R22738 two_stage_opamp_dummy_magic_26_0.Vb2_2.n3 two_stage_opamp_dummy_magic_26_0.Vb2_2.t5 76.2576
R22739 two_stage_opamp_dummy_magic_26_0.Vb2_2.n7 two_stage_opamp_dummy_magic_26_0.Vb2_2.n6 66.4414
R22740 two_stage_opamp_dummy_magic_26_0.Vb2_2.n1 two_stage_opamp_dummy_magic_26_0.Vb2_2.t9 21.8894
R22741 two_stage_opamp_dummy_magic_26_0.Vb2_2.n1 two_stage_opamp_dummy_magic_26_0.Vb2_2.t2 21.8894
R22742 two_stage_opamp_dummy_magic_26_0.Vb2_2.t8 two_stage_opamp_dummy_magic_26_0.Vb2_2.n7 11.2576
R22743 two_stage_opamp_dummy_magic_26_0.Vb2_2.n7 two_stage_opamp_dummy_magic_26_0.Vb2_2.t1 11.2576
R22744 two_stage_opamp_dummy_magic_26_0.Vb2_2.n5 two_stage_opamp_dummy_magic_26_0.Vb2_2.n4 5.1255
R22745 two_stage_opamp_dummy_magic_26_0.Vb2_2.n6 two_stage_opamp_dummy_magic_26_0.Vb2_2.n5 4.9214
R22746 two_stage_opamp_dummy_magic_26_0.Vb2_2.n5 two_stage_opamp_dummy_magic_26_0.Vb2_2.n2 4.7505
R22747 two_stage_opamp_dummy_magic_26_0.Vb2_2.n4 two_stage_opamp_dummy_magic_26_0.Vb2_2.n3 1.888
R22748 two_stage_opamp_dummy_magic_26_0.Vb2_2.n2 two_stage_opamp_dummy_magic_26_0.Vb2_2.n0 1.888
R22749 two_stage_opamp_dummy_magic_26_0.Vb3.n16 two_stage_opamp_dummy_magic_26_0.Vb3.t19 793.28
R22750 two_stage_opamp_dummy_magic_26_0.Vb3.n9 two_stage_opamp_dummy_magic_26_0.Vb3.t20 752.422
R22751 two_stage_opamp_dummy_magic_26_0.Vb3.n0 two_stage_opamp_dummy_magic_26_0.Vb3.t26 752.422
R22752 two_stage_opamp_dummy_magic_26_0.Vb3.n9 two_stage_opamp_dummy_magic_26_0.Vb3.t16 752.234
R22753 two_stage_opamp_dummy_magic_26_0.Vb3.n9 two_stage_opamp_dummy_magic_26_0.Vb3.t23 752.234
R22754 two_stage_opamp_dummy_magic_26_0.Vb3.n8 two_stage_opamp_dummy_magic_26_0.Vb3.t9 752.234
R22755 two_stage_opamp_dummy_magic_26_0.Vb3.n6 two_stage_opamp_dummy_magic_26_0.Vb3.t12 752.234
R22756 two_stage_opamp_dummy_magic_26_0.Vb3.n7 two_stage_opamp_dummy_magic_26_0.Vb3.t17 752.234
R22757 two_stage_opamp_dummy_magic_26_0.Vb3.n7 two_stage_opamp_dummy_magic_26_0.Vb3.t24 752.234
R22758 two_stage_opamp_dummy_magic_26_0.Vb3.n20 two_stage_opamp_dummy_magic_26_0.Vb3.t27 752.234
R22759 two_stage_opamp_dummy_magic_26_0.Vb3.n5 two_stage_opamp_dummy_magic_26_0.Vb3.t15 752.234
R22760 two_stage_opamp_dummy_magic_26_0.Vb3.n5 two_stage_opamp_dummy_magic_26_0.Vb3.t22 752.234
R22761 two_stage_opamp_dummy_magic_26_0.Vb3.n4 two_stage_opamp_dummy_magic_26_0.Vb3.t18 752.234
R22762 two_stage_opamp_dummy_magic_26_0.Vb3.n4 two_stage_opamp_dummy_magic_26_0.Vb3.t25 752.234
R22763 two_stage_opamp_dummy_magic_26_0.Vb3.n1 two_stage_opamp_dummy_magic_26_0.Vb3.t10 752.234
R22764 two_stage_opamp_dummy_magic_26_0.Vb3.n1 two_stage_opamp_dummy_magic_26_0.Vb3.t13 752.234
R22765 two_stage_opamp_dummy_magic_26_0.Vb3.n0 two_stage_opamp_dummy_magic_26_0.Vb3.t21 752.234
R22766 two_stage_opamp_dummy_magic_26_0.Vb3.n18 two_stage_opamp_dummy_magic_26_0.Vb3.t11 747.734
R22767 two_stage_opamp_dummy_magic_26_0.Vb3.n19 two_stage_opamp_dummy_magic_26_0.Vb3.t14 747.734
R22768 two_stage_opamp_dummy_magic_26_0.Vb3.n3 two_stage_opamp_dummy_magic_26_0.Vb3.t8 747.827
R22769 two_stage_opamp_dummy_magic_26_0.Vb3.n12 two_stage_opamp_dummy_magic_26_0.Vb3.n10 139.639
R22770 two_stage_opamp_dummy_magic_26_0.Vb3.n12 two_stage_opamp_dummy_magic_26_0.Vb3.n11 139.638
R22771 two_stage_opamp_dummy_magic_26_0.Vb3.n14 two_stage_opamp_dummy_magic_26_0.Vb3.n13 134.577
R22772 two_stage_opamp_dummy_magic_26_0.Vb3.n16 two_stage_opamp_dummy_magic_26_0.Vb3.n15 72.612
R22773 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_26_0.Vb3.n21 44.5943
R22774 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_26_0.Vb3.n14 43.0317
R22775 two_stage_opamp_dummy_magic_26_0.Vb3.n11 two_stage_opamp_dummy_magic_26_0.Vb3.t2 24.0005
R22776 two_stage_opamp_dummy_magic_26_0.Vb3.n11 two_stage_opamp_dummy_magic_26_0.Vb3.t3 24.0005
R22777 two_stage_opamp_dummy_magic_26_0.Vb3.n10 two_stage_opamp_dummy_magic_26_0.Vb3.t1 24.0005
R22778 two_stage_opamp_dummy_magic_26_0.Vb3.n10 two_stage_opamp_dummy_magic_26_0.Vb3.t4 24.0005
R22779 two_stage_opamp_dummy_magic_26_0.Vb3.n13 two_stage_opamp_dummy_magic_26_0.Vb3.t6 24.0005
R22780 two_stage_opamp_dummy_magic_26_0.Vb3.n13 two_stage_opamp_dummy_magic_26_0.Vb3.t5 24.0005
R22781 two_stage_opamp_dummy_magic_26_0.Vb3.n15 two_stage_opamp_dummy_magic_26_0.Vb3.t7 11.2576
R22782 two_stage_opamp_dummy_magic_26_0.Vb3.n15 two_stage_opamp_dummy_magic_26_0.Vb3.t0 11.2576
R22783 two_stage_opamp_dummy_magic_26_0.Vb3.n17 two_stage_opamp_dummy_magic_26_0.Vb3.n16 11.2036
R22784 two_stage_opamp_dummy_magic_26_0.Vb3.n21 two_stage_opamp_dummy_magic_26_0.Vb3.n17 6.14112
R22785 two_stage_opamp_dummy_magic_26_0.Vb3.n2 two_stage_opamp_dummy_magic_26_0.Vb3.n3 2.20508
R22786 two_stage_opamp_dummy_magic_26_0.Vb3.n6 two_stage_opamp_dummy_magic_26_0.Vb3.n19 4.5005
R22787 two_stage_opamp_dummy_magic_26_0.Vb3.n18 two_stage_opamp_dummy_magic_26_0.Vb3.n8 4.5005
R22788 two_stage_opamp_dummy_magic_26_0.Vb3.n14 two_stage_opamp_dummy_magic_26_0.Vb3.n12 4.5005
R22789 two_stage_opamp_dummy_magic_26_0.Vb3.n17 two_stage_opamp_dummy_magic_26_0.Vb3.n5 3.21925
R22790 two_stage_opamp_dummy_magic_26_0.Vb3.n21 two_stage_opamp_dummy_magic_26_0.Vb3.n20 0.641125
R22791 two_stage_opamp_dummy_magic_26_0.Vb3.n8 two_stage_opamp_dummy_magic_26_0.Vb3.n9 0.3755
R22792 two_stage_opamp_dummy_magic_26_0.Vb3.n6 two_stage_opamp_dummy_magic_26_0.Vb3.n8 0.3755
R22793 two_stage_opamp_dummy_magic_26_0.Vb3.n7 two_stage_opamp_dummy_magic_26_0.Vb3.n6 0.3755
R22794 two_stage_opamp_dummy_magic_26_0.Vb3.n20 two_stage_opamp_dummy_magic_26_0.Vb3.n7 0.3755
R22795 two_stage_opamp_dummy_magic_26_0.Vb3.n5 two_stage_opamp_dummy_magic_26_0.Vb3.n4 0.3755
R22796 two_stage_opamp_dummy_magic_26_0.Vb3.n4 two_stage_opamp_dummy_magic_26_0.Vb3.n2 0.3755
R22797 two_stage_opamp_dummy_magic_26_0.Vb3.n2 two_stage_opamp_dummy_magic_26_0.Vb3.n1 0.3755
R22798 two_stage_opamp_dummy_magic_26_0.Vb3.n19 two_stage_opamp_dummy_magic_26_0.Vb3.n18 0.188
R22799 two_stage_opamp_dummy_magic_26_0.Vb3.t28 two_stage_opamp_dummy_magic_26_0.Vb3.n3 747.827
R22800 two_stage_opamp_dummy_magic_26_0.Vb3.n1 two_stage_opamp_dummy_magic_26_0.Vb3.n0 0.3755
R22801 a_6350_30238.t0 a_6350_30238.t1 178.133
R22802 bgr_11_0.Vin+ bgr_11_0.Vin+.t6 529.879
R22803 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t0 148.653
R22804 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t1 125.418
R22805 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n1 106.609
R22806 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n2 104.484
R22807 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n0 25.0809
R22808 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n3 18.7817
R22809 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t4 13.1338
R22810 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t3 13.1338
R22811 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t2 13.1338
R22812 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t5 13.1338
R22813 bgr_11_0.Vin+ bgr_11_0.Vin+.n4 6.53175
R22814 a_6540_22450.n11 a_6540_22450.t18 310.488
R22815 a_6540_22450.n5 a_6540_22450.t13 310.488
R22816 a_6540_22450.n0 a_6540_22450.t14 310.488
R22817 a_6540_22450.n9 a_6540_22450.n8 297.433
R22818 a_6540_22450.n4 a_6540_22450.n3 297.433
R22819 a_6540_22450.n15 a_6540_22450.n14 297.433
R22820 a_6540_22450.n13 a_6540_22450.t7 184.097
R22821 a_6540_22450.n7 a_6540_22450.t5 184.097
R22822 a_6540_22450.n2 a_6540_22450.t3 184.097
R22823 a_6540_22450.n12 a_6540_22450.n11 167.094
R22824 a_6540_22450.n6 a_6540_22450.n5 167.094
R22825 a_6540_22450.n1 a_6540_22450.n0 167.094
R22826 a_6540_22450.n14 a_6540_22450.n13 161.3
R22827 a_6540_22450.n9 a_6540_22450.n7 161.3
R22828 a_6540_22450.n4 a_6540_22450.n2 161.3
R22829 a_6540_22450.n11 a_6540_22450.t15 120.501
R22830 a_6540_22450.n12 a_6540_22450.t11 120.501
R22831 a_6540_22450.n5 a_6540_22450.t17 120.501
R22832 a_6540_22450.n6 a_6540_22450.t1 120.501
R22833 a_6540_22450.n0 a_6540_22450.t16 120.501
R22834 a_6540_22450.n1 a_6540_22450.t9 120.501
R22835 a_6540_22450.n9 a_6540_22450.t0 50.2004
R22836 a_6540_22450.n13 a_6540_22450.n12 40.7027
R22837 a_6540_22450.n7 a_6540_22450.n6 40.7027
R22838 a_6540_22450.n2 a_6540_22450.n1 40.7027
R22839 a_6540_22450.n8 a_6540_22450.t2 39.4005
R22840 a_6540_22450.n8 a_6540_22450.t6 39.4005
R22841 a_6540_22450.n3 a_6540_22450.t10 39.4005
R22842 a_6540_22450.n3 a_6540_22450.t4 39.4005
R22843 a_6540_22450.t12 a_6540_22450.n15 39.4005
R22844 a_6540_22450.n15 a_6540_22450.t8 39.4005
R22845 a_6540_22450.n10 a_6540_22450.n4 6.6255
R22846 a_6540_22450.n14 a_6540_22450.n10 6.6255
R22847 a_6540_22450.n10 a_6540_22450.n9 4.5005
R22848 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t5 447.279
R22849 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t7 446.967
R22850 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t2 446.967
R22851 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t3 446.967
R22852 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t8 344.772
R22853 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n8 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t9 281.168
R22854 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t4 281.168
R22855 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t6 281.168
R22856 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n8 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n7 205.946
R22857 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n6 205.946
R22858 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n4 165.8
R22859 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n9 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n8 165.8
R22860 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t1 108.615
R22861 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n10 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t0 108.615
R22862 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n5 63.4857
R22863 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n4 51.5193
R22864 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n10 15.6567
R22865 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n3 10.5317
R22866 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n2 6.0005
R22867 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n10 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n9 6.0005
R22868 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n1 0.313
R22869 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n0 0.313
R22870 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n9 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n4 0.313
R22871 bgr_11_0.cap_res2.t0 bgr_11_0.cap_res2.t15 121.931
R22872 bgr_11_0.cap_res2.t10 bgr_11_0.cap_res2.t4 0.1603
R22873 bgr_11_0.cap_res2.t14 bgr_11_0.cap_res2.t9 0.1603
R22874 bgr_11_0.cap_res2.t8 bgr_11_0.cap_res2.t3 0.1603
R22875 bgr_11_0.cap_res2.t2 bgr_11_0.cap_res2.t16 0.1603
R22876 bgr_11_0.cap_res2.t6 bgr_11_0.cap_res2.t1 0.1603
R22877 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t11 0.159278
R22878 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t7 0.159278
R22879 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t13 0.159278
R22880 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t19 0.159278
R22881 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t20 0.1368
R22882 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t10 0.1368
R22883 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t5 0.1368
R22884 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t14 0.1368
R22885 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t18 0.1368
R22886 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t8 0.1368
R22887 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t12 0.1368
R22888 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t2 0.1368
R22889 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t17 0.1368
R22890 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t6 0.1368
R22891 bgr_11_0.cap_res2.t11 bgr_11_0.cap_res2.n0 0.00152174
R22892 bgr_11_0.cap_res2.t7 bgr_11_0.cap_res2.n1 0.00152174
R22893 bgr_11_0.cap_res2.t13 bgr_11_0.cap_res2.n2 0.00152174
R22894 bgr_11_0.cap_res2.t19 bgr_11_0.cap_res2.n3 0.00152174
R22895 bgr_11_0.cap_res2.t15 bgr_11_0.cap_res2.n4 0.00152174
R22896 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 172.969
R22897 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R22898 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R22899 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R22900 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R22901 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R22902 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R22903 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R22904 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R22905 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R22906 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R22907 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R22908 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R22909 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R22910 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R22911 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R22912 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R22913 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R22914 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R22915 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R22916 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R22917 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R22918 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R22919 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R22920 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R22921 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R22922 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R22923 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R22924 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R22925 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R22926 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R22927 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R22928 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R22929 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R22930 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R22931 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R22932 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R22933 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 65.0299
R22934 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 65.0299
R22935 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R22936 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R22937 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R22938 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R22939 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R22940 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R22941 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R22942 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R22943 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R22944 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R22945 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 25.7843
R22946 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R22947 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R22948 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R22949 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R22950 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R22951 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R22952 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R22953 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R22954 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R22955 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R22956 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R22957 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R22958 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R22959 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R22960 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R22961 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R22962 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R22963 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R22964 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R22965 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R22966 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R22967 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R22968 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R22969 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R22970 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R22971 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R22972 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R22973 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R22974 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R22975 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R22976 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R22977 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R22978 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R22979 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R22980 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R22981 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R22982 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R22983 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R22984 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R22985 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R22986 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R22987 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R22988 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R22989 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R22990 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R22991 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R22992 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R22993 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R22994 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R22995 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R22996 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R22997 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R22998 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R22999 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R23000 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R23001 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R23002 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R23003 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R23004 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R23005 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R23006 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R23007 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R23008 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R23009 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R23010 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R23011 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R23012 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R23013 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R23014 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R23015 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R23016 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R23017 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R23018 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R23019 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R23020 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R23021 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R23022 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R23023 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R23024 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R23025 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R23026 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R23027 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R23028 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R23029 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R23030 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R23031 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R23032 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R23033 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R23034 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R23035 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R23036 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R23037 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R23038 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R23039 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R23040 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R23041 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R23042 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R23043 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R23044 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R23045 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R23046 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R23047 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R23048 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R23049 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R23050 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R23051 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R23052 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R23053 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R23054 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R23055 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R23056 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R23057 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R23058 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R23059 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R23060 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R23061 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R23062 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R23063 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R23064 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R23065 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R23066 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R23067 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R23068 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R23069 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R23070 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R23071 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R23072 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R23073 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R23074 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R23075 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R23076 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R23077 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R23078 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R23079 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R23080 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R23081 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R23082 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R23083 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R23084 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R23085 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R23086 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R23087 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R23088 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R23089 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R23090 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R23091 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R23092 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R23093 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R23094 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R23095 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R23096 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R23097 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R23098 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R23099 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R23100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R23101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R23102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R23103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R23104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 0.290206
R23105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 0.290206
R23106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R23107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R23108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R23109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R23110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 0.290206
R23111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R23112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R23113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R23114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R23115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R23116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R23117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R23118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R23119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R23120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R23121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R23122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R23123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R23124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R23125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R23126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R23127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R23128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R23129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R23130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R23131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R23132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R23133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R23134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R23135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R23136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R23137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R23138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R23139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R23140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R23141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R23142 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R23143 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R23144 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R23145 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R23146 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R23147 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R23148 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R23149 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R23150 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R23151 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R23152 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R23153 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R23154 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R23155 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R23156 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R23157 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R23158 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R23159 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R23160 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R23161 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R23162 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R23163 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R23164 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R23165 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R23166 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R23167 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R23168 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R23169 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R23170 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t10 119.785
R23171 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n0 107.121
R23172 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n1 97.4332
R23173 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n20 68.5317
R23174 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n2 39.4067
R23175 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n5 24.288
R23176 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n7 24.288
R23177 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n11 24.288
R23178 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n14 24.288
R23179 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n17 24.288
R23180 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t11 24.0005
R23181 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t14 24.0005
R23182 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t13 24.0005
R23183 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t12 24.0005
R23184 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t0 8.0005
R23185 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t3 8.0005
R23186 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t7 8.0005
R23187 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t2 8.0005
R23188 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t6 8.0005
R23189 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t1 8.0005
R23190 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t9 8.0005
R23191 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t5 8.0005
R23192 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t8 8.0005
R23193 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t4 8.0005
R23194 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n16 5.7505
R23195 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n4 5.7505
R23196 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n6 5.7505
R23197 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n19 5.6255
R23198 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n8 5.188
R23199 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n4 5.188
R23200 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n10 5.188
R23201 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n12 5.188
R23202 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n3 5.188
R23203 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n15 5.188
R23204 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n18 5.188
R23205 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n13 0.563
R23206 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n4 0.563
R23207 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n9 0.563
R23208 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n3 0.563
R23209 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n3 0.563
R23210 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t1 119.785
R23211 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n0 107.121
R23212 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n1 97.4332
R23213 bgr_11_0.V_CMFB_S2 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n20 64.4067
R23214 bgr_11_0.V_CMFB_S2 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n2 30.9724
R23215 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n5 24.288
R23216 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n7 24.288
R23217 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n11 24.288
R23218 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n14 24.288
R23219 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n17 24.288
R23220 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t4 24.0005
R23221 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t0 24.0005
R23222 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t2 24.0005
R23223 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t3 24.0005
R23224 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t10 8.0005
R23225 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t5 8.0005
R23226 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t11 8.0005
R23227 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t6 8.0005
R23228 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t13 8.0005
R23229 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t7 8.0005
R23230 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t12 8.0005
R23231 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t9 8.0005
R23232 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t14 8.0005
R23233 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t8 8.0005
R23234 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n16 5.7505
R23235 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n4 5.7505
R23236 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n6 5.7505
R23237 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n19 5.6255
R23238 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n8 5.188
R23239 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n4 5.188
R23240 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n10 5.188
R23241 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n12 5.188
R23242 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n3 5.188
R23243 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n15 5.188
R23244 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n18 5.188
R23245 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n13 0.563
R23246 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n4 0.563
R23247 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n9 0.563
R23248 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n3 0.563
R23249 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n3 0.563
R23250 two_stage_opamp_dummy_magic_26_0.Vb1_2 two_stage_opamp_dummy_magic_26_0.Vb1_2.t0 74.8571
R23251 two_stage_opamp_dummy_magic_26_0.Vb1_2 two_stage_opamp_dummy_magic_26_0.Vb1_2.n0 54.689
R23252 two_stage_opamp_dummy_magic_26_0.Vb1_2 two_stage_opamp_dummy_magic_26_0.Vb1_2.n1 54.689
R23253 two_stage_opamp_dummy_magic_26_0.Vb1_2.n1 two_stage_opamp_dummy_magic_26_0.Vb1_2.t4 16.0005
R23254 two_stage_opamp_dummy_magic_26_0.Vb1_2.n1 two_stage_opamp_dummy_magic_26_0.Vb1_2.t2 16.0005
R23255 two_stage_opamp_dummy_magic_26_0.Vb1_2.n0 two_stage_opamp_dummy_magic_26_0.Vb1_2.t1 16.0005
R23256 two_stage_opamp_dummy_magic_26_0.Vb1_2.n0 two_stage_opamp_dummy_magic_26_0.Vb1_2.t3 16.0005
R23257 VIN-.n0 VIN-.t7 1097.62
R23258 VIN- VIN-.n9 433.019
R23259 VIN-.n9 VIN-.t10 273.134
R23260 VIN-.n0 VIN-.t9 273.134
R23261 VIN-.n1 VIN-.t3 273.134
R23262 VIN-.n2 VIN-.t8 273.134
R23263 VIN-.n3 VIN-.t1 273.134
R23264 VIN-.n4 VIN-.t5 273.134
R23265 VIN-.n5 VIN-.t2 273.134
R23266 VIN-.n6 VIN-.t6 273.134
R23267 VIN-.n7 VIN-.t0 273.134
R23268 VIN-.n8 VIN-.t4 273.134
R23269 VIN-.n9 VIN-.n8 176.733
R23270 VIN-.n8 VIN-.n7 176.733
R23271 VIN-.n7 VIN-.n6 176.733
R23272 VIN-.n6 VIN-.n5 176.733
R23273 VIN-.n5 VIN-.n4 176.733
R23274 VIN-.n4 VIN-.n3 176.733
R23275 VIN-.n3 VIN-.n2 176.733
R23276 VIN-.n2 VIN-.n1 176.733
R23277 VIN-.n1 VIN-.n0 176.733
R23278 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t6 661.375
R23279 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t3 661.375
R23280 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n6 213.131
R23281 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t7 213.131
R23282 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t4 146.155
R23283 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t0 146.155
R23284 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t5 76.2576
R23285 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t9 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n7 76.2576
R23286 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n1 72.4541
R23287 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n2 66.4525
R23288 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t1 11.2576
R23289 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t8 11.2576
R23290 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t2 11.2576
R23291 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t10 11.2576
R23292 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n4 5.1255
R23293 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n3 4.91035
R23294 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n0 4.7505
R23295 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n5 1.888
R23296 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n0 1.888
R23297 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t7 238.322
R23298 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t6 238.322
R23299 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n4 167.332
R23300 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t1 130.001
R23301 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n1 111.796
R23302 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n2 105.171
R23303 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t0 81.7074
R23304 bgr_11_0.START_UP bgr_11_0.START_UP.n0 36.8552
R23305 bgr_11_0.START_UP bgr_11_0.START_UP.n5 15.3755
R23306 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t2 13.1338
R23307 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t4 13.1338
R23308 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t3 13.1338
R23309 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t5 13.1338
R23310 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n3 4.21925
R23311 two_stage_opamp_dummy_magic_26_0.V_p_mir.n8 two_stage_opamp_dummy_magic_26_0.V_p_mir.n7 36.3346
R23312 two_stage_opamp_dummy_magic_26_0.V_p_mir.n6 two_stage_opamp_dummy_magic_26_0.V_p_mir.t0 16.0005
R23313 two_stage_opamp_dummy_magic_26_0.V_p_mir.n6 two_stage_opamp_dummy_magic_26_0.V_p_mir.t3 16.0005
R23314 two_stage_opamp_dummy_magic_26_0.V_p_mir.t2 two_stage_opamp_dummy_magic_26_0.V_p_mir.n8 9.6005
R23315 two_stage_opamp_dummy_magic_26_0.V_p_mir.n8 two_stage_opamp_dummy_magic_26_0.V_p_mir.t1 9.6005
R23316 two_stage_opamp_dummy_magic_26_0.V_p_mir.n7 two_stage_opamp_dummy_magic_26_0.V_p_mir.n0 2.24299
R23317 two_stage_opamp_dummy_magic_26_0.V_p_mir.n1 two_stage_opamp_dummy_magic_26_0.V_p_mir.n0 0.0273195
R23318 two_stage_opamp_dummy_magic_26_0.V_p_mir.n5 two_stage_opamp_dummy_magic_26_0.V_p_mir.n4 1.49085
R23319 two_stage_opamp_dummy_magic_26_0.V_p_mir.n1 two_stage_opamp_dummy_magic_26_0.V_p_mir.n3 0.913285
R23320 two_stage_opamp_dummy_magic_26_0.V_p_mir.n2 two_stage_opamp_dummy_magic_26_0.V_p_mir.n0 2.24321
R23321 two_stage_opamp_dummy_magic_26_0.V_p_mir.n7 two_stage_opamp_dummy_magic_26_0.V_p_mir.n4 0.0113462
R23322 two_stage_opamp_dummy_magic_26_0.V_p_mir.n5 two_stage_opamp_dummy_magic_26_0.V_p_mir.n3 1.13081
R23323 two_stage_opamp_dummy_magic_26_0.V_p_mir.n3 two_stage_opamp_dummy_magic_26_0.V_p_mir.n2 0.0253185
R23324 two_stage_opamp_dummy_magic_26_0.V_p_mir.n4 two_stage_opamp_dummy_magic_26_0.V_p_mir.n2 0.0378306
R23325 two_stage_opamp_dummy_magic_26_0.V_p_mir.n5 two_stage_opamp_dummy_magic_26_0.V_p_mir.n0 0.0326419
R23326 two_stage_opamp_dummy_magic_26_0.V_p_mir.n1 two_stage_opamp_dummy_magic_26_0.V_p_mir.n6 54.0327
R23327 a_11420_30238.t0 a_11420_30238.t1 178.133
R23328 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.t8 539.797
R23329 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.n6 351.865
R23330 bgr_11_0.Vin-.n18 bgr_11_0.Vin-.n17 141.667
R23331 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.t7 117.817
R23332 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.n3 109.204
R23333 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.n4 104.829
R23334 bgr_11_0.Vin-.n19 bgr_11_0.Vin-.n18 84.0884
R23335 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.n13 83.5719
R23336 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n0 83.5719
R23337 bgr_11_0.Vin-.n16 bgr_11_0.Vin-.n1 83.5719
R23338 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.t2 65.0299
R23339 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.t1 39.4005
R23340 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.t0 39.4005
R23341 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n14 26.074
R23342 bgr_11_0.Vin-.n16 bgr_11_0.Vin-.n15 26.074
R23343 bgr_11_0.Vin-.n18 bgr_11_0.Vin-.n16 26.074
R23344 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.n9 24.3755
R23345 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.n8 17.6255
R23346 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.t4 13.1338
R23347 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.t5 13.1338
R23348 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t6 13.1338
R23349 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t3 13.1338
R23350 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.n7 11.6567
R23351 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.n5 3.8755
R23352 bgr_11_0.Vin-.n20 bgr_11_0.Vin-.n19 1.56836
R23353 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n11 1.56363
R23354 bgr_11_0.Vin-.n21 bgr_11_0.Vin-.n20 1.5505
R23355 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n2 1.5505
R23356 bgr_11_0.Vin-.n19 bgr_11_0.Vin-.n1 1.14402
R23357 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n0 0.885803
R23358 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n12 0.77514
R23359 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n0 0.756696
R23360 bgr_11_0.Vin-.n21 bgr_11_0.Vin-.n1 0.701365
R23361 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.n10 0.530034
R23362 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.t2 0.290206
R23363 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n21 0.203382
R23364 bgr_11_0.Vin-.n20 bgr_11_0.Vin-.n2 0.0183571
R23365 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.n2 0.00817857
R23366 a_11950_28880.t0 a_11950_28880.t1 178.133
R23367 a_3810_3908.t0 a_3810_3908.t1 169.905
R23368 two_stage_opamp_dummy_magic_26_0.V_tot.n2 two_stage_opamp_dummy_magic_26_0.V_tot.t5 648.343
R23369 two_stage_opamp_dummy_magic_26_0.V_tot.n1 two_stage_opamp_dummy_magic_26_0.V_tot.t4 648.343
R23370 two_stage_opamp_dummy_magic_26_0.V_tot.n3 two_stage_opamp_dummy_magic_26_0.V_tot.t1 117.591
R23371 two_stage_opamp_dummy_magic_26_0.V_tot.n0 two_stage_opamp_dummy_magic_26_0.V_tot.t3 117.591
R23372 two_stage_opamp_dummy_magic_26_0.V_tot.n0 two_stage_opamp_dummy_magic_26_0.V_tot.t2 108.424
R23373 two_stage_opamp_dummy_magic_26_0.V_tot.t0 two_stage_opamp_dummy_magic_26_0.V_tot.n3 108.424
R23374 two_stage_opamp_dummy_magic_26_0.V_tot.n3 two_stage_opamp_dummy_magic_26_0.V_tot.n2 46.5809
R23375 two_stage_opamp_dummy_magic_26_0.V_tot.n1 two_stage_opamp_dummy_magic_26_0.V_tot.n0 46.5184
R23376 two_stage_opamp_dummy_magic_26_0.V_tot.n2 two_stage_opamp_dummy_magic_26_0.V_tot.n1 1.563
R23377 a_13840_3908.t0 a_13840_3908.t1 294.339
R23378 two_stage_opamp_dummy_magic_26_0.err_amp_out.n0 two_stage_opamp_dummy_magic_26_0.err_amp_out.t4 610.534
R23379 two_stage_opamp_dummy_magic_26_0.err_amp_out.n0 two_stage_opamp_dummy_magic_26_0.err_amp_out.t5 433.8
R23380 two_stage_opamp_dummy_magic_26_0.err_amp_out.n2 two_stage_opamp_dummy_magic_26_0.err_amp_out.n0 278.06
R23381 two_stage_opamp_dummy_magic_26_0.err_amp_out.n2 two_stage_opamp_dummy_magic_26_0.err_amp_out.n1 178.829
R23382 two_stage_opamp_dummy_magic_26_0.err_amp_out.n3 two_stage_opamp_dummy_magic_26_0.err_amp_out.n2 39.3422
R23383 two_stage_opamp_dummy_magic_26_0.err_amp_out.n1 two_stage_opamp_dummy_magic_26_0.err_amp_out.t3 15.7605
R23384 two_stage_opamp_dummy_magic_26_0.err_amp_out.n1 two_stage_opamp_dummy_magic_26_0.err_amp_out.t0 15.7605
R23385 two_stage_opamp_dummy_magic_26_0.err_amp_out.t1 two_stage_opamp_dummy_magic_26_0.err_amp_out.n3 9.6005
R23386 two_stage_opamp_dummy_magic_26_0.err_amp_out.n3 two_stage_opamp_dummy_magic_26_0.err_amp_out.t2 9.6005
R23387 two_stage_opamp_dummy_magic_26_0.V_err_p.n1 two_stage_opamp_dummy_magic_26_0.V_err_p.n0 363.962
R23388 two_stage_opamp_dummy_magic_26_0.V_err_p.n0 two_stage_opamp_dummy_magic_26_0.V_err_p.t3 15.7605
R23389 two_stage_opamp_dummy_magic_26_0.V_err_p.n0 two_stage_opamp_dummy_magic_26_0.V_err_p.t1 15.7605
R23390 two_stage_opamp_dummy_magic_26_0.V_err_p.n1 two_stage_opamp_dummy_magic_26_0.V_err_p.t0 15.7605
R23391 two_stage_opamp_dummy_magic_26_0.V_err_p.t2 two_stage_opamp_dummy_magic_26_0.V_err_p.n1 15.7605
R23392 a_3690_3908.t0 a_3690_3908.t1 294.339
R23393 a_11300_28630.t0 a_11300_28630.t1 178.133
R23394 a_13960_3908.t0 a_13960_3908.t1 169.905
R23395 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t2 99.8322
R23396 bgr_11_0.V_p_1.t0 bgr_11_0.V_p_1.n0 9.6005
R23397 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t1 9.6005
R23398 a_13940_106.t0 a_13940_106.t1 169.905
R23399 a_5700_30088.t0 a_5700_30088.t1 178.133
R23400 a_5820_28824.t0 a_5820_28824.t1 178.133
R23401 a_3830_106.t0 a_3830_106.t1 169.905
R23402 a_6470_28630.t0 a_6470_28630.t1 178.133
R23403 a_12070_30088.t0 a_12070_30088.t1 178.133
R23404 bgr_11_0.V_CUR_REF_REG bgr_11_0.V_CUR_REF_REG.t3 701.501
R23405 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.n0 357.647
R23406 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.t0 135.239
R23407 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t1 39.4005
R23408 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t2 39.4005
R23409 bgr_11_0.V_CUR_REF_REG bgr_11_0.V_CUR_REF_REG.n1 5.79738
R23410 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t2 142.558
R23411 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t1 9.6005
R23412 bgr_11_0.V_p_2.t0 bgr_11_0.V_p_2.n0 9.6005
C0 bgr_11_0.Vin+ bgr_11_0.1st_Vout_1 0.275724f
C1 two_stage_opamp_dummy_magic_26_0.V_tail_gate two_stage_opamp_dummy_magic_26_0.Y 0.031497f
C2 two_stage_opamp_dummy_magic_26_0.Y VOUT+ 3.93988f
C3 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP 0.145663f
C4 two_stage_opamp_dummy_magic_26_0.cap_res_X two_stage_opamp_dummy_magic_26_0.V_source 0.069737f
C5 bgr_11_0.START_UP VDDA 2.28936f
C6 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref two_stage_opamp_dummy_magic_26_0.cap_res_Y 0.143247f
C7 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage 0.157302f
C8 two_stage_opamp_dummy_magic_26_0.V_tail_gate VOUT+ 1.3695f
C9 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_26_0.V_tail_gate 0.403953f
C10 bgr_11_0.V_TOP bgr_11_0.1st_Vout_1 2.6266f
C11 two_stage_opamp_dummy_magic_26_0.Y two_stage_opamp_dummy_magic_26_0.cap_res_Y 0.06758f
C12 two_stage_opamp_dummy_magic_26_0.V_tail_gate VOUT- 1.37075f
C13 VOUT+ VOUT- 0.213277f
C14 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref VDDA 6.26984f
C15 two_stage_opamp_dummy_magic_26_0.Y two_stage_opamp_dummy_magic_26_0.X 0.097316f
C16 two_stage_opamp_dummy_magic_26_0.V_err_gate bgr_11_0.1st_Vout_1 0.134861f
C17 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_26_0.V_err_amp_ref 0.808133f
C18 two_stage_opamp_dummy_magic_26_0.Y two_stage_opamp_dummy_magic_26_0.VD2 4.14841f
C19 bgr_11_0.Vin+ bgr_11_0.V_TOP 1.8967f
C20 two_stage_opamp_dummy_magic_26_0.V_tail_gate two_stage_opamp_dummy_magic_26_0.cap_res_Y 2.01462f
C21 two_stage_opamp_dummy_magic_26_0.cap_res_Y VOUT+ 51.1048f
C22 two_stage_opamp_dummy_magic_26_0.V_tail_gate two_stage_opamp_dummy_magic_26_0.VD1 0.01191f
C23 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.cap_res_X 0.185404f
C24 bgr_11_0.Vin+ bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 1.06291f
C25 two_stage_opamp_dummy_magic_26_0.V_err_mir_p VDDA 0.661231f
C26 two_stage_opamp_dummy_magic_26_0.V_tail_gate two_stage_opamp_dummy_magic_26_0.X 0.031497f
C27 two_stage_opamp_dummy_magic_26_0.V_tail_gate two_stage_opamp_dummy_magic_26_0.VD2 0.01191f
C28 bgr_11_0.START_UP bgr_11_0.1st_Vout_1 0.13011f
C29 two_stage_opamp_dummy_magic_26_0.V_tail_gate VIN+ 0.04837f
C30 two_stage_opamp_dummy_magic_26_0.VD4 two_stage_opamp_dummy_magic_26_0.Y 7.95637f
C31 two_stage_opamp_dummy_magic_26_0.V_err_gate two_stage_opamp_dummy_magic_26_0.Vb1 2.4413f
C32 bgr_11_0.Vin+ two_stage_opamp_dummy_magic_26_0.V_err_gate 0.066808f
C33 two_stage_opamp_dummy_magic_26_0.Y VDDA 7.52341f
C34 two_stage_opamp_dummy_magic_26_0.cap_res_Y VOUT- 0.02055f
C35 two_stage_opamp_dummy_magic_26_0.VD4 VOUT+ 0.034338f
C36 two_stage_opamp_dummy_magic_26_0.X VOUT- 3.93988f
C37 two_stage_opamp_dummy_magic_26_0.V_tail_gate VDDA 8.026971f
C38 VDDA VOUT+ 15.0814f
C39 bgr_11_0.V_CUR_REF_REG VDDA 3.77153f
C40 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_26_0.V_tail_gate 0.582654f
C41 bgr_11_0.Vin+ bgr_11_0.START_UP 0.170134f
C42 two_stage_opamp_dummy_magic_26_0.V_tail_gate VIN- 0.04837f
C43 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.V_TOP 0.04106f
C44 bgr_11_0.PFET_GATE_10uA bgr_11_0.V_CUR_REF_REG 0.347737f
C45 two_stage_opamp_dummy_magic_26_0.VD3 VOUT- 0.027349f
C46 two_stage_opamp_dummy_magic_26_0.X two_stage_opamp_dummy_magic_26_0.VD1 4.14841f
C47 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_26_0.V_err_gate 0.104556f
C48 two_stage_opamp_dummy_magic_26_0.VD2 two_stage_opamp_dummy_magic_26_0.VD1 0.024929f
C49 VDDA VOUT- 15.089801f
C50 two_stage_opamp_dummy_magic_26_0.V_tail_gate two_stage_opamp_dummy_magic_26_0.V_source 3.23984f
C51 two_stage_opamp_dummy_magic_26_0.VD2 VIN+ 0.533699f
C52 two_stage_opamp_dummy_magic_26_0.V_err_gate two_stage_opamp_dummy_magic_26_0.cap_res_X 0.161526f
C53 two_stage_opamp_dummy_magic_26_0.V_source VOUT+ 0.052413f
C54 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref two_stage_opamp_dummy_magic_26_0.Vb1 2.49082f
C55 two_stage_opamp_dummy_magic_26_0.VD3 two_stage_opamp_dummy_magic_26_0.X 7.95637f
C56 two_stage_opamp_dummy_magic_26_0.VD4 two_stage_opamp_dummy_magic_26_0.cap_res_Y 0.168036f
C57 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref bgr_11_0.Vin+ 0.25235f
C58 bgr_11_0.V_TOP bgr_11_0.START_UP 1.37378f
C59 two_stage_opamp_dummy_magic_26_0.cap_res_Y VDDA 7.24871f
C60 two_stage_opamp_dummy_magic_26_0.VD1 VIN- 0.533699f
C61 two_stage_opamp_dummy_magic_26_0.X VDDA 7.53665f
C62 two_stage_opamp_dummy_magic_26_0.V_source VOUT- 0.054425f
C63 VIN+ VIN- 0.075694f
C64 two_stage_opamp_dummy_magic_26_0.V_err_gate bgr_11_0.START_UP 0.743841f
C65 two_stage_opamp_dummy_magic_26_0.VD3 VDDA 8.707911f
C66 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.Y 3.11678f
C67 bgr_11_0.START_UP_NFET1 VDDA 0.18791f
C68 two_stage_opamp_dummy_magic_26_0.cap_res_Y two_stage_opamp_dummy_magic_26_0.V_source 0.062141f
C69 bgr_11_0.PFET_GATE_10uA bgr_11_0.START_UP_NFET1 0.010791f
C70 two_stage_opamp_dummy_magic_26_0.VD4 VDDA 8.70788f
C71 two_stage_opamp_dummy_magic_26_0.VD1 two_stage_opamp_dummy_magic_26_0.V_source 5.034379f
C72 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref bgr_11_0.V_TOP 0.939477f
C73 two_stage_opamp_dummy_magic_26_0.VD2 two_stage_opamp_dummy_magic_26_0.V_source 5.034379f
C74 bgr_11_0.PFET_GATE_10uA VDDA 10.121f
C75 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.V_tail_gate 3.67457f
C76 two_stage_opamp_dummy_magic_26_0.Vb1 VOUT+ 0.066228f
C77 two_stage_opamp_dummy_magic_26_0.V_tail_gate two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage 5.9387f
C78 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage VOUT+ 4.74661f
C79 two_stage_opamp_dummy_magic_26_0.V_source VIN+ 0.52651f
C80 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_26_0.Vb1 0.051702f
C81 bgr_11_0.Vin+ two_stage_opamp_dummy_magic_26_0.V_tail_gate 0.014649f
C82 bgr_11_0.Vin+ bgr_11_0.V_CUR_REF_REG 1.57077f
C83 two_stage_opamp_dummy_magic_26_0.V_source two_stage_opamp_dummy_magic_26_0.Vb1_2 0.143523f
C84 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref two_stage_opamp_dummy_magic_26_0.V_err_gate 0.804531f
C85 two_stage_opamp_dummy_magic_26_0.Vb1 VOUT- 0.04853f
C86 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage VOUT- 4.720799f
C87 two_stage_opamp_dummy_magic_26_0.V_source VIN- 0.52651f
C88 two_stage_opamp_dummy_magic_26_0.V_err_gate two_stage_opamp_dummy_magic_26_0.V_err_mir_p 0.429395f
C89 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref bgr_11_0.START_UP 1.39993f
C90 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_26_0.V_tail_gate 0.028061f
C91 bgr_11_0.V_CUR_REF_REG bgr_11_0.V_TOP 0.308375f
C92 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.cap_res_Y 0.23639f
C93 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.VD1 0.560747f
C94 two_stage_opamp_dummy_magic_26_0.V_tail_gate two_stage_opamp_dummy_magic_26_0.cap_res_X 2.01375f
C95 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.X 3.10888f
C96 two_stage_opamp_dummy_magic_26_0.cap_res_X VOUT+ 0.02055f
C97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.V_CUR_REF_REG 0.779503f
C98 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.VD2 0.561266f
C99 bgr_11_0.1st_Vout_1 VDDA 2.67125f
C100 two_stage_opamp_dummy_magic_26_0.V_err_gate two_stage_opamp_dummy_magic_26_0.V_tail_gate 0.124028f
C101 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.Vb1_2 2.01461f
C102 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_26_0.V_err_gate 0.375039f
C103 two_stage_opamp_dummy_magic_26_0.cap_res_X VOUT- 51.0064f
C104 two_stage_opamp_dummy_magic_26_0.Vb1 VDDA 12.443901f
C105 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage VDDA 0.015355f
C106 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_26_0.Vb1 0.091782f
C107 bgr_11_0.Vin+ VDDA 1.72765f
C108 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref two_stage_opamp_dummy_magic_26_0.V_err_mir_p 0.047283f
C109 two_stage_opamp_dummy_magic_26_0.V_err_gate VOUT- 0.022499f
C110 two_stage_opamp_dummy_magic_26_0.cap_res_Y two_stage_opamp_dummy_magic_26_0.cap_res_X 0.477735f
C111 two_stage_opamp_dummy_magic_26_0.X two_stage_opamp_dummy_magic_26_0.cap_res_X 0.06758f
C112 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref two_stage_opamp_dummy_magic_26_0.Y 0.051178f
C113 two_stage_opamp_dummy_magic_26_0.Vb1 two_stage_opamp_dummy_magic_26_0.V_source 1.01323f
C114 two_stage_opamp_dummy_magic_26_0.V_source two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage 1.19158f
C115 two_stage_opamp_dummy_magic_26_0.VD3 two_stage_opamp_dummy_magic_26_0.cap_res_X 0.167874f
C116 bgr_11_0.V_TOP VDDA 16.3436f
C117 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref two_stage_opamp_dummy_magic_26_0.V_tail_gate 0.130865f
C118 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref VOUT+ 0.022455f
C119 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref bgr_11_0.V_CUR_REF_REG 2.48242f
C120 bgr_11_0.PFET_GATE_10uA bgr_11_0.V_TOP 0.198568f
C121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter VDDA 0.023423f
C122 two_stage_opamp_dummy_magic_26_0.cap_res_X VDDA 7.27094f
C123 two_stage_opamp_dummy_magic_26_0.V_err_gate VDDA 2.4908f
C124 VIN- GNDA 1.83462f
C125 VIN+ GNDA 1.91203f
C126 VOUT- GNDA 25.749157f
C127 VOUT+ GNDA 25.751154f
C128 VDDA GNDA 0.37242p
C129 two_stage_opamp_dummy_magic_26_0.Vb1_2 GNDA 2.64849f
C130 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage GNDA 10.040009f
C131 two_stage_opamp_dummy_magic_26_0.V_source GNDA 26.762749f
C132 two_stage_opamp_dummy_magic_26_0.VD1 GNDA 3.421288f
C133 two_stage_opamp_dummy_magic_26_0.VD2 GNDA 3.585048f
C134 two_stage_opamp_dummy_magic_26_0.cap_res_X GNDA 41.339092f
C135 two_stage_opamp_dummy_magic_26_0.cap_res_Y GNDA 41.325703f
C136 two_stage_opamp_dummy_magic_26_0.X GNDA 11.94217f
C137 two_stage_opamp_dummy_magic_26_0.V_err_mir_p GNDA 0.118015f
C138 two_stage_opamp_dummy_magic_26_0.Y GNDA 12.05367f
C139 two_stage_opamp_dummy_magic_26_0.V_tail_gate GNDA 31.59499f
C140 two_stage_opamp_dummy_magic_26_0.Vb1 GNDA 35.87373f
C141 bgr_11_0.1st_Vout_1 GNDA 12.039672f
C142 bgr_11_0.START_UP GNDA 6.621171f
C143 bgr_11_0.START_UP_NFET1 GNDA 5.23862f
C144 two_stage_opamp_dummy_magic_26_0.V_err_gate GNDA 12.120259f
C145 bgr_11_0.V_TOP GNDA 11.594524f
C146 bgr_11_0.V_CUR_REF_REG GNDA 4.878339f
C147 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 16.8453f
C148 bgr_11_0.Vin+ GNDA 4.647517f
C149 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref GNDA 10.83651f
C150 bgr_11_0.PFET_GATE_10uA GNDA 8.898517f
C151 two_stage_opamp_dummy_magic_26_0.VD3 GNDA 5.849802f
C152 two_stage_opamp_dummy_magic_26_0.VD4 GNDA 5.854362f
C153 bgr_11_0.V_CUR_REF_REG.t3 GNDA 0.066747f
C154 bgr_11_0.V_CUR_REF_REG.t0 GNDA 0.452298f
C155 bgr_11_0.V_CUR_REF_REG.t1 GNDA 0.013056f
C156 bgr_11_0.V_CUR_REF_REG.t2 GNDA 0.013056f
C157 bgr_11_0.V_CUR_REF_REG.n0 GNDA 0.100023f
C158 bgr_11_0.V_CUR_REF_REG.n1 GNDA 5.13907f
C159 two_stage_opamp_dummy_magic_26_0.err_amp_out.t2 GNDA 0.079082f
C160 two_stage_opamp_dummy_magic_26_0.err_amp_out.t5 GNDA 0.084222f
C161 two_stage_opamp_dummy_magic_26_0.err_amp_out.t4 GNDA 0.098301f
C162 two_stage_opamp_dummy_magic_26_0.err_amp_out.n0 GNDA 0.325914f
C163 two_stage_opamp_dummy_magic_26_0.err_amp_out.t3 GNDA 0.079082f
C164 two_stage_opamp_dummy_magic_26_0.err_amp_out.t0 GNDA 0.079082f
C165 two_stage_opamp_dummy_magic_26_0.err_amp_out.n1 GNDA 0.256269f
C166 two_stage_opamp_dummy_magic_26_0.err_amp_out.n2 GNDA 3.75447f
C167 two_stage_opamp_dummy_magic_26_0.err_amp_out.n3 GNDA 0.264493f
C168 two_stage_opamp_dummy_magic_26_0.err_amp_out.t1 GNDA 0.079082f
C169 two_stage_opamp_dummy_magic_26_0.V_tot.t1 GNDA 0.289866f
C170 two_stage_opamp_dummy_magic_26_0.V_tot.t3 GNDA 0.289866f
C171 two_stage_opamp_dummy_magic_26_0.V_tot.t2 GNDA 0.272113f
C172 two_stage_opamp_dummy_magic_26_0.V_tot.n0 GNDA 1.77089f
C173 two_stage_opamp_dummy_magic_26_0.V_tot.t4 GNDA 0.08245f
C174 two_stage_opamp_dummy_magic_26_0.V_tot.n1 GNDA 1.68226f
C175 two_stage_opamp_dummy_magic_26_0.V_tot.t5 GNDA 0.08245f
C176 two_stage_opamp_dummy_magic_26_0.V_tot.n2 GNDA 1.68519f
C177 two_stage_opamp_dummy_magic_26_0.V_tot.n3 GNDA 1.7728f
C178 two_stage_opamp_dummy_magic_26_0.V_tot.t0 GNDA 0.272113f
C179 bgr_11_0.Vin-.n0 GNDA 0.07858f
C180 bgr_11_0.Vin-.n1 GNDA 0.088293f
C181 bgr_11_0.Vin-.n2 GNDA 0.12735f
C182 bgr_11_0.Vin-.t2 GNDA 0.294736f
C183 bgr_11_0.Vin-.t6 GNDA 0.030534f
C184 bgr_11_0.Vin-.t3 GNDA 0.030534f
C185 bgr_11_0.Vin-.n3 GNDA 0.085799f
C186 bgr_11_0.Vin-.t4 GNDA 0.030534f
C187 bgr_11_0.Vin-.t5 GNDA 0.030534f
C188 bgr_11_0.Vin-.n4 GNDA 0.074088f
C189 bgr_11_0.Vin-.n5 GNDA 0.633984f
C190 bgr_11_0.Vin-.t1 GNDA 0.010178f
C191 bgr_11_0.Vin-.t0 GNDA 0.010178f
C192 bgr_11_0.Vin-.n6 GNDA 0.031534f
C193 bgr_11_0.Vin-.n7 GNDA 0.428495f
C194 bgr_11_0.Vin-.t8 GNDA 0.049457f
C195 bgr_11_0.Vin-.n8 GNDA 0.623119f
C196 bgr_11_0.Vin-.t7 GNDA 0.128901f
C197 bgr_11_0.Vin-.n9 GNDA 0.734405f
C198 bgr_11_0.Vin-.n10 GNDA 1.36082f
C199 bgr_11_0.Vin-.n11 GNDA 0.531118f
C200 bgr_11_0.Vin-.n12 GNDA 0.079463f
C201 bgr_11_0.Vin-.n13 GNDA 0.13464f
C202 bgr_11_0.Vin-.n14 GNDA 0.078726f
C203 bgr_11_0.Vin-.n15 GNDA 0.155721f
C204 bgr_11_0.Vin-.n16 GNDA 0.155721f
C205 bgr_11_0.Vin-.n17 GNDA -0.303656f
C206 bgr_11_0.Vin-.n18 GNDA 0.501878f
C207 bgr_11_0.Vin-.n19 GNDA 0.240599f
C208 bgr_11_0.Vin-.n20 GNDA 0.454563f
C209 bgr_11_0.Vin-.n21 GNDA 0.043263f
C210 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.045912f
C211 two_stage_opamp_dummy_magic_26_0.V_p_mir.n0 GNDA 0.041422f
C212 two_stage_opamp_dummy_magic_26_0.V_p_mir.n1 GNDA 3.34407f
C213 two_stage_opamp_dummy_magic_26_0.V_p_mir.n2 GNDA 0.083146f
C214 two_stage_opamp_dummy_magic_26_0.V_p_mir.n3 GNDA 0.040904f
C215 two_stage_opamp_dummy_magic_26_0.V_p_mir.n5 GNDA 0.08194f
C216 two_stage_opamp_dummy_magic_26_0.V_p_mir.t1 GNDA 0.01618f
C217 two_stage_opamp_dummy_magic_26_0.V_p_mir.n6 GNDA 0.109281f
C218 two_stage_opamp_dummy_magic_26_0.V_p_mir.n7 GNDA 1.86634f
C219 two_stage_opamp_dummy_magic_26_0.V_p_mir.n8 GNDA 0.081126f
C220 two_stage_opamp_dummy_magic_26_0.V_p_mir.t2 GNDA 0.01618f
C221 bgr_11_0.START_UP.t0 GNDA 1.72724f
C222 bgr_11_0.START_UP.t1 GNDA 0.045404f
C223 bgr_11_0.START_UP.n0 GNDA 1.15615f
C224 bgr_11_0.START_UP.t2 GNDA 0.04333f
C225 bgr_11_0.START_UP.t4 GNDA 0.04333f
C226 bgr_11_0.START_UP.n1 GNDA 0.135247f
C227 bgr_11_0.START_UP.t3 GNDA 0.04333f
C228 bgr_11_0.START_UP.t5 GNDA 0.04333f
C229 bgr_11_0.START_UP.n2 GNDA 0.106737f
C230 bgr_11_0.START_UP.n3 GNDA 1.0283f
C231 bgr_11_0.START_UP.t6 GNDA 0.016282f
C232 bgr_11_0.START_UP.t7 GNDA 0.016282f
C233 bgr_11_0.START_UP.n4 GNDA 0.046713f
C234 bgr_11_0.START_UP.n5 GNDA 0.477587f
C235 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t6 GNDA 0.03776f
C236 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n0 GNDA 0.079757f
C237 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t5 GNDA 0.075848f
C238 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t3 GNDA 0.03776f
C239 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t2 GNDA 0.021323f
C240 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t10 GNDA 0.021323f
C241 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n1 GNDA 0.065225f
C242 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t1 GNDA 0.021323f
C243 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t8 GNDA 0.021323f
C244 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n2 GNDA 0.044611f
C245 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n3 GNDA 0.477605f
C246 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n4 GNDA 0.048057f
C247 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n5 GNDA 0.080962f
C248 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n6 GNDA 0.242604f
C249 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t4 GNDA 0.181754f
C250 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t0 GNDA 0.142559f
C251 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t7 GNDA 0.181754f
C252 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.n7 GNDA 0.242604f
C253 two_stage_opamp_dummy_magic_26_0.Vb2_Vb3.t9 GNDA 0.075848f
C254 two_stage_opamp_dummy_magic_26_0.Vb1_2.t1 GNDA 0.029732f
C255 two_stage_opamp_dummy_magic_26_0.Vb1_2.t3 GNDA 0.029732f
C256 two_stage_opamp_dummy_magic_26_0.Vb1_2.n0 GNDA 0.087151f
C257 two_stage_opamp_dummy_magic_26_0.Vb1_2.t0 GNDA 0.189479f
C258 two_stage_opamp_dummy_magic_26_0.Vb1_2.t4 GNDA 0.029732f
C259 two_stage_opamp_dummy_magic_26_0.Vb1_2.t2 GNDA 0.029732f
C260 two_stage_opamp_dummy_magic_26_0.Vb1_2.n1 GNDA 0.086354f
C261 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t4 GNDA 0.028726f
C262 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t0 GNDA 0.028726f
C263 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n0 GNDA 0.090339f
C264 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t2 GNDA 0.028726f
C265 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t3 GNDA 0.028726f
C266 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n1 GNDA 0.06162f
C267 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n2 GNDA 2.72441f
C268 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t1 GNDA 0.352049f
C269 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n3 GNDA 0.099919f
C270 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n4 GNDA 0.171922f
C271 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t10 GNDA 0.086179f
C272 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t5 GNDA 0.086179f
C273 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n5 GNDA 0.184319f
C274 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n6 GNDA 0.57655f
C275 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t11 GNDA 0.086179f
C276 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t6 GNDA 0.086179f
C277 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n7 GNDA 0.184319f
C278 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n8 GNDA 0.560935f
C279 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n9 GNDA 0.171922f
C280 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n10 GNDA 0.099919f
C281 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t13 GNDA 0.086179f
C282 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t7 GNDA 0.086179f
C283 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n11 GNDA 0.184319f
C284 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n12 GNDA 0.560935f
C285 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n13 GNDA 0.099919f
C286 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t12 GNDA 0.086179f
C287 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t9 GNDA 0.086179f
C288 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n14 GNDA 0.184319f
C289 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n15 GNDA 0.560935f
C290 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n16 GNDA 0.171922f
C291 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t14 GNDA 0.086179f
C292 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.t8 GNDA 0.086179f
C293 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n17 GNDA 0.184319f
C294 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n18 GNDA 0.568743f
C295 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n19 GNDA 0.199311f
C296 two_stage_opamp_dummy_magic_26_0.V_CMFB_S2.n20 GNDA 2.93837f
C297 bgr_11_0.V_CMFB_S2 GNDA 5.592f
C298 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t11 GNDA 0.027303f
C299 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t14 GNDA 0.027303f
C300 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n0 GNDA 0.085864f
C301 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t13 GNDA 0.027303f
C302 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t12 GNDA 0.027303f
C303 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n1 GNDA 0.058568f
C304 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n2 GNDA 1.80711f
C305 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t10 GNDA 0.334608f
C306 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n3 GNDA 0.094969f
C307 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n4 GNDA 0.163405f
C308 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t0 GNDA 0.081909f
C309 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t3 GNDA 0.081909f
C310 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n5 GNDA 0.175188f
C311 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n6 GNDA 0.547989f
C312 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t7 GNDA 0.081909f
C313 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t2 GNDA 0.081909f
C314 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n7 GNDA 0.175188f
C315 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n8 GNDA 0.533147f
C316 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n9 GNDA 0.163405f
C317 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n10 GNDA 0.094969f
C318 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t6 GNDA 0.081909f
C319 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t1 GNDA 0.081909f
C320 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n11 GNDA 0.175188f
C321 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n12 GNDA 0.533147f
C322 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n13 GNDA 0.094969f
C323 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t9 GNDA 0.081909f
C324 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t5 GNDA 0.081909f
C325 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n14 GNDA 0.175188f
C326 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n15 GNDA 0.533147f
C327 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n16 GNDA 0.163405f
C328 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t8 GNDA 0.081909f
C329 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.t4 GNDA 0.081909f
C330 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n17 GNDA 0.175188f
C331 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n18 GNDA 0.540568f
C332 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n19 GNDA 0.189438f
C333 two_stage_opamp_dummy_magic_26_0.V_CMFB_S4.n20 GNDA 2.85233f
C334 bgr_11_0.V_CMFB_S4 GNDA 4.30471f
C335 bgr_11_0.cap_res2.t4 GNDA 0.334798f
C336 bgr_11_0.cap_res2.t10 GNDA 0.336011f
C337 bgr_11_0.cap_res2.t20 GNDA 0.318043f
C338 bgr_11_0.cap_res2.t9 GNDA 0.334798f
C339 bgr_11_0.cap_res2.t14 GNDA 0.336011f
C340 bgr_11_0.cap_res2.t5 GNDA 0.318043f
C341 bgr_11_0.cap_res2.t3 GNDA 0.334798f
C342 bgr_11_0.cap_res2.t8 GNDA 0.336011f
C343 bgr_11_0.cap_res2.t18 GNDA 0.318043f
C344 bgr_11_0.cap_res2.t16 GNDA 0.334798f
C345 bgr_11_0.cap_res2.t2 GNDA 0.336011f
C346 bgr_11_0.cap_res2.t12 GNDA 0.318043f
C347 bgr_11_0.cap_res2.t1 GNDA 0.334798f
C348 bgr_11_0.cap_res2.t6 GNDA 0.336011f
C349 bgr_11_0.cap_res2.t17 GNDA 0.318043f
C350 bgr_11_0.cap_res2.n0 GNDA 0.224415f
C351 bgr_11_0.cap_res2.t11 GNDA 0.178714f
C352 bgr_11_0.cap_res2.n1 GNDA 0.243496f
C353 bgr_11_0.cap_res2.t7 GNDA 0.178714f
C354 bgr_11_0.cap_res2.n2 GNDA 0.243496f
C355 bgr_11_0.cap_res2.t13 GNDA 0.178714f
C356 bgr_11_0.cap_res2.n3 GNDA 0.243496f
C357 bgr_11_0.cap_res2.t19 GNDA 0.178714f
C358 bgr_11_0.cap_res2.n4 GNDA 0.243496f
C359 bgr_11_0.cap_res2.t15 GNDA 0.360089f
C360 bgr_11_0.cap_res2.t0 GNDA 0.082395f
C361 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t1 GNDA 0.245842f
C362 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t5 GNDA 0.773204f
C363 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t7 GNDA 0.772991f
C364 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n0 GNDA 0.636556f
C365 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t2 GNDA 0.772991f
C366 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n1 GNDA 0.331481f
C367 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t3 GNDA 0.772991f
C368 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n2 GNDA 0.667625f
C369 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n3 GNDA 0.790892f
C370 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t0 GNDA 0.245842f
C371 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n4 GNDA 0.431779f
C372 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t9 GNDA 0.667922f
C373 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t4 GNDA 0.667922f
C374 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t6 GNDA 0.667922f
C375 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.t8 GNDA 0.722234f
C376 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n5 GNDA 0.241787f
C377 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n6 GNDA 0.300709f
C378 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n7 GNDA 0.300709f
C379 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n8 GNDA 0.294161f
C380 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n9 GNDA 0.489447f
C381 two_stage_opamp_dummy_magic_26_0.V_b_2nd_stage.n10 GNDA 1.39879f
C382 bgr_11_0.Vin+.t1 GNDA 0.221779f
C383 bgr_11_0.Vin+.t0 GNDA 0.096124f
C384 bgr_11_0.Vin+.n0 GNDA 1.46352f
C385 bgr_11_0.Vin+.t2 GNDA 0.033039f
C386 bgr_11_0.Vin+.t5 GNDA 0.033039f
C387 bgr_11_0.Vin+.n1 GNDA 0.084276f
C388 bgr_11_0.Vin+.t4 GNDA 0.033039f
C389 bgr_11_0.Vin+.t3 GNDA 0.033039f
C390 bgr_11_0.Vin+.n2 GNDA 0.078979f
C391 bgr_11_0.Vin+.n3 GNDA 0.79622f
C392 bgr_11_0.Vin+.n4 GNDA 0.652102f
C393 bgr_11_0.Vin+.t6 GNDA 0.052809f
C394 two_stage_opamp_dummy_magic_26_0.Vb3.n0 GNDA 0.203603f
C395 two_stage_opamp_dummy_magic_26_0.Vb3.n1 GNDA 0.212245f
C396 two_stage_opamp_dummy_magic_26_0.Vb3.n2 GNDA 0.068945f
C397 two_stage_opamp_dummy_magic_26_0.Vb3.n3 GNDA 0.161379f
C398 two_stage_opamp_dummy_magic_26_0.Vb3.n4 GNDA 0.212245f
C399 two_stage_opamp_dummy_magic_26_0.Vb3.n5 GNDA 0.490899f
C400 two_stage_opamp_dummy_magic_26_0.Vb3.n6 GNDA 0.140595f
C401 two_stage_opamp_dummy_magic_26_0.Vb3.n7 GNDA 0.212245f
C402 two_stage_opamp_dummy_magic_26_0.Vb3.n8 GNDA 0.140595f
C403 two_stage_opamp_dummy_magic_26_0.Vb3.n9 GNDA 0.309725f
C404 two_stage_opamp_dummy_magic_26_0.Vb3.t1 GNDA 0.014364f
C405 two_stage_opamp_dummy_magic_26_0.Vb3.t4 GNDA 0.014364f
C406 two_stage_opamp_dummy_magic_26_0.Vb3.n10 GNDA 0.046266f
C407 two_stage_opamp_dummy_magic_26_0.Vb3.t2 GNDA 0.014364f
C408 two_stage_opamp_dummy_magic_26_0.Vb3.t3 GNDA 0.014364f
C409 two_stage_opamp_dummy_magic_26_0.Vb3.n11 GNDA 0.046267f
C410 two_stage_opamp_dummy_magic_26_0.Vb3.n12 GNDA 0.255066f
C411 two_stage_opamp_dummy_magic_26_0.Vb3.t6 GNDA 0.014364f
C412 two_stage_opamp_dummy_magic_26_0.Vb3.t5 GNDA 0.014364f
C413 two_stage_opamp_dummy_magic_26_0.Vb3.n13 GNDA 0.043384f
C414 two_stage_opamp_dummy_magic_26_0.Vb3.n14 GNDA 0.8142f
C415 two_stage_opamp_dummy_magic_26_0.Vb3.t26 GNDA 0.092119f
C416 two_stage_opamp_dummy_magic_26_0.Vb3.t21 GNDA 0.092095f
C417 two_stage_opamp_dummy_magic_26_0.Vb3.t13 GNDA 0.092095f
C418 two_stage_opamp_dummy_magic_26_0.Vb3.t10 GNDA 0.092095f
C419 two_stage_opamp_dummy_magic_26_0.Vb3.t8 GNDA 0.091674f
C420 two_stage_opamp_dummy_magic_26_0.Vb3.t28 GNDA 0.091674f
C421 two_stage_opamp_dummy_magic_26_0.Vb3.t25 GNDA 0.092095f
C422 two_stage_opamp_dummy_magic_26_0.Vb3.t18 GNDA 0.092095f
C423 two_stage_opamp_dummy_magic_26_0.Vb3.t22 GNDA 0.092095f
C424 two_stage_opamp_dummy_magic_26_0.Vb3.t15 GNDA 0.092095f
C425 two_stage_opamp_dummy_magic_26_0.Vb3.t7 GNDA 0.050273f
C426 two_stage_opamp_dummy_magic_26_0.Vb3.t0 GNDA 0.050273f
C427 two_stage_opamp_dummy_magic_26_0.Vb3.n15 GNDA 0.135351f
C428 two_stage_opamp_dummy_magic_26_0.Vb3.t19 GNDA 0.094402f
C429 two_stage_opamp_dummy_magic_26_0.Vb3.n16 GNDA 0.945548f
C430 two_stage_opamp_dummy_magic_26_0.Vb3.n17 GNDA 1.0744f
C431 two_stage_opamp_dummy_magic_26_0.Vb3.t20 GNDA 0.092119f
C432 two_stage_opamp_dummy_magic_26_0.Vb3.t16 GNDA 0.092095f
C433 two_stage_opamp_dummy_magic_26_0.Vb3.t23 GNDA 0.092095f
C434 two_stage_opamp_dummy_magic_26_0.Vb3.t9 GNDA 0.092095f
C435 two_stage_opamp_dummy_magic_26_0.Vb3.t14 GNDA 0.091664f
C436 two_stage_opamp_dummy_magic_26_0.Vb3.t11 GNDA 0.091664f
C437 two_stage_opamp_dummy_magic_26_0.Vb3.n18 GNDA 0.080699f
C438 two_stage_opamp_dummy_magic_26_0.Vb3.n19 GNDA 0.080699f
C439 two_stage_opamp_dummy_magic_26_0.Vb3.t12 GNDA 0.092095f
C440 two_stage_opamp_dummy_magic_26_0.Vb3.t17 GNDA 0.092095f
C441 two_stage_opamp_dummy_magic_26_0.Vb3.t24 GNDA 0.092095f
C442 two_stage_opamp_dummy_magic_26_0.Vb3.t27 GNDA 0.092095f
C443 two_stage_opamp_dummy_magic_26_0.Vb3.n20 GNDA 0.147777f
C444 two_stage_opamp_dummy_magic_26_0.Vb3.n21 GNDA 1.26883f
C445 bgr_11_0.VB3_CUR_BIAS GNDA 1.78766f
C446 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t15 GNDA 0.020643f
C447 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t14 GNDA 0.020643f
C448 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n0 GNDA 0.051768f
C449 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t12 GNDA 0.020643f
C450 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t11 GNDA 0.020643f
C451 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n1 GNDA 0.051495f
C452 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n2 GNDA 0.457775f
C453 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t13 GNDA 0.020643f
C454 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t16 GNDA 0.020643f
C455 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n3 GNDA 0.041287f
C456 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n4 GNDA 0.077381f
C457 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t10 GNDA 0.26037f
C458 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n5 GNDA 0.065212f
C459 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n6 GNDA 0.115348f
C460 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t5 GNDA 0.041287f
C461 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t8 GNDA 0.041287f
C462 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n7 GNDA 0.084415f
C463 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n8 GNDA 0.283547f
C464 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t2 GNDA 0.041287f
C465 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t7 GNDA 0.041287f
C466 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n9 GNDA 0.084415f
C467 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n10 GNDA 0.273057f
C468 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n11 GNDA 0.110879f
C469 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n12 GNDA 0.065212f
C470 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t1 GNDA 0.041287f
C471 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t6 GNDA 0.041287f
C472 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n13 GNDA 0.084415f
C473 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n14 GNDA 0.273057f
C474 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n15 GNDA 0.067596f
C475 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t4 GNDA 0.041287f
C476 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t0 GNDA 0.041287f
C477 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n16 GNDA 0.084415f
C478 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n17 GNDA 0.273057f
C479 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n18 GNDA 0.115348f
C480 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t3 GNDA 0.041287f
C481 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.t9 GNDA 0.041287f
C482 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n19 GNDA 0.084415f
C483 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n20 GNDA 0.278452f
C484 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n21 GNDA 0.150489f
C485 two_stage_opamp_dummy_magic_26_0.V_CMFB_S3.n22 GNDA 2.44046f
C486 bgr_11_0.V_CMFB_S3 GNDA 2.58941f
C487 two_stage_opamp_dummy_magic_26_0.V_err_gate.t2 GNDA 0.026355f
C488 two_stage_opamp_dummy_magic_26_0.V_err_gate.t3 GNDA 0.026355f
C489 two_stage_opamp_dummy_magic_26_0.V_err_gate.n0 GNDA 0.322787f
C490 two_stage_opamp_dummy_magic_26_0.V_err_gate.t0 GNDA 0.065888f
C491 two_stage_opamp_dummy_magic_26_0.V_err_gate.t5 GNDA 0.065888f
C492 two_stage_opamp_dummy_magic_26_0.V_err_gate.n1 GNDA 0.208826f
C493 two_stage_opamp_dummy_magic_26_0.V_err_gate.t6 GNDA 0.073575f
C494 two_stage_opamp_dummy_magic_26_0.V_err_gate.t8 GNDA 0.073575f
C495 two_stage_opamp_dummy_magic_26_0.V_err_gate.n2 GNDA 0.110515f
C496 two_stage_opamp_dummy_magic_26_0.V_err_gate.n3 GNDA 0.400917f
C497 two_stage_opamp_dummy_magic_26_0.V_err_gate.t4 GNDA 0.065888f
C498 two_stage_opamp_dummy_magic_26_0.V_err_gate.t1 GNDA 0.065888f
C499 two_stage_opamp_dummy_magic_26_0.V_err_gate.n4 GNDA 0.207973f
C500 two_stage_opamp_dummy_magic_26_0.V_err_gate.n5 GNDA 0.3051f
C501 two_stage_opamp_dummy_magic_26_0.V_err_gate.t9 GNDA 0.073575f
C502 two_stage_opamp_dummy_magic_26_0.V_err_gate.t7 GNDA 0.073575f
C503 two_stage_opamp_dummy_magic_26_0.V_err_gate.n6 GNDA 0.110515f
C504 two_stage_opamp_dummy_magic_26_0.VD2.t18 GNDA 0.03895f
C505 two_stage_opamp_dummy_magic_26_0.VD2.t13 GNDA 0.03895f
C506 two_stage_opamp_dummy_magic_26_0.VD2.n0 GNDA 0.086232f
C507 two_stage_opamp_dummy_magic_26_0.VD2.n1 GNDA 0.502457f
C508 two_stage_opamp_dummy_magic_26_0.VD2.n2 GNDA 0.058446f
C509 two_stage_opamp_dummy_magic_26_0.VD2.n3 GNDA 0.153053f
C510 two_stage_opamp_dummy_magic_26_0.VD2.t2 GNDA 0.03895f
C511 two_stage_opamp_dummy_magic_26_0.VD2.t1 GNDA 0.03895f
C512 two_stage_opamp_dummy_magic_26_0.VD2.n4 GNDA 0.084751f
C513 two_stage_opamp_dummy_magic_26_0.VD2.n5 GNDA 0.326538f
C514 two_stage_opamp_dummy_magic_26_0.VD2.n6 GNDA 0.082835f
C515 two_stage_opamp_dummy_magic_26_0.VD2.t4 GNDA 0.03895f
C516 two_stage_opamp_dummy_magic_26_0.VD2.t6 GNDA 0.03895f
C517 two_stage_opamp_dummy_magic_26_0.VD2.n7 GNDA 0.084751f
C518 two_stage_opamp_dummy_magic_26_0.VD2.n8 GNDA 0.335643f
C519 two_stage_opamp_dummy_magic_26_0.VD2.t15 GNDA 0.03895f
C520 two_stage_opamp_dummy_magic_26_0.VD2.t11 GNDA 0.03895f
C521 two_stage_opamp_dummy_magic_26_0.VD2.n9 GNDA 0.086232f
C522 two_stage_opamp_dummy_magic_26_0.VD2.t19 GNDA 0.03895f
C523 two_stage_opamp_dummy_magic_26_0.VD2.t14 GNDA 0.03895f
C524 two_stage_opamp_dummy_magic_26_0.VD2.n10 GNDA 0.086232f
C525 two_stage_opamp_dummy_magic_26_0.VD2.n11 GNDA 0.690983f
C526 two_stage_opamp_dummy_magic_26_0.VD2.t17 GNDA 0.03895f
C527 two_stage_opamp_dummy_magic_26_0.VD2.t10 GNDA 0.03895f
C528 two_stage_opamp_dummy_magic_26_0.VD2.n12 GNDA 0.086232f
C529 two_stage_opamp_dummy_magic_26_0.VD2.n13 GNDA 0.205447f
C530 two_stage_opamp_dummy_magic_26_0.VD2.t5 GNDA 0.03895f
C531 two_stage_opamp_dummy_magic_26_0.VD2.t8 GNDA 0.03895f
C532 two_stage_opamp_dummy_magic_26_0.VD2.n14 GNDA 0.084751f
C533 two_stage_opamp_dummy_magic_26_0.VD2.n15 GNDA 0.335643f
C534 two_stage_opamp_dummy_magic_26_0.VD2.n16 GNDA 0.140805f
C535 two_stage_opamp_dummy_magic_26_0.VD2.t7 GNDA 0.03895f
C536 two_stage_opamp_dummy_magic_26_0.VD2.t0 GNDA 0.03895f
C537 two_stage_opamp_dummy_magic_26_0.VD2.n17 GNDA 0.084751f
C538 two_stage_opamp_dummy_magic_26_0.VD2.n18 GNDA 0.326538f
C539 two_stage_opamp_dummy_magic_26_0.VD2.n19 GNDA 0.058446f
C540 two_stage_opamp_dummy_magic_26_0.VD2.n20 GNDA 0.153053f
C541 two_stage_opamp_dummy_magic_26_0.VD2.n21 GNDA 0.684347f
C542 two_stage_opamp_dummy_magic_26_0.VD2.n22 GNDA 0.130987f
C543 two_stage_opamp_dummy_magic_26_0.VD2.n23 GNDA 0.0779f
C544 two_stage_opamp_dummy_magic_26_0.VD2.t16 GNDA 0.03895f
C545 two_stage_opamp_dummy_magic_26_0.VD2.t12 GNDA 0.03895f
C546 two_stage_opamp_dummy_magic_26_0.VD2.n24 GNDA 0.086232f
C547 two_stage_opamp_dummy_magic_26_0.VD2.n25 GNDA 0.684347f
C548 two_stage_opamp_dummy_magic_26_0.VD2.n26 GNDA 0.130987f
C549 two_stage_opamp_dummy_magic_26_0.VD2.n27 GNDA 0.690983f
C550 two_stage_opamp_dummy_magic_26_0.VD2.n28 GNDA 0.205447f
C551 two_stage_opamp_dummy_magic_26_0.VD2.n29 GNDA 0.058446f
C552 two_stage_opamp_dummy_magic_26_0.VD2.t21 GNDA 0.03895f
C553 two_stage_opamp_dummy_magic_26_0.VD2.t9 GNDA 0.03895f
C554 two_stage_opamp_dummy_magic_26_0.VD2.n30 GNDA 0.084751f
C555 two_stage_opamp_dummy_magic_26_0.VD2.n31 GNDA 0.326538f
C556 two_stage_opamp_dummy_magic_26_0.VD2.n32 GNDA 0.140805f
C557 two_stage_opamp_dummy_magic_26_0.VD2.n33 GNDA 0.082835f
C558 two_stage_opamp_dummy_magic_26_0.VD2.t20 GNDA 0.03895f
C559 two_stage_opamp_dummy_magic_26_0.VD2.t3 GNDA 0.03895f
C560 two_stage_opamp_dummy_magic_26_0.VD2.n34 GNDA 0.084751f
C561 two_stage_opamp_dummy_magic_26_0.VD2.n35 GNDA 0.326538f
C562 two_stage_opamp_dummy_magic_26_0.VD2.n36 GNDA 0.058446f
C563 two_stage_opamp_dummy_magic_26_0.VD2.n37 GNDA 0.045235f
C564 bgr_11_0.cap_res1.t5 GNDA 0.339883f
C565 bgr_11_0.cap_res1.t17 GNDA 0.357788f
C566 bgr_11_0.cap_res1.t9 GNDA 0.359085f
C567 bgr_11_0.cap_res1.t12 GNDA 0.339883f
C568 bgr_11_0.cap_res1.t19 GNDA 0.357788f
C569 bgr_11_0.cap_res1.t16 GNDA 0.359085f
C570 bgr_11_0.cap_res1.t4 GNDA 0.339883f
C571 bgr_11_0.cap_res1.t15 GNDA 0.357788f
C572 bgr_11_0.cap_res1.t8 GNDA 0.359085f
C573 bgr_11_0.cap_res1.t0 GNDA 0.339883f
C574 bgr_11_0.cap_res1.t7 GNDA 0.357788f
C575 bgr_11_0.cap_res1.t1 GNDA 0.359085f
C576 bgr_11_0.cap_res1.t2 GNDA 0.339883f
C577 bgr_11_0.cap_res1.t14 GNDA 0.357788f
C578 bgr_11_0.cap_res1.t6 GNDA 0.359085f
C579 bgr_11_0.cap_res1.n0 GNDA 0.239826f
C580 bgr_11_0.cap_res1.t10 GNDA 0.190986f
C581 bgr_11_0.cap_res1.n1 GNDA 0.260216f
C582 bgr_11_0.cap_res1.t3 GNDA 0.190986f
C583 bgr_11_0.cap_res1.n2 GNDA 0.260216f
C584 bgr_11_0.cap_res1.t11 GNDA 0.190986f
C585 bgr_11_0.cap_res1.n3 GNDA 0.260216f
C586 bgr_11_0.cap_res1.t18 GNDA 0.190986f
C587 bgr_11_0.cap_res1.n4 GNDA 0.260216f
C588 bgr_11_0.cap_res1.t13 GNDA 0.383393f
C589 bgr_11_0.cap_res1.t20 GNDA 0.088196f
C590 bgr_11_0.1st_Vout_1.n0 GNDA 0.191219f
C591 bgr_11_0.1st_Vout_1.t27 GNDA 0.240974f
C592 bgr_11_0.1st_Vout_1.t18 GNDA 0.236938f
C593 bgr_11_0.1st_Vout_1.t14 GNDA 0.240974f
C594 bgr_11_0.1st_Vout_1.t23 GNDA 0.236938f
C595 bgr_11_0.1st_Vout_1.n1 GNDA 0.158859f
C596 bgr_11_0.1st_Vout_1.n2 GNDA 0.203285f
C597 bgr_11_0.1st_Vout_1.t32 GNDA 0.240974f
C598 bgr_11_0.1st_Vout_1.t26 GNDA 0.236938f
C599 bgr_11_0.1st_Vout_1.t22 GNDA 0.240974f
C600 bgr_11_0.1st_Vout_1.t31 GNDA 0.236938f
C601 bgr_11_0.1st_Vout_1.n3 GNDA 0.158859f
C602 bgr_11_0.1st_Vout_1.n4 GNDA 0.247711f
C603 bgr_11_0.1st_Vout_1.t25 GNDA 0.240974f
C604 bgr_11_0.1st_Vout_1.t17 GNDA 0.236938f
C605 bgr_11_0.1st_Vout_1.t12 GNDA 0.240974f
C606 bgr_11_0.1st_Vout_1.t21 GNDA 0.236938f
C607 bgr_11_0.1st_Vout_1.n5 GNDA 0.158859f
C608 bgr_11_0.1st_Vout_1.n6 GNDA 0.247711f
C609 bgr_11_0.1st_Vout_1.t16 GNDA 0.240974f
C610 bgr_11_0.1st_Vout_1.t8 GNDA 0.236938f
C611 bgr_11_0.1st_Vout_1.t7 GNDA 0.240974f
C612 bgr_11_0.1st_Vout_1.t11 GNDA 0.236938f
C613 bgr_11_0.1st_Vout_1.n7 GNDA 0.158859f
C614 bgr_11_0.1st_Vout_1.n8 GNDA 0.247711f
C615 bgr_11_0.1st_Vout_1.t24 GNDA 0.240974f
C616 bgr_11_0.1st_Vout_1.t15 GNDA 0.236938f
C617 bgr_11_0.1st_Vout_1.n9 GNDA 0.203285f
C618 bgr_11_0.1st_Vout_1.t20 GNDA 0.236938f
C619 bgr_11_0.1st_Vout_1.n10 GNDA 0.10366f
C620 bgr_11_0.1st_Vout_1.t9 GNDA 0.236938f
C621 bgr_11_0.1st_Vout_1.n11 GNDA 2.00975f
C622 bgr_11_0.1st_Vout_1.t29 GNDA 0.01424f
C623 bgr_11_0.1st_Vout_1.n12 GNDA 3.07165f
C624 bgr_11_0.1st_Vout_1.n13 GNDA 0.012548f
C625 bgr_11_0.1st_Vout_1.n14 GNDA 0.191219f
C626 bgr_11_0.1st_Vout_1.n15 GNDA 0.017467f
C627 bgr_11_0.1st_Vout_1.n16 GNDA 0.173289f
C628 bgr_11_0.1st_Vout_1.n17 GNDA 0.012189f
C629 bgr_11_0.1st_Vout_1.t3 GNDA 0.054022f
C630 bgr_11_0.1st_Vout_1.n18 GNDA 0.173688f
C631 bgr_11_0.1st_Vout_1.n19 GNDA 0.127946f
C632 bgr_11_0.1st_Vout_1.n20 GNDA 0.017467f
C633 bgr_11_0.1st_Vout_1.n21 GNDA 0.173289f
C634 bgr_11_0.1st_Vout_1.n22 GNDA 0.012548f
C635 bgr_11_0.1st_Vout_1.t13 GNDA 0.013988f
C636 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t0 GNDA 0.347912f
C637 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t9 GNDA 0.110048f
C638 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n0 GNDA 3.57839f
C639 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t5 GNDA 0.065833f
C640 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t2 GNDA 0.065833f
C641 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n1 GNDA 0.183642f
C642 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t4 GNDA 0.065833f
C643 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t1 GNDA 0.065833f
C644 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n2 GNDA 0.16529f
C645 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n3 GNDA 2.02985f
C646 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t3 GNDA 0.065833f
C647 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t6 GNDA 0.065833f
C648 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n4 GNDA 0.16529f
C649 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n5 GNDA 1.5092f
C650 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n6 GNDA 0.96323f
C651 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t7 GNDA 0.075599f
C652 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.t8 GNDA 0.074327f
C653 two_stage_opamp_dummy_magic_26_0.V_err_amp_ref.n7 GNDA 0.538641f
C654 bgr_11_0.V_TOP.n0 GNDA 0.016831f
C655 bgr_11_0.V_TOP.t29 GNDA 0.128711f
C656 bgr_11_0.V_TOP.t37 GNDA 0.128973f
C657 bgr_11_0.V_TOP.t38 GNDA 0.129529f
C658 bgr_11_0.V_TOP.n1 GNDA 0.162971f
C659 bgr_11_0.V_TOP.t23 GNDA 0.129529f
C660 bgr_11_0.V_TOP.n2 GNDA 0.089272f
C661 bgr_11_0.V_TOP.t48 GNDA 0.129529f
C662 bgr_11_0.V_TOP.n3 GNDA 0.089272f
C663 bgr_11_0.V_TOP.t39 GNDA 0.129529f
C664 bgr_11_0.V_TOP.n4 GNDA 0.089272f
C665 bgr_11_0.V_TOP.t27 GNDA 0.129529f
C666 bgr_11_0.V_TOP.n5 GNDA 0.089272f
C667 bgr_11_0.V_TOP.n6 GNDA 0.025246f
C668 bgr_11_0.V_TOP.n7 GNDA 0.057364f
C669 bgr_11_0.V_TOP.t6 GNDA 0.129887f
C670 bgr_11_0.V_TOP.t20 GNDA 0.374019f
C671 bgr_11_0.V_TOP.t24 GNDA 0.38039f
C672 bgr_11_0.V_TOP.t32 GNDA 0.374019f
C673 bgr_11_0.V_TOP.n8 GNDA 0.250768f
C674 bgr_11_0.V_TOP.t19 GNDA 0.374019f
C675 bgr_11_0.V_TOP.t46 GNDA 0.38039f
C676 bgr_11_0.V_TOP.n9 GNDA 0.320897f
C677 bgr_11_0.V_TOP.t34 GNDA 0.38039f
C678 bgr_11_0.V_TOP.t40 GNDA 0.374019f
C679 bgr_11_0.V_TOP.n10 GNDA 0.250768f
C680 bgr_11_0.V_TOP.t31 GNDA 0.374019f
C681 bgr_11_0.V_TOP.t18 GNDA 0.38039f
C682 bgr_11_0.V_TOP.n11 GNDA 0.391025f
C683 bgr_11_0.V_TOP.t22 GNDA 0.38039f
C684 bgr_11_0.V_TOP.t30 GNDA 0.374019f
C685 bgr_11_0.V_TOP.n12 GNDA 0.250768f
C686 bgr_11_0.V_TOP.t17 GNDA 0.374019f
C687 bgr_11_0.V_TOP.t44 GNDA 0.38039f
C688 bgr_11_0.V_TOP.n13 GNDA 0.391025f
C689 bgr_11_0.V_TOP.t47 GNDA 0.38039f
C690 bgr_11_0.V_TOP.t16 GNDA 0.374019f
C691 bgr_11_0.V_TOP.n14 GNDA 0.250768f
C692 bgr_11_0.V_TOP.t43 GNDA 0.374019f
C693 bgr_11_0.V_TOP.t35 GNDA 0.38039f
C694 bgr_11_0.V_TOP.n15 GNDA 0.391025f
C695 bgr_11_0.V_TOP.t41 GNDA 0.38039f
C696 bgr_11_0.V_TOP.t15 GNDA 0.374019f
C697 bgr_11_0.V_TOP.n16 GNDA 0.320897f
C698 bgr_11_0.V_TOP.t28 GNDA 0.374019f
C699 bgr_11_0.V_TOP.n17 GNDA 0.163634f
C700 bgr_11_0.V_TOP.n18 GNDA 0.875119f
C701 bgr_11_0.V_TOP.t12 GNDA 0.105245f
C702 bgr_11_0.V_TOP.n19 GNDA 1.42428f
C703 bgr_11_0.V_TOP.n20 GNDA 0.019145f
C704 bgr_11_0.V_TOP.n21 GNDA 0.024925f
C705 bgr_11_0.V_TOP.n22 GNDA 0.022551f
C706 bgr_11_0.V_TOP.n23 GNDA 0.25922f
C707 bgr_11_0.V_TOP.n24 GNDA 0.158514f
C708 bgr_11_0.V_TOP.n25 GNDA 0.655866f
C709 bgr_11_0.V_TOP.n26 GNDA 0.020198f
C710 bgr_11_0.V_TOP.n27 GNDA 0.198604f
C711 bgr_11_0.V_TOP.n28 GNDA 0.020198f
C712 bgr_11_0.V_TOP.n29 GNDA 0.204214f
C713 bgr_11_0.V_TOP.n30 GNDA 0.020198f
C714 bgr_11_0.V_TOP.n31 GNDA 0.190361f
C715 bgr_11_0.V_TOP.n32 GNDA 0.391697f
C716 bgr_11_0.V_TOP.n33 GNDA 0.089765f
C717 bgr_11_0.V_TOP.t14 GNDA 0.127788f
C718 bgr_11_0.V_TOP.n34 GNDA 0.052677f
C719 bgr_11_0.V_TOP.n35 GNDA 0.025246f
C720 bgr_11_0.V_TOP.t45 GNDA 0.128533f
C721 bgr_11_0.V_TOP.n36 GNDA 0.084658f
C722 bgr_11_0.V_TOP.t36 GNDA 0.129529f
C723 bgr_11_0.V_TOP.n37 GNDA 0.089272f
C724 bgr_11_0.V_TOP.t25 GNDA 0.129529f
C725 bgr_11_0.V_TOP.n38 GNDA 0.089272f
C726 bgr_11_0.V_TOP.t26 GNDA 0.129529f
C727 bgr_11_0.V_TOP.n39 GNDA 0.089272f
C728 bgr_11_0.V_TOP.t49 GNDA 0.129529f
C729 bgr_11_0.V_TOP.n40 GNDA 0.089272f
C730 bgr_11_0.V_TOP.t42 GNDA 0.129529f
C731 bgr_11_0.V_TOP.n41 GNDA 0.089272f
C732 bgr_11_0.V_TOP.t33 GNDA 0.129529f
C733 bgr_11_0.V_TOP.n42 GNDA 0.080857f
C734 bgr_11_0.V_TOP.t21 GNDA 0.128562f
C735 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t11 GNDA 0.019824f
C736 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t16 GNDA 0.019824f
C737 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n0 GNDA 0.049693f
C738 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t14 GNDA 0.019824f
C739 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t13 GNDA 0.019824f
C740 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n1 GNDA 0.04943f
C741 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n2 GNDA 0.439335f
C742 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t15 GNDA 0.019824f
C743 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t12 GNDA 0.019824f
C744 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n3 GNDA 0.039648f
C745 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n4 GNDA 0.074337f
C746 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t0 GNDA 0.250301f
C747 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n5 GNDA 0.062624f
C748 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n6 GNDA 0.11077f
C749 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t1 GNDA 0.039648f
C750 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t6 GNDA 0.039648f
C751 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n7 GNDA 0.081065f
C752 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n8 GNDA 0.272294f
C753 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t2 GNDA 0.039648f
C754 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t7 GNDA 0.039648f
C755 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n9 GNDA 0.081065f
C756 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n10 GNDA 0.262221f
C757 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n11 GNDA 0.106479f
C758 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n12 GNDA 0.062624f
C759 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t4 GNDA 0.039648f
C760 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t8 GNDA 0.039648f
C761 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n13 GNDA 0.081065f
C762 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n14 GNDA 0.262221f
C763 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n15 GNDA 0.064914f
C764 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t3 GNDA 0.039648f
C765 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t10 GNDA 0.039648f
C766 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n16 GNDA 0.081065f
C767 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n17 GNDA 0.262221f
C768 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n18 GNDA 0.11077f
C769 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t5 GNDA 0.039648f
C770 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.t9 GNDA 0.039648f
C771 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n19 GNDA 0.081065f
C772 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n20 GNDA 0.267402f
C773 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n21 GNDA 0.144517f
C774 two_stage_opamp_dummy_magic_26_0.V_CMFB_S1.n22 GNDA 2.31344f
C775 bgr_11_0.V_CMFB_S1 GNDA 2.274f
C776 two_stage_opamp_dummy_magic_26_0.VD3.n0 GNDA 1.11096f
C777 two_stage_opamp_dummy_magic_26_0.VD3.n1 GNDA 0.20151f
C778 two_stage_opamp_dummy_magic_26_0.VD3.n2 GNDA 0.378259f
C779 two_stage_opamp_dummy_magic_26_0.VD3.t22 GNDA 0.078836f
C780 two_stage_opamp_dummy_magic_26_0.VD3.n3 GNDA 0.149757f
C781 two_stage_opamp_dummy_magic_26_0.VD3.t32 GNDA 0.045031f
C782 two_stage_opamp_dummy_magic_26_0.VD3.t36 GNDA 0.045031f
C783 two_stage_opamp_dummy_magic_26_0.VD3.n4 GNDA 0.092115f
C784 two_stage_opamp_dummy_magic_26_0.VD3.n5 GNDA 0.260153f
C785 two_stage_opamp_dummy_magic_26_0.VD3.t1 GNDA 0.045031f
C786 two_stage_opamp_dummy_magic_26_0.VD3.t17 GNDA 0.045031f
C787 two_stage_opamp_dummy_magic_26_0.VD3.n6 GNDA 0.095624f
C788 two_stage_opamp_dummy_magic_26_0.VD3.t21 GNDA 0.045031f
C789 two_stage_opamp_dummy_magic_26_0.VD3.t33 GNDA 0.045031f
C790 two_stage_opamp_dummy_magic_26_0.VD3.n7 GNDA 0.092115f
C791 two_stage_opamp_dummy_magic_26_0.VD3.n8 GNDA 0.25692f
C792 two_stage_opamp_dummy_magic_26_0.VD3.t11 GNDA 0.045031f
C793 two_stage_opamp_dummy_magic_26_0.VD3.t15 GNDA 0.045031f
C794 two_stage_opamp_dummy_magic_26_0.VD3.n9 GNDA 0.095624f
C795 two_stage_opamp_dummy_magic_26_0.VD3.t20 GNDA 0.045031f
C796 two_stage_opamp_dummy_magic_26_0.VD3.t29 GNDA 0.045031f
C797 two_stage_opamp_dummy_magic_26_0.VD3.n10 GNDA 0.092115f
C798 two_stage_opamp_dummy_magic_26_0.VD3.n11 GNDA 0.25692f
C799 two_stage_opamp_dummy_magic_26_0.VD3.t5 GNDA 0.045031f
C800 two_stage_opamp_dummy_magic_26_0.VD3.t7 GNDA 0.045031f
C801 two_stage_opamp_dummy_magic_26_0.VD3.n12 GNDA 0.095624f
C802 two_stage_opamp_dummy_magic_26_0.VD3.n13 GNDA 0.76157f
C803 two_stage_opamp_dummy_magic_26_0.VD3.t24 GNDA 0.160181f
C804 two_stage_opamp_dummy_magic_26_0.VD3.n14 GNDA 0.51334f
C805 two_stage_opamp_dummy_magic_26_0.VD3.t23 GNDA 0.383839f
C806 two_stage_opamp_dummy_magic_26_0.VD3.t16 GNDA 0.301063f
C807 two_stage_opamp_dummy_magic_26_0.VD3.t0 GNDA 0.301063f
C808 two_stage_opamp_dummy_magic_26_0.VD3.t14 GNDA 0.301063f
C809 two_stage_opamp_dummy_magic_26_0.VD3.t10 GNDA 0.301063f
C810 two_stage_opamp_dummy_magic_26_0.VD3.t6 GNDA 0.301063f
C811 two_stage_opamp_dummy_magic_26_0.VD3.t4 GNDA 0.301063f
C812 two_stage_opamp_dummy_magic_26_0.VD3.t2 GNDA 0.301063f
C813 two_stage_opamp_dummy_magic_26_0.VD3.t18 GNDA 0.301063f
C814 two_stage_opamp_dummy_magic_26_0.VD3.t12 GNDA 0.301063f
C815 two_stage_opamp_dummy_magic_26_0.VD3.t8 GNDA 0.301063f
C816 two_stage_opamp_dummy_magic_26_0.VD3.t26 GNDA 0.383839f
C817 two_stage_opamp_dummy_magic_26_0.VD3.t27 GNDA 0.160181f
C818 two_stage_opamp_dummy_magic_26_0.VD3.n15 GNDA 0.51334f
C819 two_stage_opamp_dummy_magic_26_0.VD3.t25 GNDA 0.078836f
C820 two_stage_opamp_dummy_magic_26_0.VD3.n16 GNDA 0.215181f
C821 two_stage_opamp_dummy_magic_26_0.VD3.t31 GNDA 0.045031f
C822 two_stage_opamp_dummy_magic_26_0.VD3.t30 GNDA 0.045031f
C823 two_stage_opamp_dummy_magic_26_0.VD3.n17 GNDA 0.092115f
C824 two_stage_opamp_dummy_magic_26_0.VD3.n18 GNDA 0.25692f
C825 two_stage_opamp_dummy_magic_26_0.VD3.t9 GNDA 0.045031f
C826 two_stage_opamp_dummy_magic_26_0.VD3.t13 GNDA 0.045031f
C827 two_stage_opamp_dummy_magic_26_0.VD3.n19 GNDA 0.095624f
C828 two_stage_opamp_dummy_magic_26_0.VD3.n20 GNDA 0.115041f
C829 two_stage_opamp_dummy_magic_26_0.VD3.n21 GNDA 0.069429f
C830 two_stage_opamp_dummy_magic_26_0.VD3.t34 GNDA 0.045031f
C831 two_stage_opamp_dummy_magic_26_0.VD3.t37 GNDA 0.045031f
C832 two_stage_opamp_dummy_magic_26_0.VD3.n22 GNDA 0.092115f
C833 two_stage_opamp_dummy_magic_26_0.VD3.n23 GNDA 0.25692f
C834 two_stage_opamp_dummy_magic_26_0.VD3.n24 GNDA 0.069429f
C835 two_stage_opamp_dummy_magic_26_0.VD3.n25 GNDA 0.115041f
C836 two_stage_opamp_dummy_magic_26_0.VD3.t35 GNDA 0.045031f
C837 two_stage_opamp_dummy_magic_26_0.VD3.t28 GNDA 0.045031f
C838 two_stage_opamp_dummy_magic_26_0.VD3.n26 GNDA 0.092115f
C839 two_stage_opamp_dummy_magic_26_0.VD3.n27 GNDA 0.260153f
C840 two_stage_opamp_dummy_magic_26_0.VD3.t19 GNDA 0.045031f
C841 two_stage_opamp_dummy_magic_26_0.VD3.t3 GNDA 0.045031f
C842 two_stage_opamp_dummy_magic_26_0.VD3.n28 GNDA 0.095624f
C843 two_stage_opamp_dummy_magic_26_0.VD3.n29 GNDA 0.76157f
C844 two_stage_opamp_dummy_magic_26_0.VD3.n30 GNDA 1.26178f
C845 two_stage_opamp_dummy_magic_26_0.VD3.n31 GNDA 0.432296f
C846 two_stage_opamp_dummy_magic_26_0.VD3.n32 GNDA 0.76157f
C847 two_stage_opamp_dummy_magic_26_0.VD3.n33 GNDA 0.76157f
C848 two_stage_opamp_dummy_magic_26_0.VD3.n34 GNDA 0.342878f
C849 two_stage_opamp_dummy_magic_26_0.VD4.n0 GNDA 1.1096f
C850 two_stage_opamp_dummy_magic_26_0.VD4.n1 GNDA 0.201538f
C851 two_stage_opamp_dummy_magic_26_0.VD4.n2 GNDA 0.342878f
C852 two_stage_opamp_dummy_magic_26_0.VD4.n3 GNDA 0.432296f
C853 two_stage_opamp_dummy_magic_26_0.VD4.t15 GNDA 0.045031f
C854 two_stage_opamp_dummy_magic_26_0.VD4.t1 GNDA 0.045031f
C855 two_stage_opamp_dummy_magic_26_0.VD4.n4 GNDA 0.095624f
C856 two_stage_opamp_dummy_magic_26_0.VD4.t31 GNDA 0.045031f
C857 two_stage_opamp_dummy_magic_26_0.VD4.t22 GNDA 0.045031f
C858 two_stage_opamp_dummy_magic_26_0.VD4.n5 GNDA 0.092115f
C859 two_stage_opamp_dummy_magic_26_0.VD4.n6 GNDA 0.25692f
C860 two_stage_opamp_dummy_magic_26_0.VD4.t9 GNDA 0.045031f
C861 two_stage_opamp_dummy_magic_26_0.VD4.t5 GNDA 0.045031f
C862 two_stage_opamp_dummy_magic_26_0.VD4.n7 GNDA 0.095624f
C863 two_stage_opamp_dummy_magic_26_0.VD4.t33 GNDA 0.045031f
C864 two_stage_opamp_dummy_magic_26_0.VD4.t20 GNDA 0.045031f
C865 two_stage_opamp_dummy_magic_26_0.VD4.n8 GNDA 0.092115f
C866 two_stage_opamp_dummy_magic_26_0.VD4.n9 GNDA 0.25692f
C867 two_stage_opamp_dummy_magic_26_0.VD4.t11 GNDA 0.045031f
C868 two_stage_opamp_dummy_magic_26_0.VD4.t13 GNDA 0.045031f
C869 two_stage_opamp_dummy_magic_26_0.VD4.n10 GNDA 0.095624f
C870 two_stage_opamp_dummy_magic_26_0.VD4.t23 GNDA 0.045031f
C871 two_stage_opamp_dummy_magic_26_0.VD4.t32 GNDA 0.045031f
C872 two_stage_opamp_dummy_magic_26_0.VD4.n11 GNDA 0.092115f
C873 two_stage_opamp_dummy_magic_26_0.VD4.n12 GNDA 0.25692f
C874 two_stage_opamp_dummy_magic_26_0.VD4.t17 GNDA 0.045031f
C875 two_stage_opamp_dummy_magic_26_0.VD4.t3 GNDA 0.045031f
C876 two_stage_opamp_dummy_magic_26_0.VD4.n13 GNDA 0.095624f
C877 two_stage_opamp_dummy_magic_26_0.VD4.n14 GNDA 0.76157f
C878 two_stage_opamp_dummy_magic_26_0.VD4.t26 GNDA 0.160181f
C879 two_stage_opamp_dummy_magic_26_0.VD4.t27 GNDA 0.078836f
C880 two_stage_opamp_dummy_magic_26_0.VD4.n15 GNDA 0.149757f
C881 two_stage_opamp_dummy_magic_26_0.VD4.t29 GNDA 0.160181f
C882 two_stage_opamp_dummy_magic_26_0.VD4.n16 GNDA 0.51334f
C883 two_stage_opamp_dummy_magic_26_0.VD4.t28 GNDA 0.383839f
C884 two_stage_opamp_dummy_magic_26_0.VD4.t14 GNDA 0.301063f
C885 two_stage_opamp_dummy_magic_26_0.VD4.t0 GNDA 0.301063f
C886 two_stage_opamp_dummy_magic_26_0.VD4.t8 GNDA 0.301063f
C887 two_stage_opamp_dummy_magic_26_0.VD4.t4 GNDA 0.301063f
C888 two_stage_opamp_dummy_magic_26_0.VD4.t10 GNDA 0.301063f
C889 two_stage_opamp_dummy_magic_26_0.VD4.t12 GNDA 0.301063f
C890 two_stage_opamp_dummy_magic_26_0.VD4.t16 GNDA 0.301063f
C891 two_stage_opamp_dummy_magic_26_0.VD4.t2 GNDA 0.301063f
C892 two_stage_opamp_dummy_magic_26_0.VD4.t18 GNDA 0.301063f
C893 two_stage_opamp_dummy_magic_26_0.VD4.t6 GNDA 0.301063f
C894 two_stage_opamp_dummy_magic_26_0.VD4.t25 GNDA 0.383839f
C895 two_stage_opamp_dummy_magic_26_0.VD4.n17 GNDA 0.51334f
C896 two_stage_opamp_dummy_magic_26_0.VD4.t24 GNDA 0.078836f
C897 two_stage_opamp_dummy_magic_26_0.VD4.n18 GNDA 0.216535f
C898 two_stage_opamp_dummy_magic_26_0.VD4.t35 GNDA 0.045031f
C899 two_stage_opamp_dummy_magic_26_0.VD4.t30 GNDA 0.045031f
C900 two_stage_opamp_dummy_magic_26_0.VD4.n19 GNDA 0.092115f
C901 two_stage_opamp_dummy_magic_26_0.VD4.n20 GNDA 0.260153f
C902 two_stage_opamp_dummy_magic_26_0.VD4.n21 GNDA 0.115041f
C903 two_stage_opamp_dummy_magic_26_0.VD4.n22 GNDA 0.069429f
C904 two_stage_opamp_dummy_magic_26_0.VD4.n23 GNDA 0.069429f
C905 two_stage_opamp_dummy_magic_26_0.VD4.t36 GNDA 0.045031f
C906 two_stage_opamp_dummy_magic_26_0.VD4.t37 GNDA 0.045031f
C907 two_stage_opamp_dummy_magic_26_0.VD4.n24 GNDA 0.092115f
C908 two_stage_opamp_dummy_magic_26_0.VD4.n25 GNDA 0.25692f
C909 two_stage_opamp_dummy_magic_26_0.VD4.n26 GNDA 0.115041f
C910 two_stage_opamp_dummy_magic_26_0.VD4.t21 GNDA 0.045031f
C911 two_stage_opamp_dummy_magic_26_0.VD4.t34 GNDA 0.045031f
C912 two_stage_opamp_dummy_magic_26_0.VD4.n27 GNDA 0.092115f
C913 two_stage_opamp_dummy_magic_26_0.VD4.n28 GNDA 0.260153f
C914 two_stage_opamp_dummy_magic_26_0.VD4.t19 GNDA 0.045031f
C915 two_stage_opamp_dummy_magic_26_0.VD4.t7 GNDA 0.045031f
C916 two_stage_opamp_dummy_magic_26_0.VD4.n29 GNDA 0.095624f
C917 two_stage_opamp_dummy_magic_26_0.VD4.n30 GNDA 1.26176f
C918 two_stage_opamp_dummy_magic_26_0.VD4.n31 GNDA 0.76157f
C919 two_stage_opamp_dummy_magic_26_0.VD4.n32 GNDA 0.76157f
C920 two_stage_opamp_dummy_magic_26_0.VD4.n33 GNDA 0.76157f
C921 two_stage_opamp_dummy_magic_26_0.VD4.n34 GNDA 0.378259f
C922 two_stage_opamp_dummy_magic_26_0.Vb2.n0 GNDA 0.473604f
C923 two_stage_opamp_dummy_magic_26_0.Vb2.n1 GNDA 0.478939f
C924 two_stage_opamp_dummy_magic_26_0.Vb2.n2 GNDA 0.473604f
C925 two_stage_opamp_dummy_magic_26_0.Vb2.n3 GNDA 0.478939f
C926 two_stage_opamp_dummy_magic_26_0.Vb2.n4 GNDA 0.530034f
C927 two_stage_opamp_dummy_magic_26_0.Vb2.n5 GNDA 0.504815f
C928 two_stage_opamp_dummy_magic_26_0.Vb2.t5 GNDA 0.061734f
C929 two_stage_opamp_dummy_magic_26_0.Vb2.t19 GNDA 0.113135f
C930 two_stage_opamp_dummy_magic_26_0.Vb2.t17 GNDA 0.113092f
C931 two_stage_opamp_dummy_magic_26_0.Vb2.t12 GNDA 0.113092f
C932 two_stage_opamp_dummy_magic_26_0.Vb2.t27 GNDA 0.113092f
C933 two_stage_opamp_dummy_magic_26_0.Vb2.t23 GNDA 0.113092f
C934 two_stage_opamp_dummy_magic_26_0.Vb2.t21 GNDA 0.113092f
C935 two_stage_opamp_dummy_magic_26_0.Vb2.t18 GNDA 0.113092f
C936 two_stage_opamp_dummy_magic_26_0.Vb2.t16 GNDA 0.113092f
C937 two_stage_opamp_dummy_magic_26_0.Vb2.t32 GNDA 0.113092f
C938 two_stage_opamp_dummy_magic_26_0.Vb2.t13 GNDA 0.113092f
C939 two_stage_opamp_dummy_magic_26_0.Vb2.t2 GNDA 0.017638f
C940 two_stage_opamp_dummy_magic_26_0.Vb2.t3 GNDA 0.017638f
C941 two_stage_opamp_dummy_magic_26_0.Vb2.n6 GNDA 0.059139f
C942 two_stage_opamp_dummy_magic_26_0.Vb2.t9 GNDA 0.017638f
C943 two_stage_opamp_dummy_magic_26_0.Vb2.t8 GNDA 0.017638f
C944 two_stage_opamp_dummy_magic_26_0.Vb2.n7 GNDA 0.057517f
C945 two_stage_opamp_dummy_magic_26_0.Vb2.n8 GNDA 0.535082f
C946 two_stage_opamp_dummy_magic_26_0.Vb2.t7 GNDA 0.017638f
C947 two_stage_opamp_dummy_magic_26_0.Vb2.t6 GNDA 0.017638f
C948 two_stage_opamp_dummy_magic_26_0.Vb2.n9 GNDA 0.057517f
C949 two_stage_opamp_dummy_magic_26_0.Vb2.n10 GNDA 0.354339f
C950 two_stage_opamp_dummy_magic_26_0.Vb2.t4 GNDA 0.017638f
C951 two_stage_opamp_dummy_magic_26_0.Vb2.t10 GNDA 0.017638f
C952 two_stage_opamp_dummy_magic_26_0.Vb2.n11 GNDA 0.057517f
C953 two_stage_opamp_dummy_magic_26_0.Vb2.n12 GNDA 2.23443f
C954 two_stage_opamp_dummy_magic_26_0.Vb2.n13 GNDA 2.02851f
C955 two_stage_opamp_dummy_magic_26_0.Vb2.t20 GNDA 0.113464f
C956 two_stage_opamp_dummy_magic_26_0.Vb2.n14 GNDA 0.357216f
C957 two_stage_opamp_dummy_magic_26_0.Vb2.t28 GNDA 0.070909f
C958 two_stage_opamp_dummy_magic_26_0.Vb2.n15 GNDA 0.370277f
C959 two_stage_opamp_dummy_magic_26_0.Vb2.t26 GNDA 0.113135f
C960 two_stage_opamp_dummy_magic_26_0.Vb2.t11 GNDA 0.113092f
C961 two_stage_opamp_dummy_magic_26_0.Vb2.t30 GNDA 0.113092f
C962 two_stage_opamp_dummy_magic_26_0.Vb2.t14 GNDA 0.113092f
C963 two_stage_opamp_dummy_magic_26_0.Vb2.t22 GNDA 0.113092f
C964 two_stage_opamp_dummy_magic_26_0.Vb2.t24 GNDA 0.113092f
C965 two_stage_opamp_dummy_magic_26_0.Vb2.t29 GNDA 0.113092f
C966 two_stage_opamp_dummy_magic_26_0.Vb2.t25 GNDA 0.113092f
C967 two_stage_opamp_dummy_magic_26_0.Vb2.t31 GNDA 0.113092f
C968 two_stage_opamp_dummy_magic_26_0.Vb2.t15 GNDA 0.113092f
C969 two_stage_opamp_dummy_magic_26_0.Vb2.n16 GNDA 0.389785f
C970 two_stage_opamp_dummy_magic_26_0.Vb2.t0 GNDA 0.116811f
C971 two_stage_opamp_dummy_magic_26_0.Vb2.n17 GNDA 0.499716f
C972 two_stage_opamp_dummy_magic_26_0.Vb2.n18 GNDA 0.131339f
C973 two_stage_opamp_dummy_magic_26_0.Vb2.t1 GNDA 0.061734f
C974 two_stage_opamp_dummy_magic_26_0.Y.n0 GNDA 0.090278f
C975 two_stage_opamp_dummy_magic_26_0.Y.n1 GNDA 0.106905f
C976 two_stage_opamp_dummy_magic_26_0.Y.n2 GNDA 0.110339f
C977 two_stage_opamp_dummy_magic_26_0.Y.n3 GNDA 0.378191f
C978 two_stage_opamp_dummy_magic_26_0.Y.n4 GNDA 0.106905f
C979 two_stage_opamp_dummy_magic_26_0.Y.n5 GNDA 0.106905f
C980 two_stage_opamp_dummy_magic_26_0.Y.t20 GNDA 0.025077f
C981 two_stage_opamp_dummy_magic_26_0.Y.t3 GNDA 0.025077f
C982 two_stage_opamp_dummy_magic_26_0.Y.n6 GNDA 0.073693f
C983 two_stage_opamp_dummy_magic_26_0.Y.t17 GNDA 0.025077f
C984 two_stage_opamp_dummy_magic_26_0.Y.t14 GNDA 0.025077f
C985 two_stage_opamp_dummy_magic_26_0.Y.n7 GNDA 0.072264f
C986 two_stage_opamp_dummy_magic_26_0.Y.n8 GNDA 0.477627f
C987 two_stage_opamp_dummy_magic_26_0.Y.t15 GNDA 0.025077f
C988 two_stage_opamp_dummy_magic_26_0.Y.t18 GNDA 0.025077f
C989 two_stage_opamp_dummy_magic_26_0.Y.n9 GNDA 0.072264f
C990 two_stage_opamp_dummy_magic_26_0.Y.n10 GNDA 0.251231f
C991 two_stage_opamp_dummy_magic_26_0.Y.t16 GNDA 0.025077f
C992 two_stage_opamp_dummy_magic_26_0.Y.t11 GNDA 0.025077f
C993 two_stage_opamp_dummy_magic_26_0.Y.n11 GNDA 0.072264f
C994 two_stage_opamp_dummy_magic_26_0.Y.n12 GNDA 0.251231f
C995 two_stage_opamp_dummy_magic_26_0.Y.t12 GNDA 0.025077f
C996 two_stage_opamp_dummy_magic_26_0.Y.t19 GNDA 0.025077f
C997 two_stage_opamp_dummy_magic_26_0.Y.n13 GNDA 0.072264f
C998 two_stage_opamp_dummy_magic_26_0.Y.n14 GNDA 0.251231f
C999 two_stage_opamp_dummy_magic_26_0.Y.t2 GNDA 0.025077f
C1000 two_stage_opamp_dummy_magic_26_0.Y.t13 GNDA 0.025077f
C1001 two_stage_opamp_dummy_magic_26_0.Y.n15 GNDA 0.072264f
C1002 two_stage_opamp_dummy_magic_26_0.Y.n16 GNDA 0.446833f
C1003 two_stage_opamp_dummy_magic_26_0.Y.n17 GNDA 0.306485f
C1004 two_stage_opamp_dummy_magic_26_0.Y.n18 GNDA 0.467678f
C1005 two_stage_opamp_dummy_magic_26_0.Y.n19 GNDA 0.400848f
C1006 two_stage_opamp_dummy_magic_26_0.Y.n20 GNDA 0.110339f
C1007 two_stage_opamp_dummy_magic_26_0.Y.n21 GNDA 0.364545f
C1008 two_stage_opamp_dummy_magic_26_0.Y.n22 GNDA 0.110339f
C1009 two_stage_opamp_dummy_magic_26_0.Y.n23 GNDA 0.110339f
C1010 two_stage_opamp_dummy_magic_26_0.Y.n24 GNDA 0.110339f
C1011 two_stage_opamp_dummy_magic_26_0.Y.n25 GNDA 0.185719f
C1012 two_stage_opamp_dummy_magic_26_0.Y.n27 GNDA 0.080247f
C1013 two_stage_opamp_dummy_magic_26_0.Y.n28 GNDA 0.090217f
C1014 two_stage_opamp_dummy_magic_26_0.Y.n29 GNDA 0.090217f
C1015 two_stage_opamp_dummy_magic_26_0.Y.t10 GNDA 0.058513f
C1016 two_stage_opamp_dummy_magic_26_0.Y.t22 GNDA 0.058513f
C1017 two_stage_opamp_dummy_magic_26_0.Y.n30 GNDA 0.119695f
C1018 two_stage_opamp_dummy_magic_26_0.Y.n31 GNDA 0.385354f
C1019 two_stage_opamp_dummy_magic_26_0.Y.n32 GNDA 0.149485f
C1020 two_stage_opamp_dummy_magic_26_0.Y.t23 GNDA 0.058513f
C1021 two_stage_opamp_dummy_magic_26_0.Y.t5 GNDA 0.058513f
C1022 two_stage_opamp_dummy_magic_26_0.Y.n33 GNDA 0.119695f
C1023 two_stage_opamp_dummy_magic_26_0.Y.n34 GNDA 0.376954f
C1024 two_stage_opamp_dummy_magic_26_0.Y.n35 GNDA 0.149485f
C1025 two_stage_opamp_dummy_magic_26_0.Y.t4 GNDA 0.058513f
C1026 two_stage_opamp_dummy_magic_26_0.Y.t1 GNDA 0.058513f
C1027 two_stage_opamp_dummy_magic_26_0.Y.n36 GNDA 0.119695f
C1028 two_stage_opamp_dummy_magic_26_0.Y.n37 GNDA 0.376954f
C1029 two_stage_opamp_dummy_magic_26_0.Y.n38 GNDA 0.090217f
C1030 two_stage_opamp_dummy_magic_26_0.Y.n39 GNDA 0.090217f
C1031 two_stage_opamp_dummy_magic_26_0.Y.t21 GNDA 0.058513f
C1032 two_stage_opamp_dummy_magic_26_0.Y.t0 GNDA 0.058513f
C1033 two_stage_opamp_dummy_magic_26_0.Y.n40 GNDA 0.119695f
C1034 two_stage_opamp_dummy_magic_26_0.Y.n41 GNDA 0.376954f
C1035 two_stage_opamp_dummy_magic_26_0.Y.n42 GNDA 0.090217f
C1036 two_stage_opamp_dummy_magic_26_0.Y.t7 GNDA 0.058513f
C1037 two_stage_opamp_dummy_magic_26_0.Y.t8 GNDA 0.058513f
C1038 two_stage_opamp_dummy_magic_26_0.Y.n43 GNDA 0.119695f
C1039 two_stage_opamp_dummy_magic_26_0.Y.n44 GNDA 0.376954f
C1040 two_stage_opamp_dummy_magic_26_0.Y.n45 GNDA 0.149485f
C1041 two_stage_opamp_dummy_magic_26_0.Y.t6 GNDA 0.058513f
C1042 two_stage_opamp_dummy_magic_26_0.Y.t9 GNDA 0.058513f
C1043 two_stage_opamp_dummy_magic_26_0.Y.n46 GNDA 0.119695f
C1044 two_stage_opamp_dummy_magic_26_0.Y.n47 GNDA 0.381154f
C1045 two_stage_opamp_dummy_magic_26_0.Y.n48 GNDA 0.238347f
C1046 two_stage_opamp_dummy_magic_26_0.Y.n49 GNDA 0.080247f
C1047 two_stage_opamp_dummy_magic_26_0.Y.n51 GNDA 0.080247f
C1048 two_stage_opamp_dummy_magic_26_0.Y.n52 GNDA 0.080247f
C1049 two_stage_opamp_dummy_magic_26_0.Y.n53 GNDA 0.079493f
C1050 two_stage_opamp_dummy_magic_26_0.Y.n54 GNDA 0.080247f
C1051 two_stage_opamp_dummy_magic_26_0.Y.t24 GNDA 0.693898f
C1052 two_stage_opamp_dummy_magic_26_0.Y.n55 GNDA 0.080247f
C1053 two_stage_opamp_dummy_magic_26_0.Y.n56 GNDA 0.080247f
C1054 two_stage_opamp_dummy_magic_26_0.Y.n58 GNDA 0.744527f
C1055 two_stage_opamp_dummy_magic_26_0.Y.n60 GNDA 0.697145f
C1056 two_stage_opamp_dummy_magic_26_0.Y.n61 GNDA 0.026571f
C1057 two_stage_opamp_dummy_magic_26_0.Y.n62 GNDA 0.026749f
C1058 two_stage_opamp_dummy_magic_26_0.Y.n63 GNDA 0.026749f
C1059 two_stage_opamp_dummy_magic_26_0.Y.t35 GNDA 0.110339f
C1060 two_stage_opamp_dummy_magic_26_0.Y.t41 GNDA 0.110339f
C1061 two_stage_opamp_dummy_magic_26_0.Y.t25 GNDA 0.110339f
C1062 two_stage_opamp_dummy_magic_26_0.Y.t43 GNDA 0.110339f
C1063 two_stage_opamp_dummy_magic_26_0.Y.t28 GNDA 0.117519f
C1064 two_stage_opamp_dummy_magic_26_0.Y.n64 GNDA 0.093129f
C1065 two_stage_opamp_dummy_magic_26_0.Y.n65 GNDA 0.052662f
C1066 two_stage_opamp_dummy_magic_26_0.Y.n66 GNDA 0.052662f
C1067 two_stage_opamp_dummy_magic_26_0.Y.n67 GNDA 0.047333f
C1068 two_stage_opamp_dummy_magic_26_0.Y.t48 GNDA 0.110339f
C1069 two_stage_opamp_dummy_magic_26_0.Y.t32 GNDA 0.110339f
C1070 two_stage_opamp_dummy_magic_26_0.Y.t45 GNDA 0.110339f
C1071 two_stage_opamp_dummy_magic_26_0.Y.t29 GNDA 0.110339f
C1072 two_stage_opamp_dummy_magic_26_0.Y.t38 GNDA 0.117519f
C1073 two_stage_opamp_dummy_magic_26_0.Y.n68 GNDA 0.093129f
C1074 two_stage_opamp_dummy_magic_26_0.Y.n69 GNDA 0.052662f
C1075 two_stage_opamp_dummy_magic_26_0.Y.n70 GNDA 0.052662f
C1076 two_stage_opamp_dummy_magic_26_0.Y.n71 GNDA 0.047333f
C1077 two_stage_opamp_dummy_magic_26_0.Y.n72 GNDA 0.011366f
C1078 two_stage_opamp_dummy_magic_26_0.Y.n73 GNDA 0.026927f
C1079 two_stage_opamp_dummy_magic_26_0.Y.n74 GNDA 0.063383f
C1080 two_stage_opamp_dummy_magic_26_0.Y.n75 GNDA 0.036151f
C1081 two_stage_opamp_dummy_magic_26_0.Y.n76 GNDA 0.041026f
C1082 two_stage_opamp_dummy_magic_26_0.Y.n77 GNDA 1.10841f
C1083 two_stage_opamp_dummy_magic_26_0.Y.t37 GNDA 0.053916f
C1084 two_stage_opamp_dummy_magic_26_0.Y.t51 GNDA 0.053916f
C1085 two_stage_opamp_dummy_magic_26_0.Y.t39 GNDA 0.053916f
C1086 two_stage_opamp_dummy_magic_26_0.Y.t52 GNDA 0.053916f
C1087 two_stage_opamp_dummy_magic_26_0.Y.t30 GNDA 0.053916f
C1088 two_stage_opamp_dummy_magic_26_0.Y.t46 GNDA 0.053916f
C1089 two_stage_opamp_dummy_magic_26_0.Y.t33 GNDA 0.053916f
C1090 two_stage_opamp_dummy_magic_26_0.Y.t49 GNDA 0.061293f
C1091 two_stage_opamp_dummy_magic_26_0.Y.n79 GNDA 0.055315f
C1092 two_stage_opamp_dummy_magic_26_0.Y.n80 GNDA 0.033854f
C1093 two_stage_opamp_dummy_magic_26_0.Y.n81 GNDA 0.033854f
C1094 two_stage_opamp_dummy_magic_26_0.Y.n82 GNDA 0.033854f
C1095 two_stage_opamp_dummy_magic_26_0.Y.n83 GNDA 0.033854f
C1096 two_stage_opamp_dummy_magic_26_0.Y.n84 GNDA 0.033854f
C1097 two_stage_opamp_dummy_magic_26_0.Y.n85 GNDA 0.028525f
C1098 two_stage_opamp_dummy_magic_26_0.Y.t50 GNDA 0.053916f
C1099 two_stage_opamp_dummy_magic_26_0.Y.t53 GNDA 0.061293f
C1100 two_stage_opamp_dummy_magic_26_0.Y.n86 GNDA 0.049987f
C1101 two_stage_opamp_dummy_magic_26_0.Y.n87 GNDA 0.013852f
C1102 two_stage_opamp_dummy_magic_26_0.Y.t44 GNDA 0.035108f
C1103 two_stage_opamp_dummy_magic_26_0.Y.t31 GNDA 0.035108f
C1104 two_stage_opamp_dummy_magic_26_0.Y.t47 GNDA 0.035108f
C1105 two_stage_opamp_dummy_magic_26_0.Y.t34 GNDA 0.035108f
C1106 two_stage_opamp_dummy_magic_26_0.Y.t40 GNDA 0.035108f
C1107 two_stage_opamp_dummy_magic_26_0.Y.t54 GNDA 0.035108f
C1108 two_stage_opamp_dummy_magic_26_0.Y.t42 GNDA 0.035108f
C1109 two_stage_opamp_dummy_magic_26_0.Y.t26 GNDA 0.042631f
C1110 two_stage_opamp_dummy_magic_26_0.Y.n88 GNDA 0.042631f
C1111 two_stage_opamp_dummy_magic_26_0.Y.n89 GNDA 0.027585f
C1112 two_stage_opamp_dummy_magic_26_0.Y.n90 GNDA 0.027585f
C1113 two_stage_opamp_dummy_magic_26_0.Y.n91 GNDA 0.027585f
C1114 two_stage_opamp_dummy_magic_26_0.Y.n92 GNDA 0.027585f
C1115 two_stage_opamp_dummy_magic_26_0.Y.n93 GNDA 0.027585f
C1116 two_stage_opamp_dummy_magic_26_0.Y.n94 GNDA 0.022256f
C1117 two_stage_opamp_dummy_magic_26_0.Y.t27 GNDA 0.035108f
C1118 two_stage_opamp_dummy_magic_26_0.Y.t36 GNDA 0.042631f
C1119 two_stage_opamp_dummy_magic_26_0.Y.n95 GNDA 0.037302f
C1120 two_stage_opamp_dummy_magic_26_0.Y.n96 GNDA 0.013852f
C1121 two_stage_opamp_dummy_magic_26_0.Y.n97 GNDA 0.068968f
C1122 two_stage_opamp_dummy_magic_26_0.Y.n98 GNDA 0.079493f
C1123 two_stage_opamp_dummy_magic_26_0.Y.n99 GNDA 0.080247f
C1124 two_stage_opamp_dummy_magic_26_0.Y.n100 GNDA 0.080247f
C1125 two_stage_opamp_dummy_magic_26_0.Y.n101 GNDA 0.080247f
C1126 two_stage_opamp_dummy_magic_26_0.Y.n102 GNDA 0.080247f
C1127 two_stage_opamp_dummy_magic_26_0.Y.n104 GNDA 0.403211f
C1128 two_stage_opamp_dummy_magic_26_0.Y.n105 GNDA 1.80902f
C1129 two_stage_opamp_dummy_magic_26_0.Y.n106 GNDA 0.080247f
C1130 two_stage_opamp_dummy_magic_26_0.Y.n107 GNDA 0.858763f
C1131 two_stage_opamp_dummy_magic_26_0.Y.n108 GNDA 0.491512f
C1132 two_stage_opamp_dummy_magic_26_0.Y.n110 GNDA 0.662037f
C1133 two_stage_opamp_dummy_magic_26_0.Y.n111 GNDA 0.662037f
C1134 two_stage_opamp_dummy_magic_26_0.Y.n112 GNDA 0.079493f
C1135 two_stage_opamp_dummy_magic_26_0.Y.n114 GNDA 0.671057f
C1136 two_stage_opamp_dummy_magic_26_0.Y.n116 GNDA 0.64699f
C1137 two_stage_opamp_dummy_magic_26_0.Y.n117 GNDA 0.662037f
C1138 two_stage_opamp_dummy_magic_26_0.Y.n118 GNDA 0.354185f
C1139 two_stage_opamp_dummy_magic_26_0.Y.n119 GNDA 0.110339f
C1140 two_stage_opamp_dummy_magic_26_0.Y.n120 GNDA 0.364545f
C1141 two_stage_opamp_dummy_magic_26_0.Y.n121 GNDA 0.110339f
C1142 two_stage_opamp_dummy_magic_26_0.Y.n122 GNDA 0.110339f
C1143 two_stage_opamp_dummy_magic_26_0.Y.n123 GNDA 0.110339f
C1144 two_stage_opamp_dummy_magic_26_0.Y.n124 GNDA 0.329437f
C1145 two_stage_opamp_dummy_magic_26_0.V_source.n0 GNDA 0.041641f
C1146 two_stage_opamp_dummy_magic_26_0.V_source.n1 GNDA 1.0922f
C1147 two_stage_opamp_dummy_magic_26_0.V_source.n2 GNDA 1.1386f
C1148 two_stage_opamp_dummy_magic_26_0.V_source.n3 GNDA 0.889198f
C1149 two_stage_opamp_dummy_magic_26_0.V_source.n4 GNDA 0.306665f
C1150 two_stage_opamp_dummy_magic_26_0.V_source.t7 GNDA 0.021688f
C1151 two_stage_opamp_dummy_magic_26_0.V_source.t31 GNDA 0.021688f
C1152 two_stage_opamp_dummy_magic_26_0.V_source.n5 GNDA 0.046365f
C1153 two_stage_opamp_dummy_magic_26_0.V_source.n6 GNDA 0.18241f
C1154 two_stage_opamp_dummy_magic_26_0.V_source.n7 GNDA 0.04232f
C1155 two_stage_opamp_dummy_magic_26_0.V_source.t25 GNDA 0.021688f
C1156 two_stage_opamp_dummy_magic_26_0.V_source.t16 GNDA 0.021688f
C1157 two_stage_opamp_dummy_magic_26_0.V_source.n8 GNDA 0.046365f
C1158 two_stage_opamp_dummy_magic_26_0.V_source.n9 GNDA 0.146965f
C1159 two_stage_opamp_dummy_magic_26_0.V_source.n10 GNDA 0.138926f
C1160 two_stage_opamp_dummy_magic_26_0.V_source.n11 GNDA 0.138926f
C1161 two_stage_opamp_dummy_magic_26_0.V_source.n12 GNDA 0.148924f
C1162 two_stage_opamp_dummy_magic_26_0.V_source.n13 GNDA 0.070236f
C1163 two_stage_opamp_dummy_magic_26_0.V_source.n14 GNDA 0.047311f
C1164 two_stage_opamp_dummy_magic_26_0.V_source.t38 GNDA 0.013013f
C1165 two_stage_opamp_dummy_magic_26_0.V_source.t27 GNDA 0.013013f
C1166 two_stage_opamp_dummy_magic_26_0.V_source.n15 GNDA 0.028314f
C1167 two_stage_opamp_dummy_magic_26_0.V_source.n16 GNDA 0.118832f
C1168 two_stage_opamp_dummy_magic_26_0.V_source.t29 GNDA 0.013013f
C1169 two_stage_opamp_dummy_magic_26_0.V_source.t4 GNDA 0.013013f
C1170 two_stage_opamp_dummy_magic_26_0.V_source.n17 GNDA 0.028314f
C1171 two_stage_opamp_dummy_magic_26_0.V_source.n18 GNDA 0.114722f
C1172 two_stage_opamp_dummy_magic_26_0.V_source.n19 GNDA 0.070236f
C1173 two_stage_opamp_dummy_magic_26_0.V_source.n20 GNDA 0.054559f
C1174 two_stage_opamp_dummy_magic_26_0.V_source.t30 GNDA 0.013013f
C1175 two_stage_opamp_dummy_magic_26_0.V_source.t37 GNDA 0.013013f
C1176 two_stage_opamp_dummy_magic_26_0.V_source.n21 GNDA 0.028314f
C1177 two_stage_opamp_dummy_magic_26_0.V_source.n22 GNDA 0.114722f
C1178 two_stage_opamp_dummy_magic_26_0.V_source.n23 GNDA 0.027812f
C1179 two_stage_opamp_dummy_magic_26_0.V_source.n24 GNDA 0.027812f
C1180 two_stage_opamp_dummy_magic_26_0.V_source.t6 GNDA 0.013013f
C1181 two_stage_opamp_dummy_magic_26_0.V_source.t40 GNDA 0.013013f
C1182 two_stage_opamp_dummy_magic_26_0.V_source.n25 GNDA 0.028314f
C1183 two_stage_opamp_dummy_magic_26_0.V_source.n26 GNDA 0.085929f
C1184 two_stage_opamp_dummy_magic_26_0.V_source.t5 GNDA 0.013013f
C1185 two_stage_opamp_dummy_magic_26_0.V_source.t28 GNDA 0.013013f
C1186 two_stage_opamp_dummy_magic_26_0.V_source.n27 GNDA 0.028314f
C1187 two_stage_opamp_dummy_magic_26_0.V_source.n28 GNDA 0.085929f
C1188 two_stage_opamp_dummy_magic_26_0.V_source.n29 GNDA 0.07032f
C1189 two_stage_opamp_dummy_magic_26_0.V_source.t33 GNDA 0.013013f
C1190 two_stage_opamp_dummy_magic_26_0.V_source.t32 GNDA 0.013013f
C1191 two_stage_opamp_dummy_magic_26_0.V_source.n30 GNDA 0.028314f
C1192 two_stage_opamp_dummy_magic_26_0.V_source.n31 GNDA 0.085929f
C1193 two_stage_opamp_dummy_magic_26_0.V_source.n32 GNDA 0.07032f
C1194 two_stage_opamp_dummy_magic_26_0.V_source.t0 GNDA 0.013013f
C1195 two_stage_opamp_dummy_magic_26_0.V_source.t2 GNDA 0.013013f
C1196 two_stage_opamp_dummy_magic_26_0.V_source.n33 GNDA 0.028314f
C1197 two_stage_opamp_dummy_magic_26_0.V_source.n34 GNDA 0.085929f
C1198 two_stage_opamp_dummy_magic_26_0.V_source.n35 GNDA 0.027812f
C1199 two_stage_opamp_dummy_magic_26_0.V_source.t34 GNDA 0.013013f
C1200 two_stage_opamp_dummy_magic_26_0.V_source.t8 GNDA 0.013013f
C1201 two_stage_opamp_dummy_magic_26_0.V_source.n36 GNDA 0.028314f
C1202 two_stage_opamp_dummy_magic_26_0.V_source.n37 GNDA 0.118832f
C1203 two_stage_opamp_dummy_magic_26_0.V_source.t3 GNDA 0.013013f
C1204 two_stage_opamp_dummy_magic_26_0.V_source.t39 GNDA 0.013013f
C1205 two_stage_opamp_dummy_magic_26_0.V_source.n38 GNDA 0.028314f
C1206 two_stage_opamp_dummy_magic_26_0.V_source.n39 GNDA 0.114722f
C1207 two_stage_opamp_dummy_magic_26_0.V_source.n40 GNDA 0.047311f
C1208 two_stage_opamp_dummy_magic_26_0.V_source.n41 GNDA 0.027812f
C1209 two_stage_opamp_dummy_magic_26_0.V_source.t1 GNDA 0.013013f
C1210 two_stage_opamp_dummy_magic_26_0.V_source.t36 GNDA 0.013013f
C1211 two_stage_opamp_dummy_magic_26_0.V_source.n42 GNDA 0.028314f
C1212 two_stage_opamp_dummy_magic_26_0.V_source.n43 GNDA 0.114722f
C1213 two_stage_opamp_dummy_magic_26_0.V_source.n44 GNDA 0.054559f
C1214 two_stage_opamp_dummy_magic_26_0.V_source.n45 GNDA 0.148924f
C1215 two_stage_opamp_dummy_magic_26_0.V_source.t22 GNDA 0.021688f
C1216 two_stage_opamp_dummy_magic_26_0.V_source.t12 GNDA 0.021688f
C1217 two_stage_opamp_dummy_magic_26_0.V_source.n46 GNDA 0.046365f
C1218 two_stage_opamp_dummy_magic_26_0.V_source.n47 GNDA 0.146965f
C1219 two_stage_opamp_dummy_magic_26_0.V_source.t21 GNDA 0.021688f
C1220 two_stage_opamp_dummy_magic_26_0.V_source.t11 GNDA 0.021688f
C1221 two_stage_opamp_dummy_magic_26_0.V_source.n48 GNDA 0.046365f
C1222 two_stage_opamp_dummy_magic_26_0.V_source.n49 GNDA 0.146965f
C1223 two_stage_opamp_dummy_magic_26_0.V_source.n50 GNDA 0.138926f
C1224 two_stage_opamp_dummy_magic_26_0.V_source.n51 GNDA 0.041641f
C1225 two_stage_opamp_dummy_magic_26_0.V_source.t10 GNDA 0.021688f
C1226 two_stage_opamp_dummy_magic_26_0.V_source.t17 GNDA 0.021688f
C1227 two_stage_opamp_dummy_magic_26_0.V_source.n53 GNDA 0.046365f
C1228 two_stage_opamp_dummy_magic_26_0.V_source.n54 GNDA 0.146965f
C1229 two_stage_opamp_dummy_magic_26_0.V_source.n55 GNDA 0.138926f
C1230 two_stage_opamp_dummy_magic_26_0.V_source.t15 GNDA 0.021688f
C1231 two_stage_opamp_dummy_magic_26_0.V_source.t19 GNDA 0.021688f
C1232 two_stage_opamp_dummy_magic_26_0.V_source.n56 GNDA 0.046365f
C1233 two_stage_opamp_dummy_magic_26_0.V_source.n57 GNDA 0.146965f
C1234 two_stage_opamp_dummy_magic_26_0.V_source.n58 GNDA 0.138926f
C1235 two_stage_opamp_dummy_magic_26_0.V_source.n59 GNDA 1.01369f
C1236 two_stage_opamp_dummy_magic_26_0.V_source.t35 GNDA 0.047819f
C1237 two_stage_opamp_dummy_magic_26_0.V_source.n60 GNDA 1.62399f
C1238 two_stage_opamp_dummy_magic_26_0.V_source.n61 GNDA 0.481468f
C1239 two_stage_opamp_dummy_magic_26_0.V_source.n62 GNDA 0.041641f
C1240 two_stage_opamp_dummy_magic_26_0.V_source.n63 GNDA 0.041641f
C1241 two_stage_opamp_dummy_magic_26_0.V_source.n65 GNDA 0.726854f
C1242 two_stage_opamp_dummy_magic_26_0.V_source.n66 GNDA 0.682106f
C1243 two_stage_opamp_dummy_magic_26_0.V_source.t18 GNDA 0.021688f
C1244 two_stage_opamp_dummy_magic_26_0.V_source.t26 GNDA 0.021688f
C1245 two_stage_opamp_dummy_magic_26_0.V_source.n67 GNDA 0.046365f
C1246 two_stage_opamp_dummy_magic_26_0.V_source.n68 GNDA 0.146966f
C1247 two_stage_opamp_dummy_magic_26_0.V_source.n69 GNDA 0.119105f
C1248 two_stage_opamp_dummy_magic_26_0.V_source.t9 GNDA 0.021688f
C1249 two_stage_opamp_dummy_magic_26_0.V_source.t13 GNDA 0.021688f
C1250 two_stage_opamp_dummy_magic_26_0.V_source.n70 GNDA 0.046365f
C1251 two_stage_opamp_dummy_magic_26_0.V_source.n71 GNDA 0.176215f
C1252 two_stage_opamp_dummy_magic_26_0.V_source.n72 GNDA 0.138926f
C1253 two_stage_opamp_dummy_magic_26_0.V_source.t23 GNDA 0.021688f
C1254 two_stage_opamp_dummy_magic_26_0.V_source.t20 GNDA 0.021688f
C1255 two_stage_opamp_dummy_magic_26_0.V_source.n73 GNDA 0.046365f
C1256 two_stage_opamp_dummy_magic_26_0.V_source.n74 GNDA 0.176215f
C1257 two_stage_opamp_dummy_magic_26_0.V_source.n75 GNDA 0.138926f
C1258 two_stage_opamp_dummy_magic_26_0.V_source.n76 GNDA 0.138926f
C1259 two_stage_opamp_dummy_magic_26_0.V_source.t24 GNDA 0.021688f
C1260 two_stage_opamp_dummy_magic_26_0.V_source.t14 GNDA 0.021688f
C1261 two_stage_opamp_dummy_magic_26_0.V_source.n77 GNDA 0.046365f
C1262 two_stage_opamp_dummy_magic_26_0.V_source.n78 GNDA 0.176215f
C1263 two_stage_opamp_dummy_magic_26_0.V_source.n79 GNDA 0.066721f
C1264 two_stage_opamp_dummy_magic_26_0.V_source.n80 GNDA 0.114089f
C1265 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n0 GNDA 7.1978f
C1266 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n1 GNDA 10.9345f
C1267 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n2 GNDA 0.174244f
C1268 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n3 GNDA 6.78312f
C1269 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t1 GNDA 0.011902f
C1270 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t11 GNDA 0.011902f
C1271 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n4 GNDA 0.026342f
C1272 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n5 GNDA 0.200994f
C1273 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t25 GNDA 0.021127f
C1274 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t14 GNDA 0.021127f
C1275 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t23 GNDA 0.021127f
C1276 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t13 GNDA 0.021127f
C1277 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t22 GNDA 0.021127f
C1278 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t30 GNDA 0.021127f
C1279 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t20 GNDA 0.021127f
C1280 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t24 GNDA 0.024658f
C1281 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n6 GNDA 0.023249f
C1282 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n7 GNDA 0.01458f
C1283 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n8 GNDA 0.01458f
C1284 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n9 GNDA 0.01458f
C1285 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n10 GNDA 0.01458f
C1286 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n11 GNDA 0.01458f
C1287 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n12 GNDA 0.013644f
C1288 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n13 GNDA 0.012355f
C1289 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n14 GNDA 0.01587f
C1290 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n15 GNDA 0.01587f
C1291 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n16 GNDA 0.028817f
C1292 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n17 GNDA 0.090862f
C1293 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n18 GNDA 0.01587f
C1294 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n19 GNDA 0.173786f
C1295 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n20 GNDA 0.090862f
C1296 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n21 GNDA 0.01587f
C1297 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n22 GNDA 0.174254f
C1298 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t2 GNDA 0.011902f
C1299 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t0 GNDA 0.011902f
C1300 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n23 GNDA 0.026342f
C1301 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n24 GNDA 0.209834f
C1302 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t19 GNDA 0.021127f
C1303 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t16 GNDA 0.021127f
C1304 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n25 GNDA 0.013644f
C1305 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n26 GNDA 0.013644f
C1306 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t31 GNDA 0.021127f
C1307 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t27 GNDA 0.021127f
C1308 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t17 GNDA 0.021127f
C1309 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t28 GNDA 0.021127f
C1310 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t18 GNDA 0.021127f
C1311 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t29 GNDA 0.021127f
C1312 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t21 GNDA 0.021127f
C1313 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t12 GNDA 0.021127f
C1314 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t15 GNDA 0.021127f
C1315 two_stage_opamp_dummy_magic_26_0.V_tail_gate.t26 GNDA 0.024658f
C1316 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n27 GNDA 0.023249f
C1317 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n28 GNDA 0.01458f
C1318 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n29 GNDA 0.01458f
C1319 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n30 GNDA 0.01458f
C1320 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n31 GNDA 0.01458f
C1321 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n32 GNDA 0.01458f
C1322 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n33 GNDA 0.01458f
C1323 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n34 GNDA 0.01458f
C1324 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n35 GNDA 0.013644f
C1325 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n36 GNDA 0.012355f
C1326 two_stage_opamp_dummy_magic_26_0.V_tail_gate.n37 GNDA 0.207617f
C1327 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t13 GNDA 0.408922f
C1328 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t43 GNDA 0.428972f
C1329 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t46 GNDA 0.408922f
C1330 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t86 GNDA 0.21964f
C1331 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n0 GNDA 0.235069f
C1332 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t32 GNDA 0.408922f
C1333 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t62 GNDA 0.21964f
C1334 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n1 GNDA 0.233173f
C1335 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t67 GNDA 0.408922f
C1336 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t100 GNDA 0.21964f
C1337 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n2 GNDA 0.233173f
C1338 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t102 GNDA 0.408922f
C1339 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t0 GNDA 0.21964f
C1340 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n3 GNDA 0.233173f
C1341 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t5 GNDA 0.408922f
C1342 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t36 GNDA 0.21964f
C1343 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n4 GNDA 0.233173f
C1344 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t128 GNDA 0.408922f
C1345 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t17 GNDA 0.21964f
C1346 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n5 GNDA 0.233173f
C1347 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t12 GNDA 0.408922f
C1348 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t81 GNDA 0.410404f
C1349 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t34 GNDA 0.408922f
C1350 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t75 GNDA 0.410404f
C1351 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t124 GNDA 0.408922f
C1352 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t40 GNDA 0.410404f
C1353 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t18 GNDA 0.408922f
C1354 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t48 GNDA 0.410404f
C1355 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t130 GNDA 0.408922f
C1356 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t77 GNDA 0.410404f
C1357 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t52 GNDA 0.408922f
C1358 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t91 GNDA 0.410404f
C1359 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t25 GNDA 0.408922f
C1360 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t120 GNDA 0.410404f
C1361 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t24 GNDA 0.408922f
C1362 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t54 GNDA 0.410404f
C1363 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t135 GNDA 0.408922f
C1364 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t82 GNDA 0.410404f
C1365 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t60 GNDA 0.408922f
C1366 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t96 GNDA 0.410404f
C1367 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t31 GNDA 0.408922f
C1368 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t126 GNDA 0.410404f
C1369 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t98 GNDA 0.408922f
C1370 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t137 GNDA 0.410404f
C1371 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t68 GNDA 0.408922f
C1372 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t22 GNDA 0.410404f
C1373 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t66 GNDA 0.408922f
C1374 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t99 GNDA 0.410404f
C1375 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t33 GNDA 0.408922f
C1376 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t131 GNDA 0.410404f
C1377 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t108 GNDA 0.408922f
C1378 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t4 GNDA 0.410404f
C1379 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t76 GNDA 0.408922f
C1380 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t29 GNDA 0.410404f
C1381 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t7 GNDA 0.408922f
C1382 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t39 GNDA 0.410404f
C1383 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t118 GNDA 0.408922f
C1384 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t63 GNDA 0.410404f
C1385 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t41 GNDA 0.408922f
C1386 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t84 GNDA 0.410404f
C1387 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t14 GNDA 0.408922f
C1388 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t103 GNDA 0.410404f
C1389 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t11 GNDA 0.408922f
C1390 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t42 GNDA 0.410404f
C1391 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t125 GNDA 0.408922f
C1392 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t71 GNDA 0.410404f
C1393 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t47 GNDA 0.408922f
C1394 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t87 GNDA 0.410404f
C1395 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t20 GNDA 0.408922f
C1396 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t113 GNDA 0.410404f
C1397 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t90 GNDA 0.408922f
C1398 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t133 GNDA 0.410404f
C1399 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t57 GNDA 0.408922f
C1400 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t9 GNDA 0.410404f
C1401 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t53 GNDA 0.408922f
C1402 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t92 GNDA 0.410404f
C1403 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t26 GNDA 0.408922f
C1404 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t121 GNDA 0.410404f
C1405 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t116 GNDA 0.408922f
C1406 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t61 GNDA 0.410404f
C1407 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t109 GNDA 0.408922f
C1408 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t44 GNDA 0.410404f
C1409 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t106 GNDA 0.408922f
C1410 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t2 GNDA 0.410404f
C1411 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t74 GNDA 0.408922f
C1412 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t27 GNDA 0.410404f
C1413 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t1 GNDA 0.408922f
C1414 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t35 GNDA 0.410404f
C1415 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t110 GNDA 0.408922f
C1416 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t58 GNDA 0.410404f
C1417 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t45 GNDA 0.408922f
C1418 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t89 GNDA 0.428972f
C1419 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t88 GNDA 0.408922f
C1420 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t134 GNDA 0.21964f
C1421 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n6 GNDA 0.235069f
C1422 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t64 GNDA 0.408922f
C1423 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t104 GNDA 0.21964f
C1424 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n7 GNDA 0.233173f
C1425 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t101 GNDA 0.408922f
C1426 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t6 GNDA 0.21964f
C1427 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n8 GNDA 0.233173f
C1428 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t3 GNDA 0.408922f
C1429 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t38 GNDA 0.21964f
C1430 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n9 GNDA 0.233173f
C1431 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t37 GNDA 0.408922f
C1432 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t80 GNDA 0.21964f
C1433 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n10 GNDA 0.233173f
C1434 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t19 GNDA 0.408922f
C1435 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t56 GNDA 0.21964f
C1436 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n11 GNDA 0.233173f
C1437 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t51 GNDA 0.408922f
C1438 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t95 GNDA 0.21964f
C1439 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n12 GNDA 0.233173f
C1440 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t94 GNDA 0.408922f
C1441 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t136 GNDA 0.21964f
C1442 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n13 GNDA 0.233173f
C1443 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t73 GNDA 0.408922f
C1444 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t115 GNDA 0.21964f
C1445 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n14 GNDA 0.233173f
C1446 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t112 GNDA 0.408922f
C1447 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t8 GNDA 0.21964f
C1448 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n15 GNDA 0.233173f
C1449 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t49 GNDA 0.408922f
C1450 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t129 GNDA 0.410404f
C1451 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t15 GNDA 0.408922f
C1452 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t85 GNDA 0.410404f
C1453 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t119 GNDA 0.197694f
C1454 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n16 GNDA 0.254996f
C1455 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t16 GNDA 0.218281f
C1456 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n17 GNDA 0.276942f
C1457 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t59 GNDA 0.218281f
C1458 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n18 GNDA 0.297406f
C1459 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t28 GNDA 0.218281f
C1460 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n19 GNDA 0.297406f
C1461 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t97 GNDA 0.218281f
C1462 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n20 GNDA 0.297406f
C1463 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t123 GNDA 0.218281f
C1464 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n21 GNDA 0.297406f
C1465 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t10 GNDA 0.218281f
C1466 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n22 GNDA 0.297406f
C1467 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t114 GNDA 0.218281f
C1468 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n23 GNDA 0.297406f
C1469 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t72 GNDA 0.218281f
C1470 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n24 GNDA 0.297406f
C1471 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t107 GNDA 0.218281f
C1472 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n25 GNDA 0.297406f
C1473 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t65 GNDA 0.218281f
C1474 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n26 GNDA 0.297406f
C1475 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t30 GNDA 0.218281f
C1476 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n27 GNDA 0.297406f
C1477 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t132 GNDA 0.218281f
C1478 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n28 GNDA 0.297406f
C1479 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t23 GNDA 0.218281f
C1480 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n29 GNDA 0.297406f
C1481 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t127 GNDA 0.218281f
C1482 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n30 GNDA 0.297406f
C1483 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t83 GNDA 0.218281f
C1484 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n31 GNDA 0.297406f
C1485 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t122 GNDA 0.218281f
C1486 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n32 GNDA 0.297406f
C1487 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t78 GNDA 0.218281f
C1488 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n33 GNDA 0.297406f
C1489 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t79 GNDA 0.218281f
C1490 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n34 GNDA 0.297406f
C1491 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t117 GNDA 0.218281f
C1492 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n35 GNDA 0.257642f
C1493 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t111 GNDA 0.410404f
C1494 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t69 GNDA 0.410404f
C1495 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t105 GNDA 0.408922f
C1496 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t55 GNDA 0.430868f
C1497 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t93 GNDA 0.21964f
C1498 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n36 GNDA 0.253637f
C1499 two_stage_opamp_dummy_magic_26_0.cap_res_Y.n37 GNDA 0.233173f
C1500 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t50 GNDA 0.21964f
C1501 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t21 GNDA 0.430868f
C1502 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t70 GNDA 0.517768f
C1503 two_stage_opamp_dummy_magic_26_0.cap_res_Y.t138 GNDA 0.362101f
C1504 VOUT+.n0 GNDA 0.037009f
C1505 VOUT+.t11 GNDA 0.053972f
C1506 VOUT+.t5 GNDA 0.053972f
C1507 VOUT+.n1 GNDA 0.115965f
C1508 VOUT+.n2 GNDA 0.284675f
C1509 VOUT+.n3 GNDA 0.037009f
C1510 VOUT+.n4 GNDA 0.245545f
C1511 VOUT+.t6 GNDA 0.053972f
C1512 VOUT+.t3 GNDA 0.053972f
C1513 VOUT+.n5 GNDA 0.115965f
C1514 VOUT+.n6 GNDA 0.293651f
C1515 VOUT+.n7 GNDA 0.164981f
C1516 VOUT+.t15 GNDA 0.053972f
C1517 VOUT+.t0 GNDA 0.053972f
C1518 VOUT+.n8 GNDA 0.115965f
C1519 VOUT+.n9 GNDA 0.279983f
C1520 VOUT+.n10 GNDA 0.13162f
C1521 VOUT+.n11 GNDA 0.037009f
C1522 VOUT+.n12 GNDA 0.190971f
C1523 VOUT+.n13 GNDA 0.037009f
C1524 VOUT+.n14 GNDA 0.037009f
C1525 VOUT+.n15 GNDA 0.037009f
C1526 VOUT+.n16 GNDA 0.037009f
C1527 VOUT+.n17 GNDA 0.085005f
C1528 VOUT+.n18 GNDA 0.099462f
C1529 VOUT+.n19 GNDA 0.077102f
C1530 VOUT+.n22 GNDA 0.039322f
C1531 VOUT+.n24 GNDA 0.039322f
C1532 VOUT+.n27 GNDA 0.057827f
C1533 VOUT+.n28 GNDA 0.096378f
C1534 VOUT+.n29 GNDA 0.061265f
C1535 VOUT+.n30 GNDA 0.057827f
C1536 VOUT+.n32 GNDA 0.039322f
C1537 VOUT+.n33 GNDA 0.036662f
C1538 VOUT+.n34 GNDA 0.039322f
C1539 VOUT+.n35 GNDA 0.050888f
C1540 VOUT+.n36 GNDA 0.073419f
C1541 VOUT+.n37 GNDA 0.071448f
C1542 VOUT+.n38 GNDA 0.050888f
C1543 VOUT+.n39 GNDA 0.050888f
C1544 VOUT+.n40 GNDA 0.071448f
C1545 VOUT+.n41 GNDA 0.071448f
C1546 VOUT+.n42 GNDA 0.050888f
C1547 VOUT+.n43 GNDA 0.081467f
C1548 VOUT+.t13 GNDA 0.046262f
C1549 VOUT+.t9 GNDA 0.046262f
C1550 VOUT+.n44 GNDA 0.09479f
C1551 VOUT+.n45 GNDA 0.24468f
C1552 VOUT+.t2 GNDA 0.046262f
C1553 VOUT+.t14 GNDA 0.046262f
C1554 VOUT+.n46 GNDA 0.09479f
C1555 VOUT+.n47 GNDA 0.24468f
C1556 VOUT+.t17 GNDA 0.046262f
C1557 VOUT+.t16 GNDA 0.046262f
C1558 VOUT+.n48 GNDA 0.09479f
C1559 VOUT+.n49 GNDA 0.242214f
C1560 VOUT+.n50 GNDA 0.058826f
C1561 VOUT+.t10 GNDA 0.046262f
C1562 VOUT+.t18 GNDA 0.046262f
C1563 VOUT+.n51 GNDA 0.09479f
C1564 VOUT+.n52 GNDA 0.242214f
C1565 VOUT+.n53 GNDA 0.033345f
C1566 VOUT+.t12 GNDA 0.046262f
C1567 VOUT+.t1 GNDA 0.046262f
C1568 VOUT+.n54 GNDA 0.09479f
C1569 VOUT+.n55 GNDA 0.242214f
C1570 VOUT+.n56 GNDA 0.033345f
C1571 VOUT+.n57 GNDA 0.058826f
C1572 VOUT+.t4 GNDA 0.046262f
C1573 VOUT+.t8 GNDA 0.046262f
C1574 VOUT+.n58 GNDA 0.09479f
C1575 VOUT+.n59 GNDA 0.242214f
C1576 VOUT+.n60 GNDA 0.038894f
C1577 VOUT+.n61 GNDA 0.023131f
C1578 VOUT+.n62 GNDA 0.023131f
C1579 VOUT+.n63 GNDA 0.038894f
C1580 VOUT+.n64 GNDA 0.071448f
C1581 VOUT+.n65 GNDA 0.100013f
C1582 VOUT+.n66 GNDA 0.124621f
C1583 VOUT+.n67 GNDA 0.174419f
C1584 VOUT+.n68 GNDA 0.050888f
C1585 VOUT+.n69 GNDA 0.083271f
C1586 VOUT+.n70 GNDA 0.050888f
C1587 VOUT+.n71 GNDA 0.083271f
C1588 VOUT+.n72 GNDA 0.050888f
C1589 VOUT+.n73 GNDA 0.050888f
C1590 VOUT+.n74 GNDA 0.050888f
C1591 VOUT+.n75 GNDA 0.083271f
C1592 VOUT+.n76 GNDA 0.050888f
C1593 VOUT+.n77 GNDA 0.076331f
C1594 VOUT+.n78 GNDA 0.245186f
C1595 VOUT+.n80 GNDA 0.077102f
C1596 VOUT+.n81 GNDA 0.039322f
C1597 VOUT+.n83 GNDA 0.039322f
C1598 VOUT+.n86 GNDA 0.077102f
C1599 VOUT+.n87 GNDA 0.238247f
C1600 VOUT+.n88 GNDA 0.510804f
C1601 VOUT+.n91 GNDA 0.057827f
C1602 VOUT+.n92 GNDA 0.057827f
C1603 VOUT+.n93 GNDA 0.057827f
C1604 VOUT+.n94 GNDA 0.057827f
C1605 VOUT+.n95 GNDA 0.169615f
C1606 VOUT+.n96 GNDA 0.057827f
C1607 VOUT+.t37 GNDA 0.30841f
C1608 VOUT+.t141 GNDA 0.313663f
C1609 VOUT+.t71 GNDA 0.30841f
C1610 VOUT+.n97 GNDA 0.206779f
C1611 VOUT+.n98 GNDA 0.134929f
C1612 VOUT+.t44 GNDA 0.313005f
C1613 VOUT+.t83 GNDA 0.313005f
C1614 VOUT+.t62 GNDA 0.313005f
C1615 VOUT+.t105 GNDA 0.313005f
C1616 VOUT+.t137 GNDA 0.313005f
C1617 VOUT+.t119 GNDA 0.313005f
C1618 VOUT+.t153 GNDA 0.313005f
C1619 VOUT+.t55 GNDA 0.313005f
C1620 VOUT+.t92 GNDA 0.313005f
C1621 VOUT+.t68 GNDA 0.313005f
C1622 VOUT+.t111 GNDA 0.313005f
C1623 VOUT+.t67 GNDA 0.30841f
C1624 VOUT+.n99 GNDA 0.207436f
C1625 VOUT+.t22 GNDA 0.30841f
C1626 VOUT+.n100 GNDA 0.265263f
C1627 VOUT+.t52 GNDA 0.30841f
C1628 VOUT+.n101 GNDA 0.265263f
C1629 VOUT+.t150 GNDA 0.30841f
C1630 VOUT+.n102 GNDA 0.265263f
C1631 VOUT+.t118 GNDA 0.30841f
C1632 VOUT+.n103 GNDA 0.265263f
C1633 VOUT+.t76 GNDA 0.30841f
C1634 VOUT+.n104 GNDA 0.265263f
C1635 VOUT+.t100 GNDA 0.30841f
C1636 VOUT+.n105 GNDA 0.265263f
C1637 VOUT+.t61 GNDA 0.30841f
C1638 VOUT+.n106 GNDA 0.265263f
C1639 VOUT+.t20 GNDA 0.30841f
C1640 VOUT+.n107 GNDA 0.265263f
C1641 VOUT+.t41 GNDA 0.30841f
C1642 VOUT+.n108 GNDA 0.265263f
C1643 VOUT+.t148 GNDA 0.30841f
C1644 VOUT+.n109 GNDA 0.265263f
C1645 VOUT+.t140 GNDA 0.30841f
C1646 VOUT+.t107 GNDA 0.313663f
C1647 VOUT+.t27 GNDA 0.30841f
C1648 VOUT+.n110 GNDA 0.206779f
C1649 VOUT+.n111 GNDA 0.250583f
C1650 VOUT+.t155 GNDA 0.313663f
C1651 VOUT+.t121 GNDA 0.30841f
C1652 VOUT+.n112 GNDA 0.206779f
C1653 VOUT+.t97 GNDA 0.30841f
C1654 VOUT+.t46 GNDA 0.313663f
C1655 VOUT+.t98 GNDA 0.30841f
C1656 VOUT+.n113 GNDA 0.206779f
C1657 VOUT+.n114 GNDA 0.250583f
C1658 VOUT+.t50 GNDA 0.313663f
C1659 VOUT+.t154 GNDA 0.30841f
C1660 VOUT+.n115 GNDA 0.206779f
C1661 VOUT+.t128 GNDA 0.30841f
C1662 VOUT+.t82 GNDA 0.313663f
C1663 VOUT+.t129 GNDA 0.30841f
C1664 VOUT+.n116 GNDA 0.206779f
C1665 VOUT+.n117 GNDA 0.250583f
C1666 VOUT+.t40 GNDA 0.313663f
C1667 VOUT+.t95 GNDA 0.30841f
C1668 VOUT+.n118 GNDA 0.206779f
C1669 VOUT+.t59 GNDA 0.30841f
C1670 VOUT+.t47 GNDA 0.313663f
C1671 VOUT+.t112 GNDA 0.30841f
C1672 VOUT+.n119 GNDA 0.206779f
C1673 VOUT+.n120 GNDA 0.250583f
C1674 VOUT+.t103 GNDA 0.313663f
C1675 VOUT+.t64 GNDA 0.30841f
C1676 VOUT+.n121 GNDA 0.206779f
C1677 VOUT+.t33 GNDA 0.30841f
C1678 VOUT+.t130 GNDA 0.313663f
C1679 VOUT+.t35 GNDA 0.30841f
C1680 VOUT+.n122 GNDA 0.206779f
C1681 VOUT+.n123 GNDA 0.250583f
C1682 VOUT+.t66 GNDA 0.313663f
C1683 VOUT+.t23 GNDA 0.30841f
C1684 VOUT+.n124 GNDA 0.206779f
C1685 VOUT+.t146 GNDA 0.30841f
C1686 VOUT+.t99 GNDA 0.313663f
C1687 VOUT+.t147 GNDA 0.30841f
C1688 VOUT+.n125 GNDA 0.206779f
C1689 VOUT+.n126 GNDA 0.250583f
C1690 VOUT+.t109 GNDA 0.313663f
C1691 VOUT+.t69 GNDA 0.30841f
C1692 VOUT+.n127 GNDA 0.206779f
C1693 VOUT+.t42 GNDA 0.30841f
C1694 VOUT+.t136 GNDA 0.313663f
C1695 VOUT+.t43 GNDA 0.30841f
C1696 VOUT+.n128 GNDA 0.206779f
C1697 VOUT+.n129 GNDA 0.250583f
C1698 VOUT+.t145 GNDA 0.313663f
C1699 VOUT+.t114 GNDA 0.30841f
C1700 VOUT+.n130 GNDA 0.206779f
C1701 VOUT+.t84 GNDA 0.30841f
C1702 VOUT+.t31 GNDA 0.313663f
C1703 VOUT+.t85 GNDA 0.30841f
C1704 VOUT+.n131 GNDA 0.206779f
C1705 VOUT+.n132 GNDA 0.250583f
C1706 VOUT+.t51 GNDA 0.313663f
C1707 VOUT+.t101 GNDA 0.30841f
C1708 VOUT+.n133 GNDA 0.20196f
C1709 VOUT+.t86 GNDA 0.313663f
C1710 VOUT+.t135 GNDA 0.30841f
C1711 VOUT+.n134 GNDA 0.20196f
C1712 VOUT+.t28 GNDA 0.31325f
C1713 VOUT+.t151 GNDA 0.31325f
C1714 VOUT+.t54 GNDA 0.313263f
C1715 VOUT+.t89 GNDA 0.313263f
C1716 VOUT+.t124 GNDA 0.31325f
C1717 VOUT+.t110 GNDA 0.313263f
C1718 VOUT+.t143 GNDA 0.313263f
C1719 VOUT+.t113 GNDA 0.30841f
C1720 VOUT+.n135 GNDA 0.211033f
C1721 VOUT+.t70 GNDA 0.30841f
C1722 VOUT+.n136 GNDA 0.26886f
C1723 VOUT+.t94 GNDA 0.30841f
C1724 VOUT+.n137 GNDA 0.268873f
C1725 VOUT+.t56 GNDA 0.30841f
C1726 VOUT+.n138 GNDA 0.26886f
C1727 VOUT+.t156 GNDA 0.30841f
C1728 VOUT+.n139 GNDA 0.26886f
C1729 VOUT+.t120 GNDA 0.30841f
C1730 VOUT+.n140 GNDA 0.268873f
C1731 VOUT+.t139 GNDA 0.30841f
C1732 VOUT+.n141 GNDA 0.268873f
C1733 VOUT+.t106 GNDA 0.30841f
C1734 VOUT+.n142 GNDA 0.197575f
C1735 VOUT+.t63 GNDA 0.30841f
C1736 VOUT+.n143 GNDA 0.197575f
C1737 VOUT+.t87 GNDA 0.30841f
C1738 VOUT+.n144 GNDA 0.134929f
C1739 VOUT+.t45 GNDA 0.30841f
C1740 VOUT+.n145 GNDA 0.134929f
C1741 VOUT+.t39 GNDA 0.30841f
C1742 VOUT+.t144 GNDA 0.313663f
C1743 VOUT+.t75 GNDA 0.30841f
C1744 VOUT+.n146 GNDA 0.206779f
C1745 VOUT+.n147 GNDA 0.14264f
C1746 VOUT+.t122 GNDA 0.313663f
C1747 VOUT+.t81 GNDA 0.30841f
C1748 VOUT+.n148 GNDA 0.206779f
C1749 VOUT+.t77 GNDA 0.30841f
C1750 VOUT+.t32 GNDA 0.313663f
C1751 VOUT+.t116 GNDA 0.30841f
C1752 VOUT+.n149 GNDA 0.206779f
C1753 VOUT+.n150 GNDA 0.250583f
C1754 VOUT+.t138 GNDA 0.313663f
C1755 VOUT+.t108 GNDA 0.30841f
C1756 VOUT+.n151 GNDA 0.206779f
C1757 VOUT+.t78 GNDA 0.30841f
C1758 VOUT+.t26 GNDA 0.313663f
C1759 VOUT+.t79 GNDA 0.30841f
C1760 VOUT+.n152 GNDA 0.206779f
C1761 VOUT+.n153 GNDA 0.250583f
C1762 VOUT+.t104 GNDA 0.313663f
C1763 VOUT+.t65 GNDA 0.30841f
C1764 VOUT+.n154 GNDA 0.206779f
C1765 VOUT+.t34 GNDA 0.30841f
C1766 VOUT+.t131 GNDA 0.313663f
C1767 VOUT+.t36 GNDA 0.30841f
C1768 VOUT+.n155 GNDA 0.206779f
C1769 VOUT+.n156 GNDA 0.250583f
C1770 VOUT+.t132 GNDA 0.313663f
C1771 VOUT+.t102 GNDA 0.30841f
C1772 VOUT+.n157 GNDA 0.206779f
C1773 VOUT+.t73 GNDA 0.30841f
C1774 VOUT+.t21 GNDA 0.313663f
C1775 VOUT+.t74 GNDA 0.30841f
C1776 VOUT+.n158 GNDA 0.206779f
C1777 VOUT+.n159 GNDA 0.250583f
C1778 VOUT+.t96 GNDA 0.313663f
C1779 VOUT+.t60 GNDA 0.30841f
C1780 VOUT+.n160 GNDA 0.206779f
C1781 VOUT+.t29 GNDA 0.30841f
C1782 VOUT+.t125 GNDA 0.313663f
C1783 VOUT+.t30 GNDA 0.30841f
C1784 VOUT+.n161 GNDA 0.206779f
C1785 VOUT+.n162 GNDA 0.250583f
C1786 VOUT+.t58 GNDA 0.313663f
C1787 VOUT+.t19 GNDA 0.30841f
C1788 VOUT+.n163 GNDA 0.206779f
C1789 VOUT+.t133 GNDA 0.30841f
C1790 VOUT+.t88 GNDA 0.313663f
C1791 VOUT+.t134 GNDA 0.30841f
C1792 VOUT+.n164 GNDA 0.206779f
C1793 VOUT+.n165 GNDA 0.250583f
C1794 VOUT+.t90 GNDA 0.313663f
C1795 VOUT+.t57 GNDA 0.30841f
C1796 VOUT+.n166 GNDA 0.206779f
C1797 VOUT+.t24 GNDA 0.30841f
C1798 VOUT+.t123 GNDA 0.313663f
C1799 VOUT+.t25 GNDA 0.30841f
C1800 VOUT+.n167 GNDA 0.206779f
C1801 VOUT+.n168 GNDA 0.250583f
C1802 VOUT+.t48 GNDA 0.313663f
C1803 VOUT+.t152 GNDA 0.30841f
C1804 VOUT+.n169 GNDA 0.206779f
C1805 VOUT+.t126 GNDA 0.30841f
C1806 VOUT+.t80 GNDA 0.313663f
C1807 VOUT+.t127 GNDA 0.30841f
C1808 VOUT+.n170 GNDA 0.206779f
C1809 VOUT+.n171 GNDA 0.250583f
C1810 VOUT+.t149 GNDA 0.313663f
C1811 VOUT+.t117 GNDA 0.30841f
C1812 VOUT+.n172 GNDA 0.206779f
C1813 VOUT+.t91 GNDA 0.30841f
C1814 VOUT+.t38 GNDA 0.313663f
C1815 VOUT+.t93 GNDA 0.30841f
C1816 VOUT+.n173 GNDA 0.206779f
C1817 VOUT+.n174 GNDA 0.250583f
C1818 VOUT+.t142 GNDA 0.313663f
C1819 VOUT+.t53 GNDA 0.30841f
C1820 VOUT+.n175 GNDA 0.206779f
C1821 VOUT+.t49 GNDA 0.30841f
C1822 VOUT+.n176 GNDA 0.250583f
C1823 VOUT+.t72 GNDA 0.30841f
C1824 VOUT+.n177 GNDA 0.132038f
C1825 VOUT+.t115 GNDA 0.30841f
C1826 VOUT+.n178 GNDA 0.34407f
C1827 VOUT+.n179 GNDA 0.283352f
C1828 VOUT+.n180 GNDA 0.057827f
C1829 VOUT+.n181 GNDA 0.057827f
C1830 VOUT+.n183 GNDA 0.520442f
C1831 VOUT+.n184 GNDA 0.058253f
C1832 VOUT+.n185 GNDA 1.09871f
C1833 VOUT+.n186 GNDA 0.039322f
C1834 VOUT+.n188 GNDA 0.037009f
C1835 VOUT+.n189 GNDA 1.08907f
C1836 VOUT+.n191 GNDA 0.039322f
C1837 VOUT+.n192 GNDA 0.077102f
C1838 VOUT+.n193 GNDA 0.104088f
C1839 VOUT+.t7 GNDA 0.088348f
C1840 VOUT+.n194 GNDA 0.271914f
C1841 two_stage_opamp_dummy_magic_26_0.cap_res_X.t57 GNDA 0.40891f
C1842 two_stage_opamp_dummy_magic_26_0.cap_res_X.t92 GNDA 0.410391f
C1843 two_stage_opamp_dummy_magic_26_0.cap_res_X.t26 GNDA 0.40891f
C1844 two_stage_opamp_dummy_magic_26_0.cap_res_X.t62 GNDA 0.410391f
C1845 two_stage_opamp_dummy_magic_26_0.cap_res_X.t114 GNDA 0.40891f
C1846 two_stage_opamp_dummy_magic_26_0.cap_res_X.t79 GNDA 0.410391f
C1847 two_stage_opamp_dummy_magic_26_0.cap_res_X.t54 GNDA 0.40891f
C1848 two_stage_opamp_dummy_magic_26_0.cap_res_X.t87 GNDA 0.410391f
C1849 two_stage_opamp_dummy_magic_26_0.cap_res_X.t71 GNDA 0.40891f
C1850 two_stage_opamp_dummy_magic_26_0.cap_res_X.t38 GNDA 0.410391f
C1851 two_stage_opamp_dummy_magic_26_0.cap_res_X.t89 GNDA 0.40891f
C1852 two_stage_opamp_dummy_magic_26_0.cap_res_X.t130 GNDA 0.410391f
C1853 two_stage_opamp_dummy_magic_26_0.cap_res_X.t108 GNDA 0.40891f
C1854 two_stage_opamp_dummy_magic_26_0.cap_res_X.t75 GNDA 0.410391f
C1855 two_stage_opamp_dummy_magic_26_0.cap_res_X.t59 GNDA 0.40891f
C1856 two_stage_opamp_dummy_magic_26_0.cap_res_X.t91 GNDA 0.410391f
C1857 two_stage_opamp_dummy_magic_26_0.cap_res_X.t77 GNDA 0.40891f
C1858 two_stage_opamp_dummy_magic_26_0.cap_res_X.t45 GNDA 0.410391f
C1859 two_stage_opamp_dummy_magic_26_0.cap_res_X.t95 GNDA 0.40891f
C1860 two_stage_opamp_dummy_magic_26_0.cap_res_X.t133 GNDA 0.410391f
C1861 two_stage_opamp_dummy_magic_26_0.cap_res_X.t113 GNDA 0.40891f
C1862 two_stage_opamp_dummy_magic_26_0.cap_res_X.t81 GNDA 0.410391f
C1863 two_stage_opamp_dummy_magic_26_0.cap_res_X.t138 GNDA 0.40891f
C1864 two_stage_opamp_dummy_magic_26_0.cap_res_X.t35 GNDA 0.410391f
C1865 two_stage_opamp_dummy_magic_26_0.cap_res_X.t16 GNDA 0.40891f
C1866 two_stage_opamp_dummy_magic_26_0.cap_res_X.t120 GNDA 0.410391f
C1867 two_stage_opamp_dummy_magic_26_0.cap_res_X.t101 GNDA 0.40891f
C1868 two_stage_opamp_dummy_magic_26_0.cap_res_X.t1 GNDA 0.410391f
C1869 two_stage_opamp_dummy_magic_26_0.cap_res_X.t121 GNDA 0.40891f
C1870 two_stage_opamp_dummy_magic_26_0.cap_res_X.t85 GNDA 0.410391f
C1871 two_stage_opamp_dummy_magic_26_0.cap_res_X.t7 GNDA 0.40891f
C1872 two_stage_opamp_dummy_magic_26_0.cap_res_X.t43 GNDA 0.410391f
C1873 two_stage_opamp_dummy_magic_26_0.cap_res_X.t24 GNDA 0.40891f
C1874 two_stage_opamp_dummy_magic_26_0.cap_res_X.t126 GNDA 0.410391f
C1875 two_stage_opamp_dummy_magic_26_0.cap_res_X.t47 GNDA 0.40891f
C1876 two_stage_opamp_dummy_magic_26_0.cap_res_X.t80 GNDA 0.410391f
C1877 two_stage_opamp_dummy_magic_26_0.cap_res_X.t60 GNDA 0.40891f
C1878 two_stage_opamp_dummy_magic_26_0.cap_res_X.t29 GNDA 0.410391f
C1879 two_stage_opamp_dummy_magic_26_0.cap_res_X.t83 GNDA 0.40891f
C1880 two_stage_opamp_dummy_magic_26_0.cap_res_X.t117 GNDA 0.410391f
C1881 two_stage_opamp_dummy_magic_26_0.cap_res_X.t97 GNDA 0.40891f
C1882 two_stage_opamp_dummy_magic_26_0.cap_res_X.t64 GNDA 0.410391f
C1883 two_stage_opamp_dummy_magic_26_0.cap_res_X.t50 GNDA 0.40891f
C1884 two_stage_opamp_dummy_magic_26_0.cap_res_X.t84 GNDA 0.410391f
C1885 two_stage_opamp_dummy_magic_26_0.cap_res_X.t65 GNDA 0.40891f
C1886 two_stage_opamp_dummy_magic_26_0.cap_res_X.t34 GNDA 0.410391f
C1887 two_stage_opamp_dummy_magic_26_0.cap_res_X.t86 GNDA 0.40891f
C1888 two_stage_opamp_dummy_magic_26_0.cap_res_X.t123 GNDA 0.410391f
C1889 two_stage_opamp_dummy_magic_26_0.cap_res_X.t103 GNDA 0.40891f
C1890 two_stage_opamp_dummy_magic_26_0.cap_res_X.t70 GNDA 0.410391f
C1891 two_stage_opamp_dummy_magic_26_0.cap_res_X.t128 GNDA 0.40891f
C1892 two_stage_opamp_dummy_magic_26_0.cap_res_X.t25 GNDA 0.410391f
C1893 two_stage_opamp_dummy_magic_26_0.cap_res_X.t8 GNDA 0.40891f
C1894 two_stage_opamp_dummy_magic_26_0.cap_res_X.t107 GNDA 0.410391f
C1895 two_stage_opamp_dummy_magic_26_0.cap_res_X.t90 GNDA 0.40891f
C1896 two_stage_opamp_dummy_magic_26_0.cap_res_X.t129 GNDA 0.410391f
C1897 two_stage_opamp_dummy_magic_26_0.cap_res_X.t109 GNDA 0.40891f
C1898 two_stage_opamp_dummy_magic_26_0.cap_res_X.t76 GNDA 0.410391f
C1899 two_stage_opamp_dummy_magic_26_0.cap_res_X.t94 GNDA 0.40891f
C1900 two_stage_opamp_dummy_magic_26_0.cap_res_X.t48 GNDA 0.410391f
C1901 two_stage_opamp_dummy_magic_26_0.cap_res_X.t127 GNDA 0.40891f
C1902 two_stage_opamp_dummy_magic_26_0.cap_res_X.t44 GNDA 0.410391f
C1903 two_stage_opamp_dummy_magic_26_0.cap_res_X.t5 GNDA 0.40891f
C1904 two_stage_opamp_dummy_magic_26_0.cap_res_X.t42 GNDA 0.410391f
C1905 two_stage_opamp_dummy_magic_26_0.cap_res_X.t22 GNDA 0.40891f
C1906 two_stage_opamp_dummy_magic_26_0.cap_res_X.t124 GNDA 0.410391f
C1907 two_stage_opamp_dummy_magic_26_0.cap_res_X.t41 GNDA 0.40891f
C1908 two_stage_opamp_dummy_magic_26_0.cap_res_X.t72 GNDA 0.410391f
C1909 two_stage_opamp_dummy_magic_26_0.cap_res_X.t55 GNDA 0.40891f
C1910 two_stage_opamp_dummy_magic_26_0.cap_res_X.t21 GNDA 0.410391f
C1911 two_stage_opamp_dummy_magic_26_0.cap_res_X.t98 GNDA 0.40891f
C1912 two_stage_opamp_dummy_magic_26_0.cap_res_X.t137 GNDA 0.410391f
C1913 two_stage_opamp_dummy_magic_26_0.cap_res_X.t12 GNDA 0.40891f
C1914 two_stage_opamp_dummy_magic_26_0.cap_res_X.t53 GNDA 0.428959f
C1915 two_stage_opamp_dummy_magic_26_0.cap_res_X.t39 GNDA 0.40891f
C1916 two_stage_opamp_dummy_magic_26_0.cap_res_X.t78 GNDA 0.219633f
C1917 two_stage_opamp_dummy_magic_26_0.cap_res_X.n0 GNDA 0.235062f
C1918 two_stage_opamp_dummy_magic_26_0.cap_res_X.t19 GNDA 0.40891f
C1919 two_stage_opamp_dummy_magic_26_0.cap_res_X.t56 GNDA 0.219633f
C1920 two_stage_opamp_dummy_magic_26_0.cap_res_X.n1 GNDA 0.233166f
C1921 two_stage_opamp_dummy_magic_26_0.cap_res_X.t119 GNDA 0.40891f
C1922 two_stage_opamp_dummy_magic_26_0.cap_res_X.t23 GNDA 0.219633f
C1923 two_stage_opamp_dummy_magic_26_0.cap_res_X.n2 GNDA 0.233166f
C1924 two_stage_opamp_dummy_magic_26_0.cap_res_X.t4 GNDA 0.40891f
C1925 two_stage_opamp_dummy_magic_26_0.cap_res_X.t46 GNDA 0.219633f
C1926 two_stage_opamp_dummy_magic_26_0.cap_res_X.n3 GNDA 0.233166f
C1927 two_stage_opamp_dummy_magic_26_0.cap_res_X.t100 GNDA 0.40891f
C1928 two_stage_opamp_dummy_magic_26_0.cap_res_X.t6 GNDA 0.219633f
C1929 two_stage_opamp_dummy_magic_26_0.cap_res_X.n4 GNDA 0.233166f
C1930 two_stage_opamp_dummy_magic_26_0.cap_res_X.t66 GNDA 0.40891f
C1931 two_stage_opamp_dummy_magic_26_0.cap_res_X.t105 GNDA 0.219633f
C1932 two_stage_opamp_dummy_magic_26_0.cap_res_X.n5 GNDA 0.233166f
C1933 two_stage_opamp_dummy_magic_26_0.cap_res_X.t31 GNDA 0.40891f
C1934 two_stage_opamp_dummy_magic_26_0.cap_res_X.t68 GNDA 0.219633f
C1935 two_stage_opamp_dummy_magic_26_0.cap_res_X.n6 GNDA 0.233166f
C1936 two_stage_opamp_dummy_magic_26_0.cap_res_X.t51 GNDA 0.40891f
C1937 two_stage_opamp_dummy_magic_26_0.cap_res_X.t88 GNDA 0.219633f
C1938 two_stage_opamp_dummy_magic_26_0.cap_res_X.n7 GNDA 0.233166f
C1939 two_stage_opamp_dummy_magic_26_0.cap_res_X.t10 GNDA 0.40891f
C1940 two_stage_opamp_dummy_magic_26_0.cap_res_X.t52 GNDA 0.219633f
C1941 two_stage_opamp_dummy_magic_26_0.cap_res_X.n8 GNDA 0.233166f
C1942 two_stage_opamp_dummy_magic_26_0.cap_res_X.t111 GNDA 0.40891f
C1943 two_stage_opamp_dummy_magic_26_0.cap_res_X.t14 GNDA 0.219633f
C1944 two_stage_opamp_dummy_magic_26_0.cap_res_X.n9 GNDA 0.233166f
C1945 two_stage_opamp_dummy_magic_26_0.cap_res_X.t61 GNDA 0.40891f
C1946 two_stage_opamp_dummy_magic_26_0.cap_res_X.t93 GNDA 0.410391f
C1947 two_stage_opamp_dummy_magic_26_0.cap_res_X.t135 GNDA 0.197688f
C1948 two_stage_opamp_dummy_magic_26_0.cap_res_X.n10 GNDA 0.254989f
C1949 two_stage_opamp_dummy_magic_26_0.cap_res_X.t40 GNDA 0.218274f
C1950 two_stage_opamp_dummy_magic_26_0.cap_res_X.n11 GNDA 0.276934f
C1951 two_stage_opamp_dummy_magic_26_0.cap_res_X.t106 GNDA 0.218274f
C1952 two_stage_opamp_dummy_magic_26_0.cap_res_X.n12 GNDA 0.297397f
C1953 two_stage_opamp_dummy_magic_26_0.cap_res_X.t73 GNDA 0.218274f
C1954 two_stage_opamp_dummy_magic_26_0.cap_res_X.n13 GNDA 0.297397f
C1955 two_stage_opamp_dummy_magic_26_0.cap_res_X.t136 GNDA 0.218274f
C1956 two_stage_opamp_dummy_magic_26_0.cap_res_X.n14 GNDA 0.297397f
C1957 two_stage_opamp_dummy_magic_26_0.cap_res_X.t28 GNDA 0.218274f
C1958 two_stage_opamp_dummy_magic_26_0.cap_res_X.n15 GNDA 0.297397f
C1959 two_stage_opamp_dummy_magic_26_0.cap_res_X.t58 GNDA 0.218274f
C1960 two_stage_opamp_dummy_magic_26_0.cap_res_X.n16 GNDA 0.297397f
C1961 two_stage_opamp_dummy_magic_26_0.cap_res_X.t20 GNDA 0.218274f
C1962 two_stage_opamp_dummy_magic_26_0.cap_res_X.n17 GNDA 0.297397f
C1963 two_stage_opamp_dummy_magic_26_0.cap_res_X.t118 GNDA 0.218274f
C1964 two_stage_opamp_dummy_magic_26_0.cap_res_X.n18 GNDA 0.297397f
C1965 two_stage_opamp_dummy_magic_26_0.cap_res_X.t15 GNDA 0.218274f
C1966 two_stage_opamp_dummy_magic_26_0.cap_res_X.n19 GNDA 0.297397f
C1967 two_stage_opamp_dummy_magic_26_0.cap_res_X.t112 GNDA 0.218274f
C1968 two_stage_opamp_dummy_magic_26_0.cap_res_X.n20 GNDA 0.297397f
C1969 two_stage_opamp_dummy_magic_26_0.cap_res_X.t74 GNDA 0.218274f
C1970 two_stage_opamp_dummy_magic_26_0.cap_res_X.n21 GNDA 0.297397f
C1971 two_stage_opamp_dummy_magic_26_0.cap_res_X.t37 GNDA 0.218274f
C1972 two_stage_opamp_dummy_magic_26_0.cap_res_X.n22 GNDA 0.297397f
C1973 two_stage_opamp_dummy_magic_26_0.cap_res_X.t69 GNDA 0.218274f
C1974 two_stage_opamp_dummy_magic_26_0.cap_res_X.n23 GNDA 0.297397f
C1975 two_stage_opamp_dummy_magic_26_0.cap_res_X.t32 GNDA 0.218274f
C1976 two_stage_opamp_dummy_magic_26_0.cap_res_X.n24 GNDA 0.297397f
C1977 two_stage_opamp_dummy_magic_26_0.cap_res_X.t131 GNDA 0.218274f
C1978 two_stage_opamp_dummy_magic_26_0.cap_res_X.n25 GNDA 0.297397f
C1979 two_stage_opamp_dummy_magic_26_0.cap_res_X.t27 GNDA 0.218274f
C1980 two_stage_opamp_dummy_magic_26_0.cap_res_X.n26 GNDA 0.297397f
C1981 two_stage_opamp_dummy_magic_26_0.cap_res_X.t125 GNDA 0.218274f
C1982 two_stage_opamp_dummy_magic_26_0.cap_res_X.n27 GNDA 0.297397f
C1983 two_stage_opamp_dummy_magic_26_0.cap_res_X.t96 GNDA 0.218274f
C1984 two_stage_opamp_dummy_magic_26_0.cap_res_X.n28 GNDA 0.297397f
C1985 two_stage_opamp_dummy_magic_26_0.cap_res_X.t134 GNDA 0.218274f
C1986 two_stage_opamp_dummy_magic_26_0.cap_res_X.n29 GNDA 0.259462f
C1987 two_stage_opamp_dummy_magic_26_0.cap_res_X.t110 GNDA 0.410391f
C1988 two_stage_opamp_dummy_magic_26_0.cap_res_X.t9 GNDA 0.410391f
C1989 two_stage_opamp_dummy_magic_26_0.cap_res_X.t102 GNDA 0.40891f
C1990 two_stage_opamp_dummy_magic_26_0.cap_res_X.t13 GNDA 0.430855f
C1991 two_stage_opamp_dummy_magic_26_0.cap_res_X.t49 GNDA 0.219633f
C1992 two_stage_opamp_dummy_magic_26_0.cap_res_X.n30 GNDA 0.253629f
C1993 two_stage_opamp_dummy_magic_26_0.cap_res_X.t115 GNDA 0.40891f
C1994 two_stage_opamp_dummy_magic_26_0.cap_res_X.t11 GNDA 0.428959f
C1995 two_stage_opamp_dummy_magic_26_0.cap_res_X.t2 GNDA 0.40891f
C1996 two_stage_opamp_dummy_magic_26_0.cap_res_X.t36 GNDA 0.219633f
C1997 two_stage_opamp_dummy_magic_26_0.cap_res_X.n31 GNDA 0.235062f
C1998 two_stage_opamp_dummy_magic_26_0.cap_res_X.t122 GNDA 0.40891f
C1999 two_stage_opamp_dummy_magic_26_0.cap_res_X.t18 GNDA 0.219633f
C2000 two_stage_opamp_dummy_magic_26_0.cap_res_X.n32 GNDA 0.233166f
C2001 two_stage_opamp_dummy_magic_26_0.cap_res_X.t82 GNDA 0.40891f
C2002 two_stage_opamp_dummy_magic_26_0.cap_res_X.t116 GNDA 0.219633f
C2003 two_stage_opamp_dummy_magic_26_0.cap_res_X.n33 GNDA 0.233166f
C2004 two_stage_opamp_dummy_magic_26_0.cap_res_X.t104 GNDA 0.40891f
C2005 two_stage_opamp_dummy_magic_26_0.cap_res_X.t3 GNDA 0.219633f
C2006 two_stage_opamp_dummy_magic_26_0.cap_res_X.n34 GNDA 0.233166f
C2007 two_stage_opamp_dummy_magic_26_0.cap_res_X.t67 GNDA 0.40891f
C2008 two_stage_opamp_dummy_magic_26_0.cap_res_X.t99 GNDA 0.219633f
C2009 two_stage_opamp_dummy_magic_26_0.cap_res_X.n35 GNDA 0.233166f
C2010 two_stage_opamp_dummy_magic_26_0.cap_res_X.t33 GNDA 0.40891f
C2011 two_stage_opamp_dummy_magic_26_0.cap_res_X.t63 GNDA 0.219633f
C2012 two_stage_opamp_dummy_magic_26_0.cap_res_X.n36 GNDA 0.233166f
C2013 two_stage_opamp_dummy_magic_26_0.cap_res_X.n37 GNDA 0.233166f
C2014 two_stage_opamp_dummy_magic_26_0.cap_res_X.t30 GNDA 0.219633f
C2015 two_stage_opamp_dummy_magic_26_0.cap_res_X.t132 GNDA 0.430855f
C2016 two_stage_opamp_dummy_magic_26_0.cap_res_X.t17 GNDA 0.517753f
C2017 two_stage_opamp_dummy_magic_26_0.cap_res_X.t0 GNDA 0.362088f
C2018 VOUT-.n1 GNDA 0.077013f
C2019 VOUT-.n4 GNDA 0.05776f
C2020 VOUT-.n5 GNDA 0.096267f
C2021 VOUT-.n6 GNDA 0.05776f
C2022 VOUT-.n7 GNDA 0.05776f
C2023 VOUT-.n9 GNDA 0.039277f
C2024 VOUT-.n11 GNDA 0.039277f
C2025 VOUT-.n13 GNDA 0.077013f
C2026 VOUT-.n14 GNDA 0.039277f
C2027 VOUT-.n16 GNDA 0.039277f
C2028 VOUT-.n18 GNDA 0.050829f
C2029 VOUT-.n19 GNDA 0.073334f
C2030 VOUT-.n20 GNDA 0.071366f
C2031 VOUT-.n21 GNDA 0.050829f
C2032 VOUT-.n22 GNDA 0.050829f
C2033 VOUT-.n23 GNDA 0.071366f
C2034 VOUT-.n24 GNDA 0.071366f
C2035 VOUT-.n25 GNDA 0.050829f
C2036 VOUT-.n26 GNDA 0.081373f
C2037 VOUT-.t16 GNDA 0.046208f
C2038 VOUT-.t9 GNDA 0.046208f
C2039 VOUT-.n27 GNDA 0.09468f
C2040 VOUT-.n28 GNDA 0.244397f
C2041 VOUT-.t13 GNDA 0.046208f
C2042 VOUT-.t7 GNDA 0.046208f
C2043 VOUT-.n29 GNDA 0.09468f
C2044 VOUT-.n30 GNDA 0.241934f
C2045 VOUT-.n31 GNDA 0.058758f
C2046 VOUT-.t14 GNDA 0.046208f
C2047 VOUT-.t8 GNDA 0.046208f
C2048 VOUT-.n32 GNDA 0.09468f
C2049 VOUT-.n33 GNDA 0.241934f
C2050 VOUT-.n34 GNDA 0.033306f
C2051 VOUT-.t12 GNDA 0.046208f
C2052 VOUT-.t6 GNDA 0.046208f
C2053 VOUT-.n35 GNDA 0.09468f
C2054 VOUT-.n36 GNDA 0.241934f
C2055 VOUT-.n37 GNDA 0.033306f
C2056 VOUT-.t10 GNDA 0.046208f
C2057 VOUT-.t17 GNDA 0.046208f
C2058 VOUT-.n38 GNDA 0.09468f
C2059 VOUT-.n39 GNDA 0.244397f
C2060 VOUT-.n40 GNDA 0.058758f
C2061 VOUT-.t11 GNDA 0.046208f
C2062 VOUT-.t5 GNDA 0.046208f
C2063 VOUT-.n41 GNDA 0.09468f
C2064 VOUT-.n42 GNDA 0.241934f
C2065 VOUT-.n43 GNDA 0.038849f
C2066 VOUT-.n44 GNDA 0.023104f
C2067 VOUT-.n45 GNDA 0.023104f
C2068 VOUT-.n46 GNDA 0.038849f
C2069 VOUT-.n47 GNDA 0.071366f
C2070 VOUT-.n48 GNDA 0.099897f
C2071 VOUT-.n49 GNDA 0.124477f
C2072 VOUT-.n50 GNDA 0.174217f
C2073 VOUT-.n51 GNDA 0.050829f
C2074 VOUT-.n52 GNDA 0.083174f
C2075 VOUT-.n53 GNDA 0.050829f
C2076 VOUT-.n54 GNDA 0.083174f
C2077 VOUT-.n55 GNDA 0.050829f
C2078 VOUT-.n56 GNDA 0.050829f
C2079 VOUT-.n57 GNDA 0.050829f
C2080 VOUT-.n58 GNDA 0.083174f
C2081 VOUT-.n59 GNDA 0.050829f
C2082 VOUT-.n60 GNDA 0.076243f
C2083 VOUT-.n61 GNDA 0.244902f
C2084 VOUT-.n62 GNDA 0.237971f
C2085 VOUT-.n64 GNDA 0.077013f
C2086 VOUT-.n65 GNDA 0.036966f
C2087 VOUT-.n66 GNDA 0.510213f
C2088 VOUT-.n69 GNDA 0.05776f
C2089 VOUT-.n70 GNDA 0.05776f
C2090 VOUT-.t96 GNDA 0.3133f
C2091 VOUT-.t64 GNDA 0.308053f
C2092 VOUT-.n71 GNDA 0.20654f
C2093 VOUT-.t22 GNDA 0.308053f
C2094 VOUT-.n72 GNDA 0.134773f
C2095 VOUT-.t59 GNDA 0.3133f
C2096 VOUT-.t20 GNDA 0.308053f
C2097 VOUT-.n73 GNDA 0.20654f
C2098 VOUT-.t117 GNDA 0.308053f
C2099 VOUT-.t46 GNDA 0.312643f
C2100 VOUT-.t147 GNDA 0.312643f
C2101 VOUT-.t106 GNDA 0.312643f
C2102 VOUT-.t126 GNDA 0.312643f
C2103 VOUT-.t91 GNDA 0.312643f
C2104 VOUT-.t57 GNDA 0.312643f
C2105 VOUT-.t153 GNDA 0.312643f
C2106 VOUT-.t38 GNDA 0.312643f
C2107 VOUT-.t138 GNDA 0.312643f
C2108 VOUT-.t118 GNDA 0.312643f
C2109 VOUT-.t145 GNDA 0.312643f
C2110 VOUT-.t104 GNDA 0.308053f
C2111 VOUT-.n74 GNDA 0.207197f
C2112 VOUT-.t79 GNDA 0.308053f
C2113 VOUT-.n75 GNDA 0.264956f
C2114 VOUT-.t101 GNDA 0.308053f
C2115 VOUT-.n76 GNDA 0.264956f
C2116 VOUT-.t134 GNDA 0.308053f
C2117 VOUT-.n77 GNDA 0.264956f
C2118 VOUT-.t111 GNDA 0.308053f
C2119 VOUT-.n78 GNDA 0.264956f
C2120 VOUT-.t151 GNDA 0.308053f
C2121 VOUT-.n79 GNDA 0.264956f
C2122 VOUT-.t52 GNDA 0.308053f
C2123 VOUT-.n80 GNDA 0.264956f
C2124 VOUT-.t89 GNDA 0.308053f
C2125 VOUT-.n81 GNDA 0.264956f
C2126 VOUT-.t69 GNDA 0.308053f
C2127 VOUT-.n82 GNDA 0.264956f
C2128 VOUT-.t105 GNDA 0.308053f
C2129 VOUT-.n83 GNDA 0.264956f
C2130 VOUT-.t143 GNDA 0.308053f
C2131 VOUT-.n84 GNDA 0.264956f
C2132 VOUT-.n85 GNDA 0.250293f
C2133 VOUT-.t116 GNDA 0.3133f
C2134 VOUT-.t85 GNDA 0.308053f
C2135 VOUT-.n86 GNDA 0.20654f
C2136 VOUT-.t51 GNDA 0.308053f
C2137 VOUT-.t102 GNDA 0.3133f
C2138 VOUT-.t136 GNDA 0.308053f
C2139 VOUT-.n87 GNDA 0.20654f
C2140 VOUT-.n88 GNDA 0.250293f
C2141 VOUT-.t152 GNDA 0.3133f
C2142 VOUT-.t115 GNDA 0.308053f
C2143 VOUT-.n89 GNDA 0.20654f
C2144 VOUT-.t84 GNDA 0.308053f
C2145 VOUT-.t135 GNDA 0.3133f
C2146 VOUT-.t33 GNDA 0.308053f
C2147 VOUT-.n90 GNDA 0.20654f
C2148 VOUT-.n91 GNDA 0.250293f
C2149 VOUT-.t63 GNDA 0.3133f
C2150 VOUT-.t109 GNDA 0.308053f
C2151 VOUT-.n92 GNDA 0.20654f
C2152 VOUT-.t21 GNDA 0.308053f
C2153 VOUT-.t30 GNDA 0.3133f
C2154 VOUT-.t113 GNDA 0.308053f
C2155 VOUT-.n93 GNDA 0.20654f
C2156 VOUT-.n94 GNDA 0.250293f
C2157 VOUT-.t67 GNDA 0.3133f
C2158 VOUT-.t28 GNDA 0.308053f
C2159 VOUT-.n95 GNDA 0.20654f
C2160 VOUT-.t129 GNDA 0.308053f
C2161 VOUT-.t48 GNDA 0.3133f
C2162 VOUT-.t81 GNDA 0.308053f
C2163 VOUT-.n96 GNDA 0.20654f
C2164 VOUT-.n97 GNDA 0.250293f
C2165 VOUT-.t29 GNDA 0.3133f
C2166 VOUT-.t132 GNDA 0.308053f
C2167 VOUT-.n98 GNDA 0.20654f
C2168 VOUT-.t99 GNDA 0.308053f
C2169 VOUT-.t149 GNDA 0.3133f
C2170 VOUT-.t50 GNDA 0.308053f
C2171 VOUT-.n99 GNDA 0.20654f
C2172 VOUT-.n100 GNDA 0.250293f
C2173 VOUT-.t71 GNDA 0.3133f
C2174 VOUT-.t34 GNDA 0.308053f
C2175 VOUT-.n101 GNDA 0.20654f
C2176 VOUT-.t137 GNDA 0.308053f
C2177 VOUT-.t54 GNDA 0.3133f
C2178 VOUT-.t87 GNDA 0.308053f
C2179 VOUT-.n102 GNDA 0.20654f
C2180 VOUT-.n103 GNDA 0.250293f
C2181 VOUT-.t107 GNDA 0.3133f
C2182 VOUT-.t73 GNDA 0.308053f
C2183 VOUT-.n104 GNDA 0.20654f
C2184 VOUT-.t39 GNDA 0.308053f
C2185 VOUT-.t92 GNDA 0.3133f
C2186 VOUT-.t123 GNDA 0.308053f
C2187 VOUT-.n105 GNDA 0.20654f
C2188 VOUT-.n106 GNDA 0.250293f
C2189 VOUT-.t100 GNDA 0.3133f
C2190 VOUT-.t65 GNDA 0.308053f
C2191 VOUT-.n107 GNDA 0.20654f
C2192 VOUT-.t23 GNDA 0.308053f
C2193 VOUT-.t55 GNDA 0.3133f
C2194 VOUT-.t144 GNDA 0.308053f
C2195 VOUT-.n108 GNDA 0.201726f
C2196 VOUT-.t140 GNDA 0.3133f
C2197 VOUT-.t25 GNDA 0.308053f
C2198 VOUT-.n109 GNDA 0.201726f
C2199 VOUT-.t124 GNDA 0.312643f
C2200 VOUT-.t90 GNDA 0.312643f
C2201 VOUT-.t53 GNDA 0.312648f
C2202 VOUT-.t75 GNDA 0.312901f
C2203 VOUT-.t35 GNDA 0.312643f
C2204 VOUT-.t155 GNDA 0.312648f
C2205 VOUT-.t42 GNDA 0.312901f
C2206 VOUT-.t146 GNDA 0.308053f
C2207 VOUT-.n110 GNDA 0.210789f
C2208 VOUT-.t121 GNDA 0.308053f
C2209 VOUT-.n111 GNDA 0.264951f
C2210 VOUT-.t139 GNDA 0.308053f
C2211 VOUT-.n112 GNDA 0.264956f
C2212 VOUT-.t41 GNDA 0.308053f
C2213 VOUT-.n113 GNDA 0.268549f
C2214 VOUT-.t154 GNDA 0.308053f
C2215 VOUT-.n114 GNDA 0.264951f
C2216 VOUT-.t58 GNDA 0.308053f
C2217 VOUT-.n115 GNDA 0.264956f
C2218 VOUT-.t94 GNDA 0.308053f
C2219 VOUT-.n116 GNDA 0.264956f
C2220 VOUT-.t127 GNDA 0.308053f
C2221 VOUT-.n117 GNDA 0.197347f
C2222 VOUT-.t108 GNDA 0.308053f
C2223 VOUT-.n118 GNDA 0.197347f
C2224 VOUT-.t148 GNDA 0.308053f
C2225 VOUT-.n119 GNDA 0.134773f
C2226 VOUT-.t47 GNDA 0.308053f
C2227 VOUT-.n120 GNDA 0.134773f
C2228 VOUT-.n121 GNDA 0.1444f
C2229 VOUT-.t131 GNDA 0.3133f
C2230 VOUT-.t95 GNDA 0.308053f
C2231 VOUT-.n122 GNDA 0.20654f
C2232 VOUT-.t61 GNDA 0.308053f
C2233 VOUT-.t43 GNDA 0.3133f
C2234 VOUT-.t78 GNDA 0.308053f
C2235 VOUT-.n123 GNDA 0.20654f
C2236 VOUT-.n124 GNDA 0.250293f
C2237 VOUT-.t103 GNDA 0.3133f
C2238 VOUT-.t70 GNDA 0.308053f
C2239 VOUT-.n125 GNDA 0.20654f
C2240 VOUT-.t32 GNDA 0.308053f
C2241 VOUT-.t86 GNDA 0.3133f
C2242 VOUT-.t119 GNDA 0.308053f
C2243 VOUT-.n126 GNDA 0.20654f
C2244 VOUT-.n127 GNDA 0.250293f
C2245 VOUT-.t68 GNDA 0.3133f
C2246 VOUT-.t27 GNDA 0.308053f
C2247 VOUT-.n128 GNDA 0.20654f
C2248 VOUT-.t130 GNDA 0.308053f
C2249 VOUT-.t49 GNDA 0.3133f
C2250 VOUT-.t82 GNDA 0.308053f
C2251 VOUT-.n129 GNDA 0.20654f
C2252 VOUT-.n130 GNDA 0.250293f
C2253 VOUT-.t98 GNDA 0.3133f
C2254 VOUT-.t66 GNDA 0.308053f
C2255 VOUT-.n131 GNDA 0.20654f
C2256 VOUT-.t26 GNDA 0.308053f
C2257 VOUT-.t80 GNDA 0.3133f
C2258 VOUT-.t112 GNDA 0.308053f
C2259 VOUT-.n132 GNDA 0.20654f
C2260 VOUT-.n133 GNDA 0.250293f
C2261 VOUT-.t62 GNDA 0.3133f
C2262 VOUT-.t24 GNDA 0.308053f
C2263 VOUT-.n134 GNDA 0.20654f
C2264 VOUT-.t125 GNDA 0.308053f
C2265 VOUT-.t44 GNDA 0.3133f
C2266 VOUT-.t76 GNDA 0.308053f
C2267 VOUT-.n135 GNDA 0.20654f
C2268 VOUT-.n136 GNDA 0.250293f
C2269 VOUT-.t19 GNDA 0.3133f
C2270 VOUT-.t122 GNDA 0.308053f
C2271 VOUT-.n137 GNDA 0.20654f
C2272 VOUT-.t88 GNDA 0.308053f
C2273 VOUT-.t141 GNDA 0.3133f
C2274 VOUT-.t37 GNDA 0.308053f
C2275 VOUT-.n138 GNDA 0.20654f
C2276 VOUT-.n139 GNDA 0.250293f
C2277 VOUT-.t56 GNDA 0.3133f
C2278 VOUT-.t156 GNDA 0.308053f
C2279 VOUT-.n140 GNDA 0.20654f
C2280 VOUT-.t120 GNDA 0.308053f
C2281 VOUT-.t36 GNDA 0.3133f
C2282 VOUT-.t72 GNDA 0.308053f
C2283 VOUT-.n141 GNDA 0.20654f
C2284 VOUT-.n142 GNDA 0.250293f
C2285 VOUT-.t150 GNDA 0.3133f
C2286 VOUT-.t114 GNDA 0.308053f
C2287 VOUT-.n143 GNDA 0.20654f
C2288 VOUT-.t83 GNDA 0.308053f
C2289 VOUT-.t133 GNDA 0.3133f
C2290 VOUT-.t31 GNDA 0.308053f
C2291 VOUT-.n144 GNDA 0.20654f
C2292 VOUT-.n145 GNDA 0.250293f
C2293 VOUT-.t110 GNDA 0.3133f
C2294 VOUT-.t77 GNDA 0.308053f
C2295 VOUT-.n146 GNDA 0.20654f
C2296 VOUT-.t45 GNDA 0.308053f
C2297 VOUT-.t97 GNDA 0.3133f
C2298 VOUT-.t128 GNDA 0.308053f
C2299 VOUT-.n147 GNDA 0.20654f
C2300 VOUT-.n148 GNDA 0.250293f
C2301 VOUT-.t74 GNDA 0.3133f
C2302 VOUT-.t40 GNDA 0.308053f
C2303 VOUT-.n149 GNDA 0.20654f
C2304 VOUT-.t142 GNDA 0.308053f
C2305 VOUT-.n150 GNDA 0.250293f
C2306 VOUT-.t93 GNDA 0.308053f
C2307 VOUT-.n151 GNDA 0.131389f
C2308 VOUT-.t60 GNDA 0.308053f
C2309 VOUT-.n152 GNDA 0.348018f
C2310 VOUT-.n153 GNDA 0.283024f
C2311 VOUT-.n154 GNDA 0.05776f
C2312 VOUT-.n155 GNDA 0.05776f
C2313 VOUT-.n156 GNDA 0.05776f
C2314 VOUT-.n157 GNDA 0.169419f
C2315 VOUT-.n158 GNDA 0.061194f
C2316 VOUT-.n159 GNDA 0.058186f
C2317 VOUT-.n161 GNDA 0.51984f
C2318 VOUT-.n162 GNDA 0.05776f
C2319 VOUT-.n163 GNDA 1.09744f
C2320 VOUT-.n167 GNDA 0.039277f
C2321 VOUT-.n168 GNDA 0.039277f
C2322 VOUT-.n169 GNDA 0.036966f
C2323 VOUT-.n170 GNDA 0.077013f
C2324 VOUT-.n171 GNDA 0.039277f
C2325 VOUT-.n172 GNDA 0.039277f
C2326 VOUT-.n174 GNDA 1.08781f
C2327 VOUT-.n175 GNDA 0.103968f
C2328 VOUT-.t1 GNDA 0.088245f
C2329 VOUT-.n176 GNDA 0.271599f
C2330 VOUT-.n177 GNDA 0.036966f
C2331 VOUT-.t3 GNDA 0.053909f
C2332 VOUT-.t4 GNDA 0.053909f
C2333 VOUT-.n178 GNDA 0.11583f
C2334 VOUT-.n179 GNDA 0.284346f
C2335 VOUT-.n180 GNDA 0.036966f
C2336 VOUT-.n181 GNDA 0.245261f
C2337 VOUT-.t0 GNDA 0.053909f
C2338 VOUT-.t2 GNDA 0.053909f
C2339 VOUT-.n182 GNDA 0.11583f
C2340 VOUT-.n183 GNDA 0.293311f
C2341 VOUT-.n184 GNDA 0.16479f
C2342 VOUT-.t15 GNDA 0.053909f
C2343 VOUT-.t18 GNDA 0.053909f
C2344 VOUT-.n185 GNDA 0.11583f
C2345 VOUT-.n186 GNDA 0.279659f
C2346 VOUT-.n187 GNDA 0.131468f
C2347 VOUT-.n188 GNDA 0.036966f
C2348 VOUT-.n189 GNDA 0.19075f
C2349 VOUT-.n190 GNDA 0.036966f
C2350 VOUT-.n191 GNDA 0.036966f
C2351 VOUT-.n192 GNDA 0.036966f
C2352 VOUT-.n193 GNDA 0.036966f
C2353 VOUT-.n194 GNDA 0.084907f
C2354 VOUT-.n195 GNDA 0.099347f
C2355 two_stage_opamp_dummy_magic_26_0.VD1.t14 GNDA 0.03895f
C2356 two_stage_opamp_dummy_magic_26_0.VD1.t11 GNDA 0.03895f
C2357 two_stage_opamp_dummy_magic_26_0.VD1.n0 GNDA 0.086232f
C2358 two_stage_opamp_dummy_magic_26_0.VD1.n1 GNDA 0.502457f
C2359 two_stage_opamp_dummy_magic_26_0.VD1.n2 GNDA 0.058446f
C2360 two_stage_opamp_dummy_magic_26_0.VD1.n3 GNDA 0.153053f
C2361 two_stage_opamp_dummy_magic_26_0.VD1.t0 GNDA 0.03895f
C2362 two_stage_opamp_dummy_magic_26_0.VD1.t8 GNDA 0.03895f
C2363 two_stage_opamp_dummy_magic_26_0.VD1.n4 GNDA 0.084751f
C2364 two_stage_opamp_dummy_magic_26_0.VD1.n5 GNDA 0.326538f
C2365 two_stage_opamp_dummy_magic_26_0.VD1.n6 GNDA 0.082835f
C2366 two_stage_opamp_dummy_magic_26_0.VD1.t4 GNDA 0.03895f
C2367 two_stage_opamp_dummy_magic_26_0.VD1.t6 GNDA 0.03895f
C2368 two_stage_opamp_dummy_magic_26_0.VD1.n7 GNDA 0.084751f
C2369 two_stage_opamp_dummy_magic_26_0.VD1.n8 GNDA 0.335643f
C2370 two_stage_opamp_dummy_magic_26_0.VD1.t13 GNDA 0.03895f
C2371 two_stage_opamp_dummy_magic_26_0.VD1.t18 GNDA 0.03895f
C2372 two_stage_opamp_dummy_magic_26_0.VD1.n9 GNDA 0.086232f
C2373 two_stage_opamp_dummy_magic_26_0.VD1.t17 GNDA 0.03895f
C2374 two_stage_opamp_dummy_magic_26_0.VD1.t12 GNDA 0.03895f
C2375 two_stage_opamp_dummy_magic_26_0.VD1.n10 GNDA 0.086232f
C2376 two_stage_opamp_dummy_magic_26_0.VD1.n11 GNDA 0.690983f
C2377 two_stage_opamp_dummy_magic_26_0.VD1.t16 GNDA 0.03895f
C2378 two_stage_opamp_dummy_magic_26_0.VD1.t10 GNDA 0.03895f
C2379 two_stage_opamp_dummy_magic_26_0.VD1.n12 GNDA 0.086232f
C2380 two_stage_opamp_dummy_magic_26_0.VD1.n13 GNDA 0.205447f
C2381 two_stage_opamp_dummy_magic_26_0.VD1.t5 GNDA 0.03895f
C2382 two_stage_opamp_dummy_magic_26_0.VD1.t20 GNDA 0.03895f
C2383 two_stage_opamp_dummy_magic_26_0.VD1.n14 GNDA 0.084751f
C2384 two_stage_opamp_dummy_magic_26_0.VD1.n15 GNDA 0.335643f
C2385 two_stage_opamp_dummy_magic_26_0.VD1.n16 GNDA 0.140805f
C2386 two_stage_opamp_dummy_magic_26_0.VD1.t3 GNDA 0.03895f
C2387 two_stage_opamp_dummy_magic_26_0.VD1.t7 GNDA 0.03895f
C2388 two_stage_opamp_dummy_magic_26_0.VD1.n17 GNDA 0.084751f
C2389 two_stage_opamp_dummy_magic_26_0.VD1.n18 GNDA 0.326538f
C2390 two_stage_opamp_dummy_magic_26_0.VD1.n19 GNDA 0.058446f
C2391 two_stage_opamp_dummy_magic_26_0.VD1.n20 GNDA 0.153053f
C2392 two_stage_opamp_dummy_magic_26_0.VD1.n21 GNDA 0.684347f
C2393 two_stage_opamp_dummy_magic_26_0.VD1.n22 GNDA 0.130987f
C2394 two_stage_opamp_dummy_magic_26_0.VD1.n23 GNDA 0.0779f
C2395 two_stage_opamp_dummy_magic_26_0.VD1.t15 GNDA 0.03895f
C2396 two_stage_opamp_dummy_magic_26_0.VD1.t9 GNDA 0.03895f
C2397 two_stage_opamp_dummy_magic_26_0.VD1.n24 GNDA 0.086232f
C2398 two_stage_opamp_dummy_magic_26_0.VD1.n25 GNDA 0.684347f
C2399 two_stage_opamp_dummy_magic_26_0.VD1.n26 GNDA 0.130987f
C2400 two_stage_opamp_dummy_magic_26_0.VD1.n27 GNDA 0.690983f
C2401 two_stage_opamp_dummy_magic_26_0.VD1.n28 GNDA 0.205447f
C2402 two_stage_opamp_dummy_magic_26_0.VD1.n29 GNDA 0.058446f
C2403 two_stage_opamp_dummy_magic_26_0.VD1.t21 GNDA 0.03895f
C2404 two_stage_opamp_dummy_magic_26_0.VD1.t1 GNDA 0.03895f
C2405 two_stage_opamp_dummy_magic_26_0.VD1.n30 GNDA 0.084751f
C2406 two_stage_opamp_dummy_magic_26_0.VD1.n31 GNDA 0.326538f
C2407 two_stage_opamp_dummy_magic_26_0.VD1.n32 GNDA 0.140805f
C2408 two_stage_opamp_dummy_magic_26_0.VD1.n33 GNDA 0.082835f
C2409 two_stage_opamp_dummy_magic_26_0.VD1.t19 GNDA 0.03895f
C2410 two_stage_opamp_dummy_magic_26_0.VD1.t2 GNDA 0.03895f
C2411 two_stage_opamp_dummy_magic_26_0.VD1.n34 GNDA 0.084751f
C2412 two_stage_opamp_dummy_magic_26_0.VD1.n35 GNDA 0.326538f
C2413 two_stage_opamp_dummy_magic_26_0.VD1.n36 GNDA 0.058446f
C2414 two_stage_opamp_dummy_magic_26_0.VD1.n37 GNDA 0.045235f
C2415 two_stage_opamp_dummy_magic_26_0.X.n0 GNDA 0.075231f
C2416 two_stage_opamp_dummy_magic_26_0.X.n1 GNDA 0.110339f
C2417 two_stage_opamp_dummy_magic_26_0.X.n2 GNDA 0.364545f
C2418 two_stage_opamp_dummy_magic_26_0.X.n3 GNDA 0.354185f
C2419 two_stage_opamp_dummy_magic_26_0.X.n4 GNDA 0.110339f
C2420 two_stage_opamp_dummy_magic_26_0.X.n5 GNDA 0.110339f
C2421 two_stage_opamp_dummy_magic_26_0.X.n7 GNDA 0.080247f
C2422 two_stage_opamp_dummy_magic_26_0.X.n8 GNDA 0.090217f
C2423 two_stage_opamp_dummy_magic_26_0.X.n9 GNDA 0.090217f
C2424 two_stage_opamp_dummy_magic_26_0.X.t23 GNDA 0.058513f
C2425 two_stage_opamp_dummy_magic_26_0.X.t24 GNDA 0.058513f
C2426 two_stage_opamp_dummy_magic_26_0.X.n10 GNDA 0.119695f
C2427 two_stage_opamp_dummy_magic_26_0.X.n11 GNDA 0.385354f
C2428 two_stage_opamp_dummy_magic_26_0.X.n12 GNDA 0.149485f
C2429 two_stage_opamp_dummy_magic_26_0.X.t6 GNDA 0.058513f
C2430 two_stage_opamp_dummy_magic_26_0.X.t1 GNDA 0.058513f
C2431 two_stage_opamp_dummy_magic_26_0.X.n13 GNDA 0.119695f
C2432 two_stage_opamp_dummy_magic_26_0.X.n14 GNDA 0.376954f
C2433 two_stage_opamp_dummy_magic_26_0.X.n15 GNDA 0.149485f
C2434 two_stage_opamp_dummy_magic_26_0.X.t0 GNDA 0.058513f
C2435 two_stage_opamp_dummy_magic_26_0.X.t20 GNDA 0.058513f
C2436 two_stage_opamp_dummy_magic_26_0.X.n16 GNDA 0.119695f
C2437 two_stage_opamp_dummy_magic_26_0.X.n17 GNDA 0.376954f
C2438 two_stage_opamp_dummy_magic_26_0.X.n18 GNDA 0.090217f
C2439 two_stage_opamp_dummy_magic_26_0.X.n19 GNDA 0.090217f
C2440 two_stage_opamp_dummy_magic_26_0.X.t5 GNDA 0.058513f
C2441 two_stage_opamp_dummy_magic_26_0.X.t21 GNDA 0.058513f
C2442 two_stage_opamp_dummy_magic_26_0.X.n20 GNDA 0.119695f
C2443 two_stage_opamp_dummy_magic_26_0.X.n21 GNDA 0.376954f
C2444 two_stage_opamp_dummy_magic_26_0.X.n22 GNDA 0.090217f
C2445 two_stage_opamp_dummy_magic_26_0.X.t8 GNDA 0.058513f
C2446 two_stage_opamp_dummy_magic_26_0.X.t19 GNDA 0.058513f
C2447 two_stage_opamp_dummy_magic_26_0.X.n23 GNDA 0.119695f
C2448 two_stage_opamp_dummy_magic_26_0.X.n24 GNDA 0.376954f
C2449 two_stage_opamp_dummy_magic_26_0.X.n25 GNDA 0.149485f
C2450 two_stage_opamp_dummy_magic_26_0.X.t22 GNDA 0.058513f
C2451 two_stage_opamp_dummy_magic_26_0.X.t7 GNDA 0.058513f
C2452 two_stage_opamp_dummy_magic_26_0.X.n26 GNDA 0.119695f
C2453 two_stage_opamp_dummy_magic_26_0.X.n27 GNDA 0.381154f
C2454 two_stage_opamp_dummy_magic_26_0.X.n28 GNDA 0.238369f
C2455 two_stage_opamp_dummy_magic_26_0.X.n29 GNDA 0.080247f
C2456 two_stage_opamp_dummy_magic_26_0.X.n31 GNDA 0.080247f
C2457 two_stage_opamp_dummy_magic_26_0.X.n32 GNDA 0.080247f
C2458 two_stage_opamp_dummy_magic_26_0.X.t39 GNDA 0.053916f
C2459 two_stage_opamp_dummy_magic_26_0.X.t54 GNDA 0.061293f
C2460 two_stage_opamp_dummy_magic_26_0.X.n34 GNDA 0.049987f
C2461 two_stage_opamp_dummy_magic_26_0.X.t53 GNDA 0.053916f
C2462 two_stage_opamp_dummy_magic_26_0.X.t38 GNDA 0.053916f
C2463 two_stage_opamp_dummy_magic_26_0.X.t52 GNDA 0.053916f
C2464 two_stage_opamp_dummy_magic_26_0.X.t34 GNDA 0.053916f
C2465 two_stage_opamp_dummy_magic_26_0.X.t48 GNDA 0.053916f
C2466 two_stage_opamp_dummy_magic_26_0.X.t35 GNDA 0.053916f
C2467 two_stage_opamp_dummy_magic_26_0.X.t49 GNDA 0.053916f
C2468 two_stage_opamp_dummy_magic_26_0.X.t31 GNDA 0.061293f
C2469 two_stage_opamp_dummy_magic_26_0.X.n35 GNDA 0.055315f
C2470 two_stage_opamp_dummy_magic_26_0.X.n36 GNDA 0.033854f
C2471 two_stage_opamp_dummy_magic_26_0.X.n37 GNDA 0.033854f
C2472 two_stage_opamp_dummy_magic_26_0.X.n38 GNDA 0.033854f
C2473 two_stage_opamp_dummy_magic_26_0.X.n39 GNDA 0.033854f
C2474 two_stage_opamp_dummy_magic_26_0.X.n40 GNDA 0.033854f
C2475 two_stage_opamp_dummy_magic_26_0.X.n41 GNDA 0.028525f
C2476 two_stage_opamp_dummy_magic_26_0.X.n42 GNDA 0.013852f
C2477 two_stage_opamp_dummy_magic_26_0.X.t50 GNDA 0.035108f
C2478 two_stage_opamp_dummy_magic_26_0.X.t36 GNDA 0.042631f
C2479 two_stage_opamp_dummy_magic_26_0.X.n43 GNDA 0.037302f
C2480 two_stage_opamp_dummy_magic_26_0.X.t32 GNDA 0.035108f
C2481 two_stage_opamp_dummy_magic_26_0.X.t46 GNDA 0.035108f
C2482 two_stage_opamp_dummy_magic_26_0.X.t29 GNDA 0.035108f
C2483 two_stage_opamp_dummy_magic_26_0.X.t42 GNDA 0.035108f
C2484 two_stage_opamp_dummy_magic_26_0.X.t25 GNDA 0.035108f
C2485 two_stage_opamp_dummy_magic_26_0.X.t43 GNDA 0.035108f
C2486 two_stage_opamp_dummy_magic_26_0.X.t26 GNDA 0.035108f
C2487 two_stage_opamp_dummy_magic_26_0.X.t40 GNDA 0.042631f
C2488 two_stage_opamp_dummy_magic_26_0.X.n44 GNDA 0.042631f
C2489 two_stage_opamp_dummy_magic_26_0.X.n45 GNDA 0.027585f
C2490 two_stage_opamp_dummy_magic_26_0.X.n46 GNDA 0.027585f
C2491 two_stage_opamp_dummy_magic_26_0.X.n47 GNDA 0.027585f
C2492 two_stage_opamp_dummy_magic_26_0.X.n48 GNDA 0.027585f
C2493 two_stage_opamp_dummy_magic_26_0.X.n49 GNDA 0.027585f
C2494 two_stage_opamp_dummy_magic_26_0.X.n50 GNDA 0.022256f
C2495 two_stage_opamp_dummy_magic_26_0.X.n51 GNDA 0.013852f
C2496 two_stage_opamp_dummy_magic_26_0.X.n52 GNDA 0.068964f
C2497 two_stage_opamp_dummy_magic_26_0.X.n53 GNDA 0.079493f
C2498 two_stage_opamp_dummy_magic_26_0.X.n54 GNDA 0.080247f
C2499 two_stage_opamp_dummy_magic_26_0.X.n55 GNDA 0.080247f
C2500 two_stage_opamp_dummy_magic_26_0.X.n56 GNDA 0.080247f
C2501 two_stage_opamp_dummy_magic_26_0.X.n57 GNDA 0.080247f
C2502 two_stage_opamp_dummy_magic_26_0.X.n59 GNDA 0.403512f
C2503 two_stage_opamp_dummy_magic_26_0.X.n60 GNDA 1.80807f
C2504 two_stage_opamp_dummy_magic_26_0.X.n62 GNDA 0.080247f
C2505 two_stage_opamp_dummy_magic_26_0.X.t2 GNDA 0.693898f
C2506 two_stage_opamp_dummy_magic_26_0.X.n63 GNDA 0.080247f
C2507 two_stage_opamp_dummy_magic_26_0.X.n64 GNDA 0.080247f
C2508 two_stage_opamp_dummy_magic_26_0.X.n65 GNDA 0.079493f
C2509 two_stage_opamp_dummy_magic_26_0.X.n66 GNDA 0.744527f
C2510 two_stage_opamp_dummy_magic_26_0.X.n68 GNDA 0.697145f
C2511 two_stage_opamp_dummy_magic_26_0.X.n69 GNDA 0.026571f
C2512 two_stage_opamp_dummy_magic_26_0.X.n70 GNDA 0.026749f
C2513 two_stage_opamp_dummy_magic_26_0.X.n71 GNDA 0.026749f
C2514 two_stage_opamp_dummy_magic_26_0.X.t30 GNDA 0.110339f
C2515 two_stage_opamp_dummy_magic_26_0.X.t47 GNDA 0.110339f
C2516 two_stage_opamp_dummy_magic_26_0.X.t33 GNDA 0.110339f
C2517 two_stage_opamp_dummy_magic_26_0.X.t51 GNDA 0.110339f
C2518 two_stage_opamp_dummy_magic_26_0.X.t37 GNDA 0.117519f
C2519 two_stage_opamp_dummy_magic_26_0.X.n72 GNDA 0.093129f
C2520 two_stage_opamp_dummy_magic_26_0.X.n73 GNDA 0.052662f
C2521 two_stage_opamp_dummy_magic_26_0.X.n74 GNDA 0.052662f
C2522 two_stage_opamp_dummy_magic_26_0.X.n75 GNDA 0.047333f
C2523 two_stage_opamp_dummy_magic_26_0.X.t44 GNDA 0.110339f
C2524 two_stage_opamp_dummy_magic_26_0.X.t27 GNDA 0.110339f
C2525 two_stage_opamp_dummy_magic_26_0.X.t45 GNDA 0.110339f
C2526 two_stage_opamp_dummy_magic_26_0.X.t28 GNDA 0.110339f
C2527 two_stage_opamp_dummy_magic_26_0.X.t41 GNDA 0.117519f
C2528 two_stage_opamp_dummy_magic_26_0.X.n76 GNDA 0.093129f
C2529 two_stage_opamp_dummy_magic_26_0.X.n77 GNDA 0.052662f
C2530 two_stage_opamp_dummy_magic_26_0.X.n78 GNDA 0.052662f
C2531 two_stage_opamp_dummy_magic_26_0.X.n79 GNDA 0.047333f
C2532 two_stage_opamp_dummy_magic_26_0.X.n80 GNDA 0.011366f
C2533 two_stage_opamp_dummy_magic_26_0.X.n81 GNDA 0.026927f
C2534 two_stage_opamp_dummy_magic_26_0.X.n82 GNDA 0.063383f
C2535 two_stage_opamp_dummy_magic_26_0.X.n83 GNDA 0.036151f
C2536 two_stage_opamp_dummy_magic_26_0.X.n84 GNDA 0.041026f
C2537 two_stage_opamp_dummy_magic_26_0.X.n85 GNDA 1.10841f
C2538 two_stage_opamp_dummy_magic_26_0.X.n86 GNDA 0.491512f
C2539 two_stage_opamp_dummy_magic_26_0.X.n87 GNDA 0.859415f
C2540 two_stage_opamp_dummy_magic_26_0.X.n88 GNDA 0.080247f
C2541 two_stage_opamp_dummy_magic_26_0.X.n90 GNDA 0.662037f
C2542 two_stage_opamp_dummy_magic_26_0.X.n91 GNDA 0.662037f
C2543 two_stage_opamp_dummy_magic_26_0.X.n93 GNDA 0.079493f
C2544 two_stage_opamp_dummy_magic_26_0.X.n94 GNDA 0.671035f
C2545 two_stage_opamp_dummy_magic_26_0.X.n96 GNDA 0.64699f
C2546 two_stage_opamp_dummy_magic_26_0.X.n97 GNDA 0.662037f
C2547 two_stage_opamp_dummy_magic_26_0.X.n98 GNDA 0.110339f
C2548 two_stage_opamp_dummy_magic_26_0.X.n99 GNDA 0.110339f
C2549 two_stage_opamp_dummy_magic_26_0.X.n100 GNDA 0.110339f
C2550 two_stage_opamp_dummy_magic_26_0.X.n101 GNDA 0.364545f
C2551 two_stage_opamp_dummy_magic_26_0.X.n102 GNDA 0.185719f
C2552 two_stage_opamp_dummy_magic_26_0.X.n103 GNDA 0.106905f
C2553 two_stage_opamp_dummy_magic_26_0.X.n104 GNDA 0.106905f
C2554 two_stage_opamp_dummy_magic_26_0.X.n105 GNDA 0.400848f
C2555 two_stage_opamp_dummy_magic_26_0.X.n106 GNDA 0.106905f
C2556 two_stage_opamp_dummy_magic_26_0.X.t3 GNDA 0.025077f
C2557 two_stage_opamp_dummy_magic_26_0.X.t9 GNDA 0.025077f
C2558 two_stage_opamp_dummy_magic_26_0.X.n107 GNDA 0.073693f
C2559 two_stage_opamp_dummy_magic_26_0.X.t12 GNDA 0.025077f
C2560 two_stage_opamp_dummy_magic_26_0.X.t14 GNDA 0.025077f
C2561 two_stage_opamp_dummy_magic_26_0.X.n108 GNDA 0.072264f
C2562 two_stage_opamp_dummy_magic_26_0.X.n109 GNDA 0.477627f
C2563 two_stage_opamp_dummy_magic_26_0.X.t18 GNDA 0.025077f
C2564 two_stage_opamp_dummy_magic_26_0.X.t13 GNDA 0.025077f
C2565 two_stage_opamp_dummy_magic_26_0.X.n110 GNDA 0.072264f
C2566 two_stage_opamp_dummy_magic_26_0.X.n111 GNDA 0.251231f
C2567 two_stage_opamp_dummy_magic_26_0.X.t11 GNDA 0.025077f
C2568 two_stage_opamp_dummy_magic_26_0.X.t17 GNDA 0.025077f
C2569 two_stage_opamp_dummy_magic_26_0.X.n112 GNDA 0.072264f
C2570 two_stage_opamp_dummy_magic_26_0.X.n113 GNDA 0.251231f
C2571 two_stage_opamp_dummy_magic_26_0.X.t10 GNDA 0.025077f
C2572 two_stage_opamp_dummy_magic_26_0.X.t15 GNDA 0.025077f
C2573 two_stage_opamp_dummy_magic_26_0.X.n114 GNDA 0.072264f
C2574 two_stage_opamp_dummy_magic_26_0.X.n115 GNDA 0.251231f
C2575 two_stage_opamp_dummy_magic_26_0.X.t16 GNDA 0.025077f
C2576 two_stage_opamp_dummy_magic_26_0.X.t4 GNDA 0.025077f
C2577 two_stage_opamp_dummy_magic_26_0.X.n116 GNDA 0.072264f
C2578 two_stage_opamp_dummy_magic_26_0.X.n117 GNDA 0.446833f
C2579 two_stage_opamp_dummy_magic_26_0.X.n118 GNDA 0.306485f
C2580 two_stage_opamp_dummy_magic_26_0.X.n119 GNDA 0.467678f
C2581 two_stage_opamp_dummy_magic_26_0.X.n120 GNDA 0.378191f
C2582 two_stage_opamp_dummy_magic_26_0.X.n121 GNDA 0.110339f
C2583 two_stage_opamp_dummy_magic_26_0.X.n122 GNDA 0.364545f
C2584 two_stage_opamp_dummy_magic_26_0.X.n123 GNDA 0.110339f
C2585 two_stage_opamp_dummy_magic_26_0.X.n124 GNDA 0.090278f
C2586 two_stage_opamp_dummy_magic_26_0.Vb1.n0 GNDA 5.32092f
C2587 two_stage_opamp_dummy_magic_26_0.Vb1.n1 GNDA 2.85762f
C2588 two_stage_opamp_dummy_magic_26_0.Vb1.n2 GNDA 1.17864f
C2589 two_stage_opamp_dummy_magic_26_0.Vb1.n3 GNDA 0.827858f
C2590 two_stage_opamp_dummy_magic_26_0.Vb1.n4 GNDA 3.26269f
C2591 two_stage_opamp_dummy_magic_26_0.Vb1.n5 GNDA 0.339027f
C2592 two_stage_opamp_dummy_magic_26_0.Vb1.t3 GNDA 0.058064f
C2593 two_stage_opamp_dummy_magic_26_0.Vb1.t2 GNDA 0.058064f
C2594 two_stage_opamp_dummy_magic_26_0.Vb1.n6 GNDA 0.132099f
C2595 two_stage_opamp_dummy_magic_26_0.Vb1.t12 GNDA 0.068766f
C2596 two_stage_opamp_dummy_magic_26_0.Vb1.t6 GNDA 0.044637f
C2597 two_stage_opamp_dummy_magic_26_0.Vb1.t10 GNDA 0.057895f
C2598 two_stage_opamp_dummy_magic_26_0.Vb1.n7 GNDA 0.059524f
C2599 two_stage_opamp_dummy_magic_26_0.Vb1.t4 GNDA 0.044637f
C2600 two_stage_opamp_dummy_magic_26_0.Vb1.t8 GNDA 0.057895f
C2601 two_stage_opamp_dummy_magic_26_0.Vb1.n8 GNDA 0.059524f
C2602 two_stage_opamp_dummy_magic_26_0.Vb1.n9 GNDA 0.044369f
C2603 two_stage_opamp_dummy_magic_26_0.Vb1.t7 GNDA 0.043548f
C2604 two_stage_opamp_dummy_magic_26_0.Vb1.t5 GNDA 0.043548f
C2605 two_stage_opamp_dummy_magic_26_0.Vb1.n10 GNDA 0.094755f
C2606 two_stage_opamp_dummy_magic_26_0.Vb1.t23 GNDA 1.3556f
C2607 two_stage_opamp_dummy_magic_26_0.Vb1.n11 GNDA 0.15936f
C2608 two_stage_opamp_dummy_magic_26_0.Vb1.t22 GNDA 0.068766f
C2609 two_stage_opamp_dummy_magic_26_0.Vb1.t32 GNDA 0.068766f
C2610 two_stage_opamp_dummy_magic_26_0.Vb1.t20 GNDA 0.068766f
C2611 two_stage_opamp_dummy_magic_26_0.Vb1.t29 GNDA 0.068766f
C2612 two_stage_opamp_dummy_magic_26_0.Vb1.t21 GNDA 0.068766f
C2613 two_stage_opamp_dummy_magic_26_0.Vb1.t30 GNDA 0.068766f
C2614 two_stage_opamp_dummy_magic_26_0.Vb1.t19 GNDA 0.068766f
C2615 two_stage_opamp_dummy_magic_26_0.Vb1.t27 GNDA 0.068766f
C2616 two_stage_opamp_dummy_magic_26_0.Vb1.t13 GNDA 0.068766f
C2617 two_stage_opamp_dummy_magic_26_0.Vb1.t1 GNDA 0.043548f
C2618 two_stage_opamp_dummy_magic_26_0.Vb1.t11 GNDA 0.043548f
C2619 two_stage_opamp_dummy_magic_26_0.Vb1.n12 GNDA 0.094755f
C2620 two_stage_opamp_dummy_magic_26_0.Vb1.n13 GNDA 0.356178f
C2621 two_stage_opamp_dummy_magic_26_0.Vb1.n14 GNDA 0.349554f
C2622 two_stage_opamp_dummy_magic_26_0.Vb1.t9 GNDA 0.043548f
C2623 two_stage_opamp_dummy_magic_26_0.Vb1.t0 GNDA 0.043548f
C2624 two_stage_opamp_dummy_magic_26_0.Vb1.n15 GNDA 0.094755f
C2625 two_stage_opamp_dummy_magic_26_0.Vb1.n16 GNDA 0.356178f
C2626 two_stage_opamp_dummy_magic_26_0.Vb1.t28 GNDA 0.068766f
C2627 two_stage_opamp_dummy_magic_26_0.Vb1.t18 GNDA 0.068766f
C2628 two_stage_opamp_dummy_magic_26_0.Vb1.t26 GNDA 0.068766f
C2629 two_stage_opamp_dummy_magic_26_0.Vb1.t17 GNDA 0.068766f
C2630 two_stage_opamp_dummy_magic_26_0.Vb1.t25 GNDA 0.068766f
C2631 two_stage_opamp_dummy_magic_26_0.Vb1.t15 GNDA 0.068766f
C2632 two_stage_opamp_dummy_magic_26_0.Vb1.t31 GNDA 0.068766f
C2633 two_stage_opamp_dummy_magic_26_0.Vb1.t16 GNDA 0.068766f
C2634 two_stage_opamp_dummy_magic_26_0.Vb1.t24 GNDA 0.068766f
C2635 two_stage_opamp_dummy_magic_26_0.Vb1.t14 GNDA 0.068766f
C2636 VDDA.n16 GNDA 0.135311f
C2637 VDDA.n17 GNDA 0.165381f
C2638 VDDA.n18 GNDA 0.135311f
C2639 VDDA.n19 GNDA 1.05242f
C2640 VDDA.n93 GNDA 0.021987f
C2641 VDDA.n192 GNDA 0.017478f
C2642 VDDA.n197 GNDA 1.91691f
C2643 VDDA.n271 GNDA 0.021987f
C2644 VDDA.n409 GNDA 0.021987f
C2645 VDDA.n529 GNDA 0.10092f
C2646 VDDA.n535 GNDA 0.014555f
C2647 VDDA.n536 GNDA 0.049717f
C2648 VDDA.t308 GNDA 0.019841f
C2649 VDDA.n542 GNDA 0.027643f
C2650 VDDA.t332 GNDA 0.016691f
C2651 VDDA.n548 GNDA 0.024063f
C2652 VDDA.t269 GNDA 0.011699f
C2653 VDDA.n550 GNDA 0.024063f
C2654 VDDA.n552 GNDA 0.024063f
C2655 VDDA.n554 GNDA 0.024063f
C2656 VDDA.n556 GNDA 0.026838f
C2657 VDDA.n557 GNDA 0.012444f
C2658 VDDA.n558 GNDA 0.037419f
C2659 VDDA.t268 GNDA 0.028034f
C2660 VDDA.t91 GNDA 0.021988f
C2661 VDDA.t155 GNDA 0.021988f
C2662 VDDA.t153 GNDA 0.021988f
C2663 VDDA.t179 GNDA 0.021988f
C2664 VDDA.t410 GNDA 0.021988f
C2665 VDDA.t66 GNDA 0.021988f
C2666 VDDA.t141 GNDA 0.021988f
C2667 VDDA.t85 GNDA 0.021988f
C2668 VDDA.t177 GNDA 0.021988f
C2669 VDDA.t160 GNDA 0.021988f
C2670 VDDA.t347 GNDA 0.028034f
C2671 VDDA.t348 GNDA 0.011699f
C2672 VDDA.n559 GNDA 0.037419f
C2673 VDDA.n560 GNDA 0.012212f
C2674 VDDA.n561 GNDA 0.013112f
C2675 VDDA.n575 GNDA 0.061458f
C2676 VDDA.n577 GNDA 0.032764f
C2677 VDDA.n579 GNDA 0.032764f
C2678 VDDA.n581 GNDA 0.032764f
C2679 VDDA.n583 GNDA 0.04404f
C2680 VDDA.n584 GNDA 0.019733f
C2681 VDDA.n588 GNDA 0.060044f
C2682 VDDA.n589 GNDA 0.024417f
C2683 VDDA.n590 GNDA 0.020598f
C2684 VDDA.t271 GNDA 0.016704f
C2685 VDDA.t391 GNDA 0.012404f
C2686 VDDA.t56 GNDA 0.012404f
C2687 VDDA.t19 GNDA 0.012404f
C2688 VDDA.t387 GNDA 0.012404f
C2689 VDDA.t84 GNDA 0.012404f
C2690 VDDA.t22 GNDA 0.012404f
C2691 VDDA.t54 GNDA 0.012404f
C2692 VDDA.t207 GNDA 0.012404f
C2693 VDDA.t4 GNDA 0.012404f
C2694 VDDA.t98 GNDA 0.012404f
C2695 VDDA.t295 GNDA 0.016704f
C2696 VDDA.n591 GNDA 0.020598f
C2697 VDDA.n592 GNDA 0.014764f
C2698 VDDA.n593 GNDA 0.085694f
C2699 VDDA.n594 GNDA 0.016632f
C2700 VDDA.n596 GNDA 0.060044f
C2701 VDDA.n599 GNDA 0.064273f
C2702 VDDA.n600 GNDA 0.014555f
C2703 VDDA.n601 GNDA 0.049717f
C2704 VDDA.t263 GNDA 0.019841f
C2705 VDDA.n606 GNDA 0.037211f
C2706 VDDA.n612 GNDA 1.05242f
C2707 VDDA.n686 GNDA 0.021987f
C2708 VDDA.n784 GNDA 0.017478f
C2709 VDDA.n840 GNDA 0.021987f
C2710 VDDA.n957 GNDA 0.09951f
C2711 VDDA.n958 GNDA 0.10092f
C2712 VDDA.n961 GNDA 0.706627f
C2713 VDDA.n1027 GNDA 0.021987f
C2714 VDDA.n1121 GNDA 1.05242f
C2715 VDDA.n1124 GNDA 0.10092f
C2716 VDDA.n1125 GNDA 0.09951f
C2717 VDDA.n1127 GNDA 0.017478f
C2718 VDDA.n1129 GNDA 0.017478f
C2719 VDDA.n1175 GNDA 0.021987f
C2720 VDDA.n1295 GNDA 0.10092f
C2721 VDDA.n1296 GNDA 0.09951f
C2722 VDDA.n1298 GNDA 0.017478f
C2723 VDDA.n1300 GNDA 0.017478f
C2724 VDDA.n1302 GNDA 0.017478f
C2725 VDDA.n1305 GNDA 0.09951f
C2726 VDDA.n1306 GNDA 0.10092f
C2727 VDDA.n1309 GNDA 1.57863f
C2728 VDDA.n1375 GNDA 0.021987f
C2729 VDDA.n1516 GNDA 0.255588f
C2730 VDDA.n1541 GNDA 0.022825f
C2731 VDDA.n1552 GNDA 0.025706f
C2732 VDDA.t414 GNDA 0.052527f
C2733 VDDA.t117 GNDA 0.052717f
C2734 VDDA.t171 GNDA 0.049898f
C2735 VDDA.t76 GNDA 0.052527f
C2736 VDDA.t30 GNDA 0.052717f
C2737 VDDA.t380 GNDA 0.049898f
C2738 VDDA.t55 GNDA 0.052527f
C2739 VDDA.t49 GNDA 0.052717f
C2740 VDDA.t103 GNDA 0.049898f
C2741 VDDA.t379 GNDA 0.052527f
C2742 VDDA.t170 GNDA 0.052717f
C2743 VDDA.t57 GNDA 0.049898f
C2744 VDDA.t42 GNDA 0.052527f
C2745 VDDA.t27 GNDA 0.052717f
C2746 VDDA.t75 GNDA 0.049898f
C2747 VDDA.n1606 GNDA 0.035209f
C2748 VDDA.t53 GNDA 0.028039f
C2749 VDDA.n1607 GNDA 0.038203f
C2750 VDDA.t50 GNDA 0.028039f
C2751 VDDA.n1608 GNDA 0.038203f
C2752 VDDA.t188 GNDA 0.028039f
C2753 VDDA.n1609 GNDA 0.038203f
C2754 VDDA.t169 GNDA 0.028039f
C2755 VDDA.n1610 GNDA 0.038203f
C2756 VDDA.t46 GNDA 0.150237f
C2757 VDDA.n1611 GNDA 0.63619f
C2758 VDDA.n1725 GNDA 0.021987f
C2759 VDDA.n1728 GNDA 2.26271f
C2760 VDDA.n1729 GNDA 1.48843f
C2761 VDDA.n1801 GNDA 0.02053f
C2762 VDDA.n1914 GNDA 0.029271f
C2763 VDDA.n1915 GNDA 0.01429f
C2764 VDDA.n1925 GNDA 0.016632f
C2765 VDDA.t363 GNDA 0.013813f
C2766 VDDA.t224 GNDA 0.012404f
C2767 VDDA.t329 GNDA 0.013813f
C2768 VDDA.n1933 GNDA 0.016632f
C2769 VDDA.n1938 GNDA 0.015099f
C2770 VDDA.n1939 GNDA 0.016634f
C2771 VDDA.n2056 GNDA 5.20949f
C2772 VDDA.t421 GNDA 0.111005f
C2773 VDDA.t423 GNDA 0.111005f
C2774 VDDA.t424 GNDA 0.10546f
C2775 VDDA.n2089 GNDA 0.204113f
C2776 VDDA.n2090 GNDA 0.107772f
C2777 VDDA.t422 GNDA 0.104174f
C2778 VDDA.n2091 GNDA 0.139848f
C2779 VDDA.n2092 GNDA 0.073953f
C2780 VDDA.n2097 GNDA 0.053279f
C2781 VDDA.n2098 GNDA 0.053279f
C2782 VDDA.n2100 GNDA 0.02512f
C2783 VDDA.n2104 GNDA 0.02512f
C2784 VDDA.n2106 GNDA 0.02512f
C2785 VDDA.n2108 GNDA 0.02512f
C2786 VDDA.n2110 GNDA 0.02512f
C2787 VDDA.n2112 GNDA 0.02512f
C2788 VDDA.n2114 GNDA 0.02512f
C2789 VDDA.n2116 GNDA 0.02512f
C2790 VDDA.n2118 GNDA 0.02512f
C2791 VDDA.n2120 GNDA 0.02512f
C2792 VDDA.n2124 GNDA 0.02512f
C2793 VDDA.n2126 GNDA 0.02512f
C2794 VDDA.n2128 GNDA 0.02512f
C2795 VDDA.n2130 GNDA 0.02512f
C2796 VDDA.n2132 GNDA 0.02512f
C2797 VDDA.n2134 GNDA 0.02512f
C2798 VDDA.n2136 GNDA 0.02512f
C2799 VDDA.n2138 GNDA 0.03423f
C2800 VDDA.n2139 GNDA 0.010985f
C2801 VDDA.n2142 GNDA 0.011583f
C2802 VDDA.t301 GNDA 0.011994f
C2803 VDDA.n2147 GNDA 0.025536f
C2804 VDDA.n2148 GNDA 0.025536f
C2805 VDDA.n2149 GNDA 0.010345f
C2806 VDDA.n2152 GNDA 0.012161f
C2807 VDDA.t353 GNDA 0.011811f
C2808 VDDA.n2157 GNDA 0.05429f
C2809 VDDA.n2158 GNDA 0.04905f
C2810 VDDA.n2163 GNDA 0.03862f
C2811 VDDA.n2164 GNDA 0.03862f
C2812 VDDA.t282 GNDA 0.013442f
C2813 VDDA.n2166 GNDA 0.010968f
C2814 VDDA.n2167 GNDA 0.010968f
C2815 VDDA.n2168 GNDA 0.010968f
C2816 VDDA.n2169 GNDA 0.010968f
C2817 VDDA.n2170 GNDA 0.010968f
C2818 VDDA.n2171 GNDA 0.010968f
C2819 VDDA.n2172 GNDA 0.010968f
C2820 VDDA.n2173 GNDA 0.010968f
C2821 VDDA.n2199 GNDA 0.026357f
C2822 VDDA.t283 GNDA 0.027955f
C2823 VDDA.t64 GNDA 0.028754f
C2824 VDDA.t77 GNDA 0.028754f
C2825 VDDA.t193 GNDA 0.028754f
C2826 VDDA.t99 GNDA 0.028754f
C2827 VDDA.t79 GNDA 0.028754f
C2828 VDDA.t182 GNDA 0.028754f
C2829 VDDA.t118 GNDA 0.028754f
C2830 VDDA.t51 GNDA 0.028754f
C2831 VDDA.t104 GNDA 0.028754f
C2832 VDDA.t62 GNDA 0.028754f
C2833 VDDA.t149 GNDA 0.028754f
C2834 VDDA.t7 GNDA 0.028754f
C2835 VDDA.t101 GNDA 0.028754f
C2836 VDDA.t167 GNDA 0.028754f
C2837 VDDA.t28 GNDA 0.028754f
C2838 VDDA.t60 GNDA 0.028754f
C2839 VDDA.t370 GNDA 0.027955f
C2840 VDDA.n2216 GNDA 0.026357f
C2841 VDDA.t369 GNDA 0.013442f
C2842 VDDA.n2220 GNDA 0.053721f
C2843 VDDA.n2221 GNDA 0.037706f
C2844 VDDA.n2222 GNDA 0.037706f
C2845 VDDA.n2223 GNDA 0.037706f
C2846 VDDA.n2224 GNDA 0.037706f
C2847 VDDA.n2225 GNDA 0.037706f
C2848 VDDA.n2226 GNDA 0.037706f
C2849 VDDA.n2227 GNDA 0.037706f
C2850 VDDA.n2228 GNDA 0.031795f
C2851 VDDA.n2229 GNDA 0.036255f
C2852 VDDA.n2231 GNDA 0.017245f
C2853 VDDA.t367 GNDA 0.011653f
C2854 VDDA.t286 GNDA 0.011402f
C2855 VDDA.n2232 GNDA 0.016466f
C2856 VDDA.n2234 GNDA 0.066136f
C2857 VDDA.n2235 GNDA 0.049896f
C2858 VDDA.n2240 GNDA 0.018042f
C2859 VDDA.n2241 GNDA 0.018042f
C2860 VDDA.n2244 GNDA 0.016375f
C2861 VDDA.t350 GNDA 0.011401f
C2862 VDDA.t259 GNDA 0.011401f
C2863 VDDA.n2245 GNDA 0.016375f
C2864 VDDA.t292 GNDA 0.010308f
C2865 VDDA.t360 GNDA 0.010308f
C2866 VDDA.n2259 GNDA 0.016375f
C2867 VDDA.t338 GNDA 0.011401f
C2868 VDDA.t356 GNDA 0.011401f
C2869 VDDA.n2260 GNDA 0.016375f
C2870 VDDA.t313 GNDA 0.010308f
C2871 VDDA.t344 GNDA 0.010308f
C2872 VDDA.n2268 GNDA 0.033115f
C2873 VDDA.n2269 GNDA 0.0209f
C2874 VDDA.n2270 GNDA 0.025876f
C2875 VDDA.n2271 GNDA 0.023338f
C2876 VDDA.n2272 GNDA 0.018367f
C2877 VDDA.n2273 GNDA 0.020904f
C2878 VDDA.n2274 GNDA 0.020904f
C2879 VDDA.n2275 GNDA 0.020904f
C2880 VDDA.n2276 GNDA 0.018367f
C2881 VDDA.n2277 GNDA 0.023338f
C2882 VDDA.n2278 GNDA 0.025876f
C2883 VDDA.n2279 GNDA 0.020899f
C2884 VDDA.n2280 GNDA 0.020899f
C2885 VDDA.n2281 GNDA 0.025876f
C2886 VDDA.n2282 GNDA 0.026439f
C2887 VDDA.n2283 GNDA 0.022032f
C2888 VDDA.n2284 GNDA 0.054347f
C2889 VDDA.n2285 GNDA 0.04595f
C2890 VDDA.n2290 GNDA 0.026499f
C2891 VDDA.n2292 GNDA 0.02819f
C2892 VDDA.n2402 GNDA 0.021987f
C2893 VDDA.n2405 GNDA 5.90111f
C2894 VDDA.n2406 GNDA 1.9094f
C2895 VDDA.n2409 GNDA 0.10092f
C2896 VDDA.n2411 GNDA 0.09951f
C2897 VDDA.n2413 GNDA 0.037211f
C2898 VDDA.n2414 GNDA 0.053843f
C2899 VDDA.n2418 GNDA 0.053843f
C2900 VDDA.n2420 GNDA 0.030445f
C2901 VDDA.n2421 GNDA 0.014555f
C2902 VDDA.n2422 GNDA 0.049717f
C2903 VDDA.n2423 GNDA 0.014555f
C2904 VDDA.n2424 GNDA 0.049717f
C2905 VDDA.n2425 GNDA 0.014555f
C2906 VDDA.n2426 GNDA 0.049717f
C2907 VDDA.n2427 GNDA 0.014555f
C2908 VDDA.n2428 GNDA 0.049717f
C2909 VDDA.n2429 GNDA 0.035404f
C2910 VDDA.n2430 GNDA 0.017898f
C2911 VDDA.n2431 GNDA 0.066371f
C2912 VDDA.t262 GNDA 0.042987f
C2913 VDDA.t383 GNDA 0.033076f
C2914 VDDA.t205 GNDA 0.032867f
C2915 VDDA.t20 GNDA 0.032628f
C2916 VDDA.t44 GNDA 0.033076f
C2917 VDDA.t96 GNDA 0.033076f
C2918 VDDA.t175 GNDA 0.033076f
C2919 VDDA.t392 GNDA 0.033076f
C2920 VDDA.t89 GNDA 0.033076f
C2921 VDDA.t385 GNDA 0.033076f
C2922 VDDA.t58 GNDA 0.033076f
C2923 VDDA.t289 GNDA 0.042987f
C2924 VDDA.t290 GNDA 0.019841f
C2925 VDDA.n2432 GNDA 0.066371f
C2926 VDDA.n2433 GNDA 0.017898f
C2927 VDDA.n2434 GNDA 0.021591f
C2928 VDDA.n2435 GNDA 0.016632f
C2929 VDDA.n2436 GNDA 0.064273f
C2930 VDDA.n2439 GNDA 0.029036f
C2931 VDDA.n2440 GNDA 0.029036f
C2932 VDDA.n2443 GNDA 0.037442f
C2933 VDDA.n2445 GNDA 0.052715f
C2934 VDDA.t166 GNDA 0.014988f
C2935 VDDA.t0 GNDA 0.014988f
C2936 VDDA.t70 GNDA 0.014988f
C2937 VDDA.t181 GNDA 0.014988f
C2938 VDDA.t304 GNDA 0.020049f
C2939 VDDA.n2446 GNDA 0.023741f
C2940 VDDA.n2448 GNDA 0.06365f
C2941 VDDA.n2450 GNDA 0.027643f
C2942 VDDA.n2451 GNDA 0.013813f
C2943 VDDA.n2456 GNDA 0.039091f
C2944 VDDA.t311 GNDA 0.014988f
C2945 VDDA.n2458 GNDA 0.015247f
C2946 VDDA.n2459 GNDA 0.037419f
C2947 VDDA.t310 GNDA 0.028034f
C2948 VDDA.t412 GNDA 0.021988f
C2949 VDDA.t341 GNDA 0.028034f
C2950 VDDA.t342 GNDA 0.011699f
C2951 VDDA.n2460 GNDA 0.037419f
C2952 VDDA.n2461 GNDA 0.015024f
C2953 VDDA.n2462 GNDA 0.018519f
C2954 VDDA.n2466 GNDA 0.013813f
C2955 VDDA.n2470 GNDA 0.030163f
C2956 VDDA.n2471 GNDA 0.012304f
C2957 VDDA.n2472 GNDA 0.018381f
C2958 VDDA.t319 GNDA 0.016364f
C2959 VDDA.t16 GNDA 0.012404f
C2960 VDDA.t298 GNDA 0.016364f
C2961 VDDA.n2473 GNDA 0.018381f
C2962 VDDA.n2474 GNDA 0.01208f
C2963 VDDA.n2475 GNDA 0.018519f
C2964 VDDA.n2476 GNDA 0.013813f
C2965 VDDA.n2482 GNDA 0.024807f
C2966 VDDA.n2483 GNDA 0.024807f
C2967 VDDA.n2485 GNDA 0.013813f
C2968 VDDA.n2489 GNDA 0.015868f
C2969 VDDA.n2490 GNDA 0.013696f
C2970 VDDA.t265 GNDA 0.016691f
C2971 VDDA.t33 GNDA 0.014988f
C2972 VDDA.t2 GNDA 0.014988f
C2973 VDDA.t5 GNDA 0.014988f
C2974 VDDA.t120 GNDA 0.014988f
C2975 VDDA.t277 GNDA 0.020049f
C2976 VDDA.n2491 GNDA 0.023741f
C2977 VDDA.n2493 GNDA 0.06365f
C2978 VDDA.n2497 GNDA 0.024063f
C2979 VDDA.n2499 GNDA 0.024063f
C2980 VDDA.n2501 GNDA 0.024063f
C2981 VDDA.n2503 GNDA 0.024063f
C2982 VDDA.n2505 GNDA 0.026838f
C2983 VDDA.n2506 GNDA 0.012444f
C2984 VDDA.t336 GNDA 0.011699f
C2985 VDDA.n2507 GNDA 0.037419f
C2986 VDDA.t335 GNDA 0.028034f
C2987 VDDA.t31 GNDA 0.021988f
C2988 VDDA.t418 GNDA 0.021988f
C2989 VDDA.t394 GNDA 0.021988f
C2990 VDDA.t191 GNDA 0.021988f
C2991 VDDA.t81 GNDA 0.021988f
C2992 VDDA.t25 GNDA 0.021988f
C2993 VDDA.t199 GNDA 0.021988f
C2994 VDDA.t40 GNDA 0.021988f
C2995 VDDA.t139 GNDA 0.021988f
C2996 VDDA.t113 GNDA 0.021988f
C2997 VDDA.t373 GNDA 0.028034f
C2998 VDDA.t374 GNDA 0.011699f
C2999 VDDA.n2508 GNDA 0.037419f
C3000 VDDA.n2509 GNDA 0.012212f
C3001 VDDA.n2510 GNDA 0.013111f
C3002 VDDA.n2512 GNDA 0.037443f
C3003 VDDA.n2514 GNDA 0.052715f
C3004 VDDA.n2515 GNDA 0.029036f
C3005 VDDA.n2527 GNDA 0.061458f
C3006 VDDA.n2529 GNDA 0.032764f
C3007 VDDA.n2531 GNDA 0.032764f
C3008 VDDA.n2533 GNDA 0.032764f
C3009 VDDA.n2535 GNDA 0.04404f
C3010 VDDA.n2536 GNDA 0.019733f
C3011 VDDA.n2538 GNDA 0.060044f
C3012 VDDA.n2540 GNDA 0.060044f
C3013 VDDA.n2542 GNDA 0.024417f
C3014 VDDA.n2543 GNDA 0.020598f
C3015 VDDA.t326 GNDA 0.016704f
C3016 VDDA.t116 GNDA 0.012404f
C3017 VDDA.t129 GNDA 0.012404f
C3018 VDDA.t34 GNDA 0.012404f
C3019 VDDA.t400 GNDA 0.012404f
C3020 VDDA.t37 GNDA 0.012404f
C3021 VDDA.t389 GNDA 0.012404f
C3022 VDDA.t132 GNDA 0.012404f
C3023 VDDA.t406 GNDA 0.012404f
C3024 VDDA.t390 GNDA 0.012404f
C3025 VDDA.t401 GNDA 0.012404f
C3026 VDDA.t316 GNDA 0.016704f
C3027 VDDA.n2544 GNDA 0.020598f
C3028 VDDA.n2545 GNDA 0.014764f
C3029 VDDA.n2546 GNDA 0.085694f
C3030 VDDA.n2547 GNDA 0.016632f
C3031 VDDA.n2549 GNDA 0.064273f
C3032 VDDA.n2550 GNDA 0.064273f
C3033 VDDA.n2553 GNDA 0.029036f
C3034 VDDA.n2555 GNDA 0.016632f
C3035 VDDA.n2556 GNDA 0.014555f
C3036 VDDA.n2557 GNDA 0.049717f
C3037 VDDA.n2558 GNDA 0.014555f
C3038 VDDA.n2559 GNDA 0.049717f
C3039 VDDA.n2560 GNDA 0.014555f
C3040 VDDA.n2561 GNDA 0.049717f
C3041 VDDA.n2562 GNDA 0.014555f
C3042 VDDA.n2563 GNDA 0.049717f
C3043 VDDA.n2564 GNDA 0.021591f
C3044 VDDA.n2565 GNDA 0.017898f
C3045 VDDA.n2566 GNDA 0.066371f
C3046 VDDA.t307 GNDA 0.042987f
C3047 VDDA.t130 GNDA 0.033076f
C3048 VDDA.t73 GNDA 0.033076f
C3049 VDDA.t111 GNDA 0.033076f
C3050 VDDA.t173 GNDA 0.033076f
C3051 VDDA.t35 GNDA 0.033076f
C3052 VDDA.t145 GNDA 0.033076f
C3053 VDDA.t415 GNDA 0.033076f
C3054 VDDA.t407 GNDA 0.033076f
C3055 VDDA.t398 GNDA 0.033076f
C3056 VDDA.t38 GNDA 0.033076f
C3057 VDDA.t323 GNDA 0.042987f
C3058 VDDA.t324 GNDA 0.019841f
C3059 VDDA.n2567 GNDA 0.066371f
C3060 VDDA.n2568 GNDA 0.017898f
C3061 VDDA.n2569 GNDA 0.035404f
C3062 VDDA.n2570 GNDA 0.030445f
C3063 VDDA.n2574 GNDA 0.053843f
C3064 VDDA.n2575 GNDA 0.053843f
C3065 VDDA.n2578 GNDA 0.09951f
C3066 VDDA.n2580 GNDA 0.037211f
C3067 VDDA.n2582 GNDA 0.037211f
C3068 VDDA.n2585 GNDA 0.09951f
C3069 VDDA.n2586 GNDA 0.10092f
C3070 VDDA.n2589 GNDA 1.57863f
C3071 VDDA.n2655 GNDA 0.021987f
C3072 VDDA.n2749 GNDA 1.05242f
C3073 VDDA.n2752 GNDA 0.10092f
C3074 VDDA.n2753 GNDA 0.09951f
C3075 VDDA.n2755 GNDA 0.017478f
C3076 VDDA.n2757 GNDA 0.017478f
C3077 VDDA.n2803 GNDA 0.021987f
C3078 VDDA.n2923 GNDA 0.10092f
C3079 VDDA.n2924 GNDA 0.09951f
C3080 VDDA.n2926 GNDA 0.017478f
C3081 VDDA.n2928 GNDA 0.017478f
C3082 VDDA.n2929 GNDA 0.017478f
C3083 VDDA.n2933 GNDA 0.09951f
C3084 VDDA.n2934 GNDA 0.10092f
C3085 VDDA.n2937 GNDA 56.376f
C3086 VDDA.n2938 GNDA 0.067656f
C3087 VDDA.n2939 GNDA 0.067656f
C3088 VDDA.n2940 GNDA 0.067656f
C3089 VDDA.n2941 GNDA 0.067656f
C3090 VDDA.n2942 GNDA 0.067656f
C3091 VDDA.n2943 GNDA 0.067656f
C3092 VDDA.n2944 GNDA 0.067656f
C3093 VDDA.n2945 GNDA 0.067656f
C3094 VDDA.n2946 GNDA 0.067656f
C3095 VDDA.n2947 GNDA 0.067656f
C3096 VDDA.n2948 GNDA 0.067656f
C3097 VDDA.n2949 GNDA 0.067656f
C3098 VDDA.n2950 GNDA 0.067656f
C3099 VDDA.n2951 GNDA 0.067656f
C3100 VDDA.n2952 GNDA 0.067656f
C3101 VDDA.n2953 GNDA 0.067656f
C3102 VDDA.n2954 GNDA 0.067656f
C3103 VDDA.n2955 GNDA 0.086449f
C3104 VDDA.n2956 GNDA 0.067656f
C3105 VDDA.n2957 GNDA 0.067656f
C3106 VDDA.n2958 GNDA 0.067656f
C3107 VDDA.n2959 GNDA 0.067656f
C3108 VDDA.n2960 GNDA 0.067656f
C3109 VDDA.n2961 GNDA 0.067656f
C3110 VDDA.n2962 GNDA 0.067656f
C3111 VDDA.n2963 GNDA 0.067656f
C3112 VDDA.n2964 GNDA 0.067656f
C3113 VDDA.n2965 GNDA 0.067656f
C3114 VDDA.n2966 GNDA 0.067656f
C3115 VDDA.n2967 GNDA 0.067656f
C3116 VDDA.n2968 GNDA 0.067656f
C3117 VDDA.n2969 GNDA 0.067656f
C3118 VDDA.n2970 GNDA 0.067656f
C3119 VDDA.n2971 GNDA 0.067656f
C3120 VDDA.n2972 GNDA 0.135311f
C3121 VDDA.n2974 GNDA 0.067656f
C3122 VDDA.n2977 GNDA 0.067656f
C3123 VDDA.n2980 GNDA 0.067656f
C3124 VDDA.n2983 GNDA 0.067656f
C3125 VDDA.n2986 GNDA 0.067656f
C3126 VDDA.n2989 GNDA 0.067656f
C3127 VDDA.n2992 GNDA 0.067656f
C3128 VDDA.n2995 GNDA 0.067656f
C3129 VDDA.n2998 GNDA 0.067656f
C3130 VDDA.n3001 GNDA 0.067656f
C3131 VDDA.n3004 GNDA 0.067656f
C3132 VDDA.n3007 GNDA 0.067656f
C3133 VDDA.n3010 GNDA 0.067656f
C3134 VDDA.n3013 GNDA 0.067656f
C3135 VDDA.n3016 GNDA 0.067656f
C3136 VDDA.n3019 GNDA 0.067656f
C3137 VDDA.n3022 GNDA 0.067656f
C3138 VDDA.n3025 GNDA 0.086449f
C3139 VDDA.n3028 GNDA 0.067656f
C3140 VDDA.n3031 GNDA 0.067656f
C3141 VDDA.n3034 GNDA 0.067656f
C3142 VDDA.n3037 GNDA 0.067656f
C3143 VDDA.n3040 GNDA 0.067656f
C3144 VDDA.n3043 GNDA 0.067656f
C3145 VDDA.n3046 GNDA 0.067656f
C3146 VDDA.n3049 GNDA 0.067656f
C3147 VDDA.n3052 GNDA 0.067656f
C3148 VDDA.n3055 GNDA 0.067656f
C3149 VDDA.n3058 GNDA 0.067656f
C3150 VDDA.n3061 GNDA 0.067656f
C3151 VDDA.n3064 GNDA 0.067656f
C3152 VDDA.n3067 GNDA 0.067656f
C3153 VDDA.n3070 GNDA 0.067656f
C3154 VDDA.n3073 GNDA 0.067656f
C3155 VDDA.n3076 GNDA 0.135311f
C3156 VDDA.n3077 GNDA 0.135311f
C3157 VDDA.n3078 GNDA 0.135311f
C3158 VDDA.n3079 GNDA 0.135311f
C3159 VDDA.n3080 GNDA 0.135311f
C3160 VDDA.n3081 GNDA 0.135311f
C3161 VDDA.n3082 GNDA 0.135311f
C3162 VDDA.n3083 GNDA 0.135311f
C3163 VDDA.n3084 GNDA 0.135311f
C3164 VDDA.n3085 GNDA 0.135311f
C3165 VDDA.n3086 GNDA 0.135311f
C3166 VDDA.n3087 GNDA 0.135311f
C3167 VDDA.n3088 GNDA 0.135311f
C3168 VDDA.n3089 GNDA 0.135311f
C3169 VDDA.n3090 GNDA 0.135311f
C3170 VDDA.n3093 GNDA 0.135311f
C3171 VDDA.n3095 GNDA 0.135311f
C3172 VDDA.n3097 GNDA 0.135311f
C3173 VDDA.n3099 GNDA 0.135311f
C3174 VDDA.n3101 GNDA 0.135311f
C3175 VDDA.n3103 GNDA 0.135311f
C3176 VDDA.n3105 GNDA 0.135311f
C3177 VDDA.n3107 GNDA 0.135311f
C3178 VDDA.n3109 GNDA 0.135311f
C3179 VDDA.n3111 GNDA 0.135311f
C3180 VDDA.n3113 GNDA 0.135311f
C3181 VDDA.n3115 GNDA 0.135311f
C3182 VDDA.n3117 GNDA 0.135311f
C3183 VDDA.n3119 GNDA 0.135311f
C3184 VDDA.n3121 GNDA 0.135311f
C3185 VDDA.n3122 GNDA 0.08269f
C3186 VDDA.n3123 GNDA 55.9175f
C3187 VDDA.n3124 GNDA 0.441642f
C3188 bgr_11_0.PFET_GATE_10uA.t28 GNDA 0.023614f
C3189 bgr_11_0.PFET_GATE_10uA.t20 GNDA 0.023614f
C3190 bgr_11_0.PFET_GATE_10uA.n0 GNDA 0.082684f
C3191 bgr_11_0.PFET_GATE_10uA.t13 GNDA 0.020346f
C3192 bgr_11_0.PFET_GATE_10uA.t24 GNDA 0.030076f
C3193 bgr_11_0.PFET_GATE_10uA.n1 GNDA 0.03314f
C3194 bgr_11_0.PFET_GATE_10uA.t17 GNDA 0.020346f
C3195 bgr_11_0.PFET_GATE_10uA.t25 GNDA 0.030076f
C3196 bgr_11_0.PFET_GATE_10uA.n2 GNDA 0.03314f
C3197 bgr_11_0.PFET_GATE_10uA.n3 GNDA 0.032464f
C3198 bgr_11_0.PFET_GATE_10uA.n4 GNDA 1.03417f
C3199 bgr_11_0.PFET_GATE_10uA.t1 GNDA 0.363431f
C3200 bgr_11_0.PFET_GATE_10uA.t0 GNDA 0.324056f
C3201 bgr_11_0.PFET_GATE_10uA.t3 GNDA 0.020867f
C3202 bgr_11_0.PFET_GATE_10uA.t7 GNDA 0.020867f
C3203 bgr_11_0.PFET_GATE_10uA.n5 GNDA 0.045075f
C3204 bgr_11_0.PFET_GATE_10uA.n6 GNDA 1.1187f
C3205 bgr_11_0.PFET_GATE_10uA.t9 GNDA 0.020867f
C3206 bgr_11_0.PFET_GATE_10uA.t5 GNDA 0.020867f
C3207 bgr_11_0.PFET_GATE_10uA.n7 GNDA 0.045075f
C3208 bgr_11_0.PFET_GATE_10uA.n8 GNDA 0.455737f
C3209 bgr_11_0.PFET_GATE_10uA.t8 GNDA 0.020867f
C3210 bgr_11_0.PFET_GATE_10uA.t4 GNDA 0.020867f
C3211 bgr_11_0.PFET_GATE_10uA.n9 GNDA 0.045075f
C3212 bgr_11_0.PFET_GATE_10uA.n10 GNDA 0.446347f
C3213 bgr_11_0.PFET_GATE_10uA.t6 GNDA 0.020867f
C3214 bgr_11_0.PFET_GATE_10uA.t2 GNDA 0.020867f
C3215 bgr_11_0.PFET_GATE_10uA.n11 GNDA 0.045075f
C3216 bgr_11_0.PFET_GATE_10uA.n12 GNDA 0.700571f
C3217 bgr_11_0.PFET_GATE_10uA.n13 GNDA 2.98162f
C3218 bgr_11_0.PFET_GATE_10uA.t26 GNDA 0.074194f
C3219 bgr_11_0.PFET_GATE_10uA.n14 GNDA 1.61003f
C3220 bgr_11_0.PFET_GATE_10uA.t15 GNDA 0.020346f
C3221 bgr_11_0.PFET_GATE_10uA.t10 GNDA 0.030076f
C3222 bgr_11_0.PFET_GATE_10uA.n15 GNDA 0.03314f
C3223 bgr_11_0.PFET_GATE_10uA.t21 GNDA 0.020346f
C3224 bgr_11_0.PFET_GATE_10uA.t11 GNDA 0.030076f
C3225 bgr_11_0.PFET_GATE_10uA.n16 GNDA 0.03314f
C3226 bgr_11_0.PFET_GATE_10uA.n17 GNDA 0.031974f
C3227 bgr_11_0.PFET_GATE_10uA.n18 GNDA 1.29057f
C3228 bgr_11_0.PFET_GATE_10uA.t14 GNDA 0.020346f
C3229 bgr_11_0.PFET_GATE_10uA.t19 GNDA 0.020346f
C3230 bgr_11_0.PFET_GATE_10uA.t18 GNDA 0.020346f
C3231 bgr_11_0.PFET_GATE_10uA.t27 GNDA 0.030076f
C3232 bgr_11_0.PFET_GATE_10uA.n19 GNDA 0.037221f
C3233 bgr_11_0.PFET_GATE_10uA.n20 GNDA 0.026606f
C3234 bgr_11_0.PFET_GATE_10uA.n21 GNDA 0.020737f
C3235 bgr_11_0.PFET_GATE_10uA.t23 GNDA 0.020346f
C3236 bgr_11_0.PFET_GATE_10uA.t16 GNDA 0.020346f
C3237 bgr_11_0.PFET_GATE_10uA.t12 GNDA 0.020346f
C3238 bgr_11_0.PFET_GATE_10uA.t22 GNDA 0.030076f
C3239 bgr_11_0.PFET_GATE_10uA.n22 GNDA 0.037221f
C3240 bgr_11_0.PFET_GATE_10uA.n23 GNDA 0.026606f
C3241 bgr_11_0.PFET_GATE_10uA.n24 GNDA 0.020737f
C3242 bgr_11_0.PFET_GATE_10uA.n25 GNDA 0.059033f
C3243 bgr_11_0.1st_Vout_2.n0 GNDA 1.07305f
C3244 bgr_11_0.1st_Vout_2.n1 GNDA 0.297625f
C3245 bgr_11_0.1st_Vout_2.n2 GNDA 0.668271f
C3246 bgr_11_0.1st_Vout_2.n3 GNDA 0.091542f
C3247 bgr_11_0.1st_Vout_2.n4 GNDA 0.158156f
C3248 bgr_11_0.1st_Vout_2.t14 GNDA 0.011681f
C3249 bgr_11_0.1st_Vout_2.n6 GNDA 0.010675f
C3250 bgr_11_0.1st_Vout_2.n7 GNDA 0.115898f
C3251 bgr_11_0.1st_Vout_2.n8 GNDA 0.0146f
C3252 bgr_11_0.1st_Vout_2.t15 GNDA 0.011528f
C3253 bgr_11_0.1st_Vout_2.t29 GNDA 0.194725f
C3254 bgr_11_0.1st_Vout_2.t32 GNDA 0.198042f
C3255 bgr_11_0.1st_Vout_2.t27 GNDA 0.194725f
C3256 bgr_11_0.1st_Vout_2.t20 GNDA 0.194725f
C3257 bgr_11_0.1st_Vout_2.t12 GNDA 0.198042f
C3258 bgr_11_0.1st_Vout_2.t13 GNDA 0.198042f
C3259 bgr_11_0.1st_Vout_2.t31 GNDA 0.194725f
C3260 bgr_11_0.1st_Vout_2.t25 GNDA 0.194725f
C3261 bgr_11_0.1st_Vout_2.t19 GNDA 0.198042f
C3262 bgr_11_0.1st_Vout_2.t30 GNDA 0.198042f
C3263 bgr_11_0.1st_Vout_2.t24 GNDA 0.194725f
C3264 bgr_11_0.1st_Vout_2.t18 GNDA 0.194725f
C3265 bgr_11_0.1st_Vout_2.t11 GNDA 0.198042f
C3266 bgr_11_0.1st_Vout_2.t23 GNDA 0.198042f
C3267 bgr_11_0.1st_Vout_2.t17 GNDA 0.194725f
C3268 bgr_11_0.1st_Vout_2.t10 GNDA 0.194725f
C3269 bgr_11_0.1st_Vout_2.t28 GNDA 0.198042f
C3270 bgr_11_0.1st_Vout_2.t8 GNDA 0.198042f
C3271 bgr_11_0.1st_Vout_2.t16 GNDA 0.194725f
C3272 bgr_11_0.1st_Vout_2.t22 GNDA 0.194725f
C3273 bgr_11_0.1st_Vout_2.n9 GNDA 0.641071f
C3274 bgr_11_0.1st_Vout_2.n10 GNDA 0.010675f
C3275 bgr_11_0.1st_Vout_2.n11 GNDA 0.0146f
C3276 bgr_11_0.1st_Vout_2.n12 GNDA 0.14235f
C3277 bgr_11_0.1st_Vout_2.t0 GNDA 0.044569f
.ends

