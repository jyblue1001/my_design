magic
tech sky130A
timestamp 1752398240
<< error_s >>
rect 4150 2460 4170 2480
rect 4175 2460 4184 2480
rect 4150 2240 4170 2260
<< metal1 >>
rect 2950 6685 2990 6690
rect 2950 6655 2955 6685
rect 2985 6655 2990 6685
rect 2950 6650 2990 6655
rect 3030 6685 3070 6690
rect 3030 6655 3035 6685
rect 3065 6655 3070 6685
rect 6095 6685 6135 6690
rect 6095 6655 6100 6685
rect 6130 6655 6135 6685
rect 3030 6650 3070 6655
rect 2905 6580 2945 6585
rect 2905 6550 2910 6580
rect 2940 6550 2945 6580
rect 2905 6545 2945 6550
rect 2915 3090 2935 6545
rect 2960 3140 2980 6650
rect 3280 6525 3300 6650
rect 3400 6645 3440 6650
rect 3400 6615 3405 6645
rect 3435 6615 3440 6645
rect 3400 6610 3440 6615
rect 3270 6520 3310 6525
rect 3270 6490 3275 6520
rect 3305 6490 3310 6520
rect 3270 6485 3310 6490
rect 3555 6480 3575 6655
rect 3955 6645 3995 6650
rect 3955 6615 3960 6645
rect 3990 6615 3995 6645
rect 3955 6610 3995 6615
rect 3545 6475 3585 6480
rect 3545 6445 3550 6475
rect 3580 6445 3585 6475
rect 3545 6440 3585 6445
rect 3965 3780 3985 6610
rect 4340 6585 4360 6655
rect 4330 6580 4370 6585
rect 4330 6550 4335 6580
rect 4365 6550 4370 6580
rect 4330 6545 4370 6550
rect 4000 6475 4040 6480
rect 4000 6445 4005 6475
rect 4035 6445 4040 6475
rect 4000 6440 4040 6445
rect 4010 5405 4030 6440
rect 4000 5400 4040 5405
rect 4000 5370 4005 5400
rect 4035 5370 4040 5400
rect 4000 5365 4040 5370
rect 4090 5400 4130 5405
rect 4090 5370 4095 5400
rect 4125 5370 4130 5400
rect 4090 5365 4130 5370
rect 3965 3775 4030 3780
rect 3965 3745 3985 3775
rect 4015 3745 4030 3775
rect 3965 3740 4030 3745
rect 4010 3640 4030 3740
rect 4000 3635 4040 3640
rect 4000 3605 4005 3635
rect 4035 3605 4040 3635
rect 2950 3135 2990 3140
rect 2950 3105 2955 3135
rect 2985 3105 2990 3135
rect 3055 3135 3095 3140
rect 3055 3105 3060 3135
rect 3090 3105 3095 3135
rect 2905 3085 2945 3090
rect 2905 3055 2910 3085
rect 2940 3055 2945 3085
rect 2905 3050 2945 3055
rect 3010 3085 3050 3090
rect 3010 3055 3015 3085
rect 3045 3055 3050 3085
rect 3010 3050 3050 3055
rect 3020 2865 3040 3050
rect 3065 2755 3085 3105
rect 4100 2890 4120 5365
rect 5085 5340 5105 6655
rect 5730 6585 5750 6655
rect 6095 6650 6135 6655
rect 6700 6685 6740 6690
rect 6700 6655 6705 6685
rect 6735 6655 6740 6685
rect 7020 6685 7060 6690
rect 7020 6655 7025 6685
rect 7055 6655 7060 6685
rect 6700 6650 6740 6655
rect 5720 6580 5760 6585
rect 5720 6550 5725 6580
rect 5755 6550 5760 6580
rect 5720 6545 5760 6550
rect 5375 6520 5415 6525
rect 5375 6490 5380 6520
rect 5410 6490 5415 6520
rect 5375 6485 5415 6490
rect 5385 5420 5405 6485
rect 5375 5415 5415 5420
rect 5375 5385 5380 5415
rect 5410 5385 5415 5415
rect 5375 5380 5415 5385
rect 5495 5415 5535 5420
rect 5495 5385 5500 5415
rect 5530 5385 5535 5415
rect 5495 5380 5535 5385
rect 5075 5335 5115 5340
rect 5075 5305 5080 5335
rect 5110 5305 5115 5335
rect 5075 5300 5115 5305
rect 5505 4720 5525 5380
rect 5960 5335 6000 5340
rect 5960 5305 5965 5335
rect 5995 5305 6000 5335
rect 5960 5300 6000 5305
rect 5495 4715 5535 4720
rect 5495 4685 5500 4715
rect 5530 4685 5535 4715
rect 5495 4680 5535 4685
rect 5970 3530 5990 5300
rect 6105 3685 6125 6650
rect 6785 5090 6805 6655
rect 7020 6650 7060 6655
rect 7100 6685 7140 6690
rect 7100 6655 7105 6685
rect 7135 6655 7140 6685
rect 7100 6650 7140 6655
rect 6410 5085 6450 5090
rect 6410 5055 6415 5085
rect 6445 5055 6450 5085
rect 6410 5050 6450 5055
rect 6775 5085 6815 5090
rect 6775 5055 6780 5085
rect 6810 5055 6815 5085
rect 6775 5050 6815 5055
rect 6420 4775 6440 5050
rect 6410 4770 6450 4775
rect 6410 4740 6415 4770
rect 6445 4740 6450 4770
rect 6410 4735 6450 4740
rect 6095 3680 6135 3685
rect 6095 3650 6100 3680
rect 6130 3650 6135 3680
rect 6095 3645 6135 3650
rect 5885 3525 5925 3530
rect 5885 3495 5890 3525
rect 5920 3495 5925 3525
rect 5885 3490 5925 3495
rect 5960 3525 6000 3530
rect 5960 3495 5965 3525
rect 5995 3495 6000 3525
rect 5960 3490 6000 3495
rect 5895 3030 5915 3490
rect 7110 3140 7130 6650
rect 7145 6580 7185 6585
rect 7145 6550 7150 6580
rect 7180 6550 7185 6580
rect 7145 6545 7185 6550
rect 6995 3135 7035 3140
rect 6995 3105 7000 3135
rect 7030 3105 7035 3135
rect 7100 3135 7140 3140
rect 7100 3105 7105 3135
rect 7135 3105 7140 3135
rect 5095 3025 5135 3030
rect 5095 2995 5100 3025
rect 5130 2995 5135 3025
rect 5095 2990 5135 2995
rect 5885 3025 5925 3030
rect 5885 2995 5890 3025
rect 5920 2995 5925 3025
rect 5885 2990 5925 2995
rect 5105 2700 5125 2990
rect 7005 2755 7025 3105
rect 7155 3090 7175 6545
rect 7040 3085 7080 3090
rect 7040 3055 7045 3085
rect 7075 3055 7080 3085
rect 7040 3050 7080 3055
rect 7145 3085 7185 3090
rect 7145 3055 7150 3085
rect 7180 3055 7185 3085
rect 7145 3050 7185 3055
rect 7050 2865 7070 3050
rect 2440 1800 2480 1830
<< via1 >>
rect 2955 6655 2985 6685
rect 3035 6655 3065 6685
rect 6100 6655 6130 6685
rect 2910 6550 2940 6580
rect 3405 6615 3435 6645
rect 3275 6490 3305 6520
rect 3960 6615 3990 6645
rect 3550 6445 3580 6475
rect 4335 6550 4365 6580
rect 4005 6445 4035 6475
rect 4005 5370 4035 5400
rect 4095 5370 4125 5400
rect 3985 3745 4015 3775
rect 4005 3605 4035 3635
rect 2955 3105 2985 3135
rect 3060 3105 3090 3135
rect 2910 3055 2940 3085
rect 3015 3055 3045 3085
rect 6705 6655 6735 6685
rect 7025 6655 7055 6685
rect 5725 6550 5755 6580
rect 5380 6490 5410 6520
rect 5380 5385 5410 5415
rect 5500 5385 5530 5415
rect 5080 5305 5110 5335
rect 5965 5305 5995 5335
rect 5500 4685 5530 4715
rect 7105 6655 7135 6685
rect 6415 5055 6445 5085
rect 6780 5055 6810 5085
rect 6415 4740 6445 4770
rect 6100 3650 6130 3680
rect 5890 3495 5920 3525
rect 5965 3495 5995 3525
rect 7150 6550 7180 6580
rect 7000 3105 7030 3135
rect 7105 3105 7135 3135
rect 5100 2995 5130 3025
rect 5890 2995 5920 3025
rect 7045 3055 7075 3085
rect 7150 3055 7180 3085
<< metal2 >>
rect 2950 6685 2990 6690
rect 2950 6655 2955 6685
rect 2985 6680 2990 6685
rect 3030 6685 3070 6690
rect 3030 6680 3035 6685
rect 2985 6660 3035 6680
rect 2985 6655 2990 6660
rect 2950 6650 2990 6655
rect 3030 6655 3035 6660
rect 3065 6655 3070 6685
rect 3030 6650 3070 6655
rect 6095 6685 6135 6690
rect 6095 6655 6100 6685
rect 6130 6680 6135 6685
rect 6700 6685 6740 6690
rect 6700 6680 6705 6685
rect 6130 6660 6705 6680
rect 6130 6655 6135 6660
rect 6095 6650 6135 6655
rect 6700 6655 6705 6660
rect 6735 6655 6740 6685
rect 6700 6650 6740 6655
rect 7020 6685 7060 6690
rect 7020 6655 7025 6685
rect 7055 6680 7060 6685
rect 7100 6685 7140 6690
rect 7100 6680 7105 6685
rect 7055 6660 7105 6680
rect 7055 6655 7060 6660
rect 7020 6650 7060 6655
rect 7100 6655 7105 6660
rect 7135 6655 7140 6685
rect 7100 6650 7140 6655
rect 3400 6645 3440 6650
rect 3400 6615 3405 6645
rect 3435 6640 3440 6645
rect 3955 6645 3995 6650
rect 3955 6640 3960 6645
rect 3435 6620 3960 6640
rect 3435 6615 3440 6620
rect 3400 6610 3440 6615
rect 3955 6615 3960 6620
rect 3990 6615 3995 6645
rect 3955 6610 3995 6615
rect 2905 6580 2945 6585
rect 2905 6550 2910 6580
rect 2940 6575 2945 6580
rect 4330 6580 4370 6585
rect 4330 6575 4335 6580
rect 2940 6555 4335 6575
rect 2940 6550 2945 6555
rect 2905 6545 2945 6550
rect 4330 6550 4335 6555
rect 4365 6550 4370 6580
rect 4330 6545 4370 6550
rect 5720 6580 5760 6585
rect 5720 6550 5725 6580
rect 5755 6575 5760 6580
rect 7145 6580 7185 6585
rect 7145 6575 7150 6580
rect 5755 6555 7150 6575
rect 5755 6550 5760 6555
rect 5720 6545 5760 6550
rect 7145 6550 7150 6555
rect 7180 6550 7185 6580
rect 7145 6545 7185 6550
rect 3270 6520 3310 6525
rect 3270 6490 3275 6520
rect 3305 6515 3310 6520
rect 5375 6520 5415 6525
rect 5375 6515 5380 6520
rect 3305 6495 5380 6515
rect 3305 6490 3310 6495
rect 3270 6485 3310 6490
rect 5375 6490 5380 6495
rect 5410 6490 5415 6520
rect 5375 6485 5415 6490
rect 3545 6475 3585 6480
rect 3545 6445 3550 6475
rect 3580 6470 3585 6475
rect 4000 6475 4040 6480
rect 4000 6470 4005 6475
rect 3580 6450 4005 6470
rect 3580 6445 3585 6450
rect 3545 6440 3585 6445
rect 4000 6445 4005 6450
rect 4035 6445 4040 6475
rect 4000 6440 4040 6445
rect 5375 5415 5415 5420
rect 4000 5400 4040 5405
rect 4000 5370 4005 5400
rect 4035 5395 4040 5400
rect 4090 5400 4130 5405
rect 4090 5395 4095 5400
rect 4035 5375 4095 5395
rect 4035 5370 4040 5375
rect 4000 5365 4040 5370
rect 4090 5370 4095 5375
rect 4125 5370 4130 5400
rect 5375 5385 5380 5415
rect 5410 5410 5415 5415
rect 5495 5415 5535 5420
rect 5495 5410 5500 5415
rect 5410 5390 5500 5410
rect 5410 5385 5415 5390
rect 5375 5380 5415 5385
rect 5495 5385 5500 5390
rect 5530 5385 5535 5415
rect 5495 5380 5535 5385
rect 4090 5365 4130 5370
rect 5075 5335 5115 5340
rect 5075 5305 5080 5335
rect 5110 5330 5115 5335
rect 5960 5335 6000 5340
rect 5960 5330 5965 5335
rect 5110 5310 5965 5330
rect 5110 5305 5115 5310
rect 5075 5300 5115 5305
rect 5960 5305 5965 5310
rect 5995 5305 6000 5335
rect 5960 5300 6000 5305
rect 6410 5085 6450 5090
rect 6410 5055 6415 5085
rect 6445 5080 6450 5085
rect 6775 5085 6815 5090
rect 6775 5080 6780 5085
rect 6445 5060 6780 5080
rect 6445 5055 6450 5060
rect 6410 5050 6450 5055
rect 6775 5055 6780 5060
rect 6810 5055 6815 5085
rect 6775 5050 6815 5055
rect 6410 4770 6450 4775
rect 6410 4765 6415 4770
rect 5745 4745 6415 4765
rect 6410 4740 6415 4745
rect 6445 4740 6450 4770
rect 6410 4735 6450 4740
rect 5495 4715 5535 4720
rect 5495 4685 5500 4715
rect 5530 4685 5535 4715
rect 5495 4680 5535 4685
rect 3980 3775 4020 3780
rect 3980 3745 3985 3775
rect 4015 3745 4020 3775
rect 3980 3740 4020 3745
rect 6095 3680 6135 3685
rect 6095 3675 6100 3680
rect 5270 3655 6100 3675
rect 6095 3650 6100 3655
rect 6130 3650 6135 3680
rect 6095 3645 6135 3650
rect 4000 3635 4040 3640
rect 4000 3605 4005 3635
rect 4035 3630 4040 3635
rect 4035 3610 4110 3630
rect 4035 3605 4040 3610
rect 5885 3525 5925 3530
rect 5885 3495 5890 3525
rect 5920 3520 5925 3525
rect 5960 3525 6000 3530
rect 5960 3520 5965 3525
rect 5920 3500 5965 3520
rect 5920 3495 5925 3500
rect 5885 3490 5925 3495
rect 5960 3495 5965 3500
rect 5995 3495 6000 3525
rect 5960 3490 6000 3495
rect 2950 3135 2990 3140
rect 2950 3105 2955 3135
rect 2985 3130 2990 3135
rect 3055 3135 3095 3140
rect 3055 3130 3060 3135
rect 2985 3110 3060 3130
rect 2985 3105 2990 3110
rect 3055 3105 3060 3110
rect 3090 3105 3095 3135
rect 6995 3135 7035 3140
rect 6995 3105 7000 3135
rect 7030 3130 7035 3135
rect 7100 3135 7140 3140
rect 7100 3130 7105 3135
rect 7030 3110 7105 3130
rect 7030 3105 7035 3110
rect 7100 3105 7105 3110
rect 7135 3105 7140 3135
rect 2905 3085 2945 3090
rect 2905 3055 2910 3085
rect 2940 3080 2945 3085
rect 3010 3085 3050 3090
rect 3010 3080 3015 3085
rect 2940 3060 3015 3080
rect 2940 3055 2945 3060
rect 2905 3050 2945 3055
rect 3010 3055 3015 3060
rect 3045 3055 3050 3085
rect 3010 3050 3050 3055
rect 7040 3085 7080 3090
rect 7040 3055 7045 3085
rect 7075 3080 7080 3085
rect 7145 3085 7185 3090
rect 7145 3080 7150 3085
rect 7075 3060 7150 3080
rect 7075 3055 7080 3060
rect 7040 3050 7080 3055
rect 7145 3055 7150 3060
rect 7180 3055 7185 3085
rect 7145 3050 7185 3055
rect 5095 3025 5135 3030
rect 5095 2995 5100 3025
rect 5130 3020 5135 3025
rect 5885 3025 5925 3030
rect 5885 3020 5890 3025
rect 5130 3000 5890 3020
rect 5130 2995 5135 3000
rect 5095 2990 5135 2995
rect 5885 2995 5890 3000
rect 5920 2995 5925 3025
rect 5885 2990 5925 2995
rect 4150 2460 4170 2480
rect 4150 2240 4170 2260
rect 2815 2140 2835 2160
rect 7220 2140 7240 2160
rect 2440 1800 2480 1830
<< metal3 >>
rect 9335 14460 9385 14465
rect 9335 14420 9340 14460
rect 9380 14420 9385 14460
rect 9335 14415 9385 14420
rect 9340 50 9380 14415
rect 9335 45 9385 50
rect 9335 5 9340 45
rect 9380 5 9385 45
rect 9335 0 9385 5
<< via3 >>
rect 9340 14420 9380 14460
rect 9340 5 9380 45
<< metal4 >>
rect 7255 14460 9385 14465
rect 7255 14420 9340 14460
rect 9380 14420 9385 14460
rect 7255 14415 9385 14420
rect 540 6700 590 6750
rect 540 0 590 50
rect 9325 45 9385 50
rect 9325 5 9340 45
rect 9380 5 9385 45
rect 9325 0 9385 5
use bgr  bgr_0
timestamp 1752209448
transform -1 0 22845 0 -1 8250
box 15505 -6295 20095 1600
use two_stage_opamp_dummy_magic_14  two_stage_opamp_dummy_magic_14_0
timestamp 1752398166
transform 1 0 4200 0 1 2465
box -3850 -2465 5140 4285
<< labels >>
flabel metal4 565 6750 565 6750 1 FreeSans 800 0 0 320 VDDA
port 1 n
flabel metal4 565 0 565 0 5 FreeSans 800 0 0 -320 GNDA
port 2 s
flabel metal2 2825 2140 2825 2140 5 FreeSans 800 0 0 -320 VOUT+
port 3 s
flabel metal2 7230 2140 7230 2140 5 FreeSans 800 0 0 -320 VOUT-
port 4 s
flabel metal2 4150 2470 4150 2470 7 FreeSans 800 0 -320 0 VIN-
port 6 w
flabel metal2 4150 2250 4150 2250 7 FreeSans 800 0 -320 0 VIN+
port 5 w
<< end >>
