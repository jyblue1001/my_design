magic
tech sky130A
timestamp 1737911406
<< nmos >>
rect 1070 460 1120 710
rect 1170 460 1220 710
rect 1270 460 1320 710
rect 1370 460 1420 710
rect 1470 460 1520 710
rect 1570 460 1620 710
rect 1670 460 1720 710
rect 1770 460 1820 710
rect 1050 245 1065 345
rect 1115 245 1130 345
rect 1180 245 1195 345
rect 1245 245 1260 345
rect 1410 245 1425 345
rect 1475 245 1490 345
rect 1540 245 1555 345
rect 1605 245 1620 345
rect 1790 245 1805 345
rect 1855 245 1870 345
rect 1920 245 1935 345
rect 1985 245 2000 345
rect 1050 50 1065 100
rect 1115 50 1130 100
rect 1180 50 1195 100
rect 1245 50 1260 100
rect 1410 50 1425 100
rect 1475 50 1490 100
rect 1540 50 1555 100
rect 1605 50 1620 100
rect 1790 50 1805 100
rect 1855 50 1870 100
rect 1920 50 1935 100
rect 1985 50 2000 100
rect 1615 -345 1665 -95
rect 1715 -345 1765 -95
rect 1815 -345 1865 -95
rect 1915 -345 1965 -95
<< ndiff >>
rect 1020 695 1070 710
rect 1020 475 1035 695
rect 1055 475 1070 695
rect 1020 460 1070 475
rect 1120 695 1170 710
rect 1120 475 1135 695
rect 1155 475 1170 695
rect 1120 460 1170 475
rect 1220 695 1270 710
rect 1220 475 1235 695
rect 1255 475 1270 695
rect 1220 460 1270 475
rect 1320 695 1370 710
rect 1320 475 1335 695
rect 1355 475 1370 695
rect 1320 460 1370 475
rect 1420 695 1470 710
rect 1420 475 1435 695
rect 1455 475 1470 695
rect 1420 460 1470 475
rect 1520 695 1570 710
rect 1520 475 1535 695
rect 1555 475 1570 695
rect 1520 460 1570 475
rect 1620 695 1670 710
rect 1620 475 1635 695
rect 1655 475 1670 695
rect 1620 460 1670 475
rect 1720 695 1770 710
rect 1720 475 1735 695
rect 1755 475 1770 695
rect 1720 460 1770 475
rect 1820 695 1870 710
rect 1820 475 1835 695
rect 1855 475 1870 695
rect 1820 460 1870 475
rect 1000 330 1050 345
rect 1000 260 1015 330
rect 1035 260 1050 330
rect 1000 245 1050 260
rect 1065 330 1115 345
rect 1065 260 1080 330
rect 1100 260 1115 330
rect 1065 245 1115 260
rect 1130 330 1180 345
rect 1130 260 1145 330
rect 1165 260 1180 330
rect 1130 245 1180 260
rect 1195 330 1245 345
rect 1195 260 1210 330
rect 1230 260 1245 330
rect 1195 245 1245 260
rect 1260 330 1310 345
rect 1360 330 1410 345
rect 1260 260 1275 330
rect 1295 260 1310 330
rect 1360 260 1375 330
rect 1395 260 1410 330
rect 1260 245 1310 260
rect 1360 245 1410 260
rect 1425 330 1475 345
rect 1425 260 1440 330
rect 1460 260 1475 330
rect 1425 245 1475 260
rect 1490 330 1540 345
rect 1490 260 1505 330
rect 1525 260 1540 330
rect 1490 245 1540 260
rect 1555 330 1605 345
rect 1555 260 1570 330
rect 1590 260 1605 330
rect 1555 245 1605 260
rect 1620 330 1670 345
rect 1620 260 1635 330
rect 1655 260 1670 330
rect 1620 245 1670 260
rect 1740 330 1790 345
rect 1740 260 1755 330
rect 1775 260 1790 330
rect 1740 245 1790 260
rect 1805 330 1855 345
rect 1805 260 1820 330
rect 1840 260 1855 330
rect 1805 245 1855 260
rect 1870 330 1920 345
rect 1870 260 1885 330
rect 1905 260 1920 330
rect 1870 245 1920 260
rect 1935 330 1985 345
rect 1935 260 1950 330
rect 1970 260 1985 330
rect 1935 245 1985 260
rect 2000 330 2050 345
rect 2000 260 2015 330
rect 2035 260 2050 330
rect 2000 245 2050 260
rect 1000 85 1050 100
rect 1000 65 1015 85
rect 1035 65 1050 85
rect 1000 50 1050 65
rect 1065 85 1115 100
rect 1065 65 1080 85
rect 1100 65 1115 85
rect 1065 50 1115 65
rect 1130 85 1180 100
rect 1130 65 1145 85
rect 1165 65 1180 85
rect 1130 50 1180 65
rect 1195 85 1245 100
rect 1195 65 1210 85
rect 1230 65 1245 85
rect 1195 50 1245 65
rect 1260 85 1310 100
rect 1360 85 1410 100
rect 1260 65 1275 85
rect 1295 65 1310 85
rect 1360 65 1375 85
rect 1395 65 1410 85
rect 1260 50 1310 65
rect 1360 50 1410 65
rect 1425 85 1475 100
rect 1425 65 1440 85
rect 1460 65 1475 85
rect 1425 50 1475 65
rect 1490 85 1540 100
rect 1490 65 1505 85
rect 1525 65 1540 85
rect 1490 50 1540 65
rect 1555 85 1605 100
rect 1555 65 1570 85
rect 1590 65 1605 85
rect 1555 50 1605 65
rect 1620 85 1670 100
rect 1620 65 1635 85
rect 1655 65 1670 85
rect 1620 50 1670 65
rect 1740 85 1790 100
rect 1740 65 1755 85
rect 1775 65 1790 85
rect 1740 50 1790 65
rect 1805 85 1855 100
rect 1805 65 1820 85
rect 1840 65 1855 85
rect 1805 50 1855 65
rect 1870 85 1920 100
rect 1870 65 1885 85
rect 1905 65 1920 85
rect 1870 50 1920 65
rect 1935 85 1985 100
rect 1935 65 1950 85
rect 1970 65 1985 85
rect 1935 50 1985 65
rect 2000 85 2050 100
rect 2000 65 2015 85
rect 2035 65 2050 85
rect 2000 50 2050 65
rect 1565 -110 1615 -95
rect 1565 -330 1580 -110
rect 1600 -330 1615 -110
rect 1565 -345 1615 -330
rect 1665 -110 1715 -95
rect 1665 -330 1680 -110
rect 1700 -330 1715 -110
rect 1665 -345 1715 -330
rect 1765 -110 1815 -95
rect 1765 -330 1780 -110
rect 1800 -330 1815 -110
rect 1765 -345 1815 -330
rect 1865 -110 1915 -95
rect 1865 -330 1880 -110
rect 1900 -330 1915 -110
rect 1865 -345 1915 -330
rect 1965 -110 2015 -95
rect 1965 -330 1980 -110
rect 2000 -330 2015 -110
rect 1965 -345 2015 -330
<< ndiffc >>
rect 1035 475 1055 695
rect 1135 475 1155 695
rect 1235 475 1255 695
rect 1335 475 1355 695
rect 1435 475 1455 695
rect 1535 475 1555 695
rect 1635 475 1655 695
rect 1735 475 1755 695
rect 1835 475 1855 695
rect 1015 260 1035 330
rect 1080 260 1100 330
rect 1145 260 1165 330
rect 1210 260 1230 330
rect 1275 260 1295 330
rect 1375 260 1395 330
rect 1440 260 1460 330
rect 1505 260 1525 330
rect 1570 260 1590 330
rect 1635 260 1655 330
rect 1755 260 1775 330
rect 1820 260 1840 330
rect 1885 260 1905 330
rect 1950 260 1970 330
rect 2015 260 2035 330
rect 1015 65 1035 85
rect 1080 65 1100 85
rect 1145 65 1165 85
rect 1210 65 1230 85
rect 1275 65 1295 85
rect 1375 65 1395 85
rect 1440 65 1460 85
rect 1505 65 1525 85
rect 1570 65 1590 85
rect 1635 65 1655 85
rect 1755 65 1775 85
rect 1820 65 1840 85
rect 1885 65 1905 85
rect 1950 65 1970 85
rect 2015 65 2035 85
rect 1580 -330 1600 -110
rect 1680 -330 1700 -110
rect 1780 -330 1800 -110
rect 1880 -330 1900 -110
rect 1980 -330 2000 -110
<< psubdiff >>
rect 1310 330 1360 345
rect 1310 260 1325 330
rect 1345 260 1360 330
rect 1310 245 1360 260
rect 1310 85 1360 100
rect 1310 65 1325 85
rect 1345 65 1360 85
rect 1310 50 1360 65
<< psubdiffcont >>
rect 1325 260 1345 330
rect 1325 65 1345 85
<< poly >>
rect 1075 755 1115 765
rect 1075 740 1085 755
rect 1070 735 1085 740
rect 1105 740 1115 755
rect 1425 755 1465 765
rect 1425 740 1435 755
rect 1105 735 1435 740
rect 1455 740 1465 755
rect 1775 755 1815 765
rect 1775 740 1785 755
rect 1455 735 1785 740
rect 1805 740 1815 755
rect 1805 735 1820 740
rect 1070 725 1820 735
rect 1070 710 1120 725
rect 1170 710 1220 725
rect 1270 710 1320 725
rect 1370 710 1420 725
rect 1470 710 1520 725
rect 1570 710 1620 725
rect 1670 710 1720 725
rect 1770 710 1820 725
rect 1070 445 1120 460
rect 1170 445 1220 460
rect 1270 445 1320 460
rect 1370 445 1420 460
rect 1470 445 1520 460
rect 1570 445 1620 460
rect 1670 445 1720 460
rect 1770 445 1820 460
rect 855 385 1195 400
rect 1050 345 1065 360
rect 1115 345 1130 360
rect 1180 345 1195 385
rect 1400 390 1440 400
rect 1400 370 1410 390
rect 1430 370 1440 390
rect 1585 390 1625 400
rect 1585 370 1595 390
rect 1615 370 1625 390
rect 1400 360 1625 370
rect 1245 345 1260 360
rect 1410 355 1620 360
rect 1410 345 1425 355
rect 1475 345 1490 355
rect 1540 345 1555 355
rect 1605 345 1620 355
rect 1790 345 1805 360
rect 1855 345 1870 360
rect 1920 345 1935 360
rect 1985 345 2000 360
rect 1050 235 1065 245
rect 1115 235 1130 245
rect 975 220 1130 235
rect 1180 235 1195 245
rect 1245 235 1260 245
rect 1180 220 1300 235
rect 1410 230 1425 245
rect 1475 230 1490 245
rect 1540 230 1555 245
rect 1605 230 1620 245
rect 1685 240 1725 250
rect 2065 250 2105 260
rect 975 -30 990 220
rect 1285 125 1300 220
rect 1685 220 1695 240
rect 1715 235 1725 240
rect 1790 235 1805 245
rect 1855 235 1870 245
rect 1920 235 1935 245
rect 1985 235 2000 245
rect 2065 235 2075 250
rect 1715 230 2075 235
rect 2095 230 2105 250
rect 1715 220 2105 230
rect 1685 210 1725 220
rect 1380 180 1420 190
rect 1380 160 1390 180
rect 1410 165 1490 180
rect 1410 160 1420 165
rect 1380 150 1420 160
rect 1475 155 1490 165
rect 1475 140 1725 155
rect 1050 100 1065 115
rect 1115 100 1130 115
rect 1180 100 1195 115
rect 1245 100 1260 115
rect 1285 110 1425 125
rect 1685 120 1695 140
rect 1715 125 1725 140
rect 1715 120 2105 125
rect 1685 115 2105 120
rect 1410 100 1425 110
rect 1475 100 1490 115
rect 1540 100 1555 115
rect 1605 100 1620 115
rect 1685 110 2075 115
rect 1790 100 1805 110
rect 1855 100 1870 110
rect 1920 100 1935 110
rect 1985 100 2000 110
rect 2065 95 2075 110
rect 2095 95 2105 115
rect 2065 85 2105 95
rect 1050 40 1065 50
rect 1115 40 1130 50
rect 1180 40 1195 50
rect 1245 40 1260 50
rect 1040 35 1260 40
rect 1410 40 1425 50
rect 1475 40 1490 50
rect 1040 25 1270 35
rect 1410 25 1490 40
rect 1540 40 1555 50
rect 1605 40 1620 50
rect 1540 25 1620 40
rect 1790 35 1805 50
rect 1855 35 1870 50
rect 1920 35 1935 50
rect 1985 35 2000 50
rect 1040 5 1050 25
rect 1070 20 1240 25
rect 1070 5 1080 20
rect 1040 -5 1080 5
rect 1230 5 1240 20
rect 1260 5 1270 25
rect 1230 -5 1270 5
rect 1540 -30 1555 25
rect 860 -45 1555 -30
rect 1615 -95 1665 -80
rect 1715 -95 1765 -80
rect 1815 -95 1865 -80
rect 1915 -95 1965 -80
rect 1615 -360 1665 -345
rect 1715 -360 1765 -345
rect 1815 -360 1865 -345
rect 1915 -360 1965 -345
rect 1615 -370 1965 -360
rect 1615 -375 1630 -370
rect 1620 -390 1630 -375
rect 1650 -375 1930 -370
rect 1650 -390 1660 -375
rect 1620 -400 1660 -390
rect 1920 -390 1930 -375
rect 1950 -375 1965 -370
rect 1950 -390 1960 -375
rect 1920 -400 1960 -390
<< polycont >>
rect 1085 735 1105 755
rect 1435 735 1455 755
rect 1785 735 1805 755
rect 1410 370 1430 390
rect 1595 370 1615 390
rect 1695 220 1715 240
rect 2075 230 2095 250
rect 1390 160 1410 180
rect 1695 120 1715 140
rect 2075 95 2095 115
rect 1050 5 1070 25
rect 1240 5 1260 25
rect 1630 -390 1650 -370
rect 1930 -390 1950 -370
<< xpolycontact >>
rect 2070 745 2105 965
rect 2070 410 2105 630
rect 1020 -380 1240 -95
rect 1290 -380 1510 -95
rect 2070 -230 2105 -10
rect 2070 -535 2105 -315
<< xpolyres >>
rect 2070 630 2105 745
rect 1240 -380 1290 -95
rect 2070 -315 2105 -230
<< locali >>
rect 2125 1070 2165 1080
rect 2085 1050 2135 1070
rect 2155 1050 2165 1070
rect 2085 965 2105 1050
rect 2125 1040 2165 1050
rect 1075 755 1115 765
rect 1075 745 1085 755
rect 965 735 1085 745
rect 1105 745 1115 755
rect 1425 755 1465 765
rect 1425 745 1435 755
rect 1105 735 1435 745
rect 1455 745 1465 755
rect 1775 755 1815 765
rect 1775 745 1785 755
rect 1455 735 1785 745
rect 1805 745 1815 755
rect 1805 735 1855 745
rect 965 725 1855 735
rect 965 -95 985 725
rect 1035 705 1055 725
rect 1435 705 1455 725
rect 1835 705 1855 725
rect 1025 695 1065 705
rect 1025 475 1035 695
rect 1055 475 1065 695
rect 1025 465 1065 475
rect 1125 695 1165 705
rect 1125 475 1135 695
rect 1155 475 1165 695
rect 1125 465 1165 475
rect 1225 695 1265 705
rect 1225 475 1235 695
rect 1255 475 1265 695
rect 1225 465 1265 475
rect 1325 695 1365 705
rect 1325 475 1335 695
rect 1355 475 1365 695
rect 1325 465 1365 475
rect 1425 695 1465 705
rect 1425 475 1435 695
rect 1455 475 1465 695
rect 1425 465 1465 475
rect 1525 695 1565 705
rect 1525 475 1535 695
rect 1555 475 1565 695
rect 1525 465 1565 475
rect 1625 695 1665 705
rect 1625 475 1635 695
rect 1655 475 1665 695
rect 1625 465 1665 475
rect 1725 695 1765 705
rect 1725 475 1735 695
rect 1755 475 1765 695
rect 1725 465 1765 475
rect 1825 695 1865 705
rect 1825 475 1835 695
rect 1855 475 1865 695
rect 1825 465 1865 475
rect 1235 440 1255 465
rect 1635 440 1655 465
rect 1235 420 1655 440
rect 1235 380 1255 420
rect 1400 390 1440 400
rect 1400 380 1410 390
rect 1015 360 1295 380
rect 1015 340 1035 360
rect 1145 340 1165 360
rect 1275 340 1295 360
rect 1375 370 1410 380
rect 1430 380 1440 390
rect 1585 390 1625 400
rect 1585 380 1595 390
rect 1430 370 1595 380
rect 1615 380 1625 390
rect 2085 380 2105 410
rect 1615 370 1655 380
rect 1375 360 1655 370
rect 1375 340 1395 360
rect 1635 340 1655 360
rect 1820 360 2105 380
rect 1820 340 1840 360
rect 1950 340 1970 360
rect 1005 330 1045 340
rect 1005 260 1015 330
rect 1035 260 1045 330
rect 1005 250 1045 260
rect 1070 330 1110 340
rect 1070 260 1080 330
rect 1100 260 1110 330
rect 1070 250 1110 260
rect 1135 330 1175 340
rect 1135 260 1145 330
rect 1165 260 1175 330
rect 1135 250 1175 260
rect 1200 330 1240 340
rect 1200 260 1210 330
rect 1230 260 1240 330
rect 1200 250 1240 260
rect 1265 330 1405 340
rect 1265 260 1275 330
rect 1295 260 1325 330
rect 1345 260 1375 330
rect 1395 260 1405 330
rect 1265 250 1405 260
rect 1430 330 1470 340
rect 1430 260 1440 330
rect 1460 260 1470 330
rect 1430 250 1470 260
rect 1495 330 1535 340
rect 1495 260 1505 330
rect 1525 260 1535 330
rect 1495 250 1535 260
rect 1560 330 1600 340
rect 1560 260 1570 330
rect 1590 260 1600 330
rect 1560 250 1600 260
rect 1625 330 1665 340
rect 1625 260 1635 330
rect 1655 260 1665 330
rect 1625 250 1665 260
rect 1745 330 1785 340
rect 1745 260 1755 330
rect 1775 260 1785 330
rect 1745 250 1785 260
rect 1810 330 1850 340
rect 1810 260 1820 330
rect 1840 260 1850 330
rect 1810 250 1850 260
rect 1875 330 1915 340
rect 1875 260 1885 330
rect 1905 260 1915 330
rect 1875 250 1915 260
rect 1940 330 1980 340
rect 1940 260 1950 330
rect 1970 260 1980 330
rect 1940 250 1980 260
rect 2005 330 2045 340
rect 2005 260 2015 330
rect 2035 260 2045 330
rect 2085 260 2105 360
rect 2005 250 2045 260
rect 2065 250 2105 260
rect 1080 230 1100 250
rect 1210 230 1230 250
rect 1015 210 1100 230
rect 1145 210 1230 230
rect 1375 230 1395 250
rect 1505 230 1525 250
rect 1685 240 1725 250
rect 1685 230 1695 240
rect 1375 210 1460 230
rect 1505 220 1695 230
rect 1715 220 1725 240
rect 2065 230 2075 250
rect 2095 240 2105 250
rect 2125 305 2165 315
rect 2125 285 2135 305
rect 2155 285 2165 305
rect 2125 275 2165 285
rect 2125 240 2145 275
rect 2095 230 2145 240
rect 2065 220 2145 230
rect 1505 210 1725 220
rect 1015 95 1035 210
rect 1145 180 1165 210
rect 1380 180 1420 190
rect 1145 160 1390 180
rect 1410 160 1420 180
rect 1145 95 1165 160
rect 1380 150 1420 160
rect 1440 95 1460 210
rect 1570 95 1590 210
rect 2125 195 2145 220
rect 2125 175 3055 195
rect 1685 140 1725 155
rect 1685 120 1695 140
rect 1715 120 1725 140
rect 2125 125 2145 175
rect 1685 110 1725 120
rect 2065 115 2145 125
rect 2065 95 2075 115
rect 2095 105 2145 115
rect 2095 95 2105 105
rect 1005 85 1045 95
rect 1005 65 1015 85
rect 1035 65 1045 85
rect 1005 55 1045 65
rect 1070 85 1110 95
rect 1070 65 1080 85
rect 1100 65 1110 85
rect 1070 55 1110 65
rect 1135 85 1175 95
rect 1135 65 1145 85
rect 1165 65 1175 85
rect 1135 55 1175 65
rect 1200 85 1240 95
rect 1200 65 1210 85
rect 1230 65 1240 85
rect 1200 55 1240 65
rect 1265 85 1405 95
rect 1265 65 1275 85
rect 1295 65 1325 85
rect 1345 65 1375 85
rect 1395 65 1405 85
rect 1265 55 1405 65
rect 1430 85 1470 95
rect 1430 65 1440 85
rect 1460 65 1470 85
rect 1430 55 1470 65
rect 1495 85 1535 95
rect 1495 65 1505 85
rect 1525 65 1535 85
rect 1495 55 1535 65
rect 1560 85 1600 95
rect 1560 65 1570 85
rect 1590 65 1600 85
rect 1560 55 1600 65
rect 1625 85 1665 95
rect 1625 65 1635 85
rect 1655 65 1665 85
rect 1625 55 1665 65
rect 1745 85 1785 95
rect 1745 65 1755 85
rect 1775 65 1785 85
rect 1745 55 1785 65
rect 1810 85 1850 95
rect 1810 65 1820 85
rect 1840 65 1850 85
rect 1810 55 1850 65
rect 1875 85 1915 95
rect 1875 65 1885 85
rect 1905 65 1915 85
rect 1875 55 1915 65
rect 1940 85 1980 95
rect 1940 65 1950 85
rect 1970 65 1980 85
rect 1940 55 1980 65
rect 2005 85 2045 95
rect 2065 85 2105 95
rect 2005 65 2015 85
rect 2035 65 2045 85
rect 2005 55 2045 65
rect 1015 35 1035 55
rect 1275 35 1295 55
rect 1015 25 1295 35
rect 1015 15 1050 25
rect 1040 5 1050 15
rect 1070 15 1240 25
rect 1070 5 1080 15
rect 1040 -5 1080 5
rect 1230 5 1240 15
rect 1260 15 1295 25
rect 1375 35 1395 55
rect 1505 35 1525 55
rect 1635 35 1655 55
rect 1820 35 1840 55
rect 1950 35 1970 55
rect 2085 35 2105 85
rect 1375 15 1700 35
rect 1820 15 2105 35
rect 2125 70 2145 105
rect 2125 60 2165 70
rect 2125 40 2135 60
rect 2155 40 2165 60
rect 2125 30 2165 40
rect 1260 5 1270 15
rect 1230 -5 1270 5
rect 1680 -20 1700 15
rect 2085 -10 2105 15
rect 1680 -45 1800 -20
rect 965 -115 1020 -95
rect 1780 -100 1800 -45
rect 1570 -110 1610 -100
rect 1570 -330 1580 -110
rect 1600 -330 1610 -110
rect 1570 -340 1610 -330
rect 1670 -110 1710 -100
rect 1670 -330 1680 -110
rect 1700 -330 1710 -110
rect 1670 -340 1710 -330
rect 1770 -110 1810 -100
rect 1770 -330 1780 -110
rect 1800 -330 1810 -110
rect 1770 -340 1810 -330
rect 1870 -110 1910 -100
rect 1870 -330 1880 -110
rect 1900 -330 1910 -110
rect 1870 -340 1910 -330
rect 1970 -110 2010 -100
rect 1970 -330 1980 -110
rect 2000 -330 2010 -110
rect 1970 -340 2010 -330
rect 1580 -360 1600 -340
rect 1980 -360 2000 -340
rect 1510 -370 2000 -360
rect 1510 -380 1630 -370
rect 1620 -390 1630 -380
rect 1650 -380 1930 -370
rect 1650 -390 1660 -380
rect 1620 -400 1660 -390
rect 1920 -390 1930 -380
rect 1950 -380 2000 -370
rect 1950 -390 1960 -380
rect 1920 -400 1960 -390
rect 2085 -705 2105 -535
rect 2125 -705 2165 -695
rect 2085 -725 2135 -705
rect 2155 -725 2165 -705
rect 2125 -735 2165 -725
<< viali >>
rect 2135 1050 2155 1070
rect 2135 285 2155 305
rect 2135 40 2155 60
rect 2135 -725 2155 -705
<< metal1 >>
rect 2125 1070 2165 1080
rect 2125 1050 2135 1070
rect 2155 1050 2165 1070
rect 2125 1040 2165 1050
rect 2125 305 2165 315
rect 2125 285 2135 305
rect 2155 285 2165 305
rect 2125 275 2165 285
rect 2125 60 2165 70
rect 2125 40 2135 60
rect 2155 40 2165 60
rect 2125 30 2165 40
rect 2125 -705 2165 -695
rect 2125 -725 2135 -705
rect 2155 -725 2165 -705
rect 2125 -735 2165 -725
<< metal3 >>
rect 2125 1040 3010 1085
rect 2180 255 3010 1040
rect 2180 -695 3010 90
rect 2125 -740 3010 -695
<< mimcap >>
rect 2195 315 2995 1070
rect 2195 280 2205 315
rect 2240 280 2995 315
rect 2195 270 2995 280
rect 2195 65 2995 75
rect 2195 30 2205 65
rect 2240 30 2995 65
rect 2195 -725 2995 30
<< mimcapcontact >>
rect 2205 280 2240 315
rect 2205 30 2240 65
<< metal4 >>
rect 2125 315 2245 320
rect 2125 280 2205 315
rect 2240 280 2245 315
rect 2125 275 2245 280
rect 2125 65 2245 70
rect 2125 30 2205 65
rect 2240 30 2245 65
rect 2125 25 2245 30
<< end >>
