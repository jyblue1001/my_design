magic
tech sky130A
timestamp 1739892886
<< nwell >>
rect 455 105 2380 210
<< nmos >>
rect 515 -35 530 15
rect 740 -35 755 15
rect 795 -35 810 15
rect 920 -35 935 15
rect 975 -35 990 15
rect 1030 -35 1045 15
rect 1085 -35 1100 15
rect 1260 -35 1275 15
rect 1315 -35 1330 15
rect 1370 -35 1385 15
rect 1425 -35 1440 15
rect 1590 -35 1605 15
rect 1645 -35 1660 15
rect 1700 -35 1715 15
rect 1755 -35 1770 15
rect 1925 -35 1940 15
rect 1980 -35 1995 15
rect 2105 -35 2120 15
rect 2160 -35 2175 15
rect 2215 -35 2230 15
rect 2270 -35 2285 15
<< pmos >>
rect 515 125 530 175
rect 570 125 585 175
rect 740 125 755 175
rect 795 125 810 175
rect 1005 125 1020 175
rect 1315 125 1330 175
rect 1370 125 1385 175
rect 1425 125 1440 175
rect 1590 125 1605 175
rect 1645 125 1660 175
rect 1925 125 1940 175
rect 1980 125 1995 175
rect 2190 125 2205 175
<< ndiff >>
rect 475 0 515 15
rect 475 -20 485 0
rect 505 -20 515 0
rect 475 -35 515 -20
rect 530 0 570 15
rect 530 -20 540 0
rect 560 -20 570 0
rect 530 -35 570 -20
rect 700 0 740 15
rect 700 -20 710 0
rect 730 -20 740 0
rect 700 -35 740 -20
rect 755 0 795 15
rect 755 -20 765 0
rect 785 -20 795 0
rect 755 -35 795 -20
rect 810 0 850 15
rect 810 -20 820 0
rect 840 -20 850 0
rect 810 -35 850 -20
rect 880 0 920 15
rect 880 -20 890 0
rect 910 -20 920 0
rect 880 -35 920 -20
rect 935 0 975 15
rect 935 -20 945 0
rect 965 -20 975 0
rect 935 -35 975 -20
rect 990 0 1030 15
rect 990 -20 1000 0
rect 1020 -20 1030 0
rect 990 -35 1030 -20
rect 1045 0 1085 15
rect 1045 -20 1055 0
rect 1075 -20 1085 0
rect 1045 -35 1085 -20
rect 1100 0 1140 15
rect 1100 -20 1110 0
rect 1130 -20 1140 0
rect 1100 -35 1140 -20
rect 1220 0 1260 15
rect 1220 -20 1230 0
rect 1250 -20 1260 0
rect 1220 -35 1260 -20
rect 1275 0 1315 15
rect 1275 -20 1285 0
rect 1305 -20 1315 0
rect 1275 -35 1315 -20
rect 1330 0 1370 15
rect 1330 -20 1340 0
rect 1360 -20 1370 0
rect 1330 -35 1370 -20
rect 1385 0 1425 15
rect 1385 -20 1395 0
rect 1415 -20 1425 0
rect 1385 -35 1425 -20
rect 1440 0 1480 15
rect 1440 -20 1450 0
rect 1470 -20 1480 0
rect 1440 -35 1480 -20
rect 1550 0 1590 15
rect 1550 -20 1560 0
rect 1580 -20 1590 0
rect 1550 -35 1590 -20
rect 1605 0 1645 15
rect 1605 -20 1615 0
rect 1635 -20 1645 0
rect 1605 -35 1645 -20
rect 1660 0 1700 15
rect 1660 -20 1670 0
rect 1690 -20 1700 0
rect 1660 -35 1700 -20
rect 1715 0 1755 15
rect 1715 -20 1725 0
rect 1745 -20 1755 0
rect 1715 -35 1755 -20
rect 1770 0 1810 15
rect 1770 -20 1780 0
rect 1800 -20 1810 0
rect 1770 -35 1810 -20
rect 1885 0 1925 15
rect 1885 -20 1895 0
rect 1915 -20 1925 0
rect 1885 -35 1925 -20
rect 1940 0 1980 15
rect 1940 -20 1950 0
rect 1970 -20 1980 0
rect 1940 -35 1980 -20
rect 1995 0 2035 15
rect 1995 -20 2005 0
rect 2025 -20 2035 0
rect 1995 -35 2035 -20
rect 2065 0 2105 15
rect 2065 -20 2075 0
rect 2095 -20 2105 0
rect 2065 -35 2105 -20
rect 2120 0 2160 15
rect 2120 -20 2130 0
rect 2150 -20 2160 0
rect 2120 -35 2160 -20
rect 2175 0 2215 15
rect 2175 -20 2185 0
rect 2205 -20 2215 0
rect 2175 -35 2215 -20
rect 2230 0 2270 15
rect 2230 -20 2240 0
rect 2260 -20 2270 0
rect 2230 -35 2270 -20
rect 2285 0 2325 15
rect 2285 -20 2295 0
rect 2315 -20 2325 0
rect 2285 -35 2325 -20
<< pdiff >>
rect 475 160 515 175
rect 475 140 485 160
rect 505 140 515 160
rect 475 125 515 140
rect 530 160 570 175
rect 530 140 540 160
rect 560 140 570 160
rect 530 125 570 140
rect 585 160 625 175
rect 585 140 595 160
rect 615 140 625 160
rect 585 125 625 140
rect 700 160 740 175
rect 700 140 710 160
rect 730 140 740 160
rect 700 125 740 140
rect 755 160 795 175
rect 755 140 765 160
rect 785 140 795 160
rect 755 125 795 140
rect 810 160 850 175
rect 810 140 820 160
rect 840 140 850 160
rect 810 125 850 140
rect 965 160 1005 175
rect 965 140 975 160
rect 995 140 1005 160
rect 965 125 1005 140
rect 1020 160 1060 175
rect 1020 140 1030 160
rect 1050 140 1060 160
rect 1020 125 1060 140
rect 1275 160 1315 175
rect 1275 140 1285 160
rect 1305 140 1315 160
rect 1275 125 1315 140
rect 1330 160 1370 175
rect 1330 140 1340 160
rect 1360 140 1370 160
rect 1330 125 1370 140
rect 1385 160 1425 175
rect 1385 140 1395 160
rect 1415 140 1425 160
rect 1385 125 1425 140
rect 1440 160 1480 175
rect 1440 140 1450 160
rect 1470 140 1480 160
rect 1440 125 1480 140
rect 1550 160 1590 175
rect 1550 140 1560 160
rect 1580 140 1590 160
rect 1550 125 1590 140
rect 1605 160 1645 175
rect 1605 140 1615 160
rect 1635 140 1645 160
rect 1605 125 1645 140
rect 1660 160 1700 175
rect 1660 140 1670 160
rect 1690 140 1700 160
rect 1660 125 1700 140
rect 1885 160 1925 175
rect 1885 140 1895 160
rect 1915 140 1925 160
rect 1885 125 1925 140
rect 1940 160 1980 175
rect 1940 140 1950 160
rect 1970 140 1980 160
rect 1940 125 1980 140
rect 1995 160 2035 175
rect 1995 140 2005 160
rect 2025 140 2035 160
rect 1995 125 2035 140
rect 2150 160 2190 175
rect 2150 140 2160 160
rect 2180 140 2190 160
rect 2150 125 2190 140
rect 2205 160 2245 175
rect 2205 140 2215 160
rect 2235 140 2245 160
rect 2205 125 2245 140
<< ndiffc >>
rect 485 -20 505 0
rect 540 -20 560 0
rect 710 -20 730 0
rect 765 -20 785 0
rect 820 -20 840 0
rect 890 -20 910 0
rect 945 -20 965 0
rect 1000 -20 1020 0
rect 1055 -20 1075 0
rect 1110 -20 1130 0
rect 1230 -20 1250 0
rect 1285 -20 1305 0
rect 1340 -20 1360 0
rect 1395 -20 1415 0
rect 1450 -20 1470 0
rect 1560 -20 1580 0
rect 1615 -20 1635 0
rect 1670 -20 1690 0
rect 1725 -20 1745 0
rect 1780 -20 1800 0
rect 1895 -20 1915 0
rect 1950 -20 1970 0
rect 2005 -20 2025 0
rect 2075 -20 2095 0
rect 2130 -20 2150 0
rect 2185 -20 2205 0
rect 2240 -20 2260 0
rect 2295 -20 2315 0
<< pdiffc >>
rect 485 140 505 160
rect 540 140 560 160
rect 595 140 615 160
rect 710 140 730 160
rect 765 140 785 160
rect 820 140 840 160
rect 975 140 995 160
rect 1030 140 1050 160
rect 1285 140 1305 160
rect 1340 140 1360 160
rect 1395 140 1415 160
rect 1450 140 1470 160
rect 1560 140 1580 160
rect 1615 140 1635 160
rect 1670 140 1690 160
rect 1895 140 1915 160
rect 1950 140 1970 160
rect 2005 140 2025 160
rect 2160 140 2180 160
rect 2215 140 2235 160
<< psubdiff >>
rect 660 0 700 15
rect 660 -20 670 0
rect 690 -20 700 0
rect 660 -35 700 -20
<< nsubdiff >>
rect 925 160 965 175
rect 925 140 935 160
rect 955 140 965 160
rect 925 125 965 140
rect 2110 160 2150 175
rect 2110 140 2120 160
rect 2140 140 2150 160
rect 2110 125 2150 140
<< psubdiffcont >>
rect 670 -20 690 0
<< nsubdiffcont >>
rect 935 140 955 160
rect 2120 140 2140 160
<< poly >>
rect 795 220 840 230
rect 795 200 810 220
rect 830 200 840 220
rect 795 190 840 200
rect 1370 220 1400 230
rect 1370 200 1375 220
rect 1395 200 1400 220
rect 1370 190 1400 200
rect 1425 220 1470 230
rect 1980 220 2030 230
rect 1425 200 1440 220
rect 1460 200 1470 220
rect 1425 190 1470 200
rect 1835 210 1875 220
rect 1835 190 1845 210
rect 1865 190 1875 210
rect 1980 200 2000 220
rect 2020 200 2030 220
rect 1980 190 2030 200
rect 515 175 530 190
rect 570 175 585 190
rect 740 175 755 190
rect 795 175 810 190
rect 1005 175 1020 190
rect 1315 175 1330 190
rect 1370 175 1385 190
rect 1425 175 1440 190
rect 1590 175 1605 190
rect 1645 175 1660 190
rect 1835 180 1875 190
rect 515 115 530 125
rect 570 115 585 125
rect 515 100 585 115
rect 645 120 685 130
rect 645 100 655 120
rect 675 105 685 120
rect 740 105 755 125
rect 795 110 810 125
rect 675 100 755 105
rect 515 15 530 100
rect 645 90 755 100
rect 555 60 595 70
rect 675 60 715 65
rect 555 40 565 60
rect 585 45 685 60
rect 585 40 595 45
rect 555 30 595 40
rect 675 40 685 45
rect 705 40 715 60
rect 675 30 715 40
rect 740 15 755 90
rect 1005 105 1020 125
rect 1005 90 1185 105
rect 780 60 820 70
rect 780 40 790 60
rect 810 40 820 60
rect 1005 40 1020 90
rect 1070 60 1110 65
rect 1070 40 1080 60
rect 1100 40 1110 60
rect 780 30 1045 40
rect 1070 30 1110 40
rect 1170 45 1185 90
rect 1245 60 1285 65
rect 1245 45 1255 60
rect 1170 40 1255 45
rect 1275 40 1285 60
rect 1170 30 1285 40
rect 795 25 1045 30
rect 795 15 810 25
rect 920 15 935 25
rect 975 15 990 25
rect 1030 15 1045 25
rect 1085 15 1100 30
rect 1260 15 1275 30
rect 1315 15 1330 125
rect 1370 15 1385 125
rect 1425 15 1440 125
rect 1495 120 1535 130
rect 1495 100 1505 120
rect 1525 110 1535 120
rect 1590 110 1605 125
rect 1525 100 1605 110
rect 1495 95 1605 100
rect 1495 90 1535 95
rect 1505 60 1545 65
rect 1505 40 1515 60
rect 1535 45 1545 60
rect 1645 45 1660 125
rect 1695 100 1735 110
rect 1695 80 1705 100
rect 1725 85 1735 100
rect 1860 95 1875 180
rect 1925 175 1940 190
rect 1980 175 1995 190
rect 2190 175 2205 190
rect 2320 160 2360 170
rect 2320 140 2330 160
rect 2350 140 2360 160
rect 2320 130 2360 140
rect 1925 95 1940 125
rect 1980 110 1995 125
rect 1725 80 1770 85
rect 1695 70 1770 80
rect 1860 80 1940 95
rect 1535 40 1715 45
rect 1505 30 1715 40
rect 1590 15 1605 30
rect 1645 15 1660 30
rect 1700 15 1715 30
rect 1755 15 1770 70
rect 1795 60 1835 70
rect 1795 40 1805 60
rect 1825 40 1835 60
rect 1795 30 1835 40
rect 515 -50 530 -35
rect 740 -50 755 -35
rect 795 -50 810 -35
rect 920 -50 935 -35
rect 975 -50 990 -35
rect 1030 -50 1045 -35
rect 1085 -50 1100 -35
rect 1260 -50 1275 -35
rect 1315 -50 1330 -35
rect 1370 -50 1385 -35
rect 1425 -50 1440 -35
rect 1590 -50 1605 -35
rect 1645 -50 1660 -35
rect 1700 -50 1715 -35
rect 1755 -50 1770 -35
rect 1860 -40 1875 80
rect 1925 15 1940 80
rect 1965 60 2005 70
rect 1965 40 1975 60
rect 1995 40 2005 60
rect 2190 40 2205 125
rect 2255 60 2295 70
rect 2255 40 2265 60
rect 2285 40 2295 60
rect 1965 30 2230 40
rect 2255 30 2295 40
rect 1980 25 2230 30
rect 1980 15 1995 25
rect 2105 15 2120 25
rect 2160 15 2175 25
rect 2215 15 2230 25
rect 2270 15 2285 30
rect 1835 -50 1875 -40
rect 1925 -50 1940 -35
rect 1980 -50 1995 -35
rect 2105 -50 2120 -35
rect 2160 -50 2175 -35
rect 2215 -50 2230 -35
rect 2270 -50 2285 -35
rect 515 -55 560 -50
rect 515 -75 530 -55
rect 550 -75 560 -55
rect 515 -85 560 -75
rect 1300 -55 1340 -50
rect 1300 -75 1310 -55
rect 1330 -75 1340 -55
rect 1300 -85 1340 -75
rect 1835 -70 1845 -50
rect 1865 -70 1875 -50
rect 1835 -80 1875 -70
rect 2310 -60 2350 -50
rect 2310 -80 2320 -60
rect 2340 -80 2350 -60
rect 2310 -90 2350 -80
<< polycont >>
rect 810 200 830 220
rect 1375 200 1395 220
rect 1440 200 1460 220
rect 1845 190 1865 210
rect 2000 200 2020 220
rect 655 100 675 120
rect 565 40 585 60
rect 685 40 705 60
rect 790 40 810 60
rect 1080 40 1100 60
rect 1255 40 1275 60
rect 1505 100 1525 120
rect 1515 40 1535 60
rect 1705 80 1725 100
rect 2330 140 2350 160
rect 1805 40 1825 60
rect 1975 40 1995 60
rect 2265 40 2285 60
rect 530 -75 550 -55
rect 1310 -75 1330 -55
rect 1845 -70 1865 -50
rect 2320 -80 2340 -60
<< locali >>
rect 455 255 485 275
rect 505 255 535 275
rect 555 255 585 275
rect 605 255 635 275
rect 655 255 685 275
rect 705 255 735 275
rect 755 255 785 275
rect 805 255 835 275
rect 855 255 885 275
rect 905 255 935 275
rect 955 255 985 275
rect 1005 255 1035 275
rect 1055 255 1085 275
rect 1105 255 1135 275
rect 1155 255 1185 275
rect 1205 255 1235 275
rect 1255 255 1285 275
rect 1305 255 1335 275
rect 1355 255 1385 275
rect 1405 255 1435 275
rect 1455 255 1485 275
rect 1505 255 1535 275
rect 1555 255 1585 275
rect 1605 255 1635 275
rect 1655 255 1685 275
rect 1705 255 1735 275
rect 1755 255 1785 275
rect 1805 255 1835 275
rect 1855 255 1885 275
rect 1905 255 1935 275
rect 1955 255 1985 275
rect 2005 255 2035 275
rect 2055 255 2085 275
rect 2105 255 2135 275
rect 2155 255 2185 275
rect 2205 255 2235 275
rect 2255 255 2285 275
rect 2305 255 2335 275
rect 2355 255 2380 275
rect 540 170 560 255
rect 690 220 730 230
rect 690 200 700 220
rect 720 200 730 220
rect 690 190 730 200
rect 710 170 730 190
rect 760 170 780 255
rect 800 220 840 230
rect 800 200 810 220
rect 830 200 840 220
rect 800 190 840 200
rect 975 170 995 255
rect 1330 170 1350 255
rect 1370 220 1400 230
rect 1370 200 1375 220
rect 1395 200 1400 220
rect 1370 190 1400 200
rect 1430 220 1470 230
rect 1430 200 1440 220
rect 1460 200 1470 220
rect 1430 190 1470 200
rect 1615 170 1635 255
rect 1895 220 1930 230
rect 1835 210 1875 220
rect 1835 190 1845 210
rect 1865 190 1875 210
rect 1835 180 1875 190
rect 1895 200 1905 220
rect 1925 200 1930 220
rect 1895 190 1930 200
rect 1895 170 1915 190
rect 1950 170 1970 255
rect 1990 220 2030 230
rect 1990 200 2000 220
rect 2020 200 2030 220
rect 1990 190 2030 200
rect 2160 170 2180 255
rect 480 160 510 170
rect 480 140 485 160
rect 505 140 510 160
rect 480 130 510 140
rect 535 160 565 170
rect 535 140 540 160
rect 560 140 565 160
rect 535 130 565 140
rect 590 160 620 170
rect 590 140 595 160
rect 615 140 620 160
rect 590 130 620 140
rect 705 160 735 170
rect 705 140 710 160
rect 730 140 735 160
rect 705 130 735 140
rect 760 160 790 170
rect 760 140 765 160
rect 785 140 790 160
rect 760 130 790 140
rect 815 160 845 170
rect 930 160 1000 170
rect 815 140 820 160
rect 840 140 910 160
rect 815 130 845 140
rect 485 110 505 130
rect 595 110 615 130
rect 645 120 685 130
rect 645 110 655 120
rect 485 100 655 110
rect 675 100 685 120
rect 485 90 685 100
rect 710 110 730 130
rect 710 90 865 110
rect 455 60 595 70
rect 455 50 565 60
rect 555 40 565 50
rect 585 40 595 60
rect 555 30 595 40
rect 480 0 510 10
rect 480 -20 485 0
rect 505 -20 510 0
rect 480 -30 510 -20
rect 535 0 565 10
rect 625 0 645 90
rect 675 60 715 65
rect 780 60 820 70
rect 675 40 685 60
rect 705 40 790 60
rect 810 40 820 60
rect 675 30 715 40
rect 780 30 820 40
rect 845 10 865 90
rect 890 50 910 140
rect 930 140 935 160
rect 955 140 975 160
rect 995 140 1000 160
rect 930 130 1000 140
rect 1025 160 1055 170
rect 1135 160 1175 170
rect 1025 140 1030 160
rect 1050 140 1145 160
rect 1165 140 1175 160
rect 1025 130 1055 140
rect 1135 130 1175 140
rect 1280 160 1310 170
rect 1280 140 1285 160
rect 1305 140 1310 160
rect 1280 130 1310 140
rect 1330 160 1365 170
rect 1330 140 1340 160
rect 1360 140 1365 160
rect 1330 130 1365 140
rect 1390 160 1420 170
rect 1390 140 1395 160
rect 1415 140 1420 160
rect 1390 130 1420 140
rect 1445 160 1475 170
rect 1445 140 1450 160
rect 1470 140 1475 160
rect 1445 130 1475 140
rect 1555 160 1585 170
rect 1555 140 1560 160
rect 1580 140 1585 160
rect 1555 130 1585 140
rect 1610 160 1640 170
rect 1610 140 1615 160
rect 1635 140 1640 160
rect 1610 130 1640 140
rect 1665 160 1695 170
rect 1890 160 1920 170
rect 1665 140 1670 160
rect 1690 140 1805 160
rect 1665 130 1695 140
rect 1070 60 1110 65
rect 1070 50 1080 60
rect 890 40 1080 50
rect 1100 40 1110 60
rect 890 30 1110 40
rect 890 10 910 30
rect 1000 10 1020 30
rect 1135 10 1155 130
rect 1285 110 1305 130
rect 1450 110 1470 130
rect 1495 120 1535 130
rect 1495 110 1505 120
rect 535 -20 540 0
rect 560 -20 645 0
rect 665 0 735 10
rect 665 -20 670 0
rect 690 -20 710 0
rect 730 -20 735 0
rect 535 -30 565 -20
rect 665 -30 735 -20
rect 760 0 790 10
rect 760 -20 765 0
rect 785 -20 790 0
rect 760 -30 790 -20
rect 815 0 865 10
rect 815 -20 820 0
rect 840 -20 865 0
rect 885 0 915 10
rect 885 -20 890 0
rect 910 -20 915 0
rect 815 -30 845 -20
rect 885 -30 915 -20
rect 940 0 970 10
rect 940 -20 945 0
rect 965 -20 970 0
rect 940 -30 970 -20
rect 995 0 1025 10
rect 995 -20 1000 0
rect 1020 -20 1025 0
rect 995 -30 1025 -20
rect 1050 0 1080 10
rect 1050 -20 1055 0
rect 1075 -20 1080 0
rect 1050 -30 1080 -20
rect 1105 0 1155 10
rect 1105 -20 1110 0
rect 1130 -20 1155 0
rect 1205 100 1505 110
rect 1525 100 1535 120
rect 1205 90 1535 100
rect 1205 10 1225 90
rect 1245 60 1285 65
rect 1245 40 1255 60
rect 1275 40 1285 60
rect 1505 60 1545 65
rect 1245 30 1285 40
rect 1340 30 1470 50
rect 1505 40 1515 60
rect 1535 40 1545 60
rect 1505 30 1545 40
rect 1565 50 1585 130
rect 1695 100 1735 110
rect 1695 80 1705 100
rect 1725 80 1735 100
rect 1695 70 1735 80
rect 1785 70 1805 140
rect 1890 140 1895 160
rect 1915 140 1920 160
rect 1890 130 1920 140
rect 1945 160 1975 170
rect 1945 140 1950 160
rect 1970 140 1975 160
rect 1945 130 1975 140
rect 2000 160 2030 170
rect 2115 160 2185 170
rect 2000 140 2005 160
rect 2025 140 2095 160
rect 2000 130 2030 140
rect 1895 110 1915 130
rect 1895 90 2050 110
rect 1695 50 1715 70
rect 1565 30 1715 50
rect 1785 60 1835 70
rect 1965 60 2005 70
rect 1785 40 1805 60
rect 1825 40 1975 60
rect 1995 40 2005 60
rect 1785 30 1835 40
rect 1965 30 2005 40
rect 1340 10 1360 30
rect 1450 10 1470 30
rect 1565 10 1585 30
rect 1675 10 1695 30
rect 1785 10 1805 30
rect 2030 10 2050 90
rect 2075 50 2095 140
rect 2115 140 2120 160
rect 2140 140 2160 160
rect 2180 140 2185 160
rect 2115 130 2185 140
rect 2210 160 2240 170
rect 2320 160 2360 170
rect 2210 140 2215 160
rect 2235 140 2330 160
rect 2350 140 2360 160
rect 2210 130 2240 140
rect 2320 130 2360 140
rect 2320 85 2340 130
rect 2255 60 2295 70
rect 2255 50 2265 60
rect 2075 40 2265 50
rect 2285 40 2295 60
rect 2075 30 2295 40
rect 2320 65 2380 85
rect 2075 10 2095 30
rect 2185 10 2205 30
rect 2320 10 2340 65
rect 1205 0 1255 10
rect 1205 -20 1230 0
rect 1250 -20 1255 0
rect 1105 -30 1135 -20
rect 1225 -30 1255 -20
rect 1280 0 1310 10
rect 1280 -20 1285 0
rect 1305 -20 1310 0
rect 1280 -30 1310 -20
rect 1335 0 1365 10
rect 1335 -20 1340 0
rect 1360 -20 1365 0
rect 1335 -30 1365 -20
rect 1390 0 1420 10
rect 1390 -20 1395 0
rect 1415 -20 1420 0
rect 1390 -30 1420 -20
rect 1445 0 1475 10
rect 1445 -20 1450 0
rect 1470 -20 1475 0
rect 1445 -30 1475 -20
rect 1555 0 1585 10
rect 1555 -20 1560 0
rect 1580 -20 1585 0
rect 1555 -30 1585 -20
rect 1610 0 1640 10
rect 1610 -20 1615 0
rect 1635 -20 1640 0
rect 1610 -30 1640 -20
rect 1665 0 1695 10
rect 1665 -20 1670 0
rect 1690 -20 1695 0
rect 1665 -30 1695 -20
rect 1720 0 1750 10
rect 1720 -20 1725 0
rect 1745 -20 1750 0
rect 1720 -30 1750 -20
rect 1775 0 1805 10
rect 1775 -20 1780 0
rect 1800 -20 1805 0
rect 1775 -30 1805 -20
rect 1890 0 1920 10
rect 1890 -20 1895 0
rect 1915 -20 1920 0
rect 1890 -30 1920 -20
rect 1945 0 1975 10
rect 1945 -20 1950 0
rect 1970 -20 1975 0
rect 1945 -30 1975 -20
rect 2000 0 2050 10
rect 2000 -20 2005 0
rect 2025 -20 2050 0
rect 2070 0 2100 10
rect 2070 -20 2075 0
rect 2095 -20 2100 0
rect 2000 -30 2030 -20
rect 2070 -30 2100 -20
rect 2125 0 2155 10
rect 2125 -20 2130 0
rect 2150 -20 2155 0
rect 2125 -30 2155 -20
rect 2180 0 2210 10
rect 2180 -20 2185 0
rect 2205 -20 2210 0
rect 2180 -30 2210 -20
rect 2235 0 2265 10
rect 2235 -20 2240 0
rect 2260 -20 2265 0
rect 2235 -30 2265 -20
rect 2290 0 2340 10
rect 2290 -20 2295 0
rect 2315 -20 2340 0
rect 2290 -30 2340 -20
rect 480 -115 500 -30
rect 520 -55 560 -50
rect 520 -75 530 -55
rect 550 -75 560 -55
rect 520 -85 560 -75
rect 710 -115 730 -30
rect 945 -115 965 -30
rect 1055 -115 1075 -30
rect 1300 -55 1340 -50
rect 1300 -75 1310 -55
rect 1330 -75 1340 -55
rect 1300 -85 1340 -75
rect 1395 -115 1415 -30
rect 1615 -115 1635 -30
rect 1725 -115 1745 -30
rect 1780 -50 1800 -30
rect 1835 -50 1875 -40
rect 1770 -55 1810 -50
rect 1770 -75 1780 -55
rect 1800 -75 1810 -55
rect 1770 -85 1810 -75
rect 1835 -70 1845 -50
rect 1865 -70 1875 -50
rect 1835 -80 1875 -70
rect 1895 -115 1915 -30
rect 2130 -115 2150 -30
rect 2240 -115 2260 -30
rect 2320 -50 2340 -30
rect 2310 -60 2350 -50
rect 2310 -80 2320 -60
rect 2340 -80 2350 -60
rect 2310 -90 2350 -80
rect 455 -135 485 -115
rect 505 -135 535 -115
rect 555 -135 585 -115
rect 605 -135 635 -115
rect 655 -135 685 -115
rect 705 -135 735 -115
rect 755 -135 785 -115
rect 805 -135 835 -115
rect 855 -135 885 -115
rect 905 -135 935 -115
rect 955 -135 985 -115
rect 1005 -135 1035 -115
rect 1055 -135 1085 -115
rect 1105 -135 1135 -115
rect 1155 -135 1185 -115
rect 1205 -135 1235 -115
rect 1255 -135 1285 -115
rect 1305 -135 1335 -115
rect 1355 -135 1385 -115
rect 1405 -135 1435 -115
rect 1455 -135 1485 -115
rect 1505 -135 1535 -115
rect 1555 -135 1585 -115
rect 1605 -135 1635 -115
rect 1655 -135 1685 -115
rect 1705 -135 1735 -115
rect 1755 -135 1785 -115
rect 1805 -135 1835 -115
rect 1855 -135 1885 -115
rect 1905 -135 1935 -115
rect 1955 -135 1985 -115
rect 2005 -135 2035 -115
rect 2055 -135 2085 -115
rect 2105 -135 2135 -115
rect 2155 -135 2185 -115
rect 2205 -135 2235 -115
rect 2255 -135 2285 -115
rect 2305 -135 2335 -115
rect 2355 -135 2380 -115
<< viali >>
rect 485 255 505 275
rect 535 255 555 275
rect 585 255 605 275
rect 635 255 655 275
rect 685 255 705 275
rect 735 255 755 275
rect 785 255 805 275
rect 835 255 855 275
rect 885 255 905 275
rect 935 255 955 275
rect 985 255 1005 275
rect 1035 255 1055 275
rect 1085 255 1105 275
rect 1135 255 1155 275
rect 1185 255 1205 275
rect 1235 255 1255 275
rect 1285 255 1305 275
rect 1335 255 1355 275
rect 1385 255 1405 275
rect 1435 255 1455 275
rect 1485 255 1505 275
rect 1535 255 1555 275
rect 1585 255 1605 275
rect 1635 255 1655 275
rect 1685 255 1705 275
rect 1735 255 1755 275
rect 1785 255 1805 275
rect 1835 255 1855 275
rect 1885 255 1905 275
rect 1935 255 1955 275
rect 1985 255 2005 275
rect 2035 255 2055 275
rect 2085 255 2105 275
rect 2135 255 2155 275
rect 2185 255 2205 275
rect 2235 255 2255 275
rect 2285 255 2305 275
rect 2335 255 2355 275
rect 700 200 720 220
rect 810 200 830 220
rect 1375 200 1395 220
rect 1440 200 1460 220
rect 1845 190 1865 210
rect 1905 200 1925 220
rect 2000 200 2020 220
rect 1145 140 1165 160
rect 1255 40 1275 60
rect 1515 40 1535 60
rect 530 -75 550 -55
rect 1310 -75 1330 -55
rect 1780 -75 1800 -55
rect 1845 -70 1865 -50
rect 2320 -80 2340 -60
rect 485 -135 505 -115
rect 535 -135 555 -115
rect 585 -135 605 -115
rect 635 -135 655 -115
rect 685 -135 705 -115
rect 735 -135 755 -115
rect 785 -135 805 -115
rect 835 -135 855 -115
rect 885 -135 905 -115
rect 935 -135 955 -115
rect 985 -135 1005 -115
rect 1035 -135 1055 -115
rect 1085 -135 1105 -115
rect 1135 -135 1155 -115
rect 1185 -135 1205 -115
rect 1235 -135 1255 -115
rect 1285 -135 1305 -115
rect 1335 -135 1355 -115
rect 1385 -135 1405 -115
rect 1435 -135 1455 -115
rect 1485 -135 1505 -115
rect 1535 -135 1555 -115
rect 1585 -135 1605 -115
rect 1635 -135 1655 -115
rect 1685 -135 1705 -115
rect 1735 -135 1755 -115
rect 1785 -135 1805 -115
rect 1835 -135 1855 -115
rect 1885 -135 1905 -115
rect 1935 -135 1955 -115
rect 1985 -135 2005 -115
rect 2035 -135 2055 -115
rect 2085 -135 2105 -115
rect 2135 -135 2155 -115
rect 2185 -135 2205 -115
rect 2235 -135 2255 -115
rect 2285 -135 2305 -115
rect 2335 -135 2355 -115
<< metal1 >>
rect 455 275 2380 285
rect 455 255 485 275
rect 505 255 535 275
rect 555 255 585 275
rect 605 255 635 275
rect 655 255 685 275
rect 705 255 735 275
rect 755 255 785 275
rect 805 255 835 275
rect 855 255 885 275
rect 905 255 935 275
rect 955 255 985 275
rect 1005 255 1035 275
rect 1055 255 1085 275
rect 1105 255 1135 275
rect 1155 255 1185 275
rect 1205 255 1235 275
rect 1255 255 1285 275
rect 1305 255 1335 275
rect 1355 255 1385 275
rect 1405 255 1435 275
rect 1455 255 1485 275
rect 1505 255 1535 275
rect 1555 255 1585 275
rect 1605 255 1635 275
rect 1655 255 1685 275
rect 1705 255 1735 275
rect 1755 255 1785 275
rect 1805 255 1835 275
rect 1855 255 1885 275
rect 1905 255 1935 275
rect 1955 255 1985 275
rect 2005 255 2035 275
rect 2055 255 2085 275
rect 2105 255 2135 275
rect 2155 255 2185 275
rect 2205 255 2235 275
rect 2255 255 2285 275
rect 2305 255 2335 275
rect 2355 255 2380 275
rect 455 245 2380 255
rect 690 220 730 230
rect 690 200 700 220
rect 720 210 730 220
rect 800 220 840 230
rect 800 210 810 220
rect 720 200 810 210
rect 830 200 840 220
rect 1370 220 1400 230
rect 1370 210 1375 220
rect 690 190 840 200
rect 1155 200 1375 210
rect 1395 200 1400 220
rect 1155 190 1400 200
rect 1430 220 1470 230
rect 1895 220 1930 230
rect 1430 200 1440 220
rect 1460 210 1470 220
rect 1835 210 1875 220
rect 1460 200 1845 210
rect 1430 190 1845 200
rect 1865 190 1875 210
rect 1895 200 1905 220
rect 1925 210 1930 220
rect 1990 220 2030 230
rect 1990 210 2000 220
rect 1925 200 2000 210
rect 2020 200 2030 220
rect 1895 190 2030 200
rect 1155 170 1175 190
rect 1835 180 1875 190
rect 1135 160 1175 170
rect 1135 140 1145 160
rect 1165 140 1175 160
rect 1135 130 1175 140
rect 1245 60 1545 65
rect 1245 40 1255 60
rect 1275 45 1515 60
rect 1275 40 1285 45
rect 1245 30 1285 40
rect 1505 40 1515 45
rect 1535 40 1545 60
rect 1505 30 1545 40
rect 1835 -50 1875 -40
rect 520 -55 560 -50
rect 520 -75 530 -55
rect 550 -65 560 -55
rect 1300 -55 1340 -50
rect 1300 -65 1310 -55
rect 550 -75 1310 -65
rect 1330 -65 1340 -55
rect 1770 -55 1810 -50
rect 1770 -65 1780 -55
rect 1330 -75 1780 -65
rect 1800 -75 1810 -55
rect 520 -85 1810 -75
rect 1835 -70 1845 -50
rect 1865 -60 1875 -50
rect 2310 -60 2350 -50
rect 1865 -70 2320 -60
rect 1835 -80 2320 -70
rect 2340 -80 2350 -60
rect 2310 -90 2350 -80
rect 455 -115 2380 -105
rect 455 -135 485 -115
rect 505 -135 535 -115
rect 555 -135 585 -115
rect 605 -135 635 -115
rect 655 -135 685 -115
rect 705 -135 735 -115
rect 755 -135 785 -115
rect 805 -135 835 -115
rect 855 -135 885 -115
rect 905 -135 935 -115
rect 955 -135 985 -115
rect 1005 -135 1035 -115
rect 1055 -135 1085 -115
rect 1105 -135 1135 -115
rect 1155 -135 1185 -115
rect 1205 -135 1235 -115
rect 1255 -135 1285 -115
rect 1305 -135 1335 -115
rect 1355 -135 1385 -115
rect 1405 -135 1435 -115
rect 1455 -135 1485 -115
rect 1505 -135 1535 -115
rect 1555 -135 1585 -115
rect 1605 -135 1635 -115
rect 1655 -135 1685 -115
rect 1705 -135 1735 -115
rect 1755 -135 1785 -115
rect 1805 -135 1835 -115
rect 1855 -135 1885 -115
rect 1905 -135 1935 -115
rect 1955 -135 1985 -115
rect 2005 -135 2035 -115
rect 2055 -135 2085 -115
rect 2105 -135 2135 -115
rect 2155 -135 2185 -115
rect 2205 -135 2235 -115
rect 2255 -135 2285 -115
rect 2305 -135 2335 -115
rect 2355 -135 2380 -115
rect 455 -145 2380 -135
<< labels >>
flabel locali 775 -30 775 -30 5 FreeSans 160 0 0 -80 C
flabel locali 845 80 845 80 7 FreeSans 160 0 -80 0 B
flabel locali 910 80 910 80 3 FreeSans 160 0 80 0 D
flabel locali 1175 150 1175 150 3 FreeSans 160 0 80 0 E
flabel locali 1405 170 1405 170 1 FreeSans 160 0 0 80 F
flabel locali 1475 150 1475 150 3 FreeSans 160 0 80 0 G
flabel locali 1295 -30 1295 -30 5 FreeSans 160 0 0 -80 H
flabel locali 1585 70 1585 70 3 FreeSans 160 0 80 0 J
flabel locali 1755 160 1755 160 1 FreeSans 160 0 0 80 Q2_b
flabel locali 1960 -30 1960 -30 5 FreeSans 160 0 0 -80 L
flabel locali 2050 70 2050 70 3 FreeSans 160 0 80 0 K
flabel locali 2095 85 2095 85 3 FreeSans 160 0 80 0 M
flabel locali 2380 75 2380 75 3 FreeSans 160 0 80 0 VOUT
port 1 e
flabel locali 455 60 455 60 7 FreeSans 160 0 -80 0 VIN
port 2 w
flabel locali 625 -20 625 -20 5 FreeSans 160 0 0 -80 A
flabel locali 1470 25 1470 25 3 FreeSans 160 0 80 0 I
flabel metal1 455 265 455 265 7 FreeSans 160 0 -80 0 VDDA
port 3 w
flabel metal1 455 -125 455 -125 7 FreeSans 160 0 -80 0 GNDA
port 4 w
<< end >>
