* PEX produced on Mon Feb 17 06:40:05 AM CET 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from pfd_8.ext - technology: sky130A

.subckt pfd_cp_input_magic DOWN_input VDDA GNDA UP_input opamp_out F_REF I_IN F_VCO UP_b DOWN
X0 GNDA.t43 E.t3 QA.t2 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X1 a_4210_n7910.t1 before_Reset.t3 GNDA.t58 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X2 UP_PFD_b.t1 QA.t3 GNDA.t48 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X3 F.t0 QB_b.t3 GNDA.t17 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X4 GNDA.t46 QA.t4 QA_b.t1 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X5 GNDA.t11 Reset.t2 E_b.t0 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X6 DOWN_input.t2 DOWN.t2 I_IN.t1 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X7 VDDA.t29 E.t4 a_2350_n7910.t1 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X8 a_4210_n7910.t0 before_Reset.t4 VDDA.t34 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X9 UP_PFD_b.t0 QA.t5 VDDA.t32 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X10 GNDA.t34 E_b.t3 E.t2 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X11 before_Reset.t1 QA.t6 a_3770_n7290.t1 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X12 VDDA.t21 F.t3 a_2350_n8670.t1 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X13 GNDA.t19 a_4060_n9120.t2 a_3730_n9120.t0 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X14 GNDA.t21 a_4390_n9120.t2 a_4060_n9120.t0 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X15 QA_b.t0 QA.t7 a_1830_n7910.t0 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X16 VDDA.t25 Reset.t3 a_3250_n7910.t0 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X17 DOWN_PFD_b.t1 QB.t3 VDDA.t9 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X18 QB_b.t0 QB.t4 a_1830_n8670.t0 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X19 DOWN.t0 DOWN_b.t2 GNDA.t28 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X20 E.t1 E_b.t4 a_2730_n7910.t1 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X21 VDDA.t31 QA.t8 before_Reset.t2 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X22 VDDA.t24 Reset.t4 a_3250_n8670.t1 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X23 F.t2 F_b.t3 a_2730_n8670.t1 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X24 GNDA.t7 a_3730_n9120.t2 Reset.t1 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X25 QA.t1 QA_b.t3 GNDA.t15 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X26 DOWN_b.t1 VDDA.t41 DOWN_PFD_b.t3 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X27 a_4390_n9120.t0 a_4210_n7910.t2 GNDA.t30 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X28 QA_b.t2 F_REF.t0 GNDA.t56 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X29 E_b.t2 E.t5 GNDA.t41 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X30 E.t0 QA_b.t4 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X31 a_3770_n7290.t0 QB.t5 GNDA.t23 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X32 a_2350_n7910.t0 QA_b.t5 QA.t0 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X33 a_4390_n9120.t1 a_4210_n7910.t3 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X34 a_1830_n7910.t1 F_REF.t1 VDDA.t38 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X35 a_2350_n8670.t0 QB_b.t4 QB.t0 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X36 UP_input.t0 UP.t2 opamp_out.t0 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X37 a_3250_n7910.t1 E.t6 E_b.t1 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X38 UP_input.t1 UP.t3 VDDA.t37 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X39 a_2730_n7910.t0 QA_b.t6 VDDA.t22 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X40 a_1830_n8670.t1 F_VCO.t0 VDDA.t15 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X41 a_3250_n8670.t0 F.t4 F_b.t0 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X42 GNDA.t3 F.t5 QB.t2 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X43 before_Reset.t0 QB.t6 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X44 DOWN_PFD_b.t0 QB.t7 GNDA.t9 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X45 UP_input.t2 UP_b.t2 opamp_out.t1 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X46 a_2730_n8670.t0 QB_b.t5 VDDA.t17 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X47 GNDA.t32 QB.t8 QB_b.t1 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X48 GNDA.t39 Reset.t5 F_b.t2 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X49 UP_b.t0 UP.t4 GNDA.t54 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X50 DOWN_input.t0 DOWN_b.t3 I_IN.t0 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X51 GNDA.t52 F_b.t4 F.t1 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X52 VDDA.t4 a_4060_n9120.t3 a_3730_n9120.t1 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X53 VDDA.t7 a_4390_n9120.t3 a_4060_n9120.t1 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X54 UP_b.t1 UP.t5 VDDA.t35 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X55 UP.t0 UP_PFD_b.t2 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X56 DOWN.t1 DOWN_b.t4 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X57 VDDA.t1 a_3730_n9120.t3 Reset.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X58 UP.t1 UP_PFD_b.t3 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X59 QB.t1 QB_b.t6 GNDA.t13 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X60 DOWN_b.t0 GNDA.t60 DOWN_PFD_b.t2 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X61 QB_b.t2 F_VCO.t1 GNDA.t50 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X62 F_b.t1 F.t6 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X63 DOWN_input.t1 DOWN_b.t5 GNDA.t26 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
R0 E.n4 E.n0 1319.38
R1 E.n0 E.t6 562.333
R2 E.n2 E.t4 388.813
R3 E.n2 E.t3 356.68
R4 E.n3 E.n2 232
R5 E.n0 E.t5 224.934
R6 E.t1 E.n4 221.411
R7 E.n3 E.n1 157.278
R8 E.n4 E.n3 90.64
R9 E.n1 E.t2 24.0005
R10 E.n1 E.t0 24.0005
R11 QA.t6 QA.t8 835.467
R12 QA.n2 QA.t7 517.347
R13 QA.n0 QA.t5 465.933
R14 QA.n1 QA.n0 454.031
R15 QA.n1 QA.t6 394.267
R16 QA.n0 QA.t3 321.334
R17 QA.n4 QA.n3 244.715
R18 QA.n2 QA.t4 228.148
R19 QA.n4 QA.t0 221.411
R20 QA.n5 QA.n2 216
R21 QA.n5 QA.n4 201.573
R22 QA QA.n5 60.8005
R23 QA QA.n1 56.1505
R24 QA.n3 QA.t2 24.0005
R25 QA.n3 QA.t1 24.0005
R26 GNDA.n155 GNDA.n154 21560
R27 GNDA.t40 GNDA.t33 3006.67
R28 GNDA.t14 GNDA.t45 3006.67
R29 GNDA.t35 GNDA.t51 3006.67
R30 GNDA.t12 GNDA.t31 3006.67
R31 GNDA.t37 GNDA.t8 2860
R32 GNDA.t53 GNDA.t59 2126.67
R33 GNDA.t24 GNDA.t27 2126.67
R34 GNDA.n82 GNDA.t29 2090
R35 GNDA.t6 GNDA.n158 1943.33
R36 GNDA.n161 GNDA.n52 1906.67
R37 GNDA.t4 GNDA.n77 1723.33
R38 GNDA.n83 GNDA.t47 1723.33
R39 GNDA.n30 GNDA.t24 1650
R40 GNDA.n29 GNDA.t37 1650
R41 GNDA.n81 GNDA.t57 1430
R42 GNDA.n79 GNDA.t44 1430
R43 GNDA.t20 GNDA.n160 1430
R44 GNDA.t18 GNDA.n159 1430
R45 GNDA.n30 GNDA.t25 1210
R46 GNDA.t27 GNDA.n29 1210
R47 GNDA.n52 GNDA.t8 1210
R48 GNDA.n77 GNDA.t53 1136.67
R49 GNDA.n83 GNDA.t4 1136.67
R50 GNDA.t47 GNDA.n82 1136.67
R51 GNDA.n120 GNDA.n116 1026.67
R52 GNDA.t29 GNDA.n81 990
R53 GNDA.t57 GNDA.n79 990
R54 GNDA.n116 GNDA.t22 990
R55 GNDA.n120 GNDA.t10 990
R56 GNDA.t0 GNDA.n119 990
R57 GNDA.n119 GNDA.t42 990
R58 GNDA.n154 GNDA.t55 990
R59 GNDA.n161 GNDA.t20 990
R60 GNDA.n160 GNDA.t18 990
R61 GNDA.n159 GNDA.t6 990
R62 GNDA.n158 GNDA.t38 990
R63 GNDA.t16 GNDA.n157 990
R64 GNDA.n157 GNDA.t2 990
R65 GNDA.t49 GNDA.n155 990
R66 GNDA.t44 GNDA.t22 806.668
R67 GNDA.t10 GNDA.t40 806.668
R68 GNDA.t33 GNDA.t0 806.668
R69 GNDA.t42 GNDA.t14 806.668
R70 GNDA.t45 GNDA.t55 806.668
R71 GNDA.t38 GNDA.t35 806.668
R72 GNDA.t51 GNDA.t16 806.668
R73 GNDA.t2 GNDA.t12 806.668
R74 GNDA.t31 GNDA.t49 806.668
R75 GNDA.n157 GNDA.n156 585.003
R76 GNDA.n119 GNDA.n118 585.003
R77 GNDA.n121 GNDA.n120 585.001
R78 GNDA.n116 GNDA.n115 585.001
R79 GNDA.n79 GNDA.n78 585.001
R80 GNDA.n81 GNDA.n80 585.001
R81 GNDA.n77 GNDA.n76 585.001
R82 GNDA.n84 GNDA.n83 585.001
R83 GNDA.n82 GNDA.n73 585.001
R84 GNDA.n154 GNDA.n153 585.001
R85 GNDA.n31 GNDA.n30 585.001
R86 GNDA.n29 GNDA.n28 585.001
R87 GNDA.n52 GNDA.n51 585.001
R88 GNDA.n162 GNDA.n161 585.001
R89 GNDA.n160 GNDA.n19 585.001
R90 GNDA.n159 GNDA.n16 585.001
R91 GNDA.n158 GNDA.n13 585.001
R92 GNDA.n155 GNDA.n2 585.001
R93 GNDA.n38 GNDA.t60 566.966
R94 GNDA.n3 GNDA.t32 198.058
R95 GNDA.n203 GNDA.t13 198.058
R96 GNDA.n191 GNDA.t52 198.058
R97 GNDA.n11 GNDA.t36 198.058
R98 GNDA.n147 GNDA.t46 198.058
R99 GNDA.n55 GNDA.t15 198.058
R100 GNDA.n133 GNDA.t34 198.058
R101 GNDA.n128 GNDA.t41 198.058
R102 GNDA.n7 GNDA.t3 130.713
R103 GNDA.n13 GNDA.t39 130.001
R104 GNDA.n16 GNDA.t7 130.001
R105 GNDA.n19 GNDA.t19 130.001
R106 GNDA.n162 GNDA.t21 130.001
R107 GNDA.n153 GNDA.t56 130.001
R108 GNDA.n121 GNDA.t11 130.001
R109 GNDA.n115 GNDA.t23 130.001
R110 GNDA.n78 GNDA.t58 130.001
R111 GNDA.n80 GNDA.t30 130.001
R112 GNDA.n2 GNDA.t50 130.001
R113 GNDA.n8 GNDA.t17 130.001
R114 GNDA.n117 GNDA.t1 130.001
R115 GNDA.n57 GNDA.t43 130.001
R116 GNDA.n51 GNDA.t9 122.501
R117 GNDA.n28 GNDA.t28 122.501
R118 GNDA.n31 GNDA.t26 122.501
R119 GNDA.n73 GNDA.t48 122.501
R120 GNDA.n84 GNDA.t5 122.501
R121 GNDA.n76 GNDA.t54 122.501
R122 GNDA.n32 GNDA.n31 69.7785
R123 GNDA.n76 GNDA.n75 66.2006
R124 GNDA.n183 GNDA.n13 60.29
R125 GNDA.n176 GNDA.n16 60.29
R126 GNDA.n170 GNDA.n19 60.29
R127 GNDA.n163 GNDA.n162 60.29
R128 GNDA.n153 GNDA.n152 60.29
R129 GNDA.n122 GNDA.n121 60.29
R130 GNDA.n115 GNDA.n114 60.29
R131 GNDA.n78 GNDA.n67 60.29
R132 GNDA.n80 GNDA.n69 60.29
R133 GNDA.n211 GNDA.n2 60.29
R134 GNDA.n92 GNDA.n73 59.5478
R135 GNDA.n85 GNDA.n84 59.5478
R136 GNDA.n51 GNDA.n50 58.9809
R137 GNDA.n33 GNDA.n28 58.9809
R138 GNDA.n196 GNDA.n8 54.4005
R139 GNDA.n198 GNDA.n7 54.4005
R140 GNDA.n139 GNDA.n57 54.4005
R141 GNDA.n117 GNDA.n58 54.4005
R142 GNDA.n85 GNDA.n75 36.2476
R143 GNDA.n152 GNDA.n0 33.0991
R144 GNDA.n212 GNDA.n211 33.0991
R145 GNDA.n86 GNDA.n74 32.0005
R146 GNDA.n90 GNDA.n74 32.0005
R147 GNDA.n91 GNDA.n90 32.0005
R148 GNDA.n93 GNDA.n71 32.0005
R149 GNDA.n97 GNDA.n71 32.0005
R150 GNDA.n98 GNDA.n97 32.0005
R151 GNDA.n99 GNDA.n98 32.0005
R152 GNDA.n103 GNDA.n102 32.0005
R153 GNDA.n104 GNDA.n103 32.0005
R154 GNDA.n108 GNDA.n107 32.0005
R155 GNDA.n109 GNDA.n108 32.0005
R156 GNDA.n109 GNDA.n65 32.0005
R157 GNDA.n113 GNDA.n64 32.0005
R158 GNDA.n123 GNDA.n64 32.0005
R159 GNDA.n127 GNDA.n62 32.0005
R160 GNDA.n128 GNDA.n127 32.0005
R161 GNDA.n129 GNDA.n128 32.0005
R162 GNDA.n129 GNDA.n60 32.0005
R163 GNDA.n133 GNDA.n60 32.0005
R164 GNDA.n134 GNDA.n133 32.0005
R165 GNDA.n135 GNDA.n134 32.0005
R166 GNDA.n141 GNDA.n140 32.0005
R167 GNDA.n141 GNDA.n55 32.0005
R168 GNDA.n145 GNDA.n55 32.0005
R169 GNDA.n146 GNDA.n145 32.0005
R170 GNDA.n147 GNDA.n146 32.0005
R171 GNDA.n147 GNDA.n53 32.0005
R172 GNDA.n151 GNDA.n53 32.0005
R173 GNDA.n34 GNDA.n33 32.0005
R174 GNDA.n35 GNDA.n34 32.0005
R175 GNDA.n35 GNDA.n26 32.0005
R176 GNDA.n40 GNDA.n26 32.0005
R177 GNDA.n41 GNDA.n40 32.0005
R178 GNDA.n42 GNDA.n41 32.0005
R179 GNDA.n42 GNDA.n23 32.0005
R180 GNDA.n49 GNDA.n24 32.0005
R181 GNDA.n45 GNDA.n24 32.0005
R182 GNDA.n45 GNDA.n22 32.0005
R183 GNDA.n164 GNDA.n22 32.0005
R184 GNDA.n168 GNDA.n20 32.0005
R185 GNDA.n169 GNDA.n168 32.0005
R186 GNDA.n171 GNDA.n17 32.0005
R187 GNDA.n175 GNDA.n17 32.0005
R188 GNDA.n178 GNDA.n177 32.0005
R189 GNDA.n178 GNDA.n14 32.0005
R190 GNDA.n182 GNDA.n14 32.0005
R191 GNDA.n185 GNDA.n184 32.0005
R192 GNDA.n185 GNDA.n11 32.0005
R193 GNDA.n189 GNDA.n11 32.0005
R194 GNDA.n190 GNDA.n189 32.0005
R195 GNDA.n191 GNDA.n190 32.0005
R196 GNDA.n191 GNDA.n9 32.0005
R197 GNDA.n195 GNDA.n9 32.0005
R198 GNDA.n199 GNDA.n5 32.0005
R199 GNDA.n203 GNDA.n5 32.0005
R200 GNDA.n204 GNDA.n203 32.0005
R201 GNDA.n205 GNDA.n204 32.0005
R202 GNDA.n205 GNDA.n3 32.0005
R203 GNDA.n209 GNDA.n3 32.0005
R204 GNDA.n210 GNDA.n209 32.0005
R205 GNDA.n102 GNDA.n69 28.8005
R206 GNDA.n92 GNDA.n91 25.6005
R207 GNDA.n114 GNDA.n65 25.6005
R208 GNDA.n123 GNDA.n122 25.6005
R209 GNDA.n138 GNDA.n58 25.6005
R210 GNDA.n139 GNDA.n138 25.6005
R211 GNDA.n50 GNDA.n23 25.6005
R212 GNDA.n163 GNDA.n20 25.6005
R213 GNDA.n176 GNDA.n175 25.6005
R214 GNDA.n183 GNDA.n182 25.6005
R215 GNDA.n197 GNDA.n196 25.6005
R216 GNDA.n198 GNDA.n197 22.4005
R217 GNDA.n107 GNDA.n67 19.2005
R218 GNDA.n170 GNDA.n169 16.0005
R219 GNDA.n171 GNDA.n170 16.0005
R220 GNDA.n104 GNDA.n67 12.8005
R221 GNDA GNDA.n0 12.7806
R222 GNDA GNDA.n212 11.8876
R223 GNDA.n199 GNDA.n198 9.6005
R224 GNDA.n87 GNDA.n86 9.3005
R225 GNDA.n88 GNDA.n74 9.3005
R226 GNDA.n90 GNDA.n89 9.3005
R227 GNDA.n91 GNDA.n72 9.3005
R228 GNDA.n94 GNDA.n93 9.3005
R229 GNDA.n95 GNDA.n71 9.3005
R230 GNDA.n97 GNDA.n96 9.3005
R231 GNDA.n98 GNDA.n70 9.3005
R232 GNDA.n100 GNDA.n99 9.3005
R233 GNDA.n102 GNDA.n101 9.3005
R234 GNDA.n103 GNDA.n68 9.3005
R235 GNDA.n105 GNDA.n104 9.3005
R236 GNDA.n107 GNDA.n106 9.3005
R237 GNDA.n108 GNDA.n66 9.3005
R238 GNDA.n110 GNDA.n109 9.3005
R239 GNDA.n111 GNDA.n65 9.3005
R240 GNDA.n113 GNDA.n112 9.3005
R241 GNDA.n64 GNDA.n63 9.3005
R242 GNDA.n124 GNDA.n123 9.3005
R243 GNDA.n125 GNDA.n62 9.3005
R244 GNDA.n127 GNDA.n126 9.3005
R245 GNDA.n128 GNDA.n61 9.3005
R246 GNDA.n130 GNDA.n129 9.3005
R247 GNDA.n131 GNDA.n60 9.3005
R248 GNDA.n133 GNDA.n132 9.3005
R249 GNDA.n134 GNDA.n59 9.3005
R250 GNDA.n136 GNDA.n135 9.3005
R251 GNDA.n138 GNDA.n137 9.3005
R252 GNDA.n140 GNDA.n56 9.3005
R253 GNDA.n142 GNDA.n141 9.3005
R254 GNDA.n143 GNDA.n55 9.3005
R255 GNDA.n145 GNDA.n144 9.3005
R256 GNDA.n146 GNDA.n54 9.3005
R257 GNDA.n148 GNDA.n147 9.3005
R258 GNDA.n149 GNDA.n53 9.3005
R259 GNDA.n151 GNDA.n150 9.3005
R260 GNDA.n34 GNDA.n27 9.3005
R261 GNDA.n36 GNDA.n35 9.3005
R262 GNDA.n37 GNDA.n26 9.3005
R263 GNDA.n40 GNDA.n39 9.3005
R264 GNDA.n41 GNDA.n25 9.3005
R265 GNDA.n43 GNDA.n42 9.3005
R266 GNDA.n44 GNDA.n23 9.3005
R267 GNDA.n49 GNDA.n48 9.3005
R268 GNDA.n47 GNDA.n24 9.3005
R269 GNDA.n46 GNDA.n45 9.3005
R270 GNDA.n22 GNDA.n21 9.3005
R271 GNDA.n165 GNDA.n164 9.3005
R272 GNDA.n166 GNDA.n20 9.3005
R273 GNDA.n168 GNDA.n167 9.3005
R274 GNDA.n169 GNDA.n18 9.3005
R275 GNDA.n172 GNDA.n171 9.3005
R276 GNDA.n173 GNDA.n17 9.3005
R277 GNDA.n175 GNDA.n174 9.3005
R278 GNDA.n177 GNDA.n15 9.3005
R279 GNDA.n179 GNDA.n178 9.3005
R280 GNDA.n180 GNDA.n14 9.3005
R281 GNDA.n182 GNDA.n181 9.3005
R282 GNDA.n184 GNDA.n12 9.3005
R283 GNDA.n186 GNDA.n185 9.3005
R284 GNDA.n187 GNDA.n11 9.3005
R285 GNDA.n189 GNDA.n188 9.3005
R286 GNDA.n190 GNDA.n10 9.3005
R287 GNDA.n192 GNDA.n191 9.3005
R288 GNDA.n193 GNDA.n9 9.3005
R289 GNDA.n195 GNDA.n194 9.3005
R290 GNDA.n197 GNDA.n6 9.3005
R291 GNDA.n200 GNDA.n199 9.3005
R292 GNDA.n201 GNDA.n5 9.3005
R293 GNDA.n203 GNDA.n202 9.3005
R294 GNDA.n204 GNDA.n4 9.3005
R295 GNDA.n206 GNDA.n205 9.3005
R296 GNDA.n207 GNDA.n3 9.3005
R297 GNDA.n209 GNDA.n208 9.3005
R298 GNDA.n210 GNDA.n1 9.3005
R299 GNDA.n33 GNDA.n32 7.49875
R300 GNDA.n93 GNDA.n92 6.4005
R301 GNDA.n114 GNDA.n113 6.4005
R302 GNDA.n122 GNDA.n62 6.4005
R303 GNDA.n135 GNDA.n58 6.4005
R304 GNDA.n140 GNDA.n139 6.4005
R305 GNDA.n152 GNDA.n151 6.4005
R306 GNDA.n50 GNDA.n49 6.4005
R307 GNDA.n164 GNDA.n163 6.4005
R308 GNDA.n177 GNDA.n176 6.4005
R309 GNDA.n184 GNDA.n183 6.4005
R310 GNDA.n196 GNDA.n195 6.4005
R311 GNDA.n211 GNDA.n210 6.4005
R312 GNDA.n156 GNDA.n8 5.68939
R313 GNDA.n118 GNDA.n117 5.68939
R314 GNDA.n118 GNDA.n57 5.68939
R315 GNDA.n156 GNDA.n7 4.97828
R316 GNDA.n86 GNDA.n85 3.2005
R317 GNDA.n99 GNDA.n69 3.2005
R318 GNDA.n87 GNDA.n75 0.245263
R319 GNDA.n32 GNDA.n27 0.194101
R320 GNDA.n150 GNDA.n0 0.193881
R321 GNDA.n212 GNDA.n1 0.193881
R322 GNDA.n88 GNDA.n87 0.15675
R323 GNDA.n89 GNDA.n88 0.15675
R324 GNDA.n89 GNDA.n72 0.15675
R325 GNDA.n94 GNDA.n72 0.15675
R326 GNDA.n95 GNDA.n94 0.15675
R327 GNDA.n96 GNDA.n95 0.15675
R328 GNDA.n96 GNDA.n70 0.15675
R329 GNDA.n100 GNDA.n70 0.15675
R330 GNDA.n101 GNDA.n100 0.15675
R331 GNDA.n101 GNDA.n68 0.15675
R332 GNDA.n105 GNDA.n68 0.15675
R333 GNDA.n106 GNDA.n105 0.15675
R334 GNDA.n106 GNDA.n66 0.15675
R335 GNDA.n110 GNDA.n66 0.15675
R336 GNDA.n111 GNDA.n110 0.15675
R337 GNDA.n112 GNDA.n111 0.15675
R338 GNDA.n112 GNDA.n63 0.15675
R339 GNDA.n124 GNDA.n63 0.15675
R340 GNDA.n125 GNDA.n124 0.15675
R341 GNDA.n126 GNDA.n125 0.15675
R342 GNDA.n126 GNDA.n61 0.15675
R343 GNDA.n130 GNDA.n61 0.15675
R344 GNDA.n131 GNDA.n130 0.15675
R345 GNDA.n132 GNDA.n131 0.15675
R346 GNDA.n132 GNDA.n59 0.15675
R347 GNDA.n136 GNDA.n59 0.15675
R348 GNDA.n137 GNDA.n136 0.15675
R349 GNDA.n137 GNDA.n56 0.15675
R350 GNDA.n142 GNDA.n56 0.15675
R351 GNDA.n143 GNDA.n142 0.15675
R352 GNDA.n144 GNDA.n143 0.15675
R353 GNDA.n144 GNDA.n54 0.15675
R354 GNDA.n148 GNDA.n54 0.15675
R355 GNDA.n149 GNDA.n148 0.15675
R356 GNDA.n150 GNDA.n149 0.15675
R357 GNDA.n36 GNDA.n27 0.15675
R358 GNDA.n37 GNDA.n36 0.15675
R359 GNDA.n39 GNDA.n25 0.15675
R360 GNDA.n43 GNDA.n25 0.15675
R361 GNDA.n44 GNDA.n43 0.15675
R362 GNDA.n48 GNDA.n44 0.15675
R363 GNDA.n48 GNDA.n47 0.15675
R364 GNDA.n47 GNDA.n46 0.15675
R365 GNDA.n46 GNDA.n21 0.15675
R366 GNDA.n165 GNDA.n21 0.15675
R367 GNDA.n166 GNDA.n165 0.15675
R368 GNDA.n167 GNDA.n166 0.15675
R369 GNDA.n167 GNDA.n18 0.15675
R370 GNDA.n172 GNDA.n18 0.15675
R371 GNDA.n173 GNDA.n172 0.15675
R372 GNDA.n174 GNDA.n173 0.15675
R373 GNDA.n174 GNDA.n15 0.15675
R374 GNDA.n179 GNDA.n15 0.15675
R375 GNDA.n180 GNDA.n179 0.15675
R376 GNDA.n181 GNDA.n180 0.15675
R377 GNDA.n181 GNDA.n12 0.15675
R378 GNDA.n186 GNDA.n12 0.15675
R379 GNDA.n187 GNDA.n186 0.15675
R380 GNDA.n188 GNDA.n187 0.15675
R381 GNDA.n188 GNDA.n10 0.15675
R382 GNDA.n192 GNDA.n10 0.15675
R383 GNDA.n193 GNDA.n192 0.15675
R384 GNDA.n194 GNDA.n193 0.15675
R385 GNDA.n194 GNDA.n6 0.15675
R386 GNDA.n200 GNDA.n6 0.15675
R387 GNDA.n201 GNDA.n200 0.15675
R388 GNDA.n202 GNDA.n201 0.15675
R389 GNDA.n202 GNDA.n4 0.15675
R390 GNDA.n206 GNDA.n4 0.15675
R391 GNDA.n207 GNDA.n206 0.15675
R392 GNDA.n208 GNDA.n207 0.15675
R393 GNDA.n208 GNDA.n1 0.15675
R394 GNDA.n38 GNDA.n37 0.109875
R395 GNDA.n39 GNDA.n38 0.047375
R396 before_Reset.n1 before_Reset.n0 481.334
R397 before_Reset.n0 before_Reset.t4 465.933
R398 before_Reset.n0 before_Reset.t3 321.334
R399 before_Reset.n2 before_Reset.n1 226.889
R400 before_Reset.n1 before_Reset.t1 172.458
R401 before_Reset.n2 before_Reset.t2 19.7005
R402 before_Reset.t0 before_Reset.n2 19.7005
R403 a_4210_n7910.t0 a_4210_n7910.n2 500.086
R404 a_4210_n7910.n1 a_4210_n7910.n0 473.334
R405 a_4210_n7910.n0 a_4210_n7910.t3 465.933
R406 a_4210_n7910.t0 a_4210_n7910.n2 461.389
R407 a_4210_n7910.n0 a_4210_n7910.t2 321.334
R408 a_4210_n7910.n1 a_4210_n7910.t1 177.577
R409 a_4210_n7910.n2 a_4210_n7910.n1 48.3899
R410 UP_PFD_b.n0 UP_PFD_b.t3 441.834
R411 UP_PFD_b.n0 UP_PFD_b.t2 313.3
R412 UP_PFD_b.n1 UP_PFD_b.n0 235.201
R413 UP_PFD_b.t0 UP_PFD_b.n1 219.528
R414 UP_PFD_b.n1 UP_PFD_b.t1 167.935
R415 QB_b.t6 QB_b.t3 1188.93
R416 QB_b QB_b.n2 899.734
R417 QB_b.t3 QB_b.t5 835.467
R418 QB_b.n2 QB_b.t4 562.333
R419 QB_b QB_b.n1 419.647
R420 QB_b.n1 QB_b.n0 247.917
R421 QB_b.n2 QB_b.t6 224.934
R422 QB_b.n1 QB_b.t0 221.411
R423 QB_b.n0 QB_b.t1 24.0005
R424 QB_b.n0 QB_b.t2 24.0005
R425 F.n4 F.n0 1319.38
R426 F.n0 F.t4 562.333
R427 F.n2 F.t3 388.813
R428 F.n2 F.t5 356.68
R429 F.n3 F.n2 232
R430 F.n0 F.t6 224.934
R431 F.t2 F.n4 221.411
R432 F.n3 F.n1 157.278
R433 F.n4 F.n3 90.64
R434 F.n1 F.t1 24.0005
R435 F.n1 F.t0 24.0005
R436 QA_b.t3 QA_b.t4 1188.93
R437 QA_b QA_b.n2 837.38
R438 QA_b.t4 QA_b.t6 835.467
R439 QA_b.n0 QA_b.t5 562.333
R440 QA_b QA_b.n0 482
R441 QA_b.n2 QA_b.n1 247.917
R442 QA_b.n0 QA_b.t3 224.934
R443 QA_b.n2 QA_b.t0 221.411
R444 QA_b.n1 QA_b.t1 24.0005
R445 QA_b.n1 QA_b.t2 24.0005
R446 Reset.n1 Reset.t3 562.333
R447 Reset.n2 Reset.n1 480.45
R448 Reset.n0 Reset.t4 417.733
R449 Reset.n0 Reset.t5 369.534
R450 Reset.n3 Reset.n2 328.733
R451 Reset.t0 Reset.n3 288.37
R452 Reset.n1 Reset.t2 224.934
R453 Reset.n3 Reset.t1 177.577
R454 Reset.n2 Reset.n0 176.733
R455 E_b.n0 E_b.t4 517.347
R456 E_b.n2 E_b.n0 417.574
R457 E_b.n2 E_b.n1 244.716
R458 E_b.n0 E_b.t3 228.148
R459 E_b.t1 E_b.n2 221.411
R460 E_b.n1 E_b.t0 24.0005
R461 E_b.n1 E_b.t2 24.0005
R462 DOWN.n0 DOWN.t2 605.311
R463 DOWN DOWN.t1 222.727
R464 DOWN.n0 DOWN.t0 148.736
R465 DOWN DOWN.n0 17.6005
R466 I_IN I_IN.t0 241.928
R467 I_IN I_IN.t1 158.335
R468 DOWN_input.n0 DOWN_input.t0 229.127
R469 DOWN_input.n0 DOWN_input.t2 158.335
R470 DOWN_input.n2 DOWN_input.t1 158.335
R471 DOWN_input.n2 DOWN_input.n0 124.8
R472 DOWN_input DOWN_input.n2 6.4005
R473 DOWN_input.n2 DOWN_input.n1 6.4005
R474 a_2350_n7910.t0 a_2350_n7910.t1 39.4005
R475 VDDA.n222 VDDA.n214 831.25
R476 VDDA.n217 VDDA.n216 831.25
R477 VDDA.n211 VDDA.n203 831.25
R478 VDDA.n206 VDDA.n205 831.25
R479 VDDA.n215 VDDA.n214 585
R480 VDDA.n219 VDDA.n217 585
R481 VDDA.n109 VDDA.n104 585
R482 VDDA.n104 VDDA.n41 585
R483 VDDA.n118 VDDA.n113 585
R484 VDDA.n113 VDDA.n45 585
R485 VDDA.n132 VDDA.n127 585
R486 VDDA.n127 VDDA.n48 585
R487 VDDA.n60 VDDA.n54 585
R488 VDDA.n55 VDDA.n54 585
R489 VDDA.n204 VDDA.n203 585
R490 VDDA.n208 VDDA.n206 585
R491 VDDA.n98 VDDA.n42 585
R492 VDDA.n98 VDDA.n97 585
R493 VDDA.n136 VDDA.n49 585
R494 VDDA.n121 VDDA.n49 585
R495 VDDA.n221 VDDA.t22 465.079
R496 VDDA.t22 VDDA.n220 465.079
R497 VDDA.n210 VDDA.t17 465.079
R498 VDDA.t17 VDDA.n209 465.079
R499 VDDA.t7 VDDA.n86 464.281
R500 VDDA.n88 VDDA.t7 464.281
R501 VDDA.t38 VDDA.n195 464.281
R502 VDDA.n196 VDDA.t38 464.281
R503 VDDA.n238 VDDA.t25 464.281
R504 VDDA.t25 VDDA.n237 464.281
R505 VDDA.n244 VDDA.t11 464.281
R506 VDDA.t11 VDDA.n18 464.281
R507 VDDA.n29 VDDA.t34 464.281
R508 VDDA.t34 VDDA.n26 464.281
R509 VDDA.n83 VDDA.t40 464.281
R510 VDDA.t40 VDDA.n82 464.281
R511 VDDA.t15 VDDA.n187 464.281
R512 VDDA.n188 VDDA.t15 464.281
R513 VDDA.t24 VDDA.n227 464.281
R514 VDDA.n228 VDDA.t24 464.281
R515 VDDA.n178 VDDA.t1 464.281
R516 VDDA.t1 VDDA.n177 464.281
R517 VDDA.t4 VDDA.n71 464.281
R518 VDDA.n72 VDDA.t4 464.281
R519 VDDA.n141 VDDA.t41 415.336
R520 VDDA.n23 VDDA.t31 315.25
R521 VDDA.t19 VDDA.t26 314.113
R522 VDDA.t18 VDDA.t5 314.113
R523 VDDA.n107 VDDA.n104 290.733
R524 VDDA.n116 VDDA.n113 290.733
R525 VDDA.n130 VDDA.n127 290.733
R526 VDDA.n58 VDDA.n54 290.733
R527 VDDA.n99 VDDA.n98 290.733
R528 VDDA.n122 VDDA.n49 290.733
R529 VDDA.n195 VDDA.n184 243.698
R530 VDDA.n239 VDDA.n238 243.698
R531 VDDA.n245 VDDA.n244 243.698
R532 VDDA.n29 VDDA.n28 243.698
R533 VDDA.n84 VDDA.n83 243.698
R534 VDDA.n188 VDDA.n185 243.698
R535 VDDA.n228 VDDA.n225 243.698
R536 VDDA.n177 VDDA.n21 243.698
R537 VDDA.n72 VDDA.n69 243.698
R538 VDDA.n223 VDDA.n222 238.367
R539 VDDA.n216 VDDA.n183 238.367
R540 VDDA.n182 VDDA.n13 238.367
R541 VDDA.n248 VDDA.n247 238.367
R542 VDDA.n34 VDDA.n33 238.367
R543 VDDA.n68 VDDA.n38 238.367
R544 VDDA.n192 VDDA.n2 238.367
R545 VDDA.n212 VDDA.n211 238.367
R546 VDDA.n232 VDDA.n14 238.367
R547 VDDA.n180 VDDA.n179 238.367
R548 VDDA.n76 VDDA.n25 238.367
R549 VDDA.n205 VDDA.n201 238.367
R550 VDDA.n199 VDDA.n1 238.367
R551 VDDA.n110 VDDA.n109 230.308
R552 VDDA.n65 VDDA.n41 230.308
R553 VDDA.n119 VDDA.n118 230.308
R554 VDDA.n64 VDDA.n45 230.308
R555 VDDA.n133 VDDA.n132 230.308
R556 VDDA.n63 VDDA.n48 230.308
R557 VDDA.n61 VDDA.n60 230.308
R558 VDDA.n55 VDDA.n52 230.308
R559 VDDA.n102 VDDA.n42 230.308
R560 VDDA.n136 VDDA.n135 230.308
R561 VDDA.n125 VDDA.n121 230.308
R562 VDDA.n97 VDDA.n94 230.308
R563 VDDA.t12 VDDA.t2 222.178
R564 VDDA.n111 VDDA.n93 199.195
R565 VDDA.n88 VDDA.n67 190.333
R566 VDDA.n51 VDDA.n50 185
R567 VDDA.n124 VDDA.n123 185
R568 VDDA.n101 VDDA.n100 185
R569 VDDA.n96 VDDA.n95 185
R570 VDDA.n75 VDDA.n74 185
R571 VDDA.n73 VDDA.n70 185
R572 VDDA.n174 VDDA.n22 185
R573 VDDA.n176 VDDA.n175 185
R574 VDDA.n231 VDDA.n230 185
R575 VDDA.n229 VDDA.n226 185
R576 VDDA.n204 VDDA.n202 185
R577 VDDA.n208 VDDA.n207 185
R578 VDDA.n191 VDDA.n190 185
R579 VDDA.n189 VDDA.n186 185
R580 VDDA.n59 VDDA.n53 185
R581 VDDA.n57 VDDA.n56 185
R582 VDDA.n131 VDDA.n126 185
R583 VDDA.n129 VDDA.n128 185
R584 VDDA.n117 VDDA.n112 185
R585 VDDA.n115 VDDA.n114 185
R586 VDDA.n108 VDDA.n103 185
R587 VDDA.n106 VDDA.n105 185
R588 VDDA.n79 VDDA.n78 185
R589 VDDA.n81 VDDA.n80 185
R590 VDDA.n30 VDDA.n27 185
R591 VDDA.n32 VDDA.n31 185
R592 VDDA.n243 VDDA.n241 185
R593 VDDA.n242 VDDA.n19 185
R594 VDDA.n234 VDDA.n233 185
R595 VDDA.n236 VDDA.n235 185
R596 VDDA.n215 VDDA.n213 185
R597 VDDA.n219 VDDA.n218 185
R598 VDDA.n194 VDDA.n193 185
R599 VDDA.n198 VDDA.n197 185
R600 VDDA.n92 VDDA.n37 185
R601 VDDA.n93 VDDA.n92 185
R602 VDDA.n91 VDDA.n90 185
R603 VDDA.n89 VDDA.n87 185
R604 VDDA.n93 VDDA.n67 185
R605 VDDA.t2 VDDA.n62 172.38
R606 VDDA.n134 VDDA.t27 172.38
R607 VDDA.n120 VDDA.t8 172.38
R608 VDDA.n198 VDDA.n193 150
R609 VDDA.n218 VDDA.n213 150
R610 VDDA.n235 VDDA.n233 150
R611 VDDA.n241 VDDA.n19 150
R612 VDDA.n32 VDDA.n27 150
R613 VDDA.n80 VDDA.n78 150
R614 VDDA.n191 VDDA.n186 150
R615 VDDA.n207 VDDA.n202 150
R616 VDDA.n231 VDDA.n226 150
R617 VDDA.n175 VDDA.n22 150
R618 VDDA.n75 VDDA.n70 150
R619 VDDA.n92 VDDA.n91 150
R620 VDDA.n87 VDDA.n67 150
R621 VDDA.n85 VDDA.n77 137.904
R622 VDDA.n181 VDDA.n20 137.904
R623 VDDA.n62 VDDA.t36 126.412
R624 VDDA.n134 VDDA.t12 126.412
R625 VDDA.t27 VDDA.n120 126.412
R626 VDDA.t8 VDDA.n111 126.412
R627 VDDA.t29 VDDA.n214 123.126
R628 VDDA.n217 VDDA.t29 123.126
R629 VDDA.t21 VDDA.n203 123.126
R630 VDDA.n206 VDDA.t21 123.126
R631 VDDA.n105 VDDA.n103 120.001
R632 VDDA.n114 VDDA.n112 120.001
R633 VDDA.n128 VDDA.n126 120.001
R634 VDDA.n56 VDDA.n53 120.001
R635 VDDA.n101 VDDA.n95 120.001
R636 VDDA.n124 VDDA.n51 120.001
R637 VDDA.n246 VDDA.n240 107.258
R638 VDDA.n240 VDDA.t23 103.427
R639 VDDA.t16 VDDA.n224 103.427
R640 VDDA.n224 VDDA.t20 103.427
R641 VDDA.t14 VDDA.n200 103.427
R642 VDDA.n246 VDDA.t0 95.7666
R643 VDDA.t39 VDDA.t6 91.936
R644 VDDA.t33 VDDA.t3 91.936
R645 VDDA.t10 VDDA.t30 84.2747
R646 VDDA.t23 VDDA.t19 84.2747
R647 VDDA.t26 VDDA.t16 84.2747
R648 VDDA.t20 VDDA.t18 84.2747
R649 VDDA.t5 VDDA.t14 84.2747
R650 VDDA.n135 VDDA.n134 69.8479
R651 VDDA.n134 VDDA.n125 69.8479
R652 VDDA.n111 VDDA.n102 69.8479
R653 VDDA.n111 VDDA.n94 69.8479
R654 VDDA.n62 VDDA.n61 69.8479
R655 VDDA.n62 VDDA.n52 69.8479
R656 VDDA.n134 VDDA.n133 69.8479
R657 VDDA.n134 VDDA.n63 69.8479
R658 VDDA.n120 VDDA.n119 69.8479
R659 VDDA.n120 VDDA.n64 69.8479
R660 VDDA.n111 VDDA.n110 69.8479
R661 VDDA.n111 VDDA.n65 69.8479
R662 VDDA.n55 VDDA.n47 68.0425
R663 VDDA.n77 VDDA.n76 65.8183
R664 VDDA.n77 VDDA.n69 65.8183
R665 VDDA.n181 VDDA.n180 65.8183
R666 VDDA.n181 VDDA.n21 65.8183
R667 VDDA.n240 VDDA.n232 65.8183
R668 VDDA.n240 VDDA.n225 65.8183
R669 VDDA.n224 VDDA.n212 65.8183
R670 VDDA.n224 VDDA.n201 65.8183
R671 VDDA.n200 VDDA.n192 65.8183
R672 VDDA.n200 VDDA.n185 65.8183
R673 VDDA.n85 VDDA.n84 65.8183
R674 VDDA.n85 VDDA.n68 65.8183
R675 VDDA.n28 VDDA.n20 65.8183
R676 VDDA.n33 VDDA.n20 65.8183
R677 VDDA.n246 VDDA.n245 65.8183
R678 VDDA.n247 VDDA.n246 65.8183
R679 VDDA.n240 VDDA.n239 65.8183
R680 VDDA.n240 VDDA.n182 65.8183
R681 VDDA.n224 VDDA.n223 65.8183
R682 VDDA.n224 VDDA.n183 65.8183
R683 VDDA.n200 VDDA.n184 65.8183
R684 VDDA.n200 VDDA.n199 65.8183
R685 VDDA.n93 VDDA.n66 65.8183
R686 VDDA.n283 VDDA.n1 58.0576
R687 VDDA.n255 VDDA.n13 58.0576
R688 VDDA.n249 VDDA.n248 58.0576
R689 VDDA.n166 VDDA.n34 58.0576
R690 VDDA.n159 VDDA.n38 58.0576
R691 VDDA.n283 VDDA.n2 58.0576
R692 VDDA.n255 VDDA.n14 58.0576
R693 VDDA.n179 VDDA.n173 58.0576
R694 VDDA.n167 VDDA.n25 58.0576
R695 VDDA.n160 VDDA.n37 58.0576
R696 VDDA.n151 VDDA.n41 57.2449
R697 VDDA.n144 VDDA.n45 57.2449
R698 VDDA.n137 VDDA.n48 57.2449
R699 VDDA.n151 VDDA.n42 57.2449
R700 VDDA.n137 VDDA.n136 57.2449
R701 VDDA.n270 VDDA.n7 54.4005
R702 VDDA.n268 VDDA.n7 54.4005
R703 VDDA.n268 VDDA.n8 54.4005
R704 VDDA.n270 VDDA.n8 54.4005
R705 VDDA.n193 VDDA.n184 53.3664
R706 VDDA.n199 VDDA.n198 53.3664
R707 VDDA.n186 VDDA.n185 53.3664
R708 VDDA.n207 VDDA.n201 53.3664
R709 VDDA.n226 VDDA.n225 53.3664
R710 VDDA.n76 VDDA.n75 53.3664
R711 VDDA.n70 VDDA.n69 53.3664
R712 VDDA.n180 VDDA.n22 53.3664
R713 VDDA.n175 VDDA.n21 53.3664
R714 VDDA.n232 VDDA.n231 53.3664
R715 VDDA.n212 VDDA.n202 53.3664
R716 VDDA.n192 VDDA.n191 53.3664
R717 VDDA.n84 VDDA.n78 53.3664
R718 VDDA.n80 VDDA.n68 53.3664
R719 VDDA.n28 VDDA.n27 53.3664
R720 VDDA.n33 VDDA.n32 53.3664
R721 VDDA.n245 VDDA.n241 53.3664
R722 VDDA.n247 VDDA.n19 53.3664
R723 VDDA.n239 VDDA.n233 53.3664
R724 VDDA.n235 VDDA.n182 53.3664
R725 VDDA.n223 VDDA.n213 53.3664
R726 VDDA.n218 VDDA.n183 53.3664
R727 VDDA.n91 VDDA.n66 53.3664
R728 VDDA.n87 VDDA.n66 53.3664
R729 VDDA.n95 VDDA.n94 45.3071
R730 VDDA.n125 VDDA.n124 45.3071
R731 VDDA.n135 VDDA.n51 45.3071
R732 VDDA.n102 VDDA.n101 45.3071
R733 VDDA.n61 VDDA.n53 45.3071
R734 VDDA.n56 VDDA.n52 45.3071
R735 VDDA.n133 VDDA.n126 45.3071
R736 VDDA.n128 VDDA.n63 45.3071
R737 VDDA.n119 VDDA.n112 45.3071
R738 VDDA.n114 VDDA.n64 45.3071
R739 VDDA.n110 VDDA.n103 45.3071
R740 VDDA.n105 VDDA.n65 45.3071
R741 VDDA.n284 VDDA.n283 34.9005
R742 VDDA.n138 VDDA.n137 32.0005
R743 VDDA.n138 VDDA.n46 32.0005
R744 VDDA.n143 VDDA.n46 32.0005
R745 VDDA.n146 VDDA.n145 32.0005
R746 VDDA.n146 VDDA.n43 32.0005
R747 VDDA.n150 VDDA.n43 32.0005
R748 VDDA.n153 VDDA.n152 32.0005
R749 VDDA.n153 VDDA.n39 32.0005
R750 VDDA.n157 VDDA.n39 32.0005
R751 VDDA.n158 VDDA.n157 32.0005
R752 VDDA.n161 VDDA.n35 32.0005
R753 VDDA.n165 VDDA.n35 32.0005
R754 VDDA.n169 VDDA.n168 32.0005
R755 VDDA.n250 VDDA.n17 32.0005
R756 VDDA.n254 VDDA.n15 32.0005
R757 VDDA.n257 VDDA.n256 32.0005
R758 VDDA.n257 VDDA.n11 32.0005
R759 VDDA.n261 VDDA.n11 32.0005
R760 VDDA.n262 VDDA.n261 32.0005
R761 VDDA.n263 VDDA.n262 32.0005
R762 VDDA.n263 VDDA.n9 32.0005
R763 VDDA.n267 VDDA.n9 32.0005
R764 VDDA.n271 VDDA.n5 32.0005
R765 VDDA.n275 VDDA.n5 32.0005
R766 VDDA.n276 VDDA.n275 32.0005
R767 VDDA.n277 VDDA.n276 32.0005
R768 VDDA.n277 VDDA.n3 32.0005
R769 VDDA.n281 VDDA.n3 32.0005
R770 VDDA.n282 VDDA.n281 32.0005
R771 VDDA.n144 VDDA.n143 28.8005
R772 VDDA.n151 VDDA.n150 25.6005
R773 VDDA.n161 VDDA.n160 25.6005
R774 VDDA.n173 VDDA.n172 25.6005
R775 VDDA.n249 VDDA.n15 25.6005
R776 VDDA.n255 VDDA.n254 25.6005
R777 VDDA.n269 VDDA.n268 25.6005
R778 VDDA.n270 VDDA.n269 25.6005
R779 VDDA.n104 VDDA.t32 24.6255
R780 VDDA.n113 VDDA.t28 24.6255
R781 VDDA.n127 VDDA.t35 24.6255
R782 VDDA.n54 VDDA.t37 24.6255
R783 VDDA.n98 VDDA.t9 24.6255
R784 VDDA.n49 VDDA.t13 24.6255
R785 VDDA.n169 VDDA.n23 19.2005
R786 VDDA.n168 VDDA.n167 16.0005
R787 VDDA.n166 VDDA.n165 12.8005
R788 VDDA.n172 VDDA.n23 12.8005
R789 VDDA.n93 VDDA.t39 11.4924
R790 VDDA.t6 VDDA.n85 11.4924
R791 VDDA.n77 VDDA.t33 11.4924
R792 VDDA.t3 VDDA.n20 11.4924
R793 VDDA.t30 VDDA.n181 11.4924
R794 VDDA.n139 VDDA.n138 9.3005
R795 VDDA.n140 VDDA.n46 9.3005
R796 VDDA.n143 VDDA.n142 9.3005
R797 VDDA.n145 VDDA.n44 9.3005
R798 VDDA.n147 VDDA.n146 9.3005
R799 VDDA.n148 VDDA.n43 9.3005
R800 VDDA.n150 VDDA.n149 9.3005
R801 VDDA.n152 VDDA.n40 9.3005
R802 VDDA.n154 VDDA.n153 9.3005
R803 VDDA.n155 VDDA.n39 9.3005
R804 VDDA.n157 VDDA.n156 9.3005
R805 VDDA.n158 VDDA.n36 9.3005
R806 VDDA.n162 VDDA.n161 9.3005
R807 VDDA.n163 VDDA.n35 9.3005
R808 VDDA.n165 VDDA.n164 9.3005
R809 VDDA.n168 VDDA.n24 9.3005
R810 VDDA.n170 VDDA.n169 9.3005
R811 VDDA.n172 VDDA.n171 9.3005
R812 VDDA.n17 VDDA.n16 9.3005
R813 VDDA.n251 VDDA.n250 9.3005
R814 VDDA.n252 VDDA.n15 9.3005
R815 VDDA.n254 VDDA.n253 9.3005
R816 VDDA.n256 VDDA.n12 9.3005
R817 VDDA.n258 VDDA.n257 9.3005
R818 VDDA.n259 VDDA.n11 9.3005
R819 VDDA.n261 VDDA.n260 9.3005
R820 VDDA.n262 VDDA.n10 9.3005
R821 VDDA.n264 VDDA.n263 9.3005
R822 VDDA.n265 VDDA.n9 9.3005
R823 VDDA.n267 VDDA.n266 9.3005
R824 VDDA.n269 VDDA.n6 9.3005
R825 VDDA.n272 VDDA.n271 9.3005
R826 VDDA.n273 VDDA.n5 9.3005
R827 VDDA.n275 VDDA.n274 9.3005
R828 VDDA.n276 VDDA.n4 9.3005
R829 VDDA.n278 VDDA.n277 9.3005
R830 VDDA.n279 VDDA.n3 9.3005
R831 VDDA.n281 VDDA.n280 9.3005
R832 VDDA.n282 VDDA.n0 9.3005
R833 VDDA.n197 VDDA.n194 9.14336
R834 VDDA.n236 VDDA.n234 9.14336
R835 VDDA.n243 VDDA.n242 9.14336
R836 VDDA.n31 VDDA.n30 9.14336
R837 VDDA.n81 VDDA.n79 9.14336
R838 VDDA.n190 VDDA.n189 9.14336
R839 VDDA.n230 VDDA.n229 9.14336
R840 VDDA.n176 VDDA.n174 9.14336
R841 VDDA.n74 VDDA.n73 9.14336
R842 VDDA.n90 VDDA.n89 9.14336
R843 VDDA.t0 VDDA.t10 7.66179
R844 VDDA.n137 VDDA.n47 7.49875
R845 VDDA.n109 VDDA.n108 7.11161
R846 VDDA.n106 VDDA.n41 7.11161
R847 VDDA.n118 VDDA.n117 7.11161
R848 VDDA.n115 VDDA.n45 7.11161
R849 VDDA.n132 VDDA.n131 7.11161
R850 VDDA.n129 VDDA.n48 7.11161
R851 VDDA.n60 VDDA.n59 7.11161
R852 VDDA.n57 VDDA.n55 7.11161
R853 VDDA.n100 VDDA.n42 7.11161
R854 VDDA.n97 VDDA.n96 7.11161
R855 VDDA.n136 VDDA.n50 7.11161
R856 VDDA.n123 VDDA.n121 7.11161
R857 VDDA.n152 VDDA.n151 6.4005
R858 VDDA.n173 VDDA.n17 6.4005
R859 VDDA.n250 VDDA.n249 6.4005
R860 VDDA.n256 VDDA.n255 6.4005
R861 VDDA.n268 VDDA.n267 6.4005
R862 VDDA.n271 VDDA.n270 6.4005
R863 VDDA.n283 VDDA.n282 6.4005
R864 VDDA.n219 VDDA.n215 5.81868
R865 VDDA.n208 VDDA.n204 5.81868
R866 VDDA.n86 VDDA.n37 5.33286
R867 VDDA.n196 VDDA.n1 5.33286
R868 VDDA.n237 VDDA.n13 5.33286
R869 VDDA.n248 VDDA.n18 5.33286
R870 VDDA.n34 VDDA.n26 5.33286
R871 VDDA.n82 VDDA.n38 5.33286
R872 VDDA.n187 VDDA.n2 5.33286
R873 VDDA.n227 VDDA.n14 5.33286
R874 VDDA.n179 VDDA.n178 5.33286
R875 VDDA.n71 VDDA.n25 5.33286
R876 VDDA.n195 VDDA.n194 3.75335
R877 VDDA.n197 VDDA.n196 3.75335
R878 VDDA.n238 VDDA.n234 3.75335
R879 VDDA.n237 VDDA.n236 3.75335
R880 VDDA.n244 VDDA.n243 3.75335
R881 VDDA.n242 VDDA.n18 3.75335
R882 VDDA.n30 VDDA.n29 3.75335
R883 VDDA.n31 VDDA.n26 3.75335
R884 VDDA.n83 VDDA.n79 3.75335
R885 VDDA.n82 VDDA.n81 3.75335
R886 VDDA.n190 VDDA.n187 3.75335
R887 VDDA.n189 VDDA.n188 3.75335
R888 VDDA.n230 VDDA.n227 3.75335
R889 VDDA.n229 VDDA.n228 3.75335
R890 VDDA.n178 VDDA.n174 3.75335
R891 VDDA.n177 VDDA.n176 3.75335
R892 VDDA.n74 VDDA.n71 3.75335
R893 VDDA.n73 VDDA.n72 3.75335
R894 VDDA.n90 VDDA.n86 3.75335
R895 VDDA.n89 VDDA.n88 3.75335
R896 VDDA.n108 VDDA.n107 3.53508
R897 VDDA.n107 VDDA.n106 3.53508
R898 VDDA.n117 VDDA.n116 3.53508
R899 VDDA.n116 VDDA.n115 3.53508
R900 VDDA.n131 VDDA.n130 3.53508
R901 VDDA.n130 VDDA.n129 3.53508
R902 VDDA.n59 VDDA.n58 3.53508
R903 VDDA.n58 VDDA.n57 3.53508
R904 VDDA.n100 VDDA.n99 3.53508
R905 VDDA.n99 VDDA.n96 3.53508
R906 VDDA.n122 VDDA.n50 3.53508
R907 VDDA.n123 VDDA.n122 3.53508
R908 VDDA.n222 VDDA.n221 3.40194
R909 VDDA.n220 VDDA.n216 3.40194
R910 VDDA.n211 VDDA.n210 3.40194
R911 VDDA.n209 VDDA.n205 3.40194
R912 VDDA.n145 VDDA.n144 3.2005
R913 VDDA.n159 VDDA.n158 3.2005
R914 VDDA.n160 VDDA.n159 3.2005
R915 VDDA.n167 VDDA.n166 3.2005
R916 VDDA.n221 VDDA.n215 2.39444
R917 VDDA.n220 VDDA.n219 2.39444
R918 VDDA.n210 VDDA.n204 2.39444
R919 VDDA.n209 VDDA.n208 2.39444
R920 VDDA.n216 VDDA.n7 2.32777
R921 VDDA.n211 VDDA.n8 2.32777
R922 VDDA.n139 VDDA.n47 0.194101
R923 VDDA.n140 VDDA.n139 0.15675
R924 VDDA.n142 VDDA.n44 0.15675
R925 VDDA.n147 VDDA.n44 0.15675
R926 VDDA.n148 VDDA.n147 0.15675
R927 VDDA.n149 VDDA.n148 0.15675
R928 VDDA.n149 VDDA.n40 0.15675
R929 VDDA.n154 VDDA.n40 0.15675
R930 VDDA.n155 VDDA.n154 0.15675
R931 VDDA.n156 VDDA.n155 0.15675
R932 VDDA.n156 VDDA.n36 0.15675
R933 VDDA.n162 VDDA.n36 0.15675
R934 VDDA.n163 VDDA.n162 0.15675
R935 VDDA.n164 VDDA.n163 0.15675
R936 VDDA.n164 VDDA.n24 0.15675
R937 VDDA.n170 VDDA.n24 0.15675
R938 VDDA.n171 VDDA.n170 0.15675
R939 VDDA.n171 VDDA.n16 0.15675
R940 VDDA.n251 VDDA.n16 0.15675
R941 VDDA.n252 VDDA.n251 0.15675
R942 VDDA.n253 VDDA.n252 0.15675
R943 VDDA.n253 VDDA.n12 0.15675
R944 VDDA.n258 VDDA.n12 0.15675
R945 VDDA.n259 VDDA.n258 0.15675
R946 VDDA.n260 VDDA.n259 0.15675
R947 VDDA.n260 VDDA.n10 0.15675
R948 VDDA.n264 VDDA.n10 0.15675
R949 VDDA.n265 VDDA.n264 0.15675
R950 VDDA.n266 VDDA.n265 0.15675
R951 VDDA.n266 VDDA.n6 0.15675
R952 VDDA.n272 VDDA.n6 0.15675
R953 VDDA.n273 VDDA.n272 0.15675
R954 VDDA.n274 VDDA.n273 0.15675
R955 VDDA.n274 VDDA.n4 0.15675
R956 VDDA.n278 VDDA.n4 0.15675
R957 VDDA.n279 VDDA.n278 0.15675
R958 VDDA.n280 VDDA.n279 0.15675
R959 VDDA.n280 VDDA.n0 0.15675
R960 VDDA.n284 VDDA.n0 0.15675
R961 VDDA VDDA.n284 0.1255
R962 VDDA.n141 VDDA.n140 0.078625
R963 VDDA.n142 VDDA.n141 0.078625
R964 a_3770_n7290.t0 a_3770_n7290.t1 48.0005
R965 a_2350_n8670.t0 a_2350_n8670.t1 39.4005
R966 a_4060_n9120.t1 a_4060_n9120.n2 500.086
R967 a_4060_n9120.n1 a_4060_n9120.n0 473.334
R968 a_4060_n9120.n0 a_4060_n9120.t3 465.933
R969 a_4060_n9120.t1 a_4060_n9120.n2 461.389
R970 a_4060_n9120.n0 a_4060_n9120.t2 321.334
R971 a_4060_n9120.n1 a_4060_n9120.t0 177.577
R972 a_4060_n9120.n2 a_4060_n9120.n1 48.3898
R973 a_3730_n9120.t1 a_3730_n9120.n2 500.086
R974 a_3730_n9120.n1 a_3730_n9120.n0 473.334
R975 a_3730_n9120.n0 a_3730_n9120.t3 465.933
R976 a_3730_n9120.t1 a_3730_n9120.n2 461.389
R977 a_3730_n9120.n0 a_3730_n9120.t2 321.334
R978 a_3730_n9120.n1 a_3730_n9120.t0 177.577
R979 a_3730_n9120.n2 a_3730_n9120.n1 48.3898
R980 a_4390_n9120.t1 a_4390_n9120.n2 500.086
R981 a_4390_n9120.n0 a_4390_n9120.t3 465.933
R982 a_4390_n9120.t1 a_4390_n9120.n2 461.389
R983 a_4390_n9120.n1 a_4390_n9120.n0 392.623
R984 a_4390_n9120.n0 a_4390_n9120.t2 321.334
R985 a_4390_n9120.n1 a_4390_n9120.t0 177.577
R986 a_4390_n9120.n2 a_4390_n9120.n1 48.3899
R987 a_1830_n7910.t0 a_1830_n7910.t1 39.4005
R988 a_3250_n7910.t0 a_3250_n7910.t1 39.4005
R989 QB.t6 QB.t5 835.467
R990 QB.n1 QB.t6 564.496
R991 QB.n2 QB.t4 517.347
R992 QB.n0 QB.t3 514.134
R993 QB.n1 QB.n0 455.219
R994 QB.n5 QB.n2 363.2
R995 QB.n0 QB.t7 273.134
R996 QB.n4 QB.n3 244.716
R997 QB.n2 QB.t8 228.148
R998 QB.n4 QB.t0 221.411
R999 QB.n5 QB.n4 54.3734
R1000 QB QB.n1 26.7568
R1001 QB.n3 QB.t2 24.0005
R1002 QB.n3 QB.t1 24.0005
R1003 QB QB.n5 6.4005
R1004 DOWN_PFD_b.t1 DOWN_PFD_b.n1 203.528
R1005 DOWN_PFD_b.n0 DOWN_PFD_b.t2 203.528
R1006 DOWN_PFD_b.n1 DOWN_PFD_b.t0 183.935
R1007 DOWN_PFD_b.n0 DOWN_PFD_b.t3 183.935
R1008 DOWN_PFD_b.n1 DOWN_PFD_b.n0 83.2005
R1009 a_1830_n8670.t0 a_1830_n8670.t1 39.4005
R1010 DOWN_b.n0 DOWN_b.t5 1028.27
R1011 DOWN_b.n2 DOWN_b.n1 569.734
R1012 DOWN_b.n1 DOWN_b.n0 465.933
R1013 DOWN_b.n1 DOWN_b.t2 401.668
R1014 DOWN_b.n0 DOWN_b.t3 385.601
R1015 DOWN_b.n1 DOWN_b.t4 385.601
R1016 DOWN_b.t0 DOWN_b.n2 211.847
R1017 DOWN_b.n2 DOWN_b.t1 173.055
R1018 a_2730_n7910.t0 a_2730_n7910.t1 39.4005
R1019 a_3250_n8670.t0 a_3250_n8670.t1 39.4005
R1020 F_b.n0 F_b.t3 517.347
R1021 F_b.n2 F_b.n0 417.574
R1022 F_b.n2 F_b.n1 244.716
R1023 F_b.n0 F_b.t4 228.148
R1024 F_b.t0 F_b.n2 221.411
R1025 F_b.n1 F_b.t2 24.0005
R1026 F_b.n1 F_b.t1 24.0005
R1027 a_2730_n8670.t0 a_2730_n8670.t1 39.4005
R1028 F_REF.n0 F_REF.t1 514.134
R1029 F_REF.n0 F_REF.t0 273.134
R1030 F_REF F_REF.n0 216.9
R1031 UP.n0 UP.t3 1205
R1032 UP.n2 UP.t5 522.168
R1033 UP.n1 UP.n0 441.834
R1034 UP.n3 UP.n2 235.201
R1035 UP.t1 UP.n3 229.127
R1036 UP.n1 UP.t4 217.905
R1037 UP.n0 UP.t2 208.868
R1038 UP.n3 UP.t0 158.335
R1039 UP.n2 UP.n1 15.063
R1040 opamp_out opamp_out.t1 225.928
R1041 opamp_out opamp_out.t0 174.335
R1042 UP_input.n0 UP_input.t2 241.928
R1043 UP_input.n2 UP_input.t1 241.928
R1044 UP_input.n0 UP_input.t0 145.536
R1045 UP_input.n2 UP_input.n0 124.8
R1046 UP_input UP_input.n2 6.4005
R1047 UP_input.n2 UP_input.n1 6.4005
R1048 F_VCO.n0 F_VCO.t0 514.134
R1049 F_VCO.n0 F_VCO.t1 273.134
R1050 F_VCO F_VCO.n0 216.9
R1051 UP_b.n0 UP_b.t2 778.601
R1052 UP_b.n0 UP_b.t1 209.928
R1053 UP_b UP_b.t0 161.536
R1054 UP_b UP_b.n0 16.0005
C0 F_REF QA_b 0.026369f
C1 VDDA QA 0.550605f
C2 I_IN VDDA 0.051398f
C3 VDDA opamp_out 0.042251f
C4 VDDA DOWN_input 0.153934f
C5 F_REF VDDA 0.085173f
C6 I_IN DOWN_input 0.243956f
C7 F_REF QA 0.056f
C8 VDDA UP_input 0.356612f
C9 UP_input opamp_out 0.243956f
C10 VDDA DOWN 0.197633f
C11 QB_b QB 0.388258f
C12 I_IN DOWN 0.2232f
C13 QB_b F_VCO 0.026369f
C14 DOWN_input DOWN 0.013059f
C15 VDDA UP_b 0.293124f
C16 QB_b VDDA 0.511838f
C17 UP_b opamp_out 0.234797f
C18 VDDA QA_b 0.52066f
C19 QB F_VCO 0.056153f
C20 QA_b QA 0.422694f
C21 UP_b UP_input 0.022182f
C22 VDDA QB 2.75002f
C23 VDDA F_VCO 0.085127f
C24 QB QA 0.074487f
C25 DOWN_input GNDA 0.391369f
C26 I_IN GNDA 0.049563f
C27 DOWN GNDA 0.327262f
C28 F_VCO GNDA 0.236218f
C29 UP_input GNDA 0.317125f
C30 opamp_out GNDA 0.050519f
C31 UP_b GNDA 0.218542f
C32 F_REF GNDA 0.236218f
C33 VDDA GNDA 20.080345f
C34 QB_b GNDA 1.06408f
C35 QB GNDA 1.310209f
C36 QA GNDA 3.10607f
C37 QA_b GNDA 1.05212f
C38 QB.t3 GNDA 0.069179f
C39 QB.t7 GNDA 0.032493f
C40 QB.n0 GNDA 0.099932f
C41 QB.t5 GNDA 0.069179f
C42 QB.t6 GNDA 0.104293f
C43 QB.n1 GNDA 1.25065f
C44 QB.t4 GNDA 0.069862f
C45 QB.t8 GNDA 0.030633f
C46 QB.n2 GNDA 0.176466f
C47 QB.t0 GNDA 0.147114f
C48 QB.t2 GNDA 0.027951f
C49 QB.t1 GNDA 0.027951f
C50 QB.n3 GNDA 0.149246f
C51 QB.n4 GNDA 0.265156f
C52 QB.n5 GNDA 0.226459f
C53 VDDA.n20 GNDA 0.035733f
C54 VDDA.n47 GNDA 0.032081f
C55 VDDA.t36 GNDA 0.087042f
C56 VDDA.n62 GNDA 0.071466f
C57 VDDA.t2 GNDA 0.094372f
C58 VDDA.t12 GNDA 0.083377f
C59 VDDA.t3 GNDA 0.024738f
C60 VDDA.t33 GNDA 0.024738f
C61 VDDA.n77 GNDA 0.035733f
C62 VDDA.n85 GNDA 0.035733f
C63 VDDA.t6 GNDA 0.024738f
C64 VDDA.t39 GNDA 0.024738f
C65 VDDA.n93 GNDA 0.050393f
C66 VDDA.n111 GNDA 0.07788f
C67 VDDA.t8 GNDA 0.071466f
C68 VDDA.n120 GNDA 0.071466f
C69 VDDA.t27 GNDA 0.071466f
C70 VDDA.n134 GNDA 0.071466f
C71 VDDA.n141 GNDA 0.022763f
C72 VDDA.n181 GNDA 0.035733f
C73 VDDA.t30 GNDA 0.022906f
C74 VDDA.t10 GNDA 0.02199f
C75 VDDA.t0 GNDA 0.024738f
C76 VDDA.n200 GNDA 0.054058f
C77 VDDA.t14 GNDA 0.044895f
C78 VDDA.t5 GNDA 0.095288f
C79 VDDA.t18 GNDA 0.095288f
C80 VDDA.t20 GNDA 0.044895f
C81 VDDA.n224 GNDA 0.049476f
C82 VDDA.t16 GNDA 0.044895f
C83 VDDA.t26 GNDA 0.095288f
C84 VDDA.t19 GNDA 0.095288f
C85 VDDA.t23 GNDA 0.044895f
C86 VDDA.n240 GNDA 0.050393f
C87 VDDA.n246 GNDA 0.04856f
.ends

