magic
tech sky130A
timestamp 1739812843
<< nwell >>
rect 3005 1875 4725 2070
rect 3005 900 4645 1875
rect 2340 610 3055 900
rect 3265 640 3325 655
<< poly >>
rect 2645 2790 3005 2800
rect 2645 2770 2655 2790
rect 2675 2785 3005 2790
rect 2675 2770 2685 2785
rect 2645 2760 2685 2770
rect -130 960 -90 975
rect 2180 945 2220 955
rect 2180 930 2190 945
rect 2090 925 2190 930
rect 2210 925 2220 945
rect 2090 915 2220 925
rect 3030 650 3070 660
rect 3030 630 3040 650
rect 3060 640 3070 650
rect 3265 640 3325 655
rect 3060 630 3325 640
rect 3030 620 3325 630
rect 4025 640 4065 650
rect 4025 620 4035 640
rect 4055 620 4065 640
rect 4025 610 4065 620
rect 4245 455 4285 465
rect 4245 435 4255 455
rect 4275 435 4285 455
rect 4245 425 4285 435
rect -130 245 -90 260
rect 2075 85 2115 95
rect 2075 65 2085 85
rect 2105 65 2115 85
rect 2075 55 2115 65
<< polycont >>
rect 2655 2770 2675 2790
rect 2190 925 2210 945
rect 3040 630 3060 650
rect 4035 620 4055 640
rect 4255 435 4275 455
rect 2085 65 2105 85
<< locali >>
rect 2865 3045 2915 3060
rect 2865 3025 2880 3045
rect 2900 3025 2915 3045
rect 2865 3010 2915 3025
rect 2705 2810 2745 2820
rect 2645 2790 2685 2800
rect 2645 2770 2655 2790
rect 2675 2770 2685 2790
rect 2645 1575 2685 2770
rect 2645 1555 2655 1575
rect 2675 1555 2685 1575
rect 2645 1545 2685 1555
rect 2705 2790 2715 2810
rect 2735 2790 2745 2810
rect 2380 1210 2430 1220
rect 2355 1190 2390 1210
rect 2380 1180 2390 1190
rect 2420 1180 2430 1210
rect 2380 1170 2430 1180
rect 2040 1130 2680 1150
rect 2040 1105 2060 1130
rect 2180 945 2220 955
rect 2180 925 2190 945
rect 2210 925 2220 945
rect 2180 915 2220 925
rect 2300 945 2340 955
rect 2300 925 2310 945
rect 2330 925 2340 945
rect 2300 915 2340 925
rect 2660 660 2680 1130
rect 2640 650 2680 660
rect 2500 625 2550 640
rect 2500 620 2515 625
rect 2370 600 2400 620
rect 2420 600 2450 620
rect 2470 605 2515 620
rect 2535 605 2550 625
rect 2640 630 2650 650
rect 2670 630 2680 650
rect 2640 620 2680 630
rect 2470 600 2550 605
rect 2500 590 2550 600
rect 2705 585 2745 2790
rect 4910 2755 5950 2775
rect 2865 2450 2915 2465
rect 2865 2430 2880 2450
rect 2900 2430 2915 2450
rect 2865 2415 2915 2430
rect 5930 1625 5950 2755
rect 2785 1605 5950 1625
rect 2785 660 2805 1605
rect 2910 975 2960 990
rect 2910 955 2925 975
rect 2945 955 2960 975
rect 2910 940 2960 955
rect 2765 650 2805 660
rect 2765 630 2775 650
rect 2795 640 2805 650
rect 3030 650 3070 660
rect 3030 640 3040 650
rect 2795 630 3040 640
rect 3060 630 3070 650
rect 2765 620 3070 630
rect 4025 640 4065 650
rect 3330 585 3370 625
rect 4025 620 4035 640
rect 4055 620 4065 640
rect 4025 610 4065 620
rect 2040 540 2200 560
rect 2705 545 3370 585
rect 4625 555 4665 565
rect 2040 505 2060 540
rect 2180 520 2200 540
rect 4625 535 4635 555
rect 4655 535 4665 555
rect 4625 525 4665 535
rect 2180 500 2900 520
rect 2650 455 2690 465
rect 2650 435 2660 455
rect 2680 435 2690 455
rect 2650 425 2690 435
rect 4245 455 4285 465
rect 4245 435 4255 455
rect 4275 435 4285 455
rect 4245 425 4285 435
rect 2650 265 2670 425
rect 2320 245 2670 265
rect 2910 135 2960 150
rect 2910 115 2925 135
rect 2945 115 2960 135
rect 2910 100 2960 115
rect 2075 85 2115 95
rect 2075 65 2085 85
rect 2105 65 2115 85
rect 2075 55 2115 65
rect 2380 40 2430 50
rect 2380 30 2390 40
rect 2355 10 2390 30
rect 2420 10 2430 40
rect 2380 0 2430 10
rect 2380 -125 2430 -115
rect 2380 -155 2390 -125
rect 2420 -135 2430 -125
rect 7080 -135 7130 -105
rect 2420 -155 2460 -135
rect 2480 -155 2510 -135
rect 2530 -155 2560 -135
rect 2580 -155 2610 -135
rect 2630 -155 2660 -135
rect 2680 -155 2710 -135
rect 2730 -155 2760 -135
rect 2780 -155 2810 -135
rect 2830 -155 2860 -135
rect 2880 -155 2910 -135
rect 2930 -155 2960 -135
rect 2980 -155 3010 -135
rect 3030 -155 3060 -135
rect 3080 -155 3110 -135
rect 3130 -155 3160 -135
rect 3180 -155 3210 -135
rect 3230 -155 3260 -135
rect 3280 -155 3310 -135
rect 3330 -155 3360 -135
rect 3380 -155 3410 -135
rect 3430 -155 3460 -135
rect 3480 -155 3510 -135
rect 3530 -155 3560 -135
rect 3580 -155 3610 -135
rect 3630 -155 3660 -135
rect 3680 -155 3710 -135
rect 3730 -155 3760 -135
rect 3780 -155 3810 -135
rect 3830 -155 3860 -135
rect 3880 -155 3910 -135
rect 3930 -155 3960 -135
rect 3980 -155 4010 -135
rect 4030 -155 4060 -135
rect 4080 -155 4110 -135
rect 4130 -155 4160 -135
rect 4180 -155 4210 -135
rect 4230 -155 4260 -135
rect 4280 -155 4310 -135
rect 4330 -155 4360 -135
rect 4380 -155 4410 -135
rect 4430 -155 4460 -135
rect 4480 -155 4510 -135
rect 4530 -155 4560 -135
rect 4580 -155 4610 -135
rect 4630 -155 4660 -135
rect 4680 -155 4710 -135
rect 4730 -155 4760 -135
rect 4780 -155 4810 -135
rect 4830 -155 4860 -135
rect 4880 -155 4910 -135
rect 4930 -155 4960 -135
rect 4980 -155 5010 -135
rect 5030 -155 5060 -135
rect 5080 -155 5110 -135
rect 5130 -155 5160 -135
rect 5180 -155 5210 -135
rect 5230 -155 5260 -135
rect 5280 -155 5310 -135
rect 5330 -155 5360 -135
rect 5380 -155 5410 -135
rect 5430 -155 5460 -135
rect 5480 -155 5510 -135
rect 5530 -155 5560 -135
rect 5580 -155 5610 -135
rect 5630 -155 5660 -135
rect 5680 -155 5710 -135
rect 5730 -155 5760 -135
rect 5780 -155 5810 -135
rect 5830 -155 5860 -135
rect 5880 -155 5910 -135
rect 5930 -155 5960 -135
rect 5980 -155 6010 -135
rect 6030 -155 6060 -135
rect 6080 -155 6110 -135
rect 6130 -155 6160 -135
rect 6180 -155 6210 -135
rect 6230 -155 6260 -135
rect 6280 -155 6310 -135
rect 6330 -155 6360 -135
rect 6380 -155 6410 -135
rect 6430 -155 6460 -135
rect 6480 -155 6510 -135
rect 6530 -155 6560 -135
rect 6580 -155 6610 -135
rect 6630 -155 6660 -135
rect 6680 -155 6710 -135
rect 6730 -155 6760 -135
rect 6780 -155 6810 -135
rect 6830 -155 6860 -135
rect 6880 -155 6910 -135
rect 6930 -155 6960 -135
rect 6980 -155 7010 -135
rect 7030 -155 7060 -135
rect 7080 -155 7100 -135
rect 7120 -155 7130 -135
rect 2380 -165 2430 -155
<< viali >>
rect 2880 3025 2900 3045
rect 2655 1555 2675 1575
rect 2715 2790 2735 2810
rect 2390 1180 2420 1210
rect 2190 925 2210 945
rect 2310 925 2330 945
rect 2350 600 2370 620
rect 2400 600 2420 620
rect 2450 600 2470 620
rect 2515 605 2535 625
rect 2650 630 2670 650
rect 2880 2430 2900 2450
rect 2925 955 2945 975
rect 2775 630 2795 650
rect 4035 620 4055 640
rect 4635 535 4655 555
rect 2660 435 2680 455
rect 4255 435 4275 455
rect 2925 115 2945 135
rect 2085 65 2105 85
rect 2390 10 2420 40
rect 2390 -155 2420 -125
rect 2460 -155 2480 -135
rect 2510 -155 2530 -135
rect 2560 -155 2580 -135
rect 2610 -155 2630 -135
rect 2660 -155 2680 -135
rect 2710 -155 2730 -135
rect 2760 -155 2780 -135
rect 2810 -155 2830 -135
rect 2860 -155 2880 -135
rect 2910 -155 2930 -135
rect 2960 -155 2980 -135
rect 3010 -155 3030 -135
rect 3060 -155 3080 -135
rect 3110 -155 3130 -135
rect 3160 -155 3180 -135
rect 3210 -155 3230 -135
rect 3260 -155 3280 -135
rect 3310 -155 3330 -135
rect 3360 -155 3380 -135
rect 3410 -155 3430 -135
rect 3460 -155 3480 -135
rect 3510 -155 3530 -135
rect 3560 -155 3580 -135
rect 3610 -155 3630 -135
rect 3660 -155 3680 -135
rect 3710 -155 3730 -135
rect 3760 -155 3780 -135
rect 3810 -155 3830 -135
rect 3860 -155 3880 -135
rect 3910 -155 3930 -135
rect 3960 -155 3980 -135
rect 4010 -155 4030 -135
rect 4060 -155 4080 -135
rect 4110 -155 4130 -135
rect 4160 -155 4180 -135
rect 4210 -155 4230 -135
rect 4260 -155 4280 -135
rect 4310 -155 4330 -135
rect 4360 -155 4380 -135
rect 4410 -155 4430 -135
rect 4460 -155 4480 -135
rect 4510 -155 4530 -135
rect 4560 -155 4580 -135
rect 4610 -155 4630 -135
rect 4660 -155 4680 -135
rect 4710 -155 4730 -135
rect 4760 -155 4780 -135
rect 4810 -155 4830 -135
rect 4860 -155 4880 -135
rect 4910 -155 4930 -135
rect 4960 -155 4980 -135
rect 5010 -155 5030 -135
rect 5060 -155 5080 -135
rect 5110 -155 5130 -135
rect 5160 -155 5180 -135
rect 5210 -155 5230 -135
rect 5260 -155 5280 -135
rect 5310 -155 5330 -135
rect 5360 -155 5380 -135
rect 5410 -155 5430 -135
rect 5460 -155 5480 -135
rect 5510 -155 5530 -135
rect 5560 -155 5580 -135
rect 5610 -155 5630 -135
rect 5660 -155 5680 -135
rect 5710 -155 5730 -135
rect 5760 -155 5780 -135
rect 5810 -155 5830 -135
rect 5860 -155 5880 -135
rect 5910 -155 5930 -135
rect 5960 -155 5980 -135
rect 6010 -155 6030 -135
rect 6060 -155 6080 -135
rect 6110 -155 6130 -135
rect 6160 -155 6180 -135
rect 6210 -155 6230 -135
rect 6260 -155 6280 -135
rect 6310 -155 6330 -135
rect 6360 -155 6380 -135
rect 6410 -155 6430 -135
rect 6460 -155 6480 -135
rect 6510 -155 6530 -135
rect 6560 -155 6580 -135
rect 6610 -155 6630 -135
rect 6660 -155 6680 -135
rect 6710 -155 6730 -135
rect 6760 -155 6780 -135
rect 6810 -155 6830 -135
rect 6860 -155 6880 -135
rect 6910 -155 6930 -135
rect 6960 -155 6980 -135
rect 7010 -155 7030 -135
rect 7060 -155 7080 -135
rect 7100 -155 7120 -135
<< metal1 >>
rect 2865 3050 2915 3060
rect 2865 3020 2875 3050
rect 2905 3020 2915 3050
rect 2865 3010 2915 3020
rect 2705 2810 3005 2820
rect 2705 2790 2715 2810
rect 2735 2805 3005 2810
rect 2735 2790 2745 2805
rect 2705 2780 2745 2790
rect 2865 2455 2915 2465
rect 2865 2425 2875 2455
rect 2905 2425 2915 2455
rect 2865 2415 2915 2425
rect 2645 1575 5650 1585
rect 2645 1555 2655 1575
rect 2675 1555 5650 1575
rect 2645 1545 5650 1555
rect 2520 1445 2910 1500
rect 2355 1210 2430 1220
rect 2355 1180 2390 1210
rect 2420 1180 2430 1210
rect 2380 1170 2430 1180
rect 2520 1020 2565 1445
rect 2180 980 2565 1020
rect 2910 980 2960 990
rect 2180 945 2220 980
rect 2180 925 2190 945
rect 2210 925 2220 945
rect 2180 915 2220 925
rect 2300 945 2340 955
rect 2300 925 2310 945
rect 2330 935 2340 945
rect 2910 950 2920 980
rect 2950 950 2960 980
rect 2910 940 2960 950
rect 2330 925 2595 935
rect 2300 915 2595 925
rect 2500 630 2550 640
rect -140 590 -115 630
rect 2355 620 2510 630
rect 2370 600 2400 620
rect 2420 600 2450 620
rect 2470 600 2510 620
rect 2540 600 2550 630
rect 2355 590 2550 600
rect 2575 605 2595 915
rect 2640 650 2680 660
rect 2640 630 2650 650
rect 2670 640 2680 650
rect 2765 650 2805 660
rect 2765 640 2775 650
rect 2670 630 2775 640
rect 2795 630 2805 650
rect 2640 620 2805 630
rect 4025 640 4065 650
rect 4025 620 4035 640
rect 4055 620 4065 640
rect 4025 605 4065 620
rect 2575 585 4065 605
rect 5610 565 5650 1545
rect 4625 555 5650 565
rect 4625 535 4635 555
rect 4655 535 5650 555
rect 4625 525 5650 535
rect 2650 455 4285 465
rect 2650 435 2660 455
rect 2680 445 4255 455
rect 2680 435 2690 445
rect 2650 425 2690 435
rect 4245 435 4255 445
rect 4275 435 4285 455
rect 4245 425 4285 435
rect 2910 140 2960 150
rect 2910 110 2920 140
rect 2950 110 2960 140
rect 2910 100 2960 110
rect 2075 85 2775 95
rect 2075 65 2085 85
rect 2105 75 2775 85
rect 2105 65 2115 75
rect 2075 55 2115 65
rect 2380 40 2430 50
rect 2355 10 2390 40
rect 2420 10 2430 40
rect 2355 0 2430 10
rect 2735 5 2775 75
rect 5610 65 5650 525
rect 2735 -50 2910 5
rect 2380 -125 2430 -115
rect 2380 -155 2390 -125
rect 2420 -135 7130 -125
rect 2420 -155 2460 -135
rect 2480 -155 2510 -135
rect 2530 -155 2560 -135
rect 2580 -155 2610 -135
rect 2630 -155 2660 -135
rect 2680 -155 2710 -135
rect 2730 -155 2760 -135
rect 2780 -155 2810 -135
rect 2830 -155 2860 -135
rect 2880 -155 2910 -135
rect 2930 -155 2960 -135
rect 2980 -155 3010 -135
rect 3030 -155 3060 -135
rect 3080 -155 3110 -135
rect 3130 -155 3160 -135
rect 3180 -155 3210 -135
rect 3230 -155 3260 -135
rect 3280 -155 3310 -135
rect 3330 -155 3360 -135
rect 3380 -155 3410 -135
rect 3430 -155 3460 -135
rect 3480 -155 3510 -135
rect 3530 -155 3560 -135
rect 3580 -155 3610 -135
rect 3630 -155 3660 -135
rect 3680 -155 3710 -135
rect 3730 -155 3760 -135
rect 3780 -155 3810 -135
rect 3830 -155 3860 -135
rect 3880 -155 3910 -135
rect 3930 -155 3960 -135
rect 3980 -155 4010 -135
rect 4030 -155 4060 -135
rect 4080 -155 4110 -135
rect 4130 -155 4160 -135
rect 4180 -155 4210 -135
rect 4230 -155 4260 -135
rect 4280 -155 4310 -135
rect 4330 -155 4360 -135
rect 4380 -155 4410 -135
rect 4430 -155 4460 -135
rect 4480 -155 4510 -135
rect 4530 -155 4560 -135
rect 4580 -155 4610 -135
rect 4630 -155 4660 -135
rect 4680 -155 4710 -135
rect 4730 -155 4760 -135
rect 4780 -155 4810 -135
rect 4830 -155 4860 -135
rect 4880 -155 4910 -135
rect 4930 -155 4960 -135
rect 4980 -155 5010 -135
rect 5030 -155 5060 -135
rect 5080 -155 5110 -135
rect 5130 -155 5160 -135
rect 5180 -155 5210 -135
rect 5230 -155 5260 -135
rect 5280 -155 5310 -135
rect 5330 -155 5360 -135
rect 5380 -155 5410 -135
rect 5430 -155 5460 -135
rect 5480 -155 5510 -135
rect 5530 -155 5560 -135
rect 5580 -155 5610 -135
rect 5630 -155 5660 -135
rect 5680 -155 5710 -135
rect 5730 -155 5760 -135
rect 5780 -155 5810 -135
rect 5830 -155 5860 -135
rect 5880 -155 5910 -135
rect 5930 -155 5960 -135
rect 5980 -155 6010 -135
rect 6030 -155 6060 -135
rect 6080 -155 6110 -135
rect 6130 -155 6160 -135
rect 6180 -155 6210 -135
rect 6230 -155 6260 -135
rect 6280 -155 6310 -135
rect 6330 -155 6360 -135
rect 6380 -155 6410 -135
rect 6430 -155 6460 -135
rect 6480 -155 6510 -135
rect 6530 -155 6560 -135
rect 6580 -155 6610 -135
rect 6630 -155 6660 -135
rect 6680 -155 6710 -135
rect 6730 -155 6760 -135
rect 6780 -155 6810 -135
rect 6830 -155 6860 -135
rect 6880 -155 6910 -135
rect 6930 -155 6960 -135
rect 6980 -155 7010 -135
rect 7030 -155 7060 -135
rect 7080 -155 7100 -135
rect 7120 -155 7130 -135
rect 2380 -165 7130 -155
<< via1 >>
rect 2875 3045 2905 3050
rect 2875 3025 2880 3045
rect 2880 3025 2900 3045
rect 2900 3025 2905 3045
rect 2875 3020 2905 3025
rect 2875 2450 2905 2455
rect 2875 2430 2880 2450
rect 2880 2430 2900 2450
rect 2900 2430 2905 2450
rect 2875 2425 2905 2430
rect 2390 1180 2420 1210
rect 2920 975 2950 980
rect 2920 955 2925 975
rect 2925 955 2945 975
rect 2945 955 2950 975
rect 2920 950 2950 955
rect 2510 625 2540 630
rect 2510 605 2515 625
rect 2515 605 2535 625
rect 2535 605 2540 625
rect 2510 600 2540 605
rect 2920 135 2950 140
rect 2920 115 2925 135
rect 2925 115 2945 135
rect 2945 115 2950 135
rect 2920 110 2950 115
rect 2390 10 2420 40
rect 2390 -155 2420 -125
<< metal2 >>
rect 2865 3050 2915 3060
rect 2865 3020 2875 3050
rect 2905 3020 2915 3050
rect 2865 3010 2915 3020
rect 2865 2455 2915 2465
rect 2865 2425 2875 2455
rect 2905 2425 2915 2455
rect 2865 2415 2915 2425
rect 2380 1210 2430 1220
rect 2380 1180 2390 1210
rect 2420 1180 2430 1210
rect 2380 1170 2430 1180
rect 2910 980 2960 990
rect 2910 950 2920 980
rect 2950 950 2960 980
rect 2910 940 2960 950
rect 2500 630 2550 640
rect 2500 600 2510 630
rect 2540 600 2550 630
rect 2500 590 2550 600
rect 2910 140 2960 150
rect 2910 110 2920 140
rect 2950 110 2960 140
rect 2910 100 2960 110
rect 2380 40 2430 50
rect 2380 10 2390 40
rect 2420 10 2430 40
rect 2380 0 2430 10
rect 2380 -125 2430 -115
rect 2380 -155 2390 -125
rect 2420 -155 2430 -125
rect 2380 -165 2430 -155
<< via2 >>
rect 2875 3020 2905 3050
rect 2875 2425 2905 2455
rect 2390 1180 2420 1210
rect 2920 950 2950 980
rect 2510 600 2540 630
rect 2920 110 2950 140
rect 2390 10 2420 40
rect 2390 -155 2420 -125
<< metal3 >>
rect 2380 3055 2915 3060
rect 2380 3015 2385 3055
rect 2425 3050 2915 3055
rect 2425 3020 2875 3050
rect 2905 3020 2915 3050
rect 2425 3015 2915 3020
rect 2380 3010 2915 3015
rect 2500 2460 2915 2465
rect 2500 2420 2505 2460
rect 2545 2455 2915 2460
rect 2545 2425 2875 2455
rect 2905 2425 2915 2455
rect 2545 2420 2915 2425
rect 2500 2415 2915 2420
rect 2380 1215 2430 1220
rect 2380 1175 2385 1215
rect 2425 1175 2430 1215
rect 2380 1170 2430 1175
rect 2500 985 2960 990
rect 2500 945 2505 985
rect 2545 980 2960 985
rect 2545 950 2920 980
rect 2950 950 2960 980
rect 2545 945 2960 950
rect 2500 940 2960 945
rect 2500 635 2550 640
rect 2500 595 2505 635
rect 2545 595 2550 635
rect 2500 590 2550 595
rect 2380 145 2960 150
rect 2380 105 2385 145
rect 2425 140 2960 145
rect 2425 110 2920 140
rect 2950 110 2960 140
rect 2425 105 2960 110
rect 2380 100 2960 105
rect 2380 45 2430 50
rect 2380 5 2385 45
rect 2425 5 2430 45
rect 2380 0 2430 5
rect 2380 -120 2430 -115
rect 2380 -160 2385 -120
rect 2425 -160 2430 -120
rect 2380 -165 2430 -160
<< via3 >>
rect 2385 3015 2425 3055
rect 2505 2420 2545 2460
rect 2385 1210 2425 1215
rect 2385 1180 2390 1210
rect 2390 1180 2420 1210
rect 2420 1180 2425 1210
rect 2385 1175 2425 1180
rect 2505 945 2545 985
rect 2505 630 2545 635
rect 2505 600 2510 630
rect 2510 600 2540 630
rect 2540 600 2545 630
rect 2505 595 2545 600
rect 2385 105 2425 145
rect 2385 40 2425 45
rect 2385 10 2390 40
rect 2390 10 2420 40
rect 2420 10 2425 40
rect 2385 5 2425 10
rect 2385 -125 2425 -120
rect 2385 -155 2390 -125
rect 2390 -155 2420 -125
rect 2420 -155 2425 -125
rect 2385 -160 2425 -155
<< metal4 >>
rect 2380 3055 2430 3060
rect 2380 3015 2385 3055
rect 2425 3015 2430 3055
rect 2380 1215 2430 3015
rect 2380 1175 2385 1215
rect 2425 1175 2430 1215
rect -280 105 -230 155
rect 2380 145 2430 1175
rect 2500 2460 2550 2465
rect 2500 2420 2505 2460
rect 2545 2420 2550 2460
rect 2500 985 2550 2420
rect 2500 945 2505 985
rect 2545 945 2550 985
rect 2500 635 2550 945
rect 2500 595 2505 635
rect 2545 595 2550 635
rect 2500 590 2550 595
rect 2380 105 2385 145
rect 2425 105 2430 145
rect 2380 45 2430 105
rect 2380 5 2385 45
rect 2425 5 2430 45
rect 2380 -120 2430 5
rect 2380 -160 2385 -120
rect 2425 -160 2430 -120
rect 2380 -165 2430 -160
use charge_pump_cell_6  charge_pump_cell_6_0
timestamp 1739811829
transform 1 0 -6195 0 1 -1605
box 9095 1555 11620 3105
use loop_filter_2  loop_filter_2_0
timestamp 1739812747
transform 1 0 4475 0 1 -265
box 1135 -5975 9720 330
use opamp_cell_4  opamp_cell_4_0
timestamp 1739772381
transform 1 0 -335 0 -1 4855
box 3110 897 6365 3205
use pfd_8  pfd_8_0
timestamp 1739770731
transform 1 0 -930 0 1 4655
box 650 -4655 3290 -3435
<< labels >>
flabel locali 2880 510 2880 510 5 FreeSans 400 0 0 -200 I_IN
port 6 s
flabel metal1 -140 610 -140 610 7 FreeSans 400 0 -200 0 VDDA
port 2 w
flabel metal4 -280 130 -280 130 7 FreeSans 400 0 -200 0 GNDA
port 3 w
flabel poly -130 250 -130 250 7 FreeSans 400 0 -200 0 F_VCO
port 5 w
flabel poly -130 965 -130 965 7 FreeSans 400 0 -200 0 F_REF
port 4 w
flabel metal1 5650 545 5650 545 3 FreeSans 400 0 200 0 V_OUT
port 1 e
<< end >>
