magic
tech sky130A
magscale 1 2
timestamp 1748919360
<< xpolycontact >>
rect -69 64 69 496
rect -69 -496 69 -64
<< xpolyres >>
rect -69 -64 69 64
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.69 l 0.8 m 1 nx 1 wmin 0.690 lmin 0.50 class resistor rho 2000 val 2.864k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 0 glc 0 grc 0 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 0 n_guard 0 hv_guard 0 vias 0 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
