magic
tech sky130A
timestamp 1740145811
<< nwell >>
rect 3340 2185 5060 2840
rect 4265 2175 4640 2185
<< nmos >>
rect 3460 1925 3475 1975
rect 3525 1925 3540 1975
rect 3590 1925 3605 1975
rect 3655 1925 3670 1975
rect 3720 1925 3735 1975
rect 3785 1925 3800 1975
rect 4030 1925 4045 1975
rect 4095 1925 4110 1975
rect 4160 1925 4175 1975
rect 4225 1925 4240 1975
rect 4290 1925 4305 1975
rect 4355 1925 4370 1975
rect 4600 1925 4615 1975
rect 4665 1925 4680 1975
rect 4730 1925 4745 1975
rect 4795 1925 4810 1975
rect 4860 1925 4875 1975
rect 4925 1925 4940 1975
rect 3435 1580 3485 1705
rect 3535 1580 3585 1705
rect 3635 1580 3685 1705
rect 3735 1580 3785 1705
rect 3835 1580 3885 1705
rect 3935 1580 3985 1705
rect 4035 1580 4085 1705
rect 4135 1580 4185 1705
rect 4235 1580 4285 1705
rect 4335 1580 4385 1705
<< pmos >>
rect 3495 2535 3545 2785
rect 3595 2535 3645 2785
rect 3695 2535 3745 2785
rect 3795 2535 3845 2785
rect 3895 2535 3945 2785
rect 3995 2535 4045 2785
rect 4095 2535 4145 2785
rect 4195 2535 4245 2785
rect 4295 2535 4345 2785
rect 4395 2535 4445 2785
rect 3460 2210 3475 2310
rect 3525 2210 3540 2310
rect 3590 2210 3605 2310
rect 3655 2210 3670 2310
rect 3720 2210 3735 2310
rect 3785 2210 3800 2310
rect 4030 2210 4045 2310
rect 4095 2210 4110 2310
rect 4160 2210 4175 2310
rect 4225 2210 4240 2310
rect 4290 2210 4305 2310
rect 4355 2210 4370 2310
rect 4600 2210 4615 2310
rect 4665 2210 4680 2310
rect 4730 2210 4745 2310
rect 4795 2210 4810 2310
rect 4860 2210 4875 2310
rect 4925 2210 4940 2310
<< ndiff >>
rect 3410 1960 3460 1975
rect 3410 1940 3425 1960
rect 3445 1940 3460 1960
rect 3410 1925 3460 1940
rect 3475 1960 3525 1975
rect 3475 1940 3490 1960
rect 3510 1940 3525 1960
rect 3475 1925 3525 1940
rect 3540 1960 3590 1975
rect 3540 1940 3555 1960
rect 3575 1940 3590 1960
rect 3540 1925 3590 1940
rect 3605 1960 3655 1975
rect 3605 1940 3620 1960
rect 3640 1940 3655 1960
rect 3605 1925 3655 1940
rect 3670 1960 3720 1975
rect 3670 1940 3685 1960
rect 3705 1940 3720 1960
rect 3670 1925 3720 1940
rect 3735 1960 3785 1975
rect 3735 1940 3750 1960
rect 3770 1940 3785 1960
rect 3735 1925 3785 1940
rect 3800 1960 3850 1975
rect 3800 1940 3815 1960
rect 3835 1940 3850 1960
rect 3800 1925 3850 1940
rect 3980 1960 4030 1975
rect 3980 1940 3995 1960
rect 4015 1940 4030 1960
rect 3980 1925 4030 1940
rect 4045 1960 4095 1975
rect 4045 1940 4060 1960
rect 4080 1940 4095 1960
rect 4045 1925 4095 1940
rect 4110 1960 4160 1975
rect 4110 1940 4125 1960
rect 4145 1940 4160 1960
rect 4110 1925 4160 1940
rect 4175 1960 4225 1975
rect 4175 1940 4190 1960
rect 4210 1940 4225 1960
rect 4175 1925 4225 1940
rect 4240 1960 4290 1975
rect 4240 1940 4255 1960
rect 4275 1940 4290 1960
rect 4240 1925 4290 1940
rect 4305 1960 4355 1975
rect 4305 1940 4320 1960
rect 4340 1940 4355 1960
rect 4305 1925 4355 1940
rect 4370 1960 4420 1975
rect 4370 1940 4385 1960
rect 4405 1940 4420 1960
rect 4370 1925 4420 1940
rect 4550 1960 4600 1975
rect 4550 1940 4565 1960
rect 4585 1940 4600 1960
rect 4550 1925 4600 1940
rect 4615 1960 4665 1975
rect 4615 1940 4630 1960
rect 4650 1940 4665 1960
rect 4615 1925 4665 1940
rect 4680 1960 4730 1975
rect 4680 1940 4695 1960
rect 4715 1940 4730 1960
rect 4680 1925 4730 1940
rect 4745 1960 4795 1975
rect 4745 1940 4760 1960
rect 4780 1940 4795 1960
rect 4745 1925 4795 1940
rect 4810 1960 4860 1975
rect 4810 1940 4825 1960
rect 4845 1940 4860 1960
rect 4810 1925 4860 1940
rect 4875 1960 4925 1975
rect 4875 1940 4890 1960
rect 4910 1940 4925 1960
rect 4875 1925 4925 1940
rect 4940 1960 4990 1975
rect 4940 1940 4955 1960
rect 4975 1940 4990 1960
rect 4940 1925 4990 1940
rect 3385 1690 3435 1705
rect 3385 1665 3400 1690
rect 3420 1665 3435 1690
rect 3385 1620 3435 1665
rect 3385 1595 3400 1620
rect 3420 1595 3435 1620
rect 3385 1580 3435 1595
rect 3485 1690 3535 1705
rect 3485 1665 3500 1690
rect 3520 1665 3535 1690
rect 3485 1620 3535 1665
rect 3485 1595 3500 1620
rect 3520 1595 3535 1620
rect 3485 1580 3535 1595
rect 3585 1690 3635 1705
rect 3585 1665 3600 1690
rect 3620 1665 3635 1690
rect 3585 1620 3635 1665
rect 3585 1595 3600 1620
rect 3620 1595 3635 1620
rect 3585 1580 3635 1595
rect 3685 1690 3735 1705
rect 3685 1665 3700 1690
rect 3720 1665 3735 1690
rect 3685 1620 3735 1665
rect 3685 1595 3700 1620
rect 3720 1595 3735 1620
rect 3685 1580 3735 1595
rect 3785 1690 3835 1705
rect 3785 1665 3800 1690
rect 3820 1665 3835 1690
rect 3785 1620 3835 1665
rect 3785 1595 3800 1620
rect 3820 1595 3835 1620
rect 3785 1580 3835 1595
rect 3885 1690 3935 1705
rect 3885 1665 3900 1690
rect 3920 1665 3935 1690
rect 3885 1620 3935 1665
rect 3885 1595 3900 1620
rect 3920 1595 3935 1620
rect 3885 1580 3935 1595
rect 3985 1690 4035 1705
rect 3985 1665 4000 1690
rect 4020 1665 4035 1690
rect 3985 1620 4035 1665
rect 3985 1595 4000 1620
rect 4020 1595 4035 1620
rect 3985 1580 4035 1595
rect 4085 1690 4135 1705
rect 4085 1665 4100 1690
rect 4120 1665 4135 1690
rect 4085 1620 4135 1665
rect 4085 1595 4100 1620
rect 4120 1595 4135 1620
rect 4085 1580 4135 1595
rect 4185 1690 4235 1705
rect 4185 1665 4200 1690
rect 4220 1665 4235 1690
rect 4185 1620 4235 1665
rect 4185 1595 4200 1620
rect 4220 1595 4235 1620
rect 4185 1580 4235 1595
rect 4285 1690 4335 1705
rect 4285 1665 4300 1690
rect 4320 1665 4335 1690
rect 4285 1620 4335 1665
rect 4285 1595 4300 1620
rect 4320 1595 4335 1620
rect 4285 1580 4335 1595
rect 4385 1690 4435 1705
rect 4385 1665 4400 1690
rect 4420 1665 4435 1690
rect 4385 1620 4435 1665
rect 4385 1595 4400 1620
rect 4420 1595 4435 1620
rect 4385 1580 4435 1595
<< pdiff >>
rect 3445 2770 3495 2785
rect 3445 2750 3460 2770
rect 3480 2750 3495 2770
rect 3445 2720 3495 2750
rect 3445 2700 3460 2720
rect 3480 2700 3495 2720
rect 3445 2670 3495 2700
rect 3445 2650 3460 2670
rect 3480 2650 3495 2670
rect 3445 2620 3495 2650
rect 3445 2600 3460 2620
rect 3480 2600 3495 2620
rect 3445 2570 3495 2600
rect 3445 2550 3460 2570
rect 3480 2550 3495 2570
rect 3445 2535 3495 2550
rect 3545 2770 3595 2785
rect 3545 2750 3560 2770
rect 3580 2750 3595 2770
rect 3545 2720 3595 2750
rect 3545 2700 3560 2720
rect 3580 2700 3595 2720
rect 3545 2670 3595 2700
rect 3545 2650 3560 2670
rect 3580 2650 3595 2670
rect 3545 2620 3595 2650
rect 3545 2600 3560 2620
rect 3580 2600 3595 2620
rect 3545 2570 3595 2600
rect 3545 2550 3560 2570
rect 3580 2550 3595 2570
rect 3545 2535 3595 2550
rect 3645 2770 3695 2785
rect 3645 2750 3660 2770
rect 3680 2750 3695 2770
rect 3645 2720 3695 2750
rect 3645 2700 3660 2720
rect 3680 2700 3695 2720
rect 3645 2670 3695 2700
rect 3645 2650 3660 2670
rect 3680 2650 3695 2670
rect 3645 2620 3695 2650
rect 3645 2600 3660 2620
rect 3680 2600 3695 2620
rect 3645 2570 3695 2600
rect 3645 2550 3660 2570
rect 3680 2550 3695 2570
rect 3645 2535 3695 2550
rect 3745 2770 3795 2785
rect 3745 2750 3760 2770
rect 3780 2750 3795 2770
rect 3745 2720 3795 2750
rect 3745 2700 3760 2720
rect 3780 2700 3795 2720
rect 3745 2670 3795 2700
rect 3745 2650 3760 2670
rect 3780 2650 3795 2670
rect 3745 2620 3795 2650
rect 3745 2600 3760 2620
rect 3780 2600 3795 2620
rect 3745 2570 3795 2600
rect 3745 2550 3760 2570
rect 3780 2550 3795 2570
rect 3745 2535 3795 2550
rect 3845 2770 3895 2785
rect 3845 2750 3860 2770
rect 3880 2750 3895 2770
rect 3845 2720 3895 2750
rect 3845 2700 3860 2720
rect 3880 2700 3895 2720
rect 3845 2670 3895 2700
rect 3845 2650 3860 2670
rect 3880 2650 3895 2670
rect 3845 2620 3895 2650
rect 3845 2600 3860 2620
rect 3880 2600 3895 2620
rect 3845 2570 3895 2600
rect 3845 2550 3860 2570
rect 3880 2550 3895 2570
rect 3845 2535 3895 2550
rect 3945 2770 3995 2785
rect 3945 2750 3960 2770
rect 3980 2750 3995 2770
rect 3945 2720 3995 2750
rect 3945 2700 3960 2720
rect 3980 2700 3995 2720
rect 3945 2670 3995 2700
rect 3945 2650 3960 2670
rect 3980 2650 3995 2670
rect 3945 2620 3995 2650
rect 3945 2600 3960 2620
rect 3980 2600 3995 2620
rect 3945 2570 3995 2600
rect 3945 2550 3960 2570
rect 3980 2550 3995 2570
rect 3945 2535 3995 2550
rect 4045 2770 4095 2785
rect 4045 2750 4060 2770
rect 4080 2750 4095 2770
rect 4045 2720 4095 2750
rect 4045 2700 4060 2720
rect 4080 2700 4095 2720
rect 4045 2670 4095 2700
rect 4045 2650 4060 2670
rect 4080 2650 4095 2670
rect 4045 2620 4095 2650
rect 4045 2600 4060 2620
rect 4080 2600 4095 2620
rect 4045 2570 4095 2600
rect 4045 2550 4060 2570
rect 4080 2550 4095 2570
rect 4045 2535 4095 2550
rect 4145 2770 4195 2785
rect 4145 2750 4160 2770
rect 4180 2750 4195 2770
rect 4145 2720 4195 2750
rect 4145 2700 4160 2720
rect 4180 2700 4195 2720
rect 4145 2670 4195 2700
rect 4145 2650 4160 2670
rect 4180 2650 4195 2670
rect 4145 2620 4195 2650
rect 4145 2600 4160 2620
rect 4180 2600 4195 2620
rect 4145 2570 4195 2600
rect 4145 2550 4160 2570
rect 4180 2550 4195 2570
rect 4145 2535 4195 2550
rect 4245 2770 4295 2785
rect 4245 2750 4260 2770
rect 4280 2750 4295 2770
rect 4245 2720 4295 2750
rect 4245 2700 4260 2720
rect 4280 2700 4295 2720
rect 4245 2670 4295 2700
rect 4245 2650 4260 2670
rect 4280 2650 4295 2670
rect 4245 2620 4295 2650
rect 4245 2600 4260 2620
rect 4280 2600 4295 2620
rect 4245 2570 4295 2600
rect 4245 2550 4260 2570
rect 4280 2550 4295 2570
rect 4245 2535 4295 2550
rect 4345 2770 4395 2785
rect 4345 2750 4360 2770
rect 4380 2750 4395 2770
rect 4345 2720 4395 2750
rect 4345 2700 4360 2720
rect 4380 2700 4395 2720
rect 4345 2670 4395 2700
rect 4345 2650 4360 2670
rect 4380 2650 4395 2670
rect 4345 2620 4395 2650
rect 4345 2600 4360 2620
rect 4380 2600 4395 2620
rect 4345 2570 4395 2600
rect 4345 2550 4360 2570
rect 4380 2550 4395 2570
rect 4345 2535 4395 2550
rect 4445 2770 4495 2785
rect 4445 2750 4460 2770
rect 4480 2750 4495 2770
rect 4445 2720 4495 2750
rect 4445 2700 4460 2720
rect 4480 2700 4495 2720
rect 4445 2670 4495 2700
rect 4445 2650 4460 2670
rect 4480 2650 4495 2670
rect 4445 2620 4495 2650
rect 4445 2600 4460 2620
rect 4480 2600 4495 2620
rect 4445 2570 4495 2600
rect 4445 2550 4460 2570
rect 4480 2550 4495 2570
rect 4445 2535 4495 2550
rect 3410 2295 3460 2310
rect 3410 2275 3425 2295
rect 3445 2275 3460 2295
rect 3410 2245 3460 2275
rect 3410 2225 3425 2245
rect 3445 2225 3460 2245
rect 3410 2210 3460 2225
rect 3475 2295 3525 2310
rect 3475 2275 3490 2295
rect 3510 2275 3525 2295
rect 3475 2245 3525 2275
rect 3475 2225 3490 2245
rect 3510 2225 3525 2245
rect 3475 2210 3525 2225
rect 3540 2295 3590 2310
rect 3540 2275 3555 2295
rect 3575 2275 3590 2295
rect 3540 2245 3590 2275
rect 3540 2225 3555 2245
rect 3575 2225 3590 2245
rect 3540 2210 3590 2225
rect 3605 2295 3655 2310
rect 3605 2275 3620 2295
rect 3640 2275 3655 2295
rect 3605 2245 3655 2275
rect 3605 2225 3620 2245
rect 3640 2225 3655 2245
rect 3605 2210 3655 2225
rect 3670 2295 3720 2310
rect 3670 2275 3685 2295
rect 3705 2275 3720 2295
rect 3670 2245 3720 2275
rect 3670 2225 3685 2245
rect 3705 2225 3720 2245
rect 3670 2210 3720 2225
rect 3735 2295 3785 2310
rect 3735 2275 3750 2295
rect 3770 2275 3785 2295
rect 3735 2245 3785 2275
rect 3735 2225 3750 2245
rect 3770 2225 3785 2245
rect 3735 2210 3785 2225
rect 3800 2295 3850 2310
rect 3800 2275 3815 2295
rect 3835 2275 3850 2295
rect 3800 2245 3850 2275
rect 3800 2225 3815 2245
rect 3835 2225 3850 2245
rect 3800 2210 3850 2225
rect 3980 2295 4030 2310
rect 3980 2275 3995 2295
rect 4015 2275 4030 2295
rect 3980 2245 4030 2275
rect 3980 2225 3995 2245
rect 4015 2225 4030 2245
rect 3980 2210 4030 2225
rect 4045 2295 4095 2310
rect 4045 2275 4060 2295
rect 4080 2275 4095 2295
rect 4045 2245 4095 2275
rect 4045 2225 4060 2245
rect 4080 2225 4095 2245
rect 4045 2210 4095 2225
rect 4110 2295 4160 2310
rect 4110 2275 4125 2295
rect 4145 2275 4160 2295
rect 4110 2245 4160 2275
rect 4110 2225 4125 2245
rect 4145 2225 4160 2245
rect 4110 2210 4160 2225
rect 4175 2295 4225 2310
rect 4175 2275 4190 2295
rect 4210 2275 4225 2295
rect 4175 2245 4225 2275
rect 4175 2225 4190 2245
rect 4210 2225 4225 2245
rect 4175 2210 4225 2225
rect 4240 2295 4290 2310
rect 4240 2275 4255 2295
rect 4275 2275 4290 2295
rect 4240 2245 4290 2275
rect 4240 2225 4255 2245
rect 4275 2225 4290 2245
rect 4240 2210 4290 2225
rect 4305 2295 4355 2310
rect 4305 2275 4320 2295
rect 4340 2275 4355 2295
rect 4305 2245 4355 2275
rect 4305 2225 4320 2245
rect 4340 2225 4355 2245
rect 4305 2210 4355 2225
rect 4370 2295 4420 2310
rect 4370 2275 4385 2295
rect 4405 2275 4420 2295
rect 4370 2245 4420 2275
rect 4370 2225 4385 2245
rect 4405 2225 4420 2245
rect 4370 2210 4420 2225
rect 4550 2295 4600 2310
rect 4550 2275 4565 2295
rect 4585 2275 4600 2295
rect 4550 2245 4600 2275
rect 4550 2225 4565 2245
rect 4585 2225 4600 2245
rect 4550 2210 4600 2225
rect 4615 2295 4665 2310
rect 4615 2275 4630 2295
rect 4650 2275 4665 2295
rect 4615 2245 4665 2275
rect 4615 2225 4630 2245
rect 4650 2225 4665 2245
rect 4615 2210 4665 2225
rect 4680 2295 4730 2310
rect 4680 2275 4695 2295
rect 4715 2275 4730 2295
rect 4680 2245 4730 2275
rect 4680 2225 4695 2245
rect 4715 2225 4730 2245
rect 4680 2210 4730 2225
rect 4745 2295 4795 2310
rect 4745 2275 4760 2295
rect 4780 2275 4795 2295
rect 4745 2245 4795 2275
rect 4745 2225 4760 2245
rect 4780 2225 4795 2245
rect 4745 2210 4795 2225
rect 4810 2295 4860 2310
rect 4810 2275 4825 2295
rect 4845 2275 4860 2295
rect 4810 2245 4860 2275
rect 4810 2225 4825 2245
rect 4845 2225 4860 2245
rect 4810 2210 4860 2225
rect 4875 2295 4925 2310
rect 4875 2275 4890 2295
rect 4910 2275 4925 2295
rect 4875 2245 4925 2275
rect 4875 2225 4890 2245
rect 4910 2225 4925 2245
rect 4875 2210 4925 2225
rect 4940 2295 4990 2310
rect 4940 2275 4955 2295
rect 4975 2275 4990 2295
rect 4940 2245 4990 2275
rect 4940 2225 4955 2245
rect 4975 2225 4990 2245
rect 4940 2210 4990 2225
<< ndiffc >>
rect 3425 1940 3445 1960
rect 3490 1940 3510 1960
rect 3555 1940 3575 1960
rect 3620 1940 3640 1960
rect 3685 1940 3705 1960
rect 3750 1940 3770 1960
rect 3815 1940 3835 1960
rect 3995 1940 4015 1960
rect 4060 1940 4080 1960
rect 4125 1940 4145 1960
rect 4190 1940 4210 1960
rect 4255 1940 4275 1960
rect 4320 1940 4340 1960
rect 4385 1940 4405 1960
rect 4565 1940 4585 1960
rect 4630 1940 4650 1960
rect 4695 1940 4715 1960
rect 4760 1940 4780 1960
rect 4825 1940 4845 1960
rect 4890 1940 4910 1960
rect 4955 1940 4975 1960
rect 3400 1665 3420 1690
rect 3400 1595 3420 1620
rect 3500 1665 3520 1690
rect 3500 1595 3520 1620
rect 3600 1665 3620 1690
rect 3600 1595 3620 1620
rect 3700 1665 3720 1690
rect 3700 1595 3720 1620
rect 3800 1665 3820 1690
rect 3800 1595 3820 1620
rect 3900 1665 3920 1690
rect 3900 1595 3920 1620
rect 4000 1665 4020 1690
rect 4000 1595 4020 1620
rect 4100 1665 4120 1690
rect 4100 1595 4120 1620
rect 4200 1665 4220 1690
rect 4200 1595 4220 1620
rect 4300 1665 4320 1690
rect 4300 1595 4320 1620
rect 4400 1665 4420 1690
rect 4400 1595 4420 1620
<< pdiffc >>
rect 3460 2750 3480 2770
rect 3460 2700 3480 2720
rect 3460 2650 3480 2670
rect 3460 2600 3480 2620
rect 3460 2550 3480 2570
rect 3560 2750 3580 2770
rect 3560 2700 3580 2720
rect 3560 2650 3580 2670
rect 3560 2600 3580 2620
rect 3560 2550 3580 2570
rect 3660 2750 3680 2770
rect 3660 2700 3680 2720
rect 3660 2650 3680 2670
rect 3660 2600 3680 2620
rect 3660 2550 3680 2570
rect 3760 2750 3780 2770
rect 3760 2700 3780 2720
rect 3760 2650 3780 2670
rect 3760 2600 3780 2620
rect 3760 2550 3780 2570
rect 3860 2750 3880 2770
rect 3860 2700 3880 2720
rect 3860 2650 3880 2670
rect 3860 2600 3880 2620
rect 3860 2550 3880 2570
rect 3960 2750 3980 2770
rect 3960 2700 3980 2720
rect 3960 2650 3980 2670
rect 3960 2600 3980 2620
rect 3960 2550 3980 2570
rect 4060 2750 4080 2770
rect 4060 2700 4080 2720
rect 4060 2650 4080 2670
rect 4060 2600 4080 2620
rect 4060 2550 4080 2570
rect 4160 2750 4180 2770
rect 4160 2700 4180 2720
rect 4160 2650 4180 2670
rect 4160 2600 4180 2620
rect 4160 2550 4180 2570
rect 4260 2750 4280 2770
rect 4260 2700 4280 2720
rect 4260 2650 4280 2670
rect 4260 2600 4280 2620
rect 4260 2550 4280 2570
rect 4360 2750 4380 2770
rect 4360 2700 4380 2720
rect 4360 2650 4380 2670
rect 4360 2600 4380 2620
rect 4360 2550 4380 2570
rect 4460 2750 4480 2770
rect 4460 2700 4480 2720
rect 4460 2650 4480 2670
rect 4460 2600 4480 2620
rect 4460 2550 4480 2570
rect 3425 2275 3445 2295
rect 3425 2225 3445 2245
rect 3490 2275 3510 2295
rect 3490 2225 3510 2245
rect 3555 2275 3575 2295
rect 3555 2225 3575 2245
rect 3620 2275 3640 2295
rect 3620 2225 3640 2245
rect 3685 2275 3705 2295
rect 3685 2225 3705 2245
rect 3750 2275 3770 2295
rect 3750 2225 3770 2245
rect 3815 2275 3835 2295
rect 3815 2225 3835 2245
rect 3995 2275 4015 2295
rect 3995 2225 4015 2245
rect 4060 2275 4080 2295
rect 4060 2225 4080 2245
rect 4125 2275 4145 2295
rect 4125 2225 4145 2245
rect 4190 2275 4210 2295
rect 4190 2225 4210 2245
rect 4255 2275 4275 2295
rect 4255 2225 4275 2245
rect 4320 2275 4340 2295
rect 4320 2225 4340 2245
rect 4385 2275 4405 2295
rect 4385 2225 4405 2245
rect 4565 2275 4585 2295
rect 4565 2225 4585 2245
rect 4630 2275 4650 2295
rect 4630 2225 4650 2245
rect 4695 2275 4715 2295
rect 4695 2225 4715 2245
rect 4760 2275 4780 2295
rect 4760 2225 4780 2245
rect 4825 2275 4845 2295
rect 4825 2225 4845 2245
rect 4890 2275 4910 2295
rect 4890 2225 4910 2245
rect 4955 2275 4975 2295
rect 4955 2225 4975 2245
<< psubdiff >>
rect 3360 1960 3410 1975
rect 3360 1940 3375 1960
rect 3395 1940 3410 1960
rect 3360 1925 3410 1940
rect 3850 1960 3900 1975
rect 3850 1940 3865 1960
rect 3885 1940 3900 1960
rect 3850 1925 3900 1940
rect 4500 1960 4550 1975
rect 4500 1940 4515 1960
rect 4535 1940 4550 1960
rect 4500 1925 4550 1940
rect 4990 1960 5040 1975
rect 4990 1940 5005 1960
rect 5025 1940 5040 1960
rect 4990 1925 5040 1940
rect 3335 1690 3385 1705
rect 3335 1665 3350 1690
rect 3370 1665 3385 1690
rect 3335 1620 3385 1665
rect 3335 1595 3350 1620
rect 3370 1595 3385 1620
rect 3335 1580 3385 1595
rect 4435 1690 4485 1705
rect 4435 1665 4450 1690
rect 4470 1665 4485 1690
rect 4435 1620 4485 1665
rect 4435 1595 4450 1620
rect 4470 1595 4485 1620
rect 4435 1580 4485 1595
<< nsubdiff >>
rect 3395 2770 3445 2785
rect 3395 2750 3410 2770
rect 3430 2750 3445 2770
rect 3395 2720 3445 2750
rect 3395 2700 3410 2720
rect 3430 2700 3445 2720
rect 3395 2670 3445 2700
rect 3395 2650 3410 2670
rect 3430 2650 3445 2670
rect 3395 2620 3445 2650
rect 3395 2600 3410 2620
rect 3430 2600 3445 2620
rect 3395 2570 3445 2600
rect 3395 2550 3410 2570
rect 3430 2550 3445 2570
rect 3395 2535 3445 2550
rect 4495 2770 4545 2785
rect 4495 2750 4510 2770
rect 4530 2750 4545 2770
rect 4495 2720 4545 2750
rect 4495 2700 4510 2720
rect 4530 2700 4545 2720
rect 4495 2670 4545 2700
rect 4495 2650 4510 2670
rect 4530 2650 4545 2670
rect 4495 2620 4545 2650
rect 4495 2600 4510 2620
rect 4530 2600 4545 2620
rect 4495 2570 4545 2600
rect 4495 2550 4510 2570
rect 4530 2550 4545 2570
rect 4495 2535 4545 2550
rect 3930 2295 3980 2310
rect 3930 2275 3945 2295
rect 3965 2275 3980 2295
rect 3930 2245 3980 2275
rect 3930 2225 3945 2245
rect 3965 2225 3980 2245
rect 3930 2210 3980 2225
rect 4420 2295 4470 2310
rect 4420 2275 4435 2295
rect 4455 2275 4470 2295
rect 4420 2245 4470 2275
rect 4420 2225 4435 2245
rect 4455 2225 4470 2245
rect 4420 2210 4470 2225
rect 4500 2295 4550 2310
rect 4500 2275 4515 2295
rect 4535 2275 4550 2295
rect 4500 2245 4550 2275
rect 4500 2225 4515 2245
rect 4535 2225 4550 2245
rect 4500 2210 4550 2225
rect 4990 2295 5040 2310
rect 4990 2275 5005 2295
rect 5025 2275 5040 2295
rect 4990 2245 5040 2275
rect 4990 2225 5005 2245
rect 5025 2225 5040 2245
rect 4990 2210 5040 2225
<< psubdiffcont >>
rect 3375 1940 3395 1960
rect 3865 1940 3885 1960
rect 4515 1940 4535 1960
rect 5005 1940 5025 1960
rect 3350 1665 3370 1690
rect 3350 1595 3370 1620
rect 4450 1665 4470 1690
rect 4450 1595 4470 1620
<< nsubdiffcont >>
rect 3410 2750 3430 2770
rect 3410 2700 3430 2720
rect 3410 2650 3430 2670
rect 3410 2600 3430 2620
rect 3410 2550 3430 2570
rect 4510 2750 4530 2770
rect 4510 2700 4530 2720
rect 4510 2650 4530 2670
rect 4510 2600 4530 2620
rect 4510 2550 4530 2570
rect 3945 2275 3965 2295
rect 3945 2225 3965 2245
rect 4435 2275 4455 2295
rect 4435 2225 4455 2245
rect 4515 2275 4535 2295
rect 4515 2225 4535 2245
rect 5005 2275 5025 2295
rect 5005 2225 5025 2245
<< poly >>
rect 3850 2830 3890 2840
rect 3850 2810 3860 2830
rect 3880 2810 3890 2830
rect 4050 2830 4090 2840
rect 4050 2810 4060 2830
rect 4080 2810 4090 2830
rect 3495 2785 3545 2800
rect 3595 2795 4345 2810
rect 3595 2785 3645 2795
rect 3695 2785 3745 2795
rect 3795 2785 3845 2795
rect 3895 2785 3945 2795
rect 3995 2785 4045 2795
rect 4095 2785 4145 2795
rect 4195 2785 4245 2795
rect 4295 2785 4345 2795
rect 4395 2785 4445 2800
rect 3495 2520 3545 2535
rect 3595 2520 3645 2535
rect 3695 2520 3745 2535
rect 3795 2520 3845 2535
rect 3895 2520 3945 2535
rect 3995 2520 4045 2535
rect 4095 2520 4145 2535
rect 4195 2520 4245 2535
rect 4295 2520 4345 2535
rect 4395 2520 4445 2535
rect 3450 2510 3545 2520
rect 3450 2490 3460 2510
rect 3480 2505 3545 2510
rect 4395 2510 4490 2520
rect 4395 2505 4460 2510
rect 3480 2490 3490 2505
rect 3450 2480 3490 2490
rect 4450 2490 4460 2505
rect 4480 2490 4490 2510
rect 4450 2480 4490 2490
rect 3445 2355 3485 2365
rect 3445 2335 3455 2355
rect 3475 2335 3485 2355
rect 3445 2325 3485 2335
rect 3775 2355 3815 2365
rect 3775 2335 3785 2355
rect 3805 2335 3815 2355
rect 3775 2325 3815 2335
rect 4015 2355 4055 2365
rect 4015 2335 4025 2355
rect 4045 2335 4055 2355
rect 4015 2325 4055 2335
rect 4345 2355 4385 2365
rect 4345 2335 4355 2355
rect 4375 2335 4385 2355
rect 4345 2325 4385 2335
rect 4585 2355 4625 2365
rect 4585 2335 4595 2355
rect 4615 2335 4625 2355
rect 4585 2325 4625 2335
rect 4915 2355 4955 2365
rect 4915 2335 4925 2355
rect 4945 2335 4955 2355
rect 4915 2325 4955 2335
rect 3460 2310 3475 2325
rect 3525 2310 3540 2325
rect 3590 2310 3605 2325
rect 3655 2310 3670 2325
rect 3720 2310 3735 2325
rect 3785 2310 3800 2325
rect 4030 2310 4045 2325
rect 4095 2310 4110 2325
rect 4160 2310 4175 2325
rect 4225 2310 4240 2325
rect 4290 2310 4305 2325
rect 4355 2310 4370 2325
rect 4600 2310 4615 2325
rect 4665 2310 4680 2325
rect 4730 2310 4745 2325
rect 4795 2310 4810 2325
rect 4860 2310 4875 2325
rect 4925 2310 4940 2325
rect 3460 2195 3475 2210
rect 3525 2200 3540 2210
rect 3590 2200 3605 2210
rect 3525 2195 3605 2200
rect 3500 2185 3605 2195
rect 3655 2200 3670 2210
rect 3720 2200 3735 2210
rect 3655 2195 3735 2200
rect 3785 2195 3800 2210
rect 4030 2195 4045 2210
rect 4095 2200 4110 2210
rect 4160 2200 4175 2210
rect 4225 2200 4240 2210
rect 4290 2200 4305 2210
rect 3655 2185 3760 2195
rect 4095 2185 4305 2200
rect 4355 2195 4370 2210
rect 4600 2195 4615 2210
rect 4665 2195 4680 2210
rect 3500 2165 3510 2185
rect 3530 2165 3540 2185
rect 3500 2155 3540 2165
rect 3720 2165 3730 2185
rect 3750 2165 3760 2185
rect 3720 2155 3760 2165
rect 4115 2180 4155 2185
rect 4115 2160 4125 2180
rect 4145 2160 4155 2180
rect 4265 2175 4305 2185
rect 4640 2185 4680 2195
rect 4115 2150 4155 2160
rect 4640 2165 4650 2185
rect 4670 2170 4680 2185
rect 4730 2170 4745 2210
rect 4795 2170 4810 2210
rect 4860 2170 4875 2210
rect 4925 2195 4940 2210
rect 5060 2185 5100 2195
rect 5060 2170 5070 2185
rect 4670 2165 5070 2170
rect 5090 2165 5100 2185
rect 4640 2155 5100 2165
rect 4640 2080 4680 2090
rect 4640 2060 4650 2080
rect 4670 2060 4680 2080
rect 4640 2050 4680 2060
rect 4290 2030 4330 2040
rect 3545 2020 3585 2030
rect 3545 2000 3555 2020
rect 3575 2000 3585 2020
rect 4070 2020 4110 2030
rect 4070 2000 4080 2020
rect 4100 2000 4110 2020
rect 4290 2010 4300 2030
rect 4320 2010 4330 2030
rect 4290 2000 4330 2010
rect 4665 2030 4680 2050
rect 4665 2020 5100 2030
rect 4665 2015 5070 2020
rect 3460 1975 3475 1990
rect 3525 1985 3735 2000
rect 4070 1990 4175 2000
rect 3525 1975 3540 1985
rect 3590 1975 3605 1985
rect 3655 1975 3670 1985
rect 3720 1975 3735 1985
rect 3785 1975 3800 1990
rect 4030 1975 4045 1990
rect 4095 1985 4175 1990
rect 4095 1975 4110 1985
rect 4160 1975 4175 1985
rect 4225 1985 4305 2000
rect 4225 1975 4240 1985
rect 4290 1975 4305 1985
rect 4355 1975 4370 1990
rect 4600 1975 4615 1990
rect 4665 1975 4680 2015
rect 4730 1975 4745 2015
rect 4795 1975 4810 2015
rect 4860 1975 4875 2015
rect 5060 2000 5070 2015
rect 5090 2000 5100 2020
rect 5060 1990 5100 2000
rect 4925 1975 4940 1990
rect 3460 1910 3475 1925
rect 3525 1910 3540 1925
rect 3590 1910 3605 1925
rect 3655 1910 3670 1925
rect 3720 1910 3735 1925
rect 3785 1910 3800 1925
rect 4030 1910 4045 1925
rect 4095 1910 4110 1925
rect 4160 1910 4175 1925
rect 4225 1910 4240 1925
rect 4290 1910 4305 1925
rect 4355 1910 4370 1925
rect 4600 1910 4615 1925
rect 4665 1910 4680 1925
rect 4730 1910 4745 1925
rect 4795 1910 4810 1925
rect 4860 1910 4875 1925
rect 4925 1910 4940 1925
rect 3445 1900 3490 1910
rect 3445 1875 3455 1900
rect 3480 1875 3490 1900
rect 3445 1865 3490 1875
rect 3770 1900 3815 1910
rect 3770 1875 3780 1900
rect 3805 1875 3815 1900
rect 3770 1865 3815 1875
rect 4015 1900 4055 1910
rect 4015 1880 4025 1900
rect 4045 1880 4055 1900
rect 4015 1870 4055 1880
rect 4345 1900 4385 1910
rect 4345 1880 4355 1900
rect 4375 1880 4385 1900
rect 4345 1870 4385 1880
rect 4585 1900 4625 1910
rect 4585 1880 4595 1900
rect 4615 1880 4625 1900
rect 4585 1870 4625 1880
rect 4915 1900 4955 1910
rect 4915 1880 4925 1900
rect 4945 1880 4955 1900
rect 4915 1870 4955 1880
rect 3390 1750 3430 1760
rect 3390 1730 3400 1750
rect 3420 1735 3430 1750
rect 4390 1750 4430 1760
rect 4390 1735 4400 1750
rect 3420 1730 3485 1735
rect 3390 1720 3485 1730
rect 4335 1730 4400 1735
rect 4420 1730 4430 1750
rect 4335 1720 4430 1730
rect 3435 1705 3485 1720
rect 3535 1705 3585 1720
rect 3635 1705 3685 1720
rect 3735 1705 3785 1720
rect 3835 1705 3885 1720
rect 3935 1705 3985 1720
rect 4035 1705 4085 1720
rect 4135 1705 4185 1720
rect 4235 1705 4285 1720
rect 4335 1705 4385 1720
rect 3435 1565 3485 1580
rect 3535 1570 3585 1580
rect 3635 1570 3685 1580
rect 3735 1570 3785 1580
rect 3835 1570 3885 1580
rect 3935 1570 3985 1580
rect 4035 1570 4085 1580
rect 4135 1570 4185 1580
rect 4235 1570 4285 1580
rect 3535 1555 4285 1570
rect 4335 1565 4385 1580
rect 3790 1535 3800 1555
rect 3820 1535 3830 1555
rect 3790 1525 3830 1535
rect 3990 1535 4000 1555
rect 4020 1535 4030 1555
rect 3990 1525 4030 1535
<< polycont >>
rect 3860 2810 3880 2830
rect 4060 2810 4080 2830
rect 3460 2490 3480 2510
rect 4460 2490 4480 2510
rect 3455 2335 3475 2355
rect 3785 2335 3805 2355
rect 4025 2335 4045 2355
rect 4355 2335 4375 2355
rect 4595 2335 4615 2355
rect 4925 2335 4945 2355
rect 3510 2165 3530 2185
rect 3730 2165 3750 2185
rect 4125 2160 4145 2180
rect 4650 2165 4670 2185
rect 5070 2165 5090 2185
rect 4650 2060 4670 2080
rect 3555 2000 3575 2020
rect 4080 2000 4100 2020
rect 4300 2010 4320 2030
rect 5070 2000 5090 2020
rect 3455 1875 3480 1900
rect 3780 1875 3805 1900
rect 4025 1880 4045 1900
rect 4355 1880 4375 1900
rect 4595 1880 4615 1900
rect 4925 1880 4945 1900
rect 3400 1730 3420 1750
rect 4400 1730 4420 1750
rect 3800 1535 3820 1555
rect 4000 1535 4020 1555
<< xpolycontact >>
rect 5105 2648 5140 2868
rect 5105 2330 5140 2550
rect 5105 1475 5140 1695
rect 3286 897 3506 1470
rect 3590 897 3810 1470
rect 5105 1185 5140 1405
<< xpolyres >>
rect 5105 2550 5140 2648
rect 3506 897 3590 1470
rect 5105 1405 5140 1475
<< locali >>
rect 5160 3195 5210 3205
rect 5160 3185 5170 3195
rect 5120 3165 5170 3185
rect 5200 3165 5210 3195
rect 5120 2868 5140 3165
rect 5160 3155 5210 3165
rect 3850 2830 3890 2840
rect 3850 2825 3860 2830
rect 3110 2810 3860 2825
rect 3880 2825 3890 2830
rect 4050 2830 4090 2840
rect 4050 2825 4060 2830
rect 3880 2810 4060 2825
rect 4080 2810 4090 2830
rect 3110 2805 4090 2810
rect 3110 1470 3130 2805
rect 3850 2800 3890 2805
rect 4050 2800 4090 2805
rect 3860 2780 3880 2800
rect 4060 2780 4080 2800
rect 3400 2770 3490 2780
rect 3400 2750 3410 2770
rect 3430 2750 3460 2770
rect 3480 2750 3490 2770
rect 3400 2720 3490 2750
rect 3400 2700 3410 2720
rect 3430 2700 3460 2720
rect 3480 2700 3490 2720
rect 3400 2670 3490 2700
rect 3400 2650 3410 2670
rect 3430 2650 3460 2670
rect 3480 2650 3490 2670
rect 3400 2620 3490 2650
rect 3400 2600 3410 2620
rect 3430 2600 3460 2620
rect 3480 2600 3490 2620
rect 3400 2570 3490 2600
rect 3400 2550 3410 2570
rect 3430 2550 3460 2570
rect 3480 2550 3490 2570
rect 3400 2540 3490 2550
rect 3550 2770 3590 2780
rect 3550 2750 3560 2770
rect 3580 2750 3590 2770
rect 3550 2720 3590 2750
rect 3550 2700 3560 2720
rect 3580 2700 3590 2720
rect 3550 2670 3590 2700
rect 3550 2650 3560 2670
rect 3580 2650 3590 2670
rect 3550 2620 3590 2650
rect 3550 2600 3560 2620
rect 3580 2600 3590 2620
rect 3550 2570 3590 2600
rect 3550 2550 3560 2570
rect 3580 2550 3590 2570
rect 3550 2540 3590 2550
rect 3650 2770 3690 2780
rect 3650 2750 3660 2770
rect 3680 2750 3690 2770
rect 3650 2720 3690 2750
rect 3650 2700 3660 2720
rect 3680 2700 3690 2720
rect 3650 2670 3690 2700
rect 3650 2650 3660 2670
rect 3680 2650 3690 2670
rect 3650 2620 3690 2650
rect 3650 2600 3660 2620
rect 3680 2600 3690 2620
rect 3650 2570 3690 2600
rect 3650 2550 3660 2570
rect 3680 2550 3690 2570
rect 3650 2540 3690 2550
rect 3750 2770 3790 2780
rect 3750 2750 3760 2770
rect 3780 2750 3790 2770
rect 3750 2720 3790 2750
rect 3750 2700 3760 2720
rect 3780 2700 3790 2720
rect 3750 2670 3790 2700
rect 3750 2650 3760 2670
rect 3780 2650 3790 2670
rect 3750 2620 3790 2650
rect 3750 2600 3760 2620
rect 3780 2600 3790 2620
rect 3750 2570 3790 2600
rect 3750 2550 3760 2570
rect 3780 2550 3790 2570
rect 3750 2540 3790 2550
rect 3850 2770 3890 2780
rect 3850 2750 3860 2770
rect 3880 2750 3890 2770
rect 3850 2720 3890 2750
rect 3850 2700 3860 2720
rect 3880 2700 3890 2720
rect 3850 2670 3890 2700
rect 3850 2650 3860 2670
rect 3880 2650 3890 2670
rect 3850 2620 3890 2650
rect 3850 2600 3860 2620
rect 3880 2600 3890 2620
rect 3850 2570 3890 2600
rect 3850 2550 3860 2570
rect 3880 2550 3890 2570
rect 3850 2540 3890 2550
rect 3950 2770 3990 2780
rect 3950 2750 3960 2770
rect 3980 2750 3990 2770
rect 3950 2720 3990 2750
rect 3950 2700 3960 2720
rect 3980 2700 3990 2720
rect 3950 2670 3990 2700
rect 3950 2650 3960 2670
rect 3980 2650 3990 2670
rect 3950 2620 3990 2650
rect 3950 2600 3960 2620
rect 3980 2600 3990 2620
rect 3950 2570 3990 2600
rect 3950 2550 3960 2570
rect 3980 2550 3990 2570
rect 3950 2540 3990 2550
rect 4050 2770 4090 2780
rect 4050 2750 4060 2770
rect 4080 2750 4090 2770
rect 4050 2720 4090 2750
rect 4050 2700 4060 2720
rect 4080 2700 4090 2720
rect 4050 2670 4090 2700
rect 4050 2650 4060 2670
rect 4080 2650 4090 2670
rect 4050 2620 4090 2650
rect 4050 2600 4060 2620
rect 4080 2600 4090 2620
rect 4050 2570 4090 2600
rect 4050 2550 4060 2570
rect 4080 2550 4090 2570
rect 4050 2540 4090 2550
rect 4150 2770 4190 2780
rect 4150 2750 4160 2770
rect 4180 2750 4190 2770
rect 4150 2720 4190 2750
rect 4150 2700 4160 2720
rect 4180 2700 4190 2720
rect 4150 2670 4190 2700
rect 4150 2650 4160 2670
rect 4180 2650 4190 2670
rect 4150 2620 4190 2650
rect 4150 2600 4160 2620
rect 4180 2600 4190 2620
rect 4150 2570 4190 2600
rect 4150 2550 4160 2570
rect 4180 2550 4190 2570
rect 4150 2540 4190 2550
rect 4250 2770 4290 2780
rect 4250 2750 4260 2770
rect 4280 2750 4290 2770
rect 4250 2720 4290 2750
rect 4250 2700 4260 2720
rect 4280 2700 4290 2720
rect 4250 2670 4290 2700
rect 4250 2650 4260 2670
rect 4280 2650 4290 2670
rect 4250 2620 4290 2650
rect 4250 2600 4260 2620
rect 4280 2600 4290 2620
rect 4250 2570 4290 2600
rect 4250 2550 4260 2570
rect 4280 2550 4290 2570
rect 4250 2540 4290 2550
rect 4350 2770 4390 2780
rect 4350 2750 4360 2770
rect 4380 2750 4390 2770
rect 4350 2720 4390 2750
rect 4350 2700 4360 2720
rect 4380 2700 4390 2720
rect 4350 2670 4390 2700
rect 4350 2650 4360 2670
rect 4380 2650 4390 2670
rect 4350 2620 4390 2650
rect 4350 2600 4360 2620
rect 4380 2600 4390 2620
rect 4350 2570 4390 2600
rect 4350 2550 4360 2570
rect 4380 2550 4390 2570
rect 4350 2540 4390 2550
rect 4450 2770 4540 2780
rect 4450 2750 4460 2770
rect 4480 2750 4510 2770
rect 4530 2750 4540 2770
rect 4450 2720 4540 2750
rect 4450 2700 4460 2720
rect 4480 2700 4510 2720
rect 4530 2700 4540 2720
rect 4450 2670 4540 2700
rect 4450 2650 4460 2670
rect 4480 2650 4510 2670
rect 4530 2650 4540 2670
rect 4450 2620 4540 2650
rect 4450 2600 4460 2620
rect 4480 2600 4510 2620
rect 4530 2600 4540 2620
rect 4450 2570 4540 2600
rect 4450 2550 4460 2570
rect 4480 2550 4510 2570
rect 4530 2550 4540 2570
rect 4450 2540 4540 2550
rect 3460 2520 3480 2540
rect 3450 2510 3490 2520
rect 3450 2490 3460 2510
rect 3480 2490 3490 2510
rect 3450 2480 3490 2490
rect 3660 2515 3680 2540
rect 4260 2515 4280 2540
rect 4460 2520 4480 2540
rect 3660 2495 4280 2515
rect 4450 2510 4490 2520
rect 3660 2485 3700 2495
rect 3660 2465 3670 2485
rect 3690 2465 3700 2485
rect 4450 2490 4460 2510
rect 4480 2490 4490 2510
rect 4450 2480 4490 2490
rect 3660 2455 3700 2465
rect 3250 2410 3280 2430
rect 3300 2410 3330 2430
rect 3350 2410 3380 2430
rect 3400 2410 3430 2430
rect 3450 2410 3480 2430
rect 3500 2410 3530 2430
rect 3550 2410 3580 2430
rect 3600 2410 3630 2430
rect 3650 2410 3680 2430
rect 3700 2410 3730 2430
rect 3750 2410 3780 2430
rect 3800 2410 3830 2430
rect 3850 2410 3880 2430
rect 3900 2410 3930 2430
rect 3950 2410 3980 2430
rect 4000 2410 4030 2430
rect 4050 2410 4080 2430
rect 4100 2410 4130 2430
rect 4150 2410 4180 2430
rect 4200 2410 4230 2430
rect 4250 2410 4280 2430
rect 4300 2410 4330 2430
rect 4350 2410 4380 2430
rect 4400 2410 4430 2430
rect 4450 2410 4480 2430
rect 4500 2410 4530 2430
rect 4550 2410 4580 2430
rect 4600 2410 4630 2430
rect 4650 2410 4680 2430
rect 4700 2410 4730 2430
rect 4750 2410 4780 2430
rect 3660 2375 3700 2385
rect 3445 2355 3485 2365
rect 3445 2345 3455 2355
rect 3425 2335 3455 2345
rect 3475 2345 3485 2355
rect 3660 2355 3670 2375
rect 3690 2355 3700 2375
rect 3660 2345 3700 2355
rect 3775 2355 3815 2365
rect 3775 2345 3785 2355
rect 3475 2335 3785 2345
rect 3805 2345 3815 2355
rect 4015 2355 4055 2365
rect 4015 2345 4025 2355
rect 3805 2335 3835 2345
rect 3425 2325 3835 2335
rect 3425 2305 3445 2325
rect 3490 2305 3510 2325
rect 3620 2305 3640 2325
rect 3750 2305 3770 2325
rect 3815 2305 3835 2325
rect 3995 2335 4025 2345
rect 4045 2345 4055 2355
rect 4190 2345 4210 2410
rect 4345 2355 4385 2365
rect 4345 2345 4355 2355
rect 4045 2335 4355 2345
rect 4375 2345 4385 2355
rect 4585 2355 4625 2365
rect 4585 2345 4595 2355
rect 4375 2335 4405 2345
rect 3995 2325 4405 2335
rect 3995 2305 4015 2325
rect 4060 2305 4080 2325
rect 4190 2305 4210 2325
rect 4320 2305 4340 2325
rect 4385 2305 4405 2325
rect 4565 2335 4595 2345
rect 4615 2345 4625 2355
rect 4760 2345 4780 2410
rect 4915 2355 4955 2365
rect 4915 2345 4925 2355
rect 4615 2335 4925 2345
rect 4945 2345 4955 2355
rect 4945 2335 4975 2345
rect 4565 2325 4975 2335
rect 4565 2305 4585 2325
rect 4630 2305 4650 2325
rect 4760 2305 4780 2325
rect 4890 2305 4910 2325
rect 4955 2305 4975 2325
rect 3410 2295 3455 2305
rect 3410 2275 3425 2295
rect 3445 2275 3455 2295
rect 3410 2245 3455 2275
rect 3410 2225 3425 2245
rect 3445 2225 3455 2245
rect 3410 2215 3455 2225
rect 3480 2295 3520 2305
rect 3480 2275 3490 2295
rect 3510 2275 3520 2295
rect 3480 2245 3520 2275
rect 3480 2225 3490 2245
rect 3510 2225 3520 2245
rect 3480 2215 3520 2225
rect 3545 2295 3585 2305
rect 3545 2275 3555 2295
rect 3575 2275 3585 2295
rect 3545 2245 3585 2275
rect 3545 2225 3555 2245
rect 3575 2225 3585 2245
rect 3545 2215 3585 2225
rect 3610 2295 3650 2305
rect 3610 2275 3620 2295
rect 3640 2275 3650 2295
rect 3610 2245 3650 2275
rect 3610 2225 3620 2245
rect 3640 2225 3650 2245
rect 3610 2215 3650 2225
rect 3675 2295 3715 2305
rect 3675 2275 3685 2295
rect 3705 2275 3715 2295
rect 3675 2245 3715 2275
rect 3675 2225 3685 2245
rect 3705 2225 3715 2245
rect 3675 2215 3715 2225
rect 3740 2295 3785 2305
rect 3740 2275 3750 2295
rect 3770 2275 3785 2295
rect 3740 2245 3785 2275
rect 3740 2225 3750 2245
rect 3770 2225 3785 2245
rect 3740 2215 3785 2225
rect 3805 2295 3850 2305
rect 3805 2275 3815 2295
rect 3835 2275 3850 2295
rect 3805 2245 3850 2275
rect 3805 2225 3815 2245
rect 3835 2225 3850 2245
rect 3805 2215 3850 2225
rect 3935 2295 4025 2305
rect 3935 2275 3945 2295
rect 3965 2275 3995 2295
rect 4015 2275 4025 2295
rect 3935 2245 4025 2275
rect 3935 2225 3945 2245
rect 3965 2225 3995 2245
rect 4015 2225 4025 2245
rect 3935 2215 4025 2225
rect 4050 2295 4090 2305
rect 4050 2275 4060 2295
rect 4080 2275 4090 2295
rect 4050 2245 4090 2275
rect 4050 2225 4060 2245
rect 4080 2225 4090 2245
rect 4050 2215 4090 2225
rect 4115 2295 4155 2305
rect 4115 2275 4125 2295
rect 4145 2275 4155 2295
rect 4115 2245 4155 2275
rect 4115 2225 4125 2245
rect 4145 2225 4155 2245
rect 4115 2215 4155 2225
rect 4180 2295 4220 2305
rect 4180 2275 4190 2295
rect 4210 2275 4220 2295
rect 4180 2245 4220 2275
rect 4180 2225 4190 2245
rect 4210 2225 4220 2245
rect 4180 2215 4220 2225
rect 4245 2295 4285 2305
rect 4245 2275 4255 2295
rect 4275 2275 4285 2295
rect 4245 2245 4285 2275
rect 4245 2225 4255 2245
rect 4275 2225 4285 2245
rect 4245 2215 4285 2225
rect 4310 2295 4350 2305
rect 4310 2275 4320 2295
rect 4340 2275 4350 2295
rect 4310 2245 4350 2275
rect 4310 2225 4320 2245
rect 4340 2225 4350 2245
rect 4310 2215 4350 2225
rect 4375 2295 4465 2305
rect 4375 2275 4385 2295
rect 4405 2275 4435 2295
rect 4455 2275 4465 2295
rect 4375 2245 4465 2275
rect 4375 2225 4385 2245
rect 4405 2225 4435 2245
rect 4455 2225 4465 2245
rect 4375 2215 4465 2225
rect 4505 2295 4595 2305
rect 4505 2275 4515 2295
rect 4535 2275 4565 2295
rect 4585 2275 4595 2295
rect 4505 2245 4595 2275
rect 4505 2225 4515 2245
rect 4535 2225 4565 2245
rect 4585 2225 4595 2245
rect 4505 2215 4595 2225
rect 4620 2295 4660 2305
rect 4620 2275 4630 2295
rect 4650 2275 4660 2295
rect 4620 2245 4660 2275
rect 4620 2225 4630 2245
rect 4650 2225 4660 2245
rect 4620 2215 4660 2225
rect 4685 2295 4725 2305
rect 4685 2275 4695 2295
rect 4715 2275 4725 2295
rect 4685 2245 4725 2275
rect 4685 2225 4695 2245
rect 4715 2225 4725 2245
rect 4685 2215 4725 2225
rect 4750 2295 4790 2305
rect 4750 2275 4760 2295
rect 4780 2275 4790 2295
rect 4750 2245 4790 2275
rect 4750 2225 4760 2245
rect 4780 2225 4790 2245
rect 4750 2215 4790 2225
rect 4815 2295 4855 2305
rect 4815 2275 4825 2295
rect 4845 2275 4855 2295
rect 4815 2245 4855 2275
rect 4815 2225 4825 2245
rect 4845 2225 4855 2245
rect 4815 2215 4855 2225
rect 4880 2295 4920 2305
rect 4880 2275 4890 2295
rect 4910 2275 4920 2295
rect 4880 2245 4920 2275
rect 4880 2225 4890 2245
rect 4910 2225 4920 2245
rect 4880 2215 4920 2225
rect 4945 2295 5035 2305
rect 4945 2275 4955 2295
rect 4975 2275 5005 2295
rect 5025 2275 5035 2295
rect 4945 2245 5035 2275
rect 4945 2225 4955 2245
rect 4975 2225 5005 2245
rect 5025 2225 5035 2245
rect 4945 2215 5035 2225
rect 3500 2185 3540 2195
rect 3500 2165 3510 2185
rect 3530 2165 3540 2185
rect 3500 2155 3540 2165
rect 3565 2030 3585 2215
rect 3545 2020 3585 2030
rect 3545 2000 3555 2020
rect 3575 2000 3585 2020
rect 3545 1990 3585 2000
rect 3565 1970 3585 1990
rect 3675 2095 3695 2215
rect 3720 2185 3760 2195
rect 4125 2190 4145 2215
rect 3720 2165 3730 2185
rect 3750 2165 3760 2185
rect 3720 2155 3760 2165
rect 4115 2180 4155 2190
rect 4115 2160 4125 2180
rect 4145 2160 4155 2180
rect 4115 2150 4155 2160
rect 3950 2105 3990 2110
rect 3950 2095 3960 2105
rect 3675 2085 3960 2095
rect 3980 2085 3990 2105
rect 3675 2075 3990 2085
rect 3675 1970 3695 2075
rect 4070 2020 4110 2030
rect 4070 2000 4080 2020
rect 4100 2000 4110 2020
rect 4070 1990 4110 2000
rect 4135 1970 4155 2150
rect 4245 2185 4265 2215
rect 4640 2185 4680 2195
rect 4245 2165 4650 2185
rect 4670 2165 4680 2185
rect 4245 1970 4265 2165
rect 4640 2155 4680 2165
rect 4705 2135 4725 2215
rect 4815 2135 4835 2215
rect 5060 2185 5100 2195
rect 5060 2165 5070 2185
rect 5090 2175 5100 2185
rect 5120 2175 5140 2330
rect 5090 2165 5140 2175
rect 5060 2155 5140 2165
rect 5160 2230 5215 2240
rect 5160 2195 5170 2230
rect 5205 2195 5215 2230
rect 5160 2185 5215 2195
rect 5160 2135 5180 2185
rect 4705 2115 5265 2135
rect 4640 2080 4680 2090
rect 4640 2060 4650 2080
rect 4670 2060 4680 2080
rect 5245 2070 5265 2115
rect 4640 2050 4680 2060
rect 4705 2050 5265 2070
rect 4290 2030 4330 2040
rect 4290 2010 4300 2030
rect 4320 2010 4330 2030
rect 4290 2000 4330 2010
rect 4705 1970 4725 2050
rect 4815 1970 4835 2050
rect 5060 2020 5140 2030
rect 5060 2000 5070 2020
rect 5090 2010 5140 2020
rect 5090 2000 5100 2010
rect 5060 1990 5100 2000
rect 3365 1960 3455 1970
rect 3365 1940 3375 1960
rect 3395 1940 3425 1960
rect 3445 1940 3455 1960
rect 3365 1930 3455 1940
rect 3480 1960 3520 1970
rect 3480 1940 3490 1960
rect 3510 1940 3520 1960
rect 3480 1930 3520 1940
rect 3545 1960 3585 1970
rect 3545 1940 3555 1960
rect 3575 1940 3585 1960
rect 3545 1930 3585 1940
rect 3610 1960 3650 1970
rect 3610 1940 3620 1960
rect 3640 1940 3650 1960
rect 3610 1930 3650 1940
rect 3675 1960 3715 1970
rect 3675 1940 3685 1960
rect 3705 1940 3715 1960
rect 3675 1930 3715 1940
rect 3740 1960 3780 1970
rect 3740 1940 3750 1960
rect 3770 1940 3780 1960
rect 3740 1930 3780 1940
rect 3805 1960 3895 1970
rect 3805 1940 3815 1960
rect 3835 1940 3865 1960
rect 3885 1940 3895 1960
rect 3805 1930 3895 1940
rect 3980 1960 4025 1970
rect 3980 1940 3995 1960
rect 4015 1940 4025 1960
rect 3980 1930 4025 1940
rect 4050 1960 4090 1970
rect 4050 1940 4060 1960
rect 4080 1940 4090 1960
rect 4050 1930 4090 1940
rect 4115 1960 4155 1970
rect 4115 1940 4125 1960
rect 4145 1940 4155 1960
rect 4115 1930 4155 1940
rect 4180 1960 4220 1970
rect 4180 1940 4190 1960
rect 4210 1940 4220 1960
rect 4180 1930 4220 1940
rect 4245 1960 4285 1970
rect 4245 1940 4255 1960
rect 4275 1940 4285 1960
rect 4245 1930 4285 1940
rect 4310 1960 4350 1970
rect 4310 1940 4320 1960
rect 4340 1940 4350 1960
rect 4310 1930 4350 1940
rect 4375 1960 4420 1970
rect 4375 1940 4385 1960
rect 4405 1940 4420 1960
rect 4375 1930 4420 1940
rect 4505 1960 4595 1970
rect 4505 1940 4515 1960
rect 4535 1940 4565 1960
rect 4585 1940 4595 1960
rect 4505 1930 4595 1940
rect 4620 1960 4660 1970
rect 4620 1940 4630 1960
rect 4650 1940 4660 1960
rect 4620 1930 4660 1940
rect 4685 1960 4725 1970
rect 4685 1940 4695 1960
rect 4715 1940 4725 1960
rect 4685 1930 4725 1940
rect 4750 1960 4790 1970
rect 4750 1940 4760 1960
rect 4780 1940 4790 1960
rect 4750 1930 4790 1940
rect 4815 1960 4855 1970
rect 4815 1940 4825 1960
rect 4845 1940 4855 1960
rect 4815 1930 4855 1940
rect 4880 1960 4920 1970
rect 4880 1940 4890 1960
rect 4910 1940 4920 1960
rect 4880 1930 4920 1940
rect 4945 1960 5035 1970
rect 4945 1940 4955 1960
rect 4975 1940 5005 1960
rect 5025 1940 5035 1960
rect 4945 1930 5035 1940
rect 3425 1910 3445 1930
rect 3490 1910 3510 1930
rect 3620 1910 3640 1930
rect 3750 1910 3770 1930
rect 3815 1910 3835 1930
rect 3425 1900 3835 1910
rect 3425 1890 3455 1900
rect 3445 1875 3455 1890
rect 3480 1890 3780 1900
rect 3480 1875 3490 1890
rect 3445 1865 3490 1875
rect 3620 1825 3640 1890
rect 3770 1875 3780 1890
rect 3805 1890 3835 1900
rect 3995 1910 4015 1930
rect 4060 1910 4080 1930
rect 4190 1910 4210 1930
rect 4320 1910 4340 1930
rect 4385 1910 4405 1930
rect 3995 1900 4405 1910
rect 3995 1890 4025 1900
rect 3805 1875 3815 1890
rect 3770 1865 3815 1875
rect 4015 1880 4025 1890
rect 4045 1890 4355 1900
rect 4045 1880 4055 1890
rect 4015 1870 4055 1880
rect 4180 1880 4220 1890
rect 4180 1860 4190 1880
rect 4210 1860 4220 1880
rect 4345 1880 4355 1890
rect 4375 1890 4405 1900
rect 4565 1910 4585 1930
rect 4630 1910 4650 1930
rect 4760 1910 4780 1930
rect 4890 1910 4910 1930
rect 4955 1910 4975 1930
rect 4565 1900 4975 1910
rect 4375 1880 4385 1890
rect 4565 1885 4595 1900
rect 4345 1870 4385 1880
rect 4585 1880 4595 1885
rect 4615 1885 4925 1900
rect 4615 1880 4625 1885
rect 4585 1870 4625 1880
rect 4180 1850 4220 1860
rect 4760 1825 4780 1885
rect 4915 1880 4925 1885
rect 4945 1885 4975 1900
rect 4945 1880 4955 1885
rect 4915 1870 4955 1880
rect 3250 1805 3280 1825
rect 3300 1805 3330 1825
rect 3350 1805 3380 1825
rect 3400 1805 3430 1825
rect 3450 1805 3480 1825
rect 3500 1805 3530 1825
rect 3550 1805 3580 1825
rect 3600 1805 3630 1825
rect 3650 1805 3680 1825
rect 3700 1805 3730 1825
rect 3750 1805 3780 1825
rect 3800 1805 3830 1825
rect 3850 1805 3880 1825
rect 3900 1805 3930 1825
rect 3950 1805 3980 1825
rect 4000 1805 4030 1825
rect 4050 1805 4080 1825
rect 4100 1805 4130 1825
rect 4150 1805 4180 1825
rect 4200 1805 4230 1825
rect 4250 1805 4280 1825
rect 4300 1805 4330 1825
rect 4350 1805 4380 1825
rect 4400 1805 4430 1825
rect 4450 1805 4480 1825
rect 4500 1805 4530 1825
rect 4550 1805 4580 1825
rect 4600 1805 4630 1825
rect 4650 1805 4680 1825
rect 4700 1805 4730 1825
rect 4750 1805 4780 1825
rect 4180 1770 4220 1780
rect 3390 1750 3430 1760
rect 3390 1730 3400 1750
rect 3420 1730 3430 1750
rect 4180 1750 4190 1770
rect 4210 1750 4220 1770
rect 4180 1740 4220 1750
rect 3390 1720 3430 1730
rect 3600 1720 4220 1740
rect 4390 1750 4430 1760
rect 4390 1730 4400 1750
rect 4420 1730 4430 1750
rect 4390 1720 4430 1730
rect 3400 1700 3420 1720
rect 3600 1700 3620 1720
rect 4200 1700 4220 1720
rect 4400 1700 4420 1720
rect 3340 1690 3430 1700
rect 3340 1665 3350 1690
rect 3370 1665 3400 1690
rect 3420 1665 3430 1690
rect 3340 1620 3430 1665
rect 3340 1595 3350 1620
rect 3370 1595 3400 1620
rect 3420 1595 3430 1620
rect 3340 1585 3430 1595
rect 3490 1690 3530 1700
rect 3490 1665 3500 1690
rect 3520 1665 3530 1690
rect 3490 1620 3530 1665
rect 3490 1595 3500 1620
rect 3520 1595 3530 1620
rect 3490 1585 3530 1595
rect 3590 1690 3630 1700
rect 3590 1665 3600 1690
rect 3620 1665 3630 1690
rect 3590 1620 3630 1665
rect 3590 1595 3600 1620
rect 3620 1595 3630 1620
rect 3590 1585 3630 1595
rect 3690 1690 3730 1700
rect 3690 1665 3700 1690
rect 3720 1665 3730 1690
rect 3690 1620 3730 1665
rect 3690 1595 3700 1620
rect 3720 1595 3730 1620
rect 3690 1585 3730 1595
rect 3790 1690 3830 1700
rect 3790 1665 3800 1690
rect 3820 1665 3830 1690
rect 3790 1620 3830 1665
rect 3790 1595 3800 1620
rect 3820 1595 3830 1620
rect 3790 1585 3830 1595
rect 3890 1690 3930 1700
rect 3890 1665 3900 1690
rect 3920 1665 3930 1690
rect 3890 1620 3930 1665
rect 3890 1595 3900 1620
rect 3920 1595 3930 1620
rect 3890 1585 3930 1595
rect 3990 1690 4030 1700
rect 3990 1665 4000 1690
rect 4020 1665 4030 1690
rect 3990 1620 4030 1665
rect 3990 1595 4000 1620
rect 4020 1595 4030 1620
rect 3990 1585 4030 1595
rect 4090 1690 4130 1700
rect 4090 1665 4100 1690
rect 4120 1665 4130 1690
rect 4090 1620 4130 1665
rect 4090 1595 4100 1620
rect 4120 1595 4130 1620
rect 4090 1585 4130 1595
rect 4190 1690 4230 1700
rect 4190 1665 4200 1690
rect 4220 1665 4230 1690
rect 4190 1620 4230 1665
rect 4190 1595 4200 1620
rect 4220 1595 4230 1620
rect 4190 1585 4230 1595
rect 4290 1690 4330 1700
rect 4290 1665 4300 1690
rect 4320 1665 4330 1690
rect 4290 1620 4330 1665
rect 4290 1595 4300 1620
rect 4320 1595 4330 1620
rect 4290 1585 4330 1595
rect 4390 1690 4480 1700
rect 5120 1695 5140 2010
rect 5160 1990 5180 2050
rect 5160 1980 5215 1990
rect 5160 1945 5170 1980
rect 5205 1945 5215 1980
rect 5160 1935 5215 1945
rect 4390 1665 4400 1690
rect 4420 1665 4450 1690
rect 4470 1665 4480 1690
rect 4390 1620 4480 1665
rect 4390 1595 4400 1620
rect 4420 1595 4450 1620
rect 4470 1595 4480 1620
rect 4390 1585 4480 1595
rect 3800 1565 3820 1585
rect 4000 1565 4020 1585
rect 3790 1555 4030 1565
rect 3790 1535 3800 1555
rect 3820 1545 4000 1555
rect 3820 1535 3830 1545
rect 3790 1525 3830 1535
rect 3990 1535 4000 1545
rect 4020 1535 4030 1555
rect 3990 1525 4030 1535
rect 4000 1470 4020 1525
rect 3110 1450 3286 1470
rect 3810 1450 4020 1470
rect 5120 1010 5140 1185
rect 5160 1010 5210 1020
rect 5120 990 5170 1010
rect 5160 980 5170 990
rect 5200 980 5210 1010
rect 5160 970 5210 980
<< viali >>
rect 5170 3165 5200 3195
rect 3560 2750 3580 2770
rect 3560 2700 3580 2720
rect 3560 2650 3580 2670
rect 3560 2600 3580 2620
rect 3560 2550 3580 2570
rect 3760 2750 3780 2770
rect 3760 2700 3780 2720
rect 3760 2650 3780 2670
rect 3760 2600 3780 2620
rect 3760 2550 3780 2570
rect 3960 2750 3980 2770
rect 3960 2700 3980 2720
rect 3960 2650 3980 2670
rect 3960 2600 3980 2620
rect 3960 2550 3980 2570
rect 4160 2750 4180 2770
rect 4160 2700 4180 2720
rect 4160 2650 4180 2670
rect 4160 2600 4180 2620
rect 4160 2550 4180 2570
rect 4360 2750 4380 2770
rect 4360 2700 4380 2720
rect 4360 2650 4380 2670
rect 4360 2600 4380 2620
rect 4360 2550 4380 2570
rect 3460 2490 3480 2510
rect 3670 2465 3690 2485
rect 3280 2410 3300 2430
rect 3330 2410 3350 2430
rect 3380 2410 3400 2430
rect 3430 2410 3450 2430
rect 3480 2410 3500 2430
rect 3530 2410 3550 2430
rect 3580 2410 3600 2430
rect 3630 2410 3650 2430
rect 3680 2410 3700 2430
rect 3730 2410 3750 2430
rect 3780 2410 3800 2430
rect 3830 2410 3850 2430
rect 3880 2410 3900 2430
rect 3930 2410 3950 2430
rect 3980 2410 4000 2430
rect 4030 2410 4050 2430
rect 4080 2410 4100 2430
rect 4130 2410 4150 2430
rect 4180 2410 4200 2430
rect 4230 2410 4250 2430
rect 4280 2410 4300 2430
rect 4330 2410 4350 2430
rect 4380 2410 4400 2430
rect 4430 2410 4450 2430
rect 4480 2410 4500 2430
rect 4530 2410 4550 2430
rect 4580 2410 4600 2430
rect 4630 2410 4650 2430
rect 4680 2410 4700 2430
rect 4730 2410 4750 2430
rect 3670 2355 3690 2375
rect 3510 2165 3530 2185
rect 3730 2165 3750 2185
rect 3960 2085 3980 2105
rect 4080 2000 4100 2020
rect 5170 2195 5205 2230
rect 4650 2060 4670 2080
rect 4300 2010 4320 2030
rect 4190 1860 4210 1880
rect 3280 1805 3300 1825
rect 3330 1805 3350 1825
rect 3380 1805 3400 1825
rect 3430 1805 3450 1825
rect 3480 1805 3500 1825
rect 3530 1805 3550 1825
rect 3580 1805 3600 1825
rect 3630 1805 3650 1825
rect 3680 1805 3700 1825
rect 3730 1805 3750 1825
rect 3780 1805 3800 1825
rect 3830 1805 3850 1825
rect 3880 1805 3900 1825
rect 3930 1805 3950 1825
rect 3980 1805 4000 1825
rect 4030 1805 4050 1825
rect 4080 1805 4100 1825
rect 4130 1805 4150 1825
rect 4180 1805 4200 1825
rect 4230 1805 4250 1825
rect 4280 1805 4300 1825
rect 4330 1805 4350 1825
rect 4380 1805 4400 1825
rect 4430 1805 4450 1825
rect 4480 1805 4500 1825
rect 4530 1805 4550 1825
rect 4580 1805 4600 1825
rect 4630 1805 4650 1825
rect 4680 1805 4700 1825
rect 4730 1805 4750 1825
rect 3400 1730 3420 1750
rect 4190 1750 4210 1770
rect 4400 1730 4420 1750
rect 3500 1665 3520 1690
rect 3500 1595 3520 1620
rect 3700 1665 3720 1690
rect 3700 1595 3720 1620
rect 3900 1665 3920 1690
rect 3900 1595 3920 1620
rect 4100 1665 4120 1690
rect 4100 1595 4120 1620
rect 4300 1665 4320 1690
rect 4300 1595 4320 1620
rect 5170 1945 5205 1980
rect 5170 980 5200 1010
<< metal1 >>
rect 5160 3195 5210 3205
rect 5160 3165 5170 3195
rect 5200 3165 5210 3195
rect 5160 3155 5210 3165
rect 3550 2770 3590 2780
rect 3550 2750 3560 2770
rect 3580 2750 3590 2770
rect 3550 2720 3590 2750
rect 3550 2700 3560 2720
rect 3580 2700 3590 2720
rect 3550 2670 3590 2700
rect 3550 2650 3560 2670
rect 3580 2650 3590 2670
rect 3550 2620 3590 2650
rect 3550 2600 3560 2620
rect 3580 2600 3590 2620
rect 3550 2570 3590 2600
rect 3550 2550 3560 2570
rect 3580 2550 3590 2570
rect 3550 2540 3590 2550
rect 3750 2770 3790 2780
rect 3750 2750 3760 2770
rect 3780 2750 3790 2770
rect 3750 2720 3790 2750
rect 3750 2700 3760 2720
rect 3780 2700 3790 2720
rect 3750 2670 3790 2700
rect 3750 2650 3760 2670
rect 3780 2650 3790 2670
rect 3750 2620 3790 2650
rect 3750 2600 3760 2620
rect 3780 2600 3790 2620
rect 3750 2570 3790 2600
rect 3750 2550 3760 2570
rect 3780 2550 3790 2570
rect 3750 2540 3790 2550
rect 3950 2770 3990 2780
rect 3950 2750 3960 2770
rect 3980 2750 3990 2770
rect 3950 2720 3990 2750
rect 3950 2700 3960 2720
rect 3980 2700 3990 2720
rect 3950 2670 3990 2700
rect 3950 2650 3960 2670
rect 3980 2650 3990 2670
rect 3950 2620 3990 2650
rect 3950 2600 3960 2620
rect 3980 2600 3990 2620
rect 3950 2570 3990 2600
rect 3950 2550 3960 2570
rect 3980 2550 3990 2570
rect 3950 2540 3990 2550
rect 4150 2770 4190 2780
rect 4150 2750 4160 2770
rect 4180 2750 4190 2770
rect 4150 2720 4190 2750
rect 4150 2700 4160 2720
rect 4180 2700 4190 2720
rect 4150 2670 4190 2700
rect 4150 2650 4160 2670
rect 4180 2650 4190 2670
rect 4150 2620 4190 2650
rect 4150 2600 4160 2620
rect 4180 2600 4190 2620
rect 4150 2570 4190 2600
rect 4150 2550 4160 2570
rect 4180 2550 4190 2570
rect 4150 2540 4190 2550
rect 4350 2770 4390 2780
rect 4350 2750 4360 2770
rect 4380 2750 4390 2770
rect 4350 2720 4390 2750
rect 4350 2700 4360 2720
rect 4380 2700 4390 2720
rect 4350 2670 4390 2700
rect 4350 2650 4360 2670
rect 4380 2650 4390 2670
rect 4350 2620 4390 2650
rect 4350 2600 4360 2620
rect 4380 2600 4390 2620
rect 4350 2570 4390 2600
rect 4350 2550 4360 2570
rect 4380 2550 4390 2570
rect 4350 2540 4390 2550
rect 3450 2510 3490 2520
rect 3450 2490 3460 2510
rect 3480 2490 3490 2510
rect 3450 2480 3490 2490
rect 3460 2440 3480 2480
rect 3560 2440 3580 2540
rect 3660 2490 3700 2495
rect 3660 2460 3665 2490
rect 3695 2460 3700 2490
rect 3660 2455 3700 2460
rect 3760 2440 3780 2540
rect 3960 2440 3980 2540
rect 4160 2440 4180 2540
rect 4360 2440 4380 2540
rect 4450 2480 4490 2520
rect 4460 2440 4480 2480
rect 3250 2430 4780 2440
rect 3250 2410 3280 2430
rect 3300 2410 3330 2430
rect 3350 2410 3380 2430
rect 3400 2410 3430 2430
rect 3450 2410 3480 2430
rect 3500 2410 3530 2430
rect 3550 2410 3580 2430
rect 3600 2410 3630 2430
rect 3650 2410 3680 2430
rect 3700 2410 3730 2430
rect 3750 2410 3780 2430
rect 3800 2410 3830 2430
rect 3850 2410 3880 2430
rect 3900 2410 3930 2430
rect 3950 2410 3980 2430
rect 4000 2410 4030 2430
rect 4050 2410 4080 2430
rect 4100 2410 4130 2430
rect 4150 2410 4180 2430
rect 4200 2410 4230 2430
rect 4250 2410 4280 2430
rect 4300 2410 4330 2430
rect 4350 2410 4380 2430
rect 4400 2410 4430 2430
rect 4450 2410 4480 2430
rect 4500 2410 4530 2430
rect 4550 2410 4580 2430
rect 4600 2410 4630 2430
rect 4650 2410 4680 2430
rect 4700 2410 4730 2430
rect 4750 2410 4780 2430
rect 3250 2400 4780 2410
rect 3660 2380 3700 2385
rect 3660 2350 3665 2380
rect 3695 2350 3700 2380
rect 3660 2345 3700 2350
rect 5160 2230 5215 2240
rect 5160 2195 5170 2230
rect 5205 2195 5215 2230
rect 3500 2190 3540 2195
rect 3500 2160 3505 2190
rect 3535 2160 3540 2190
rect 3500 2155 3540 2160
rect 3720 2190 3760 2195
rect 3720 2160 3725 2190
rect 3755 2160 3760 2190
rect 5160 2185 5215 2195
rect 3720 2155 3760 2160
rect 4070 2140 4110 2145
rect 3340 2135 4075 2140
rect 3340 2125 3505 2135
rect 3500 2105 3505 2125
rect 3535 2125 4075 2135
rect 3535 2105 3540 2125
rect 4070 2110 4075 2125
rect 4105 2110 4110 2140
rect 3500 2100 3540 2105
rect 3950 2105 3990 2110
rect 4070 2105 4110 2110
rect 3950 2085 3960 2105
rect 3980 2090 3990 2105
rect 3980 2085 4680 2090
rect 3950 2080 4680 2085
rect 3950 2075 4650 2080
rect 4640 2060 4650 2075
rect 4670 2060 4680 2080
rect 3340 2055 4330 2060
rect 3340 2045 3735 2055
rect 3730 2025 3735 2045
rect 3765 2045 4330 2055
rect 4640 2050 4680 2060
rect 3765 2025 3770 2045
rect 4290 2030 4330 2045
rect 3730 2020 3770 2025
rect 4070 2025 4110 2030
rect 4070 1995 4075 2025
rect 4105 1995 4110 2025
rect 4290 2010 4300 2030
rect 4320 2010 4330 2030
rect 4290 2000 4330 2010
rect 4070 1990 4110 1995
rect 5160 1980 5215 1990
rect 5160 1945 5170 1980
rect 5205 1945 5215 1980
rect 5160 1935 5215 1945
rect 4180 1885 4220 1890
rect 4180 1855 4185 1885
rect 4215 1855 4220 1885
rect 4180 1850 4220 1855
rect 3250 1825 4780 1835
rect 3250 1805 3280 1825
rect 3300 1805 3330 1825
rect 3350 1805 3380 1825
rect 3400 1805 3430 1825
rect 3450 1805 3480 1825
rect 3500 1805 3530 1825
rect 3550 1805 3580 1825
rect 3600 1805 3630 1825
rect 3650 1805 3680 1825
rect 3700 1805 3730 1825
rect 3750 1805 3780 1825
rect 3800 1805 3830 1825
rect 3850 1805 3880 1825
rect 3900 1805 3930 1825
rect 3950 1805 3980 1825
rect 4000 1805 4030 1825
rect 4050 1805 4080 1825
rect 4100 1805 4130 1825
rect 4150 1805 4180 1825
rect 4200 1805 4230 1825
rect 4250 1805 4280 1825
rect 4300 1805 4330 1825
rect 4350 1805 4380 1825
rect 4400 1805 4430 1825
rect 4450 1805 4480 1825
rect 4500 1805 4530 1825
rect 4550 1805 4580 1825
rect 4600 1805 4630 1825
rect 4650 1805 4680 1825
rect 4700 1805 4730 1825
rect 4750 1805 4780 1825
rect 3250 1795 4780 1805
rect 3400 1760 3420 1795
rect 3390 1750 3430 1760
rect 3390 1730 3400 1750
rect 3420 1730 3430 1750
rect 3390 1720 3430 1730
rect 3500 1700 3520 1795
rect 3700 1700 3720 1795
rect 3900 1700 3920 1795
rect 4100 1700 4120 1795
rect 4180 1775 4220 1780
rect 4180 1745 4185 1775
rect 4215 1745 4220 1775
rect 4180 1740 4220 1745
rect 4300 1700 4320 1795
rect 4400 1760 4420 1795
rect 4390 1750 4430 1760
rect 4390 1730 4400 1750
rect 4420 1730 4430 1750
rect 4390 1720 4430 1730
rect 3490 1690 3530 1700
rect 3490 1665 3500 1690
rect 3520 1665 3530 1690
rect 3490 1620 3530 1665
rect 3490 1595 3500 1620
rect 3520 1595 3530 1620
rect 3490 1585 3530 1595
rect 3690 1690 3730 1700
rect 3690 1665 3700 1690
rect 3720 1665 3730 1690
rect 3690 1620 3730 1665
rect 3690 1595 3700 1620
rect 3720 1595 3730 1620
rect 3690 1585 3730 1595
rect 3890 1690 3930 1700
rect 3890 1665 3900 1690
rect 3920 1665 3930 1690
rect 3890 1620 3930 1665
rect 3890 1595 3900 1620
rect 3920 1595 3930 1620
rect 3890 1585 3930 1595
rect 4090 1690 4130 1700
rect 4090 1665 4100 1690
rect 4120 1665 4130 1690
rect 4090 1620 4130 1665
rect 4090 1595 4100 1620
rect 4120 1595 4130 1620
rect 4090 1585 4130 1595
rect 4290 1690 4330 1700
rect 4290 1665 4300 1690
rect 4320 1665 4330 1690
rect 4290 1620 4330 1665
rect 4290 1595 4300 1620
rect 4320 1595 4330 1620
rect 4290 1585 4330 1595
rect 5160 1010 5210 1020
rect 5160 980 5170 1010
rect 5200 980 5210 1010
rect 5160 970 5210 980
<< via1 >>
rect 5170 3165 5200 3195
rect 3665 2485 3695 2490
rect 3665 2465 3670 2485
rect 3670 2465 3690 2485
rect 3690 2465 3695 2485
rect 3665 2460 3695 2465
rect 3665 2375 3695 2380
rect 3665 2355 3670 2375
rect 3670 2355 3690 2375
rect 3690 2355 3695 2375
rect 3665 2350 3695 2355
rect 5170 2195 5205 2230
rect 3505 2185 3535 2190
rect 3505 2165 3510 2185
rect 3510 2165 3530 2185
rect 3530 2165 3535 2185
rect 3505 2160 3535 2165
rect 3725 2185 3755 2190
rect 3725 2165 3730 2185
rect 3730 2165 3750 2185
rect 3750 2165 3755 2185
rect 3725 2160 3755 2165
rect 3505 2105 3535 2135
rect 4075 2110 4105 2140
rect 3735 2025 3765 2055
rect 4075 2020 4105 2025
rect 4075 2000 4080 2020
rect 4080 2000 4100 2020
rect 4100 2000 4105 2020
rect 4075 1995 4105 2000
rect 5170 1945 5205 1980
rect 4185 1880 4215 1885
rect 4185 1860 4190 1880
rect 4190 1860 4210 1880
rect 4210 1860 4215 1880
rect 4185 1855 4215 1860
rect 4185 1770 4215 1775
rect 4185 1750 4190 1770
rect 4190 1750 4210 1770
rect 4210 1750 4215 1770
rect 4185 1745 4215 1750
rect 5170 980 5200 1010
<< metal2 >>
rect 5160 3195 5210 3205
rect 5160 3165 5170 3195
rect 5200 3165 5210 3195
rect 5160 3155 5210 3165
rect 3660 2490 3700 2495
rect 3660 2460 3665 2490
rect 3695 2460 3700 2490
rect 3660 2455 3700 2460
rect 3670 2385 3690 2455
rect 3660 2380 3700 2385
rect 3660 2350 3665 2380
rect 3695 2350 3700 2380
rect 3660 2345 3700 2350
rect 5160 2230 5215 2240
rect 5160 2195 5170 2230
rect 5205 2195 5215 2230
rect 3500 2190 3540 2195
rect 3500 2160 3505 2190
rect 3535 2160 3540 2190
rect 3500 2155 3540 2160
rect 3720 2190 3760 2195
rect 3720 2160 3725 2190
rect 3755 2160 3760 2190
rect 5160 2185 5215 2195
rect 3720 2155 3760 2160
rect 3510 2140 3525 2155
rect 3500 2135 3540 2140
rect 3500 2105 3505 2135
rect 3535 2105 3540 2135
rect 3500 2100 3540 2105
rect 3730 2060 3745 2155
rect 4070 2140 4110 2145
rect 4070 2110 4075 2140
rect 4105 2110 4110 2140
rect 4070 2105 4110 2110
rect 3730 2055 3770 2060
rect 3730 2025 3735 2055
rect 3765 2025 3770 2055
rect 4080 2030 4095 2105
rect 3730 2020 3770 2025
rect 4070 2025 4110 2030
rect 4070 1995 4075 2025
rect 4105 1995 4110 2025
rect 4070 1990 4110 1995
rect 5160 1980 5215 1990
rect 5160 1945 5170 1980
rect 5205 1945 5215 1980
rect 5160 1935 5215 1945
rect 4180 1885 4220 1890
rect 4180 1855 4185 1885
rect 4215 1855 4220 1885
rect 4180 1850 4220 1855
rect 4190 1780 4210 1850
rect 4180 1775 4220 1780
rect 4180 1745 4185 1775
rect 4215 1745 4220 1775
rect 4180 1740 4220 1745
rect 5160 1010 5210 1020
rect 5160 980 5170 1010
rect 5200 980 5210 1010
rect 5160 970 5210 980
<< via2 >>
rect 5170 3165 5200 3195
rect 5170 2195 5205 2230
rect 5170 1945 5205 1980
rect 5170 980 5200 1010
<< metal3 >>
rect 5160 3200 5210 3205
rect 5160 3195 6365 3200
rect 5160 3165 5170 3195
rect 5200 3165 6365 3195
rect 5160 3155 6365 3165
rect 5160 2230 5215 2240
rect 5160 2195 5170 2230
rect 5205 2195 5215 2230
rect 5160 2185 5215 2195
rect 5335 2170 6365 3155
rect 5160 1980 5215 1990
rect 5160 1945 5170 1980
rect 5205 1945 5215 1980
rect 5160 1935 5215 1945
rect 5335 1020 6365 2005
rect 5160 1010 6365 1020
rect 5160 980 5170 1010
rect 5200 980 6365 1010
rect 5160 975 6365 980
rect 5160 970 5210 975
<< via3 >>
rect 5170 2195 5205 2230
rect 5170 1945 5205 1980
<< mimcap >>
rect 5350 2230 6350 3185
rect 5350 2195 5360 2230
rect 5395 2195 6350 2230
rect 5350 2185 6350 2195
rect 5350 1980 6350 1990
rect 5350 1945 5360 1980
rect 5395 1945 6350 1980
rect 5350 990 6350 1945
<< mimcapcontact >>
rect 5360 2195 5395 2230
rect 5360 1945 5395 1980
<< metal4 >>
rect 5160 2230 5400 2240
rect 5160 2195 5170 2230
rect 5205 2195 5360 2230
rect 5395 2195 5400 2230
rect 5160 2185 5400 2195
rect 5160 1980 5400 1990
rect 5160 1945 5170 1980
rect 5205 1945 5360 1980
rect 5395 1945 5400 1980
rect 5160 1935 5400 1945
<< labels >>
flabel locali 3250 2420 3250 2420 7 FreeSans 400 0 -200 0 VDDA
port 1 w
flabel locali 3250 1815 3250 1815 7 FreeSans 400 0 -200 0 GNDA
port 5 w
flabel locali 5265 2090 5265 2090 3 FreeSans 400 0 200 0 VOUT
port 4 e
flabel locali 3110 2700 3110 2700 7 FreeSans 160 0 -80 0 p_bias
flabel locali 4265 2185 4265 2185 3 FreeSans 160 0 80 0 n_right
flabel locali 4155 2130 4155 2130 3 FreeSans 160 0 80 0 n_left
flabel metal1 3340 2050 3340 2050 7 FreeSans 400 0 -200 -200 VIN+
port 2 w
flabel metal1 3340 2130 3340 2130 7 FreeSans 400 0 -200 0 VIN-
port 3 w
<< end >>
