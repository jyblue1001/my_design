magic
tech sky130A
timestamp 1754401177
<< nwell >>
rect 56025 4510 56365 4900
rect 56495 4510 56835 4730
rect 56965 4510 57305 4900
rect 57435 4510 57775 4900
rect 54530 3645 55410 4035
rect 55945 3645 56825 4035
rect 56975 3645 57855 4035
rect 58390 3645 59270 4035
rect 54560 2535 55380 3175
rect 56450 2900 57350 3190
rect 58420 2535 59240 3175
rect 58915 2530 59055 2535
rect 54560 1660 55380 1900
rect 58420 1660 59240 1900
<< nmos >>
rect 56810 2315 56825 2565
rect 56865 2315 56880 2565
rect 56920 2315 56935 2565
rect 56975 2315 56990 2565
rect 56070 1745 56085 1895
rect 56125 1745 56140 1895
rect 56180 1745 56195 1895
rect 56235 1745 56250 1895
rect 56290 1745 56305 1895
rect 56345 1745 56360 1895
rect 56400 1745 56415 1895
rect 56455 1745 56470 1895
rect 56510 1745 56525 1895
rect 56565 1745 56580 1895
rect 56620 1745 56635 1895
rect 56675 1745 56690 1895
rect 57110 1745 57125 1895
rect 57165 1745 57180 1895
rect 57220 1745 57235 1895
rect 57275 1745 57290 1895
rect 57330 1745 57345 1895
rect 57385 1745 57400 1895
rect 57440 1745 57455 1895
rect 57495 1745 57510 1895
rect 57550 1745 57565 1895
rect 57605 1745 57620 1895
rect 57660 1745 57675 1895
rect 57715 1745 57730 1895
rect 54660 1140 54675 1440
rect 54715 1140 54730 1440
rect 54770 1140 54785 1440
rect 54825 1140 54840 1440
rect 54880 1140 54895 1440
rect 54935 1140 54950 1440
rect 54990 1140 55005 1440
rect 55045 1140 55060 1440
rect 55100 1140 55115 1440
rect 55155 1140 55170 1440
rect 55210 1140 55225 1440
rect 55265 1140 55280 1440
rect 56070 1070 56085 1220
rect 56125 1070 56140 1220
rect 56180 1070 56195 1220
rect 56235 1070 56250 1220
rect 56290 1070 56305 1220
rect 56345 1070 56360 1220
rect 56400 1070 56415 1220
rect 56455 1070 56470 1220
rect 56510 1070 56525 1220
rect 56565 1070 56580 1220
rect 56620 1070 56635 1220
rect 56675 1070 56690 1220
rect 56810 1070 56825 1220
rect 56865 1070 56880 1220
rect 56920 1070 56935 1220
rect 56975 1070 56990 1220
rect 57110 1070 57125 1220
rect 57165 1070 57180 1220
rect 57220 1070 57235 1220
rect 57275 1070 57290 1220
rect 57330 1070 57345 1220
rect 57385 1070 57400 1220
rect 57440 1070 57455 1220
rect 57495 1070 57510 1220
rect 57550 1070 57565 1220
rect 57605 1070 57620 1220
rect 57660 1070 57675 1220
rect 57715 1070 57730 1220
rect 58520 1140 58535 1440
rect 58575 1140 58590 1440
rect 58630 1140 58645 1440
rect 58685 1140 58700 1440
rect 58740 1140 58755 1440
rect 58795 1140 58810 1440
rect 58850 1140 58865 1440
rect 58905 1140 58920 1440
rect 58960 1140 58975 1440
rect 59015 1140 59030 1440
rect 59070 1140 59085 1440
rect 59125 1140 59140 1440
rect 54690 -360 54750 340
rect 54790 -360 54850 340
rect 54890 -360 54950 340
rect 54990 -360 55050 340
rect 55090 -360 55150 340
rect 55190 -360 55250 340
rect 56260 170 56275 420
rect 56315 170 56330 420
rect 56370 170 56385 420
rect 56425 170 56440 420
rect 56480 170 56495 420
rect 56535 170 56550 420
rect 56590 170 56605 420
rect 56645 170 56660 420
rect 56700 170 56715 420
rect 56755 170 56770 420
rect 56810 170 56825 420
rect 56865 170 56880 420
rect 56920 170 56935 420
rect 56975 170 56990 420
rect 57030 170 57045 420
rect 57085 170 57100 420
rect 57140 170 57155 420
rect 57195 170 57210 420
rect 57250 170 57265 420
rect 57305 170 57320 420
rect 57360 170 57375 420
rect 57415 170 57430 420
rect 57470 170 57485 420
rect 56470 -450 56485 -300
rect 56525 -450 56540 -300
rect 56580 -450 56595 -300
rect 56635 -450 56650 -300
rect 56690 -450 56705 -300
rect 56745 -450 56760 -300
rect 56910 -450 57210 -300
rect 58550 -360 58610 340
rect 58650 -360 58710 340
rect 58750 -360 58810 340
rect 58850 -360 58910 340
rect 58950 -360 59010 340
rect 59050 -360 59110 340
<< pmos >>
rect 56125 4530 56145 4880
rect 56185 4530 56205 4880
rect 56245 4530 56265 4880
rect 56595 4530 56615 4710
rect 56655 4530 56675 4710
rect 56715 4530 56735 4710
rect 57065 4530 57085 4880
rect 57125 4530 57145 4880
rect 57185 4530 57205 4880
rect 57535 4530 57555 4880
rect 57595 4530 57615 4880
rect 57655 4530 57675 4880
rect 54630 3665 54650 4015
rect 54690 3665 54710 4015
rect 54750 3665 54770 4015
rect 54810 3665 54830 4015
rect 54870 3665 54890 4015
rect 54930 3665 54950 4015
rect 54990 3665 55010 4015
rect 55050 3665 55070 4015
rect 55110 3665 55130 4015
rect 55170 3665 55190 4015
rect 55230 3665 55250 4015
rect 55290 3665 55310 4015
rect 56045 3665 56065 4015
rect 56105 3665 56125 4015
rect 56165 3665 56185 4015
rect 56225 3665 56245 4015
rect 56285 3665 56305 4015
rect 56345 3665 56365 4015
rect 56405 3665 56425 4015
rect 56465 3665 56485 4015
rect 56525 3665 56545 4015
rect 56585 3665 56605 4015
rect 56645 3665 56665 4015
rect 56705 3665 56725 4015
rect 57075 3665 57095 4015
rect 57135 3665 57155 4015
rect 57195 3665 57215 4015
rect 57255 3665 57275 4015
rect 57315 3665 57335 4015
rect 57375 3665 57395 4015
rect 57435 3665 57455 4015
rect 57495 3665 57515 4015
rect 57555 3665 57575 4015
rect 57615 3665 57635 4015
rect 57675 3665 57695 4015
rect 57735 3665 57755 4015
rect 58490 3665 58510 4015
rect 58550 3665 58570 4015
rect 58610 3665 58630 4015
rect 58670 3665 58690 4015
rect 58730 3665 58750 4015
rect 58790 3665 58810 4015
rect 58850 3665 58870 4015
rect 58910 3665 58930 4015
rect 58970 3665 58990 4015
rect 59030 3665 59050 4015
rect 59090 3665 59110 4015
rect 59150 3665 59170 4015
rect 54660 2555 54675 3155
rect 54715 2555 54730 3155
rect 54770 2555 54785 3155
rect 54825 2555 54840 3155
rect 54880 2555 54895 3155
rect 54935 2555 54950 3155
rect 54990 2555 55005 3155
rect 55045 2555 55060 3155
rect 55100 2555 55115 3155
rect 55155 2555 55170 3155
rect 55210 2555 55225 3155
rect 55265 2555 55280 3155
rect 56550 2920 56565 3170
rect 56605 2920 56620 3170
rect 56660 2920 56675 3170
rect 56715 2920 56730 3170
rect 56770 2920 56785 3170
rect 56825 2920 56840 3170
rect 56960 2920 56975 3170
rect 57015 2920 57030 3170
rect 57070 2920 57085 3170
rect 57125 2920 57140 3170
rect 57180 2920 57195 3170
rect 57235 2920 57250 3170
rect 58520 2555 58535 3155
rect 58575 2555 58590 3155
rect 58630 2555 58645 3155
rect 58685 2555 58700 3155
rect 58740 2555 58755 3155
rect 58795 2555 58810 3155
rect 58850 2555 58865 3155
rect 58905 2555 58920 3155
rect 58960 2555 58975 3155
rect 59015 2555 59030 3155
rect 59070 2555 59085 3155
rect 59125 2555 59140 3155
rect 54660 1680 54675 1880
rect 54715 1680 54730 1880
rect 54770 1680 54785 1880
rect 54825 1680 54840 1880
rect 54880 1680 54895 1880
rect 54935 1680 54950 1880
rect 54990 1680 55005 1880
rect 55045 1680 55060 1880
rect 55100 1680 55115 1880
rect 55155 1680 55170 1880
rect 55210 1680 55225 1880
rect 55265 1680 55280 1880
rect 58520 1680 58535 1880
rect 58575 1680 58590 1880
rect 58630 1680 58645 1880
rect 58685 1680 58700 1880
rect 58740 1680 58755 1880
rect 58795 1680 58810 1880
rect 58850 1680 58865 1880
rect 58905 1680 58920 1880
rect 58960 1680 58975 1880
rect 59015 1680 59030 1880
rect 59070 1680 59085 1880
rect 59125 1680 59140 1880
<< ndiff >>
rect 56770 2550 56810 2565
rect 56770 2330 56780 2550
rect 56800 2330 56810 2550
rect 56770 2315 56810 2330
rect 56825 2550 56865 2565
rect 56825 2330 56835 2550
rect 56855 2330 56865 2550
rect 56825 2315 56865 2330
rect 56880 2550 56920 2565
rect 56880 2330 56890 2550
rect 56910 2330 56920 2550
rect 56880 2315 56920 2330
rect 56935 2550 56975 2565
rect 56935 2330 56945 2550
rect 56965 2330 56975 2550
rect 56935 2315 56975 2330
rect 56990 2550 57030 2565
rect 56990 2330 57000 2550
rect 57020 2330 57030 2550
rect 56990 2315 57030 2330
rect 56030 1880 56070 1895
rect 56030 1760 56040 1880
rect 56060 1760 56070 1880
rect 56030 1745 56070 1760
rect 56085 1880 56125 1895
rect 56085 1760 56095 1880
rect 56115 1760 56125 1880
rect 56085 1745 56125 1760
rect 56140 1880 56180 1895
rect 56140 1760 56150 1880
rect 56170 1760 56180 1880
rect 56140 1745 56180 1760
rect 56195 1880 56235 1895
rect 56195 1760 56205 1880
rect 56225 1760 56235 1880
rect 56195 1745 56235 1760
rect 56250 1880 56290 1895
rect 56250 1760 56260 1880
rect 56280 1760 56290 1880
rect 56250 1745 56290 1760
rect 56305 1880 56345 1895
rect 56305 1760 56315 1880
rect 56335 1760 56345 1880
rect 56305 1745 56345 1760
rect 56360 1880 56400 1895
rect 56360 1760 56370 1880
rect 56390 1760 56400 1880
rect 56360 1745 56400 1760
rect 56415 1880 56455 1895
rect 56415 1760 56425 1880
rect 56445 1760 56455 1880
rect 56415 1745 56455 1760
rect 56470 1880 56510 1895
rect 56470 1760 56480 1880
rect 56500 1760 56510 1880
rect 56470 1745 56510 1760
rect 56525 1880 56565 1895
rect 56525 1760 56535 1880
rect 56555 1760 56565 1880
rect 56525 1745 56565 1760
rect 56580 1880 56620 1895
rect 56580 1760 56590 1880
rect 56610 1760 56620 1880
rect 56580 1745 56620 1760
rect 56635 1880 56675 1895
rect 56635 1760 56645 1880
rect 56665 1760 56675 1880
rect 56635 1745 56675 1760
rect 56690 1880 56730 1895
rect 56690 1760 56700 1880
rect 56720 1760 56730 1880
rect 56690 1745 56730 1760
rect 57070 1880 57110 1895
rect 57070 1760 57080 1880
rect 57100 1760 57110 1880
rect 57070 1745 57110 1760
rect 57125 1880 57165 1895
rect 57125 1760 57135 1880
rect 57155 1760 57165 1880
rect 57125 1745 57165 1760
rect 57180 1880 57220 1895
rect 57180 1760 57190 1880
rect 57210 1760 57220 1880
rect 57180 1745 57220 1760
rect 57235 1880 57275 1895
rect 57235 1760 57245 1880
rect 57265 1760 57275 1880
rect 57235 1745 57275 1760
rect 57290 1880 57330 1895
rect 57290 1760 57300 1880
rect 57320 1760 57330 1880
rect 57290 1745 57330 1760
rect 57345 1880 57385 1895
rect 57345 1760 57355 1880
rect 57375 1760 57385 1880
rect 57345 1745 57385 1760
rect 57400 1880 57440 1895
rect 57400 1760 57410 1880
rect 57430 1760 57440 1880
rect 57400 1745 57440 1760
rect 57455 1880 57495 1895
rect 57455 1760 57465 1880
rect 57485 1760 57495 1880
rect 57455 1745 57495 1760
rect 57510 1880 57550 1895
rect 57510 1760 57520 1880
rect 57540 1760 57550 1880
rect 57510 1745 57550 1760
rect 57565 1880 57605 1895
rect 57565 1760 57575 1880
rect 57595 1760 57605 1880
rect 57565 1745 57605 1760
rect 57620 1880 57660 1895
rect 57620 1760 57630 1880
rect 57650 1760 57660 1880
rect 57620 1745 57660 1760
rect 57675 1880 57715 1895
rect 57675 1760 57685 1880
rect 57705 1760 57715 1880
rect 57675 1745 57715 1760
rect 57730 1880 57770 1895
rect 57730 1760 57740 1880
rect 57760 1760 57770 1880
rect 57730 1745 57770 1760
rect 54620 1425 54660 1440
rect 54620 1155 54630 1425
rect 54650 1155 54660 1425
rect 54620 1140 54660 1155
rect 54675 1425 54715 1440
rect 54675 1155 54685 1425
rect 54705 1155 54715 1425
rect 54675 1140 54715 1155
rect 54730 1425 54770 1440
rect 54730 1155 54740 1425
rect 54760 1155 54770 1425
rect 54730 1140 54770 1155
rect 54785 1425 54825 1440
rect 54785 1155 54795 1425
rect 54815 1155 54825 1425
rect 54785 1140 54825 1155
rect 54840 1425 54880 1440
rect 54840 1155 54850 1425
rect 54870 1155 54880 1425
rect 54840 1140 54880 1155
rect 54895 1425 54935 1440
rect 54895 1155 54905 1425
rect 54925 1155 54935 1425
rect 54895 1140 54935 1155
rect 54950 1425 54990 1440
rect 54950 1155 54960 1425
rect 54980 1155 54990 1425
rect 54950 1140 54990 1155
rect 55005 1425 55045 1440
rect 55005 1155 55015 1425
rect 55035 1155 55045 1425
rect 55005 1140 55045 1155
rect 55060 1425 55100 1440
rect 55060 1155 55070 1425
rect 55090 1155 55100 1425
rect 55060 1140 55100 1155
rect 55115 1425 55155 1440
rect 55115 1155 55125 1425
rect 55145 1155 55155 1425
rect 55115 1140 55155 1155
rect 55170 1425 55210 1440
rect 55170 1155 55180 1425
rect 55200 1155 55210 1425
rect 55170 1140 55210 1155
rect 55225 1425 55265 1440
rect 55225 1155 55235 1425
rect 55255 1155 55265 1425
rect 55225 1140 55265 1155
rect 55280 1425 55320 1440
rect 55280 1155 55290 1425
rect 55310 1155 55320 1425
rect 58480 1425 58520 1440
rect 55280 1140 55320 1155
rect 56030 1205 56070 1220
rect 56030 1085 56040 1205
rect 56060 1085 56070 1205
rect 56030 1070 56070 1085
rect 56085 1205 56125 1220
rect 56085 1085 56095 1205
rect 56115 1085 56125 1205
rect 56085 1070 56125 1085
rect 56140 1205 56180 1220
rect 56140 1085 56150 1205
rect 56170 1085 56180 1205
rect 56140 1070 56180 1085
rect 56195 1205 56235 1220
rect 56195 1085 56205 1205
rect 56225 1085 56235 1205
rect 56195 1070 56235 1085
rect 56250 1205 56290 1220
rect 56250 1085 56260 1205
rect 56280 1085 56290 1205
rect 56250 1070 56290 1085
rect 56305 1205 56345 1220
rect 56305 1085 56315 1205
rect 56335 1085 56345 1205
rect 56305 1070 56345 1085
rect 56360 1205 56400 1220
rect 56360 1085 56370 1205
rect 56390 1085 56400 1205
rect 56360 1070 56400 1085
rect 56415 1205 56455 1220
rect 56415 1085 56425 1205
rect 56445 1085 56455 1205
rect 56415 1070 56455 1085
rect 56470 1205 56510 1220
rect 56470 1085 56480 1205
rect 56500 1085 56510 1205
rect 56470 1070 56510 1085
rect 56525 1205 56565 1220
rect 56525 1085 56535 1205
rect 56555 1085 56565 1205
rect 56525 1070 56565 1085
rect 56580 1205 56620 1220
rect 56580 1085 56590 1205
rect 56610 1085 56620 1205
rect 56580 1070 56620 1085
rect 56635 1205 56675 1220
rect 56635 1085 56645 1205
rect 56665 1085 56675 1205
rect 56635 1070 56675 1085
rect 56690 1205 56730 1220
rect 56770 1205 56810 1220
rect 56690 1085 56700 1205
rect 56720 1085 56730 1205
rect 56770 1085 56780 1205
rect 56800 1085 56810 1205
rect 56690 1070 56730 1085
rect 56770 1070 56810 1085
rect 56825 1205 56865 1220
rect 56825 1085 56835 1205
rect 56855 1085 56865 1205
rect 56825 1070 56865 1085
rect 56880 1205 56920 1220
rect 56880 1085 56890 1205
rect 56910 1085 56920 1205
rect 56880 1070 56920 1085
rect 56935 1205 56975 1220
rect 56935 1085 56945 1205
rect 56965 1085 56975 1205
rect 56935 1070 56975 1085
rect 56990 1205 57030 1220
rect 57070 1205 57110 1220
rect 56990 1085 57000 1205
rect 57020 1085 57030 1205
rect 57070 1085 57080 1205
rect 57100 1085 57110 1205
rect 56990 1070 57030 1085
rect 57070 1070 57110 1085
rect 57125 1205 57165 1220
rect 57125 1085 57135 1205
rect 57155 1085 57165 1205
rect 57125 1070 57165 1085
rect 57180 1205 57220 1220
rect 57180 1085 57190 1205
rect 57210 1085 57220 1205
rect 57180 1070 57220 1085
rect 57235 1205 57275 1220
rect 57235 1085 57245 1205
rect 57265 1085 57275 1205
rect 57235 1070 57275 1085
rect 57290 1205 57330 1220
rect 57290 1085 57300 1205
rect 57320 1085 57330 1205
rect 57290 1070 57330 1085
rect 57345 1205 57385 1220
rect 57345 1085 57355 1205
rect 57375 1085 57385 1205
rect 57345 1070 57385 1085
rect 57400 1205 57440 1220
rect 57400 1085 57410 1205
rect 57430 1085 57440 1205
rect 57400 1070 57440 1085
rect 57455 1205 57495 1220
rect 57455 1085 57465 1205
rect 57485 1085 57495 1205
rect 57455 1070 57495 1085
rect 57510 1205 57550 1220
rect 57510 1085 57520 1205
rect 57540 1085 57550 1205
rect 57510 1070 57550 1085
rect 57565 1205 57605 1220
rect 57565 1085 57575 1205
rect 57595 1085 57605 1205
rect 57565 1070 57605 1085
rect 57620 1205 57660 1220
rect 57620 1085 57630 1205
rect 57650 1085 57660 1205
rect 57620 1070 57660 1085
rect 57675 1205 57715 1220
rect 57675 1085 57685 1205
rect 57705 1085 57715 1205
rect 57675 1070 57715 1085
rect 57730 1205 57770 1220
rect 57730 1085 57740 1205
rect 57760 1085 57770 1205
rect 58480 1155 58490 1425
rect 58510 1155 58520 1425
rect 58480 1140 58520 1155
rect 58535 1425 58575 1440
rect 58535 1155 58545 1425
rect 58565 1155 58575 1425
rect 58535 1140 58575 1155
rect 58590 1425 58630 1440
rect 58590 1155 58600 1425
rect 58620 1155 58630 1425
rect 58590 1140 58630 1155
rect 58645 1425 58685 1440
rect 58645 1155 58655 1425
rect 58675 1155 58685 1425
rect 58645 1140 58685 1155
rect 58700 1425 58740 1440
rect 58700 1155 58710 1425
rect 58730 1155 58740 1425
rect 58700 1140 58740 1155
rect 58755 1425 58795 1440
rect 58755 1155 58765 1425
rect 58785 1155 58795 1425
rect 58755 1140 58795 1155
rect 58810 1425 58850 1440
rect 58810 1155 58820 1425
rect 58840 1155 58850 1425
rect 58810 1140 58850 1155
rect 58865 1425 58905 1440
rect 58865 1155 58875 1425
rect 58895 1155 58905 1425
rect 58865 1140 58905 1155
rect 58920 1425 58960 1440
rect 58920 1155 58930 1425
rect 58950 1155 58960 1425
rect 58920 1140 58960 1155
rect 58975 1425 59015 1440
rect 58975 1155 58985 1425
rect 59005 1155 59015 1425
rect 58975 1140 59015 1155
rect 59030 1425 59070 1440
rect 59030 1155 59040 1425
rect 59060 1155 59070 1425
rect 59030 1140 59070 1155
rect 59085 1425 59125 1440
rect 59085 1155 59095 1425
rect 59115 1155 59125 1425
rect 59085 1140 59125 1155
rect 59140 1425 59180 1440
rect 59140 1155 59150 1425
rect 59170 1155 59180 1425
rect 59140 1140 59180 1155
rect 57730 1070 57770 1085
rect 56220 405 56260 420
rect 54650 325 54690 340
rect 54650 -345 54660 325
rect 54680 -345 54690 325
rect 54650 -360 54690 -345
rect 54750 325 54790 340
rect 54750 -345 54760 325
rect 54780 -345 54790 325
rect 54750 -360 54790 -345
rect 54850 325 54890 340
rect 54850 -345 54860 325
rect 54880 -345 54890 325
rect 54850 -360 54890 -345
rect 54950 325 54990 340
rect 54950 -345 54960 325
rect 54980 -345 54990 325
rect 54950 -360 54990 -345
rect 55050 325 55090 340
rect 55050 -345 55060 325
rect 55080 -345 55090 325
rect 55050 -360 55090 -345
rect 55150 325 55190 340
rect 55150 -345 55160 325
rect 55180 -345 55190 325
rect 55150 -360 55190 -345
rect 55250 325 55290 340
rect 55250 -345 55260 325
rect 55280 -345 55290 325
rect 56220 185 56230 405
rect 56250 185 56260 405
rect 56220 170 56260 185
rect 56275 405 56315 420
rect 56275 185 56285 405
rect 56305 185 56315 405
rect 56275 170 56315 185
rect 56330 405 56370 420
rect 56330 185 56340 405
rect 56360 185 56370 405
rect 56330 170 56370 185
rect 56385 405 56425 420
rect 56385 185 56395 405
rect 56415 185 56425 405
rect 56385 170 56425 185
rect 56440 405 56480 420
rect 56440 185 56450 405
rect 56470 185 56480 405
rect 56440 170 56480 185
rect 56495 405 56535 420
rect 56495 185 56505 405
rect 56525 185 56535 405
rect 56495 170 56535 185
rect 56550 405 56590 420
rect 56550 185 56560 405
rect 56580 185 56590 405
rect 56550 170 56590 185
rect 56605 405 56645 420
rect 56605 185 56615 405
rect 56635 185 56645 405
rect 56605 170 56645 185
rect 56660 405 56700 420
rect 56660 185 56670 405
rect 56690 185 56700 405
rect 56660 170 56700 185
rect 56715 405 56755 420
rect 56715 185 56725 405
rect 56745 185 56755 405
rect 56715 170 56755 185
rect 56770 405 56810 420
rect 56770 185 56780 405
rect 56800 185 56810 405
rect 56770 170 56810 185
rect 56825 405 56865 420
rect 56825 185 56835 405
rect 56855 185 56865 405
rect 56825 170 56865 185
rect 56880 405 56920 420
rect 56880 185 56890 405
rect 56910 185 56920 405
rect 56880 170 56920 185
rect 56935 405 56975 420
rect 56935 185 56945 405
rect 56965 185 56975 405
rect 56935 170 56975 185
rect 56990 405 57030 420
rect 56990 185 57000 405
rect 57020 185 57030 405
rect 56990 170 57030 185
rect 57045 405 57085 420
rect 57045 185 57055 405
rect 57075 185 57085 405
rect 57045 170 57085 185
rect 57100 405 57140 420
rect 57100 185 57110 405
rect 57130 185 57140 405
rect 57100 170 57140 185
rect 57155 405 57195 420
rect 57155 185 57165 405
rect 57185 185 57195 405
rect 57155 170 57195 185
rect 57210 405 57250 420
rect 57210 185 57220 405
rect 57240 185 57250 405
rect 57210 170 57250 185
rect 57265 405 57305 420
rect 57265 185 57275 405
rect 57295 185 57305 405
rect 57265 170 57305 185
rect 57320 405 57360 420
rect 57320 185 57330 405
rect 57350 185 57360 405
rect 57320 170 57360 185
rect 57375 405 57415 420
rect 57375 185 57385 405
rect 57405 185 57415 405
rect 57375 170 57415 185
rect 57430 405 57470 420
rect 57430 185 57440 405
rect 57460 185 57470 405
rect 57430 170 57470 185
rect 57485 405 57525 420
rect 57485 185 57495 405
rect 57515 185 57525 405
rect 57485 170 57525 185
rect 58510 325 58550 340
rect 55250 -360 55290 -345
rect 56430 -315 56470 -300
rect 56430 -435 56440 -315
rect 56460 -435 56470 -315
rect 56430 -450 56470 -435
rect 56485 -315 56525 -300
rect 56485 -435 56495 -315
rect 56515 -435 56525 -315
rect 56485 -450 56525 -435
rect 56540 -315 56580 -300
rect 56540 -435 56550 -315
rect 56570 -435 56580 -315
rect 56540 -450 56580 -435
rect 56595 -315 56635 -300
rect 56595 -435 56605 -315
rect 56625 -435 56635 -315
rect 56595 -450 56635 -435
rect 56650 -315 56690 -300
rect 56650 -435 56660 -315
rect 56680 -435 56690 -315
rect 56650 -450 56690 -435
rect 56705 -315 56745 -300
rect 56705 -435 56715 -315
rect 56735 -435 56745 -315
rect 56705 -450 56745 -435
rect 56760 -315 56800 -300
rect 56760 -435 56770 -315
rect 56790 -435 56800 -315
rect 56760 -450 56800 -435
rect 56870 -315 56910 -300
rect 56870 -435 56880 -315
rect 56900 -435 56910 -315
rect 56870 -450 56910 -435
rect 57210 -325 57250 -300
rect 57210 -425 57220 -325
rect 57240 -425 57250 -325
rect 58510 -345 58520 325
rect 58540 -345 58550 325
rect 58510 -360 58550 -345
rect 58610 325 58650 340
rect 58610 -345 58620 325
rect 58640 -345 58650 325
rect 58610 -360 58650 -345
rect 58710 325 58750 340
rect 58710 -345 58720 325
rect 58740 -345 58750 325
rect 58710 -360 58750 -345
rect 58810 325 58850 340
rect 58810 -345 58820 325
rect 58840 -345 58850 325
rect 58810 -360 58850 -345
rect 58910 325 58950 340
rect 58910 -345 58920 325
rect 58940 -345 58950 325
rect 58910 -360 58950 -345
rect 59010 325 59050 340
rect 59010 -345 59020 325
rect 59040 -345 59050 325
rect 59010 -360 59050 -345
rect 59110 325 59150 340
rect 59110 -345 59120 325
rect 59140 -345 59150 325
rect 59110 -360 59150 -345
rect 57210 -450 57250 -425
<< pdiff >>
rect 56085 4865 56125 4880
rect 56085 4545 56095 4865
rect 56115 4545 56125 4865
rect 56085 4530 56125 4545
rect 56145 4865 56185 4880
rect 56145 4545 56155 4865
rect 56175 4545 56185 4865
rect 56145 4530 56185 4545
rect 56205 4865 56245 4880
rect 56205 4545 56215 4865
rect 56235 4545 56245 4865
rect 56205 4530 56245 4545
rect 56265 4865 56305 4880
rect 56265 4545 56275 4865
rect 56295 4545 56305 4865
rect 57025 4865 57065 4880
rect 56265 4530 56305 4545
rect 56555 4695 56595 4710
rect 56555 4545 56565 4695
rect 56585 4545 56595 4695
rect 56555 4530 56595 4545
rect 56615 4695 56655 4710
rect 56615 4545 56625 4695
rect 56645 4545 56655 4695
rect 56615 4530 56655 4545
rect 56675 4695 56715 4710
rect 56675 4545 56685 4695
rect 56705 4545 56715 4695
rect 56675 4530 56715 4545
rect 56735 4695 56775 4710
rect 56735 4545 56745 4695
rect 56765 4545 56775 4695
rect 56735 4530 56775 4545
rect 57025 4545 57035 4865
rect 57055 4545 57065 4865
rect 57025 4530 57065 4545
rect 57085 4865 57125 4880
rect 57085 4545 57095 4865
rect 57115 4545 57125 4865
rect 57085 4530 57125 4545
rect 57145 4865 57185 4880
rect 57145 4545 57155 4865
rect 57175 4545 57185 4865
rect 57145 4530 57185 4545
rect 57205 4865 57245 4880
rect 57205 4545 57215 4865
rect 57235 4545 57245 4865
rect 57205 4530 57245 4545
rect 57495 4865 57535 4880
rect 57495 4545 57505 4865
rect 57525 4545 57535 4865
rect 57495 4530 57535 4545
rect 57555 4865 57595 4880
rect 57555 4545 57565 4865
rect 57585 4545 57595 4865
rect 57555 4530 57595 4545
rect 57615 4865 57655 4880
rect 57615 4545 57625 4865
rect 57645 4545 57655 4865
rect 57615 4530 57655 4545
rect 57675 4865 57715 4880
rect 57675 4545 57685 4865
rect 57705 4545 57715 4865
rect 57675 4530 57715 4545
rect 54590 4000 54630 4015
rect 54590 3680 54600 4000
rect 54620 3680 54630 4000
rect 54590 3665 54630 3680
rect 54650 4000 54690 4015
rect 54650 3680 54660 4000
rect 54680 3680 54690 4000
rect 54650 3665 54690 3680
rect 54710 4000 54750 4015
rect 54710 3680 54720 4000
rect 54740 3680 54750 4000
rect 54710 3665 54750 3680
rect 54770 4000 54810 4015
rect 54770 3680 54780 4000
rect 54800 3680 54810 4000
rect 54770 3665 54810 3680
rect 54830 4000 54870 4015
rect 54830 3680 54840 4000
rect 54860 3680 54870 4000
rect 54830 3665 54870 3680
rect 54890 4000 54930 4015
rect 54890 3680 54900 4000
rect 54920 3680 54930 4000
rect 54890 3665 54930 3680
rect 54950 4000 54990 4015
rect 54950 3680 54960 4000
rect 54980 3680 54990 4000
rect 54950 3665 54990 3680
rect 55010 4000 55050 4015
rect 55010 3680 55020 4000
rect 55040 3680 55050 4000
rect 55010 3665 55050 3680
rect 55070 4000 55110 4015
rect 55070 3680 55080 4000
rect 55100 3680 55110 4000
rect 55070 3665 55110 3680
rect 55130 4000 55170 4015
rect 55130 3680 55140 4000
rect 55160 3680 55170 4000
rect 55130 3665 55170 3680
rect 55190 4000 55230 4015
rect 55190 3680 55200 4000
rect 55220 3680 55230 4000
rect 55190 3665 55230 3680
rect 55250 4000 55290 4015
rect 55250 3680 55260 4000
rect 55280 3680 55290 4000
rect 55250 3665 55290 3680
rect 55310 4000 55350 4015
rect 55310 3680 55320 4000
rect 55340 3680 55350 4000
rect 55310 3665 55350 3680
rect 56005 4000 56045 4015
rect 56005 3680 56015 4000
rect 56035 3680 56045 4000
rect 56005 3665 56045 3680
rect 56065 4000 56105 4015
rect 56065 3680 56075 4000
rect 56095 3680 56105 4000
rect 56065 3665 56105 3680
rect 56125 4000 56165 4015
rect 56125 3680 56135 4000
rect 56155 3680 56165 4000
rect 56125 3665 56165 3680
rect 56185 4000 56225 4015
rect 56185 3680 56195 4000
rect 56215 3680 56225 4000
rect 56185 3665 56225 3680
rect 56245 4000 56285 4015
rect 56245 3680 56255 4000
rect 56275 3680 56285 4000
rect 56245 3665 56285 3680
rect 56305 4000 56345 4015
rect 56305 3680 56315 4000
rect 56335 3680 56345 4000
rect 56305 3665 56345 3680
rect 56365 4000 56405 4015
rect 56365 3680 56375 4000
rect 56395 3680 56405 4000
rect 56365 3665 56405 3680
rect 56425 4000 56465 4015
rect 56425 3680 56435 4000
rect 56455 3680 56465 4000
rect 56425 3665 56465 3680
rect 56485 4000 56525 4015
rect 56485 3680 56495 4000
rect 56515 3680 56525 4000
rect 56485 3665 56525 3680
rect 56545 4000 56585 4015
rect 56545 3680 56555 4000
rect 56575 3680 56585 4000
rect 56545 3665 56585 3680
rect 56605 4000 56645 4015
rect 56605 3680 56615 4000
rect 56635 3680 56645 4000
rect 56605 3665 56645 3680
rect 56665 4000 56705 4015
rect 56665 3680 56675 4000
rect 56695 3680 56705 4000
rect 56665 3665 56705 3680
rect 56725 4000 56765 4015
rect 56725 3680 56735 4000
rect 56755 3680 56765 4000
rect 56725 3665 56765 3680
rect 57035 4000 57075 4015
rect 57035 3680 57045 4000
rect 57065 3680 57075 4000
rect 57035 3665 57075 3680
rect 57095 4000 57135 4015
rect 57095 3680 57105 4000
rect 57125 3680 57135 4000
rect 57095 3665 57135 3680
rect 57155 4000 57195 4015
rect 57155 3680 57165 4000
rect 57185 3680 57195 4000
rect 57155 3665 57195 3680
rect 57215 4000 57255 4015
rect 57215 3680 57225 4000
rect 57245 3680 57255 4000
rect 57215 3665 57255 3680
rect 57275 4000 57315 4015
rect 57275 3680 57285 4000
rect 57305 3680 57315 4000
rect 57275 3665 57315 3680
rect 57335 4000 57375 4015
rect 57335 3680 57345 4000
rect 57365 3680 57375 4000
rect 57335 3665 57375 3680
rect 57395 4000 57435 4015
rect 57395 3680 57405 4000
rect 57425 3680 57435 4000
rect 57395 3665 57435 3680
rect 57455 4000 57495 4015
rect 57455 3680 57465 4000
rect 57485 3680 57495 4000
rect 57455 3665 57495 3680
rect 57515 4000 57555 4015
rect 57515 3680 57525 4000
rect 57545 3680 57555 4000
rect 57515 3665 57555 3680
rect 57575 4000 57615 4015
rect 57575 3680 57585 4000
rect 57605 3680 57615 4000
rect 57575 3665 57615 3680
rect 57635 4000 57675 4015
rect 57635 3680 57645 4000
rect 57665 3680 57675 4000
rect 57635 3665 57675 3680
rect 57695 4000 57735 4015
rect 57695 3680 57705 4000
rect 57725 3680 57735 4000
rect 57695 3665 57735 3680
rect 57755 4000 57795 4015
rect 57755 3680 57765 4000
rect 57785 3680 57795 4000
rect 57755 3665 57795 3680
rect 58450 4000 58490 4015
rect 58450 3680 58460 4000
rect 58480 3680 58490 4000
rect 58450 3665 58490 3680
rect 58510 4000 58550 4015
rect 58510 3680 58520 4000
rect 58540 3680 58550 4000
rect 58510 3665 58550 3680
rect 58570 4000 58610 4015
rect 58570 3680 58580 4000
rect 58600 3680 58610 4000
rect 58570 3665 58610 3680
rect 58630 4000 58670 4015
rect 58630 3680 58640 4000
rect 58660 3680 58670 4000
rect 58630 3665 58670 3680
rect 58690 4000 58730 4015
rect 58690 3680 58700 4000
rect 58720 3680 58730 4000
rect 58690 3665 58730 3680
rect 58750 4000 58790 4015
rect 58750 3680 58760 4000
rect 58780 3680 58790 4000
rect 58750 3665 58790 3680
rect 58810 4000 58850 4015
rect 58810 3680 58820 4000
rect 58840 3680 58850 4000
rect 58810 3665 58850 3680
rect 58870 4000 58910 4015
rect 58870 3680 58880 4000
rect 58900 3680 58910 4000
rect 58870 3665 58910 3680
rect 58930 4000 58970 4015
rect 58930 3680 58940 4000
rect 58960 3680 58970 4000
rect 58930 3665 58970 3680
rect 58990 4000 59030 4015
rect 58990 3680 59000 4000
rect 59020 3680 59030 4000
rect 58990 3665 59030 3680
rect 59050 4000 59090 4015
rect 59050 3680 59060 4000
rect 59080 3680 59090 4000
rect 59050 3665 59090 3680
rect 59110 4000 59150 4015
rect 59110 3680 59120 4000
rect 59140 3680 59150 4000
rect 59110 3665 59150 3680
rect 59170 4000 59210 4015
rect 59170 3680 59180 4000
rect 59200 3680 59210 4000
rect 59170 3665 59210 3680
rect 56510 3155 56550 3170
rect 54620 3140 54660 3155
rect 54620 2570 54630 3140
rect 54650 2570 54660 3140
rect 54620 2555 54660 2570
rect 54675 3140 54715 3155
rect 54675 2570 54685 3140
rect 54705 2570 54715 3140
rect 54675 2555 54715 2570
rect 54730 3140 54770 3155
rect 54730 2570 54740 3140
rect 54760 2570 54770 3140
rect 54730 2555 54770 2570
rect 54785 3140 54825 3155
rect 54785 2570 54795 3140
rect 54815 2570 54825 3140
rect 54785 2555 54825 2570
rect 54840 3140 54880 3155
rect 54840 2570 54850 3140
rect 54870 2570 54880 3140
rect 54840 2555 54880 2570
rect 54895 3140 54935 3155
rect 54895 2570 54905 3140
rect 54925 2570 54935 3140
rect 54895 2555 54935 2570
rect 54950 3140 54990 3155
rect 54950 2570 54960 3140
rect 54980 2570 54990 3140
rect 54950 2555 54990 2570
rect 55005 3140 55045 3155
rect 55005 2570 55015 3140
rect 55035 2570 55045 3140
rect 55005 2555 55045 2570
rect 55060 3140 55100 3155
rect 55060 2570 55070 3140
rect 55090 2570 55100 3140
rect 55060 2555 55100 2570
rect 55115 3140 55155 3155
rect 55115 2570 55125 3140
rect 55145 2570 55155 3140
rect 55115 2555 55155 2570
rect 55170 3140 55210 3155
rect 55170 2570 55180 3140
rect 55200 2570 55210 3140
rect 55170 2555 55210 2570
rect 55225 3140 55265 3155
rect 55225 2570 55235 3140
rect 55255 2570 55265 3140
rect 55225 2555 55265 2570
rect 55280 3140 55320 3155
rect 55280 2570 55290 3140
rect 55310 2570 55320 3140
rect 56510 3135 56520 3155
rect 56540 3135 56550 3155
rect 56510 3105 56550 3135
rect 56510 3085 56520 3105
rect 56540 3085 56550 3105
rect 56510 3055 56550 3085
rect 56510 3035 56520 3055
rect 56540 3035 56550 3055
rect 56510 3005 56550 3035
rect 56510 2985 56520 3005
rect 56540 2985 56550 3005
rect 56510 2955 56550 2985
rect 56510 2935 56520 2955
rect 56540 2935 56550 2955
rect 56510 2920 56550 2935
rect 56565 3155 56605 3170
rect 56565 3135 56575 3155
rect 56595 3135 56605 3155
rect 56565 3105 56605 3135
rect 56565 3085 56575 3105
rect 56595 3085 56605 3105
rect 56565 3055 56605 3085
rect 56565 3035 56575 3055
rect 56595 3035 56605 3055
rect 56565 3005 56605 3035
rect 56565 2985 56575 3005
rect 56595 2985 56605 3005
rect 56565 2955 56605 2985
rect 56565 2935 56575 2955
rect 56595 2935 56605 2955
rect 56565 2920 56605 2935
rect 56620 3155 56660 3170
rect 56620 3135 56630 3155
rect 56650 3135 56660 3155
rect 56620 3105 56660 3135
rect 56620 3085 56630 3105
rect 56650 3085 56660 3105
rect 56620 3055 56660 3085
rect 56620 3035 56630 3055
rect 56650 3035 56660 3055
rect 56620 3005 56660 3035
rect 56620 2985 56630 3005
rect 56650 2985 56660 3005
rect 56620 2955 56660 2985
rect 56620 2935 56630 2955
rect 56650 2935 56660 2955
rect 56620 2920 56660 2935
rect 56675 3155 56715 3170
rect 56675 3135 56685 3155
rect 56705 3135 56715 3155
rect 56675 3105 56715 3135
rect 56675 3085 56685 3105
rect 56705 3085 56715 3105
rect 56675 3055 56715 3085
rect 56675 3035 56685 3055
rect 56705 3035 56715 3055
rect 56675 3005 56715 3035
rect 56675 2985 56685 3005
rect 56705 2985 56715 3005
rect 56675 2955 56715 2985
rect 56675 2935 56685 2955
rect 56705 2935 56715 2955
rect 56675 2920 56715 2935
rect 56730 3155 56770 3170
rect 56730 3135 56740 3155
rect 56760 3135 56770 3155
rect 56730 3105 56770 3135
rect 56730 3085 56740 3105
rect 56760 3085 56770 3105
rect 56730 3055 56770 3085
rect 56730 3035 56740 3055
rect 56760 3035 56770 3055
rect 56730 3005 56770 3035
rect 56730 2985 56740 3005
rect 56760 2985 56770 3005
rect 56730 2955 56770 2985
rect 56730 2935 56740 2955
rect 56760 2935 56770 2955
rect 56730 2920 56770 2935
rect 56785 3155 56825 3170
rect 56785 3135 56795 3155
rect 56815 3135 56825 3155
rect 56785 3105 56825 3135
rect 56785 3085 56795 3105
rect 56815 3085 56825 3105
rect 56785 3055 56825 3085
rect 56785 3035 56795 3055
rect 56815 3035 56825 3055
rect 56785 3005 56825 3035
rect 56785 2985 56795 3005
rect 56815 2985 56825 3005
rect 56785 2955 56825 2985
rect 56785 2935 56795 2955
rect 56815 2935 56825 2955
rect 56785 2920 56825 2935
rect 56840 3155 56880 3170
rect 56920 3155 56960 3170
rect 56840 3135 56850 3155
rect 56870 3135 56880 3155
rect 56920 3135 56930 3155
rect 56950 3135 56960 3155
rect 56840 3105 56880 3135
rect 56920 3105 56960 3135
rect 56840 3085 56850 3105
rect 56870 3085 56880 3105
rect 56920 3085 56930 3105
rect 56950 3085 56960 3105
rect 56840 3055 56880 3085
rect 56920 3055 56960 3085
rect 56840 3035 56850 3055
rect 56870 3035 56880 3055
rect 56920 3035 56930 3055
rect 56950 3035 56960 3055
rect 56840 3005 56880 3035
rect 56920 3005 56960 3035
rect 56840 2985 56850 3005
rect 56870 2985 56880 3005
rect 56920 2985 56930 3005
rect 56950 2985 56960 3005
rect 56840 2955 56880 2985
rect 56920 2955 56960 2985
rect 56840 2935 56850 2955
rect 56870 2935 56880 2955
rect 56920 2935 56930 2955
rect 56950 2935 56960 2955
rect 56840 2920 56880 2935
rect 56920 2920 56960 2935
rect 56975 3155 57015 3170
rect 56975 3135 56985 3155
rect 57005 3135 57015 3155
rect 56975 3105 57015 3135
rect 56975 3085 56985 3105
rect 57005 3085 57015 3105
rect 56975 3055 57015 3085
rect 56975 3035 56985 3055
rect 57005 3035 57015 3055
rect 56975 3005 57015 3035
rect 56975 2985 56985 3005
rect 57005 2985 57015 3005
rect 56975 2955 57015 2985
rect 56975 2935 56985 2955
rect 57005 2935 57015 2955
rect 56975 2920 57015 2935
rect 57030 3155 57070 3170
rect 57030 3135 57040 3155
rect 57060 3135 57070 3155
rect 57030 3105 57070 3135
rect 57030 3085 57040 3105
rect 57060 3085 57070 3105
rect 57030 3055 57070 3085
rect 57030 3035 57040 3055
rect 57060 3035 57070 3055
rect 57030 3005 57070 3035
rect 57030 2985 57040 3005
rect 57060 2985 57070 3005
rect 57030 2955 57070 2985
rect 57030 2935 57040 2955
rect 57060 2935 57070 2955
rect 57030 2920 57070 2935
rect 57085 3155 57125 3170
rect 57085 3135 57095 3155
rect 57115 3135 57125 3155
rect 57085 3105 57125 3135
rect 57085 3085 57095 3105
rect 57115 3085 57125 3105
rect 57085 3055 57125 3085
rect 57085 3035 57095 3055
rect 57115 3035 57125 3055
rect 57085 3005 57125 3035
rect 57085 2985 57095 3005
rect 57115 2985 57125 3005
rect 57085 2955 57125 2985
rect 57085 2935 57095 2955
rect 57115 2935 57125 2955
rect 57085 2920 57125 2935
rect 57140 3155 57180 3170
rect 57140 3135 57150 3155
rect 57170 3135 57180 3155
rect 57140 3105 57180 3135
rect 57140 3085 57150 3105
rect 57170 3085 57180 3105
rect 57140 3055 57180 3085
rect 57140 3035 57150 3055
rect 57170 3035 57180 3055
rect 57140 3005 57180 3035
rect 57140 2985 57150 3005
rect 57170 2985 57180 3005
rect 57140 2955 57180 2985
rect 57140 2935 57150 2955
rect 57170 2935 57180 2955
rect 57140 2920 57180 2935
rect 57195 3155 57235 3170
rect 57195 3135 57205 3155
rect 57225 3135 57235 3155
rect 57195 3105 57235 3135
rect 57195 3085 57205 3105
rect 57225 3085 57235 3105
rect 57195 3055 57235 3085
rect 57195 3035 57205 3055
rect 57225 3035 57235 3055
rect 57195 3005 57235 3035
rect 57195 2985 57205 3005
rect 57225 2985 57235 3005
rect 57195 2955 57235 2985
rect 57195 2935 57205 2955
rect 57225 2935 57235 2955
rect 57195 2920 57235 2935
rect 57250 3155 57290 3170
rect 57250 3135 57260 3155
rect 57280 3135 57290 3155
rect 57250 3105 57290 3135
rect 57250 3085 57260 3105
rect 57280 3085 57290 3105
rect 57250 3055 57290 3085
rect 57250 3035 57260 3055
rect 57280 3035 57290 3055
rect 57250 3005 57290 3035
rect 57250 2985 57260 3005
rect 57280 2985 57290 3005
rect 57250 2955 57290 2985
rect 57250 2935 57260 2955
rect 57280 2935 57290 2955
rect 57250 2920 57290 2935
rect 58480 3140 58520 3155
rect 55280 2555 55320 2570
rect 58480 2570 58490 3140
rect 58510 2570 58520 3140
rect 58480 2555 58520 2570
rect 58535 3140 58575 3155
rect 58535 2570 58545 3140
rect 58565 2570 58575 3140
rect 58535 2555 58575 2570
rect 58590 3140 58630 3155
rect 58590 2570 58600 3140
rect 58620 2570 58630 3140
rect 58590 2555 58630 2570
rect 58645 3140 58685 3155
rect 58645 2570 58655 3140
rect 58675 2570 58685 3140
rect 58645 2555 58685 2570
rect 58700 3140 58740 3155
rect 58700 2570 58710 3140
rect 58730 2570 58740 3140
rect 58700 2555 58740 2570
rect 58755 3140 58795 3155
rect 58755 2570 58765 3140
rect 58785 2570 58795 3140
rect 58755 2555 58795 2570
rect 58810 3140 58850 3155
rect 58810 2570 58820 3140
rect 58840 2570 58850 3140
rect 58810 2555 58850 2570
rect 58865 3140 58905 3155
rect 58865 2570 58875 3140
rect 58895 2570 58905 3140
rect 58865 2555 58905 2570
rect 58920 3140 58960 3155
rect 58920 2570 58930 3140
rect 58950 2570 58960 3140
rect 58920 2555 58960 2570
rect 58975 3140 59015 3155
rect 58975 2570 58985 3140
rect 59005 2570 59015 3140
rect 58975 2555 59015 2570
rect 59030 3140 59070 3155
rect 59030 2570 59040 3140
rect 59060 2570 59070 3140
rect 59030 2555 59070 2570
rect 59085 3140 59125 3155
rect 59085 2570 59095 3140
rect 59115 2570 59125 3140
rect 59085 2555 59125 2570
rect 59140 3140 59180 3155
rect 59140 2570 59150 3140
rect 59170 2570 59180 3140
rect 59140 2555 59180 2570
rect 54620 1865 54660 1880
rect 54620 1695 54630 1865
rect 54650 1695 54660 1865
rect 54620 1680 54660 1695
rect 54675 1865 54715 1880
rect 54675 1695 54685 1865
rect 54705 1695 54715 1865
rect 54675 1680 54715 1695
rect 54730 1865 54770 1880
rect 54730 1695 54740 1865
rect 54760 1695 54770 1865
rect 54730 1680 54770 1695
rect 54785 1865 54825 1880
rect 54785 1695 54795 1865
rect 54815 1695 54825 1865
rect 54785 1680 54825 1695
rect 54840 1865 54880 1880
rect 54840 1695 54850 1865
rect 54870 1695 54880 1865
rect 54840 1680 54880 1695
rect 54895 1865 54935 1880
rect 54895 1695 54905 1865
rect 54925 1695 54935 1865
rect 54895 1680 54935 1695
rect 54950 1865 54990 1880
rect 54950 1695 54960 1865
rect 54980 1695 54990 1865
rect 54950 1680 54990 1695
rect 55005 1865 55045 1880
rect 55005 1695 55015 1865
rect 55035 1695 55045 1865
rect 55005 1680 55045 1695
rect 55060 1865 55100 1880
rect 55060 1695 55070 1865
rect 55090 1695 55100 1865
rect 55060 1680 55100 1695
rect 55115 1865 55155 1880
rect 55115 1695 55125 1865
rect 55145 1695 55155 1865
rect 55115 1680 55155 1695
rect 55170 1865 55210 1880
rect 55170 1695 55180 1865
rect 55200 1695 55210 1865
rect 55170 1680 55210 1695
rect 55225 1865 55265 1880
rect 55225 1695 55235 1865
rect 55255 1695 55265 1865
rect 55225 1680 55265 1695
rect 55280 1865 55320 1880
rect 55280 1695 55290 1865
rect 55310 1695 55320 1865
rect 58480 1865 58520 1880
rect 55280 1680 55320 1695
rect 58480 1695 58490 1865
rect 58510 1695 58520 1865
rect 58480 1680 58520 1695
rect 58535 1865 58575 1880
rect 58535 1695 58545 1865
rect 58565 1695 58575 1865
rect 58535 1680 58575 1695
rect 58590 1865 58630 1880
rect 58590 1695 58600 1865
rect 58620 1695 58630 1865
rect 58590 1680 58630 1695
rect 58645 1865 58685 1880
rect 58645 1695 58655 1865
rect 58675 1695 58685 1865
rect 58645 1680 58685 1695
rect 58700 1865 58740 1880
rect 58700 1695 58710 1865
rect 58730 1695 58740 1865
rect 58700 1680 58740 1695
rect 58755 1865 58795 1880
rect 58755 1695 58765 1865
rect 58785 1695 58795 1865
rect 58755 1680 58795 1695
rect 58810 1865 58850 1880
rect 58810 1695 58820 1865
rect 58840 1695 58850 1865
rect 58810 1680 58850 1695
rect 58865 1865 58905 1880
rect 58865 1695 58875 1865
rect 58895 1695 58905 1865
rect 58865 1680 58905 1695
rect 58920 1865 58960 1880
rect 58920 1695 58930 1865
rect 58950 1695 58960 1865
rect 58920 1680 58960 1695
rect 58975 1865 59015 1880
rect 58975 1695 58985 1865
rect 59005 1695 59015 1865
rect 58975 1680 59015 1695
rect 59030 1865 59070 1880
rect 59030 1695 59040 1865
rect 59060 1695 59070 1865
rect 59030 1680 59070 1695
rect 59085 1865 59125 1880
rect 59085 1695 59095 1865
rect 59115 1695 59125 1865
rect 59085 1680 59125 1695
rect 59140 1865 59180 1880
rect 59140 1695 59150 1865
rect 59170 1695 59180 1865
rect 59140 1680 59180 1695
<< ndiffc >>
rect 56780 2330 56800 2550
rect 56835 2330 56855 2550
rect 56890 2330 56910 2550
rect 56945 2330 56965 2550
rect 57000 2330 57020 2550
rect 56040 1760 56060 1880
rect 56095 1760 56115 1880
rect 56150 1760 56170 1880
rect 56205 1760 56225 1880
rect 56260 1760 56280 1880
rect 56315 1760 56335 1880
rect 56370 1760 56390 1880
rect 56425 1760 56445 1880
rect 56480 1760 56500 1880
rect 56535 1760 56555 1880
rect 56590 1760 56610 1880
rect 56645 1760 56665 1880
rect 56700 1760 56720 1880
rect 57080 1760 57100 1880
rect 57135 1760 57155 1880
rect 57190 1760 57210 1880
rect 57245 1760 57265 1880
rect 57300 1760 57320 1880
rect 57355 1760 57375 1880
rect 57410 1760 57430 1880
rect 57465 1760 57485 1880
rect 57520 1760 57540 1880
rect 57575 1760 57595 1880
rect 57630 1760 57650 1880
rect 57685 1760 57705 1880
rect 57740 1760 57760 1880
rect 54630 1155 54650 1425
rect 54685 1155 54705 1425
rect 54740 1155 54760 1425
rect 54795 1155 54815 1425
rect 54850 1155 54870 1425
rect 54905 1155 54925 1425
rect 54960 1155 54980 1425
rect 55015 1155 55035 1425
rect 55070 1155 55090 1425
rect 55125 1155 55145 1425
rect 55180 1155 55200 1425
rect 55235 1155 55255 1425
rect 55290 1155 55310 1425
rect 56040 1085 56060 1205
rect 56095 1085 56115 1205
rect 56150 1085 56170 1205
rect 56205 1085 56225 1205
rect 56260 1085 56280 1205
rect 56315 1085 56335 1205
rect 56370 1085 56390 1205
rect 56425 1085 56445 1205
rect 56480 1085 56500 1205
rect 56535 1085 56555 1205
rect 56590 1085 56610 1205
rect 56645 1085 56665 1205
rect 56700 1085 56720 1205
rect 56780 1085 56800 1205
rect 56835 1085 56855 1205
rect 56890 1085 56910 1205
rect 56945 1085 56965 1205
rect 57000 1085 57020 1205
rect 57080 1085 57100 1205
rect 57135 1085 57155 1205
rect 57190 1085 57210 1205
rect 57245 1085 57265 1205
rect 57300 1085 57320 1205
rect 57355 1085 57375 1205
rect 57410 1085 57430 1205
rect 57465 1085 57485 1205
rect 57520 1085 57540 1205
rect 57575 1085 57595 1205
rect 57630 1085 57650 1205
rect 57685 1085 57705 1205
rect 57740 1085 57760 1205
rect 58490 1155 58510 1425
rect 58545 1155 58565 1425
rect 58600 1155 58620 1425
rect 58655 1155 58675 1425
rect 58710 1155 58730 1425
rect 58765 1155 58785 1425
rect 58820 1155 58840 1425
rect 58875 1155 58895 1425
rect 58930 1155 58950 1425
rect 58985 1155 59005 1425
rect 59040 1155 59060 1425
rect 59095 1155 59115 1425
rect 59150 1155 59170 1425
rect 54660 -345 54680 325
rect 54760 -345 54780 325
rect 54860 -345 54880 325
rect 54960 -345 54980 325
rect 55060 -345 55080 325
rect 55160 -345 55180 325
rect 55260 -345 55280 325
rect 56230 185 56250 405
rect 56285 185 56305 405
rect 56340 185 56360 405
rect 56395 185 56415 405
rect 56450 185 56470 405
rect 56505 185 56525 405
rect 56560 185 56580 405
rect 56615 185 56635 405
rect 56670 185 56690 405
rect 56725 185 56745 405
rect 56780 185 56800 405
rect 56835 185 56855 405
rect 56890 185 56910 405
rect 56945 185 56965 405
rect 57000 185 57020 405
rect 57055 185 57075 405
rect 57110 185 57130 405
rect 57165 185 57185 405
rect 57220 185 57240 405
rect 57275 185 57295 405
rect 57330 185 57350 405
rect 57385 185 57405 405
rect 57440 185 57460 405
rect 57495 185 57515 405
rect 56440 -435 56460 -315
rect 56495 -435 56515 -315
rect 56550 -435 56570 -315
rect 56605 -435 56625 -315
rect 56660 -435 56680 -315
rect 56715 -435 56735 -315
rect 56770 -435 56790 -315
rect 56880 -435 56900 -315
rect 57220 -425 57240 -325
rect 58520 -345 58540 325
rect 58620 -345 58640 325
rect 58720 -345 58740 325
rect 58820 -345 58840 325
rect 58920 -345 58940 325
rect 59020 -345 59040 325
rect 59120 -345 59140 325
<< pdiffc >>
rect 56095 4545 56115 4865
rect 56155 4545 56175 4865
rect 56215 4545 56235 4865
rect 56275 4545 56295 4865
rect 56565 4545 56585 4695
rect 56625 4545 56645 4695
rect 56685 4545 56705 4695
rect 56745 4545 56765 4695
rect 57035 4545 57055 4865
rect 57095 4545 57115 4865
rect 57155 4545 57175 4865
rect 57215 4545 57235 4865
rect 57505 4545 57525 4865
rect 57565 4545 57585 4865
rect 57625 4545 57645 4865
rect 57685 4545 57705 4865
rect 54600 3680 54620 4000
rect 54660 3680 54680 4000
rect 54720 3680 54740 4000
rect 54780 3680 54800 4000
rect 54840 3680 54860 4000
rect 54900 3680 54920 4000
rect 54960 3680 54980 4000
rect 55020 3680 55040 4000
rect 55080 3680 55100 4000
rect 55140 3680 55160 4000
rect 55200 3680 55220 4000
rect 55260 3680 55280 4000
rect 55320 3680 55340 4000
rect 56015 3680 56035 4000
rect 56075 3680 56095 4000
rect 56135 3680 56155 4000
rect 56195 3680 56215 4000
rect 56255 3680 56275 4000
rect 56315 3680 56335 4000
rect 56375 3680 56395 4000
rect 56435 3680 56455 4000
rect 56495 3680 56515 4000
rect 56555 3680 56575 4000
rect 56615 3680 56635 4000
rect 56675 3680 56695 4000
rect 56735 3680 56755 4000
rect 57045 3680 57065 4000
rect 57105 3680 57125 4000
rect 57165 3680 57185 4000
rect 57225 3680 57245 4000
rect 57285 3680 57305 4000
rect 57345 3680 57365 4000
rect 57405 3680 57425 4000
rect 57465 3680 57485 4000
rect 57525 3680 57545 4000
rect 57585 3680 57605 4000
rect 57645 3680 57665 4000
rect 57705 3680 57725 4000
rect 57765 3680 57785 4000
rect 58460 3680 58480 4000
rect 58520 3680 58540 4000
rect 58580 3680 58600 4000
rect 58640 3680 58660 4000
rect 58700 3680 58720 4000
rect 58760 3680 58780 4000
rect 58820 3680 58840 4000
rect 58880 3680 58900 4000
rect 58940 3680 58960 4000
rect 59000 3680 59020 4000
rect 59060 3680 59080 4000
rect 59120 3680 59140 4000
rect 59180 3680 59200 4000
rect 54630 2570 54650 3140
rect 54685 2570 54705 3140
rect 54740 2570 54760 3140
rect 54795 2570 54815 3140
rect 54850 2570 54870 3140
rect 54905 2570 54925 3140
rect 54960 2570 54980 3140
rect 55015 2570 55035 3140
rect 55070 2570 55090 3140
rect 55125 2570 55145 3140
rect 55180 2570 55200 3140
rect 55235 2570 55255 3140
rect 55290 2570 55310 3140
rect 56520 3135 56540 3155
rect 56520 3085 56540 3105
rect 56520 3035 56540 3055
rect 56520 2985 56540 3005
rect 56520 2935 56540 2955
rect 56575 3135 56595 3155
rect 56575 3085 56595 3105
rect 56575 3035 56595 3055
rect 56575 2985 56595 3005
rect 56575 2935 56595 2955
rect 56630 3135 56650 3155
rect 56630 3085 56650 3105
rect 56630 3035 56650 3055
rect 56630 2985 56650 3005
rect 56630 2935 56650 2955
rect 56685 3135 56705 3155
rect 56685 3085 56705 3105
rect 56685 3035 56705 3055
rect 56685 2985 56705 3005
rect 56685 2935 56705 2955
rect 56740 3135 56760 3155
rect 56740 3085 56760 3105
rect 56740 3035 56760 3055
rect 56740 2985 56760 3005
rect 56740 2935 56760 2955
rect 56795 3135 56815 3155
rect 56795 3085 56815 3105
rect 56795 3035 56815 3055
rect 56795 2985 56815 3005
rect 56795 2935 56815 2955
rect 56850 3135 56870 3155
rect 56930 3135 56950 3155
rect 56850 3085 56870 3105
rect 56930 3085 56950 3105
rect 56850 3035 56870 3055
rect 56930 3035 56950 3055
rect 56850 2985 56870 3005
rect 56930 2985 56950 3005
rect 56850 2935 56870 2955
rect 56930 2935 56950 2955
rect 56985 3135 57005 3155
rect 56985 3085 57005 3105
rect 56985 3035 57005 3055
rect 56985 2985 57005 3005
rect 56985 2935 57005 2955
rect 57040 3135 57060 3155
rect 57040 3085 57060 3105
rect 57040 3035 57060 3055
rect 57040 2985 57060 3005
rect 57040 2935 57060 2955
rect 57095 3135 57115 3155
rect 57095 3085 57115 3105
rect 57095 3035 57115 3055
rect 57095 2985 57115 3005
rect 57095 2935 57115 2955
rect 57150 3135 57170 3155
rect 57150 3085 57170 3105
rect 57150 3035 57170 3055
rect 57150 2985 57170 3005
rect 57150 2935 57170 2955
rect 57205 3135 57225 3155
rect 57205 3085 57225 3105
rect 57205 3035 57225 3055
rect 57205 2985 57225 3005
rect 57205 2935 57225 2955
rect 57260 3135 57280 3155
rect 57260 3085 57280 3105
rect 57260 3035 57280 3055
rect 57260 2985 57280 3005
rect 57260 2935 57280 2955
rect 58490 2570 58510 3140
rect 58545 2570 58565 3140
rect 58600 2570 58620 3140
rect 58655 2570 58675 3140
rect 58710 2570 58730 3140
rect 58765 2570 58785 3140
rect 58820 2570 58840 3140
rect 58875 2570 58895 3140
rect 58930 2570 58950 3140
rect 58985 2570 59005 3140
rect 59040 2570 59060 3140
rect 59095 2570 59115 3140
rect 59150 2570 59170 3140
rect 54630 1695 54650 1865
rect 54685 1695 54705 1865
rect 54740 1695 54760 1865
rect 54795 1695 54815 1865
rect 54850 1695 54870 1865
rect 54905 1695 54925 1865
rect 54960 1695 54980 1865
rect 55015 1695 55035 1865
rect 55070 1695 55090 1865
rect 55125 1695 55145 1865
rect 55180 1695 55200 1865
rect 55235 1695 55255 1865
rect 55290 1695 55310 1865
rect 58490 1695 58510 1865
rect 58545 1695 58565 1865
rect 58600 1695 58620 1865
rect 58655 1695 58675 1865
rect 58710 1695 58730 1865
rect 58765 1695 58785 1865
rect 58820 1695 58840 1865
rect 58875 1695 58895 1865
rect 58930 1695 58950 1865
rect 58985 1695 59005 1865
rect 59040 1695 59060 1865
rect 59095 1695 59115 1865
rect 59150 1695 59170 1865
<< psubdiff >>
rect 56730 2550 56770 2565
rect 56730 2330 56740 2550
rect 56760 2330 56770 2550
rect 56730 2315 56770 2330
rect 57030 2550 57070 2565
rect 57030 2330 57040 2550
rect 57060 2330 57070 2550
rect 57030 2315 57070 2330
rect 55990 1880 56030 1895
rect 55990 1760 56000 1880
rect 56020 1760 56030 1880
rect 55990 1745 56030 1760
rect 56730 1880 56770 1895
rect 56730 1760 56740 1880
rect 56760 1760 56770 1880
rect 56730 1745 56770 1760
rect 57030 1880 57070 1895
rect 57030 1760 57040 1880
rect 57060 1760 57070 1880
rect 57030 1745 57070 1760
rect 57770 1880 57810 1895
rect 57770 1760 57780 1880
rect 57800 1760 57810 1880
rect 57770 1745 57810 1760
rect 54580 1425 54620 1440
rect 54580 1155 54590 1425
rect 54610 1155 54620 1425
rect 54580 1140 54620 1155
rect 55320 1425 55360 1440
rect 55320 1155 55330 1425
rect 55350 1155 55360 1425
rect 58440 1425 58480 1440
rect 55320 1140 55360 1155
rect 55990 1205 56030 1220
rect 55990 1085 56000 1205
rect 56020 1085 56030 1205
rect 55990 1070 56030 1085
rect 56730 1205 56770 1220
rect 56730 1085 56740 1205
rect 56760 1085 56770 1205
rect 56730 1070 56770 1085
rect 57030 1205 57070 1220
rect 57030 1085 57040 1205
rect 57060 1085 57070 1205
rect 57030 1070 57070 1085
rect 57770 1205 57810 1220
rect 57770 1085 57780 1205
rect 57800 1085 57810 1205
rect 58440 1155 58450 1425
rect 58470 1155 58480 1425
rect 58440 1140 58480 1155
rect 59180 1425 59220 1440
rect 59180 1155 59190 1425
rect 59210 1155 59220 1425
rect 59180 1140 59220 1155
rect 57770 1070 57810 1085
rect 56180 405 56220 420
rect 54610 325 54650 340
rect 54610 -345 54620 325
rect 54640 -345 54650 325
rect 54610 -360 54650 -345
rect 55290 325 55330 340
rect 55290 -345 55300 325
rect 55320 -345 55330 325
rect 56180 185 56190 405
rect 56210 185 56220 405
rect 56180 170 56220 185
rect 57525 405 57565 420
rect 57525 185 57535 405
rect 57555 185 57565 405
rect 57525 170 57565 185
rect 58470 325 58510 340
rect 55290 -360 55330 -345
rect 56390 -315 56430 -300
rect 56390 -435 56400 -315
rect 56420 -435 56430 -315
rect 56390 -450 56430 -435
rect 56800 -315 56840 -300
rect 56800 -435 56810 -315
rect 56830 -435 56840 -315
rect 56800 -450 56840 -435
rect 58470 -345 58480 325
rect 58500 -345 58510 325
rect 58470 -360 58510 -345
rect 59150 325 59190 340
rect 59150 -345 59160 325
rect 59180 -345 59190 325
rect 59150 -360 59190 -345
<< nsubdiff >>
rect 56045 4865 56085 4880
rect 56045 4545 56055 4865
rect 56075 4545 56085 4865
rect 56045 4530 56085 4545
rect 56305 4865 56345 4880
rect 56305 4545 56315 4865
rect 56335 4545 56345 4865
rect 56985 4865 57025 4880
rect 56305 4530 56345 4545
rect 56515 4695 56555 4710
rect 56515 4545 56525 4695
rect 56545 4545 56555 4695
rect 56515 4530 56555 4545
rect 56775 4695 56815 4710
rect 56775 4545 56785 4695
rect 56805 4545 56815 4695
rect 56775 4530 56815 4545
rect 56985 4545 56995 4865
rect 57015 4545 57025 4865
rect 56985 4530 57025 4545
rect 57245 4865 57285 4880
rect 57245 4545 57255 4865
rect 57275 4545 57285 4865
rect 57245 4530 57285 4545
rect 57455 4865 57495 4880
rect 57455 4545 57465 4865
rect 57485 4545 57495 4865
rect 57455 4530 57495 4545
rect 57715 4865 57755 4880
rect 57715 4545 57725 4865
rect 57745 4545 57755 4865
rect 57715 4530 57755 4545
rect 54550 4000 54590 4015
rect 54550 3680 54560 4000
rect 54580 3680 54590 4000
rect 54550 3665 54590 3680
rect 55350 4000 55390 4015
rect 55350 3680 55360 4000
rect 55380 3680 55390 4000
rect 55350 3665 55390 3680
rect 55965 4000 56005 4015
rect 55965 3680 55975 4000
rect 55995 3680 56005 4000
rect 55965 3665 56005 3680
rect 56765 4000 56805 4015
rect 56765 3680 56775 4000
rect 56795 3680 56805 4000
rect 56765 3665 56805 3680
rect 56995 4000 57035 4015
rect 56995 3680 57005 4000
rect 57025 3680 57035 4000
rect 56995 3665 57035 3680
rect 57795 4000 57835 4015
rect 57795 3680 57805 4000
rect 57825 3680 57835 4000
rect 57795 3665 57835 3680
rect 58410 4000 58450 4015
rect 58410 3680 58420 4000
rect 58440 3680 58450 4000
rect 58410 3665 58450 3680
rect 59210 4000 59250 4015
rect 59210 3680 59220 4000
rect 59240 3680 59250 4000
rect 59210 3665 59250 3680
rect 56470 3155 56510 3170
rect 54580 3140 54620 3155
rect 54580 2570 54590 3140
rect 54610 2570 54620 3140
rect 54580 2555 54620 2570
rect 55320 3140 55360 3155
rect 55320 2570 55330 3140
rect 55350 2570 55360 3140
rect 56470 3135 56480 3155
rect 56500 3135 56510 3155
rect 56470 3105 56510 3135
rect 56470 3085 56480 3105
rect 56500 3085 56510 3105
rect 56470 3055 56510 3085
rect 56470 3035 56480 3055
rect 56500 3035 56510 3055
rect 56470 3005 56510 3035
rect 56470 2985 56480 3005
rect 56500 2985 56510 3005
rect 56470 2955 56510 2985
rect 56470 2935 56480 2955
rect 56500 2935 56510 2955
rect 56470 2920 56510 2935
rect 56880 3155 56920 3170
rect 56880 3135 56890 3155
rect 56910 3135 56920 3155
rect 56880 3105 56920 3135
rect 56880 3085 56890 3105
rect 56910 3085 56920 3105
rect 56880 3055 56920 3085
rect 56880 3035 56890 3055
rect 56910 3035 56920 3055
rect 56880 3005 56920 3035
rect 56880 2985 56890 3005
rect 56910 2985 56920 3005
rect 56880 2955 56920 2985
rect 56880 2935 56890 2955
rect 56910 2935 56920 2955
rect 56880 2920 56920 2935
rect 57290 3155 57330 3170
rect 57290 3135 57300 3155
rect 57320 3135 57330 3155
rect 57290 3105 57330 3135
rect 57290 3085 57300 3105
rect 57320 3085 57330 3105
rect 57290 3055 57330 3085
rect 57290 3035 57300 3055
rect 57320 3035 57330 3055
rect 57290 3005 57330 3035
rect 57290 2985 57300 3005
rect 57320 2985 57330 3005
rect 57290 2955 57330 2985
rect 57290 2935 57300 2955
rect 57320 2935 57330 2955
rect 57290 2920 57330 2935
rect 58440 3140 58480 3155
rect 55320 2555 55360 2570
rect 58440 2570 58450 3140
rect 58470 2570 58480 3140
rect 58440 2555 58480 2570
rect 59180 3140 59220 3155
rect 59180 2570 59190 3140
rect 59210 2570 59220 3140
rect 59180 2555 59220 2570
rect 54580 1865 54620 1880
rect 54580 1695 54590 1865
rect 54610 1695 54620 1865
rect 54580 1680 54620 1695
rect 55320 1865 55360 1880
rect 55320 1695 55330 1865
rect 55350 1695 55360 1865
rect 58440 1865 58480 1880
rect 55320 1680 55360 1695
rect 58440 1695 58450 1865
rect 58470 1695 58480 1865
rect 58440 1680 58480 1695
rect 59180 1865 59220 1880
rect 59180 1695 59190 1865
rect 59210 1695 59220 1865
rect 59180 1680 59220 1695
<< psubdiffcont >>
rect 56740 2330 56760 2550
rect 57040 2330 57060 2550
rect 56000 1760 56020 1880
rect 56740 1760 56760 1880
rect 57040 1760 57060 1880
rect 57780 1760 57800 1880
rect 54590 1155 54610 1425
rect 55330 1155 55350 1425
rect 56000 1085 56020 1205
rect 56740 1085 56760 1205
rect 57040 1085 57060 1205
rect 57780 1085 57800 1205
rect 58450 1155 58470 1425
rect 59190 1155 59210 1425
rect 54620 -345 54640 325
rect 55300 -345 55320 325
rect 56190 185 56210 405
rect 57535 185 57555 405
rect 56400 -435 56420 -315
rect 56810 -435 56830 -315
rect 58480 -345 58500 325
rect 59160 -345 59180 325
<< nsubdiffcont >>
rect 56055 4545 56075 4865
rect 56315 4545 56335 4865
rect 56525 4545 56545 4695
rect 56785 4545 56805 4695
rect 56995 4545 57015 4865
rect 57255 4545 57275 4865
rect 57465 4545 57485 4865
rect 57725 4545 57745 4865
rect 54560 3680 54580 4000
rect 55360 3680 55380 4000
rect 55975 3680 55995 4000
rect 56775 3680 56795 4000
rect 57005 3680 57025 4000
rect 57805 3680 57825 4000
rect 58420 3680 58440 4000
rect 59220 3680 59240 4000
rect 54590 2570 54610 3140
rect 55330 2570 55350 3140
rect 56480 3135 56500 3155
rect 56480 3085 56500 3105
rect 56480 3035 56500 3055
rect 56480 2985 56500 3005
rect 56480 2935 56500 2955
rect 56890 3135 56910 3155
rect 56890 3085 56910 3105
rect 56890 3035 56910 3055
rect 56890 2985 56910 3005
rect 56890 2935 56910 2955
rect 57300 3135 57320 3155
rect 57300 3085 57320 3105
rect 57300 3035 57320 3055
rect 57300 2985 57320 3005
rect 57300 2935 57320 2955
rect 58450 2570 58470 3140
rect 59190 2570 59210 3140
rect 54590 1695 54610 1865
rect 55330 1695 55350 1865
rect 58450 1695 58470 1865
rect 59190 1695 59210 1865
<< poly >>
rect 56085 4925 56125 4935
rect 56085 4905 56095 4925
rect 56115 4910 56125 4925
rect 56265 4925 56305 4935
rect 56265 4910 56275 4925
rect 56115 4905 56145 4910
rect 56085 4895 56145 4905
rect 56245 4905 56275 4910
rect 56295 4905 56305 4925
rect 56245 4895 56305 4905
rect 57025 4925 57065 4935
rect 57025 4905 57035 4925
rect 57055 4910 57065 4925
rect 57205 4925 57245 4935
rect 57205 4910 57215 4925
rect 57055 4905 57085 4910
rect 57025 4895 57085 4905
rect 57185 4905 57215 4910
rect 57235 4905 57245 4925
rect 57185 4895 57245 4905
rect 57495 4925 57535 4935
rect 57495 4905 57505 4925
rect 57525 4910 57535 4925
rect 57675 4925 57715 4935
rect 57675 4910 57685 4925
rect 57525 4905 57555 4910
rect 57495 4895 57555 4905
rect 57655 4905 57685 4910
rect 57705 4905 57715 4925
rect 57655 4895 57715 4905
rect 56125 4880 56145 4895
rect 56185 4880 56205 4895
rect 56245 4880 56265 4895
rect 57065 4880 57085 4895
rect 57125 4880 57145 4895
rect 57185 4880 57205 4895
rect 57535 4880 57555 4895
rect 57595 4880 57615 4895
rect 57655 4880 57675 4895
rect 56555 4755 56595 4765
rect 56555 4735 56565 4755
rect 56585 4740 56595 4755
rect 56735 4755 56775 4765
rect 56735 4740 56745 4755
rect 56585 4735 56615 4740
rect 56555 4725 56615 4735
rect 56715 4735 56745 4740
rect 56765 4735 56775 4755
rect 56715 4725 56775 4735
rect 56595 4710 56615 4725
rect 56655 4710 56675 4725
rect 56715 4710 56735 4725
rect 56125 4515 56145 4530
rect 56185 4485 56205 4530
rect 56245 4515 56265 4530
rect 56595 4515 56615 4530
rect 56655 4485 56675 4530
rect 56715 4515 56735 4530
rect 57065 4515 57085 4530
rect 56150 4475 56205 4485
rect 56150 4455 56160 4475
rect 56180 4455 56205 4475
rect 56150 4445 56205 4455
rect 56630 4475 56675 4485
rect 56630 4455 56635 4475
rect 56655 4470 56675 4475
rect 57125 4485 57145 4530
rect 57185 4515 57205 4530
rect 57535 4515 57555 4530
rect 57125 4475 57170 4485
rect 57595 4475 57615 4530
rect 57655 4515 57675 4530
rect 57125 4470 57145 4475
rect 56655 4455 56660 4470
rect 56630 4445 56660 4455
rect 57140 4455 57145 4470
rect 57165 4455 57170 4475
rect 57140 4445 57170 4455
rect 57576 4465 57615 4475
rect 57576 4445 57581 4465
rect 57601 4460 57615 4465
rect 57601 4445 57606 4460
rect 57576 4435 57606 4445
rect 54630 4015 54650 4030
rect 54690 4015 54710 4030
rect 54750 4015 54770 4030
rect 54810 4015 54830 4030
rect 54870 4015 54890 4030
rect 54930 4015 54950 4030
rect 54990 4015 55010 4030
rect 55050 4015 55070 4030
rect 55110 4015 55130 4030
rect 55170 4015 55190 4030
rect 55230 4015 55250 4030
rect 55290 4015 55310 4030
rect 56045 4015 56065 4030
rect 56105 4015 56125 4030
rect 56165 4015 56185 4030
rect 56225 4015 56245 4030
rect 56285 4015 56305 4030
rect 56345 4015 56365 4030
rect 56405 4015 56425 4030
rect 56465 4015 56485 4030
rect 56525 4015 56545 4030
rect 56585 4015 56605 4030
rect 56645 4015 56665 4030
rect 56705 4015 56725 4030
rect 57075 4015 57095 4030
rect 57135 4015 57155 4030
rect 57195 4015 57215 4030
rect 57255 4015 57275 4030
rect 57315 4015 57335 4030
rect 57375 4015 57395 4030
rect 57435 4015 57455 4030
rect 57495 4015 57515 4030
rect 57555 4015 57575 4030
rect 57615 4015 57635 4030
rect 57675 4015 57695 4030
rect 57735 4015 57755 4030
rect 58490 4015 58510 4030
rect 58550 4015 58570 4030
rect 58610 4015 58630 4030
rect 58670 4015 58690 4030
rect 58730 4015 58750 4030
rect 58790 4015 58810 4030
rect 58850 4015 58870 4030
rect 58910 4015 58930 4030
rect 58970 4015 58990 4030
rect 59030 4015 59050 4030
rect 59090 4015 59110 4030
rect 59150 4015 59170 4030
rect 54630 3650 54650 3665
rect 54595 3640 54650 3650
rect 54690 3655 54710 3665
rect 54750 3655 54770 3665
rect 54810 3655 54830 3665
rect 54870 3655 54890 3665
rect 54930 3655 54950 3665
rect 54990 3655 55010 3665
rect 55050 3655 55070 3665
rect 55110 3655 55130 3665
rect 55170 3655 55190 3665
rect 55230 3655 55250 3665
rect 54690 3640 55250 3655
rect 55290 3650 55310 3665
rect 56045 3650 56065 3665
rect 55290 3640 55345 3650
rect 54595 3620 54600 3640
rect 54620 3635 54650 3640
rect 54620 3620 54625 3635
rect 54595 3610 54625 3620
rect 54955 3620 54960 3640
rect 54980 3620 54985 3640
rect 55290 3635 55320 3640
rect 54955 3610 54985 3620
rect 55315 3620 55320 3635
rect 55340 3620 55345 3640
rect 55315 3610 55345 3620
rect 56010 3640 56065 3650
rect 56105 3655 56125 3665
rect 56165 3655 56185 3665
rect 56225 3655 56245 3665
rect 56285 3655 56305 3665
rect 56345 3655 56365 3665
rect 56405 3655 56425 3665
rect 56465 3655 56485 3665
rect 56525 3655 56545 3665
rect 56585 3655 56605 3665
rect 56645 3655 56665 3665
rect 56105 3640 56665 3655
rect 56705 3650 56725 3665
rect 57075 3650 57095 3665
rect 56705 3640 56760 3650
rect 56010 3620 56015 3640
rect 56035 3635 56065 3640
rect 56035 3620 56040 3635
rect 56010 3610 56040 3620
rect 56370 3620 56375 3640
rect 56395 3620 56400 3640
rect 56705 3635 56735 3640
rect 56370 3610 56400 3620
rect 56730 3620 56735 3635
rect 56755 3620 56760 3640
rect 56730 3610 56760 3620
rect 57040 3640 57095 3650
rect 57135 3655 57155 3665
rect 57195 3655 57215 3665
rect 57255 3655 57275 3665
rect 57315 3655 57335 3665
rect 57375 3655 57395 3665
rect 57435 3655 57455 3665
rect 57495 3655 57515 3665
rect 57555 3655 57575 3665
rect 57615 3655 57635 3665
rect 57675 3655 57695 3665
rect 57135 3640 57695 3655
rect 57735 3650 57755 3665
rect 58490 3650 58510 3665
rect 57735 3640 57790 3650
rect 57040 3620 57045 3640
rect 57065 3635 57095 3640
rect 57065 3620 57070 3635
rect 57040 3610 57070 3620
rect 57400 3620 57405 3640
rect 57425 3620 57430 3640
rect 57735 3635 57765 3640
rect 57400 3610 57430 3620
rect 57760 3620 57765 3635
rect 57785 3620 57790 3640
rect 57760 3610 57790 3620
rect 58455 3640 58510 3650
rect 58550 3655 58570 3665
rect 58610 3655 58630 3665
rect 58670 3655 58690 3665
rect 58730 3655 58750 3665
rect 58790 3655 58810 3665
rect 58850 3655 58870 3665
rect 58910 3655 58930 3665
rect 58970 3655 58990 3665
rect 59030 3655 59050 3665
rect 59090 3655 59110 3665
rect 58550 3640 59110 3655
rect 59150 3650 59170 3665
rect 59150 3640 59205 3650
rect 58455 3620 58460 3640
rect 58480 3635 58510 3640
rect 58480 3620 58485 3635
rect 58455 3610 58485 3620
rect 58815 3620 58820 3640
rect 58840 3620 58845 3640
rect 59150 3635 59180 3640
rect 58815 3610 58845 3620
rect 59175 3620 59180 3635
rect 59200 3620 59205 3640
rect 59175 3610 59205 3620
rect 54960 3540 54980 3610
rect 56375 3585 56395 3610
rect 57405 3585 57425 3610
rect 56365 3575 56405 3585
rect 56365 3555 56375 3575
rect 56395 3555 56405 3575
rect 56365 3545 56405 3555
rect 57395 3575 57435 3585
rect 57395 3555 57405 3575
rect 57425 3555 57435 3575
rect 57395 3545 57435 3555
rect 58820 3540 58840 3610
rect 54950 3530 54990 3540
rect 54950 3510 54960 3530
rect 54980 3510 54990 3530
rect 54950 3500 54990 3510
rect 58810 3530 58850 3540
rect 58810 3510 58820 3530
rect 58840 3510 58850 3530
rect 58810 3500 58850 3510
rect 56510 3270 56550 3280
rect 56510 3250 56520 3270
rect 56540 3255 56550 3270
rect 56840 3270 56880 3280
rect 56840 3255 56850 3270
rect 56540 3250 56565 3255
rect 56510 3240 56565 3250
rect 54625 3200 54655 3210
rect 54625 3180 54630 3200
rect 54650 3185 54655 3200
rect 55285 3200 55315 3210
rect 55285 3185 55290 3200
rect 54650 3180 54675 3185
rect 54625 3170 54675 3180
rect 55265 3180 55290 3185
rect 55310 3180 55315 3200
rect 55265 3170 55315 3180
rect 56550 3170 56565 3240
rect 56825 3250 56850 3255
rect 56870 3250 56880 3270
rect 56825 3240 56880 3250
rect 56920 3270 56960 3280
rect 56920 3250 56930 3270
rect 56950 3255 56960 3270
rect 57250 3270 57290 3280
rect 57250 3255 57260 3270
rect 56950 3250 56975 3255
rect 56920 3240 56975 3250
rect 56605 3170 56620 3185
rect 56660 3170 56675 3185
rect 56715 3170 56730 3185
rect 56770 3170 56785 3185
rect 56825 3170 56840 3240
rect 56960 3170 56975 3240
rect 57235 3250 57260 3255
rect 57280 3250 57290 3270
rect 57235 3240 57290 3250
rect 57015 3170 57030 3185
rect 57070 3170 57085 3185
rect 57125 3170 57140 3185
rect 57180 3170 57195 3185
rect 57235 3170 57250 3240
rect 58485 3200 58515 3210
rect 58485 3180 58490 3200
rect 58510 3185 58515 3200
rect 59145 3200 59175 3210
rect 59145 3185 59150 3200
rect 58510 3180 58535 3185
rect 58485 3170 58535 3180
rect 59125 3180 59150 3185
rect 59170 3180 59175 3200
rect 59125 3170 59175 3180
rect 54660 3155 54675 3170
rect 54715 3155 54730 3170
rect 54770 3155 54785 3170
rect 54825 3155 54840 3170
rect 54880 3155 54895 3170
rect 54935 3155 54950 3170
rect 54990 3155 55005 3170
rect 55045 3155 55060 3170
rect 55100 3155 55115 3170
rect 55155 3155 55170 3170
rect 55210 3155 55225 3170
rect 55265 3155 55280 3170
rect 58520 3155 58535 3170
rect 58575 3155 58590 3170
rect 58630 3155 58645 3170
rect 58685 3155 58700 3170
rect 58740 3155 58755 3170
rect 58795 3155 58810 3170
rect 58850 3155 58865 3170
rect 58905 3155 58920 3170
rect 58960 3155 58975 3170
rect 59015 3155 59030 3170
rect 59070 3155 59085 3170
rect 59125 3155 59140 3170
rect 56550 2905 56565 2920
rect 56605 2905 56620 2920
rect 56660 2910 56675 2920
rect 56715 2910 56730 2920
rect 56605 2895 56637 2905
rect 56660 2895 56730 2910
rect 56770 2905 56785 2920
rect 56825 2905 56840 2920
rect 56960 2905 56975 2920
rect 57015 2905 57030 2920
rect 57070 2910 57085 2920
rect 57125 2910 57140 2920
rect 56753 2895 56785 2905
rect 57015 2895 57047 2905
rect 57070 2895 57140 2910
rect 57180 2905 57195 2920
rect 57235 2905 57250 2920
rect 57163 2895 57195 2905
rect 56607 2875 56612 2895
rect 56632 2875 56637 2895
rect 56607 2865 56637 2875
rect 56675 2875 56685 2895
rect 56705 2875 56715 2895
rect 56675 2865 56715 2875
rect 56753 2875 56758 2895
rect 56778 2875 56783 2895
rect 56753 2865 56783 2875
rect 57017 2875 57022 2895
rect 57042 2875 57047 2895
rect 57017 2865 57047 2875
rect 57085 2875 57095 2895
rect 57115 2875 57125 2895
rect 57085 2865 57125 2875
rect 57163 2875 57168 2895
rect 57188 2875 57193 2895
rect 57163 2865 57193 2875
rect 56850 2610 56890 2620
rect 56850 2590 56860 2610
rect 56880 2590 56890 2610
rect 56850 2580 56935 2590
rect 56810 2565 56825 2580
rect 56865 2575 56935 2580
rect 56865 2565 56880 2575
rect 56920 2565 56935 2575
rect 56975 2565 56990 2580
rect 54660 2540 54675 2555
rect 54715 2545 54730 2555
rect 54770 2545 54785 2555
rect 54825 2545 54840 2555
rect 54880 2545 54895 2555
rect 54935 2545 54950 2555
rect 54990 2545 55005 2555
rect 55045 2545 55060 2555
rect 55100 2545 55115 2555
rect 55155 2545 55170 2555
rect 55210 2545 55225 2555
rect 54715 2530 55225 2545
rect 55265 2540 55280 2555
rect 54955 2510 54960 2530
rect 54980 2510 54985 2530
rect 54955 2475 54985 2510
rect 54950 2465 54990 2475
rect 54950 2445 54960 2465
rect 54980 2445 54990 2465
rect 54950 2425 54990 2445
rect 54950 2405 54960 2425
rect 54980 2405 54990 2425
rect 54950 2385 54990 2405
rect 54950 2365 54960 2385
rect 54980 2365 54990 2385
rect 54950 2355 54990 2365
rect 58520 2540 58535 2555
rect 58575 2545 58590 2555
rect 58630 2545 58645 2555
rect 58685 2545 58700 2555
rect 58740 2545 58755 2555
rect 58795 2545 58810 2555
rect 58850 2545 58865 2555
rect 58905 2545 58920 2555
rect 58960 2545 58975 2555
rect 59015 2545 59030 2555
rect 59070 2545 59085 2555
rect 58575 2530 59085 2545
rect 59125 2540 59140 2555
rect 58815 2510 58820 2530
rect 58840 2510 58845 2530
rect 58815 2475 58845 2510
rect 58810 2465 58850 2475
rect 58810 2445 58820 2465
rect 58840 2445 58850 2465
rect 58810 2425 58850 2445
rect 58810 2405 58820 2425
rect 58840 2405 58850 2425
rect 58810 2385 58850 2405
rect 58810 2365 58820 2385
rect 58840 2365 58850 2385
rect 58810 2355 58850 2365
rect 56810 2300 56825 2315
rect 56865 2300 56880 2315
rect 56920 2300 56935 2315
rect 56975 2300 56990 2315
rect 56770 2290 56825 2300
rect 56770 2270 56780 2290
rect 56800 2285 56825 2290
rect 56975 2290 57030 2300
rect 56975 2285 57000 2290
rect 56800 2270 56810 2285
rect 56770 2260 56810 2270
rect 56990 2270 57000 2285
rect 57020 2270 57030 2290
rect 56990 2260 57030 2270
rect 56040 1980 56070 1990
rect 56040 1960 56045 1980
rect 56065 1965 56070 1980
rect 56690 1980 56720 1990
rect 56690 1965 56695 1980
rect 56065 1960 56140 1965
rect 56040 1950 56140 1960
rect 54625 1925 54655 1935
rect 54625 1905 54630 1925
rect 54650 1910 54655 1925
rect 55285 1925 55315 1935
rect 55285 1910 55290 1925
rect 54650 1905 54675 1910
rect 54625 1895 54675 1905
rect 55265 1905 55290 1910
rect 55310 1905 55315 1925
rect 56125 1920 56140 1950
rect 56620 1960 56695 1965
rect 56715 1960 56720 1980
rect 56620 1950 56720 1960
rect 57080 1980 57110 1990
rect 57080 1960 57085 1980
rect 57105 1965 57110 1980
rect 57730 1980 57760 1990
rect 57730 1965 57735 1980
rect 57105 1960 57180 1965
rect 57080 1950 57180 1960
rect 56620 1920 56635 1950
rect 55265 1895 55315 1905
rect 56070 1895 56085 1910
rect 56125 1905 56635 1920
rect 57165 1920 57180 1950
rect 57660 1960 57735 1965
rect 57755 1960 57760 1980
rect 57660 1950 57760 1960
rect 57660 1920 57675 1950
rect 56125 1895 56140 1905
rect 56180 1895 56195 1905
rect 56235 1895 56250 1905
rect 56290 1895 56305 1905
rect 56345 1895 56360 1905
rect 56400 1895 56415 1905
rect 56455 1895 56470 1905
rect 56510 1895 56525 1905
rect 56565 1895 56580 1905
rect 56620 1895 56635 1905
rect 56675 1895 56690 1910
rect 57110 1895 57125 1910
rect 57165 1905 57675 1920
rect 58485 1925 58515 1935
rect 57165 1895 57180 1905
rect 57220 1895 57235 1905
rect 57275 1895 57290 1905
rect 57330 1895 57345 1905
rect 57385 1895 57400 1905
rect 57440 1895 57455 1905
rect 57495 1895 57510 1905
rect 57550 1895 57565 1905
rect 57605 1895 57620 1905
rect 57660 1895 57675 1905
rect 57715 1895 57730 1910
rect 58485 1905 58490 1925
rect 58510 1910 58515 1925
rect 59145 1925 59175 1935
rect 59145 1910 59150 1925
rect 58510 1905 58535 1910
rect 58485 1895 58535 1905
rect 59125 1905 59150 1910
rect 59170 1905 59175 1925
rect 59125 1895 59175 1905
rect 54660 1880 54675 1895
rect 54715 1880 54730 1895
rect 54770 1880 54785 1895
rect 54825 1880 54840 1895
rect 54880 1880 54895 1895
rect 54935 1880 54950 1895
rect 54990 1880 55005 1895
rect 55045 1880 55060 1895
rect 55100 1880 55115 1895
rect 55155 1880 55170 1895
rect 55210 1880 55225 1895
rect 55265 1880 55280 1895
rect 58520 1880 58535 1895
rect 58575 1880 58590 1895
rect 58630 1880 58645 1895
rect 58685 1880 58700 1895
rect 58740 1880 58755 1895
rect 58795 1880 58810 1895
rect 58850 1880 58865 1895
rect 58905 1880 58920 1895
rect 58960 1880 58975 1895
rect 59015 1880 59030 1895
rect 59070 1880 59085 1895
rect 59125 1880 59140 1895
rect 56070 1730 56085 1745
rect 56125 1730 56140 1745
rect 56180 1730 56195 1745
rect 56235 1730 56250 1745
rect 56290 1730 56305 1745
rect 56345 1730 56360 1745
rect 56400 1730 56415 1745
rect 56455 1730 56470 1745
rect 56510 1730 56525 1745
rect 56565 1730 56580 1745
rect 56620 1730 56635 1745
rect 56675 1730 56690 1745
rect 57110 1730 57125 1745
rect 57165 1730 57180 1745
rect 57220 1730 57235 1745
rect 57275 1730 57290 1745
rect 57330 1730 57345 1745
rect 57385 1730 57400 1745
rect 57440 1730 57455 1745
rect 57495 1730 57510 1745
rect 57550 1730 57565 1745
rect 57605 1730 57620 1745
rect 57660 1730 57675 1745
rect 57715 1730 57730 1745
rect 56035 1720 56085 1730
rect 56035 1700 56040 1720
rect 56060 1715 56085 1720
rect 56675 1720 56725 1730
rect 56675 1715 56700 1720
rect 56060 1700 56065 1715
rect 56035 1690 56065 1700
rect 56695 1700 56700 1715
rect 56720 1700 56725 1720
rect 56695 1690 56725 1700
rect 57075 1720 57125 1730
rect 57075 1700 57080 1720
rect 57100 1715 57125 1720
rect 57715 1720 57765 1730
rect 57715 1715 57740 1720
rect 57100 1700 57105 1715
rect 57075 1690 57105 1700
rect 57735 1700 57740 1715
rect 57760 1700 57765 1720
rect 57735 1690 57765 1700
rect 54660 1665 54675 1680
rect 54715 1670 54730 1680
rect 54770 1670 54785 1680
rect 54825 1670 54840 1680
rect 54880 1670 54895 1680
rect 54935 1670 54950 1680
rect 54990 1670 55005 1680
rect 55045 1670 55060 1680
rect 55100 1670 55115 1680
rect 55155 1670 55170 1680
rect 55210 1670 55225 1680
rect 54715 1655 55225 1670
rect 55265 1665 55280 1680
rect 58520 1665 58535 1680
rect 58575 1670 58590 1680
rect 58630 1670 58645 1680
rect 58685 1670 58700 1680
rect 58740 1670 58755 1680
rect 58795 1670 58810 1680
rect 58850 1670 58865 1680
rect 58905 1670 58920 1680
rect 58960 1670 58975 1680
rect 59015 1670 59030 1680
rect 59070 1670 59085 1680
rect 58575 1655 59085 1670
rect 59125 1665 59140 1680
rect 55120 1635 55125 1655
rect 55145 1635 55150 1655
rect 55120 1625 55150 1635
rect 58650 1635 58655 1655
rect 58675 1635 58680 1655
rect 58650 1625 58680 1635
rect 55125 1600 55145 1625
rect 58655 1600 58675 1625
rect 55115 1590 55155 1600
rect 55115 1570 55125 1590
rect 55145 1570 55155 1590
rect 55115 1550 55155 1570
rect 55115 1530 55125 1550
rect 55145 1530 55155 1550
rect 55115 1520 55155 1530
rect 58645 1590 58685 1600
rect 58645 1570 58655 1590
rect 58675 1570 58685 1590
rect 58645 1550 58685 1570
rect 58645 1530 58655 1550
rect 58675 1530 58685 1550
rect 58645 1520 58685 1530
rect 55125 1495 55145 1520
rect 58655 1495 58675 1520
rect 55120 1485 55150 1495
rect 55120 1465 55125 1485
rect 55145 1465 55150 1485
rect 58650 1485 58680 1495
rect 58650 1465 58655 1485
rect 58675 1465 58680 1485
rect 54660 1440 54675 1455
rect 54715 1450 55225 1465
rect 54715 1440 54730 1450
rect 54770 1440 54785 1450
rect 54825 1440 54840 1450
rect 54880 1440 54895 1450
rect 54935 1440 54950 1450
rect 54990 1440 55005 1450
rect 55045 1440 55060 1450
rect 55100 1440 55115 1450
rect 55155 1440 55170 1450
rect 55210 1440 55225 1450
rect 55265 1440 55280 1455
rect 58520 1440 58535 1455
rect 58575 1450 59085 1465
rect 58575 1440 58590 1450
rect 58630 1440 58645 1450
rect 58685 1440 58700 1450
rect 58740 1440 58755 1450
rect 58795 1440 58810 1450
rect 58850 1440 58865 1450
rect 58905 1440 58920 1450
rect 58960 1440 58975 1450
rect 59015 1440 59030 1450
rect 59070 1440 59085 1450
rect 59125 1440 59140 1455
rect 56690 1300 56720 1310
rect 56040 1290 56070 1300
rect 56040 1270 56045 1290
rect 56065 1275 56070 1290
rect 56690 1285 56695 1300
rect 56620 1280 56695 1285
rect 56715 1280 56720 1300
rect 56065 1270 56140 1275
rect 56040 1260 56140 1270
rect 56125 1245 56140 1260
rect 56620 1270 56720 1280
rect 56840 1300 56870 1310
rect 56840 1280 56845 1300
rect 56865 1285 56870 1300
rect 56930 1300 56960 1310
rect 56930 1285 56935 1300
rect 56865 1280 56880 1285
rect 56840 1270 56880 1280
rect 56620 1245 56635 1270
rect 56070 1220 56085 1235
rect 56125 1230 56635 1245
rect 56125 1220 56140 1230
rect 56180 1220 56195 1230
rect 56235 1220 56250 1230
rect 56290 1220 56305 1230
rect 56345 1220 56360 1230
rect 56400 1220 56415 1230
rect 56455 1220 56470 1230
rect 56510 1220 56525 1230
rect 56565 1220 56580 1230
rect 56620 1220 56635 1230
rect 56675 1220 56690 1235
rect 56810 1220 56825 1235
rect 56865 1220 56880 1270
rect 56920 1280 56935 1285
rect 56955 1280 56960 1300
rect 56920 1270 56960 1280
rect 57080 1300 57110 1310
rect 57080 1280 57085 1300
rect 57105 1285 57110 1300
rect 57730 1290 57760 1300
rect 57105 1280 57180 1285
rect 57080 1270 57180 1280
rect 57730 1275 57735 1290
rect 56920 1220 56935 1270
rect 57165 1245 57180 1270
rect 57660 1270 57735 1275
rect 57755 1270 57760 1290
rect 57660 1260 57760 1270
rect 57660 1245 57675 1260
rect 56975 1220 56990 1235
rect 57110 1220 57125 1235
rect 57165 1230 57675 1245
rect 57165 1220 57180 1230
rect 57220 1220 57235 1230
rect 57275 1220 57290 1230
rect 57330 1220 57345 1230
rect 57385 1220 57400 1230
rect 57440 1220 57455 1230
rect 57495 1220 57510 1230
rect 57550 1220 57565 1230
rect 57605 1220 57620 1230
rect 57660 1220 57675 1230
rect 57715 1220 57730 1235
rect 54660 1125 54675 1140
rect 54715 1125 54730 1140
rect 54770 1125 54785 1140
rect 54825 1125 54840 1140
rect 54880 1125 54895 1140
rect 54935 1125 54950 1140
rect 54990 1125 55005 1140
rect 55045 1125 55060 1140
rect 55100 1125 55115 1140
rect 55155 1125 55170 1140
rect 55210 1125 55225 1140
rect 55265 1125 55280 1140
rect 54625 1115 54675 1125
rect 54625 1095 54630 1115
rect 54650 1110 54675 1115
rect 55265 1115 55315 1125
rect 55265 1110 55290 1115
rect 54650 1095 54655 1110
rect 54625 1080 54655 1095
rect 55285 1095 55290 1110
rect 55310 1095 55315 1115
rect 55285 1080 55315 1095
rect 58520 1125 58535 1140
rect 58575 1125 58590 1140
rect 58630 1125 58645 1140
rect 58685 1125 58700 1140
rect 58740 1125 58755 1140
rect 58795 1125 58810 1140
rect 58850 1125 58865 1140
rect 58905 1125 58920 1140
rect 58960 1125 58975 1140
rect 59015 1125 59030 1140
rect 59070 1125 59085 1140
rect 59125 1125 59140 1140
rect 58485 1115 58535 1125
rect 58485 1095 58490 1115
rect 58510 1110 58535 1115
rect 59125 1115 59175 1125
rect 59125 1110 59150 1115
rect 58510 1095 58515 1110
rect 58485 1080 58515 1095
rect 59145 1095 59150 1110
rect 59170 1095 59175 1115
rect 59145 1085 59175 1095
rect 56070 1055 56085 1070
rect 56125 1055 56140 1070
rect 56180 1055 56195 1070
rect 56235 1055 56250 1070
rect 56290 1055 56305 1070
rect 56345 1055 56360 1070
rect 56400 1055 56415 1070
rect 56455 1055 56470 1070
rect 56510 1055 56525 1070
rect 56565 1055 56580 1070
rect 56620 1055 56635 1070
rect 56675 1055 56690 1070
rect 56810 1055 56825 1070
rect 56865 1055 56880 1070
rect 56920 1055 56935 1070
rect 56975 1055 56990 1070
rect 57110 1055 57125 1070
rect 57165 1055 57180 1070
rect 57220 1055 57235 1070
rect 57275 1055 57290 1070
rect 57330 1055 57345 1070
rect 57385 1055 57400 1070
rect 57440 1055 57455 1070
rect 57495 1055 57510 1070
rect 57550 1055 57565 1070
rect 57605 1055 57620 1070
rect 57660 1055 57675 1070
rect 57715 1055 57730 1070
rect 56035 1045 56085 1055
rect 56035 1025 56040 1045
rect 56060 1040 56085 1045
rect 56675 1045 56825 1055
rect 56675 1040 56740 1045
rect 56060 1025 56065 1040
rect 56035 1015 56065 1025
rect 56735 1025 56740 1040
rect 56760 1040 56825 1045
rect 56975 1045 57125 1055
rect 56975 1040 57040 1045
rect 56760 1025 56765 1040
rect 56735 1015 56765 1025
rect 57035 1025 57040 1040
rect 57060 1040 57125 1045
rect 57715 1045 57765 1055
rect 57715 1040 57740 1045
rect 57060 1025 57065 1040
rect 57035 1015 57065 1025
rect 57735 1025 57740 1040
rect 57760 1025 57765 1045
rect 57735 1015 57765 1025
rect 55000 520 55040 530
rect 55000 500 55010 520
rect 55030 500 55040 520
rect 55000 490 55040 500
rect 58760 520 58800 530
rect 58760 500 58770 520
rect 58790 500 58800 520
rect 58760 490 58800 500
rect 55010 365 55030 490
rect 56825 465 56865 475
rect 56825 445 56835 465
rect 56855 445 56865 465
rect 56935 465 56975 475
rect 56935 445 56945 465
rect 56965 445 56975 465
rect 56260 420 56275 435
rect 56315 430 57375 445
rect 56315 420 56330 430
rect 56370 420 56385 430
rect 56425 420 56440 430
rect 56480 420 56495 430
rect 56535 420 56550 430
rect 56590 420 56605 430
rect 56645 420 56660 430
rect 56700 420 56715 430
rect 56755 420 56770 430
rect 56810 420 56825 430
rect 56865 420 56880 430
rect 56920 420 56935 430
rect 56975 420 56990 430
rect 57030 420 57045 430
rect 57085 420 57100 430
rect 57140 420 57155 430
rect 57195 420 57210 430
rect 57250 420 57265 430
rect 57305 420 57320 430
rect 57360 420 57375 430
rect 57415 420 57430 435
rect 57470 420 57485 435
rect 54690 340 54750 355
rect 54790 350 55150 365
rect 54790 340 54850 350
rect 54890 340 54950 350
rect 54990 340 55050 350
rect 55090 340 55150 350
rect 55190 340 55250 355
rect 58770 365 58790 490
rect 58550 340 58610 355
rect 58650 350 59010 365
rect 58650 340 58710 350
rect 58750 340 58810 350
rect 58850 340 58910 350
rect 58950 340 59010 350
rect 59050 340 59110 355
rect 56260 155 56275 170
rect 56315 155 56330 170
rect 56370 155 56385 170
rect 56425 155 56440 170
rect 56480 155 56495 170
rect 56535 155 56550 170
rect 56590 155 56605 170
rect 56645 155 56660 170
rect 56700 155 56715 170
rect 56755 155 56770 170
rect 56810 155 56825 170
rect 56865 155 56880 170
rect 56920 155 56935 170
rect 56975 155 56990 170
rect 57030 155 57045 170
rect 57085 155 57100 170
rect 57140 155 57155 170
rect 57195 155 57210 170
rect 57250 155 57265 170
rect 57305 155 57320 170
rect 57360 155 57375 170
rect 56220 145 56275 155
rect 56220 125 56230 145
rect 56250 140 56275 145
rect 56250 125 56260 140
rect 56220 115 56260 125
rect 57415 45 57430 170
rect 57470 155 57485 170
rect 57470 145 57525 155
rect 57470 140 57495 145
rect 57485 125 57495 140
rect 57515 125 57525 145
rect 57485 115 57525 125
rect 57415 35 57455 45
rect 57415 15 57425 35
rect 57445 15 57455 35
rect 57415 5 57455 15
rect 56595 -255 56635 -245
rect 56595 -275 56605 -255
rect 56625 -275 56635 -255
rect 56920 -255 56960 -245
rect 56920 -275 56930 -255
rect 56950 -275 56960 -255
rect 56470 -300 56485 -285
rect 56525 -290 56705 -275
rect 56920 -285 56960 -275
rect 57040 -255 57080 -245
rect 57040 -275 57050 -255
rect 57070 -275 57080 -255
rect 57040 -285 57080 -275
rect 57160 -255 57200 -245
rect 57160 -275 57170 -255
rect 57190 -275 57200 -255
rect 57160 -285 57200 -275
rect 56525 -300 56540 -290
rect 56580 -300 56595 -290
rect 56635 -300 56650 -290
rect 56690 -300 56705 -290
rect 56745 -300 56760 -285
rect 56910 -300 57210 -285
rect 54690 -375 54750 -360
rect 54790 -375 54850 -360
rect 54890 -375 54950 -360
rect 54990 -375 55050 -360
rect 55090 -375 55150 -360
rect 55190 -375 55250 -360
rect 54655 -385 54750 -375
rect 54655 -405 54660 -385
rect 54680 -390 54750 -385
rect 55190 -385 55285 -375
rect 55190 -390 55260 -385
rect 54680 -405 54685 -390
rect 54655 -415 54685 -405
rect 55255 -405 55260 -390
rect 55280 -405 55285 -385
rect 55255 -415 55285 -405
rect 58550 -375 58610 -360
rect 58650 -375 58710 -360
rect 58750 -375 58810 -360
rect 58850 -375 58910 -360
rect 58950 -375 59010 -360
rect 59050 -375 59110 -360
rect 58515 -385 58610 -375
rect 58515 -405 58520 -385
rect 58540 -390 58610 -385
rect 59050 -385 59145 -375
rect 59050 -390 59120 -385
rect 58540 -405 58545 -390
rect 58515 -415 58545 -405
rect 59115 -405 59120 -390
rect 59140 -405 59145 -385
rect 59115 -415 59145 -405
rect 56470 -465 56485 -450
rect 56525 -465 56540 -450
rect 56580 -465 56595 -450
rect 56635 -465 56650 -450
rect 56690 -465 56705 -450
rect 56745 -465 56760 -450
rect 56910 -465 57210 -450
rect 56435 -475 56485 -465
rect 56435 -495 56440 -475
rect 56460 -480 56485 -475
rect 56745 -475 56795 -465
rect 56745 -480 56770 -475
rect 56460 -495 56465 -480
rect 56435 -505 56465 -495
rect 56765 -495 56770 -480
rect 56790 -495 56795 -475
rect 56765 -505 56795 -495
rect 56920 -475 56960 -465
rect 56920 -495 56930 -475
rect 56950 -495 56960 -475
rect 56920 -505 56960 -495
rect 57040 -475 57080 -465
rect 57040 -495 57050 -475
rect 57070 -495 57080 -475
rect 57040 -505 57080 -495
rect 57160 -475 57200 -465
rect 57160 -495 57170 -475
rect 57190 -495 57200 -475
rect 57160 -505 57200 -495
<< polycont >>
rect 56095 4905 56115 4925
rect 56275 4905 56295 4925
rect 57035 4905 57055 4925
rect 57215 4905 57235 4925
rect 57505 4905 57525 4925
rect 57685 4905 57705 4925
rect 56565 4735 56585 4755
rect 56745 4735 56765 4755
rect 56160 4455 56180 4475
rect 56635 4455 56655 4475
rect 57145 4455 57165 4475
rect 57581 4445 57601 4465
rect 54600 3620 54620 3640
rect 54960 3620 54980 3640
rect 55320 3620 55340 3640
rect 56015 3620 56035 3640
rect 56375 3620 56395 3640
rect 56735 3620 56755 3640
rect 57045 3620 57065 3640
rect 57405 3620 57425 3640
rect 57765 3620 57785 3640
rect 58460 3620 58480 3640
rect 58820 3620 58840 3640
rect 59180 3620 59200 3640
rect 56375 3555 56395 3575
rect 57405 3555 57425 3575
rect 54960 3510 54980 3530
rect 58820 3510 58840 3530
rect 56520 3250 56540 3270
rect 54630 3180 54650 3200
rect 55290 3180 55310 3200
rect 56850 3250 56870 3270
rect 56930 3250 56950 3270
rect 57260 3250 57280 3270
rect 58490 3180 58510 3200
rect 59150 3180 59170 3200
rect 56612 2875 56632 2895
rect 56685 2875 56705 2895
rect 56758 2875 56778 2895
rect 57022 2875 57042 2895
rect 57095 2875 57115 2895
rect 57168 2875 57188 2895
rect 56860 2590 56880 2610
rect 54960 2510 54980 2530
rect 54960 2445 54980 2465
rect 54960 2405 54980 2425
rect 54960 2365 54980 2385
rect 58820 2510 58840 2530
rect 58820 2445 58840 2465
rect 58820 2405 58840 2425
rect 58820 2365 58840 2385
rect 56780 2270 56800 2290
rect 57000 2270 57020 2290
rect 56045 1960 56065 1980
rect 54630 1905 54650 1925
rect 55290 1905 55310 1925
rect 56695 1960 56715 1980
rect 57085 1960 57105 1980
rect 57735 1960 57755 1980
rect 58490 1905 58510 1925
rect 59150 1905 59170 1925
rect 56040 1700 56060 1720
rect 56700 1700 56720 1720
rect 57080 1700 57100 1720
rect 57740 1700 57760 1720
rect 55125 1635 55145 1655
rect 58655 1635 58675 1655
rect 55125 1570 55145 1590
rect 55125 1530 55145 1550
rect 58655 1570 58675 1590
rect 58655 1530 58675 1550
rect 55125 1465 55145 1485
rect 58655 1465 58675 1485
rect 56045 1270 56065 1290
rect 56695 1280 56715 1300
rect 56845 1280 56865 1300
rect 56935 1280 56955 1300
rect 57085 1280 57105 1300
rect 57735 1270 57755 1290
rect 54630 1095 54650 1115
rect 55290 1095 55310 1115
rect 58490 1095 58510 1115
rect 59150 1095 59170 1115
rect 56040 1025 56060 1045
rect 56740 1025 56760 1045
rect 57040 1025 57060 1045
rect 57740 1025 57760 1045
rect 55010 500 55030 520
rect 58770 500 58790 520
rect 56835 445 56855 465
rect 56945 445 56965 465
rect 56230 125 56250 145
rect 57495 125 57515 145
rect 57425 15 57445 35
rect 56605 -275 56625 -255
rect 56930 -275 56950 -255
rect 57050 -275 57070 -255
rect 57170 -275 57190 -255
rect 54660 -405 54680 -385
rect 55260 -405 55280 -385
rect 58520 -405 58540 -385
rect 59120 -405 59140 -385
rect 56440 -495 56460 -475
rect 56770 -495 56790 -475
rect 56930 -495 56950 -475
rect 57050 -495 57070 -475
rect 57170 -495 57190 -475
<< xpolycontact >>
rect 54204 2940 54345 3160
rect 54204 2595 54345 2815
rect 59455 2940 59596 3160
rect 59455 2595 59596 2815
rect 54255 1544 54290 1764
rect 54255 1165 54290 1385
rect 54315 1544 54350 1764
rect 54315 1165 54350 1385
rect 54375 1544 54410 1764
rect 54375 1165 54410 1385
rect 54435 1544 54470 1764
rect 59330 1544 59365 1764
rect 54435 1165 54470 1385
rect 59330 1165 59365 1385
rect 59390 1544 59425 1764
rect 59390 1165 59425 1385
rect 59450 1544 59485 1764
rect 59450 1165 59485 1385
rect 59510 1544 59545 1764
rect 59510 1165 59545 1385
rect 54325 75 54360 295
rect 54325 -392 54360 -172
rect 54385 75 54420 295
rect 54385 -392 54420 -172
rect 59380 75 59415 295
rect 59380 -392 59415 -172
rect 59440 75 59475 295
rect 59440 -392 59475 -172
<< ppolyres >>
rect 54204 2815 54345 2940
rect 59455 2815 59596 2940
<< xpolyres >>
rect 54255 1385 54290 1544
rect 54315 1385 54350 1544
rect 54375 1385 54410 1544
rect 54435 1385 54470 1544
rect 59330 1385 59365 1544
rect 59390 1385 59425 1544
rect 59450 1385 59485 1544
rect 59510 1385 59545 1544
rect 54325 -172 54360 75
rect 54385 -172 54420 75
rect 59380 -172 59415 75
rect 59440 -172 59475 75
<< locali >>
rect 56085 4925 56125 4935
rect 56085 4905 56095 4925
rect 56115 4905 56125 4925
rect 56085 4895 56125 4905
rect 56265 4925 56305 4935
rect 56265 4905 56275 4925
rect 56295 4905 56305 4925
rect 56265 4895 56305 4905
rect 57025 4925 57065 4935
rect 57025 4905 57035 4925
rect 57055 4905 57065 4925
rect 57025 4895 57065 4905
rect 57205 4925 57245 4935
rect 57205 4905 57215 4925
rect 57235 4905 57245 4925
rect 57205 4895 57245 4905
rect 57495 4925 57535 4935
rect 57495 4905 57505 4925
rect 57525 4905 57535 4925
rect 57495 4895 57535 4905
rect 57675 4925 57715 4935
rect 57675 4905 57685 4925
rect 57705 4905 57715 4925
rect 57675 4895 57715 4905
rect 56050 4865 56120 4875
rect 56050 4545 56055 4865
rect 56075 4545 56095 4865
rect 56115 4545 56120 4865
rect 56050 4535 56120 4545
rect 56150 4865 56180 4875
rect 56150 4545 56155 4865
rect 56175 4545 56180 4865
rect 56150 4535 56180 4545
rect 56210 4865 56240 4875
rect 56210 4545 56215 4865
rect 56235 4545 56240 4865
rect 56210 4535 56240 4545
rect 56270 4865 56340 4875
rect 56270 4545 56275 4865
rect 56295 4545 56315 4865
rect 56335 4545 56340 4865
rect 56990 4865 57060 4875
rect 56555 4755 56595 4765
rect 56555 4735 56565 4755
rect 56585 4735 56595 4755
rect 56555 4725 56595 4735
rect 56735 4755 56775 4765
rect 56735 4735 56745 4755
rect 56765 4735 56775 4755
rect 56735 4725 56775 4735
rect 56270 4535 56340 4545
rect 56520 4695 56590 4705
rect 56520 4545 56525 4695
rect 56545 4545 56565 4695
rect 56585 4545 56590 4695
rect 56520 4535 56590 4545
rect 56620 4695 56650 4705
rect 56620 4545 56625 4695
rect 56645 4545 56650 4695
rect 56620 4535 56650 4545
rect 56680 4695 56710 4705
rect 56680 4545 56685 4695
rect 56705 4545 56710 4695
rect 56680 4535 56710 4545
rect 56740 4695 56810 4705
rect 56740 4545 56745 4695
rect 56765 4545 56785 4695
rect 56805 4545 56810 4695
rect 56740 4535 56810 4545
rect 56990 4545 56995 4865
rect 57015 4545 57035 4865
rect 57055 4545 57060 4865
rect 56990 4535 57060 4545
rect 57090 4865 57120 4875
rect 57090 4545 57095 4865
rect 57115 4545 57120 4865
rect 57090 4535 57120 4545
rect 57150 4865 57180 4875
rect 57150 4545 57155 4865
rect 57175 4545 57180 4865
rect 57150 4535 57180 4545
rect 57210 4865 57280 4875
rect 57210 4545 57215 4865
rect 57235 4545 57255 4865
rect 57275 4545 57280 4865
rect 57210 4535 57280 4545
rect 57460 4865 57530 4875
rect 57460 4545 57465 4865
rect 57485 4545 57505 4865
rect 57525 4545 57530 4865
rect 57460 4535 57530 4545
rect 57560 4865 57590 4875
rect 57560 4545 57565 4865
rect 57585 4545 57590 4865
rect 57560 4535 57590 4545
rect 57620 4865 57650 4875
rect 57620 4545 57625 4865
rect 57645 4545 57650 4865
rect 57620 4535 57650 4545
rect 57680 4865 57750 4875
rect 57680 4545 57685 4865
rect 57705 4545 57725 4865
rect 57745 4545 57750 4865
rect 57680 4535 57750 4545
rect 56150 4475 56190 4485
rect 56150 4455 56160 4475
rect 56180 4455 56190 4475
rect 56150 4445 56190 4455
rect 56630 4475 56660 4485
rect 56630 4455 56635 4475
rect 56655 4455 56660 4475
rect 56630 4445 56660 4455
rect 57140 4475 57170 4485
rect 57140 4455 57145 4475
rect 57165 4455 57170 4475
rect 57140 4445 57170 4455
rect 57576 4465 57606 4475
rect 57576 4445 57581 4465
rect 57601 4445 57606 4465
rect 57576 4435 57606 4445
rect 54555 4000 54625 4010
rect 54555 3680 54560 4000
rect 54580 3680 54600 4000
rect 54620 3680 54625 4000
rect 54555 3670 54625 3680
rect 54655 4000 54685 4010
rect 54655 3680 54660 4000
rect 54680 3680 54685 4000
rect 54655 3670 54685 3680
rect 54715 4000 54745 4010
rect 54715 3680 54720 4000
rect 54740 3680 54745 4000
rect 54715 3670 54745 3680
rect 54775 4000 54805 4010
rect 54775 3680 54780 4000
rect 54800 3680 54805 4000
rect 54775 3670 54805 3680
rect 54835 4000 54865 4010
rect 54835 3680 54840 4000
rect 54860 3680 54865 4000
rect 54835 3670 54865 3680
rect 54895 4000 54925 4010
rect 54895 3680 54900 4000
rect 54920 3680 54925 4000
rect 54895 3670 54925 3680
rect 54955 4000 54985 4010
rect 54955 3680 54960 4000
rect 54980 3680 54985 4000
rect 54955 3670 54985 3680
rect 55015 4000 55045 4010
rect 55015 3680 55020 4000
rect 55040 3680 55045 4000
rect 55015 3670 55045 3680
rect 55075 4000 55105 4010
rect 55075 3680 55080 4000
rect 55100 3680 55105 4000
rect 55075 3670 55105 3680
rect 55135 4000 55165 4010
rect 55135 3680 55140 4000
rect 55160 3680 55165 4000
rect 55135 3670 55165 3680
rect 55195 4000 55225 4010
rect 55195 3680 55200 4000
rect 55220 3680 55225 4000
rect 55195 3670 55225 3680
rect 55255 4000 55285 4010
rect 55255 3680 55260 4000
rect 55280 3680 55285 4000
rect 55255 3670 55285 3680
rect 55315 4000 55385 4010
rect 55315 3680 55320 4000
rect 55340 3680 55360 4000
rect 55380 3680 55385 4000
rect 55315 3670 55385 3680
rect 55970 4000 56040 4010
rect 55970 3680 55975 4000
rect 55995 3680 56015 4000
rect 56035 3680 56040 4000
rect 55970 3670 56040 3680
rect 56070 4000 56100 4010
rect 56070 3680 56075 4000
rect 56095 3680 56100 4000
rect 56070 3670 56100 3680
rect 56130 4000 56160 4010
rect 56130 3680 56135 4000
rect 56155 3680 56160 4000
rect 56130 3670 56160 3680
rect 56190 4000 56220 4010
rect 56190 3680 56195 4000
rect 56215 3680 56220 4000
rect 56190 3670 56220 3680
rect 56250 4000 56280 4010
rect 56250 3680 56255 4000
rect 56275 3680 56280 4000
rect 56250 3670 56280 3680
rect 56310 4000 56340 4010
rect 56310 3680 56315 4000
rect 56335 3680 56340 4000
rect 56310 3670 56340 3680
rect 56370 4000 56400 4010
rect 56370 3680 56375 4000
rect 56395 3680 56400 4000
rect 56370 3670 56400 3680
rect 56430 4000 56460 4010
rect 56430 3680 56435 4000
rect 56455 3680 56460 4000
rect 56430 3670 56460 3680
rect 56490 4000 56520 4010
rect 56490 3680 56495 4000
rect 56515 3680 56520 4000
rect 56490 3670 56520 3680
rect 56550 4000 56580 4010
rect 56550 3680 56555 4000
rect 56575 3680 56580 4000
rect 56550 3670 56580 3680
rect 56610 4000 56640 4010
rect 56610 3680 56615 4000
rect 56635 3680 56640 4000
rect 56610 3670 56640 3680
rect 56670 4000 56700 4010
rect 56670 3680 56675 4000
rect 56695 3680 56700 4000
rect 56670 3670 56700 3680
rect 56730 4000 56800 4010
rect 56730 3680 56735 4000
rect 56755 3680 56775 4000
rect 56795 3680 56800 4000
rect 56730 3670 56800 3680
rect 57000 4000 57070 4010
rect 57000 3680 57005 4000
rect 57025 3680 57045 4000
rect 57065 3680 57070 4000
rect 57000 3670 57070 3680
rect 57100 4000 57130 4010
rect 57100 3680 57105 4000
rect 57125 3680 57130 4000
rect 57100 3670 57130 3680
rect 57160 4000 57190 4010
rect 57160 3680 57165 4000
rect 57185 3680 57190 4000
rect 57160 3670 57190 3680
rect 57220 4000 57250 4010
rect 57220 3680 57225 4000
rect 57245 3680 57250 4000
rect 57220 3670 57250 3680
rect 57280 4000 57310 4010
rect 57280 3680 57285 4000
rect 57305 3680 57310 4000
rect 57280 3670 57310 3680
rect 57340 4000 57370 4010
rect 57340 3680 57345 4000
rect 57365 3680 57370 4000
rect 57340 3670 57370 3680
rect 57400 4000 57430 4010
rect 57400 3680 57405 4000
rect 57425 3680 57430 4000
rect 57400 3670 57430 3680
rect 57460 4000 57490 4010
rect 57460 3680 57465 4000
rect 57485 3680 57490 4000
rect 57460 3670 57490 3680
rect 57520 4000 57550 4010
rect 57520 3680 57525 4000
rect 57545 3680 57550 4000
rect 57520 3670 57550 3680
rect 57580 4000 57610 4010
rect 57580 3680 57585 4000
rect 57605 3680 57610 4000
rect 57580 3670 57610 3680
rect 57640 4000 57670 4010
rect 57640 3680 57645 4000
rect 57665 3680 57670 4000
rect 57640 3670 57670 3680
rect 57700 4000 57730 4010
rect 57700 3680 57705 4000
rect 57725 3680 57730 4000
rect 57700 3670 57730 3680
rect 57760 4000 57830 4010
rect 57760 3680 57765 4000
rect 57785 3680 57805 4000
rect 57825 3680 57830 4000
rect 57760 3670 57830 3680
rect 58415 4000 58485 4010
rect 58415 3680 58420 4000
rect 58440 3680 58460 4000
rect 58480 3680 58485 4000
rect 58415 3670 58485 3680
rect 58515 4000 58545 4010
rect 58515 3680 58520 4000
rect 58540 3680 58545 4000
rect 58515 3670 58545 3680
rect 58575 4000 58605 4010
rect 58575 3680 58580 4000
rect 58600 3680 58605 4000
rect 58575 3670 58605 3680
rect 58635 4000 58665 4010
rect 58635 3680 58640 4000
rect 58660 3680 58665 4000
rect 58635 3670 58665 3680
rect 58695 4000 58725 4010
rect 58695 3680 58700 4000
rect 58720 3680 58725 4000
rect 58695 3670 58725 3680
rect 58755 4000 58785 4010
rect 58755 3680 58760 4000
rect 58780 3680 58785 4000
rect 58755 3670 58785 3680
rect 58815 4000 58845 4010
rect 58815 3680 58820 4000
rect 58840 3680 58845 4000
rect 58815 3670 58845 3680
rect 58875 4000 58905 4010
rect 58875 3680 58880 4000
rect 58900 3680 58905 4000
rect 58875 3670 58905 3680
rect 58935 4000 58965 4010
rect 58935 3680 58940 4000
rect 58960 3680 58965 4000
rect 58935 3670 58965 3680
rect 58995 4000 59025 4010
rect 58995 3680 59000 4000
rect 59020 3680 59025 4000
rect 58995 3670 59025 3680
rect 59055 4000 59085 4010
rect 59055 3680 59060 4000
rect 59080 3680 59085 4000
rect 59055 3670 59085 3680
rect 59115 4000 59145 4010
rect 59115 3680 59120 4000
rect 59140 3680 59145 4000
rect 59115 3670 59145 3680
rect 59175 4000 59245 4010
rect 59175 3680 59180 4000
rect 59200 3680 59220 4000
rect 59240 3680 59245 4000
rect 59175 3670 59245 3680
rect 54595 3640 54625 3650
rect 54595 3620 54600 3640
rect 54620 3620 54625 3640
rect 54595 3610 54625 3620
rect 54955 3640 54985 3650
rect 54955 3620 54960 3640
rect 54980 3620 54985 3640
rect 54955 3610 54985 3620
rect 55315 3640 55345 3650
rect 55315 3620 55320 3640
rect 55340 3620 55345 3640
rect 55315 3610 55345 3620
rect 56010 3640 56040 3650
rect 56010 3620 56015 3640
rect 56035 3620 56040 3640
rect 56010 3610 56040 3620
rect 56370 3640 56400 3650
rect 56370 3620 56375 3640
rect 56395 3620 56400 3640
rect 56370 3610 56400 3620
rect 56730 3640 56760 3650
rect 56730 3620 56735 3640
rect 56755 3620 56760 3640
rect 56730 3610 56760 3620
rect 57040 3640 57070 3650
rect 57040 3620 57045 3640
rect 57065 3620 57070 3640
rect 57040 3610 57070 3620
rect 57400 3640 57430 3650
rect 57400 3620 57405 3640
rect 57425 3620 57430 3640
rect 57400 3610 57430 3620
rect 57760 3640 57790 3650
rect 57760 3620 57765 3640
rect 57785 3620 57790 3640
rect 57760 3610 57790 3620
rect 58455 3640 58485 3650
rect 58455 3620 58460 3640
rect 58480 3620 58485 3640
rect 58455 3610 58485 3620
rect 58815 3640 58845 3650
rect 58815 3620 58820 3640
rect 58840 3620 58845 3640
rect 58815 3610 58845 3620
rect 59175 3640 59205 3650
rect 59175 3620 59180 3640
rect 59200 3620 59205 3640
rect 59175 3610 59205 3620
rect 56365 3575 56405 3585
rect 56365 3555 56375 3575
rect 56395 3555 56405 3575
rect 56365 3545 56405 3555
rect 57395 3575 57435 3585
rect 57395 3555 57405 3575
rect 57425 3555 57435 3575
rect 57395 3545 57435 3555
rect 54950 3530 54990 3540
rect 54950 3510 54960 3530
rect 54980 3510 54990 3530
rect 54950 3500 54990 3510
rect 58810 3530 58850 3540
rect 58810 3510 58820 3530
rect 58840 3510 58850 3530
rect 58810 3500 58850 3510
rect 56510 3270 56550 3280
rect 56510 3250 56520 3270
rect 56540 3250 56550 3270
rect 56510 3240 56550 3250
rect 56680 3270 56710 3280
rect 56680 3250 56685 3270
rect 56705 3250 56710 3270
rect 56680 3240 56710 3250
rect 56840 3270 56880 3280
rect 56840 3250 56850 3270
rect 56870 3250 56880 3270
rect 56840 3240 56880 3250
rect 56920 3270 56960 3280
rect 56920 3250 56930 3270
rect 56950 3250 56960 3270
rect 56920 3240 56960 3250
rect 57090 3270 57120 3280
rect 57090 3250 57095 3270
rect 57115 3250 57120 3270
rect 57090 3240 57120 3250
rect 57250 3270 57290 3280
rect 57250 3250 57260 3270
rect 57280 3250 57290 3270
rect 57250 3240 57290 3250
rect 54625 3200 54655 3210
rect 54204 3190 54345 3200
rect 54204 3170 54210 3190
rect 54230 3170 54265 3190
rect 54285 3170 54320 3190
rect 54340 3170 54345 3190
rect 54625 3180 54630 3200
rect 54650 3180 54655 3200
rect 54625 3170 54655 3180
rect 55285 3200 55315 3210
rect 55285 3180 55290 3200
rect 55310 3180 55315 3200
rect 55285 3170 55315 3180
rect 54204 3160 54345 3170
rect 56520 3165 56540 3240
rect 56620 3215 56660 3225
rect 56620 3195 56630 3215
rect 56650 3195 56660 3215
rect 56620 3185 56660 3195
rect 56630 3165 56650 3185
rect 56685 3165 56705 3240
rect 56730 3215 56770 3225
rect 56730 3195 56740 3215
rect 56760 3195 56770 3215
rect 56730 3185 56770 3195
rect 56740 3165 56760 3185
rect 56850 3165 56870 3240
rect 56930 3165 56950 3240
rect 57030 3215 57070 3225
rect 57030 3195 57040 3215
rect 57060 3195 57070 3215
rect 57030 3185 57070 3195
rect 57040 3165 57060 3185
rect 57095 3165 57115 3240
rect 57140 3215 57180 3225
rect 57140 3195 57150 3215
rect 57170 3195 57180 3215
rect 57140 3185 57180 3195
rect 57150 3165 57170 3185
rect 57260 3165 57280 3240
rect 58485 3200 58515 3210
rect 58485 3180 58490 3200
rect 58510 3180 58515 3200
rect 58485 3170 58515 3180
rect 59145 3200 59175 3210
rect 59145 3180 59150 3200
rect 59170 3180 59175 3200
rect 59145 3170 59175 3180
rect 59455 3190 59596 3200
rect 59455 3170 59460 3190
rect 59480 3170 59515 3190
rect 59535 3170 59570 3190
rect 59590 3170 59596 3190
rect 56475 3155 56545 3165
rect 54585 3140 54655 3150
rect 54204 2585 54345 2595
rect 54204 2565 54210 2585
rect 54230 2565 54265 2585
rect 54285 2565 54320 2585
rect 54340 2565 54345 2585
rect 54204 2555 54345 2565
rect 54585 2570 54590 3140
rect 54610 2570 54630 3140
rect 54650 2570 54655 3140
rect 54585 2560 54655 2570
rect 54680 3140 54710 3150
rect 54680 2570 54685 3140
rect 54705 2570 54710 3140
rect 54680 2560 54710 2570
rect 54735 3140 54765 3150
rect 54735 2570 54740 3140
rect 54760 2570 54765 3140
rect 54735 2560 54765 2570
rect 54790 3140 54820 3150
rect 54790 2570 54795 3140
rect 54815 2570 54820 3140
rect 54790 2560 54820 2570
rect 54845 3140 54875 3150
rect 54845 2570 54850 3140
rect 54870 2570 54875 3140
rect 54845 2560 54875 2570
rect 54900 3140 54930 3150
rect 54900 2570 54905 3140
rect 54925 2570 54930 3140
rect 54900 2560 54930 2570
rect 54955 3140 54985 3150
rect 54955 2570 54960 3140
rect 54980 2570 54985 3140
rect 54955 2560 54985 2570
rect 55010 3140 55040 3150
rect 55010 2570 55015 3140
rect 55035 2570 55040 3140
rect 55010 2560 55040 2570
rect 55065 3140 55095 3150
rect 55065 2570 55070 3140
rect 55090 2570 55095 3140
rect 55065 2560 55095 2570
rect 55120 3140 55150 3150
rect 55120 2570 55125 3140
rect 55145 2570 55150 3140
rect 55120 2560 55150 2570
rect 55175 3140 55205 3150
rect 55175 2570 55180 3140
rect 55200 2570 55205 3140
rect 55175 2560 55205 2570
rect 55230 3140 55260 3150
rect 55230 2570 55235 3140
rect 55255 2570 55260 3140
rect 55230 2560 55260 2570
rect 55285 3140 55355 3150
rect 55285 2570 55290 3140
rect 55310 2570 55330 3140
rect 55350 2570 55355 3140
rect 56475 3135 56480 3155
rect 56500 3135 56520 3155
rect 56540 3135 56545 3155
rect 56475 3105 56545 3135
rect 56475 3085 56480 3105
rect 56500 3085 56520 3105
rect 56540 3085 56545 3105
rect 56475 3055 56545 3085
rect 56475 3035 56480 3055
rect 56500 3035 56520 3055
rect 56540 3035 56545 3055
rect 56475 3005 56545 3035
rect 56475 2985 56480 3005
rect 56500 2985 56520 3005
rect 56540 2985 56545 3005
rect 56475 2955 56545 2985
rect 56475 2935 56480 2955
rect 56500 2935 56520 2955
rect 56540 2935 56545 2955
rect 56475 2925 56545 2935
rect 56570 3155 56600 3165
rect 56570 3135 56575 3155
rect 56595 3135 56600 3155
rect 56570 3105 56600 3135
rect 56570 3085 56575 3105
rect 56595 3085 56600 3105
rect 56570 3055 56600 3085
rect 56570 3035 56575 3055
rect 56595 3035 56600 3055
rect 56570 3005 56600 3035
rect 56570 2985 56575 3005
rect 56595 2985 56600 3005
rect 56570 2955 56600 2985
rect 56570 2935 56575 2955
rect 56595 2935 56600 2955
rect 56570 2925 56600 2935
rect 56625 3155 56655 3165
rect 56625 3135 56630 3155
rect 56650 3135 56655 3155
rect 56625 3105 56655 3135
rect 56625 3085 56630 3105
rect 56650 3085 56655 3105
rect 56625 3055 56655 3085
rect 56625 3035 56630 3055
rect 56650 3035 56655 3055
rect 56625 3005 56655 3035
rect 56625 2985 56630 3005
rect 56650 2985 56655 3005
rect 56625 2955 56655 2985
rect 56625 2935 56630 2955
rect 56650 2935 56655 2955
rect 56625 2925 56655 2935
rect 56680 3155 56710 3165
rect 56680 3135 56685 3155
rect 56705 3135 56710 3155
rect 56680 3105 56710 3135
rect 56680 3085 56685 3105
rect 56705 3085 56710 3105
rect 56680 3055 56710 3085
rect 56680 3035 56685 3055
rect 56705 3035 56710 3055
rect 56680 3005 56710 3035
rect 56680 2985 56685 3005
rect 56705 2985 56710 3005
rect 56680 2955 56710 2985
rect 56680 2935 56685 2955
rect 56705 2935 56710 2955
rect 56680 2925 56710 2935
rect 56735 3155 56765 3165
rect 56735 3135 56740 3155
rect 56760 3135 56765 3155
rect 56735 3105 56765 3135
rect 56735 3085 56740 3105
rect 56760 3085 56765 3105
rect 56735 3055 56765 3085
rect 56735 3035 56740 3055
rect 56760 3035 56765 3055
rect 56735 3005 56765 3035
rect 56735 2985 56740 3005
rect 56760 2985 56765 3005
rect 56735 2955 56765 2985
rect 56735 2935 56740 2955
rect 56760 2935 56765 2955
rect 56735 2925 56765 2935
rect 56790 3155 56820 3165
rect 56790 3135 56795 3155
rect 56815 3135 56820 3155
rect 56790 3105 56820 3135
rect 56790 3085 56795 3105
rect 56815 3085 56820 3105
rect 56790 3055 56820 3085
rect 56790 3035 56795 3055
rect 56815 3035 56820 3055
rect 56790 3005 56820 3035
rect 56790 2985 56795 3005
rect 56815 2985 56820 3005
rect 56790 2955 56820 2985
rect 56790 2935 56795 2955
rect 56815 2935 56820 2955
rect 56790 2925 56820 2935
rect 56845 3155 56955 3165
rect 56845 3135 56850 3155
rect 56870 3135 56890 3155
rect 56910 3135 56930 3155
rect 56950 3135 56955 3155
rect 56845 3105 56955 3135
rect 56845 3085 56850 3105
rect 56870 3085 56890 3105
rect 56910 3085 56930 3105
rect 56950 3085 56955 3105
rect 56845 3055 56955 3085
rect 56845 3035 56850 3055
rect 56870 3035 56890 3055
rect 56910 3035 56930 3055
rect 56950 3035 56955 3055
rect 56845 3005 56955 3035
rect 56845 2985 56850 3005
rect 56870 2985 56890 3005
rect 56910 2985 56930 3005
rect 56950 2985 56955 3005
rect 56845 2955 56955 2985
rect 56845 2935 56850 2955
rect 56870 2935 56890 2955
rect 56910 2935 56930 2955
rect 56950 2935 56955 2955
rect 56845 2925 56955 2935
rect 56980 3155 57010 3165
rect 56980 3135 56985 3155
rect 57005 3135 57010 3155
rect 56980 3105 57010 3135
rect 56980 3085 56985 3105
rect 57005 3085 57010 3105
rect 56980 3055 57010 3085
rect 56980 3035 56985 3055
rect 57005 3035 57010 3055
rect 56980 3005 57010 3035
rect 56980 2985 56985 3005
rect 57005 2985 57010 3005
rect 56980 2955 57010 2985
rect 56980 2935 56985 2955
rect 57005 2935 57010 2955
rect 56980 2925 57010 2935
rect 57035 3155 57065 3165
rect 57035 3135 57040 3155
rect 57060 3135 57065 3155
rect 57035 3105 57065 3135
rect 57035 3085 57040 3105
rect 57060 3085 57065 3105
rect 57035 3055 57065 3085
rect 57035 3035 57040 3055
rect 57060 3035 57065 3055
rect 57035 3005 57065 3035
rect 57035 2985 57040 3005
rect 57060 2985 57065 3005
rect 57035 2955 57065 2985
rect 57035 2935 57040 2955
rect 57060 2935 57065 2955
rect 57035 2925 57065 2935
rect 57090 3155 57120 3165
rect 57090 3135 57095 3155
rect 57115 3135 57120 3155
rect 57090 3105 57120 3135
rect 57090 3085 57095 3105
rect 57115 3085 57120 3105
rect 57090 3055 57120 3085
rect 57090 3035 57095 3055
rect 57115 3035 57120 3055
rect 57090 3005 57120 3035
rect 57090 2985 57095 3005
rect 57115 2985 57120 3005
rect 57090 2955 57120 2985
rect 57090 2935 57095 2955
rect 57115 2935 57120 2955
rect 57090 2925 57120 2935
rect 57145 3155 57175 3165
rect 57145 3135 57150 3155
rect 57170 3135 57175 3155
rect 57145 3105 57175 3135
rect 57145 3085 57150 3105
rect 57170 3085 57175 3105
rect 57145 3055 57175 3085
rect 57145 3035 57150 3055
rect 57170 3035 57175 3055
rect 57145 3005 57175 3035
rect 57145 2985 57150 3005
rect 57170 2985 57175 3005
rect 57145 2955 57175 2985
rect 57145 2935 57150 2955
rect 57170 2935 57175 2955
rect 57145 2925 57175 2935
rect 57200 3155 57230 3165
rect 57200 3135 57205 3155
rect 57225 3135 57230 3155
rect 57200 3105 57230 3135
rect 57200 3085 57205 3105
rect 57225 3085 57230 3105
rect 57200 3055 57230 3085
rect 57200 3035 57205 3055
rect 57225 3035 57230 3055
rect 57200 3005 57230 3035
rect 57200 2985 57205 3005
rect 57225 2985 57230 3005
rect 57200 2955 57230 2985
rect 57200 2935 57205 2955
rect 57225 2935 57230 2955
rect 57200 2925 57230 2935
rect 57255 3155 57325 3165
rect 57255 3135 57260 3155
rect 57280 3135 57300 3155
rect 57320 3135 57325 3155
rect 59455 3160 59596 3170
rect 57255 3105 57325 3135
rect 57255 3085 57260 3105
rect 57280 3085 57300 3105
rect 57320 3085 57325 3105
rect 57255 3055 57325 3085
rect 57255 3035 57260 3055
rect 57280 3035 57300 3055
rect 57320 3035 57325 3055
rect 57255 3005 57325 3035
rect 57255 2985 57260 3005
rect 57280 2985 57300 3005
rect 57320 2985 57325 3005
rect 57255 2955 57325 2985
rect 57255 2935 57260 2955
rect 57280 2935 57300 2955
rect 57320 2935 57325 2955
rect 57255 2925 57325 2935
rect 58445 3140 58515 3150
rect 56570 2915 56590 2925
rect 56560 2905 56590 2915
rect 56800 2915 56820 2925
rect 56980 2915 57000 2925
rect 56800 2905 56830 2915
rect 56560 2885 56565 2905
rect 56585 2885 56590 2905
rect 56560 2875 56590 2885
rect 56607 2895 56637 2905
rect 56607 2875 56612 2895
rect 56632 2875 56637 2895
rect 56607 2865 56637 2875
rect 56675 2895 56715 2905
rect 56675 2875 56685 2895
rect 56705 2875 56715 2895
rect 56675 2865 56715 2875
rect 56753 2895 56783 2905
rect 56753 2875 56758 2895
rect 56778 2875 56783 2895
rect 56800 2885 56805 2905
rect 56825 2885 56830 2905
rect 56800 2875 56830 2885
rect 56970 2905 57000 2915
rect 57210 2915 57230 2925
rect 57210 2905 57240 2915
rect 56970 2885 56975 2905
rect 56995 2885 57000 2905
rect 56970 2875 57000 2885
rect 57017 2895 57047 2905
rect 57017 2875 57022 2895
rect 57042 2875 57047 2895
rect 56753 2865 56783 2875
rect 57017 2865 57047 2875
rect 57085 2895 57125 2905
rect 57085 2875 57095 2895
rect 57115 2875 57125 2895
rect 57085 2865 57125 2875
rect 57163 2895 57193 2905
rect 57163 2875 57168 2895
rect 57188 2875 57193 2895
rect 57210 2885 57215 2905
rect 57235 2885 57240 2905
rect 57210 2875 57240 2885
rect 57163 2865 57193 2875
rect 56600 2825 56640 2835
rect 56600 2805 56610 2825
rect 56630 2805 56640 2825
rect 56600 2795 56640 2805
rect 57160 2825 57200 2835
rect 57160 2805 57170 2825
rect 57190 2805 57200 2825
rect 57160 2795 57200 2805
rect 56850 2610 56890 2620
rect 56850 2590 56860 2610
rect 56880 2590 56890 2610
rect 56850 2580 56890 2590
rect 56935 2610 56975 2620
rect 56935 2590 56945 2610
rect 56965 2590 56975 2610
rect 56935 2580 56975 2590
rect 55285 2560 55355 2570
rect 58445 2570 58450 3140
rect 58470 2570 58490 3140
rect 58510 2570 58515 3140
rect 58445 2560 58515 2570
rect 58540 3140 58570 3150
rect 58540 2570 58545 3140
rect 58565 2570 58570 3140
rect 58540 2560 58570 2570
rect 58595 3140 58625 3150
rect 58595 2570 58600 3140
rect 58620 2570 58625 3140
rect 58595 2560 58625 2570
rect 58650 3140 58680 3150
rect 58650 2570 58655 3140
rect 58675 2570 58680 3140
rect 58650 2560 58680 2570
rect 58705 3140 58735 3150
rect 58705 2570 58710 3140
rect 58730 2570 58735 3140
rect 58705 2560 58735 2570
rect 58760 3140 58790 3150
rect 58760 2570 58765 3140
rect 58785 2570 58790 3140
rect 58760 2560 58790 2570
rect 58815 3140 58845 3150
rect 58815 2570 58820 3140
rect 58840 2570 58845 3140
rect 58815 2560 58845 2570
rect 58870 3140 58900 3150
rect 58870 2570 58875 3140
rect 58895 2570 58900 3140
rect 58870 2560 58900 2570
rect 58925 3140 58955 3150
rect 58925 2570 58930 3140
rect 58950 2570 58955 3140
rect 58925 2560 58955 2570
rect 58980 3140 59010 3150
rect 58980 2570 58985 3140
rect 59005 2570 59010 3140
rect 58980 2560 59010 2570
rect 59035 3140 59065 3150
rect 59035 2570 59040 3140
rect 59060 2570 59065 3140
rect 59035 2560 59065 2570
rect 59090 3140 59120 3150
rect 59090 2570 59095 3140
rect 59115 2570 59120 3140
rect 59090 2560 59120 2570
rect 59145 3140 59215 3150
rect 59145 2570 59150 3140
rect 59170 2570 59190 3140
rect 59210 2570 59215 3140
rect 59145 2560 59215 2570
rect 59455 2585 59596 2595
rect 59455 2565 59460 2585
rect 59480 2565 59515 2585
rect 59535 2565 59570 2585
rect 59590 2565 59596 2585
rect 56735 2550 56805 2560
rect 54955 2530 54985 2540
rect 54955 2510 54960 2530
rect 54980 2510 54985 2530
rect 54955 2500 54985 2510
rect 54950 2465 54990 2475
rect 54950 2445 54960 2465
rect 54980 2445 54990 2465
rect 54950 2425 54990 2445
rect 54950 2405 54960 2425
rect 54980 2405 54990 2425
rect 54950 2385 54990 2405
rect 54950 2365 54960 2385
rect 54980 2365 54990 2385
rect 54950 2355 54990 2365
rect 56735 2330 56740 2550
rect 56760 2330 56780 2550
rect 56800 2330 56805 2550
rect 56735 2320 56805 2330
rect 56830 2550 56860 2560
rect 56830 2330 56835 2550
rect 56855 2330 56860 2550
rect 56830 2320 56860 2330
rect 56885 2550 56915 2560
rect 56885 2330 56890 2550
rect 56910 2330 56915 2550
rect 56885 2320 56915 2330
rect 56940 2550 56970 2560
rect 56940 2330 56945 2550
rect 56965 2330 56970 2550
rect 56940 2320 56970 2330
rect 56995 2550 57065 2560
rect 59455 2555 59596 2565
rect 56995 2330 57000 2550
rect 57020 2330 57040 2550
rect 57060 2330 57065 2550
rect 58815 2530 58845 2540
rect 58815 2510 58820 2530
rect 58840 2510 58845 2530
rect 58815 2500 58845 2510
rect 58810 2465 58850 2475
rect 58810 2445 58820 2465
rect 58840 2445 58850 2465
rect 58810 2425 58850 2445
rect 58810 2405 58820 2425
rect 58840 2405 58850 2425
rect 58810 2385 58850 2405
rect 58810 2365 58820 2385
rect 58840 2365 58850 2385
rect 58810 2355 58850 2365
rect 56995 2320 57065 2330
rect 56770 2290 56810 2300
rect 56770 2270 56780 2290
rect 56800 2270 56810 2290
rect 56770 2260 56810 2270
rect 56990 2290 57030 2300
rect 56990 2270 57000 2290
rect 57020 2270 57030 2290
rect 56990 2260 57030 2270
rect 56040 1980 56070 1990
rect 56040 1960 56045 1980
rect 56065 1960 56070 1980
rect 56040 1950 56070 1960
rect 56690 1980 56720 1990
rect 56690 1960 56695 1980
rect 56715 1960 56720 1980
rect 56690 1950 56720 1960
rect 57080 1980 57110 1990
rect 57080 1960 57085 1980
rect 57105 1960 57110 1980
rect 57080 1950 57110 1960
rect 57730 1980 57760 1990
rect 57730 1960 57735 1980
rect 57755 1960 57760 1980
rect 57730 1950 57760 1960
rect 54625 1925 54655 1935
rect 54625 1905 54630 1925
rect 54650 1905 54655 1925
rect 54625 1895 54655 1905
rect 55285 1925 55315 1935
rect 55285 1905 55290 1925
rect 55310 1905 55315 1925
rect 55285 1895 55315 1905
rect 58485 1925 58515 1935
rect 58485 1905 58490 1925
rect 58510 1905 58515 1925
rect 58485 1895 58515 1905
rect 59145 1925 59175 1935
rect 59145 1905 59150 1925
rect 59170 1905 59175 1925
rect 59145 1895 59175 1905
rect 55995 1880 56065 1890
rect 54585 1865 54655 1875
rect 54255 1781 54470 1801
rect 54255 1764 54290 1781
rect 54435 1764 54470 1781
rect 54350 1714 54375 1764
rect 54585 1695 54590 1865
rect 54610 1695 54630 1865
rect 54650 1695 54655 1865
rect 54585 1685 54655 1695
rect 54680 1865 54710 1875
rect 54680 1695 54685 1865
rect 54705 1695 54710 1865
rect 54680 1685 54710 1695
rect 54735 1865 54765 1875
rect 54735 1695 54740 1865
rect 54760 1695 54765 1865
rect 54735 1685 54765 1695
rect 54790 1865 54820 1875
rect 54790 1695 54795 1865
rect 54815 1695 54820 1865
rect 54790 1685 54820 1695
rect 54845 1865 54875 1875
rect 54845 1695 54850 1865
rect 54870 1695 54875 1865
rect 54845 1685 54875 1695
rect 54900 1865 54930 1875
rect 54900 1695 54905 1865
rect 54925 1695 54930 1865
rect 54900 1685 54930 1695
rect 54955 1865 54985 1875
rect 54955 1695 54960 1865
rect 54980 1695 54985 1865
rect 54955 1685 54985 1695
rect 55010 1865 55040 1875
rect 55010 1695 55015 1865
rect 55035 1695 55040 1865
rect 55010 1685 55040 1695
rect 55065 1865 55095 1875
rect 55065 1695 55070 1865
rect 55090 1695 55095 1865
rect 55065 1685 55095 1695
rect 55120 1865 55150 1875
rect 55120 1695 55125 1865
rect 55145 1695 55150 1865
rect 55120 1685 55150 1695
rect 55175 1865 55205 1875
rect 55175 1695 55180 1865
rect 55200 1695 55205 1865
rect 55175 1685 55205 1695
rect 55230 1865 55260 1875
rect 55230 1695 55235 1865
rect 55255 1695 55260 1865
rect 55230 1685 55260 1695
rect 55285 1865 55355 1875
rect 55285 1695 55290 1865
rect 55310 1695 55330 1865
rect 55350 1695 55355 1865
rect 55995 1760 56000 1880
rect 56020 1760 56040 1880
rect 56060 1760 56065 1880
rect 55995 1750 56065 1760
rect 56090 1880 56120 1890
rect 56090 1760 56095 1880
rect 56115 1760 56120 1880
rect 56090 1750 56120 1760
rect 56145 1880 56175 1890
rect 56145 1760 56150 1880
rect 56170 1760 56175 1880
rect 56145 1750 56175 1760
rect 56200 1880 56230 1890
rect 56200 1760 56205 1880
rect 56225 1760 56230 1880
rect 56200 1750 56230 1760
rect 56255 1880 56285 1890
rect 56255 1760 56260 1880
rect 56280 1760 56285 1880
rect 56255 1750 56285 1760
rect 56310 1880 56340 1890
rect 56310 1760 56315 1880
rect 56335 1760 56340 1880
rect 56310 1750 56340 1760
rect 56365 1880 56395 1890
rect 56365 1760 56370 1880
rect 56390 1760 56395 1880
rect 56365 1750 56395 1760
rect 56420 1880 56450 1890
rect 56420 1760 56425 1880
rect 56445 1760 56450 1880
rect 56420 1750 56450 1760
rect 56475 1880 56505 1890
rect 56475 1760 56480 1880
rect 56500 1760 56505 1880
rect 56475 1750 56505 1760
rect 56530 1880 56560 1890
rect 56530 1760 56535 1880
rect 56555 1760 56560 1880
rect 56530 1750 56560 1760
rect 56585 1880 56615 1890
rect 56585 1760 56590 1880
rect 56610 1760 56615 1880
rect 56585 1750 56615 1760
rect 56640 1880 56670 1890
rect 56640 1760 56645 1880
rect 56665 1760 56670 1880
rect 56640 1750 56670 1760
rect 56695 1880 56765 1890
rect 56695 1760 56700 1880
rect 56720 1760 56740 1880
rect 56760 1760 56765 1880
rect 56695 1750 56765 1760
rect 57035 1880 57105 1890
rect 57035 1760 57040 1880
rect 57060 1760 57080 1880
rect 57100 1760 57105 1880
rect 57035 1750 57105 1760
rect 57130 1880 57160 1890
rect 57130 1760 57135 1880
rect 57155 1760 57160 1880
rect 57130 1750 57160 1760
rect 57185 1880 57215 1890
rect 57185 1760 57190 1880
rect 57210 1760 57215 1880
rect 57185 1750 57215 1760
rect 57240 1880 57270 1890
rect 57240 1760 57245 1880
rect 57265 1760 57270 1880
rect 57240 1750 57270 1760
rect 57295 1880 57325 1890
rect 57295 1760 57300 1880
rect 57320 1760 57325 1880
rect 57295 1750 57325 1760
rect 57350 1880 57380 1890
rect 57350 1760 57355 1880
rect 57375 1760 57380 1880
rect 57350 1750 57380 1760
rect 57405 1880 57435 1890
rect 57405 1760 57410 1880
rect 57430 1760 57435 1880
rect 57405 1750 57435 1760
rect 57460 1880 57490 1890
rect 57460 1760 57465 1880
rect 57485 1760 57490 1880
rect 57460 1750 57490 1760
rect 57515 1880 57545 1890
rect 57515 1760 57520 1880
rect 57540 1760 57545 1880
rect 57515 1750 57545 1760
rect 57570 1880 57600 1890
rect 57570 1760 57575 1880
rect 57595 1760 57600 1880
rect 57570 1750 57600 1760
rect 57625 1880 57655 1890
rect 57625 1760 57630 1880
rect 57650 1760 57655 1880
rect 57625 1750 57655 1760
rect 57680 1880 57710 1890
rect 57680 1760 57685 1880
rect 57705 1760 57710 1880
rect 57680 1750 57710 1760
rect 57735 1880 57805 1890
rect 57735 1760 57740 1880
rect 57760 1760 57780 1880
rect 57800 1760 57805 1880
rect 57735 1750 57805 1760
rect 58445 1865 58515 1875
rect 55285 1685 55355 1695
rect 56035 1720 56065 1750
rect 56035 1700 56040 1720
rect 56060 1700 56065 1720
rect 56035 1690 56065 1700
rect 56695 1720 56725 1730
rect 56695 1700 56700 1720
rect 56720 1700 56725 1720
rect 56695 1690 56725 1700
rect 57075 1720 57105 1730
rect 57075 1700 57080 1720
rect 57100 1700 57105 1720
rect 57075 1690 57105 1700
rect 57735 1720 57765 1750
rect 57735 1700 57740 1720
rect 57760 1700 57765 1720
rect 57735 1690 57765 1700
rect 58445 1695 58450 1865
rect 58470 1695 58490 1865
rect 58510 1695 58515 1865
rect 58445 1685 58515 1695
rect 58540 1865 58570 1875
rect 58540 1695 58545 1865
rect 58565 1695 58570 1865
rect 58540 1685 58570 1695
rect 58595 1865 58625 1875
rect 58595 1695 58600 1865
rect 58620 1695 58625 1865
rect 58595 1685 58625 1695
rect 58650 1865 58680 1875
rect 58650 1695 58655 1865
rect 58675 1695 58680 1865
rect 58650 1685 58680 1695
rect 58705 1865 58735 1875
rect 58705 1695 58710 1865
rect 58730 1695 58735 1865
rect 58705 1685 58735 1695
rect 58760 1865 58790 1875
rect 58760 1695 58765 1865
rect 58785 1695 58790 1865
rect 58760 1685 58790 1695
rect 58815 1865 58845 1875
rect 58815 1695 58820 1865
rect 58840 1695 58845 1865
rect 58815 1685 58845 1695
rect 58870 1865 58900 1875
rect 58870 1695 58875 1865
rect 58895 1695 58900 1865
rect 58870 1685 58900 1695
rect 58925 1865 58955 1875
rect 58925 1695 58930 1865
rect 58950 1695 58955 1865
rect 58925 1685 58955 1695
rect 58980 1865 59010 1875
rect 58980 1695 58985 1865
rect 59005 1695 59010 1865
rect 58980 1685 59010 1695
rect 59035 1865 59065 1875
rect 59035 1695 59040 1865
rect 59060 1695 59065 1865
rect 59035 1685 59065 1695
rect 59090 1865 59120 1875
rect 59090 1695 59095 1865
rect 59115 1695 59120 1865
rect 59090 1685 59120 1695
rect 59145 1865 59215 1875
rect 59145 1695 59150 1865
rect 59170 1695 59190 1865
rect 59210 1695 59215 1865
rect 59145 1685 59215 1695
rect 59330 1781 59545 1801
rect 59330 1764 59365 1781
rect 59510 1764 59545 1781
rect 54730 1655 54770 1665
rect 54730 1635 54740 1655
rect 54760 1635 54770 1655
rect 54730 1625 54770 1635
rect 54840 1655 54880 1665
rect 54840 1635 54850 1655
rect 54870 1635 54880 1655
rect 54840 1625 54880 1635
rect 54950 1655 54990 1665
rect 54950 1635 54960 1655
rect 54980 1635 54990 1655
rect 54950 1625 54990 1635
rect 55060 1655 55100 1665
rect 55060 1635 55070 1655
rect 55090 1635 55100 1655
rect 55060 1625 55100 1635
rect 55120 1655 55150 1665
rect 55120 1635 55125 1655
rect 55145 1635 55150 1655
rect 55120 1625 55150 1635
rect 55170 1655 55210 1665
rect 55170 1635 55180 1655
rect 55200 1635 55210 1655
rect 55170 1625 55210 1635
rect 58590 1655 58630 1665
rect 58590 1635 58600 1655
rect 58620 1635 58630 1655
rect 58590 1625 58630 1635
rect 58650 1655 58680 1665
rect 58650 1635 58655 1655
rect 58675 1635 58680 1655
rect 58650 1625 58680 1635
rect 58700 1655 58740 1665
rect 58700 1635 58710 1655
rect 58730 1635 58740 1655
rect 58700 1625 58740 1635
rect 58810 1655 58850 1665
rect 58810 1635 58820 1655
rect 58840 1635 58850 1655
rect 58810 1625 58850 1635
rect 58920 1655 58960 1665
rect 58920 1635 58930 1655
rect 58950 1635 58960 1655
rect 58920 1625 58960 1635
rect 59030 1655 59070 1665
rect 59030 1635 59040 1655
rect 59060 1635 59070 1655
rect 59030 1625 59070 1635
rect 55115 1590 55155 1600
rect 55115 1570 55125 1590
rect 55145 1570 55155 1590
rect 55115 1550 55155 1570
rect 55115 1530 55125 1550
rect 55145 1530 55155 1550
rect 55115 1520 55155 1530
rect 58645 1590 58685 1600
rect 58645 1570 58655 1590
rect 58675 1570 58685 1590
rect 58645 1550 58685 1570
rect 58645 1530 58655 1550
rect 58675 1530 58685 1550
rect 59425 1714 59450 1764
rect 58645 1520 58685 1530
rect 55120 1485 55150 1495
rect 55120 1465 55125 1485
rect 55145 1465 55150 1485
rect 55120 1455 55150 1465
rect 58650 1485 58680 1495
rect 58650 1465 58655 1485
rect 58675 1465 58680 1485
rect 58650 1455 58680 1465
rect 54585 1425 54655 1435
rect 54255 1155 54290 1165
rect 54255 1130 54260 1155
rect 54285 1130 54290 1155
rect 54255 1120 54290 1130
rect 54315 1155 54350 1165
rect 54315 1130 54320 1155
rect 54345 1130 54350 1155
rect 54315 1120 54350 1130
rect 54375 1155 54410 1165
rect 54375 1130 54380 1155
rect 54405 1130 54410 1155
rect 54375 1120 54410 1130
rect 54435 1155 54470 1165
rect 54435 1130 54440 1155
rect 54465 1130 54470 1155
rect 54585 1155 54590 1425
rect 54610 1155 54630 1425
rect 54650 1155 54655 1425
rect 54585 1145 54655 1155
rect 54680 1425 54710 1435
rect 54680 1155 54685 1425
rect 54705 1155 54710 1425
rect 54680 1145 54710 1155
rect 54735 1425 54765 1435
rect 54735 1155 54740 1425
rect 54760 1155 54765 1425
rect 54735 1145 54765 1155
rect 54790 1425 54820 1435
rect 54790 1155 54795 1425
rect 54815 1155 54820 1425
rect 54790 1145 54820 1155
rect 54845 1425 54875 1435
rect 54845 1155 54850 1425
rect 54870 1155 54875 1425
rect 54845 1145 54875 1155
rect 54900 1425 54930 1435
rect 54900 1155 54905 1425
rect 54925 1155 54930 1425
rect 54900 1145 54930 1155
rect 54955 1425 54985 1435
rect 54955 1155 54960 1425
rect 54980 1155 54985 1425
rect 54955 1145 54985 1155
rect 55010 1425 55040 1435
rect 55010 1155 55015 1425
rect 55035 1155 55040 1425
rect 55010 1145 55040 1155
rect 55065 1425 55095 1435
rect 55065 1155 55070 1425
rect 55090 1155 55095 1425
rect 55065 1145 55095 1155
rect 55120 1425 55150 1435
rect 55120 1155 55125 1425
rect 55145 1155 55150 1425
rect 55120 1145 55150 1155
rect 55175 1425 55205 1435
rect 55175 1155 55180 1425
rect 55200 1155 55205 1425
rect 55175 1145 55205 1155
rect 55230 1425 55260 1435
rect 55230 1155 55235 1425
rect 55255 1155 55260 1425
rect 55230 1145 55260 1155
rect 55285 1425 55355 1435
rect 55285 1155 55290 1425
rect 55310 1155 55330 1425
rect 55350 1155 55355 1425
rect 58445 1425 58515 1435
rect 56690 1300 56720 1310
rect 56040 1290 56070 1300
rect 56040 1270 56045 1290
rect 56065 1270 56070 1290
rect 56690 1280 56695 1300
rect 56715 1280 56720 1300
rect 56690 1270 56720 1280
rect 56840 1300 56870 1310
rect 56840 1280 56845 1300
rect 56865 1280 56870 1300
rect 56840 1270 56870 1280
rect 56930 1300 56960 1310
rect 56930 1280 56935 1300
rect 56955 1280 56960 1300
rect 56930 1270 56960 1280
rect 57080 1300 57110 1310
rect 57080 1280 57085 1300
rect 57105 1280 57110 1300
rect 57080 1270 57110 1280
rect 57730 1290 57760 1300
rect 57730 1270 57735 1290
rect 57755 1270 57760 1290
rect 56040 1260 56070 1270
rect 57730 1260 57760 1270
rect 55285 1145 55355 1155
rect 55995 1205 56065 1215
rect 54435 1120 54470 1130
rect 54625 1115 54655 1125
rect 54625 1095 54630 1115
rect 54650 1095 54655 1115
rect 54625 1080 54655 1095
rect 55285 1115 55315 1125
rect 55285 1095 55290 1115
rect 55310 1095 55315 1115
rect 55285 1080 55315 1095
rect 55995 1085 56000 1205
rect 56020 1085 56040 1205
rect 56060 1085 56065 1205
rect 55995 1075 56065 1085
rect 56090 1205 56120 1215
rect 56090 1085 56095 1205
rect 56115 1085 56120 1205
rect 56090 1075 56120 1085
rect 56145 1205 56175 1215
rect 56145 1085 56150 1205
rect 56170 1085 56175 1205
rect 56145 1075 56175 1085
rect 56200 1205 56230 1215
rect 56200 1085 56205 1205
rect 56225 1085 56230 1205
rect 56200 1075 56230 1085
rect 56255 1205 56285 1215
rect 56255 1085 56260 1205
rect 56280 1085 56285 1205
rect 56255 1075 56285 1085
rect 56310 1205 56340 1215
rect 56310 1085 56315 1205
rect 56335 1085 56340 1205
rect 56310 1075 56340 1085
rect 56365 1205 56395 1215
rect 56365 1085 56370 1205
rect 56390 1085 56395 1205
rect 56365 1075 56395 1085
rect 56420 1205 56450 1215
rect 56420 1085 56425 1205
rect 56445 1085 56450 1205
rect 56420 1075 56450 1085
rect 56475 1205 56505 1215
rect 56475 1085 56480 1205
rect 56500 1085 56505 1205
rect 56475 1075 56505 1085
rect 56530 1205 56560 1215
rect 56530 1085 56535 1205
rect 56555 1085 56560 1205
rect 56530 1075 56560 1085
rect 56585 1205 56615 1215
rect 56585 1085 56590 1205
rect 56610 1085 56615 1205
rect 56585 1075 56615 1085
rect 56640 1205 56670 1215
rect 56640 1085 56645 1205
rect 56665 1085 56670 1205
rect 56640 1075 56670 1085
rect 56695 1205 56805 1215
rect 56695 1085 56700 1205
rect 56720 1085 56740 1205
rect 56760 1085 56780 1205
rect 56800 1085 56805 1205
rect 56695 1075 56805 1085
rect 56830 1205 56860 1215
rect 56830 1085 56835 1205
rect 56855 1085 56860 1205
rect 56830 1075 56860 1085
rect 56885 1205 56915 1215
rect 56885 1085 56890 1205
rect 56910 1085 56915 1205
rect 56885 1075 56915 1085
rect 56940 1205 56970 1215
rect 56940 1085 56945 1205
rect 56965 1085 56970 1205
rect 56940 1075 56970 1085
rect 56995 1205 57105 1215
rect 56995 1085 57000 1205
rect 57020 1085 57040 1205
rect 57060 1085 57080 1205
rect 57100 1085 57105 1205
rect 56995 1075 57105 1085
rect 57130 1205 57160 1215
rect 57130 1085 57135 1205
rect 57155 1085 57160 1205
rect 57130 1075 57160 1085
rect 57185 1205 57215 1215
rect 57185 1085 57190 1205
rect 57210 1085 57215 1205
rect 57185 1075 57215 1085
rect 57240 1205 57270 1215
rect 57240 1085 57245 1205
rect 57265 1085 57270 1205
rect 57240 1075 57270 1085
rect 57295 1205 57325 1215
rect 57295 1085 57300 1205
rect 57320 1085 57325 1205
rect 57295 1075 57325 1085
rect 57350 1205 57380 1215
rect 57350 1085 57355 1205
rect 57375 1085 57380 1205
rect 57350 1075 57380 1085
rect 57405 1205 57435 1215
rect 57405 1085 57410 1205
rect 57430 1085 57435 1205
rect 57405 1075 57435 1085
rect 57460 1205 57490 1215
rect 57460 1085 57465 1205
rect 57485 1085 57490 1205
rect 57460 1075 57490 1085
rect 57515 1205 57545 1215
rect 57515 1085 57520 1205
rect 57540 1085 57545 1205
rect 57515 1075 57545 1085
rect 57570 1205 57600 1215
rect 57570 1085 57575 1205
rect 57595 1085 57600 1205
rect 57570 1075 57600 1085
rect 57625 1205 57655 1215
rect 57625 1085 57630 1205
rect 57650 1085 57655 1205
rect 57625 1075 57655 1085
rect 57680 1205 57710 1215
rect 57680 1085 57685 1205
rect 57705 1085 57710 1205
rect 57680 1075 57710 1085
rect 57735 1205 57805 1215
rect 57735 1085 57740 1205
rect 57760 1085 57780 1205
rect 57800 1085 57805 1205
rect 58445 1155 58450 1425
rect 58470 1155 58490 1425
rect 58510 1155 58515 1425
rect 58445 1145 58515 1155
rect 58540 1425 58570 1435
rect 58540 1155 58545 1425
rect 58565 1155 58570 1425
rect 58540 1145 58570 1155
rect 58595 1425 58625 1435
rect 58595 1155 58600 1425
rect 58620 1155 58625 1425
rect 58595 1145 58625 1155
rect 58650 1425 58680 1435
rect 58650 1155 58655 1425
rect 58675 1155 58680 1425
rect 58650 1145 58680 1155
rect 58705 1425 58735 1435
rect 58705 1155 58710 1425
rect 58730 1155 58735 1425
rect 58705 1145 58735 1155
rect 58760 1425 58790 1435
rect 58760 1155 58765 1425
rect 58785 1155 58790 1425
rect 58760 1145 58790 1155
rect 58815 1425 58845 1435
rect 58815 1155 58820 1425
rect 58840 1155 58845 1425
rect 58815 1145 58845 1155
rect 58870 1425 58900 1435
rect 58870 1155 58875 1425
rect 58895 1155 58900 1425
rect 58870 1145 58900 1155
rect 58925 1425 58955 1435
rect 58925 1155 58930 1425
rect 58950 1155 58955 1425
rect 58925 1145 58955 1155
rect 58980 1425 59010 1435
rect 58980 1155 58985 1425
rect 59005 1155 59010 1425
rect 58980 1145 59010 1155
rect 59035 1425 59065 1435
rect 59035 1155 59040 1425
rect 59060 1155 59065 1425
rect 59035 1145 59065 1155
rect 59090 1425 59120 1435
rect 59090 1155 59095 1425
rect 59115 1155 59120 1425
rect 59090 1145 59120 1155
rect 59145 1425 59215 1435
rect 59145 1155 59150 1425
rect 59170 1155 59190 1425
rect 59210 1155 59215 1425
rect 59145 1145 59215 1155
rect 59330 1155 59365 1165
rect 59330 1130 59335 1155
rect 59360 1130 59365 1155
rect 57735 1075 57805 1085
rect 58485 1115 58515 1125
rect 58485 1095 58490 1115
rect 58510 1095 58515 1115
rect 58485 1080 58515 1095
rect 59145 1115 59175 1125
rect 59330 1120 59365 1130
rect 59390 1155 59425 1165
rect 59390 1130 59395 1155
rect 59420 1130 59425 1155
rect 59390 1120 59425 1130
rect 59450 1155 59485 1165
rect 59450 1130 59455 1155
rect 59480 1130 59485 1155
rect 59450 1120 59485 1130
rect 59510 1155 59545 1165
rect 59510 1130 59515 1155
rect 59540 1130 59545 1155
rect 59510 1120 59545 1130
rect 59145 1095 59150 1115
rect 59170 1095 59175 1115
rect 59145 1085 59175 1095
rect 56040 1055 56065 1075
rect 56035 1045 56065 1055
rect 56035 1025 56040 1045
rect 56060 1025 56065 1045
rect 56035 1015 56065 1025
rect 56735 1045 56765 1055
rect 56735 1025 56740 1045
rect 56760 1025 56765 1045
rect 56735 1015 56765 1025
rect 57035 1045 57065 1055
rect 57035 1025 57040 1045
rect 57060 1025 57065 1045
rect 57035 1015 57065 1025
rect 57735 1045 57765 1075
rect 57735 1025 57740 1045
rect 57760 1025 57765 1045
rect 57735 1015 57765 1025
rect 55000 520 55040 530
rect 55000 500 55010 520
rect 55030 500 55040 520
rect 55000 490 55040 500
rect 58760 520 58800 530
rect 58760 500 58770 520
rect 58790 500 58800 520
rect 58760 490 58800 500
rect 56825 465 56865 475
rect 56825 445 56835 465
rect 56855 445 56865 465
rect 56825 435 56865 445
rect 56935 465 56975 475
rect 56935 445 56945 465
rect 56965 445 56975 465
rect 56935 435 56975 445
rect 56185 405 56255 415
rect 54325 330 54360 340
rect 54325 305 54330 330
rect 54355 305 54360 330
rect 54325 295 54360 305
rect 54385 330 54420 340
rect 54385 305 54390 330
rect 54415 305 54420 330
rect 54385 295 54420 305
rect 54615 325 54685 335
rect 54360 -392 54385 -342
rect 54615 -345 54620 325
rect 54640 -345 54660 325
rect 54680 -345 54685 325
rect 54615 -355 54685 -345
rect 54755 325 54785 335
rect 54755 -345 54760 325
rect 54780 -345 54785 325
rect 54755 -355 54785 -345
rect 54855 325 54885 335
rect 54855 -345 54860 325
rect 54880 -345 54885 325
rect 54855 -355 54885 -345
rect 54955 325 54985 335
rect 54955 -345 54960 325
rect 54980 -345 54985 325
rect 54955 -355 54985 -345
rect 55055 325 55085 335
rect 55055 -345 55060 325
rect 55080 -345 55085 325
rect 55055 -355 55085 -345
rect 55155 325 55185 335
rect 55155 -345 55160 325
rect 55180 -345 55185 325
rect 55155 -355 55185 -345
rect 55255 325 55325 335
rect 55255 -345 55260 325
rect 55280 -345 55300 325
rect 55320 -345 55325 325
rect 56185 185 56190 405
rect 56210 185 56230 405
rect 56250 185 56255 405
rect 56185 175 56255 185
rect 56280 405 56310 415
rect 56280 185 56285 405
rect 56305 185 56310 405
rect 56280 175 56310 185
rect 56335 405 56365 415
rect 56335 185 56340 405
rect 56360 185 56365 405
rect 56335 175 56365 185
rect 56390 405 56420 415
rect 56390 185 56395 405
rect 56415 185 56420 405
rect 56390 175 56420 185
rect 56445 405 56475 415
rect 56445 185 56450 405
rect 56470 185 56475 405
rect 56445 175 56475 185
rect 56500 405 56530 415
rect 56500 185 56505 405
rect 56525 185 56530 405
rect 56500 175 56530 185
rect 56555 405 56585 415
rect 56555 185 56560 405
rect 56580 185 56585 405
rect 56555 175 56585 185
rect 56610 405 56640 415
rect 56610 185 56615 405
rect 56635 185 56640 405
rect 56610 175 56640 185
rect 56665 405 56695 415
rect 56665 185 56670 405
rect 56690 185 56695 405
rect 56665 175 56695 185
rect 56720 405 56750 415
rect 56720 185 56725 405
rect 56745 185 56750 405
rect 56720 175 56750 185
rect 56775 405 56805 415
rect 56775 185 56780 405
rect 56800 185 56805 405
rect 56775 175 56805 185
rect 56830 405 56860 415
rect 56830 185 56835 405
rect 56855 185 56860 405
rect 56830 175 56860 185
rect 56885 405 56915 415
rect 56885 185 56890 405
rect 56910 185 56915 405
rect 56885 175 56915 185
rect 56940 405 56970 415
rect 56940 185 56945 405
rect 56965 185 56970 405
rect 56940 175 56970 185
rect 56995 405 57025 415
rect 56995 185 57000 405
rect 57020 185 57025 405
rect 56995 175 57025 185
rect 57050 405 57080 415
rect 57050 185 57055 405
rect 57075 185 57080 405
rect 57050 175 57080 185
rect 57105 405 57135 415
rect 57105 185 57110 405
rect 57130 185 57135 405
rect 57105 175 57135 185
rect 57160 405 57190 415
rect 57160 185 57165 405
rect 57185 185 57190 405
rect 57160 175 57190 185
rect 57215 405 57245 415
rect 57215 185 57220 405
rect 57240 185 57245 405
rect 57215 175 57245 185
rect 57270 405 57300 415
rect 57270 185 57275 405
rect 57295 185 57300 405
rect 57270 175 57300 185
rect 57325 405 57355 415
rect 57325 185 57330 405
rect 57350 185 57355 405
rect 57325 175 57355 185
rect 57380 405 57410 415
rect 57380 185 57385 405
rect 57405 185 57410 405
rect 57380 175 57410 185
rect 57435 405 57465 415
rect 57435 185 57440 405
rect 57460 185 57465 405
rect 57435 175 57465 185
rect 57490 405 57560 415
rect 57490 185 57495 405
rect 57515 185 57535 405
rect 57555 185 57560 405
rect 57490 175 57560 185
rect 58475 325 58545 335
rect 56220 145 56260 155
rect 56220 125 56230 145
rect 56250 125 56260 145
rect 56220 115 56260 125
rect 57485 145 57525 155
rect 57485 125 57495 145
rect 57515 125 57525 145
rect 57485 115 57525 125
rect 57415 35 57455 45
rect 57415 15 57425 35
rect 57445 15 57455 35
rect 57415 5 57455 15
rect 56595 -255 56635 -245
rect 56595 -275 56605 -255
rect 56625 -275 56635 -255
rect 56595 -285 56635 -275
rect 56920 -255 56960 -245
rect 56920 -275 56930 -255
rect 56950 -275 56960 -255
rect 56920 -285 56960 -275
rect 57040 -255 57080 -245
rect 57040 -275 57050 -255
rect 57070 -275 57080 -255
rect 57040 -285 57080 -275
rect 57160 -255 57200 -245
rect 57160 -275 57170 -255
rect 57190 -275 57200 -255
rect 57160 -285 57200 -275
rect 55255 -355 55325 -345
rect 56395 -315 56465 -305
rect 54655 -385 54685 -375
rect 54655 -405 54660 -385
rect 54680 -405 54685 -385
rect 54655 -415 54685 -405
rect 55255 -385 55285 -375
rect 55255 -405 55260 -385
rect 55280 -405 55285 -385
rect 55255 -415 55285 -405
rect 56395 -435 56400 -315
rect 56420 -435 56440 -315
rect 56460 -435 56465 -315
rect 56395 -445 56465 -435
rect 56490 -315 56520 -305
rect 56490 -435 56495 -315
rect 56515 -435 56520 -315
rect 56490 -445 56520 -435
rect 56545 -315 56575 -305
rect 56545 -435 56550 -315
rect 56570 -435 56575 -315
rect 56545 -445 56575 -435
rect 56600 -315 56630 -305
rect 56600 -435 56605 -315
rect 56625 -435 56630 -315
rect 56600 -445 56630 -435
rect 56655 -315 56685 -305
rect 56655 -435 56660 -315
rect 56680 -435 56685 -315
rect 56655 -445 56685 -435
rect 56710 -315 56740 -305
rect 56710 -435 56715 -315
rect 56735 -435 56740 -315
rect 56710 -445 56740 -435
rect 56765 -315 56835 -305
rect 56765 -435 56770 -315
rect 56790 -435 56810 -315
rect 56830 -435 56835 -315
rect 56765 -445 56835 -435
rect 56875 -315 56905 -305
rect 56875 -435 56880 -315
rect 56900 -435 56905 -315
rect 57215 -325 57245 -315
rect 57215 -425 57220 -325
rect 57240 -425 57245 -325
rect 58475 -345 58480 325
rect 58500 -345 58520 325
rect 58540 -345 58545 325
rect 58475 -355 58545 -345
rect 58615 325 58645 335
rect 58615 -345 58620 325
rect 58640 -345 58645 325
rect 58615 -355 58645 -345
rect 58715 325 58745 335
rect 58715 -345 58720 325
rect 58740 -345 58745 325
rect 58715 -355 58745 -345
rect 58815 325 58845 335
rect 58815 -345 58820 325
rect 58840 -345 58845 325
rect 58815 -355 58845 -345
rect 58915 325 58945 335
rect 58915 -345 58920 325
rect 58940 -345 58945 325
rect 58915 -355 58945 -345
rect 59015 325 59045 335
rect 59015 -345 59020 325
rect 59040 -345 59045 325
rect 59015 -355 59045 -345
rect 59115 325 59185 335
rect 59115 -345 59120 325
rect 59140 -345 59160 325
rect 59180 -345 59185 325
rect 59380 330 59415 340
rect 59380 305 59385 330
rect 59410 305 59415 330
rect 59380 295 59415 305
rect 59440 330 59475 340
rect 59440 305 59445 330
rect 59470 305 59475 330
rect 59440 295 59475 305
rect 59115 -355 59185 -345
rect 58515 -385 58545 -375
rect 58515 -405 58520 -385
rect 58540 -405 58545 -385
rect 58515 -415 58545 -405
rect 59115 -385 59145 -375
rect 59115 -405 59120 -385
rect 59140 -405 59145 -385
rect 59415 -392 59440 -342
rect 59115 -415 59145 -405
rect 57215 -435 57245 -425
rect 56875 -445 56905 -435
rect 56435 -475 56465 -465
rect 56435 -495 56440 -475
rect 56460 -495 56465 -475
rect 56435 -505 56465 -495
rect 56765 -475 56795 -465
rect 56765 -495 56770 -475
rect 56790 -495 56795 -475
rect 56765 -505 56795 -495
rect 56920 -475 56960 -465
rect 56920 -495 56930 -475
rect 56950 -495 56960 -475
rect 56920 -505 56960 -495
rect 57040 -475 57080 -465
rect 57040 -495 57050 -475
rect 57070 -495 57080 -475
rect 57040 -505 57080 -495
rect 57160 -475 57200 -465
rect 57160 -495 57170 -475
rect 57190 -495 57200 -475
rect 57160 -505 57200 -495
<< viali >>
rect 56095 4905 56115 4925
rect 56275 4905 56295 4925
rect 57035 4905 57055 4925
rect 57215 4905 57235 4925
rect 57505 4905 57525 4925
rect 57685 4905 57705 4925
rect 56095 4545 56115 4865
rect 56155 4545 56175 4865
rect 56215 4545 56235 4865
rect 56275 4545 56295 4865
rect 56565 4735 56585 4755
rect 56745 4735 56765 4755
rect 56565 4545 56585 4695
rect 56625 4545 56645 4695
rect 56685 4545 56705 4695
rect 56745 4545 56765 4695
rect 57035 4545 57055 4865
rect 57095 4545 57115 4865
rect 57155 4545 57175 4865
rect 57215 4545 57235 4865
rect 57505 4545 57525 4865
rect 57565 4545 57585 4865
rect 57625 4545 57645 4865
rect 57685 4545 57705 4865
rect 56160 4455 56180 4475
rect 56635 4455 56655 4475
rect 57145 4455 57165 4475
rect 57581 4445 57601 4465
rect 54600 3680 54620 4000
rect 54660 3680 54680 4000
rect 54720 3680 54740 4000
rect 54780 3680 54800 4000
rect 54840 3680 54860 4000
rect 54900 3680 54920 4000
rect 54960 3680 54980 4000
rect 55020 3680 55040 4000
rect 55080 3680 55100 4000
rect 55140 3680 55160 4000
rect 55200 3680 55220 4000
rect 55260 3680 55280 4000
rect 55320 3680 55340 4000
rect 56015 3680 56035 4000
rect 56075 3680 56095 4000
rect 56135 3680 56155 4000
rect 56195 3680 56215 4000
rect 56255 3680 56275 4000
rect 56315 3680 56335 4000
rect 56375 3680 56395 4000
rect 56435 3680 56455 4000
rect 56495 3680 56515 4000
rect 56555 3680 56575 4000
rect 56615 3680 56635 4000
rect 56675 3680 56695 4000
rect 56735 3680 56755 4000
rect 57045 3680 57065 4000
rect 57105 3680 57125 4000
rect 57165 3680 57185 4000
rect 57225 3680 57245 4000
rect 57285 3680 57305 4000
rect 57345 3680 57365 4000
rect 57405 3680 57425 4000
rect 57465 3680 57485 4000
rect 57525 3680 57545 4000
rect 57585 3680 57605 4000
rect 57645 3680 57665 4000
rect 57705 3680 57725 4000
rect 57765 3680 57785 4000
rect 58460 3680 58480 4000
rect 58520 3680 58540 4000
rect 58580 3680 58600 4000
rect 58640 3680 58660 4000
rect 58700 3680 58720 4000
rect 58760 3680 58780 4000
rect 58820 3680 58840 4000
rect 58880 3680 58900 4000
rect 58940 3680 58960 4000
rect 59000 3680 59020 4000
rect 59060 3680 59080 4000
rect 59120 3680 59140 4000
rect 59180 3680 59200 4000
rect 54600 3620 54620 3640
rect 55320 3620 55340 3640
rect 56015 3620 56035 3640
rect 56735 3620 56755 3640
rect 57045 3620 57065 3640
rect 57765 3620 57785 3640
rect 58460 3620 58480 3640
rect 59180 3620 59200 3640
rect 56375 3555 56395 3575
rect 57405 3555 57425 3575
rect 54960 3510 54980 3530
rect 58820 3510 58840 3530
rect 56520 3250 56540 3270
rect 56685 3250 56705 3270
rect 56850 3250 56870 3270
rect 56930 3250 56950 3270
rect 57095 3250 57115 3270
rect 57260 3250 57280 3270
rect 54210 3170 54230 3190
rect 54265 3170 54285 3190
rect 54320 3170 54340 3190
rect 54630 3180 54650 3200
rect 55290 3180 55310 3200
rect 56630 3195 56650 3215
rect 56740 3195 56760 3215
rect 57040 3195 57060 3215
rect 57150 3195 57170 3215
rect 58490 3180 58510 3200
rect 59150 3180 59170 3200
rect 59460 3170 59480 3190
rect 59515 3170 59535 3190
rect 59570 3170 59590 3190
rect 54210 2565 54230 2585
rect 54265 2565 54285 2585
rect 54320 2565 54340 2585
rect 54630 2570 54650 3140
rect 54685 2570 54705 3140
rect 54740 2570 54760 3140
rect 54795 2570 54815 3140
rect 54850 2570 54870 3140
rect 54905 2570 54925 3140
rect 54960 2570 54980 3140
rect 55015 2570 55035 3140
rect 55070 2570 55090 3140
rect 55125 2570 55145 3140
rect 55180 2570 55200 3140
rect 55235 2570 55255 3140
rect 55290 2570 55310 3140
rect 56565 2885 56585 2905
rect 56612 2875 56632 2895
rect 56685 2875 56705 2895
rect 56758 2875 56778 2895
rect 56805 2885 56825 2905
rect 56975 2885 56995 2905
rect 57022 2875 57042 2895
rect 57095 2875 57115 2895
rect 57168 2875 57188 2895
rect 57215 2885 57235 2905
rect 56610 2805 56630 2825
rect 57170 2805 57190 2825
rect 56860 2590 56880 2610
rect 56945 2590 56965 2610
rect 58490 2570 58510 3140
rect 58545 2570 58565 3140
rect 58600 2570 58620 3140
rect 58655 2570 58675 3140
rect 58710 2570 58730 3140
rect 58765 2570 58785 3140
rect 58820 2570 58840 3140
rect 58875 2570 58895 3140
rect 58930 2570 58950 3140
rect 58985 2570 59005 3140
rect 59040 2570 59060 3140
rect 59095 2570 59115 3140
rect 59150 2570 59170 3140
rect 59460 2565 59480 2585
rect 59515 2565 59535 2585
rect 59570 2565 59590 2585
rect 54960 2445 54980 2465
rect 54960 2405 54980 2425
rect 54960 2365 54980 2385
rect 56780 2330 56800 2550
rect 56835 2330 56855 2550
rect 56890 2330 56910 2550
rect 56945 2330 56965 2550
rect 57000 2330 57020 2550
rect 58820 2445 58840 2465
rect 58820 2405 58840 2425
rect 58820 2365 58840 2385
rect 56780 2270 56800 2290
rect 57000 2270 57020 2290
rect 56045 1960 56065 1980
rect 56695 1960 56715 1980
rect 57085 1960 57105 1980
rect 57735 1960 57755 1980
rect 54630 1905 54650 1925
rect 55290 1905 55310 1925
rect 58490 1905 58510 1925
rect 59150 1905 59170 1925
rect 54630 1695 54650 1865
rect 54685 1695 54705 1865
rect 54740 1695 54760 1865
rect 54795 1695 54815 1865
rect 54850 1695 54870 1865
rect 54905 1695 54925 1865
rect 54960 1695 54980 1865
rect 55015 1695 55035 1865
rect 55070 1695 55090 1865
rect 55125 1695 55145 1865
rect 55180 1695 55200 1865
rect 55235 1695 55255 1865
rect 55290 1695 55310 1865
rect 56040 1760 56060 1880
rect 56095 1760 56115 1880
rect 56150 1760 56170 1880
rect 56205 1760 56225 1880
rect 56260 1760 56280 1880
rect 56315 1760 56335 1880
rect 56370 1760 56390 1880
rect 56425 1760 56445 1880
rect 56480 1760 56500 1880
rect 56535 1760 56555 1880
rect 56590 1760 56610 1880
rect 56645 1760 56665 1880
rect 56700 1760 56720 1880
rect 57080 1760 57100 1880
rect 57135 1760 57155 1880
rect 57190 1760 57210 1880
rect 57245 1760 57265 1880
rect 57300 1760 57320 1880
rect 57355 1760 57375 1880
rect 57410 1760 57430 1880
rect 57465 1760 57485 1880
rect 57520 1760 57540 1880
rect 57575 1760 57595 1880
rect 57630 1760 57650 1880
rect 57685 1760 57705 1880
rect 57740 1760 57760 1880
rect 56040 1700 56060 1720
rect 56700 1700 56720 1720
rect 57080 1700 57100 1720
rect 57740 1700 57760 1720
rect 58490 1695 58510 1865
rect 58545 1695 58565 1865
rect 58600 1695 58620 1865
rect 58655 1695 58675 1865
rect 58710 1695 58730 1865
rect 58765 1695 58785 1865
rect 58820 1695 58840 1865
rect 58875 1695 58895 1865
rect 58930 1695 58950 1865
rect 58985 1695 59005 1865
rect 59040 1695 59060 1865
rect 59095 1695 59115 1865
rect 59150 1695 59170 1865
rect 54740 1635 54760 1655
rect 54850 1635 54870 1655
rect 54960 1635 54980 1655
rect 55070 1635 55090 1655
rect 55180 1635 55200 1655
rect 58600 1635 58620 1655
rect 58710 1635 58730 1655
rect 58820 1635 58840 1655
rect 58930 1635 58950 1655
rect 59040 1635 59060 1655
rect 55125 1570 55145 1590
rect 55125 1530 55145 1550
rect 58655 1570 58675 1590
rect 58655 1530 58675 1550
rect 54260 1130 54285 1155
rect 54320 1130 54345 1155
rect 54380 1130 54405 1155
rect 54440 1130 54465 1155
rect 54630 1155 54650 1425
rect 54685 1155 54705 1425
rect 54740 1155 54760 1425
rect 54795 1155 54815 1425
rect 54850 1155 54870 1425
rect 54905 1155 54925 1425
rect 54960 1155 54980 1425
rect 55015 1155 55035 1425
rect 55070 1155 55090 1425
rect 55125 1155 55145 1425
rect 55180 1155 55200 1425
rect 55235 1155 55255 1425
rect 55290 1155 55310 1425
rect 56045 1270 56065 1290
rect 56695 1280 56715 1300
rect 56845 1280 56865 1300
rect 56935 1280 56955 1300
rect 57085 1280 57105 1300
rect 57735 1270 57755 1290
rect 54630 1095 54650 1115
rect 55290 1095 55310 1115
rect 56040 1085 56060 1205
rect 56095 1085 56115 1205
rect 56150 1085 56170 1205
rect 56205 1085 56225 1205
rect 56260 1085 56280 1205
rect 56315 1085 56335 1205
rect 56370 1085 56390 1205
rect 56425 1085 56445 1205
rect 56480 1085 56500 1205
rect 56535 1085 56555 1205
rect 56590 1085 56610 1205
rect 56645 1085 56665 1205
rect 56700 1085 56720 1205
rect 56780 1085 56800 1205
rect 56835 1085 56855 1205
rect 56890 1085 56910 1205
rect 56945 1085 56965 1205
rect 57000 1085 57020 1205
rect 57080 1085 57100 1205
rect 57135 1085 57155 1205
rect 57190 1085 57210 1205
rect 57245 1085 57265 1205
rect 57300 1085 57320 1205
rect 57355 1085 57375 1205
rect 57410 1085 57430 1205
rect 57465 1085 57485 1205
rect 57520 1085 57540 1205
rect 57575 1085 57595 1205
rect 57630 1085 57650 1205
rect 57685 1085 57705 1205
rect 57740 1085 57760 1205
rect 58490 1155 58510 1425
rect 58545 1155 58565 1425
rect 58600 1155 58620 1425
rect 58655 1155 58675 1425
rect 58710 1155 58730 1425
rect 58765 1155 58785 1425
rect 58820 1155 58840 1425
rect 58875 1155 58895 1425
rect 58930 1155 58950 1425
rect 58985 1155 59005 1425
rect 59040 1155 59060 1425
rect 59095 1155 59115 1425
rect 59150 1155 59170 1425
rect 59335 1130 59360 1155
rect 58490 1095 58510 1115
rect 59395 1130 59420 1155
rect 59455 1130 59480 1155
rect 59515 1130 59540 1155
rect 59150 1095 59170 1115
rect 56040 1025 56060 1045
rect 56740 1025 56760 1045
rect 57040 1025 57060 1045
rect 57740 1025 57760 1045
rect 55010 500 55030 520
rect 58770 500 58790 520
rect 56835 445 56855 465
rect 56945 445 56965 465
rect 54330 305 54355 330
rect 54390 305 54415 330
rect 54660 -345 54680 325
rect 54760 -345 54780 325
rect 54860 -345 54880 325
rect 54960 -345 54980 325
rect 55060 -345 55080 325
rect 55160 -345 55180 325
rect 55260 -345 55280 325
rect 56230 185 56250 405
rect 56285 185 56305 405
rect 56340 185 56360 405
rect 56395 185 56415 405
rect 56450 185 56470 405
rect 56505 185 56525 405
rect 56560 185 56580 405
rect 56615 185 56635 405
rect 56670 185 56690 405
rect 56725 185 56745 405
rect 56780 185 56800 405
rect 56835 185 56855 405
rect 56890 185 56910 405
rect 56945 185 56965 405
rect 57000 185 57020 405
rect 57055 185 57075 405
rect 57110 185 57130 405
rect 57165 185 57185 405
rect 57220 185 57240 405
rect 57275 185 57295 405
rect 57330 185 57350 405
rect 57385 185 57405 405
rect 57440 185 57460 405
rect 57495 185 57515 405
rect 56230 125 56250 145
rect 57495 125 57515 145
rect 57425 15 57445 35
rect 56605 -275 56625 -255
rect 56930 -275 56950 -255
rect 57050 -275 57070 -255
rect 57170 -275 57190 -255
rect 54660 -405 54680 -385
rect 55260 -405 55280 -385
rect 56440 -435 56460 -315
rect 56495 -435 56515 -315
rect 56550 -435 56570 -315
rect 56605 -435 56625 -315
rect 56660 -435 56680 -315
rect 56715 -435 56735 -315
rect 56770 -435 56790 -315
rect 56880 -435 56900 -315
rect 57220 -425 57240 -325
rect 58520 -345 58540 325
rect 58620 -345 58640 325
rect 58720 -345 58740 325
rect 58820 -345 58840 325
rect 58920 -345 58940 325
rect 59020 -345 59040 325
rect 59120 -345 59140 325
rect 59385 305 59410 330
rect 59445 305 59470 330
rect 58520 -405 58540 -385
rect 59120 -405 59140 -385
rect 56440 -495 56460 -475
rect 56770 -495 56790 -475
rect 56930 -495 56950 -475
rect 57050 -495 57070 -475
rect 57170 -495 57190 -475
<< metal1 >>
rect 52290 4320 52410 6110
rect 52290 4290 52295 4320
rect 52325 4290 52335 4320
rect 52365 4290 52375 4320
rect 52405 4290 52410 4320
rect 52290 4280 52410 4290
rect 52290 4250 52295 4280
rect 52325 4250 52335 4280
rect 52365 4250 52375 4280
rect 52405 4250 52410 4280
rect 52290 4240 52410 4250
rect 52290 4210 52295 4240
rect 52325 4210 52335 4240
rect 52365 4210 52375 4240
rect 52405 4210 52410 4240
rect 52290 4205 52410 4210
rect 52640 4320 52760 6110
rect 52640 4290 52645 4320
rect 52675 4290 52685 4320
rect 52715 4290 52725 4320
rect 52755 4290 52760 4320
rect 52640 4280 52760 4290
rect 52640 4250 52645 4280
rect 52675 4250 52685 4280
rect 52715 4250 52725 4280
rect 52755 4250 52760 4280
rect 52640 4240 52760 4250
rect 52640 4210 52645 4240
rect 52675 4210 52685 4240
rect 52715 4210 52725 4240
rect 52755 4210 52760 4240
rect 52640 4205 52760 4210
rect 52990 4320 53110 6110
rect 52990 4290 52995 4320
rect 53025 4290 53035 4320
rect 53065 4290 53075 4320
rect 53105 4290 53110 4320
rect 52990 4280 53110 4290
rect 52990 4250 52995 4280
rect 53025 4250 53035 4280
rect 53065 4250 53075 4280
rect 53105 4250 53110 4280
rect 52990 4240 53110 4250
rect 52990 4210 52995 4240
rect 53025 4210 53035 4240
rect 53065 4210 53075 4240
rect 53105 4210 53110 4240
rect 52990 4205 53110 4210
rect 53340 4320 53460 6110
rect 53340 4290 53345 4320
rect 53375 4290 53385 4320
rect 53415 4290 53425 4320
rect 53455 4290 53460 4320
rect 53340 4280 53460 4290
rect 53340 4250 53345 4280
rect 53375 4250 53385 4280
rect 53415 4250 53425 4280
rect 53455 4250 53460 4280
rect 53340 4240 53460 4250
rect 53340 4210 53345 4240
rect 53375 4210 53385 4240
rect 53415 4210 53425 4240
rect 53455 4210 53460 4240
rect 53340 4205 53460 4210
rect 54040 4320 54160 6110
rect 56205 5065 56245 5070
rect 56205 5035 56210 5065
rect 56240 5035 56245 5065
rect 56085 4930 56125 4935
rect 56085 4900 56090 4930
rect 56120 4900 56125 4930
rect 56085 4895 56125 4900
rect 56205 4930 56245 5035
rect 56675 5065 56715 5070
rect 56675 5035 56680 5065
rect 56710 5035 56715 5065
rect 56675 5030 56715 5035
rect 57085 5065 57125 5070
rect 57085 5035 57090 5065
rect 57120 5035 57125 5065
rect 57085 5030 57125 5035
rect 57555 5065 57595 5070
rect 57555 5035 57560 5065
rect 57590 5035 57595 5065
rect 56205 4900 56210 4930
rect 56240 4900 56245 4930
rect 56205 4895 56245 4900
rect 56265 4930 56305 4935
rect 56265 4900 56270 4930
rect 56300 4900 56305 4930
rect 56265 4895 56305 4900
rect 56090 4865 56120 4895
rect 56090 4545 56095 4865
rect 56115 4545 56120 4865
rect 56090 4535 56120 4545
rect 56150 4865 56180 4875
rect 56150 4545 56155 4865
rect 56175 4545 56180 4865
rect 56150 4485 56180 4545
rect 56210 4865 56240 4895
rect 56210 4545 56215 4865
rect 56235 4545 56240 4865
rect 56210 4530 56240 4545
rect 56270 4865 56300 4895
rect 56270 4545 56275 4865
rect 56295 4545 56300 4865
rect 56555 4840 56595 4845
rect 56555 4810 56560 4840
rect 56590 4810 56595 4840
rect 56555 4800 56595 4810
rect 56555 4770 56560 4800
rect 56590 4770 56595 4800
rect 56555 4760 56595 4770
rect 56555 4730 56560 4760
rect 56590 4730 56595 4760
rect 56555 4725 56595 4730
rect 56615 4840 56655 4845
rect 56615 4810 56620 4840
rect 56650 4810 56655 4840
rect 56615 4800 56655 4810
rect 56615 4770 56620 4800
rect 56650 4770 56655 4800
rect 56615 4760 56655 4770
rect 56615 4730 56620 4760
rect 56650 4730 56655 4760
rect 56615 4725 56655 4730
rect 56270 4535 56300 4545
rect 56560 4695 56590 4725
rect 56560 4545 56565 4695
rect 56585 4545 56590 4695
rect 56560 4535 56590 4545
rect 56620 4695 56650 4725
rect 56620 4545 56625 4695
rect 56645 4545 56650 4695
rect 56620 4535 56650 4545
rect 56680 4695 56710 5030
rect 56880 5010 56920 5015
rect 56880 4980 56885 5010
rect 56915 4980 56920 5010
rect 56880 4970 56920 4980
rect 56880 4940 56885 4970
rect 56915 4940 56920 4970
rect 56880 4930 56920 4940
rect 56880 4900 56885 4930
rect 56915 4900 56920 4930
rect 56735 4840 56775 4845
rect 56735 4810 56740 4840
rect 56770 4810 56775 4840
rect 56735 4800 56775 4810
rect 56735 4770 56740 4800
rect 56770 4770 56775 4800
rect 56735 4760 56775 4770
rect 56735 4730 56740 4760
rect 56770 4730 56775 4760
rect 56735 4725 56775 4730
rect 56880 4840 56920 4900
rect 57025 5010 57065 5015
rect 57025 4980 57030 5010
rect 57060 4980 57065 5010
rect 57025 4970 57065 4980
rect 57025 4940 57030 4970
rect 57060 4940 57065 4970
rect 57025 4930 57065 4940
rect 57025 4900 57030 4930
rect 57060 4900 57065 4930
rect 57025 4895 57065 4900
rect 56880 4810 56885 4840
rect 56915 4810 56920 4840
rect 56880 4800 56920 4810
rect 56880 4770 56885 4800
rect 56915 4770 56920 4800
rect 56880 4760 56920 4770
rect 56880 4730 56885 4760
rect 56915 4730 56920 4760
rect 56680 4545 56685 4695
rect 56705 4545 56710 4695
rect 56680 4530 56710 4545
rect 56740 4695 56770 4725
rect 56740 4545 56745 4695
rect 56765 4545 56770 4695
rect 56740 4535 56770 4545
rect 56205 4525 56245 4530
rect 56205 4495 56210 4525
rect 56240 4495 56245 4525
rect 56205 4490 56245 4495
rect 56675 4525 56715 4530
rect 56675 4495 56680 4525
rect 56710 4495 56715 4525
rect 56675 4490 56715 4495
rect 56150 4480 56190 4485
rect 56150 4450 56155 4480
rect 56185 4450 56190 4480
rect 56150 4445 56190 4450
rect 56630 4480 56660 4485
rect 56630 4445 56660 4450
rect 56825 4480 56865 4485
rect 56825 4450 56830 4480
rect 56860 4450 56865 4480
rect 56825 4445 56865 4450
rect 54040 4290 54045 4320
rect 54075 4290 54085 4320
rect 54115 4290 54125 4320
rect 54155 4290 54160 4320
rect 54040 4280 54160 4290
rect 54040 4250 54045 4280
rect 54075 4250 54085 4280
rect 54115 4250 54125 4280
rect 54155 4250 54160 4280
rect 54040 4240 54160 4250
rect 54040 4210 54045 4240
rect 54075 4210 54085 4240
rect 54115 4210 54125 4240
rect 54155 4210 54160 4240
rect 54040 4205 54160 4210
rect 54590 4320 54630 4325
rect 54590 4290 54595 4320
rect 54625 4290 54630 4320
rect 54590 4280 54630 4290
rect 54590 4250 54595 4280
rect 54625 4250 54630 4280
rect 54590 4240 54630 4250
rect 54590 4210 54595 4240
rect 54625 4210 54630 4240
rect 54590 4050 54630 4210
rect 54950 4320 54990 4325
rect 54950 4290 54955 4320
rect 54985 4290 54990 4320
rect 54950 4280 54990 4290
rect 54950 4250 54955 4280
rect 54985 4250 54990 4280
rect 54950 4240 54990 4250
rect 54950 4210 54955 4240
rect 54985 4210 54990 4240
rect 54650 4185 54930 4190
rect 54650 4155 54655 4185
rect 54685 4155 54695 4185
rect 54725 4155 54735 4185
rect 54765 4155 54775 4185
rect 54805 4155 54815 4185
rect 54845 4155 54855 4185
rect 54885 4155 54895 4185
rect 54925 4155 54930 4185
rect 54650 4145 54930 4155
rect 54650 4115 54655 4145
rect 54685 4115 54695 4145
rect 54725 4115 54735 4145
rect 54765 4115 54775 4145
rect 54805 4115 54815 4145
rect 54845 4115 54855 4145
rect 54885 4115 54895 4145
rect 54925 4115 54930 4145
rect 54650 4105 54930 4115
rect 54650 4075 54655 4105
rect 54685 4075 54695 4105
rect 54725 4075 54735 4105
rect 54765 4075 54775 4105
rect 54805 4075 54815 4105
rect 54845 4075 54855 4105
rect 54885 4075 54895 4105
rect 54925 4075 54930 4105
rect 54650 4070 54930 4075
rect 54590 4020 54595 4050
rect 54625 4020 54630 4050
rect 54590 4015 54630 4020
rect 54595 4000 54625 4015
rect 54595 3680 54600 4000
rect 54620 3680 54625 4000
rect 54595 3640 54625 3680
rect 54655 4000 54685 4070
rect 54710 4050 54750 4055
rect 54710 4020 54715 4050
rect 54745 4020 54750 4050
rect 54710 4015 54750 4020
rect 54655 3680 54660 4000
rect 54680 3680 54685 4000
rect 54655 3665 54685 3680
rect 54715 4000 54745 4015
rect 54715 3680 54720 4000
rect 54740 3680 54745 4000
rect 54715 3670 54745 3680
rect 54775 4000 54805 4070
rect 54830 4050 54870 4055
rect 54830 4020 54835 4050
rect 54865 4020 54870 4050
rect 54830 4015 54870 4020
rect 54775 3680 54780 4000
rect 54800 3680 54805 4000
rect 54775 3665 54805 3680
rect 54835 4000 54865 4015
rect 54835 3680 54840 4000
rect 54860 3680 54865 4000
rect 54835 3670 54865 3680
rect 54895 4000 54925 4070
rect 54950 4050 54990 4210
rect 55310 4320 55350 4325
rect 55310 4290 55315 4320
rect 55345 4290 55350 4320
rect 55310 4280 55350 4290
rect 55310 4250 55315 4280
rect 55345 4250 55350 4280
rect 55310 4240 55350 4250
rect 55310 4210 55315 4240
rect 55345 4210 55350 4240
rect 55010 4185 55290 4190
rect 55010 4155 55015 4185
rect 55045 4155 55055 4185
rect 55085 4155 55095 4185
rect 55125 4155 55135 4185
rect 55165 4155 55175 4185
rect 55205 4155 55215 4185
rect 55245 4155 55255 4185
rect 55285 4155 55290 4185
rect 55010 4145 55290 4155
rect 55010 4115 55015 4145
rect 55045 4115 55055 4145
rect 55085 4115 55095 4145
rect 55125 4115 55135 4145
rect 55165 4115 55175 4145
rect 55205 4115 55215 4145
rect 55245 4115 55255 4145
rect 55285 4115 55290 4145
rect 55010 4105 55290 4115
rect 55010 4075 55015 4105
rect 55045 4075 55055 4105
rect 55085 4075 55095 4105
rect 55125 4075 55135 4105
rect 55165 4075 55175 4105
rect 55205 4075 55215 4105
rect 55245 4075 55255 4105
rect 55285 4075 55290 4105
rect 55010 4070 55290 4075
rect 54950 4020 54955 4050
rect 54985 4020 54990 4050
rect 54950 4015 54990 4020
rect 54895 3680 54900 4000
rect 54920 3680 54925 4000
rect 54895 3665 54925 3680
rect 54955 4000 54985 4015
rect 54955 3680 54960 4000
rect 54980 3680 54985 4000
rect 54955 3670 54985 3680
rect 55015 4000 55045 4070
rect 55070 4050 55110 4055
rect 55070 4020 55075 4050
rect 55105 4020 55110 4050
rect 55070 4015 55110 4020
rect 55015 3680 55020 4000
rect 55040 3680 55045 4000
rect 55015 3665 55045 3680
rect 55075 4000 55105 4015
rect 55075 3680 55080 4000
rect 55100 3680 55105 4000
rect 55075 3670 55105 3680
rect 55135 4000 55165 4070
rect 55190 4050 55230 4055
rect 55190 4020 55195 4050
rect 55225 4020 55230 4050
rect 55190 4015 55230 4020
rect 55135 3680 55140 4000
rect 55160 3680 55165 4000
rect 55135 3665 55165 3680
rect 55195 4000 55225 4015
rect 55195 3680 55200 4000
rect 55220 3680 55225 4000
rect 55195 3670 55225 3680
rect 55255 4000 55285 4070
rect 55310 4050 55350 4210
rect 55310 4020 55315 4050
rect 55345 4020 55350 4050
rect 55310 4015 55350 4020
rect 55535 4320 55655 4325
rect 55535 4290 55540 4320
rect 55570 4290 55580 4320
rect 55610 4290 55620 4320
rect 55650 4290 55655 4320
rect 55535 4280 55655 4290
rect 55535 4250 55540 4280
rect 55570 4250 55580 4280
rect 55610 4250 55620 4280
rect 55650 4250 55655 4280
rect 55535 4240 55655 4250
rect 55535 4210 55540 4240
rect 55570 4210 55580 4240
rect 55610 4210 55620 4240
rect 55650 4210 55655 4240
rect 55255 3680 55260 4000
rect 55280 3680 55285 4000
rect 55255 3665 55285 3680
rect 55315 4000 55345 4015
rect 55315 3680 55320 4000
rect 55340 3680 55345 4000
rect 54595 3620 54600 3640
rect 54620 3620 54625 3640
rect 54650 3660 54690 3665
rect 54650 3630 54655 3660
rect 54685 3630 54690 3660
rect 54650 3625 54690 3630
rect 54770 3660 54810 3665
rect 54770 3630 54775 3660
rect 54805 3630 54810 3660
rect 54770 3625 54810 3630
rect 54890 3660 54930 3665
rect 54890 3630 54895 3660
rect 54925 3630 54930 3660
rect 54890 3625 54930 3630
rect 55010 3660 55050 3665
rect 55010 3630 55015 3660
rect 55045 3630 55050 3660
rect 55010 3625 55050 3630
rect 55130 3660 55170 3665
rect 55130 3630 55135 3660
rect 55165 3630 55170 3660
rect 55130 3625 55170 3630
rect 55250 3660 55290 3665
rect 55250 3630 55255 3660
rect 55285 3630 55290 3660
rect 55250 3625 55290 3630
rect 55315 3640 55345 3680
rect 54595 3610 54625 3620
rect 55315 3620 55320 3640
rect 55340 3620 55345 3640
rect 55315 3610 55345 3620
rect 54950 3535 54990 3540
rect 54950 3505 54955 3535
rect 54985 3505 54990 3535
rect 54950 3500 54990 3505
rect 55400 3490 55520 3495
rect 55400 3460 55405 3490
rect 55435 3460 55445 3490
rect 55475 3460 55485 3490
rect 55515 3460 55520 3490
rect 55400 3450 55520 3460
rect 55400 3420 55405 3450
rect 55435 3420 55445 3450
rect 55475 3420 55485 3450
rect 55515 3420 55520 3450
rect 55400 3410 55520 3420
rect 55400 3380 55405 3410
rect 55435 3380 55445 3410
rect 55475 3380 55485 3410
rect 55515 3380 55520 3410
rect 54255 3375 54295 3380
rect 54255 3345 54260 3375
rect 54290 3345 54295 3375
rect 54255 3200 54295 3345
rect 54620 3355 54660 3360
rect 54620 3325 54625 3355
rect 54655 3325 54660 3355
rect 54620 3315 54660 3325
rect 54620 3285 54625 3315
rect 54655 3285 54660 3315
rect 54620 3275 54660 3285
rect 54620 3245 54625 3275
rect 54655 3245 54660 3275
rect 54620 3240 54660 3245
rect 54730 3355 54770 3360
rect 54730 3325 54735 3355
rect 54765 3325 54770 3355
rect 54730 3315 54770 3325
rect 54730 3285 54735 3315
rect 54765 3285 54770 3315
rect 54730 3275 54770 3285
rect 54730 3245 54735 3275
rect 54765 3245 54770 3275
rect 54730 3240 54770 3245
rect 54840 3355 54880 3360
rect 54840 3325 54845 3355
rect 54875 3325 54880 3355
rect 54840 3315 54880 3325
rect 54840 3285 54845 3315
rect 54875 3285 54880 3315
rect 54840 3275 54880 3285
rect 54840 3245 54845 3275
rect 54875 3245 54880 3275
rect 54840 3240 54880 3245
rect 54950 3355 54990 3360
rect 54950 3325 54955 3355
rect 54985 3325 54990 3355
rect 54950 3315 54990 3325
rect 54950 3285 54955 3315
rect 54985 3285 54990 3315
rect 54950 3275 54990 3285
rect 54950 3245 54955 3275
rect 54985 3245 54990 3275
rect 54950 3240 54990 3245
rect 55060 3355 55100 3360
rect 55060 3325 55065 3355
rect 55095 3325 55100 3355
rect 55060 3315 55100 3325
rect 55060 3285 55065 3315
rect 55095 3285 55100 3315
rect 55060 3275 55100 3285
rect 55060 3245 55065 3275
rect 55095 3245 55100 3275
rect 55060 3240 55100 3245
rect 55170 3355 55210 3360
rect 55170 3325 55175 3355
rect 55205 3325 55210 3355
rect 55170 3315 55210 3325
rect 55170 3285 55175 3315
rect 55205 3285 55210 3315
rect 55170 3275 55210 3285
rect 55170 3245 55175 3275
rect 55205 3245 55210 3275
rect 55170 3240 55210 3245
rect 55280 3355 55320 3360
rect 55280 3325 55285 3355
rect 55315 3325 55320 3355
rect 55280 3315 55320 3325
rect 55280 3285 55285 3315
rect 55315 3285 55320 3315
rect 55280 3275 55320 3285
rect 55280 3245 55285 3275
rect 55315 3245 55320 3275
rect 55280 3240 55320 3245
rect 54625 3200 54655 3240
rect 54204 3190 54345 3200
rect 54204 3170 54210 3190
rect 54230 3170 54265 3190
rect 54285 3170 54320 3190
rect 54340 3170 54345 3190
rect 54204 3160 54345 3170
rect 54625 3180 54630 3200
rect 54650 3180 54655 3200
rect 54625 3140 54655 3180
rect 54675 3190 54715 3195
rect 54675 3160 54680 3190
rect 54710 3160 54715 3190
rect 54675 3155 54715 3160
rect 54204 2585 54345 2595
rect 54204 2565 54210 2585
rect 54230 2565 54265 2585
rect 54285 2565 54320 2585
rect 54340 2565 54345 2585
rect 54204 2555 54345 2565
rect 54625 2570 54630 3140
rect 54650 2570 54655 3140
rect 54625 2560 54655 2570
rect 54680 3140 54710 3155
rect 54680 2570 54685 3140
rect 54705 2570 54710 3140
rect 54680 2555 54710 2570
rect 54735 3140 54765 3240
rect 54785 3190 54825 3195
rect 54785 3160 54790 3190
rect 54820 3160 54825 3190
rect 54785 3155 54825 3160
rect 54735 2570 54740 3140
rect 54760 2570 54765 3140
rect 54735 2560 54765 2570
rect 54790 3140 54820 3155
rect 54790 2570 54795 3140
rect 54815 2570 54820 3140
rect 54790 2555 54820 2570
rect 54845 3140 54875 3240
rect 54895 3190 54935 3195
rect 54895 3160 54900 3190
rect 54930 3160 54935 3190
rect 54895 3155 54935 3160
rect 54845 2570 54850 3140
rect 54870 2570 54875 3140
rect 54845 2560 54875 2570
rect 54900 3140 54930 3155
rect 54900 2570 54905 3140
rect 54925 2570 54930 3140
rect 54900 2555 54930 2570
rect 54955 3140 54985 3240
rect 55005 3190 55045 3195
rect 55005 3160 55010 3190
rect 55040 3160 55045 3190
rect 55005 3155 55045 3160
rect 54955 2570 54960 3140
rect 54980 2570 54985 3140
rect 54955 2560 54985 2570
rect 55010 3140 55040 3155
rect 55010 2570 55015 3140
rect 55035 2570 55040 3140
rect 55010 2555 55040 2570
rect 55065 3140 55095 3240
rect 55115 3190 55155 3195
rect 55115 3160 55120 3190
rect 55150 3160 55155 3190
rect 55115 3155 55155 3160
rect 55065 2570 55070 3140
rect 55090 2570 55095 3140
rect 55065 2560 55095 2570
rect 55120 3140 55150 3155
rect 55120 2570 55125 3140
rect 55145 2570 55150 3140
rect 55120 2555 55150 2570
rect 55175 3140 55205 3240
rect 55285 3200 55315 3240
rect 55225 3190 55265 3195
rect 55225 3160 55230 3190
rect 55260 3160 55265 3190
rect 55225 3155 55265 3160
rect 55285 3180 55290 3200
rect 55310 3180 55315 3200
rect 55175 2570 55180 3140
rect 55200 2570 55205 3140
rect 55175 2560 55205 2570
rect 55230 3140 55260 3155
rect 55230 2570 55235 3140
rect 55255 2570 55260 3140
rect 55230 2555 55260 2570
rect 55285 3140 55315 3180
rect 55285 2570 55290 3140
rect 55310 2570 55315 3140
rect 55285 2560 55315 2570
rect 54215 2470 54335 2555
rect 54215 2440 54220 2470
rect 54250 2440 54260 2470
rect 54290 2440 54300 2470
rect 54330 2440 54335 2470
rect 54215 2430 54335 2440
rect 54215 2400 54220 2430
rect 54250 2400 54260 2430
rect 54290 2400 54300 2430
rect 54330 2400 54335 2430
rect 54215 2390 54335 2400
rect 54215 2360 54220 2390
rect 54250 2360 54260 2390
rect 54290 2360 54300 2390
rect 54330 2360 54335 2390
rect 54215 2355 54335 2360
rect 54675 2550 54715 2555
rect 54675 2520 54680 2550
rect 54710 2520 54715 2550
rect 54675 2325 54715 2520
rect 54785 2550 54825 2555
rect 54785 2520 54790 2550
rect 54820 2520 54825 2550
rect 54785 2325 54825 2520
rect 54895 2550 54935 2555
rect 54895 2520 54900 2550
rect 54930 2520 54935 2550
rect 54895 2325 54935 2520
rect 55005 2550 55045 2555
rect 55005 2520 55010 2550
rect 55040 2520 55045 2550
rect 54950 2470 54990 2475
rect 54950 2440 54955 2470
rect 54985 2440 54990 2470
rect 54950 2430 54990 2440
rect 54950 2400 54955 2430
rect 54985 2400 54990 2430
rect 54950 2390 54990 2400
rect 54950 2360 54955 2390
rect 54985 2360 54990 2390
rect 54950 2355 54990 2360
rect 55005 2325 55045 2520
rect 55115 2550 55155 2555
rect 55115 2520 55120 2550
rect 55150 2520 55155 2550
rect 55115 2325 55155 2520
rect 55225 2550 55265 2555
rect 55225 2520 55230 2550
rect 55260 2520 55265 2550
rect 55225 2325 55265 2520
rect 53990 2320 54240 2325
rect 53990 2290 53995 2320
rect 54025 2290 54035 2320
rect 54065 2290 54080 2320
rect 54110 2290 54120 2320
rect 54150 2290 54165 2320
rect 54195 2290 54205 2320
rect 54235 2290 54240 2320
rect 53990 2280 54240 2290
rect 53990 2250 53995 2280
rect 54025 2250 54035 2280
rect 54065 2250 54080 2280
rect 54110 2250 54120 2280
rect 54150 2250 54165 2280
rect 54195 2250 54205 2280
rect 54235 2250 54240 2280
rect 53990 2240 54240 2250
rect 53990 2210 53995 2240
rect 54025 2210 54035 2240
rect 54065 2210 54080 2240
rect 54110 2210 54120 2240
rect 54150 2210 54165 2240
rect 54195 2210 54205 2240
rect 54235 2210 54240 2240
rect 53840 2050 53960 2055
rect 53840 2020 53845 2050
rect 53875 2020 53885 2050
rect 53915 2020 53925 2050
rect 53955 2020 53960 2050
rect 53840 2010 53960 2020
rect 53840 1980 53845 2010
rect 53875 1980 53885 2010
rect 53915 1980 53925 2010
rect 53955 1980 53960 2010
rect 53840 1970 53960 1980
rect 53840 1940 53845 1970
rect 53875 1940 53885 1970
rect 53915 1940 53925 1970
rect 53955 1940 53960 1970
rect 53840 940 53960 1940
rect 53840 910 53845 940
rect 53875 910 53885 940
rect 53915 910 53925 940
rect 53955 910 53960 940
rect 53840 900 53960 910
rect 53840 870 53845 900
rect 53875 870 53885 900
rect 53915 870 53925 900
rect 53955 870 53960 900
rect 53840 860 53960 870
rect 53840 830 53845 860
rect 53875 830 53885 860
rect 53915 830 53925 860
rect 53955 830 53960 860
rect 52290 -580 52410 -575
rect 52290 -610 52295 -580
rect 52325 -610 52335 -580
rect 52365 -610 52375 -580
rect 52405 -610 52410 -580
rect 52290 -620 52410 -610
rect 52290 -650 52295 -620
rect 52325 -650 52335 -620
rect 52365 -650 52375 -620
rect 52405 -650 52410 -620
rect 52290 -660 52410 -650
rect 52290 -690 52295 -660
rect 52325 -690 52335 -660
rect 52365 -690 52375 -660
rect 52405 -690 52410 -660
rect 52290 -1500 52410 -690
rect 52640 -580 52760 -575
rect 52640 -610 52645 -580
rect 52675 -610 52685 -580
rect 52715 -610 52725 -580
rect 52755 -610 52760 -580
rect 52640 -620 52760 -610
rect 52640 -650 52645 -620
rect 52675 -650 52685 -620
rect 52715 -650 52725 -620
rect 52755 -650 52760 -620
rect 52640 -660 52760 -650
rect 52640 -690 52645 -660
rect 52675 -690 52685 -660
rect 52715 -690 52725 -660
rect 52755 -690 52760 -660
rect 52640 -1500 52760 -690
rect 52990 -580 53110 -575
rect 52990 -610 52995 -580
rect 53025 -610 53035 -580
rect 53065 -610 53075 -580
rect 53105 -610 53110 -580
rect 52990 -620 53110 -610
rect 52990 -650 52995 -620
rect 53025 -650 53035 -620
rect 53065 -650 53075 -620
rect 53105 -650 53110 -620
rect 52990 -660 53110 -650
rect 52990 -690 52995 -660
rect 53025 -690 53035 -660
rect 53065 -690 53075 -660
rect 53105 -690 53110 -660
rect 52990 -1500 53110 -690
rect 53340 -580 53460 -575
rect 53340 -610 53345 -580
rect 53375 -610 53385 -580
rect 53415 -610 53425 -580
rect 53455 -610 53460 -580
rect 53340 -620 53460 -610
rect 53340 -650 53345 -620
rect 53375 -650 53385 -620
rect 53415 -650 53425 -620
rect 53455 -650 53460 -620
rect 53340 -660 53460 -650
rect 53340 -690 53345 -660
rect 53375 -690 53385 -660
rect 53415 -690 53425 -660
rect 53455 -690 53460 -660
rect 53340 -1500 53460 -690
rect 53690 -580 53810 -575
rect 53690 -610 53695 -580
rect 53725 -610 53735 -580
rect 53765 -610 53775 -580
rect 53805 -610 53810 -580
rect 53690 -620 53810 -610
rect 53690 -650 53695 -620
rect 53725 -650 53735 -620
rect 53765 -650 53775 -620
rect 53805 -650 53810 -620
rect 53690 -660 53810 -650
rect 53690 -690 53695 -660
rect 53725 -690 53735 -660
rect 53765 -690 53775 -660
rect 53805 -690 53810 -660
rect 53690 -1500 53810 -690
rect 53840 -580 53960 830
rect 53990 1710 54240 2210
rect 54675 2320 55265 2325
rect 54675 2290 54680 2320
rect 54710 2290 54735 2320
rect 54765 2290 54790 2320
rect 54820 2290 54845 2320
rect 54875 2290 54900 2320
rect 54930 2290 54955 2320
rect 54985 2290 55010 2320
rect 55040 2290 55065 2320
rect 55095 2290 55120 2320
rect 55150 2290 55175 2320
rect 55205 2290 55230 2320
rect 55260 2290 55265 2320
rect 54675 2280 55265 2290
rect 54675 2250 54680 2280
rect 54710 2250 54735 2280
rect 54765 2250 54790 2280
rect 54820 2250 54845 2280
rect 54875 2250 54900 2280
rect 54930 2250 54955 2280
rect 54985 2250 55010 2280
rect 55040 2250 55065 2280
rect 55095 2250 55120 2280
rect 55150 2250 55175 2280
rect 55205 2250 55230 2280
rect 55260 2250 55265 2280
rect 54675 2240 55265 2250
rect 54675 2210 54680 2240
rect 54710 2210 54735 2240
rect 54765 2210 54790 2240
rect 54820 2210 54845 2240
rect 54875 2210 54900 2240
rect 54930 2210 54955 2240
rect 54985 2210 55010 2240
rect 55040 2210 55065 2240
rect 55095 2210 55120 2240
rect 55150 2210 55175 2240
rect 55205 2210 55230 2240
rect 55260 2210 55265 2240
rect 54675 2205 55265 2210
rect 55400 2470 55520 3380
rect 55400 2440 55405 2470
rect 55435 2440 55445 2470
rect 55475 2440 55485 2470
rect 55515 2440 55520 2470
rect 55400 2430 55520 2440
rect 55400 2400 55405 2430
rect 55435 2400 55445 2430
rect 55475 2400 55485 2430
rect 55515 2400 55520 2430
rect 55400 2390 55520 2400
rect 55400 2360 55405 2390
rect 55435 2360 55445 2390
rect 55475 2360 55485 2390
rect 55515 2360 55520 2390
rect 54620 2185 54660 2190
rect 54620 2155 54625 2185
rect 54655 2155 54660 2185
rect 54620 2145 54660 2155
rect 54620 2115 54625 2145
rect 54655 2115 54660 2145
rect 54620 2105 54660 2115
rect 54620 2075 54625 2105
rect 54655 2075 54660 2105
rect 54620 2070 54660 2075
rect 55280 2185 55320 2190
rect 55280 2155 55285 2185
rect 55315 2155 55320 2185
rect 55280 2145 55320 2155
rect 55280 2115 55285 2145
rect 55315 2115 55320 2145
rect 55280 2105 55320 2115
rect 55280 2075 55285 2105
rect 55315 2075 55320 2105
rect 55280 2070 55320 2075
rect 53990 1680 54000 1710
rect 54030 1680 54050 1710
rect 54080 1680 54100 1710
rect 54130 1680 54150 1710
rect 54180 1680 54200 1710
rect 54230 1680 54240 1710
rect 54625 1925 54655 2070
rect 54675 2050 54715 2055
rect 54675 2020 54680 2050
rect 54710 2020 54715 2050
rect 54675 2010 54715 2020
rect 54675 1980 54680 2010
rect 54710 1980 54715 2010
rect 54675 1970 54715 1980
rect 54675 1940 54680 1970
rect 54710 1940 54715 1970
rect 54675 1935 54715 1940
rect 54785 2050 54825 2055
rect 54785 2020 54790 2050
rect 54820 2020 54825 2050
rect 54785 2010 54825 2020
rect 54785 1980 54790 2010
rect 54820 1980 54825 2010
rect 54785 1970 54825 1980
rect 54785 1940 54790 1970
rect 54820 1940 54825 1970
rect 54785 1935 54825 1940
rect 54895 2050 54935 2055
rect 54895 2020 54900 2050
rect 54930 2020 54935 2050
rect 54895 2010 54935 2020
rect 54895 1980 54900 2010
rect 54930 1980 54935 2010
rect 54895 1970 54935 1980
rect 54895 1940 54900 1970
rect 54930 1940 54935 1970
rect 54895 1935 54935 1940
rect 55005 2050 55045 2055
rect 55005 2020 55010 2050
rect 55040 2020 55045 2050
rect 55005 2010 55045 2020
rect 55005 1980 55010 2010
rect 55040 1980 55045 2010
rect 55005 1970 55045 1980
rect 55005 1940 55010 1970
rect 55040 1940 55045 1970
rect 55005 1935 55045 1940
rect 55115 2050 55155 2055
rect 55115 2020 55120 2050
rect 55150 2020 55155 2050
rect 55115 2010 55155 2020
rect 55115 1980 55120 2010
rect 55150 1980 55155 2010
rect 55115 1970 55155 1980
rect 55115 1940 55120 1970
rect 55150 1940 55155 1970
rect 55115 1935 55155 1940
rect 55225 2050 55265 2055
rect 55225 2020 55230 2050
rect 55260 2020 55265 2050
rect 55225 2010 55265 2020
rect 55225 1980 55230 2010
rect 55260 1980 55265 2010
rect 55225 1970 55265 1980
rect 55225 1940 55230 1970
rect 55260 1940 55265 1970
rect 55225 1935 55265 1940
rect 54625 1905 54630 1925
rect 54650 1905 54655 1925
rect 54625 1865 54655 1905
rect 54625 1695 54630 1865
rect 54650 1695 54655 1865
rect 54625 1685 54655 1695
rect 54680 1865 54710 1935
rect 54730 1915 54770 1920
rect 54730 1885 54735 1915
rect 54765 1885 54770 1915
rect 54730 1880 54770 1885
rect 54680 1695 54685 1865
rect 54705 1695 54710 1865
rect 54680 1685 54710 1695
rect 54735 1865 54765 1880
rect 54735 1695 54740 1865
rect 54760 1695 54765 1865
rect 53990 1660 54240 1680
rect 54735 1665 54765 1695
rect 54790 1865 54820 1935
rect 54840 1915 54880 1920
rect 54840 1885 54845 1915
rect 54875 1885 54880 1915
rect 54840 1880 54880 1885
rect 54790 1695 54795 1865
rect 54815 1695 54820 1865
rect 54790 1685 54820 1695
rect 54845 1865 54875 1880
rect 54845 1695 54850 1865
rect 54870 1695 54875 1865
rect 54845 1665 54875 1695
rect 54900 1865 54930 1935
rect 54950 1915 54990 1920
rect 54950 1885 54955 1915
rect 54985 1885 54990 1915
rect 54950 1880 54990 1885
rect 54900 1695 54905 1865
rect 54925 1695 54930 1865
rect 54900 1685 54930 1695
rect 54955 1865 54985 1880
rect 54955 1695 54960 1865
rect 54980 1695 54985 1865
rect 54955 1665 54985 1695
rect 55010 1865 55040 1935
rect 55060 1915 55100 1920
rect 55060 1885 55065 1915
rect 55095 1885 55100 1915
rect 55060 1880 55100 1885
rect 55010 1695 55015 1865
rect 55035 1695 55040 1865
rect 55010 1685 55040 1695
rect 55065 1865 55095 1880
rect 55065 1695 55070 1865
rect 55090 1695 55095 1865
rect 55065 1665 55095 1695
rect 55120 1865 55150 1935
rect 55170 1915 55210 1920
rect 55170 1885 55175 1915
rect 55205 1885 55210 1915
rect 55170 1880 55210 1885
rect 55120 1695 55125 1865
rect 55145 1695 55150 1865
rect 55120 1685 55150 1695
rect 55175 1865 55205 1880
rect 55175 1695 55180 1865
rect 55200 1695 55205 1865
rect 55175 1665 55205 1695
rect 55230 1865 55260 1935
rect 55230 1695 55235 1865
rect 55255 1695 55260 1865
rect 55230 1685 55260 1695
rect 55285 1925 55315 2070
rect 55285 1905 55290 1925
rect 55310 1905 55315 1925
rect 55285 1865 55315 1905
rect 55285 1695 55290 1865
rect 55310 1695 55315 1865
rect 55285 1685 55315 1695
rect 53990 1630 54000 1660
rect 54030 1630 54050 1660
rect 54080 1630 54100 1660
rect 54130 1630 54150 1660
rect 54180 1630 54200 1660
rect 54230 1630 54240 1660
rect 53990 1610 54240 1630
rect 54485 1660 54525 1665
rect 54485 1630 54490 1660
rect 54520 1630 54525 1660
rect 54485 1625 54525 1630
rect 54730 1660 54770 1665
rect 54730 1630 54735 1660
rect 54765 1630 54770 1660
rect 54730 1625 54770 1630
rect 54840 1660 54880 1665
rect 54840 1630 54845 1660
rect 54875 1630 54880 1660
rect 54840 1625 54880 1630
rect 54950 1660 54990 1665
rect 54950 1630 54955 1660
rect 54985 1630 54990 1660
rect 54950 1625 54990 1630
rect 55060 1660 55100 1665
rect 55060 1630 55065 1660
rect 55095 1630 55100 1660
rect 55060 1625 55100 1630
rect 55170 1660 55210 1665
rect 55170 1630 55175 1660
rect 55205 1630 55210 1660
rect 55170 1625 55210 1630
rect 53990 1580 54000 1610
rect 54030 1580 54050 1610
rect 54080 1580 54100 1610
rect 54130 1580 54150 1610
rect 54180 1580 54200 1610
rect 54230 1580 54240 1610
rect 53990 470 54240 1580
rect 54255 1160 54290 1166
rect 54255 1120 54290 1125
rect 54315 1160 54350 1165
rect 54315 1120 54350 1125
rect 54375 1160 54410 1165
rect 54375 1120 54410 1125
rect 54435 1160 54470 1165
rect 54435 1120 54470 1125
rect 54265 810 54285 1120
rect 54385 1090 54405 1120
rect 54495 1090 54515 1625
rect 55115 1595 55155 1600
rect 55115 1565 55120 1595
rect 55150 1565 55155 1595
rect 55115 1555 55155 1565
rect 55115 1525 55120 1555
rect 55150 1525 55155 1555
rect 55115 1520 55155 1525
rect 55400 1595 55520 2360
rect 55400 1565 55405 1595
rect 55435 1565 55445 1595
rect 55475 1565 55485 1595
rect 55515 1565 55520 1595
rect 55400 1555 55520 1565
rect 55400 1525 55405 1555
rect 55435 1525 55445 1555
rect 55475 1525 55485 1555
rect 55515 1525 55520 1555
rect 55400 1520 55520 1525
rect 55535 3355 55655 4210
rect 56005 4185 56765 4190
rect 56005 4155 56010 4185
rect 56040 4155 56050 4185
rect 56080 4155 56090 4185
rect 56120 4155 56130 4185
rect 56160 4155 56170 4185
rect 56200 4155 56210 4185
rect 56240 4155 56250 4185
rect 56280 4155 56290 4185
rect 56320 4155 56330 4185
rect 56360 4155 56370 4185
rect 56400 4155 56410 4185
rect 56440 4155 56450 4185
rect 56480 4155 56490 4185
rect 56520 4155 56530 4185
rect 56560 4155 56570 4185
rect 56600 4155 56610 4185
rect 56640 4155 56650 4185
rect 56680 4155 56690 4185
rect 56720 4155 56730 4185
rect 56760 4155 56765 4185
rect 56005 4145 56765 4155
rect 56005 4115 56010 4145
rect 56040 4115 56050 4145
rect 56080 4115 56090 4145
rect 56120 4115 56130 4145
rect 56160 4115 56170 4145
rect 56200 4115 56210 4145
rect 56240 4115 56250 4145
rect 56280 4115 56290 4145
rect 56320 4115 56330 4145
rect 56360 4115 56370 4145
rect 56400 4115 56410 4145
rect 56440 4115 56450 4145
rect 56480 4115 56490 4145
rect 56520 4115 56530 4145
rect 56560 4115 56570 4145
rect 56600 4115 56610 4145
rect 56640 4115 56650 4145
rect 56680 4115 56690 4145
rect 56720 4115 56730 4145
rect 56760 4115 56765 4145
rect 56005 4105 56765 4115
rect 56005 4075 56010 4105
rect 56040 4075 56050 4105
rect 56080 4075 56090 4105
rect 56120 4075 56130 4105
rect 56160 4075 56170 4105
rect 56200 4075 56210 4105
rect 56240 4075 56250 4105
rect 56280 4075 56290 4105
rect 56320 4075 56330 4105
rect 56360 4075 56370 4105
rect 56400 4075 56410 4105
rect 56440 4075 56450 4105
rect 56480 4075 56490 4105
rect 56520 4075 56530 4105
rect 56560 4075 56570 4105
rect 56600 4075 56610 4105
rect 56640 4075 56650 4105
rect 56680 4075 56690 4105
rect 56720 4075 56730 4105
rect 56760 4075 56765 4105
rect 56005 4070 56765 4075
rect 56010 4000 56040 4070
rect 56065 4050 56105 4055
rect 56065 4020 56070 4050
rect 56100 4020 56105 4050
rect 56065 4015 56105 4020
rect 56010 3680 56015 4000
rect 56035 3680 56040 4000
rect 56010 3640 56040 3680
rect 56070 4000 56100 4015
rect 56070 3680 56075 4000
rect 56095 3680 56100 4000
rect 56070 3665 56100 3680
rect 56130 4000 56160 4070
rect 56185 4050 56225 4055
rect 56185 4020 56190 4050
rect 56220 4020 56225 4050
rect 56185 4015 56225 4020
rect 56130 3680 56135 4000
rect 56155 3680 56160 4000
rect 56130 3670 56160 3680
rect 56190 4000 56220 4015
rect 56190 3680 56195 4000
rect 56215 3680 56220 4000
rect 56190 3665 56220 3680
rect 56250 4000 56280 4070
rect 56305 4050 56345 4055
rect 56305 4020 56310 4050
rect 56340 4020 56345 4050
rect 56305 4015 56345 4020
rect 56250 3680 56255 4000
rect 56275 3680 56280 4000
rect 56250 3670 56280 3680
rect 56310 4000 56340 4015
rect 56310 3680 56315 4000
rect 56335 3680 56340 4000
rect 56310 3665 56340 3680
rect 56370 4000 56400 4070
rect 56425 4050 56465 4055
rect 56425 4020 56430 4050
rect 56460 4020 56465 4050
rect 56425 4015 56465 4020
rect 56370 3680 56375 4000
rect 56395 3680 56400 4000
rect 56370 3670 56400 3680
rect 56430 4000 56460 4015
rect 56430 3680 56435 4000
rect 56455 3680 56460 4000
rect 56430 3665 56460 3680
rect 56490 4000 56520 4070
rect 56545 4050 56585 4055
rect 56545 4020 56550 4050
rect 56580 4020 56585 4050
rect 56545 4015 56585 4020
rect 56490 3680 56495 4000
rect 56515 3680 56520 4000
rect 56490 3670 56520 3680
rect 56550 4000 56580 4015
rect 56550 3680 56555 4000
rect 56575 3680 56580 4000
rect 56550 3665 56580 3680
rect 56610 4000 56640 4070
rect 56665 4050 56705 4055
rect 56665 4020 56670 4050
rect 56700 4020 56705 4050
rect 56665 4015 56705 4020
rect 56610 3680 56615 4000
rect 56635 3680 56640 4000
rect 56610 3670 56640 3680
rect 56670 4000 56700 4015
rect 56670 3680 56675 4000
rect 56695 3680 56700 4000
rect 56670 3665 56700 3680
rect 56730 4000 56760 4070
rect 56730 3680 56735 4000
rect 56755 3680 56760 4000
rect 56010 3620 56015 3640
rect 56035 3620 56040 3640
rect 56010 3610 56040 3620
rect 56065 3660 56105 3665
rect 56065 3630 56070 3660
rect 56100 3630 56105 3660
rect 56065 3495 56105 3630
rect 56185 3660 56225 3665
rect 56185 3630 56190 3660
rect 56220 3630 56225 3660
rect 56185 3495 56225 3630
rect 56305 3660 56345 3665
rect 56305 3630 56310 3660
rect 56340 3630 56345 3660
rect 56305 3495 56345 3630
rect 56425 3660 56465 3665
rect 56425 3630 56430 3660
rect 56460 3630 56465 3660
rect 56365 3580 56405 3585
rect 56365 3550 56370 3580
rect 56400 3550 56405 3580
rect 56365 3545 56405 3550
rect 56425 3495 56465 3630
rect 56545 3660 56585 3665
rect 56545 3630 56550 3660
rect 56580 3630 56585 3660
rect 56545 3495 56585 3630
rect 56665 3660 56705 3665
rect 56665 3630 56670 3660
rect 56700 3630 56705 3660
rect 56665 3495 56705 3630
rect 56730 3640 56760 3680
rect 56730 3620 56735 3640
rect 56755 3620 56760 3640
rect 56730 3610 56760 3620
rect 56845 3585 56865 4445
rect 56880 4320 56920 4730
rect 57030 4865 57060 4895
rect 57030 4545 57035 4865
rect 57055 4545 57060 4865
rect 57030 4535 57060 4545
rect 57090 4865 57120 5030
rect 57145 5010 57185 5015
rect 57145 4980 57150 5010
rect 57180 4980 57185 5010
rect 57145 4970 57185 4980
rect 57145 4940 57150 4970
rect 57180 4940 57185 4970
rect 57145 4930 57185 4940
rect 57145 4900 57150 4930
rect 57180 4900 57185 4930
rect 57145 4895 57185 4900
rect 57205 5010 57245 5015
rect 57205 4980 57210 5010
rect 57240 4980 57245 5010
rect 57205 4970 57245 4980
rect 57205 4940 57210 4970
rect 57240 4940 57245 4970
rect 57205 4930 57245 4940
rect 57205 4900 57210 4930
rect 57240 4900 57245 4930
rect 57205 4895 57245 4900
rect 57495 4930 57535 4935
rect 57495 4900 57500 4930
rect 57530 4900 57535 4930
rect 57495 4895 57535 4900
rect 57555 4930 57595 5035
rect 57555 4900 57560 4930
rect 57590 4900 57595 4930
rect 57555 4895 57595 4900
rect 57675 4930 57715 4935
rect 57675 4900 57680 4930
rect 57710 4900 57715 4930
rect 57675 4895 57715 4900
rect 57090 4545 57095 4865
rect 57115 4545 57120 4865
rect 57090 4530 57120 4545
rect 57150 4865 57180 4895
rect 57150 4545 57155 4865
rect 57175 4545 57180 4865
rect 57150 4535 57180 4545
rect 57210 4865 57240 4895
rect 57210 4545 57215 4865
rect 57235 4545 57240 4865
rect 57210 4535 57240 4545
rect 57500 4865 57530 4895
rect 57500 4545 57505 4865
rect 57525 4545 57530 4865
rect 57500 4535 57530 4545
rect 57560 4865 57590 4895
rect 57560 4545 57565 4865
rect 57585 4545 57590 4865
rect 57560 4530 57590 4545
rect 57620 4865 57650 4875
rect 57620 4545 57625 4865
rect 57645 4545 57650 4865
rect 57085 4525 57125 4530
rect 57085 4495 57090 4525
rect 57120 4495 57125 4525
rect 57085 4490 57125 4495
rect 57555 4525 57595 4530
rect 57555 4495 57560 4525
rect 57590 4495 57595 4525
rect 57555 4490 57595 4495
rect 57140 4475 57170 4485
rect 57140 4455 57145 4475
rect 57165 4455 57170 4475
rect 56880 4290 56885 4320
rect 56915 4290 56920 4320
rect 56880 4280 56920 4290
rect 56880 4250 56885 4280
rect 56915 4250 56920 4280
rect 56880 4240 56920 4250
rect 56880 4210 56885 4240
rect 56915 4210 56920 4240
rect 56880 4205 56920 4210
rect 56935 4425 56975 4430
rect 56935 4395 56940 4425
rect 56970 4395 56975 4425
rect 57140 4420 57170 4455
rect 57576 4470 57606 4475
rect 57576 4435 57606 4440
rect 57620 4420 57650 4545
rect 57680 4865 57710 4895
rect 57680 4545 57685 4865
rect 57705 4545 57710 4865
rect 57680 4535 57710 4545
rect 56935 4390 56975 4395
rect 57135 4415 57175 4420
rect 56835 3580 56875 3585
rect 56835 3550 56840 3580
rect 56870 3550 56875 3580
rect 56835 3545 56875 3550
rect 56935 3540 56955 4390
rect 57135 4385 57140 4415
rect 57170 4385 57175 4415
rect 57135 4380 57175 4385
rect 57615 4415 57655 4420
rect 57615 4385 57620 4415
rect 57650 4385 57655 4415
rect 57615 4380 57655 4385
rect 58145 4320 58265 4325
rect 58145 4290 58150 4320
rect 58180 4290 58190 4320
rect 58220 4290 58230 4320
rect 58260 4290 58265 4320
rect 58145 4280 58265 4290
rect 58145 4250 58150 4280
rect 58180 4250 58190 4280
rect 58220 4250 58230 4280
rect 58260 4250 58265 4280
rect 58145 4240 58265 4250
rect 58145 4210 58150 4240
rect 58180 4210 58190 4240
rect 58220 4210 58230 4240
rect 58260 4210 58265 4240
rect 57035 4185 57795 4190
rect 57035 4155 57040 4185
rect 57070 4155 57080 4185
rect 57110 4155 57120 4185
rect 57150 4155 57160 4185
rect 57190 4155 57200 4185
rect 57230 4155 57240 4185
rect 57270 4155 57280 4185
rect 57310 4155 57320 4185
rect 57350 4155 57360 4185
rect 57390 4155 57400 4185
rect 57430 4155 57440 4185
rect 57470 4155 57480 4185
rect 57510 4155 57520 4185
rect 57550 4155 57560 4185
rect 57590 4155 57600 4185
rect 57630 4155 57640 4185
rect 57670 4155 57680 4185
rect 57710 4155 57720 4185
rect 57750 4155 57760 4185
rect 57790 4155 57795 4185
rect 57035 4145 57795 4155
rect 57035 4115 57040 4145
rect 57070 4115 57080 4145
rect 57110 4115 57120 4145
rect 57150 4115 57160 4145
rect 57190 4115 57200 4145
rect 57230 4115 57240 4145
rect 57270 4115 57280 4145
rect 57310 4115 57320 4145
rect 57350 4115 57360 4145
rect 57390 4115 57400 4145
rect 57430 4115 57440 4145
rect 57470 4115 57480 4145
rect 57510 4115 57520 4145
rect 57550 4115 57560 4145
rect 57590 4115 57600 4145
rect 57630 4115 57640 4145
rect 57670 4115 57680 4145
rect 57710 4115 57720 4145
rect 57750 4115 57760 4145
rect 57790 4115 57795 4145
rect 57035 4105 57795 4115
rect 57035 4075 57040 4105
rect 57070 4075 57080 4105
rect 57110 4075 57120 4105
rect 57150 4075 57160 4105
rect 57190 4075 57200 4105
rect 57230 4075 57240 4105
rect 57270 4075 57280 4105
rect 57310 4075 57320 4105
rect 57350 4075 57360 4105
rect 57390 4075 57400 4105
rect 57430 4075 57440 4105
rect 57470 4075 57480 4105
rect 57510 4075 57520 4105
rect 57550 4075 57560 4105
rect 57590 4075 57600 4105
rect 57630 4075 57640 4105
rect 57670 4075 57680 4105
rect 57710 4075 57720 4105
rect 57750 4075 57760 4105
rect 57790 4075 57795 4105
rect 57035 4070 57795 4075
rect 57040 4000 57070 4070
rect 57095 4050 57135 4055
rect 57095 4020 57100 4050
rect 57130 4020 57135 4050
rect 57095 4015 57135 4020
rect 57040 3680 57045 4000
rect 57065 3680 57070 4000
rect 57040 3640 57070 3680
rect 57100 4000 57130 4015
rect 57100 3680 57105 4000
rect 57125 3680 57130 4000
rect 57100 3665 57130 3680
rect 57160 4000 57190 4070
rect 57215 4050 57255 4055
rect 57215 4020 57220 4050
rect 57250 4020 57255 4050
rect 57215 4015 57255 4020
rect 57160 3680 57165 4000
rect 57185 3680 57190 4000
rect 57160 3670 57190 3680
rect 57220 4000 57250 4015
rect 57220 3680 57225 4000
rect 57245 3680 57250 4000
rect 57220 3665 57250 3680
rect 57280 4000 57310 4070
rect 57335 4050 57375 4055
rect 57335 4020 57340 4050
rect 57370 4020 57375 4050
rect 57335 4015 57375 4020
rect 57280 3680 57285 4000
rect 57305 3680 57310 4000
rect 57280 3670 57310 3680
rect 57340 4000 57370 4015
rect 57340 3680 57345 4000
rect 57365 3680 57370 4000
rect 57340 3665 57370 3680
rect 57400 4000 57430 4070
rect 57455 4050 57495 4055
rect 57455 4020 57460 4050
rect 57490 4020 57495 4050
rect 57455 4015 57495 4020
rect 57400 3680 57405 4000
rect 57425 3680 57430 4000
rect 57400 3670 57430 3680
rect 57460 4000 57490 4015
rect 57460 3680 57465 4000
rect 57485 3680 57490 4000
rect 57460 3665 57490 3680
rect 57520 4000 57550 4070
rect 57575 4050 57615 4055
rect 57575 4020 57580 4050
rect 57610 4020 57615 4050
rect 57575 4015 57615 4020
rect 57520 3680 57525 4000
rect 57545 3680 57550 4000
rect 57520 3670 57550 3680
rect 57580 4000 57610 4015
rect 57580 3680 57585 4000
rect 57605 3680 57610 4000
rect 57580 3665 57610 3680
rect 57640 4000 57670 4070
rect 57695 4050 57735 4055
rect 57695 4020 57700 4050
rect 57730 4020 57735 4050
rect 57695 4015 57735 4020
rect 57640 3680 57645 4000
rect 57665 3680 57670 4000
rect 57640 3670 57670 3680
rect 57700 4000 57730 4015
rect 57700 3680 57705 4000
rect 57725 3680 57730 4000
rect 57700 3665 57730 3680
rect 57760 4000 57790 4070
rect 57760 3680 57765 4000
rect 57785 3680 57790 4000
rect 57040 3620 57045 3640
rect 57065 3620 57070 3640
rect 57040 3610 57070 3620
rect 57095 3660 57135 3665
rect 57095 3630 57100 3660
rect 57130 3630 57135 3660
rect 56925 3535 56965 3540
rect 56925 3505 56930 3535
rect 56960 3505 56965 3535
rect 56925 3500 56965 3505
rect 56065 3490 56705 3495
rect 56065 3460 56070 3490
rect 56100 3460 56110 3490
rect 56140 3460 56150 3490
rect 56180 3460 56190 3490
rect 56220 3460 56230 3490
rect 56260 3460 56270 3490
rect 56300 3460 56310 3490
rect 56340 3460 56350 3490
rect 56380 3460 56390 3490
rect 56420 3460 56430 3490
rect 56460 3460 56470 3490
rect 56500 3460 56510 3490
rect 56540 3460 56550 3490
rect 56580 3460 56590 3490
rect 56620 3460 56630 3490
rect 56660 3460 56670 3490
rect 56700 3460 56705 3490
rect 56065 3450 56705 3460
rect 56065 3420 56070 3450
rect 56100 3420 56110 3450
rect 56140 3420 56150 3450
rect 56180 3420 56190 3450
rect 56220 3420 56230 3450
rect 56260 3420 56270 3450
rect 56300 3420 56310 3450
rect 56340 3420 56350 3450
rect 56380 3420 56390 3450
rect 56420 3420 56430 3450
rect 56460 3420 56470 3450
rect 56500 3420 56510 3450
rect 56540 3420 56550 3450
rect 56580 3420 56590 3450
rect 56620 3420 56630 3450
rect 56660 3420 56670 3450
rect 56700 3420 56705 3450
rect 56065 3410 56705 3420
rect 56065 3380 56070 3410
rect 56100 3380 56110 3410
rect 56140 3380 56150 3410
rect 56180 3380 56190 3410
rect 56220 3380 56230 3410
rect 56260 3380 56270 3410
rect 56300 3380 56310 3410
rect 56340 3380 56350 3410
rect 56380 3380 56390 3410
rect 56420 3380 56430 3410
rect 56460 3380 56470 3410
rect 56500 3380 56510 3410
rect 56540 3380 56550 3410
rect 56580 3380 56590 3410
rect 56620 3380 56630 3410
rect 56660 3380 56670 3410
rect 56700 3380 56705 3410
rect 56065 3375 56705 3380
rect 57095 3495 57135 3630
rect 57215 3660 57255 3665
rect 57215 3630 57220 3660
rect 57250 3630 57255 3660
rect 57215 3495 57255 3630
rect 57335 3660 57375 3665
rect 57335 3630 57340 3660
rect 57370 3630 57375 3660
rect 57335 3495 57375 3630
rect 57455 3660 57495 3665
rect 57455 3630 57460 3660
rect 57490 3630 57495 3660
rect 57395 3580 57435 3585
rect 57395 3550 57400 3580
rect 57430 3550 57435 3580
rect 57395 3545 57435 3550
rect 57455 3495 57495 3630
rect 57575 3660 57615 3665
rect 57575 3630 57580 3660
rect 57610 3630 57615 3660
rect 57575 3495 57615 3630
rect 57695 3660 57735 3665
rect 57695 3630 57700 3660
rect 57730 3630 57735 3660
rect 57695 3495 57735 3630
rect 57760 3640 57790 3680
rect 57760 3620 57765 3640
rect 57785 3620 57790 3640
rect 57760 3610 57790 3620
rect 57095 3490 57735 3495
rect 57095 3460 57100 3490
rect 57130 3460 57140 3490
rect 57170 3460 57180 3490
rect 57210 3460 57220 3490
rect 57250 3460 57260 3490
rect 57290 3460 57300 3490
rect 57330 3460 57340 3490
rect 57370 3460 57380 3490
rect 57410 3460 57420 3490
rect 57450 3460 57460 3490
rect 57490 3460 57500 3490
rect 57530 3460 57540 3490
rect 57570 3460 57580 3490
rect 57610 3460 57620 3490
rect 57650 3460 57660 3490
rect 57690 3460 57700 3490
rect 57730 3460 57735 3490
rect 57095 3450 57735 3460
rect 57095 3420 57100 3450
rect 57130 3420 57140 3450
rect 57170 3420 57180 3450
rect 57210 3420 57220 3450
rect 57250 3420 57260 3450
rect 57290 3420 57300 3450
rect 57330 3420 57340 3450
rect 57370 3420 57380 3450
rect 57410 3420 57420 3450
rect 57450 3420 57460 3450
rect 57490 3420 57500 3450
rect 57530 3420 57540 3450
rect 57570 3420 57580 3450
rect 57610 3420 57620 3450
rect 57650 3420 57660 3450
rect 57690 3420 57700 3450
rect 57730 3420 57735 3450
rect 57095 3410 57735 3420
rect 57095 3380 57100 3410
rect 57130 3380 57140 3410
rect 57170 3380 57180 3410
rect 57210 3380 57220 3410
rect 57250 3380 57260 3410
rect 57290 3380 57300 3410
rect 57330 3380 57340 3410
rect 57370 3380 57380 3410
rect 57410 3380 57420 3410
rect 57450 3380 57460 3410
rect 57490 3380 57500 3410
rect 57530 3380 57540 3410
rect 57570 3380 57580 3410
rect 57610 3380 57620 3410
rect 57650 3380 57660 3410
rect 57690 3380 57700 3410
rect 57730 3380 57735 3410
rect 57095 3375 57735 3380
rect 55535 3325 55540 3355
rect 55570 3325 55580 3355
rect 55610 3325 55620 3355
rect 55650 3325 55655 3355
rect 55535 3315 55655 3325
rect 55535 3285 55540 3315
rect 55570 3285 55580 3315
rect 55610 3285 55620 3315
rect 55650 3285 55655 3315
rect 55535 3275 55655 3285
rect 55535 3245 55540 3275
rect 55570 3245 55580 3275
rect 55610 3245 55620 3275
rect 55650 3245 55655 3275
rect 55535 2185 55655 3245
rect 56510 3355 56550 3360
rect 56510 3325 56515 3355
rect 56545 3325 56550 3355
rect 56510 3315 56550 3325
rect 56510 3285 56515 3315
rect 56545 3285 56550 3315
rect 56510 3275 56550 3285
rect 56510 3245 56515 3275
rect 56545 3245 56550 3275
rect 56510 3240 56550 3245
rect 56680 3355 56710 3360
rect 56680 3315 56710 3325
rect 56680 3275 56710 3285
rect 56680 3240 56710 3245
rect 56840 3355 56880 3360
rect 56840 3325 56845 3355
rect 56875 3325 56880 3355
rect 56840 3315 56880 3325
rect 56840 3285 56845 3315
rect 56875 3285 56880 3315
rect 56840 3275 56880 3285
rect 56840 3245 56845 3275
rect 56875 3245 56880 3275
rect 56840 3240 56880 3245
rect 56920 3355 56960 3360
rect 56920 3325 56925 3355
rect 56955 3325 56960 3355
rect 56920 3315 56960 3325
rect 56920 3285 56925 3315
rect 56955 3285 56960 3315
rect 56920 3275 56960 3285
rect 56920 3245 56925 3275
rect 56955 3245 56960 3275
rect 56920 3240 56960 3245
rect 57090 3355 57120 3360
rect 57090 3315 57120 3325
rect 57090 3275 57120 3285
rect 57090 3240 57120 3245
rect 57250 3355 57290 3360
rect 57250 3325 57255 3355
rect 57285 3325 57290 3355
rect 57250 3315 57290 3325
rect 57250 3285 57255 3315
rect 57285 3285 57290 3315
rect 57250 3275 57290 3285
rect 57250 3245 57255 3275
rect 57285 3245 57290 3275
rect 57250 3240 57290 3245
rect 58145 3355 58265 4210
rect 58450 4320 58490 4325
rect 58450 4290 58455 4320
rect 58485 4290 58490 4320
rect 58450 4280 58490 4290
rect 58450 4250 58455 4280
rect 58485 4250 58490 4280
rect 58450 4240 58490 4250
rect 58450 4210 58455 4240
rect 58485 4210 58490 4240
rect 58450 4050 58490 4210
rect 58810 4320 58850 4325
rect 58810 4290 58815 4320
rect 58845 4290 58850 4320
rect 58810 4280 58850 4290
rect 58810 4250 58815 4280
rect 58845 4250 58850 4280
rect 58810 4240 58850 4250
rect 58810 4210 58815 4240
rect 58845 4210 58850 4240
rect 58510 4185 58790 4190
rect 58510 4155 58515 4185
rect 58545 4155 58555 4185
rect 58585 4155 58595 4185
rect 58625 4155 58635 4185
rect 58665 4155 58675 4185
rect 58705 4155 58715 4185
rect 58745 4155 58755 4185
rect 58785 4155 58790 4185
rect 58510 4145 58790 4155
rect 58510 4115 58515 4145
rect 58545 4115 58555 4145
rect 58585 4115 58595 4145
rect 58625 4115 58635 4145
rect 58665 4115 58675 4145
rect 58705 4115 58715 4145
rect 58745 4115 58755 4145
rect 58785 4115 58790 4145
rect 58510 4105 58790 4115
rect 58510 4075 58515 4105
rect 58545 4075 58555 4105
rect 58585 4075 58595 4105
rect 58625 4075 58635 4105
rect 58665 4075 58675 4105
rect 58705 4075 58715 4105
rect 58745 4075 58755 4105
rect 58785 4075 58790 4105
rect 58510 4070 58790 4075
rect 58450 4020 58455 4050
rect 58485 4020 58490 4050
rect 58450 4015 58490 4020
rect 58455 4000 58485 4015
rect 58455 3680 58460 4000
rect 58480 3680 58485 4000
rect 58455 3640 58485 3680
rect 58515 4000 58545 4070
rect 58570 4050 58610 4055
rect 58570 4020 58575 4050
rect 58605 4020 58610 4050
rect 58570 4015 58610 4020
rect 58515 3680 58520 4000
rect 58540 3680 58545 4000
rect 58515 3665 58545 3680
rect 58575 4000 58605 4015
rect 58575 3680 58580 4000
rect 58600 3680 58605 4000
rect 58575 3670 58605 3680
rect 58635 4000 58665 4070
rect 58690 4050 58730 4055
rect 58690 4020 58695 4050
rect 58725 4020 58730 4050
rect 58690 4015 58730 4020
rect 58635 3680 58640 4000
rect 58660 3680 58665 4000
rect 58635 3665 58665 3680
rect 58695 4000 58725 4015
rect 58695 3680 58700 4000
rect 58720 3680 58725 4000
rect 58695 3670 58725 3680
rect 58755 4000 58785 4070
rect 58810 4050 58850 4210
rect 59170 4320 59210 4325
rect 59170 4290 59175 4320
rect 59205 4290 59210 4320
rect 59170 4280 59210 4290
rect 59170 4250 59175 4280
rect 59205 4250 59210 4280
rect 59170 4240 59210 4250
rect 59170 4210 59175 4240
rect 59205 4210 59210 4240
rect 58870 4185 59150 4190
rect 58870 4155 58875 4185
rect 58905 4155 58915 4185
rect 58945 4155 58955 4185
rect 58985 4155 58995 4185
rect 59025 4155 59035 4185
rect 59065 4155 59075 4185
rect 59105 4155 59115 4185
rect 59145 4155 59150 4185
rect 58870 4145 59150 4155
rect 58870 4115 58875 4145
rect 58905 4115 58915 4145
rect 58945 4115 58955 4145
rect 58985 4115 58995 4145
rect 59025 4115 59035 4145
rect 59065 4115 59075 4145
rect 59105 4115 59115 4145
rect 59145 4115 59150 4145
rect 58870 4105 59150 4115
rect 58870 4075 58875 4105
rect 58905 4075 58915 4105
rect 58945 4075 58955 4105
rect 58985 4075 58995 4105
rect 59025 4075 59035 4105
rect 59065 4075 59075 4105
rect 59105 4075 59115 4105
rect 59145 4075 59150 4105
rect 58870 4070 59150 4075
rect 58810 4020 58815 4050
rect 58845 4020 58850 4050
rect 58810 4015 58850 4020
rect 58755 3680 58760 4000
rect 58780 3680 58785 4000
rect 58755 3665 58785 3680
rect 58815 4000 58845 4015
rect 58815 3680 58820 4000
rect 58840 3680 58845 4000
rect 58815 3670 58845 3680
rect 58875 4000 58905 4070
rect 58930 4050 58970 4055
rect 58930 4020 58935 4050
rect 58965 4020 58970 4050
rect 58930 4015 58970 4020
rect 58875 3680 58880 4000
rect 58900 3680 58905 4000
rect 58875 3665 58905 3680
rect 58935 4000 58965 4015
rect 58935 3680 58940 4000
rect 58960 3680 58965 4000
rect 58935 3670 58965 3680
rect 58995 4000 59025 4070
rect 59050 4050 59090 4055
rect 59050 4020 59055 4050
rect 59085 4020 59090 4050
rect 59050 4015 59090 4020
rect 58995 3680 59000 4000
rect 59020 3680 59025 4000
rect 58995 3665 59025 3680
rect 59055 4000 59085 4015
rect 59055 3680 59060 4000
rect 59080 3680 59085 4000
rect 59055 3670 59085 3680
rect 59115 4000 59145 4070
rect 59170 4050 59210 4210
rect 59640 4320 59760 6110
rect 59640 4290 59645 4320
rect 59675 4290 59685 4320
rect 59715 4290 59725 4320
rect 59755 4290 59760 4320
rect 59640 4280 59760 4290
rect 59640 4250 59645 4280
rect 59675 4250 59685 4280
rect 59715 4250 59725 4280
rect 59755 4250 59760 4280
rect 59640 4240 59760 4250
rect 59640 4210 59645 4240
rect 59675 4210 59685 4240
rect 59715 4210 59725 4240
rect 59755 4210 59760 4240
rect 59640 4205 59760 4210
rect 60340 4320 60460 6110
rect 60340 4290 60345 4320
rect 60375 4290 60385 4320
rect 60415 4290 60425 4320
rect 60455 4290 60460 4320
rect 60340 4280 60460 4290
rect 60340 4250 60345 4280
rect 60375 4250 60385 4280
rect 60415 4250 60425 4280
rect 60455 4250 60460 4280
rect 60340 4240 60460 4250
rect 60340 4210 60345 4240
rect 60375 4210 60385 4240
rect 60415 4210 60425 4240
rect 60455 4210 60460 4240
rect 60340 4205 60460 4210
rect 60690 4320 60810 6110
rect 60690 4290 60695 4320
rect 60725 4290 60735 4320
rect 60765 4290 60775 4320
rect 60805 4290 60810 4320
rect 60690 4280 60810 4290
rect 60690 4250 60695 4280
rect 60725 4250 60735 4280
rect 60765 4250 60775 4280
rect 60805 4250 60810 4280
rect 60690 4240 60810 4250
rect 60690 4210 60695 4240
rect 60725 4210 60735 4240
rect 60765 4210 60775 4240
rect 60805 4210 60810 4240
rect 60690 4205 60810 4210
rect 61040 4320 61160 6110
rect 61040 4290 61045 4320
rect 61075 4290 61085 4320
rect 61115 4290 61125 4320
rect 61155 4290 61160 4320
rect 61040 4280 61160 4290
rect 61040 4250 61045 4280
rect 61075 4250 61085 4280
rect 61115 4250 61125 4280
rect 61155 4250 61160 4280
rect 61040 4240 61160 4250
rect 61040 4210 61045 4240
rect 61075 4210 61085 4240
rect 61115 4210 61125 4240
rect 61155 4210 61160 4240
rect 61040 4205 61160 4210
rect 61390 4320 61510 6110
rect 61390 4290 61395 4320
rect 61425 4290 61435 4320
rect 61465 4290 61475 4320
rect 61505 4290 61510 4320
rect 61390 4280 61510 4290
rect 61390 4250 61395 4280
rect 61425 4250 61435 4280
rect 61465 4250 61475 4280
rect 61505 4250 61510 4280
rect 61390 4240 61510 4250
rect 61390 4210 61395 4240
rect 61425 4210 61435 4240
rect 61465 4210 61475 4240
rect 61505 4210 61510 4240
rect 61390 4205 61510 4210
rect 59170 4020 59175 4050
rect 59205 4020 59210 4050
rect 59170 4015 59210 4020
rect 59115 3680 59120 4000
rect 59140 3680 59145 4000
rect 59115 3665 59145 3680
rect 59175 4000 59205 4015
rect 59175 3680 59180 4000
rect 59200 3680 59205 4000
rect 58455 3620 58460 3640
rect 58480 3620 58485 3640
rect 58510 3660 58550 3665
rect 58510 3630 58515 3660
rect 58545 3630 58550 3660
rect 58510 3625 58550 3630
rect 58630 3660 58670 3665
rect 58630 3630 58635 3660
rect 58665 3630 58670 3660
rect 58630 3625 58670 3630
rect 58750 3660 58790 3665
rect 58750 3630 58755 3660
rect 58785 3630 58790 3660
rect 58750 3625 58790 3630
rect 58870 3660 58910 3665
rect 58870 3630 58875 3660
rect 58905 3630 58910 3660
rect 58870 3625 58910 3630
rect 58990 3660 59030 3665
rect 58990 3630 58995 3660
rect 59025 3630 59030 3660
rect 58990 3625 59030 3630
rect 59110 3660 59150 3665
rect 59110 3630 59115 3660
rect 59145 3630 59150 3660
rect 59110 3625 59150 3630
rect 59175 3640 59205 3680
rect 58455 3610 58485 3620
rect 59175 3620 59180 3640
rect 59200 3620 59205 3640
rect 59175 3610 59205 3620
rect 58810 3535 58850 3540
rect 58810 3505 58815 3535
rect 58845 3505 58850 3535
rect 58810 3500 58850 3505
rect 58145 3325 58150 3355
rect 58180 3325 58190 3355
rect 58220 3325 58230 3355
rect 58260 3325 58265 3355
rect 58145 3315 58265 3325
rect 58145 3285 58150 3315
rect 58180 3285 58190 3315
rect 58220 3285 58230 3315
rect 58260 3285 58265 3315
rect 58145 3275 58265 3285
rect 58145 3245 58150 3275
rect 58180 3245 58190 3275
rect 58220 3245 58230 3275
rect 58260 3245 58265 3275
rect 56620 3220 56660 3225
rect 56620 3190 56625 3220
rect 56655 3190 56660 3220
rect 56620 3185 56660 3190
rect 56730 3220 56770 3225
rect 56730 3190 56735 3220
rect 56765 3190 56770 3220
rect 56730 3185 56770 3190
rect 57030 3220 57070 3225
rect 57030 3190 57035 3220
rect 57065 3190 57070 3220
rect 57030 3185 57070 3190
rect 57140 3220 57180 3225
rect 57140 3190 57145 3220
rect 57175 3190 57180 3220
rect 57140 3185 57180 3190
rect 56560 2910 56590 2915
rect 56800 2910 56830 2915
rect 56560 2875 56590 2880
rect 56607 2895 56637 2905
rect 56607 2875 56612 2895
rect 56632 2875 56637 2895
rect 56607 2865 56637 2875
rect 56675 2900 56715 2905
rect 56675 2870 56680 2900
rect 56710 2870 56715 2900
rect 56675 2865 56715 2870
rect 56753 2895 56783 2905
rect 56753 2875 56758 2895
rect 56778 2875 56783 2895
rect 56800 2875 56830 2880
rect 56970 2905 57000 2915
rect 57210 2905 57240 2915
rect 56970 2885 56975 2905
rect 56995 2885 57000 2905
rect 56970 2875 57000 2885
rect 57017 2895 57047 2905
rect 57017 2875 57022 2895
rect 57042 2875 57047 2895
rect 56753 2865 56783 2875
rect 56610 2835 56630 2865
rect 56600 2830 56640 2835
rect 56600 2800 56605 2830
rect 56635 2800 56640 2830
rect 56600 2795 56640 2800
rect 56760 2785 56780 2865
rect 55950 2780 55990 2785
rect 55950 2750 55955 2780
rect 55985 2750 55990 2780
rect 55950 2745 55990 2750
rect 56745 2780 56785 2785
rect 56745 2750 56750 2780
rect 56780 2750 56785 2780
rect 56745 2745 56785 2750
rect 55535 2155 55540 2185
rect 55570 2155 55580 2185
rect 55610 2155 55620 2185
rect 55650 2155 55655 2185
rect 55535 2145 55655 2155
rect 55535 2115 55540 2145
rect 55570 2115 55580 2145
rect 55610 2115 55620 2145
rect 55650 2115 55655 2145
rect 55535 2105 55655 2115
rect 55535 2075 55540 2105
rect 55570 2075 55580 2105
rect 55610 2075 55620 2105
rect 55650 2075 55655 2105
rect 54530 1475 54570 1480
rect 54530 1445 54535 1475
rect 54565 1445 54570 1475
rect 54530 1440 54570 1445
rect 54730 1475 54770 1480
rect 54730 1445 54735 1475
rect 54765 1445 54770 1475
rect 54730 1440 54770 1445
rect 54840 1475 54880 1480
rect 54840 1445 54845 1475
rect 54875 1445 54880 1475
rect 54840 1440 54880 1445
rect 54950 1475 54990 1480
rect 54950 1445 54955 1475
rect 54985 1445 54990 1475
rect 54950 1440 54990 1445
rect 55060 1475 55100 1480
rect 55060 1445 55065 1475
rect 55095 1445 55100 1475
rect 55060 1440 55100 1445
rect 55170 1475 55210 1480
rect 55170 1445 55175 1475
rect 55205 1445 55210 1475
rect 55170 1440 55210 1445
rect 54540 1160 54560 1440
rect 54625 1425 54655 1435
rect 54530 1155 54570 1160
rect 54530 1125 54535 1155
rect 54565 1125 54570 1155
rect 54530 1120 54570 1125
rect 54625 1155 54630 1425
rect 54650 1155 54655 1425
rect 54625 1115 54655 1155
rect 54625 1095 54630 1115
rect 54650 1095 54655 1115
rect 54375 1085 54415 1090
rect 54375 1055 54380 1085
rect 54410 1055 54415 1085
rect 54375 1050 54415 1055
rect 54485 1085 54525 1090
rect 54485 1055 54490 1085
rect 54520 1055 54525 1085
rect 54485 1050 54525 1055
rect 54625 945 54655 1095
rect 54680 1425 54710 1435
rect 54680 1155 54685 1425
rect 54705 1155 54710 1425
rect 54680 1080 54710 1155
rect 54735 1425 54765 1440
rect 54735 1155 54740 1425
rect 54760 1155 54765 1425
rect 54735 1140 54765 1155
rect 54790 1425 54820 1435
rect 54790 1155 54795 1425
rect 54815 1155 54820 1425
rect 54730 1135 54770 1140
rect 54730 1105 54735 1135
rect 54765 1105 54770 1135
rect 54730 1100 54770 1105
rect 54790 1080 54820 1155
rect 54845 1425 54875 1440
rect 54845 1155 54850 1425
rect 54870 1155 54875 1425
rect 54845 1140 54875 1155
rect 54900 1425 54930 1435
rect 54900 1155 54905 1425
rect 54925 1155 54930 1425
rect 54840 1135 54880 1140
rect 54840 1105 54845 1135
rect 54875 1105 54880 1135
rect 54840 1100 54880 1105
rect 54900 1080 54930 1155
rect 54955 1425 54985 1440
rect 54955 1155 54960 1425
rect 54980 1155 54985 1425
rect 54955 1140 54985 1155
rect 55010 1425 55040 1435
rect 55010 1155 55015 1425
rect 55035 1155 55040 1425
rect 54950 1135 54990 1140
rect 54950 1105 54955 1135
rect 54985 1105 54990 1135
rect 54950 1100 54990 1105
rect 55010 1080 55040 1155
rect 55065 1425 55095 1440
rect 55065 1155 55070 1425
rect 55090 1155 55095 1425
rect 55065 1140 55095 1155
rect 55120 1425 55150 1435
rect 55120 1155 55125 1425
rect 55145 1155 55150 1425
rect 55060 1135 55100 1140
rect 55060 1105 55065 1135
rect 55095 1105 55100 1135
rect 55060 1100 55100 1105
rect 55120 1080 55150 1155
rect 55175 1425 55205 1440
rect 55175 1155 55180 1425
rect 55200 1155 55205 1425
rect 55175 1140 55205 1155
rect 55230 1425 55260 1435
rect 55230 1155 55235 1425
rect 55255 1155 55260 1425
rect 55170 1135 55210 1140
rect 55170 1105 55175 1135
rect 55205 1105 55210 1135
rect 55170 1100 55210 1105
rect 55230 1080 55260 1155
rect 55285 1425 55315 1435
rect 55285 1155 55290 1425
rect 55310 1155 55315 1425
rect 55285 1115 55315 1155
rect 55285 1095 55290 1115
rect 55310 1095 55315 1115
rect 54675 1075 54715 1080
rect 54675 1045 54680 1075
rect 54710 1045 54715 1075
rect 54675 1035 54715 1045
rect 54675 1005 54680 1035
rect 54710 1005 54715 1035
rect 54675 995 54715 1005
rect 54675 965 54680 995
rect 54710 965 54715 995
rect 54675 960 54715 965
rect 54785 1075 54825 1080
rect 54785 1045 54790 1075
rect 54820 1045 54825 1075
rect 54785 1035 54825 1045
rect 54785 1005 54790 1035
rect 54820 1005 54825 1035
rect 54785 995 54825 1005
rect 54785 965 54790 995
rect 54820 965 54825 995
rect 54785 960 54825 965
rect 54895 1075 54935 1080
rect 54895 1045 54900 1075
rect 54930 1045 54935 1075
rect 54895 1035 54935 1045
rect 54895 1005 54900 1035
rect 54930 1005 54935 1035
rect 54895 995 54935 1005
rect 54895 965 54900 995
rect 54930 965 54935 995
rect 54895 960 54935 965
rect 55005 1075 55045 1080
rect 55005 1045 55010 1075
rect 55040 1045 55045 1075
rect 55005 1035 55045 1045
rect 55005 1005 55010 1035
rect 55040 1005 55045 1035
rect 55005 995 55045 1005
rect 55005 965 55010 995
rect 55040 965 55045 995
rect 55005 960 55045 965
rect 55115 1075 55155 1080
rect 55115 1045 55120 1075
rect 55150 1045 55155 1075
rect 55115 1035 55155 1045
rect 55115 1005 55120 1035
rect 55150 1005 55155 1035
rect 55115 995 55155 1005
rect 55115 965 55120 995
rect 55150 965 55155 995
rect 55115 960 55155 965
rect 55225 1075 55265 1080
rect 55225 1045 55230 1075
rect 55260 1045 55265 1075
rect 55225 1035 55265 1045
rect 55225 1005 55230 1035
rect 55260 1005 55265 1035
rect 55225 995 55265 1005
rect 55225 965 55230 995
rect 55260 965 55265 995
rect 55225 960 55265 965
rect 55285 945 55315 1095
rect 55535 1075 55655 2075
rect 55670 2295 55790 2300
rect 55670 2265 55675 2295
rect 55705 2265 55715 2295
rect 55745 2265 55755 2295
rect 55785 2265 55790 2295
rect 55670 2255 55790 2265
rect 55670 2225 55675 2255
rect 55705 2225 55715 2255
rect 55745 2225 55755 2255
rect 55785 2225 55790 2255
rect 55670 2215 55790 2225
rect 55670 2185 55675 2215
rect 55705 2185 55715 2215
rect 55745 2185 55755 2215
rect 55785 2185 55790 2215
rect 55670 2050 55790 2185
rect 55670 2020 55675 2050
rect 55705 2020 55715 2050
rect 55745 2020 55755 2050
rect 55785 2020 55790 2050
rect 55670 2010 55790 2020
rect 55670 1980 55675 2010
rect 55705 1980 55715 2010
rect 55745 1980 55755 2010
rect 55785 1980 55790 2010
rect 55670 1970 55790 1980
rect 55670 1940 55675 1970
rect 55705 1940 55715 1970
rect 55745 1940 55755 1970
rect 55785 1940 55790 1970
rect 55885 1985 55925 1990
rect 55885 1955 55890 1985
rect 55920 1955 55925 1985
rect 55885 1950 55925 1955
rect 55670 1640 55790 1940
rect 55670 1610 55675 1640
rect 55705 1610 55715 1640
rect 55745 1610 55755 1640
rect 55785 1610 55790 1640
rect 55670 1600 55790 1610
rect 55670 1570 55675 1600
rect 55705 1570 55715 1600
rect 55745 1570 55755 1600
rect 55785 1570 55790 1600
rect 55670 1560 55790 1570
rect 55670 1530 55675 1560
rect 55705 1530 55715 1560
rect 55745 1530 55755 1560
rect 55785 1530 55790 1560
rect 55670 1525 55790 1530
rect 55535 1045 55540 1075
rect 55570 1045 55580 1075
rect 55610 1045 55620 1075
rect 55650 1045 55655 1075
rect 55535 1035 55655 1045
rect 55535 1005 55540 1035
rect 55570 1005 55580 1035
rect 55610 1005 55620 1035
rect 55650 1005 55655 1035
rect 55535 995 55655 1005
rect 55535 965 55540 995
rect 55570 965 55580 995
rect 55610 965 55620 995
rect 55650 965 55655 995
rect 55535 960 55655 965
rect 55670 1485 55790 1490
rect 55670 1455 55675 1485
rect 55705 1455 55715 1485
rect 55745 1455 55755 1485
rect 55785 1455 55790 1485
rect 55670 1445 55790 1455
rect 55670 1415 55675 1445
rect 55705 1415 55715 1445
rect 55745 1415 55755 1445
rect 55785 1415 55790 1445
rect 55670 1405 55790 1415
rect 55670 1375 55675 1405
rect 55705 1375 55715 1405
rect 55745 1375 55755 1405
rect 55785 1375 55790 1405
rect 54620 940 54660 945
rect 54620 910 54625 940
rect 54655 910 54660 940
rect 54620 900 54660 910
rect 54620 870 54625 900
rect 54655 870 54660 900
rect 54620 860 54660 870
rect 54620 830 54625 860
rect 54655 830 54660 860
rect 54620 825 54660 830
rect 55280 940 55320 945
rect 55280 910 55285 940
rect 55315 910 55320 940
rect 55280 900 55320 910
rect 55280 870 55285 900
rect 55315 870 55320 900
rect 55280 860 55320 870
rect 55280 830 55285 860
rect 55315 830 55320 860
rect 55280 825 55320 830
rect 54255 805 54295 810
rect 54255 775 54260 805
rect 54290 775 54295 805
rect 54255 770 54295 775
rect 54320 525 54360 530
rect 54320 495 54325 525
rect 54355 495 54360 525
rect 54320 490 54360 495
rect 55000 525 55040 530
rect 55000 495 55005 525
rect 55035 495 55040 525
rect 55000 490 55040 495
rect 53990 440 53995 470
rect 54025 440 54035 470
rect 54065 440 54080 470
rect 54110 440 54120 470
rect 54150 440 54165 470
rect 54195 440 54205 470
rect 54235 440 54240 470
rect 53990 430 54240 440
rect 53990 400 53995 430
rect 54025 400 54035 430
rect 54065 400 54080 430
rect 54110 400 54120 430
rect 54150 400 54165 430
rect 54195 400 54205 430
rect 54235 400 54240 430
rect 53990 390 54240 400
rect 53990 360 53995 390
rect 54025 360 54035 390
rect 54065 360 54080 390
rect 54110 360 54120 390
rect 54150 360 54165 390
rect 54195 360 54205 390
rect 54235 360 54240 390
rect 53990 355 54240 360
rect 54330 340 54350 490
rect 54385 470 54425 475
rect 54385 440 54390 470
rect 54420 440 54425 470
rect 54385 430 54425 440
rect 54385 400 54390 430
rect 54420 400 54425 430
rect 54385 390 54425 400
rect 54385 360 54390 390
rect 54420 360 54425 390
rect 54385 355 54425 360
rect 54750 470 55190 475
rect 54750 440 54755 470
rect 54785 440 54795 470
rect 54825 440 54835 470
rect 54865 440 54875 470
rect 54905 440 54915 470
rect 54945 440 54955 470
rect 54985 440 54995 470
rect 55025 440 55035 470
rect 55065 440 55075 470
rect 55105 440 55115 470
rect 55145 440 55155 470
rect 55185 440 55190 470
rect 54750 430 55190 440
rect 54750 400 54755 430
rect 54785 400 54795 430
rect 54825 400 54835 430
rect 54865 400 54875 430
rect 54905 400 54915 430
rect 54945 400 54955 430
rect 54985 400 54995 430
rect 55025 400 55035 430
rect 55065 400 55075 430
rect 55105 400 55115 430
rect 55145 400 55155 430
rect 55185 400 55190 430
rect 54750 390 55190 400
rect 54750 360 54755 390
rect 54785 360 54795 390
rect 54825 360 54835 390
rect 54865 360 54875 390
rect 54905 360 54915 390
rect 54945 360 54955 390
rect 54985 360 54995 390
rect 55025 360 55035 390
rect 55065 360 55075 390
rect 55105 360 55115 390
rect 55145 360 55155 390
rect 55185 360 55190 390
rect 54750 355 55190 360
rect 54325 335 54360 340
rect 54325 295 54360 300
rect 54385 335 54420 355
rect 54385 295 54420 300
rect 54655 325 54685 335
rect 54655 -345 54660 325
rect 54680 -345 54685 325
rect 54655 -385 54685 -345
rect 54755 325 54785 355
rect 54755 -345 54760 325
rect 54780 -345 54785 325
rect 54755 -360 54785 -345
rect 54855 325 54885 335
rect 54855 -345 54860 325
rect 54880 -345 54885 325
rect 54655 -405 54660 -385
rect 54680 -405 54685 -385
rect 54750 -365 54790 -360
rect 54750 -395 54755 -365
rect 54785 -395 54790 -365
rect 54750 -400 54790 -395
rect 54655 -575 54685 -405
rect 54855 -575 54885 -345
rect 54955 325 54985 355
rect 54955 -345 54960 325
rect 54980 -345 54985 325
rect 54955 -360 54985 -345
rect 55055 325 55085 335
rect 55055 -345 55060 325
rect 55080 -345 55085 325
rect 54950 -365 54990 -360
rect 54950 -395 54955 -365
rect 54985 -395 54990 -365
rect 54950 -400 54990 -395
rect 53840 -610 53845 -580
rect 53875 -610 53885 -580
rect 53915 -610 53925 -580
rect 53955 -610 53960 -580
rect 53840 -620 53960 -610
rect 53840 -650 53845 -620
rect 53875 -650 53885 -620
rect 53915 -650 53925 -620
rect 53955 -650 53960 -620
rect 53840 -660 53960 -650
rect 53840 -690 53845 -660
rect 53875 -690 53885 -660
rect 53915 -690 53925 -660
rect 53955 -690 53960 -660
rect 53840 -695 53960 -690
rect 54040 -580 54160 -575
rect 54040 -610 54045 -580
rect 54075 -610 54085 -580
rect 54115 -610 54125 -580
rect 54155 -610 54160 -580
rect 54040 -620 54160 -610
rect 54040 -650 54045 -620
rect 54075 -650 54085 -620
rect 54115 -650 54125 -620
rect 54155 -650 54160 -620
rect 54040 -660 54160 -650
rect 54040 -690 54045 -660
rect 54075 -690 54085 -660
rect 54115 -690 54125 -660
rect 54155 -690 54160 -660
rect 54040 -1500 54160 -690
rect 54390 -580 54510 -575
rect 54390 -610 54395 -580
rect 54425 -610 54435 -580
rect 54465 -610 54475 -580
rect 54505 -610 54510 -580
rect 54390 -620 54510 -610
rect 54390 -650 54395 -620
rect 54425 -650 54435 -620
rect 54465 -650 54475 -620
rect 54505 -650 54510 -620
rect 54390 -660 54510 -650
rect 54390 -690 54395 -660
rect 54425 -690 54435 -660
rect 54465 -690 54475 -660
rect 54505 -690 54510 -660
rect 54390 -1500 54510 -690
rect 54650 -580 54690 -575
rect 54650 -610 54655 -580
rect 54685 -610 54690 -580
rect 54650 -620 54690 -610
rect 54650 -650 54655 -620
rect 54685 -650 54690 -620
rect 54650 -660 54690 -650
rect 54650 -690 54655 -660
rect 54685 -690 54690 -660
rect 54650 -695 54690 -690
rect 54740 -580 54885 -575
rect 54740 -610 54745 -580
rect 54775 -610 54785 -580
rect 54815 -610 54825 -580
rect 54855 -610 54885 -580
rect 54740 -620 54885 -610
rect 54740 -650 54745 -620
rect 54775 -650 54785 -620
rect 54815 -650 54825 -620
rect 54855 -650 54885 -620
rect 54740 -660 54885 -650
rect 54740 -690 54745 -660
rect 54775 -690 54785 -660
rect 54815 -690 54825 -660
rect 54855 -690 54885 -660
rect 54740 -695 54885 -690
rect 55055 -575 55085 -345
rect 55155 325 55185 355
rect 55155 -345 55160 325
rect 55180 -345 55185 325
rect 55155 -360 55185 -345
rect 55255 325 55285 335
rect 55255 -345 55260 325
rect 55280 -345 55285 325
rect 55670 -60 55790 1375
rect 55670 -90 55675 -60
rect 55705 -90 55715 -60
rect 55745 -90 55755 -60
rect 55785 -90 55790 -60
rect 55670 -100 55790 -90
rect 55670 -130 55675 -100
rect 55705 -130 55715 -100
rect 55745 -130 55755 -100
rect 55785 -130 55790 -100
rect 55670 -140 55790 -130
rect 55670 -170 55675 -140
rect 55705 -170 55715 -140
rect 55745 -170 55755 -140
rect 55785 -170 55790 -140
rect 55670 -175 55790 -170
rect 55895 -245 55915 1950
rect 55950 810 55970 2745
rect 56970 2730 56990 2875
rect 57017 2865 57047 2875
rect 57085 2900 57125 2905
rect 57085 2870 57090 2900
rect 57120 2870 57125 2900
rect 57085 2865 57125 2870
rect 57163 2895 57193 2905
rect 57163 2875 57168 2895
rect 57188 2875 57193 2895
rect 57210 2885 57215 2905
rect 57235 2885 57240 2905
rect 57210 2875 57240 2885
rect 57163 2865 57193 2875
rect 57020 2785 57040 2865
rect 57170 2835 57190 2865
rect 57160 2830 57200 2835
rect 57160 2800 57165 2830
rect 57195 2800 57200 2830
rect 57160 2795 57200 2800
rect 57015 2780 57055 2785
rect 57015 2750 57020 2780
rect 57050 2750 57055 2780
rect 57015 2745 57055 2750
rect 56850 2725 56890 2730
rect 56850 2695 56855 2725
rect 56885 2695 56890 2725
rect 56850 2690 56890 2695
rect 56960 2725 57000 2730
rect 56960 2695 56965 2725
rect 56995 2695 57000 2725
rect 56960 2690 57000 2695
rect 56860 2620 56880 2690
rect 57220 2675 57240 2875
rect 57810 2780 57850 2785
rect 57810 2750 57815 2780
rect 57845 2750 57850 2780
rect 57810 2745 57850 2750
rect 56935 2670 56975 2675
rect 56935 2640 56940 2670
rect 56970 2640 56975 2670
rect 56935 2635 56975 2640
rect 57210 2670 57250 2675
rect 57210 2640 57215 2670
rect 57245 2640 57250 2670
rect 57210 2635 57250 2640
rect 56945 2620 56965 2635
rect 56830 2615 56890 2620
rect 56830 2585 56855 2615
rect 56885 2585 56890 2615
rect 56830 2580 56890 2585
rect 56935 2610 56975 2620
rect 56935 2590 56945 2610
rect 56965 2590 56975 2610
rect 56935 2580 56975 2590
rect 56775 2550 56805 2560
rect 56085 2470 56675 2475
rect 56085 2440 56090 2470
rect 56120 2440 56145 2470
rect 56175 2440 56200 2470
rect 56230 2440 56255 2470
rect 56285 2440 56310 2470
rect 56340 2440 56365 2470
rect 56395 2440 56420 2470
rect 56450 2440 56475 2470
rect 56505 2440 56530 2470
rect 56560 2440 56585 2470
rect 56615 2440 56640 2470
rect 56670 2440 56675 2470
rect 56085 2430 56675 2440
rect 56085 2400 56090 2430
rect 56120 2400 56145 2430
rect 56175 2400 56200 2430
rect 56230 2400 56255 2430
rect 56285 2400 56310 2430
rect 56340 2400 56365 2430
rect 56395 2400 56420 2430
rect 56450 2400 56475 2430
rect 56505 2400 56530 2430
rect 56560 2400 56585 2430
rect 56615 2400 56640 2430
rect 56670 2400 56675 2430
rect 56085 2390 56675 2400
rect 56085 2360 56090 2390
rect 56120 2360 56145 2390
rect 56175 2360 56200 2390
rect 56230 2360 56255 2390
rect 56285 2360 56310 2390
rect 56340 2360 56365 2390
rect 56395 2360 56420 2390
rect 56450 2360 56475 2390
rect 56505 2360 56530 2390
rect 56560 2360 56585 2390
rect 56615 2360 56640 2390
rect 56670 2360 56675 2390
rect 56085 2355 56675 2360
rect 56040 1985 56070 1990
rect 56040 1950 56070 1955
rect 56085 1930 56125 2355
rect 56140 1975 56180 1980
rect 56140 1945 56145 1975
rect 56175 1945 56180 1975
rect 56140 1940 56180 1945
rect 56085 1900 56090 1930
rect 56120 1900 56125 1930
rect 56085 1895 56125 1900
rect 56030 1880 56065 1890
rect 56030 1760 56040 1880
rect 56060 1760 56065 1880
rect 56030 1750 56065 1760
rect 56035 1745 56065 1750
rect 56090 1880 56120 1895
rect 56090 1760 56095 1880
rect 56115 1760 56120 1880
rect 56035 1720 56065 1730
rect 56035 1700 56040 1720
rect 56060 1700 56065 1720
rect 56090 1700 56120 1760
rect 56145 1880 56175 1940
rect 56195 1930 56235 2355
rect 56250 1975 56290 1980
rect 56250 1945 56255 1975
rect 56285 1945 56290 1975
rect 56250 1940 56290 1945
rect 56195 1900 56200 1930
rect 56230 1900 56235 1930
rect 56195 1895 56235 1900
rect 56145 1760 56150 1880
rect 56170 1760 56175 1880
rect 56145 1745 56175 1760
rect 56200 1880 56230 1895
rect 56200 1760 56205 1880
rect 56225 1760 56230 1880
rect 56140 1740 56180 1745
rect 56140 1710 56145 1740
rect 56175 1710 56180 1740
rect 56140 1705 56180 1710
rect 56035 1645 56065 1700
rect 56085 1695 56125 1700
rect 56085 1665 56090 1695
rect 56120 1665 56125 1695
rect 56085 1660 56125 1665
rect 56030 1640 56070 1645
rect 56030 1610 56035 1640
rect 56065 1610 56070 1640
rect 56030 1600 56070 1610
rect 56030 1570 56035 1600
rect 56065 1570 56070 1600
rect 56030 1560 56070 1570
rect 56030 1530 56035 1560
rect 56065 1530 56070 1560
rect 56030 1525 56070 1530
rect 56145 1315 56175 1705
rect 56200 1700 56230 1760
rect 56255 1880 56285 1940
rect 56305 1930 56345 2355
rect 56360 1975 56400 1980
rect 56360 1945 56365 1975
rect 56395 1945 56400 1975
rect 56360 1940 56400 1945
rect 56305 1900 56310 1930
rect 56340 1900 56345 1930
rect 56305 1895 56345 1900
rect 56255 1760 56260 1880
rect 56280 1760 56285 1880
rect 56255 1745 56285 1760
rect 56310 1880 56340 1895
rect 56310 1760 56315 1880
rect 56335 1760 56340 1880
rect 56250 1740 56290 1745
rect 56250 1710 56255 1740
rect 56285 1710 56290 1740
rect 56250 1705 56290 1710
rect 56195 1695 56235 1700
rect 56195 1665 56200 1695
rect 56230 1665 56235 1695
rect 56195 1660 56235 1665
rect 56085 1305 56125 1310
rect 56040 1295 56070 1300
rect 56085 1275 56090 1305
rect 56120 1275 56125 1305
rect 56255 1315 56285 1705
rect 56310 1700 56340 1760
rect 56365 1880 56395 1940
rect 56415 1930 56455 2355
rect 56470 1975 56510 1980
rect 56470 1945 56475 1975
rect 56505 1945 56510 1975
rect 56470 1940 56510 1945
rect 56415 1900 56420 1930
rect 56450 1900 56455 1930
rect 56415 1895 56455 1900
rect 56365 1760 56370 1880
rect 56390 1760 56395 1880
rect 56365 1745 56395 1760
rect 56420 1880 56450 1895
rect 56420 1760 56425 1880
rect 56445 1760 56450 1880
rect 56360 1740 56400 1745
rect 56360 1710 56365 1740
rect 56395 1710 56400 1740
rect 56360 1705 56400 1710
rect 56305 1695 56345 1700
rect 56305 1665 56310 1695
rect 56340 1665 56345 1695
rect 56305 1660 56345 1665
rect 56145 1280 56175 1285
rect 56195 1305 56235 1310
rect 56085 1270 56125 1275
rect 56195 1275 56200 1305
rect 56230 1275 56235 1305
rect 56365 1315 56395 1705
rect 56420 1700 56450 1760
rect 56475 1880 56505 1940
rect 56525 1930 56565 2355
rect 56580 1975 56620 1980
rect 56580 1945 56585 1975
rect 56615 1945 56620 1975
rect 56580 1940 56620 1945
rect 56525 1900 56530 1930
rect 56560 1900 56565 1930
rect 56525 1895 56565 1900
rect 56475 1760 56480 1880
rect 56500 1760 56505 1880
rect 56475 1745 56505 1760
rect 56530 1880 56560 1895
rect 56530 1760 56535 1880
rect 56555 1760 56560 1880
rect 56470 1740 56510 1745
rect 56470 1710 56475 1740
rect 56505 1710 56510 1740
rect 56470 1705 56510 1710
rect 56415 1695 56455 1700
rect 56415 1665 56420 1695
rect 56450 1665 56455 1695
rect 56415 1660 56455 1665
rect 56255 1280 56285 1285
rect 56305 1305 56345 1310
rect 56195 1270 56235 1275
rect 56305 1275 56310 1305
rect 56340 1275 56345 1305
rect 56475 1315 56505 1705
rect 56530 1700 56560 1760
rect 56585 1880 56615 1940
rect 56635 1930 56675 2355
rect 56775 2330 56780 2550
rect 56800 2330 56805 2550
rect 56775 2300 56805 2330
rect 56830 2550 56860 2580
rect 56830 2330 56835 2550
rect 56855 2330 56860 2550
rect 56830 2320 56860 2330
rect 56885 2550 56915 2560
rect 56885 2330 56890 2550
rect 56910 2330 56915 2550
rect 56885 2300 56915 2330
rect 56940 2550 56970 2580
rect 56940 2330 56945 2550
rect 56965 2330 56970 2550
rect 56940 2320 56970 2330
rect 56995 2550 57025 2560
rect 56995 2330 57000 2550
rect 57020 2330 57025 2550
rect 56995 2300 57025 2330
rect 57125 2470 57715 2475
rect 57125 2440 57130 2470
rect 57160 2440 57185 2470
rect 57215 2440 57240 2470
rect 57270 2440 57295 2470
rect 57325 2440 57350 2470
rect 57380 2440 57405 2470
rect 57435 2440 57460 2470
rect 57490 2440 57515 2470
rect 57545 2440 57570 2470
rect 57600 2440 57625 2470
rect 57655 2440 57680 2470
rect 57710 2440 57715 2470
rect 57125 2430 57715 2440
rect 57125 2400 57130 2430
rect 57160 2400 57185 2430
rect 57215 2400 57240 2430
rect 57270 2400 57295 2430
rect 57325 2400 57350 2430
rect 57380 2400 57405 2430
rect 57435 2400 57460 2430
rect 57490 2400 57515 2430
rect 57545 2400 57570 2430
rect 57600 2400 57625 2430
rect 57655 2400 57680 2430
rect 57710 2400 57715 2430
rect 57125 2390 57715 2400
rect 57125 2360 57130 2390
rect 57160 2360 57185 2390
rect 57215 2360 57240 2390
rect 57270 2360 57295 2390
rect 57325 2360 57350 2390
rect 57380 2360 57405 2390
rect 57435 2360 57460 2390
rect 57490 2360 57515 2390
rect 57545 2360 57570 2390
rect 57600 2360 57625 2390
rect 57655 2360 57680 2390
rect 57710 2360 57715 2390
rect 57125 2355 57715 2360
rect 56770 2295 56810 2300
rect 56770 2265 56775 2295
rect 56805 2265 56810 2295
rect 56770 2255 56810 2265
rect 56770 2225 56775 2255
rect 56805 2225 56810 2255
rect 56770 2215 56810 2225
rect 56770 2185 56775 2215
rect 56805 2185 56810 2215
rect 56770 2180 56810 2185
rect 56880 2295 56920 2300
rect 56880 2265 56885 2295
rect 56915 2265 56920 2295
rect 56880 2255 56920 2265
rect 56880 2225 56885 2255
rect 56915 2225 56920 2255
rect 56880 2215 56920 2225
rect 56880 2185 56885 2215
rect 56915 2185 56920 2215
rect 56880 2180 56920 2185
rect 56990 2295 57030 2300
rect 56990 2265 56995 2295
rect 57025 2265 57030 2295
rect 56990 2255 57030 2265
rect 56990 2225 56995 2255
rect 57025 2225 57030 2255
rect 56990 2215 57030 2225
rect 56990 2185 56995 2215
rect 57025 2185 57030 2215
rect 56990 2180 57030 2185
rect 56690 1985 56720 1990
rect 56690 1950 56720 1955
rect 57080 1985 57110 1990
rect 57080 1950 57110 1955
rect 56635 1900 56640 1930
rect 56670 1900 56675 1930
rect 56635 1895 56675 1900
rect 57125 1930 57165 2355
rect 57180 1975 57220 1980
rect 57180 1945 57185 1975
rect 57215 1945 57220 1975
rect 57180 1940 57220 1945
rect 57125 1900 57130 1930
rect 57160 1900 57165 1930
rect 57125 1895 57165 1900
rect 56585 1760 56590 1880
rect 56610 1760 56615 1880
rect 56585 1745 56615 1760
rect 56640 1880 56670 1895
rect 56640 1760 56645 1880
rect 56665 1760 56670 1880
rect 56580 1740 56620 1745
rect 56580 1710 56585 1740
rect 56615 1710 56620 1740
rect 56580 1705 56620 1710
rect 56525 1695 56565 1700
rect 56525 1665 56530 1695
rect 56560 1665 56565 1695
rect 56525 1660 56565 1665
rect 56365 1280 56395 1285
rect 56415 1305 56455 1310
rect 56305 1270 56345 1275
rect 56415 1275 56420 1305
rect 56450 1275 56455 1305
rect 56585 1315 56615 1705
rect 56640 1700 56670 1760
rect 56695 1880 56765 1890
rect 56695 1760 56700 1880
rect 56720 1760 56765 1880
rect 56695 1750 56765 1760
rect 57035 1880 57105 1890
rect 57035 1760 57080 1880
rect 57100 1760 57105 1880
rect 57035 1750 57105 1760
rect 56695 1720 56725 1750
rect 56695 1700 56700 1720
rect 56720 1700 56725 1720
rect 56635 1695 56675 1700
rect 56635 1665 56640 1695
rect 56670 1665 56675 1695
rect 56635 1660 56675 1665
rect 56695 1645 56725 1700
rect 57075 1720 57105 1750
rect 57075 1700 57080 1720
rect 57100 1700 57105 1720
rect 57130 1880 57160 1895
rect 57130 1760 57135 1880
rect 57155 1760 57160 1880
rect 57130 1700 57160 1760
rect 57185 1880 57215 1940
rect 57235 1930 57275 2355
rect 57290 1975 57330 1980
rect 57290 1945 57295 1975
rect 57325 1945 57330 1975
rect 57290 1940 57330 1945
rect 57235 1900 57240 1930
rect 57270 1900 57275 1930
rect 57235 1895 57275 1900
rect 57185 1760 57190 1880
rect 57210 1760 57215 1880
rect 57185 1745 57215 1760
rect 57240 1880 57270 1895
rect 57240 1760 57245 1880
rect 57265 1760 57270 1880
rect 57180 1740 57220 1745
rect 57180 1710 57185 1740
rect 57215 1710 57220 1740
rect 57180 1705 57220 1710
rect 57075 1645 57105 1700
rect 57125 1695 57165 1700
rect 57125 1665 57130 1695
rect 57160 1665 57165 1695
rect 57125 1660 57165 1665
rect 56690 1640 56730 1645
rect 56690 1610 56695 1640
rect 56725 1610 56730 1640
rect 56690 1600 56730 1610
rect 56690 1570 56695 1600
rect 56725 1570 56730 1600
rect 56690 1560 56730 1570
rect 56690 1530 56695 1560
rect 56725 1530 56730 1560
rect 56690 1525 56730 1530
rect 57070 1640 57110 1645
rect 57070 1610 57075 1640
rect 57105 1610 57110 1640
rect 57070 1600 57110 1610
rect 57070 1570 57075 1600
rect 57105 1570 57110 1600
rect 57070 1560 57110 1570
rect 57070 1530 57075 1560
rect 57105 1530 57110 1560
rect 57070 1525 57110 1530
rect 56880 1485 56920 1490
rect 56880 1455 56885 1485
rect 56915 1455 56920 1485
rect 56880 1445 56920 1455
rect 56880 1415 56885 1445
rect 56915 1415 56920 1445
rect 56880 1405 56920 1415
rect 56880 1375 56885 1405
rect 56915 1375 56920 1405
rect 56880 1370 56920 1375
rect 56475 1280 56505 1285
rect 56525 1305 56565 1310
rect 56415 1270 56455 1275
rect 56525 1275 56530 1305
rect 56560 1275 56565 1305
rect 56585 1280 56615 1285
rect 56635 1305 56675 1310
rect 56525 1270 56565 1275
rect 56635 1275 56640 1305
rect 56670 1275 56675 1305
rect 56635 1270 56675 1275
rect 56690 1305 56720 1310
rect 56690 1270 56720 1275
rect 56840 1305 56870 1310
rect 56840 1270 56870 1275
rect 56040 1260 56070 1265
rect 56035 1205 56065 1215
rect 56035 1085 56040 1205
rect 56060 1085 56065 1205
rect 56035 1075 56065 1085
rect 56090 1205 56120 1270
rect 56140 1260 56180 1265
rect 56140 1230 56145 1260
rect 56175 1230 56180 1260
rect 56140 1225 56180 1230
rect 56090 1085 56095 1205
rect 56115 1085 56120 1205
rect 56090 1070 56120 1085
rect 56145 1205 56175 1225
rect 56145 1085 56150 1205
rect 56170 1085 56175 1205
rect 56085 1065 56125 1070
rect 56035 1045 56065 1055
rect 56035 1025 56040 1045
rect 56060 1025 56065 1045
rect 56085 1035 56090 1065
rect 56120 1035 56125 1065
rect 56085 1030 56125 1035
rect 56035 1015 56065 1025
rect 56040 945 56060 1015
rect 56145 1000 56175 1085
rect 56200 1205 56230 1270
rect 56250 1260 56290 1265
rect 56250 1230 56255 1260
rect 56285 1230 56290 1260
rect 56250 1225 56290 1230
rect 56200 1085 56205 1205
rect 56225 1085 56230 1205
rect 56200 1070 56230 1085
rect 56255 1205 56285 1225
rect 56255 1085 56260 1205
rect 56280 1085 56285 1205
rect 56195 1065 56235 1070
rect 56195 1035 56200 1065
rect 56230 1035 56235 1065
rect 56195 1030 56235 1035
rect 56255 1000 56285 1085
rect 56310 1205 56340 1270
rect 56360 1260 56400 1265
rect 56360 1230 56365 1260
rect 56395 1230 56400 1260
rect 56360 1225 56400 1230
rect 56310 1085 56315 1205
rect 56335 1085 56340 1205
rect 56310 1070 56340 1085
rect 56365 1205 56395 1225
rect 56365 1085 56370 1205
rect 56390 1085 56395 1205
rect 56305 1065 56345 1070
rect 56305 1035 56310 1065
rect 56340 1035 56345 1065
rect 56305 1030 56345 1035
rect 56365 1000 56395 1085
rect 56420 1205 56450 1270
rect 56470 1260 56510 1265
rect 56470 1230 56475 1260
rect 56505 1230 56510 1260
rect 56470 1225 56510 1230
rect 56420 1085 56425 1205
rect 56445 1085 56450 1205
rect 56420 1070 56450 1085
rect 56475 1205 56505 1225
rect 56475 1085 56480 1205
rect 56500 1085 56505 1205
rect 56415 1065 56455 1070
rect 56415 1035 56420 1065
rect 56450 1035 56455 1065
rect 56415 1030 56455 1035
rect 56475 1000 56505 1085
rect 56530 1205 56560 1270
rect 56580 1260 56620 1265
rect 56580 1230 56585 1260
rect 56615 1230 56620 1260
rect 56580 1225 56620 1230
rect 56530 1085 56535 1205
rect 56555 1085 56560 1205
rect 56530 1070 56560 1085
rect 56585 1205 56615 1225
rect 56585 1085 56590 1205
rect 56610 1085 56615 1205
rect 56525 1065 56565 1070
rect 56525 1035 56530 1065
rect 56560 1035 56565 1065
rect 56525 1030 56565 1035
rect 56585 1000 56615 1085
rect 56640 1205 56670 1270
rect 56640 1085 56645 1205
rect 56665 1085 56670 1205
rect 56640 1070 56670 1085
rect 56695 1205 56805 1215
rect 56695 1085 56700 1205
rect 56720 1085 56780 1205
rect 56800 1085 56805 1205
rect 56695 1075 56805 1085
rect 56830 1205 56860 1215
rect 56830 1085 56835 1205
rect 56855 1085 56860 1205
rect 56635 1065 56675 1070
rect 56635 1035 56640 1065
rect 56670 1035 56675 1065
rect 56740 1055 56760 1075
rect 56830 1070 56860 1085
rect 56885 1205 56915 1370
rect 57185 1315 57215 1705
rect 57240 1700 57270 1760
rect 57295 1880 57325 1940
rect 57345 1930 57385 2355
rect 57400 1975 57440 1980
rect 57400 1945 57405 1975
rect 57435 1945 57440 1975
rect 57400 1940 57440 1945
rect 57345 1900 57350 1930
rect 57380 1900 57385 1930
rect 57345 1895 57385 1900
rect 57295 1760 57300 1880
rect 57320 1760 57325 1880
rect 57295 1745 57325 1760
rect 57350 1880 57380 1895
rect 57350 1760 57355 1880
rect 57375 1760 57380 1880
rect 57290 1740 57330 1745
rect 57290 1710 57295 1740
rect 57325 1710 57330 1740
rect 57290 1705 57330 1710
rect 57235 1695 57275 1700
rect 57235 1665 57240 1695
rect 57270 1665 57275 1695
rect 57235 1660 57275 1665
rect 56930 1305 56960 1310
rect 56930 1270 56960 1275
rect 57080 1305 57110 1310
rect 57080 1270 57110 1275
rect 57125 1305 57165 1310
rect 57125 1275 57130 1305
rect 57160 1275 57165 1305
rect 57295 1315 57325 1705
rect 57350 1700 57380 1760
rect 57405 1880 57435 1940
rect 57455 1930 57495 2355
rect 57510 1975 57550 1980
rect 57510 1945 57515 1975
rect 57545 1945 57550 1975
rect 57510 1940 57550 1945
rect 57455 1900 57460 1930
rect 57490 1900 57495 1930
rect 57455 1895 57495 1900
rect 57405 1760 57410 1880
rect 57430 1760 57435 1880
rect 57405 1745 57435 1760
rect 57460 1880 57490 1895
rect 57460 1760 57465 1880
rect 57485 1760 57490 1880
rect 57400 1740 57440 1745
rect 57400 1710 57405 1740
rect 57435 1710 57440 1740
rect 57400 1705 57440 1710
rect 57345 1695 57385 1700
rect 57345 1665 57350 1695
rect 57380 1665 57385 1695
rect 57345 1660 57385 1665
rect 57185 1280 57215 1285
rect 57235 1305 57275 1310
rect 57125 1270 57165 1275
rect 57235 1275 57240 1305
rect 57270 1275 57275 1305
rect 57405 1315 57435 1705
rect 57460 1700 57490 1760
rect 57515 1880 57545 1940
rect 57565 1930 57605 2355
rect 57620 1975 57660 1980
rect 57620 1945 57625 1975
rect 57655 1945 57660 1975
rect 57620 1940 57660 1945
rect 57565 1900 57570 1930
rect 57600 1900 57605 1930
rect 57565 1895 57605 1900
rect 57515 1760 57520 1880
rect 57540 1760 57545 1880
rect 57515 1745 57545 1760
rect 57570 1880 57600 1895
rect 57570 1760 57575 1880
rect 57595 1760 57600 1880
rect 57510 1740 57550 1745
rect 57510 1710 57515 1740
rect 57545 1710 57550 1740
rect 57510 1705 57550 1710
rect 57455 1695 57495 1700
rect 57455 1665 57460 1695
rect 57490 1665 57495 1695
rect 57455 1660 57495 1665
rect 57295 1280 57325 1285
rect 57345 1305 57385 1310
rect 57235 1270 57275 1275
rect 57345 1275 57350 1305
rect 57380 1275 57385 1305
rect 57515 1315 57545 1705
rect 57570 1700 57600 1760
rect 57625 1880 57655 1940
rect 57675 1930 57715 2355
rect 57730 1985 57760 1990
rect 57730 1950 57760 1955
rect 57675 1900 57680 1930
rect 57710 1900 57715 1930
rect 57675 1895 57715 1900
rect 57625 1760 57630 1880
rect 57650 1760 57655 1880
rect 57625 1745 57655 1760
rect 57680 1880 57710 1895
rect 57680 1760 57685 1880
rect 57705 1760 57710 1880
rect 57620 1740 57660 1745
rect 57620 1710 57625 1740
rect 57655 1710 57660 1740
rect 57620 1705 57660 1710
rect 57565 1695 57605 1700
rect 57565 1665 57570 1695
rect 57600 1665 57605 1695
rect 57565 1660 57605 1665
rect 57405 1280 57435 1285
rect 57455 1305 57495 1310
rect 57345 1270 57385 1275
rect 57455 1275 57460 1305
rect 57490 1275 57495 1305
rect 57625 1315 57655 1705
rect 57680 1700 57710 1760
rect 57735 1880 57765 1890
rect 57735 1760 57740 1880
rect 57760 1760 57765 1880
rect 57735 1750 57765 1760
rect 57735 1720 57765 1730
rect 57735 1700 57740 1720
rect 57760 1700 57765 1720
rect 57675 1695 57715 1700
rect 57675 1665 57680 1695
rect 57710 1665 57715 1695
rect 57675 1660 57715 1665
rect 57735 1645 57765 1700
rect 57730 1640 57770 1645
rect 57730 1610 57735 1640
rect 57765 1610 57770 1640
rect 57730 1600 57770 1610
rect 57730 1570 57735 1600
rect 57765 1570 57770 1600
rect 57730 1560 57770 1570
rect 57730 1530 57735 1560
rect 57765 1530 57770 1560
rect 57730 1525 57770 1530
rect 57515 1280 57545 1285
rect 57565 1305 57605 1310
rect 57455 1270 57495 1275
rect 57565 1275 57570 1305
rect 57600 1275 57605 1305
rect 57625 1280 57655 1285
rect 57675 1305 57715 1310
rect 57565 1270 57605 1275
rect 57675 1275 57680 1305
rect 57710 1275 57715 1305
rect 57675 1270 57715 1275
rect 57730 1295 57760 1300
rect 56885 1085 56890 1205
rect 56910 1085 56915 1205
rect 56885 1075 56915 1085
rect 56940 1205 56970 1215
rect 56940 1085 56945 1205
rect 56965 1085 56970 1205
rect 56940 1070 56970 1085
rect 56995 1205 57105 1215
rect 56995 1085 57000 1205
rect 57020 1085 57080 1205
rect 57100 1085 57105 1205
rect 56995 1075 57105 1085
rect 57130 1205 57160 1270
rect 57180 1260 57220 1265
rect 57180 1230 57185 1260
rect 57215 1230 57220 1260
rect 57180 1225 57220 1230
rect 57130 1085 57135 1205
rect 57155 1085 57160 1205
rect 56825 1065 56865 1070
rect 56635 1030 56675 1035
rect 56735 1045 56765 1055
rect 56735 1025 56740 1045
rect 56760 1025 56765 1045
rect 56735 1015 56765 1025
rect 56825 1035 56830 1065
rect 56860 1035 56865 1065
rect 56140 995 56180 1000
rect 56140 965 56145 995
rect 56175 965 56180 995
rect 56140 960 56180 965
rect 56250 995 56290 1000
rect 56250 965 56255 995
rect 56285 965 56290 995
rect 56250 960 56290 965
rect 56360 995 56400 1000
rect 56360 965 56365 995
rect 56395 965 56400 995
rect 56360 960 56400 965
rect 56440 995 56700 1000
rect 56440 965 56475 995
rect 56505 965 56585 995
rect 56615 965 56700 995
rect 56030 940 56070 945
rect 56030 910 56035 940
rect 56065 910 56070 940
rect 56030 900 56070 910
rect 56030 870 56035 900
rect 56065 870 56070 900
rect 56030 860 56070 870
rect 56030 830 56035 860
rect 56065 830 56070 860
rect 56030 825 56070 830
rect 55940 805 55980 810
rect 55940 775 55945 805
rect 55975 775 55980 805
rect 55940 770 55980 775
rect 56440 480 56700 965
rect 56740 945 56760 1015
rect 56730 940 56770 945
rect 56730 910 56735 940
rect 56765 910 56770 940
rect 56730 900 56770 910
rect 56730 870 56735 900
rect 56765 870 56770 900
rect 56730 860 56770 870
rect 56730 830 56735 860
rect 56765 830 56770 860
rect 56730 825 56770 830
rect 56440 450 56445 480
rect 56475 450 56555 480
rect 56585 450 56665 480
rect 56695 450 56700 480
rect 56440 445 56700 450
rect 56770 480 56810 485
rect 56770 450 56775 480
rect 56805 450 56810 480
rect 56770 445 56810 450
rect 56825 465 56865 1035
rect 56935 1065 56975 1070
rect 56935 1035 56940 1065
rect 56970 1035 56975 1065
rect 57040 1055 57060 1075
rect 57130 1070 57160 1085
rect 57185 1205 57215 1225
rect 57185 1085 57190 1205
rect 57210 1085 57215 1205
rect 57125 1065 57165 1070
rect 56825 445 56835 465
rect 56855 445 56865 465
rect 56880 480 56920 485
rect 56880 450 56885 480
rect 56915 450 56920 480
rect 56880 445 56920 450
rect 56935 465 56975 1035
rect 57035 1045 57065 1055
rect 57035 1025 57040 1045
rect 57060 1025 57065 1045
rect 57125 1035 57130 1065
rect 57160 1035 57165 1065
rect 57125 1030 57165 1035
rect 57035 1015 57065 1025
rect 57040 945 57060 1015
rect 57185 1000 57215 1085
rect 57240 1205 57270 1270
rect 57290 1260 57330 1265
rect 57290 1230 57295 1260
rect 57325 1230 57330 1260
rect 57290 1225 57330 1230
rect 57240 1085 57245 1205
rect 57265 1085 57270 1205
rect 57240 1070 57270 1085
rect 57295 1205 57325 1225
rect 57295 1085 57300 1205
rect 57320 1085 57325 1205
rect 57235 1065 57275 1070
rect 57235 1035 57240 1065
rect 57270 1035 57275 1065
rect 57235 1030 57275 1035
rect 57295 1000 57325 1085
rect 57350 1205 57380 1270
rect 57400 1260 57440 1265
rect 57400 1230 57405 1260
rect 57435 1230 57440 1260
rect 57400 1225 57440 1230
rect 57350 1085 57355 1205
rect 57375 1085 57380 1205
rect 57350 1070 57380 1085
rect 57405 1205 57435 1225
rect 57405 1085 57410 1205
rect 57430 1085 57435 1205
rect 57345 1065 57385 1070
rect 57345 1035 57350 1065
rect 57380 1035 57385 1065
rect 57345 1030 57385 1035
rect 57405 1000 57435 1085
rect 57460 1205 57490 1270
rect 57510 1260 57550 1265
rect 57510 1230 57515 1260
rect 57545 1230 57550 1260
rect 57510 1225 57550 1230
rect 57460 1085 57465 1205
rect 57485 1085 57490 1205
rect 57460 1070 57490 1085
rect 57515 1205 57545 1225
rect 57515 1085 57520 1205
rect 57540 1085 57545 1205
rect 57455 1065 57495 1070
rect 57455 1035 57460 1065
rect 57490 1035 57495 1065
rect 57455 1030 57495 1035
rect 57515 1000 57545 1085
rect 57570 1205 57600 1270
rect 57620 1260 57660 1265
rect 57620 1230 57625 1260
rect 57655 1230 57660 1260
rect 57620 1225 57660 1230
rect 57570 1085 57575 1205
rect 57595 1085 57600 1205
rect 57570 1070 57600 1085
rect 57625 1205 57655 1225
rect 57625 1085 57630 1205
rect 57650 1085 57655 1205
rect 57565 1065 57605 1070
rect 57565 1035 57570 1065
rect 57600 1035 57605 1065
rect 57565 1030 57605 1035
rect 57625 1000 57655 1085
rect 57680 1205 57710 1270
rect 57730 1260 57760 1265
rect 57680 1085 57685 1205
rect 57705 1085 57710 1205
rect 57680 1070 57710 1085
rect 57735 1205 57765 1215
rect 57735 1085 57740 1205
rect 57760 1085 57765 1205
rect 57735 1075 57765 1085
rect 57675 1065 57715 1070
rect 57675 1035 57680 1065
rect 57710 1035 57715 1065
rect 57675 1030 57715 1035
rect 57735 1045 57765 1055
rect 57735 1025 57740 1045
rect 57760 1025 57765 1045
rect 57735 1015 57765 1025
rect 57100 995 57360 1000
rect 57100 965 57185 995
rect 57215 965 57295 995
rect 57325 965 57360 995
rect 57030 940 57070 945
rect 57030 910 57035 940
rect 57065 910 57070 940
rect 57030 900 57070 910
rect 57030 870 57035 900
rect 57065 870 57070 900
rect 57030 860 57070 870
rect 57030 830 57035 860
rect 57065 830 57070 860
rect 57030 825 57070 830
rect 56935 445 56945 465
rect 56965 445 56975 465
rect 56990 480 57030 485
rect 56990 450 56995 480
rect 57025 450 57030 480
rect 56990 445 57030 450
rect 57100 480 57360 965
rect 57400 995 57440 1000
rect 57400 965 57405 995
rect 57435 965 57440 995
rect 57400 960 57440 965
rect 57510 995 57550 1000
rect 57510 965 57515 995
rect 57545 965 57550 995
rect 57510 960 57550 965
rect 57620 995 57660 1000
rect 57620 965 57625 995
rect 57655 965 57660 995
rect 57620 960 57660 965
rect 57740 945 57760 1015
rect 57730 940 57770 945
rect 57730 910 57735 940
rect 57765 910 57770 940
rect 57730 900 57770 910
rect 57730 870 57735 900
rect 57765 870 57770 900
rect 57730 860 57770 870
rect 57730 830 57735 860
rect 57765 830 57770 860
rect 57730 825 57770 830
rect 57830 810 57850 2745
rect 57865 2670 57905 2675
rect 57865 2640 57870 2670
rect 57900 2640 57905 2670
rect 57865 2635 57905 2640
rect 57820 805 57860 810
rect 57820 775 57825 805
rect 57855 775 57860 805
rect 57820 770 57860 775
rect 57100 450 57105 480
rect 57135 450 57215 480
rect 57245 450 57325 480
rect 57355 450 57360 480
rect 57100 445 57360 450
rect 57430 480 57470 485
rect 57430 450 57435 480
rect 57465 450 57470 480
rect 57430 445 57470 450
rect 56185 405 56255 415
rect 56185 185 56230 405
rect 56250 185 56255 405
rect 56185 175 56255 185
rect 56225 155 56255 175
rect 56280 405 56310 415
rect 56280 185 56285 405
rect 56305 185 56310 405
rect 56280 155 56310 185
rect 56335 405 56365 415
rect 56335 185 56340 405
rect 56360 185 56365 405
rect 56220 150 56260 155
rect 56220 120 56225 150
rect 56255 120 56260 150
rect 55885 -250 55925 -245
rect 55885 -280 55890 -250
rect 55920 -280 55925 -250
rect 55885 -285 55925 -280
rect 55150 -365 55190 -360
rect 55150 -395 55155 -365
rect 55185 -395 55190 -365
rect 55150 -400 55190 -395
rect 55255 -385 55285 -345
rect 55255 -405 55260 -385
rect 55280 -405 55285 -385
rect 55255 -575 55285 -405
rect 56220 -575 56260 120
rect 56275 150 56315 155
rect 56275 120 56280 150
rect 56310 120 56315 150
rect 56275 115 56315 120
rect 56335 -55 56365 185
rect 56390 405 56420 415
rect 56390 185 56395 405
rect 56415 185 56420 405
rect 56390 155 56420 185
rect 56445 405 56475 445
rect 56445 185 56450 405
rect 56470 185 56475 405
rect 56385 150 56425 155
rect 56385 120 56390 150
rect 56420 120 56425 150
rect 56385 115 56425 120
rect 56445 100 56475 185
rect 56500 405 56530 415
rect 56500 185 56505 405
rect 56525 185 56530 405
rect 56500 155 56530 185
rect 56555 405 56585 445
rect 56555 185 56560 405
rect 56580 185 56585 405
rect 56495 150 56535 155
rect 56495 120 56500 150
rect 56530 120 56535 150
rect 56495 115 56535 120
rect 56555 100 56585 185
rect 56610 405 56640 415
rect 56610 185 56615 405
rect 56635 185 56640 405
rect 56610 155 56640 185
rect 56665 405 56695 445
rect 56665 185 56670 405
rect 56690 185 56695 405
rect 56605 150 56645 155
rect 56605 120 56610 150
rect 56640 120 56645 150
rect 56605 115 56645 120
rect 56665 100 56695 185
rect 56720 405 56750 415
rect 56720 185 56725 405
rect 56745 185 56750 405
rect 56720 155 56750 185
rect 56775 405 56805 445
rect 56825 435 56865 445
rect 56775 185 56780 405
rect 56800 185 56805 405
rect 56715 150 56755 155
rect 56715 120 56720 150
rect 56750 120 56755 150
rect 56715 115 56755 120
rect 56775 100 56805 185
rect 56830 405 56860 415
rect 56830 185 56835 405
rect 56855 185 56860 405
rect 56830 155 56860 185
rect 56885 405 56915 445
rect 56935 435 56975 445
rect 56885 185 56890 405
rect 56910 185 56915 405
rect 56825 150 56865 155
rect 56825 120 56830 150
rect 56860 120 56865 150
rect 56825 115 56865 120
rect 56885 100 56915 185
rect 56940 405 56970 415
rect 56940 185 56945 405
rect 56965 185 56970 405
rect 56940 155 56970 185
rect 56995 405 57025 445
rect 56995 185 57000 405
rect 57020 185 57025 405
rect 56935 150 56975 155
rect 56935 120 56940 150
rect 56970 120 56975 150
rect 56935 115 56975 120
rect 56995 100 57025 185
rect 57050 405 57080 415
rect 57050 185 57055 405
rect 57075 185 57080 405
rect 57050 155 57080 185
rect 57105 405 57135 445
rect 57105 185 57110 405
rect 57130 185 57135 405
rect 57045 150 57085 155
rect 57045 120 57050 150
rect 57080 120 57085 150
rect 57045 115 57085 120
rect 57105 100 57135 185
rect 57160 405 57190 415
rect 57160 185 57165 405
rect 57185 185 57190 405
rect 57160 155 57190 185
rect 57215 405 57245 445
rect 57215 185 57220 405
rect 57240 185 57245 405
rect 57155 150 57195 155
rect 57155 120 57160 150
rect 57190 120 57195 150
rect 57155 115 57195 120
rect 57215 100 57245 185
rect 57270 405 57300 415
rect 57270 185 57275 405
rect 57295 185 57300 405
rect 57270 155 57300 185
rect 57325 405 57355 445
rect 57325 185 57330 405
rect 57350 185 57355 405
rect 57265 150 57305 155
rect 57265 120 57270 150
rect 57300 120 57305 150
rect 57265 115 57305 120
rect 57325 100 57355 185
rect 57380 405 57410 415
rect 57380 185 57385 405
rect 57405 185 57410 405
rect 57380 155 57410 185
rect 57435 405 57465 445
rect 57435 185 57440 405
rect 57460 185 57465 405
rect 57375 150 57415 155
rect 57375 120 57380 150
rect 57410 120 57415 150
rect 57375 115 57415 120
rect 57435 100 57465 185
rect 57490 405 57520 415
rect 57490 185 57495 405
rect 57515 185 57520 405
rect 57490 155 57520 185
rect 57485 150 57525 155
rect 57485 120 57490 150
rect 57520 120 57525 150
rect 56440 95 56480 100
rect 56440 65 56445 95
rect 56475 65 56480 95
rect 56440 60 56480 65
rect 56550 95 56590 100
rect 56550 65 56555 95
rect 56585 65 56590 95
rect 56550 60 56590 65
rect 56660 95 56700 100
rect 56660 65 56665 95
rect 56695 65 56700 95
rect 56660 60 56700 65
rect 56770 95 56810 100
rect 56770 65 56775 95
rect 56805 65 56810 95
rect 56770 60 56810 65
rect 56880 95 56920 100
rect 56880 65 56885 95
rect 56915 65 56920 95
rect 56880 60 56920 65
rect 56990 95 57030 100
rect 56990 65 56995 95
rect 57025 65 57030 95
rect 56990 60 57030 65
rect 57100 95 57140 100
rect 57100 65 57105 95
rect 57135 65 57140 95
rect 57100 60 57140 65
rect 57210 95 57250 100
rect 57210 65 57215 95
rect 57245 65 57250 95
rect 57210 60 57250 65
rect 57320 95 57360 100
rect 57320 65 57325 95
rect 57355 65 57360 95
rect 57320 60 57360 65
rect 57430 95 57470 100
rect 57430 65 57435 95
rect 57465 65 57470 95
rect 57430 60 57470 65
rect 56330 -60 56370 -55
rect 56330 -90 56335 -60
rect 56365 -90 56370 -60
rect 56330 -100 56370 -90
rect 56330 -130 56335 -100
rect 56365 -130 56370 -100
rect 56330 -140 56370 -130
rect 56330 -170 56335 -140
rect 56365 -170 56370 -140
rect 56330 -175 56370 -170
rect 56540 -195 56580 -190
rect 56540 -225 56545 -195
rect 56575 -225 56580 -195
rect 56540 -230 56580 -225
rect 56650 -195 56690 -190
rect 56650 -225 56655 -195
rect 56685 -225 56690 -195
rect 56650 -230 56690 -225
rect 56870 -195 56910 -190
rect 56870 -225 56875 -195
rect 56905 -225 56910 -195
rect 56870 -230 56910 -225
rect 56485 -250 56525 -245
rect 56485 -280 56490 -250
rect 56520 -280 56525 -250
rect 56485 -285 56525 -280
rect 56395 -315 56465 -305
rect 56395 -435 56440 -315
rect 56460 -435 56465 -315
rect 56395 -445 56465 -435
rect 56435 -475 56465 -445
rect 56490 -315 56520 -285
rect 56490 -435 56495 -315
rect 56515 -435 56520 -315
rect 56490 -465 56520 -435
rect 56545 -315 56575 -230
rect 56595 -250 56635 -245
rect 56595 -280 56600 -250
rect 56630 -280 56635 -250
rect 56595 -285 56635 -280
rect 56545 -435 56550 -315
rect 56570 -435 56575 -315
rect 56435 -495 56440 -475
rect 56460 -495 56465 -475
rect 56435 -575 56465 -495
rect 56485 -470 56525 -465
rect 56485 -500 56490 -470
rect 56520 -500 56525 -470
rect 56485 -505 56525 -500
rect 56545 -520 56575 -435
rect 56600 -315 56630 -285
rect 56600 -435 56605 -315
rect 56625 -435 56630 -315
rect 56600 -465 56630 -435
rect 56655 -315 56685 -230
rect 56705 -250 56745 -245
rect 56705 -280 56710 -250
rect 56740 -280 56745 -250
rect 56705 -285 56745 -280
rect 56655 -435 56660 -315
rect 56680 -435 56685 -315
rect 56595 -470 56635 -465
rect 56595 -500 56600 -470
rect 56630 -500 56635 -470
rect 56595 -505 56635 -500
rect 56655 -520 56685 -435
rect 56710 -315 56740 -285
rect 56710 -435 56715 -315
rect 56735 -435 56740 -315
rect 56710 -465 56740 -435
rect 56765 -315 56835 -305
rect 56765 -435 56770 -315
rect 56790 -435 56835 -315
rect 56765 -445 56835 -435
rect 56875 -315 56905 -230
rect 56920 -250 56960 -245
rect 56920 -280 56925 -250
rect 56955 -280 56960 -250
rect 56920 -285 56960 -280
rect 57040 -250 57080 -245
rect 57040 -280 57045 -250
rect 57075 -280 57080 -250
rect 57040 -285 57080 -280
rect 57160 -250 57200 -245
rect 57160 -280 57165 -250
rect 57195 -280 57200 -250
rect 57160 -285 57200 -280
rect 56875 -435 56880 -315
rect 56900 -435 56905 -315
rect 56705 -470 56745 -465
rect 56705 -500 56710 -470
rect 56740 -500 56745 -470
rect 56705 -505 56745 -500
rect 56765 -475 56795 -445
rect 56765 -495 56770 -475
rect 56790 -495 56795 -475
rect 56540 -525 56580 -520
rect 56540 -555 56545 -525
rect 56575 -555 56580 -525
rect 56540 -560 56580 -555
rect 56650 -525 56690 -520
rect 56650 -555 56655 -525
rect 56685 -555 56690 -525
rect 56650 -560 56690 -555
rect 56765 -575 56795 -495
rect 56875 -520 56905 -435
rect 57215 -325 57245 60
rect 57415 40 57455 45
rect 57415 10 57420 40
rect 57450 10 57455 40
rect 57415 5 57455 10
rect 57215 -425 57220 -325
rect 57240 -425 57245 -325
rect 57215 -445 57245 -425
rect 56920 -470 56960 -465
rect 56920 -500 56925 -470
rect 56955 -500 56960 -470
rect 56920 -505 56960 -500
rect 57040 -470 57080 -465
rect 57040 -500 57045 -470
rect 57075 -500 57080 -470
rect 57040 -505 57080 -500
rect 57160 -470 57200 -465
rect 57160 -500 57165 -470
rect 57195 -500 57200 -470
rect 57160 -505 57200 -500
rect 56870 -525 56910 -520
rect 56870 -555 56875 -525
rect 56905 -555 56910 -525
rect 56870 -560 56910 -555
rect 55055 -580 55210 -575
rect 55055 -610 55095 -580
rect 55125 -610 55135 -580
rect 55165 -610 55175 -580
rect 55205 -610 55210 -580
rect 55055 -620 55210 -610
rect 55055 -650 55095 -620
rect 55125 -650 55135 -620
rect 55165 -650 55175 -620
rect 55205 -650 55210 -620
rect 55055 -660 55210 -650
rect 55055 -690 55095 -660
rect 55125 -690 55135 -660
rect 55165 -690 55175 -660
rect 55205 -690 55210 -660
rect 55055 -695 55210 -690
rect 55250 -580 55290 -575
rect 55250 -610 55255 -580
rect 55285 -610 55290 -580
rect 55250 -620 55290 -610
rect 55250 -650 55255 -620
rect 55285 -650 55290 -620
rect 55250 -660 55290 -650
rect 55250 -690 55255 -660
rect 55285 -690 55290 -660
rect 55250 -695 55290 -690
rect 55440 -580 55560 -575
rect 55440 -610 55445 -580
rect 55475 -610 55485 -580
rect 55515 -610 55525 -580
rect 55555 -610 55560 -580
rect 55440 -620 55560 -610
rect 55440 -650 55445 -620
rect 55475 -650 55485 -620
rect 55515 -650 55525 -620
rect 55555 -650 55560 -620
rect 55440 -660 55560 -650
rect 55440 -690 55445 -660
rect 55475 -690 55485 -660
rect 55515 -690 55525 -660
rect 55555 -690 55560 -660
rect 54740 -1500 54860 -695
rect 55090 -1500 55210 -695
rect 55440 -1500 55560 -690
rect 55790 -580 55910 -575
rect 55790 -610 55795 -580
rect 55825 -610 55835 -580
rect 55865 -610 55875 -580
rect 55905 -610 55910 -580
rect 55790 -620 55910 -610
rect 55790 -650 55795 -620
rect 55825 -650 55835 -620
rect 55865 -650 55875 -620
rect 55905 -650 55910 -620
rect 55790 -660 55910 -650
rect 55790 -690 55795 -660
rect 55825 -690 55835 -660
rect 55865 -690 55875 -660
rect 55905 -690 55910 -660
rect 55790 -1500 55910 -690
rect 56140 -580 56260 -575
rect 56140 -610 56145 -580
rect 56175 -610 56185 -580
rect 56215 -610 56225 -580
rect 56255 -610 56260 -580
rect 56140 -620 56260 -610
rect 56140 -650 56145 -620
rect 56175 -650 56185 -620
rect 56215 -650 56225 -620
rect 56255 -650 56260 -620
rect 56140 -660 56260 -650
rect 56140 -690 56145 -660
rect 56175 -690 56185 -660
rect 56215 -690 56225 -660
rect 56255 -690 56260 -660
rect 56140 -1500 56260 -690
rect 56430 -580 56470 -575
rect 56430 -610 56435 -580
rect 56465 -610 56470 -580
rect 56430 -620 56470 -610
rect 56430 -650 56435 -620
rect 56465 -650 56470 -620
rect 56430 -660 56470 -650
rect 56430 -690 56435 -660
rect 56465 -690 56470 -660
rect 56430 -695 56470 -690
rect 56490 -580 56610 -575
rect 56490 -610 56495 -580
rect 56525 -610 56535 -580
rect 56565 -610 56575 -580
rect 56605 -610 56610 -580
rect 56490 -620 56610 -610
rect 56490 -650 56495 -620
rect 56525 -650 56535 -620
rect 56565 -650 56575 -620
rect 56605 -650 56610 -620
rect 56490 -660 56610 -650
rect 56490 -690 56495 -660
rect 56525 -690 56535 -660
rect 56565 -690 56575 -660
rect 56605 -690 56610 -660
rect 56490 -1500 56610 -690
rect 56760 -580 56800 -575
rect 56760 -610 56765 -580
rect 56795 -610 56800 -580
rect 56760 -620 56800 -610
rect 56760 -650 56765 -620
rect 56795 -650 56800 -620
rect 56760 -660 56800 -650
rect 56760 -690 56765 -660
rect 56795 -690 56800 -660
rect 56760 -695 56800 -690
rect 56840 -580 56960 -575
rect 56840 -610 56845 -580
rect 56875 -610 56885 -580
rect 56915 -610 56925 -580
rect 56955 -610 56960 -580
rect 56840 -620 56960 -610
rect 56840 -650 56845 -620
rect 56875 -650 56885 -620
rect 56915 -650 56925 -620
rect 56955 -650 56960 -620
rect 56840 -660 56960 -650
rect 56840 -690 56845 -660
rect 56875 -690 56885 -660
rect 56915 -690 56925 -660
rect 56955 -690 56960 -660
rect 56840 -1500 56960 -690
rect 57190 -580 57310 -575
rect 57190 -610 57195 -580
rect 57225 -610 57235 -580
rect 57265 -610 57275 -580
rect 57305 -610 57310 -580
rect 57190 -620 57310 -610
rect 57190 -650 57195 -620
rect 57225 -650 57235 -620
rect 57265 -650 57275 -620
rect 57305 -650 57310 -620
rect 57190 -660 57310 -650
rect 57190 -690 57195 -660
rect 57225 -690 57235 -660
rect 57265 -690 57275 -660
rect 57305 -690 57310 -660
rect 57190 -1500 57310 -690
rect 57485 -580 57525 120
rect 57875 45 57895 2635
rect 58010 2295 58130 2300
rect 58010 2265 58015 2295
rect 58045 2265 58055 2295
rect 58085 2265 58095 2295
rect 58125 2265 58130 2295
rect 58010 2255 58130 2265
rect 58010 2225 58015 2255
rect 58045 2225 58055 2255
rect 58085 2225 58095 2255
rect 58125 2225 58130 2255
rect 58010 2215 58130 2225
rect 58010 2185 58015 2215
rect 58045 2185 58055 2215
rect 58085 2185 58095 2215
rect 58125 2185 58130 2215
rect 58010 2050 58130 2185
rect 58010 2020 58015 2050
rect 58045 2020 58055 2050
rect 58085 2020 58095 2050
rect 58125 2020 58130 2050
rect 58010 2010 58130 2020
rect 58010 1980 58015 2010
rect 58045 1980 58055 2010
rect 58085 1980 58095 2010
rect 58125 1980 58130 2010
rect 58010 1970 58130 1980
rect 58010 1940 58015 1970
rect 58045 1940 58055 1970
rect 58085 1940 58095 1970
rect 58125 1940 58130 1970
rect 58010 1640 58130 1940
rect 58010 1610 58015 1640
rect 58045 1610 58055 1640
rect 58085 1610 58095 1640
rect 58125 1610 58130 1640
rect 58010 1600 58130 1610
rect 58010 1570 58015 1600
rect 58045 1570 58055 1600
rect 58085 1570 58095 1600
rect 58125 1570 58130 1600
rect 58010 1560 58130 1570
rect 58010 1530 58015 1560
rect 58045 1530 58055 1560
rect 58085 1530 58095 1560
rect 58125 1530 58130 1560
rect 58010 1525 58130 1530
rect 58145 2185 58265 3245
rect 58145 2155 58150 2185
rect 58180 2155 58190 2185
rect 58220 2155 58230 2185
rect 58260 2155 58265 2185
rect 58145 2145 58265 2155
rect 58145 2115 58150 2145
rect 58180 2115 58190 2145
rect 58220 2115 58230 2145
rect 58260 2115 58265 2145
rect 58145 2105 58265 2115
rect 58145 2075 58150 2105
rect 58180 2075 58190 2105
rect 58220 2075 58230 2105
rect 58260 2075 58265 2105
rect 58010 1485 58130 1490
rect 58010 1455 58015 1485
rect 58045 1455 58055 1485
rect 58085 1455 58095 1485
rect 58125 1455 58130 1485
rect 58010 1445 58130 1455
rect 58010 1415 58015 1445
rect 58045 1415 58055 1445
rect 58085 1415 58095 1445
rect 58125 1415 58130 1445
rect 58010 1405 58130 1415
rect 58010 1375 58015 1405
rect 58045 1375 58055 1405
rect 58085 1375 58095 1405
rect 58125 1375 58130 1405
rect 57865 40 57905 45
rect 57865 10 57870 40
rect 57900 10 57905 40
rect 57865 5 57905 10
rect 58010 -60 58130 1375
rect 58145 1080 58265 2075
rect 58280 3490 58400 3495
rect 58280 3460 58285 3490
rect 58315 3460 58325 3490
rect 58355 3460 58365 3490
rect 58395 3460 58400 3490
rect 58280 3450 58400 3460
rect 58280 3420 58285 3450
rect 58315 3420 58325 3450
rect 58355 3420 58365 3450
rect 58395 3420 58400 3450
rect 58280 3410 58400 3420
rect 58280 3380 58285 3410
rect 58315 3380 58325 3410
rect 58355 3380 58365 3410
rect 58395 3380 58400 3410
rect 58280 2470 58400 3380
rect 59505 3375 59545 3380
rect 58480 3355 58520 3360
rect 58480 3325 58485 3355
rect 58515 3325 58520 3355
rect 58480 3315 58520 3325
rect 58480 3285 58485 3315
rect 58515 3285 58520 3315
rect 58480 3275 58520 3285
rect 58480 3245 58485 3275
rect 58515 3245 58520 3275
rect 58480 3240 58520 3245
rect 58590 3355 58630 3360
rect 58590 3325 58595 3355
rect 58625 3325 58630 3355
rect 58590 3315 58630 3325
rect 58590 3285 58595 3315
rect 58625 3285 58630 3315
rect 58590 3275 58630 3285
rect 58590 3245 58595 3275
rect 58625 3245 58630 3275
rect 58590 3240 58630 3245
rect 58700 3355 58740 3360
rect 58700 3325 58705 3355
rect 58735 3325 58740 3355
rect 58700 3315 58740 3325
rect 58700 3285 58705 3315
rect 58735 3285 58740 3315
rect 58700 3275 58740 3285
rect 58700 3245 58705 3275
rect 58735 3245 58740 3275
rect 58700 3240 58740 3245
rect 58810 3355 58850 3360
rect 58810 3325 58815 3355
rect 58845 3325 58850 3355
rect 58810 3315 58850 3325
rect 58810 3285 58815 3315
rect 58845 3285 58850 3315
rect 58810 3275 58850 3285
rect 58810 3245 58815 3275
rect 58845 3245 58850 3275
rect 58810 3240 58850 3245
rect 58920 3355 58960 3360
rect 58920 3325 58925 3355
rect 58955 3325 58960 3355
rect 58920 3315 58960 3325
rect 58920 3285 58925 3315
rect 58955 3285 58960 3315
rect 58920 3275 58960 3285
rect 58920 3245 58925 3275
rect 58955 3245 58960 3275
rect 58920 3240 58960 3245
rect 59030 3355 59070 3360
rect 59030 3325 59035 3355
rect 59065 3325 59070 3355
rect 59030 3315 59070 3325
rect 59030 3285 59035 3315
rect 59065 3285 59070 3315
rect 59030 3275 59070 3285
rect 59030 3245 59035 3275
rect 59065 3245 59070 3275
rect 59030 3240 59070 3245
rect 59140 3355 59180 3360
rect 59140 3325 59145 3355
rect 59175 3325 59180 3355
rect 59140 3315 59180 3325
rect 59140 3285 59145 3315
rect 59175 3285 59180 3315
rect 59140 3275 59180 3285
rect 59140 3245 59145 3275
rect 59175 3245 59180 3275
rect 59140 3240 59180 3245
rect 59505 3345 59510 3375
rect 59540 3345 59545 3375
rect 58485 3200 58515 3240
rect 58485 3180 58490 3200
rect 58510 3180 58515 3200
rect 58485 3140 58515 3180
rect 58535 3190 58575 3195
rect 58535 3160 58540 3190
rect 58570 3160 58575 3190
rect 58535 3155 58575 3160
rect 58485 2570 58490 3140
rect 58510 2570 58515 3140
rect 58485 2560 58515 2570
rect 58540 3140 58570 3155
rect 58540 2570 58545 3140
rect 58565 2570 58570 3140
rect 58540 2555 58570 2570
rect 58595 3140 58625 3240
rect 58645 3190 58685 3195
rect 58645 3160 58650 3190
rect 58680 3160 58685 3190
rect 58645 3155 58685 3160
rect 58595 2570 58600 3140
rect 58620 2570 58625 3140
rect 58595 2560 58625 2570
rect 58650 3140 58680 3155
rect 58650 2570 58655 3140
rect 58675 2570 58680 3140
rect 58650 2555 58680 2570
rect 58705 3140 58735 3240
rect 58755 3190 58795 3195
rect 58755 3160 58760 3190
rect 58790 3160 58795 3190
rect 58755 3155 58795 3160
rect 58705 2570 58710 3140
rect 58730 2570 58735 3140
rect 58705 2560 58735 2570
rect 58760 3140 58790 3155
rect 58760 2570 58765 3140
rect 58785 2570 58790 3140
rect 58760 2555 58790 2570
rect 58815 3140 58845 3240
rect 58865 3190 58905 3195
rect 58865 3160 58870 3190
rect 58900 3160 58905 3190
rect 58865 3155 58905 3160
rect 58815 2570 58820 3140
rect 58840 2570 58845 3140
rect 58815 2560 58845 2570
rect 58870 3140 58900 3155
rect 58870 2570 58875 3140
rect 58895 2570 58900 3140
rect 58870 2555 58900 2570
rect 58925 3140 58955 3240
rect 58975 3190 59015 3195
rect 58975 3160 58980 3190
rect 59010 3160 59015 3190
rect 58975 3155 59015 3160
rect 58925 2570 58930 3140
rect 58950 2570 58955 3140
rect 58925 2560 58955 2570
rect 58980 3140 59010 3155
rect 58980 2570 58985 3140
rect 59005 2570 59010 3140
rect 58980 2555 59010 2570
rect 59035 3140 59065 3240
rect 59145 3200 59175 3240
rect 59505 3200 59545 3345
rect 59085 3190 59125 3195
rect 59085 3160 59090 3190
rect 59120 3160 59125 3190
rect 59085 3155 59125 3160
rect 59145 3180 59150 3200
rect 59170 3180 59175 3200
rect 59035 2570 59040 3140
rect 59060 2570 59065 3140
rect 59035 2560 59065 2570
rect 59090 3140 59120 3155
rect 59090 2570 59095 3140
rect 59115 2570 59120 3140
rect 59090 2555 59120 2570
rect 59145 3140 59175 3180
rect 59455 3190 59596 3200
rect 59455 3170 59460 3190
rect 59480 3170 59515 3190
rect 59535 3170 59570 3190
rect 59590 3170 59596 3190
rect 59455 3160 59596 3170
rect 59145 2570 59150 3140
rect 59170 2570 59175 3140
rect 59145 2560 59175 2570
rect 59455 2585 59596 2595
rect 59455 2565 59460 2585
rect 59480 2565 59515 2585
rect 59535 2565 59570 2585
rect 59590 2565 59596 2585
rect 59455 2555 59596 2565
rect 58280 2440 58285 2470
rect 58315 2440 58325 2470
rect 58355 2440 58365 2470
rect 58395 2440 58400 2470
rect 58280 2430 58400 2440
rect 58280 2400 58285 2430
rect 58315 2400 58325 2430
rect 58355 2400 58365 2430
rect 58395 2400 58400 2430
rect 58280 2390 58400 2400
rect 58280 2360 58285 2390
rect 58315 2360 58325 2390
rect 58355 2360 58365 2390
rect 58395 2360 58400 2390
rect 58280 1595 58400 2360
rect 58535 2550 58575 2555
rect 58535 2520 58540 2550
rect 58570 2520 58575 2550
rect 58535 2325 58575 2520
rect 58645 2550 58685 2555
rect 58645 2520 58650 2550
rect 58680 2520 58685 2550
rect 58645 2325 58685 2520
rect 58755 2550 58795 2555
rect 58755 2520 58760 2550
rect 58790 2520 58795 2550
rect 58755 2325 58795 2520
rect 58865 2550 58905 2555
rect 58865 2520 58870 2550
rect 58900 2520 58905 2550
rect 58810 2470 58850 2475
rect 58810 2440 58815 2470
rect 58845 2440 58850 2470
rect 58810 2430 58850 2440
rect 58810 2400 58815 2430
rect 58845 2400 58850 2430
rect 58810 2390 58850 2400
rect 58810 2360 58815 2390
rect 58845 2360 58850 2390
rect 58810 2355 58850 2360
rect 58865 2325 58905 2520
rect 58975 2550 59015 2555
rect 58975 2520 58980 2550
rect 59010 2520 59015 2550
rect 58975 2325 59015 2520
rect 59085 2550 59125 2555
rect 59085 2520 59090 2550
rect 59120 2520 59125 2550
rect 59085 2325 59125 2520
rect 59465 2470 59585 2555
rect 59465 2440 59470 2470
rect 59500 2440 59510 2470
rect 59540 2440 59550 2470
rect 59580 2440 59585 2470
rect 59465 2430 59585 2440
rect 59465 2400 59470 2430
rect 59500 2400 59510 2430
rect 59540 2400 59550 2430
rect 59580 2400 59585 2430
rect 59465 2390 59585 2400
rect 59465 2360 59470 2390
rect 59500 2360 59510 2390
rect 59540 2360 59550 2390
rect 59580 2360 59585 2390
rect 59465 2355 59585 2360
rect 58535 2320 59125 2325
rect 58535 2290 58540 2320
rect 58570 2290 58595 2320
rect 58625 2290 58650 2320
rect 58680 2290 58705 2320
rect 58735 2290 58760 2320
rect 58790 2290 58815 2320
rect 58845 2290 58870 2320
rect 58900 2290 58925 2320
rect 58955 2290 58980 2320
rect 59010 2290 59035 2320
rect 59065 2290 59090 2320
rect 59120 2290 59125 2320
rect 58535 2280 59125 2290
rect 58535 2250 58540 2280
rect 58570 2250 58595 2280
rect 58625 2250 58650 2280
rect 58680 2250 58705 2280
rect 58735 2250 58760 2280
rect 58790 2250 58815 2280
rect 58845 2250 58870 2280
rect 58900 2250 58925 2280
rect 58955 2250 58980 2280
rect 59010 2250 59035 2280
rect 59065 2250 59090 2280
rect 59120 2250 59125 2280
rect 58535 2240 59125 2250
rect 58535 2210 58540 2240
rect 58570 2210 58595 2240
rect 58625 2210 58650 2240
rect 58680 2210 58705 2240
rect 58735 2210 58760 2240
rect 58790 2210 58815 2240
rect 58845 2210 58870 2240
rect 58900 2210 58925 2240
rect 58955 2210 58980 2240
rect 59010 2210 59035 2240
rect 59065 2210 59090 2240
rect 59120 2210 59125 2240
rect 58535 2205 59125 2210
rect 59560 2320 59810 2325
rect 59560 2290 59565 2320
rect 59595 2290 59605 2320
rect 59635 2290 59650 2320
rect 59680 2290 59690 2320
rect 59720 2290 59735 2320
rect 59765 2290 59775 2320
rect 59805 2290 59810 2320
rect 59560 2280 59810 2290
rect 59560 2250 59565 2280
rect 59595 2250 59605 2280
rect 59635 2250 59650 2280
rect 59680 2250 59690 2280
rect 59720 2250 59735 2280
rect 59765 2250 59775 2280
rect 59805 2250 59810 2280
rect 59560 2240 59810 2250
rect 59560 2210 59565 2240
rect 59595 2210 59605 2240
rect 59635 2210 59650 2240
rect 59680 2210 59690 2240
rect 59720 2210 59735 2240
rect 59765 2210 59775 2240
rect 59805 2210 59810 2240
rect 58480 2185 58520 2190
rect 58480 2155 58485 2185
rect 58515 2155 58520 2185
rect 58480 2145 58520 2155
rect 58480 2115 58485 2145
rect 58515 2115 58520 2145
rect 58480 2105 58520 2115
rect 58480 2075 58485 2105
rect 58515 2075 58520 2105
rect 58480 2070 58520 2075
rect 59140 2185 59180 2190
rect 59140 2155 59145 2185
rect 59175 2155 59180 2185
rect 59140 2145 59180 2155
rect 59140 2115 59145 2145
rect 59175 2115 59180 2145
rect 59140 2105 59180 2115
rect 59140 2075 59145 2105
rect 59175 2075 59180 2105
rect 59140 2070 59180 2075
rect 58485 1925 58515 2070
rect 58535 2050 58575 2055
rect 58535 2020 58540 2050
rect 58570 2020 58575 2050
rect 58535 2010 58575 2020
rect 58535 1980 58540 2010
rect 58570 1980 58575 2010
rect 58535 1970 58575 1980
rect 58535 1940 58540 1970
rect 58570 1940 58575 1970
rect 58535 1935 58575 1940
rect 58645 2050 58685 2055
rect 58645 2020 58650 2050
rect 58680 2020 58685 2050
rect 58645 2010 58685 2020
rect 58645 1980 58650 2010
rect 58680 1980 58685 2010
rect 58645 1970 58685 1980
rect 58645 1940 58650 1970
rect 58680 1940 58685 1970
rect 58645 1935 58685 1940
rect 58755 2050 58795 2055
rect 58755 2020 58760 2050
rect 58790 2020 58795 2050
rect 58755 2010 58795 2020
rect 58755 1980 58760 2010
rect 58790 1980 58795 2010
rect 58755 1970 58795 1980
rect 58755 1940 58760 1970
rect 58790 1940 58795 1970
rect 58755 1935 58795 1940
rect 58865 2050 58905 2055
rect 58865 2020 58870 2050
rect 58900 2020 58905 2050
rect 58865 2010 58905 2020
rect 58865 1980 58870 2010
rect 58900 1980 58905 2010
rect 58865 1970 58905 1980
rect 58865 1940 58870 1970
rect 58900 1940 58905 1970
rect 58865 1935 58905 1940
rect 58975 2050 59015 2055
rect 58975 2020 58980 2050
rect 59010 2020 59015 2050
rect 58975 2010 59015 2020
rect 58975 1980 58980 2010
rect 59010 1980 59015 2010
rect 58975 1970 59015 1980
rect 58975 1940 58980 1970
rect 59010 1940 59015 1970
rect 58975 1935 59015 1940
rect 59085 2050 59125 2055
rect 59085 2020 59090 2050
rect 59120 2020 59125 2050
rect 59085 2010 59125 2020
rect 59085 1980 59090 2010
rect 59120 1980 59125 2010
rect 59085 1970 59125 1980
rect 59085 1940 59090 1970
rect 59120 1940 59125 1970
rect 59085 1935 59125 1940
rect 58485 1905 58490 1925
rect 58510 1905 58515 1925
rect 58485 1865 58515 1905
rect 58485 1695 58490 1865
rect 58510 1695 58515 1865
rect 58485 1685 58515 1695
rect 58540 1865 58570 1935
rect 58590 1915 58630 1920
rect 58590 1885 58595 1915
rect 58625 1885 58630 1915
rect 58590 1880 58630 1885
rect 58540 1695 58545 1865
rect 58565 1695 58570 1865
rect 58540 1685 58570 1695
rect 58595 1865 58625 1880
rect 58595 1695 58600 1865
rect 58620 1695 58625 1865
rect 58595 1665 58625 1695
rect 58650 1865 58680 1935
rect 58700 1915 58740 1920
rect 58700 1885 58705 1915
rect 58735 1885 58740 1915
rect 58700 1880 58740 1885
rect 58650 1695 58655 1865
rect 58675 1695 58680 1865
rect 58650 1685 58680 1695
rect 58705 1865 58735 1880
rect 58705 1695 58710 1865
rect 58730 1695 58735 1865
rect 58705 1665 58735 1695
rect 58760 1865 58790 1935
rect 58810 1915 58850 1920
rect 58810 1885 58815 1915
rect 58845 1885 58850 1915
rect 58810 1880 58850 1885
rect 58760 1695 58765 1865
rect 58785 1695 58790 1865
rect 58760 1685 58790 1695
rect 58815 1865 58845 1880
rect 58815 1695 58820 1865
rect 58840 1695 58845 1865
rect 58815 1665 58845 1695
rect 58870 1865 58900 1935
rect 58920 1915 58960 1920
rect 58920 1885 58925 1915
rect 58955 1885 58960 1915
rect 58920 1880 58960 1885
rect 58870 1695 58875 1865
rect 58895 1695 58900 1865
rect 58870 1685 58900 1695
rect 58925 1865 58955 1880
rect 58925 1695 58930 1865
rect 58950 1695 58955 1865
rect 58925 1665 58955 1695
rect 58980 1865 59010 1935
rect 59030 1915 59070 1920
rect 59030 1885 59035 1915
rect 59065 1885 59070 1915
rect 59030 1880 59070 1885
rect 58980 1695 58985 1865
rect 59005 1695 59010 1865
rect 58980 1685 59010 1695
rect 59035 1865 59065 1880
rect 59035 1695 59040 1865
rect 59060 1695 59065 1865
rect 59035 1665 59065 1695
rect 59090 1865 59120 1935
rect 59090 1695 59095 1865
rect 59115 1695 59120 1865
rect 59090 1685 59120 1695
rect 59145 1925 59175 2070
rect 59145 1905 59150 1925
rect 59170 1905 59175 1925
rect 59145 1865 59175 1905
rect 59145 1695 59150 1865
rect 59170 1695 59175 1865
rect 59145 1685 59175 1695
rect 59560 1710 59810 2210
rect 59560 1680 59570 1710
rect 59600 1680 59620 1710
rect 59650 1680 59670 1710
rect 59700 1680 59720 1710
rect 59750 1680 59770 1710
rect 59800 1680 59810 1710
rect 58590 1660 58630 1665
rect 58590 1630 58595 1660
rect 58625 1630 58630 1660
rect 58590 1625 58630 1630
rect 58700 1660 58740 1665
rect 58700 1630 58705 1660
rect 58735 1630 58740 1660
rect 58700 1625 58740 1630
rect 58810 1660 58850 1665
rect 58810 1630 58815 1660
rect 58845 1630 58850 1660
rect 58810 1625 58850 1630
rect 58920 1660 58960 1665
rect 58920 1630 58925 1660
rect 58955 1630 58960 1660
rect 58920 1625 58960 1630
rect 59030 1660 59070 1665
rect 59030 1630 59035 1660
rect 59065 1630 59070 1660
rect 59030 1625 59070 1630
rect 59275 1660 59315 1665
rect 59275 1630 59280 1660
rect 59310 1630 59315 1660
rect 59275 1625 59315 1630
rect 59560 1660 59810 1680
rect 59560 1630 59570 1660
rect 59600 1630 59620 1660
rect 59650 1630 59670 1660
rect 59700 1630 59720 1660
rect 59750 1630 59770 1660
rect 59800 1630 59810 1660
rect 58280 1565 58285 1595
rect 58315 1565 58325 1595
rect 58355 1565 58365 1595
rect 58395 1565 58400 1595
rect 58280 1555 58400 1565
rect 58280 1525 58285 1555
rect 58315 1525 58325 1555
rect 58355 1525 58365 1555
rect 58395 1525 58400 1555
rect 58280 1520 58400 1525
rect 58645 1595 58685 1600
rect 58645 1565 58650 1595
rect 58680 1565 58685 1595
rect 58645 1555 58685 1565
rect 58645 1525 58650 1555
rect 58680 1525 58685 1555
rect 58645 1520 58685 1525
rect 58590 1475 58630 1480
rect 58590 1445 58595 1475
rect 58625 1445 58630 1475
rect 58590 1440 58630 1445
rect 58700 1475 58740 1480
rect 58700 1445 58705 1475
rect 58735 1445 58740 1475
rect 58700 1440 58740 1445
rect 58810 1475 58850 1480
rect 58810 1445 58815 1475
rect 58845 1445 58850 1475
rect 58810 1440 58850 1445
rect 58920 1475 58960 1480
rect 58920 1445 58925 1475
rect 58955 1445 58960 1475
rect 58920 1440 58960 1445
rect 59030 1475 59070 1480
rect 59030 1445 59035 1475
rect 59065 1445 59070 1475
rect 59030 1440 59070 1445
rect 59230 1475 59270 1480
rect 59230 1445 59235 1475
rect 59265 1445 59270 1475
rect 59230 1440 59270 1445
rect 58145 1050 58150 1080
rect 58180 1050 58190 1080
rect 58220 1050 58230 1080
rect 58260 1050 58265 1080
rect 58145 1040 58265 1050
rect 58145 1010 58150 1040
rect 58180 1010 58190 1040
rect 58220 1010 58230 1040
rect 58260 1010 58265 1040
rect 58145 1000 58265 1010
rect 58145 970 58150 1000
rect 58180 970 58190 1000
rect 58220 970 58230 1000
rect 58260 970 58265 1000
rect 58145 965 58265 970
rect 58485 1425 58515 1435
rect 58485 1155 58490 1425
rect 58510 1155 58515 1425
rect 58485 1115 58515 1155
rect 58485 1095 58490 1115
rect 58510 1095 58515 1115
rect 58485 945 58515 1095
rect 58540 1425 58570 1435
rect 58540 1155 58545 1425
rect 58565 1155 58570 1425
rect 58540 1085 58570 1155
rect 58595 1425 58625 1440
rect 58595 1155 58600 1425
rect 58620 1155 58625 1425
rect 58595 1140 58625 1155
rect 58650 1425 58680 1435
rect 58650 1155 58655 1425
rect 58675 1155 58680 1425
rect 58590 1135 58630 1140
rect 58590 1105 58595 1135
rect 58625 1105 58630 1135
rect 58590 1100 58630 1105
rect 58650 1085 58680 1155
rect 58705 1425 58735 1440
rect 58705 1155 58710 1425
rect 58730 1155 58735 1425
rect 58705 1140 58735 1155
rect 58760 1425 58790 1435
rect 58760 1155 58765 1425
rect 58785 1155 58790 1425
rect 58700 1135 58740 1140
rect 58700 1105 58705 1135
rect 58735 1105 58740 1135
rect 58700 1100 58740 1105
rect 58760 1085 58790 1155
rect 58815 1425 58845 1440
rect 58815 1155 58820 1425
rect 58840 1155 58845 1425
rect 58815 1140 58845 1155
rect 58870 1425 58900 1435
rect 58870 1155 58875 1425
rect 58895 1155 58900 1425
rect 58810 1135 58850 1140
rect 58810 1105 58815 1135
rect 58845 1105 58850 1135
rect 58810 1100 58850 1105
rect 58870 1085 58900 1155
rect 58925 1425 58955 1440
rect 58925 1155 58930 1425
rect 58950 1155 58955 1425
rect 58925 1140 58955 1155
rect 58980 1425 59010 1435
rect 58980 1155 58985 1425
rect 59005 1155 59010 1425
rect 58920 1135 58960 1140
rect 58920 1105 58925 1135
rect 58955 1105 58960 1135
rect 58920 1100 58960 1105
rect 58980 1085 59010 1155
rect 59035 1425 59065 1440
rect 59035 1155 59040 1425
rect 59060 1155 59065 1425
rect 59035 1140 59065 1155
rect 59090 1425 59120 1435
rect 59090 1155 59095 1425
rect 59115 1155 59120 1425
rect 59030 1135 59070 1140
rect 59030 1105 59035 1135
rect 59065 1105 59070 1135
rect 59030 1100 59070 1105
rect 59090 1085 59120 1155
rect 59145 1425 59175 1435
rect 59145 1155 59150 1425
rect 59170 1155 59175 1425
rect 59240 1160 59260 1440
rect 59145 1115 59175 1155
rect 59230 1155 59270 1160
rect 59230 1125 59235 1155
rect 59265 1125 59270 1155
rect 59230 1120 59270 1125
rect 59145 1095 59150 1115
rect 59170 1095 59175 1115
rect 58535 1080 58575 1085
rect 58535 1050 58540 1080
rect 58570 1050 58575 1080
rect 58535 1040 58575 1050
rect 58535 1010 58540 1040
rect 58570 1010 58575 1040
rect 58535 1000 58575 1010
rect 58535 970 58540 1000
rect 58570 970 58575 1000
rect 58535 965 58575 970
rect 58645 1080 58685 1085
rect 58645 1050 58650 1080
rect 58680 1050 58685 1080
rect 58645 1040 58685 1050
rect 58645 1010 58650 1040
rect 58680 1010 58685 1040
rect 58645 1000 58685 1010
rect 58645 970 58650 1000
rect 58680 970 58685 1000
rect 58645 965 58685 970
rect 58755 1080 58795 1085
rect 58755 1050 58760 1080
rect 58790 1050 58795 1080
rect 58755 1040 58795 1050
rect 58755 1010 58760 1040
rect 58790 1010 58795 1040
rect 58755 1000 58795 1010
rect 58755 970 58760 1000
rect 58790 970 58795 1000
rect 58755 965 58795 970
rect 58865 1080 58905 1085
rect 58865 1050 58870 1080
rect 58900 1050 58905 1080
rect 58865 1040 58905 1050
rect 58865 1010 58870 1040
rect 58900 1010 58905 1040
rect 58865 1000 58905 1010
rect 58865 970 58870 1000
rect 58900 970 58905 1000
rect 58865 965 58905 970
rect 58975 1080 59015 1085
rect 58975 1050 58980 1080
rect 59010 1050 59015 1080
rect 58975 1040 59015 1050
rect 58975 1010 58980 1040
rect 59010 1010 59015 1040
rect 58975 1000 59015 1010
rect 58975 970 58980 1000
rect 59010 970 59015 1000
rect 58975 965 59015 970
rect 59085 1080 59125 1085
rect 59085 1050 59090 1080
rect 59120 1050 59125 1080
rect 59085 1040 59125 1050
rect 59085 1010 59090 1040
rect 59120 1010 59125 1040
rect 59085 1000 59125 1010
rect 59085 970 59090 1000
rect 59120 970 59125 1000
rect 59085 965 59125 970
rect 59145 945 59175 1095
rect 59285 1090 59305 1625
rect 59560 1610 59810 1630
rect 59560 1580 59570 1610
rect 59600 1580 59620 1610
rect 59650 1580 59670 1610
rect 59700 1580 59720 1610
rect 59750 1580 59770 1610
rect 59800 1580 59810 1610
rect 59330 1160 59365 1165
rect 59330 1120 59365 1125
rect 59390 1160 59425 1165
rect 59390 1120 59425 1125
rect 59450 1160 59485 1165
rect 59450 1120 59485 1125
rect 59510 1160 59545 1166
rect 59510 1120 59545 1125
rect 59395 1090 59415 1120
rect 59275 1085 59315 1090
rect 59275 1055 59280 1085
rect 59310 1055 59315 1085
rect 59275 1050 59315 1055
rect 59385 1085 59425 1090
rect 59385 1055 59390 1085
rect 59420 1055 59425 1085
rect 59385 1050 59425 1055
rect 58480 940 58520 945
rect 58480 910 58485 940
rect 58515 910 58520 940
rect 58480 900 58520 910
rect 58480 870 58485 900
rect 58515 870 58520 900
rect 58480 860 58520 870
rect 58480 830 58485 860
rect 58515 830 58520 860
rect 58480 825 58520 830
rect 59140 940 59180 945
rect 59140 910 59145 940
rect 59175 910 59180 940
rect 59140 900 59180 910
rect 59140 870 59145 900
rect 59175 870 59180 900
rect 59140 860 59180 870
rect 59140 830 59145 860
rect 59175 830 59180 860
rect 59140 825 59180 830
rect 59515 810 59535 1120
rect 59505 805 59545 810
rect 59505 775 59510 805
rect 59540 775 59545 805
rect 59505 770 59545 775
rect 58760 525 58800 530
rect 58760 495 58765 525
rect 58795 495 58800 525
rect 58760 490 58800 495
rect 59440 525 59480 530
rect 59440 495 59445 525
rect 59475 495 59480 525
rect 59440 490 59480 495
rect 58610 470 59050 475
rect 58610 440 58615 470
rect 58645 440 58655 470
rect 58685 440 58695 470
rect 58725 440 58735 470
rect 58765 440 58775 470
rect 58805 440 58815 470
rect 58845 440 58855 470
rect 58885 440 58895 470
rect 58925 440 58935 470
rect 58965 440 58975 470
rect 59005 440 59015 470
rect 59045 440 59050 470
rect 58610 430 59050 440
rect 58610 400 58615 430
rect 58645 400 58655 430
rect 58685 400 58695 430
rect 58725 400 58735 430
rect 58765 400 58775 430
rect 58805 400 58815 430
rect 58845 400 58855 430
rect 58885 400 58895 430
rect 58925 400 58935 430
rect 58965 400 58975 430
rect 59005 400 59015 430
rect 59045 400 59050 430
rect 58610 390 59050 400
rect 58610 360 58615 390
rect 58645 360 58655 390
rect 58685 360 58695 390
rect 58725 360 58735 390
rect 58765 360 58775 390
rect 58805 360 58815 390
rect 58845 360 58855 390
rect 58885 360 58895 390
rect 58925 360 58935 390
rect 58965 360 58975 390
rect 59005 360 59015 390
rect 59045 360 59050 390
rect 58610 355 59050 360
rect 59375 470 59415 475
rect 59375 440 59380 470
rect 59410 440 59415 470
rect 59375 430 59415 440
rect 59375 400 59380 430
rect 59410 400 59415 430
rect 59375 390 59415 400
rect 59375 360 59380 390
rect 59410 360 59415 390
rect 59375 355 59415 360
rect 58010 -90 58015 -60
rect 58045 -90 58055 -60
rect 58085 -90 58095 -60
rect 58125 -90 58130 -60
rect 58010 -100 58130 -90
rect 58010 -130 58015 -100
rect 58045 -130 58055 -100
rect 58085 -130 58095 -100
rect 58125 -130 58130 -100
rect 58010 -140 58130 -130
rect 58010 -170 58015 -140
rect 58045 -170 58055 -140
rect 58085 -170 58095 -140
rect 58125 -170 58130 -140
rect 58010 -175 58130 -170
rect 58515 325 58545 335
rect 58515 -345 58520 325
rect 58540 -345 58545 325
rect 58515 -385 58545 -345
rect 58615 325 58645 355
rect 58615 -345 58620 325
rect 58640 -345 58645 325
rect 58615 -360 58645 -345
rect 58715 325 58745 335
rect 58715 -345 58720 325
rect 58740 -345 58745 325
rect 58515 -405 58520 -385
rect 58540 -405 58545 -385
rect 58610 -365 58650 -360
rect 58610 -395 58615 -365
rect 58645 -395 58650 -365
rect 58610 -400 58650 -395
rect 58515 -575 58545 -405
rect 58715 -575 58745 -345
rect 58815 325 58845 355
rect 58815 -345 58820 325
rect 58840 -345 58845 325
rect 58815 -360 58845 -345
rect 58915 325 58945 335
rect 58915 -345 58920 325
rect 58940 -345 58945 325
rect 58810 -365 58850 -360
rect 58810 -395 58815 -365
rect 58845 -395 58850 -365
rect 58810 -400 58850 -395
rect 57485 -610 57490 -580
rect 57520 -610 57525 -580
rect 57485 -620 57525 -610
rect 57485 -650 57490 -620
rect 57520 -650 57525 -620
rect 57485 -660 57525 -650
rect 57485 -690 57490 -660
rect 57520 -690 57525 -660
rect 57485 -695 57525 -690
rect 57540 -580 57660 -575
rect 57540 -610 57545 -580
rect 57575 -610 57585 -580
rect 57615 -610 57625 -580
rect 57655 -610 57660 -580
rect 57540 -620 57660 -610
rect 57540 -650 57545 -620
rect 57575 -650 57585 -620
rect 57615 -650 57625 -620
rect 57655 -650 57660 -620
rect 57540 -660 57660 -650
rect 57540 -690 57545 -660
rect 57575 -690 57585 -660
rect 57615 -690 57625 -660
rect 57655 -690 57660 -660
rect 57540 -1500 57660 -690
rect 57890 -580 58010 -575
rect 57890 -610 57895 -580
rect 57925 -610 57935 -580
rect 57965 -610 57975 -580
rect 58005 -610 58010 -580
rect 57890 -620 58010 -610
rect 57890 -650 57895 -620
rect 57925 -650 57935 -620
rect 57965 -650 57975 -620
rect 58005 -650 58010 -620
rect 57890 -660 58010 -650
rect 57890 -690 57895 -660
rect 57925 -690 57935 -660
rect 57965 -690 57975 -660
rect 58005 -690 58010 -660
rect 57890 -1500 58010 -690
rect 58240 -580 58360 -575
rect 58240 -610 58245 -580
rect 58275 -610 58285 -580
rect 58315 -610 58325 -580
rect 58355 -610 58360 -580
rect 58240 -620 58360 -610
rect 58240 -650 58245 -620
rect 58275 -650 58285 -620
rect 58315 -650 58325 -620
rect 58355 -650 58360 -620
rect 58240 -660 58360 -650
rect 58240 -690 58245 -660
rect 58275 -690 58285 -660
rect 58315 -690 58325 -660
rect 58355 -690 58360 -660
rect 58240 -1500 58360 -690
rect 58510 -580 58550 -575
rect 58510 -610 58515 -580
rect 58545 -610 58550 -580
rect 58510 -620 58550 -610
rect 58510 -650 58515 -620
rect 58545 -650 58550 -620
rect 58510 -660 58550 -650
rect 58510 -690 58515 -660
rect 58545 -690 58550 -660
rect 58510 -695 58550 -690
rect 58590 -580 58745 -575
rect 58590 -610 58595 -580
rect 58625 -610 58635 -580
rect 58665 -610 58675 -580
rect 58705 -610 58745 -580
rect 58590 -620 58745 -610
rect 58590 -650 58595 -620
rect 58625 -650 58635 -620
rect 58665 -650 58675 -620
rect 58705 -650 58745 -620
rect 58590 -660 58745 -650
rect 58590 -690 58595 -660
rect 58625 -690 58635 -660
rect 58665 -690 58675 -660
rect 58705 -690 58745 -660
rect 58590 -695 58745 -690
rect 58915 -575 58945 -345
rect 59015 325 59045 355
rect 59380 335 59415 355
rect 59450 340 59470 490
rect 59560 470 59810 1580
rect 59560 440 59565 470
rect 59595 440 59605 470
rect 59635 440 59650 470
rect 59680 440 59690 470
rect 59720 440 59735 470
rect 59765 440 59775 470
rect 59805 440 59810 470
rect 59560 430 59810 440
rect 59560 400 59565 430
rect 59595 400 59605 430
rect 59635 400 59650 430
rect 59680 400 59690 430
rect 59720 400 59735 430
rect 59765 400 59775 430
rect 59805 400 59810 430
rect 59560 390 59810 400
rect 59560 360 59565 390
rect 59595 360 59605 390
rect 59635 360 59650 390
rect 59680 360 59690 390
rect 59720 360 59735 390
rect 59765 360 59775 390
rect 59805 360 59810 390
rect 59560 355 59810 360
rect 59840 2050 59960 2055
rect 59840 2020 59845 2050
rect 59875 2020 59885 2050
rect 59915 2020 59925 2050
rect 59955 2020 59960 2050
rect 59840 2010 59960 2020
rect 59840 1980 59845 2010
rect 59875 1980 59885 2010
rect 59915 1980 59925 2010
rect 59955 1980 59960 2010
rect 59840 1970 59960 1980
rect 59840 1940 59845 1970
rect 59875 1940 59885 1970
rect 59915 1940 59925 1970
rect 59955 1940 59960 1970
rect 59840 940 59960 1940
rect 59840 910 59845 940
rect 59875 910 59885 940
rect 59915 910 59925 940
rect 59955 910 59960 940
rect 59840 900 59960 910
rect 59840 870 59845 900
rect 59875 870 59885 900
rect 59915 870 59925 900
rect 59955 870 59960 900
rect 59840 860 59960 870
rect 59840 830 59845 860
rect 59875 830 59885 860
rect 59915 830 59925 860
rect 59955 830 59960 860
rect 59015 -345 59020 325
rect 59040 -345 59045 325
rect 59015 -360 59045 -345
rect 59115 325 59145 335
rect 59115 -345 59120 325
rect 59140 -345 59145 325
rect 59380 295 59415 300
rect 59440 335 59475 340
rect 59440 295 59475 300
rect 59010 -365 59050 -360
rect 59010 -395 59015 -365
rect 59045 -395 59050 -365
rect 59010 -400 59050 -395
rect 59115 -385 59145 -345
rect 59115 -405 59120 -385
rect 59140 -405 59145 -385
rect 59115 -575 59145 -405
rect 58915 -580 59060 -575
rect 58915 -610 58945 -580
rect 58975 -610 58985 -580
rect 59015 -610 59025 -580
rect 59055 -610 59060 -580
rect 58915 -620 59060 -610
rect 58915 -650 58945 -620
rect 58975 -650 58985 -620
rect 59015 -650 59025 -620
rect 59055 -650 59060 -620
rect 58915 -660 59060 -650
rect 58915 -690 58945 -660
rect 58975 -690 58985 -660
rect 59015 -690 59025 -660
rect 59055 -690 59060 -660
rect 58915 -695 59060 -690
rect 59110 -580 59150 -575
rect 59110 -610 59115 -580
rect 59145 -610 59150 -580
rect 59110 -620 59150 -610
rect 59110 -650 59115 -620
rect 59145 -650 59150 -620
rect 59110 -660 59150 -650
rect 59110 -690 59115 -660
rect 59145 -690 59150 -660
rect 59110 -695 59150 -690
rect 59370 -580 59490 -575
rect 59370 -610 59375 -580
rect 59405 -610 59415 -580
rect 59445 -610 59455 -580
rect 59485 -610 59490 -580
rect 59370 -620 59490 -610
rect 59370 -650 59375 -620
rect 59405 -650 59415 -620
rect 59445 -650 59455 -620
rect 59485 -650 59490 -620
rect 59370 -660 59490 -650
rect 59370 -690 59375 -660
rect 59405 -690 59415 -660
rect 59445 -690 59455 -660
rect 59485 -690 59490 -660
rect 59370 -695 59490 -690
rect 59640 -580 59760 -575
rect 59640 -610 59645 -580
rect 59675 -610 59685 -580
rect 59715 -610 59725 -580
rect 59755 -610 59760 -580
rect 59640 -620 59760 -610
rect 59640 -650 59645 -620
rect 59675 -650 59685 -620
rect 59715 -650 59725 -620
rect 59755 -650 59760 -620
rect 59640 -660 59760 -650
rect 59640 -690 59645 -660
rect 59675 -690 59685 -660
rect 59715 -690 59725 -660
rect 59755 -690 59760 -660
rect 58590 -1500 58710 -695
rect 58940 -1500 59060 -695
rect 59290 -1500 59410 -695
rect 59640 -1500 59760 -690
rect 59840 -580 59960 830
rect 59840 -610 59845 -580
rect 59875 -610 59885 -580
rect 59915 -610 59925 -580
rect 59955 -610 59960 -580
rect 59840 -620 59960 -610
rect 59840 -650 59845 -620
rect 59875 -650 59885 -620
rect 59915 -650 59925 -620
rect 59955 -650 59960 -620
rect 59840 -660 59960 -650
rect 59840 -690 59845 -660
rect 59875 -690 59885 -660
rect 59915 -690 59925 -660
rect 59955 -690 59960 -660
rect 59840 -695 59960 -690
rect 59990 -580 60110 -575
rect 59990 -610 59995 -580
rect 60025 -610 60035 -580
rect 60065 -610 60075 -580
rect 60105 -610 60110 -580
rect 59990 -620 60110 -610
rect 59990 -650 59995 -620
rect 60025 -650 60035 -620
rect 60065 -650 60075 -620
rect 60105 -650 60110 -620
rect 59990 -660 60110 -650
rect 59990 -690 59995 -660
rect 60025 -690 60035 -660
rect 60065 -690 60075 -660
rect 60105 -690 60110 -660
rect 59990 -1500 60110 -690
rect 60340 -580 60460 -575
rect 60340 -610 60345 -580
rect 60375 -610 60385 -580
rect 60415 -610 60425 -580
rect 60455 -610 60460 -580
rect 60340 -620 60460 -610
rect 60340 -650 60345 -620
rect 60375 -650 60385 -620
rect 60415 -650 60425 -620
rect 60455 -650 60460 -620
rect 60340 -660 60460 -650
rect 60340 -690 60345 -660
rect 60375 -690 60385 -660
rect 60415 -690 60425 -660
rect 60455 -690 60460 -660
rect 60340 -1500 60460 -690
rect 60690 -580 60810 -575
rect 60690 -610 60695 -580
rect 60725 -610 60735 -580
rect 60765 -610 60775 -580
rect 60805 -610 60810 -580
rect 60690 -620 60810 -610
rect 60690 -650 60695 -620
rect 60725 -650 60735 -620
rect 60765 -650 60775 -620
rect 60805 -650 60810 -620
rect 60690 -660 60810 -650
rect 60690 -690 60695 -660
rect 60725 -690 60735 -660
rect 60765 -690 60775 -660
rect 60805 -690 60810 -660
rect 60690 -1500 60810 -690
rect 61040 -580 61160 -575
rect 61040 -610 61045 -580
rect 61075 -610 61085 -580
rect 61115 -610 61125 -580
rect 61155 -610 61160 -580
rect 61040 -620 61160 -610
rect 61040 -650 61045 -620
rect 61075 -650 61085 -620
rect 61115 -650 61125 -620
rect 61155 -650 61160 -620
rect 61040 -660 61160 -650
rect 61040 -690 61045 -660
rect 61075 -690 61085 -660
rect 61115 -690 61125 -660
rect 61155 -690 61160 -660
rect 61040 -1500 61160 -690
rect 61390 -580 61510 -575
rect 61390 -610 61395 -580
rect 61425 -610 61435 -580
rect 61465 -610 61475 -580
rect 61505 -610 61510 -580
rect 61390 -620 61510 -610
rect 61390 -650 61395 -620
rect 61425 -650 61435 -620
rect 61465 -650 61475 -620
rect 61505 -650 61510 -620
rect 61390 -660 61510 -650
rect 61390 -690 61395 -660
rect 61425 -690 61435 -660
rect 61465 -690 61475 -660
rect 61505 -690 61510 -660
rect 61390 -1500 61510 -690
<< via1 >>
rect 52295 4290 52325 4320
rect 52335 4290 52365 4320
rect 52375 4290 52405 4320
rect 52295 4250 52325 4280
rect 52335 4250 52365 4280
rect 52375 4250 52405 4280
rect 52295 4210 52325 4240
rect 52335 4210 52365 4240
rect 52375 4210 52405 4240
rect 52645 4290 52675 4320
rect 52685 4290 52715 4320
rect 52725 4290 52755 4320
rect 52645 4250 52675 4280
rect 52685 4250 52715 4280
rect 52725 4250 52755 4280
rect 52645 4210 52675 4240
rect 52685 4210 52715 4240
rect 52725 4210 52755 4240
rect 52995 4290 53025 4320
rect 53035 4290 53065 4320
rect 53075 4290 53105 4320
rect 52995 4250 53025 4280
rect 53035 4250 53065 4280
rect 53075 4250 53105 4280
rect 52995 4210 53025 4240
rect 53035 4210 53065 4240
rect 53075 4210 53105 4240
rect 53345 4290 53375 4320
rect 53385 4290 53415 4320
rect 53425 4290 53455 4320
rect 53345 4250 53375 4280
rect 53385 4250 53415 4280
rect 53425 4250 53455 4280
rect 53345 4210 53375 4240
rect 53385 4210 53415 4240
rect 53425 4210 53455 4240
rect 56210 5035 56240 5065
rect 56090 4925 56120 4930
rect 56090 4905 56095 4925
rect 56095 4905 56115 4925
rect 56115 4905 56120 4925
rect 56090 4900 56120 4905
rect 56680 5035 56710 5065
rect 57090 5035 57120 5065
rect 57560 5035 57590 5065
rect 56210 4900 56240 4930
rect 56270 4925 56300 4930
rect 56270 4905 56275 4925
rect 56275 4905 56295 4925
rect 56295 4905 56300 4925
rect 56270 4900 56300 4905
rect 56560 4810 56590 4840
rect 56560 4770 56590 4800
rect 56560 4755 56590 4760
rect 56560 4735 56565 4755
rect 56565 4735 56585 4755
rect 56585 4735 56590 4755
rect 56560 4730 56590 4735
rect 56620 4810 56650 4840
rect 56620 4770 56650 4800
rect 56620 4730 56650 4760
rect 56885 4980 56915 5010
rect 56885 4940 56915 4970
rect 56885 4900 56915 4930
rect 56740 4810 56770 4840
rect 56740 4770 56770 4800
rect 56740 4755 56770 4760
rect 56740 4735 56745 4755
rect 56745 4735 56765 4755
rect 56765 4735 56770 4755
rect 56740 4730 56770 4735
rect 57030 4980 57060 5010
rect 57030 4940 57060 4970
rect 57030 4925 57060 4930
rect 57030 4905 57035 4925
rect 57035 4905 57055 4925
rect 57055 4905 57060 4925
rect 57030 4900 57060 4905
rect 56885 4810 56915 4840
rect 56885 4770 56915 4800
rect 56885 4730 56915 4760
rect 56210 4495 56240 4525
rect 56680 4495 56710 4525
rect 56155 4475 56185 4480
rect 56155 4455 56160 4475
rect 56160 4455 56180 4475
rect 56180 4455 56185 4475
rect 56155 4450 56185 4455
rect 56630 4475 56660 4480
rect 56630 4455 56635 4475
rect 56635 4455 56655 4475
rect 56655 4455 56660 4475
rect 56630 4450 56660 4455
rect 56830 4450 56860 4480
rect 54045 4290 54075 4320
rect 54085 4290 54115 4320
rect 54125 4290 54155 4320
rect 54045 4250 54075 4280
rect 54085 4250 54115 4280
rect 54125 4250 54155 4280
rect 54045 4210 54075 4240
rect 54085 4210 54115 4240
rect 54125 4210 54155 4240
rect 54595 4290 54625 4320
rect 54595 4250 54625 4280
rect 54595 4210 54625 4240
rect 54955 4290 54985 4320
rect 54955 4250 54985 4280
rect 54955 4210 54985 4240
rect 54655 4155 54685 4185
rect 54695 4155 54725 4185
rect 54735 4155 54765 4185
rect 54775 4155 54805 4185
rect 54815 4155 54845 4185
rect 54855 4155 54885 4185
rect 54895 4155 54925 4185
rect 54655 4115 54685 4145
rect 54695 4115 54725 4145
rect 54735 4115 54765 4145
rect 54775 4115 54805 4145
rect 54815 4115 54845 4145
rect 54855 4115 54885 4145
rect 54895 4115 54925 4145
rect 54655 4075 54685 4105
rect 54695 4075 54725 4105
rect 54735 4075 54765 4105
rect 54775 4075 54805 4105
rect 54815 4075 54845 4105
rect 54855 4075 54885 4105
rect 54895 4075 54925 4105
rect 54595 4020 54625 4050
rect 54715 4020 54745 4050
rect 54835 4020 54865 4050
rect 55315 4290 55345 4320
rect 55315 4250 55345 4280
rect 55315 4210 55345 4240
rect 55015 4155 55045 4185
rect 55055 4155 55085 4185
rect 55095 4155 55125 4185
rect 55135 4155 55165 4185
rect 55175 4155 55205 4185
rect 55215 4155 55245 4185
rect 55255 4155 55285 4185
rect 55015 4115 55045 4145
rect 55055 4115 55085 4145
rect 55095 4115 55125 4145
rect 55135 4115 55165 4145
rect 55175 4115 55205 4145
rect 55215 4115 55245 4145
rect 55255 4115 55285 4145
rect 55015 4075 55045 4105
rect 55055 4075 55085 4105
rect 55095 4075 55125 4105
rect 55135 4075 55165 4105
rect 55175 4075 55205 4105
rect 55215 4075 55245 4105
rect 55255 4075 55285 4105
rect 54955 4020 54985 4050
rect 55075 4020 55105 4050
rect 55195 4020 55225 4050
rect 55315 4020 55345 4050
rect 55540 4290 55570 4320
rect 55580 4290 55610 4320
rect 55620 4290 55650 4320
rect 55540 4250 55570 4280
rect 55580 4250 55610 4280
rect 55620 4250 55650 4280
rect 55540 4210 55570 4240
rect 55580 4210 55610 4240
rect 55620 4210 55650 4240
rect 54655 3630 54685 3660
rect 54775 3630 54805 3660
rect 54895 3630 54925 3660
rect 55015 3630 55045 3660
rect 55135 3630 55165 3660
rect 55255 3630 55285 3660
rect 54955 3530 54985 3535
rect 54955 3510 54960 3530
rect 54960 3510 54980 3530
rect 54980 3510 54985 3530
rect 54955 3505 54985 3510
rect 55405 3460 55435 3490
rect 55445 3460 55475 3490
rect 55485 3460 55515 3490
rect 55405 3420 55435 3450
rect 55445 3420 55475 3450
rect 55485 3420 55515 3450
rect 55405 3380 55435 3410
rect 55445 3380 55475 3410
rect 55485 3380 55515 3410
rect 54260 3345 54290 3375
rect 54625 3325 54655 3355
rect 54625 3285 54655 3315
rect 54625 3245 54655 3275
rect 54735 3325 54765 3355
rect 54735 3285 54765 3315
rect 54735 3245 54765 3275
rect 54845 3325 54875 3355
rect 54845 3285 54875 3315
rect 54845 3245 54875 3275
rect 54955 3325 54985 3355
rect 54955 3285 54985 3315
rect 54955 3245 54985 3275
rect 55065 3325 55095 3355
rect 55065 3285 55095 3315
rect 55065 3245 55095 3275
rect 55175 3325 55205 3355
rect 55175 3285 55205 3315
rect 55175 3245 55205 3275
rect 55285 3325 55315 3355
rect 55285 3285 55315 3315
rect 55285 3245 55315 3275
rect 54680 3160 54710 3190
rect 54790 3160 54820 3190
rect 54900 3160 54930 3190
rect 55010 3160 55040 3190
rect 55120 3160 55150 3190
rect 55230 3160 55260 3190
rect 54220 2440 54250 2470
rect 54260 2440 54290 2470
rect 54300 2440 54330 2470
rect 54220 2400 54250 2430
rect 54260 2400 54290 2430
rect 54300 2400 54330 2430
rect 54220 2360 54250 2390
rect 54260 2360 54290 2390
rect 54300 2360 54330 2390
rect 54680 2520 54710 2550
rect 54790 2520 54820 2550
rect 54900 2520 54930 2550
rect 55010 2520 55040 2550
rect 54955 2465 54985 2470
rect 54955 2445 54960 2465
rect 54960 2445 54980 2465
rect 54980 2445 54985 2465
rect 54955 2440 54985 2445
rect 54955 2425 54985 2430
rect 54955 2405 54960 2425
rect 54960 2405 54980 2425
rect 54980 2405 54985 2425
rect 54955 2400 54985 2405
rect 54955 2385 54985 2390
rect 54955 2365 54960 2385
rect 54960 2365 54980 2385
rect 54980 2365 54985 2385
rect 54955 2360 54985 2365
rect 55120 2520 55150 2550
rect 55230 2520 55260 2550
rect 53995 2290 54025 2320
rect 54035 2290 54065 2320
rect 54080 2290 54110 2320
rect 54120 2290 54150 2320
rect 54165 2290 54195 2320
rect 54205 2290 54235 2320
rect 53995 2250 54025 2280
rect 54035 2250 54065 2280
rect 54080 2250 54110 2280
rect 54120 2250 54150 2280
rect 54165 2250 54195 2280
rect 54205 2250 54235 2280
rect 53995 2210 54025 2240
rect 54035 2210 54065 2240
rect 54080 2210 54110 2240
rect 54120 2210 54150 2240
rect 54165 2210 54195 2240
rect 54205 2210 54235 2240
rect 53845 2020 53875 2050
rect 53885 2020 53915 2050
rect 53925 2020 53955 2050
rect 53845 1980 53875 2010
rect 53885 1980 53915 2010
rect 53925 1980 53955 2010
rect 53845 1940 53875 1970
rect 53885 1940 53915 1970
rect 53925 1940 53955 1970
rect 53845 910 53875 940
rect 53885 910 53915 940
rect 53925 910 53955 940
rect 53845 870 53875 900
rect 53885 870 53915 900
rect 53925 870 53955 900
rect 53845 830 53875 860
rect 53885 830 53915 860
rect 53925 830 53955 860
rect 52295 -610 52325 -580
rect 52335 -610 52365 -580
rect 52375 -610 52405 -580
rect 52295 -650 52325 -620
rect 52335 -650 52365 -620
rect 52375 -650 52405 -620
rect 52295 -690 52325 -660
rect 52335 -690 52365 -660
rect 52375 -690 52405 -660
rect 52645 -610 52675 -580
rect 52685 -610 52715 -580
rect 52725 -610 52755 -580
rect 52645 -650 52675 -620
rect 52685 -650 52715 -620
rect 52725 -650 52755 -620
rect 52645 -690 52675 -660
rect 52685 -690 52715 -660
rect 52725 -690 52755 -660
rect 52995 -610 53025 -580
rect 53035 -610 53065 -580
rect 53075 -610 53105 -580
rect 52995 -650 53025 -620
rect 53035 -650 53065 -620
rect 53075 -650 53105 -620
rect 52995 -690 53025 -660
rect 53035 -690 53065 -660
rect 53075 -690 53105 -660
rect 53345 -610 53375 -580
rect 53385 -610 53415 -580
rect 53425 -610 53455 -580
rect 53345 -650 53375 -620
rect 53385 -650 53415 -620
rect 53425 -650 53455 -620
rect 53345 -690 53375 -660
rect 53385 -690 53415 -660
rect 53425 -690 53455 -660
rect 53695 -610 53725 -580
rect 53735 -610 53765 -580
rect 53775 -610 53805 -580
rect 53695 -650 53725 -620
rect 53735 -650 53765 -620
rect 53775 -650 53805 -620
rect 53695 -690 53725 -660
rect 53735 -690 53765 -660
rect 53775 -690 53805 -660
rect 54680 2290 54710 2320
rect 54735 2290 54765 2320
rect 54790 2290 54820 2320
rect 54845 2290 54875 2320
rect 54900 2290 54930 2320
rect 54955 2290 54985 2320
rect 55010 2290 55040 2320
rect 55065 2290 55095 2320
rect 55120 2290 55150 2320
rect 55175 2290 55205 2320
rect 55230 2290 55260 2320
rect 54680 2250 54710 2280
rect 54735 2250 54765 2280
rect 54790 2250 54820 2280
rect 54845 2250 54875 2280
rect 54900 2250 54930 2280
rect 54955 2250 54985 2280
rect 55010 2250 55040 2280
rect 55065 2250 55095 2280
rect 55120 2250 55150 2280
rect 55175 2250 55205 2280
rect 55230 2250 55260 2280
rect 54680 2210 54710 2240
rect 54735 2210 54765 2240
rect 54790 2210 54820 2240
rect 54845 2210 54875 2240
rect 54900 2210 54930 2240
rect 54955 2210 54985 2240
rect 55010 2210 55040 2240
rect 55065 2210 55095 2240
rect 55120 2210 55150 2240
rect 55175 2210 55205 2240
rect 55230 2210 55260 2240
rect 55405 2440 55435 2470
rect 55445 2440 55475 2470
rect 55485 2440 55515 2470
rect 55405 2400 55435 2430
rect 55445 2400 55475 2430
rect 55485 2400 55515 2430
rect 55405 2360 55435 2390
rect 55445 2360 55475 2390
rect 55485 2360 55515 2390
rect 54625 2155 54655 2185
rect 54625 2115 54655 2145
rect 54625 2075 54655 2105
rect 55285 2155 55315 2185
rect 55285 2115 55315 2145
rect 55285 2075 55315 2105
rect 54000 1680 54030 1710
rect 54050 1680 54080 1710
rect 54100 1680 54130 1710
rect 54150 1680 54180 1710
rect 54200 1680 54230 1710
rect 54680 2020 54710 2050
rect 54680 1980 54710 2010
rect 54680 1940 54710 1970
rect 54790 2020 54820 2050
rect 54790 1980 54820 2010
rect 54790 1940 54820 1970
rect 54900 2020 54930 2050
rect 54900 1980 54930 2010
rect 54900 1940 54930 1970
rect 55010 2020 55040 2050
rect 55010 1980 55040 2010
rect 55010 1940 55040 1970
rect 55120 2020 55150 2050
rect 55120 1980 55150 2010
rect 55120 1940 55150 1970
rect 55230 2020 55260 2050
rect 55230 1980 55260 2010
rect 55230 1940 55260 1970
rect 54735 1885 54765 1915
rect 54845 1885 54875 1915
rect 54955 1885 54985 1915
rect 55065 1885 55095 1915
rect 55175 1885 55205 1915
rect 54000 1630 54030 1660
rect 54050 1630 54080 1660
rect 54100 1630 54130 1660
rect 54150 1630 54180 1660
rect 54200 1630 54230 1660
rect 54490 1630 54520 1660
rect 54735 1655 54765 1660
rect 54735 1635 54740 1655
rect 54740 1635 54760 1655
rect 54760 1635 54765 1655
rect 54735 1630 54765 1635
rect 54845 1655 54875 1660
rect 54845 1635 54850 1655
rect 54850 1635 54870 1655
rect 54870 1635 54875 1655
rect 54845 1630 54875 1635
rect 54955 1655 54985 1660
rect 54955 1635 54960 1655
rect 54960 1635 54980 1655
rect 54980 1635 54985 1655
rect 54955 1630 54985 1635
rect 55065 1655 55095 1660
rect 55065 1635 55070 1655
rect 55070 1635 55090 1655
rect 55090 1635 55095 1655
rect 55065 1630 55095 1635
rect 55175 1655 55205 1660
rect 55175 1635 55180 1655
rect 55180 1635 55200 1655
rect 55200 1635 55205 1655
rect 55175 1630 55205 1635
rect 54000 1580 54030 1610
rect 54050 1580 54080 1610
rect 54100 1580 54130 1610
rect 54150 1580 54180 1610
rect 54200 1580 54230 1610
rect 54255 1155 54290 1160
rect 54255 1130 54260 1155
rect 54260 1130 54285 1155
rect 54285 1130 54290 1155
rect 54255 1125 54290 1130
rect 54315 1155 54350 1160
rect 54315 1130 54320 1155
rect 54320 1130 54345 1155
rect 54345 1130 54350 1155
rect 54315 1125 54350 1130
rect 54375 1155 54410 1160
rect 54375 1130 54380 1155
rect 54380 1130 54405 1155
rect 54405 1130 54410 1155
rect 54375 1125 54410 1130
rect 54435 1155 54470 1160
rect 54435 1130 54440 1155
rect 54440 1130 54465 1155
rect 54465 1130 54470 1155
rect 54435 1125 54470 1130
rect 55120 1590 55150 1595
rect 55120 1570 55125 1590
rect 55125 1570 55145 1590
rect 55145 1570 55150 1590
rect 55120 1565 55150 1570
rect 55120 1550 55150 1555
rect 55120 1530 55125 1550
rect 55125 1530 55145 1550
rect 55145 1530 55150 1550
rect 55120 1525 55150 1530
rect 55405 1565 55435 1595
rect 55445 1565 55475 1595
rect 55485 1565 55515 1595
rect 55405 1525 55435 1555
rect 55445 1525 55475 1555
rect 55485 1525 55515 1555
rect 56010 4155 56040 4185
rect 56050 4155 56080 4185
rect 56090 4155 56120 4185
rect 56130 4155 56160 4185
rect 56170 4155 56200 4185
rect 56210 4155 56240 4185
rect 56250 4155 56280 4185
rect 56290 4155 56320 4185
rect 56330 4155 56360 4185
rect 56370 4155 56400 4185
rect 56410 4155 56440 4185
rect 56450 4155 56480 4185
rect 56490 4155 56520 4185
rect 56530 4155 56560 4185
rect 56570 4155 56600 4185
rect 56610 4155 56640 4185
rect 56650 4155 56680 4185
rect 56690 4155 56720 4185
rect 56730 4155 56760 4185
rect 56010 4115 56040 4145
rect 56050 4115 56080 4145
rect 56090 4115 56120 4145
rect 56130 4115 56160 4145
rect 56170 4115 56200 4145
rect 56210 4115 56240 4145
rect 56250 4115 56280 4145
rect 56290 4115 56320 4145
rect 56330 4115 56360 4145
rect 56370 4115 56400 4145
rect 56410 4115 56440 4145
rect 56450 4115 56480 4145
rect 56490 4115 56520 4145
rect 56530 4115 56560 4145
rect 56570 4115 56600 4145
rect 56610 4115 56640 4145
rect 56650 4115 56680 4145
rect 56690 4115 56720 4145
rect 56730 4115 56760 4145
rect 56010 4075 56040 4105
rect 56050 4075 56080 4105
rect 56090 4075 56120 4105
rect 56130 4075 56160 4105
rect 56170 4075 56200 4105
rect 56210 4075 56240 4105
rect 56250 4075 56280 4105
rect 56290 4075 56320 4105
rect 56330 4075 56360 4105
rect 56370 4075 56400 4105
rect 56410 4075 56440 4105
rect 56450 4075 56480 4105
rect 56490 4075 56520 4105
rect 56530 4075 56560 4105
rect 56570 4075 56600 4105
rect 56610 4075 56640 4105
rect 56650 4075 56680 4105
rect 56690 4075 56720 4105
rect 56730 4075 56760 4105
rect 56070 4020 56100 4050
rect 56190 4020 56220 4050
rect 56310 4020 56340 4050
rect 56430 4020 56460 4050
rect 56550 4020 56580 4050
rect 56670 4020 56700 4050
rect 56070 3630 56100 3660
rect 56190 3630 56220 3660
rect 56310 3630 56340 3660
rect 56430 3630 56460 3660
rect 56370 3575 56400 3580
rect 56370 3555 56375 3575
rect 56375 3555 56395 3575
rect 56395 3555 56400 3575
rect 56370 3550 56400 3555
rect 56550 3630 56580 3660
rect 56670 3630 56700 3660
rect 57150 4980 57180 5010
rect 57150 4940 57180 4970
rect 57150 4900 57180 4930
rect 57210 4980 57240 5010
rect 57210 4940 57240 4970
rect 57210 4925 57240 4930
rect 57210 4905 57215 4925
rect 57215 4905 57235 4925
rect 57235 4905 57240 4925
rect 57210 4900 57240 4905
rect 57500 4925 57530 4930
rect 57500 4905 57505 4925
rect 57505 4905 57525 4925
rect 57525 4905 57530 4925
rect 57500 4900 57530 4905
rect 57560 4900 57590 4930
rect 57680 4925 57710 4930
rect 57680 4905 57685 4925
rect 57685 4905 57705 4925
rect 57705 4905 57710 4925
rect 57680 4900 57710 4905
rect 57090 4495 57120 4525
rect 57560 4495 57590 4525
rect 56885 4290 56915 4320
rect 56885 4250 56915 4280
rect 56885 4210 56915 4240
rect 56940 4395 56970 4425
rect 57576 4465 57606 4470
rect 57576 4445 57581 4465
rect 57581 4445 57601 4465
rect 57601 4445 57606 4465
rect 57576 4440 57606 4445
rect 56840 3550 56870 3580
rect 57140 4385 57170 4415
rect 57620 4385 57650 4415
rect 58150 4290 58180 4320
rect 58190 4290 58220 4320
rect 58230 4290 58260 4320
rect 58150 4250 58180 4280
rect 58190 4250 58220 4280
rect 58230 4250 58260 4280
rect 58150 4210 58180 4240
rect 58190 4210 58220 4240
rect 58230 4210 58260 4240
rect 57040 4155 57070 4185
rect 57080 4155 57110 4185
rect 57120 4155 57150 4185
rect 57160 4155 57190 4185
rect 57200 4155 57230 4185
rect 57240 4155 57270 4185
rect 57280 4155 57310 4185
rect 57320 4155 57350 4185
rect 57360 4155 57390 4185
rect 57400 4155 57430 4185
rect 57440 4155 57470 4185
rect 57480 4155 57510 4185
rect 57520 4155 57550 4185
rect 57560 4155 57590 4185
rect 57600 4155 57630 4185
rect 57640 4155 57670 4185
rect 57680 4155 57710 4185
rect 57720 4155 57750 4185
rect 57760 4155 57790 4185
rect 57040 4115 57070 4145
rect 57080 4115 57110 4145
rect 57120 4115 57150 4145
rect 57160 4115 57190 4145
rect 57200 4115 57230 4145
rect 57240 4115 57270 4145
rect 57280 4115 57310 4145
rect 57320 4115 57350 4145
rect 57360 4115 57390 4145
rect 57400 4115 57430 4145
rect 57440 4115 57470 4145
rect 57480 4115 57510 4145
rect 57520 4115 57550 4145
rect 57560 4115 57590 4145
rect 57600 4115 57630 4145
rect 57640 4115 57670 4145
rect 57680 4115 57710 4145
rect 57720 4115 57750 4145
rect 57760 4115 57790 4145
rect 57040 4075 57070 4105
rect 57080 4075 57110 4105
rect 57120 4075 57150 4105
rect 57160 4075 57190 4105
rect 57200 4075 57230 4105
rect 57240 4075 57270 4105
rect 57280 4075 57310 4105
rect 57320 4075 57350 4105
rect 57360 4075 57390 4105
rect 57400 4075 57430 4105
rect 57440 4075 57470 4105
rect 57480 4075 57510 4105
rect 57520 4075 57550 4105
rect 57560 4075 57590 4105
rect 57600 4075 57630 4105
rect 57640 4075 57670 4105
rect 57680 4075 57710 4105
rect 57720 4075 57750 4105
rect 57760 4075 57790 4105
rect 57100 4020 57130 4050
rect 57220 4020 57250 4050
rect 57340 4020 57370 4050
rect 57460 4020 57490 4050
rect 57580 4020 57610 4050
rect 57700 4020 57730 4050
rect 57100 3630 57130 3660
rect 56930 3505 56960 3535
rect 56070 3460 56100 3490
rect 56110 3460 56140 3490
rect 56150 3460 56180 3490
rect 56190 3460 56220 3490
rect 56230 3460 56260 3490
rect 56270 3460 56300 3490
rect 56310 3460 56340 3490
rect 56350 3460 56380 3490
rect 56390 3460 56420 3490
rect 56430 3460 56460 3490
rect 56470 3460 56500 3490
rect 56510 3460 56540 3490
rect 56550 3460 56580 3490
rect 56590 3460 56620 3490
rect 56630 3460 56660 3490
rect 56670 3460 56700 3490
rect 56070 3420 56100 3450
rect 56110 3420 56140 3450
rect 56150 3420 56180 3450
rect 56190 3420 56220 3450
rect 56230 3420 56260 3450
rect 56270 3420 56300 3450
rect 56310 3420 56340 3450
rect 56350 3420 56380 3450
rect 56390 3420 56420 3450
rect 56430 3420 56460 3450
rect 56470 3420 56500 3450
rect 56510 3420 56540 3450
rect 56550 3420 56580 3450
rect 56590 3420 56620 3450
rect 56630 3420 56660 3450
rect 56670 3420 56700 3450
rect 56070 3380 56100 3410
rect 56110 3380 56140 3410
rect 56150 3380 56180 3410
rect 56190 3380 56220 3410
rect 56230 3380 56260 3410
rect 56270 3380 56300 3410
rect 56310 3380 56340 3410
rect 56350 3380 56380 3410
rect 56390 3380 56420 3410
rect 56430 3380 56460 3410
rect 56470 3380 56500 3410
rect 56510 3380 56540 3410
rect 56550 3380 56580 3410
rect 56590 3380 56620 3410
rect 56630 3380 56660 3410
rect 56670 3380 56700 3410
rect 57220 3630 57250 3660
rect 57340 3630 57370 3660
rect 57460 3630 57490 3660
rect 57400 3575 57430 3580
rect 57400 3555 57405 3575
rect 57405 3555 57425 3575
rect 57425 3555 57430 3575
rect 57400 3550 57430 3555
rect 57580 3630 57610 3660
rect 57700 3630 57730 3660
rect 57100 3460 57130 3490
rect 57140 3460 57170 3490
rect 57180 3460 57210 3490
rect 57220 3460 57250 3490
rect 57260 3460 57290 3490
rect 57300 3460 57330 3490
rect 57340 3460 57370 3490
rect 57380 3460 57410 3490
rect 57420 3460 57450 3490
rect 57460 3460 57490 3490
rect 57500 3460 57530 3490
rect 57540 3460 57570 3490
rect 57580 3460 57610 3490
rect 57620 3460 57650 3490
rect 57660 3460 57690 3490
rect 57700 3460 57730 3490
rect 57100 3420 57130 3450
rect 57140 3420 57170 3450
rect 57180 3420 57210 3450
rect 57220 3420 57250 3450
rect 57260 3420 57290 3450
rect 57300 3420 57330 3450
rect 57340 3420 57370 3450
rect 57380 3420 57410 3450
rect 57420 3420 57450 3450
rect 57460 3420 57490 3450
rect 57500 3420 57530 3450
rect 57540 3420 57570 3450
rect 57580 3420 57610 3450
rect 57620 3420 57650 3450
rect 57660 3420 57690 3450
rect 57700 3420 57730 3450
rect 57100 3380 57130 3410
rect 57140 3380 57170 3410
rect 57180 3380 57210 3410
rect 57220 3380 57250 3410
rect 57260 3380 57290 3410
rect 57300 3380 57330 3410
rect 57340 3380 57370 3410
rect 57380 3380 57410 3410
rect 57420 3380 57450 3410
rect 57460 3380 57490 3410
rect 57500 3380 57530 3410
rect 57540 3380 57570 3410
rect 57580 3380 57610 3410
rect 57620 3380 57650 3410
rect 57660 3380 57690 3410
rect 57700 3380 57730 3410
rect 55540 3325 55570 3355
rect 55580 3325 55610 3355
rect 55620 3325 55650 3355
rect 55540 3285 55570 3315
rect 55580 3285 55610 3315
rect 55620 3285 55650 3315
rect 55540 3245 55570 3275
rect 55580 3245 55610 3275
rect 55620 3245 55650 3275
rect 56515 3325 56545 3355
rect 56515 3285 56545 3315
rect 56515 3270 56545 3275
rect 56515 3250 56520 3270
rect 56520 3250 56540 3270
rect 56540 3250 56545 3270
rect 56515 3245 56545 3250
rect 56680 3325 56710 3355
rect 56680 3285 56710 3315
rect 56680 3270 56710 3275
rect 56680 3250 56685 3270
rect 56685 3250 56705 3270
rect 56705 3250 56710 3270
rect 56680 3245 56710 3250
rect 56845 3325 56875 3355
rect 56845 3285 56875 3315
rect 56845 3270 56875 3275
rect 56845 3250 56850 3270
rect 56850 3250 56870 3270
rect 56870 3250 56875 3270
rect 56845 3245 56875 3250
rect 56925 3325 56955 3355
rect 56925 3285 56955 3315
rect 56925 3270 56955 3275
rect 56925 3250 56930 3270
rect 56930 3250 56950 3270
rect 56950 3250 56955 3270
rect 56925 3245 56955 3250
rect 57090 3325 57120 3355
rect 57090 3285 57120 3315
rect 57090 3270 57120 3275
rect 57090 3250 57095 3270
rect 57095 3250 57115 3270
rect 57115 3250 57120 3270
rect 57090 3245 57120 3250
rect 57255 3325 57285 3355
rect 57255 3285 57285 3315
rect 57255 3270 57285 3275
rect 57255 3250 57260 3270
rect 57260 3250 57280 3270
rect 57280 3250 57285 3270
rect 57255 3245 57285 3250
rect 58455 4290 58485 4320
rect 58455 4250 58485 4280
rect 58455 4210 58485 4240
rect 58815 4290 58845 4320
rect 58815 4250 58845 4280
rect 58815 4210 58845 4240
rect 58515 4155 58545 4185
rect 58555 4155 58585 4185
rect 58595 4155 58625 4185
rect 58635 4155 58665 4185
rect 58675 4155 58705 4185
rect 58715 4155 58745 4185
rect 58755 4155 58785 4185
rect 58515 4115 58545 4145
rect 58555 4115 58585 4145
rect 58595 4115 58625 4145
rect 58635 4115 58665 4145
rect 58675 4115 58705 4145
rect 58715 4115 58745 4145
rect 58755 4115 58785 4145
rect 58515 4075 58545 4105
rect 58555 4075 58585 4105
rect 58595 4075 58625 4105
rect 58635 4075 58665 4105
rect 58675 4075 58705 4105
rect 58715 4075 58745 4105
rect 58755 4075 58785 4105
rect 58455 4020 58485 4050
rect 58575 4020 58605 4050
rect 58695 4020 58725 4050
rect 59175 4290 59205 4320
rect 59175 4250 59205 4280
rect 59175 4210 59205 4240
rect 58875 4155 58905 4185
rect 58915 4155 58945 4185
rect 58955 4155 58985 4185
rect 58995 4155 59025 4185
rect 59035 4155 59065 4185
rect 59075 4155 59105 4185
rect 59115 4155 59145 4185
rect 58875 4115 58905 4145
rect 58915 4115 58945 4145
rect 58955 4115 58985 4145
rect 58995 4115 59025 4145
rect 59035 4115 59065 4145
rect 59075 4115 59105 4145
rect 59115 4115 59145 4145
rect 58875 4075 58905 4105
rect 58915 4075 58945 4105
rect 58955 4075 58985 4105
rect 58995 4075 59025 4105
rect 59035 4075 59065 4105
rect 59075 4075 59105 4105
rect 59115 4075 59145 4105
rect 58815 4020 58845 4050
rect 58935 4020 58965 4050
rect 59055 4020 59085 4050
rect 59645 4290 59675 4320
rect 59685 4290 59715 4320
rect 59725 4290 59755 4320
rect 59645 4250 59675 4280
rect 59685 4250 59715 4280
rect 59725 4250 59755 4280
rect 59645 4210 59675 4240
rect 59685 4210 59715 4240
rect 59725 4210 59755 4240
rect 60345 4290 60375 4320
rect 60385 4290 60415 4320
rect 60425 4290 60455 4320
rect 60345 4250 60375 4280
rect 60385 4250 60415 4280
rect 60425 4250 60455 4280
rect 60345 4210 60375 4240
rect 60385 4210 60415 4240
rect 60425 4210 60455 4240
rect 60695 4290 60725 4320
rect 60735 4290 60765 4320
rect 60775 4290 60805 4320
rect 60695 4250 60725 4280
rect 60735 4250 60765 4280
rect 60775 4250 60805 4280
rect 60695 4210 60725 4240
rect 60735 4210 60765 4240
rect 60775 4210 60805 4240
rect 61045 4290 61075 4320
rect 61085 4290 61115 4320
rect 61125 4290 61155 4320
rect 61045 4250 61075 4280
rect 61085 4250 61115 4280
rect 61125 4250 61155 4280
rect 61045 4210 61075 4240
rect 61085 4210 61115 4240
rect 61125 4210 61155 4240
rect 61395 4290 61425 4320
rect 61435 4290 61465 4320
rect 61475 4290 61505 4320
rect 61395 4250 61425 4280
rect 61435 4250 61465 4280
rect 61475 4250 61505 4280
rect 61395 4210 61425 4240
rect 61435 4210 61465 4240
rect 61475 4210 61505 4240
rect 59175 4020 59205 4050
rect 58515 3630 58545 3660
rect 58635 3630 58665 3660
rect 58755 3630 58785 3660
rect 58875 3630 58905 3660
rect 58995 3630 59025 3660
rect 59115 3630 59145 3660
rect 58815 3530 58845 3535
rect 58815 3510 58820 3530
rect 58820 3510 58840 3530
rect 58840 3510 58845 3530
rect 58815 3505 58845 3510
rect 58150 3325 58180 3355
rect 58190 3325 58220 3355
rect 58230 3325 58260 3355
rect 58150 3285 58180 3315
rect 58190 3285 58220 3315
rect 58230 3285 58260 3315
rect 58150 3245 58180 3275
rect 58190 3245 58220 3275
rect 58230 3245 58260 3275
rect 56625 3215 56655 3220
rect 56625 3195 56630 3215
rect 56630 3195 56650 3215
rect 56650 3195 56655 3215
rect 56625 3190 56655 3195
rect 56735 3215 56765 3220
rect 56735 3195 56740 3215
rect 56740 3195 56760 3215
rect 56760 3195 56765 3215
rect 56735 3190 56765 3195
rect 57035 3215 57065 3220
rect 57035 3195 57040 3215
rect 57040 3195 57060 3215
rect 57060 3195 57065 3215
rect 57035 3190 57065 3195
rect 57145 3215 57175 3220
rect 57145 3195 57150 3215
rect 57150 3195 57170 3215
rect 57170 3195 57175 3215
rect 57145 3190 57175 3195
rect 56560 2905 56590 2910
rect 56800 2905 56830 2910
rect 56560 2885 56565 2905
rect 56565 2885 56585 2905
rect 56585 2885 56590 2905
rect 56560 2880 56590 2885
rect 56680 2895 56710 2900
rect 56680 2875 56685 2895
rect 56685 2875 56705 2895
rect 56705 2875 56710 2895
rect 56680 2870 56710 2875
rect 56800 2885 56805 2905
rect 56805 2885 56825 2905
rect 56825 2885 56830 2905
rect 56800 2880 56830 2885
rect 56605 2825 56635 2830
rect 56605 2805 56610 2825
rect 56610 2805 56630 2825
rect 56630 2805 56635 2825
rect 56605 2800 56635 2805
rect 55955 2750 55985 2780
rect 56750 2750 56780 2780
rect 55540 2155 55570 2185
rect 55580 2155 55610 2185
rect 55620 2155 55650 2185
rect 55540 2115 55570 2145
rect 55580 2115 55610 2145
rect 55620 2115 55650 2145
rect 55540 2075 55570 2105
rect 55580 2075 55610 2105
rect 55620 2075 55650 2105
rect 54535 1445 54565 1475
rect 54735 1445 54765 1475
rect 54845 1445 54875 1475
rect 54955 1445 54985 1475
rect 55065 1445 55095 1475
rect 55175 1445 55205 1475
rect 54535 1125 54565 1155
rect 54380 1055 54410 1085
rect 54490 1055 54520 1085
rect 54735 1105 54765 1135
rect 54845 1105 54875 1135
rect 54955 1105 54985 1135
rect 55065 1105 55095 1135
rect 55175 1105 55205 1135
rect 54680 1045 54710 1075
rect 54680 1005 54710 1035
rect 54680 965 54710 995
rect 54790 1045 54820 1075
rect 54790 1005 54820 1035
rect 54790 965 54820 995
rect 54900 1045 54930 1075
rect 54900 1005 54930 1035
rect 54900 965 54930 995
rect 55010 1045 55040 1075
rect 55010 1005 55040 1035
rect 55010 965 55040 995
rect 55120 1045 55150 1075
rect 55120 1005 55150 1035
rect 55120 965 55150 995
rect 55230 1045 55260 1075
rect 55230 1005 55260 1035
rect 55230 965 55260 995
rect 55675 2265 55705 2295
rect 55715 2265 55745 2295
rect 55755 2265 55785 2295
rect 55675 2225 55705 2255
rect 55715 2225 55745 2255
rect 55755 2225 55785 2255
rect 55675 2185 55705 2215
rect 55715 2185 55745 2215
rect 55755 2185 55785 2215
rect 55675 2020 55705 2050
rect 55715 2020 55745 2050
rect 55755 2020 55785 2050
rect 55675 1980 55705 2010
rect 55715 1980 55745 2010
rect 55755 1980 55785 2010
rect 55675 1940 55705 1970
rect 55715 1940 55745 1970
rect 55755 1940 55785 1970
rect 55890 1955 55920 1985
rect 55675 1610 55705 1640
rect 55715 1610 55745 1640
rect 55755 1610 55785 1640
rect 55675 1570 55705 1600
rect 55715 1570 55745 1600
rect 55755 1570 55785 1600
rect 55675 1530 55705 1560
rect 55715 1530 55745 1560
rect 55755 1530 55785 1560
rect 55540 1045 55570 1075
rect 55580 1045 55610 1075
rect 55620 1045 55650 1075
rect 55540 1005 55570 1035
rect 55580 1005 55610 1035
rect 55620 1005 55650 1035
rect 55540 965 55570 995
rect 55580 965 55610 995
rect 55620 965 55650 995
rect 55675 1455 55705 1485
rect 55715 1455 55745 1485
rect 55755 1455 55785 1485
rect 55675 1415 55705 1445
rect 55715 1415 55745 1445
rect 55755 1415 55785 1445
rect 55675 1375 55705 1405
rect 55715 1375 55745 1405
rect 55755 1375 55785 1405
rect 54625 910 54655 940
rect 54625 870 54655 900
rect 54625 830 54655 860
rect 55285 910 55315 940
rect 55285 870 55315 900
rect 55285 830 55315 860
rect 54260 775 54290 805
rect 54325 495 54355 525
rect 55005 520 55035 525
rect 55005 500 55010 520
rect 55010 500 55030 520
rect 55030 500 55035 520
rect 55005 495 55035 500
rect 53995 440 54025 470
rect 54035 440 54065 470
rect 54080 440 54110 470
rect 54120 440 54150 470
rect 54165 440 54195 470
rect 54205 440 54235 470
rect 53995 400 54025 430
rect 54035 400 54065 430
rect 54080 400 54110 430
rect 54120 400 54150 430
rect 54165 400 54195 430
rect 54205 400 54235 430
rect 53995 360 54025 390
rect 54035 360 54065 390
rect 54080 360 54110 390
rect 54120 360 54150 390
rect 54165 360 54195 390
rect 54205 360 54235 390
rect 54390 440 54420 470
rect 54390 400 54420 430
rect 54390 360 54420 390
rect 54755 440 54785 470
rect 54795 440 54825 470
rect 54835 440 54865 470
rect 54875 440 54905 470
rect 54915 440 54945 470
rect 54955 440 54985 470
rect 54995 440 55025 470
rect 55035 440 55065 470
rect 55075 440 55105 470
rect 55115 440 55145 470
rect 55155 440 55185 470
rect 54755 400 54785 430
rect 54795 400 54825 430
rect 54835 400 54865 430
rect 54875 400 54905 430
rect 54915 400 54945 430
rect 54955 400 54985 430
rect 54995 400 55025 430
rect 55035 400 55065 430
rect 55075 400 55105 430
rect 55115 400 55145 430
rect 55155 400 55185 430
rect 54755 360 54785 390
rect 54795 360 54825 390
rect 54835 360 54865 390
rect 54875 360 54905 390
rect 54915 360 54945 390
rect 54955 360 54985 390
rect 54995 360 55025 390
rect 55035 360 55065 390
rect 55075 360 55105 390
rect 55115 360 55145 390
rect 55155 360 55185 390
rect 54325 330 54360 335
rect 54325 305 54330 330
rect 54330 305 54355 330
rect 54355 305 54360 330
rect 54325 300 54360 305
rect 54385 330 54420 335
rect 54385 305 54390 330
rect 54390 305 54415 330
rect 54415 305 54420 330
rect 54385 300 54420 305
rect 54755 -395 54785 -365
rect 54955 -395 54985 -365
rect 53845 -610 53875 -580
rect 53885 -610 53915 -580
rect 53925 -610 53955 -580
rect 53845 -650 53875 -620
rect 53885 -650 53915 -620
rect 53925 -650 53955 -620
rect 53845 -690 53875 -660
rect 53885 -690 53915 -660
rect 53925 -690 53955 -660
rect 54045 -610 54075 -580
rect 54085 -610 54115 -580
rect 54125 -610 54155 -580
rect 54045 -650 54075 -620
rect 54085 -650 54115 -620
rect 54125 -650 54155 -620
rect 54045 -690 54075 -660
rect 54085 -690 54115 -660
rect 54125 -690 54155 -660
rect 54395 -610 54425 -580
rect 54435 -610 54465 -580
rect 54475 -610 54505 -580
rect 54395 -650 54425 -620
rect 54435 -650 54465 -620
rect 54475 -650 54505 -620
rect 54395 -690 54425 -660
rect 54435 -690 54465 -660
rect 54475 -690 54505 -660
rect 54655 -610 54685 -580
rect 54655 -650 54685 -620
rect 54655 -690 54685 -660
rect 54745 -610 54775 -580
rect 54785 -610 54815 -580
rect 54825 -610 54855 -580
rect 54745 -650 54775 -620
rect 54785 -650 54815 -620
rect 54825 -650 54855 -620
rect 54745 -690 54775 -660
rect 54785 -690 54815 -660
rect 54825 -690 54855 -660
rect 55675 -90 55705 -60
rect 55715 -90 55745 -60
rect 55755 -90 55785 -60
rect 55675 -130 55705 -100
rect 55715 -130 55745 -100
rect 55755 -130 55785 -100
rect 55675 -170 55705 -140
rect 55715 -170 55745 -140
rect 55755 -170 55785 -140
rect 57090 2895 57120 2900
rect 57090 2875 57095 2895
rect 57095 2875 57115 2895
rect 57115 2875 57120 2895
rect 57090 2870 57120 2875
rect 57165 2825 57195 2830
rect 57165 2805 57170 2825
rect 57170 2805 57190 2825
rect 57190 2805 57195 2825
rect 57165 2800 57195 2805
rect 57020 2750 57050 2780
rect 56855 2695 56885 2725
rect 56965 2695 56995 2725
rect 57815 2750 57845 2780
rect 56940 2640 56970 2670
rect 57215 2640 57245 2670
rect 56855 2610 56885 2615
rect 56855 2590 56860 2610
rect 56860 2590 56880 2610
rect 56880 2590 56885 2610
rect 56855 2585 56885 2590
rect 56090 2440 56120 2470
rect 56145 2440 56175 2470
rect 56200 2440 56230 2470
rect 56255 2440 56285 2470
rect 56310 2440 56340 2470
rect 56365 2440 56395 2470
rect 56420 2440 56450 2470
rect 56475 2440 56505 2470
rect 56530 2440 56560 2470
rect 56585 2440 56615 2470
rect 56640 2440 56670 2470
rect 56090 2400 56120 2430
rect 56145 2400 56175 2430
rect 56200 2400 56230 2430
rect 56255 2400 56285 2430
rect 56310 2400 56340 2430
rect 56365 2400 56395 2430
rect 56420 2400 56450 2430
rect 56475 2400 56505 2430
rect 56530 2400 56560 2430
rect 56585 2400 56615 2430
rect 56640 2400 56670 2430
rect 56090 2360 56120 2390
rect 56145 2360 56175 2390
rect 56200 2360 56230 2390
rect 56255 2360 56285 2390
rect 56310 2360 56340 2390
rect 56365 2360 56395 2390
rect 56420 2360 56450 2390
rect 56475 2360 56505 2390
rect 56530 2360 56560 2390
rect 56585 2360 56615 2390
rect 56640 2360 56670 2390
rect 56040 1980 56070 1985
rect 56040 1960 56045 1980
rect 56045 1960 56065 1980
rect 56065 1960 56070 1980
rect 56040 1955 56070 1960
rect 56145 1945 56175 1975
rect 56090 1900 56120 1930
rect 56255 1945 56285 1975
rect 56200 1900 56230 1930
rect 56145 1710 56175 1740
rect 56090 1665 56120 1695
rect 56035 1610 56065 1640
rect 56035 1570 56065 1600
rect 56035 1530 56065 1560
rect 56365 1945 56395 1975
rect 56310 1900 56340 1930
rect 56255 1710 56285 1740
rect 56200 1665 56230 1695
rect 56040 1290 56070 1295
rect 56040 1270 56045 1290
rect 56045 1270 56065 1290
rect 56065 1270 56070 1290
rect 56090 1275 56120 1305
rect 56145 1285 56175 1315
rect 56475 1945 56505 1975
rect 56420 1900 56450 1930
rect 56365 1710 56395 1740
rect 56310 1665 56340 1695
rect 56200 1275 56230 1305
rect 56255 1285 56285 1315
rect 56585 1945 56615 1975
rect 56530 1900 56560 1930
rect 56475 1710 56505 1740
rect 56420 1665 56450 1695
rect 56310 1275 56340 1305
rect 56365 1285 56395 1315
rect 57130 2440 57160 2470
rect 57185 2440 57215 2470
rect 57240 2440 57270 2470
rect 57295 2440 57325 2470
rect 57350 2440 57380 2470
rect 57405 2440 57435 2470
rect 57460 2440 57490 2470
rect 57515 2440 57545 2470
rect 57570 2440 57600 2470
rect 57625 2440 57655 2470
rect 57680 2440 57710 2470
rect 57130 2400 57160 2430
rect 57185 2400 57215 2430
rect 57240 2400 57270 2430
rect 57295 2400 57325 2430
rect 57350 2400 57380 2430
rect 57405 2400 57435 2430
rect 57460 2400 57490 2430
rect 57515 2400 57545 2430
rect 57570 2400 57600 2430
rect 57625 2400 57655 2430
rect 57680 2400 57710 2430
rect 57130 2360 57160 2390
rect 57185 2360 57215 2390
rect 57240 2360 57270 2390
rect 57295 2360 57325 2390
rect 57350 2360 57380 2390
rect 57405 2360 57435 2390
rect 57460 2360 57490 2390
rect 57515 2360 57545 2390
rect 57570 2360 57600 2390
rect 57625 2360 57655 2390
rect 57680 2360 57710 2390
rect 56775 2290 56805 2295
rect 56775 2270 56780 2290
rect 56780 2270 56800 2290
rect 56800 2270 56805 2290
rect 56775 2265 56805 2270
rect 56775 2225 56805 2255
rect 56775 2185 56805 2215
rect 56885 2265 56915 2295
rect 56885 2225 56915 2255
rect 56885 2185 56915 2215
rect 56995 2290 57025 2295
rect 56995 2270 57000 2290
rect 57000 2270 57020 2290
rect 57020 2270 57025 2290
rect 56995 2265 57025 2270
rect 56995 2225 57025 2255
rect 56995 2185 57025 2215
rect 56690 1980 56720 1985
rect 56690 1960 56695 1980
rect 56695 1960 56715 1980
rect 56715 1960 56720 1980
rect 56690 1955 56720 1960
rect 57080 1980 57110 1985
rect 57080 1960 57085 1980
rect 57085 1960 57105 1980
rect 57105 1960 57110 1980
rect 57080 1955 57110 1960
rect 56640 1900 56670 1930
rect 57185 1945 57215 1975
rect 57130 1900 57160 1930
rect 56585 1710 56615 1740
rect 56530 1665 56560 1695
rect 56420 1275 56450 1305
rect 56475 1285 56505 1315
rect 56640 1665 56670 1695
rect 57295 1945 57325 1975
rect 57240 1900 57270 1930
rect 57185 1710 57215 1740
rect 57130 1665 57160 1695
rect 56695 1610 56725 1640
rect 56695 1570 56725 1600
rect 56695 1530 56725 1560
rect 57075 1610 57105 1640
rect 57075 1570 57105 1600
rect 57075 1530 57105 1560
rect 56885 1455 56915 1485
rect 56885 1415 56915 1445
rect 56885 1375 56915 1405
rect 56530 1275 56560 1305
rect 56585 1285 56615 1315
rect 56640 1275 56670 1305
rect 56690 1300 56720 1305
rect 56690 1280 56695 1300
rect 56695 1280 56715 1300
rect 56715 1280 56720 1300
rect 56690 1275 56720 1280
rect 56840 1300 56870 1305
rect 56840 1280 56845 1300
rect 56845 1280 56865 1300
rect 56865 1280 56870 1300
rect 56840 1275 56870 1280
rect 56040 1265 56070 1270
rect 56145 1230 56175 1260
rect 56090 1035 56120 1065
rect 56255 1230 56285 1260
rect 56200 1035 56230 1065
rect 56365 1230 56395 1260
rect 56310 1035 56340 1065
rect 56475 1230 56505 1260
rect 56420 1035 56450 1065
rect 56585 1230 56615 1260
rect 56530 1035 56560 1065
rect 56640 1035 56670 1065
rect 57405 1945 57435 1975
rect 57350 1900 57380 1930
rect 57295 1710 57325 1740
rect 57240 1665 57270 1695
rect 56930 1300 56960 1305
rect 56930 1280 56935 1300
rect 56935 1280 56955 1300
rect 56955 1280 56960 1300
rect 56930 1275 56960 1280
rect 57080 1300 57110 1305
rect 57080 1280 57085 1300
rect 57085 1280 57105 1300
rect 57105 1280 57110 1300
rect 57080 1275 57110 1280
rect 57130 1275 57160 1305
rect 57185 1285 57215 1315
rect 57515 1945 57545 1975
rect 57460 1900 57490 1930
rect 57405 1710 57435 1740
rect 57350 1665 57380 1695
rect 57240 1275 57270 1305
rect 57295 1285 57325 1315
rect 57625 1945 57655 1975
rect 57570 1900 57600 1930
rect 57515 1710 57545 1740
rect 57460 1665 57490 1695
rect 57350 1275 57380 1305
rect 57405 1285 57435 1315
rect 57730 1980 57760 1985
rect 57730 1960 57735 1980
rect 57735 1960 57755 1980
rect 57755 1960 57760 1980
rect 57730 1955 57760 1960
rect 57680 1900 57710 1930
rect 57625 1710 57655 1740
rect 57570 1665 57600 1695
rect 57460 1275 57490 1305
rect 57515 1285 57545 1315
rect 57680 1665 57710 1695
rect 57735 1610 57765 1640
rect 57735 1570 57765 1600
rect 57735 1530 57765 1560
rect 57570 1275 57600 1305
rect 57625 1285 57655 1315
rect 57680 1275 57710 1305
rect 57730 1290 57760 1295
rect 57730 1270 57735 1290
rect 57735 1270 57755 1290
rect 57755 1270 57760 1290
rect 57185 1230 57215 1260
rect 56830 1035 56860 1065
rect 56145 965 56175 995
rect 56255 965 56285 995
rect 56365 965 56395 995
rect 56475 965 56505 995
rect 56585 965 56615 995
rect 56035 910 56065 940
rect 56035 870 56065 900
rect 56035 830 56065 860
rect 55945 775 55975 805
rect 56735 910 56765 940
rect 56735 870 56765 900
rect 56735 830 56765 860
rect 56445 450 56475 480
rect 56555 450 56585 480
rect 56665 450 56695 480
rect 56775 450 56805 480
rect 56940 1035 56970 1065
rect 56885 450 56915 480
rect 57130 1035 57160 1065
rect 57295 1230 57325 1260
rect 57240 1035 57270 1065
rect 57405 1230 57435 1260
rect 57350 1035 57380 1065
rect 57515 1230 57545 1260
rect 57460 1035 57490 1065
rect 57625 1230 57655 1260
rect 57570 1035 57600 1065
rect 57730 1265 57760 1270
rect 57680 1035 57710 1065
rect 57185 965 57215 995
rect 57295 965 57325 995
rect 57035 910 57065 940
rect 57035 870 57065 900
rect 57035 830 57065 860
rect 56995 450 57025 480
rect 57405 965 57435 995
rect 57515 965 57545 995
rect 57625 965 57655 995
rect 57735 910 57765 940
rect 57735 870 57765 900
rect 57735 830 57765 860
rect 57870 2640 57900 2670
rect 57825 775 57855 805
rect 57105 450 57135 480
rect 57215 450 57245 480
rect 57325 450 57355 480
rect 57435 450 57465 480
rect 56225 145 56255 150
rect 56225 125 56230 145
rect 56230 125 56250 145
rect 56250 125 56255 145
rect 56225 120 56255 125
rect 55890 -280 55920 -250
rect 55155 -395 55185 -365
rect 56280 120 56310 150
rect 56390 120 56420 150
rect 56500 120 56530 150
rect 56610 120 56640 150
rect 56720 120 56750 150
rect 56830 120 56860 150
rect 56940 120 56970 150
rect 57050 120 57080 150
rect 57160 120 57190 150
rect 57270 120 57300 150
rect 57380 120 57410 150
rect 57490 145 57520 150
rect 57490 125 57495 145
rect 57495 125 57515 145
rect 57515 125 57520 145
rect 57490 120 57520 125
rect 56445 65 56475 95
rect 56555 65 56585 95
rect 56665 65 56695 95
rect 56775 65 56805 95
rect 56885 65 56915 95
rect 56995 65 57025 95
rect 57105 65 57135 95
rect 57215 65 57245 95
rect 57325 65 57355 95
rect 57435 65 57465 95
rect 56335 -90 56365 -60
rect 56335 -130 56365 -100
rect 56335 -170 56365 -140
rect 56545 -225 56575 -195
rect 56655 -225 56685 -195
rect 56875 -225 56905 -195
rect 56490 -280 56520 -250
rect 56600 -255 56630 -250
rect 56600 -275 56605 -255
rect 56605 -275 56625 -255
rect 56625 -275 56630 -255
rect 56600 -280 56630 -275
rect 56490 -500 56520 -470
rect 56710 -280 56740 -250
rect 56600 -500 56630 -470
rect 56925 -255 56955 -250
rect 56925 -275 56930 -255
rect 56930 -275 56950 -255
rect 56950 -275 56955 -255
rect 56925 -280 56955 -275
rect 57045 -255 57075 -250
rect 57045 -275 57050 -255
rect 57050 -275 57070 -255
rect 57070 -275 57075 -255
rect 57045 -280 57075 -275
rect 57165 -255 57195 -250
rect 57165 -275 57170 -255
rect 57170 -275 57190 -255
rect 57190 -275 57195 -255
rect 57165 -280 57195 -275
rect 56710 -500 56740 -470
rect 56545 -555 56575 -525
rect 56655 -555 56685 -525
rect 57420 35 57450 40
rect 57420 15 57425 35
rect 57425 15 57445 35
rect 57445 15 57450 35
rect 57420 10 57450 15
rect 56925 -475 56955 -470
rect 56925 -495 56930 -475
rect 56930 -495 56950 -475
rect 56950 -495 56955 -475
rect 56925 -500 56955 -495
rect 57045 -475 57075 -470
rect 57045 -495 57050 -475
rect 57050 -495 57070 -475
rect 57070 -495 57075 -475
rect 57045 -500 57075 -495
rect 57165 -475 57195 -470
rect 57165 -495 57170 -475
rect 57170 -495 57190 -475
rect 57190 -495 57195 -475
rect 57165 -500 57195 -495
rect 56875 -555 56905 -525
rect 55095 -610 55125 -580
rect 55135 -610 55165 -580
rect 55175 -610 55205 -580
rect 55095 -650 55125 -620
rect 55135 -650 55165 -620
rect 55175 -650 55205 -620
rect 55095 -690 55125 -660
rect 55135 -690 55165 -660
rect 55175 -690 55205 -660
rect 55255 -610 55285 -580
rect 55255 -650 55285 -620
rect 55255 -690 55285 -660
rect 55445 -610 55475 -580
rect 55485 -610 55515 -580
rect 55525 -610 55555 -580
rect 55445 -650 55475 -620
rect 55485 -650 55515 -620
rect 55525 -650 55555 -620
rect 55445 -690 55475 -660
rect 55485 -690 55515 -660
rect 55525 -690 55555 -660
rect 55795 -610 55825 -580
rect 55835 -610 55865 -580
rect 55875 -610 55905 -580
rect 55795 -650 55825 -620
rect 55835 -650 55865 -620
rect 55875 -650 55905 -620
rect 55795 -690 55825 -660
rect 55835 -690 55865 -660
rect 55875 -690 55905 -660
rect 56145 -610 56175 -580
rect 56185 -610 56215 -580
rect 56225 -610 56255 -580
rect 56145 -650 56175 -620
rect 56185 -650 56215 -620
rect 56225 -650 56255 -620
rect 56145 -690 56175 -660
rect 56185 -690 56215 -660
rect 56225 -690 56255 -660
rect 56435 -610 56465 -580
rect 56435 -650 56465 -620
rect 56435 -690 56465 -660
rect 56495 -610 56525 -580
rect 56535 -610 56565 -580
rect 56575 -610 56605 -580
rect 56495 -650 56525 -620
rect 56535 -650 56565 -620
rect 56575 -650 56605 -620
rect 56495 -690 56525 -660
rect 56535 -690 56565 -660
rect 56575 -690 56605 -660
rect 56765 -610 56795 -580
rect 56765 -650 56795 -620
rect 56765 -690 56795 -660
rect 56845 -610 56875 -580
rect 56885 -610 56915 -580
rect 56925 -610 56955 -580
rect 56845 -650 56875 -620
rect 56885 -650 56915 -620
rect 56925 -650 56955 -620
rect 56845 -690 56875 -660
rect 56885 -690 56915 -660
rect 56925 -690 56955 -660
rect 57195 -610 57225 -580
rect 57235 -610 57265 -580
rect 57275 -610 57305 -580
rect 57195 -650 57225 -620
rect 57235 -650 57265 -620
rect 57275 -650 57305 -620
rect 57195 -690 57225 -660
rect 57235 -690 57265 -660
rect 57275 -690 57305 -660
rect 58015 2265 58045 2295
rect 58055 2265 58085 2295
rect 58095 2265 58125 2295
rect 58015 2225 58045 2255
rect 58055 2225 58085 2255
rect 58095 2225 58125 2255
rect 58015 2185 58045 2215
rect 58055 2185 58085 2215
rect 58095 2185 58125 2215
rect 58015 2020 58045 2050
rect 58055 2020 58085 2050
rect 58095 2020 58125 2050
rect 58015 1980 58045 2010
rect 58055 1980 58085 2010
rect 58095 1980 58125 2010
rect 58015 1940 58045 1970
rect 58055 1940 58085 1970
rect 58095 1940 58125 1970
rect 58015 1610 58045 1640
rect 58055 1610 58085 1640
rect 58095 1610 58125 1640
rect 58015 1570 58045 1600
rect 58055 1570 58085 1600
rect 58095 1570 58125 1600
rect 58015 1530 58045 1560
rect 58055 1530 58085 1560
rect 58095 1530 58125 1560
rect 58150 2155 58180 2185
rect 58190 2155 58220 2185
rect 58230 2155 58260 2185
rect 58150 2115 58180 2145
rect 58190 2115 58220 2145
rect 58230 2115 58260 2145
rect 58150 2075 58180 2105
rect 58190 2075 58220 2105
rect 58230 2075 58260 2105
rect 58015 1455 58045 1485
rect 58055 1455 58085 1485
rect 58095 1455 58125 1485
rect 58015 1415 58045 1445
rect 58055 1415 58085 1445
rect 58095 1415 58125 1445
rect 58015 1375 58045 1405
rect 58055 1375 58085 1405
rect 58095 1375 58125 1405
rect 57870 10 57900 40
rect 58285 3460 58315 3490
rect 58325 3460 58355 3490
rect 58365 3460 58395 3490
rect 58285 3420 58315 3450
rect 58325 3420 58355 3450
rect 58365 3420 58395 3450
rect 58285 3380 58315 3410
rect 58325 3380 58355 3410
rect 58365 3380 58395 3410
rect 58485 3325 58515 3355
rect 58485 3285 58515 3315
rect 58485 3245 58515 3275
rect 58595 3325 58625 3355
rect 58595 3285 58625 3315
rect 58595 3245 58625 3275
rect 58705 3325 58735 3355
rect 58705 3285 58735 3315
rect 58705 3245 58735 3275
rect 58815 3325 58845 3355
rect 58815 3285 58845 3315
rect 58815 3245 58845 3275
rect 58925 3325 58955 3355
rect 58925 3285 58955 3315
rect 58925 3245 58955 3275
rect 59035 3325 59065 3355
rect 59035 3285 59065 3315
rect 59035 3245 59065 3275
rect 59145 3325 59175 3355
rect 59145 3285 59175 3315
rect 59145 3245 59175 3275
rect 59510 3345 59540 3375
rect 58540 3160 58570 3190
rect 58650 3160 58680 3190
rect 58760 3160 58790 3190
rect 58870 3160 58900 3190
rect 58980 3160 59010 3190
rect 59090 3160 59120 3190
rect 58285 2440 58315 2470
rect 58325 2440 58355 2470
rect 58365 2440 58395 2470
rect 58285 2400 58315 2430
rect 58325 2400 58355 2430
rect 58365 2400 58395 2430
rect 58285 2360 58315 2390
rect 58325 2360 58355 2390
rect 58365 2360 58395 2390
rect 58540 2520 58570 2550
rect 58650 2520 58680 2550
rect 58760 2520 58790 2550
rect 58870 2520 58900 2550
rect 58815 2465 58845 2470
rect 58815 2445 58820 2465
rect 58820 2445 58840 2465
rect 58840 2445 58845 2465
rect 58815 2440 58845 2445
rect 58815 2425 58845 2430
rect 58815 2405 58820 2425
rect 58820 2405 58840 2425
rect 58840 2405 58845 2425
rect 58815 2400 58845 2405
rect 58815 2385 58845 2390
rect 58815 2365 58820 2385
rect 58820 2365 58840 2385
rect 58840 2365 58845 2385
rect 58815 2360 58845 2365
rect 58980 2520 59010 2550
rect 59090 2520 59120 2550
rect 59470 2440 59500 2470
rect 59510 2440 59540 2470
rect 59550 2440 59580 2470
rect 59470 2400 59500 2430
rect 59510 2400 59540 2430
rect 59550 2400 59580 2430
rect 59470 2360 59500 2390
rect 59510 2360 59540 2390
rect 59550 2360 59580 2390
rect 58540 2290 58570 2320
rect 58595 2290 58625 2320
rect 58650 2290 58680 2320
rect 58705 2290 58735 2320
rect 58760 2290 58790 2320
rect 58815 2290 58845 2320
rect 58870 2290 58900 2320
rect 58925 2290 58955 2320
rect 58980 2290 59010 2320
rect 59035 2290 59065 2320
rect 59090 2290 59120 2320
rect 58540 2250 58570 2280
rect 58595 2250 58625 2280
rect 58650 2250 58680 2280
rect 58705 2250 58735 2280
rect 58760 2250 58790 2280
rect 58815 2250 58845 2280
rect 58870 2250 58900 2280
rect 58925 2250 58955 2280
rect 58980 2250 59010 2280
rect 59035 2250 59065 2280
rect 59090 2250 59120 2280
rect 58540 2210 58570 2240
rect 58595 2210 58625 2240
rect 58650 2210 58680 2240
rect 58705 2210 58735 2240
rect 58760 2210 58790 2240
rect 58815 2210 58845 2240
rect 58870 2210 58900 2240
rect 58925 2210 58955 2240
rect 58980 2210 59010 2240
rect 59035 2210 59065 2240
rect 59090 2210 59120 2240
rect 59565 2290 59595 2320
rect 59605 2290 59635 2320
rect 59650 2290 59680 2320
rect 59690 2290 59720 2320
rect 59735 2290 59765 2320
rect 59775 2290 59805 2320
rect 59565 2250 59595 2280
rect 59605 2250 59635 2280
rect 59650 2250 59680 2280
rect 59690 2250 59720 2280
rect 59735 2250 59765 2280
rect 59775 2250 59805 2280
rect 59565 2210 59595 2240
rect 59605 2210 59635 2240
rect 59650 2210 59680 2240
rect 59690 2210 59720 2240
rect 59735 2210 59765 2240
rect 59775 2210 59805 2240
rect 58485 2155 58515 2185
rect 58485 2115 58515 2145
rect 58485 2075 58515 2105
rect 59145 2155 59175 2185
rect 59145 2115 59175 2145
rect 59145 2075 59175 2105
rect 58540 2020 58570 2050
rect 58540 1980 58570 2010
rect 58540 1940 58570 1970
rect 58650 2020 58680 2050
rect 58650 1980 58680 2010
rect 58650 1940 58680 1970
rect 58760 2020 58790 2050
rect 58760 1980 58790 2010
rect 58760 1940 58790 1970
rect 58870 2020 58900 2050
rect 58870 1980 58900 2010
rect 58870 1940 58900 1970
rect 58980 2020 59010 2050
rect 58980 1980 59010 2010
rect 58980 1940 59010 1970
rect 59090 2020 59120 2050
rect 59090 1980 59120 2010
rect 59090 1940 59120 1970
rect 58595 1885 58625 1915
rect 58705 1885 58735 1915
rect 58815 1885 58845 1915
rect 58925 1885 58955 1915
rect 59035 1885 59065 1915
rect 59570 1680 59600 1710
rect 59620 1680 59650 1710
rect 59670 1680 59700 1710
rect 59720 1680 59750 1710
rect 59770 1680 59800 1710
rect 58595 1655 58625 1660
rect 58595 1635 58600 1655
rect 58600 1635 58620 1655
rect 58620 1635 58625 1655
rect 58595 1630 58625 1635
rect 58705 1655 58735 1660
rect 58705 1635 58710 1655
rect 58710 1635 58730 1655
rect 58730 1635 58735 1655
rect 58705 1630 58735 1635
rect 58815 1655 58845 1660
rect 58815 1635 58820 1655
rect 58820 1635 58840 1655
rect 58840 1635 58845 1655
rect 58815 1630 58845 1635
rect 58925 1655 58955 1660
rect 58925 1635 58930 1655
rect 58930 1635 58950 1655
rect 58950 1635 58955 1655
rect 58925 1630 58955 1635
rect 59035 1655 59065 1660
rect 59035 1635 59040 1655
rect 59040 1635 59060 1655
rect 59060 1635 59065 1655
rect 59035 1630 59065 1635
rect 59280 1630 59310 1660
rect 59570 1630 59600 1660
rect 59620 1630 59650 1660
rect 59670 1630 59700 1660
rect 59720 1630 59750 1660
rect 59770 1630 59800 1660
rect 58285 1565 58315 1595
rect 58325 1565 58355 1595
rect 58365 1565 58395 1595
rect 58285 1525 58315 1555
rect 58325 1525 58355 1555
rect 58365 1525 58395 1555
rect 58650 1590 58680 1595
rect 58650 1570 58655 1590
rect 58655 1570 58675 1590
rect 58675 1570 58680 1590
rect 58650 1565 58680 1570
rect 58650 1550 58680 1555
rect 58650 1530 58655 1550
rect 58655 1530 58675 1550
rect 58675 1530 58680 1550
rect 58650 1525 58680 1530
rect 58595 1445 58625 1475
rect 58705 1445 58735 1475
rect 58815 1445 58845 1475
rect 58925 1445 58955 1475
rect 59035 1445 59065 1475
rect 59235 1445 59265 1475
rect 58150 1050 58180 1080
rect 58190 1050 58220 1080
rect 58230 1050 58260 1080
rect 58150 1010 58180 1040
rect 58190 1010 58220 1040
rect 58230 1010 58260 1040
rect 58150 970 58180 1000
rect 58190 970 58220 1000
rect 58230 970 58260 1000
rect 58595 1105 58625 1135
rect 58705 1105 58735 1135
rect 58815 1105 58845 1135
rect 58925 1105 58955 1135
rect 59035 1105 59065 1135
rect 59235 1125 59265 1155
rect 58540 1050 58570 1080
rect 58540 1010 58570 1040
rect 58540 970 58570 1000
rect 58650 1050 58680 1080
rect 58650 1010 58680 1040
rect 58650 970 58680 1000
rect 58760 1050 58790 1080
rect 58760 1010 58790 1040
rect 58760 970 58790 1000
rect 58870 1050 58900 1080
rect 58870 1010 58900 1040
rect 58870 970 58900 1000
rect 58980 1050 59010 1080
rect 58980 1010 59010 1040
rect 58980 970 59010 1000
rect 59090 1050 59120 1080
rect 59090 1010 59120 1040
rect 59090 970 59120 1000
rect 59570 1580 59600 1610
rect 59620 1580 59650 1610
rect 59670 1580 59700 1610
rect 59720 1580 59750 1610
rect 59770 1580 59800 1610
rect 59330 1155 59365 1160
rect 59330 1130 59335 1155
rect 59335 1130 59360 1155
rect 59360 1130 59365 1155
rect 59330 1125 59365 1130
rect 59390 1155 59425 1160
rect 59390 1130 59395 1155
rect 59395 1130 59420 1155
rect 59420 1130 59425 1155
rect 59390 1125 59425 1130
rect 59450 1155 59485 1160
rect 59450 1130 59455 1155
rect 59455 1130 59480 1155
rect 59480 1130 59485 1155
rect 59450 1125 59485 1130
rect 59510 1155 59545 1160
rect 59510 1130 59515 1155
rect 59515 1130 59540 1155
rect 59540 1130 59545 1155
rect 59510 1125 59545 1130
rect 59280 1055 59310 1085
rect 59390 1055 59420 1085
rect 58485 910 58515 940
rect 58485 870 58515 900
rect 58485 830 58515 860
rect 59145 910 59175 940
rect 59145 870 59175 900
rect 59145 830 59175 860
rect 59510 775 59540 805
rect 58765 520 58795 525
rect 58765 500 58770 520
rect 58770 500 58790 520
rect 58790 500 58795 520
rect 58765 495 58795 500
rect 59445 495 59475 525
rect 58615 440 58645 470
rect 58655 440 58685 470
rect 58695 440 58725 470
rect 58735 440 58765 470
rect 58775 440 58805 470
rect 58815 440 58845 470
rect 58855 440 58885 470
rect 58895 440 58925 470
rect 58935 440 58965 470
rect 58975 440 59005 470
rect 59015 440 59045 470
rect 58615 400 58645 430
rect 58655 400 58685 430
rect 58695 400 58725 430
rect 58735 400 58765 430
rect 58775 400 58805 430
rect 58815 400 58845 430
rect 58855 400 58885 430
rect 58895 400 58925 430
rect 58935 400 58965 430
rect 58975 400 59005 430
rect 59015 400 59045 430
rect 58615 360 58645 390
rect 58655 360 58685 390
rect 58695 360 58725 390
rect 58735 360 58765 390
rect 58775 360 58805 390
rect 58815 360 58845 390
rect 58855 360 58885 390
rect 58895 360 58925 390
rect 58935 360 58965 390
rect 58975 360 59005 390
rect 59015 360 59045 390
rect 59380 440 59410 470
rect 59380 400 59410 430
rect 59380 360 59410 390
rect 58015 -90 58045 -60
rect 58055 -90 58085 -60
rect 58095 -90 58125 -60
rect 58015 -130 58045 -100
rect 58055 -130 58085 -100
rect 58095 -130 58125 -100
rect 58015 -170 58045 -140
rect 58055 -170 58085 -140
rect 58095 -170 58125 -140
rect 58615 -395 58645 -365
rect 58815 -395 58845 -365
rect 57490 -610 57520 -580
rect 57490 -650 57520 -620
rect 57490 -690 57520 -660
rect 57545 -610 57575 -580
rect 57585 -610 57615 -580
rect 57625 -610 57655 -580
rect 57545 -650 57575 -620
rect 57585 -650 57615 -620
rect 57625 -650 57655 -620
rect 57545 -690 57575 -660
rect 57585 -690 57615 -660
rect 57625 -690 57655 -660
rect 57895 -610 57925 -580
rect 57935 -610 57965 -580
rect 57975 -610 58005 -580
rect 57895 -650 57925 -620
rect 57935 -650 57965 -620
rect 57975 -650 58005 -620
rect 57895 -690 57925 -660
rect 57935 -690 57965 -660
rect 57975 -690 58005 -660
rect 58245 -610 58275 -580
rect 58285 -610 58315 -580
rect 58325 -610 58355 -580
rect 58245 -650 58275 -620
rect 58285 -650 58315 -620
rect 58325 -650 58355 -620
rect 58245 -690 58275 -660
rect 58285 -690 58315 -660
rect 58325 -690 58355 -660
rect 58515 -610 58545 -580
rect 58515 -650 58545 -620
rect 58515 -690 58545 -660
rect 58595 -610 58625 -580
rect 58635 -610 58665 -580
rect 58675 -610 58705 -580
rect 58595 -650 58625 -620
rect 58635 -650 58665 -620
rect 58675 -650 58705 -620
rect 58595 -690 58625 -660
rect 58635 -690 58665 -660
rect 58675 -690 58705 -660
rect 59565 440 59595 470
rect 59605 440 59635 470
rect 59650 440 59680 470
rect 59690 440 59720 470
rect 59735 440 59765 470
rect 59775 440 59805 470
rect 59565 400 59595 430
rect 59605 400 59635 430
rect 59650 400 59680 430
rect 59690 400 59720 430
rect 59735 400 59765 430
rect 59775 400 59805 430
rect 59565 360 59595 390
rect 59605 360 59635 390
rect 59650 360 59680 390
rect 59690 360 59720 390
rect 59735 360 59765 390
rect 59775 360 59805 390
rect 59845 2020 59875 2050
rect 59885 2020 59915 2050
rect 59925 2020 59955 2050
rect 59845 1980 59875 2010
rect 59885 1980 59915 2010
rect 59925 1980 59955 2010
rect 59845 1940 59875 1970
rect 59885 1940 59915 1970
rect 59925 1940 59955 1970
rect 59845 910 59875 940
rect 59885 910 59915 940
rect 59925 910 59955 940
rect 59845 870 59875 900
rect 59885 870 59915 900
rect 59925 870 59955 900
rect 59845 830 59875 860
rect 59885 830 59915 860
rect 59925 830 59955 860
rect 59380 330 59415 335
rect 59380 305 59385 330
rect 59385 305 59410 330
rect 59410 305 59415 330
rect 59380 300 59415 305
rect 59440 330 59475 335
rect 59440 305 59445 330
rect 59445 305 59470 330
rect 59470 305 59475 330
rect 59440 300 59475 305
rect 59015 -395 59045 -365
rect 58945 -610 58975 -580
rect 58985 -610 59015 -580
rect 59025 -610 59055 -580
rect 58945 -650 58975 -620
rect 58985 -650 59015 -620
rect 59025 -650 59055 -620
rect 58945 -690 58975 -660
rect 58985 -690 59015 -660
rect 59025 -690 59055 -660
rect 59115 -610 59145 -580
rect 59115 -650 59145 -620
rect 59115 -690 59145 -660
rect 59375 -610 59405 -580
rect 59415 -610 59445 -580
rect 59455 -610 59485 -580
rect 59375 -650 59405 -620
rect 59415 -650 59445 -620
rect 59455 -650 59485 -620
rect 59375 -690 59405 -660
rect 59415 -690 59445 -660
rect 59455 -690 59485 -660
rect 59645 -610 59675 -580
rect 59685 -610 59715 -580
rect 59725 -610 59755 -580
rect 59645 -650 59675 -620
rect 59685 -650 59715 -620
rect 59725 -650 59755 -620
rect 59645 -690 59675 -660
rect 59685 -690 59715 -660
rect 59725 -690 59755 -660
rect 59845 -610 59875 -580
rect 59885 -610 59915 -580
rect 59925 -610 59955 -580
rect 59845 -650 59875 -620
rect 59885 -650 59915 -620
rect 59925 -650 59955 -620
rect 59845 -690 59875 -660
rect 59885 -690 59915 -660
rect 59925 -690 59955 -660
rect 59995 -610 60025 -580
rect 60035 -610 60065 -580
rect 60075 -610 60105 -580
rect 59995 -650 60025 -620
rect 60035 -650 60065 -620
rect 60075 -650 60105 -620
rect 59995 -690 60025 -660
rect 60035 -690 60065 -660
rect 60075 -690 60105 -660
rect 60345 -610 60375 -580
rect 60385 -610 60415 -580
rect 60425 -610 60455 -580
rect 60345 -650 60375 -620
rect 60385 -650 60415 -620
rect 60425 -650 60455 -620
rect 60345 -690 60375 -660
rect 60385 -690 60415 -660
rect 60425 -690 60455 -660
rect 60695 -610 60725 -580
rect 60735 -610 60765 -580
rect 60775 -610 60805 -580
rect 60695 -650 60725 -620
rect 60735 -650 60765 -620
rect 60775 -650 60805 -620
rect 60695 -690 60725 -660
rect 60735 -690 60765 -660
rect 60775 -690 60805 -660
rect 61045 -610 61075 -580
rect 61085 -610 61115 -580
rect 61125 -610 61155 -580
rect 61045 -650 61075 -620
rect 61085 -650 61115 -620
rect 61125 -650 61155 -620
rect 61045 -690 61075 -660
rect 61085 -690 61115 -660
rect 61125 -690 61155 -660
rect 61395 -610 61425 -580
rect 61435 -610 61465 -580
rect 61475 -610 61505 -580
rect 61395 -650 61425 -620
rect 61435 -650 61465 -620
rect 61475 -650 61505 -620
rect 61395 -690 61425 -660
rect 61435 -690 61465 -660
rect 61475 -690 61505 -660
<< metal2 >>
rect 56205 5065 56245 5070
rect 56205 5035 56210 5065
rect 56240 5060 56245 5065
rect 56675 5065 56715 5070
rect 56675 5060 56680 5065
rect 56240 5040 56680 5060
rect 56240 5035 56245 5040
rect 56205 5030 56245 5035
rect 56675 5035 56680 5040
rect 56710 5035 56715 5065
rect 56675 5030 56715 5035
rect 57085 5065 57125 5070
rect 57085 5035 57090 5065
rect 57120 5060 57125 5065
rect 57555 5065 57595 5070
rect 57555 5060 57560 5065
rect 57120 5040 57560 5060
rect 57120 5035 57125 5040
rect 57085 5030 57125 5035
rect 57555 5035 57560 5040
rect 57590 5035 57595 5065
rect 57555 5030 57595 5035
rect 56880 5010 57245 5015
rect 56880 4980 56885 5010
rect 56915 4980 57030 5010
rect 57060 4980 57150 5010
rect 57180 4980 57210 5010
rect 57240 4980 57245 5010
rect 56880 4970 57245 4980
rect 56880 4940 56885 4970
rect 56915 4940 57030 4970
rect 57060 4940 57150 4970
rect 57180 4940 57210 4970
rect 57240 4940 57245 4970
rect 56085 4930 56125 4935
rect 56085 4900 56090 4930
rect 56120 4925 56125 4930
rect 56205 4930 56245 4935
rect 56205 4925 56210 4930
rect 56120 4905 56210 4925
rect 56120 4900 56125 4905
rect 56085 4895 56125 4900
rect 56205 4900 56210 4905
rect 56240 4925 56245 4930
rect 56265 4930 56305 4935
rect 56265 4925 56270 4930
rect 56240 4905 56270 4925
rect 56240 4900 56245 4905
rect 56205 4895 56245 4900
rect 56265 4900 56270 4905
rect 56300 4900 56305 4930
rect 56265 4895 56305 4900
rect 56880 4930 57245 4940
rect 56880 4900 56885 4930
rect 56915 4900 57030 4930
rect 57060 4900 57150 4930
rect 57180 4900 57210 4930
rect 57240 4900 57245 4930
rect 56880 4895 57245 4900
rect 57495 4930 57535 4935
rect 57495 4900 57500 4930
rect 57530 4925 57535 4930
rect 57555 4930 57595 4935
rect 57555 4925 57560 4930
rect 57530 4905 57560 4925
rect 57530 4900 57535 4905
rect 57495 4895 57535 4900
rect 57555 4900 57560 4905
rect 57590 4925 57595 4930
rect 57675 4930 57715 4935
rect 57675 4925 57680 4930
rect 57590 4905 57680 4925
rect 57590 4900 57595 4905
rect 57555 4895 57595 4900
rect 57675 4900 57680 4905
rect 57710 4900 57715 4930
rect 57675 4895 57715 4900
rect 56555 4840 56920 4845
rect 56555 4810 56560 4840
rect 56590 4810 56620 4840
rect 56650 4810 56740 4840
rect 56770 4810 56885 4840
rect 56915 4810 56920 4840
rect 56555 4800 56920 4810
rect 56555 4770 56560 4800
rect 56590 4770 56620 4800
rect 56650 4770 56740 4800
rect 56770 4770 56885 4800
rect 56915 4770 56920 4800
rect 56555 4760 56920 4770
rect 56555 4730 56560 4760
rect 56590 4730 56620 4760
rect 56650 4730 56740 4760
rect 56770 4730 56885 4760
rect 56915 4730 56920 4760
rect 56555 4725 56920 4730
rect 56205 4525 56245 4530
rect 56205 4495 56210 4525
rect 56240 4520 56245 4525
rect 56675 4525 56715 4530
rect 56675 4520 56680 4525
rect 56240 4500 56680 4520
rect 56240 4495 56245 4500
rect 56205 4490 56245 4495
rect 56675 4495 56680 4500
rect 56710 4495 56715 4525
rect 56675 4490 56715 4495
rect 57085 4525 57125 4530
rect 57085 4495 57090 4525
rect 57120 4520 57125 4525
rect 57555 4525 57595 4530
rect 57555 4520 57560 4525
rect 57120 4500 57560 4520
rect 57120 4495 57125 4500
rect 57085 4490 57125 4495
rect 57555 4495 57560 4500
rect 57590 4495 57595 4525
rect 57555 4490 57595 4495
rect 56150 4480 56190 4485
rect 56150 4450 56155 4480
rect 56185 4475 56190 4480
rect 56630 4480 56660 4485
rect 56185 4455 56630 4475
rect 56185 4450 56190 4455
rect 56150 4445 56190 4450
rect 56825 4480 56865 4485
rect 56825 4475 56830 4480
rect 56660 4455 56830 4475
rect 56630 4445 56660 4450
rect 56825 4450 56830 4455
rect 56860 4475 56865 4480
rect 56860 4470 57606 4475
rect 56860 4455 57576 4470
rect 56860 4450 56865 4455
rect 56825 4445 56865 4450
rect 57576 4435 57606 4440
rect 56935 4425 56975 4430
rect 56935 4395 56940 4425
rect 56970 4410 56975 4425
rect 57135 4415 57175 4420
rect 57135 4410 57140 4415
rect 56970 4395 57140 4410
rect 56935 4390 57140 4395
rect 57135 4385 57140 4390
rect 57170 4410 57175 4415
rect 57615 4415 57655 4420
rect 57615 4410 57620 4415
rect 57170 4390 57620 4410
rect 57170 4385 57175 4390
rect 57135 4380 57175 4385
rect 57615 4385 57620 4390
rect 57650 4385 57655 4415
rect 57615 4380 57655 4385
rect 52290 4320 61510 4325
rect 52290 4290 52295 4320
rect 52325 4290 52335 4320
rect 52365 4290 52375 4320
rect 52405 4290 52645 4320
rect 52675 4290 52685 4320
rect 52715 4290 52725 4320
rect 52755 4290 52995 4320
rect 53025 4290 53035 4320
rect 53065 4290 53075 4320
rect 53105 4290 53345 4320
rect 53375 4290 53385 4320
rect 53415 4290 53425 4320
rect 53455 4290 54045 4320
rect 54075 4290 54085 4320
rect 54115 4290 54125 4320
rect 54155 4290 54595 4320
rect 54625 4290 54955 4320
rect 54985 4290 55315 4320
rect 55345 4290 55540 4320
rect 55570 4290 55580 4320
rect 55610 4290 55620 4320
rect 55650 4290 56885 4320
rect 56915 4290 58150 4320
rect 58180 4290 58190 4320
rect 58220 4290 58230 4320
rect 58260 4290 58455 4320
rect 58485 4290 58815 4320
rect 58845 4290 59175 4320
rect 59205 4290 59645 4320
rect 59675 4290 59685 4320
rect 59715 4290 59725 4320
rect 59755 4290 60345 4320
rect 60375 4290 60385 4320
rect 60415 4290 60425 4320
rect 60455 4290 60695 4320
rect 60725 4290 60735 4320
rect 60765 4290 60775 4320
rect 60805 4290 61045 4320
rect 61075 4290 61085 4320
rect 61115 4290 61125 4320
rect 61155 4290 61395 4320
rect 61425 4290 61435 4320
rect 61465 4290 61475 4320
rect 61505 4290 61510 4320
rect 52290 4280 61510 4290
rect 52290 4250 52295 4280
rect 52325 4250 52335 4280
rect 52365 4250 52375 4280
rect 52405 4250 52645 4280
rect 52675 4250 52685 4280
rect 52715 4250 52725 4280
rect 52755 4250 52995 4280
rect 53025 4250 53035 4280
rect 53065 4250 53075 4280
rect 53105 4250 53345 4280
rect 53375 4250 53385 4280
rect 53415 4250 53425 4280
rect 53455 4250 54045 4280
rect 54075 4250 54085 4280
rect 54115 4250 54125 4280
rect 54155 4250 54595 4280
rect 54625 4250 54955 4280
rect 54985 4250 55315 4280
rect 55345 4250 55540 4280
rect 55570 4250 55580 4280
rect 55610 4250 55620 4280
rect 55650 4250 56885 4280
rect 56915 4250 58150 4280
rect 58180 4250 58190 4280
rect 58220 4250 58230 4280
rect 58260 4250 58455 4280
rect 58485 4250 58815 4280
rect 58845 4250 59175 4280
rect 59205 4250 59645 4280
rect 59675 4250 59685 4280
rect 59715 4250 59725 4280
rect 59755 4250 60345 4280
rect 60375 4250 60385 4280
rect 60415 4250 60425 4280
rect 60455 4250 60695 4280
rect 60725 4250 60735 4280
rect 60765 4250 60775 4280
rect 60805 4250 61045 4280
rect 61075 4250 61085 4280
rect 61115 4250 61125 4280
rect 61155 4250 61395 4280
rect 61425 4250 61435 4280
rect 61465 4250 61475 4280
rect 61505 4250 61510 4280
rect 52290 4240 61510 4250
rect 52290 4210 52295 4240
rect 52325 4210 52335 4240
rect 52365 4210 52375 4240
rect 52405 4210 52645 4240
rect 52675 4210 52685 4240
rect 52715 4210 52725 4240
rect 52755 4210 52995 4240
rect 53025 4210 53035 4240
rect 53065 4210 53075 4240
rect 53105 4210 53345 4240
rect 53375 4210 53385 4240
rect 53415 4210 53425 4240
rect 53455 4210 54045 4240
rect 54075 4210 54085 4240
rect 54115 4210 54125 4240
rect 54155 4210 54595 4240
rect 54625 4210 54955 4240
rect 54985 4210 55315 4240
rect 55345 4210 55540 4240
rect 55570 4210 55580 4240
rect 55610 4210 55620 4240
rect 55650 4210 56885 4240
rect 56915 4210 58150 4240
rect 58180 4210 58190 4240
rect 58220 4210 58230 4240
rect 58260 4210 58455 4240
rect 58485 4210 58815 4240
rect 58845 4210 59175 4240
rect 59205 4210 59645 4240
rect 59675 4210 59685 4240
rect 59715 4210 59725 4240
rect 59755 4210 60345 4240
rect 60375 4210 60385 4240
rect 60415 4210 60425 4240
rect 60455 4210 60695 4240
rect 60725 4210 60735 4240
rect 60765 4210 60775 4240
rect 60805 4210 61045 4240
rect 61075 4210 61085 4240
rect 61115 4210 61125 4240
rect 61155 4210 61395 4240
rect 61425 4210 61435 4240
rect 61465 4210 61475 4240
rect 61505 4210 61510 4240
rect 52290 4205 61510 4210
rect 54650 4185 56765 4190
rect 54650 4155 54655 4185
rect 54685 4155 54695 4185
rect 54725 4155 54735 4185
rect 54765 4155 54775 4185
rect 54805 4155 54815 4185
rect 54845 4155 54855 4185
rect 54885 4155 54895 4185
rect 54925 4155 55015 4185
rect 55045 4155 55055 4185
rect 55085 4155 55095 4185
rect 55125 4155 55135 4185
rect 55165 4155 55175 4185
rect 55205 4155 55215 4185
rect 55245 4155 55255 4185
rect 55285 4155 56010 4185
rect 56040 4155 56050 4185
rect 56080 4155 56090 4185
rect 56120 4155 56130 4185
rect 56160 4155 56170 4185
rect 56200 4155 56210 4185
rect 56240 4155 56250 4185
rect 56280 4155 56290 4185
rect 56320 4155 56330 4185
rect 56360 4155 56370 4185
rect 56400 4155 56410 4185
rect 56440 4155 56450 4185
rect 56480 4155 56490 4185
rect 56520 4155 56530 4185
rect 56560 4155 56570 4185
rect 56600 4155 56610 4185
rect 56640 4155 56650 4185
rect 56680 4155 56690 4185
rect 56720 4155 56730 4185
rect 56760 4155 56765 4185
rect 54650 4145 56765 4155
rect 54650 4115 54655 4145
rect 54685 4115 54695 4145
rect 54725 4115 54735 4145
rect 54765 4115 54775 4145
rect 54805 4115 54815 4145
rect 54845 4115 54855 4145
rect 54885 4115 54895 4145
rect 54925 4115 55015 4145
rect 55045 4115 55055 4145
rect 55085 4115 55095 4145
rect 55125 4115 55135 4145
rect 55165 4115 55175 4145
rect 55205 4115 55215 4145
rect 55245 4115 55255 4145
rect 55285 4115 56010 4145
rect 56040 4115 56050 4145
rect 56080 4115 56090 4145
rect 56120 4115 56130 4145
rect 56160 4115 56170 4145
rect 56200 4115 56210 4145
rect 56240 4115 56250 4145
rect 56280 4115 56290 4145
rect 56320 4115 56330 4145
rect 56360 4115 56370 4145
rect 56400 4115 56410 4145
rect 56440 4115 56450 4145
rect 56480 4115 56490 4145
rect 56520 4115 56530 4145
rect 56560 4115 56570 4145
rect 56600 4115 56610 4145
rect 56640 4115 56650 4145
rect 56680 4115 56690 4145
rect 56720 4115 56730 4145
rect 56760 4115 56765 4145
rect 54650 4105 56765 4115
rect 54650 4075 54655 4105
rect 54685 4075 54695 4105
rect 54725 4075 54735 4105
rect 54765 4075 54775 4105
rect 54805 4075 54815 4105
rect 54845 4075 54855 4105
rect 54885 4075 54895 4105
rect 54925 4075 55015 4105
rect 55045 4075 55055 4105
rect 55085 4075 55095 4105
rect 55125 4075 55135 4105
rect 55165 4075 55175 4105
rect 55205 4075 55215 4105
rect 55245 4075 55255 4105
rect 55285 4075 56010 4105
rect 56040 4075 56050 4105
rect 56080 4075 56090 4105
rect 56120 4075 56130 4105
rect 56160 4075 56170 4105
rect 56200 4075 56210 4105
rect 56240 4075 56250 4105
rect 56280 4075 56290 4105
rect 56320 4075 56330 4105
rect 56360 4075 56370 4105
rect 56400 4075 56410 4105
rect 56440 4075 56450 4105
rect 56480 4075 56490 4105
rect 56520 4075 56530 4105
rect 56560 4075 56570 4105
rect 56600 4075 56610 4105
rect 56640 4075 56650 4105
rect 56680 4075 56690 4105
rect 56720 4075 56730 4105
rect 56760 4075 56765 4105
rect 54650 4070 56765 4075
rect 57035 4185 59150 4190
rect 57035 4155 57040 4185
rect 57070 4155 57080 4185
rect 57110 4155 57120 4185
rect 57150 4155 57160 4185
rect 57190 4155 57200 4185
rect 57230 4155 57240 4185
rect 57270 4155 57280 4185
rect 57310 4155 57320 4185
rect 57350 4155 57360 4185
rect 57390 4155 57400 4185
rect 57430 4155 57440 4185
rect 57470 4155 57480 4185
rect 57510 4155 57520 4185
rect 57550 4155 57560 4185
rect 57590 4155 57600 4185
rect 57630 4155 57640 4185
rect 57670 4155 57680 4185
rect 57710 4155 57720 4185
rect 57750 4155 57760 4185
rect 57790 4155 58515 4185
rect 58545 4155 58555 4185
rect 58585 4155 58595 4185
rect 58625 4155 58635 4185
rect 58665 4155 58675 4185
rect 58705 4155 58715 4185
rect 58745 4155 58755 4185
rect 58785 4155 58875 4185
rect 58905 4155 58915 4185
rect 58945 4155 58955 4185
rect 58985 4155 58995 4185
rect 59025 4155 59035 4185
rect 59065 4155 59075 4185
rect 59105 4155 59115 4185
rect 59145 4155 59150 4185
rect 57035 4145 59150 4155
rect 57035 4115 57040 4145
rect 57070 4115 57080 4145
rect 57110 4115 57120 4145
rect 57150 4115 57160 4145
rect 57190 4115 57200 4145
rect 57230 4115 57240 4145
rect 57270 4115 57280 4145
rect 57310 4115 57320 4145
rect 57350 4115 57360 4145
rect 57390 4115 57400 4145
rect 57430 4115 57440 4145
rect 57470 4115 57480 4145
rect 57510 4115 57520 4145
rect 57550 4115 57560 4145
rect 57590 4115 57600 4145
rect 57630 4115 57640 4145
rect 57670 4115 57680 4145
rect 57710 4115 57720 4145
rect 57750 4115 57760 4145
rect 57790 4115 58515 4145
rect 58545 4115 58555 4145
rect 58585 4115 58595 4145
rect 58625 4115 58635 4145
rect 58665 4115 58675 4145
rect 58705 4115 58715 4145
rect 58745 4115 58755 4145
rect 58785 4115 58875 4145
rect 58905 4115 58915 4145
rect 58945 4115 58955 4145
rect 58985 4115 58995 4145
rect 59025 4115 59035 4145
rect 59065 4115 59075 4145
rect 59105 4115 59115 4145
rect 59145 4115 59150 4145
rect 57035 4105 59150 4115
rect 57035 4075 57040 4105
rect 57070 4075 57080 4105
rect 57110 4075 57120 4105
rect 57150 4075 57160 4105
rect 57190 4075 57200 4105
rect 57230 4075 57240 4105
rect 57270 4075 57280 4105
rect 57310 4075 57320 4105
rect 57350 4075 57360 4105
rect 57390 4075 57400 4105
rect 57430 4075 57440 4105
rect 57470 4075 57480 4105
rect 57510 4075 57520 4105
rect 57550 4075 57560 4105
rect 57590 4075 57600 4105
rect 57630 4075 57640 4105
rect 57670 4075 57680 4105
rect 57710 4075 57720 4105
rect 57750 4075 57760 4105
rect 57790 4075 58515 4105
rect 58545 4075 58555 4105
rect 58585 4075 58595 4105
rect 58625 4075 58635 4105
rect 58665 4075 58675 4105
rect 58705 4075 58715 4105
rect 58745 4075 58755 4105
rect 58785 4075 58875 4105
rect 58905 4075 58915 4105
rect 58945 4075 58955 4105
rect 58985 4075 58995 4105
rect 59025 4075 59035 4105
rect 59065 4075 59075 4105
rect 59105 4075 59115 4105
rect 59145 4075 59150 4105
rect 57035 4070 59150 4075
rect 54590 4050 54630 4055
rect 54590 4020 54595 4050
rect 54625 4045 54630 4050
rect 54710 4050 54750 4055
rect 54710 4045 54715 4050
rect 54625 4025 54715 4045
rect 54625 4020 54630 4025
rect 54590 4015 54630 4020
rect 54710 4020 54715 4025
rect 54745 4045 54750 4050
rect 54830 4050 54870 4055
rect 54830 4045 54835 4050
rect 54745 4025 54835 4045
rect 54745 4020 54750 4025
rect 54710 4015 54750 4020
rect 54830 4020 54835 4025
rect 54865 4045 54870 4050
rect 54950 4050 54990 4055
rect 54950 4045 54955 4050
rect 54865 4025 54955 4045
rect 54865 4020 54870 4025
rect 54830 4015 54870 4020
rect 54950 4020 54955 4025
rect 54985 4045 54990 4050
rect 55070 4050 55110 4055
rect 55070 4045 55075 4050
rect 54985 4025 55075 4045
rect 54985 4020 54990 4025
rect 54950 4015 54990 4020
rect 55070 4020 55075 4025
rect 55105 4045 55110 4050
rect 55190 4050 55230 4055
rect 55190 4045 55195 4050
rect 55105 4025 55195 4045
rect 55105 4020 55110 4025
rect 55070 4015 55110 4020
rect 55190 4020 55195 4025
rect 55225 4045 55230 4050
rect 55310 4050 55350 4055
rect 55310 4045 55315 4050
rect 55225 4025 55315 4045
rect 55225 4020 55230 4025
rect 55190 4015 55230 4020
rect 55310 4020 55315 4025
rect 55345 4020 55350 4050
rect 55310 4015 55350 4020
rect 56065 4050 56105 4055
rect 56065 4020 56070 4050
rect 56100 4045 56105 4050
rect 56185 4050 56225 4055
rect 56185 4045 56190 4050
rect 56100 4025 56190 4045
rect 56100 4020 56105 4025
rect 56065 4015 56105 4020
rect 56185 4020 56190 4025
rect 56220 4045 56225 4050
rect 56305 4050 56345 4055
rect 56305 4045 56310 4050
rect 56220 4025 56310 4045
rect 56220 4020 56225 4025
rect 56185 4015 56225 4020
rect 56305 4020 56310 4025
rect 56340 4045 56345 4050
rect 56425 4050 56465 4055
rect 56425 4045 56430 4050
rect 56340 4025 56430 4045
rect 56340 4020 56345 4025
rect 56305 4015 56345 4020
rect 56425 4020 56430 4025
rect 56460 4045 56465 4050
rect 56545 4050 56585 4055
rect 56545 4045 56550 4050
rect 56460 4025 56550 4045
rect 56460 4020 56465 4025
rect 56425 4015 56465 4020
rect 56545 4020 56550 4025
rect 56580 4045 56585 4050
rect 56665 4050 56705 4055
rect 56665 4045 56670 4050
rect 56580 4025 56670 4045
rect 56580 4020 56585 4025
rect 56545 4015 56585 4020
rect 56665 4020 56670 4025
rect 56700 4020 56705 4050
rect 56665 4015 56705 4020
rect 57095 4050 57135 4055
rect 57095 4020 57100 4050
rect 57130 4045 57135 4050
rect 57215 4050 57255 4055
rect 57215 4045 57220 4050
rect 57130 4025 57220 4045
rect 57130 4020 57135 4025
rect 57095 4015 57135 4020
rect 57215 4020 57220 4025
rect 57250 4045 57255 4050
rect 57335 4050 57375 4055
rect 57335 4045 57340 4050
rect 57250 4025 57340 4045
rect 57250 4020 57255 4025
rect 57215 4015 57255 4020
rect 57335 4020 57340 4025
rect 57370 4045 57375 4050
rect 57455 4050 57495 4055
rect 57455 4045 57460 4050
rect 57370 4025 57460 4045
rect 57370 4020 57375 4025
rect 57335 4015 57375 4020
rect 57455 4020 57460 4025
rect 57490 4045 57495 4050
rect 57575 4050 57615 4055
rect 57575 4045 57580 4050
rect 57490 4025 57580 4045
rect 57490 4020 57495 4025
rect 57455 4015 57495 4020
rect 57575 4020 57580 4025
rect 57610 4045 57615 4050
rect 57695 4050 57735 4055
rect 57695 4045 57700 4050
rect 57610 4025 57700 4045
rect 57610 4020 57615 4025
rect 57575 4015 57615 4020
rect 57695 4020 57700 4025
rect 57730 4020 57735 4050
rect 57695 4015 57735 4020
rect 58450 4050 58490 4055
rect 58450 4020 58455 4050
rect 58485 4045 58490 4050
rect 58570 4050 58610 4055
rect 58570 4045 58575 4050
rect 58485 4025 58575 4045
rect 58485 4020 58490 4025
rect 58450 4015 58490 4020
rect 58570 4020 58575 4025
rect 58605 4045 58610 4050
rect 58690 4050 58730 4055
rect 58690 4045 58695 4050
rect 58605 4025 58695 4045
rect 58605 4020 58610 4025
rect 58570 4015 58610 4020
rect 58690 4020 58695 4025
rect 58725 4045 58730 4050
rect 58810 4050 58850 4055
rect 58810 4045 58815 4050
rect 58725 4025 58815 4045
rect 58725 4020 58730 4025
rect 58690 4015 58730 4020
rect 58810 4020 58815 4025
rect 58845 4045 58850 4050
rect 58930 4050 58970 4055
rect 58930 4045 58935 4050
rect 58845 4025 58935 4045
rect 58845 4020 58850 4025
rect 58810 4015 58850 4020
rect 58930 4020 58935 4025
rect 58965 4045 58970 4050
rect 59050 4050 59090 4055
rect 59050 4045 59055 4050
rect 58965 4025 59055 4045
rect 58965 4020 58970 4025
rect 58930 4015 58970 4020
rect 59050 4020 59055 4025
rect 59085 4045 59090 4050
rect 59170 4050 59210 4055
rect 59170 4045 59175 4050
rect 59085 4025 59175 4045
rect 59085 4020 59090 4025
rect 59050 4015 59090 4020
rect 59170 4020 59175 4025
rect 59205 4020 59210 4050
rect 59170 4015 59210 4020
rect 54650 3660 54690 3665
rect 54650 3630 54655 3660
rect 54685 3655 54690 3660
rect 54770 3660 54810 3665
rect 54770 3655 54775 3660
rect 54685 3635 54775 3655
rect 54685 3630 54690 3635
rect 54650 3625 54690 3630
rect 54770 3630 54775 3635
rect 54805 3655 54810 3660
rect 54890 3660 54930 3665
rect 54890 3655 54895 3660
rect 54805 3635 54895 3655
rect 54805 3630 54810 3635
rect 54770 3625 54810 3630
rect 54890 3630 54895 3635
rect 54925 3655 54930 3660
rect 55010 3660 55050 3665
rect 55010 3655 55015 3660
rect 54925 3635 55015 3655
rect 54925 3630 54930 3635
rect 54890 3625 54930 3630
rect 55010 3630 55015 3635
rect 55045 3655 55050 3660
rect 55130 3660 55170 3665
rect 55130 3655 55135 3660
rect 55045 3635 55135 3655
rect 55045 3630 55050 3635
rect 55010 3625 55050 3630
rect 55130 3630 55135 3635
rect 55165 3655 55170 3660
rect 55250 3660 55290 3665
rect 55250 3655 55255 3660
rect 55165 3635 55255 3655
rect 55165 3630 55170 3635
rect 55130 3625 55170 3630
rect 55250 3630 55255 3635
rect 55285 3630 55290 3660
rect 55250 3625 55290 3630
rect 56065 3660 56105 3665
rect 56065 3630 56070 3660
rect 56100 3655 56105 3660
rect 56185 3660 56225 3665
rect 56185 3655 56190 3660
rect 56100 3635 56190 3655
rect 56100 3630 56105 3635
rect 56065 3625 56105 3630
rect 56185 3630 56190 3635
rect 56220 3655 56225 3660
rect 56305 3660 56345 3665
rect 56305 3655 56310 3660
rect 56220 3635 56310 3655
rect 56220 3630 56225 3635
rect 56185 3625 56225 3630
rect 56305 3630 56310 3635
rect 56340 3655 56345 3660
rect 56425 3660 56465 3665
rect 56425 3655 56430 3660
rect 56340 3635 56430 3655
rect 56340 3630 56345 3635
rect 56305 3625 56345 3630
rect 56425 3630 56430 3635
rect 56460 3655 56465 3660
rect 56545 3660 56585 3665
rect 56545 3655 56550 3660
rect 56460 3635 56550 3655
rect 56460 3630 56465 3635
rect 56425 3625 56465 3630
rect 56545 3630 56550 3635
rect 56580 3655 56585 3660
rect 56665 3660 56705 3665
rect 56665 3655 56670 3660
rect 56580 3635 56670 3655
rect 56580 3630 56585 3635
rect 56545 3625 56585 3630
rect 56665 3630 56670 3635
rect 56700 3630 56705 3660
rect 56665 3625 56705 3630
rect 57095 3660 57135 3665
rect 57095 3630 57100 3660
rect 57130 3655 57135 3660
rect 57215 3660 57255 3665
rect 57215 3655 57220 3660
rect 57130 3635 57220 3655
rect 57130 3630 57135 3635
rect 57095 3625 57135 3630
rect 57215 3630 57220 3635
rect 57250 3655 57255 3660
rect 57335 3660 57375 3665
rect 57335 3655 57340 3660
rect 57250 3635 57340 3655
rect 57250 3630 57255 3635
rect 57215 3625 57255 3630
rect 57335 3630 57340 3635
rect 57370 3655 57375 3660
rect 57455 3660 57495 3665
rect 57455 3655 57460 3660
rect 57370 3635 57460 3655
rect 57370 3630 57375 3635
rect 57335 3625 57375 3630
rect 57455 3630 57460 3635
rect 57490 3655 57495 3660
rect 57575 3660 57615 3665
rect 57575 3655 57580 3660
rect 57490 3635 57580 3655
rect 57490 3630 57495 3635
rect 57455 3625 57495 3630
rect 57575 3630 57580 3635
rect 57610 3655 57615 3660
rect 57695 3660 57735 3665
rect 57695 3655 57700 3660
rect 57610 3635 57700 3655
rect 57610 3630 57615 3635
rect 57575 3625 57615 3630
rect 57695 3630 57700 3635
rect 57730 3630 57735 3660
rect 57695 3625 57735 3630
rect 58510 3660 58550 3665
rect 58510 3630 58515 3660
rect 58545 3655 58550 3660
rect 58630 3660 58670 3665
rect 58630 3655 58635 3660
rect 58545 3635 58635 3655
rect 58545 3630 58550 3635
rect 58510 3625 58550 3630
rect 58630 3630 58635 3635
rect 58665 3655 58670 3660
rect 58750 3660 58790 3665
rect 58750 3655 58755 3660
rect 58665 3635 58755 3655
rect 58665 3630 58670 3635
rect 58630 3625 58670 3630
rect 58750 3630 58755 3635
rect 58785 3655 58790 3660
rect 58870 3660 58910 3665
rect 58870 3655 58875 3660
rect 58785 3635 58875 3655
rect 58785 3630 58790 3635
rect 58750 3625 58790 3630
rect 58870 3630 58875 3635
rect 58905 3655 58910 3660
rect 58990 3660 59030 3665
rect 58990 3655 58995 3660
rect 58905 3635 58995 3655
rect 58905 3630 58910 3635
rect 58870 3625 58910 3630
rect 58990 3630 58995 3635
rect 59025 3655 59030 3660
rect 59110 3660 59150 3665
rect 59110 3655 59115 3660
rect 59025 3635 59115 3655
rect 59025 3630 59030 3635
rect 58990 3625 59030 3630
rect 59110 3630 59115 3635
rect 59145 3630 59150 3660
rect 59110 3625 59150 3630
rect 56365 3580 56405 3585
rect 56365 3550 56370 3580
rect 56400 3575 56405 3580
rect 56835 3580 56875 3585
rect 56835 3575 56840 3580
rect 56400 3555 56840 3575
rect 56400 3550 56405 3555
rect 56365 3545 56405 3550
rect 56835 3550 56840 3555
rect 56870 3575 56875 3580
rect 57395 3580 57435 3585
rect 57395 3575 57400 3580
rect 56870 3555 57400 3575
rect 56870 3550 56875 3555
rect 56835 3545 56875 3550
rect 57395 3550 57400 3555
rect 57430 3550 57435 3580
rect 57395 3545 57435 3550
rect 54950 3535 54990 3540
rect 54950 3505 54955 3535
rect 54985 3530 54990 3535
rect 56925 3535 56965 3540
rect 56925 3530 56930 3535
rect 54985 3510 56930 3530
rect 54985 3505 54990 3510
rect 54950 3500 54990 3505
rect 56925 3505 56930 3510
rect 56960 3530 56965 3535
rect 58810 3535 58850 3540
rect 58810 3530 58815 3535
rect 56960 3510 58815 3530
rect 56960 3505 56965 3510
rect 56925 3500 56965 3505
rect 58810 3505 58815 3510
rect 58845 3505 58850 3535
rect 58810 3500 58850 3505
rect 55400 3490 56705 3495
rect 55400 3460 55405 3490
rect 55435 3460 55445 3490
rect 55475 3460 55485 3490
rect 55515 3460 56070 3490
rect 56100 3460 56110 3490
rect 56140 3460 56150 3490
rect 56180 3460 56190 3490
rect 56220 3460 56230 3490
rect 56260 3460 56270 3490
rect 56300 3460 56310 3490
rect 56340 3460 56350 3490
rect 56380 3460 56390 3490
rect 56420 3460 56430 3490
rect 56460 3460 56470 3490
rect 56500 3460 56510 3490
rect 56540 3460 56550 3490
rect 56580 3460 56590 3490
rect 56620 3460 56630 3490
rect 56660 3460 56670 3490
rect 56700 3460 56705 3490
rect 55400 3450 56705 3460
rect 55400 3420 55405 3450
rect 55435 3420 55445 3450
rect 55475 3420 55485 3450
rect 55515 3420 56070 3450
rect 56100 3420 56110 3450
rect 56140 3420 56150 3450
rect 56180 3420 56190 3450
rect 56220 3420 56230 3450
rect 56260 3420 56270 3450
rect 56300 3420 56310 3450
rect 56340 3420 56350 3450
rect 56380 3420 56390 3450
rect 56420 3420 56430 3450
rect 56460 3420 56470 3450
rect 56500 3420 56510 3450
rect 56540 3420 56550 3450
rect 56580 3420 56590 3450
rect 56620 3420 56630 3450
rect 56660 3420 56670 3450
rect 56700 3420 56705 3450
rect 55400 3410 56705 3420
rect 55400 3380 55405 3410
rect 55435 3380 55445 3410
rect 55475 3380 55485 3410
rect 55515 3380 56070 3410
rect 56100 3380 56110 3410
rect 56140 3380 56150 3410
rect 56180 3380 56190 3410
rect 56220 3380 56230 3410
rect 56260 3380 56270 3410
rect 56300 3380 56310 3410
rect 56340 3380 56350 3410
rect 56380 3380 56390 3410
rect 56420 3380 56430 3410
rect 56460 3380 56470 3410
rect 56500 3380 56510 3410
rect 56540 3380 56550 3410
rect 56580 3380 56590 3410
rect 56620 3380 56630 3410
rect 56660 3380 56670 3410
rect 56700 3380 56705 3410
rect 54255 3375 54295 3380
rect 55400 3375 56705 3380
rect 57095 3490 58400 3495
rect 57095 3460 57100 3490
rect 57130 3460 57140 3490
rect 57170 3460 57180 3490
rect 57210 3460 57220 3490
rect 57250 3460 57260 3490
rect 57290 3460 57300 3490
rect 57330 3460 57340 3490
rect 57370 3460 57380 3490
rect 57410 3460 57420 3490
rect 57450 3460 57460 3490
rect 57490 3460 57500 3490
rect 57530 3460 57540 3490
rect 57570 3460 57580 3490
rect 57610 3460 57620 3490
rect 57650 3460 57660 3490
rect 57690 3460 57700 3490
rect 57730 3460 58285 3490
rect 58315 3460 58325 3490
rect 58355 3460 58365 3490
rect 58395 3460 58400 3490
rect 57095 3450 58400 3460
rect 57095 3420 57100 3450
rect 57130 3420 57140 3450
rect 57170 3420 57180 3450
rect 57210 3420 57220 3450
rect 57250 3420 57260 3450
rect 57290 3420 57300 3450
rect 57330 3420 57340 3450
rect 57370 3420 57380 3450
rect 57410 3420 57420 3450
rect 57450 3420 57460 3450
rect 57490 3420 57500 3450
rect 57530 3420 57540 3450
rect 57570 3420 57580 3450
rect 57610 3420 57620 3450
rect 57650 3420 57660 3450
rect 57690 3420 57700 3450
rect 57730 3420 58285 3450
rect 58315 3420 58325 3450
rect 58355 3420 58365 3450
rect 58395 3420 58400 3450
rect 57095 3410 58400 3420
rect 57095 3380 57100 3410
rect 57130 3380 57140 3410
rect 57170 3380 57180 3410
rect 57210 3380 57220 3410
rect 57250 3380 57260 3410
rect 57290 3380 57300 3410
rect 57330 3380 57340 3410
rect 57370 3380 57380 3410
rect 57410 3380 57420 3410
rect 57450 3380 57460 3410
rect 57490 3380 57500 3410
rect 57530 3380 57540 3410
rect 57570 3380 57580 3410
rect 57610 3380 57620 3410
rect 57650 3380 57660 3410
rect 57690 3380 57700 3410
rect 57730 3380 58285 3410
rect 58315 3380 58325 3410
rect 58355 3380 58365 3410
rect 58395 3380 58400 3410
rect 57095 3375 58400 3380
rect 59505 3375 59545 3380
rect 54255 3345 54260 3375
rect 54290 3345 54295 3375
rect 54255 3340 54295 3345
rect 54620 3355 59180 3360
rect 54620 3325 54625 3355
rect 54655 3325 54735 3355
rect 54765 3325 54845 3355
rect 54875 3325 54955 3355
rect 54985 3325 55065 3355
rect 55095 3325 55175 3355
rect 55205 3325 55285 3355
rect 55315 3325 55540 3355
rect 55570 3325 55580 3355
rect 55610 3325 55620 3355
rect 55650 3325 56515 3355
rect 56545 3325 56680 3355
rect 56710 3325 56845 3355
rect 56875 3325 56925 3355
rect 56955 3325 57090 3355
rect 57120 3325 57255 3355
rect 57285 3325 58150 3355
rect 58180 3325 58190 3355
rect 58220 3325 58230 3355
rect 58260 3325 58485 3355
rect 58515 3325 58595 3355
rect 58625 3325 58705 3355
rect 58735 3325 58815 3355
rect 58845 3325 58925 3355
rect 58955 3325 59035 3355
rect 59065 3325 59145 3355
rect 59175 3325 59180 3355
rect 59505 3345 59510 3375
rect 59540 3345 59545 3375
rect 59505 3340 59545 3345
rect 54620 3315 59180 3325
rect 54620 3285 54625 3315
rect 54655 3285 54735 3315
rect 54765 3285 54845 3315
rect 54875 3285 54955 3315
rect 54985 3285 55065 3315
rect 55095 3285 55175 3315
rect 55205 3285 55285 3315
rect 55315 3285 55540 3315
rect 55570 3285 55580 3315
rect 55610 3285 55620 3315
rect 55650 3285 56515 3315
rect 56545 3285 56680 3315
rect 56710 3285 56845 3315
rect 56875 3285 56925 3315
rect 56955 3285 57090 3315
rect 57120 3285 57255 3315
rect 57285 3285 58150 3315
rect 58180 3285 58190 3315
rect 58220 3285 58230 3315
rect 58260 3285 58485 3315
rect 58515 3285 58595 3315
rect 58625 3285 58705 3315
rect 58735 3285 58815 3315
rect 58845 3285 58925 3315
rect 58955 3285 59035 3315
rect 59065 3285 59145 3315
rect 59175 3285 59180 3315
rect 54620 3275 59180 3285
rect 54620 3245 54625 3275
rect 54655 3245 54735 3275
rect 54765 3245 54845 3275
rect 54875 3245 54955 3275
rect 54985 3245 55065 3275
rect 55095 3245 55175 3275
rect 55205 3245 55285 3275
rect 55315 3245 55540 3275
rect 55570 3245 55580 3275
rect 55610 3245 55620 3275
rect 55650 3245 56515 3275
rect 56545 3245 56680 3275
rect 56710 3245 56845 3275
rect 56875 3245 56925 3275
rect 56955 3245 57090 3275
rect 57120 3245 57255 3275
rect 57285 3245 58150 3275
rect 58180 3245 58190 3275
rect 58220 3245 58230 3275
rect 58260 3245 58485 3275
rect 58515 3245 58595 3275
rect 58625 3245 58705 3275
rect 58735 3245 58815 3275
rect 58845 3245 58925 3275
rect 58955 3245 59035 3275
rect 59065 3245 59145 3275
rect 59175 3245 59180 3275
rect 54620 3240 59180 3245
rect 56620 3220 56660 3225
rect 54675 3190 54715 3195
rect 54675 3160 54680 3190
rect 54710 3185 54715 3190
rect 54785 3190 54825 3195
rect 54785 3185 54790 3190
rect 54710 3165 54790 3185
rect 54710 3160 54715 3165
rect 54675 3155 54715 3160
rect 54785 3160 54790 3165
rect 54820 3185 54825 3190
rect 54895 3190 54935 3195
rect 54895 3185 54900 3190
rect 54820 3165 54900 3185
rect 54820 3160 54825 3165
rect 54785 3155 54825 3160
rect 54895 3160 54900 3165
rect 54930 3185 54935 3190
rect 55005 3190 55045 3195
rect 55005 3185 55010 3190
rect 54930 3165 55010 3185
rect 54930 3160 54935 3165
rect 54895 3155 54935 3160
rect 55005 3160 55010 3165
rect 55040 3185 55045 3190
rect 55115 3190 55155 3195
rect 55115 3185 55120 3190
rect 55040 3165 55120 3185
rect 55040 3160 55045 3165
rect 55005 3155 55045 3160
rect 55115 3160 55120 3165
rect 55150 3185 55155 3190
rect 55225 3190 55265 3195
rect 55225 3185 55230 3190
rect 55150 3165 55230 3185
rect 55150 3160 55155 3165
rect 55115 3155 55155 3160
rect 55225 3160 55230 3165
rect 55260 3160 55265 3190
rect 56620 3190 56625 3220
rect 56655 3215 56660 3220
rect 56730 3220 56770 3225
rect 56730 3215 56735 3220
rect 56655 3195 56735 3215
rect 56655 3190 56660 3195
rect 56620 3185 56660 3190
rect 56730 3190 56735 3195
rect 56765 3190 56770 3220
rect 56730 3185 56770 3190
rect 57030 3220 57070 3225
rect 57030 3190 57035 3220
rect 57065 3215 57070 3220
rect 57140 3220 57180 3225
rect 57140 3215 57145 3220
rect 57065 3195 57145 3215
rect 57065 3190 57070 3195
rect 57030 3185 57070 3190
rect 57140 3190 57145 3195
rect 57175 3190 57180 3220
rect 57140 3185 57180 3190
rect 58535 3190 58575 3195
rect 55225 3155 55265 3160
rect 58535 3160 58540 3190
rect 58570 3185 58575 3190
rect 58645 3190 58685 3195
rect 58645 3185 58650 3190
rect 58570 3165 58650 3185
rect 58570 3160 58575 3165
rect 58535 3155 58575 3160
rect 58645 3160 58650 3165
rect 58680 3185 58685 3190
rect 58755 3190 58795 3195
rect 58755 3185 58760 3190
rect 58680 3165 58760 3185
rect 58680 3160 58685 3165
rect 58645 3155 58685 3160
rect 58755 3160 58760 3165
rect 58790 3185 58795 3190
rect 58865 3190 58905 3195
rect 58865 3185 58870 3190
rect 58790 3165 58870 3185
rect 58790 3160 58795 3165
rect 58755 3155 58795 3160
rect 58865 3160 58870 3165
rect 58900 3185 58905 3190
rect 58975 3190 59015 3195
rect 58975 3185 58980 3190
rect 58900 3165 58980 3185
rect 58900 3160 58905 3165
rect 58865 3155 58905 3160
rect 58975 3160 58980 3165
rect 59010 3185 59015 3190
rect 59085 3190 59125 3195
rect 59085 3185 59090 3190
rect 59010 3165 59090 3185
rect 59010 3160 59015 3165
rect 58975 3155 59015 3160
rect 59085 3160 59090 3165
rect 59120 3160 59125 3190
rect 59085 3155 59125 3160
rect 56560 2910 56590 2915
rect 56800 2910 56830 2915
rect 56675 2900 56715 2905
rect 56675 2895 56680 2900
rect 56590 2880 56680 2895
rect 56560 2875 56680 2880
rect 56675 2870 56680 2875
rect 56710 2895 56715 2900
rect 56710 2880 56800 2895
rect 57085 2900 57125 2905
rect 57085 2895 57090 2900
rect 56830 2880 57090 2895
rect 56710 2875 57090 2880
rect 56710 2870 56715 2875
rect 56675 2865 56715 2870
rect 57085 2870 57090 2875
rect 57120 2895 57125 2900
rect 57120 2875 57130 2895
rect 57120 2870 57125 2875
rect 57085 2865 57125 2870
rect 56600 2830 56640 2835
rect 56600 2825 56605 2830
rect 56365 2805 56605 2825
rect 56600 2800 56605 2805
rect 56635 2825 56640 2830
rect 57160 2830 57200 2835
rect 57160 2825 57165 2830
rect 56635 2805 57165 2825
rect 56635 2800 56640 2805
rect 56600 2795 56640 2800
rect 57160 2800 57165 2805
rect 57195 2800 57200 2830
rect 57160 2795 57200 2800
rect 55950 2780 55990 2785
rect 55950 2750 55955 2780
rect 55985 2775 55990 2780
rect 56745 2780 56785 2785
rect 56745 2775 56750 2780
rect 55985 2755 56750 2775
rect 55985 2750 55990 2755
rect 55950 2745 55990 2750
rect 56745 2750 56750 2755
rect 56780 2775 56785 2780
rect 57015 2780 57055 2785
rect 57015 2775 57020 2780
rect 56780 2755 57020 2775
rect 56780 2750 56785 2755
rect 56745 2745 56785 2750
rect 57015 2750 57020 2755
rect 57050 2775 57055 2780
rect 57810 2780 57850 2785
rect 57810 2775 57815 2780
rect 57050 2755 57815 2775
rect 57050 2750 57055 2755
rect 57015 2745 57055 2750
rect 57810 2750 57815 2755
rect 57845 2750 57850 2780
rect 57810 2745 57850 2750
rect 56850 2725 56890 2730
rect 56850 2695 56855 2725
rect 56885 2720 56890 2725
rect 56960 2725 57000 2730
rect 56960 2720 56965 2725
rect 56885 2700 56965 2720
rect 56885 2695 56890 2700
rect 56850 2690 56890 2695
rect 56960 2695 56965 2700
rect 56995 2695 57000 2725
rect 56960 2690 57000 2695
rect 56935 2670 56975 2675
rect 56935 2640 56940 2670
rect 56970 2665 56975 2670
rect 57210 2670 57250 2675
rect 57210 2665 57215 2670
rect 56970 2645 57215 2665
rect 56970 2640 56975 2645
rect 56935 2635 56975 2640
rect 57210 2640 57215 2645
rect 57245 2665 57250 2670
rect 57865 2670 57905 2675
rect 57865 2665 57870 2670
rect 57245 2645 57870 2665
rect 57245 2640 57250 2645
rect 57210 2635 57250 2640
rect 57865 2640 57870 2645
rect 57900 2640 57905 2670
rect 57865 2635 57905 2640
rect 56850 2615 56890 2620
rect 56850 2585 56855 2615
rect 56885 2585 56890 2615
rect 56850 2580 56890 2585
rect 54675 2550 54715 2555
rect 54675 2520 54680 2550
rect 54710 2545 54715 2550
rect 54785 2550 54825 2555
rect 54785 2545 54790 2550
rect 54710 2525 54790 2545
rect 54710 2520 54715 2525
rect 54675 2515 54715 2520
rect 54785 2520 54790 2525
rect 54820 2545 54825 2550
rect 54895 2550 54935 2555
rect 54895 2545 54900 2550
rect 54820 2525 54900 2545
rect 54820 2520 54825 2525
rect 54785 2515 54825 2520
rect 54895 2520 54900 2525
rect 54930 2545 54935 2550
rect 55005 2550 55045 2555
rect 55005 2545 55010 2550
rect 54930 2525 55010 2545
rect 54930 2520 54935 2525
rect 54895 2515 54935 2520
rect 55005 2520 55010 2525
rect 55040 2545 55045 2550
rect 55115 2550 55155 2555
rect 55115 2545 55120 2550
rect 55040 2525 55120 2545
rect 55040 2520 55045 2525
rect 55005 2515 55045 2520
rect 55115 2520 55120 2525
rect 55150 2545 55155 2550
rect 55225 2550 55265 2555
rect 55225 2545 55230 2550
rect 55150 2525 55230 2545
rect 55150 2520 55155 2525
rect 55115 2515 55155 2520
rect 55225 2520 55230 2525
rect 55260 2520 55265 2550
rect 55225 2515 55265 2520
rect 58535 2550 58575 2555
rect 58535 2520 58540 2550
rect 58570 2545 58575 2550
rect 58645 2550 58685 2555
rect 58645 2545 58650 2550
rect 58570 2525 58650 2545
rect 58570 2520 58575 2525
rect 58535 2515 58575 2520
rect 58645 2520 58650 2525
rect 58680 2545 58685 2550
rect 58755 2550 58795 2555
rect 58755 2545 58760 2550
rect 58680 2525 58760 2545
rect 58680 2520 58685 2525
rect 58645 2515 58685 2520
rect 58755 2520 58760 2525
rect 58790 2545 58795 2550
rect 58865 2550 58905 2555
rect 58865 2545 58870 2550
rect 58790 2525 58870 2545
rect 58790 2520 58795 2525
rect 58755 2515 58795 2520
rect 58865 2520 58870 2525
rect 58900 2545 58905 2550
rect 58975 2550 59015 2555
rect 58975 2545 58980 2550
rect 58900 2525 58980 2545
rect 58900 2520 58905 2525
rect 58865 2515 58905 2520
rect 58975 2520 58980 2525
rect 59010 2545 59015 2550
rect 59085 2550 59125 2555
rect 59085 2545 59090 2550
rect 59010 2525 59090 2545
rect 59010 2520 59015 2525
rect 58975 2515 59015 2520
rect 59085 2520 59090 2525
rect 59120 2520 59125 2550
rect 59085 2515 59125 2520
rect 54215 2470 56675 2475
rect 54215 2440 54220 2470
rect 54250 2440 54260 2470
rect 54290 2440 54300 2470
rect 54330 2440 54955 2470
rect 54985 2440 55405 2470
rect 55435 2440 55445 2470
rect 55475 2440 55485 2470
rect 55515 2440 56090 2470
rect 56120 2440 56145 2470
rect 56175 2440 56200 2470
rect 56230 2440 56255 2470
rect 56285 2440 56310 2470
rect 56340 2440 56365 2470
rect 56395 2440 56420 2470
rect 56450 2440 56475 2470
rect 56505 2440 56530 2470
rect 56560 2440 56585 2470
rect 56615 2440 56640 2470
rect 56670 2440 56675 2470
rect 54215 2430 56675 2440
rect 54215 2400 54220 2430
rect 54250 2400 54260 2430
rect 54290 2400 54300 2430
rect 54330 2400 54955 2430
rect 54985 2400 55405 2430
rect 55435 2400 55445 2430
rect 55475 2400 55485 2430
rect 55515 2400 56090 2430
rect 56120 2400 56145 2430
rect 56175 2400 56200 2430
rect 56230 2400 56255 2430
rect 56285 2400 56310 2430
rect 56340 2400 56365 2430
rect 56395 2400 56420 2430
rect 56450 2400 56475 2430
rect 56505 2400 56530 2430
rect 56560 2400 56585 2430
rect 56615 2400 56640 2430
rect 56670 2400 56675 2430
rect 54215 2390 56675 2400
rect 54215 2360 54220 2390
rect 54250 2360 54260 2390
rect 54290 2360 54300 2390
rect 54330 2360 54955 2390
rect 54985 2360 55405 2390
rect 55435 2360 55445 2390
rect 55475 2360 55485 2390
rect 55515 2360 56090 2390
rect 56120 2360 56145 2390
rect 56175 2360 56200 2390
rect 56230 2360 56255 2390
rect 56285 2360 56310 2390
rect 56340 2360 56365 2390
rect 56395 2360 56420 2390
rect 56450 2360 56475 2390
rect 56505 2360 56530 2390
rect 56560 2360 56585 2390
rect 56615 2360 56640 2390
rect 56670 2360 56675 2390
rect 54215 2355 56675 2360
rect 57125 2470 59585 2475
rect 57125 2440 57130 2470
rect 57160 2440 57185 2470
rect 57215 2440 57240 2470
rect 57270 2440 57295 2470
rect 57325 2440 57350 2470
rect 57380 2440 57405 2470
rect 57435 2440 57460 2470
rect 57490 2440 57515 2470
rect 57545 2440 57570 2470
rect 57600 2440 57625 2470
rect 57655 2440 57680 2470
rect 57710 2440 58285 2470
rect 58315 2440 58325 2470
rect 58355 2440 58365 2470
rect 58395 2440 58815 2470
rect 58845 2440 59470 2470
rect 59500 2440 59510 2470
rect 59540 2440 59550 2470
rect 59580 2440 59585 2470
rect 57125 2430 59585 2440
rect 57125 2400 57130 2430
rect 57160 2400 57185 2430
rect 57215 2400 57240 2430
rect 57270 2400 57295 2430
rect 57325 2400 57350 2430
rect 57380 2400 57405 2430
rect 57435 2400 57460 2430
rect 57490 2400 57515 2430
rect 57545 2400 57570 2430
rect 57600 2400 57625 2430
rect 57655 2400 57680 2430
rect 57710 2400 58285 2430
rect 58315 2400 58325 2430
rect 58355 2400 58365 2430
rect 58395 2400 58815 2430
rect 58845 2400 59470 2430
rect 59500 2400 59510 2430
rect 59540 2400 59550 2430
rect 59580 2400 59585 2430
rect 57125 2390 59585 2400
rect 57125 2360 57130 2390
rect 57160 2360 57185 2390
rect 57215 2360 57240 2390
rect 57270 2360 57295 2390
rect 57325 2360 57350 2390
rect 57380 2360 57405 2390
rect 57435 2360 57460 2390
rect 57490 2360 57515 2390
rect 57545 2360 57570 2390
rect 57600 2360 57625 2390
rect 57655 2360 57680 2390
rect 57710 2360 58285 2390
rect 58315 2360 58325 2390
rect 58355 2360 58365 2390
rect 58395 2360 58815 2390
rect 58845 2360 59470 2390
rect 59500 2360 59510 2390
rect 59540 2360 59550 2390
rect 59580 2360 59585 2390
rect 57125 2355 59585 2360
rect 53990 2320 55265 2325
rect 53990 2290 53995 2320
rect 54025 2290 54035 2320
rect 54065 2290 54080 2320
rect 54110 2290 54120 2320
rect 54150 2290 54165 2320
rect 54195 2290 54205 2320
rect 54235 2290 54680 2320
rect 54710 2290 54735 2320
rect 54765 2290 54790 2320
rect 54820 2290 54845 2320
rect 54875 2290 54900 2320
rect 54930 2290 54955 2320
rect 54985 2290 55010 2320
rect 55040 2290 55065 2320
rect 55095 2290 55120 2320
rect 55150 2290 55175 2320
rect 55205 2290 55230 2320
rect 55260 2290 55265 2320
rect 58535 2320 59810 2325
rect 53990 2280 55265 2290
rect 53990 2250 53995 2280
rect 54025 2250 54035 2280
rect 54065 2250 54080 2280
rect 54110 2250 54120 2280
rect 54150 2250 54165 2280
rect 54195 2250 54205 2280
rect 54235 2250 54680 2280
rect 54710 2250 54735 2280
rect 54765 2250 54790 2280
rect 54820 2250 54845 2280
rect 54875 2250 54900 2280
rect 54930 2250 54955 2280
rect 54985 2250 55010 2280
rect 55040 2250 55065 2280
rect 55095 2250 55120 2280
rect 55150 2250 55175 2280
rect 55205 2250 55230 2280
rect 55260 2250 55265 2280
rect 53990 2240 55265 2250
rect 53990 2210 53995 2240
rect 54025 2210 54035 2240
rect 54065 2210 54080 2240
rect 54110 2210 54120 2240
rect 54150 2210 54165 2240
rect 54195 2210 54205 2240
rect 54235 2210 54680 2240
rect 54710 2210 54735 2240
rect 54765 2210 54790 2240
rect 54820 2210 54845 2240
rect 54875 2210 54900 2240
rect 54930 2210 54955 2240
rect 54985 2210 55010 2240
rect 55040 2210 55065 2240
rect 55095 2210 55120 2240
rect 55150 2210 55175 2240
rect 55205 2210 55230 2240
rect 55260 2210 55265 2240
rect 53990 2205 55265 2210
rect 55670 2295 58130 2300
rect 55670 2265 55675 2295
rect 55705 2265 55715 2295
rect 55745 2265 55755 2295
rect 55785 2265 56775 2295
rect 56805 2265 56885 2295
rect 56915 2265 56995 2295
rect 57025 2265 58015 2295
rect 58045 2265 58055 2295
rect 58085 2265 58095 2295
rect 58125 2265 58130 2295
rect 55670 2255 58130 2265
rect 55670 2225 55675 2255
rect 55705 2225 55715 2255
rect 55745 2225 55755 2255
rect 55785 2225 56775 2255
rect 56805 2225 56885 2255
rect 56915 2225 56995 2255
rect 57025 2225 58015 2255
rect 58045 2225 58055 2255
rect 58085 2225 58095 2255
rect 58125 2225 58130 2255
rect 55670 2215 58130 2225
rect 54620 2185 55655 2190
rect 54620 2155 54625 2185
rect 54655 2155 55285 2185
rect 55315 2155 55540 2185
rect 55570 2155 55580 2185
rect 55610 2155 55620 2185
rect 55650 2155 55655 2185
rect 55670 2185 55675 2215
rect 55705 2185 55715 2215
rect 55745 2185 55755 2215
rect 55785 2185 56775 2215
rect 56805 2185 56885 2215
rect 56915 2185 56995 2215
rect 57025 2185 58015 2215
rect 58045 2185 58055 2215
rect 58085 2185 58095 2215
rect 58125 2185 58130 2215
rect 58535 2290 58540 2320
rect 58570 2290 58595 2320
rect 58625 2290 58650 2320
rect 58680 2290 58705 2320
rect 58735 2290 58760 2320
rect 58790 2290 58815 2320
rect 58845 2290 58870 2320
rect 58900 2290 58925 2320
rect 58955 2290 58980 2320
rect 59010 2290 59035 2320
rect 59065 2290 59090 2320
rect 59120 2290 59565 2320
rect 59595 2290 59605 2320
rect 59635 2290 59650 2320
rect 59680 2290 59690 2320
rect 59720 2290 59735 2320
rect 59765 2290 59775 2320
rect 59805 2290 59810 2320
rect 58535 2280 59810 2290
rect 58535 2250 58540 2280
rect 58570 2250 58595 2280
rect 58625 2250 58650 2280
rect 58680 2250 58705 2280
rect 58735 2250 58760 2280
rect 58790 2250 58815 2280
rect 58845 2250 58870 2280
rect 58900 2250 58925 2280
rect 58955 2250 58980 2280
rect 59010 2250 59035 2280
rect 59065 2250 59090 2280
rect 59120 2250 59565 2280
rect 59595 2250 59605 2280
rect 59635 2250 59650 2280
rect 59680 2250 59690 2280
rect 59720 2250 59735 2280
rect 59765 2250 59775 2280
rect 59805 2250 59810 2280
rect 58535 2240 59810 2250
rect 58535 2210 58540 2240
rect 58570 2210 58595 2240
rect 58625 2210 58650 2240
rect 58680 2210 58705 2240
rect 58735 2210 58760 2240
rect 58790 2210 58815 2240
rect 58845 2210 58870 2240
rect 58900 2210 58925 2240
rect 58955 2210 58980 2240
rect 59010 2210 59035 2240
rect 59065 2210 59090 2240
rect 59120 2210 59565 2240
rect 59595 2210 59605 2240
rect 59635 2210 59650 2240
rect 59680 2210 59690 2240
rect 59720 2210 59735 2240
rect 59765 2210 59775 2240
rect 59805 2210 59810 2240
rect 58535 2205 59810 2210
rect 55670 2180 58130 2185
rect 58145 2185 59180 2190
rect 54620 2145 55655 2155
rect 54620 2115 54625 2145
rect 54655 2115 55285 2145
rect 55315 2115 55540 2145
rect 55570 2115 55580 2145
rect 55610 2115 55620 2145
rect 55650 2115 55655 2145
rect 54620 2105 55655 2115
rect 54620 2075 54625 2105
rect 54655 2075 55285 2105
rect 55315 2075 55540 2105
rect 55570 2075 55580 2105
rect 55610 2075 55620 2105
rect 55650 2075 55655 2105
rect 54620 2070 55655 2075
rect 58145 2155 58150 2185
rect 58180 2155 58190 2185
rect 58220 2155 58230 2185
rect 58260 2155 58485 2185
rect 58515 2155 59145 2185
rect 59175 2155 59180 2185
rect 58145 2145 59180 2155
rect 58145 2115 58150 2145
rect 58180 2115 58190 2145
rect 58220 2115 58230 2145
rect 58260 2115 58485 2145
rect 58515 2115 59145 2145
rect 59175 2115 59180 2145
rect 58145 2105 59180 2115
rect 58145 2075 58150 2105
rect 58180 2075 58190 2105
rect 58220 2075 58230 2105
rect 58260 2075 58485 2105
rect 58515 2075 59145 2105
rect 59175 2075 59180 2105
rect 58145 2070 59180 2075
rect 53840 2050 55265 2055
rect 53840 2020 53845 2050
rect 53875 2020 53885 2050
rect 53915 2020 53925 2050
rect 53955 2020 54680 2050
rect 54710 2020 54790 2050
rect 54820 2020 54900 2050
rect 54930 2020 55010 2050
rect 55040 2020 55120 2050
rect 55150 2020 55230 2050
rect 55260 2020 55265 2050
rect 53840 2010 55265 2020
rect 53840 1980 53845 2010
rect 53875 1980 53885 2010
rect 53915 1980 53925 2010
rect 53955 1980 54680 2010
rect 54710 1980 54790 2010
rect 54820 1980 54900 2010
rect 54930 1980 55010 2010
rect 55040 1980 55120 2010
rect 55150 1980 55230 2010
rect 55260 1980 55265 2010
rect 53840 1970 55265 1980
rect 53840 1940 53845 1970
rect 53875 1940 53885 1970
rect 53915 1940 53925 1970
rect 53955 1940 54680 1970
rect 54710 1940 54790 1970
rect 54820 1940 54900 1970
rect 54930 1940 55010 1970
rect 55040 1940 55120 1970
rect 55150 1940 55230 1970
rect 55260 1940 55265 1970
rect 53840 1935 55265 1940
rect 55670 2050 55790 2055
rect 55670 2020 55675 2050
rect 55705 2020 55715 2050
rect 55745 2020 55755 2050
rect 55785 2020 55790 2050
rect 55670 2010 55790 2020
rect 55670 1980 55675 2010
rect 55705 1980 55715 2010
rect 55745 1980 55755 2010
rect 55785 1980 55790 2010
rect 58010 2050 59960 2055
rect 58010 2020 58015 2050
rect 58045 2020 58055 2050
rect 58085 2020 58095 2050
rect 58125 2020 58540 2050
rect 58570 2020 58650 2050
rect 58680 2020 58760 2050
rect 58790 2020 58870 2050
rect 58900 2020 58980 2050
rect 59010 2020 59090 2050
rect 59120 2020 59845 2050
rect 59875 2020 59885 2050
rect 59915 2020 59925 2050
rect 59955 2020 59960 2050
rect 58010 2010 59960 2020
rect 55670 1970 55790 1980
rect 55670 1940 55675 1970
rect 55705 1940 55715 1970
rect 55745 1940 55755 1970
rect 55785 1940 55790 1970
rect 55885 1985 55925 1990
rect 55885 1955 55890 1985
rect 55920 1980 55925 1985
rect 56040 1985 56070 1990
rect 55920 1960 56040 1980
rect 55920 1955 55925 1960
rect 55885 1950 55925 1955
rect 56690 1985 56720 1990
rect 56040 1950 56070 1955
rect 56140 1975 56180 1980
rect 56140 1945 56145 1975
rect 56175 1970 56180 1975
rect 56250 1975 56290 1980
rect 56250 1970 56255 1975
rect 56175 1950 56255 1970
rect 56175 1945 56180 1950
rect 56140 1940 56180 1945
rect 56250 1945 56255 1950
rect 56285 1970 56290 1975
rect 56360 1975 56400 1980
rect 56360 1970 56365 1975
rect 56285 1950 56365 1970
rect 56285 1945 56290 1950
rect 56250 1940 56290 1945
rect 56360 1945 56365 1950
rect 56395 1970 56400 1975
rect 56470 1975 56510 1980
rect 56470 1970 56475 1975
rect 56395 1950 56475 1970
rect 56395 1945 56400 1950
rect 56360 1940 56400 1945
rect 56470 1945 56475 1950
rect 56505 1970 56510 1975
rect 56580 1975 56620 1980
rect 56580 1970 56585 1975
rect 56505 1950 56585 1970
rect 56505 1945 56510 1950
rect 56470 1940 56510 1945
rect 56580 1945 56585 1950
rect 56615 1945 56620 1975
rect 57080 1985 57110 1990
rect 56720 1960 57080 1980
rect 56690 1950 56720 1955
rect 57730 1985 57760 1990
rect 57080 1950 57110 1955
rect 57180 1975 57220 1980
rect 56580 1940 56620 1945
rect 57180 1945 57185 1975
rect 57215 1970 57220 1975
rect 57290 1975 57330 1980
rect 57290 1970 57295 1975
rect 57215 1950 57295 1970
rect 57215 1945 57220 1950
rect 57180 1940 57220 1945
rect 57290 1945 57295 1950
rect 57325 1970 57330 1975
rect 57400 1975 57440 1980
rect 57400 1970 57405 1975
rect 57325 1950 57405 1970
rect 57325 1945 57330 1950
rect 57290 1940 57330 1945
rect 57400 1945 57405 1950
rect 57435 1970 57440 1975
rect 57510 1975 57550 1980
rect 57510 1970 57515 1975
rect 57435 1950 57515 1970
rect 57435 1945 57440 1950
rect 57400 1940 57440 1945
rect 57510 1945 57515 1950
rect 57545 1970 57550 1975
rect 57620 1975 57660 1980
rect 57620 1970 57625 1975
rect 57545 1950 57625 1970
rect 57545 1945 57550 1950
rect 57510 1940 57550 1945
rect 57620 1945 57625 1950
rect 57655 1945 57660 1975
rect 57730 1950 57760 1955
rect 58010 1980 58015 2010
rect 58045 1980 58055 2010
rect 58085 1980 58095 2010
rect 58125 1980 58540 2010
rect 58570 1980 58650 2010
rect 58680 1980 58760 2010
rect 58790 1980 58870 2010
rect 58900 1980 58980 2010
rect 59010 1980 59090 2010
rect 59120 1980 59845 2010
rect 59875 1980 59885 2010
rect 59915 1980 59925 2010
rect 59955 1980 59960 2010
rect 58010 1970 59960 1980
rect 57620 1940 57660 1945
rect 58010 1940 58015 1970
rect 58045 1940 58055 1970
rect 58085 1940 58095 1970
rect 58125 1940 58540 1970
rect 58570 1940 58650 1970
rect 58680 1940 58760 1970
rect 58790 1940 58870 1970
rect 58900 1940 58980 1970
rect 59010 1940 59090 1970
rect 59120 1940 59845 1970
rect 59875 1940 59885 1970
rect 59915 1940 59925 1970
rect 59955 1940 59960 1970
rect 55670 1935 55790 1940
rect 58010 1935 59960 1940
rect 54625 1930 54655 1935
rect 56085 1930 56125 1935
rect 54730 1915 54770 1920
rect 54730 1885 54735 1915
rect 54765 1910 54770 1915
rect 54840 1915 54880 1920
rect 54840 1910 54845 1915
rect 54765 1890 54845 1910
rect 54765 1885 54770 1890
rect 54730 1880 54770 1885
rect 54840 1885 54845 1890
rect 54875 1910 54880 1915
rect 54950 1915 54990 1920
rect 54950 1910 54955 1915
rect 54875 1890 54955 1910
rect 54875 1885 54880 1890
rect 54840 1880 54880 1885
rect 54950 1885 54955 1890
rect 54985 1910 54990 1915
rect 55060 1915 55100 1920
rect 55060 1910 55065 1915
rect 54985 1890 55065 1910
rect 54985 1885 54990 1890
rect 54950 1880 54990 1885
rect 55060 1885 55065 1890
rect 55095 1910 55100 1915
rect 55170 1915 55210 1920
rect 55170 1910 55175 1915
rect 55095 1890 55175 1910
rect 55095 1885 55100 1890
rect 55060 1880 55100 1885
rect 55170 1885 55175 1890
rect 55205 1885 55210 1915
rect 56085 1900 56090 1930
rect 56120 1925 56125 1930
rect 56195 1930 56235 1935
rect 56195 1925 56200 1930
rect 56120 1905 56200 1925
rect 56120 1900 56125 1905
rect 56085 1895 56125 1900
rect 56195 1900 56200 1905
rect 56230 1925 56235 1930
rect 56305 1930 56345 1935
rect 56305 1925 56310 1930
rect 56230 1905 56310 1925
rect 56230 1900 56235 1905
rect 56195 1895 56235 1900
rect 56305 1900 56310 1905
rect 56340 1925 56345 1930
rect 56415 1930 56455 1935
rect 56415 1925 56420 1930
rect 56340 1905 56420 1925
rect 56340 1900 56345 1905
rect 56305 1895 56345 1900
rect 56415 1900 56420 1905
rect 56450 1925 56455 1930
rect 56525 1930 56565 1935
rect 56525 1925 56530 1930
rect 56450 1905 56530 1925
rect 56450 1900 56455 1905
rect 56415 1895 56455 1900
rect 56525 1900 56530 1905
rect 56560 1925 56565 1930
rect 56635 1930 56675 1935
rect 56635 1925 56640 1930
rect 56560 1905 56640 1925
rect 56560 1900 56565 1905
rect 56525 1895 56565 1900
rect 56635 1900 56640 1905
rect 56670 1900 56675 1930
rect 56635 1895 56675 1900
rect 57125 1930 57165 1935
rect 57125 1900 57130 1930
rect 57160 1925 57165 1930
rect 57235 1930 57275 1935
rect 57235 1925 57240 1930
rect 57160 1905 57240 1925
rect 57160 1900 57165 1905
rect 57125 1895 57165 1900
rect 57235 1900 57240 1905
rect 57270 1925 57275 1930
rect 57345 1930 57385 1935
rect 57345 1925 57350 1930
rect 57270 1905 57350 1925
rect 57270 1900 57275 1905
rect 57235 1895 57275 1900
rect 57345 1900 57350 1905
rect 57380 1925 57385 1930
rect 57455 1930 57495 1935
rect 57455 1925 57460 1930
rect 57380 1905 57460 1925
rect 57380 1900 57385 1905
rect 57345 1895 57385 1900
rect 57455 1900 57460 1905
rect 57490 1925 57495 1930
rect 57565 1930 57605 1935
rect 57565 1925 57570 1930
rect 57490 1905 57570 1925
rect 57490 1900 57495 1905
rect 57455 1895 57495 1900
rect 57565 1900 57570 1905
rect 57600 1925 57605 1930
rect 57675 1930 57715 1935
rect 58485 1930 58515 1935
rect 59145 1930 59175 1935
rect 57675 1925 57680 1930
rect 57600 1905 57680 1925
rect 57600 1900 57605 1905
rect 57565 1895 57605 1900
rect 57675 1900 57680 1905
rect 57710 1900 57715 1930
rect 57675 1895 57715 1900
rect 58590 1915 58630 1920
rect 55170 1880 55210 1885
rect 58590 1885 58595 1915
rect 58625 1910 58630 1915
rect 58700 1915 58740 1920
rect 58700 1910 58705 1915
rect 58625 1890 58705 1910
rect 58625 1885 58630 1890
rect 58590 1880 58630 1885
rect 58700 1885 58705 1890
rect 58735 1910 58740 1915
rect 58810 1915 58850 1920
rect 58810 1910 58815 1915
rect 58735 1890 58815 1910
rect 58735 1885 58740 1890
rect 58700 1880 58740 1885
rect 58810 1885 58815 1890
rect 58845 1910 58850 1915
rect 58920 1915 58960 1920
rect 58920 1910 58925 1915
rect 58845 1890 58925 1910
rect 58845 1885 58850 1890
rect 58810 1880 58850 1885
rect 58920 1885 58925 1890
rect 58955 1910 58960 1915
rect 59030 1915 59070 1920
rect 59030 1910 59035 1915
rect 58955 1890 59035 1910
rect 58955 1885 58960 1890
rect 58920 1880 58960 1885
rect 59030 1885 59035 1890
rect 59065 1885 59070 1915
rect 59030 1880 59070 1885
rect 56140 1740 56180 1745
rect 53990 1710 54240 1720
rect 53990 1680 54000 1710
rect 54030 1680 54050 1710
rect 54080 1680 54100 1710
rect 54130 1680 54150 1710
rect 54180 1680 54200 1710
rect 54230 1680 54240 1710
rect 56140 1710 56145 1740
rect 56175 1735 56180 1740
rect 56250 1740 56290 1745
rect 56250 1735 56255 1740
rect 56175 1715 56255 1735
rect 56175 1710 56180 1715
rect 56140 1705 56180 1710
rect 56250 1710 56255 1715
rect 56285 1735 56290 1740
rect 56360 1740 56400 1745
rect 56360 1735 56365 1740
rect 56285 1715 56365 1735
rect 56285 1710 56290 1715
rect 56250 1705 56290 1710
rect 56360 1710 56365 1715
rect 56395 1735 56400 1740
rect 56470 1740 56510 1745
rect 56470 1735 56475 1740
rect 56395 1715 56475 1735
rect 56395 1710 56400 1715
rect 56360 1705 56400 1710
rect 56470 1710 56475 1715
rect 56505 1735 56510 1740
rect 56580 1740 56620 1745
rect 56580 1735 56585 1740
rect 56505 1715 56585 1735
rect 56505 1710 56510 1715
rect 56470 1705 56510 1710
rect 56580 1710 56585 1715
rect 56615 1710 56620 1740
rect 56580 1705 56620 1710
rect 57180 1740 57220 1745
rect 57180 1710 57185 1740
rect 57215 1735 57220 1740
rect 57290 1740 57330 1745
rect 57290 1735 57295 1740
rect 57215 1715 57295 1735
rect 57215 1710 57220 1715
rect 57180 1705 57220 1710
rect 57290 1710 57295 1715
rect 57325 1735 57330 1740
rect 57400 1740 57440 1745
rect 57400 1735 57405 1740
rect 57325 1715 57405 1735
rect 57325 1710 57330 1715
rect 57290 1705 57330 1710
rect 57400 1710 57405 1715
rect 57435 1735 57440 1740
rect 57510 1740 57550 1745
rect 57510 1735 57515 1740
rect 57435 1715 57515 1735
rect 57435 1710 57440 1715
rect 57400 1705 57440 1710
rect 57510 1710 57515 1715
rect 57545 1735 57550 1740
rect 57620 1740 57660 1745
rect 57620 1735 57625 1740
rect 57545 1715 57625 1735
rect 57545 1710 57550 1715
rect 57510 1705 57550 1710
rect 57620 1710 57625 1715
rect 57655 1710 57660 1740
rect 57620 1705 57660 1710
rect 59560 1710 59810 1720
rect 53990 1660 54240 1680
rect 56085 1695 56125 1700
rect 56085 1665 56090 1695
rect 56120 1690 56125 1695
rect 56195 1695 56235 1700
rect 56195 1690 56200 1695
rect 56120 1670 56200 1690
rect 56120 1665 56125 1670
rect 53990 1630 54000 1660
rect 54030 1630 54050 1660
rect 54080 1630 54100 1660
rect 54130 1630 54150 1660
rect 54180 1630 54200 1660
rect 54230 1630 54240 1660
rect 53990 1610 54240 1630
rect 54485 1660 54525 1665
rect 54485 1630 54490 1660
rect 54520 1655 54525 1660
rect 54730 1660 54770 1665
rect 54730 1655 54735 1660
rect 54520 1635 54735 1655
rect 54520 1630 54525 1635
rect 54485 1625 54525 1630
rect 54730 1630 54735 1635
rect 54765 1655 54770 1660
rect 54840 1660 54880 1665
rect 54840 1655 54845 1660
rect 54765 1635 54845 1655
rect 54765 1630 54770 1635
rect 54730 1625 54770 1630
rect 54840 1630 54845 1635
rect 54875 1655 54880 1660
rect 54950 1660 54990 1665
rect 54950 1655 54955 1660
rect 54875 1635 54955 1655
rect 54875 1630 54880 1635
rect 54840 1625 54880 1630
rect 54950 1630 54955 1635
rect 54985 1655 54990 1660
rect 55060 1660 55100 1665
rect 55060 1655 55065 1660
rect 54985 1635 55065 1655
rect 54985 1630 54990 1635
rect 54950 1625 54990 1630
rect 55060 1630 55065 1635
rect 55095 1655 55100 1660
rect 55170 1660 55210 1665
rect 56085 1660 56125 1665
rect 56195 1665 56200 1670
rect 56230 1690 56235 1695
rect 56305 1695 56345 1700
rect 56305 1690 56310 1695
rect 56230 1670 56310 1690
rect 56230 1665 56235 1670
rect 56195 1660 56235 1665
rect 56305 1665 56310 1670
rect 56340 1690 56345 1695
rect 56415 1695 56455 1700
rect 56415 1690 56420 1695
rect 56340 1670 56420 1690
rect 56340 1665 56345 1670
rect 56305 1660 56345 1665
rect 56415 1665 56420 1670
rect 56450 1690 56455 1695
rect 56525 1695 56565 1700
rect 56525 1690 56530 1695
rect 56450 1670 56530 1690
rect 56450 1665 56455 1670
rect 56415 1660 56455 1665
rect 56525 1665 56530 1670
rect 56560 1690 56565 1695
rect 56635 1695 56675 1700
rect 56635 1690 56640 1695
rect 56560 1670 56640 1690
rect 56560 1665 56565 1670
rect 56525 1660 56565 1665
rect 56635 1665 56640 1670
rect 56670 1665 56675 1695
rect 56635 1660 56675 1665
rect 57125 1695 57165 1700
rect 57125 1665 57130 1695
rect 57160 1690 57165 1695
rect 57235 1695 57275 1700
rect 57235 1690 57240 1695
rect 57160 1670 57240 1690
rect 57160 1665 57165 1670
rect 57125 1660 57165 1665
rect 57235 1665 57240 1670
rect 57270 1690 57275 1695
rect 57345 1695 57385 1700
rect 57345 1690 57350 1695
rect 57270 1670 57350 1690
rect 57270 1665 57275 1670
rect 57235 1660 57275 1665
rect 57345 1665 57350 1670
rect 57380 1690 57385 1695
rect 57455 1695 57495 1700
rect 57455 1690 57460 1695
rect 57380 1670 57460 1690
rect 57380 1665 57385 1670
rect 57345 1660 57385 1665
rect 57455 1665 57460 1670
rect 57490 1690 57495 1695
rect 57565 1695 57605 1700
rect 57565 1690 57570 1695
rect 57490 1670 57570 1690
rect 57490 1665 57495 1670
rect 57455 1660 57495 1665
rect 57565 1665 57570 1670
rect 57600 1690 57605 1695
rect 57675 1695 57715 1700
rect 57675 1690 57680 1695
rect 57600 1670 57680 1690
rect 57600 1665 57605 1670
rect 57565 1660 57605 1665
rect 57675 1665 57680 1670
rect 57710 1665 57715 1695
rect 59560 1680 59570 1710
rect 59600 1680 59620 1710
rect 59650 1680 59670 1710
rect 59700 1680 59720 1710
rect 59750 1680 59770 1710
rect 59800 1680 59810 1710
rect 57675 1660 57715 1665
rect 58590 1660 58630 1665
rect 55170 1655 55175 1660
rect 55095 1635 55175 1655
rect 55095 1630 55100 1635
rect 55060 1625 55100 1630
rect 55170 1630 55175 1635
rect 55205 1630 55210 1660
rect 55170 1625 55210 1630
rect 55670 1640 58130 1645
rect 53990 1580 54000 1610
rect 54030 1580 54050 1610
rect 54080 1580 54100 1610
rect 54130 1580 54150 1610
rect 54180 1580 54200 1610
rect 54230 1580 54240 1610
rect 55670 1610 55675 1640
rect 55705 1610 55715 1640
rect 55745 1610 55755 1640
rect 55785 1610 56035 1640
rect 56065 1610 56695 1640
rect 56725 1610 57075 1640
rect 57105 1610 57735 1640
rect 57765 1610 58015 1640
rect 58045 1610 58055 1640
rect 58085 1610 58095 1640
rect 58125 1610 58130 1640
rect 58590 1630 58595 1660
rect 58625 1655 58630 1660
rect 58700 1660 58740 1665
rect 58700 1655 58705 1660
rect 58625 1635 58705 1655
rect 58625 1630 58630 1635
rect 58590 1625 58630 1630
rect 58700 1630 58705 1635
rect 58735 1655 58740 1660
rect 58810 1660 58850 1665
rect 58810 1655 58815 1660
rect 58735 1635 58815 1655
rect 58735 1630 58740 1635
rect 58700 1625 58740 1630
rect 58810 1630 58815 1635
rect 58845 1655 58850 1660
rect 58920 1660 58960 1665
rect 58920 1655 58925 1660
rect 58845 1635 58925 1655
rect 58845 1630 58850 1635
rect 58810 1625 58850 1630
rect 58920 1630 58925 1635
rect 58955 1655 58960 1660
rect 59030 1660 59070 1665
rect 59030 1655 59035 1660
rect 58955 1635 59035 1655
rect 58955 1630 58960 1635
rect 58920 1625 58960 1630
rect 59030 1630 59035 1635
rect 59065 1655 59070 1660
rect 59275 1660 59315 1665
rect 59275 1655 59280 1660
rect 59065 1635 59280 1655
rect 59065 1630 59070 1635
rect 59030 1625 59070 1630
rect 59275 1630 59280 1635
rect 59310 1630 59315 1660
rect 59275 1625 59315 1630
rect 59560 1660 59810 1680
rect 59560 1630 59570 1660
rect 59600 1630 59620 1660
rect 59650 1630 59670 1660
rect 59700 1630 59720 1660
rect 59750 1630 59770 1660
rect 59800 1630 59810 1660
rect 55670 1600 58130 1610
rect 59560 1610 59810 1630
rect 53990 1570 54240 1580
rect 55115 1595 55520 1600
rect 55115 1565 55120 1595
rect 55150 1565 55405 1595
rect 55435 1565 55445 1595
rect 55475 1565 55485 1595
rect 55515 1565 55520 1595
rect 55115 1555 55520 1565
rect 55115 1525 55120 1555
rect 55150 1525 55405 1555
rect 55435 1525 55445 1555
rect 55475 1525 55485 1555
rect 55515 1525 55520 1555
rect 55670 1570 55675 1600
rect 55705 1570 55715 1600
rect 55745 1570 55755 1600
rect 55785 1570 56035 1600
rect 56065 1570 56695 1600
rect 56725 1570 57075 1600
rect 57105 1570 57735 1600
rect 57765 1570 58015 1600
rect 58045 1570 58055 1600
rect 58085 1570 58095 1600
rect 58125 1570 58130 1600
rect 55670 1560 58130 1570
rect 55670 1530 55675 1560
rect 55705 1530 55715 1560
rect 55745 1530 55755 1560
rect 55785 1530 56035 1560
rect 56065 1530 56695 1560
rect 56725 1530 57075 1560
rect 57105 1530 57735 1560
rect 57765 1530 58015 1560
rect 58045 1530 58055 1560
rect 58085 1530 58095 1560
rect 58125 1530 58130 1560
rect 55670 1525 58130 1530
rect 58280 1595 58685 1600
rect 58280 1565 58285 1595
rect 58315 1565 58325 1595
rect 58355 1565 58365 1595
rect 58395 1565 58650 1595
rect 58680 1565 58685 1595
rect 59560 1580 59570 1610
rect 59600 1580 59620 1610
rect 59650 1580 59670 1610
rect 59700 1580 59720 1610
rect 59750 1580 59770 1610
rect 59800 1580 59810 1610
rect 59560 1570 59810 1580
rect 58280 1555 58685 1565
rect 58280 1525 58285 1555
rect 58315 1525 58325 1555
rect 58355 1525 58365 1555
rect 58395 1525 58650 1555
rect 58680 1525 58685 1555
rect 55115 1520 55520 1525
rect 58280 1520 58685 1525
rect 55670 1485 58130 1490
rect 54530 1475 54570 1480
rect 54530 1445 54535 1475
rect 54565 1470 54570 1475
rect 54730 1475 54770 1480
rect 54730 1470 54735 1475
rect 54565 1450 54735 1470
rect 54565 1445 54570 1450
rect 54530 1440 54570 1445
rect 54730 1445 54735 1450
rect 54765 1470 54770 1475
rect 54840 1475 54880 1480
rect 54840 1470 54845 1475
rect 54765 1450 54845 1470
rect 54765 1445 54770 1450
rect 54730 1440 54770 1445
rect 54840 1445 54845 1450
rect 54875 1470 54880 1475
rect 54950 1475 54990 1480
rect 54950 1470 54955 1475
rect 54875 1450 54955 1470
rect 54875 1445 54880 1450
rect 54840 1440 54880 1445
rect 54950 1445 54955 1450
rect 54985 1470 54990 1475
rect 55060 1475 55100 1480
rect 55060 1470 55065 1475
rect 54985 1450 55065 1470
rect 54985 1445 54990 1450
rect 54950 1440 54990 1445
rect 55060 1445 55065 1450
rect 55095 1470 55100 1475
rect 55170 1475 55210 1480
rect 55170 1470 55175 1475
rect 55095 1450 55175 1470
rect 55095 1445 55100 1450
rect 55060 1440 55100 1445
rect 55170 1445 55175 1450
rect 55205 1445 55210 1475
rect 55170 1440 55210 1445
rect 55670 1455 55675 1485
rect 55705 1455 55715 1485
rect 55745 1455 55755 1485
rect 55785 1455 56885 1485
rect 56915 1455 58015 1485
rect 58045 1455 58055 1485
rect 58085 1455 58095 1485
rect 58125 1455 58130 1485
rect 55670 1445 58130 1455
rect 55670 1415 55675 1445
rect 55705 1415 55715 1445
rect 55745 1415 55755 1445
rect 55785 1415 56885 1445
rect 56915 1415 58015 1445
rect 58045 1415 58055 1445
rect 58085 1415 58095 1445
rect 58125 1415 58130 1445
rect 58590 1475 58630 1480
rect 58590 1445 58595 1475
rect 58625 1470 58630 1475
rect 58700 1475 58740 1480
rect 58700 1470 58705 1475
rect 58625 1450 58705 1470
rect 58625 1445 58630 1450
rect 58590 1440 58630 1445
rect 58700 1445 58705 1450
rect 58735 1470 58740 1475
rect 58810 1475 58850 1480
rect 58810 1470 58815 1475
rect 58735 1450 58815 1470
rect 58735 1445 58740 1450
rect 58700 1440 58740 1445
rect 58810 1445 58815 1450
rect 58845 1470 58850 1475
rect 58920 1475 58960 1480
rect 58920 1470 58925 1475
rect 58845 1450 58925 1470
rect 58845 1445 58850 1450
rect 58810 1440 58850 1445
rect 58920 1445 58925 1450
rect 58955 1470 58960 1475
rect 59030 1475 59070 1480
rect 59030 1470 59035 1475
rect 58955 1450 59035 1470
rect 58955 1445 58960 1450
rect 58920 1440 58960 1445
rect 59030 1445 59035 1450
rect 59065 1470 59070 1475
rect 59230 1475 59270 1480
rect 59230 1470 59235 1475
rect 59065 1450 59235 1470
rect 59065 1445 59070 1450
rect 59030 1440 59070 1445
rect 59230 1445 59235 1450
rect 59265 1445 59270 1475
rect 59230 1440 59270 1445
rect 55670 1405 58130 1415
rect 55670 1375 55675 1405
rect 55705 1375 55715 1405
rect 55745 1375 55755 1405
rect 55785 1375 56885 1405
rect 56915 1375 58015 1405
rect 58045 1375 58055 1405
rect 58085 1375 58095 1405
rect 58125 1375 58130 1405
rect 55670 1370 58130 1375
rect 56145 1315 56175 1320
rect 56085 1305 56125 1310
rect 56040 1295 56070 1300
rect 56030 1270 56040 1290
rect 56085 1275 56090 1305
rect 56120 1300 56125 1305
rect 56120 1285 56145 1300
rect 56255 1315 56285 1320
rect 56195 1305 56235 1310
rect 56195 1300 56200 1305
rect 56175 1285 56200 1300
rect 56120 1280 56200 1285
rect 56120 1275 56125 1280
rect 56085 1270 56125 1275
rect 56195 1275 56200 1280
rect 56230 1300 56235 1305
rect 56230 1285 56255 1300
rect 56365 1315 56395 1320
rect 56305 1305 56345 1310
rect 56305 1300 56310 1305
rect 56285 1285 56310 1300
rect 56230 1280 56310 1285
rect 56230 1275 56235 1280
rect 56195 1270 56235 1275
rect 56305 1275 56310 1280
rect 56340 1300 56345 1305
rect 56340 1285 56365 1300
rect 56475 1315 56505 1320
rect 56415 1305 56455 1310
rect 56415 1300 56420 1305
rect 56395 1285 56420 1300
rect 56340 1280 56420 1285
rect 56340 1275 56345 1280
rect 56305 1270 56345 1275
rect 56415 1275 56420 1280
rect 56450 1300 56455 1305
rect 56450 1285 56475 1300
rect 56585 1315 56615 1320
rect 56525 1305 56565 1310
rect 56525 1300 56530 1305
rect 56505 1285 56530 1300
rect 56450 1280 56530 1285
rect 56450 1275 56455 1280
rect 56415 1270 56455 1275
rect 56525 1275 56530 1280
rect 56560 1300 56565 1305
rect 56560 1285 56585 1300
rect 57185 1315 57215 1320
rect 56635 1305 56675 1310
rect 56635 1300 56640 1305
rect 56615 1285 56640 1300
rect 56560 1280 56640 1285
rect 56560 1275 56565 1280
rect 56525 1270 56565 1275
rect 56635 1275 56640 1280
rect 56670 1275 56675 1305
rect 56635 1270 56675 1275
rect 56690 1305 56720 1310
rect 56840 1305 56870 1310
rect 56720 1280 56840 1300
rect 56690 1270 56720 1275
rect 56840 1270 56870 1275
rect 56930 1305 56960 1310
rect 57080 1305 57110 1310
rect 56960 1280 57080 1300
rect 56930 1270 56960 1275
rect 57080 1270 57110 1275
rect 57125 1305 57165 1310
rect 57125 1275 57130 1305
rect 57160 1300 57165 1305
rect 57160 1285 57185 1300
rect 57295 1315 57325 1320
rect 57235 1305 57275 1310
rect 57235 1300 57240 1305
rect 57215 1285 57240 1300
rect 57160 1280 57240 1285
rect 57160 1275 57165 1280
rect 57125 1270 57165 1275
rect 57235 1275 57240 1280
rect 57270 1300 57275 1305
rect 57270 1285 57295 1300
rect 57405 1315 57435 1320
rect 57345 1305 57385 1310
rect 57345 1300 57350 1305
rect 57325 1285 57350 1300
rect 57270 1280 57350 1285
rect 57270 1275 57275 1280
rect 57235 1270 57275 1275
rect 57345 1275 57350 1280
rect 57380 1300 57385 1305
rect 57380 1285 57405 1300
rect 57515 1315 57545 1320
rect 57455 1305 57495 1310
rect 57455 1300 57460 1305
rect 57435 1285 57460 1300
rect 57380 1280 57460 1285
rect 57380 1275 57385 1280
rect 57345 1270 57385 1275
rect 57455 1275 57460 1280
rect 57490 1300 57495 1305
rect 57490 1285 57515 1300
rect 57625 1315 57655 1320
rect 57565 1305 57605 1310
rect 57565 1300 57570 1305
rect 57545 1285 57570 1300
rect 57490 1280 57570 1285
rect 57490 1275 57495 1280
rect 57455 1270 57495 1275
rect 57565 1275 57570 1280
rect 57600 1300 57605 1305
rect 57600 1285 57625 1300
rect 57675 1305 57715 1310
rect 57675 1300 57680 1305
rect 57655 1285 57680 1300
rect 57600 1280 57680 1285
rect 57600 1275 57605 1280
rect 57565 1270 57605 1275
rect 57675 1275 57680 1280
rect 57710 1275 57715 1305
rect 57675 1270 57715 1275
rect 57730 1295 57760 1300
rect 57760 1270 57770 1290
rect 56040 1260 56070 1265
rect 56140 1260 56180 1265
rect 56140 1230 56145 1260
rect 56175 1255 56180 1260
rect 56250 1260 56290 1265
rect 56250 1255 56255 1260
rect 56175 1235 56255 1255
rect 56175 1230 56180 1235
rect 56140 1225 56180 1230
rect 56250 1230 56255 1235
rect 56285 1255 56290 1260
rect 56360 1260 56400 1265
rect 56360 1255 56365 1260
rect 56285 1235 56365 1255
rect 56285 1230 56290 1235
rect 56250 1225 56290 1230
rect 56360 1230 56365 1235
rect 56395 1255 56400 1260
rect 56470 1260 56510 1265
rect 56470 1255 56475 1260
rect 56395 1235 56475 1255
rect 56395 1230 56400 1235
rect 56360 1225 56400 1230
rect 56470 1230 56475 1235
rect 56505 1255 56510 1260
rect 56580 1260 56620 1265
rect 56580 1255 56585 1260
rect 56505 1235 56585 1255
rect 56505 1230 56510 1235
rect 56470 1225 56510 1230
rect 56580 1230 56585 1235
rect 56615 1255 56620 1260
rect 57180 1260 57220 1265
rect 57180 1255 57185 1260
rect 56615 1235 57185 1255
rect 56615 1230 56620 1235
rect 56580 1225 56620 1230
rect 57180 1230 57185 1235
rect 57215 1255 57220 1260
rect 57290 1260 57330 1265
rect 57290 1255 57295 1260
rect 57215 1235 57295 1255
rect 57215 1230 57220 1235
rect 57180 1225 57220 1230
rect 57290 1230 57295 1235
rect 57325 1255 57330 1260
rect 57400 1260 57440 1265
rect 57400 1255 57405 1260
rect 57325 1235 57405 1255
rect 57325 1230 57330 1235
rect 57290 1225 57330 1230
rect 57400 1230 57405 1235
rect 57435 1255 57440 1260
rect 57510 1260 57550 1265
rect 57510 1255 57515 1260
rect 57435 1235 57515 1255
rect 57435 1230 57440 1235
rect 57400 1225 57440 1230
rect 57510 1230 57515 1235
rect 57545 1255 57550 1260
rect 57620 1260 57660 1265
rect 57730 1260 57760 1265
rect 57620 1255 57625 1260
rect 57545 1235 57625 1255
rect 57545 1230 57550 1235
rect 57510 1225 57550 1230
rect 57620 1230 57625 1235
rect 57655 1230 57660 1260
rect 57620 1225 57660 1230
rect 54255 1165 54290 1166
rect 59510 1165 59545 1166
rect 54255 1160 54350 1165
rect 54290 1125 54315 1160
rect 54255 1120 54350 1125
rect 54375 1160 54410 1165
rect 54375 1120 54410 1125
rect 54435 1160 54470 1165
rect 59330 1160 59365 1165
rect 54530 1155 54570 1160
rect 54530 1150 54535 1155
rect 54470 1130 54535 1150
rect 54435 1120 54470 1125
rect 54530 1125 54535 1130
rect 54565 1125 54570 1155
rect 59230 1155 59270 1160
rect 54530 1120 54570 1125
rect 54730 1135 54770 1140
rect 54730 1105 54735 1135
rect 54765 1130 54770 1135
rect 54840 1135 54880 1140
rect 54840 1130 54845 1135
rect 54765 1110 54845 1130
rect 54765 1105 54770 1110
rect 54730 1100 54770 1105
rect 54840 1105 54845 1110
rect 54875 1130 54880 1135
rect 54950 1135 54990 1140
rect 54950 1130 54955 1135
rect 54875 1110 54955 1130
rect 54875 1105 54880 1110
rect 54840 1100 54880 1105
rect 54950 1105 54955 1110
rect 54985 1130 54990 1135
rect 55060 1135 55100 1140
rect 55060 1130 55065 1135
rect 54985 1110 55065 1130
rect 54985 1105 54990 1110
rect 54950 1100 54990 1105
rect 55060 1105 55065 1110
rect 55095 1130 55100 1135
rect 55170 1135 55210 1140
rect 55170 1130 55175 1135
rect 55095 1110 55175 1130
rect 55095 1105 55100 1110
rect 55060 1100 55100 1105
rect 55170 1105 55175 1110
rect 55205 1105 55210 1135
rect 55170 1100 55210 1105
rect 58590 1135 58630 1140
rect 58590 1105 58595 1135
rect 58625 1130 58630 1135
rect 58700 1135 58740 1140
rect 58700 1130 58705 1135
rect 58625 1110 58705 1130
rect 58625 1105 58630 1110
rect 58590 1100 58630 1105
rect 58700 1105 58705 1110
rect 58735 1130 58740 1135
rect 58810 1135 58850 1140
rect 58810 1130 58815 1135
rect 58735 1110 58815 1130
rect 58735 1105 58740 1110
rect 58700 1100 58740 1105
rect 58810 1105 58815 1110
rect 58845 1130 58850 1135
rect 58920 1135 58960 1140
rect 58920 1130 58925 1135
rect 58845 1110 58925 1130
rect 58845 1105 58850 1110
rect 58810 1100 58850 1105
rect 58920 1105 58925 1110
rect 58955 1130 58960 1135
rect 59030 1135 59070 1140
rect 59030 1130 59035 1135
rect 58955 1110 59035 1130
rect 58955 1105 58960 1110
rect 58920 1100 58960 1105
rect 59030 1105 59035 1110
rect 59065 1105 59070 1135
rect 59230 1125 59235 1155
rect 59265 1150 59270 1155
rect 59265 1130 59330 1150
rect 59265 1125 59270 1130
rect 59230 1120 59270 1125
rect 59330 1120 59365 1125
rect 59390 1160 59425 1165
rect 59390 1120 59425 1125
rect 59450 1160 59545 1165
rect 59485 1125 59510 1160
rect 59450 1120 59545 1125
rect 59030 1100 59070 1105
rect 54375 1085 54415 1090
rect 54375 1055 54380 1085
rect 54410 1075 54415 1085
rect 54485 1085 54525 1090
rect 59275 1085 59315 1090
rect 54485 1075 54490 1085
rect 54410 1060 54490 1075
rect 54410 1055 54415 1060
rect 54375 1050 54415 1055
rect 54485 1055 54490 1060
rect 54520 1055 54525 1085
rect 58145 1080 59125 1085
rect 54485 1050 54525 1055
rect 54675 1075 55655 1080
rect 54675 1045 54680 1075
rect 54710 1045 54790 1075
rect 54820 1045 54900 1075
rect 54930 1045 55010 1075
rect 55040 1045 55120 1075
rect 55150 1045 55230 1075
rect 55260 1045 55540 1075
rect 55570 1045 55580 1075
rect 55610 1045 55620 1075
rect 55650 1045 55655 1075
rect 54675 1035 55655 1045
rect 54675 1005 54680 1035
rect 54710 1005 54790 1035
rect 54820 1005 54900 1035
rect 54930 1005 55010 1035
rect 55040 1005 55120 1035
rect 55150 1005 55230 1035
rect 55260 1005 55540 1035
rect 55570 1005 55580 1035
rect 55610 1005 55620 1035
rect 55650 1005 55655 1035
rect 56085 1065 56125 1070
rect 56085 1035 56090 1065
rect 56120 1060 56125 1065
rect 56195 1065 56235 1070
rect 56195 1060 56200 1065
rect 56120 1040 56200 1060
rect 56120 1035 56125 1040
rect 56085 1030 56125 1035
rect 56195 1035 56200 1040
rect 56230 1060 56235 1065
rect 56305 1065 56345 1070
rect 56305 1060 56310 1065
rect 56230 1040 56310 1060
rect 56230 1035 56235 1040
rect 56195 1030 56235 1035
rect 56305 1035 56310 1040
rect 56340 1060 56345 1065
rect 56415 1065 56455 1070
rect 56415 1060 56420 1065
rect 56340 1040 56420 1060
rect 56340 1035 56345 1040
rect 56305 1030 56345 1035
rect 56415 1035 56420 1040
rect 56450 1060 56455 1065
rect 56525 1065 56565 1070
rect 56525 1060 56530 1065
rect 56450 1040 56530 1060
rect 56450 1035 56455 1040
rect 56415 1030 56455 1035
rect 56525 1035 56530 1040
rect 56560 1060 56565 1065
rect 56635 1065 56675 1070
rect 56635 1060 56640 1065
rect 56560 1040 56640 1060
rect 56560 1035 56565 1040
rect 56525 1030 56565 1035
rect 56635 1035 56640 1040
rect 56670 1035 56675 1065
rect 56635 1030 56675 1035
rect 56825 1065 56865 1070
rect 56825 1035 56830 1065
rect 56860 1060 56865 1065
rect 56935 1065 56975 1070
rect 56935 1060 56940 1065
rect 56860 1040 56940 1060
rect 56860 1035 56865 1040
rect 56825 1030 56865 1035
rect 56935 1035 56940 1040
rect 56970 1035 56975 1065
rect 56935 1030 56975 1035
rect 57125 1065 57165 1070
rect 57125 1035 57130 1065
rect 57160 1060 57165 1065
rect 57235 1065 57275 1070
rect 57235 1060 57240 1065
rect 57160 1040 57240 1060
rect 57160 1035 57165 1040
rect 57125 1030 57165 1035
rect 57235 1035 57240 1040
rect 57270 1060 57275 1065
rect 57345 1065 57385 1070
rect 57345 1060 57350 1065
rect 57270 1040 57350 1060
rect 57270 1035 57275 1040
rect 57235 1030 57275 1035
rect 57345 1035 57350 1040
rect 57380 1060 57385 1065
rect 57455 1065 57495 1070
rect 57455 1060 57460 1065
rect 57380 1040 57460 1060
rect 57380 1035 57385 1040
rect 57345 1030 57385 1035
rect 57455 1035 57460 1040
rect 57490 1060 57495 1065
rect 57565 1065 57605 1070
rect 57565 1060 57570 1065
rect 57490 1040 57570 1060
rect 57490 1035 57495 1040
rect 57455 1030 57495 1035
rect 57565 1035 57570 1040
rect 57600 1060 57605 1065
rect 57675 1065 57715 1070
rect 57675 1060 57680 1065
rect 57600 1040 57680 1060
rect 57600 1035 57605 1040
rect 57565 1030 57605 1035
rect 57675 1035 57680 1040
rect 57710 1035 57715 1065
rect 57675 1030 57715 1035
rect 58145 1050 58150 1080
rect 58180 1050 58190 1080
rect 58220 1050 58230 1080
rect 58260 1050 58540 1080
rect 58570 1050 58650 1080
rect 58680 1050 58760 1080
rect 58790 1050 58870 1080
rect 58900 1050 58980 1080
rect 59010 1050 59090 1080
rect 59120 1050 59125 1080
rect 59275 1055 59280 1085
rect 59310 1080 59315 1085
rect 59385 1085 59425 1090
rect 59385 1080 59390 1085
rect 59310 1060 59390 1080
rect 59310 1055 59315 1060
rect 59275 1050 59315 1055
rect 59385 1055 59390 1060
rect 59420 1055 59425 1085
rect 59385 1050 59425 1055
rect 58145 1040 59125 1050
rect 54675 995 55655 1005
rect 58145 1010 58150 1040
rect 58180 1010 58190 1040
rect 58220 1010 58230 1040
rect 58260 1010 58540 1040
rect 58570 1010 58650 1040
rect 58680 1010 58760 1040
rect 58790 1010 58870 1040
rect 58900 1010 58980 1040
rect 59010 1010 59090 1040
rect 59120 1010 59125 1040
rect 58145 1000 59125 1010
rect 54675 965 54680 995
rect 54710 965 54790 995
rect 54820 965 54900 995
rect 54930 965 55010 995
rect 55040 965 55120 995
rect 55150 965 55230 995
rect 55260 965 55540 995
rect 55570 965 55580 995
rect 55610 965 55620 995
rect 55650 965 55655 995
rect 54675 960 55655 965
rect 56140 995 57660 1000
rect 56140 965 56145 995
rect 56175 965 56255 995
rect 56285 965 56365 995
rect 56395 965 56475 995
rect 56505 965 56585 995
rect 56615 965 57185 995
rect 57215 965 57295 995
rect 57325 965 57405 995
rect 57435 965 57515 995
rect 57545 965 57625 995
rect 57655 965 57660 995
rect 58145 970 58150 1000
rect 58180 970 58190 1000
rect 58220 970 58230 1000
rect 58260 970 58540 1000
rect 58570 970 58650 1000
rect 58680 970 58760 1000
rect 58790 970 58870 1000
rect 58900 970 58980 1000
rect 59010 970 59090 1000
rect 59120 970 59125 1000
rect 58145 965 59125 970
rect 56140 960 57660 965
rect 53840 940 59960 945
rect 53840 910 53845 940
rect 53875 910 53885 940
rect 53915 910 53925 940
rect 53955 910 54625 940
rect 54655 910 55285 940
rect 55315 910 56035 940
rect 56065 910 56735 940
rect 56765 910 57035 940
rect 57065 910 57735 940
rect 57765 910 58485 940
rect 58515 910 59145 940
rect 59175 910 59845 940
rect 59875 910 59885 940
rect 59915 910 59925 940
rect 59955 910 59960 940
rect 53840 900 59960 910
rect 53840 870 53845 900
rect 53875 870 53885 900
rect 53915 870 53925 900
rect 53955 870 54625 900
rect 54655 870 55285 900
rect 55315 870 56035 900
rect 56065 870 56735 900
rect 56765 870 57035 900
rect 57065 870 57735 900
rect 57765 870 58485 900
rect 58515 870 59145 900
rect 59175 870 59845 900
rect 59875 870 59885 900
rect 59915 870 59925 900
rect 59955 870 59960 900
rect 53840 860 59960 870
rect 53840 830 53845 860
rect 53875 830 53885 860
rect 53915 830 53925 860
rect 53955 830 54625 860
rect 54655 830 55285 860
rect 55315 830 56035 860
rect 56065 830 56735 860
rect 56765 830 57035 860
rect 57065 830 57735 860
rect 57765 830 58485 860
rect 58515 830 59145 860
rect 59175 830 59845 860
rect 59875 830 59885 860
rect 59915 830 59925 860
rect 59955 830 59960 860
rect 53840 825 59960 830
rect 54255 805 54295 810
rect 54255 775 54260 805
rect 54290 800 54295 805
rect 55940 805 55980 810
rect 55940 800 55945 805
rect 54290 780 55945 800
rect 54290 775 54295 780
rect 54255 770 54295 775
rect 55940 775 55945 780
rect 55975 775 55980 805
rect 55940 770 55980 775
rect 57820 805 57860 810
rect 57820 775 57825 805
rect 57855 800 57860 805
rect 59505 805 59545 810
rect 59505 800 59510 805
rect 57855 780 59510 800
rect 57855 775 57860 780
rect 57820 770 57860 775
rect 59505 775 59510 780
rect 59540 775 59545 805
rect 59505 770 59545 775
rect 54320 525 54360 530
rect 54320 495 54325 525
rect 54355 520 54360 525
rect 55000 525 55040 530
rect 55000 520 55005 525
rect 54355 500 55005 520
rect 54355 495 54360 500
rect 54320 490 54360 495
rect 55000 495 55005 500
rect 55035 520 55040 525
rect 58760 525 58800 530
rect 58760 520 58765 525
rect 55035 500 58765 520
rect 55035 495 55040 500
rect 55000 490 55040 495
rect 58760 495 58765 500
rect 58795 520 58800 525
rect 59440 525 59480 530
rect 59440 520 59445 525
rect 58795 500 59445 520
rect 58795 495 58800 500
rect 58760 490 58800 495
rect 59440 495 59445 500
rect 59475 495 59480 525
rect 59440 490 59480 495
rect 56440 480 57470 485
rect 53990 470 55190 475
rect 53990 440 53995 470
rect 54025 440 54035 470
rect 54065 440 54080 470
rect 54110 440 54120 470
rect 54150 440 54165 470
rect 54195 440 54205 470
rect 54235 440 54390 470
rect 54420 440 54755 470
rect 54785 440 54795 470
rect 54825 440 54835 470
rect 54865 440 54875 470
rect 54905 440 54915 470
rect 54945 440 54955 470
rect 54985 440 54995 470
rect 55025 440 55035 470
rect 55065 440 55075 470
rect 55105 440 55115 470
rect 55145 440 55155 470
rect 55185 440 55190 470
rect 56440 450 56445 480
rect 56475 450 56555 480
rect 56585 450 56665 480
rect 56695 450 56775 480
rect 56805 450 56885 480
rect 56915 450 56995 480
rect 57025 450 57105 480
rect 57135 450 57215 480
rect 57245 450 57325 480
rect 57355 450 57435 480
rect 57465 450 57470 480
rect 56440 445 57470 450
rect 58610 470 59810 475
rect 53990 430 55190 440
rect 53990 400 53995 430
rect 54025 400 54035 430
rect 54065 400 54080 430
rect 54110 400 54120 430
rect 54150 400 54165 430
rect 54195 400 54205 430
rect 54235 400 54390 430
rect 54420 400 54755 430
rect 54785 400 54795 430
rect 54825 400 54835 430
rect 54865 400 54875 430
rect 54905 400 54915 430
rect 54945 400 54955 430
rect 54985 400 54995 430
rect 55025 400 55035 430
rect 55065 400 55075 430
rect 55105 400 55115 430
rect 55145 400 55155 430
rect 55185 400 55190 430
rect 53990 390 55190 400
rect 53990 360 53995 390
rect 54025 360 54035 390
rect 54065 360 54080 390
rect 54110 360 54120 390
rect 54150 360 54165 390
rect 54195 360 54205 390
rect 54235 360 54390 390
rect 54420 360 54755 390
rect 54785 360 54795 390
rect 54825 360 54835 390
rect 54865 360 54875 390
rect 54905 360 54915 390
rect 54945 360 54955 390
rect 54985 360 54995 390
rect 55025 360 55035 390
rect 55065 360 55075 390
rect 55105 360 55115 390
rect 55145 360 55155 390
rect 55185 360 55190 390
rect 53990 355 55190 360
rect 58610 440 58615 470
rect 58645 440 58655 470
rect 58685 440 58695 470
rect 58725 440 58735 470
rect 58765 440 58775 470
rect 58805 440 58815 470
rect 58845 440 58855 470
rect 58885 440 58895 470
rect 58925 440 58935 470
rect 58965 440 58975 470
rect 59005 440 59015 470
rect 59045 440 59380 470
rect 59410 440 59565 470
rect 59595 440 59605 470
rect 59635 440 59650 470
rect 59680 440 59690 470
rect 59720 440 59735 470
rect 59765 440 59775 470
rect 59805 440 59810 470
rect 58610 430 59810 440
rect 58610 400 58615 430
rect 58645 400 58655 430
rect 58685 400 58695 430
rect 58725 400 58735 430
rect 58765 400 58775 430
rect 58805 400 58815 430
rect 58845 400 58855 430
rect 58885 400 58895 430
rect 58925 400 58935 430
rect 58965 400 58975 430
rect 59005 400 59015 430
rect 59045 400 59380 430
rect 59410 400 59565 430
rect 59595 400 59605 430
rect 59635 400 59650 430
rect 59680 400 59690 430
rect 59720 400 59735 430
rect 59765 400 59775 430
rect 59805 400 59810 430
rect 58610 390 59810 400
rect 58610 360 58615 390
rect 58645 360 58655 390
rect 58685 360 58695 390
rect 58725 360 58735 390
rect 58765 360 58775 390
rect 58805 360 58815 390
rect 58845 360 58855 390
rect 58885 360 58895 390
rect 58925 360 58935 390
rect 58965 360 58975 390
rect 59005 360 59015 390
rect 59045 360 59380 390
rect 59410 360 59565 390
rect 59595 360 59605 390
rect 59635 360 59650 390
rect 59680 360 59690 390
rect 59720 360 59735 390
rect 59765 360 59775 390
rect 59805 360 59810 390
rect 58610 355 59810 360
rect 54325 335 54360 340
rect 54325 295 54360 300
rect 54385 335 54420 340
rect 54385 295 54420 300
rect 59380 335 59415 340
rect 59380 295 59415 300
rect 59440 335 59475 340
rect 59440 295 59475 300
rect 56220 150 56260 155
rect 56220 120 56225 150
rect 56255 145 56260 150
rect 56275 150 56315 155
rect 56275 145 56280 150
rect 56255 125 56280 145
rect 56255 120 56260 125
rect 56220 115 56260 120
rect 56275 120 56280 125
rect 56310 145 56315 150
rect 56385 150 56425 155
rect 56385 145 56390 150
rect 56310 125 56390 145
rect 56310 120 56315 125
rect 56275 115 56315 120
rect 56385 120 56390 125
rect 56420 145 56425 150
rect 56495 150 56535 155
rect 56495 145 56500 150
rect 56420 125 56500 145
rect 56420 120 56425 125
rect 56385 115 56425 120
rect 56495 120 56500 125
rect 56530 145 56535 150
rect 56605 150 56645 155
rect 56605 145 56610 150
rect 56530 125 56610 145
rect 56530 120 56535 125
rect 56495 115 56535 120
rect 56605 120 56610 125
rect 56640 145 56645 150
rect 56715 150 56755 155
rect 56715 145 56720 150
rect 56640 125 56720 145
rect 56640 120 56645 125
rect 56605 115 56645 120
rect 56715 120 56720 125
rect 56750 145 56755 150
rect 56825 150 56865 155
rect 56825 145 56830 150
rect 56750 125 56830 145
rect 56750 120 56755 125
rect 56715 115 56755 120
rect 56825 120 56830 125
rect 56860 145 56865 150
rect 56935 150 56975 155
rect 56935 145 56940 150
rect 56860 125 56940 145
rect 56860 120 56865 125
rect 56825 115 56865 120
rect 56935 120 56940 125
rect 56970 145 56975 150
rect 57045 150 57085 155
rect 57045 145 57050 150
rect 56970 125 57050 145
rect 56970 120 56975 125
rect 56935 115 56975 120
rect 57045 120 57050 125
rect 57080 145 57085 150
rect 57155 150 57195 155
rect 57155 145 57160 150
rect 57080 125 57160 145
rect 57080 120 57085 125
rect 57045 115 57085 120
rect 57155 120 57160 125
rect 57190 145 57195 150
rect 57265 150 57305 155
rect 57265 145 57270 150
rect 57190 125 57270 145
rect 57190 120 57195 125
rect 57155 115 57195 120
rect 57265 120 57270 125
rect 57300 145 57305 150
rect 57375 150 57415 155
rect 57375 145 57380 150
rect 57300 125 57380 145
rect 57300 120 57305 125
rect 57265 115 57305 120
rect 57375 120 57380 125
rect 57410 145 57415 150
rect 57485 150 57525 155
rect 57485 145 57490 150
rect 57410 125 57490 145
rect 57410 120 57415 125
rect 57375 115 57415 120
rect 57485 120 57490 125
rect 57520 120 57525 150
rect 57485 115 57525 120
rect 56440 95 57470 100
rect 56440 65 56445 95
rect 56475 65 56555 95
rect 56585 65 56665 95
rect 56695 65 56775 95
rect 56805 65 56885 95
rect 56915 65 56995 95
rect 57025 65 57105 95
rect 57135 65 57215 95
rect 57245 65 57325 95
rect 57355 65 57435 95
rect 57465 65 57470 95
rect 56440 60 57470 65
rect 57415 40 57455 45
rect 57415 10 57420 40
rect 57450 35 57455 40
rect 57865 40 57905 45
rect 57865 35 57870 40
rect 57450 15 57870 35
rect 57450 10 57455 15
rect 57415 5 57455 10
rect 57865 10 57870 15
rect 57900 10 57905 40
rect 57865 5 57905 10
rect 55670 -60 58130 -55
rect 55670 -90 55675 -60
rect 55705 -90 55715 -60
rect 55745 -90 55755 -60
rect 55785 -90 56335 -60
rect 56365 -90 58015 -60
rect 58045 -90 58055 -60
rect 58085 -90 58095 -60
rect 58125 -90 58130 -60
rect 55670 -100 58130 -90
rect 55670 -130 55675 -100
rect 55705 -130 55715 -100
rect 55745 -130 55755 -100
rect 55785 -130 56335 -100
rect 56365 -130 58015 -100
rect 58045 -130 58055 -100
rect 58085 -130 58095 -100
rect 58125 -130 58130 -100
rect 55670 -140 58130 -130
rect 55670 -170 55675 -140
rect 55705 -170 55715 -140
rect 55745 -170 55755 -140
rect 55785 -170 56335 -140
rect 56365 -170 58015 -140
rect 58045 -170 58055 -140
rect 58085 -170 58095 -140
rect 58125 -170 58130 -140
rect 55670 -175 58130 -170
rect 56540 -195 56580 -190
rect 56540 -225 56545 -195
rect 56575 -200 56580 -195
rect 56650 -195 56690 -190
rect 56650 -200 56655 -195
rect 56575 -220 56655 -200
rect 56575 -225 56580 -220
rect 56540 -230 56580 -225
rect 56650 -225 56655 -220
rect 56685 -200 56690 -195
rect 56870 -195 56910 -190
rect 56870 -200 56875 -195
rect 56685 -220 56875 -200
rect 56685 -225 56690 -220
rect 56650 -230 56690 -225
rect 56870 -225 56875 -220
rect 56905 -225 56910 -195
rect 56870 -230 56910 -225
rect 55885 -250 55925 -245
rect 55885 -280 55890 -250
rect 55920 -255 55925 -250
rect 56485 -250 57200 -245
rect 56485 -255 56490 -250
rect 55920 -270 56490 -255
rect 55920 -280 55925 -270
rect 55885 -285 55925 -280
rect 56485 -280 56490 -270
rect 56520 -280 56600 -250
rect 56630 -280 56710 -250
rect 56740 -280 56925 -250
rect 56955 -280 57045 -250
rect 57075 -280 57165 -250
rect 57195 -280 57200 -250
rect 56485 -285 57200 -280
rect 54750 -365 55190 -360
rect 54750 -395 54755 -365
rect 54785 -395 54955 -365
rect 54985 -395 55155 -365
rect 55185 -395 55190 -365
rect 54750 -400 55190 -395
rect 58610 -365 59050 -360
rect 58610 -395 58615 -365
rect 58645 -395 58815 -365
rect 58845 -395 59015 -365
rect 59045 -395 59050 -365
rect 58610 -400 59050 -395
rect 56485 -470 57200 -465
rect 56485 -500 56490 -470
rect 56520 -500 56600 -470
rect 56630 -500 56710 -470
rect 56740 -500 56925 -470
rect 56955 -500 57045 -470
rect 57075 -500 57165 -470
rect 57195 -500 57200 -470
rect 56485 -505 57200 -500
rect 56540 -525 56910 -520
rect 56540 -555 56545 -525
rect 56575 -555 56655 -525
rect 56685 -555 56875 -525
rect 56905 -555 56910 -525
rect 56540 -560 56910 -555
rect 52290 -580 61510 -575
rect 52290 -610 52295 -580
rect 52325 -610 52335 -580
rect 52365 -610 52375 -580
rect 52405 -610 52645 -580
rect 52675 -610 52685 -580
rect 52715 -610 52725 -580
rect 52755 -610 52995 -580
rect 53025 -610 53035 -580
rect 53065 -610 53075 -580
rect 53105 -610 53345 -580
rect 53375 -610 53385 -580
rect 53415 -610 53425 -580
rect 53455 -610 53695 -580
rect 53725 -610 53735 -580
rect 53765 -610 53775 -580
rect 53805 -610 53845 -580
rect 53875 -610 53885 -580
rect 53915 -610 53925 -580
rect 53955 -610 54045 -580
rect 54075 -610 54085 -580
rect 54115 -610 54125 -580
rect 54155 -610 54395 -580
rect 54425 -610 54435 -580
rect 54465 -610 54475 -580
rect 54505 -610 54655 -580
rect 54685 -610 54745 -580
rect 54775 -610 54785 -580
rect 54815 -610 54825 -580
rect 54855 -610 55095 -580
rect 55125 -610 55135 -580
rect 55165 -610 55175 -580
rect 55205 -610 55255 -580
rect 55285 -610 55445 -580
rect 55475 -610 55485 -580
rect 55515 -610 55525 -580
rect 55555 -610 55795 -580
rect 55825 -610 55835 -580
rect 55865 -610 55875 -580
rect 55905 -610 56145 -580
rect 56175 -610 56185 -580
rect 56215 -610 56225 -580
rect 56255 -610 56435 -580
rect 56465 -610 56495 -580
rect 56525 -610 56535 -580
rect 56565 -610 56575 -580
rect 56605 -610 56765 -580
rect 56795 -610 56845 -580
rect 56875 -610 56885 -580
rect 56915 -610 56925 -580
rect 56955 -610 57195 -580
rect 57225 -610 57235 -580
rect 57265 -610 57275 -580
rect 57305 -610 57490 -580
rect 57520 -610 57545 -580
rect 57575 -610 57585 -580
rect 57615 -610 57625 -580
rect 57655 -610 57895 -580
rect 57925 -610 57935 -580
rect 57965 -610 57975 -580
rect 58005 -610 58245 -580
rect 58275 -610 58285 -580
rect 58315 -610 58325 -580
rect 58355 -610 58515 -580
rect 58545 -610 58595 -580
rect 58625 -610 58635 -580
rect 58665 -610 58675 -580
rect 58705 -610 58945 -580
rect 58975 -610 58985 -580
rect 59015 -610 59025 -580
rect 59055 -610 59115 -580
rect 59145 -610 59375 -580
rect 59405 -610 59415 -580
rect 59445 -610 59455 -580
rect 59485 -610 59645 -580
rect 59675 -610 59685 -580
rect 59715 -610 59725 -580
rect 59755 -610 59845 -580
rect 59875 -610 59885 -580
rect 59915 -610 59925 -580
rect 59955 -610 59995 -580
rect 60025 -610 60035 -580
rect 60065 -610 60075 -580
rect 60105 -610 60345 -580
rect 60375 -610 60385 -580
rect 60415 -610 60425 -580
rect 60455 -610 60695 -580
rect 60725 -610 60735 -580
rect 60765 -610 60775 -580
rect 60805 -610 61045 -580
rect 61075 -610 61085 -580
rect 61115 -610 61125 -580
rect 61155 -610 61395 -580
rect 61425 -610 61435 -580
rect 61465 -610 61475 -580
rect 61505 -610 61510 -580
rect 52290 -620 61510 -610
rect 52290 -650 52295 -620
rect 52325 -650 52335 -620
rect 52365 -650 52375 -620
rect 52405 -650 52645 -620
rect 52675 -650 52685 -620
rect 52715 -650 52725 -620
rect 52755 -650 52995 -620
rect 53025 -650 53035 -620
rect 53065 -650 53075 -620
rect 53105 -650 53345 -620
rect 53375 -650 53385 -620
rect 53415 -650 53425 -620
rect 53455 -650 53695 -620
rect 53725 -650 53735 -620
rect 53765 -650 53775 -620
rect 53805 -650 53845 -620
rect 53875 -650 53885 -620
rect 53915 -650 53925 -620
rect 53955 -650 54045 -620
rect 54075 -650 54085 -620
rect 54115 -650 54125 -620
rect 54155 -650 54395 -620
rect 54425 -650 54435 -620
rect 54465 -650 54475 -620
rect 54505 -650 54655 -620
rect 54685 -650 54745 -620
rect 54775 -650 54785 -620
rect 54815 -650 54825 -620
rect 54855 -650 55095 -620
rect 55125 -650 55135 -620
rect 55165 -650 55175 -620
rect 55205 -650 55255 -620
rect 55285 -650 55445 -620
rect 55475 -650 55485 -620
rect 55515 -650 55525 -620
rect 55555 -650 55795 -620
rect 55825 -650 55835 -620
rect 55865 -650 55875 -620
rect 55905 -650 56145 -620
rect 56175 -650 56185 -620
rect 56215 -650 56225 -620
rect 56255 -650 56435 -620
rect 56465 -650 56495 -620
rect 56525 -650 56535 -620
rect 56565 -650 56575 -620
rect 56605 -650 56765 -620
rect 56795 -650 56845 -620
rect 56875 -650 56885 -620
rect 56915 -650 56925 -620
rect 56955 -650 57195 -620
rect 57225 -650 57235 -620
rect 57265 -650 57275 -620
rect 57305 -650 57490 -620
rect 57520 -650 57545 -620
rect 57575 -650 57585 -620
rect 57615 -650 57625 -620
rect 57655 -650 57895 -620
rect 57925 -650 57935 -620
rect 57965 -650 57975 -620
rect 58005 -650 58245 -620
rect 58275 -650 58285 -620
rect 58315 -650 58325 -620
rect 58355 -650 58515 -620
rect 58545 -650 58595 -620
rect 58625 -650 58635 -620
rect 58665 -650 58675 -620
rect 58705 -650 58945 -620
rect 58975 -650 58985 -620
rect 59015 -650 59025 -620
rect 59055 -650 59115 -620
rect 59145 -650 59375 -620
rect 59405 -650 59415 -620
rect 59445 -650 59455 -620
rect 59485 -650 59645 -620
rect 59675 -650 59685 -620
rect 59715 -650 59725 -620
rect 59755 -650 59845 -620
rect 59875 -650 59885 -620
rect 59915 -650 59925 -620
rect 59955 -650 59995 -620
rect 60025 -650 60035 -620
rect 60065 -650 60075 -620
rect 60105 -650 60345 -620
rect 60375 -650 60385 -620
rect 60415 -650 60425 -620
rect 60455 -650 60695 -620
rect 60725 -650 60735 -620
rect 60765 -650 60775 -620
rect 60805 -650 61045 -620
rect 61075 -650 61085 -620
rect 61115 -650 61125 -620
rect 61155 -650 61395 -620
rect 61425 -650 61435 -620
rect 61465 -650 61475 -620
rect 61505 -650 61510 -620
rect 52290 -660 61510 -650
rect 52290 -690 52295 -660
rect 52325 -690 52335 -660
rect 52365 -690 52375 -660
rect 52405 -690 52645 -660
rect 52675 -690 52685 -660
rect 52715 -690 52725 -660
rect 52755 -690 52995 -660
rect 53025 -690 53035 -660
rect 53065 -690 53075 -660
rect 53105 -690 53345 -660
rect 53375 -690 53385 -660
rect 53415 -690 53425 -660
rect 53455 -690 53695 -660
rect 53725 -690 53735 -660
rect 53765 -690 53775 -660
rect 53805 -690 53845 -660
rect 53875 -690 53885 -660
rect 53915 -690 53925 -660
rect 53955 -690 54045 -660
rect 54075 -690 54085 -660
rect 54115 -690 54125 -660
rect 54155 -690 54395 -660
rect 54425 -690 54435 -660
rect 54465 -690 54475 -660
rect 54505 -690 54655 -660
rect 54685 -690 54745 -660
rect 54775 -690 54785 -660
rect 54815 -690 54825 -660
rect 54855 -690 55095 -660
rect 55125 -690 55135 -660
rect 55165 -690 55175 -660
rect 55205 -690 55255 -660
rect 55285 -690 55445 -660
rect 55475 -690 55485 -660
rect 55515 -690 55525 -660
rect 55555 -690 55795 -660
rect 55825 -690 55835 -660
rect 55865 -690 55875 -660
rect 55905 -690 56145 -660
rect 56175 -690 56185 -660
rect 56215 -690 56225 -660
rect 56255 -690 56435 -660
rect 56465 -690 56495 -660
rect 56525 -690 56535 -660
rect 56565 -690 56575 -660
rect 56605 -690 56765 -660
rect 56795 -690 56845 -660
rect 56875 -690 56885 -660
rect 56915 -690 56925 -660
rect 56955 -690 57195 -660
rect 57225 -690 57235 -660
rect 57265 -690 57275 -660
rect 57305 -690 57490 -660
rect 57520 -690 57545 -660
rect 57575 -690 57585 -660
rect 57615 -690 57625 -660
rect 57655 -690 57895 -660
rect 57925 -690 57935 -660
rect 57965 -690 57975 -660
rect 58005 -690 58245 -660
rect 58275 -690 58285 -660
rect 58315 -690 58325 -660
rect 58355 -690 58515 -660
rect 58545 -690 58595 -660
rect 58625 -690 58635 -660
rect 58665 -690 58675 -660
rect 58705 -690 58945 -660
rect 58975 -690 58985 -660
rect 59015 -690 59025 -660
rect 59055 -690 59115 -660
rect 59145 -690 59375 -660
rect 59405 -690 59415 -660
rect 59445 -690 59455 -660
rect 59485 -690 59645 -660
rect 59675 -690 59685 -660
rect 59715 -690 59725 -660
rect 59755 -690 59845 -660
rect 59875 -690 59885 -660
rect 59915 -690 59925 -660
rect 59955 -690 59995 -660
rect 60025 -690 60035 -660
rect 60065 -690 60075 -660
rect 60105 -690 60345 -660
rect 60375 -690 60385 -660
rect 60415 -690 60425 -660
rect 60455 -690 60695 -660
rect 60725 -690 60735 -660
rect 60765 -690 60775 -660
rect 60805 -690 61045 -660
rect 61075 -690 61085 -660
rect 61115 -690 61125 -660
rect 61155 -690 61395 -660
rect 61425 -690 61435 -660
rect 61465 -690 61475 -660
rect 61505 -690 61510 -660
rect 52290 -695 61510 -690
<< via2 >>
rect 54260 3345 54290 3375
rect 59510 3345 59540 3375
rect 54000 1680 54030 1710
rect 54050 1680 54080 1710
rect 54100 1680 54130 1710
rect 54150 1680 54180 1710
rect 54200 1680 54230 1710
rect 54000 1630 54030 1660
rect 54050 1630 54080 1660
rect 54100 1630 54130 1660
rect 54150 1630 54180 1660
rect 54200 1630 54230 1660
rect 59570 1680 59600 1710
rect 59620 1680 59650 1710
rect 59670 1680 59700 1710
rect 59720 1680 59750 1710
rect 59770 1680 59800 1710
rect 54000 1580 54030 1610
rect 54050 1580 54080 1610
rect 54100 1580 54130 1610
rect 54150 1580 54180 1610
rect 54200 1580 54230 1610
rect 59570 1630 59600 1660
rect 59620 1630 59650 1660
rect 59670 1630 59700 1660
rect 59720 1630 59750 1660
rect 59770 1630 59800 1660
rect 59570 1580 59600 1610
rect 59620 1580 59650 1610
rect 59670 1580 59700 1610
rect 59720 1580 59750 1610
rect 59770 1580 59800 1610
<< metal3 >>
rect 52060 5520 52290 5605
rect 52410 5520 52640 5605
rect 52760 5520 52990 5605
rect 53110 5520 53340 5605
rect 53460 5520 53690 5605
rect 53810 5520 54040 5605
rect 54160 5520 54390 5605
rect 54510 5520 54740 5605
rect 54860 5520 55090 5605
rect 55210 5520 55440 5605
rect 55560 5520 55790 5605
rect 55910 5520 56140 5605
rect 56260 5520 56490 5605
rect 56610 5520 56840 5605
rect 52060 5470 56840 5520
rect 52060 5375 52290 5470
rect 52410 5375 52640 5470
rect 52760 5375 52990 5470
rect 53110 5375 53340 5470
rect 53460 5375 53690 5470
rect 53810 5375 54040 5470
rect 54160 5375 54390 5470
rect 54510 5375 54740 5470
rect 54860 5375 55090 5470
rect 55210 5375 55440 5470
rect 55560 5375 55790 5470
rect 55910 5375 56140 5470
rect 56260 5375 56490 5470
rect 56610 5375 56840 5470
rect 56960 5520 57190 5605
rect 57310 5520 57540 5605
rect 57660 5520 57890 5605
rect 58010 5520 58240 5605
rect 58360 5520 58590 5605
rect 58710 5520 58940 5605
rect 59060 5520 59290 5605
rect 59410 5520 59640 5605
rect 59760 5520 59990 5605
rect 60110 5520 60340 5605
rect 60460 5520 60690 5605
rect 60810 5520 61040 5605
rect 61160 5520 61390 5605
rect 61510 5520 61740 5605
rect 56960 5470 61740 5520
rect 56960 5375 57190 5470
rect 57310 5375 57540 5470
rect 57660 5375 57890 5470
rect 58010 5375 58240 5470
rect 58360 5375 58590 5470
rect 58710 5375 58940 5470
rect 59060 5375 59290 5470
rect 59410 5375 59640 5470
rect 59760 5375 59990 5470
rect 60110 5375 60340 5470
rect 60460 5375 60690 5470
rect 60810 5375 61040 5470
rect 61160 5375 61390 5470
rect 61510 5375 61740 5470
rect 52850 5255 52900 5375
rect 53900 5255 53950 5375
rect 54250 5255 54300 5375
rect 54600 5255 54650 5375
rect 54950 5255 55000 5375
rect 55300 5255 55350 5375
rect 55650 5255 55700 5375
rect 58100 5255 58150 5375
rect 58450 5255 58500 5375
rect 58800 5255 58850 5375
rect 59150 5255 59200 5375
rect 59500 5255 59550 5375
rect 59850 5255 59900 5375
rect 60900 5255 60950 5375
rect 52060 5170 52290 5255
rect 52410 5170 52640 5255
rect 52760 5170 52990 5255
rect 53110 5170 53340 5255
rect 53460 5170 53690 5255
rect 52060 5120 53690 5170
rect 52060 5025 52290 5120
rect 52410 5025 52640 5120
rect 52760 5025 52990 5120
rect 53110 5025 53340 5120
rect 53460 5025 53690 5120
rect 53810 5025 54040 5255
rect 54160 5025 54390 5255
rect 54510 5025 54740 5255
rect 54860 5025 55090 5255
rect 55210 5025 55440 5255
rect 55560 5025 55790 5255
rect 58010 5025 58240 5255
rect 58360 5025 58590 5255
rect 58710 5025 58940 5255
rect 59060 5025 59290 5255
rect 59410 5025 59640 5255
rect 59760 5025 59990 5255
rect 60110 5170 60340 5255
rect 60460 5170 60690 5255
rect 60810 5170 61040 5255
rect 61160 5170 61390 5255
rect 61510 5170 61740 5255
rect 60110 5120 61740 5170
rect 60110 5025 60340 5120
rect 60460 5025 60690 5120
rect 60810 5025 61040 5120
rect 61160 5025 61390 5120
rect 61510 5025 61740 5120
rect 52850 4905 52900 5025
rect 53900 4905 53950 5025
rect 54250 4905 54300 5025
rect 54600 4905 54650 5025
rect 54950 4905 55000 5025
rect 55300 4905 55350 5025
rect 58450 4905 58500 5025
rect 58800 4905 58850 5025
rect 59150 4905 59200 5025
rect 59500 4905 59550 5025
rect 59850 4905 59900 5025
rect 60900 4905 60950 5025
rect 52060 4820 52290 4905
rect 52410 4820 52640 4905
rect 52760 4820 52990 4905
rect 53110 4820 53340 4905
rect 53460 4820 53690 4905
rect 52060 4770 53690 4820
rect 52060 4675 52290 4770
rect 52410 4675 52640 4770
rect 52760 4675 52990 4770
rect 53110 4675 53340 4770
rect 53460 4675 53690 4770
rect 53810 4675 54040 4905
rect 54160 4675 54390 4905
rect 54510 4675 54740 4905
rect 54860 4675 55090 4905
rect 55210 4675 55440 4905
rect 58360 4675 58590 4905
rect 58710 4675 58940 4905
rect 59060 4675 59290 4905
rect 59410 4675 59640 4905
rect 59760 4675 59990 4905
rect 60110 4820 60340 4905
rect 60460 4820 60690 4905
rect 60810 4820 61040 4905
rect 61160 4820 61390 4905
rect 61510 4820 61740 4905
rect 60110 4770 61740 4820
rect 60110 4675 60340 4770
rect 60460 4675 60690 4770
rect 60810 4675 61040 4770
rect 61160 4675 61390 4770
rect 61510 4675 61740 4770
rect 52850 4555 52900 4675
rect 52060 4470 52290 4555
rect 52410 4470 52640 4555
rect 52760 4470 52990 4555
rect 53110 4470 53340 4555
rect 53460 4470 53690 4555
rect 52060 4420 53690 4470
rect 52060 4325 52290 4420
rect 52410 4325 52640 4420
rect 52760 4325 52990 4420
rect 53110 4325 53340 4420
rect 53460 4325 53690 4420
rect 52850 4205 52900 4325
rect 52060 4120 52290 4205
rect 52410 4120 52640 4205
rect 52760 4120 52990 4205
rect 53110 4120 53340 4205
rect 53460 4120 53690 4205
rect 52060 4070 53690 4120
rect 52060 3975 52290 4070
rect 52410 3975 52640 4070
rect 52760 3975 52990 4070
rect 53110 3975 53340 4070
rect 53460 3975 53690 4070
rect 52850 3855 52900 3975
rect 52060 3770 52290 3855
rect 52410 3770 52640 3855
rect 52760 3770 52990 3855
rect 53110 3770 53340 3855
rect 53460 3770 53690 3855
rect 52060 3720 53690 3770
rect 52060 3625 52290 3720
rect 52410 3625 52640 3720
rect 52760 3625 52990 3720
rect 53110 3625 53340 3720
rect 53460 3625 53690 3720
rect 52850 3505 52900 3625
rect 52060 3420 52290 3505
rect 52410 3420 52640 3505
rect 52760 3420 52990 3505
rect 53110 3420 53340 3505
rect 53460 3420 53690 3505
rect 52060 3370 53690 3420
rect 52060 3275 52290 3370
rect 52410 3275 52640 3370
rect 52760 3275 52990 3370
rect 53110 3275 53340 3370
rect 53460 3275 53690 3370
rect 54255 3375 54295 4675
rect 54255 3345 54260 3375
rect 54290 3345 54295 3375
rect 54255 3340 54295 3345
rect 59505 3375 59545 4675
rect 60900 4555 60950 4675
rect 60110 4470 60340 4555
rect 60460 4470 60690 4555
rect 60810 4470 61040 4555
rect 61160 4470 61390 4555
rect 61510 4470 61740 4555
rect 60110 4420 61740 4470
rect 60110 4325 60340 4420
rect 60460 4325 60690 4420
rect 60810 4325 61040 4420
rect 61160 4325 61390 4420
rect 61510 4325 61740 4420
rect 60900 4205 60950 4325
rect 60110 4120 60340 4205
rect 60460 4120 60690 4205
rect 60810 4120 61040 4205
rect 61160 4120 61390 4205
rect 61510 4120 61740 4205
rect 60110 4070 61740 4120
rect 60110 3975 60340 4070
rect 60460 3975 60690 4070
rect 60810 3975 61040 4070
rect 61160 3975 61390 4070
rect 61510 3975 61740 4070
rect 60900 3855 60950 3975
rect 60110 3770 60340 3855
rect 60460 3770 60690 3855
rect 60810 3770 61040 3855
rect 61160 3770 61390 3855
rect 61510 3770 61740 3855
rect 60110 3720 61740 3770
rect 60110 3625 60340 3720
rect 60460 3625 60690 3720
rect 60810 3625 61040 3720
rect 61160 3625 61390 3720
rect 61510 3625 61740 3720
rect 60900 3505 60950 3625
rect 59505 3345 59510 3375
rect 59540 3345 59545 3375
rect 59505 3340 59545 3345
rect 60110 3420 60340 3505
rect 60460 3420 60690 3505
rect 60810 3420 61040 3505
rect 61160 3420 61390 3505
rect 61510 3420 61740 3505
rect 60110 3370 61740 3420
rect 60110 3275 60340 3370
rect 60460 3275 60690 3370
rect 60810 3275 61040 3370
rect 61160 3275 61390 3370
rect 61510 3275 61740 3370
rect 52850 3155 52900 3275
rect 60900 3155 60950 3275
rect 52060 3070 52290 3155
rect 52410 3070 52640 3155
rect 52760 3070 52990 3155
rect 53110 3070 53340 3155
rect 53460 3070 53690 3155
rect 52060 3020 53690 3070
rect 52060 2925 52290 3020
rect 52410 2925 52640 3020
rect 52760 2925 52990 3020
rect 53110 2925 53340 3020
rect 53460 2925 53690 3020
rect 60110 3070 60340 3155
rect 60460 3070 60690 3155
rect 60810 3070 61040 3155
rect 61160 3070 61390 3155
rect 61510 3070 61740 3155
rect 60110 3020 61740 3070
rect 60110 2925 60340 3020
rect 60460 2925 60690 3020
rect 60810 2925 61040 3020
rect 61160 2925 61390 3020
rect 61510 2925 61740 3020
rect 52850 2805 52900 2925
rect 60900 2805 60950 2925
rect 52060 2720 52290 2805
rect 52410 2720 52640 2805
rect 52760 2720 52990 2805
rect 53110 2720 53340 2805
rect 53460 2720 53690 2805
rect 52060 2670 53690 2720
rect 52060 2575 52290 2670
rect 52410 2575 52640 2670
rect 52760 2575 52990 2670
rect 53110 2575 53340 2670
rect 53460 2575 53690 2670
rect 60110 2720 60340 2805
rect 60460 2720 60690 2805
rect 60810 2720 61040 2805
rect 61160 2720 61390 2805
rect 61510 2720 61740 2805
rect 60110 2670 61740 2720
rect 60110 2575 60340 2670
rect 60460 2575 60690 2670
rect 60810 2575 61040 2670
rect 61160 2575 61390 2670
rect 61510 2575 61740 2670
rect 52850 2455 52900 2575
rect 60900 2455 60950 2575
rect 52060 2370 52290 2455
rect 52410 2370 52640 2455
rect 52760 2370 52990 2455
rect 53110 2370 53340 2455
rect 53460 2370 53690 2455
rect 52060 2320 53690 2370
rect 52060 2225 52290 2320
rect 52410 2225 52640 2320
rect 52760 2225 52990 2320
rect 53110 2225 53340 2320
rect 53460 2225 53690 2320
rect 60110 2370 60340 2455
rect 60460 2370 60690 2455
rect 60810 2370 61040 2455
rect 61160 2370 61390 2455
rect 61510 2370 61740 2455
rect 60110 2320 61740 2370
rect 60110 2225 60340 2320
rect 60460 2225 60690 2320
rect 60810 2225 61040 2320
rect 61160 2225 61390 2320
rect 61510 2225 61740 2320
rect 52850 2105 52900 2225
rect 60900 2105 60950 2225
rect 52060 2020 52290 2105
rect 52410 2020 52640 2105
rect 52760 2020 52990 2105
rect 53110 2020 53340 2105
rect 53460 2020 53690 2105
rect 52060 1970 53690 2020
rect 52060 1875 52290 1970
rect 52410 1875 52640 1970
rect 52760 1875 52990 1970
rect 53110 1875 53340 1970
rect 53460 1875 53690 1970
rect 60110 2020 60340 2105
rect 60460 2020 60690 2105
rect 60810 2020 61040 2105
rect 61160 2020 61390 2105
rect 61510 2020 61740 2105
rect 60110 1970 61740 2020
rect 60110 1875 60340 1970
rect 60460 1875 60690 1970
rect 60810 1875 61040 1970
rect 61160 1875 61390 1970
rect 61510 1875 61740 1970
rect 52850 1755 52900 1875
rect 60900 1755 60950 1875
rect 52060 1670 52290 1755
rect 52410 1670 52640 1755
rect 52760 1670 52990 1755
rect 53110 1670 53340 1755
rect 53460 1670 53690 1755
rect 52060 1620 53690 1670
rect 52060 1525 52290 1620
rect 52410 1525 52640 1620
rect 52760 1525 52990 1620
rect 53110 1525 53340 1620
rect 53460 1525 53690 1620
rect 53990 1715 54240 1720
rect 53990 1675 53995 1715
rect 54035 1675 54045 1715
rect 54085 1675 54095 1715
rect 54135 1675 54145 1715
rect 54185 1675 54195 1715
rect 54235 1675 54240 1715
rect 53990 1665 54240 1675
rect 53990 1625 53995 1665
rect 54035 1625 54045 1665
rect 54085 1625 54095 1665
rect 54135 1625 54145 1665
rect 54185 1625 54195 1665
rect 54235 1625 54240 1665
rect 53990 1615 54240 1625
rect 53990 1575 53995 1615
rect 54035 1575 54045 1615
rect 54085 1575 54095 1615
rect 54135 1575 54145 1615
rect 54185 1575 54195 1615
rect 54235 1575 54240 1615
rect 53990 1570 54240 1575
rect 59560 1715 59810 1720
rect 59560 1675 59565 1715
rect 59605 1675 59615 1715
rect 59655 1675 59665 1715
rect 59705 1675 59715 1715
rect 59755 1675 59765 1715
rect 59805 1675 59810 1715
rect 59560 1665 59810 1675
rect 59560 1625 59565 1665
rect 59605 1625 59615 1665
rect 59655 1625 59665 1665
rect 59705 1625 59715 1665
rect 59755 1625 59765 1665
rect 59805 1625 59810 1665
rect 59560 1615 59810 1625
rect 59560 1575 59565 1615
rect 59605 1575 59615 1615
rect 59655 1575 59665 1615
rect 59705 1575 59715 1615
rect 59755 1575 59765 1615
rect 59805 1575 59810 1615
rect 59560 1570 59810 1575
rect 60110 1670 60340 1755
rect 60460 1670 60690 1755
rect 60810 1670 61040 1755
rect 61160 1670 61390 1755
rect 61510 1670 61740 1755
rect 60110 1620 61740 1670
rect 60110 1525 60340 1620
rect 60460 1525 60690 1620
rect 60810 1525 61040 1620
rect 61160 1525 61390 1620
rect 61510 1525 61740 1620
rect 52850 1405 52900 1525
rect 60900 1405 60950 1525
rect 52060 1320 52290 1405
rect 52410 1320 52640 1405
rect 52760 1320 52990 1405
rect 53110 1320 53340 1405
rect 53460 1320 53690 1405
rect 52060 1270 53690 1320
rect 52060 1175 52290 1270
rect 52410 1175 52640 1270
rect 52760 1175 52990 1270
rect 53110 1175 53340 1270
rect 53460 1175 53690 1270
rect 60110 1320 60340 1405
rect 60460 1320 60690 1405
rect 60810 1320 61040 1405
rect 61160 1320 61390 1405
rect 61510 1320 61740 1405
rect 60110 1270 61740 1320
rect 60110 1175 60340 1270
rect 60460 1175 60690 1270
rect 60810 1175 61040 1270
rect 61160 1175 61390 1270
rect 61510 1175 61740 1270
rect 52850 1055 52900 1175
rect 60900 1055 60950 1175
rect 52060 970 52290 1055
rect 52410 970 52640 1055
rect 52760 970 52990 1055
rect 53110 970 53340 1055
rect 53460 970 53690 1055
rect 52060 920 53690 970
rect 52060 825 52290 920
rect 52410 825 52640 920
rect 52760 825 52990 920
rect 53110 825 53340 920
rect 53460 825 53690 920
rect 60110 970 60340 1055
rect 60460 970 60690 1055
rect 60810 970 61040 1055
rect 61160 970 61390 1055
rect 61510 970 61740 1055
rect 60110 920 61740 970
rect 60110 825 60340 920
rect 60460 825 60690 920
rect 60810 825 61040 920
rect 61160 825 61390 920
rect 61510 825 61740 920
rect 52850 705 52900 825
rect 60900 705 60950 825
rect 52060 620 52290 705
rect 52410 620 52640 705
rect 52760 620 52990 705
rect 53110 620 53340 705
rect 53460 620 53690 705
rect 52060 570 53690 620
rect 52060 475 52290 570
rect 52410 475 52640 570
rect 52760 475 52990 570
rect 53110 475 53340 570
rect 53460 475 53690 570
rect 60110 620 60340 705
rect 60460 620 60690 705
rect 60810 620 61040 705
rect 61160 620 61390 705
rect 61510 620 61740 705
rect 60110 570 61740 620
rect 60110 475 60340 570
rect 60460 475 60690 570
rect 60810 475 61040 570
rect 61160 475 61390 570
rect 61510 475 61740 570
rect 52850 355 52900 475
rect 60900 355 60950 475
rect 52060 270 52290 355
rect 52410 270 52640 355
rect 52760 270 52990 355
rect 53110 270 53340 355
rect 53460 270 53690 355
rect 52060 220 53690 270
rect 52060 125 52290 220
rect 52410 125 52640 220
rect 52760 125 52990 220
rect 53110 125 53340 220
rect 53460 125 53690 220
rect 60110 270 60340 355
rect 60460 270 60690 355
rect 60810 270 61040 355
rect 61160 270 61390 355
rect 61510 270 61740 355
rect 60110 220 61740 270
rect 60110 125 60340 220
rect 60460 125 60690 220
rect 60810 125 61040 220
rect 61160 125 61390 220
rect 61510 125 61740 220
rect 52850 5 52900 125
rect 60900 5 60950 125
rect 52060 -80 52290 5
rect 52410 -80 52640 5
rect 52760 -80 52990 5
rect 53110 -80 53340 5
rect 53460 -80 53690 5
rect 52060 -130 53690 -80
rect 52060 -225 52290 -130
rect 52410 -225 52640 -130
rect 52760 -225 52990 -130
rect 53110 -225 53340 -130
rect 53460 -225 53690 -130
rect 60110 -80 60340 5
rect 60460 -80 60690 5
rect 60810 -80 61040 5
rect 61160 -80 61390 5
rect 61510 -80 61740 5
rect 60110 -130 61740 -80
rect 60110 -225 60340 -130
rect 60460 -225 60690 -130
rect 60810 -225 61040 -130
rect 61160 -225 61390 -130
rect 61510 -225 61740 -130
rect 52850 -345 52900 -225
rect 60900 -345 60950 -225
rect 52060 -430 52290 -345
rect 52410 -430 52640 -345
rect 52760 -430 52990 -345
rect 53110 -430 53340 -345
rect 53460 -430 53690 -345
rect 52060 -480 53690 -430
rect 52060 -575 52290 -480
rect 52410 -575 52640 -480
rect 52760 -575 52990 -480
rect 53110 -575 53340 -480
rect 53460 -575 53690 -480
rect 60110 -430 60340 -345
rect 60460 -430 60690 -345
rect 60810 -430 61040 -345
rect 61160 -430 61390 -345
rect 61510 -430 61740 -345
rect 60110 -480 61740 -430
rect 60110 -575 60340 -480
rect 60460 -575 60690 -480
rect 60810 -575 61040 -480
rect 61160 -575 61390 -480
rect 61510 -575 61740 -480
rect 52850 -695 52900 -575
rect 60900 -695 60950 -575
rect 52060 -780 52290 -695
rect 52410 -780 52640 -695
rect 52760 -780 52990 -695
rect 53110 -780 53340 -695
rect 53460 -780 53690 -695
rect 53810 -780 54040 -695
rect 54160 -780 54390 -695
rect 54510 -780 54740 -695
rect 54860 -780 55090 -695
rect 55210 -780 55440 -695
rect 55560 -780 55790 -695
rect 55910 -780 56140 -695
rect 56260 -780 56490 -695
rect 56610 -780 56840 -695
rect 52060 -830 56840 -780
rect 52060 -925 52290 -830
rect 52410 -925 52640 -830
rect 52760 -925 52990 -830
rect 53110 -925 53340 -830
rect 53460 -925 53690 -830
rect 53810 -925 54040 -830
rect 54160 -925 54390 -830
rect 54510 -925 54740 -830
rect 54860 -925 55090 -830
rect 55210 -925 55440 -830
rect 55560 -925 55790 -830
rect 55910 -925 56140 -830
rect 56260 -925 56490 -830
rect 56610 -925 56840 -830
rect 56960 -780 57190 -695
rect 57310 -780 57540 -695
rect 57660 -780 57890 -695
rect 58010 -780 58240 -695
rect 58360 -780 58590 -695
rect 58710 -780 58940 -695
rect 59060 -780 59290 -695
rect 59410 -780 59640 -695
rect 59760 -780 59990 -695
rect 60110 -780 60340 -695
rect 60460 -780 60690 -695
rect 60810 -780 61040 -695
rect 61160 -780 61390 -695
rect 61510 -780 61740 -695
rect 56960 -830 61740 -780
rect 56960 -925 57190 -830
rect 57310 -925 57540 -830
rect 57660 -925 57890 -830
rect 58010 -925 58240 -830
rect 58360 -925 58590 -830
rect 58710 -925 58940 -830
rect 59060 -925 59290 -830
rect 59410 -925 59640 -830
rect 59760 -925 59990 -830
rect 60110 -925 60340 -830
rect 60460 -925 60690 -830
rect 60810 -925 61040 -830
rect 61160 -925 61390 -830
rect 61510 -925 61740 -830
rect 52850 -1045 52900 -925
rect 53200 -1045 53250 -925
rect 53550 -1045 53600 -925
rect 53900 -1045 53950 -925
rect 54250 -1045 54300 -925
rect 54600 -1045 54650 -925
rect 54950 -1045 55000 -925
rect 55300 -1045 55350 -925
rect 55650 -1045 55700 -925
rect 56000 -1045 56050 -925
rect 56350 -1045 56400 -925
rect 56700 -1045 56750 -925
rect 57050 -1045 57100 -925
rect 57400 -1045 57450 -925
rect 57750 -1045 57800 -925
rect 58100 -1045 58150 -925
rect 58450 -1045 58500 -925
rect 58800 -1045 58850 -925
rect 59150 -1045 59200 -925
rect 59500 -1045 59550 -925
rect 59850 -1045 59900 -925
rect 60200 -1045 60250 -925
rect 60550 -1045 60600 -925
rect 60900 -1045 60950 -925
rect 52060 -1130 52290 -1045
rect 52410 -1130 52640 -1045
rect 52760 -1130 52990 -1045
rect 52060 -1180 52990 -1130
rect 52060 -1275 52290 -1180
rect 52410 -1275 52640 -1180
rect 52760 -1275 52990 -1180
rect 53110 -1275 53340 -1045
rect 53460 -1275 53690 -1045
rect 53810 -1275 54040 -1045
rect 54160 -1275 54390 -1045
rect 54510 -1275 54740 -1045
rect 54860 -1275 55090 -1045
rect 55210 -1275 55440 -1045
rect 55560 -1275 55790 -1045
rect 55910 -1275 56140 -1045
rect 56260 -1275 56490 -1045
rect 56610 -1275 56840 -1045
rect 56960 -1275 57190 -1045
rect 57310 -1275 57540 -1045
rect 57660 -1275 57890 -1045
rect 58010 -1275 58240 -1045
rect 58360 -1275 58590 -1045
rect 58710 -1275 58940 -1045
rect 59060 -1275 59290 -1045
rect 59410 -1275 59640 -1045
rect 59760 -1275 59990 -1045
rect 60110 -1275 60340 -1045
rect 60460 -1275 60690 -1045
rect 60810 -1130 61040 -1045
rect 61160 -1130 61390 -1045
rect 61510 -1130 61740 -1045
rect 60810 -1180 61740 -1130
rect 60810 -1275 61040 -1180
rect 61160 -1275 61390 -1180
rect 61510 -1275 61740 -1180
<< via3 >>
rect 53995 1710 54035 1715
rect 53995 1680 54000 1710
rect 54000 1680 54030 1710
rect 54030 1680 54035 1710
rect 53995 1675 54035 1680
rect 54045 1710 54085 1715
rect 54045 1680 54050 1710
rect 54050 1680 54080 1710
rect 54080 1680 54085 1710
rect 54045 1675 54085 1680
rect 54095 1710 54135 1715
rect 54095 1680 54100 1710
rect 54100 1680 54130 1710
rect 54130 1680 54135 1710
rect 54095 1675 54135 1680
rect 54145 1710 54185 1715
rect 54145 1680 54150 1710
rect 54150 1680 54180 1710
rect 54180 1680 54185 1710
rect 54145 1675 54185 1680
rect 54195 1710 54235 1715
rect 54195 1680 54200 1710
rect 54200 1680 54230 1710
rect 54230 1680 54235 1710
rect 54195 1675 54235 1680
rect 53995 1660 54035 1665
rect 53995 1630 54000 1660
rect 54000 1630 54030 1660
rect 54030 1630 54035 1660
rect 53995 1625 54035 1630
rect 54045 1660 54085 1665
rect 54045 1630 54050 1660
rect 54050 1630 54080 1660
rect 54080 1630 54085 1660
rect 54045 1625 54085 1630
rect 54095 1660 54135 1665
rect 54095 1630 54100 1660
rect 54100 1630 54130 1660
rect 54130 1630 54135 1660
rect 54095 1625 54135 1630
rect 54145 1660 54185 1665
rect 54145 1630 54150 1660
rect 54150 1630 54180 1660
rect 54180 1630 54185 1660
rect 54145 1625 54185 1630
rect 54195 1660 54235 1665
rect 54195 1630 54200 1660
rect 54200 1630 54230 1660
rect 54230 1630 54235 1660
rect 54195 1625 54235 1630
rect 53995 1610 54035 1615
rect 53995 1580 54000 1610
rect 54000 1580 54030 1610
rect 54030 1580 54035 1610
rect 53995 1575 54035 1580
rect 54045 1610 54085 1615
rect 54045 1580 54050 1610
rect 54050 1580 54080 1610
rect 54080 1580 54085 1610
rect 54045 1575 54085 1580
rect 54095 1610 54135 1615
rect 54095 1580 54100 1610
rect 54100 1580 54130 1610
rect 54130 1580 54135 1610
rect 54095 1575 54135 1580
rect 54145 1610 54185 1615
rect 54145 1580 54150 1610
rect 54150 1580 54180 1610
rect 54180 1580 54185 1610
rect 54145 1575 54185 1580
rect 54195 1610 54235 1615
rect 54195 1580 54200 1610
rect 54200 1580 54230 1610
rect 54230 1580 54235 1610
rect 54195 1575 54235 1580
rect 59565 1710 59605 1715
rect 59565 1680 59570 1710
rect 59570 1680 59600 1710
rect 59600 1680 59605 1710
rect 59565 1675 59605 1680
rect 59615 1710 59655 1715
rect 59615 1680 59620 1710
rect 59620 1680 59650 1710
rect 59650 1680 59655 1710
rect 59615 1675 59655 1680
rect 59665 1710 59705 1715
rect 59665 1680 59670 1710
rect 59670 1680 59700 1710
rect 59700 1680 59705 1710
rect 59665 1675 59705 1680
rect 59715 1710 59755 1715
rect 59715 1680 59720 1710
rect 59720 1680 59750 1710
rect 59750 1680 59755 1710
rect 59715 1675 59755 1680
rect 59765 1710 59805 1715
rect 59765 1680 59770 1710
rect 59770 1680 59800 1710
rect 59800 1680 59805 1710
rect 59765 1675 59805 1680
rect 59565 1660 59605 1665
rect 59565 1630 59570 1660
rect 59570 1630 59600 1660
rect 59600 1630 59605 1660
rect 59565 1625 59605 1630
rect 59615 1660 59655 1665
rect 59615 1630 59620 1660
rect 59620 1630 59650 1660
rect 59650 1630 59655 1660
rect 59615 1625 59655 1630
rect 59665 1660 59705 1665
rect 59665 1630 59670 1660
rect 59670 1630 59700 1660
rect 59700 1630 59705 1660
rect 59665 1625 59705 1630
rect 59715 1660 59755 1665
rect 59715 1630 59720 1660
rect 59720 1630 59750 1660
rect 59750 1630 59755 1660
rect 59715 1625 59755 1630
rect 59765 1660 59805 1665
rect 59765 1630 59770 1660
rect 59770 1630 59800 1660
rect 59800 1630 59805 1660
rect 59765 1625 59805 1630
rect 59565 1610 59605 1615
rect 59565 1580 59570 1610
rect 59570 1580 59600 1610
rect 59600 1580 59605 1610
rect 59565 1575 59605 1580
rect 59615 1610 59655 1615
rect 59615 1580 59620 1610
rect 59620 1580 59650 1610
rect 59650 1580 59655 1610
rect 59615 1575 59655 1580
rect 59665 1610 59705 1615
rect 59665 1580 59670 1610
rect 59670 1580 59700 1610
rect 59700 1580 59705 1610
rect 59665 1575 59705 1580
rect 59715 1610 59755 1615
rect 59715 1580 59720 1610
rect 59720 1580 59750 1610
rect 59750 1580 59755 1610
rect 59715 1575 59755 1580
rect 59765 1610 59805 1615
rect 59765 1580 59770 1610
rect 59770 1580 59800 1610
rect 59800 1580 59805 1610
rect 59765 1575 59805 1580
<< mimcap >>
rect 52075 5515 52275 5590
rect 52075 5475 52155 5515
rect 52195 5475 52275 5515
rect 52075 5390 52275 5475
rect 52425 5515 52625 5590
rect 52425 5475 52505 5515
rect 52545 5475 52625 5515
rect 52425 5390 52625 5475
rect 52775 5515 52975 5590
rect 52775 5475 52855 5515
rect 52895 5475 52975 5515
rect 52775 5390 52975 5475
rect 53125 5515 53325 5590
rect 53125 5475 53205 5515
rect 53245 5475 53325 5515
rect 53125 5390 53325 5475
rect 53475 5515 53675 5590
rect 53475 5475 53555 5515
rect 53595 5475 53675 5515
rect 53475 5390 53675 5475
rect 53825 5515 54025 5590
rect 53825 5475 53905 5515
rect 53945 5475 54025 5515
rect 53825 5390 54025 5475
rect 54175 5515 54375 5590
rect 54175 5475 54255 5515
rect 54295 5475 54375 5515
rect 54175 5390 54375 5475
rect 54525 5515 54725 5590
rect 54525 5475 54605 5515
rect 54645 5475 54725 5515
rect 54525 5390 54725 5475
rect 54875 5515 55075 5590
rect 54875 5475 54955 5515
rect 54995 5475 55075 5515
rect 54875 5390 55075 5475
rect 55225 5515 55425 5590
rect 55225 5475 55305 5515
rect 55345 5475 55425 5515
rect 55225 5390 55425 5475
rect 55575 5515 55775 5590
rect 55575 5475 55655 5515
rect 55695 5475 55775 5515
rect 55575 5390 55775 5475
rect 55925 5515 56125 5590
rect 55925 5475 56005 5515
rect 56045 5475 56125 5515
rect 55925 5390 56125 5475
rect 56275 5515 56475 5590
rect 56275 5475 56355 5515
rect 56395 5475 56475 5515
rect 56275 5390 56475 5475
rect 56625 5515 56825 5590
rect 56625 5475 56705 5515
rect 56745 5475 56825 5515
rect 56625 5390 56825 5475
rect 56975 5515 57175 5590
rect 56975 5475 57055 5515
rect 57095 5475 57175 5515
rect 56975 5390 57175 5475
rect 57325 5515 57525 5590
rect 57325 5475 57405 5515
rect 57445 5475 57525 5515
rect 57325 5390 57525 5475
rect 57675 5515 57875 5590
rect 57675 5475 57755 5515
rect 57795 5475 57875 5515
rect 57675 5390 57875 5475
rect 58025 5515 58225 5590
rect 58025 5475 58105 5515
rect 58145 5475 58225 5515
rect 58025 5390 58225 5475
rect 58375 5515 58575 5590
rect 58375 5475 58455 5515
rect 58495 5475 58575 5515
rect 58375 5390 58575 5475
rect 58725 5515 58925 5590
rect 58725 5475 58805 5515
rect 58845 5475 58925 5515
rect 58725 5390 58925 5475
rect 59075 5515 59275 5590
rect 59075 5475 59155 5515
rect 59195 5475 59275 5515
rect 59075 5390 59275 5475
rect 59425 5515 59625 5590
rect 59425 5475 59505 5515
rect 59545 5475 59625 5515
rect 59425 5390 59625 5475
rect 59775 5515 59975 5590
rect 59775 5475 59855 5515
rect 59895 5475 59975 5515
rect 59775 5390 59975 5475
rect 60125 5515 60325 5590
rect 60125 5475 60205 5515
rect 60245 5475 60325 5515
rect 60125 5390 60325 5475
rect 60475 5515 60675 5590
rect 60475 5475 60555 5515
rect 60595 5475 60675 5515
rect 60475 5390 60675 5475
rect 60825 5515 61025 5590
rect 60825 5475 60905 5515
rect 60945 5475 61025 5515
rect 60825 5390 61025 5475
rect 61175 5515 61375 5590
rect 61175 5475 61255 5515
rect 61295 5475 61375 5515
rect 61175 5390 61375 5475
rect 61525 5515 61725 5590
rect 61525 5475 61605 5515
rect 61645 5475 61725 5515
rect 61525 5390 61725 5475
rect 52075 5165 52275 5240
rect 52075 5125 52155 5165
rect 52195 5125 52275 5165
rect 52075 5040 52275 5125
rect 52425 5165 52625 5240
rect 52425 5125 52505 5165
rect 52545 5125 52625 5165
rect 52425 5040 52625 5125
rect 52775 5165 52975 5240
rect 52775 5125 52855 5165
rect 52895 5125 52975 5165
rect 52775 5040 52975 5125
rect 53125 5165 53325 5240
rect 53125 5125 53205 5165
rect 53245 5125 53325 5165
rect 53125 5040 53325 5125
rect 53475 5165 53675 5240
rect 53475 5125 53555 5165
rect 53595 5125 53675 5165
rect 53475 5040 53675 5125
rect 53825 5165 54025 5240
rect 53825 5125 53905 5165
rect 53945 5125 54025 5165
rect 53825 5040 54025 5125
rect 54175 5165 54375 5240
rect 54175 5125 54255 5165
rect 54295 5125 54375 5165
rect 54175 5040 54375 5125
rect 54525 5165 54725 5240
rect 54525 5125 54605 5165
rect 54645 5125 54725 5165
rect 54525 5040 54725 5125
rect 54875 5165 55075 5240
rect 54875 5125 54955 5165
rect 54995 5125 55075 5165
rect 54875 5040 55075 5125
rect 55225 5155 55425 5240
rect 55225 5115 55305 5155
rect 55345 5115 55425 5155
rect 55225 5040 55425 5115
rect 55575 5155 55775 5240
rect 55575 5115 55655 5155
rect 55695 5115 55775 5155
rect 55575 5040 55775 5115
rect 58025 5155 58225 5240
rect 58025 5115 58105 5155
rect 58145 5115 58225 5155
rect 58025 5040 58225 5115
rect 58375 5155 58575 5240
rect 58375 5115 58455 5155
rect 58495 5115 58575 5155
rect 58375 5040 58575 5115
rect 58725 5165 58925 5240
rect 58725 5125 58805 5165
rect 58845 5125 58925 5165
rect 58725 5040 58925 5125
rect 59075 5165 59275 5240
rect 59075 5125 59155 5165
rect 59195 5125 59275 5165
rect 59075 5040 59275 5125
rect 59425 5165 59625 5240
rect 59425 5125 59505 5165
rect 59545 5125 59625 5165
rect 59425 5040 59625 5125
rect 59775 5165 59975 5240
rect 59775 5125 59855 5165
rect 59895 5125 59975 5165
rect 59775 5040 59975 5125
rect 60125 5165 60325 5240
rect 60125 5125 60205 5165
rect 60245 5125 60325 5165
rect 60125 5040 60325 5125
rect 60475 5165 60675 5240
rect 60475 5125 60555 5165
rect 60595 5125 60675 5165
rect 60475 5040 60675 5125
rect 60825 5165 61025 5240
rect 60825 5125 60905 5165
rect 60945 5125 61025 5165
rect 60825 5040 61025 5125
rect 61175 5165 61375 5240
rect 61175 5125 61255 5165
rect 61295 5125 61375 5165
rect 61175 5040 61375 5125
rect 61525 5165 61725 5240
rect 61525 5125 61605 5165
rect 61645 5125 61725 5165
rect 61525 5040 61725 5125
rect 52075 4815 52275 4890
rect 52075 4775 52155 4815
rect 52195 4775 52275 4815
rect 52075 4690 52275 4775
rect 52425 4815 52625 4890
rect 52425 4775 52505 4815
rect 52545 4775 52625 4815
rect 52425 4690 52625 4775
rect 52775 4815 52975 4890
rect 52775 4775 52855 4815
rect 52895 4775 52975 4815
rect 52775 4690 52975 4775
rect 53125 4815 53325 4890
rect 53125 4775 53205 4815
rect 53245 4775 53325 4815
rect 53125 4690 53325 4775
rect 53475 4815 53675 4890
rect 53475 4775 53555 4815
rect 53595 4775 53675 4815
rect 53475 4690 53675 4775
rect 53825 4815 54025 4890
rect 53825 4775 53905 4815
rect 53945 4775 54025 4815
rect 53825 4690 54025 4775
rect 54175 4815 54375 4890
rect 54175 4775 54255 4815
rect 54295 4775 54375 4815
rect 54175 4690 54375 4775
rect 54525 4815 54725 4890
rect 54525 4775 54605 4815
rect 54645 4775 54725 4815
rect 54525 4690 54725 4775
rect 54875 4815 55075 4890
rect 54875 4775 54955 4815
rect 54995 4775 55075 4815
rect 54875 4690 55075 4775
rect 55225 4805 55425 4890
rect 55225 4765 55305 4805
rect 55345 4765 55425 4805
rect 55225 4690 55425 4765
rect 58375 4805 58575 4890
rect 58375 4765 58455 4805
rect 58495 4765 58575 4805
rect 58375 4690 58575 4765
rect 58725 4815 58925 4890
rect 58725 4775 58805 4815
rect 58845 4775 58925 4815
rect 58725 4690 58925 4775
rect 59075 4815 59275 4890
rect 59075 4775 59155 4815
rect 59195 4775 59275 4815
rect 59075 4690 59275 4775
rect 59425 4815 59625 4890
rect 59425 4775 59505 4815
rect 59545 4775 59625 4815
rect 59425 4690 59625 4775
rect 59775 4815 59975 4890
rect 59775 4775 59855 4815
rect 59895 4775 59975 4815
rect 59775 4690 59975 4775
rect 60125 4815 60325 4890
rect 60125 4775 60205 4815
rect 60245 4775 60325 4815
rect 60125 4690 60325 4775
rect 60475 4815 60675 4890
rect 60475 4775 60555 4815
rect 60595 4775 60675 4815
rect 60475 4690 60675 4775
rect 60825 4815 61025 4890
rect 60825 4775 60905 4815
rect 60945 4775 61025 4815
rect 60825 4690 61025 4775
rect 61175 4815 61375 4890
rect 61175 4775 61255 4815
rect 61295 4775 61375 4815
rect 61175 4690 61375 4775
rect 61525 4815 61725 4890
rect 61525 4775 61605 4815
rect 61645 4775 61725 4815
rect 61525 4690 61725 4775
rect 52075 4465 52275 4540
rect 52075 4425 52155 4465
rect 52195 4425 52275 4465
rect 52075 4340 52275 4425
rect 52425 4465 52625 4540
rect 52425 4425 52505 4465
rect 52545 4425 52625 4465
rect 52425 4340 52625 4425
rect 52775 4465 52975 4540
rect 52775 4425 52855 4465
rect 52895 4425 52975 4465
rect 52775 4340 52975 4425
rect 53125 4465 53325 4540
rect 53125 4425 53205 4465
rect 53245 4425 53325 4465
rect 53125 4340 53325 4425
rect 53475 4465 53675 4540
rect 53475 4425 53555 4465
rect 53595 4425 53675 4465
rect 53475 4340 53675 4425
rect 60125 4465 60325 4540
rect 60125 4425 60205 4465
rect 60245 4425 60325 4465
rect 60125 4340 60325 4425
rect 60475 4465 60675 4540
rect 60475 4425 60555 4465
rect 60595 4425 60675 4465
rect 60475 4340 60675 4425
rect 60825 4465 61025 4540
rect 60825 4425 60905 4465
rect 60945 4425 61025 4465
rect 60825 4340 61025 4425
rect 61175 4465 61375 4540
rect 61175 4425 61255 4465
rect 61295 4425 61375 4465
rect 61175 4340 61375 4425
rect 61525 4465 61725 4540
rect 61525 4425 61605 4465
rect 61645 4425 61725 4465
rect 61525 4340 61725 4425
rect 52075 4115 52275 4190
rect 52075 4075 52155 4115
rect 52195 4075 52275 4115
rect 52075 3990 52275 4075
rect 52425 4115 52625 4190
rect 52425 4075 52505 4115
rect 52545 4075 52625 4115
rect 52425 3990 52625 4075
rect 52775 4115 52975 4190
rect 52775 4075 52855 4115
rect 52895 4075 52975 4115
rect 52775 3990 52975 4075
rect 53125 4115 53325 4190
rect 53125 4075 53205 4115
rect 53245 4075 53325 4115
rect 53125 3990 53325 4075
rect 53475 4115 53675 4190
rect 53475 4075 53555 4115
rect 53595 4075 53675 4115
rect 53475 3990 53675 4075
rect 60125 4115 60325 4190
rect 60125 4075 60205 4115
rect 60245 4075 60325 4115
rect 60125 3990 60325 4075
rect 60475 4115 60675 4190
rect 60475 4075 60555 4115
rect 60595 4075 60675 4115
rect 60475 3990 60675 4075
rect 60825 4115 61025 4190
rect 60825 4075 60905 4115
rect 60945 4075 61025 4115
rect 60825 3990 61025 4075
rect 61175 4115 61375 4190
rect 61175 4075 61255 4115
rect 61295 4075 61375 4115
rect 61175 3990 61375 4075
rect 61525 4115 61725 4190
rect 61525 4075 61605 4115
rect 61645 4075 61725 4115
rect 61525 3990 61725 4075
rect 52075 3765 52275 3840
rect 52075 3725 52155 3765
rect 52195 3725 52275 3765
rect 52075 3640 52275 3725
rect 52425 3765 52625 3840
rect 52425 3725 52505 3765
rect 52545 3725 52625 3765
rect 52425 3640 52625 3725
rect 52775 3765 52975 3840
rect 52775 3725 52855 3765
rect 52895 3725 52975 3765
rect 52775 3640 52975 3725
rect 53125 3765 53325 3840
rect 53125 3725 53205 3765
rect 53245 3725 53325 3765
rect 53125 3640 53325 3725
rect 53475 3765 53675 3840
rect 53475 3725 53555 3765
rect 53595 3725 53675 3765
rect 53475 3640 53675 3725
rect 60125 3765 60325 3840
rect 60125 3725 60205 3765
rect 60245 3725 60325 3765
rect 60125 3640 60325 3725
rect 60475 3765 60675 3840
rect 60475 3725 60555 3765
rect 60595 3725 60675 3765
rect 60475 3640 60675 3725
rect 60825 3765 61025 3840
rect 60825 3725 60905 3765
rect 60945 3725 61025 3765
rect 60825 3640 61025 3725
rect 61175 3765 61375 3840
rect 61175 3725 61255 3765
rect 61295 3725 61375 3765
rect 61175 3640 61375 3725
rect 61525 3765 61725 3840
rect 61525 3725 61605 3765
rect 61645 3725 61725 3765
rect 61525 3640 61725 3725
rect 52075 3415 52275 3490
rect 52075 3375 52155 3415
rect 52195 3375 52275 3415
rect 52075 3290 52275 3375
rect 52425 3415 52625 3490
rect 52425 3375 52505 3415
rect 52545 3375 52625 3415
rect 52425 3290 52625 3375
rect 52775 3415 52975 3490
rect 52775 3375 52855 3415
rect 52895 3375 52975 3415
rect 52775 3290 52975 3375
rect 53125 3415 53325 3490
rect 53125 3375 53205 3415
rect 53245 3375 53325 3415
rect 53125 3290 53325 3375
rect 53475 3415 53675 3490
rect 53475 3375 53555 3415
rect 53595 3375 53675 3415
rect 53475 3290 53675 3375
rect 60125 3415 60325 3490
rect 60125 3375 60205 3415
rect 60245 3375 60325 3415
rect 60125 3290 60325 3375
rect 60475 3415 60675 3490
rect 60475 3375 60555 3415
rect 60595 3375 60675 3415
rect 60475 3290 60675 3375
rect 60825 3415 61025 3490
rect 60825 3375 60905 3415
rect 60945 3375 61025 3415
rect 60825 3290 61025 3375
rect 61175 3415 61375 3490
rect 61175 3375 61255 3415
rect 61295 3375 61375 3415
rect 61175 3290 61375 3375
rect 61525 3415 61725 3490
rect 61525 3375 61605 3415
rect 61645 3375 61725 3415
rect 61525 3290 61725 3375
rect 52075 3065 52275 3140
rect 52075 3025 52155 3065
rect 52195 3025 52275 3065
rect 52075 2940 52275 3025
rect 52425 3065 52625 3140
rect 52425 3025 52505 3065
rect 52545 3025 52625 3065
rect 52425 2940 52625 3025
rect 52775 3065 52975 3140
rect 52775 3025 52855 3065
rect 52895 3025 52975 3065
rect 52775 2940 52975 3025
rect 53125 3065 53325 3140
rect 53125 3025 53205 3065
rect 53245 3025 53325 3065
rect 53125 2940 53325 3025
rect 53475 3065 53675 3140
rect 53475 3025 53555 3065
rect 53595 3025 53675 3065
rect 53475 2940 53675 3025
rect 60125 3065 60325 3140
rect 60125 3025 60205 3065
rect 60245 3025 60325 3065
rect 60125 2940 60325 3025
rect 60475 3065 60675 3140
rect 60475 3025 60555 3065
rect 60595 3025 60675 3065
rect 60475 2940 60675 3025
rect 60825 3065 61025 3140
rect 60825 3025 60905 3065
rect 60945 3025 61025 3065
rect 60825 2940 61025 3025
rect 61175 3065 61375 3140
rect 61175 3025 61255 3065
rect 61295 3025 61375 3065
rect 61175 2940 61375 3025
rect 61525 3065 61725 3140
rect 61525 3025 61605 3065
rect 61645 3025 61725 3065
rect 61525 2940 61725 3025
rect 52075 2715 52275 2790
rect 52075 2675 52155 2715
rect 52195 2675 52275 2715
rect 52075 2590 52275 2675
rect 52425 2715 52625 2790
rect 52425 2675 52505 2715
rect 52545 2675 52625 2715
rect 52425 2590 52625 2675
rect 52775 2715 52975 2790
rect 52775 2675 52855 2715
rect 52895 2675 52975 2715
rect 52775 2590 52975 2675
rect 53125 2715 53325 2790
rect 53125 2675 53205 2715
rect 53245 2675 53325 2715
rect 53125 2590 53325 2675
rect 53475 2715 53675 2790
rect 53475 2675 53555 2715
rect 53595 2675 53675 2715
rect 53475 2590 53675 2675
rect 60125 2715 60325 2790
rect 60125 2675 60205 2715
rect 60245 2675 60325 2715
rect 60125 2590 60325 2675
rect 60475 2715 60675 2790
rect 60475 2675 60555 2715
rect 60595 2675 60675 2715
rect 60475 2590 60675 2675
rect 60825 2715 61025 2790
rect 60825 2675 60905 2715
rect 60945 2675 61025 2715
rect 60825 2590 61025 2675
rect 61175 2715 61375 2790
rect 61175 2675 61255 2715
rect 61295 2675 61375 2715
rect 61175 2590 61375 2675
rect 61525 2715 61725 2790
rect 61525 2675 61605 2715
rect 61645 2675 61725 2715
rect 61525 2590 61725 2675
rect 52075 2365 52275 2440
rect 52075 2325 52155 2365
rect 52195 2325 52275 2365
rect 52075 2240 52275 2325
rect 52425 2365 52625 2440
rect 52425 2325 52505 2365
rect 52545 2325 52625 2365
rect 52425 2240 52625 2325
rect 52775 2365 52975 2440
rect 52775 2325 52855 2365
rect 52895 2325 52975 2365
rect 52775 2240 52975 2325
rect 53125 2365 53325 2440
rect 53125 2325 53205 2365
rect 53245 2325 53325 2365
rect 53125 2240 53325 2325
rect 53475 2365 53675 2440
rect 53475 2325 53555 2365
rect 53595 2325 53675 2365
rect 53475 2240 53675 2325
rect 60125 2365 60325 2440
rect 60125 2325 60205 2365
rect 60245 2325 60325 2365
rect 60125 2240 60325 2325
rect 60475 2365 60675 2440
rect 60475 2325 60555 2365
rect 60595 2325 60675 2365
rect 60475 2240 60675 2325
rect 60825 2365 61025 2440
rect 60825 2325 60905 2365
rect 60945 2325 61025 2365
rect 60825 2240 61025 2325
rect 61175 2365 61375 2440
rect 61175 2325 61255 2365
rect 61295 2325 61375 2365
rect 61175 2240 61375 2325
rect 61525 2365 61725 2440
rect 61525 2325 61605 2365
rect 61645 2325 61725 2365
rect 61525 2240 61725 2325
rect 52075 2015 52275 2090
rect 52075 1975 52155 2015
rect 52195 1975 52275 2015
rect 52075 1890 52275 1975
rect 52425 2015 52625 2090
rect 52425 1975 52505 2015
rect 52545 1975 52625 2015
rect 52425 1890 52625 1975
rect 52775 2015 52975 2090
rect 52775 1975 52855 2015
rect 52895 1975 52975 2015
rect 52775 1890 52975 1975
rect 53125 2015 53325 2090
rect 53125 1975 53205 2015
rect 53245 1975 53325 2015
rect 53125 1890 53325 1975
rect 53475 2015 53675 2090
rect 53475 1975 53555 2015
rect 53595 1975 53675 2015
rect 53475 1890 53675 1975
rect 60125 2015 60325 2090
rect 60125 1975 60205 2015
rect 60245 1975 60325 2015
rect 60125 1890 60325 1975
rect 60475 2015 60675 2090
rect 60475 1975 60555 2015
rect 60595 1975 60675 2015
rect 60475 1890 60675 1975
rect 60825 2015 61025 2090
rect 60825 1975 60905 2015
rect 60945 1975 61025 2015
rect 60825 1890 61025 1975
rect 61175 2015 61375 2090
rect 61175 1975 61255 2015
rect 61295 1975 61375 2015
rect 61175 1890 61375 1975
rect 61525 2015 61725 2090
rect 61525 1975 61605 2015
rect 61645 1975 61725 2015
rect 61525 1890 61725 1975
rect 52075 1665 52275 1740
rect 52075 1625 52155 1665
rect 52195 1625 52275 1665
rect 52075 1540 52275 1625
rect 52425 1665 52625 1740
rect 52425 1625 52505 1665
rect 52545 1625 52625 1665
rect 52425 1540 52625 1625
rect 52775 1665 52975 1740
rect 52775 1625 52855 1665
rect 52895 1625 52975 1665
rect 52775 1540 52975 1625
rect 53125 1665 53325 1740
rect 53125 1625 53205 1665
rect 53245 1625 53325 1665
rect 53125 1540 53325 1625
rect 53475 1665 53675 1740
rect 53475 1625 53555 1665
rect 53595 1625 53675 1665
rect 53475 1540 53675 1625
rect 60125 1665 60325 1740
rect 60125 1625 60205 1665
rect 60245 1625 60325 1665
rect 60125 1540 60325 1625
rect 60475 1665 60675 1740
rect 60475 1625 60555 1665
rect 60595 1625 60675 1665
rect 60475 1540 60675 1625
rect 60825 1665 61025 1740
rect 60825 1625 60905 1665
rect 60945 1625 61025 1665
rect 60825 1540 61025 1625
rect 61175 1665 61375 1740
rect 61175 1625 61255 1665
rect 61295 1625 61375 1665
rect 61175 1540 61375 1625
rect 61525 1665 61725 1740
rect 61525 1625 61605 1665
rect 61645 1625 61725 1665
rect 61525 1540 61725 1625
rect 52075 1315 52275 1390
rect 52075 1275 52155 1315
rect 52195 1275 52275 1315
rect 52075 1190 52275 1275
rect 52425 1315 52625 1390
rect 52425 1275 52505 1315
rect 52545 1275 52625 1315
rect 52425 1190 52625 1275
rect 52775 1315 52975 1390
rect 52775 1275 52855 1315
rect 52895 1275 52975 1315
rect 52775 1190 52975 1275
rect 53125 1315 53325 1390
rect 53125 1275 53205 1315
rect 53245 1275 53325 1315
rect 53125 1190 53325 1275
rect 53475 1315 53675 1390
rect 53475 1275 53555 1315
rect 53595 1275 53675 1315
rect 53475 1190 53675 1275
rect 60125 1315 60325 1390
rect 60125 1275 60205 1315
rect 60245 1275 60325 1315
rect 60125 1190 60325 1275
rect 60475 1315 60675 1390
rect 60475 1275 60555 1315
rect 60595 1275 60675 1315
rect 60475 1190 60675 1275
rect 60825 1315 61025 1390
rect 60825 1275 60905 1315
rect 60945 1275 61025 1315
rect 60825 1190 61025 1275
rect 61175 1315 61375 1390
rect 61175 1275 61255 1315
rect 61295 1275 61375 1315
rect 61175 1190 61375 1275
rect 61525 1315 61725 1390
rect 61525 1275 61605 1315
rect 61645 1275 61725 1315
rect 61525 1190 61725 1275
rect 52075 965 52275 1040
rect 52075 925 52155 965
rect 52195 925 52275 965
rect 52075 840 52275 925
rect 52425 965 52625 1040
rect 52425 925 52505 965
rect 52545 925 52625 965
rect 52425 840 52625 925
rect 52775 965 52975 1040
rect 52775 925 52855 965
rect 52895 925 52975 965
rect 52775 840 52975 925
rect 53125 965 53325 1040
rect 53125 925 53205 965
rect 53245 925 53325 965
rect 53125 840 53325 925
rect 53475 965 53675 1040
rect 53475 925 53555 965
rect 53595 925 53675 965
rect 53475 840 53675 925
rect 60125 965 60325 1040
rect 60125 925 60205 965
rect 60245 925 60325 965
rect 60125 840 60325 925
rect 60475 965 60675 1040
rect 60475 925 60555 965
rect 60595 925 60675 965
rect 60475 840 60675 925
rect 60825 965 61025 1040
rect 60825 925 60905 965
rect 60945 925 61025 965
rect 60825 840 61025 925
rect 61175 965 61375 1040
rect 61175 925 61255 965
rect 61295 925 61375 965
rect 61175 840 61375 925
rect 61525 965 61725 1040
rect 61525 925 61605 965
rect 61645 925 61725 965
rect 61525 840 61725 925
rect 52075 615 52275 690
rect 52075 575 52155 615
rect 52195 575 52275 615
rect 52075 490 52275 575
rect 52425 615 52625 690
rect 52425 575 52505 615
rect 52545 575 52625 615
rect 52425 490 52625 575
rect 52775 615 52975 690
rect 52775 575 52855 615
rect 52895 575 52975 615
rect 52775 490 52975 575
rect 53125 615 53325 690
rect 53125 575 53205 615
rect 53245 575 53325 615
rect 53125 490 53325 575
rect 53475 615 53675 690
rect 53475 575 53555 615
rect 53595 575 53675 615
rect 53475 490 53675 575
rect 60125 615 60325 690
rect 60125 575 60205 615
rect 60245 575 60325 615
rect 60125 490 60325 575
rect 60475 615 60675 690
rect 60475 575 60555 615
rect 60595 575 60675 615
rect 60475 490 60675 575
rect 60825 615 61025 690
rect 60825 575 60905 615
rect 60945 575 61025 615
rect 60825 490 61025 575
rect 61175 615 61375 690
rect 61175 575 61255 615
rect 61295 575 61375 615
rect 61175 490 61375 575
rect 61525 615 61725 690
rect 61525 575 61605 615
rect 61645 575 61725 615
rect 61525 490 61725 575
rect 52075 265 52275 340
rect 52075 225 52155 265
rect 52195 225 52275 265
rect 52075 140 52275 225
rect 52425 265 52625 340
rect 52425 225 52505 265
rect 52545 225 52625 265
rect 52425 140 52625 225
rect 52775 265 52975 340
rect 52775 225 52855 265
rect 52895 225 52975 265
rect 52775 140 52975 225
rect 53125 265 53325 340
rect 53125 225 53205 265
rect 53245 225 53325 265
rect 53125 140 53325 225
rect 53475 265 53675 340
rect 53475 225 53555 265
rect 53595 225 53675 265
rect 53475 140 53675 225
rect 60125 265 60325 340
rect 60125 225 60205 265
rect 60245 225 60325 265
rect 60125 140 60325 225
rect 60475 265 60675 340
rect 60475 225 60555 265
rect 60595 225 60675 265
rect 60475 140 60675 225
rect 60825 265 61025 340
rect 60825 225 60905 265
rect 60945 225 61025 265
rect 60825 140 61025 225
rect 61175 265 61375 340
rect 61175 225 61255 265
rect 61295 225 61375 265
rect 61175 140 61375 225
rect 61525 265 61725 340
rect 61525 225 61605 265
rect 61645 225 61725 265
rect 61525 140 61725 225
rect 52075 -85 52275 -10
rect 52075 -125 52155 -85
rect 52195 -125 52275 -85
rect 52075 -210 52275 -125
rect 52425 -85 52625 -10
rect 52425 -125 52505 -85
rect 52545 -125 52625 -85
rect 52425 -210 52625 -125
rect 52775 -85 52975 -10
rect 52775 -125 52855 -85
rect 52895 -125 52975 -85
rect 52775 -210 52975 -125
rect 53125 -85 53325 -10
rect 53125 -125 53205 -85
rect 53245 -125 53325 -85
rect 53125 -210 53325 -125
rect 53475 -85 53675 -10
rect 53475 -125 53555 -85
rect 53595 -125 53675 -85
rect 53475 -210 53675 -125
rect 60125 -85 60325 -10
rect 60125 -125 60205 -85
rect 60245 -125 60325 -85
rect 60125 -210 60325 -125
rect 60475 -85 60675 -10
rect 60475 -125 60555 -85
rect 60595 -125 60675 -85
rect 60475 -210 60675 -125
rect 60825 -85 61025 -10
rect 60825 -125 60905 -85
rect 60945 -125 61025 -85
rect 60825 -210 61025 -125
rect 61175 -85 61375 -10
rect 61175 -125 61255 -85
rect 61295 -125 61375 -85
rect 61175 -210 61375 -125
rect 61525 -85 61725 -10
rect 61525 -125 61605 -85
rect 61645 -125 61725 -85
rect 61525 -210 61725 -125
rect 52075 -435 52275 -360
rect 52075 -475 52155 -435
rect 52195 -475 52275 -435
rect 52075 -560 52275 -475
rect 52425 -435 52625 -360
rect 52425 -475 52505 -435
rect 52545 -475 52625 -435
rect 52425 -560 52625 -475
rect 52775 -435 52975 -360
rect 52775 -475 52855 -435
rect 52895 -475 52975 -435
rect 52775 -560 52975 -475
rect 53125 -435 53325 -360
rect 53125 -475 53205 -435
rect 53245 -475 53325 -435
rect 53125 -560 53325 -475
rect 53475 -435 53675 -360
rect 53475 -475 53555 -435
rect 53595 -475 53675 -435
rect 53475 -560 53675 -475
rect 60125 -435 60325 -360
rect 60125 -475 60205 -435
rect 60245 -475 60325 -435
rect 60125 -560 60325 -475
rect 60475 -435 60675 -360
rect 60475 -475 60555 -435
rect 60595 -475 60675 -435
rect 60475 -560 60675 -475
rect 60825 -435 61025 -360
rect 60825 -475 60905 -435
rect 60945 -475 61025 -435
rect 60825 -560 61025 -475
rect 61175 -435 61375 -360
rect 61175 -475 61255 -435
rect 61295 -475 61375 -435
rect 61175 -560 61375 -475
rect 61525 -435 61725 -360
rect 61525 -475 61605 -435
rect 61645 -475 61725 -435
rect 61525 -560 61725 -475
rect 52075 -785 52275 -710
rect 52075 -825 52155 -785
rect 52195 -825 52275 -785
rect 52075 -910 52275 -825
rect 52425 -785 52625 -710
rect 52425 -825 52505 -785
rect 52545 -825 52625 -785
rect 52425 -910 52625 -825
rect 52775 -785 52975 -710
rect 52775 -825 52855 -785
rect 52895 -825 52975 -785
rect 52775 -910 52975 -825
rect 53125 -785 53325 -710
rect 53125 -825 53205 -785
rect 53245 -825 53325 -785
rect 53125 -910 53325 -825
rect 53475 -785 53675 -710
rect 53475 -825 53555 -785
rect 53595 -825 53675 -785
rect 53475 -910 53675 -825
rect 53825 -785 54025 -710
rect 53825 -825 53905 -785
rect 53945 -825 54025 -785
rect 53825 -910 54025 -825
rect 54175 -785 54375 -710
rect 54175 -825 54255 -785
rect 54295 -825 54375 -785
rect 54175 -910 54375 -825
rect 54525 -785 54725 -710
rect 54525 -825 54605 -785
rect 54645 -825 54725 -785
rect 54525 -910 54725 -825
rect 54875 -785 55075 -710
rect 54875 -825 54955 -785
rect 54995 -825 55075 -785
rect 54875 -910 55075 -825
rect 55225 -785 55425 -710
rect 55225 -825 55305 -785
rect 55345 -825 55425 -785
rect 55225 -910 55425 -825
rect 55575 -785 55775 -710
rect 55575 -825 55655 -785
rect 55695 -825 55775 -785
rect 55575 -910 55775 -825
rect 55925 -785 56125 -710
rect 55925 -825 56005 -785
rect 56045 -825 56125 -785
rect 55925 -910 56125 -825
rect 56275 -785 56475 -710
rect 56275 -825 56355 -785
rect 56395 -825 56475 -785
rect 56275 -910 56475 -825
rect 56625 -785 56825 -710
rect 56625 -825 56705 -785
rect 56745 -825 56825 -785
rect 56625 -910 56825 -825
rect 56975 -785 57175 -710
rect 56975 -825 57055 -785
rect 57095 -825 57175 -785
rect 56975 -910 57175 -825
rect 57325 -785 57525 -710
rect 57325 -825 57405 -785
rect 57445 -825 57525 -785
rect 57325 -910 57525 -825
rect 57675 -785 57875 -710
rect 57675 -825 57755 -785
rect 57795 -825 57875 -785
rect 57675 -910 57875 -825
rect 58025 -785 58225 -710
rect 58025 -825 58105 -785
rect 58145 -825 58225 -785
rect 58025 -910 58225 -825
rect 58375 -785 58575 -710
rect 58375 -825 58455 -785
rect 58495 -825 58575 -785
rect 58375 -910 58575 -825
rect 58725 -785 58925 -710
rect 58725 -825 58805 -785
rect 58845 -825 58925 -785
rect 58725 -910 58925 -825
rect 59075 -785 59275 -710
rect 59075 -825 59155 -785
rect 59195 -825 59275 -785
rect 59075 -910 59275 -825
rect 59425 -785 59625 -710
rect 59425 -825 59505 -785
rect 59545 -825 59625 -785
rect 59425 -910 59625 -825
rect 59775 -785 59975 -710
rect 59775 -825 59855 -785
rect 59895 -825 59975 -785
rect 59775 -910 59975 -825
rect 60125 -785 60325 -710
rect 60125 -825 60205 -785
rect 60245 -825 60325 -785
rect 60125 -910 60325 -825
rect 60475 -785 60675 -710
rect 60475 -825 60555 -785
rect 60595 -825 60675 -785
rect 60475 -910 60675 -825
rect 60825 -785 61025 -710
rect 60825 -825 60905 -785
rect 60945 -825 61025 -785
rect 60825 -910 61025 -825
rect 61175 -785 61375 -710
rect 61175 -825 61255 -785
rect 61295 -825 61375 -785
rect 61175 -910 61375 -825
rect 61525 -785 61725 -710
rect 61525 -825 61605 -785
rect 61645 -825 61725 -785
rect 61525 -910 61725 -825
rect 52075 -1135 52275 -1060
rect 52075 -1175 52155 -1135
rect 52195 -1175 52275 -1135
rect 52075 -1260 52275 -1175
rect 52425 -1135 52625 -1060
rect 52425 -1175 52505 -1135
rect 52545 -1175 52625 -1135
rect 52425 -1260 52625 -1175
rect 52775 -1135 52975 -1060
rect 52775 -1175 52855 -1135
rect 52895 -1175 52975 -1135
rect 52775 -1260 52975 -1175
rect 53125 -1135 53325 -1060
rect 53125 -1175 53205 -1135
rect 53245 -1175 53325 -1135
rect 53125 -1260 53325 -1175
rect 53475 -1135 53675 -1060
rect 53475 -1175 53555 -1135
rect 53595 -1175 53675 -1135
rect 53475 -1260 53675 -1175
rect 53825 -1135 54025 -1060
rect 53825 -1175 53905 -1135
rect 53945 -1175 54025 -1135
rect 53825 -1260 54025 -1175
rect 54175 -1135 54375 -1060
rect 54175 -1175 54255 -1135
rect 54295 -1175 54375 -1135
rect 54175 -1260 54375 -1175
rect 54525 -1135 54725 -1060
rect 54525 -1175 54605 -1135
rect 54645 -1175 54725 -1135
rect 54525 -1260 54725 -1175
rect 54875 -1135 55075 -1060
rect 54875 -1175 54955 -1135
rect 54995 -1175 55075 -1135
rect 54875 -1260 55075 -1175
rect 55225 -1135 55425 -1060
rect 55225 -1175 55305 -1135
rect 55345 -1175 55425 -1135
rect 55225 -1260 55425 -1175
rect 55575 -1135 55775 -1060
rect 55575 -1175 55655 -1135
rect 55695 -1175 55775 -1135
rect 55575 -1260 55775 -1175
rect 55925 -1135 56125 -1060
rect 55925 -1175 56005 -1135
rect 56045 -1175 56125 -1135
rect 55925 -1260 56125 -1175
rect 56275 -1135 56475 -1060
rect 56275 -1175 56355 -1135
rect 56395 -1175 56475 -1135
rect 56275 -1260 56475 -1175
rect 56625 -1135 56825 -1060
rect 56625 -1175 56705 -1135
rect 56745 -1175 56825 -1135
rect 56625 -1260 56825 -1175
rect 56975 -1135 57175 -1060
rect 56975 -1175 57055 -1135
rect 57095 -1175 57175 -1135
rect 56975 -1260 57175 -1175
rect 57325 -1135 57525 -1060
rect 57325 -1175 57405 -1135
rect 57445 -1175 57525 -1135
rect 57325 -1260 57525 -1175
rect 57675 -1135 57875 -1060
rect 57675 -1175 57755 -1135
rect 57795 -1175 57875 -1135
rect 57675 -1260 57875 -1175
rect 58025 -1135 58225 -1060
rect 58025 -1175 58105 -1135
rect 58145 -1175 58225 -1135
rect 58025 -1260 58225 -1175
rect 58375 -1135 58575 -1060
rect 58375 -1175 58455 -1135
rect 58495 -1175 58575 -1135
rect 58375 -1260 58575 -1175
rect 58725 -1135 58925 -1060
rect 58725 -1175 58805 -1135
rect 58845 -1175 58925 -1135
rect 58725 -1260 58925 -1175
rect 59075 -1135 59275 -1060
rect 59075 -1175 59155 -1135
rect 59195 -1175 59275 -1135
rect 59075 -1260 59275 -1175
rect 59425 -1135 59625 -1060
rect 59425 -1175 59505 -1135
rect 59545 -1175 59625 -1135
rect 59425 -1260 59625 -1175
rect 59775 -1135 59975 -1060
rect 59775 -1175 59855 -1135
rect 59895 -1175 59975 -1135
rect 59775 -1260 59975 -1175
rect 60125 -1135 60325 -1060
rect 60125 -1175 60205 -1135
rect 60245 -1175 60325 -1135
rect 60125 -1260 60325 -1175
rect 60475 -1135 60675 -1060
rect 60475 -1175 60555 -1135
rect 60595 -1175 60675 -1135
rect 60475 -1260 60675 -1175
rect 60825 -1135 61025 -1060
rect 60825 -1175 60905 -1135
rect 60945 -1175 61025 -1135
rect 60825 -1260 61025 -1175
rect 61175 -1135 61375 -1060
rect 61175 -1175 61255 -1135
rect 61295 -1175 61375 -1135
rect 61175 -1260 61375 -1175
rect 61525 -1135 61725 -1060
rect 61525 -1175 61605 -1135
rect 61645 -1175 61725 -1135
rect 61525 -1260 61725 -1175
<< mimcapcontact >>
rect 52155 5475 52195 5515
rect 52505 5475 52545 5515
rect 52855 5475 52895 5515
rect 53205 5475 53245 5515
rect 53555 5475 53595 5515
rect 53905 5475 53945 5515
rect 54255 5475 54295 5515
rect 54605 5475 54645 5515
rect 54955 5475 54995 5515
rect 55305 5475 55345 5515
rect 55655 5475 55695 5515
rect 56005 5475 56045 5515
rect 56355 5475 56395 5515
rect 56705 5475 56745 5515
rect 57055 5475 57095 5515
rect 57405 5475 57445 5515
rect 57755 5475 57795 5515
rect 58105 5475 58145 5515
rect 58455 5475 58495 5515
rect 58805 5475 58845 5515
rect 59155 5475 59195 5515
rect 59505 5475 59545 5515
rect 59855 5475 59895 5515
rect 60205 5475 60245 5515
rect 60555 5475 60595 5515
rect 60905 5475 60945 5515
rect 61255 5475 61295 5515
rect 61605 5475 61645 5515
rect 52155 5125 52195 5165
rect 52505 5125 52545 5165
rect 52855 5125 52895 5165
rect 53205 5125 53245 5165
rect 53555 5125 53595 5165
rect 53905 5125 53945 5165
rect 54255 5125 54295 5165
rect 54605 5125 54645 5165
rect 54955 5125 54995 5165
rect 55305 5115 55345 5155
rect 55655 5115 55695 5155
rect 58105 5115 58145 5155
rect 58455 5115 58495 5155
rect 58805 5125 58845 5165
rect 59155 5125 59195 5165
rect 59505 5125 59545 5165
rect 59855 5125 59895 5165
rect 60205 5125 60245 5165
rect 60555 5125 60595 5165
rect 60905 5125 60945 5165
rect 61255 5125 61295 5165
rect 61605 5125 61645 5165
rect 52155 4775 52195 4815
rect 52505 4775 52545 4815
rect 52855 4775 52895 4815
rect 53205 4775 53245 4815
rect 53555 4775 53595 4815
rect 53905 4775 53945 4815
rect 54255 4775 54295 4815
rect 54605 4775 54645 4815
rect 54955 4775 54995 4815
rect 55305 4765 55345 4805
rect 58455 4765 58495 4805
rect 58805 4775 58845 4815
rect 59155 4775 59195 4815
rect 59505 4775 59545 4815
rect 59855 4775 59895 4815
rect 60205 4775 60245 4815
rect 60555 4775 60595 4815
rect 60905 4775 60945 4815
rect 61255 4775 61295 4815
rect 61605 4775 61645 4815
rect 52155 4425 52195 4465
rect 52505 4425 52545 4465
rect 52855 4425 52895 4465
rect 53205 4425 53245 4465
rect 53555 4425 53595 4465
rect 60205 4425 60245 4465
rect 60555 4425 60595 4465
rect 60905 4425 60945 4465
rect 61255 4425 61295 4465
rect 61605 4425 61645 4465
rect 52155 4075 52195 4115
rect 52505 4075 52545 4115
rect 52855 4075 52895 4115
rect 53205 4075 53245 4115
rect 53555 4075 53595 4115
rect 60205 4075 60245 4115
rect 60555 4075 60595 4115
rect 60905 4075 60945 4115
rect 61255 4075 61295 4115
rect 61605 4075 61645 4115
rect 52155 3725 52195 3765
rect 52505 3725 52545 3765
rect 52855 3725 52895 3765
rect 53205 3725 53245 3765
rect 53555 3725 53595 3765
rect 60205 3725 60245 3765
rect 60555 3725 60595 3765
rect 60905 3725 60945 3765
rect 61255 3725 61295 3765
rect 61605 3725 61645 3765
rect 52155 3375 52195 3415
rect 52505 3375 52545 3415
rect 52855 3375 52895 3415
rect 53205 3375 53245 3415
rect 53555 3375 53595 3415
rect 60205 3375 60245 3415
rect 60555 3375 60595 3415
rect 60905 3375 60945 3415
rect 61255 3375 61295 3415
rect 61605 3375 61645 3415
rect 52155 3025 52195 3065
rect 52505 3025 52545 3065
rect 52855 3025 52895 3065
rect 53205 3025 53245 3065
rect 53555 3025 53595 3065
rect 60205 3025 60245 3065
rect 60555 3025 60595 3065
rect 60905 3025 60945 3065
rect 61255 3025 61295 3065
rect 61605 3025 61645 3065
rect 52155 2675 52195 2715
rect 52505 2675 52545 2715
rect 52855 2675 52895 2715
rect 53205 2675 53245 2715
rect 53555 2675 53595 2715
rect 60205 2675 60245 2715
rect 60555 2675 60595 2715
rect 60905 2675 60945 2715
rect 61255 2675 61295 2715
rect 61605 2675 61645 2715
rect 52155 2325 52195 2365
rect 52505 2325 52545 2365
rect 52855 2325 52895 2365
rect 53205 2325 53245 2365
rect 53555 2325 53595 2365
rect 60205 2325 60245 2365
rect 60555 2325 60595 2365
rect 60905 2325 60945 2365
rect 61255 2325 61295 2365
rect 61605 2325 61645 2365
rect 52155 1975 52195 2015
rect 52505 1975 52545 2015
rect 52855 1975 52895 2015
rect 53205 1975 53245 2015
rect 53555 1975 53595 2015
rect 60205 1975 60245 2015
rect 60555 1975 60595 2015
rect 60905 1975 60945 2015
rect 61255 1975 61295 2015
rect 61605 1975 61645 2015
rect 52155 1625 52195 1665
rect 52505 1625 52545 1665
rect 52855 1625 52895 1665
rect 53205 1625 53245 1665
rect 53555 1625 53595 1665
rect 60205 1625 60245 1665
rect 60555 1625 60595 1665
rect 60905 1625 60945 1665
rect 61255 1625 61295 1665
rect 61605 1625 61645 1665
rect 52155 1275 52195 1315
rect 52505 1275 52545 1315
rect 52855 1275 52895 1315
rect 53205 1275 53245 1315
rect 53555 1275 53595 1315
rect 60205 1275 60245 1315
rect 60555 1275 60595 1315
rect 60905 1275 60945 1315
rect 61255 1275 61295 1315
rect 61605 1275 61645 1315
rect 52155 925 52195 965
rect 52505 925 52545 965
rect 52855 925 52895 965
rect 53205 925 53245 965
rect 53555 925 53595 965
rect 60205 925 60245 965
rect 60555 925 60595 965
rect 60905 925 60945 965
rect 61255 925 61295 965
rect 61605 925 61645 965
rect 52155 575 52195 615
rect 52505 575 52545 615
rect 52855 575 52895 615
rect 53205 575 53245 615
rect 53555 575 53595 615
rect 60205 575 60245 615
rect 60555 575 60595 615
rect 60905 575 60945 615
rect 61255 575 61295 615
rect 61605 575 61645 615
rect 52155 225 52195 265
rect 52505 225 52545 265
rect 52855 225 52895 265
rect 53205 225 53245 265
rect 53555 225 53595 265
rect 60205 225 60245 265
rect 60555 225 60595 265
rect 60905 225 60945 265
rect 61255 225 61295 265
rect 61605 225 61645 265
rect 52155 -125 52195 -85
rect 52505 -125 52545 -85
rect 52855 -125 52895 -85
rect 53205 -125 53245 -85
rect 53555 -125 53595 -85
rect 60205 -125 60245 -85
rect 60555 -125 60595 -85
rect 60905 -125 60945 -85
rect 61255 -125 61295 -85
rect 61605 -125 61645 -85
rect 52155 -475 52195 -435
rect 52505 -475 52545 -435
rect 52855 -475 52895 -435
rect 53205 -475 53245 -435
rect 53555 -475 53595 -435
rect 60205 -475 60245 -435
rect 60555 -475 60595 -435
rect 60905 -475 60945 -435
rect 61255 -475 61295 -435
rect 61605 -475 61645 -435
rect 52155 -825 52195 -785
rect 52505 -825 52545 -785
rect 52855 -825 52895 -785
rect 53205 -825 53245 -785
rect 53555 -825 53595 -785
rect 53905 -825 53945 -785
rect 54255 -825 54295 -785
rect 54605 -825 54645 -785
rect 54955 -825 54995 -785
rect 55305 -825 55345 -785
rect 55655 -825 55695 -785
rect 56005 -825 56045 -785
rect 56355 -825 56395 -785
rect 56705 -825 56745 -785
rect 57055 -825 57095 -785
rect 57405 -825 57445 -785
rect 57755 -825 57795 -785
rect 58105 -825 58145 -785
rect 58455 -825 58495 -785
rect 58805 -825 58845 -785
rect 59155 -825 59195 -785
rect 59505 -825 59545 -785
rect 59855 -825 59895 -785
rect 60205 -825 60245 -785
rect 60555 -825 60595 -785
rect 60905 -825 60945 -785
rect 61255 -825 61295 -785
rect 61605 -825 61645 -785
rect 52155 -1175 52195 -1135
rect 52505 -1175 52545 -1135
rect 52855 -1175 52895 -1135
rect 53205 -1175 53245 -1135
rect 53555 -1175 53595 -1135
rect 53905 -1175 53945 -1135
rect 54255 -1175 54295 -1135
rect 54605 -1175 54645 -1135
rect 54955 -1175 54995 -1135
rect 55305 -1175 55345 -1135
rect 55655 -1175 55695 -1135
rect 56005 -1175 56045 -1135
rect 56355 -1175 56395 -1135
rect 56705 -1175 56745 -1135
rect 57055 -1175 57095 -1135
rect 57405 -1175 57445 -1135
rect 57755 -1175 57795 -1135
rect 58105 -1175 58145 -1135
rect 58455 -1175 58495 -1135
rect 58805 -1175 58845 -1135
rect 59155 -1175 59195 -1135
rect 59505 -1175 59545 -1135
rect 59855 -1175 59895 -1135
rect 60205 -1175 60245 -1135
rect 60555 -1175 60595 -1135
rect 60905 -1175 60945 -1135
rect 61255 -1175 61295 -1135
rect 61605 -1175 61645 -1135
<< metal4 >>
rect 52150 5515 56750 5520
rect 52150 5475 52155 5515
rect 52195 5475 52505 5515
rect 52545 5475 52855 5515
rect 52895 5475 53205 5515
rect 53245 5475 53555 5515
rect 53595 5475 53905 5515
rect 53945 5475 54255 5515
rect 54295 5475 54605 5515
rect 54645 5475 54955 5515
rect 54995 5475 55305 5515
rect 55345 5475 55655 5515
rect 55695 5475 56005 5515
rect 56045 5475 56355 5515
rect 56395 5475 56705 5515
rect 56745 5475 56750 5515
rect 52150 5470 56750 5475
rect 57050 5515 61650 5520
rect 57050 5475 57055 5515
rect 57095 5475 57405 5515
rect 57445 5475 57755 5515
rect 57795 5475 58105 5515
rect 58145 5475 58455 5515
rect 58495 5475 58805 5515
rect 58845 5475 59155 5515
rect 59195 5475 59505 5515
rect 59545 5475 59855 5515
rect 59895 5475 60205 5515
rect 60245 5475 60555 5515
rect 60595 5475 60905 5515
rect 60945 5475 61255 5515
rect 61295 5475 61605 5515
rect 61645 5475 61650 5515
rect 57050 5470 61650 5475
rect 52850 5170 52900 5470
rect 52150 5165 53600 5170
rect 52150 5125 52155 5165
rect 52195 5125 52505 5165
rect 52545 5125 52855 5165
rect 52895 5125 53205 5165
rect 53245 5125 53555 5165
rect 53595 5125 53600 5165
rect 52150 5120 53600 5125
rect 53900 5165 53950 5470
rect 53900 5125 53905 5165
rect 53945 5125 53950 5165
rect 52850 4820 52900 5120
rect 52150 4815 53600 4820
rect 52150 4775 52155 4815
rect 52195 4775 52505 4815
rect 52545 4775 52855 4815
rect 52895 4775 53205 4815
rect 53245 4775 53555 4815
rect 53595 4775 53600 4815
rect 52150 4770 53600 4775
rect 53900 4815 53950 5125
rect 53900 4775 53905 4815
rect 53945 4775 53950 4815
rect 53900 4770 53950 4775
rect 54250 5165 54300 5470
rect 54250 5125 54255 5165
rect 54295 5125 54300 5165
rect 54250 4815 54300 5125
rect 54250 4775 54255 4815
rect 54295 4775 54300 4815
rect 54250 4770 54300 4775
rect 54600 5165 54650 5470
rect 54600 5125 54605 5165
rect 54645 5125 54650 5165
rect 54600 4815 54650 5125
rect 54600 4775 54605 4815
rect 54645 4775 54650 4815
rect 54600 4770 54650 4775
rect 54950 5165 55000 5470
rect 54950 5125 54955 5165
rect 54995 5125 55000 5165
rect 54950 4815 55000 5125
rect 54950 4775 54955 4815
rect 54995 4775 55000 4815
rect 54950 4770 55000 4775
rect 55300 5155 55350 5470
rect 55300 5115 55305 5155
rect 55345 5115 55350 5155
rect 55300 4805 55350 5115
rect 55650 5155 55700 5470
rect 55650 5115 55655 5155
rect 55695 5115 55700 5155
rect 55650 5110 55700 5115
rect 58100 5155 58150 5470
rect 58100 5115 58105 5155
rect 58145 5115 58150 5155
rect 58100 5110 58150 5115
rect 58450 5155 58500 5470
rect 58450 5115 58455 5155
rect 58495 5115 58500 5155
rect 52850 4470 52900 4770
rect 55300 4765 55305 4805
rect 55345 4765 55350 4805
rect 55300 4760 55350 4765
rect 58450 4805 58500 5115
rect 58450 4765 58455 4805
rect 58495 4765 58500 4805
rect 58800 5165 58850 5470
rect 58800 5125 58805 5165
rect 58845 5125 58850 5165
rect 58800 4815 58850 5125
rect 58800 4775 58805 4815
rect 58845 4775 58850 4815
rect 58800 4770 58850 4775
rect 59150 5165 59200 5470
rect 59150 5125 59155 5165
rect 59195 5125 59200 5165
rect 59150 4815 59200 5125
rect 59150 4775 59155 4815
rect 59195 4775 59200 4815
rect 59150 4770 59200 4775
rect 59500 5165 59550 5470
rect 59500 5125 59505 5165
rect 59545 5125 59550 5165
rect 59500 4815 59550 5125
rect 59500 4775 59505 4815
rect 59545 4775 59550 4815
rect 59500 4770 59550 4775
rect 59850 5165 59900 5470
rect 60900 5170 60950 5470
rect 59850 5125 59855 5165
rect 59895 5125 59900 5165
rect 59850 4815 59900 5125
rect 60200 5165 61650 5170
rect 60200 5125 60205 5165
rect 60245 5125 60555 5165
rect 60595 5125 60905 5165
rect 60945 5125 61255 5165
rect 61295 5125 61605 5165
rect 61645 5125 61650 5165
rect 60200 5120 61650 5125
rect 60900 4820 60950 5120
rect 59850 4775 59855 4815
rect 59895 4775 59900 4815
rect 59850 4770 59900 4775
rect 60200 4815 61650 4820
rect 60200 4775 60205 4815
rect 60245 4775 60555 4815
rect 60595 4775 60905 4815
rect 60945 4775 61255 4815
rect 61295 4775 61605 4815
rect 61645 4775 61650 4815
rect 60200 4770 61650 4775
rect 58450 4760 58500 4765
rect 60900 4470 60950 4770
rect 52150 4465 53600 4470
rect 52150 4425 52155 4465
rect 52195 4425 52505 4465
rect 52545 4425 52855 4465
rect 52895 4425 53205 4465
rect 53245 4425 53555 4465
rect 53595 4425 53600 4465
rect 52150 4420 53600 4425
rect 60200 4465 61650 4470
rect 60200 4425 60205 4465
rect 60245 4425 60555 4465
rect 60595 4425 60905 4465
rect 60945 4425 61255 4465
rect 61295 4425 61605 4465
rect 61645 4425 61650 4465
rect 60200 4420 61650 4425
rect 52850 4120 52900 4420
rect 60900 4120 60950 4420
rect 52150 4115 53600 4120
rect 52150 4075 52155 4115
rect 52195 4075 52505 4115
rect 52545 4075 52855 4115
rect 52895 4075 53205 4115
rect 53245 4075 53555 4115
rect 53595 4075 53600 4115
rect 52150 4070 53600 4075
rect 60200 4115 61650 4120
rect 60200 4075 60205 4115
rect 60245 4075 60555 4115
rect 60595 4075 60905 4115
rect 60945 4075 61255 4115
rect 61295 4075 61605 4115
rect 61645 4075 61650 4115
rect 60200 4070 61650 4075
rect 52850 3770 52900 4070
rect 60900 3770 60950 4070
rect 52150 3765 53600 3770
rect 52150 3725 52155 3765
rect 52195 3725 52505 3765
rect 52545 3725 52855 3765
rect 52895 3725 53205 3765
rect 53245 3725 53555 3765
rect 53595 3725 53600 3765
rect 52150 3720 53600 3725
rect 60200 3765 61650 3770
rect 60200 3725 60205 3765
rect 60245 3725 60555 3765
rect 60595 3725 60905 3765
rect 60945 3725 61255 3765
rect 61295 3725 61605 3765
rect 61645 3725 61650 3765
rect 60200 3720 61650 3725
rect 52850 3420 52900 3720
rect 60900 3420 60950 3720
rect 52150 3415 53600 3420
rect 52150 3375 52155 3415
rect 52195 3375 52505 3415
rect 52545 3375 52855 3415
rect 52895 3375 53205 3415
rect 53245 3375 53555 3415
rect 53595 3375 53600 3415
rect 52150 3370 53600 3375
rect 60200 3415 61650 3420
rect 60200 3375 60205 3415
rect 60245 3375 60555 3415
rect 60595 3375 60905 3415
rect 60945 3375 61255 3415
rect 61295 3375 61605 3415
rect 61645 3375 61650 3415
rect 60200 3370 61650 3375
rect 52850 3070 52900 3370
rect 60900 3070 60950 3370
rect 52150 3065 53600 3070
rect 52150 3025 52155 3065
rect 52195 3025 52505 3065
rect 52545 3025 52855 3065
rect 52895 3025 53205 3065
rect 53245 3025 53555 3065
rect 53595 3025 53600 3065
rect 52150 3020 53600 3025
rect 60200 3065 61650 3070
rect 60200 3025 60205 3065
rect 60245 3025 60555 3065
rect 60595 3025 60905 3065
rect 60945 3025 61255 3065
rect 61295 3025 61605 3065
rect 61645 3025 61650 3065
rect 60200 3020 61650 3025
rect 52850 2720 52900 3020
rect 60900 2720 60950 3020
rect 52150 2715 53600 2720
rect 52150 2675 52155 2715
rect 52195 2675 52505 2715
rect 52545 2675 52855 2715
rect 52895 2675 53205 2715
rect 53245 2675 53555 2715
rect 53595 2675 53600 2715
rect 52150 2670 53600 2675
rect 60200 2715 61650 2720
rect 60200 2675 60205 2715
rect 60245 2675 60555 2715
rect 60595 2675 60905 2715
rect 60945 2675 61255 2715
rect 61295 2675 61605 2715
rect 61645 2675 61650 2715
rect 60200 2670 61650 2675
rect 52850 2370 52900 2670
rect 60900 2370 60950 2670
rect 52150 2365 53600 2370
rect 52150 2325 52155 2365
rect 52195 2325 52505 2365
rect 52545 2325 52855 2365
rect 52895 2325 53205 2365
rect 53245 2325 53555 2365
rect 53595 2325 53600 2365
rect 52150 2320 53600 2325
rect 60200 2365 61650 2370
rect 60200 2325 60205 2365
rect 60245 2325 60555 2365
rect 60595 2325 60905 2365
rect 60945 2325 61255 2365
rect 61295 2325 61605 2365
rect 61645 2325 61650 2365
rect 60200 2320 61650 2325
rect 52850 2020 52900 2320
rect 60900 2020 60950 2320
rect 52150 2015 53600 2020
rect 52150 1975 52155 2015
rect 52195 1975 52505 2015
rect 52545 1975 52855 2015
rect 52895 1975 53205 2015
rect 53245 1975 53555 2015
rect 53595 1975 53600 2015
rect 52150 1970 53600 1975
rect 60200 2015 61650 2020
rect 60200 1975 60205 2015
rect 60245 1975 60555 2015
rect 60595 1975 60905 2015
rect 60945 1975 61255 2015
rect 61295 1975 61605 2015
rect 61645 1975 61650 2015
rect 60200 1970 61650 1975
rect 52850 1670 52900 1970
rect 53550 1715 54240 1720
rect 53550 1675 53995 1715
rect 54035 1675 54045 1715
rect 54085 1675 54095 1715
rect 54135 1675 54145 1715
rect 54185 1675 54195 1715
rect 54235 1675 54240 1715
rect 53550 1670 54240 1675
rect 52150 1665 54240 1670
rect 52150 1625 52155 1665
rect 52195 1625 52505 1665
rect 52545 1625 52855 1665
rect 52895 1625 53205 1665
rect 53245 1625 53555 1665
rect 53595 1625 53995 1665
rect 54035 1625 54045 1665
rect 54085 1625 54095 1665
rect 54135 1625 54145 1665
rect 54185 1625 54195 1665
rect 54235 1625 54240 1665
rect 52150 1620 54240 1625
rect 52850 1320 52900 1620
rect 53550 1615 54240 1620
rect 53550 1575 53995 1615
rect 54035 1575 54045 1615
rect 54085 1575 54095 1615
rect 54135 1575 54145 1615
rect 54185 1575 54195 1615
rect 54235 1575 54240 1615
rect 53550 1570 54240 1575
rect 59560 1715 60255 1720
rect 59560 1675 59565 1715
rect 59605 1675 59615 1715
rect 59655 1675 59665 1715
rect 59705 1675 59715 1715
rect 59755 1675 59765 1715
rect 59805 1675 60255 1715
rect 59560 1670 60255 1675
rect 60900 1670 60950 1970
rect 59560 1665 61650 1670
rect 59560 1625 59565 1665
rect 59605 1625 59615 1665
rect 59655 1625 59665 1665
rect 59705 1625 59715 1665
rect 59755 1625 59765 1665
rect 59805 1625 60205 1665
rect 60245 1625 60555 1665
rect 60595 1625 60905 1665
rect 60945 1625 61255 1665
rect 61295 1625 61605 1665
rect 61645 1625 61650 1665
rect 59560 1620 61650 1625
rect 59560 1615 60255 1620
rect 59560 1575 59565 1615
rect 59605 1575 59615 1615
rect 59655 1575 59665 1615
rect 59705 1575 59715 1615
rect 59755 1575 59765 1615
rect 59805 1575 60255 1615
rect 59560 1570 60255 1575
rect 60900 1320 60950 1620
rect 52150 1315 53600 1320
rect 52150 1275 52155 1315
rect 52195 1275 52505 1315
rect 52545 1275 52855 1315
rect 52895 1275 53205 1315
rect 53245 1275 53555 1315
rect 53595 1275 53600 1315
rect 52150 1270 53600 1275
rect 60200 1315 61650 1320
rect 60200 1275 60205 1315
rect 60245 1275 60555 1315
rect 60595 1275 60905 1315
rect 60945 1275 61255 1315
rect 61295 1275 61605 1315
rect 61645 1275 61650 1315
rect 60200 1270 61650 1275
rect 52850 970 52900 1270
rect 60900 970 60950 1270
rect 52150 965 53600 970
rect 52150 925 52155 965
rect 52195 925 52505 965
rect 52545 925 52855 965
rect 52895 925 53205 965
rect 53245 925 53555 965
rect 53595 925 53600 965
rect 52150 920 53600 925
rect 60200 965 61650 970
rect 60200 925 60205 965
rect 60245 925 60555 965
rect 60595 925 60905 965
rect 60945 925 61255 965
rect 61295 925 61605 965
rect 61645 925 61650 965
rect 60200 920 61650 925
rect 52850 620 52900 920
rect 60900 620 60950 920
rect 52150 615 53600 620
rect 52150 575 52155 615
rect 52195 575 52505 615
rect 52545 575 52855 615
rect 52895 575 53205 615
rect 53245 575 53555 615
rect 53595 575 53600 615
rect 52150 570 53600 575
rect 60200 615 61650 620
rect 60200 575 60205 615
rect 60245 575 60555 615
rect 60595 575 60905 615
rect 60945 575 61255 615
rect 61295 575 61605 615
rect 61645 575 61650 615
rect 60200 570 61650 575
rect 52850 270 52900 570
rect 60900 270 60950 570
rect 52150 265 53600 270
rect 52150 225 52155 265
rect 52195 225 52505 265
rect 52545 225 52855 265
rect 52895 225 53205 265
rect 53245 225 53555 265
rect 53595 225 53600 265
rect 52150 220 53600 225
rect 60200 265 61650 270
rect 60200 225 60205 265
rect 60245 225 60555 265
rect 60595 225 60905 265
rect 60945 225 61255 265
rect 61295 225 61605 265
rect 61645 225 61650 265
rect 60200 220 61650 225
rect 52850 -80 52900 220
rect 60900 -80 60950 220
rect 52150 -85 53600 -80
rect 52150 -125 52155 -85
rect 52195 -125 52505 -85
rect 52545 -125 52855 -85
rect 52895 -125 53205 -85
rect 53245 -125 53555 -85
rect 53595 -125 53600 -85
rect 52150 -130 53600 -125
rect 60200 -85 61650 -80
rect 60200 -125 60205 -85
rect 60245 -125 60555 -85
rect 60595 -125 60905 -85
rect 60945 -125 61255 -85
rect 61295 -125 61605 -85
rect 61645 -125 61650 -85
rect 60200 -130 61650 -125
rect 52850 -430 52900 -130
rect 60900 -430 60950 -130
rect 52150 -435 53600 -430
rect 52150 -475 52155 -435
rect 52195 -475 52505 -435
rect 52545 -475 52855 -435
rect 52895 -475 53205 -435
rect 53245 -475 53555 -435
rect 53595 -475 53600 -435
rect 52150 -480 53600 -475
rect 60200 -435 61650 -430
rect 60200 -475 60205 -435
rect 60245 -475 60555 -435
rect 60595 -475 60905 -435
rect 60945 -475 61255 -435
rect 61295 -475 61605 -435
rect 61645 -475 61650 -435
rect 60200 -480 61650 -475
rect 52850 -780 52900 -480
rect 60900 -780 60950 -480
rect 52150 -785 56750 -780
rect 52150 -825 52155 -785
rect 52195 -825 52505 -785
rect 52545 -825 52855 -785
rect 52895 -825 53205 -785
rect 53245 -825 53555 -785
rect 53595 -825 53905 -785
rect 53945 -825 54255 -785
rect 54295 -825 54605 -785
rect 54645 -825 54955 -785
rect 54995 -825 55305 -785
rect 55345 -825 55655 -785
rect 55695 -825 56005 -785
rect 56045 -825 56355 -785
rect 56395 -825 56705 -785
rect 56745 -825 56750 -785
rect 52150 -830 56750 -825
rect 52850 -1130 52900 -830
rect 52150 -1135 52900 -1130
rect 52150 -1175 52155 -1135
rect 52195 -1175 52505 -1135
rect 52545 -1175 52855 -1135
rect 52895 -1175 52900 -1135
rect 52150 -1180 52900 -1175
rect 53200 -1135 53250 -830
rect 53200 -1175 53205 -1135
rect 53245 -1175 53250 -1135
rect 53200 -1180 53250 -1175
rect 53550 -1135 53600 -830
rect 53550 -1175 53555 -1135
rect 53595 -1175 53600 -1135
rect 53550 -1180 53600 -1175
rect 53900 -1135 53950 -830
rect 53900 -1175 53905 -1135
rect 53945 -1175 53950 -1135
rect 53900 -1180 53950 -1175
rect 54250 -1135 54300 -830
rect 54250 -1175 54255 -1135
rect 54295 -1175 54300 -1135
rect 54250 -1180 54300 -1175
rect 54600 -1135 54650 -830
rect 54600 -1175 54605 -1135
rect 54645 -1175 54650 -1135
rect 54600 -1180 54650 -1175
rect 54950 -1135 55000 -830
rect 54950 -1175 54955 -1135
rect 54995 -1175 55000 -1135
rect 54950 -1180 55000 -1175
rect 55300 -1135 55350 -830
rect 55300 -1175 55305 -1135
rect 55345 -1175 55350 -1135
rect 55300 -1180 55350 -1175
rect 55650 -1135 55700 -830
rect 55650 -1175 55655 -1135
rect 55695 -1175 55700 -1135
rect 55650 -1180 55700 -1175
rect 56000 -1135 56050 -830
rect 56000 -1175 56005 -1135
rect 56045 -1175 56050 -1135
rect 56000 -1180 56050 -1175
rect 56350 -1135 56400 -830
rect 56350 -1175 56355 -1135
rect 56395 -1175 56400 -1135
rect 56350 -1180 56400 -1175
rect 56700 -1135 56750 -830
rect 56700 -1175 56705 -1135
rect 56745 -1175 56750 -1135
rect 56700 -1180 56750 -1175
rect 57050 -785 61650 -780
rect 57050 -825 57055 -785
rect 57095 -825 57405 -785
rect 57445 -825 57755 -785
rect 57795 -825 58105 -785
rect 58145 -825 58455 -785
rect 58495 -825 58805 -785
rect 58845 -825 59155 -785
rect 59195 -825 59505 -785
rect 59545 -825 59855 -785
rect 59895 -825 60205 -785
rect 60245 -825 60555 -785
rect 60595 -825 60905 -785
rect 60945 -825 61255 -785
rect 61295 -825 61605 -785
rect 61645 -825 61650 -785
rect 57050 -830 61650 -825
rect 57050 -1135 57100 -830
rect 57050 -1175 57055 -1135
rect 57095 -1175 57100 -1135
rect 57050 -1180 57100 -1175
rect 57400 -1135 57450 -830
rect 57400 -1175 57405 -1135
rect 57445 -1175 57450 -1135
rect 57400 -1180 57450 -1175
rect 57750 -1135 57800 -830
rect 57750 -1175 57755 -1135
rect 57795 -1175 57800 -1135
rect 57750 -1180 57800 -1175
rect 58100 -1135 58150 -830
rect 58100 -1175 58105 -1135
rect 58145 -1175 58150 -1135
rect 58100 -1180 58150 -1175
rect 58450 -1135 58500 -830
rect 58450 -1175 58455 -1135
rect 58495 -1175 58500 -1135
rect 58450 -1180 58500 -1175
rect 58800 -1135 58850 -830
rect 58800 -1175 58805 -1135
rect 58845 -1175 58850 -1135
rect 58800 -1180 58850 -1175
rect 59150 -1135 59200 -830
rect 59150 -1175 59155 -1135
rect 59195 -1175 59200 -1135
rect 59150 -1180 59200 -1175
rect 59500 -1135 59550 -830
rect 59500 -1175 59505 -1135
rect 59545 -1175 59550 -1135
rect 59500 -1180 59550 -1175
rect 59850 -1135 59900 -830
rect 59850 -1175 59855 -1135
rect 59895 -1175 59900 -1135
rect 59850 -1180 59900 -1175
rect 60200 -1135 60250 -830
rect 60200 -1175 60205 -1135
rect 60245 -1175 60250 -1135
rect 60200 -1180 60250 -1175
rect 60550 -1135 60600 -830
rect 60550 -1175 60555 -1135
rect 60595 -1175 60600 -1135
rect 60550 -1180 60600 -1175
rect 60900 -1130 60950 -830
rect 60900 -1135 61650 -1130
rect 60900 -1175 60905 -1135
rect 60945 -1175 61255 -1135
rect 61295 -1175 61605 -1135
rect 61645 -1175 61650 -1135
rect 60900 -1180 61650 -1175
<< labels >>
flabel metal2 57365 5060 57365 5060 1 FreeSans 240 0 0 80 Vb2_Vb3
flabel metal2 56455 5060 56455 5060 1 FreeSans 240 0 0 80 Vb2_2
flabel metal2 57000 3510 57000 3510 5 FreeSans 200 0 0 -80 Vb3
port 4 s
flabel metal1 56855 3545 56855 3545 5 FreeSans 200 0 0 -80 Vb2
port 5 s
flabel metal1 56945 655 56945 655 7 FreeSans 240 0 -80 0 V_tail_gate
port 11 w
flabel metal2 57770 1280 57770 1280 3 FreeSans 240 0 80 0 VIN-
flabel metal2 56030 1280 56030 1280 7 FreeSans 240 0 -80 0 VIN+
flabel metal1 57430 1325 57430 1325 3 FreeSans 240 0 80 0 VD1
flabel metal1 56370 1325 56370 1325 7 FreeSans 240 0 -80 0 VD2
flabel metal2 57455 2465 57455 2465 7 FreeSans 240 0 -80 0 X
flabel metal2 57525 2665 57525 2665 1 FreeSans 240 0 0 80 err_amp_out
flabel metal2 57000 2710 57000 2710 3 FreeSans 240 0 80 0 err_amp_mir
flabel metal2 56365 2815 56365 2815 7 FreeSans 240 0 -80 0 V_err_amp_ref
port 12 w
flabel metal2 57580 2775 57580 2775 1 FreeSans 240 0 0 160 V_tot
flabel metal1 56345 2455 56345 2455 3 FreeSans 240 0 80 0 Y
flabel metal2 57180 3205 57180 3205 3 FreeSans 240 0 80 0 V_err_p
flabel metal1 56620 3205 56620 3205 7 FreeSans 240 0 -80 0 V_err_mir_p
flabel metal2 57125 2885 57125 2885 3 FreeSans 240 0 80 0 V_err_gate
port 13 e
flabel metal2 57720 500 57720 500 5 FreeSans 200 0 0 -80 V_b_2nd_stage
flabel metal1 57220 530 57220 530 3 FreeSans 240 0 80 0 V_source
flabel metal2 56800 -200 56800 -200 1 FreeSans 240 0 0 80 Vb1_2
flabel metal2 56460 -55 56460 -55 1 FreeSans 240 0 0 80 V_p_mir
flabel metal2 55780 4070 55780 4070 5 FreeSans 240 0 0 -80 VD4
flabel metal2 54095 355 54095 355 5 FreeSans 240 0 0 -80 VOUT+
port 10 s
flabel metal2 54505 1665 54505 1665 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal2 54550 1480 54550 1480 1 FreeSans 240 0 0 80 V_CMFB_S4
port 8 n
flabel metal1 59705 355 59705 355 5 FreeSans 240 0 0 -80 VOUT-
port 9 s
flabel metal1 59250 1480 59250 1480 1 FreeSans 240 0 0 80 V_CMFB_S2
port 7 n
flabel metal1 59295 1665 59295 1665 1 FreeSans 240 0 0 80 V_CMFB_S1
port 2 n
flabel metal2 56900 1965 56900 1965 5 FreeSans 240 0 0 -80 Vb1
flabel metal3 54255 3435 54255 3435 7 FreeSans 240 0 -80 0 cap_res_Y
flabel metal3 59545 3435 59545 3435 3 FreeSans 240 0 80 0 cap_res_X
flabel metal2 58040 4070 58040 4070 5 FreeSans 240 0 0 -80 VD3
<< end >>
