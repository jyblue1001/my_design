magic
tech sky130A
timestamp 1754402060
<< metal1 >>
rect 2150 20910 2270 20925
rect 2150 20880 2195 20910
rect 2225 20880 2270 20910
rect 2150 20845 2270 20880
rect 2150 20815 2195 20845
rect 2225 20815 2270 20845
rect 2150 20775 2270 20815
rect 2150 20745 2195 20775
rect 2225 20745 2270 20775
rect 2150 20705 2270 20745
rect 2150 20675 2195 20705
rect 2225 20675 2270 20705
rect 2150 20635 2270 20675
rect 2150 20605 2195 20635
rect 2225 20605 2270 20635
rect 2150 20570 2270 20605
rect 2150 20540 2195 20570
rect 2225 20540 2270 20570
rect 2150 20510 2270 20540
rect 2150 20480 2195 20510
rect 2225 20480 2270 20510
rect 2150 20445 2270 20480
rect 2150 20415 2195 20445
rect 2225 20415 2270 20445
rect 2150 20375 2270 20415
rect 2150 20345 2195 20375
rect 2225 20345 2270 20375
rect 2150 20305 2270 20345
rect 2150 20275 2195 20305
rect 2225 20275 2270 20305
rect 2150 20235 2270 20275
rect 2150 20205 2195 20235
rect 2225 20205 2270 20235
rect 2150 20170 2270 20205
rect 2150 20140 2195 20170
rect 2225 20140 2270 20170
rect 2150 20110 2270 20140
rect 2150 20080 2195 20110
rect 2225 20080 2270 20110
rect 2150 20045 2270 20080
rect 2150 20015 2195 20045
rect 2225 20015 2270 20045
rect 2150 19975 2270 20015
rect 2150 19945 2195 19975
rect 2225 19945 2270 19975
rect 2150 19905 2270 19945
rect 2150 19875 2195 19905
rect 2225 19875 2270 19905
rect 2150 19835 2270 19875
rect 2150 19805 2195 19835
rect 2225 19805 2270 19835
rect 2150 19770 2270 19805
rect 2150 19740 2195 19770
rect 2225 19740 2270 19770
rect 2150 19710 2270 19740
rect 2150 19680 2195 19710
rect 2225 19680 2270 19710
rect 2150 19645 2270 19680
rect 2150 19615 2195 19645
rect 2225 19615 2270 19645
rect 2150 19575 2270 19615
rect 2150 19545 2195 19575
rect 2225 19545 2270 19575
rect 2150 19505 2270 19545
rect 2150 19475 2195 19505
rect 2225 19475 2270 19505
rect 2150 19435 2270 19475
rect 2150 19405 2195 19435
rect 2225 19405 2270 19435
rect 2150 19370 2270 19405
rect 2150 19340 2195 19370
rect 2225 19340 2270 19370
rect 2150 19310 2270 19340
rect 2150 19280 2195 19310
rect 2225 19280 2270 19310
rect 2150 19245 2270 19280
rect 2150 19215 2195 19245
rect 2225 19215 2270 19245
rect 2150 19175 2270 19215
rect 2150 19145 2195 19175
rect 2225 19145 2270 19175
rect 2150 19105 2270 19145
rect 2150 19075 2195 19105
rect 2225 19075 2270 19105
rect 2150 19035 2270 19075
rect 2150 19005 2195 19035
rect 2225 19005 2270 19035
rect 2150 18970 2270 19005
rect 2150 18940 2195 18970
rect 2225 18940 2270 18970
rect 2150 18910 2270 18940
rect 2150 18880 2195 18910
rect 2225 18880 2270 18910
rect 2150 18845 2270 18880
rect 2150 18815 2195 18845
rect 2225 18815 2270 18845
rect 2150 18775 2270 18815
rect 2150 18745 2195 18775
rect 2225 18745 2270 18775
rect 2150 18705 2270 18745
rect 2150 18675 2195 18705
rect 2225 18675 2270 18705
rect 2150 18635 2270 18675
rect 2150 18605 2195 18635
rect 2225 18605 2270 18635
rect 2150 18570 2270 18605
rect 2150 18540 2195 18570
rect 2225 18540 2270 18570
rect 2150 18510 2270 18540
rect 2150 18480 2195 18510
rect 2225 18480 2270 18510
rect 2150 18445 2270 18480
rect 2150 18415 2195 18445
rect 2225 18415 2270 18445
rect 2150 18375 2270 18415
rect 2150 18345 2195 18375
rect 2225 18345 2270 18375
rect 2150 18305 2270 18345
rect 2150 18275 2195 18305
rect 2225 18275 2270 18305
rect 2150 18235 2270 18275
rect 2150 18205 2195 18235
rect 2225 18205 2270 18235
rect 2150 18170 2270 18205
rect 2150 18140 2195 18170
rect 2225 18140 2270 18170
rect 2150 18110 2270 18140
rect 2150 18080 2195 18110
rect 2225 18080 2270 18110
rect 2150 18045 2270 18080
rect 2150 18015 2195 18045
rect 2225 18015 2270 18045
rect 2150 17975 2270 18015
rect 2150 17945 2195 17975
rect 2225 17945 2270 17975
rect 2150 17905 2270 17945
rect 2150 17875 2195 17905
rect 2225 17875 2270 17905
rect 2150 17835 2270 17875
rect 2150 17805 2195 17835
rect 2225 17805 2270 17835
rect 2150 17770 2270 17805
rect 2150 17740 2195 17770
rect 2225 17740 2270 17770
rect 2150 15780 2270 17740
rect 6650 20910 6710 20925
rect 6650 20880 6665 20910
rect 6695 20880 6710 20910
rect 6650 20845 6710 20880
rect 6650 20815 6665 20845
rect 6695 20815 6710 20845
rect 6650 20775 6710 20815
rect 6650 20745 6665 20775
rect 6695 20745 6710 20775
rect 6650 20705 6710 20745
rect 6650 20675 6665 20705
rect 6695 20675 6710 20705
rect 6650 20635 6710 20675
rect 6650 20605 6665 20635
rect 6695 20605 6710 20635
rect 6650 20570 6710 20605
rect 6650 20540 6665 20570
rect 6695 20540 6710 20570
rect 6650 20510 6710 20540
rect 6650 20480 6665 20510
rect 6695 20480 6710 20510
rect 6650 20445 6710 20480
rect 6650 20415 6665 20445
rect 6695 20415 6710 20445
rect 6650 20375 6710 20415
rect 6650 20345 6665 20375
rect 6695 20345 6710 20375
rect 6650 20305 6710 20345
rect 6650 20275 6665 20305
rect 6695 20275 6710 20305
rect 6650 20235 6710 20275
rect 6650 20205 6665 20235
rect 6695 20205 6710 20235
rect 6650 20170 6710 20205
rect 6650 20140 6665 20170
rect 6695 20140 6710 20170
rect 6650 20110 6710 20140
rect 6650 20080 6665 20110
rect 6695 20080 6710 20110
rect 6650 20045 6710 20080
rect 6650 20015 6665 20045
rect 6695 20015 6710 20045
rect 6650 19975 6710 20015
rect 6650 19945 6665 19975
rect 6695 19945 6710 19975
rect 6650 19905 6710 19945
rect 6650 19875 6665 19905
rect 6695 19875 6710 19905
rect 6650 19835 6710 19875
rect 6650 19805 6665 19835
rect 6695 19805 6710 19835
rect 6650 19770 6710 19805
rect 6650 19740 6665 19770
rect 6695 19740 6710 19770
rect 6650 19710 6710 19740
rect 6650 19680 6665 19710
rect 6695 19680 6710 19710
rect 6650 19645 6710 19680
rect 6650 19615 6665 19645
rect 6695 19615 6710 19645
rect 6650 19575 6710 19615
rect 6650 19545 6665 19575
rect 6695 19545 6710 19575
rect 6650 19505 6710 19545
rect 6650 19475 6665 19505
rect 6695 19475 6710 19505
rect 6650 19435 6710 19475
rect 6650 19405 6665 19435
rect 6695 19405 6710 19435
rect 6650 19370 6710 19405
rect 6650 19340 6665 19370
rect 6695 19340 6710 19370
rect 6650 19310 6710 19340
rect 6650 19280 6665 19310
rect 6695 19280 6710 19310
rect 6650 19245 6710 19280
rect 6650 19215 6665 19245
rect 6695 19215 6710 19245
rect 6650 19175 6710 19215
rect 6650 19145 6665 19175
rect 6695 19145 6710 19175
rect 6650 19105 6710 19145
rect 6650 19075 6665 19105
rect 6695 19075 6710 19105
rect 6650 19035 6710 19075
rect 6650 19005 6665 19035
rect 6695 19005 6710 19035
rect 6650 18970 6710 19005
rect 6650 18940 6665 18970
rect 6695 18940 6710 18970
rect 6650 18910 6710 18940
rect 6650 18880 6665 18910
rect 6695 18880 6710 18910
rect 6650 18845 6710 18880
rect 6650 18815 6665 18845
rect 6695 18815 6710 18845
rect 6650 18775 6710 18815
rect 6650 18745 6665 18775
rect 6695 18745 6710 18775
rect 6650 18705 6710 18745
rect 6650 18675 6665 18705
rect 6695 18675 6710 18705
rect 6650 18635 6710 18675
rect 6650 18605 6665 18635
rect 6695 18605 6710 18635
rect 6650 18570 6710 18605
rect 6650 18540 6665 18570
rect 6695 18540 6710 18570
rect 6650 18510 6710 18540
rect 6650 18480 6665 18510
rect 6695 18480 6710 18510
rect 6650 18445 6710 18480
rect 6650 18415 6665 18445
rect 6695 18415 6710 18445
rect 6650 18375 6710 18415
rect 6650 18345 6665 18375
rect 6695 18345 6710 18375
rect 6650 18305 6710 18345
rect 6650 18275 6665 18305
rect 6695 18275 6710 18305
rect 6650 18235 6710 18275
rect 6650 18205 6665 18235
rect 6695 18205 6710 18235
rect 6650 18170 6710 18205
rect 6650 18140 6665 18170
rect 6695 18140 6710 18170
rect 6650 18110 6710 18140
rect 6650 18080 6665 18110
rect 6695 18080 6710 18110
rect 6650 18045 6710 18080
rect 6650 18015 6665 18045
rect 6695 18015 6710 18045
rect 6650 17975 6710 18015
rect 6650 17945 6665 17975
rect 6695 17945 6710 17975
rect 6650 17905 6710 17945
rect 6650 17875 6665 17905
rect 6695 17875 6710 17905
rect 6650 17835 6710 17875
rect 6650 17805 6665 17835
rect 6695 17805 6710 17835
rect 6650 17770 6710 17805
rect 6650 17740 6665 17770
rect 6695 17740 6710 17770
rect 6650 17725 6710 17740
rect 2150 15750 2155 15780
rect 2185 15750 2195 15780
rect 2225 15750 2235 15780
rect 2265 15750 2270 15780
rect 2150 15740 2270 15750
rect 2150 15710 2155 15740
rect 2185 15710 2195 15740
rect 2225 15710 2235 15740
rect 2265 15710 2270 15740
rect 2150 15700 2270 15710
rect 2150 15670 2155 15700
rect 2185 15670 2195 15700
rect 2225 15670 2235 15700
rect 2265 15670 2270 15700
rect 2150 12720 2270 15670
rect 2150 12690 2155 12720
rect 2185 12690 2195 12720
rect 2225 12690 2235 12720
rect 2265 12690 2270 12720
rect 2150 12680 2270 12690
rect 2150 12650 2155 12680
rect 2185 12650 2195 12680
rect 2225 12650 2235 12680
rect 2265 12650 2270 12680
rect 2150 12560 2270 12650
rect 2150 12530 2155 12560
rect 2185 12530 2195 12560
rect 2225 12530 2235 12560
rect 2265 12530 2270 12560
rect 2150 12520 2270 12530
rect 2150 12490 2155 12520
rect 2185 12490 2195 12520
rect 2225 12490 2235 12520
rect 2265 12490 2270 12520
rect 2150 12480 2270 12490
rect 2150 12450 2155 12480
rect 2185 12450 2195 12480
rect 2225 12450 2235 12480
rect 2265 12450 2270 12480
rect 2150 12445 2270 12450
rect 2285 15925 2405 15930
rect 2285 15895 2290 15925
rect 2320 15895 2330 15925
rect 2360 15895 2370 15925
rect 2400 15895 2405 15925
rect -120 9635 0 9650
rect -120 9605 -75 9635
rect -45 9605 0 9635
rect -120 9570 0 9605
rect -120 9540 -75 9570
rect -45 9540 0 9570
rect -120 9500 0 9540
rect -120 9470 -75 9500
rect -45 9470 0 9500
rect -120 9430 0 9470
rect -120 9400 -75 9430
rect -45 9400 0 9430
rect -120 9360 0 9400
rect -120 9330 -75 9360
rect -45 9330 0 9360
rect -120 9295 0 9330
rect -120 9265 -75 9295
rect -45 9265 0 9295
rect -120 9235 0 9265
rect -120 9205 -75 9235
rect -45 9205 0 9235
rect -120 9170 0 9205
rect -120 9140 -75 9170
rect -45 9140 0 9170
rect -120 9100 0 9140
rect -120 9070 -75 9100
rect -45 9070 0 9100
rect -120 9030 0 9070
rect -120 9000 -75 9030
rect -45 9000 0 9030
rect -120 8960 0 9000
rect -120 8930 -75 8960
rect -45 8930 0 8960
rect -120 8895 0 8930
rect -120 8865 -75 8895
rect -45 8865 0 8895
rect -120 8835 0 8865
rect -120 8805 -75 8835
rect -45 8805 0 8835
rect -120 8770 0 8805
rect -120 8740 -75 8770
rect -45 8740 0 8770
rect -120 8700 0 8740
rect -120 8670 -75 8700
rect -45 8670 0 8700
rect -120 8630 0 8670
rect -120 8600 -75 8630
rect -45 8600 0 8630
rect -120 8560 0 8600
rect -120 8530 -75 8560
rect -45 8530 0 8560
rect -120 8495 0 8530
rect -120 8465 -75 8495
rect -45 8465 0 8495
rect -120 8435 0 8465
rect -120 8405 -75 8435
rect -45 8405 0 8435
rect -120 8370 0 8405
rect -120 8340 -75 8370
rect -45 8340 0 8370
rect -120 8300 0 8340
rect -120 8270 -75 8300
rect -45 8270 0 8300
rect -120 8230 0 8270
rect -120 8200 -75 8230
rect -45 8200 0 8230
rect -120 8160 0 8200
rect -120 8130 -75 8160
rect -45 8130 0 8160
rect -120 8095 0 8130
rect -120 8065 -75 8095
rect -45 8065 0 8095
rect -120 8035 0 8065
rect -120 8005 -75 8035
rect -45 8005 0 8035
rect -120 7970 0 8005
rect -120 7940 -75 7970
rect -45 7940 0 7970
rect -120 7900 0 7940
rect -120 7870 -75 7900
rect -45 7870 0 7900
rect -120 7830 0 7870
rect -120 7800 -75 7830
rect -45 7800 0 7830
rect -120 7760 0 7800
rect -120 7730 -75 7760
rect -45 7730 0 7760
rect -120 7695 0 7730
rect -120 7665 -75 7695
rect -45 7665 0 7695
rect -120 7635 0 7665
rect -120 7605 -75 7635
rect -45 7605 0 7635
rect -120 7570 0 7605
rect -120 7540 -75 7570
rect -45 7540 0 7570
rect -120 7500 0 7540
rect -120 7470 -75 7500
rect -45 7470 0 7500
rect -120 7430 0 7470
rect -120 7400 -75 7430
rect -45 7400 0 7430
rect -120 7360 0 7400
rect -120 7330 -75 7360
rect -45 7330 0 7360
rect -120 7295 0 7330
rect -120 7265 -75 7295
rect -45 7265 0 7295
rect -120 7235 0 7265
rect -120 7205 -75 7235
rect -45 7205 0 7235
rect -120 7170 0 7205
rect -120 7140 -75 7170
rect -45 7140 0 7170
rect -120 7100 0 7140
rect -120 7070 -75 7100
rect -45 7070 0 7100
rect -120 7030 0 7070
rect -120 7000 -75 7030
rect -45 7000 0 7030
rect -120 6960 0 7000
rect -120 6930 -75 6960
rect -45 6930 0 6960
rect -120 6895 0 6930
rect -120 6865 -75 6895
rect -45 6865 0 6895
rect -120 6835 0 6865
rect -120 6805 -75 6835
rect -45 6805 0 6835
rect -120 6770 0 6805
rect -120 6740 -75 6770
rect -45 6740 0 6770
rect -120 6700 0 6740
rect -120 6670 -75 6700
rect -45 6670 0 6700
rect -120 6630 0 6670
rect -120 6600 -75 6630
rect -45 6600 0 6630
rect -120 6560 0 6600
rect -120 6530 -75 6560
rect -45 6530 0 6560
rect -120 6495 0 6530
rect -120 6465 -75 6495
rect -45 6465 0 6495
rect -120 6210 0 6465
rect 230 9635 350 9650
rect 230 9605 275 9635
rect 305 9605 350 9635
rect 230 9570 350 9605
rect 230 9540 275 9570
rect 305 9540 350 9570
rect 230 9500 350 9540
rect 230 9470 275 9500
rect 305 9470 350 9500
rect 230 9430 350 9470
rect 230 9400 275 9430
rect 305 9400 350 9430
rect 230 9360 350 9400
rect 230 9330 275 9360
rect 305 9330 350 9360
rect 230 9295 350 9330
rect 230 9265 275 9295
rect 305 9265 350 9295
rect 230 9235 350 9265
rect 230 9205 275 9235
rect 305 9205 350 9235
rect 230 9170 350 9205
rect 230 9140 275 9170
rect 305 9140 350 9170
rect 230 9100 350 9140
rect 230 9070 275 9100
rect 305 9070 350 9100
rect 230 9030 350 9070
rect 230 9000 275 9030
rect 305 9000 350 9030
rect 230 8960 350 9000
rect 230 8930 275 8960
rect 305 8930 350 8960
rect 230 8895 350 8930
rect 230 8865 275 8895
rect 305 8865 350 8895
rect 230 8835 350 8865
rect 230 8805 275 8835
rect 305 8805 350 8835
rect 230 8770 350 8805
rect 230 8740 275 8770
rect 305 8740 350 8770
rect 230 8700 350 8740
rect 230 8670 275 8700
rect 305 8670 350 8700
rect 230 8630 350 8670
rect 230 8600 275 8630
rect 305 8600 350 8630
rect 230 8560 350 8600
rect 230 8530 275 8560
rect 305 8530 350 8560
rect 230 8495 350 8530
rect 230 8465 275 8495
rect 305 8465 350 8495
rect 230 8435 350 8465
rect 230 8405 275 8435
rect 305 8405 350 8435
rect 230 8370 350 8405
rect 230 8340 275 8370
rect 305 8340 350 8370
rect 230 8300 350 8340
rect 230 8270 275 8300
rect 305 8270 350 8300
rect 230 8230 350 8270
rect 230 8200 275 8230
rect 305 8200 350 8230
rect 230 8160 350 8200
rect 230 8130 275 8160
rect 305 8130 350 8160
rect 230 8095 350 8130
rect 230 8065 275 8095
rect 305 8065 350 8095
rect 230 8035 350 8065
rect 230 8005 275 8035
rect 305 8005 350 8035
rect 230 7970 350 8005
rect 230 7940 275 7970
rect 305 7940 350 7970
rect 230 7900 350 7940
rect 230 7870 275 7900
rect 305 7870 350 7900
rect 230 7830 350 7870
rect 230 7800 275 7830
rect 305 7800 350 7830
rect 230 7760 350 7800
rect 230 7730 275 7760
rect 305 7730 350 7760
rect 230 7695 350 7730
rect 230 7665 275 7695
rect 305 7665 350 7695
rect 230 7635 350 7665
rect 230 7605 275 7635
rect 305 7605 350 7635
rect 230 7570 350 7605
rect 230 7540 275 7570
rect 305 7540 350 7570
rect 230 7500 350 7540
rect 230 7470 275 7500
rect 305 7470 350 7500
rect 230 7430 350 7470
rect 230 7400 275 7430
rect 305 7400 350 7430
rect 230 7360 350 7400
rect 230 7330 275 7360
rect 305 7330 350 7360
rect 230 7295 350 7330
rect 230 7265 275 7295
rect 305 7265 350 7295
rect 230 7235 350 7265
rect 230 7205 275 7235
rect 305 7205 350 7235
rect 230 7170 350 7205
rect 230 7140 275 7170
rect 305 7140 350 7170
rect 230 7100 350 7140
rect 230 7070 275 7100
rect 305 7070 350 7100
rect 230 7030 350 7070
rect 230 7000 275 7030
rect 305 7000 350 7030
rect 230 6960 350 7000
rect 230 6930 275 6960
rect 305 6930 350 6960
rect 230 6895 350 6930
rect 230 6865 275 6895
rect 305 6865 350 6895
rect 230 6835 350 6865
rect 230 6805 275 6835
rect 305 6805 350 6835
rect 230 6770 350 6805
rect 230 6740 275 6770
rect 305 6740 350 6770
rect 230 6700 350 6740
rect 230 6670 275 6700
rect 305 6670 350 6700
rect 230 6630 350 6670
rect 230 6600 275 6630
rect 305 6600 350 6630
rect 230 6560 350 6600
rect 230 6530 275 6560
rect 305 6530 350 6560
rect 230 6495 350 6530
rect 230 6465 275 6495
rect 305 6465 350 6495
rect 230 6210 350 6465
rect 580 9635 700 9650
rect 580 9605 625 9635
rect 655 9605 700 9635
rect 580 9570 700 9605
rect 580 9540 625 9570
rect 655 9540 700 9570
rect 580 9500 700 9540
rect 580 9470 625 9500
rect 655 9470 700 9500
rect 580 9430 700 9470
rect 580 9400 625 9430
rect 655 9400 700 9430
rect 580 9360 700 9400
rect 580 9330 625 9360
rect 655 9330 700 9360
rect 580 9295 700 9330
rect 580 9265 625 9295
rect 655 9265 700 9295
rect 580 9235 700 9265
rect 580 9205 625 9235
rect 655 9205 700 9235
rect 580 9170 700 9205
rect 580 9140 625 9170
rect 655 9140 700 9170
rect 580 9100 700 9140
rect 580 9070 625 9100
rect 655 9070 700 9100
rect 580 9030 700 9070
rect 580 9000 625 9030
rect 655 9000 700 9030
rect 580 8960 700 9000
rect 580 8930 625 8960
rect 655 8930 700 8960
rect 580 8895 700 8930
rect 580 8865 625 8895
rect 655 8865 700 8895
rect 580 8835 700 8865
rect 580 8805 625 8835
rect 655 8805 700 8835
rect 580 8770 700 8805
rect 580 8740 625 8770
rect 655 8740 700 8770
rect 580 8700 700 8740
rect 580 8670 625 8700
rect 655 8670 700 8700
rect 580 8630 700 8670
rect 580 8600 625 8630
rect 655 8600 700 8630
rect 580 8560 700 8600
rect 580 8530 625 8560
rect 655 8530 700 8560
rect 580 8495 700 8530
rect 580 8465 625 8495
rect 655 8465 700 8495
rect 580 8435 700 8465
rect 580 8405 625 8435
rect 655 8405 700 8435
rect 580 8370 700 8405
rect 580 8340 625 8370
rect 655 8340 700 8370
rect 580 8300 700 8340
rect 580 8270 625 8300
rect 655 8270 700 8300
rect 580 8230 700 8270
rect 580 8200 625 8230
rect 655 8200 700 8230
rect 580 8160 700 8200
rect 580 8130 625 8160
rect 655 8130 700 8160
rect 580 8095 700 8130
rect 580 8065 625 8095
rect 655 8065 700 8095
rect 580 8035 700 8065
rect 580 8005 625 8035
rect 655 8005 700 8035
rect 580 7970 700 8005
rect 580 7940 625 7970
rect 655 7940 700 7970
rect 580 7900 700 7940
rect 580 7870 625 7900
rect 655 7870 700 7900
rect 580 7830 700 7870
rect 580 7800 625 7830
rect 655 7800 700 7830
rect 580 7760 700 7800
rect 580 7730 625 7760
rect 655 7730 700 7760
rect 580 7695 700 7730
rect 580 7665 625 7695
rect 655 7665 700 7695
rect 580 7635 700 7665
rect 580 7605 625 7635
rect 655 7605 700 7635
rect 580 7570 700 7605
rect 580 7540 625 7570
rect 655 7540 700 7570
rect 580 7500 700 7540
rect 580 7470 625 7500
rect 655 7470 700 7500
rect 580 7430 700 7470
rect 580 7400 625 7430
rect 655 7400 700 7430
rect 580 7360 700 7400
rect 580 7330 625 7360
rect 655 7330 700 7360
rect 580 7295 700 7330
rect 580 7265 625 7295
rect 655 7265 700 7295
rect 580 7235 700 7265
rect 580 7205 625 7235
rect 655 7205 700 7235
rect 580 7170 700 7205
rect 580 7140 625 7170
rect 655 7140 700 7170
rect 580 7100 700 7140
rect 580 7070 625 7100
rect 655 7070 700 7100
rect 580 7030 700 7070
rect 580 7000 625 7030
rect 655 7000 700 7030
rect 580 6960 700 7000
rect 580 6930 625 6960
rect 655 6930 700 6960
rect 580 6895 700 6930
rect 580 6865 625 6895
rect 655 6865 700 6895
rect 580 6835 700 6865
rect 580 6805 625 6835
rect 655 6805 700 6835
rect 580 6770 700 6805
rect 580 6740 625 6770
rect 655 6740 700 6770
rect 580 6700 700 6740
rect 580 6670 625 6700
rect 655 6670 700 6700
rect 580 6630 700 6670
rect 580 6600 625 6630
rect 655 6600 700 6630
rect 580 6560 700 6600
rect 580 6530 625 6560
rect 655 6530 700 6560
rect 580 6495 700 6530
rect 580 6465 625 6495
rect 655 6465 700 6495
rect 580 6210 700 6465
rect 930 9635 1050 9650
rect 930 9605 975 9635
rect 1005 9605 1050 9635
rect 930 9570 1050 9605
rect 930 9540 975 9570
rect 1005 9540 1050 9570
rect 930 9500 1050 9540
rect 930 9470 975 9500
rect 1005 9470 1050 9500
rect 930 9430 1050 9470
rect 930 9400 975 9430
rect 1005 9400 1050 9430
rect 930 9360 1050 9400
rect 930 9330 975 9360
rect 1005 9330 1050 9360
rect 930 9295 1050 9330
rect 930 9265 975 9295
rect 1005 9265 1050 9295
rect 930 9235 1050 9265
rect 930 9205 975 9235
rect 1005 9205 1050 9235
rect 930 9170 1050 9205
rect 930 9140 975 9170
rect 1005 9140 1050 9170
rect 930 9100 1050 9140
rect 930 9070 975 9100
rect 1005 9070 1050 9100
rect 930 9030 1050 9070
rect 930 9000 975 9030
rect 1005 9000 1050 9030
rect 930 8960 1050 9000
rect 930 8930 975 8960
rect 1005 8930 1050 8960
rect 930 8895 1050 8930
rect 930 8865 975 8895
rect 1005 8865 1050 8895
rect 930 8835 1050 8865
rect 930 8805 975 8835
rect 1005 8805 1050 8835
rect 930 8770 1050 8805
rect 930 8740 975 8770
rect 1005 8740 1050 8770
rect 930 8700 1050 8740
rect 930 8670 975 8700
rect 1005 8670 1050 8700
rect 930 8630 1050 8670
rect 930 8600 975 8630
rect 1005 8600 1050 8630
rect 930 8560 1050 8600
rect 930 8530 975 8560
rect 1005 8530 1050 8560
rect 930 8495 1050 8530
rect 930 8465 975 8495
rect 1005 8465 1050 8495
rect 930 8435 1050 8465
rect 930 8405 975 8435
rect 1005 8405 1050 8435
rect 930 8370 1050 8405
rect 930 8340 975 8370
rect 1005 8340 1050 8370
rect 930 8300 1050 8340
rect 930 8270 975 8300
rect 1005 8270 1050 8300
rect 930 8230 1050 8270
rect 930 8200 975 8230
rect 1005 8200 1050 8230
rect 930 8160 1050 8200
rect 930 8130 975 8160
rect 1005 8130 1050 8160
rect 930 8095 1050 8130
rect 930 8065 975 8095
rect 1005 8065 1050 8095
rect 930 8035 1050 8065
rect 930 8005 975 8035
rect 1005 8005 1050 8035
rect 930 7970 1050 8005
rect 930 7940 975 7970
rect 1005 7940 1050 7970
rect 930 7900 1050 7940
rect 930 7870 975 7900
rect 1005 7870 1050 7900
rect 930 7830 1050 7870
rect 930 7800 975 7830
rect 1005 7800 1050 7830
rect 930 7760 1050 7800
rect 930 7730 975 7760
rect 1005 7730 1050 7760
rect 930 7695 1050 7730
rect 930 7665 975 7695
rect 1005 7665 1050 7695
rect 930 7635 1050 7665
rect 930 7605 975 7635
rect 1005 7605 1050 7635
rect 930 7570 1050 7605
rect 930 7540 975 7570
rect 1005 7540 1050 7570
rect 930 7500 1050 7540
rect 930 7470 975 7500
rect 1005 7470 1050 7500
rect 930 7430 1050 7470
rect 930 7400 975 7430
rect 1005 7400 1050 7430
rect 930 7360 1050 7400
rect 930 7330 975 7360
rect 1005 7330 1050 7360
rect 930 7295 1050 7330
rect 930 7265 975 7295
rect 1005 7265 1050 7295
rect 930 7235 1050 7265
rect 930 7205 975 7235
rect 1005 7205 1050 7235
rect 930 7170 1050 7205
rect 930 7140 975 7170
rect 1005 7140 1050 7170
rect 930 7100 1050 7140
rect 930 7070 975 7100
rect 1005 7070 1050 7100
rect 930 7030 1050 7070
rect 930 7000 975 7030
rect 1005 7000 1050 7030
rect 930 6960 1050 7000
rect 930 6930 975 6960
rect 1005 6930 1050 6960
rect 930 6895 1050 6930
rect 930 6865 975 6895
rect 1005 6865 1050 6895
rect 930 6835 1050 6865
rect 930 6805 975 6835
rect 1005 6805 1050 6835
rect 930 6770 1050 6805
rect 930 6740 975 6770
rect 1005 6740 1050 6770
rect 930 6700 1050 6740
rect 930 6670 975 6700
rect 1005 6670 1050 6700
rect 930 6630 1050 6670
rect 930 6600 975 6630
rect 1005 6600 1050 6630
rect 930 6560 1050 6600
rect 930 6530 975 6560
rect 1005 6530 1050 6560
rect 930 6495 1050 6530
rect 930 6465 975 6495
rect 1005 6465 1050 6495
rect 930 6210 1050 6465
rect 1630 9635 1750 9650
rect 1630 9605 1675 9635
rect 1705 9605 1750 9635
rect 1630 9570 1750 9605
rect 1630 9540 1675 9570
rect 1705 9540 1750 9570
rect 1630 9500 1750 9540
rect 1630 9470 1675 9500
rect 1705 9470 1750 9500
rect 1630 9430 1750 9470
rect 1630 9400 1675 9430
rect 1705 9400 1750 9430
rect 1630 9360 1750 9400
rect 1630 9330 1675 9360
rect 1705 9330 1750 9360
rect 1630 9295 1750 9330
rect 1630 9265 1675 9295
rect 1705 9265 1750 9295
rect 1630 9235 1750 9265
rect 1630 9205 1675 9235
rect 1705 9205 1750 9235
rect 1630 9170 1750 9205
rect 1630 9140 1675 9170
rect 1705 9140 1750 9170
rect 1630 9100 1750 9140
rect 1630 9070 1675 9100
rect 1705 9070 1750 9100
rect 1630 9030 1750 9070
rect 1630 9000 1675 9030
rect 1705 9000 1750 9030
rect 1630 8960 1750 9000
rect 1630 8930 1675 8960
rect 1705 8930 1750 8960
rect 1630 8895 1750 8930
rect 1630 8865 1675 8895
rect 1705 8865 1750 8895
rect 1630 8835 1750 8865
rect 1630 8805 1675 8835
rect 1705 8805 1750 8835
rect 1630 8770 1750 8805
rect 1630 8740 1675 8770
rect 1705 8740 1750 8770
rect 1630 8700 1750 8740
rect 1630 8670 1675 8700
rect 1705 8670 1750 8700
rect 1630 8630 1750 8670
rect 1630 8600 1675 8630
rect 1705 8600 1750 8630
rect 1630 8560 1750 8600
rect 1630 8530 1675 8560
rect 1705 8530 1750 8560
rect 1630 8495 1750 8530
rect 1630 8465 1675 8495
rect 1705 8465 1750 8495
rect 1630 8435 1750 8465
rect 1630 8405 1675 8435
rect 1705 8405 1750 8435
rect 1630 8370 1750 8405
rect 1630 8340 1675 8370
rect 1705 8340 1750 8370
rect 1630 8300 1750 8340
rect 1630 8270 1675 8300
rect 1705 8270 1750 8300
rect 1630 8230 1750 8270
rect 1630 8200 1675 8230
rect 1705 8200 1750 8230
rect 1630 8160 1750 8200
rect 1630 8130 1675 8160
rect 1705 8130 1750 8160
rect 1630 8095 1750 8130
rect 1630 8065 1675 8095
rect 1705 8065 1750 8095
rect 1630 8035 1750 8065
rect 1630 8005 1675 8035
rect 1705 8005 1750 8035
rect 1630 7970 1750 8005
rect 1630 7940 1675 7970
rect 1705 7940 1750 7970
rect 1630 7900 1750 7940
rect 1630 7870 1675 7900
rect 1705 7870 1750 7900
rect 1630 7830 1750 7870
rect 1630 7800 1675 7830
rect 1705 7800 1750 7830
rect 1630 7760 1750 7800
rect 1630 7730 1675 7760
rect 1705 7730 1750 7760
rect 1630 7695 1750 7730
rect 1630 7665 1675 7695
rect 1705 7665 1750 7695
rect 1630 7635 1750 7665
rect 1630 7605 1675 7635
rect 1705 7605 1750 7635
rect 1630 7570 1750 7605
rect 1630 7540 1675 7570
rect 1705 7540 1750 7570
rect 1630 7500 1750 7540
rect 1630 7470 1675 7500
rect 1705 7470 1750 7500
rect 1630 7430 1750 7470
rect 1630 7400 1675 7430
rect 1705 7400 1750 7430
rect 1630 7360 1750 7400
rect 1630 7330 1675 7360
rect 1705 7330 1750 7360
rect 1630 7295 1750 7330
rect 1630 7265 1675 7295
rect 1705 7265 1750 7295
rect 1630 7235 1750 7265
rect 1630 7205 1675 7235
rect 1705 7205 1750 7235
rect 1630 7170 1750 7205
rect 1630 7140 1675 7170
rect 1705 7140 1750 7170
rect 1630 7100 1750 7140
rect 1630 7070 1675 7100
rect 1705 7070 1750 7100
rect 1630 7030 1750 7070
rect 1630 7000 1675 7030
rect 1705 7000 1750 7030
rect 1630 6960 1750 7000
rect 1630 6930 1675 6960
rect 1705 6930 1750 6960
rect 1630 6895 1750 6930
rect 1630 6865 1675 6895
rect 1705 6865 1750 6895
rect 1630 6835 1750 6865
rect 1630 6805 1675 6835
rect 1705 6805 1750 6835
rect 1630 6770 1750 6805
rect 1630 6740 1675 6770
rect 1705 6740 1750 6770
rect 1630 6700 1750 6740
rect 1630 6670 1675 6700
rect 1705 6670 1750 6700
rect 1630 6630 1750 6670
rect 1630 6600 1675 6630
rect 1705 6600 1750 6630
rect 1630 6560 1750 6600
rect 1630 6530 1675 6560
rect 1705 6530 1750 6560
rect 1630 6495 1750 6530
rect 1630 6465 1675 6495
rect 1705 6465 1750 6495
rect 1630 6210 1750 6465
rect 2285 9635 2405 15895
rect 2650 15665 2670 15745
rect 2970 15740 3010 15745
rect 2970 15710 2975 15740
rect 3005 15710 3010 15740
rect 2970 15700 3010 15710
rect 2970 15670 2975 15700
rect 3005 15670 3010 15700
rect 2970 15665 3010 15670
rect 3295 15740 3335 15745
rect 3295 15710 3300 15740
rect 3330 15710 3335 15740
rect 3295 15700 3335 15710
rect 3295 15670 3300 15700
rect 3330 15670 3335 15700
rect 6620 15705 6740 17725
rect 6620 15675 6625 15705
rect 6655 15675 6665 15705
rect 6695 15675 6705 15705
rect 6735 15675 6740 15705
rect 3295 15665 3335 15670
rect 5645 15665 5685 15670
rect 5645 15635 5650 15665
rect 5680 15635 5685 15665
rect 5645 15625 5685 15635
rect 5645 15595 5650 15625
rect 5680 15595 5685 15625
rect 5645 15590 5685 15595
rect 5970 15665 6010 15670
rect 5970 15635 5975 15665
rect 6005 15635 6010 15665
rect 5970 15625 6010 15635
rect 5970 15595 5975 15625
rect 6005 15595 6010 15625
rect 5970 15590 6010 15595
rect 6310 15590 6330 15670
rect 6440 15590 6460 15670
rect 6535 15590 6555 15670
rect 6620 15665 6740 15675
rect 6620 15635 6625 15665
rect 6655 15635 6665 15665
rect 6695 15635 6705 15665
rect 6735 15635 6740 15665
rect 6620 15625 6740 15635
rect 6620 15595 6625 15625
rect 6655 15595 6665 15625
rect 6695 15595 6705 15625
rect 6735 15595 6740 15625
rect 6620 13005 6740 15595
rect 6620 12975 6625 13005
rect 6655 12975 6665 13005
rect 6695 12975 6705 13005
rect 6735 12975 6740 13005
rect 6620 12965 6740 12975
rect 6620 12935 6625 12965
rect 6655 12935 6665 12965
rect 6695 12935 6705 12965
rect 6735 12935 6740 12965
rect 6620 12925 6740 12935
rect 6620 12895 6625 12925
rect 6655 12895 6665 12925
rect 6695 12895 6705 12925
rect 6735 12895 6740 12925
rect 6620 12890 6740 12895
rect 6590 12160 6710 12165
rect 6590 12130 6595 12160
rect 6625 12130 6635 12160
rect 6665 12130 6675 12160
rect 6705 12130 6710 12160
rect 6590 12120 6710 12130
rect 6590 12090 6595 12120
rect 6625 12090 6635 12120
rect 6665 12090 6675 12120
rect 6705 12090 6710 12120
rect 6590 12080 6710 12090
rect 6590 12050 6595 12080
rect 6625 12050 6635 12080
rect 6665 12050 6675 12080
rect 6705 12050 6710 12080
rect 6590 11205 6710 12050
rect 6590 11175 6595 11205
rect 6625 11175 6635 11205
rect 6665 11175 6675 11205
rect 6705 11175 6710 11205
rect 6590 11165 6710 11175
rect 6590 11135 6595 11165
rect 6625 11135 6635 11165
rect 6665 11135 6675 11165
rect 6705 11135 6710 11165
rect 6590 11125 6710 11135
rect 6590 11095 6595 11125
rect 6625 11095 6635 11125
rect 6665 11095 6675 11125
rect 6705 11095 6710 11125
rect 2285 9605 2330 9635
rect 2360 9605 2405 9635
rect 2285 9570 2405 9605
rect 2285 9540 2330 9570
rect 2360 9540 2405 9570
rect 2285 9500 2405 9540
rect 2285 9470 2330 9500
rect 2360 9470 2405 9500
rect 2285 9430 2405 9470
rect 2285 9400 2330 9430
rect 2360 9400 2405 9430
rect 2285 9360 2405 9400
rect 2285 9330 2330 9360
rect 2360 9330 2405 9360
rect 2285 9295 2405 9330
rect 2285 9265 2330 9295
rect 2360 9265 2405 9295
rect 2285 9235 2405 9265
rect 2285 9205 2330 9235
rect 2360 9205 2405 9235
rect 2285 9170 2405 9205
rect 2285 9140 2330 9170
rect 2360 9140 2405 9170
rect 2285 9100 2405 9140
rect 2285 9070 2330 9100
rect 2360 9070 2405 9100
rect 2285 9030 2405 9070
rect 2285 9000 2330 9030
rect 2360 9000 2405 9030
rect 2285 8960 2405 9000
rect 2285 8930 2330 8960
rect 2360 8930 2405 8960
rect 2285 8895 2405 8930
rect 2285 8865 2330 8895
rect 2360 8865 2405 8895
rect 2285 8835 2405 8865
rect 2285 8805 2330 8835
rect 2360 8805 2405 8835
rect 2285 8770 2405 8805
rect 2285 8740 2330 8770
rect 2360 8740 2405 8770
rect 2285 8700 2405 8740
rect 2285 8670 2330 8700
rect 2360 8670 2405 8700
rect 2285 8630 2405 8670
rect 2285 8600 2330 8630
rect 2360 8600 2405 8630
rect 2285 8560 2405 8600
rect 2285 8530 2330 8560
rect 2360 8530 2405 8560
rect 2285 8495 2405 8530
rect 2285 8465 2330 8495
rect 2360 8465 2405 8495
rect 2285 8435 2405 8465
rect 2285 8405 2330 8435
rect 2360 8405 2405 8435
rect 2285 8370 2405 8405
rect 2285 8340 2330 8370
rect 2360 8340 2405 8370
rect 2285 8300 2405 8340
rect 2285 8270 2330 8300
rect 2360 8270 2405 8300
rect 2285 8230 2405 8270
rect 2285 8200 2330 8230
rect 2360 8200 2405 8230
rect 2285 8160 2405 8200
rect 2285 8130 2330 8160
rect 2360 8130 2405 8160
rect 2285 8095 2405 8130
rect 2285 8065 2330 8095
rect 2360 8065 2405 8095
rect 2285 8035 2405 8065
rect 2285 8005 2330 8035
rect 2360 8005 2405 8035
rect 2285 7970 2405 8005
rect 2285 7940 2330 7970
rect 2360 7940 2405 7970
rect 2285 7900 2405 7940
rect 2285 7870 2330 7900
rect 2360 7870 2405 7900
rect 2285 7830 2405 7870
rect 2285 7800 2330 7830
rect 2360 7800 2405 7830
rect 2285 7760 2405 7800
rect 2285 7730 2330 7760
rect 2360 7730 2405 7760
rect 2285 7695 2405 7730
rect 2285 7665 2330 7695
rect 2360 7665 2405 7695
rect 2285 7635 2405 7665
rect 2285 7605 2330 7635
rect 2360 7605 2405 7635
rect 2285 7570 2405 7605
rect 2285 7540 2330 7570
rect 2360 7540 2405 7570
rect 2285 7500 2405 7540
rect 2285 7470 2330 7500
rect 2360 7470 2405 7500
rect 2285 7430 2405 7470
rect 2285 7400 2330 7430
rect 2360 7400 2405 7430
rect 2285 7360 2405 7400
rect 2285 7330 2330 7360
rect 2360 7330 2405 7360
rect 2285 7295 2405 7330
rect 2285 7265 2330 7295
rect 2360 7265 2405 7295
rect 2285 7235 2405 7265
rect 2285 7205 2330 7235
rect 2360 7205 2405 7235
rect 2285 7170 2405 7205
rect 2285 7140 2330 7170
rect 2360 7140 2405 7170
rect 2285 7100 2405 7140
rect 2285 7070 2330 7100
rect 2360 7070 2405 7100
rect 2285 7030 2405 7070
rect 2285 7000 2330 7030
rect 2360 7000 2405 7030
rect 2285 6960 2405 7000
rect 2285 6930 2330 6960
rect 2360 6930 2405 6960
rect 2285 6895 2405 6930
rect 2285 6865 2330 6895
rect 2360 6865 2405 6895
rect 2285 6835 2405 6865
rect 2285 6805 2330 6835
rect 2360 6805 2405 6835
rect 2285 6770 2405 6805
rect 2285 6740 2330 6770
rect 2360 6740 2405 6770
rect 2285 6700 2405 6740
rect 2285 6670 2330 6700
rect 2360 6670 2405 6700
rect 2285 6630 2405 6670
rect 2285 6600 2330 6630
rect 2360 6600 2405 6630
rect 2285 6560 2405 6600
rect 2285 6530 2330 6560
rect 2360 6530 2405 6560
rect 2285 6495 2405 6530
rect 2285 6465 2330 6495
rect 2360 6465 2405 6495
rect 2285 6450 2405 6465
rect 2485 6435 2505 9690
rect 2045 6430 2085 6435
rect 2045 6400 2050 6430
rect 2080 6400 2085 6430
rect 2045 6395 2085 6400
rect 2475 6430 2515 6435
rect 2475 6400 2480 6430
rect 2510 6400 2515 6430
rect 2475 6395 2515 6400
rect 2000 6375 2040 6380
rect 2000 6345 2005 6375
rect 2035 6345 2040 6375
rect 2000 6340 2040 6345
rect 1280 6205 1400 6210
rect 1280 6175 1285 6205
rect 1315 6175 1325 6205
rect 1355 6175 1365 6205
rect 1395 6175 1400 6205
rect 1280 6165 1400 6175
rect 1280 6135 1285 6165
rect 1315 6135 1325 6165
rect 1355 6135 1365 6165
rect 1395 6135 1400 6165
rect 1280 6125 1400 6135
rect 1280 6095 1285 6125
rect 1315 6095 1325 6125
rect 1355 6095 1365 6125
rect 1395 6095 1400 6125
rect 1280 850 1400 6095
rect 2010 1955 2030 6340
rect 2055 2010 2075 6395
rect 2725 6335 2745 9690
rect 2855 6435 2875 9690
rect 2845 6430 2885 6435
rect 2845 6400 2850 6430
rect 2880 6400 2885 6430
rect 2845 6395 2885 6400
rect 2715 6330 2755 6335
rect 2715 6300 2720 6330
rect 2750 6300 2755 6330
rect 2715 6295 2755 6300
rect 3000 6280 3020 10735
rect 6590 10500 6710 11095
rect 6590 10470 6595 10500
rect 6625 10470 6635 10500
rect 6665 10470 6675 10500
rect 6705 10470 6710 10500
rect 6590 10460 6710 10470
rect 6590 10430 6595 10460
rect 6625 10430 6635 10460
rect 6665 10430 6675 10460
rect 6705 10430 6710 10460
rect 6590 10420 6710 10430
rect 6590 10390 6595 10420
rect 6625 10390 6635 10420
rect 6665 10390 6675 10420
rect 6705 10390 6710 10420
rect 3175 9650 3215 10385
rect 3235 9650 3275 10385
rect 3345 9650 3385 10385
rect 6590 10035 6710 10390
rect 6590 10005 6595 10035
rect 6625 10005 6635 10035
rect 6665 10005 6675 10035
rect 6705 10005 6710 10035
rect 6590 9995 6710 10005
rect 6590 9965 6595 9995
rect 6625 9965 6635 9995
rect 6665 9965 6675 9995
rect 6705 9965 6710 9995
rect 6590 9955 6710 9965
rect 6590 9925 6595 9955
rect 6625 9925 6635 9955
rect 6665 9925 6675 9955
rect 6705 9925 6710 9955
rect 3165 9635 3285 9650
rect 3165 9605 3180 9635
rect 3210 9605 3240 9635
rect 3270 9605 3285 9635
rect 3165 9570 3285 9605
rect 3165 9540 3180 9570
rect 3210 9540 3240 9570
rect 3270 9540 3285 9570
rect 3165 9500 3285 9540
rect 3165 9470 3180 9500
rect 3210 9470 3240 9500
rect 3270 9470 3285 9500
rect 3165 9430 3285 9470
rect 3165 9400 3180 9430
rect 3210 9400 3240 9430
rect 3270 9400 3285 9430
rect 3165 9360 3285 9400
rect 3165 9330 3180 9360
rect 3210 9330 3240 9360
rect 3270 9330 3285 9360
rect 3165 9295 3285 9330
rect 3165 9265 3180 9295
rect 3210 9265 3240 9295
rect 3270 9265 3285 9295
rect 3165 9235 3285 9265
rect 3165 9205 3180 9235
rect 3210 9205 3240 9235
rect 3270 9205 3285 9235
rect 3165 9170 3285 9205
rect 3165 9140 3180 9170
rect 3210 9140 3240 9170
rect 3270 9140 3285 9170
rect 3165 9100 3285 9140
rect 3165 9070 3180 9100
rect 3210 9070 3240 9100
rect 3270 9070 3285 9100
rect 3165 9030 3285 9070
rect 3165 9000 3180 9030
rect 3210 9000 3240 9030
rect 3270 9000 3285 9030
rect 3165 8960 3285 9000
rect 3165 8930 3180 8960
rect 3210 8930 3240 8960
rect 3270 8930 3285 8960
rect 3165 8895 3285 8930
rect 3165 8865 3180 8895
rect 3210 8865 3240 8895
rect 3270 8865 3285 8895
rect 3165 8835 3285 8865
rect 3165 8805 3180 8835
rect 3210 8805 3240 8835
rect 3270 8805 3285 8835
rect 3165 8770 3285 8805
rect 3165 8740 3180 8770
rect 3210 8740 3240 8770
rect 3270 8740 3285 8770
rect 3165 8700 3285 8740
rect 3165 8670 3180 8700
rect 3210 8670 3240 8700
rect 3270 8670 3285 8700
rect 3165 8630 3285 8670
rect 3165 8600 3180 8630
rect 3210 8600 3240 8630
rect 3270 8600 3285 8630
rect 3165 8560 3285 8600
rect 3165 8530 3180 8560
rect 3210 8530 3240 8560
rect 3270 8530 3285 8560
rect 3165 8495 3285 8530
rect 3165 8465 3180 8495
rect 3210 8465 3240 8495
rect 3270 8465 3285 8495
rect 3165 8435 3285 8465
rect 3165 8405 3180 8435
rect 3210 8405 3240 8435
rect 3270 8405 3285 8435
rect 3165 8370 3285 8405
rect 3165 8340 3180 8370
rect 3210 8340 3240 8370
rect 3270 8340 3285 8370
rect 3165 8300 3285 8340
rect 3165 8270 3180 8300
rect 3210 8270 3240 8300
rect 3270 8270 3285 8300
rect 3165 8230 3285 8270
rect 3165 8200 3180 8230
rect 3210 8200 3240 8230
rect 3270 8200 3285 8230
rect 3165 8160 3285 8200
rect 3165 8130 3180 8160
rect 3210 8130 3240 8160
rect 3270 8130 3285 8160
rect 3165 8095 3285 8130
rect 3165 8065 3180 8095
rect 3210 8065 3240 8095
rect 3270 8065 3285 8095
rect 3165 8035 3285 8065
rect 3165 8005 3180 8035
rect 3210 8005 3240 8035
rect 3270 8005 3285 8035
rect 3165 7970 3285 8005
rect 3165 7940 3180 7970
rect 3210 7940 3240 7970
rect 3270 7940 3285 7970
rect 3165 7900 3285 7940
rect 3165 7870 3180 7900
rect 3210 7870 3240 7900
rect 3270 7870 3285 7900
rect 3165 7830 3285 7870
rect 3165 7800 3180 7830
rect 3210 7800 3240 7830
rect 3270 7800 3285 7830
rect 3165 7760 3285 7800
rect 3165 7730 3180 7760
rect 3210 7730 3240 7760
rect 3270 7730 3285 7760
rect 3165 7695 3285 7730
rect 3165 7665 3180 7695
rect 3210 7665 3240 7695
rect 3270 7665 3285 7695
rect 3165 7635 3285 7665
rect 3165 7605 3180 7635
rect 3210 7605 3240 7635
rect 3270 7605 3285 7635
rect 3165 7570 3285 7605
rect 3165 7540 3180 7570
rect 3210 7540 3240 7570
rect 3270 7540 3285 7570
rect 3165 7500 3285 7540
rect 3165 7470 3180 7500
rect 3210 7470 3240 7500
rect 3270 7470 3285 7500
rect 3165 7430 3285 7470
rect 3165 7400 3180 7430
rect 3210 7400 3240 7430
rect 3270 7400 3285 7430
rect 3165 7360 3285 7400
rect 3165 7330 3180 7360
rect 3210 7330 3240 7360
rect 3270 7330 3285 7360
rect 3165 7295 3285 7330
rect 3165 7265 3180 7295
rect 3210 7265 3240 7295
rect 3270 7265 3285 7295
rect 3165 7235 3285 7265
rect 3165 7205 3180 7235
rect 3210 7205 3240 7235
rect 3270 7205 3285 7235
rect 3165 7170 3285 7205
rect 3165 7140 3180 7170
rect 3210 7140 3240 7170
rect 3270 7140 3285 7170
rect 3165 7100 3285 7140
rect 3165 7070 3180 7100
rect 3210 7070 3240 7100
rect 3270 7070 3285 7100
rect 3165 7030 3285 7070
rect 3165 7000 3180 7030
rect 3210 7000 3240 7030
rect 3270 7000 3285 7030
rect 3165 6960 3285 7000
rect 3165 6930 3180 6960
rect 3210 6930 3240 6960
rect 3270 6930 3285 6960
rect 3165 6895 3285 6930
rect 3165 6865 3180 6895
rect 3210 6865 3240 6895
rect 3270 6865 3285 6895
rect 3165 6835 3285 6865
rect 3165 6805 3180 6835
rect 3210 6805 3240 6835
rect 3270 6805 3285 6835
rect 3165 6770 3285 6805
rect 3165 6740 3180 6770
rect 3210 6740 3240 6770
rect 3270 6740 3285 6770
rect 3165 6700 3285 6740
rect 3165 6670 3180 6700
rect 3210 6670 3240 6700
rect 3270 6670 3285 6700
rect 3165 6630 3285 6670
rect 3165 6600 3180 6630
rect 3210 6600 3240 6630
rect 3270 6600 3285 6630
rect 3165 6560 3285 6600
rect 3165 6530 3180 6560
rect 3210 6530 3240 6560
rect 3270 6530 3285 6560
rect 3165 6495 3285 6530
rect 3165 6465 3180 6495
rect 3210 6465 3240 6495
rect 3270 6465 3285 6495
rect 3165 6450 3285 6465
rect 3335 9635 3395 9650
rect 3335 9605 3350 9635
rect 3380 9605 3395 9635
rect 3335 9570 3395 9605
rect 3335 9540 3350 9570
rect 3380 9540 3395 9570
rect 3335 9500 3395 9540
rect 3335 9470 3350 9500
rect 3380 9470 3395 9500
rect 3335 9430 3395 9470
rect 3335 9400 3350 9430
rect 3380 9400 3395 9430
rect 3335 9360 3395 9400
rect 3335 9330 3350 9360
rect 3380 9330 3395 9360
rect 3335 9295 3395 9330
rect 3335 9265 3350 9295
rect 3380 9265 3395 9295
rect 3335 9235 3395 9265
rect 3335 9205 3350 9235
rect 3380 9205 3395 9235
rect 3335 9170 3395 9205
rect 3335 9140 3350 9170
rect 3380 9140 3395 9170
rect 3335 9100 3395 9140
rect 3335 9070 3350 9100
rect 3380 9070 3395 9100
rect 3335 9030 3395 9070
rect 3335 9000 3350 9030
rect 3380 9000 3395 9030
rect 3335 8960 3395 9000
rect 3335 8930 3350 8960
rect 3380 8930 3395 8960
rect 3335 8895 3395 8930
rect 3335 8865 3350 8895
rect 3380 8865 3395 8895
rect 3335 8835 3395 8865
rect 3335 8805 3350 8835
rect 3380 8805 3395 8835
rect 3335 8770 3395 8805
rect 3335 8740 3350 8770
rect 3380 8740 3395 8770
rect 3335 8700 3395 8740
rect 3335 8670 3350 8700
rect 3380 8670 3395 8700
rect 3335 8630 3395 8670
rect 3335 8600 3350 8630
rect 3380 8600 3395 8630
rect 3335 8560 3395 8600
rect 3335 8530 3350 8560
rect 3380 8530 3395 8560
rect 3335 8495 3395 8530
rect 3335 8465 3350 8495
rect 3380 8465 3395 8495
rect 3335 8435 3395 8465
rect 3335 8405 3350 8435
rect 3380 8405 3395 8435
rect 3335 8370 3395 8405
rect 3335 8340 3350 8370
rect 3380 8340 3395 8370
rect 3335 8300 3395 8340
rect 3335 8270 3350 8300
rect 3380 8270 3395 8300
rect 3335 8230 3395 8270
rect 3335 8200 3350 8230
rect 3380 8200 3395 8230
rect 3335 8160 3395 8200
rect 3335 8130 3350 8160
rect 3380 8130 3395 8160
rect 3335 8095 3395 8130
rect 3335 8065 3350 8095
rect 3380 8065 3395 8095
rect 3335 8035 3395 8065
rect 3335 8005 3350 8035
rect 3380 8005 3395 8035
rect 3335 7970 3395 8005
rect 3335 7940 3350 7970
rect 3380 7940 3395 7970
rect 3335 7900 3395 7940
rect 3335 7870 3350 7900
rect 3380 7870 3395 7900
rect 3335 7830 3395 7870
rect 3335 7800 3350 7830
rect 3380 7800 3395 7830
rect 3335 7760 3395 7800
rect 3335 7730 3350 7760
rect 3380 7730 3395 7760
rect 3335 7695 3395 7730
rect 3335 7665 3350 7695
rect 3380 7665 3395 7695
rect 3335 7635 3395 7665
rect 3335 7605 3350 7635
rect 3380 7605 3395 7635
rect 3335 7570 3395 7605
rect 3335 7540 3350 7570
rect 3380 7540 3395 7570
rect 3335 7500 3395 7540
rect 3335 7470 3350 7500
rect 3380 7470 3395 7500
rect 3335 7430 3395 7470
rect 3335 7400 3350 7430
rect 3380 7400 3395 7430
rect 3335 7360 3395 7400
rect 3335 7330 3350 7360
rect 3380 7330 3395 7360
rect 3335 7295 3395 7330
rect 3335 7265 3350 7295
rect 3380 7265 3395 7295
rect 3335 7235 3395 7265
rect 3335 7205 3350 7235
rect 3380 7205 3395 7235
rect 3335 7170 3395 7205
rect 3335 7140 3350 7170
rect 3380 7140 3395 7170
rect 3335 7100 3395 7140
rect 3335 7070 3350 7100
rect 3380 7070 3395 7100
rect 3335 7030 3395 7070
rect 3335 7000 3350 7030
rect 3380 7000 3395 7030
rect 3640 7010 3660 9690
rect 3335 6960 3395 7000
rect 3335 6930 3350 6960
rect 3380 6930 3395 6960
rect 3335 6895 3395 6930
rect 3335 6865 3350 6895
rect 3380 6865 3395 6895
rect 3335 6835 3395 6865
rect 3335 6805 3350 6835
rect 3380 6805 3395 6835
rect 3335 6770 3395 6805
rect 3335 6740 3350 6770
rect 3380 6740 3395 6770
rect 3335 6700 3395 6740
rect 3335 6670 3350 6700
rect 3380 6670 3395 6700
rect 3335 6630 3395 6670
rect 3335 6600 3350 6630
rect 3380 6600 3395 6630
rect 3335 6560 3395 6600
rect 3335 6530 3350 6560
rect 3380 6530 3395 6560
rect 3335 6495 3395 6530
rect 3335 6465 3350 6495
rect 3380 6465 3395 6495
rect 3335 6450 3395 6465
rect 3390 6430 3430 6435
rect 3390 6400 3395 6430
rect 3425 6400 3430 6430
rect 3390 6395 3430 6400
rect 2990 6275 3030 6280
rect 2990 6245 2995 6275
rect 3025 6245 3030 6275
rect 2990 6240 3030 6245
rect 3400 2935 3420 6395
rect 3630 6375 3670 7010
rect 3630 6345 3635 6375
rect 3665 6345 3670 6375
rect 3630 6340 3670 6345
rect 4310 6205 4340 9690
rect 4310 6165 4340 6175
rect 4310 6125 4340 6135
rect 4310 6090 4340 6095
rect 4420 6205 4450 9690
rect 4420 6165 4450 6175
rect 4420 6125 4450 6135
rect 4420 6090 4450 6095
rect 4530 6205 4560 9690
rect 4530 6165 4560 6175
rect 4530 6125 4560 6135
rect 4530 6090 4560 6095
rect 4640 6205 4670 9690
rect 5320 6380 5340 9690
rect 6155 6435 6175 9690
rect 5490 6430 5530 6435
rect 5490 6400 5495 6430
rect 5525 6400 5530 6430
rect 5490 6395 5530 6400
rect 6145 6430 6185 6435
rect 6145 6400 6150 6430
rect 6180 6400 6185 6430
rect 6145 6395 6185 6400
rect 5310 6375 5350 6380
rect 5310 6345 5315 6375
rect 5345 6345 5350 6375
rect 5310 6340 5350 6345
rect 4850 6330 4890 6335
rect 4850 6300 4855 6330
rect 4885 6300 4890 6330
rect 4850 6295 4890 6300
rect 4640 6165 4670 6175
rect 4640 6125 4670 6135
rect 4640 6090 4670 6095
rect 4860 5070 4880 6295
rect 4850 5065 4890 5070
rect 4850 5035 4855 5065
rect 4885 5035 4890 5065
rect 4850 5030 4890 5035
rect 4940 5065 4980 5070
rect 4940 5035 4945 5065
rect 4975 5035 4980 5065
rect 4940 5030 4980 5035
rect 4950 4505 4970 5030
rect 4940 4500 4980 4505
rect 4940 4470 4945 4500
rect 4975 4470 4980 4500
rect 4940 4465 4980 4470
rect 5500 3005 5520 6395
rect 5545 6275 5585 6280
rect 5545 6245 5550 6275
rect 5580 6245 5585 6275
rect 5545 6240 5585 6245
rect 5490 3000 5530 3005
rect 5490 2970 5495 3000
rect 5525 2970 5530 3000
rect 5490 2965 5530 2970
rect 5555 2950 5575 6240
rect 6230 5090 6250 9690
rect 6475 6435 6500 9690
rect 6590 9635 6710 9925
rect 6590 9605 6635 9635
rect 6665 9605 6710 9635
rect 6590 9570 6710 9605
rect 6590 9540 6635 9570
rect 6665 9540 6710 9570
rect 6590 9500 6710 9540
rect 6590 9470 6635 9500
rect 6665 9470 6710 9500
rect 6590 9430 6710 9470
rect 6590 9400 6635 9430
rect 6665 9400 6710 9430
rect 6590 9360 6710 9400
rect 6590 9330 6635 9360
rect 6665 9330 6710 9360
rect 6590 9295 6710 9330
rect 6590 9265 6635 9295
rect 6665 9265 6710 9295
rect 6590 9235 6710 9265
rect 6590 9205 6635 9235
rect 6665 9205 6710 9235
rect 6590 9170 6710 9205
rect 6590 9140 6635 9170
rect 6665 9140 6710 9170
rect 6590 9100 6710 9140
rect 6590 9070 6635 9100
rect 6665 9070 6710 9100
rect 6590 9030 6710 9070
rect 6590 9000 6635 9030
rect 6665 9000 6710 9030
rect 6590 8960 6710 9000
rect 6590 8930 6635 8960
rect 6665 8930 6710 8960
rect 6590 8895 6710 8930
rect 6590 8865 6635 8895
rect 6665 8865 6710 8895
rect 6590 8835 6710 8865
rect 6590 8805 6635 8835
rect 6665 8805 6710 8835
rect 6590 8770 6710 8805
rect 6590 8740 6635 8770
rect 6665 8740 6710 8770
rect 6590 8700 6710 8740
rect 6590 8670 6635 8700
rect 6665 8670 6710 8700
rect 6590 8630 6710 8670
rect 6590 8600 6635 8630
rect 6665 8600 6710 8630
rect 6590 8560 6710 8600
rect 6590 8530 6635 8560
rect 6665 8530 6710 8560
rect 6590 8495 6710 8530
rect 6590 8465 6635 8495
rect 6665 8465 6710 8495
rect 6590 8435 6710 8465
rect 6590 8405 6635 8435
rect 6665 8405 6710 8435
rect 6590 8370 6710 8405
rect 6590 8340 6635 8370
rect 6665 8340 6710 8370
rect 6590 8300 6710 8340
rect 6590 8270 6635 8300
rect 6665 8270 6710 8300
rect 6590 8230 6710 8270
rect 6590 8200 6635 8230
rect 6665 8200 6710 8230
rect 6590 8160 6710 8200
rect 6590 8130 6635 8160
rect 6665 8130 6710 8160
rect 6590 8095 6710 8130
rect 6590 8065 6635 8095
rect 6665 8065 6710 8095
rect 6590 8035 6710 8065
rect 6590 8005 6635 8035
rect 6665 8005 6710 8035
rect 6590 7970 6710 8005
rect 6590 7940 6635 7970
rect 6665 7940 6710 7970
rect 6590 7900 6710 7940
rect 6590 7870 6635 7900
rect 6665 7870 6710 7900
rect 6590 7830 6710 7870
rect 6590 7800 6635 7830
rect 6665 7800 6710 7830
rect 6590 7760 6710 7800
rect 6590 7730 6635 7760
rect 6665 7730 6710 7760
rect 6590 7695 6710 7730
rect 6590 7665 6635 7695
rect 6665 7665 6710 7695
rect 6590 7635 6710 7665
rect 6590 7605 6635 7635
rect 6665 7605 6710 7635
rect 6590 7570 6710 7605
rect 6590 7540 6635 7570
rect 6665 7540 6710 7570
rect 6590 7500 6710 7540
rect 6590 7470 6635 7500
rect 6665 7470 6710 7500
rect 6590 7430 6710 7470
rect 6590 7400 6635 7430
rect 6665 7400 6710 7430
rect 6590 7360 6710 7400
rect 6590 7330 6635 7360
rect 6665 7330 6710 7360
rect 6590 7295 6710 7330
rect 6590 7265 6635 7295
rect 6665 7265 6710 7295
rect 6590 7235 6710 7265
rect 6590 7205 6635 7235
rect 6665 7205 6710 7235
rect 6590 7170 6710 7205
rect 6590 7140 6635 7170
rect 6665 7140 6710 7170
rect 6590 7100 6710 7140
rect 6590 7070 6635 7100
rect 6665 7070 6710 7100
rect 6590 7030 6710 7070
rect 6590 7000 6635 7030
rect 6665 7000 6710 7030
rect 6590 6960 6710 7000
rect 6590 6930 6635 6960
rect 6665 6930 6710 6960
rect 6590 6895 6710 6930
rect 6590 6865 6635 6895
rect 6665 6865 6710 6895
rect 6590 6835 6710 6865
rect 6590 6805 6635 6835
rect 6665 6805 6710 6835
rect 6590 6770 6710 6805
rect 6590 6740 6635 6770
rect 6665 6740 6710 6770
rect 6590 6700 6710 6740
rect 6590 6670 6635 6700
rect 6665 6670 6710 6700
rect 6590 6630 6710 6670
rect 6590 6600 6635 6630
rect 6665 6600 6710 6630
rect 6590 6560 6710 6600
rect 6590 6530 6635 6560
rect 6665 6530 6710 6560
rect 6590 6495 6710 6530
rect 6590 6465 6635 6495
rect 6665 6465 6710 6495
rect 6590 6450 6710 6465
rect 7230 9635 7350 9650
rect 7230 9605 7275 9635
rect 7305 9605 7350 9635
rect 7230 9570 7350 9605
rect 7230 9540 7275 9570
rect 7305 9540 7350 9570
rect 7230 9500 7350 9540
rect 7230 9470 7275 9500
rect 7305 9470 7350 9500
rect 7230 9430 7350 9470
rect 7230 9400 7275 9430
rect 7305 9400 7350 9430
rect 7230 9360 7350 9400
rect 7230 9330 7275 9360
rect 7305 9330 7350 9360
rect 7230 9295 7350 9330
rect 7230 9265 7275 9295
rect 7305 9265 7350 9295
rect 7230 9235 7350 9265
rect 7230 9205 7275 9235
rect 7305 9205 7350 9235
rect 7230 9170 7350 9205
rect 7230 9140 7275 9170
rect 7305 9140 7350 9170
rect 7230 9100 7350 9140
rect 7230 9070 7275 9100
rect 7305 9070 7350 9100
rect 7230 9030 7350 9070
rect 7230 9000 7275 9030
rect 7305 9000 7350 9030
rect 7230 8960 7350 9000
rect 7230 8930 7275 8960
rect 7305 8930 7350 8960
rect 7230 8895 7350 8930
rect 7230 8865 7275 8895
rect 7305 8865 7350 8895
rect 7230 8835 7350 8865
rect 7230 8805 7275 8835
rect 7305 8805 7350 8835
rect 7230 8770 7350 8805
rect 7230 8740 7275 8770
rect 7305 8740 7350 8770
rect 7230 8700 7350 8740
rect 7230 8670 7275 8700
rect 7305 8670 7350 8700
rect 7230 8630 7350 8670
rect 7230 8600 7275 8630
rect 7305 8600 7350 8630
rect 7230 8560 7350 8600
rect 7230 8530 7275 8560
rect 7305 8530 7350 8560
rect 7230 8495 7350 8530
rect 7230 8465 7275 8495
rect 7305 8465 7350 8495
rect 7230 8435 7350 8465
rect 7230 8405 7275 8435
rect 7305 8405 7350 8435
rect 7230 8370 7350 8405
rect 7230 8340 7275 8370
rect 7305 8340 7350 8370
rect 7230 8300 7350 8340
rect 7230 8270 7275 8300
rect 7305 8270 7350 8300
rect 7230 8230 7350 8270
rect 7230 8200 7275 8230
rect 7305 8200 7350 8230
rect 7230 8160 7350 8200
rect 7230 8130 7275 8160
rect 7305 8130 7350 8160
rect 7230 8095 7350 8130
rect 7230 8065 7275 8095
rect 7305 8065 7350 8095
rect 7230 8035 7350 8065
rect 7230 8005 7275 8035
rect 7305 8005 7350 8035
rect 7230 7970 7350 8005
rect 7230 7940 7275 7970
rect 7305 7940 7350 7970
rect 7230 7900 7350 7940
rect 7230 7870 7275 7900
rect 7305 7870 7350 7900
rect 7230 7830 7350 7870
rect 7230 7800 7275 7830
rect 7305 7800 7350 7830
rect 7230 7760 7350 7800
rect 7230 7730 7275 7760
rect 7305 7730 7350 7760
rect 7230 7695 7350 7730
rect 7230 7665 7275 7695
rect 7305 7665 7350 7695
rect 7230 7635 7350 7665
rect 7230 7605 7275 7635
rect 7305 7605 7350 7635
rect 7230 7570 7350 7605
rect 7230 7540 7275 7570
rect 7305 7540 7350 7570
rect 7230 7500 7350 7540
rect 7230 7470 7275 7500
rect 7305 7470 7350 7500
rect 7230 7430 7350 7470
rect 7230 7400 7275 7430
rect 7305 7400 7350 7430
rect 7230 7360 7350 7400
rect 7230 7330 7275 7360
rect 7305 7330 7350 7360
rect 7230 7295 7350 7330
rect 7230 7265 7275 7295
rect 7305 7265 7350 7295
rect 7230 7235 7350 7265
rect 7230 7205 7275 7235
rect 7305 7205 7350 7235
rect 7230 7170 7350 7205
rect 7230 7140 7275 7170
rect 7305 7140 7350 7170
rect 7230 7100 7350 7140
rect 7230 7070 7275 7100
rect 7305 7070 7350 7100
rect 7230 7030 7350 7070
rect 7230 7000 7275 7030
rect 7305 7000 7350 7030
rect 7230 6960 7350 7000
rect 7230 6930 7275 6960
rect 7305 6930 7350 6960
rect 7230 6895 7350 6930
rect 7230 6865 7275 6895
rect 7305 6865 7350 6895
rect 7230 6835 7350 6865
rect 7230 6805 7275 6835
rect 7305 6805 7350 6835
rect 7230 6770 7350 6805
rect 7230 6740 7275 6770
rect 7305 6740 7350 6770
rect 7230 6700 7350 6740
rect 7230 6670 7275 6700
rect 7305 6670 7350 6700
rect 7230 6630 7350 6670
rect 7230 6600 7275 6630
rect 7305 6600 7350 6630
rect 7230 6560 7350 6600
rect 7230 6530 7275 6560
rect 7305 6530 7350 6560
rect 7230 6495 7350 6530
rect 7230 6465 7275 6495
rect 7305 6465 7350 6495
rect 6465 6430 6505 6435
rect 6465 6400 6470 6430
rect 6500 6400 6505 6430
rect 6465 6395 6505 6400
rect 6895 6430 6935 6435
rect 6895 6400 6900 6430
rect 6930 6400 6935 6430
rect 6895 6395 6935 6400
rect 5870 5085 5910 5090
rect 5870 5055 5875 5085
rect 5905 5055 5910 5085
rect 5870 5050 5910 5055
rect 6220 5085 6260 5090
rect 6220 5055 6225 5085
rect 6255 5055 6260 5085
rect 6220 5050 6260 5055
rect 5880 4585 5900 5050
rect 5870 4580 5910 4585
rect 5870 4550 5875 4580
rect 5905 4550 5910 4580
rect 5870 4545 5910 4550
rect 5320 2945 5350 2950
rect 3390 2930 3430 2935
rect 3390 2900 3395 2930
rect 3425 2900 3430 2930
rect 5320 2910 5350 2915
rect 5545 2945 5585 2950
rect 5545 2915 5550 2945
rect 5580 2915 5585 2945
rect 5545 2910 5585 2915
rect 3390 2895 3430 2900
rect 5325 2090 5345 2910
rect 6905 2010 6925 6395
rect 6940 6375 6980 6380
rect 6940 6345 6945 6375
rect 6975 6345 6980 6375
rect 6940 6340 6980 6345
rect 2045 2005 2085 2010
rect 2045 1975 2050 2005
rect 2080 1975 2085 2005
rect 2045 1970 2085 1975
rect 2200 2005 2240 2010
rect 2200 1975 2205 2005
rect 2235 1975 2240 2005
rect 2200 1970 2240 1975
rect 6740 2005 6780 2010
rect 6740 1975 6745 2005
rect 6775 1975 6780 2005
rect 6740 1970 6780 1975
rect 6895 2005 6935 2010
rect 6895 1975 6900 2005
rect 6930 1975 6935 2005
rect 6895 1970 6935 1975
rect 2000 1950 2040 1955
rect 2000 1920 2005 1950
rect 2035 1920 2040 1950
rect 2000 1915 2040 1920
rect 2155 1950 2195 1955
rect 2155 1920 2160 1950
rect 2190 1920 2195 1950
rect 2155 1915 2195 1920
rect 2165 1765 2185 1915
rect 2210 1580 2230 1970
rect 6750 1580 6770 1970
rect 6950 1955 6970 6340
rect 7230 6210 7350 6465
rect 7930 9635 8050 9650
rect 7930 9605 7975 9635
rect 8005 9605 8050 9635
rect 7930 9570 8050 9605
rect 7930 9540 7975 9570
rect 8005 9540 8050 9570
rect 7930 9500 8050 9540
rect 7930 9470 7975 9500
rect 8005 9470 8050 9500
rect 7930 9430 8050 9470
rect 7930 9400 7975 9430
rect 8005 9400 8050 9430
rect 7930 9360 8050 9400
rect 7930 9330 7975 9360
rect 8005 9330 8050 9360
rect 7930 9295 8050 9330
rect 7930 9265 7975 9295
rect 8005 9265 8050 9295
rect 7930 9235 8050 9265
rect 7930 9205 7975 9235
rect 8005 9205 8050 9235
rect 7930 9170 8050 9205
rect 7930 9140 7975 9170
rect 8005 9140 8050 9170
rect 7930 9100 8050 9140
rect 7930 9070 7975 9100
rect 8005 9070 8050 9100
rect 7930 9030 8050 9070
rect 7930 9000 7975 9030
rect 8005 9000 8050 9030
rect 7930 8960 8050 9000
rect 7930 8930 7975 8960
rect 8005 8930 8050 8960
rect 7930 8895 8050 8930
rect 7930 8865 7975 8895
rect 8005 8865 8050 8895
rect 7930 8835 8050 8865
rect 7930 8805 7975 8835
rect 8005 8805 8050 8835
rect 7930 8770 8050 8805
rect 7930 8740 7975 8770
rect 8005 8740 8050 8770
rect 7930 8700 8050 8740
rect 7930 8670 7975 8700
rect 8005 8670 8050 8700
rect 7930 8630 8050 8670
rect 7930 8600 7975 8630
rect 8005 8600 8050 8630
rect 7930 8560 8050 8600
rect 7930 8530 7975 8560
rect 8005 8530 8050 8560
rect 7930 8495 8050 8530
rect 7930 8465 7975 8495
rect 8005 8465 8050 8495
rect 7930 8435 8050 8465
rect 7930 8405 7975 8435
rect 8005 8405 8050 8435
rect 7930 8370 8050 8405
rect 7930 8340 7975 8370
rect 8005 8340 8050 8370
rect 7930 8300 8050 8340
rect 7930 8270 7975 8300
rect 8005 8270 8050 8300
rect 7930 8230 8050 8270
rect 7930 8200 7975 8230
rect 8005 8200 8050 8230
rect 7930 8160 8050 8200
rect 7930 8130 7975 8160
rect 8005 8130 8050 8160
rect 7930 8095 8050 8130
rect 7930 8065 7975 8095
rect 8005 8065 8050 8095
rect 7930 8035 8050 8065
rect 7930 8005 7975 8035
rect 8005 8005 8050 8035
rect 7930 7970 8050 8005
rect 7930 7940 7975 7970
rect 8005 7940 8050 7970
rect 7930 7900 8050 7940
rect 7930 7870 7975 7900
rect 8005 7870 8050 7900
rect 7930 7830 8050 7870
rect 7930 7800 7975 7830
rect 8005 7800 8050 7830
rect 7930 7760 8050 7800
rect 7930 7730 7975 7760
rect 8005 7730 8050 7760
rect 7930 7695 8050 7730
rect 7930 7665 7975 7695
rect 8005 7665 8050 7695
rect 7930 7635 8050 7665
rect 7930 7605 7975 7635
rect 8005 7605 8050 7635
rect 7930 7570 8050 7605
rect 7930 7540 7975 7570
rect 8005 7540 8050 7570
rect 7930 7500 8050 7540
rect 7930 7470 7975 7500
rect 8005 7470 8050 7500
rect 7930 7430 8050 7470
rect 7930 7400 7975 7430
rect 8005 7400 8050 7430
rect 7930 7360 8050 7400
rect 7930 7330 7975 7360
rect 8005 7330 8050 7360
rect 7930 7295 8050 7330
rect 7930 7265 7975 7295
rect 8005 7265 8050 7295
rect 7930 7235 8050 7265
rect 7930 7205 7975 7235
rect 8005 7205 8050 7235
rect 7930 7170 8050 7205
rect 7930 7140 7975 7170
rect 8005 7140 8050 7170
rect 7930 7100 8050 7140
rect 7930 7070 7975 7100
rect 8005 7070 8050 7100
rect 7930 7030 8050 7070
rect 7930 7000 7975 7030
rect 8005 7000 8050 7030
rect 7930 6960 8050 7000
rect 7930 6930 7975 6960
rect 8005 6930 8050 6960
rect 7930 6895 8050 6930
rect 7930 6865 7975 6895
rect 8005 6865 8050 6895
rect 7930 6835 8050 6865
rect 7930 6805 7975 6835
rect 8005 6805 8050 6835
rect 7930 6770 8050 6805
rect 7930 6740 7975 6770
rect 8005 6740 8050 6770
rect 7930 6700 8050 6740
rect 7930 6670 7975 6700
rect 8005 6670 8050 6700
rect 7930 6630 8050 6670
rect 7930 6600 7975 6630
rect 8005 6600 8050 6630
rect 7930 6560 8050 6600
rect 7930 6530 7975 6560
rect 8005 6530 8050 6560
rect 7930 6495 8050 6530
rect 7930 6465 7975 6495
rect 8005 6465 8050 6495
rect 7580 6205 7700 6210
rect 7580 6175 7585 6205
rect 7615 6175 7625 6205
rect 7655 6175 7665 6205
rect 7695 6175 7700 6205
rect 7930 6195 8050 6465
rect 8280 9635 8400 9650
rect 8280 9605 8325 9635
rect 8355 9605 8400 9635
rect 8280 9570 8400 9605
rect 8280 9540 8325 9570
rect 8355 9540 8400 9570
rect 8280 9500 8400 9540
rect 8280 9470 8325 9500
rect 8355 9470 8400 9500
rect 8280 9430 8400 9470
rect 8280 9400 8325 9430
rect 8355 9400 8400 9430
rect 8280 9360 8400 9400
rect 8280 9330 8325 9360
rect 8355 9330 8400 9360
rect 8280 9295 8400 9330
rect 8280 9265 8325 9295
rect 8355 9265 8400 9295
rect 8280 9235 8400 9265
rect 8280 9205 8325 9235
rect 8355 9205 8400 9235
rect 8280 9170 8400 9205
rect 8280 9140 8325 9170
rect 8355 9140 8400 9170
rect 8280 9100 8400 9140
rect 8280 9070 8325 9100
rect 8355 9070 8400 9100
rect 8280 9030 8400 9070
rect 8280 9000 8325 9030
rect 8355 9000 8400 9030
rect 8280 8960 8400 9000
rect 8280 8930 8325 8960
rect 8355 8930 8400 8960
rect 8280 8895 8400 8930
rect 8280 8865 8325 8895
rect 8355 8865 8400 8895
rect 8280 8835 8400 8865
rect 8280 8805 8325 8835
rect 8355 8805 8400 8835
rect 8280 8770 8400 8805
rect 8280 8740 8325 8770
rect 8355 8740 8400 8770
rect 8280 8700 8400 8740
rect 8280 8670 8325 8700
rect 8355 8670 8400 8700
rect 8280 8630 8400 8670
rect 8280 8600 8325 8630
rect 8355 8600 8400 8630
rect 8280 8560 8400 8600
rect 8280 8530 8325 8560
rect 8355 8530 8400 8560
rect 8280 8495 8400 8530
rect 8280 8465 8325 8495
rect 8355 8465 8400 8495
rect 8280 8435 8400 8465
rect 8280 8405 8325 8435
rect 8355 8405 8400 8435
rect 8280 8370 8400 8405
rect 8280 8340 8325 8370
rect 8355 8340 8400 8370
rect 8280 8300 8400 8340
rect 8280 8270 8325 8300
rect 8355 8270 8400 8300
rect 8280 8230 8400 8270
rect 8280 8200 8325 8230
rect 8355 8200 8400 8230
rect 8280 8160 8400 8200
rect 8280 8130 8325 8160
rect 8355 8130 8400 8160
rect 8280 8095 8400 8130
rect 8280 8065 8325 8095
rect 8355 8065 8400 8095
rect 8280 8035 8400 8065
rect 8280 8005 8325 8035
rect 8355 8005 8400 8035
rect 8280 7970 8400 8005
rect 8280 7940 8325 7970
rect 8355 7940 8400 7970
rect 8280 7900 8400 7940
rect 8280 7870 8325 7900
rect 8355 7870 8400 7900
rect 8280 7830 8400 7870
rect 8280 7800 8325 7830
rect 8355 7800 8400 7830
rect 8280 7760 8400 7800
rect 8280 7730 8325 7760
rect 8355 7730 8400 7760
rect 8280 7695 8400 7730
rect 8280 7665 8325 7695
rect 8355 7665 8400 7695
rect 8280 7635 8400 7665
rect 8280 7605 8325 7635
rect 8355 7605 8400 7635
rect 8280 7570 8400 7605
rect 8280 7540 8325 7570
rect 8355 7540 8400 7570
rect 8280 7500 8400 7540
rect 8280 7470 8325 7500
rect 8355 7470 8400 7500
rect 8280 7430 8400 7470
rect 8280 7400 8325 7430
rect 8355 7400 8400 7430
rect 8280 7360 8400 7400
rect 8280 7330 8325 7360
rect 8355 7330 8400 7360
rect 8280 7295 8400 7330
rect 8280 7265 8325 7295
rect 8355 7265 8400 7295
rect 8280 7235 8400 7265
rect 8280 7205 8325 7235
rect 8355 7205 8400 7235
rect 8280 7170 8400 7205
rect 8280 7140 8325 7170
rect 8355 7140 8400 7170
rect 8280 7100 8400 7140
rect 8280 7070 8325 7100
rect 8355 7070 8400 7100
rect 8280 7030 8400 7070
rect 8280 7000 8325 7030
rect 8355 7000 8400 7030
rect 8280 6960 8400 7000
rect 8280 6930 8325 6960
rect 8355 6930 8400 6960
rect 8280 6895 8400 6930
rect 8280 6865 8325 6895
rect 8355 6865 8400 6895
rect 8280 6835 8400 6865
rect 8280 6805 8325 6835
rect 8355 6805 8400 6835
rect 8280 6770 8400 6805
rect 8280 6740 8325 6770
rect 8355 6740 8400 6770
rect 8280 6700 8400 6740
rect 8280 6670 8325 6700
rect 8355 6670 8400 6700
rect 8280 6630 8400 6670
rect 8280 6600 8325 6630
rect 8355 6600 8400 6630
rect 8280 6560 8400 6600
rect 8280 6530 8325 6560
rect 8355 6530 8400 6560
rect 8280 6495 8400 6530
rect 8280 6465 8325 6495
rect 8355 6465 8400 6495
rect 8280 6210 8400 6465
rect 8630 9635 8750 9650
rect 8630 9605 8675 9635
rect 8705 9605 8750 9635
rect 8630 9570 8750 9605
rect 8630 9540 8675 9570
rect 8705 9540 8750 9570
rect 8630 9500 8750 9540
rect 8630 9470 8675 9500
rect 8705 9470 8750 9500
rect 8630 9430 8750 9470
rect 8630 9400 8675 9430
rect 8705 9400 8750 9430
rect 8630 9360 8750 9400
rect 8630 9330 8675 9360
rect 8705 9330 8750 9360
rect 8630 9295 8750 9330
rect 8630 9265 8675 9295
rect 8705 9265 8750 9295
rect 8630 9235 8750 9265
rect 8630 9205 8675 9235
rect 8705 9205 8750 9235
rect 8630 9170 8750 9205
rect 8630 9140 8675 9170
rect 8705 9140 8750 9170
rect 8630 9100 8750 9140
rect 8630 9070 8675 9100
rect 8705 9070 8750 9100
rect 8630 9030 8750 9070
rect 8630 9000 8675 9030
rect 8705 9000 8750 9030
rect 8630 8960 8750 9000
rect 8630 8930 8675 8960
rect 8705 8930 8750 8960
rect 8630 8895 8750 8930
rect 8630 8865 8675 8895
rect 8705 8865 8750 8895
rect 8630 8835 8750 8865
rect 8630 8805 8675 8835
rect 8705 8805 8750 8835
rect 8630 8770 8750 8805
rect 8630 8740 8675 8770
rect 8705 8740 8750 8770
rect 8630 8700 8750 8740
rect 8630 8670 8675 8700
rect 8705 8670 8750 8700
rect 8630 8630 8750 8670
rect 8630 8600 8675 8630
rect 8705 8600 8750 8630
rect 8630 8560 8750 8600
rect 8630 8530 8675 8560
rect 8705 8530 8750 8560
rect 8630 8495 8750 8530
rect 8630 8465 8675 8495
rect 8705 8465 8750 8495
rect 8630 8435 8750 8465
rect 8630 8405 8675 8435
rect 8705 8405 8750 8435
rect 8630 8370 8750 8405
rect 8630 8340 8675 8370
rect 8705 8340 8750 8370
rect 8630 8300 8750 8340
rect 8630 8270 8675 8300
rect 8705 8270 8750 8300
rect 8630 8230 8750 8270
rect 8630 8200 8675 8230
rect 8705 8200 8750 8230
rect 8630 8160 8750 8200
rect 8630 8130 8675 8160
rect 8705 8130 8750 8160
rect 8630 8095 8750 8130
rect 8630 8065 8675 8095
rect 8705 8065 8750 8095
rect 8630 8035 8750 8065
rect 8630 8005 8675 8035
rect 8705 8005 8750 8035
rect 8630 7970 8750 8005
rect 8630 7940 8675 7970
rect 8705 7940 8750 7970
rect 8630 7900 8750 7940
rect 8630 7870 8675 7900
rect 8705 7870 8750 7900
rect 8630 7830 8750 7870
rect 8630 7800 8675 7830
rect 8705 7800 8750 7830
rect 8630 7760 8750 7800
rect 8630 7730 8675 7760
rect 8705 7730 8750 7760
rect 8630 7695 8750 7730
rect 8630 7665 8675 7695
rect 8705 7665 8750 7695
rect 8630 7635 8750 7665
rect 8630 7605 8675 7635
rect 8705 7605 8750 7635
rect 8630 7570 8750 7605
rect 8630 7540 8675 7570
rect 8705 7540 8750 7570
rect 8630 7500 8750 7540
rect 8630 7470 8675 7500
rect 8705 7470 8750 7500
rect 8630 7430 8750 7470
rect 8630 7400 8675 7430
rect 8705 7400 8750 7430
rect 8630 7360 8750 7400
rect 8630 7330 8675 7360
rect 8705 7330 8750 7360
rect 8630 7295 8750 7330
rect 8630 7265 8675 7295
rect 8705 7265 8750 7295
rect 8630 7235 8750 7265
rect 8630 7205 8675 7235
rect 8705 7205 8750 7235
rect 8630 7170 8750 7205
rect 8630 7140 8675 7170
rect 8705 7140 8750 7170
rect 8630 7100 8750 7140
rect 8630 7070 8675 7100
rect 8705 7070 8750 7100
rect 8630 7030 8750 7070
rect 8630 7000 8675 7030
rect 8705 7000 8750 7030
rect 8630 6960 8750 7000
rect 8630 6930 8675 6960
rect 8705 6930 8750 6960
rect 8630 6895 8750 6930
rect 8630 6865 8675 6895
rect 8705 6865 8750 6895
rect 8630 6835 8750 6865
rect 8630 6805 8675 6835
rect 8705 6805 8750 6835
rect 8630 6770 8750 6805
rect 8630 6740 8675 6770
rect 8705 6740 8750 6770
rect 8630 6700 8750 6740
rect 8630 6670 8675 6700
rect 8705 6670 8750 6700
rect 8630 6630 8750 6670
rect 8630 6600 8675 6630
rect 8705 6600 8750 6630
rect 8630 6560 8750 6600
rect 8630 6530 8675 6560
rect 8705 6530 8750 6560
rect 8630 6495 8750 6530
rect 8630 6465 8675 6495
rect 8705 6465 8750 6495
rect 8630 6210 8750 6465
rect 8980 9635 9100 9650
rect 8980 9605 9025 9635
rect 9055 9605 9100 9635
rect 8980 9570 9100 9605
rect 8980 9540 9025 9570
rect 9055 9540 9100 9570
rect 8980 9500 9100 9540
rect 8980 9470 9025 9500
rect 9055 9470 9100 9500
rect 8980 9430 9100 9470
rect 8980 9400 9025 9430
rect 9055 9400 9100 9430
rect 8980 9360 9100 9400
rect 8980 9330 9025 9360
rect 9055 9330 9100 9360
rect 8980 9295 9100 9330
rect 8980 9265 9025 9295
rect 9055 9265 9100 9295
rect 8980 9235 9100 9265
rect 8980 9205 9025 9235
rect 9055 9205 9100 9235
rect 8980 9170 9100 9205
rect 8980 9140 9025 9170
rect 9055 9140 9100 9170
rect 8980 9100 9100 9140
rect 8980 9070 9025 9100
rect 9055 9070 9100 9100
rect 8980 9030 9100 9070
rect 8980 9000 9025 9030
rect 9055 9000 9100 9030
rect 8980 8960 9100 9000
rect 8980 8930 9025 8960
rect 9055 8930 9100 8960
rect 8980 8895 9100 8930
rect 8980 8865 9025 8895
rect 9055 8865 9100 8895
rect 8980 8835 9100 8865
rect 8980 8805 9025 8835
rect 9055 8805 9100 8835
rect 8980 8770 9100 8805
rect 8980 8740 9025 8770
rect 9055 8740 9100 8770
rect 8980 8700 9100 8740
rect 8980 8670 9025 8700
rect 9055 8670 9100 8700
rect 8980 8630 9100 8670
rect 8980 8600 9025 8630
rect 9055 8600 9100 8630
rect 8980 8560 9100 8600
rect 8980 8530 9025 8560
rect 9055 8530 9100 8560
rect 8980 8495 9100 8530
rect 8980 8465 9025 8495
rect 9055 8465 9100 8495
rect 8980 8435 9100 8465
rect 8980 8405 9025 8435
rect 9055 8405 9100 8435
rect 8980 8370 9100 8405
rect 8980 8340 9025 8370
rect 9055 8340 9100 8370
rect 8980 8300 9100 8340
rect 8980 8270 9025 8300
rect 9055 8270 9100 8300
rect 8980 8230 9100 8270
rect 8980 8200 9025 8230
rect 9055 8200 9100 8230
rect 8980 8160 9100 8200
rect 8980 8130 9025 8160
rect 9055 8130 9100 8160
rect 8980 8095 9100 8130
rect 8980 8065 9025 8095
rect 9055 8065 9100 8095
rect 8980 8035 9100 8065
rect 8980 8005 9025 8035
rect 9055 8005 9100 8035
rect 8980 7970 9100 8005
rect 8980 7940 9025 7970
rect 9055 7940 9100 7970
rect 8980 7900 9100 7940
rect 8980 7870 9025 7900
rect 9055 7870 9100 7900
rect 8980 7830 9100 7870
rect 8980 7800 9025 7830
rect 9055 7800 9100 7830
rect 8980 7760 9100 7800
rect 8980 7730 9025 7760
rect 9055 7730 9100 7760
rect 8980 7695 9100 7730
rect 8980 7665 9025 7695
rect 9055 7665 9100 7695
rect 8980 7635 9100 7665
rect 8980 7605 9025 7635
rect 9055 7605 9100 7635
rect 8980 7570 9100 7605
rect 8980 7540 9025 7570
rect 9055 7540 9100 7570
rect 8980 7500 9100 7540
rect 8980 7470 9025 7500
rect 9055 7470 9100 7500
rect 8980 7430 9100 7470
rect 8980 7400 9025 7430
rect 9055 7400 9100 7430
rect 8980 7360 9100 7400
rect 8980 7330 9025 7360
rect 9055 7330 9100 7360
rect 8980 7295 9100 7330
rect 8980 7265 9025 7295
rect 9055 7265 9100 7295
rect 8980 7235 9100 7265
rect 8980 7205 9025 7235
rect 9055 7205 9100 7235
rect 8980 7170 9100 7205
rect 8980 7140 9025 7170
rect 9055 7140 9100 7170
rect 8980 7100 9100 7140
rect 8980 7070 9025 7100
rect 9055 7070 9100 7100
rect 8980 7030 9100 7070
rect 8980 7000 9025 7030
rect 9055 7000 9100 7030
rect 8980 6960 9100 7000
rect 8980 6930 9025 6960
rect 9055 6930 9100 6960
rect 8980 6895 9100 6930
rect 8980 6865 9025 6895
rect 9055 6865 9100 6895
rect 8980 6835 9100 6865
rect 8980 6805 9025 6835
rect 9055 6805 9100 6835
rect 8980 6770 9100 6805
rect 8980 6740 9025 6770
rect 9055 6740 9100 6770
rect 8980 6700 9100 6740
rect 8980 6670 9025 6700
rect 9055 6670 9100 6700
rect 8980 6630 9100 6670
rect 8980 6600 9025 6630
rect 9055 6600 9100 6630
rect 8980 6560 9100 6600
rect 8980 6530 9025 6560
rect 9055 6530 9100 6560
rect 8980 6495 9100 6530
rect 8980 6465 9025 6495
rect 9055 6465 9100 6495
rect 8980 6210 9100 6465
rect 7580 6165 7700 6175
rect 7580 6135 7585 6165
rect 7615 6135 7625 6165
rect 7655 6135 7665 6165
rect 7695 6135 7700 6165
rect 7580 6125 7700 6135
rect 7580 6095 7585 6125
rect 7615 6095 7625 6125
rect 7655 6095 7665 6125
rect 7695 6095 7700 6125
rect 6785 1950 6825 1955
rect 6785 1920 6790 1950
rect 6820 1920 6825 1950
rect 6785 1915 6825 1920
rect 6940 1950 6980 1955
rect 6940 1920 6945 1950
rect 6975 1920 6980 1950
rect 6940 1915 6980 1920
rect 6795 1765 6815 1915
rect 1280 820 1285 850
rect 1315 820 1325 850
rect 1355 820 1365 850
rect 1395 820 1400 850
rect 1280 810 1400 820
rect 1280 780 1285 810
rect 1315 780 1325 810
rect 1355 780 1365 810
rect 1395 780 1400 810
rect 1280 770 1400 780
rect 1280 740 1285 770
rect 1315 740 1325 770
rect 1355 740 1365 770
rect 1395 740 1400 770
rect 1280 735 1400 740
rect 4415 850 4565 855
rect 4415 820 4420 850
rect 4450 820 4475 850
rect 4505 820 4530 850
rect 4560 820 4565 850
rect 4415 810 4565 820
rect 4415 780 4420 810
rect 4450 780 4475 810
rect 4505 780 4530 810
rect 4560 780 4565 810
rect 4415 770 4565 780
rect 4415 740 4420 770
rect 4450 740 4475 770
rect 4505 740 4530 770
rect 4560 740 4565 770
rect 4415 735 4565 740
rect 7580 850 7700 6095
rect 7580 820 7585 850
rect 7615 820 7625 850
rect 7655 820 7665 850
rect 7695 820 7700 850
rect 7580 810 7700 820
rect 7580 780 7585 810
rect 7615 780 7625 810
rect 7655 780 7665 810
rect 7695 780 7700 810
rect 7580 770 7700 780
rect 7580 740 7585 770
rect 7615 740 7625 770
rect 7655 740 7665 770
rect 7695 740 7700 770
rect 7580 735 7700 740
rect -120 -1305 0 -1240
rect -120 -1335 -75 -1305
rect -45 -1335 0 -1305
rect -120 -1370 0 -1335
rect -120 -1400 -75 -1370
rect -45 -1400 0 -1370
rect -120 -1440 0 -1400
rect -120 -1470 -75 -1440
rect -45 -1470 0 -1440
rect -120 -1510 0 -1470
rect -120 -1540 -75 -1510
rect -45 -1540 0 -1510
rect -120 -1580 0 -1540
rect -120 -1610 -75 -1580
rect -45 -1610 0 -1580
rect -120 -1645 0 -1610
rect -120 -1675 -75 -1645
rect -45 -1675 0 -1645
rect -120 -1705 0 -1675
rect -120 -1735 -75 -1705
rect -45 -1735 0 -1705
rect -120 -1770 0 -1735
rect -120 -1800 -75 -1770
rect -45 -1800 0 -1770
rect -120 -1840 0 -1800
rect -120 -1870 -75 -1840
rect -45 -1870 0 -1840
rect -120 -1910 0 -1870
rect -120 -1940 -75 -1910
rect -45 -1940 0 -1910
rect -120 -1980 0 -1940
rect -120 -2010 -75 -1980
rect -45 -2010 0 -1980
rect -120 -2045 0 -2010
rect -120 -2075 -75 -2045
rect -45 -2075 0 -2045
rect -120 -2105 0 -2075
rect -120 -2135 -75 -2105
rect -45 -2135 0 -2105
rect -120 -2170 0 -2135
rect -120 -2200 -75 -2170
rect -45 -2200 0 -2170
rect -120 -2240 0 -2200
rect -120 -2270 -75 -2240
rect -45 -2270 0 -2240
rect -120 -2310 0 -2270
rect -120 -2340 -75 -2310
rect -45 -2340 0 -2310
rect -120 -2380 0 -2340
rect -120 -2410 -75 -2380
rect -45 -2410 0 -2380
rect -120 -2445 0 -2410
rect -120 -2475 -75 -2445
rect -45 -2475 0 -2445
rect -120 -2505 0 -2475
rect -120 -2535 -75 -2505
rect -45 -2535 0 -2505
rect -120 -2570 0 -2535
rect -120 -2600 -75 -2570
rect -45 -2600 0 -2570
rect -120 -2640 0 -2600
rect -120 -2670 -75 -2640
rect -45 -2670 0 -2640
rect -120 -2710 0 -2670
rect -120 -2740 -75 -2710
rect -45 -2740 0 -2710
rect -120 -2780 0 -2740
rect -120 -2810 -75 -2780
rect -45 -2810 0 -2780
rect -120 -2845 0 -2810
rect -120 -2875 -75 -2845
rect -45 -2875 0 -2845
rect -120 -2905 0 -2875
rect -120 -2935 -75 -2905
rect -45 -2935 0 -2905
rect -120 -2970 0 -2935
rect -120 -3000 -75 -2970
rect -45 -3000 0 -2970
rect -120 -3040 0 -3000
rect -120 -3070 -75 -3040
rect -45 -3070 0 -3040
rect -120 -3110 0 -3070
rect -120 -3140 -75 -3110
rect -45 -3140 0 -3110
rect -120 -3180 0 -3140
rect -120 -3210 -75 -3180
rect -45 -3210 0 -3180
rect -120 -3245 0 -3210
rect -120 -3275 -75 -3245
rect -45 -3275 0 -3245
rect -120 -3305 0 -3275
rect -120 -3335 -75 -3305
rect -45 -3335 0 -3305
rect -120 -3370 0 -3335
rect -120 -3400 -75 -3370
rect -45 -3400 0 -3370
rect -120 -3440 0 -3400
rect -120 -3470 -75 -3440
rect -45 -3470 0 -3440
rect -120 -3510 0 -3470
rect -120 -3540 -75 -3510
rect -45 -3540 0 -3510
rect -120 -3580 0 -3540
rect -120 -3610 -75 -3580
rect -45 -3610 0 -3580
rect -120 -3645 0 -3610
rect -120 -3675 -75 -3645
rect -45 -3675 0 -3645
rect -120 -3705 0 -3675
rect -120 -3735 -75 -3705
rect -45 -3735 0 -3705
rect -120 -3770 0 -3735
rect -120 -3800 -75 -3770
rect -45 -3800 0 -3770
rect -120 -3840 0 -3800
rect -120 -3870 -75 -3840
rect -45 -3870 0 -3840
rect -120 -3910 0 -3870
rect -120 -3940 -75 -3910
rect -45 -3940 0 -3910
rect -120 -3980 0 -3940
rect -120 -4010 -75 -3980
rect -45 -4010 0 -3980
rect -120 -4045 0 -4010
rect -120 -4075 -75 -4045
rect -45 -4075 0 -4045
rect -120 -4105 0 -4075
rect -120 -4135 -75 -4105
rect -45 -4135 0 -4105
rect -120 -4170 0 -4135
rect -120 -4200 -75 -4170
rect -45 -4200 0 -4170
rect -120 -4240 0 -4200
rect -120 -4270 -75 -4240
rect -45 -4270 0 -4240
rect -120 -4310 0 -4270
rect -120 -4340 -75 -4310
rect -45 -4340 0 -4310
rect -120 -4380 0 -4340
rect -120 -4410 -75 -4380
rect -45 -4410 0 -4380
rect -120 -4445 0 -4410
rect -120 -4475 -75 -4445
rect -45 -4475 0 -4445
rect -120 -4490 0 -4475
rect 230 -1305 350 -1240
rect 230 -1335 275 -1305
rect 305 -1335 350 -1305
rect 230 -1370 350 -1335
rect 230 -1400 275 -1370
rect 305 -1400 350 -1370
rect 230 -1440 350 -1400
rect 230 -1470 275 -1440
rect 305 -1470 350 -1440
rect 230 -1510 350 -1470
rect 230 -1540 275 -1510
rect 305 -1540 350 -1510
rect 230 -1580 350 -1540
rect 230 -1610 275 -1580
rect 305 -1610 350 -1580
rect 230 -1645 350 -1610
rect 230 -1675 275 -1645
rect 305 -1675 350 -1645
rect 230 -1705 350 -1675
rect 230 -1735 275 -1705
rect 305 -1735 350 -1705
rect 230 -1770 350 -1735
rect 230 -1800 275 -1770
rect 305 -1800 350 -1770
rect 230 -1840 350 -1800
rect 230 -1870 275 -1840
rect 305 -1870 350 -1840
rect 230 -1910 350 -1870
rect 230 -1940 275 -1910
rect 305 -1940 350 -1910
rect 230 -1980 350 -1940
rect 230 -2010 275 -1980
rect 305 -2010 350 -1980
rect 230 -2045 350 -2010
rect 230 -2075 275 -2045
rect 305 -2075 350 -2045
rect 230 -2105 350 -2075
rect 230 -2135 275 -2105
rect 305 -2135 350 -2105
rect 230 -2170 350 -2135
rect 230 -2200 275 -2170
rect 305 -2200 350 -2170
rect 230 -2240 350 -2200
rect 230 -2270 275 -2240
rect 305 -2270 350 -2240
rect 230 -2310 350 -2270
rect 230 -2340 275 -2310
rect 305 -2340 350 -2310
rect 230 -2380 350 -2340
rect 230 -2410 275 -2380
rect 305 -2410 350 -2380
rect 230 -2445 350 -2410
rect 230 -2475 275 -2445
rect 305 -2475 350 -2445
rect 230 -2505 350 -2475
rect 230 -2535 275 -2505
rect 305 -2535 350 -2505
rect 230 -2570 350 -2535
rect 230 -2600 275 -2570
rect 305 -2600 350 -2570
rect 230 -2640 350 -2600
rect 230 -2670 275 -2640
rect 305 -2670 350 -2640
rect 230 -2710 350 -2670
rect 230 -2740 275 -2710
rect 305 -2740 350 -2710
rect 230 -2780 350 -2740
rect 230 -2810 275 -2780
rect 305 -2810 350 -2780
rect 230 -2845 350 -2810
rect 230 -2875 275 -2845
rect 305 -2875 350 -2845
rect 230 -2905 350 -2875
rect 230 -2935 275 -2905
rect 305 -2935 350 -2905
rect 230 -2970 350 -2935
rect 230 -3000 275 -2970
rect 305 -3000 350 -2970
rect 230 -3040 350 -3000
rect 230 -3070 275 -3040
rect 305 -3070 350 -3040
rect 230 -3110 350 -3070
rect 230 -3140 275 -3110
rect 305 -3140 350 -3110
rect 230 -3180 350 -3140
rect 230 -3210 275 -3180
rect 305 -3210 350 -3180
rect 230 -3245 350 -3210
rect 230 -3275 275 -3245
rect 305 -3275 350 -3245
rect 230 -3305 350 -3275
rect 230 -3335 275 -3305
rect 305 -3335 350 -3305
rect 230 -3370 350 -3335
rect 230 -3400 275 -3370
rect 305 -3400 350 -3370
rect 230 -3440 350 -3400
rect 230 -3470 275 -3440
rect 305 -3470 350 -3440
rect 230 -3510 350 -3470
rect 230 -3540 275 -3510
rect 305 -3540 350 -3510
rect 230 -3580 350 -3540
rect 230 -3610 275 -3580
rect 305 -3610 350 -3580
rect 230 -3645 350 -3610
rect 230 -3675 275 -3645
rect 305 -3675 350 -3645
rect 230 -3705 350 -3675
rect 230 -3735 275 -3705
rect 305 -3735 350 -3705
rect 230 -3770 350 -3735
rect 230 -3800 275 -3770
rect 305 -3800 350 -3770
rect 230 -3840 350 -3800
rect 230 -3870 275 -3840
rect 305 -3870 350 -3840
rect 230 -3910 350 -3870
rect 230 -3940 275 -3910
rect 305 -3940 350 -3910
rect 230 -3980 350 -3940
rect 230 -4010 275 -3980
rect 305 -4010 350 -3980
rect 230 -4045 350 -4010
rect 230 -4075 275 -4045
rect 305 -4075 350 -4045
rect 230 -4105 350 -4075
rect 230 -4135 275 -4105
rect 305 -4135 350 -4105
rect 230 -4170 350 -4135
rect 230 -4200 275 -4170
rect 305 -4200 350 -4170
rect 230 -4240 350 -4200
rect 230 -4270 275 -4240
rect 305 -4270 350 -4240
rect 230 -4310 350 -4270
rect 230 -4340 275 -4310
rect 305 -4340 350 -4310
rect 230 -4380 350 -4340
rect 230 -4410 275 -4380
rect 305 -4410 350 -4380
rect 230 -4445 350 -4410
rect 230 -4475 275 -4445
rect 305 -4475 350 -4445
rect 230 -4490 350 -4475
rect 580 -1305 700 -1240
rect 580 -1335 625 -1305
rect 655 -1335 700 -1305
rect 580 -1370 700 -1335
rect 580 -1400 625 -1370
rect 655 -1400 700 -1370
rect 580 -1440 700 -1400
rect 580 -1470 625 -1440
rect 655 -1470 700 -1440
rect 580 -1510 700 -1470
rect 580 -1540 625 -1510
rect 655 -1540 700 -1510
rect 580 -1580 700 -1540
rect 580 -1610 625 -1580
rect 655 -1610 700 -1580
rect 580 -1645 700 -1610
rect 580 -1675 625 -1645
rect 655 -1675 700 -1645
rect 580 -1705 700 -1675
rect 580 -1735 625 -1705
rect 655 -1735 700 -1705
rect 580 -1770 700 -1735
rect 580 -1800 625 -1770
rect 655 -1800 700 -1770
rect 580 -1840 700 -1800
rect 580 -1870 625 -1840
rect 655 -1870 700 -1840
rect 580 -1910 700 -1870
rect 580 -1940 625 -1910
rect 655 -1940 700 -1910
rect 580 -1980 700 -1940
rect 580 -2010 625 -1980
rect 655 -2010 700 -1980
rect 580 -2045 700 -2010
rect 580 -2075 625 -2045
rect 655 -2075 700 -2045
rect 580 -2105 700 -2075
rect 580 -2135 625 -2105
rect 655 -2135 700 -2105
rect 580 -2170 700 -2135
rect 580 -2200 625 -2170
rect 655 -2200 700 -2170
rect 580 -2240 700 -2200
rect 580 -2270 625 -2240
rect 655 -2270 700 -2240
rect 580 -2310 700 -2270
rect 580 -2340 625 -2310
rect 655 -2340 700 -2310
rect 580 -2380 700 -2340
rect 580 -2410 625 -2380
rect 655 -2410 700 -2380
rect 580 -2445 700 -2410
rect 580 -2475 625 -2445
rect 655 -2475 700 -2445
rect 580 -2505 700 -2475
rect 580 -2535 625 -2505
rect 655 -2535 700 -2505
rect 580 -2570 700 -2535
rect 580 -2600 625 -2570
rect 655 -2600 700 -2570
rect 580 -2640 700 -2600
rect 580 -2670 625 -2640
rect 655 -2670 700 -2640
rect 580 -2710 700 -2670
rect 580 -2740 625 -2710
rect 655 -2740 700 -2710
rect 580 -2780 700 -2740
rect 580 -2810 625 -2780
rect 655 -2810 700 -2780
rect 580 -2845 700 -2810
rect 580 -2875 625 -2845
rect 655 -2875 700 -2845
rect 580 -2905 700 -2875
rect 580 -2935 625 -2905
rect 655 -2935 700 -2905
rect 580 -2970 700 -2935
rect 580 -3000 625 -2970
rect 655 -3000 700 -2970
rect 580 -3040 700 -3000
rect 580 -3070 625 -3040
rect 655 -3070 700 -3040
rect 580 -3110 700 -3070
rect 580 -3140 625 -3110
rect 655 -3140 700 -3110
rect 580 -3180 700 -3140
rect 580 -3210 625 -3180
rect 655 -3210 700 -3180
rect 580 -3245 700 -3210
rect 580 -3275 625 -3245
rect 655 -3275 700 -3245
rect 580 -3305 700 -3275
rect 580 -3335 625 -3305
rect 655 -3335 700 -3305
rect 580 -3370 700 -3335
rect 580 -3400 625 -3370
rect 655 -3400 700 -3370
rect 580 -3440 700 -3400
rect 580 -3470 625 -3440
rect 655 -3470 700 -3440
rect 580 -3510 700 -3470
rect 580 -3540 625 -3510
rect 655 -3540 700 -3510
rect 580 -3580 700 -3540
rect 580 -3610 625 -3580
rect 655 -3610 700 -3580
rect 580 -3645 700 -3610
rect 580 -3675 625 -3645
rect 655 -3675 700 -3645
rect 580 -3705 700 -3675
rect 580 -3735 625 -3705
rect 655 -3735 700 -3705
rect 580 -3770 700 -3735
rect 580 -3800 625 -3770
rect 655 -3800 700 -3770
rect 580 -3840 700 -3800
rect 580 -3870 625 -3840
rect 655 -3870 700 -3840
rect 580 -3910 700 -3870
rect 580 -3940 625 -3910
rect 655 -3940 700 -3910
rect 580 -3980 700 -3940
rect 580 -4010 625 -3980
rect 655 -4010 700 -3980
rect 580 -4045 700 -4010
rect 580 -4075 625 -4045
rect 655 -4075 700 -4045
rect 580 -4105 700 -4075
rect 580 -4135 625 -4105
rect 655 -4135 700 -4105
rect 580 -4170 700 -4135
rect 580 -4200 625 -4170
rect 655 -4200 700 -4170
rect 580 -4240 700 -4200
rect 580 -4270 625 -4240
rect 655 -4270 700 -4240
rect 580 -4310 700 -4270
rect 580 -4340 625 -4310
rect 655 -4340 700 -4310
rect 580 -4380 700 -4340
rect 580 -4410 625 -4380
rect 655 -4410 700 -4380
rect 580 -4445 700 -4410
rect 580 -4475 625 -4445
rect 655 -4475 700 -4445
rect 580 -4490 700 -4475
rect 930 -1305 1050 -1240
rect 930 -1335 975 -1305
rect 1005 -1335 1050 -1305
rect 930 -1370 1050 -1335
rect 930 -1400 975 -1370
rect 1005 -1400 1050 -1370
rect 930 -1440 1050 -1400
rect 930 -1470 975 -1440
rect 1005 -1470 1050 -1440
rect 930 -1510 1050 -1470
rect 930 -1540 975 -1510
rect 1005 -1540 1050 -1510
rect 930 -1580 1050 -1540
rect 930 -1610 975 -1580
rect 1005 -1610 1050 -1580
rect 930 -1645 1050 -1610
rect 930 -1675 975 -1645
rect 1005 -1675 1050 -1645
rect 930 -1705 1050 -1675
rect 930 -1735 975 -1705
rect 1005 -1735 1050 -1705
rect 930 -1770 1050 -1735
rect 930 -1800 975 -1770
rect 1005 -1800 1050 -1770
rect 930 -1840 1050 -1800
rect 930 -1870 975 -1840
rect 1005 -1870 1050 -1840
rect 930 -1910 1050 -1870
rect 930 -1940 975 -1910
rect 1005 -1940 1050 -1910
rect 930 -1980 1050 -1940
rect 930 -2010 975 -1980
rect 1005 -2010 1050 -1980
rect 930 -2045 1050 -2010
rect 930 -2075 975 -2045
rect 1005 -2075 1050 -2045
rect 930 -2105 1050 -2075
rect 930 -2135 975 -2105
rect 1005 -2135 1050 -2105
rect 930 -2170 1050 -2135
rect 930 -2200 975 -2170
rect 1005 -2200 1050 -2170
rect 930 -2240 1050 -2200
rect 930 -2270 975 -2240
rect 1005 -2270 1050 -2240
rect 930 -2310 1050 -2270
rect 930 -2340 975 -2310
rect 1005 -2340 1050 -2310
rect 930 -2380 1050 -2340
rect 930 -2410 975 -2380
rect 1005 -2410 1050 -2380
rect 930 -2445 1050 -2410
rect 930 -2475 975 -2445
rect 1005 -2475 1050 -2445
rect 930 -2505 1050 -2475
rect 930 -2535 975 -2505
rect 1005 -2535 1050 -2505
rect 930 -2570 1050 -2535
rect 930 -2600 975 -2570
rect 1005 -2600 1050 -2570
rect 930 -2640 1050 -2600
rect 930 -2670 975 -2640
rect 1005 -2670 1050 -2640
rect 930 -2710 1050 -2670
rect 930 -2740 975 -2710
rect 1005 -2740 1050 -2710
rect 930 -2780 1050 -2740
rect 930 -2810 975 -2780
rect 1005 -2810 1050 -2780
rect 930 -2845 1050 -2810
rect 930 -2875 975 -2845
rect 1005 -2875 1050 -2845
rect 930 -2905 1050 -2875
rect 930 -2935 975 -2905
rect 1005 -2935 1050 -2905
rect 930 -2970 1050 -2935
rect 930 -3000 975 -2970
rect 1005 -3000 1050 -2970
rect 930 -3040 1050 -3000
rect 930 -3070 975 -3040
rect 1005 -3070 1050 -3040
rect 930 -3110 1050 -3070
rect 930 -3140 975 -3110
rect 1005 -3140 1050 -3110
rect 930 -3180 1050 -3140
rect 930 -3210 975 -3180
rect 1005 -3210 1050 -3180
rect 930 -3245 1050 -3210
rect 930 -3275 975 -3245
rect 1005 -3275 1050 -3245
rect 930 -3305 1050 -3275
rect 930 -3335 975 -3305
rect 1005 -3335 1050 -3305
rect 930 -3370 1050 -3335
rect 930 -3400 975 -3370
rect 1005 -3400 1050 -3370
rect 930 -3440 1050 -3400
rect 930 -3470 975 -3440
rect 1005 -3470 1050 -3440
rect 930 -3510 1050 -3470
rect 930 -3540 975 -3510
rect 1005 -3540 1050 -3510
rect 930 -3580 1050 -3540
rect 930 -3610 975 -3580
rect 1005 -3610 1050 -3580
rect 930 -3645 1050 -3610
rect 930 -3675 975 -3645
rect 1005 -3675 1050 -3645
rect 930 -3705 1050 -3675
rect 930 -3735 975 -3705
rect 1005 -3735 1050 -3705
rect 930 -3770 1050 -3735
rect 930 -3800 975 -3770
rect 1005 -3800 1050 -3770
rect 930 -3840 1050 -3800
rect 930 -3870 975 -3840
rect 1005 -3870 1050 -3840
rect 930 -3910 1050 -3870
rect 930 -3940 975 -3910
rect 1005 -3940 1050 -3910
rect 930 -3980 1050 -3940
rect 930 -4010 975 -3980
rect 1005 -4010 1050 -3980
rect 930 -4045 1050 -4010
rect 930 -4075 975 -4045
rect 1005 -4075 1050 -4045
rect 930 -4105 1050 -4075
rect 930 -4135 975 -4105
rect 1005 -4135 1050 -4105
rect 930 -4170 1050 -4135
rect 930 -4200 975 -4170
rect 1005 -4200 1050 -4170
rect 930 -4240 1050 -4200
rect 930 -4270 975 -4240
rect 1005 -4270 1050 -4240
rect 930 -4310 1050 -4270
rect 930 -4340 975 -4310
rect 1005 -4340 1050 -4310
rect 930 -4380 1050 -4340
rect 930 -4410 975 -4380
rect 1005 -4410 1050 -4380
rect 930 -4445 1050 -4410
rect 930 -4475 975 -4445
rect 1005 -4475 1050 -4445
rect 930 -4490 1050 -4475
rect 1280 -1305 1400 -1240
rect 1280 -1335 1325 -1305
rect 1355 -1335 1400 -1305
rect 1280 -1370 1400 -1335
rect 1280 -1400 1325 -1370
rect 1355 -1400 1400 -1370
rect 1280 -1440 1400 -1400
rect 1280 -1470 1325 -1440
rect 1355 -1470 1400 -1440
rect 1280 -1510 1400 -1470
rect 1280 -1540 1325 -1510
rect 1355 -1540 1400 -1510
rect 1280 -1580 1400 -1540
rect 1280 -1610 1325 -1580
rect 1355 -1610 1400 -1580
rect 1280 -1645 1400 -1610
rect 1280 -1675 1325 -1645
rect 1355 -1675 1400 -1645
rect 1280 -1705 1400 -1675
rect 1280 -1735 1325 -1705
rect 1355 -1735 1400 -1705
rect 1280 -1770 1400 -1735
rect 1280 -1800 1325 -1770
rect 1355 -1800 1400 -1770
rect 1280 -1840 1400 -1800
rect 1280 -1870 1325 -1840
rect 1355 -1870 1400 -1840
rect 1280 -1910 1400 -1870
rect 1280 -1940 1325 -1910
rect 1355 -1940 1400 -1910
rect 1280 -1980 1400 -1940
rect 1280 -2010 1325 -1980
rect 1355 -2010 1400 -1980
rect 1280 -2045 1400 -2010
rect 1280 -2075 1325 -2045
rect 1355 -2075 1400 -2045
rect 1280 -2105 1400 -2075
rect 1280 -2135 1325 -2105
rect 1355 -2135 1400 -2105
rect 1280 -2170 1400 -2135
rect 1280 -2200 1325 -2170
rect 1355 -2200 1400 -2170
rect 1280 -2240 1400 -2200
rect 1280 -2270 1325 -2240
rect 1355 -2270 1400 -2240
rect 1280 -2310 1400 -2270
rect 1280 -2340 1325 -2310
rect 1355 -2340 1400 -2310
rect 1280 -2380 1400 -2340
rect 1280 -2410 1325 -2380
rect 1355 -2410 1400 -2380
rect 1280 -2445 1400 -2410
rect 1280 -2475 1325 -2445
rect 1355 -2475 1400 -2445
rect 1280 -2505 1400 -2475
rect 1280 -2535 1325 -2505
rect 1355 -2535 1400 -2505
rect 1280 -2570 1400 -2535
rect 1280 -2600 1325 -2570
rect 1355 -2600 1400 -2570
rect 1280 -2640 1400 -2600
rect 1280 -2670 1325 -2640
rect 1355 -2670 1400 -2640
rect 1280 -2710 1400 -2670
rect 1280 -2740 1325 -2710
rect 1355 -2740 1400 -2710
rect 1280 -2780 1400 -2740
rect 1280 -2810 1325 -2780
rect 1355 -2810 1400 -2780
rect 1280 -2845 1400 -2810
rect 1280 -2875 1325 -2845
rect 1355 -2875 1400 -2845
rect 1280 -2905 1400 -2875
rect 1280 -2935 1325 -2905
rect 1355 -2935 1400 -2905
rect 1280 -2970 1400 -2935
rect 1280 -3000 1325 -2970
rect 1355 -3000 1400 -2970
rect 1280 -3040 1400 -3000
rect 1280 -3070 1325 -3040
rect 1355 -3070 1400 -3040
rect 1280 -3110 1400 -3070
rect 1280 -3140 1325 -3110
rect 1355 -3140 1400 -3110
rect 1280 -3180 1400 -3140
rect 1280 -3210 1325 -3180
rect 1355 -3210 1400 -3180
rect 1280 -3245 1400 -3210
rect 1280 -3275 1325 -3245
rect 1355 -3275 1400 -3245
rect 1280 -3305 1400 -3275
rect 1280 -3335 1325 -3305
rect 1355 -3335 1400 -3305
rect 1280 -3370 1400 -3335
rect 1280 -3400 1325 -3370
rect 1355 -3400 1400 -3370
rect 1280 -3440 1400 -3400
rect 1280 -3470 1325 -3440
rect 1355 -3470 1400 -3440
rect 1280 -3510 1400 -3470
rect 1280 -3540 1325 -3510
rect 1355 -3540 1400 -3510
rect 1280 -3580 1400 -3540
rect 1280 -3610 1325 -3580
rect 1355 -3610 1400 -3580
rect 1280 -3645 1400 -3610
rect 1280 -3675 1325 -3645
rect 1355 -3675 1400 -3645
rect 1280 -3705 1400 -3675
rect 1280 -3735 1325 -3705
rect 1355 -3735 1400 -3705
rect 1280 -3770 1400 -3735
rect 1280 -3800 1325 -3770
rect 1355 -3800 1400 -3770
rect 1280 -3840 1400 -3800
rect 1280 -3870 1325 -3840
rect 1355 -3870 1400 -3840
rect 1280 -3910 1400 -3870
rect 1280 -3940 1325 -3910
rect 1355 -3940 1400 -3910
rect 1280 -3980 1400 -3940
rect 1280 -4010 1325 -3980
rect 1355 -4010 1400 -3980
rect 1280 -4045 1400 -4010
rect 1280 -4075 1325 -4045
rect 1355 -4075 1400 -4045
rect 1280 -4105 1400 -4075
rect 1280 -4135 1325 -4105
rect 1355 -4135 1400 -4105
rect 1280 -4170 1400 -4135
rect 1280 -4200 1325 -4170
rect 1355 -4200 1400 -4170
rect 1280 -4240 1400 -4200
rect 1280 -4270 1325 -4240
rect 1355 -4270 1400 -4240
rect 1280 -4310 1400 -4270
rect 1280 -4340 1325 -4310
rect 1355 -4340 1400 -4310
rect 1280 -4380 1400 -4340
rect 1280 -4410 1325 -4380
rect 1355 -4410 1400 -4380
rect 1280 -4445 1400 -4410
rect 1280 -4475 1325 -4445
rect 1355 -4475 1400 -4445
rect 1280 -4490 1400 -4475
rect 1630 -1305 1750 -1240
rect 1630 -1335 1675 -1305
rect 1705 -1335 1750 -1305
rect 1630 -1370 1750 -1335
rect 1630 -1400 1675 -1370
rect 1705 -1400 1750 -1370
rect 1630 -1440 1750 -1400
rect 1630 -1470 1675 -1440
rect 1705 -1470 1750 -1440
rect 1630 -1510 1750 -1470
rect 1630 -1540 1675 -1510
rect 1705 -1540 1750 -1510
rect 1630 -1580 1750 -1540
rect 1630 -1610 1675 -1580
rect 1705 -1610 1750 -1580
rect 1630 -1645 1750 -1610
rect 1630 -1675 1675 -1645
rect 1705 -1675 1750 -1645
rect 1630 -1705 1750 -1675
rect 1630 -1735 1675 -1705
rect 1705 -1735 1750 -1705
rect 1630 -1770 1750 -1735
rect 1630 -1800 1675 -1770
rect 1705 -1800 1750 -1770
rect 1630 -1840 1750 -1800
rect 1630 -1870 1675 -1840
rect 1705 -1870 1750 -1840
rect 1630 -1910 1750 -1870
rect 1630 -1940 1675 -1910
rect 1705 -1940 1750 -1910
rect 1630 -1980 1750 -1940
rect 1630 -2010 1675 -1980
rect 1705 -2010 1750 -1980
rect 1630 -2045 1750 -2010
rect 1630 -2075 1675 -2045
rect 1705 -2075 1750 -2045
rect 1630 -2105 1750 -2075
rect 1630 -2135 1675 -2105
rect 1705 -2135 1750 -2105
rect 1630 -2170 1750 -2135
rect 1630 -2200 1675 -2170
rect 1705 -2200 1750 -2170
rect 1630 -2240 1750 -2200
rect 1630 -2270 1675 -2240
rect 1705 -2270 1750 -2240
rect 1630 -2310 1750 -2270
rect 1630 -2340 1675 -2310
rect 1705 -2340 1750 -2310
rect 1630 -2380 1750 -2340
rect 1630 -2410 1675 -2380
rect 1705 -2410 1750 -2380
rect 1630 -2445 1750 -2410
rect 1630 -2475 1675 -2445
rect 1705 -2475 1750 -2445
rect 1630 -2505 1750 -2475
rect 1630 -2535 1675 -2505
rect 1705 -2535 1750 -2505
rect 1630 -2570 1750 -2535
rect 1630 -2600 1675 -2570
rect 1705 -2600 1750 -2570
rect 1630 -2640 1750 -2600
rect 1630 -2670 1675 -2640
rect 1705 -2670 1750 -2640
rect 1630 -2710 1750 -2670
rect 1630 -2740 1675 -2710
rect 1705 -2740 1750 -2710
rect 1630 -2780 1750 -2740
rect 1630 -2810 1675 -2780
rect 1705 -2810 1750 -2780
rect 1630 -2845 1750 -2810
rect 1630 -2875 1675 -2845
rect 1705 -2875 1750 -2845
rect 1630 -2905 1750 -2875
rect 1630 -2935 1675 -2905
rect 1705 -2935 1750 -2905
rect 1630 -2970 1750 -2935
rect 1630 -3000 1675 -2970
rect 1705 -3000 1750 -2970
rect 1630 -3040 1750 -3000
rect 1630 -3070 1675 -3040
rect 1705 -3070 1750 -3040
rect 1630 -3110 1750 -3070
rect 1630 -3140 1675 -3110
rect 1705 -3140 1750 -3110
rect 1630 -3180 1750 -3140
rect 1630 -3210 1675 -3180
rect 1705 -3210 1750 -3180
rect 1630 -3245 1750 -3210
rect 1630 -3275 1675 -3245
rect 1705 -3275 1750 -3245
rect 1630 -3305 1750 -3275
rect 1630 -3335 1675 -3305
rect 1705 -3335 1750 -3305
rect 1630 -3370 1750 -3335
rect 1630 -3400 1675 -3370
rect 1705 -3400 1750 -3370
rect 1630 -3440 1750 -3400
rect 1630 -3470 1675 -3440
rect 1705 -3470 1750 -3440
rect 1630 -3510 1750 -3470
rect 1630 -3540 1675 -3510
rect 1705 -3540 1750 -3510
rect 1630 -3580 1750 -3540
rect 1630 -3610 1675 -3580
rect 1705 -3610 1750 -3580
rect 1630 -3645 1750 -3610
rect 1630 -3675 1675 -3645
rect 1705 -3675 1750 -3645
rect 1630 -3705 1750 -3675
rect 1630 -3735 1675 -3705
rect 1705 -3735 1750 -3705
rect 1630 -3770 1750 -3735
rect 1630 -3800 1675 -3770
rect 1705 -3800 1750 -3770
rect 1630 -3840 1750 -3800
rect 1630 -3870 1675 -3840
rect 1705 -3870 1750 -3840
rect 1630 -3910 1750 -3870
rect 1630 -3940 1675 -3910
rect 1705 -3940 1750 -3910
rect 1630 -3980 1750 -3940
rect 1630 -4010 1675 -3980
rect 1705 -4010 1750 -3980
rect 1630 -4045 1750 -4010
rect 1630 -4075 1675 -4045
rect 1705 -4075 1750 -4045
rect 1630 -4105 1750 -4075
rect 1630 -4135 1675 -4105
rect 1705 -4135 1750 -4105
rect 1630 -4170 1750 -4135
rect 1630 -4200 1675 -4170
rect 1705 -4200 1750 -4170
rect 1630 -4240 1750 -4200
rect 1630 -4270 1675 -4240
rect 1705 -4270 1750 -4240
rect 1630 -4310 1750 -4270
rect 1630 -4340 1675 -4310
rect 1705 -4340 1750 -4310
rect 1630 -4380 1750 -4340
rect 1630 -4410 1675 -4380
rect 1705 -4410 1750 -4380
rect 1630 -4445 1750 -4410
rect 1630 -4475 1675 -4445
rect 1705 -4475 1750 -4445
rect 1630 -4490 1750 -4475
rect 1980 -1305 2100 -1240
rect 1980 -1335 2025 -1305
rect 2055 -1335 2100 -1305
rect 1980 -1370 2100 -1335
rect 1980 -1400 2025 -1370
rect 2055 -1400 2100 -1370
rect 1980 -1440 2100 -1400
rect 1980 -1470 2025 -1440
rect 2055 -1470 2100 -1440
rect 1980 -1510 2100 -1470
rect 1980 -1540 2025 -1510
rect 2055 -1540 2100 -1510
rect 1980 -1580 2100 -1540
rect 1980 -1610 2025 -1580
rect 2055 -1610 2100 -1580
rect 1980 -1645 2100 -1610
rect 1980 -1675 2025 -1645
rect 2055 -1675 2100 -1645
rect 1980 -1705 2100 -1675
rect 1980 -1735 2025 -1705
rect 2055 -1735 2100 -1705
rect 1980 -1770 2100 -1735
rect 1980 -1800 2025 -1770
rect 2055 -1800 2100 -1770
rect 1980 -1840 2100 -1800
rect 1980 -1870 2025 -1840
rect 2055 -1870 2100 -1840
rect 1980 -1910 2100 -1870
rect 1980 -1940 2025 -1910
rect 2055 -1940 2100 -1910
rect 1980 -1980 2100 -1940
rect 1980 -2010 2025 -1980
rect 2055 -2010 2100 -1980
rect 1980 -2045 2100 -2010
rect 1980 -2075 2025 -2045
rect 2055 -2075 2100 -2045
rect 1980 -2105 2100 -2075
rect 1980 -2135 2025 -2105
rect 2055 -2135 2100 -2105
rect 1980 -2170 2100 -2135
rect 1980 -2200 2025 -2170
rect 2055 -2200 2100 -2170
rect 1980 -2240 2100 -2200
rect 1980 -2270 2025 -2240
rect 2055 -2270 2100 -2240
rect 1980 -2310 2100 -2270
rect 1980 -2340 2025 -2310
rect 2055 -2340 2100 -2310
rect 1980 -2380 2100 -2340
rect 1980 -2410 2025 -2380
rect 2055 -2410 2100 -2380
rect 1980 -2445 2100 -2410
rect 1980 -2475 2025 -2445
rect 2055 -2475 2100 -2445
rect 1980 -2505 2100 -2475
rect 1980 -2535 2025 -2505
rect 2055 -2535 2100 -2505
rect 1980 -2570 2100 -2535
rect 1980 -2600 2025 -2570
rect 2055 -2600 2100 -2570
rect 1980 -2640 2100 -2600
rect 1980 -2670 2025 -2640
rect 2055 -2670 2100 -2640
rect 1980 -2710 2100 -2670
rect 1980 -2740 2025 -2710
rect 2055 -2740 2100 -2710
rect 1980 -2780 2100 -2740
rect 1980 -2810 2025 -2780
rect 2055 -2810 2100 -2780
rect 1980 -2845 2100 -2810
rect 1980 -2875 2025 -2845
rect 2055 -2875 2100 -2845
rect 1980 -2905 2100 -2875
rect 1980 -2935 2025 -2905
rect 2055 -2935 2100 -2905
rect 1980 -2970 2100 -2935
rect 1980 -3000 2025 -2970
rect 2055 -3000 2100 -2970
rect 1980 -3040 2100 -3000
rect 1980 -3070 2025 -3040
rect 2055 -3070 2100 -3040
rect 1980 -3110 2100 -3070
rect 1980 -3140 2025 -3110
rect 2055 -3140 2100 -3110
rect 1980 -3180 2100 -3140
rect 1980 -3210 2025 -3180
rect 2055 -3210 2100 -3180
rect 1980 -3245 2100 -3210
rect 1980 -3275 2025 -3245
rect 2055 -3275 2100 -3245
rect 1980 -3305 2100 -3275
rect 1980 -3335 2025 -3305
rect 2055 -3335 2100 -3305
rect 1980 -3370 2100 -3335
rect 1980 -3400 2025 -3370
rect 2055 -3400 2100 -3370
rect 1980 -3440 2100 -3400
rect 1980 -3470 2025 -3440
rect 2055 -3470 2100 -3440
rect 1980 -3510 2100 -3470
rect 1980 -3540 2025 -3510
rect 2055 -3540 2100 -3510
rect 1980 -3580 2100 -3540
rect 1980 -3610 2025 -3580
rect 2055 -3610 2100 -3580
rect 1980 -3645 2100 -3610
rect 1980 -3675 2025 -3645
rect 2055 -3675 2100 -3645
rect 1980 -3705 2100 -3675
rect 1980 -3735 2025 -3705
rect 2055 -3735 2100 -3705
rect 1980 -3770 2100 -3735
rect 1980 -3800 2025 -3770
rect 2055 -3800 2100 -3770
rect 1980 -3840 2100 -3800
rect 1980 -3870 2025 -3840
rect 2055 -3870 2100 -3840
rect 1980 -3910 2100 -3870
rect 1980 -3940 2025 -3910
rect 2055 -3940 2100 -3910
rect 1980 -3980 2100 -3940
rect 1980 -4010 2025 -3980
rect 2055 -4010 2100 -3980
rect 1980 -4045 2100 -4010
rect 1980 -4075 2025 -4045
rect 2055 -4075 2100 -4045
rect 1980 -4105 2100 -4075
rect 1980 -4135 2025 -4105
rect 2055 -4135 2100 -4105
rect 1980 -4170 2100 -4135
rect 1980 -4200 2025 -4170
rect 2055 -4200 2100 -4170
rect 1980 -4240 2100 -4200
rect 1980 -4270 2025 -4240
rect 2055 -4270 2100 -4240
rect 1980 -4310 2100 -4270
rect 1980 -4340 2025 -4310
rect 2055 -4340 2100 -4310
rect 1980 -4380 2100 -4340
rect 1980 -4410 2025 -4380
rect 2055 -4410 2100 -4380
rect 1980 -4445 2100 -4410
rect 1980 -4475 2025 -4445
rect 2055 -4475 2100 -4445
rect 1980 -4490 2100 -4475
rect 2330 -1305 2450 -1240
rect 2330 -1335 2375 -1305
rect 2405 -1335 2450 -1305
rect 2330 -1370 2450 -1335
rect 2330 -1400 2375 -1370
rect 2405 -1400 2450 -1370
rect 2330 -1440 2450 -1400
rect 2330 -1470 2375 -1440
rect 2405 -1470 2450 -1440
rect 2330 -1510 2450 -1470
rect 2330 -1540 2375 -1510
rect 2405 -1540 2450 -1510
rect 2330 -1580 2450 -1540
rect 2330 -1610 2375 -1580
rect 2405 -1610 2450 -1580
rect 2330 -1645 2450 -1610
rect 2330 -1675 2375 -1645
rect 2405 -1675 2450 -1645
rect 2330 -1705 2450 -1675
rect 2330 -1735 2375 -1705
rect 2405 -1735 2450 -1705
rect 2330 -1770 2450 -1735
rect 2330 -1800 2375 -1770
rect 2405 -1800 2450 -1770
rect 2330 -1840 2450 -1800
rect 2330 -1870 2375 -1840
rect 2405 -1870 2450 -1840
rect 2330 -1910 2450 -1870
rect 2330 -1940 2375 -1910
rect 2405 -1940 2450 -1910
rect 2330 -1980 2450 -1940
rect 2330 -2010 2375 -1980
rect 2405 -2010 2450 -1980
rect 2330 -2045 2450 -2010
rect 2330 -2075 2375 -2045
rect 2405 -2075 2450 -2045
rect 2330 -2105 2450 -2075
rect 2330 -2135 2375 -2105
rect 2405 -2135 2450 -2105
rect 2330 -2170 2450 -2135
rect 2330 -2200 2375 -2170
rect 2405 -2200 2450 -2170
rect 2330 -2240 2450 -2200
rect 2330 -2270 2375 -2240
rect 2405 -2270 2450 -2240
rect 2330 -2310 2450 -2270
rect 2330 -2340 2375 -2310
rect 2405 -2340 2450 -2310
rect 2330 -2380 2450 -2340
rect 2330 -2410 2375 -2380
rect 2405 -2410 2450 -2380
rect 2330 -2445 2450 -2410
rect 2330 -2475 2375 -2445
rect 2405 -2475 2450 -2445
rect 2330 -2505 2450 -2475
rect 2330 -2535 2375 -2505
rect 2405 -2535 2450 -2505
rect 2330 -2570 2450 -2535
rect 2330 -2600 2375 -2570
rect 2405 -2600 2450 -2570
rect 2330 -2640 2450 -2600
rect 2330 -2670 2375 -2640
rect 2405 -2670 2450 -2640
rect 2330 -2710 2450 -2670
rect 2330 -2740 2375 -2710
rect 2405 -2740 2450 -2710
rect 2330 -2780 2450 -2740
rect 2330 -2810 2375 -2780
rect 2405 -2810 2450 -2780
rect 2330 -2845 2450 -2810
rect 2330 -2875 2375 -2845
rect 2405 -2875 2450 -2845
rect 2330 -2905 2450 -2875
rect 2330 -2935 2375 -2905
rect 2405 -2935 2450 -2905
rect 2330 -2970 2450 -2935
rect 2330 -3000 2375 -2970
rect 2405 -3000 2450 -2970
rect 2330 -3040 2450 -3000
rect 2330 -3070 2375 -3040
rect 2405 -3070 2450 -3040
rect 2330 -3110 2450 -3070
rect 2330 -3140 2375 -3110
rect 2405 -3140 2450 -3110
rect 2330 -3180 2450 -3140
rect 2330 -3210 2375 -3180
rect 2405 -3210 2450 -3180
rect 2330 -3245 2450 -3210
rect 2330 -3275 2375 -3245
rect 2405 -3275 2450 -3245
rect 2330 -3305 2450 -3275
rect 2330 -3335 2375 -3305
rect 2405 -3335 2450 -3305
rect 2330 -3370 2450 -3335
rect 2330 -3400 2375 -3370
rect 2405 -3400 2450 -3370
rect 2330 -3440 2450 -3400
rect 2330 -3470 2375 -3440
rect 2405 -3470 2450 -3440
rect 2330 -3510 2450 -3470
rect 2330 -3540 2375 -3510
rect 2405 -3540 2450 -3510
rect 2330 -3580 2450 -3540
rect 2330 -3610 2375 -3580
rect 2405 -3610 2450 -3580
rect 2330 -3645 2450 -3610
rect 2330 -3675 2375 -3645
rect 2405 -3675 2450 -3645
rect 2330 -3705 2450 -3675
rect 2330 -3735 2375 -3705
rect 2405 -3735 2450 -3705
rect 2330 -3770 2450 -3735
rect 2330 -3800 2375 -3770
rect 2405 -3800 2450 -3770
rect 2330 -3840 2450 -3800
rect 2330 -3870 2375 -3840
rect 2405 -3870 2450 -3840
rect 2330 -3910 2450 -3870
rect 2330 -3940 2375 -3910
rect 2405 -3940 2450 -3910
rect 2330 -3980 2450 -3940
rect 2330 -4010 2375 -3980
rect 2405 -4010 2450 -3980
rect 2330 -4045 2450 -4010
rect 2330 -4075 2375 -4045
rect 2405 -4075 2450 -4045
rect 2330 -4105 2450 -4075
rect 2330 -4135 2375 -4105
rect 2405 -4135 2450 -4105
rect 2330 -4170 2450 -4135
rect 2330 -4200 2375 -4170
rect 2405 -4200 2450 -4170
rect 2330 -4240 2450 -4200
rect 2330 -4270 2375 -4240
rect 2405 -4270 2450 -4240
rect 2330 -4310 2450 -4270
rect 2330 -4340 2375 -4310
rect 2405 -4340 2450 -4310
rect 2330 -4380 2450 -4340
rect 2330 -4410 2375 -4380
rect 2405 -4410 2450 -4380
rect 2330 -4445 2450 -4410
rect 2330 -4475 2375 -4445
rect 2405 -4475 2450 -4445
rect 2330 -4490 2450 -4475
rect 2680 -1305 2800 -1240
rect 2680 -1335 2725 -1305
rect 2755 -1335 2800 -1305
rect 2680 -1370 2800 -1335
rect 2680 -1400 2725 -1370
rect 2755 -1400 2800 -1370
rect 2680 -1440 2800 -1400
rect 2680 -1470 2725 -1440
rect 2755 -1470 2800 -1440
rect 2680 -1510 2800 -1470
rect 2680 -1540 2725 -1510
rect 2755 -1540 2800 -1510
rect 2680 -1580 2800 -1540
rect 2680 -1610 2725 -1580
rect 2755 -1610 2800 -1580
rect 2680 -1645 2800 -1610
rect 2680 -1675 2725 -1645
rect 2755 -1675 2800 -1645
rect 2680 -1705 2800 -1675
rect 2680 -1735 2725 -1705
rect 2755 -1735 2800 -1705
rect 2680 -1770 2800 -1735
rect 2680 -1800 2725 -1770
rect 2755 -1800 2800 -1770
rect 2680 -1840 2800 -1800
rect 2680 -1870 2725 -1840
rect 2755 -1870 2800 -1840
rect 2680 -1910 2800 -1870
rect 2680 -1940 2725 -1910
rect 2755 -1940 2800 -1910
rect 2680 -1980 2800 -1940
rect 2680 -2010 2725 -1980
rect 2755 -2010 2800 -1980
rect 2680 -2045 2800 -2010
rect 2680 -2075 2725 -2045
rect 2755 -2075 2800 -2045
rect 2680 -2105 2800 -2075
rect 2680 -2135 2725 -2105
rect 2755 -2135 2800 -2105
rect 2680 -2170 2800 -2135
rect 2680 -2200 2725 -2170
rect 2755 -2200 2800 -2170
rect 2680 -2240 2800 -2200
rect 2680 -2270 2725 -2240
rect 2755 -2270 2800 -2240
rect 2680 -2310 2800 -2270
rect 2680 -2340 2725 -2310
rect 2755 -2340 2800 -2310
rect 2680 -2380 2800 -2340
rect 2680 -2410 2725 -2380
rect 2755 -2410 2800 -2380
rect 2680 -2445 2800 -2410
rect 2680 -2475 2725 -2445
rect 2755 -2475 2800 -2445
rect 2680 -2505 2800 -2475
rect 2680 -2535 2725 -2505
rect 2755 -2535 2800 -2505
rect 2680 -2570 2800 -2535
rect 2680 -2600 2725 -2570
rect 2755 -2600 2800 -2570
rect 2680 -2640 2800 -2600
rect 2680 -2670 2725 -2640
rect 2755 -2670 2800 -2640
rect 2680 -2710 2800 -2670
rect 2680 -2740 2725 -2710
rect 2755 -2740 2800 -2710
rect 2680 -2780 2800 -2740
rect 2680 -2810 2725 -2780
rect 2755 -2810 2800 -2780
rect 2680 -2845 2800 -2810
rect 2680 -2875 2725 -2845
rect 2755 -2875 2800 -2845
rect 2680 -2905 2800 -2875
rect 2680 -2935 2725 -2905
rect 2755 -2935 2800 -2905
rect 2680 -2970 2800 -2935
rect 2680 -3000 2725 -2970
rect 2755 -3000 2800 -2970
rect 2680 -3040 2800 -3000
rect 2680 -3070 2725 -3040
rect 2755 -3070 2800 -3040
rect 2680 -3110 2800 -3070
rect 2680 -3140 2725 -3110
rect 2755 -3140 2800 -3110
rect 2680 -3180 2800 -3140
rect 2680 -3210 2725 -3180
rect 2755 -3210 2800 -3180
rect 2680 -3245 2800 -3210
rect 2680 -3275 2725 -3245
rect 2755 -3275 2800 -3245
rect 2680 -3305 2800 -3275
rect 2680 -3335 2725 -3305
rect 2755 -3335 2800 -3305
rect 2680 -3370 2800 -3335
rect 2680 -3400 2725 -3370
rect 2755 -3400 2800 -3370
rect 2680 -3440 2800 -3400
rect 2680 -3470 2725 -3440
rect 2755 -3470 2800 -3440
rect 2680 -3510 2800 -3470
rect 2680 -3540 2725 -3510
rect 2755 -3540 2800 -3510
rect 2680 -3580 2800 -3540
rect 2680 -3610 2725 -3580
rect 2755 -3610 2800 -3580
rect 2680 -3645 2800 -3610
rect 2680 -3675 2725 -3645
rect 2755 -3675 2800 -3645
rect 2680 -3705 2800 -3675
rect 2680 -3735 2725 -3705
rect 2755 -3735 2800 -3705
rect 2680 -3770 2800 -3735
rect 2680 -3800 2725 -3770
rect 2755 -3800 2800 -3770
rect 2680 -3840 2800 -3800
rect 2680 -3870 2725 -3840
rect 2755 -3870 2800 -3840
rect 2680 -3910 2800 -3870
rect 2680 -3940 2725 -3910
rect 2755 -3940 2800 -3910
rect 2680 -3980 2800 -3940
rect 2680 -4010 2725 -3980
rect 2755 -4010 2800 -3980
rect 2680 -4045 2800 -4010
rect 2680 -4075 2725 -4045
rect 2755 -4075 2800 -4045
rect 2680 -4105 2800 -4075
rect 2680 -4135 2725 -4105
rect 2755 -4135 2800 -4105
rect 2680 -4170 2800 -4135
rect 2680 -4200 2725 -4170
rect 2755 -4200 2800 -4170
rect 2680 -4240 2800 -4200
rect 2680 -4270 2725 -4240
rect 2755 -4270 2800 -4240
rect 2680 -4310 2800 -4270
rect 2680 -4340 2725 -4310
rect 2755 -4340 2800 -4310
rect 2680 -4380 2800 -4340
rect 2680 -4410 2725 -4380
rect 2755 -4410 2800 -4380
rect 2680 -4445 2800 -4410
rect 2680 -4475 2725 -4445
rect 2755 -4475 2800 -4445
rect 2680 -4490 2800 -4475
rect 3030 -1305 3150 -1240
rect 3030 -1335 3075 -1305
rect 3105 -1335 3150 -1305
rect 3030 -1370 3150 -1335
rect 3030 -1400 3075 -1370
rect 3105 -1400 3150 -1370
rect 3030 -1440 3150 -1400
rect 3030 -1470 3075 -1440
rect 3105 -1470 3150 -1440
rect 3030 -1510 3150 -1470
rect 3030 -1540 3075 -1510
rect 3105 -1540 3150 -1510
rect 3030 -1580 3150 -1540
rect 3030 -1610 3075 -1580
rect 3105 -1610 3150 -1580
rect 3030 -1645 3150 -1610
rect 3030 -1675 3075 -1645
rect 3105 -1675 3150 -1645
rect 3030 -1705 3150 -1675
rect 3030 -1735 3075 -1705
rect 3105 -1735 3150 -1705
rect 3030 -1770 3150 -1735
rect 3030 -1800 3075 -1770
rect 3105 -1800 3150 -1770
rect 3030 -1840 3150 -1800
rect 3030 -1870 3075 -1840
rect 3105 -1870 3150 -1840
rect 3030 -1910 3150 -1870
rect 3030 -1940 3075 -1910
rect 3105 -1940 3150 -1910
rect 3030 -1980 3150 -1940
rect 3030 -2010 3075 -1980
rect 3105 -2010 3150 -1980
rect 3030 -2045 3150 -2010
rect 3030 -2075 3075 -2045
rect 3105 -2075 3150 -2045
rect 3030 -2105 3150 -2075
rect 3030 -2135 3075 -2105
rect 3105 -2135 3150 -2105
rect 3030 -2170 3150 -2135
rect 3030 -2200 3075 -2170
rect 3105 -2200 3150 -2170
rect 3030 -2240 3150 -2200
rect 3030 -2270 3075 -2240
rect 3105 -2270 3150 -2240
rect 3030 -2310 3150 -2270
rect 3030 -2340 3075 -2310
rect 3105 -2340 3150 -2310
rect 3030 -2380 3150 -2340
rect 3030 -2410 3075 -2380
rect 3105 -2410 3150 -2380
rect 3030 -2445 3150 -2410
rect 3030 -2475 3075 -2445
rect 3105 -2475 3150 -2445
rect 3030 -2505 3150 -2475
rect 3030 -2535 3075 -2505
rect 3105 -2535 3150 -2505
rect 3030 -2570 3150 -2535
rect 3030 -2600 3075 -2570
rect 3105 -2600 3150 -2570
rect 3030 -2640 3150 -2600
rect 3030 -2670 3075 -2640
rect 3105 -2670 3150 -2640
rect 3030 -2710 3150 -2670
rect 3030 -2740 3075 -2710
rect 3105 -2740 3150 -2710
rect 3030 -2780 3150 -2740
rect 3030 -2810 3075 -2780
rect 3105 -2810 3150 -2780
rect 3030 -2845 3150 -2810
rect 3030 -2875 3075 -2845
rect 3105 -2875 3150 -2845
rect 3030 -2905 3150 -2875
rect 3030 -2935 3075 -2905
rect 3105 -2935 3150 -2905
rect 3030 -2970 3150 -2935
rect 3030 -3000 3075 -2970
rect 3105 -3000 3150 -2970
rect 3030 -3040 3150 -3000
rect 3030 -3070 3075 -3040
rect 3105 -3070 3150 -3040
rect 3030 -3110 3150 -3070
rect 3030 -3140 3075 -3110
rect 3105 -3140 3150 -3110
rect 3030 -3180 3150 -3140
rect 3030 -3210 3075 -3180
rect 3105 -3210 3150 -3180
rect 3030 -3245 3150 -3210
rect 3030 -3275 3075 -3245
rect 3105 -3275 3150 -3245
rect 3030 -3305 3150 -3275
rect 3030 -3335 3075 -3305
rect 3105 -3335 3150 -3305
rect 3030 -3370 3150 -3335
rect 3030 -3400 3075 -3370
rect 3105 -3400 3150 -3370
rect 3030 -3440 3150 -3400
rect 3030 -3470 3075 -3440
rect 3105 -3470 3150 -3440
rect 3030 -3510 3150 -3470
rect 3030 -3540 3075 -3510
rect 3105 -3540 3150 -3510
rect 3030 -3580 3150 -3540
rect 3030 -3610 3075 -3580
rect 3105 -3610 3150 -3580
rect 3030 -3645 3150 -3610
rect 3030 -3675 3075 -3645
rect 3105 -3675 3150 -3645
rect 3030 -3705 3150 -3675
rect 3030 -3735 3075 -3705
rect 3105 -3735 3150 -3705
rect 3030 -3770 3150 -3735
rect 3030 -3800 3075 -3770
rect 3105 -3800 3150 -3770
rect 3030 -3840 3150 -3800
rect 3030 -3870 3075 -3840
rect 3105 -3870 3150 -3840
rect 3030 -3910 3150 -3870
rect 3030 -3940 3075 -3910
rect 3105 -3940 3150 -3910
rect 3030 -3980 3150 -3940
rect 3030 -4010 3075 -3980
rect 3105 -4010 3150 -3980
rect 3030 -4045 3150 -4010
rect 3030 -4075 3075 -4045
rect 3105 -4075 3150 -4045
rect 3030 -4105 3150 -4075
rect 3030 -4135 3075 -4105
rect 3105 -4135 3150 -4105
rect 3030 -4170 3150 -4135
rect 3030 -4200 3075 -4170
rect 3105 -4200 3150 -4170
rect 3030 -4240 3150 -4200
rect 3030 -4270 3075 -4240
rect 3105 -4270 3150 -4240
rect 3030 -4310 3150 -4270
rect 3030 -4340 3075 -4310
rect 3105 -4340 3150 -4310
rect 3030 -4380 3150 -4340
rect 3030 -4410 3075 -4380
rect 3105 -4410 3150 -4380
rect 3030 -4445 3150 -4410
rect 3030 -4475 3075 -4445
rect 3105 -4475 3150 -4445
rect 3030 -4490 3150 -4475
rect 3380 -1305 3500 -1240
rect 3380 -1335 3425 -1305
rect 3455 -1335 3500 -1305
rect 3380 -1370 3500 -1335
rect 3380 -1400 3425 -1370
rect 3455 -1400 3500 -1370
rect 3380 -1440 3500 -1400
rect 3380 -1470 3425 -1440
rect 3455 -1470 3500 -1440
rect 3380 -1510 3500 -1470
rect 3380 -1540 3425 -1510
rect 3455 -1540 3500 -1510
rect 3380 -1580 3500 -1540
rect 3380 -1610 3425 -1580
rect 3455 -1610 3500 -1580
rect 3380 -1645 3500 -1610
rect 3380 -1675 3425 -1645
rect 3455 -1675 3500 -1645
rect 3380 -1705 3500 -1675
rect 3380 -1735 3425 -1705
rect 3455 -1735 3500 -1705
rect 3380 -1770 3500 -1735
rect 3380 -1800 3425 -1770
rect 3455 -1800 3500 -1770
rect 3380 -1840 3500 -1800
rect 3380 -1870 3425 -1840
rect 3455 -1870 3500 -1840
rect 3380 -1910 3500 -1870
rect 3380 -1940 3425 -1910
rect 3455 -1940 3500 -1910
rect 3380 -1980 3500 -1940
rect 3380 -2010 3425 -1980
rect 3455 -2010 3500 -1980
rect 3380 -2045 3500 -2010
rect 3380 -2075 3425 -2045
rect 3455 -2075 3500 -2045
rect 3380 -2105 3500 -2075
rect 3380 -2135 3425 -2105
rect 3455 -2135 3500 -2105
rect 3380 -2170 3500 -2135
rect 3380 -2200 3425 -2170
rect 3455 -2200 3500 -2170
rect 3380 -2240 3500 -2200
rect 3380 -2270 3425 -2240
rect 3455 -2270 3500 -2240
rect 3380 -2310 3500 -2270
rect 3380 -2340 3425 -2310
rect 3455 -2340 3500 -2310
rect 3380 -2380 3500 -2340
rect 3380 -2410 3425 -2380
rect 3455 -2410 3500 -2380
rect 3380 -2445 3500 -2410
rect 3380 -2475 3425 -2445
rect 3455 -2475 3500 -2445
rect 3380 -2505 3500 -2475
rect 3380 -2535 3425 -2505
rect 3455 -2535 3500 -2505
rect 3380 -2570 3500 -2535
rect 3380 -2600 3425 -2570
rect 3455 -2600 3500 -2570
rect 3380 -2640 3500 -2600
rect 3380 -2670 3425 -2640
rect 3455 -2670 3500 -2640
rect 3380 -2710 3500 -2670
rect 3380 -2740 3425 -2710
rect 3455 -2740 3500 -2710
rect 3380 -2780 3500 -2740
rect 3380 -2810 3425 -2780
rect 3455 -2810 3500 -2780
rect 3380 -2845 3500 -2810
rect 3380 -2875 3425 -2845
rect 3455 -2875 3500 -2845
rect 3380 -2905 3500 -2875
rect 3380 -2935 3425 -2905
rect 3455 -2935 3500 -2905
rect 3380 -2970 3500 -2935
rect 3380 -3000 3425 -2970
rect 3455 -3000 3500 -2970
rect 3380 -3040 3500 -3000
rect 3380 -3070 3425 -3040
rect 3455 -3070 3500 -3040
rect 3380 -3110 3500 -3070
rect 3380 -3140 3425 -3110
rect 3455 -3140 3500 -3110
rect 3380 -3180 3500 -3140
rect 3380 -3210 3425 -3180
rect 3455 -3210 3500 -3180
rect 3380 -3245 3500 -3210
rect 3380 -3275 3425 -3245
rect 3455 -3275 3500 -3245
rect 3380 -3305 3500 -3275
rect 3380 -3335 3425 -3305
rect 3455 -3335 3500 -3305
rect 3380 -3370 3500 -3335
rect 3380 -3400 3425 -3370
rect 3455 -3400 3500 -3370
rect 3380 -3440 3500 -3400
rect 3380 -3470 3425 -3440
rect 3455 -3470 3500 -3440
rect 3380 -3510 3500 -3470
rect 3380 -3540 3425 -3510
rect 3455 -3540 3500 -3510
rect 3380 -3580 3500 -3540
rect 3380 -3610 3425 -3580
rect 3455 -3610 3500 -3580
rect 3380 -3645 3500 -3610
rect 3380 -3675 3425 -3645
rect 3455 -3675 3500 -3645
rect 3380 -3705 3500 -3675
rect 3380 -3735 3425 -3705
rect 3455 -3735 3500 -3705
rect 3380 -3770 3500 -3735
rect 3380 -3800 3425 -3770
rect 3455 -3800 3500 -3770
rect 3380 -3840 3500 -3800
rect 3380 -3870 3425 -3840
rect 3455 -3870 3500 -3840
rect 3380 -3910 3500 -3870
rect 3380 -3940 3425 -3910
rect 3455 -3940 3500 -3910
rect 3380 -3980 3500 -3940
rect 3380 -4010 3425 -3980
rect 3455 -4010 3500 -3980
rect 3380 -4045 3500 -4010
rect 3380 -4075 3425 -4045
rect 3455 -4075 3500 -4045
rect 3380 -4105 3500 -4075
rect 3380 -4135 3425 -4105
rect 3455 -4135 3500 -4105
rect 3380 -4170 3500 -4135
rect 3380 -4200 3425 -4170
rect 3455 -4200 3500 -4170
rect 3380 -4240 3500 -4200
rect 3380 -4270 3425 -4240
rect 3455 -4270 3500 -4240
rect 3380 -4310 3500 -4270
rect 3380 -4340 3425 -4310
rect 3455 -4340 3500 -4310
rect 3380 -4380 3500 -4340
rect 3380 -4410 3425 -4380
rect 3455 -4410 3500 -4380
rect 3380 -4445 3500 -4410
rect 3380 -4475 3425 -4445
rect 3455 -4475 3500 -4445
rect 3380 -4490 3500 -4475
rect 3730 -1305 3850 -1240
rect 3730 -1335 3775 -1305
rect 3805 -1335 3850 -1305
rect 3730 -1370 3850 -1335
rect 3730 -1400 3775 -1370
rect 3805 -1400 3850 -1370
rect 3730 -1440 3850 -1400
rect 3730 -1470 3775 -1440
rect 3805 -1470 3850 -1440
rect 3730 -1510 3850 -1470
rect 3730 -1540 3775 -1510
rect 3805 -1540 3850 -1510
rect 3730 -1580 3850 -1540
rect 3730 -1610 3775 -1580
rect 3805 -1610 3850 -1580
rect 3730 -1645 3850 -1610
rect 3730 -1675 3775 -1645
rect 3805 -1675 3850 -1645
rect 3730 -1705 3850 -1675
rect 3730 -1735 3775 -1705
rect 3805 -1735 3850 -1705
rect 3730 -1770 3850 -1735
rect 3730 -1800 3775 -1770
rect 3805 -1800 3850 -1770
rect 3730 -1840 3850 -1800
rect 3730 -1870 3775 -1840
rect 3805 -1870 3850 -1840
rect 3730 -1910 3850 -1870
rect 3730 -1940 3775 -1910
rect 3805 -1940 3850 -1910
rect 3730 -1980 3850 -1940
rect 3730 -2010 3775 -1980
rect 3805 -2010 3850 -1980
rect 3730 -2045 3850 -2010
rect 3730 -2075 3775 -2045
rect 3805 -2075 3850 -2045
rect 3730 -2105 3850 -2075
rect 3730 -2135 3775 -2105
rect 3805 -2135 3850 -2105
rect 3730 -2170 3850 -2135
rect 3730 -2200 3775 -2170
rect 3805 -2200 3850 -2170
rect 3730 -2240 3850 -2200
rect 3730 -2270 3775 -2240
rect 3805 -2270 3850 -2240
rect 3730 -2310 3850 -2270
rect 3730 -2340 3775 -2310
rect 3805 -2340 3850 -2310
rect 3730 -2380 3850 -2340
rect 3730 -2410 3775 -2380
rect 3805 -2410 3850 -2380
rect 3730 -2445 3850 -2410
rect 3730 -2475 3775 -2445
rect 3805 -2475 3850 -2445
rect 3730 -2505 3850 -2475
rect 3730 -2535 3775 -2505
rect 3805 -2535 3850 -2505
rect 3730 -2570 3850 -2535
rect 3730 -2600 3775 -2570
rect 3805 -2600 3850 -2570
rect 3730 -2640 3850 -2600
rect 3730 -2670 3775 -2640
rect 3805 -2670 3850 -2640
rect 3730 -2710 3850 -2670
rect 3730 -2740 3775 -2710
rect 3805 -2740 3850 -2710
rect 3730 -2780 3850 -2740
rect 3730 -2810 3775 -2780
rect 3805 -2810 3850 -2780
rect 3730 -2845 3850 -2810
rect 3730 -2875 3775 -2845
rect 3805 -2875 3850 -2845
rect 3730 -2905 3850 -2875
rect 3730 -2935 3775 -2905
rect 3805 -2935 3850 -2905
rect 3730 -2970 3850 -2935
rect 3730 -3000 3775 -2970
rect 3805 -3000 3850 -2970
rect 3730 -3040 3850 -3000
rect 3730 -3070 3775 -3040
rect 3805 -3070 3850 -3040
rect 3730 -3110 3850 -3070
rect 3730 -3140 3775 -3110
rect 3805 -3140 3850 -3110
rect 3730 -3180 3850 -3140
rect 3730 -3210 3775 -3180
rect 3805 -3210 3850 -3180
rect 3730 -3245 3850 -3210
rect 3730 -3275 3775 -3245
rect 3805 -3275 3850 -3245
rect 3730 -3305 3850 -3275
rect 3730 -3335 3775 -3305
rect 3805 -3335 3850 -3305
rect 3730 -3370 3850 -3335
rect 3730 -3400 3775 -3370
rect 3805 -3400 3850 -3370
rect 3730 -3440 3850 -3400
rect 3730 -3470 3775 -3440
rect 3805 -3470 3850 -3440
rect 3730 -3510 3850 -3470
rect 3730 -3540 3775 -3510
rect 3805 -3540 3850 -3510
rect 3730 -3580 3850 -3540
rect 3730 -3610 3775 -3580
rect 3805 -3610 3850 -3580
rect 3730 -3645 3850 -3610
rect 3730 -3675 3775 -3645
rect 3805 -3675 3850 -3645
rect 3730 -3705 3850 -3675
rect 3730 -3735 3775 -3705
rect 3805 -3735 3850 -3705
rect 3730 -3770 3850 -3735
rect 3730 -3800 3775 -3770
rect 3805 -3800 3850 -3770
rect 3730 -3840 3850 -3800
rect 3730 -3870 3775 -3840
rect 3805 -3870 3850 -3840
rect 3730 -3910 3850 -3870
rect 3730 -3940 3775 -3910
rect 3805 -3940 3850 -3910
rect 3730 -3980 3850 -3940
rect 3730 -4010 3775 -3980
rect 3805 -4010 3850 -3980
rect 3730 -4045 3850 -4010
rect 3730 -4075 3775 -4045
rect 3805 -4075 3850 -4045
rect 3730 -4105 3850 -4075
rect 3730 -4135 3775 -4105
rect 3805 -4135 3850 -4105
rect 3730 -4170 3850 -4135
rect 3730 -4200 3775 -4170
rect 3805 -4200 3850 -4170
rect 3730 -4240 3850 -4200
rect 3730 -4270 3775 -4240
rect 3805 -4270 3850 -4240
rect 3730 -4310 3850 -4270
rect 3730 -4340 3775 -4310
rect 3805 -4340 3850 -4310
rect 3730 -4380 3850 -4340
rect 3730 -4410 3775 -4380
rect 3805 -4410 3850 -4380
rect 3730 -4445 3850 -4410
rect 3730 -4475 3775 -4445
rect 3805 -4475 3850 -4445
rect 3730 -4490 3850 -4475
rect 4080 -1305 4200 -1240
rect 4080 -1335 4125 -1305
rect 4155 -1335 4200 -1305
rect 4080 -1370 4200 -1335
rect 4080 -1400 4125 -1370
rect 4155 -1400 4200 -1370
rect 4080 -1440 4200 -1400
rect 4080 -1470 4125 -1440
rect 4155 -1470 4200 -1440
rect 4080 -1510 4200 -1470
rect 4080 -1540 4125 -1510
rect 4155 -1540 4200 -1510
rect 4080 -1580 4200 -1540
rect 4080 -1610 4125 -1580
rect 4155 -1610 4200 -1580
rect 4080 -1645 4200 -1610
rect 4080 -1675 4125 -1645
rect 4155 -1675 4200 -1645
rect 4080 -1705 4200 -1675
rect 4080 -1735 4125 -1705
rect 4155 -1735 4200 -1705
rect 4080 -1770 4200 -1735
rect 4080 -1800 4125 -1770
rect 4155 -1800 4200 -1770
rect 4080 -1840 4200 -1800
rect 4080 -1870 4125 -1840
rect 4155 -1870 4200 -1840
rect 4080 -1910 4200 -1870
rect 4080 -1940 4125 -1910
rect 4155 -1940 4200 -1910
rect 4080 -1980 4200 -1940
rect 4080 -2010 4125 -1980
rect 4155 -2010 4200 -1980
rect 4080 -2045 4200 -2010
rect 4080 -2075 4125 -2045
rect 4155 -2075 4200 -2045
rect 4080 -2105 4200 -2075
rect 4080 -2135 4125 -2105
rect 4155 -2135 4200 -2105
rect 4080 -2170 4200 -2135
rect 4080 -2200 4125 -2170
rect 4155 -2200 4200 -2170
rect 4080 -2240 4200 -2200
rect 4080 -2270 4125 -2240
rect 4155 -2270 4200 -2240
rect 4080 -2310 4200 -2270
rect 4080 -2340 4125 -2310
rect 4155 -2340 4200 -2310
rect 4080 -2380 4200 -2340
rect 4080 -2410 4125 -2380
rect 4155 -2410 4200 -2380
rect 4080 -2445 4200 -2410
rect 4080 -2475 4125 -2445
rect 4155 -2475 4200 -2445
rect 4080 -2505 4200 -2475
rect 4080 -2535 4125 -2505
rect 4155 -2535 4200 -2505
rect 4080 -2570 4200 -2535
rect 4080 -2600 4125 -2570
rect 4155 -2600 4200 -2570
rect 4080 -2640 4200 -2600
rect 4080 -2670 4125 -2640
rect 4155 -2670 4200 -2640
rect 4080 -2710 4200 -2670
rect 4080 -2740 4125 -2710
rect 4155 -2740 4200 -2710
rect 4080 -2780 4200 -2740
rect 4080 -2810 4125 -2780
rect 4155 -2810 4200 -2780
rect 4080 -2845 4200 -2810
rect 4080 -2875 4125 -2845
rect 4155 -2875 4200 -2845
rect 4080 -2905 4200 -2875
rect 4080 -2935 4125 -2905
rect 4155 -2935 4200 -2905
rect 4080 -2970 4200 -2935
rect 4080 -3000 4125 -2970
rect 4155 -3000 4200 -2970
rect 4080 -3040 4200 -3000
rect 4080 -3070 4125 -3040
rect 4155 -3070 4200 -3040
rect 4080 -3110 4200 -3070
rect 4080 -3140 4125 -3110
rect 4155 -3140 4200 -3110
rect 4080 -3180 4200 -3140
rect 4080 -3210 4125 -3180
rect 4155 -3210 4200 -3180
rect 4080 -3245 4200 -3210
rect 4080 -3275 4125 -3245
rect 4155 -3275 4200 -3245
rect 4080 -3305 4200 -3275
rect 4080 -3335 4125 -3305
rect 4155 -3335 4200 -3305
rect 4080 -3370 4200 -3335
rect 4080 -3400 4125 -3370
rect 4155 -3400 4200 -3370
rect 4080 -3440 4200 -3400
rect 4080 -3470 4125 -3440
rect 4155 -3470 4200 -3440
rect 4080 -3510 4200 -3470
rect 4080 -3540 4125 -3510
rect 4155 -3540 4200 -3510
rect 4080 -3580 4200 -3540
rect 4080 -3610 4125 -3580
rect 4155 -3610 4200 -3580
rect 4080 -3645 4200 -3610
rect 4080 -3675 4125 -3645
rect 4155 -3675 4200 -3645
rect 4080 -3705 4200 -3675
rect 4080 -3735 4125 -3705
rect 4155 -3735 4200 -3705
rect 4080 -3770 4200 -3735
rect 4080 -3800 4125 -3770
rect 4155 -3800 4200 -3770
rect 4080 -3840 4200 -3800
rect 4080 -3870 4125 -3840
rect 4155 -3870 4200 -3840
rect 4080 -3910 4200 -3870
rect 4080 -3940 4125 -3910
rect 4155 -3940 4200 -3910
rect 4080 -3980 4200 -3940
rect 4080 -4010 4125 -3980
rect 4155 -4010 4200 -3980
rect 4080 -4045 4200 -4010
rect 4080 -4075 4125 -4045
rect 4155 -4075 4200 -4045
rect 4080 -4105 4200 -4075
rect 4080 -4135 4125 -4105
rect 4155 -4135 4200 -4105
rect 4080 -4170 4200 -4135
rect 4080 -4200 4125 -4170
rect 4155 -4200 4200 -4170
rect 4080 -4240 4200 -4200
rect 4080 -4270 4125 -4240
rect 4155 -4270 4200 -4240
rect 4080 -4310 4200 -4270
rect 4080 -4340 4125 -4310
rect 4155 -4340 4200 -4310
rect 4080 -4380 4200 -4340
rect 4080 -4410 4125 -4380
rect 4155 -4410 4200 -4380
rect 4080 -4445 4200 -4410
rect 4080 -4475 4125 -4445
rect 4155 -4475 4200 -4445
rect 4080 -4490 4200 -4475
rect 4430 -1305 4550 -1240
rect 4430 -1335 4475 -1305
rect 4505 -1335 4550 -1305
rect 4430 -1370 4550 -1335
rect 4430 -1400 4475 -1370
rect 4505 -1400 4550 -1370
rect 4430 -1440 4550 -1400
rect 4430 -1470 4475 -1440
rect 4505 -1470 4550 -1440
rect 4430 -1510 4550 -1470
rect 4430 -1540 4475 -1510
rect 4505 -1540 4550 -1510
rect 4430 -1580 4550 -1540
rect 4430 -1610 4475 -1580
rect 4505 -1610 4550 -1580
rect 4430 -1645 4550 -1610
rect 4430 -1675 4475 -1645
rect 4505 -1675 4550 -1645
rect 4430 -1705 4550 -1675
rect 4430 -1735 4475 -1705
rect 4505 -1735 4550 -1705
rect 4430 -1770 4550 -1735
rect 4430 -1800 4475 -1770
rect 4505 -1800 4550 -1770
rect 4430 -1840 4550 -1800
rect 4430 -1870 4475 -1840
rect 4505 -1870 4550 -1840
rect 4430 -1910 4550 -1870
rect 4430 -1940 4475 -1910
rect 4505 -1940 4550 -1910
rect 4430 -1980 4550 -1940
rect 4430 -2010 4475 -1980
rect 4505 -2010 4550 -1980
rect 4430 -2045 4550 -2010
rect 4430 -2075 4475 -2045
rect 4505 -2075 4550 -2045
rect 4430 -2105 4550 -2075
rect 4430 -2135 4475 -2105
rect 4505 -2135 4550 -2105
rect 4430 -2170 4550 -2135
rect 4430 -2200 4475 -2170
rect 4505 -2200 4550 -2170
rect 4430 -2240 4550 -2200
rect 4430 -2270 4475 -2240
rect 4505 -2270 4550 -2240
rect 4430 -2310 4550 -2270
rect 4430 -2340 4475 -2310
rect 4505 -2340 4550 -2310
rect 4430 -2380 4550 -2340
rect 4430 -2410 4475 -2380
rect 4505 -2410 4550 -2380
rect 4430 -2445 4550 -2410
rect 4430 -2475 4475 -2445
rect 4505 -2475 4550 -2445
rect 4430 -2505 4550 -2475
rect 4430 -2535 4475 -2505
rect 4505 -2535 4550 -2505
rect 4430 -2570 4550 -2535
rect 4430 -2600 4475 -2570
rect 4505 -2600 4550 -2570
rect 4430 -2640 4550 -2600
rect 4430 -2670 4475 -2640
rect 4505 -2670 4550 -2640
rect 4430 -2710 4550 -2670
rect 4430 -2740 4475 -2710
rect 4505 -2740 4550 -2710
rect 4430 -2780 4550 -2740
rect 4430 -2810 4475 -2780
rect 4505 -2810 4550 -2780
rect 4430 -2845 4550 -2810
rect 4430 -2875 4475 -2845
rect 4505 -2875 4550 -2845
rect 4430 -2905 4550 -2875
rect 4430 -2935 4475 -2905
rect 4505 -2935 4550 -2905
rect 4430 -2970 4550 -2935
rect 4430 -3000 4475 -2970
rect 4505 -3000 4550 -2970
rect 4430 -3040 4550 -3000
rect 4430 -3070 4475 -3040
rect 4505 -3070 4550 -3040
rect 4430 -3110 4550 -3070
rect 4430 -3140 4475 -3110
rect 4505 -3140 4550 -3110
rect 4430 -3180 4550 -3140
rect 4430 -3210 4475 -3180
rect 4505 -3210 4550 -3180
rect 4430 -3245 4550 -3210
rect 4430 -3275 4475 -3245
rect 4505 -3275 4550 -3245
rect 4430 -3305 4550 -3275
rect 4430 -3335 4475 -3305
rect 4505 -3335 4550 -3305
rect 4430 -3370 4550 -3335
rect 4430 -3400 4475 -3370
rect 4505 -3400 4550 -3370
rect 4430 -3440 4550 -3400
rect 4430 -3470 4475 -3440
rect 4505 -3470 4550 -3440
rect 4430 -3510 4550 -3470
rect 4430 -3540 4475 -3510
rect 4505 -3540 4550 -3510
rect 4430 -3580 4550 -3540
rect 4430 -3610 4475 -3580
rect 4505 -3610 4550 -3580
rect 4430 -3645 4550 -3610
rect 4430 -3675 4475 -3645
rect 4505 -3675 4550 -3645
rect 4430 -3705 4550 -3675
rect 4430 -3735 4475 -3705
rect 4505 -3735 4550 -3705
rect 4430 -3770 4550 -3735
rect 4430 -3800 4475 -3770
rect 4505 -3800 4550 -3770
rect 4430 -3840 4550 -3800
rect 4430 -3870 4475 -3840
rect 4505 -3870 4550 -3840
rect 4430 -3910 4550 -3870
rect 4430 -3940 4475 -3910
rect 4505 -3940 4550 -3910
rect 4430 -3980 4550 -3940
rect 4430 -4010 4475 -3980
rect 4505 -4010 4550 -3980
rect 4430 -4045 4550 -4010
rect 4430 -4075 4475 -4045
rect 4505 -4075 4550 -4045
rect 4430 -4105 4550 -4075
rect 4430 -4135 4475 -4105
rect 4505 -4135 4550 -4105
rect 4430 -4170 4550 -4135
rect 4430 -4200 4475 -4170
rect 4505 -4200 4550 -4170
rect 4430 -4240 4550 -4200
rect 4430 -4270 4475 -4240
rect 4505 -4270 4550 -4240
rect 4430 -4310 4550 -4270
rect 4430 -4340 4475 -4310
rect 4505 -4340 4550 -4310
rect 4430 -4380 4550 -4340
rect 4430 -4410 4475 -4380
rect 4505 -4410 4550 -4380
rect 4430 -4445 4550 -4410
rect 4430 -4475 4475 -4445
rect 4505 -4475 4550 -4445
rect 4430 -4490 4550 -4475
rect 4780 -1305 4900 -1240
rect 4780 -1335 4825 -1305
rect 4855 -1335 4900 -1305
rect 4780 -1370 4900 -1335
rect 4780 -1400 4825 -1370
rect 4855 -1400 4900 -1370
rect 4780 -1440 4900 -1400
rect 4780 -1470 4825 -1440
rect 4855 -1470 4900 -1440
rect 4780 -1510 4900 -1470
rect 4780 -1540 4825 -1510
rect 4855 -1540 4900 -1510
rect 4780 -1580 4900 -1540
rect 4780 -1610 4825 -1580
rect 4855 -1610 4900 -1580
rect 4780 -1645 4900 -1610
rect 4780 -1675 4825 -1645
rect 4855 -1675 4900 -1645
rect 4780 -1705 4900 -1675
rect 4780 -1735 4825 -1705
rect 4855 -1735 4900 -1705
rect 4780 -1770 4900 -1735
rect 4780 -1800 4825 -1770
rect 4855 -1800 4900 -1770
rect 4780 -1840 4900 -1800
rect 4780 -1870 4825 -1840
rect 4855 -1870 4900 -1840
rect 4780 -1910 4900 -1870
rect 4780 -1940 4825 -1910
rect 4855 -1940 4900 -1910
rect 4780 -1980 4900 -1940
rect 4780 -2010 4825 -1980
rect 4855 -2010 4900 -1980
rect 4780 -2045 4900 -2010
rect 4780 -2075 4825 -2045
rect 4855 -2075 4900 -2045
rect 4780 -2105 4900 -2075
rect 4780 -2135 4825 -2105
rect 4855 -2135 4900 -2105
rect 4780 -2170 4900 -2135
rect 4780 -2200 4825 -2170
rect 4855 -2200 4900 -2170
rect 4780 -2240 4900 -2200
rect 4780 -2270 4825 -2240
rect 4855 -2270 4900 -2240
rect 4780 -2310 4900 -2270
rect 4780 -2340 4825 -2310
rect 4855 -2340 4900 -2310
rect 4780 -2380 4900 -2340
rect 4780 -2410 4825 -2380
rect 4855 -2410 4900 -2380
rect 4780 -2445 4900 -2410
rect 4780 -2475 4825 -2445
rect 4855 -2475 4900 -2445
rect 4780 -2505 4900 -2475
rect 4780 -2535 4825 -2505
rect 4855 -2535 4900 -2505
rect 4780 -2570 4900 -2535
rect 4780 -2600 4825 -2570
rect 4855 -2600 4900 -2570
rect 4780 -2640 4900 -2600
rect 4780 -2670 4825 -2640
rect 4855 -2670 4900 -2640
rect 4780 -2710 4900 -2670
rect 4780 -2740 4825 -2710
rect 4855 -2740 4900 -2710
rect 4780 -2780 4900 -2740
rect 4780 -2810 4825 -2780
rect 4855 -2810 4900 -2780
rect 4780 -2845 4900 -2810
rect 4780 -2875 4825 -2845
rect 4855 -2875 4900 -2845
rect 4780 -2905 4900 -2875
rect 4780 -2935 4825 -2905
rect 4855 -2935 4900 -2905
rect 4780 -2970 4900 -2935
rect 4780 -3000 4825 -2970
rect 4855 -3000 4900 -2970
rect 4780 -3040 4900 -3000
rect 4780 -3070 4825 -3040
rect 4855 -3070 4900 -3040
rect 4780 -3110 4900 -3070
rect 4780 -3140 4825 -3110
rect 4855 -3140 4900 -3110
rect 4780 -3180 4900 -3140
rect 4780 -3210 4825 -3180
rect 4855 -3210 4900 -3180
rect 4780 -3245 4900 -3210
rect 4780 -3275 4825 -3245
rect 4855 -3275 4900 -3245
rect 4780 -3305 4900 -3275
rect 4780 -3335 4825 -3305
rect 4855 -3335 4900 -3305
rect 4780 -3370 4900 -3335
rect 4780 -3400 4825 -3370
rect 4855 -3400 4900 -3370
rect 4780 -3440 4900 -3400
rect 4780 -3470 4825 -3440
rect 4855 -3470 4900 -3440
rect 4780 -3510 4900 -3470
rect 4780 -3540 4825 -3510
rect 4855 -3540 4900 -3510
rect 4780 -3580 4900 -3540
rect 4780 -3610 4825 -3580
rect 4855 -3610 4900 -3580
rect 4780 -3645 4900 -3610
rect 4780 -3675 4825 -3645
rect 4855 -3675 4900 -3645
rect 4780 -3705 4900 -3675
rect 4780 -3735 4825 -3705
rect 4855 -3735 4900 -3705
rect 4780 -3770 4900 -3735
rect 4780 -3800 4825 -3770
rect 4855 -3800 4900 -3770
rect 4780 -3840 4900 -3800
rect 4780 -3870 4825 -3840
rect 4855 -3870 4900 -3840
rect 4780 -3910 4900 -3870
rect 4780 -3940 4825 -3910
rect 4855 -3940 4900 -3910
rect 4780 -3980 4900 -3940
rect 4780 -4010 4825 -3980
rect 4855 -4010 4900 -3980
rect 4780 -4045 4900 -4010
rect 4780 -4075 4825 -4045
rect 4855 -4075 4900 -4045
rect 4780 -4105 4900 -4075
rect 4780 -4135 4825 -4105
rect 4855 -4135 4900 -4105
rect 4780 -4170 4900 -4135
rect 4780 -4200 4825 -4170
rect 4855 -4200 4900 -4170
rect 4780 -4240 4900 -4200
rect 4780 -4270 4825 -4240
rect 4855 -4270 4900 -4240
rect 4780 -4310 4900 -4270
rect 4780 -4340 4825 -4310
rect 4855 -4340 4900 -4310
rect 4780 -4380 4900 -4340
rect 4780 -4410 4825 -4380
rect 4855 -4410 4900 -4380
rect 4780 -4445 4900 -4410
rect 4780 -4475 4825 -4445
rect 4855 -4475 4900 -4445
rect 4780 -4490 4900 -4475
rect 5130 -1305 5250 -1240
rect 5130 -1335 5175 -1305
rect 5205 -1335 5250 -1305
rect 5130 -1370 5250 -1335
rect 5130 -1400 5175 -1370
rect 5205 -1400 5250 -1370
rect 5130 -1440 5250 -1400
rect 5130 -1470 5175 -1440
rect 5205 -1470 5250 -1440
rect 5130 -1510 5250 -1470
rect 5130 -1540 5175 -1510
rect 5205 -1540 5250 -1510
rect 5130 -1580 5250 -1540
rect 5130 -1610 5175 -1580
rect 5205 -1610 5250 -1580
rect 5130 -1645 5250 -1610
rect 5130 -1675 5175 -1645
rect 5205 -1675 5250 -1645
rect 5130 -1705 5250 -1675
rect 5130 -1735 5175 -1705
rect 5205 -1735 5250 -1705
rect 5130 -1770 5250 -1735
rect 5130 -1800 5175 -1770
rect 5205 -1800 5250 -1770
rect 5130 -1840 5250 -1800
rect 5130 -1870 5175 -1840
rect 5205 -1870 5250 -1840
rect 5130 -1910 5250 -1870
rect 5130 -1940 5175 -1910
rect 5205 -1940 5250 -1910
rect 5130 -1980 5250 -1940
rect 5130 -2010 5175 -1980
rect 5205 -2010 5250 -1980
rect 5130 -2045 5250 -2010
rect 5130 -2075 5175 -2045
rect 5205 -2075 5250 -2045
rect 5130 -2105 5250 -2075
rect 5130 -2135 5175 -2105
rect 5205 -2135 5250 -2105
rect 5130 -2170 5250 -2135
rect 5130 -2200 5175 -2170
rect 5205 -2200 5250 -2170
rect 5130 -2240 5250 -2200
rect 5130 -2270 5175 -2240
rect 5205 -2270 5250 -2240
rect 5130 -2310 5250 -2270
rect 5130 -2340 5175 -2310
rect 5205 -2340 5250 -2310
rect 5130 -2380 5250 -2340
rect 5130 -2410 5175 -2380
rect 5205 -2410 5250 -2380
rect 5130 -2445 5250 -2410
rect 5130 -2475 5175 -2445
rect 5205 -2475 5250 -2445
rect 5130 -2505 5250 -2475
rect 5130 -2535 5175 -2505
rect 5205 -2535 5250 -2505
rect 5130 -2570 5250 -2535
rect 5130 -2600 5175 -2570
rect 5205 -2600 5250 -2570
rect 5130 -2640 5250 -2600
rect 5130 -2670 5175 -2640
rect 5205 -2670 5250 -2640
rect 5130 -2710 5250 -2670
rect 5130 -2740 5175 -2710
rect 5205 -2740 5250 -2710
rect 5130 -2780 5250 -2740
rect 5130 -2810 5175 -2780
rect 5205 -2810 5250 -2780
rect 5130 -2845 5250 -2810
rect 5130 -2875 5175 -2845
rect 5205 -2875 5250 -2845
rect 5130 -2905 5250 -2875
rect 5130 -2935 5175 -2905
rect 5205 -2935 5250 -2905
rect 5130 -2970 5250 -2935
rect 5130 -3000 5175 -2970
rect 5205 -3000 5250 -2970
rect 5130 -3040 5250 -3000
rect 5130 -3070 5175 -3040
rect 5205 -3070 5250 -3040
rect 5130 -3110 5250 -3070
rect 5130 -3140 5175 -3110
rect 5205 -3140 5250 -3110
rect 5130 -3180 5250 -3140
rect 5130 -3210 5175 -3180
rect 5205 -3210 5250 -3180
rect 5130 -3245 5250 -3210
rect 5130 -3275 5175 -3245
rect 5205 -3275 5250 -3245
rect 5130 -3305 5250 -3275
rect 5130 -3335 5175 -3305
rect 5205 -3335 5250 -3305
rect 5130 -3370 5250 -3335
rect 5130 -3400 5175 -3370
rect 5205 -3400 5250 -3370
rect 5130 -3440 5250 -3400
rect 5130 -3470 5175 -3440
rect 5205 -3470 5250 -3440
rect 5130 -3510 5250 -3470
rect 5130 -3540 5175 -3510
rect 5205 -3540 5250 -3510
rect 5130 -3580 5250 -3540
rect 5130 -3610 5175 -3580
rect 5205 -3610 5250 -3580
rect 5130 -3645 5250 -3610
rect 5130 -3675 5175 -3645
rect 5205 -3675 5250 -3645
rect 5130 -3705 5250 -3675
rect 5130 -3735 5175 -3705
rect 5205 -3735 5250 -3705
rect 5130 -3770 5250 -3735
rect 5130 -3800 5175 -3770
rect 5205 -3800 5250 -3770
rect 5130 -3840 5250 -3800
rect 5130 -3870 5175 -3840
rect 5205 -3870 5250 -3840
rect 5130 -3910 5250 -3870
rect 5130 -3940 5175 -3910
rect 5205 -3940 5250 -3910
rect 5130 -3980 5250 -3940
rect 5130 -4010 5175 -3980
rect 5205 -4010 5250 -3980
rect 5130 -4045 5250 -4010
rect 5130 -4075 5175 -4045
rect 5205 -4075 5250 -4045
rect 5130 -4105 5250 -4075
rect 5130 -4135 5175 -4105
rect 5205 -4135 5250 -4105
rect 5130 -4170 5250 -4135
rect 5130 -4200 5175 -4170
rect 5205 -4200 5250 -4170
rect 5130 -4240 5250 -4200
rect 5130 -4270 5175 -4240
rect 5205 -4270 5250 -4240
rect 5130 -4310 5250 -4270
rect 5130 -4340 5175 -4310
rect 5205 -4340 5250 -4310
rect 5130 -4380 5250 -4340
rect 5130 -4410 5175 -4380
rect 5205 -4410 5250 -4380
rect 5130 -4445 5250 -4410
rect 5130 -4475 5175 -4445
rect 5205 -4475 5250 -4445
rect 5130 -4490 5250 -4475
rect 5480 -1305 5600 -1240
rect 5480 -1335 5525 -1305
rect 5555 -1335 5600 -1305
rect 5480 -1370 5600 -1335
rect 5480 -1400 5525 -1370
rect 5555 -1400 5600 -1370
rect 5480 -1440 5600 -1400
rect 5480 -1470 5525 -1440
rect 5555 -1470 5600 -1440
rect 5480 -1510 5600 -1470
rect 5480 -1540 5525 -1510
rect 5555 -1540 5600 -1510
rect 5480 -1580 5600 -1540
rect 5480 -1610 5525 -1580
rect 5555 -1610 5600 -1580
rect 5480 -1645 5600 -1610
rect 5480 -1675 5525 -1645
rect 5555 -1675 5600 -1645
rect 5480 -1705 5600 -1675
rect 5480 -1735 5525 -1705
rect 5555 -1735 5600 -1705
rect 5480 -1770 5600 -1735
rect 5480 -1800 5525 -1770
rect 5555 -1800 5600 -1770
rect 5480 -1840 5600 -1800
rect 5480 -1870 5525 -1840
rect 5555 -1870 5600 -1840
rect 5480 -1910 5600 -1870
rect 5480 -1940 5525 -1910
rect 5555 -1940 5600 -1910
rect 5480 -1980 5600 -1940
rect 5480 -2010 5525 -1980
rect 5555 -2010 5600 -1980
rect 5480 -2045 5600 -2010
rect 5480 -2075 5525 -2045
rect 5555 -2075 5600 -2045
rect 5480 -2105 5600 -2075
rect 5480 -2135 5525 -2105
rect 5555 -2135 5600 -2105
rect 5480 -2170 5600 -2135
rect 5480 -2200 5525 -2170
rect 5555 -2200 5600 -2170
rect 5480 -2240 5600 -2200
rect 5480 -2270 5525 -2240
rect 5555 -2270 5600 -2240
rect 5480 -2310 5600 -2270
rect 5480 -2340 5525 -2310
rect 5555 -2340 5600 -2310
rect 5480 -2380 5600 -2340
rect 5480 -2410 5525 -2380
rect 5555 -2410 5600 -2380
rect 5480 -2445 5600 -2410
rect 5480 -2475 5525 -2445
rect 5555 -2475 5600 -2445
rect 5480 -2505 5600 -2475
rect 5480 -2535 5525 -2505
rect 5555 -2535 5600 -2505
rect 5480 -2570 5600 -2535
rect 5480 -2600 5525 -2570
rect 5555 -2600 5600 -2570
rect 5480 -2640 5600 -2600
rect 5480 -2670 5525 -2640
rect 5555 -2670 5600 -2640
rect 5480 -2710 5600 -2670
rect 5480 -2740 5525 -2710
rect 5555 -2740 5600 -2710
rect 5480 -2780 5600 -2740
rect 5480 -2810 5525 -2780
rect 5555 -2810 5600 -2780
rect 5480 -2845 5600 -2810
rect 5480 -2875 5525 -2845
rect 5555 -2875 5600 -2845
rect 5480 -2905 5600 -2875
rect 5480 -2935 5525 -2905
rect 5555 -2935 5600 -2905
rect 5480 -2970 5600 -2935
rect 5480 -3000 5525 -2970
rect 5555 -3000 5600 -2970
rect 5480 -3040 5600 -3000
rect 5480 -3070 5525 -3040
rect 5555 -3070 5600 -3040
rect 5480 -3110 5600 -3070
rect 5480 -3140 5525 -3110
rect 5555 -3140 5600 -3110
rect 5480 -3180 5600 -3140
rect 5480 -3210 5525 -3180
rect 5555 -3210 5600 -3180
rect 5480 -3245 5600 -3210
rect 5480 -3275 5525 -3245
rect 5555 -3275 5600 -3245
rect 5480 -3305 5600 -3275
rect 5480 -3335 5525 -3305
rect 5555 -3335 5600 -3305
rect 5480 -3370 5600 -3335
rect 5480 -3400 5525 -3370
rect 5555 -3400 5600 -3370
rect 5480 -3440 5600 -3400
rect 5480 -3470 5525 -3440
rect 5555 -3470 5600 -3440
rect 5480 -3510 5600 -3470
rect 5480 -3540 5525 -3510
rect 5555 -3540 5600 -3510
rect 5480 -3580 5600 -3540
rect 5480 -3610 5525 -3580
rect 5555 -3610 5600 -3580
rect 5480 -3645 5600 -3610
rect 5480 -3675 5525 -3645
rect 5555 -3675 5600 -3645
rect 5480 -3705 5600 -3675
rect 5480 -3735 5525 -3705
rect 5555 -3735 5600 -3705
rect 5480 -3770 5600 -3735
rect 5480 -3800 5525 -3770
rect 5555 -3800 5600 -3770
rect 5480 -3840 5600 -3800
rect 5480 -3870 5525 -3840
rect 5555 -3870 5600 -3840
rect 5480 -3910 5600 -3870
rect 5480 -3940 5525 -3910
rect 5555 -3940 5600 -3910
rect 5480 -3980 5600 -3940
rect 5480 -4010 5525 -3980
rect 5555 -4010 5600 -3980
rect 5480 -4045 5600 -4010
rect 5480 -4075 5525 -4045
rect 5555 -4075 5600 -4045
rect 5480 -4105 5600 -4075
rect 5480 -4135 5525 -4105
rect 5555 -4135 5600 -4105
rect 5480 -4170 5600 -4135
rect 5480 -4200 5525 -4170
rect 5555 -4200 5600 -4170
rect 5480 -4240 5600 -4200
rect 5480 -4270 5525 -4240
rect 5555 -4270 5600 -4240
rect 5480 -4310 5600 -4270
rect 5480 -4340 5525 -4310
rect 5555 -4340 5600 -4310
rect 5480 -4380 5600 -4340
rect 5480 -4410 5525 -4380
rect 5555 -4410 5600 -4380
rect 5480 -4445 5600 -4410
rect 5480 -4475 5525 -4445
rect 5555 -4475 5600 -4445
rect 5480 -4490 5600 -4475
rect 5830 -1305 5950 -1240
rect 5830 -1335 5875 -1305
rect 5905 -1335 5950 -1305
rect 5830 -1370 5950 -1335
rect 5830 -1400 5875 -1370
rect 5905 -1400 5950 -1370
rect 5830 -1440 5950 -1400
rect 5830 -1470 5875 -1440
rect 5905 -1470 5950 -1440
rect 5830 -1510 5950 -1470
rect 5830 -1540 5875 -1510
rect 5905 -1540 5950 -1510
rect 5830 -1580 5950 -1540
rect 5830 -1610 5875 -1580
rect 5905 -1610 5950 -1580
rect 5830 -1645 5950 -1610
rect 5830 -1675 5875 -1645
rect 5905 -1675 5950 -1645
rect 5830 -1705 5950 -1675
rect 5830 -1735 5875 -1705
rect 5905 -1735 5950 -1705
rect 5830 -1770 5950 -1735
rect 5830 -1800 5875 -1770
rect 5905 -1800 5950 -1770
rect 5830 -1840 5950 -1800
rect 5830 -1870 5875 -1840
rect 5905 -1870 5950 -1840
rect 5830 -1910 5950 -1870
rect 5830 -1940 5875 -1910
rect 5905 -1940 5950 -1910
rect 5830 -1980 5950 -1940
rect 5830 -2010 5875 -1980
rect 5905 -2010 5950 -1980
rect 5830 -2045 5950 -2010
rect 5830 -2075 5875 -2045
rect 5905 -2075 5950 -2045
rect 5830 -2105 5950 -2075
rect 5830 -2135 5875 -2105
rect 5905 -2135 5950 -2105
rect 5830 -2170 5950 -2135
rect 5830 -2200 5875 -2170
rect 5905 -2200 5950 -2170
rect 5830 -2240 5950 -2200
rect 5830 -2270 5875 -2240
rect 5905 -2270 5950 -2240
rect 5830 -2310 5950 -2270
rect 5830 -2340 5875 -2310
rect 5905 -2340 5950 -2310
rect 5830 -2380 5950 -2340
rect 5830 -2410 5875 -2380
rect 5905 -2410 5950 -2380
rect 5830 -2445 5950 -2410
rect 5830 -2475 5875 -2445
rect 5905 -2475 5950 -2445
rect 5830 -2505 5950 -2475
rect 5830 -2535 5875 -2505
rect 5905 -2535 5950 -2505
rect 5830 -2570 5950 -2535
rect 5830 -2600 5875 -2570
rect 5905 -2600 5950 -2570
rect 5830 -2640 5950 -2600
rect 5830 -2670 5875 -2640
rect 5905 -2670 5950 -2640
rect 5830 -2710 5950 -2670
rect 5830 -2740 5875 -2710
rect 5905 -2740 5950 -2710
rect 5830 -2780 5950 -2740
rect 5830 -2810 5875 -2780
rect 5905 -2810 5950 -2780
rect 5830 -2845 5950 -2810
rect 5830 -2875 5875 -2845
rect 5905 -2875 5950 -2845
rect 5830 -2905 5950 -2875
rect 5830 -2935 5875 -2905
rect 5905 -2935 5950 -2905
rect 5830 -2970 5950 -2935
rect 5830 -3000 5875 -2970
rect 5905 -3000 5950 -2970
rect 5830 -3040 5950 -3000
rect 5830 -3070 5875 -3040
rect 5905 -3070 5950 -3040
rect 5830 -3110 5950 -3070
rect 5830 -3140 5875 -3110
rect 5905 -3140 5950 -3110
rect 5830 -3180 5950 -3140
rect 5830 -3210 5875 -3180
rect 5905 -3210 5950 -3180
rect 5830 -3245 5950 -3210
rect 5830 -3275 5875 -3245
rect 5905 -3275 5950 -3245
rect 5830 -3305 5950 -3275
rect 5830 -3335 5875 -3305
rect 5905 -3335 5950 -3305
rect 5830 -3370 5950 -3335
rect 5830 -3400 5875 -3370
rect 5905 -3400 5950 -3370
rect 5830 -3440 5950 -3400
rect 5830 -3470 5875 -3440
rect 5905 -3470 5950 -3440
rect 5830 -3510 5950 -3470
rect 5830 -3540 5875 -3510
rect 5905 -3540 5950 -3510
rect 5830 -3580 5950 -3540
rect 5830 -3610 5875 -3580
rect 5905 -3610 5950 -3580
rect 5830 -3645 5950 -3610
rect 5830 -3675 5875 -3645
rect 5905 -3675 5950 -3645
rect 5830 -3705 5950 -3675
rect 5830 -3735 5875 -3705
rect 5905 -3735 5950 -3705
rect 5830 -3770 5950 -3735
rect 5830 -3800 5875 -3770
rect 5905 -3800 5950 -3770
rect 5830 -3840 5950 -3800
rect 5830 -3870 5875 -3840
rect 5905 -3870 5950 -3840
rect 5830 -3910 5950 -3870
rect 5830 -3940 5875 -3910
rect 5905 -3940 5950 -3910
rect 5830 -3980 5950 -3940
rect 5830 -4010 5875 -3980
rect 5905 -4010 5950 -3980
rect 5830 -4045 5950 -4010
rect 5830 -4075 5875 -4045
rect 5905 -4075 5950 -4045
rect 5830 -4105 5950 -4075
rect 5830 -4135 5875 -4105
rect 5905 -4135 5950 -4105
rect 5830 -4170 5950 -4135
rect 5830 -4200 5875 -4170
rect 5905 -4200 5950 -4170
rect 5830 -4240 5950 -4200
rect 5830 -4270 5875 -4240
rect 5905 -4270 5950 -4240
rect 5830 -4310 5950 -4270
rect 5830 -4340 5875 -4310
rect 5905 -4340 5950 -4310
rect 5830 -4380 5950 -4340
rect 5830 -4410 5875 -4380
rect 5905 -4410 5950 -4380
rect 5830 -4445 5950 -4410
rect 5830 -4475 5875 -4445
rect 5905 -4475 5950 -4445
rect 5830 -4490 5950 -4475
rect 6180 -1305 6300 -1240
rect 6180 -1335 6225 -1305
rect 6255 -1335 6300 -1305
rect 6180 -1370 6300 -1335
rect 6180 -1400 6225 -1370
rect 6255 -1400 6300 -1370
rect 6180 -1440 6300 -1400
rect 6180 -1470 6225 -1440
rect 6255 -1470 6300 -1440
rect 6180 -1510 6300 -1470
rect 6180 -1540 6225 -1510
rect 6255 -1540 6300 -1510
rect 6180 -1580 6300 -1540
rect 6180 -1610 6225 -1580
rect 6255 -1610 6300 -1580
rect 6180 -1645 6300 -1610
rect 6180 -1675 6225 -1645
rect 6255 -1675 6300 -1645
rect 6180 -1705 6300 -1675
rect 6180 -1735 6225 -1705
rect 6255 -1735 6300 -1705
rect 6180 -1770 6300 -1735
rect 6180 -1800 6225 -1770
rect 6255 -1800 6300 -1770
rect 6180 -1840 6300 -1800
rect 6180 -1870 6225 -1840
rect 6255 -1870 6300 -1840
rect 6180 -1910 6300 -1870
rect 6180 -1940 6225 -1910
rect 6255 -1940 6300 -1910
rect 6180 -1980 6300 -1940
rect 6180 -2010 6225 -1980
rect 6255 -2010 6300 -1980
rect 6180 -2045 6300 -2010
rect 6180 -2075 6225 -2045
rect 6255 -2075 6300 -2045
rect 6180 -2105 6300 -2075
rect 6180 -2135 6225 -2105
rect 6255 -2135 6300 -2105
rect 6180 -2170 6300 -2135
rect 6180 -2200 6225 -2170
rect 6255 -2200 6300 -2170
rect 6180 -2240 6300 -2200
rect 6180 -2270 6225 -2240
rect 6255 -2270 6300 -2240
rect 6180 -2310 6300 -2270
rect 6180 -2340 6225 -2310
rect 6255 -2340 6300 -2310
rect 6180 -2380 6300 -2340
rect 6180 -2410 6225 -2380
rect 6255 -2410 6300 -2380
rect 6180 -2445 6300 -2410
rect 6180 -2475 6225 -2445
rect 6255 -2475 6300 -2445
rect 6180 -2505 6300 -2475
rect 6180 -2535 6225 -2505
rect 6255 -2535 6300 -2505
rect 6180 -2570 6300 -2535
rect 6180 -2600 6225 -2570
rect 6255 -2600 6300 -2570
rect 6180 -2640 6300 -2600
rect 6180 -2670 6225 -2640
rect 6255 -2670 6300 -2640
rect 6180 -2710 6300 -2670
rect 6180 -2740 6225 -2710
rect 6255 -2740 6300 -2710
rect 6180 -2780 6300 -2740
rect 6180 -2810 6225 -2780
rect 6255 -2810 6300 -2780
rect 6180 -2845 6300 -2810
rect 6180 -2875 6225 -2845
rect 6255 -2875 6300 -2845
rect 6180 -2905 6300 -2875
rect 6180 -2935 6225 -2905
rect 6255 -2935 6300 -2905
rect 6180 -2970 6300 -2935
rect 6180 -3000 6225 -2970
rect 6255 -3000 6300 -2970
rect 6180 -3040 6300 -3000
rect 6180 -3070 6225 -3040
rect 6255 -3070 6300 -3040
rect 6180 -3110 6300 -3070
rect 6180 -3140 6225 -3110
rect 6255 -3140 6300 -3110
rect 6180 -3180 6300 -3140
rect 6180 -3210 6225 -3180
rect 6255 -3210 6300 -3180
rect 6180 -3245 6300 -3210
rect 6180 -3275 6225 -3245
rect 6255 -3275 6300 -3245
rect 6180 -3305 6300 -3275
rect 6180 -3335 6225 -3305
rect 6255 -3335 6300 -3305
rect 6180 -3370 6300 -3335
rect 6180 -3400 6225 -3370
rect 6255 -3400 6300 -3370
rect 6180 -3440 6300 -3400
rect 6180 -3470 6225 -3440
rect 6255 -3470 6300 -3440
rect 6180 -3510 6300 -3470
rect 6180 -3540 6225 -3510
rect 6255 -3540 6300 -3510
rect 6180 -3580 6300 -3540
rect 6180 -3610 6225 -3580
rect 6255 -3610 6300 -3580
rect 6180 -3645 6300 -3610
rect 6180 -3675 6225 -3645
rect 6255 -3675 6300 -3645
rect 6180 -3705 6300 -3675
rect 6180 -3735 6225 -3705
rect 6255 -3735 6300 -3705
rect 6180 -3770 6300 -3735
rect 6180 -3800 6225 -3770
rect 6255 -3800 6300 -3770
rect 6180 -3840 6300 -3800
rect 6180 -3870 6225 -3840
rect 6255 -3870 6300 -3840
rect 6180 -3910 6300 -3870
rect 6180 -3940 6225 -3910
rect 6255 -3940 6300 -3910
rect 6180 -3980 6300 -3940
rect 6180 -4010 6225 -3980
rect 6255 -4010 6300 -3980
rect 6180 -4045 6300 -4010
rect 6180 -4075 6225 -4045
rect 6255 -4075 6300 -4045
rect 6180 -4105 6300 -4075
rect 6180 -4135 6225 -4105
rect 6255 -4135 6300 -4105
rect 6180 -4170 6300 -4135
rect 6180 -4200 6225 -4170
rect 6255 -4200 6300 -4170
rect 6180 -4240 6300 -4200
rect 6180 -4270 6225 -4240
rect 6255 -4270 6300 -4240
rect 6180 -4310 6300 -4270
rect 6180 -4340 6225 -4310
rect 6255 -4340 6300 -4310
rect 6180 -4380 6300 -4340
rect 6180 -4410 6225 -4380
rect 6255 -4410 6300 -4380
rect 6180 -4445 6300 -4410
rect 6180 -4475 6225 -4445
rect 6255 -4475 6300 -4445
rect 6180 -4490 6300 -4475
rect 6530 -1305 6650 -1240
rect 6530 -1335 6575 -1305
rect 6605 -1335 6650 -1305
rect 6530 -1370 6650 -1335
rect 6530 -1400 6575 -1370
rect 6605 -1400 6650 -1370
rect 6530 -1440 6650 -1400
rect 6530 -1470 6575 -1440
rect 6605 -1470 6650 -1440
rect 6530 -1510 6650 -1470
rect 6530 -1540 6575 -1510
rect 6605 -1540 6650 -1510
rect 6530 -1580 6650 -1540
rect 6530 -1610 6575 -1580
rect 6605 -1610 6650 -1580
rect 6530 -1645 6650 -1610
rect 6530 -1675 6575 -1645
rect 6605 -1675 6650 -1645
rect 6530 -1705 6650 -1675
rect 6530 -1735 6575 -1705
rect 6605 -1735 6650 -1705
rect 6530 -1770 6650 -1735
rect 6530 -1800 6575 -1770
rect 6605 -1800 6650 -1770
rect 6530 -1840 6650 -1800
rect 6530 -1870 6575 -1840
rect 6605 -1870 6650 -1840
rect 6530 -1910 6650 -1870
rect 6530 -1940 6575 -1910
rect 6605 -1940 6650 -1910
rect 6530 -1980 6650 -1940
rect 6530 -2010 6575 -1980
rect 6605 -2010 6650 -1980
rect 6530 -2045 6650 -2010
rect 6530 -2075 6575 -2045
rect 6605 -2075 6650 -2045
rect 6530 -2105 6650 -2075
rect 6530 -2135 6575 -2105
rect 6605 -2135 6650 -2105
rect 6530 -2170 6650 -2135
rect 6530 -2200 6575 -2170
rect 6605 -2200 6650 -2170
rect 6530 -2240 6650 -2200
rect 6530 -2270 6575 -2240
rect 6605 -2270 6650 -2240
rect 6530 -2310 6650 -2270
rect 6530 -2340 6575 -2310
rect 6605 -2340 6650 -2310
rect 6530 -2380 6650 -2340
rect 6530 -2410 6575 -2380
rect 6605 -2410 6650 -2380
rect 6530 -2445 6650 -2410
rect 6530 -2475 6575 -2445
rect 6605 -2475 6650 -2445
rect 6530 -2505 6650 -2475
rect 6530 -2535 6575 -2505
rect 6605 -2535 6650 -2505
rect 6530 -2570 6650 -2535
rect 6530 -2600 6575 -2570
rect 6605 -2600 6650 -2570
rect 6530 -2640 6650 -2600
rect 6530 -2670 6575 -2640
rect 6605 -2670 6650 -2640
rect 6530 -2710 6650 -2670
rect 6530 -2740 6575 -2710
rect 6605 -2740 6650 -2710
rect 6530 -2780 6650 -2740
rect 6530 -2810 6575 -2780
rect 6605 -2810 6650 -2780
rect 6530 -2845 6650 -2810
rect 6530 -2875 6575 -2845
rect 6605 -2875 6650 -2845
rect 6530 -2905 6650 -2875
rect 6530 -2935 6575 -2905
rect 6605 -2935 6650 -2905
rect 6530 -2970 6650 -2935
rect 6530 -3000 6575 -2970
rect 6605 -3000 6650 -2970
rect 6530 -3040 6650 -3000
rect 6530 -3070 6575 -3040
rect 6605 -3070 6650 -3040
rect 6530 -3110 6650 -3070
rect 6530 -3140 6575 -3110
rect 6605 -3140 6650 -3110
rect 6530 -3180 6650 -3140
rect 6530 -3210 6575 -3180
rect 6605 -3210 6650 -3180
rect 6530 -3245 6650 -3210
rect 6530 -3275 6575 -3245
rect 6605 -3275 6650 -3245
rect 6530 -3305 6650 -3275
rect 6530 -3335 6575 -3305
rect 6605 -3335 6650 -3305
rect 6530 -3370 6650 -3335
rect 6530 -3400 6575 -3370
rect 6605 -3400 6650 -3370
rect 6530 -3440 6650 -3400
rect 6530 -3470 6575 -3440
rect 6605 -3470 6650 -3440
rect 6530 -3510 6650 -3470
rect 6530 -3540 6575 -3510
rect 6605 -3540 6650 -3510
rect 6530 -3580 6650 -3540
rect 6530 -3610 6575 -3580
rect 6605 -3610 6650 -3580
rect 6530 -3645 6650 -3610
rect 6530 -3675 6575 -3645
rect 6605 -3675 6650 -3645
rect 6530 -3705 6650 -3675
rect 6530 -3735 6575 -3705
rect 6605 -3735 6650 -3705
rect 6530 -3770 6650 -3735
rect 6530 -3800 6575 -3770
rect 6605 -3800 6650 -3770
rect 6530 -3840 6650 -3800
rect 6530 -3870 6575 -3840
rect 6605 -3870 6650 -3840
rect 6530 -3910 6650 -3870
rect 6530 -3940 6575 -3910
rect 6605 -3940 6650 -3910
rect 6530 -3980 6650 -3940
rect 6530 -4010 6575 -3980
rect 6605 -4010 6650 -3980
rect 6530 -4045 6650 -4010
rect 6530 -4075 6575 -4045
rect 6605 -4075 6650 -4045
rect 6530 -4105 6650 -4075
rect 6530 -4135 6575 -4105
rect 6605 -4135 6650 -4105
rect 6530 -4170 6650 -4135
rect 6530 -4200 6575 -4170
rect 6605 -4200 6650 -4170
rect 6530 -4240 6650 -4200
rect 6530 -4270 6575 -4240
rect 6605 -4270 6650 -4240
rect 6530 -4310 6650 -4270
rect 6530 -4340 6575 -4310
rect 6605 -4340 6650 -4310
rect 6530 -4380 6650 -4340
rect 6530 -4410 6575 -4380
rect 6605 -4410 6650 -4380
rect 6530 -4445 6650 -4410
rect 6530 -4475 6575 -4445
rect 6605 -4475 6650 -4445
rect 6530 -4490 6650 -4475
rect 6880 -1305 7000 -1240
rect 6880 -1335 6925 -1305
rect 6955 -1335 7000 -1305
rect 6880 -1370 7000 -1335
rect 6880 -1400 6925 -1370
rect 6955 -1400 7000 -1370
rect 6880 -1440 7000 -1400
rect 6880 -1470 6925 -1440
rect 6955 -1470 7000 -1440
rect 6880 -1510 7000 -1470
rect 6880 -1540 6925 -1510
rect 6955 -1540 7000 -1510
rect 6880 -1580 7000 -1540
rect 6880 -1610 6925 -1580
rect 6955 -1610 7000 -1580
rect 6880 -1645 7000 -1610
rect 6880 -1675 6925 -1645
rect 6955 -1675 7000 -1645
rect 6880 -1705 7000 -1675
rect 6880 -1735 6925 -1705
rect 6955 -1735 7000 -1705
rect 6880 -1770 7000 -1735
rect 6880 -1800 6925 -1770
rect 6955 -1800 7000 -1770
rect 6880 -1840 7000 -1800
rect 6880 -1870 6925 -1840
rect 6955 -1870 7000 -1840
rect 6880 -1910 7000 -1870
rect 6880 -1940 6925 -1910
rect 6955 -1940 7000 -1910
rect 6880 -1980 7000 -1940
rect 6880 -2010 6925 -1980
rect 6955 -2010 7000 -1980
rect 6880 -2045 7000 -2010
rect 6880 -2075 6925 -2045
rect 6955 -2075 7000 -2045
rect 6880 -2105 7000 -2075
rect 6880 -2135 6925 -2105
rect 6955 -2135 7000 -2105
rect 6880 -2170 7000 -2135
rect 6880 -2200 6925 -2170
rect 6955 -2200 7000 -2170
rect 6880 -2240 7000 -2200
rect 6880 -2270 6925 -2240
rect 6955 -2270 7000 -2240
rect 6880 -2310 7000 -2270
rect 6880 -2340 6925 -2310
rect 6955 -2340 7000 -2310
rect 6880 -2380 7000 -2340
rect 6880 -2410 6925 -2380
rect 6955 -2410 7000 -2380
rect 6880 -2445 7000 -2410
rect 6880 -2475 6925 -2445
rect 6955 -2475 7000 -2445
rect 6880 -2505 7000 -2475
rect 6880 -2535 6925 -2505
rect 6955 -2535 7000 -2505
rect 6880 -2570 7000 -2535
rect 6880 -2600 6925 -2570
rect 6955 -2600 7000 -2570
rect 6880 -2640 7000 -2600
rect 6880 -2670 6925 -2640
rect 6955 -2670 7000 -2640
rect 6880 -2710 7000 -2670
rect 6880 -2740 6925 -2710
rect 6955 -2740 7000 -2710
rect 6880 -2780 7000 -2740
rect 6880 -2810 6925 -2780
rect 6955 -2810 7000 -2780
rect 6880 -2845 7000 -2810
rect 6880 -2875 6925 -2845
rect 6955 -2875 7000 -2845
rect 6880 -2905 7000 -2875
rect 6880 -2935 6925 -2905
rect 6955 -2935 7000 -2905
rect 6880 -2970 7000 -2935
rect 6880 -3000 6925 -2970
rect 6955 -3000 7000 -2970
rect 6880 -3040 7000 -3000
rect 6880 -3070 6925 -3040
rect 6955 -3070 7000 -3040
rect 6880 -3110 7000 -3070
rect 6880 -3140 6925 -3110
rect 6955 -3140 7000 -3110
rect 6880 -3180 7000 -3140
rect 6880 -3210 6925 -3180
rect 6955 -3210 7000 -3180
rect 6880 -3245 7000 -3210
rect 6880 -3275 6925 -3245
rect 6955 -3275 7000 -3245
rect 6880 -3305 7000 -3275
rect 6880 -3335 6925 -3305
rect 6955 -3335 7000 -3305
rect 6880 -3370 7000 -3335
rect 6880 -3400 6925 -3370
rect 6955 -3400 7000 -3370
rect 6880 -3440 7000 -3400
rect 6880 -3470 6925 -3440
rect 6955 -3470 7000 -3440
rect 6880 -3510 7000 -3470
rect 6880 -3540 6925 -3510
rect 6955 -3540 7000 -3510
rect 6880 -3580 7000 -3540
rect 6880 -3610 6925 -3580
rect 6955 -3610 7000 -3580
rect 6880 -3645 7000 -3610
rect 6880 -3675 6925 -3645
rect 6955 -3675 7000 -3645
rect 6880 -3705 7000 -3675
rect 6880 -3735 6925 -3705
rect 6955 -3735 7000 -3705
rect 6880 -3770 7000 -3735
rect 6880 -3800 6925 -3770
rect 6955 -3800 7000 -3770
rect 6880 -3840 7000 -3800
rect 6880 -3870 6925 -3840
rect 6955 -3870 7000 -3840
rect 6880 -3910 7000 -3870
rect 6880 -3940 6925 -3910
rect 6955 -3940 7000 -3910
rect 6880 -3980 7000 -3940
rect 6880 -4010 6925 -3980
rect 6955 -4010 7000 -3980
rect 6880 -4045 7000 -4010
rect 6880 -4075 6925 -4045
rect 6955 -4075 7000 -4045
rect 6880 -4105 7000 -4075
rect 6880 -4135 6925 -4105
rect 6955 -4135 7000 -4105
rect 6880 -4170 7000 -4135
rect 6880 -4200 6925 -4170
rect 6955 -4200 7000 -4170
rect 6880 -4240 7000 -4200
rect 6880 -4270 6925 -4240
rect 6955 -4270 7000 -4240
rect 6880 -4310 7000 -4270
rect 6880 -4340 6925 -4310
rect 6955 -4340 7000 -4310
rect 6880 -4380 7000 -4340
rect 6880 -4410 6925 -4380
rect 6955 -4410 7000 -4380
rect 6880 -4445 7000 -4410
rect 6880 -4475 6925 -4445
rect 6955 -4475 7000 -4445
rect 6880 -4490 7000 -4475
rect 7230 -1305 7350 -1240
rect 7230 -1335 7275 -1305
rect 7305 -1335 7350 -1305
rect 7230 -1370 7350 -1335
rect 7230 -1400 7275 -1370
rect 7305 -1400 7350 -1370
rect 7230 -1440 7350 -1400
rect 7230 -1470 7275 -1440
rect 7305 -1470 7350 -1440
rect 7230 -1510 7350 -1470
rect 7230 -1540 7275 -1510
rect 7305 -1540 7350 -1510
rect 7230 -1580 7350 -1540
rect 7230 -1610 7275 -1580
rect 7305 -1610 7350 -1580
rect 7230 -1645 7350 -1610
rect 7230 -1675 7275 -1645
rect 7305 -1675 7350 -1645
rect 7230 -1705 7350 -1675
rect 7230 -1735 7275 -1705
rect 7305 -1735 7350 -1705
rect 7230 -1770 7350 -1735
rect 7230 -1800 7275 -1770
rect 7305 -1800 7350 -1770
rect 7230 -1840 7350 -1800
rect 7230 -1870 7275 -1840
rect 7305 -1870 7350 -1840
rect 7230 -1910 7350 -1870
rect 7230 -1940 7275 -1910
rect 7305 -1940 7350 -1910
rect 7230 -1980 7350 -1940
rect 7230 -2010 7275 -1980
rect 7305 -2010 7350 -1980
rect 7230 -2045 7350 -2010
rect 7230 -2075 7275 -2045
rect 7305 -2075 7350 -2045
rect 7230 -2105 7350 -2075
rect 7230 -2135 7275 -2105
rect 7305 -2135 7350 -2105
rect 7230 -2170 7350 -2135
rect 7230 -2200 7275 -2170
rect 7305 -2200 7350 -2170
rect 7230 -2240 7350 -2200
rect 7230 -2270 7275 -2240
rect 7305 -2270 7350 -2240
rect 7230 -2310 7350 -2270
rect 7230 -2340 7275 -2310
rect 7305 -2340 7350 -2310
rect 7230 -2380 7350 -2340
rect 7230 -2410 7275 -2380
rect 7305 -2410 7350 -2380
rect 7230 -2445 7350 -2410
rect 7230 -2475 7275 -2445
rect 7305 -2475 7350 -2445
rect 7230 -2505 7350 -2475
rect 7230 -2535 7275 -2505
rect 7305 -2535 7350 -2505
rect 7230 -2570 7350 -2535
rect 7230 -2600 7275 -2570
rect 7305 -2600 7350 -2570
rect 7230 -2640 7350 -2600
rect 7230 -2670 7275 -2640
rect 7305 -2670 7350 -2640
rect 7230 -2710 7350 -2670
rect 7230 -2740 7275 -2710
rect 7305 -2740 7350 -2710
rect 7230 -2780 7350 -2740
rect 7230 -2810 7275 -2780
rect 7305 -2810 7350 -2780
rect 7230 -2845 7350 -2810
rect 7230 -2875 7275 -2845
rect 7305 -2875 7350 -2845
rect 7230 -2905 7350 -2875
rect 7230 -2935 7275 -2905
rect 7305 -2935 7350 -2905
rect 7230 -2970 7350 -2935
rect 7230 -3000 7275 -2970
rect 7305 -3000 7350 -2970
rect 7230 -3040 7350 -3000
rect 7230 -3070 7275 -3040
rect 7305 -3070 7350 -3040
rect 7230 -3110 7350 -3070
rect 7230 -3140 7275 -3110
rect 7305 -3140 7350 -3110
rect 7230 -3180 7350 -3140
rect 7230 -3210 7275 -3180
rect 7305 -3210 7350 -3180
rect 7230 -3245 7350 -3210
rect 7230 -3275 7275 -3245
rect 7305 -3275 7350 -3245
rect 7230 -3305 7350 -3275
rect 7230 -3335 7275 -3305
rect 7305 -3335 7350 -3305
rect 7230 -3370 7350 -3335
rect 7230 -3400 7275 -3370
rect 7305 -3400 7350 -3370
rect 7230 -3440 7350 -3400
rect 7230 -3470 7275 -3440
rect 7305 -3470 7350 -3440
rect 7230 -3510 7350 -3470
rect 7230 -3540 7275 -3510
rect 7305 -3540 7350 -3510
rect 7230 -3580 7350 -3540
rect 7230 -3610 7275 -3580
rect 7305 -3610 7350 -3580
rect 7230 -3645 7350 -3610
rect 7230 -3675 7275 -3645
rect 7305 -3675 7350 -3645
rect 7230 -3705 7350 -3675
rect 7230 -3735 7275 -3705
rect 7305 -3735 7350 -3705
rect 7230 -3770 7350 -3735
rect 7230 -3800 7275 -3770
rect 7305 -3800 7350 -3770
rect 7230 -3840 7350 -3800
rect 7230 -3870 7275 -3840
rect 7305 -3870 7350 -3840
rect 7230 -3910 7350 -3870
rect 7230 -3940 7275 -3910
rect 7305 -3940 7350 -3910
rect 7230 -3980 7350 -3940
rect 7230 -4010 7275 -3980
rect 7305 -4010 7350 -3980
rect 7230 -4045 7350 -4010
rect 7230 -4075 7275 -4045
rect 7305 -4075 7350 -4045
rect 7230 -4105 7350 -4075
rect 7230 -4135 7275 -4105
rect 7305 -4135 7350 -4105
rect 7230 -4170 7350 -4135
rect 7230 -4200 7275 -4170
rect 7305 -4200 7350 -4170
rect 7230 -4240 7350 -4200
rect 7230 -4270 7275 -4240
rect 7305 -4270 7350 -4240
rect 7230 -4310 7350 -4270
rect 7230 -4340 7275 -4310
rect 7305 -4340 7350 -4310
rect 7230 -4380 7350 -4340
rect 7230 -4410 7275 -4380
rect 7305 -4410 7350 -4380
rect 7230 -4445 7350 -4410
rect 7230 -4475 7275 -4445
rect 7305 -4475 7350 -4445
rect 7230 -4490 7350 -4475
rect 7580 -1305 7700 -1240
rect 7580 -1335 7625 -1305
rect 7655 -1335 7700 -1305
rect 7580 -1370 7700 -1335
rect 7580 -1400 7625 -1370
rect 7655 -1400 7700 -1370
rect 7580 -1440 7700 -1400
rect 7580 -1470 7625 -1440
rect 7655 -1470 7700 -1440
rect 7580 -1510 7700 -1470
rect 7580 -1540 7625 -1510
rect 7655 -1540 7700 -1510
rect 7580 -1580 7700 -1540
rect 7580 -1610 7625 -1580
rect 7655 -1610 7700 -1580
rect 7580 -1645 7700 -1610
rect 7580 -1675 7625 -1645
rect 7655 -1675 7700 -1645
rect 7580 -1705 7700 -1675
rect 7580 -1735 7625 -1705
rect 7655 -1735 7700 -1705
rect 7580 -1770 7700 -1735
rect 7580 -1800 7625 -1770
rect 7655 -1800 7700 -1770
rect 7580 -1840 7700 -1800
rect 7580 -1870 7625 -1840
rect 7655 -1870 7700 -1840
rect 7580 -1910 7700 -1870
rect 7580 -1940 7625 -1910
rect 7655 -1940 7700 -1910
rect 7580 -1980 7700 -1940
rect 7580 -2010 7625 -1980
rect 7655 -2010 7700 -1980
rect 7580 -2045 7700 -2010
rect 7580 -2075 7625 -2045
rect 7655 -2075 7700 -2045
rect 7580 -2105 7700 -2075
rect 7580 -2135 7625 -2105
rect 7655 -2135 7700 -2105
rect 7580 -2170 7700 -2135
rect 7580 -2200 7625 -2170
rect 7655 -2200 7700 -2170
rect 7580 -2240 7700 -2200
rect 7580 -2270 7625 -2240
rect 7655 -2270 7700 -2240
rect 7580 -2310 7700 -2270
rect 7580 -2340 7625 -2310
rect 7655 -2340 7700 -2310
rect 7580 -2380 7700 -2340
rect 7580 -2410 7625 -2380
rect 7655 -2410 7700 -2380
rect 7580 -2445 7700 -2410
rect 7580 -2475 7625 -2445
rect 7655 -2475 7700 -2445
rect 7580 -2505 7700 -2475
rect 7580 -2535 7625 -2505
rect 7655 -2535 7700 -2505
rect 7580 -2570 7700 -2535
rect 7580 -2600 7625 -2570
rect 7655 -2600 7700 -2570
rect 7580 -2640 7700 -2600
rect 7580 -2670 7625 -2640
rect 7655 -2670 7700 -2640
rect 7580 -2710 7700 -2670
rect 7580 -2740 7625 -2710
rect 7655 -2740 7700 -2710
rect 7580 -2780 7700 -2740
rect 7580 -2810 7625 -2780
rect 7655 -2810 7700 -2780
rect 7580 -2845 7700 -2810
rect 7580 -2875 7625 -2845
rect 7655 -2875 7700 -2845
rect 7580 -2905 7700 -2875
rect 7580 -2935 7625 -2905
rect 7655 -2935 7700 -2905
rect 7580 -2970 7700 -2935
rect 7580 -3000 7625 -2970
rect 7655 -3000 7700 -2970
rect 7580 -3040 7700 -3000
rect 7580 -3070 7625 -3040
rect 7655 -3070 7700 -3040
rect 7580 -3110 7700 -3070
rect 7580 -3140 7625 -3110
rect 7655 -3140 7700 -3110
rect 7580 -3180 7700 -3140
rect 7580 -3210 7625 -3180
rect 7655 -3210 7700 -3180
rect 7580 -3245 7700 -3210
rect 7580 -3275 7625 -3245
rect 7655 -3275 7700 -3245
rect 7580 -3305 7700 -3275
rect 7580 -3335 7625 -3305
rect 7655 -3335 7700 -3305
rect 7580 -3370 7700 -3335
rect 7580 -3400 7625 -3370
rect 7655 -3400 7700 -3370
rect 7580 -3440 7700 -3400
rect 7580 -3470 7625 -3440
rect 7655 -3470 7700 -3440
rect 7580 -3510 7700 -3470
rect 7580 -3540 7625 -3510
rect 7655 -3540 7700 -3510
rect 7580 -3580 7700 -3540
rect 7580 -3610 7625 -3580
rect 7655 -3610 7700 -3580
rect 7580 -3645 7700 -3610
rect 7580 -3675 7625 -3645
rect 7655 -3675 7700 -3645
rect 7580 -3705 7700 -3675
rect 7580 -3735 7625 -3705
rect 7655 -3735 7700 -3705
rect 7580 -3770 7700 -3735
rect 7580 -3800 7625 -3770
rect 7655 -3800 7700 -3770
rect 7580 -3840 7700 -3800
rect 7580 -3870 7625 -3840
rect 7655 -3870 7700 -3840
rect 7580 -3910 7700 -3870
rect 7580 -3940 7625 -3910
rect 7655 -3940 7700 -3910
rect 7580 -3980 7700 -3940
rect 7580 -4010 7625 -3980
rect 7655 -4010 7700 -3980
rect 7580 -4045 7700 -4010
rect 7580 -4075 7625 -4045
rect 7655 -4075 7700 -4045
rect 7580 -4105 7700 -4075
rect 7580 -4135 7625 -4105
rect 7655 -4135 7700 -4105
rect 7580 -4170 7700 -4135
rect 7580 -4200 7625 -4170
rect 7655 -4200 7700 -4170
rect 7580 -4240 7700 -4200
rect 7580 -4270 7625 -4240
rect 7655 -4270 7700 -4240
rect 7580 -4310 7700 -4270
rect 7580 -4340 7625 -4310
rect 7655 -4340 7700 -4310
rect 7580 -4380 7700 -4340
rect 7580 -4410 7625 -4380
rect 7655 -4410 7700 -4380
rect 7580 -4445 7700 -4410
rect 7580 -4475 7625 -4445
rect 7655 -4475 7700 -4445
rect 7580 -4490 7700 -4475
rect 7930 -1305 8050 -1240
rect 7930 -1335 7975 -1305
rect 8005 -1335 8050 -1305
rect 7930 -1370 8050 -1335
rect 7930 -1400 7975 -1370
rect 8005 -1400 8050 -1370
rect 7930 -1440 8050 -1400
rect 7930 -1470 7975 -1440
rect 8005 -1470 8050 -1440
rect 7930 -1510 8050 -1470
rect 7930 -1540 7975 -1510
rect 8005 -1540 8050 -1510
rect 7930 -1580 8050 -1540
rect 7930 -1610 7975 -1580
rect 8005 -1610 8050 -1580
rect 7930 -1645 8050 -1610
rect 7930 -1675 7975 -1645
rect 8005 -1675 8050 -1645
rect 7930 -1705 8050 -1675
rect 7930 -1735 7975 -1705
rect 8005 -1735 8050 -1705
rect 7930 -1770 8050 -1735
rect 7930 -1800 7975 -1770
rect 8005 -1800 8050 -1770
rect 7930 -1840 8050 -1800
rect 7930 -1870 7975 -1840
rect 8005 -1870 8050 -1840
rect 7930 -1910 8050 -1870
rect 7930 -1940 7975 -1910
rect 8005 -1940 8050 -1910
rect 7930 -1980 8050 -1940
rect 7930 -2010 7975 -1980
rect 8005 -2010 8050 -1980
rect 7930 -2045 8050 -2010
rect 7930 -2075 7975 -2045
rect 8005 -2075 8050 -2045
rect 7930 -2105 8050 -2075
rect 7930 -2135 7975 -2105
rect 8005 -2135 8050 -2105
rect 7930 -2170 8050 -2135
rect 7930 -2200 7975 -2170
rect 8005 -2200 8050 -2170
rect 7930 -2240 8050 -2200
rect 7930 -2270 7975 -2240
rect 8005 -2270 8050 -2240
rect 7930 -2310 8050 -2270
rect 7930 -2340 7975 -2310
rect 8005 -2340 8050 -2310
rect 7930 -2380 8050 -2340
rect 7930 -2410 7975 -2380
rect 8005 -2410 8050 -2380
rect 7930 -2445 8050 -2410
rect 7930 -2475 7975 -2445
rect 8005 -2475 8050 -2445
rect 7930 -2505 8050 -2475
rect 7930 -2535 7975 -2505
rect 8005 -2535 8050 -2505
rect 7930 -2570 8050 -2535
rect 7930 -2600 7975 -2570
rect 8005 -2600 8050 -2570
rect 7930 -2640 8050 -2600
rect 7930 -2670 7975 -2640
rect 8005 -2670 8050 -2640
rect 7930 -2710 8050 -2670
rect 7930 -2740 7975 -2710
rect 8005 -2740 8050 -2710
rect 7930 -2780 8050 -2740
rect 7930 -2810 7975 -2780
rect 8005 -2810 8050 -2780
rect 7930 -2845 8050 -2810
rect 7930 -2875 7975 -2845
rect 8005 -2875 8050 -2845
rect 7930 -2905 8050 -2875
rect 7930 -2935 7975 -2905
rect 8005 -2935 8050 -2905
rect 7930 -2970 8050 -2935
rect 7930 -3000 7975 -2970
rect 8005 -3000 8050 -2970
rect 7930 -3040 8050 -3000
rect 7930 -3070 7975 -3040
rect 8005 -3070 8050 -3040
rect 7930 -3110 8050 -3070
rect 7930 -3140 7975 -3110
rect 8005 -3140 8050 -3110
rect 7930 -3180 8050 -3140
rect 7930 -3210 7975 -3180
rect 8005 -3210 8050 -3180
rect 7930 -3245 8050 -3210
rect 7930 -3275 7975 -3245
rect 8005 -3275 8050 -3245
rect 7930 -3305 8050 -3275
rect 7930 -3335 7975 -3305
rect 8005 -3335 8050 -3305
rect 7930 -3370 8050 -3335
rect 7930 -3400 7975 -3370
rect 8005 -3400 8050 -3370
rect 7930 -3440 8050 -3400
rect 7930 -3470 7975 -3440
rect 8005 -3470 8050 -3440
rect 7930 -3510 8050 -3470
rect 7930 -3540 7975 -3510
rect 8005 -3540 8050 -3510
rect 7930 -3580 8050 -3540
rect 7930 -3610 7975 -3580
rect 8005 -3610 8050 -3580
rect 7930 -3645 8050 -3610
rect 7930 -3675 7975 -3645
rect 8005 -3675 8050 -3645
rect 7930 -3705 8050 -3675
rect 7930 -3735 7975 -3705
rect 8005 -3735 8050 -3705
rect 7930 -3770 8050 -3735
rect 7930 -3800 7975 -3770
rect 8005 -3800 8050 -3770
rect 7930 -3840 8050 -3800
rect 7930 -3870 7975 -3840
rect 8005 -3870 8050 -3840
rect 7930 -3910 8050 -3870
rect 7930 -3940 7975 -3910
rect 8005 -3940 8050 -3910
rect 7930 -3980 8050 -3940
rect 7930 -4010 7975 -3980
rect 8005 -4010 8050 -3980
rect 7930 -4045 8050 -4010
rect 7930 -4075 7975 -4045
rect 8005 -4075 8050 -4045
rect 7930 -4105 8050 -4075
rect 7930 -4135 7975 -4105
rect 8005 -4135 8050 -4105
rect 7930 -4170 8050 -4135
rect 7930 -4200 7975 -4170
rect 8005 -4200 8050 -4170
rect 7930 -4240 8050 -4200
rect 7930 -4270 7975 -4240
rect 8005 -4270 8050 -4240
rect 7930 -4310 8050 -4270
rect 7930 -4340 7975 -4310
rect 8005 -4340 8050 -4310
rect 7930 -4380 8050 -4340
rect 7930 -4410 7975 -4380
rect 8005 -4410 8050 -4380
rect 7930 -4445 8050 -4410
rect 7930 -4475 7975 -4445
rect 8005 -4475 8050 -4445
rect 7930 -4490 8050 -4475
rect 8280 -1305 8400 -1240
rect 8280 -1335 8325 -1305
rect 8355 -1335 8400 -1305
rect 8280 -1370 8400 -1335
rect 8280 -1400 8325 -1370
rect 8355 -1400 8400 -1370
rect 8280 -1440 8400 -1400
rect 8280 -1470 8325 -1440
rect 8355 -1470 8400 -1440
rect 8280 -1510 8400 -1470
rect 8280 -1540 8325 -1510
rect 8355 -1540 8400 -1510
rect 8280 -1580 8400 -1540
rect 8280 -1610 8325 -1580
rect 8355 -1610 8400 -1580
rect 8280 -1645 8400 -1610
rect 8280 -1675 8325 -1645
rect 8355 -1675 8400 -1645
rect 8280 -1705 8400 -1675
rect 8280 -1735 8325 -1705
rect 8355 -1735 8400 -1705
rect 8280 -1770 8400 -1735
rect 8280 -1800 8325 -1770
rect 8355 -1800 8400 -1770
rect 8280 -1840 8400 -1800
rect 8280 -1870 8325 -1840
rect 8355 -1870 8400 -1840
rect 8280 -1910 8400 -1870
rect 8280 -1940 8325 -1910
rect 8355 -1940 8400 -1910
rect 8280 -1980 8400 -1940
rect 8280 -2010 8325 -1980
rect 8355 -2010 8400 -1980
rect 8280 -2045 8400 -2010
rect 8280 -2075 8325 -2045
rect 8355 -2075 8400 -2045
rect 8280 -2105 8400 -2075
rect 8280 -2135 8325 -2105
rect 8355 -2135 8400 -2105
rect 8280 -2170 8400 -2135
rect 8280 -2200 8325 -2170
rect 8355 -2200 8400 -2170
rect 8280 -2240 8400 -2200
rect 8280 -2270 8325 -2240
rect 8355 -2270 8400 -2240
rect 8280 -2310 8400 -2270
rect 8280 -2340 8325 -2310
rect 8355 -2340 8400 -2310
rect 8280 -2380 8400 -2340
rect 8280 -2410 8325 -2380
rect 8355 -2410 8400 -2380
rect 8280 -2445 8400 -2410
rect 8280 -2475 8325 -2445
rect 8355 -2475 8400 -2445
rect 8280 -2505 8400 -2475
rect 8280 -2535 8325 -2505
rect 8355 -2535 8400 -2505
rect 8280 -2570 8400 -2535
rect 8280 -2600 8325 -2570
rect 8355 -2600 8400 -2570
rect 8280 -2640 8400 -2600
rect 8280 -2670 8325 -2640
rect 8355 -2670 8400 -2640
rect 8280 -2710 8400 -2670
rect 8280 -2740 8325 -2710
rect 8355 -2740 8400 -2710
rect 8280 -2780 8400 -2740
rect 8280 -2810 8325 -2780
rect 8355 -2810 8400 -2780
rect 8280 -2845 8400 -2810
rect 8280 -2875 8325 -2845
rect 8355 -2875 8400 -2845
rect 8280 -2905 8400 -2875
rect 8280 -2935 8325 -2905
rect 8355 -2935 8400 -2905
rect 8280 -2970 8400 -2935
rect 8280 -3000 8325 -2970
rect 8355 -3000 8400 -2970
rect 8280 -3040 8400 -3000
rect 8280 -3070 8325 -3040
rect 8355 -3070 8400 -3040
rect 8280 -3110 8400 -3070
rect 8280 -3140 8325 -3110
rect 8355 -3140 8400 -3110
rect 8280 -3180 8400 -3140
rect 8280 -3210 8325 -3180
rect 8355 -3210 8400 -3180
rect 8280 -3245 8400 -3210
rect 8280 -3275 8325 -3245
rect 8355 -3275 8400 -3245
rect 8280 -3305 8400 -3275
rect 8280 -3335 8325 -3305
rect 8355 -3335 8400 -3305
rect 8280 -3370 8400 -3335
rect 8280 -3400 8325 -3370
rect 8355 -3400 8400 -3370
rect 8280 -3440 8400 -3400
rect 8280 -3470 8325 -3440
rect 8355 -3470 8400 -3440
rect 8280 -3510 8400 -3470
rect 8280 -3540 8325 -3510
rect 8355 -3540 8400 -3510
rect 8280 -3580 8400 -3540
rect 8280 -3610 8325 -3580
rect 8355 -3610 8400 -3580
rect 8280 -3645 8400 -3610
rect 8280 -3675 8325 -3645
rect 8355 -3675 8400 -3645
rect 8280 -3705 8400 -3675
rect 8280 -3735 8325 -3705
rect 8355 -3735 8400 -3705
rect 8280 -3770 8400 -3735
rect 8280 -3800 8325 -3770
rect 8355 -3800 8400 -3770
rect 8280 -3840 8400 -3800
rect 8280 -3870 8325 -3840
rect 8355 -3870 8400 -3840
rect 8280 -3910 8400 -3870
rect 8280 -3940 8325 -3910
rect 8355 -3940 8400 -3910
rect 8280 -3980 8400 -3940
rect 8280 -4010 8325 -3980
rect 8355 -4010 8400 -3980
rect 8280 -4045 8400 -4010
rect 8280 -4075 8325 -4045
rect 8355 -4075 8400 -4045
rect 8280 -4105 8400 -4075
rect 8280 -4135 8325 -4105
rect 8355 -4135 8400 -4105
rect 8280 -4170 8400 -4135
rect 8280 -4200 8325 -4170
rect 8355 -4200 8400 -4170
rect 8280 -4240 8400 -4200
rect 8280 -4270 8325 -4240
rect 8355 -4270 8400 -4240
rect 8280 -4310 8400 -4270
rect 8280 -4340 8325 -4310
rect 8355 -4340 8400 -4310
rect 8280 -4380 8400 -4340
rect 8280 -4410 8325 -4380
rect 8355 -4410 8400 -4380
rect 8280 -4445 8400 -4410
rect 8280 -4475 8325 -4445
rect 8355 -4475 8400 -4445
rect 8280 -4490 8400 -4475
rect 8630 -1305 8750 -1240
rect 8630 -1335 8675 -1305
rect 8705 -1335 8750 -1305
rect 8630 -1370 8750 -1335
rect 8630 -1400 8675 -1370
rect 8705 -1400 8750 -1370
rect 8630 -1440 8750 -1400
rect 8630 -1470 8675 -1440
rect 8705 -1470 8750 -1440
rect 8630 -1510 8750 -1470
rect 8630 -1540 8675 -1510
rect 8705 -1540 8750 -1510
rect 8630 -1580 8750 -1540
rect 8630 -1610 8675 -1580
rect 8705 -1610 8750 -1580
rect 8630 -1645 8750 -1610
rect 8630 -1675 8675 -1645
rect 8705 -1675 8750 -1645
rect 8630 -1705 8750 -1675
rect 8630 -1735 8675 -1705
rect 8705 -1735 8750 -1705
rect 8630 -1770 8750 -1735
rect 8630 -1800 8675 -1770
rect 8705 -1800 8750 -1770
rect 8630 -1840 8750 -1800
rect 8630 -1870 8675 -1840
rect 8705 -1870 8750 -1840
rect 8630 -1910 8750 -1870
rect 8630 -1940 8675 -1910
rect 8705 -1940 8750 -1910
rect 8630 -1980 8750 -1940
rect 8630 -2010 8675 -1980
rect 8705 -2010 8750 -1980
rect 8630 -2045 8750 -2010
rect 8630 -2075 8675 -2045
rect 8705 -2075 8750 -2045
rect 8630 -2105 8750 -2075
rect 8630 -2135 8675 -2105
rect 8705 -2135 8750 -2105
rect 8630 -2170 8750 -2135
rect 8630 -2200 8675 -2170
rect 8705 -2200 8750 -2170
rect 8630 -2240 8750 -2200
rect 8630 -2270 8675 -2240
rect 8705 -2270 8750 -2240
rect 8630 -2310 8750 -2270
rect 8630 -2340 8675 -2310
rect 8705 -2340 8750 -2310
rect 8630 -2380 8750 -2340
rect 8630 -2410 8675 -2380
rect 8705 -2410 8750 -2380
rect 8630 -2445 8750 -2410
rect 8630 -2475 8675 -2445
rect 8705 -2475 8750 -2445
rect 8630 -2505 8750 -2475
rect 8630 -2535 8675 -2505
rect 8705 -2535 8750 -2505
rect 8630 -2570 8750 -2535
rect 8630 -2600 8675 -2570
rect 8705 -2600 8750 -2570
rect 8630 -2640 8750 -2600
rect 8630 -2670 8675 -2640
rect 8705 -2670 8750 -2640
rect 8630 -2710 8750 -2670
rect 8630 -2740 8675 -2710
rect 8705 -2740 8750 -2710
rect 8630 -2780 8750 -2740
rect 8630 -2810 8675 -2780
rect 8705 -2810 8750 -2780
rect 8630 -2845 8750 -2810
rect 8630 -2875 8675 -2845
rect 8705 -2875 8750 -2845
rect 8630 -2905 8750 -2875
rect 8630 -2935 8675 -2905
rect 8705 -2935 8750 -2905
rect 8630 -2970 8750 -2935
rect 8630 -3000 8675 -2970
rect 8705 -3000 8750 -2970
rect 8630 -3040 8750 -3000
rect 8630 -3070 8675 -3040
rect 8705 -3070 8750 -3040
rect 8630 -3110 8750 -3070
rect 8630 -3140 8675 -3110
rect 8705 -3140 8750 -3110
rect 8630 -3180 8750 -3140
rect 8630 -3210 8675 -3180
rect 8705 -3210 8750 -3180
rect 8630 -3245 8750 -3210
rect 8630 -3275 8675 -3245
rect 8705 -3275 8750 -3245
rect 8630 -3305 8750 -3275
rect 8630 -3335 8675 -3305
rect 8705 -3335 8750 -3305
rect 8630 -3370 8750 -3335
rect 8630 -3400 8675 -3370
rect 8705 -3400 8750 -3370
rect 8630 -3440 8750 -3400
rect 8630 -3470 8675 -3440
rect 8705 -3470 8750 -3440
rect 8630 -3510 8750 -3470
rect 8630 -3540 8675 -3510
rect 8705 -3540 8750 -3510
rect 8630 -3580 8750 -3540
rect 8630 -3610 8675 -3580
rect 8705 -3610 8750 -3580
rect 8630 -3645 8750 -3610
rect 8630 -3675 8675 -3645
rect 8705 -3675 8750 -3645
rect 8630 -3705 8750 -3675
rect 8630 -3735 8675 -3705
rect 8705 -3735 8750 -3705
rect 8630 -3770 8750 -3735
rect 8630 -3800 8675 -3770
rect 8705 -3800 8750 -3770
rect 8630 -3840 8750 -3800
rect 8630 -3870 8675 -3840
rect 8705 -3870 8750 -3840
rect 8630 -3910 8750 -3870
rect 8630 -3940 8675 -3910
rect 8705 -3940 8750 -3910
rect 8630 -3980 8750 -3940
rect 8630 -4010 8675 -3980
rect 8705 -4010 8750 -3980
rect 8630 -4045 8750 -4010
rect 8630 -4075 8675 -4045
rect 8705 -4075 8750 -4045
rect 8630 -4105 8750 -4075
rect 8630 -4135 8675 -4105
rect 8705 -4135 8750 -4105
rect 8630 -4170 8750 -4135
rect 8630 -4200 8675 -4170
rect 8705 -4200 8750 -4170
rect 8630 -4240 8750 -4200
rect 8630 -4270 8675 -4240
rect 8705 -4270 8750 -4240
rect 8630 -4310 8750 -4270
rect 8630 -4340 8675 -4310
rect 8705 -4340 8750 -4310
rect 8630 -4380 8750 -4340
rect 8630 -4410 8675 -4380
rect 8705 -4410 8750 -4380
rect 8630 -4445 8750 -4410
rect 8630 -4475 8675 -4445
rect 8705 -4475 8750 -4445
rect 8630 -4490 8750 -4475
rect 8980 -1305 9100 -1290
rect 8980 -1335 9025 -1305
rect 9055 -1335 9100 -1305
rect 8980 -1370 9100 -1335
rect 8980 -1400 9025 -1370
rect 9055 -1400 9100 -1370
rect 8980 -1440 9100 -1400
rect 8980 -1470 9025 -1440
rect 9055 -1470 9100 -1440
rect 8980 -1510 9100 -1470
rect 8980 -1540 9025 -1510
rect 9055 -1540 9100 -1510
rect 8980 -1580 9100 -1540
rect 8980 -1610 9025 -1580
rect 9055 -1610 9100 -1580
rect 8980 -1645 9100 -1610
rect 8980 -1675 9025 -1645
rect 9055 -1675 9100 -1645
rect 8980 -1705 9100 -1675
rect 8980 -1735 9025 -1705
rect 9055 -1735 9100 -1705
rect 8980 -1770 9100 -1735
rect 8980 -1800 9025 -1770
rect 9055 -1800 9100 -1770
rect 8980 -1840 9100 -1800
rect 8980 -1870 9025 -1840
rect 9055 -1870 9100 -1840
rect 8980 -1910 9100 -1870
rect 8980 -1940 9025 -1910
rect 9055 -1940 9100 -1910
rect 8980 -1980 9100 -1940
rect 8980 -2010 9025 -1980
rect 9055 -2010 9100 -1980
rect 8980 -2045 9100 -2010
rect 8980 -2075 9025 -2045
rect 9055 -2075 9100 -2045
rect 8980 -2105 9100 -2075
rect 8980 -2135 9025 -2105
rect 9055 -2135 9100 -2105
rect 8980 -2170 9100 -2135
rect 8980 -2200 9025 -2170
rect 9055 -2200 9100 -2170
rect 8980 -2240 9100 -2200
rect 8980 -2270 9025 -2240
rect 9055 -2270 9100 -2240
rect 8980 -2310 9100 -2270
rect 8980 -2340 9025 -2310
rect 9055 -2340 9100 -2310
rect 8980 -2380 9100 -2340
rect 8980 -2410 9025 -2380
rect 9055 -2410 9100 -2380
rect 8980 -2445 9100 -2410
rect 8980 -2475 9025 -2445
rect 9055 -2475 9100 -2445
rect 8980 -2505 9100 -2475
rect 8980 -2535 9025 -2505
rect 9055 -2535 9100 -2505
rect 8980 -2570 9100 -2535
rect 8980 -2600 9025 -2570
rect 9055 -2600 9100 -2570
rect 8980 -2640 9100 -2600
rect 8980 -2670 9025 -2640
rect 9055 -2670 9100 -2640
rect 8980 -2710 9100 -2670
rect 8980 -2740 9025 -2710
rect 9055 -2740 9100 -2710
rect 8980 -2780 9100 -2740
rect 8980 -2810 9025 -2780
rect 9055 -2810 9100 -2780
rect 8980 -2845 9100 -2810
rect 8980 -2875 9025 -2845
rect 9055 -2875 9100 -2845
rect 8980 -2905 9100 -2875
rect 8980 -2935 9025 -2905
rect 9055 -2935 9100 -2905
rect 8980 -2970 9100 -2935
rect 8980 -3000 9025 -2970
rect 9055 -3000 9100 -2970
rect 8980 -3040 9100 -3000
rect 8980 -3070 9025 -3040
rect 9055 -3070 9100 -3040
rect 8980 -3110 9100 -3070
rect 8980 -3140 9025 -3110
rect 9055 -3140 9100 -3110
rect 8980 -3180 9100 -3140
rect 8980 -3210 9025 -3180
rect 9055 -3210 9100 -3180
rect 8980 -3245 9100 -3210
rect 8980 -3275 9025 -3245
rect 9055 -3275 9100 -3245
rect 8980 -3305 9100 -3275
rect 8980 -3335 9025 -3305
rect 9055 -3335 9100 -3305
rect 8980 -3370 9100 -3335
rect 8980 -3400 9025 -3370
rect 9055 -3400 9100 -3370
rect 8980 -3440 9100 -3400
rect 8980 -3470 9025 -3440
rect 9055 -3470 9100 -3440
rect 8980 -3510 9100 -3470
rect 8980 -3540 9025 -3510
rect 9055 -3540 9100 -3510
rect 8980 -3580 9100 -3540
rect 8980 -3610 9025 -3580
rect 9055 -3610 9100 -3580
rect 8980 -3645 9100 -3610
rect 8980 -3675 9025 -3645
rect 9055 -3675 9100 -3645
rect 8980 -3705 9100 -3675
rect 8980 -3735 9025 -3705
rect 9055 -3735 9100 -3705
rect 8980 -3770 9100 -3735
rect 8980 -3800 9025 -3770
rect 9055 -3800 9100 -3770
rect 8980 -3840 9100 -3800
rect 8980 -3870 9025 -3840
rect 9055 -3870 9100 -3840
rect 8980 -3910 9100 -3870
rect 8980 -3940 9025 -3910
rect 9055 -3940 9100 -3910
rect 8980 -3980 9100 -3940
rect 8980 -4010 9025 -3980
rect 9055 -4010 9100 -3980
rect 8980 -4045 9100 -4010
rect 8980 -4075 9025 -4045
rect 9055 -4075 9100 -4045
rect 8980 -4105 9100 -4075
rect 8980 -4135 9025 -4105
rect 9055 -4135 9100 -4105
rect 8980 -4170 9100 -4135
rect 8980 -4200 9025 -4170
rect 9055 -4200 9100 -4170
rect 8980 -4240 9100 -4200
rect 8980 -4270 9025 -4240
rect 9055 -4270 9100 -4240
rect 8980 -4310 9100 -4270
rect 8980 -4340 9025 -4310
rect 9055 -4340 9100 -4310
rect 8980 -4380 9100 -4340
rect 8980 -4410 9025 -4380
rect 9055 -4410 9100 -4380
rect 8980 -4445 9100 -4410
rect 8980 -4475 9025 -4445
rect 9055 -4475 9100 -4445
rect 8980 -4490 9100 -4475
<< via1 >>
rect 2195 20880 2225 20910
rect 2195 20815 2225 20845
rect 2195 20745 2225 20775
rect 2195 20675 2225 20705
rect 2195 20605 2225 20635
rect 2195 20540 2225 20570
rect 2195 20480 2225 20510
rect 2195 20415 2225 20445
rect 2195 20345 2225 20375
rect 2195 20275 2225 20305
rect 2195 20205 2225 20235
rect 2195 20140 2225 20170
rect 2195 20080 2225 20110
rect 2195 20015 2225 20045
rect 2195 19945 2225 19975
rect 2195 19875 2225 19905
rect 2195 19805 2225 19835
rect 2195 19740 2225 19770
rect 2195 19680 2225 19710
rect 2195 19615 2225 19645
rect 2195 19545 2225 19575
rect 2195 19475 2225 19505
rect 2195 19405 2225 19435
rect 2195 19340 2225 19370
rect 2195 19280 2225 19310
rect 2195 19215 2225 19245
rect 2195 19145 2225 19175
rect 2195 19075 2225 19105
rect 2195 19005 2225 19035
rect 2195 18940 2225 18970
rect 2195 18880 2225 18910
rect 2195 18815 2225 18845
rect 2195 18745 2225 18775
rect 2195 18675 2225 18705
rect 2195 18605 2225 18635
rect 2195 18540 2225 18570
rect 2195 18480 2225 18510
rect 2195 18415 2225 18445
rect 2195 18345 2225 18375
rect 2195 18275 2225 18305
rect 2195 18205 2225 18235
rect 2195 18140 2225 18170
rect 2195 18080 2225 18110
rect 2195 18015 2225 18045
rect 2195 17945 2225 17975
rect 2195 17875 2225 17905
rect 2195 17805 2225 17835
rect 2195 17740 2225 17770
rect 6665 20880 6695 20910
rect 6665 20815 6695 20845
rect 6665 20745 6695 20775
rect 6665 20675 6695 20705
rect 6665 20605 6695 20635
rect 6665 20540 6695 20570
rect 6665 20480 6695 20510
rect 6665 20415 6695 20445
rect 6665 20345 6695 20375
rect 6665 20275 6695 20305
rect 6665 20205 6695 20235
rect 6665 20140 6695 20170
rect 6665 20080 6695 20110
rect 6665 20015 6695 20045
rect 6665 19945 6695 19975
rect 6665 19875 6695 19905
rect 6665 19805 6695 19835
rect 6665 19740 6695 19770
rect 6665 19680 6695 19710
rect 6665 19615 6695 19645
rect 6665 19545 6695 19575
rect 6665 19475 6695 19505
rect 6665 19405 6695 19435
rect 6665 19340 6695 19370
rect 6665 19280 6695 19310
rect 6665 19215 6695 19245
rect 6665 19145 6695 19175
rect 6665 19075 6695 19105
rect 6665 19005 6695 19035
rect 6665 18940 6695 18970
rect 6665 18880 6695 18910
rect 6665 18815 6695 18845
rect 6665 18745 6695 18775
rect 6665 18675 6695 18705
rect 6665 18605 6695 18635
rect 6665 18540 6695 18570
rect 6665 18480 6695 18510
rect 6665 18415 6695 18445
rect 6665 18345 6695 18375
rect 6665 18275 6695 18305
rect 6665 18205 6695 18235
rect 6665 18140 6695 18170
rect 6665 18080 6695 18110
rect 6665 18015 6695 18045
rect 6665 17945 6695 17975
rect 6665 17875 6695 17905
rect 6665 17805 6695 17835
rect 6665 17740 6695 17770
rect 2155 15750 2185 15780
rect 2195 15750 2225 15780
rect 2235 15750 2265 15780
rect 2155 15710 2185 15740
rect 2195 15710 2225 15740
rect 2235 15710 2265 15740
rect 2155 15670 2185 15700
rect 2195 15670 2225 15700
rect 2235 15670 2265 15700
rect 2155 12690 2185 12720
rect 2195 12690 2225 12720
rect 2235 12690 2265 12720
rect 2155 12650 2185 12680
rect 2195 12650 2225 12680
rect 2235 12650 2265 12680
rect 2155 12530 2185 12560
rect 2195 12530 2225 12560
rect 2235 12530 2265 12560
rect 2155 12490 2185 12520
rect 2195 12490 2225 12520
rect 2235 12490 2265 12520
rect 2155 12450 2185 12480
rect 2195 12450 2225 12480
rect 2235 12450 2265 12480
rect 2290 15895 2320 15925
rect 2330 15895 2360 15925
rect 2370 15895 2400 15925
rect -75 9605 -45 9635
rect -75 9540 -45 9570
rect -75 9470 -45 9500
rect -75 9400 -45 9430
rect -75 9330 -45 9360
rect -75 9265 -45 9295
rect -75 9205 -45 9235
rect -75 9140 -45 9170
rect -75 9070 -45 9100
rect -75 9000 -45 9030
rect -75 8930 -45 8960
rect -75 8865 -45 8895
rect -75 8805 -45 8835
rect -75 8740 -45 8770
rect -75 8670 -45 8700
rect -75 8600 -45 8630
rect -75 8530 -45 8560
rect -75 8465 -45 8495
rect -75 8405 -45 8435
rect -75 8340 -45 8370
rect -75 8270 -45 8300
rect -75 8200 -45 8230
rect -75 8130 -45 8160
rect -75 8065 -45 8095
rect -75 8005 -45 8035
rect -75 7940 -45 7970
rect -75 7870 -45 7900
rect -75 7800 -45 7830
rect -75 7730 -45 7760
rect -75 7665 -45 7695
rect -75 7605 -45 7635
rect -75 7540 -45 7570
rect -75 7470 -45 7500
rect -75 7400 -45 7430
rect -75 7330 -45 7360
rect -75 7265 -45 7295
rect -75 7205 -45 7235
rect -75 7140 -45 7170
rect -75 7070 -45 7100
rect -75 7000 -45 7030
rect -75 6930 -45 6960
rect -75 6865 -45 6895
rect -75 6805 -45 6835
rect -75 6740 -45 6770
rect -75 6670 -45 6700
rect -75 6600 -45 6630
rect -75 6530 -45 6560
rect -75 6465 -45 6495
rect 275 9605 305 9635
rect 275 9540 305 9570
rect 275 9470 305 9500
rect 275 9400 305 9430
rect 275 9330 305 9360
rect 275 9265 305 9295
rect 275 9205 305 9235
rect 275 9140 305 9170
rect 275 9070 305 9100
rect 275 9000 305 9030
rect 275 8930 305 8960
rect 275 8865 305 8895
rect 275 8805 305 8835
rect 275 8740 305 8770
rect 275 8670 305 8700
rect 275 8600 305 8630
rect 275 8530 305 8560
rect 275 8465 305 8495
rect 275 8405 305 8435
rect 275 8340 305 8370
rect 275 8270 305 8300
rect 275 8200 305 8230
rect 275 8130 305 8160
rect 275 8065 305 8095
rect 275 8005 305 8035
rect 275 7940 305 7970
rect 275 7870 305 7900
rect 275 7800 305 7830
rect 275 7730 305 7760
rect 275 7665 305 7695
rect 275 7605 305 7635
rect 275 7540 305 7570
rect 275 7470 305 7500
rect 275 7400 305 7430
rect 275 7330 305 7360
rect 275 7265 305 7295
rect 275 7205 305 7235
rect 275 7140 305 7170
rect 275 7070 305 7100
rect 275 7000 305 7030
rect 275 6930 305 6960
rect 275 6865 305 6895
rect 275 6805 305 6835
rect 275 6740 305 6770
rect 275 6670 305 6700
rect 275 6600 305 6630
rect 275 6530 305 6560
rect 275 6465 305 6495
rect 625 9605 655 9635
rect 625 9540 655 9570
rect 625 9470 655 9500
rect 625 9400 655 9430
rect 625 9330 655 9360
rect 625 9265 655 9295
rect 625 9205 655 9235
rect 625 9140 655 9170
rect 625 9070 655 9100
rect 625 9000 655 9030
rect 625 8930 655 8960
rect 625 8865 655 8895
rect 625 8805 655 8835
rect 625 8740 655 8770
rect 625 8670 655 8700
rect 625 8600 655 8630
rect 625 8530 655 8560
rect 625 8465 655 8495
rect 625 8405 655 8435
rect 625 8340 655 8370
rect 625 8270 655 8300
rect 625 8200 655 8230
rect 625 8130 655 8160
rect 625 8065 655 8095
rect 625 8005 655 8035
rect 625 7940 655 7970
rect 625 7870 655 7900
rect 625 7800 655 7830
rect 625 7730 655 7760
rect 625 7665 655 7695
rect 625 7605 655 7635
rect 625 7540 655 7570
rect 625 7470 655 7500
rect 625 7400 655 7430
rect 625 7330 655 7360
rect 625 7265 655 7295
rect 625 7205 655 7235
rect 625 7140 655 7170
rect 625 7070 655 7100
rect 625 7000 655 7030
rect 625 6930 655 6960
rect 625 6865 655 6895
rect 625 6805 655 6835
rect 625 6740 655 6770
rect 625 6670 655 6700
rect 625 6600 655 6630
rect 625 6530 655 6560
rect 625 6465 655 6495
rect 975 9605 1005 9635
rect 975 9540 1005 9570
rect 975 9470 1005 9500
rect 975 9400 1005 9430
rect 975 9330 1005 9360
rect 975 9265 1005 9295
rect 975 9205 1005 9235
rect 975 9140 1005 9170
rect 975 9070 1005 9100
rect 975 9000 1005 9030
rect 975 8930 1005 8960
rect 975 8865 1005 8895
rect 975 8805 1005 8835
rect 975 8740 1005 8770
rect 975 8670 1005 8700
rect 975 8600 1005 8630
rect 975 8530 1005 8560
rect 975 8465 1005 8495
rect 975 8405 1005 8435
rect 975 8340 1005 8370
rect 975 8270 1005 8300
rect 975 8200 1005 8230
rect 975 8130 1005 8160
rect 975 8065 1005 8095
rect 975 8005 1005 8035
rect 975 7940 1005 7970
rect 975 7870 1005 7900
rect 975 7800 1005 7830
rect 975 7730 1005 7760
rect 975 7665 1005 7695
rect 975 7605 1005 7635
rect 975 7540 1005 7570
rect 975 7470 1005 7500
rect 975 7400 1005 7430
rect 975 7330 1005 7360
rect 975 7265 1005 7295
rect 975 7205 1005 7235
rect 975 7140 1005 7170
rect 975 7070 1005 7100
rect 975 7000 1005 7030
rect 975 6930 1005 6960
rect 975 6865 1005 6895
rect 975 6805 1005 6835
rect 975 6740 1005 6770
rect 975 6670 1005 6700
rect 975 6600 1005 6630
rect 975 6530 1005 6560
rect 975 6465 1005 6495
rect 1675 9605 1705 9635
rect 1675 9540 1705 9570
rect 1675 9470 1705 9500
rect 1675 9400 1705 9430
rect 1675 9330 1705 9360
rect 1675 9265 1705 9295
rect 1675 9205 1705 9235
rect 1675 9140 1705 9170
rect 1675 9070 1705 9100
rect 1675 9000 1705 9030
rect 1675 8930 1705 8960
rect 1675 8865 1705 8895
rect 1675 8805 1705 8835
rect 1675 8740 1705 8770
rect 1675 8670 1705 8700
rect 1675 8600 1705 8630
rect 1675 8530 1705 8560
rect 1675 8465 1705 8495
rect 1675 8405 1705 8435
rect 1675 8340 1705 8370
rect 1675 8270 1705 8300
rect 1675 8200 1705 8230
rect 1675 8130 1705 8160
rect 1675 8065 1705 8095
rect 1675 8005 1705 8035
rect 1675 7940 1705 7970
rect 1675 7870 1705 7900
rect 1675 7800 1705 7830
rect 1675 7730 1705 7760
rect 1675 7665 1705 7695
rect 1675 7605 1705 7635
rect 1675 7540 1705 7570
rect 1675 7470 1705 7500
rect 1675 7400 1705 7430
rect 1675 7330 1705 7360
rect 1675 7265 1705 7295
rect 1675 7205 1705 7235
rect 1675 7140 1705 7170
rect 1675 7070 1705 7100
rect 1675 7000 1705 7030
rect 1675 6930 1705 6960
rect 1675 6865 1705 6895
rect 1675 6805 1705 6835
rect 1675 6740 1705 6770
rect 1675 6670 1705 6700
rect 1675 6600 1705 6630
rect 1675 6530 1705 6560
rect 1675 6465 1705 6495
rect 2975 15710 3005 15740
rect 2975 15670 3005 15700
rect 3300 15710 3330 15740
rect 3300 15670 3330 15700
rect 6625 15675 6655 15705
rect 6665 15675 6695 15705
rect 6705 15675 6735 15705
rect 5650 15635 5680 15665
rect 5650 15595 5680 15625
rect 5975 15635 6005 15665
rect 5975 15595 6005 15625
rect 6625 15635 6655 15665
rect 6665 15635 6695 15665
rect 6705 15635 6735 15665
rect 6625 15595 6655 15625
rect 6665 15595 6695 15625
rect 6705 15595 6735 15625
rect 6625 12975 6655 13005
rect 6665 12975 6695 13005
rect 6705 12975 6735 13005
rect 6625 12935 6655 12965
rect 6665 12935 6695 12965
rect 6705 12935 6735 12965
rect 6625 12895 6655 12925
rect 6665 12895 6695 12925
rect 6705 12895 6735 12925
rect 6595 12130 6625 12160
rect 6635 12130 6665 12160
rect 6675 12130 6705 12160
rect 6595 12090 6625 12120
rect 6635 12090 6665 12120
rect 6675 12090 6705 12120
rect 6595 12050 6625 12080
rect 6635 12050 6665 12080
rect 6675 12050 6705 12080
rect 6595 11175 6625 11205
rect 6635 11175 6665 11205
rect 6675 11175 6705 11205
rect 6595 11135 6625 11165
rect 6635 11135 6665 11165
rect 6675 11135 6705 11165
rect 6595 11095 6625 11125
rect 6635 11095 6665 11125
rect 6675 11095 6705 11125
rect 2330 9605 2360 9635
rect 2330 9540 2360 9570
rect 2330 9470 2360 9500
rect 2330 9400 2360 9430
rect 2330 9330 2360 9360
rect 2330 9265 2360 9295
rect 2330 9205 2360 9235
rect 2330 9140 2360 9170
rect 2330 9070 2360 9100
rect 2330 9000 2360 9030
rect 2330 8930 2360 8960
rect 2330 8865 2360 8895
rect 2330 8805 2360 8835
rect 2330 8740 2360 8770
rect 2330 8670 2360 8700
rect 2330 8600 2360 8630
rect 2330 8530 2360 8560
rect 2330 8465 2360 8495
rect 2330 8405 2360 8435
rect 2330 8340 2360 8370
rect 2330 8270 2360 8300
rect 2330 8200 2360 8230
rect 2330 8130 2360 8160
rect 2330 8065 2360 8095
rect 2330 8005 2360 8035
rect 2330 7940 2360 7970
rect 2330 7870 2360 7900
rect 2330 7800 2360 7830
rect 2330 7730 2360 7760
rect 2330 7665 2360 7695
rect 2330 7605 2360 7635
rect 2330 7540 2360 7570
rect 2330 7470 2360 7500
rect 2330 7400 2360 7430
rect 2330 7330 2360 7360
rect 2330 7265 2360 7295
rect 2330 7205 2360 7235
rect 2330 7140 2360 7170
rect 2330 7070 2360 7100
rect 2330 7000 2360 7030
rect 2330 6930 2360 6960
rect 2330 6865 2360 6895
rect 2330 6805 2360 6835
rect 2330 6740 2360 6770
rect 2330 6670 2360 6700
rect 2330 6600 2360 6630
rect 2330 6530 2360 6560
rect 2330 6465 2360 6495
rect 2050 6400 2080 6430
rect 2480 6400 2510 6430
rect 2005 6345 2035 6375
rect 1285 6175 1315 6205
rect 1325 6175 1355 6205
rect 1365 6175 1395 6205
rect 1285 6135 1315 6165
rect 1325 6135 1355 6165
rect 1365 6135 1395 6165
rect 1285 6095 1315 6125
rect 1325 6095 1355 6125
rect 1365 6095 1395 6125
rect 2850 6400 2880 6430
rect 2720 6300 2750 6330
rect 6595 10470 6625 10500
rect 6635 10470 6665 10500
rect 6675 10470 6705 10500
rect 6595 10430 6625 10460
rect 6635 10430 6665 10460
rect 6675 10430 6705 10460
rect 6595 10390 6625 10420
rect 6635 10390 6665 10420
rect 6675 10390 6705 10420
rect 6595 10005 6625 10035
rect 6635 10005 6665 10035
rect 6675 10005 6705 10035
rect 6595 9965 6625 9995
rect 6635 9965 6665 9995
rect 6675 9965 6705 9995
rect 6595 9925 6625 9955
rect 6635 9925 6665 9955
rect 6675 9925 6705 9955
rect 3180 9605 3210 9635
rect 3240 9605 3270 9635
rect 3180 9540 3210 9570
rect 3240 9540 3270 9570
rect 3180 9470 3210 9500
rect 3240 9470 3270 9500
rect 3180 9400 3210 9430
rect 3240 9400 3270 9430
rect 3180 9330 3210 9360
rect 3240 9330 3270 9360
rect 3180 9265 3210 9295
rect 3240 9265 3270 9295
rect 3180 9205 3210 9235
rect 3240 9205 3270 9235
rect 3180 9140 3210 9170
rect 3240 9140 3270 9170
rect 3180 9070 3210 9100
rect 3240 9070 3270 9100
rect 3180 9000 3210 9030
rect 3240 9000 3270 9030
rect 3180 8930 3210 8960
rect 3240 8930 3270 8960
rect 3180 8865 3210 8895
rect 3240 8865 3270 8895
rect 3180 8805 3210 8835
rect 3240 8805 3270 8835
rect 3180 8740 3210 8770
rect 3240 8740 3270 8770
rect 3180 8670 3210 8700
rect 3240 8670 3270 8700
rect 3180 8600 3210 8630
rect 3240 8600 3270 8630
rect 3180 8530 3210 8560
rect 3240 8530 3270 8560
rect 3180 8465 3210 8495
rect 3240 8465 3270 8495
rect 3180 8405 3210 8435
rect 3240 8405 3270 8435
rect 3180 8340 3210 8370
rect 3240 8340 3270 8370
rect 3180 8270 3210 8300
rect 3240 8270 3270 8300
rect 3180 8200 3210 8230
rect 3240 8200 3270 8230
rect 3180 8130 3210 8160
rect 3240 8130 3270 8160
rect 3180 8065 3210 8095
rect 3240 8065 3270 8095
rect 3180 8005 3210 8035
rect 3240 8005 3270 8035
rect 3180 7940 3210 7970
rect 3240 7940 3270 7970
rect 3180 7870 3210 7900
rect 3240 7870 3270 7900
rect 3180 7800 3210 7830
rect 3240 7800 3270 7830
rect 3180 7730 3210 7760
rect 3240 7730 3270 7760
rect 3180 7665 3210 7695
rect 3240 7665 3270 7695
rect 3180 7605 3210 7635
rect 3240 7605 3270 7635
rect 3180 7540 3210 7570
rect 3240 7540 3270 7570
rect 3180 7470 3210 7500
rect 3240 7470 3270 7500
rect 3180 7400 3210 7430
rect 3240 7400 3270 7430
rect 3180 7330 3210 7360
rect 3240 7330 3270 7360
rect 3180 7265 3210 7295
rect 3240 7265 3270 7295
rect 3180 7205 3210 7235
rect 3240 7205 3270 7235
rect 3180 7140 3210 7170
rect 3240 7140 3270 7170
rect 3180 7070 3210 7100
rect 3240 7070 3270 7100
rect 3180 7000 3210 7030
rect 3240 7000 3270 7030
rect 3180 6930 3210 6960
rect 3240 6930 3270 6960
rect 3180 6865 3210 6895
rect 3240 6865 3270 6895
rect 3180 6805 3210 6835
rect 3240 6805 3270 6835
rect 3180 6740 3210 6770
rect 3240 6740 3270 6770
rect 3180 6670 3210 6700
rect 3240 6670 3270 6700
rect 3180 6600 3210 6630
rect 3240 6600 3270 6630
rect 3180 6530 3210 6560
rect 3240 6530 3270 6560
rect 3180 6465 3210 6495
rect 3240 6465 3270 6495
rect 3350 9605 3380 9635
rect 3350 9540 3380 9570
rect 3350 9470 3380 9500
rect 3350 9400 3380 9430
rect 3350 9330 3380 9360
rect 3350 9265 3380 9295
rect 3350 9205 3380 9235
rect 3350 9140 3380 9170
rect 3350 9070 3380 9100
rect 3350 9000 3380 9030
rect 3350 8930 3380 8960
rect 3350 8865 3380 8895
rect 3350 8805 3380 8835
rect 3350 8740 3380 8770
rect 3350 8670 3380 8700
rect 3350 8600 3380 8630
rect 3350 8530 3380 8560
rect 3350 8465 3380 8495
rect 3350 8405 3380 8435
rect 3350 8340 3380 8370
rect 3350 8270 3380 8300
rect 3350 8200 3380 8230
rect 3350 8130 3380 8160
rect 3350 8065 3380 8095
rect 3350 8005 3380 8035
rect 3350 7940 3380 7970
rect 3350 7870 3380 7900
rect 3350 7800 3380 7830
rect 3350 7730 3380 7760
rect 3350 7665 3380 7695
rect 3350 7605 3380 7635
rect 3350 7540 3380 7570
rect 3350 7470 3380 7500
rect 3350 7400 3380 7430
rect 3350 7330 3380 7360
rect 3350 7265 3380 7295
rect 3350 7205 3380 7235
rect 3350 7140 3380 7170
rect 3350 7070 3380 7100
rect 3350 7000 3380 7030
rect 3350 6930 3380 6960
rect 3350 6865 3380 6895
rect 3350 6805 3380 6835
rect 3350 6740 3380 6770
rect 3350 6670 3380 6700
rect 3350 6600 3380 6630
rect 3350 6530 3380 6560
rect 3350 6465 3380 6495
rect 3395 6400 3425 6430
rect 2995 6245 3025 6275
rect 3635 6345 3665 6375
rect 4310 6175 4340 6205
rect 4310 6135 4340 6165
rect 4310 6095 4340 6125
rect 4420 6175 4450 6205
rect 4420 6135 4450 6165
rect 4420 6095 4450 6125
rect 4530 6175 4560 6205
rect 4530 6135 4560 6165
rect 4530 6095 4560 6125
rect 5495 6400 5525 6430
rect 6150 6400 6180 6430
rect 5315 6345 5345 6375
rect 4855 6300 4885 6330
rect 4640 6175 4670 6205
rect 4640 6135 4670 6165
rect 4640 6095 4670 6125
rect 4855 5035 4885 5065
rect 4945 5035 4975 5065
rect 4945 4470 4975 4500
rect 5550 6245 5580 6275
rect 5495 2970 5525 3000
rect 6635 9605 6665 9635
rect 6635 9540 6665 9570
rect 6635 9470 6665 9500
rect 6635 9400 6665 9430
rect 6635 9330 6665 9360
rect 6635 9265 6665 9295
rect 6635 9205 6665 9235
rect 6635 9140 6665 9170
rect 6635 9070 6665 9100
rect 6635 9000 6665 9030
rect 6635 8930 6665 8960
rect 6635 8865 6665 8895
rect 6635 8805 6665 8835
rect 6635 8740 6665 8770
rect 6635 8670 6665 8700
rect 6635 8600 6665 8630
rect 6635 8530 6665 8560
rect 6635 8465 6665 8495
rect 6635 8405 6665 8435
rect 6635 8340 6665 8370
rect 6635 8270 6665 8300
rect 6635 8200 6665 8230
rect 6635 8130 6665 8160
rect 6635 8065 6665 8095
rect 6635 8005 6665 8035
rect 6635 7940 6665 7970
rect 6635 7870 6665 7900
rect 6635 7800 6665 7830
rect 6635 7730 6665 7760
rect 6635 7665 6665 7695
rect 6635 7605 6665 7635
rect 6635 7540 6665 7570
rect 6635 7470 6665 7500
rect 6635 7400 6665 7430
rect 6635 7330 6665 7360
rect 6635 7265 6665 7295
rect 6635 7205 6665 7235
rect 6635 7140 6665 7170
rect 6635 7070 6665 7100
rect 6635 7000 6665 7030
rect 6635 6930 6665 6960
rect 6635 6865 6665 6895
rect 6635 6805 6665 6835
rect 6635 6740 6665 6770
rect 6635 6670 6665 6700
rect 6635 6600 6665 6630
rect 6635 6530 6665 6560
rect 6635 6465 6665 6495
rect 7275 9605 7305 9635
rect 7275 9540 7305 9570
rect 7275 9470 7305 9500
rect 7275 9400 7305 9430
rect 7275 9330 7305 9360
rect 7275 9265 7305 9295
rect 7275 9205 7305 9235
rect 7275 9140 7305 9170
rect 7275 9070 7305 9100
rect 7275 9000 7305 9030
rect 7275 8930 7305 8960
rect 7275 8865 7305 8895
rect 7275 8805 7305 8835
rect 7275 8740 7305 8770
rect 7275 8670 7305 8700
rect 7275 8600 7305 8630
rect 7275 8530 7305 8560
rect 7275 8465 7305 8495
rect 7275 8405 7305 8435
rect 7275 8340 7305 8370
rect 7275 8270 7305 8300
rect 7275 8200 7305 8230
rect 7275 8130 7305 8160
rect 7275 8065 7305 8095
rect 7275 8005 7305 8035
rect 7275 7940 7305 7970
rect 7275 7870 7305 7900
rect 7275 7800 7305 7830
rect 7275 7730 7305 7760
rect 7275 7665 7305 7695
rect 7275 7605 7305 7635
rect 7275 7540 7305 7570
rect 7275 7470 7305 7500
rect 7275 7400 7305 7430
rect 7275 7330 7305 7360
rect 7275 7265 7305 7295
rect 7275 7205 7305 7235
rect 7275 7140 7305 7170
rect 7275 7070 7305 7100
rect 7275 7000 7305 7030
rect 7275 6930 7305 6960
rect 7275 6865 7305 6895
rect 7275 6805 7305 6835
rect 7275 6740 7305 6770
rect 7275 6670 7305 6700
rect 7275 6600 7305 6630
rect 7275 6530 7305 6560
rect 7275 6465 7305 6495
rect 6470 6400 6500 6430
rect 6900 6400 6930 6430
rect 5875 5055 5905 5085
rect 6225 5055 6255 5085
rect 5875 4550 5905 4580
rect 3395 2900 3425 2930
rect 5320 2915 5350 2945
rect 5550 2915 5580 2945
rect 6945 6345 6975 6375
rect 2050 1975 2080 2005
rect 2205 1975 2235 2005
rect 6745 1975 6775 2005
rect 6900 1975 6930 2005
rect 2005 1920 2035 1950
rect 2160 1920 2190 1950
rect 7975 9605 8005 9635
rect 7975 9540 8005 9570
rect 7975 9470 8005 9500
rect 7975 9400 8005 9430
rect 7975 9330 8005 9360
rect 7975 9265 8005 9295
rect 7975 9205 8005 9235
rect 7975 9140 8005 9170
rect 7975 9070 8005 9100
rect 7975 9000 8005 9030
rect 7975 8930 8005 8960
rect 7975 8865 8005 8895
rect 7975 8805 8005 8835
rect 7975 8740 8005 8770
rect 7975 8670 8005 8700
rect 7975 8600 8005 8630
rect 7975 8530 8005 8560
rect 7975 8465 8005 8495
rect 7975 8405 8005 8435
rect 7975 8340 8005 8370
rect 7975 8270 8005 8300
rect 7975 8200 8005 8230
rect 7975 8130 8005 8160
rect 7975 8065 8005 8095
rect 7975 8005 8005 8035
rect 7975 7940 8005 7970
rect 7975 7870 8005 7900
rect 7975 7800 8005 7830
rect 7975 7730 8005 7760
rect 7975 7665 8005 7695
rect 7975 7605 8005 7635
rect 7975 7540 8005 7570
rect 7975 7470 8005 7500
rect 7975 7400 8005 7430
rect 7975 7330 8005 7360
rect 7975 7265 8005 7295
rect 7975 7205 8005 7235
rect 7975 7140 8005 7170
rect 7975 7070 8005 7100
rect 7975 7000 8005 7030
rect 7975 6930 8005 6960
rect 7975 6865 8005 6895
rect 7975 6805 8005 6835
rect 7975 6740 8005 6770
rect 7975 6670 8005 6700
rect 7975 6600 8005 6630
rect 7975 6530 8005 6560
rect 7975 6465 8005 6495
rect 7585 6175 7615 6205
rect 7625 6175 7655 6205
rect 7665 6175 7695 6205
rect 8325 9605 8355 9635
rect 8325 9540 8355 9570
rect 8325 9470 8355 9500
rect 8325 9400 8355 9430
rect 8325 9330 8355 9360
rect 8325 9265 8355 9295
rect 8325 9205 8355 9235
rect 8325 9140 8355 9170
rect 8325 9070 8355 9100
rect 8325 9000 8355 9030
rect 8325 8930 8355 8960
rect 8325 8865 8355 8895
rect 8325 8805 8355 8835
rect 8325 8740 8355 8770
rect 8325 8670 8355 8700
rect 8325 8600 8355 8630
rect 8325 8530 8355 8560
rect 8325 8465 8355 8495
rect 8325 8405 8355 8435
rect 8325 8340 8355 8370
rect 8325 8270 8355 8300
rect 8325 8200 8355 8230
rect 8325 8130 8355 8160
rect 8325 8065 8355 8095
rect 8325 8005 8355 8035
rect 8325 7940 8355 7970
rect 8325 7870 8355 7900
rect 8325 7800 8355 7830
rect 8325 7730 8355 7760
rect 8325 7665 8355 7695
rect 8325 7605 8355 7635
rect 8325 7540 8355 7570
rect 8325 7470 8355 7500
rect 8325 7400 8355 7430
rect 8325 7330 8355 7360
rect 8325 7265 8355 7295
rect 8325 7205 8355 7235
rect 8325 7140 8355 7170
rect 8325 7070 8355 7100
rect 8325 7000 8355 7030
rect 8325 6930 8355 6960
rect 8325 6865 8355 6895
rect 8325 6805 8355 6835
rect 8325 6740 8355 6770
rect 8325 6670 8355 6700
rect 8325 6600 8355 6630
rect 8325 6530 8355 6560
rect 8325 6465 8355 6495
rect 8675 9605 8705 9635
rect 8675 9540 8705 9570
rect 8675 9470 8705 9500
rect 8675 9400 8705 9430
rect 8675 9330 8705 9360
rect 8675 9265 8705 9295
rect 8675 9205 8705 9235
rect 8675 9140 8705 9170
rect 8675 9070 8705 9100
rect 8675 9000 8705 9030
rect 8675 8930 8705 8960
rect 8675 8865 8705 8895
rect 8675 8805 8705 8835
rect 8675 8740 8705 8770
rect 8675 8670 8705 8700
rect 8675 8600 8705 8630
rect 8675 8530 8705 8560
rect 8675 8465 8705 8495
rect 8675 8405 8705 8435
rect 8675 8340 8705 8370
rect 8675 8270 8705 8300
rect 8675 8200 8705 8230
rect 8675 8130 8705 8160
rect 8675 8065 8705 8095
rect 8675 8005 8705 8035
rect 8675 7940 8705 7970
rect 8675 7870 8705 7900
rect 8675 7800 8705 7830
rect 8675 7730 8705 7760
rect 8675 7665 8705 7695
rect 8675 7605 8705 7635
rect 8675 7540 8705 7570
rect 8675 7470 8705 7500
rect 8675 7400 8705 7430
rect 8675 7330 8705 7360
rect 8675 7265 8705 7295
rect 8675 7205 8705 7235
rect 8675 7140 8705 7170
rect 8675 7070 8705 7100
rect 8675 7000 8705 7030
rect 8675 6930 8705 6960
rect 8675 6865 8705 6895
rect 8675 6805 8705 6835
rect 8675 6740 8705 6770
rect 8675 6670 8705 6700
rect 8675 6600 8705 6630
rect 8675 6530 8705 6560
rect 8675 6465 8705 6495
rect 9025 9605 9055 9635
rect 9025 9540 9055 9570
rect 9025 9470 9055 9500
rect 9025 9400 9055 9430
rect 9025 9330 9055 9360
rect 9025 9265 9055 9295
rect 9025 9205 9055 9235
rect 9025 9140 9055 9170
rect 9025 9070 9055 9100
rect 9025 9000 9055 9030
rect 9025 8930 9055 8960
rect 9025 8865 9055 8895
rect 9025 8805 9055 8835
rect 9025 8740 9055 8770
rect 9025 8670 9055 8700
rect 9025 8600 9055 8630
rect 9025 8530 9055 8560
rect 9025 8465 9055 8495
rect 9025 8405 9055 8435
rect 9025 8340 9055 8370
rect 9025 8270 9055 8300
rect 9025 8200 9055 8230
rect 9025 8130 9055 8160
rect 9025 8065 9055 8095
rect 9025 8005 9055 8035
rect 9025 7940 9055 7970
rect 9025 7870 9055 7900
rect 9025 7800 9055 7830
rect 9025 7730 9055 7760
rect 9025 7665 9055 7695
rect 9025 7605 9055 7635
rect 9025 7540 9055 7570
rect 9025 7470 9055 7500
rect 9025 7400 9055 7430
rect 9025 7330 9055 7360
rect 9025 7265 9055 7295
rect 9025 7205 9055 7235
rect 9025 7140 9055 7170
rect 9025 7070 9055 7100
rect 9025 7000 9055 7030
rect 9025 6930 9055 6960
rect 9025 6865 9055 6895
rect 9025 6805 9055 6835
rect 9025 6740 9055 6770
rect 9025 6670 9055 6700
rect 9025 6600 9055 6630
rect 9025 6530 9055 6560
rect 9025 6465 9055 6495
rect 7585 6135 7615 6165
rect 7625 6135 7655 6165
rect 7665 6135 7695 6165
rect 7585 6095 7615 6125
rect 7625 6095 7655 6125
rect 7665 6095 7695 6125
rect 6790 1920 6820 1950
rect 6945 1920 6975 1950
rect 1285 820 1315 850
rect 1325 820 1355 850
rect 1365 820 1395 850
rect 1285 780 1315 810
rect 1325 780 1355 810
rect 1365 780 1395 810
rect 1285 740 1315 770
rect 1325 740 1355 770
rect 1365 740 1395 770
rect 4420 820 4450 850
rect 4475 820 4505 850
rect 4530 820 4560 850
rect 4420 780 4450 810
rect 4475 780 4505 810
rect 4530 780 4560 810
rect 4420 740 4450 770
rect 4475 740 4505 770
rect 4530 740 4560 770
rect 7585 820 7615 850
rect 7625 820 7655 850
rect 7665 820 7695 850
rect 7585 780 7615 810
rect 7625 780 7655 810
rect 7665 780 7695 810
rect 7585 740 7615 770
rect 7625 740 7655 770
rect 7665 740 7695 770
rect -75 -1335 -45 -1305
rect -75 -1400 -45 -1370
rect -75 -1470 -45 -1440
rect -75 -1540 -45 -1510
rect -75 -1610 -45 -1580
rect -75 -1675 -45 -1645
rect -75 -1735 -45 -1705
rect -75 -1800 -45 -1770
rect -75 -1870 -45 -1840
rect -75 -1940 -45 -1910
rect -75 -2010 -45 -1980
rect -75 -2075 -45 -2045
rect -75 -2135 -45 -2105
rect -75 -2200 -45 -2170
rect -75 -2270 -45 -2240
rect -75 -2340 -45 -2310
rect -75 -2410 -45 -2380
rect -75 -2475 -45 -2445
rect -75 -2535 -45 -2505
rect -75 -2600 -45 -2570
rect -75 -2670 -45 -2640
rect -75 -2740 -45 -2710
rect -75 -2810 -45 -2780
rect -75 -2875 -45 -2845
rect -75 -2935 -45 -2905
rect -75 -3000 -45 -2970
rect -75 -3070 -45 -3040
rect -75 -3140 -45 -3110
rect -75 -3210 -45 -3180
rect -75 -3275 -45 -3245
rect -75 -3335 -45 -3305
rect -75 -3400 -45 -3370
rect -75 -3470 -45 -3440
rect -75 -3540 -45 -3510
rect -75 -3610 -45 -3580
rect -75 -3675 -45 -3645
rect -75 -3735 -45 -3705
rect -75 -3800 -45 -3770
rect -75 -3870 -45 -3840
rect -75 -3940 -45 -3910
rect -75 -4010 -45 -3980
rect -75 -4075 -45 -4045
rect -75 -4135 -45 -4105
rect -75 -4200 -45 -4170
rect -75 -4270 -45 -4240
rect -75 -4340 -45 -4310
rect -75 -4410 -45 -4380
rect -75 -4475 -45 -4445
rect 275 -1335 305 -1305
rect 275 -1400 305 -1370
rect 275 -1470 305 -1440
rect 275 -1540 305 -1510
rect 275 -1610 305 -1580
rect 275 -1675 305 -1645
rect 275 -1735 305 -1705
rect 275 -1800 305 -1770
rect 275 -1870 305 -1840
rect 275 -1940 305 -1910
rect 275 -2010 305 -1980
rect 275 -2075 305 -2045
rect 275 -2135 305 -2105
rect 275 -2200 305 -2170
rect 275 -2270 305 -2240
rect 275 -2340 305 -2310
rect 275 -2410 305 -2380
rect 275 -2475 305 -2445
rect 275 -2535 305 -2505
rect 275 -2600 305 -2570
rect 275 -2670 305 -2640
rect 275 -2740 305 -2710
rect 275 -2810 305 -2780
rect 275 -2875 305 -2845
rect 275 -2935 305 -2905
rect 275 -3000 305 -2970
rect 275 -3070 305 -3040
rect 275 -3140 305 -3110
rect 275 -3210 305 -3180
rect 275 -3275 305 -3245
rect 275 -3335 305 -3305
rect 275 -3400 305 -3370
rect 275 -3470 305 -3440
rect 275 -3540 305 -3510
rect 275 -3610 305 -3580
rect 275 -3675 305 -3645
rect 275 -3735 305 -3705
rect 275 -3800 305 -3770
rect 275 -3870 305 -3840
rect 275 -3940 305 -3910
rect 275 -4010 305 -3980
rect 275 -4075 305 -4045
rect 275 -4135 305 -4105
rect 275 -4200 305 -4170
rect 275 -4270 305 -4240
rect 275 -4340 305 -4310
rect 275 -4410 305 -4380
rect 275 -4475 305 -4445
rect 625 -1335 655 -1305
rect 625 -1400 655 -1370
rect 625 -1470 655 -1440
rect 625 -1540 655 -1510
rect 625 -1610 655 -1580
rect 625 -1675 655 -1645
rect 625 -1735 655 -1705
rect 625 -1800 655 -1770
rect 625 -1870 655 -1840
rect 625 -1940 655 -1910
rect 625 -2010 655 -1980
rect 625 -2075 655 -2045
rect 625 -2135 655 -2105
rect 625 -2200 655 -2170
rect 625 -2270 655 -2240
rect 625 -2340 655 -2310
rect 625 -2410 655 -2380
rect 625 -2475 655 -2445
rect 625 -2535 655 -2505
rect 625 -2600 655 -2570
rect 625 -2670 655 -2640
rect 625 -2740 655 -2710
rect 625 -2810 655 -2780
rect 625 -2875 655 -2845
rect 625 -2935 655 -2905
rect 625 -3000 655 -2970
rect 625 -3070 655 -3040
rect 625 -3140 655 -3110
rect 625 -3210 655 -3180
rect 625 -3275 655 -3245
rect 625 -3335 655 -3305
rect 625 -3400 655 -3370
rect 625 -3470 655 -3440
rect 625 -3540 655 -3510
rect 625 -3610 655 -3580
rect 625 -3675 655 -3645
rect 625 -3735 655 -3705
rect 625 -3800 655 -3770
rect 625 -3870 655 -3840
rect 625 -3940 655 -3910
rect 625 -4010 655 -3980
rect 625 -4075 655 -4045
rect 625 -4135 655 -4105
rect 625 -4200 655 -4170
rect 625 -4270 655 -4240
rect 625 -4340 655 -4310
rect 625 -4410 655 -4380
rect 625 -4475 655 -4445
rect 975 -1335 1005 -1305
rect 975 -1400 1005 -1370
rect 975 -1470 1005 -1440
rect 975 -1540 1005 -1510
rect 975 -1610 1005 -1580
rect 975 -1675 1005 -1645
rect 975 -1735 1005 -1705
rect 975 -1800 1005 -1770
rect 975 -1870 1005 -1840
rect 975 -1940 1005 -1910
rect 975 -2010 1005 -1980
rect 975 -2075 1005 -2045
rect 975 -2135 1005 -2105
rect 975 -2200 1005 -2170
rect 975 -2270 1005 -2240
rect 975 -2340 1005 -2310
rect 975 -2410 1005 -2380
rect 975 -2475 1005 -2445
rect 975 -2535 1005 -2505
rect 975 -2600 1005 -2570
rect 975 -2670 1005 -2640
rect 975 -2740 1005 -2710
rect 975 -2810 1005 -2780
rect 975 -2875 1005 -2845
rect 975 -2935 1005 -2905
rect 975 -3000 1005 -2970
rect 975 -3070 1005 -3040
rect 975 -3140 1005 -3110
rect 975 -3210 1005 -3180
rect 975 -3275 1005 -3245
rect 975 -3335 1005 -3305
rect 975 -3400 1005 -3370
rect 975 -3470 1005 -3440
rect 975 -3540 1005 -3510
rect 975 -3610 1005 -3580
rect 975 -3675 1005 -3645
rect 975 -3735 1005 -3705
rect 975 -3800 1005 -3770
rect 975 -3870 1005 -3840
rect 975 -3940 1005 -3910
rect 975 -4010 1005 -3980
rect 975 -4075 1005 -4045
rect 975 -4135 1005 -4105
rect 975 -4200 1005 -4170
rect 975 -4270 1005 -4240
rect 975 -4340 1005 -4310
rect 975 -4410 1005 -4380
rect 975 -4475 1005 -4445
rect 1325 -1335 1355 -1305
rect 1325 -1400 1355 -1370
rect 1325 -1470 1355 -1440
rect 1325 -1540 1355 -1510
rect 1325 -1610 1355 -1580
rect 1325 -1675 1355 -1645
rect 1325 -1735 1355 -1705
rect 1325 -1800 1355 -1770
rect 1325 -1870 1355 -1840
rect 1325 -1940 1355 -1910
rect 1325 -2010 1355 -1980
rect 1325 -2075 1355 -2045
rect 1325 -2135 1355 -2105
rect 1325 -2200 1355 -2170
rect 1325 -2270 1355 -2240
rect 1325 -2340 1355 -2310
rect 1325 -2410 1355 -2380
rect 1325 -2475 1355 -2445
rect 1325 -2535 1355 -2505
rect 1325 -2600 1355 -2570
rect 1325 -2670 1355 -2640
rect 1325 -2740 1355 -2710
rect 1325 -2810 1355 -2780
rect 1325 -2875 1355 -2845
rect 1325 -2935 1355 -2905
rect 1325 -3000 1355 -2970
rect 1325 -3070 1355 -3040
rect 1325 -3140 1355 -3110
rect 1325 -3210 1355 -3180
rect 1325 -3275 1355 -3245
rect 1325 -3335 1355 -3305
rect 1325 -3400 1355 -3370
rect 1325 -3470 1355 -3440
rect 1325 -3540 1355 -3510
rect 1325 -3610 1355 -3580
rect 1325 -3675 1355 -3645
rect 1325 -3735 1355 -3705
rect 1325 -3800 1355 -3770
rect 1325 -3870 1355 -3840
rect 1325 -3940 1355 -3910
rect 1325 -4010 1355 -3980
rect 1325 -4075 1355 -4045
rect 1325 -4135 1355 -4105
rect 1325 -4200 1355 -4170
rect 1325 -4270 1355 -4240
rect 1325 -4340 1355 -4310
rect 1325 -4410 1355 -4380
rect 1325 -4475 1355 -4445
rect 1675 -1335 1705 -1305
rect 1675 -1400 1705 -1370
rect 1675 -1470 1705 -1440
rect 1675 -1540 1705 -1510
rect 1675 -1610 1705 -1580
rect 1675 -1675 1705 -1645
rect 1675 -1735 1705 -1705
rect 1675 -1800 1705 -1770
rect 1675 -1870 1705 -1840
rect 1675 -1940 1705 -1910
rect 1675 -2010 1705 -1980
rect 1675 -2075 1705 -2045
rect 1675 -2135 1705 -2105
rect 1675 -2200 1705 -2170
rect 1675 -2270 1705 -2240
rect 1675 -2340 1705 -2310
rect 1675 -2410 1705 -2380
rect 1675 -2475 1705 -2445
rect 1675 -2535 1705 -2505
rect 1675 -2600 1705 -2570
rect 1675 -2670 1705 -2640
rect 1675 -2740 1705 -2710
rect 1675 -2810 1705 -2780
rect 1675 -2875 1705 -2845
rect 1675 -2935 1705 -2905
rect 1675 -3000 1705 -2970
rect 1675 -3070 1705 -3040
rect 1675 -3140 1705 -3110
rect 1675 -3210 1705 -3180
rect 1675 -3275 1705 -3245
rect 1675 -3335 1705 -3305
rect 1675 -3400 1705 -3370
rect 1675 -3470 1705 -3440
rect 1675 -3540 1705 -3510
rect 1675 -3610 1705 -3580
rect 1675 -3675 1705 -3645
rect 1675 -3735 1705 -3705
rect 1675 -3800 1705 -3770
rect 1675 -3870 1705 -3840
rect 1675 -3940 1705 -3910
rect 1675 -4010 1705 -3980
rect 1675 -4075 1705 -4045
rect 1675 -4135 1705 -4105
rect 1675 -4200 1705 -4170
rect 1675 -4270 1705 -4240
rect 1675 -4340 1705 -4310
rect 1675 -4410 1705 -4380
rect 1675 -4475 1705 -4445
rect 2025 -1335 2055 -1305
rect 2025 -1400 2055 -1370
rect 2025 -1470 2055 -1440
rect 2025 -1540 2055 -1510
rect 2025 -1610 2055 -1580
rect 2025 -1675 2055 -1645
rect 2025 -1735 2055 -1705
rect 2025 -1800 2055 -1770
rect 2025 -1870 2055 -1840
rect 2025 -1940 2055 -1910
rect 2025 -2010 2055 -1980
rect 2025 -2075 2055 -2045
rect 2025 -2135 2055 -2105
rect 2025 -2200 2055 -2170
rect 2025 -2270 2055 -2240
rect 2025 -2340 2055 -2310
rect 2025 -2410 2055 -2380
rect 2025 -2475 2055 -2445
rect 2025 -2535 2055 -2505
rect 2025 -2600 2055 -2570
rect 2025 -2670 2055 -2640
rect 2025 -2740 2055 -2710
rect 2025 -2810 2055 -2780
rect 2025 -2875 2055 -2845
rect 2025 -2935 2055 -2905
rect 2025 -3000 2055 -2970
rect 2025 -3070 2055 -3040
rect 2025 -3140 2055 -3110
rect 2025 -3210 2055 -3180
rect 2025 -3275 2055 -3245
rect 2025 -3335 2055 -3305
rect 2025 -3400 2055 -3370
rect 2025 -3470 2055 -3440
rect 2025 -3540 2055 -3510
rect 2025 -3610 2055 -3580
rect 2025 -3675 2055 -3645
rect 2025 -3735 2055 -3705
rect 2025 -3800 2055 -3770
rect 2025 -3870 2055 -3840
rect 2025 -3940 2055 -3910
rect 2025 -4010 2055 -3980
rect 2025 -4075 2055 -4045
rect 2025 -4135 2055 -4105
rect 2025 -4200 2055 -4170
rect 2025 -4270 2055 -4240
rect 2025 -4340 2055 -4310
rect 2025 -4410 2055 -4380
rect 2025 -4475 2055 -4445
rect 2375 -1335 2405 -1305
rect 2375 -1400 2405 -1370
rect 2375 -1470 2405 -1440
rect 2375 -1540 2405 -1510
rect 2375 -1610 2405 -1580
rect 2375 -1675 2405 -1645
rect 2375 -1735 2405 -1705
rect 2375 -1800 2405 -1770
rect 2375 -1870 2405 -1840
rect 2375 -1940 2405 -1910
rect 2375 -2010 2405 -1980
rect 2375 -2075 2405 -2045
rect 2375 -2135 2405 -2105
rect 2375 -2200 2405 -2170
rect 2375 -2270 2405 -2240
rect 2375 -2340 2405 -2310
rect 2375 -2410 2405 -2380
rect 2375 -2475 2405 -2445
rect 2375 -2535 2405 -2505
rect 2375 -2600 2405 -2570
rect 2375 -2670 2405 -2640
rect 2375 -2740 2405 -2710
rect 2375 -2810 2405 -2780
rect 2375 -2875 2405 -2845
rect 2375 -2935 2405 -2905
rect 2375 -3000 2405 -2970
rect 2375 -3070 2405 -3040
rect 2375 -3140 2405 -3110
rect 2375 -3210 2405 -3180
rect 2375 -3275 2405 -3245
rect 2375 -3335 2405 -3305
rect 2375 -3400 2405 -3370
rect 2375 -3470 2405 -3440
rect 2375 -3540 2405 -3510
rect 2375 -3610 2405 -3580
rect 2375 -3675 2405 -3645
rect 2375 -3735 2405 -3705
rect 2375 -3800 2405 -3770
rect 2375 -3870 2405 -3840
rect 2375 -3940 2405 -3910
rect 2375 -4010 2405 -3980
rect 2375 -4075 2405 -4045
rect 2375 -4135 2405 -4105
rect 2375 -4200 2405 -4170
rect 2375 -4270 2405 -4240
rect 2375 -4340 2405 -4310
rect 2375 -4410 2405 -4380
rect 2375 -4475 2405 -4445
rect 2725 -1335 2755 -1305
rect 2725 -1400 2755 -1370
rect 2725 -1470 2755 -1440
rect 2725 -1540 2755 -1510
rect 2725 -1610 2755 -1580
rect 2725 -1675 2755 -1645
rect 2725 -1735 2755 -1705
rect 2725 -1800 2755 -1770
rect 2725 -1870 2755 -1840
rect 2725 -1940 2755 -1910
rect 2725 -2010 2755 -1980
rect 2725 -2075 2755 -2045
rect 2725 -2135 2755 -2105
rect 2725 -2200 2755 -2170
rect 2725 -2270 2755 -2240
rect 2725 -2340 2755 -2310
rect 2725 -2410 2755 -2380
rect 2725 -2475 2755 -2445
rect 2725 -2535 2755 -2505
rect 2725 -2600 2755 -2570
rect 2725 -2670 2755 -2640
rect 2725 -2740 2755 -2710
rect 2725 -2810 2755 -2780
rect 2725 -2875 2755 -2845
rect 2725 -2935 2755 -2905
rect 2725 -3000 2755 -2970
rect 2725 -3070 2755 -3040
rect 2725 -3140 2755 -3110
rect 2725 -3210 2755 -3180
rect 2725 -3275 2755 -3245
rect 2725 -3335 2755 -3305
rect 2725 -3400 2755 -3370
rect 2725 -3470 2755 -3440
rect 2725 -3540 2755 -3510
rect 2725 -3610 2755 -3580
rect 2725 -3675 2755 -3645
rect 2725 -3735 2755 -3705
rect 2725 -3800 2755 -3770
rect 2725 -3870 2755 -3840
rect 2725 -3940 2755 -3910
rect 2725 -4010 2755 -3980
rect 2725 -4075 2755 -4045
rect 2725 -4135 2755 -4105
rect 2725 -4200 2755 -4170
rect 2725 -4270 2755 -4240
rect 2725 -4340 2755 -4310
rect 2725 -4410 2755 -4380
rect 2725 -4475 2755 -4445
rect 3075 -1335 3105 -1305
rect 3075 -1400 3105 -1370
rect 3075 -1470 3105 -1440
rect 3075 -1540 3105 -1510
rect 3075 -1610 3105 -1580
rect 3075 -1675 3105 -1645
rect 3075 -1735 3105 -1705
rect 3075 -1800 3105 -1770
rect 3075 -1870 3105 -1840
rect 3075 -1940 3105 -1910
rect 3075 -2010 3105 -1980
rect 3075 -2075 3105 -2045
rect 3075 -2135 3105 -2105
rect 3075 -2200 3105 -2170
rect 3075 -2270 3105 -2240
rect 3075 -2340 3105 -2310
rect 3075 -2410 3105 -2380
rect 3075 -2475 3105 -2445
rect 3075 -2535 3105 -2505
rect 3075 -2600 3105 -2570
rect 3075 -2670 3105 -2640
rect 3075 -2740 3105 -2710
rect 3075 -2810 3105 -2780
rect 3075 -2875 3105 -2845
rect 3075 -2935 3105 -2905
rect 3075 -3000 3105 -2970
rect 3075 -3070 3105 -3040
rect 3075 -3140 3105 -3110
rect 3075 -3210 3105 -3180
rect 3075 -3275 3105 -3245
rect 3075 -3335 3105 -3305
rect 3075 -3400 3105 -3370
rect 3075 -3470 3105 -3440
rect 3075 -3540 3105 -3510
rect 3075 -3610 3105 -3580
rect 3075 -3675 3105 -3645
rect 3075 -3735 3105 -3705
rect 3075 -3800 3105 -3770
rect 3075 -3870 3105 -3840
rect 3075 -3940 3105 -3910
rect 3075 -4010 3105 -3980
rect 3075 -4075 3105 -4045
rect 3075 -4135 3105 -4105
rect 3075 -4200 3105 -4170
rect 3075 -4270 3105 -4240
rect 3075 -4340 3105 -4310
rect 3075 -4410 3105 -4380
rect 3075 -4475 3105 -4445
rect 3425 -1335 3455 -1305
rect 3425 -1400 3455 -1370
rect 3425 -1470 3455 -1440
rect 3425 -1540 3455 -1510
rect 3425 -1610 3455 -1580
rect 3425 -1675 3455 -1645
rect 3425 -1735 3455 -1705
rect 3425 -1800 3455 -1770
rect 3425 -1870 3455 -1840
rect 3425 -1940 3455 -1910
rect 3425 -2010 3455 -1980
rect 3425 -2075 3455 -2045
rect 3425 -2135 3455 -2105
rect 3425 -2200 3455 -2170
rect 3425 -2270 3455 -2240
rect 3425 -2340 3455 -2310
rect 3425 -2410 3455 -2380
rect 3425 -2475 3455 -2445
rect 3425 -2535 3455 -2505
rect 3425 -2600 3455 -2570
rect 3425 -2670 3455 -2640
rect 3425 -2740 3455 -2710
rect 3425 -2810 3455 -2780
rect 3425 -2875 3455 -2845
rect 3425 -2935 3455 -2905
rect 3425 -3000 3455 -2970
rect 3425 -3070 3455 -3040
rect 3425 -3140 3455 -3110
rect 3425 -3210 3455 -3180
rect 3425 -3275 3455 -3245
rect 3425 -3335 3455 -3305
rect 3425 -3400 3455 -3370
rect 3425 -3470 3455 -3440
rect 3425 -3540 3455 -3510
rect 3425 -3610 3455 -3580
rect 3425 -3675 3455 -3645
rect 3425 -3735 3455 -3705
rect 3425 -3800 3455 -3770
rect 3425 -3870 3455 -3840
rect 3425 -3940 3455 -3910
rect 3425 -4010 3455 -3980
rect 3425 -4075 3455 -4045
rect 3425 -4135 3455 -4105
rect 3425 -4200 3455 -4170
rect 3425 -4270 3455 -4240
rect 3425 -4340 3455 -4310
rect 3425 -4410 3455 -4380
rect 3425 -4475 3455 -4445
rect 3775 -1335 3805 -1305
rect 3775 -1400 3805 -1370
rect 3775 -1470 3805 -1440
rect 3775 -1540 3805 -1510
rect 3775 -1610 3805 -1580
rect 3775 -1675 3805 -1645
rect 3775 -1735 3805 -1705
rect 3775 -1800 3805 -1770
rect 3775 -1870 3805 -1840
rect 3775 -1940 3805 -1910
rect 3775 -2010 3805 -1980
rect 3775 -2075 3805 -2045
rect 3775 -2135 3805 -2105
rect 3775 -2200 3805 -2170
rect 3775 -2270 3805 -2240
rect 3775 -2340 3805 -2310
rect 3775 -2410 3805 -2380
rect 3775 -2475 3805 -2445
rect 3775 -2535 3805 -2505
rect 3775 -2600 3805 -2570
rect 3775 -2670 3805 -2640
rect 3775 -2740 3805 -2710
rect 3775 -2810 3805 -2780
rect 3775 -2875 3805 -2845
rect 3775 -2935 3805 -2905
rect 3775 -3000 3805 -2970
rect 3775 -3070 3805 -3040
rect 3775 -3140 3805 -3110
rect 3775 -3210 3805 -3180
rect 3775 -3275 3805 -3245
rect 3775 -3335 3805 -3305
rect 3775 -3400 3805 -3370
rect 3775 -3470 3805 -3440
rect 3775 -3540 3805 -3510
rect 3775 -3610 3805 -3580
rect 3775 -3675 3805 -3645
rect 3775 -3735 3805 -3705
rect 3775 -3800 3805 -3770
rect 3775 -3870 3805 -3840
rect 3775 -3940 3805 -3910
rect 3775 -4010 3805 -3980
rect 3775 -4075 3805 -4045
rect 3775 -4135 3805 -4105
rect 3775 -4200 3805 -4170
rect 3775 -4270 3805 -4240
rect 3775 -4340 3805 -4310
rect 3775 -4410 3805 -4380
rect 3775 -4475 3805 -4445
rect 4125 -1335 4155 -1305
rect 4125 -1400 4155 -1370
rect 4125 -1470 4155 -1440
rect 4125 -1540 4155 -1510
rect 4125 -1610 4155 -1580
rect 4125 -1675 4155 -1645
rect 4125 -1735 4155 -1705
rect 4125 -1800 4155 -1770
rect 4125 -1870 4155 -1840
rect 4125 -1940 4155 -1910
rect 4125 -2010 4155 -1980
rect 4125 -2075 4155 -2045
rect 4125 -2135 4155 -2105
rect 4125 -2200 4155 -2170
rect 4125 -2270 4155 -2240
rect 4125 -2340 4155 -2310
rect 4125 -2410 4155 -2380
rect 4125 -2475 4155 -2445
rect 4125 -2535 4155 -2505
rect 4125 -2600 4155 -2570
rect 4125 -2670 4155 -2640
rect 4125 -2740 4155 -2710
rect 4125 -2810 4155 -2780
rect 4125 -2875 4155 -2845
rect 4125 -2935 4155 -2905
rect 4125 -3000 4155 -2970
rect 4125 -3070 4155 -3040
rect 4125 -3140 4155 -3110
rect 4125 -3210 4155 -3180
rect 4125 -3275 4155 -3245
rect 4125 -3335 4155 -3305
rect 4125 -3400 4155 -3370
rect 4125 -3470 4155 -3440
rect 4125 -3540 4155 -3510
rect 4125 -3610 4155 -3580
rect 4125 -3675 4155 -3645
rect 4125 -3735 4155 -3705
rect 4125 -3800 4155 -3770
rect 4125 -3870 4155 -3840
rect 4125 -3940 4155 -3910
rect 4125 -4010 4155 -3980
rect 4125 -4075 4155 -4045
rect 4125 -4135 4155 -4105
rect 4125 -4200 4155 -4170
rect 4125 -4270 4155 -4240
rect 4125 -4340 4155 -4310
rect 4125 -4410 4155 -4380
rect 4125 -4475 4155 -4445
rect 4475 -1335 4505 -1305
rect 4475 -1400 4505 -1370
rect 4475 -1470 4505 -1440
rect 4475 -1540 4505 -1510
rect 4475 -1610 4505 -1580
rect 4475 -1675 4505 -1645
rect 4475 -1735 4505 -1705
rect 4475 -1800 4505 -1770
rect 4475 -1870 4505 -1840
rect 4475 -1940 4505 -1910
rect 4475 -2010 4505 -1980
rect 4475 -2075 4505 -2045
rect 4475 -2135 4505 -2105
rect 4475 -2200 4505 -2170
rect 4475 -2270 4505 -2240
rect 4475 -2340 4505 -2310
rect 4475 -2410 4505 -2380
rect 4475 -2475 4505 -2445
rect 4475 -2535 4505 -2505
rect 4475 -2600 4505 -2570
rect 4475 -2670 4505 -2640
rect 4475 -2740 4505 -2710
rect 4475 -2810 4505 -2780
rect 4475 -2875 4505 -2845
rect 4475 -2935 4505 -2905
rect 4475 -3000 4505 -2970
rect 4475 -3070 4505 -3040
rect 4475 -3140 4505 -3110
rect 4475 -3210 4505 -3180
rect 4475 -3275 4505 -3245
rect 4475 -3335 4505 -3305
rect 4475 -3400 4505 -3370
rect 4475 -3470 4505 -3440
rect 4475 -3540 4505 -3510
rect 4475 -3610 4505 -3580
rect 4475 -3675 4505 -3645
rect 4475 -3735 4505 -3705
rect 4475 -3800 4505 -3770
rect 4475 -3870 4505 -3840
rect 4475 -3940 4505 -3910
rect 4475 -4010 4505 -3980
rect 4475 -4075 4505 -4045
rect 4475 -4135 4505 -4105
rect 4475 -4200 4505 -4170
rect 4475 -4270 4505 -4240
rect 4475 -4340 4505 -4310
rect 4475 -4410 4505 -4380
rect 4475 -4475 4505 -4445
rect 4825 -1335 4855 -1305
rect 4825 -1400 4855 -1370
rect 4825 -1470 4855 -1440
rect 4825 -1540 4855 -1510
rect 4825 -1610 4855 -1580
rect 4825 -1675 4855 -1645
rect 4825 -1735 4855 -1705
rect 4825 -1800 4855 -1770
rect 4825 -1870 4855 -1840
rect 4825 -1940 4855 -1910
rect 4825 -2010 4855 -1980
rect 4825 -2075 4855 -2045
rect 4825 -2135 4855 -2105
rect 4825 -2200 4855 -2170
rect 4825 -2270 4855 -2240
rect 4825 -2340 4855 -2310
rect 4825 -2410 4855 -2380
rect 4825 -2475 4855 -2445
rect 4825 -2535 4855 -2505
rect 4825 -2600 4855 -2570
rect 4825 -2670 4855 -2640
rect 4825 -2740 4855 -2710
rect 4825 -2810 4855 -2780
rect 4825 -2875 4855 -2845
rect 4825 -2935 4855 -2905
rect 4825 -3000 4855 -2970
rect 4825 -3070 4855 -3040
rect 4825 -3140 4855 -3110
rect 4825 -3210 4855 -3180
rect 4825 -3275 4855 -3245
rect 4825 -3335 4855 -3305
rect 4825 -3400 4855 -3370
rect 4825 -3470 4855 -3440
rect 4825 -3540 4855 -3510
rect 4825 -3610 4855 -3580
rect 4825 -3675 4855 -3645
rect 4825 -3735 4855 -3705
rect 4825 -3800 4855 -3770
rect 4825 -3870 4855 -3840
rect 4825 -3940 4855 -3910
rect 4825 -4010 4855 -3980
rect 4825 -4075 4855 -4045
rect 4825 -4135 4855 -4105
rect 4825 -4200 4855 -4170
rect 4825 -4270 4855 -4240
rect 4825 -4340 4855 -4310
rect 4825 -4410 4855 -4380
rect 4825 -4475 4855 -4445
rect 5175 -1335 5205 -1305
rect 5175 -1400 5205 -1370
rect 5175 -1470 5205 -1440
rect 5175 -1540 5205 -1510
rect 5175 -1610 5205 -1580
rect 5175 -1675 5205 -1645
rect 5175 -1735 5205 -1705
rect 5175 -1800 5205 -1770
rect 5175 -1870 5205 -1840
rect 5175 -1940 5205 -1910
rect 5175 -2010 5205 -1980
rect 5175 -2075 5205 -2045
rect 5175 -2135 5205 -2105
rect 5175 -2200 5205 -2170
rect 5175 -2270 5205 -2240
rect 5175 -2340 5205 -2310
rect 5175 -2410 5205 -2380
rect 5175 -2475 5205 -2445
rect 5175 -2535 5205 -2505
rect 5175 -2600 5205 -2570
rect 5175 -2670 5205 -2640
rect 5175 -2740 5205 -2710
rect 5175 -2810 5205 -2780
rect 5175 -2875 5205 -2845
rect 5175 -2935 5205 -2905
rect 5175 -3000 5205 -2970
rect 5175 -3070 5205 -3040
rect 5175 -3140 5205 -3110
rect 5175 -3210 5205 -3180
rect 5175 -3275 5205 -3245
rect 5175 -3335 5205 -3305
rect 5175 -3400 5205 -3370
rect 5175 -3470 5205 -3440
rect 5175 -3540 5205 -3510
rect 5175 -3610 5205 -3580
rect 5175 -3675 5205 -3645
rect 5175 -3735 5205 -3705
rect 5175 -3800 5205 -3770
rect 5175 -3870 5205 -3840
rect 5175 -3940 5205 -3910
rect 5175 -4010 5205 -3980
rect 5175 -4075 5205 -4045
rect 5175 -4135 5205 -4105
rect 5175 -4200 5205 -4170
rect 5175 -4270 5205 -4240
rect 5175 -4340 5205 -4310
rect 5175 -4410 5205 -4380
rect 5175 -4475 5205 -4445
rect 5525 -1335 5555 -1305
rect 5525 -1400 5555 -1370
rect 5525 -1470 5555 -1440
rect 5525 -1540 5555 -1510
rect 5525 -1610 5555 -1580
rect 5525 -1675 5555 -1645
rect 5525 -1735 5555 -1705
rect 5525 -1800 5555 -1770
rect 5525 -1870 5555 -1840
rect 5525 -1940 5555 -1910
rect 5525 -2010 5555 -1980
rect 5525 -2075 5555 -2045
rect 5525 -2135 5555 -2105
rect 5525 -2200 5555 -2170
rect 5525 -2270 5555 -2240
rect 5525 -2340 5555 -2310
rect 5525 -2410 5555 -2380
rect 5525 -2475 5555 -2445
rect 5525 -2535 5555 -2505
rect 5525 -2600 5555 -2570
rect 5525 -2670 5555 -2640
rect 5525 -2740 5555 -2710
rect 5525 -2810 5555 -2780
rect 5525 -2875 5555 -2845
rect 5525 -2935 5555 -2905
rect 5525 -3000 5555 -2970
rect 5525 -3070 5555 -3040
rect 5525 -3140 5555 -3110
rect 5525 -3210 5555 -3180
rect 5525 -3275 5555 -3245
rect 5525 -3335 5555 -3305
rect 5525 -3400 5555 -3370
rect 5525 -3470 5555 -3440
rect 5525 -3540 5555 -3510
rect 5525 -3610 5555 -3580
rect 5525 -3675 5555 -3645
rect 5525 -3735 5555 -3705
rect 5525 -3800 5555 -3770
rect 5525 -3870 5555 -3840
rect 5525 -3940 5555 -3910
rect 5525 -4010 5555 -3980
rect 5525 -4075 5555 -4045
rect 5525 -4135 5555 -4105
rect 5525 -4200 5555 -4170
rect 5525 -4270 5555 -4240
rect 5525 -4340 5555 -4310
rect 5525 -4410 5555 -4380
rect 5525 -4475 5555 -4445
rect 5875 -1335 5905 -1305
rect 5875 -1400 5905 -1370
rect 5875 -1470 5905 -1440
rect 5875 -1540 5905 -1510
rect 5875 -1610 5905 -1580
rect 5875 -1675 5905 -1645
rect 5875 -1735 5905 -1705
rect 5875 -1800 5905 -1770
rect 5875 -1870 5905 -1840
rect 5875 -1940 5905 -1910
rect 5875 -2010 5905 -1980
rect 5875 -2075 5905 -2045
rect 5875 -2135 5905 -2105
rect 5875 -2200 5905 -2170
rect 5875 -2270 5905 -2240
rect 5875 -2340 5905 -2310
rect 5875 -2410 5905 -2380
rect 5875 -2475 5905 -2445
rect 5875 -2535 5905 -2505
rect 5875 -2600 5905 -2570
rect 5875 -2670 5905 -2640
rect 5875 -2740 5905 -2710
rect 5875 -2810 5905 -2780
rect 5875 -2875 5905 -2845
rect 5875 -2935 5905 -2905
rect 5875 -3000 5905 -2970
rect 5875 -3070 5905 -3040
rect 5875 -3140 5905 -3110
rect 5875 -3210 5905 -3180
rect 5875 -3275 5905 -3245
rect 5875 -3335 5905 -3305
rect 5875 -3400 5905 -3370
rect 5875 -3470 5905 -3440
rect 5875 -3540 5905 -3510
rect 5875 -3610 5905 -3580
rect 5875 -3675 5905 -3645
rect 5875 -3735 5905 -3705
rect 5875 -3800 5905 -3770
rect 5875 -3870 5905 -3840
rect 5875 -3940 5905 -3910
rect 5875 -4010 5905 -3980
rect 5875 -4075 5905 -4045
rect 5875 -4135 5905 -4105
rect 5875 -4200 5905 -4170
rect 5875 -4270 5905 -4240
rect 5875 -4340 5905 -4310
rect 5875 -4410 5905 -4380
rect 5875 -4475 5905 -4445
rect 6225 -1335 6255 -1305
rect 6225 -1400 6255 -1370
rect 6225 -1470 6255 -1440
rect 6225 -1540 6255 -1510
rect 6225 -1610 6255 -1580
rect 6225 -1675 6255 -1645
rect 6225 -1735 6255 -1705
rect 6225 -1800 6255 -1770
rect 6225 -1870 6255 -1840
rect 6225 -1940 6255 -1910
rect 6225 -2010 6255 -1980
rect 6225 -2075 6255 -2045
rect 6225 -2135 6255 -2105
rect 6225 -2200 6255 -2170
rect 6225 -2270 6255 -2240
rect 6225 -2340 6255 -2310
rect 6225 -2410 6255 -2380
rect 6225 -2475 6255 -2445
rect 6225 -2535 6255 -2505
rect 6225 -2600 6255 -2570
rect 6225 -2670 6255 -2640
rect 6225 -2740 6255 -2710
rect 6225 -2810 6255 -2780
rect 6225 -2875 6255 -2845
rect 6225 -2935 6255 -2905
rect 6225 -3000 6255 -2970
rect 6225 -3070 6255 -3040
rect 6225 -3140 6255 -3110
rect 6225 -3210 6255 -3180
rect 6225 -3275 6255 -3245
rect 6225 -3335 6255 -3305
rect 6225 -3400 6255 -3370
rect 6225 -3470 6255 -3440
rect 6225 -3540 6255 -3510
rect 6225 -3610 6255 -3580
rect 6225 -3675 6255 -3645
rect 6225 -3735 6255 -3705
rect 6225 -3800 6255 -3770
rect 6225 -3870 6255 -3840
rect 6225 -3940 6255 -3910
rect 6225 -4010 6255 -3980
rect 6225 -4075 6255 -4045
rect 6225 -4135 6255 -4105
rect 6225 -4200 6255 -4170
rect 6225 -4270 6255 -4240
rect 6225 -4340 6255 -4310
rect 6225 -4410 6255 -4380
rect 6225 -4475 6255 -4445
rect 6575 -1335 6605 -1305
rect 6575 -1400 6605 -1370
rect 6575 -1470 6605 -1440
rect 6575 -1540 6605 -1510
rect 6575 -1610 6605 -1580
rect 6575 -1675 6605 -1645
rect 6575 -1735 6605 -1705
rect 6575 -1800 6605 -1770
rect 6575 -1870 6605 -1840
rect 6575 -1940 6605 -1910
rect 6575 -2010 6605 -1980
rect 6575 -2075 6605 -2045
rect 6575 -2135 6605 -2105
rect 6575 -2200 6605 -2170
rect 6575 -2270 6605 -2240
rect 6575 -2340 6605 -2310
rect 6575 -2410 6605 -2380
rect 6575 -2475 6605 -2445
rect 6575 -2535 6605 -2505
rect 6575 -2600 6605 -2570
rect 6575 -2670 6605 -2640
rect 6575 -2740 6605 -2710
rect 6575 -2810 6605 -2780
rect 6575 -2875 6605 -2845
rect 6575 -2935 6605 -2905
rect 6575 -3000 6605 -2970
rect 6575 -3070 6605 -3040
rect 6575 -3140 6605 -3110
rect 6575 -3210 6605 -3180
rect 6575 -3275 6605 -3245
rect 6575 -3335 6605 -3305
rect 6575 -3400 6605 -3370
rect 6575 -3470 6605 -3440
rect 6575 -3540 6605 -3510
rect 6575 -3610 6605 -3580
rect 6575 -3675 6605 -3645
rect 6575 -3735 6605 -3705
rect 6575 -3800 6605 -3770
rect 6575 -3870 6605 -3840
rect 6575 -3940 6605 -3910
rect 6575 -4010 6605 -3980
rect 6575 -4075 6605 -4045
rect 6575 -4135 6605 -4105
rect 6575 -4200 6605 -4170
rect 6575 -4270 6605 -4240
rect 6575 -4340 6605 -4310
rect 6575 -4410 6605 -4380
rect 6575 -4475 6605 -4445
rect 6925 -1335 6955 -1305
rect 6925 -1400 6955 -1370
rect 6925 -1470 6955 -1440
rect 6925 -1540 6955 -1510
rect 6925 -1610 6955 -1580
rect 6925 -1675 6955 -1645
rect 6925 -1735 6955 -1705
rect 6925 -1800 6955 -1770
rect 6925 -1870 6955 -1840
rect 6925 -1940 6955 -1910
rect 6925 -2010 6955 -1980
rect 6925 -2075 6955 -2045
rect 6925 -2135 6955 -2105
rect 6925 -2200 6955 -2170
rect 6925 -2270 6955 -2240
rect 6925 -2340 6955 -2310
rect 6925 -2410 6955 -2380
rect 6925 -2475 6955 -2445
rect 6925 -2535 6955 -2505
rect 6925 -2600 6955 -2570
rect 6925 -2670 6955 -2640
rect 6925 -2740 6955 -2710
rect 6925 -2810 6955 -2780
rect 6925 -2875 6955 -2845
rect 6925 -2935 6955 -2905
rect 6925 -3000 6955 -2970
rect 6925 -3070 6955 -3040
rect 6925 -3140 6955 -3110
rect 6925 -3210 6955 -3180
rect 6925 -3275 6955 -3245
rect 6925 -3335 6955 -3305
rect 6925 -3400 6955 -3370
rect 6925 -3470 6955 -3440
rect 6925 -3540 6955 -3510
rect 6925 -3610 6955 -3580
rect 6925 -3675 6955 -3645
rect 6925 -3735 6955 -3705
rect 6925 -3800 6955 -3770
rect 6925 -3870 6955 -3840
rect 6925 -3940 6955 -3910
rect 6925 -4010 6955 -3980
rect 6925 -4075 6955 -4045
rect 6925 -4135 6955 -4105
rect 6925 -4200 6955 -4170
rect 6925 -4270 6955 -4240
rect 6925 -4340 6955 -4310
rect 6925 -4410 6955 -4380
rect 6925 -4475 6955 -4445
rect 7275 -1335 7305 -1305
rect 7275 -1400 7305 -1370
rect 7275 -1470 7305 -1440
rect 7275 -1540 7305 -1510
rect 7275 -1610 7305 -1580
rect 7275 -1675 7305 -1645
rect 7275 -1735 7305 -1705
rect 7275 -1800 7305 -1770
rect 7275 -1870 7305 -1840
rect 7275 -1940 7305 -1910
rect 7275 -2010 7305 -1980
rect 7275 -2075 7305 -2045
rect 7275 -2135 7305 -2105
rect 7275 -2200 7305 -2170
rect 7275 -2270 7305 -2240
rect 7275 -2340 7305 -2310
rect 7275 -2410 7305 -2380
rect 7275 -2475 7305 -2445
rect 7275 -2535 7305 -2505
rect 7275 -2600 7305 -2570
rect 7275 -2670 7305 -2640
rect 7275 -2740 7305 -2710
rect 7275 -2810 7305 -2780
rect 7275 -2875 7305 -2845
rect 7275 -2935 7305 -2905
rect 7275 -3000 7305 -2970
rect 7275 -3070 7305 -3040
rect 7275 -3140 7305 -3110
rect 7275 -3210 7305 -3180
rect 7275 -3275 7305 -3245
rect 7275 -3335 7305 -3305
rect 7275 -3400 7305 -3370
rect 7275 -3470 7305 -3440
rect 7275 -3540 7305 -3510
rect 7275 -3610 7305 -3580
rect 7275 -3675 7305 -3645
rect 7275 -3735 7305 -3705
rect 7275 -3800 7305 -3770
rect 7275 -3870 7305 -3840
rect 7275 -3940 7305 -3910
rect 7275 -4010 7305 -3980
rect 7275 -4075 7305 -4045
rect 7275 -4135 7305 -4105
rect 7275 -4200 7305 -4170
rect 7275 -4270 7305 -4240
rect 7275 -4340 7305 -4310
rect 7275 -4410 7305 -4380
rect 7275 -4475 7305 -4445
rect 7625 -1335 7655 -1305
rect 7625 -1400 7655 -1370
rect 7625 -1470 7655 -1440
rect 7625 -1540 7655 -1510
rect 7625 -1610 7655 -1580
rect 7625 -1675 7655 -1645
rect 7625 -1735 7655 -1705
rect 7625 -1800 7655 -1770
rect 7625 -1870 7655 -1840
rect 7625 -1940 7655 -1910
rect 7625 -2010 7655 -1980
rect 7625 -2075 7655 -2045
rect 7625 -2135 7655 -2105
rect 7625 -2200 7655 -2170
rect 7625 -2270 7655 -2240
rect 7625 -2340 7655 -2310
rect 7625 -2410 7655 -2380
rect 7625 -2475 7655 -2445
rect 7625 -2535 7655 -2505
rect 7625 -2600 7655 -2570
rect 7625 -2670 7655 -2640
rect 7625 -2740 7655 -2710
rect 7625 -2810 7655 -2780
rect 7625 -2875 7655 -2845
rect 7625 -2935 7655 -2905
rect 7625 -3000 7655 -2970
rect 7625 -3070 7655 -3040
rect 7625 -3140 7655 -3110
rect 7625 -3210 7655 -3180
rect 7625 -3275 7655 -3245
rect 7625 -3335 7655 -3305
rect 7625 -3400 7655 -3370
rect 7625 -3470 7655 -3440
rect 7625 -3540 7655 -3510
rect 7625 -3610 7655 -3580
rect 7625 -3675 7655 -3645
rect 7625 -3735 7655 -3705
rect 7625 -3800 7655 -3770
rect 7625 -3870 7655 -3840
rect 7625 -3940 7655 -3910
rect 7625 -4010 7655 -3980
rect 7625 -4075 7655 -4045
rect 7625 -4135 7655 -4105
rect 7625 -4200 7655 -4170
rect 7625 -4270 7655 -4240
rect 7625 -4340 7655 -4310
rect 7625 -4410 7655 -4380
rect 7625 -4475 7655 -4445
rect 7975 -1335 8005 -1305
rect 7975 -1400 8005 -1370
rect 7975 -1470 8005 -1440
rect 7975 -1540 8005 -1510
rect 7975 -1610 8005 -1580
rect 7975 -1675 8005 -1645
rect 7975 -1735 8005 -1705
rect 7975 -1800 8005 -1770
rect 7975 -1870 8005 -1840
rect 7975 -1940 8005 -1910
rect 7975 -2010 8005 -1980
rect 7975 -2075 8005 -2045
rect 7975 -2135 8005 -2105
rect 7975 -2200 8005 -2170
rect 7975 -2270 8005 -2240
rect 7975 -2340 8005 -2310
rect 7975 -2410 8005 -2380
rect 7975 -2475 8005 -2445
rect 7975 -2535 8005 -2505
rect 7975 -2600 8005 -2570
rect 7975 -2670 8005 -2640
rect 7975 -2740 8005 -2710
rect 7975 -2810 8005 -2780
rect 7975 -2875 8005 -2845
rect 7975 -2935 8005 -2905
rect 7975 -3000 8005 -2970
rect 7975 -3070 8005 -3040
rect 7975 -3140 8005 -3110
rect 7975 -3210 8005 -3180
rect 7975 -3275 8005 -3245
rect 7975 -3335 8005 -3305
rect 7975 -3400 8005 -3370
rect 7975 -3470 8005 -3440
rect 7975 -3540 8005 -3510
rect 7975 -3610 8005 -3580
rect 7975 -3675 8005 -3645
rect 7975 -3735 8005 -3705
rect 7975 -3800 8005 -3770
rect 7975 -3870 8005 -3840
rect 7975 -3940 8005 -3910
rect 7975 -4010 8005 -3980
rect 7975 -4075 8005 -4045
rect 7975 -4135 8005 -4105
rect 7975 -4200 8005 -4170
rect 7975 -4270 8005 -4240
rect 7975 -4340 8005 -4310
rect 7975 -4410 8005 -4380
rect 7975 -4475 8005 -4445
rect 8325 -1335 8355 -1305
rect 8325 -1400 8355 -1370
rect 8325 -1470 8355 -1440
rect 8325 -1540 8355 -1510
rect 8325 -1610 8355 -1580
rect 8325 -1675 8355 -1645
rect 8325 -1735 8355 -1705
rect 8325 -1800 8355 -1770
rect 8325 -1870 8355 -1840
rect 8325 -1940 8355 -1910
rect 8325 -2010 8355 -1980
rect 8325 -2075 8355 -2045
rect 8325 -2135 8355 -2105
rect 8325 -2200 8355 -2170
rect 8325 -2270 8355 -2240
rect 8325 -2340 8355 -2310
rect 8325 -2410 8355 -2380
rect 8325 -2475 8355 -2445
rect 8325 -2535 8355 -2505
rect 8325 -2600 8355 -2570
rect 8325 -2670 8355 -2640
rect 8325 -2740 8355 -2710
rect 8325 -2810 8355 -2780
rect 8325 -2875 8355 -2845
rect 8325 -2935 8355 -2905
rect 8325 -3000 8355 -2970
rect 8325 -3070 8355 -3040
rect 8325 -3140 8355 -3110
rect 8325 -3210 8355 -3180
rect 8325 -3275 8355 -3245
rect 8325 -3335 8355 -3305
rect 8325 -3400 8355 -3370
rect 8325 -3470 8355 -3440
rect 8325 -3540 8355 -3510
rect 8325 -3610 8355 -3580
rect 8325 -3675 8355 -3645
rect 8325 -3735 8355 -3705
rect 8325 -3800 8355 -3770
rect 8325 -3870 8355 -3840
rect 8325 -3940 8355 -3910
rect 8325 -4010 8355 -3980
rect 8325 -4075 8355 -4045
rect 8325 -4135 8355 -4105
rect 8325 -4200 8355 -4170
rect 8325 -4270 8355 -4240
rect 8325 -4340 8355 -4310
rect 8325 -4410 8355 -4380
rect 8325 -4475 8355 -4445
rect 8675 -1335 8705 -1305
rect 8675 -1400 8705 -1370
rect 8675 -1470 8705 -1440
rect 8675 -1540 8705 -1510
rect 8675 -1610 8705 -1580
rect 8675 -1675 8705 -1645
rect 8675 -1735 8705 -1705
rect 8675 -1800 8705 -1770
rect 8675 -1870 8705 -1840
rect 8675 -1940 8705 -1910
rect 8675 -2010 8705 -1980
rect 8675 -2075 8705 -2045
rect 8675 -2135 8705 -2105
rect 8675 -2200 8705 -2170
rect 8675 -2270 8705 -2240
rect 8675 -2340 8705 -2310
rect 8675 -2410 8705 -2380
rect 8675 -2475 8705 -2445
rect 8675 -2535 8705 -2505
rect 8675 -2600 8705 -2570
rect 8675 -2670 8705 -2640
rect 8675 -2740 8705 -2710
rect 8675 -2810 8705 -2780
rect 8675 -2875 8705 -2845
rect 8675 -2935 8705 -2905
rect 8675 -3000 8705 -2970
rect 8675 -3070 8705 -3040
rect 8675 -3140 8705 -3110
rect 8675 -3210 8705 -3180
rect 8675 -3275 8705 -3245
rect 8675 -3335 8705 -3305
rect 8675 -3400 8705 -3370
rect 8675 -3470 8705 -3440
rect 8675 -3540 8705 -3510
rect 8675 -3610 8705 -3580
rect 8675 -3675 8705 -3645
rect 8675 -3735 8705 -3705
rect 8675 -3800 8705 -3770
rect 8675 -3870 8705 -3840
rect 8675 -3940 8705 -3910
rect 8675 -4010 8705 -3980
rect 8675 -4075 8705 -4045
rect 8675 -4135 8705 -4105
rect 8675 -4200 8705 -4170
rect 8675 -4270 8705 -4240
rect 8675 -4340 8705 -4310
rect 8675 -4410 8705 -4380
rect 8675 -4475 8705 -4445
rect 9025 -1335 9055 -1305
rect 9025 -1400 9055 -1370
rect 9025 -1470 9055 -1440
rect 9025 -1540 9055 -1510
rect 9025 -1610 9055 -1580
rect 9025 -1675 9055 -1645
rect 9025 -1735 9055 -1705
rect 9025 -1800 9055 -1770
rect 9025 -1870 9055 -1840
rect 9025 -1940 9055 -1910
rect 9025 -2010 9055 -1980
rect 9025 -2075 9055 -2045
rect 9025 -2135 9055 -2105
rect 9025 -2200 9055 -2170
rect 9025 -2270 9055 -2240
rect 9025 -2340 9055 -2310
rect 9025 -2410 9055 -2380
rect 9025 -2475 9055 -2445
rect 9025 -2535 9055 -2505
rect 9025 -2600 9055 -2570
rect 9025 -2670 9055 -2640
rect 9025 -2740 9055 -2710
rect 9025 -2810 9055 -2780
rect 9025 -2875 9055 -2845
rect 9025 -2935 9055 -2905
rect 9025 -3000 9055 -2970
rect 9025 -3070 9055 -3040
rect 9025 -3140 9055 -3110
rect 9025 -3210 9055 -3180
rect 9025 -3275 9055 -3245
rect 9025 -3335 9055 -3305
rect 9025 -3400 9055 -3370
rect 9025 -3470 9055 -3440
rect 9025 -3540 9055 -3510
rect 9025 -3610 9055 -3580
rect 9025 -3675 9055 -3645
rect 9025 -3735 9055 -3705
rect 9025 -3800 9055 -3770
rect 9025 -3870 9055 -3840
rect 9025 -3940 9055 -3910
rect 9025 -4010 9055 -3980
rect 9025 -4075 9055 -4045
rect 9025 -4135 9055 -4105
rect 9025 -4200 9055 -4170
rect 9025 -4270 9055 -4240
rect 9025 -4340 9055 -4310
rect 9025 -4410 9055 -4380
rect 9025 -4475 9055 -4445
<< metal2 >>
rect 2180 20910 2240 20925
rect 2180 20880 2195 20910
rect 2225 20880 2240 20910
rect 2180 20845 2240 20880
rect 2180 20815 2195 20845
rect 2225 20815 2240 20845
rect 2180 20775 2240 20815
rect 2180 20745 2195 20775
rect 2225 20745 2240 20775
rect 2180 20705 2240 20745
rect 2180 20675 2195 20705
rect 2225 20675 2240 20705
rect 2180 20635 2240 20675
rect 2180 20605 2195 20635
rect 2225 20605 2240 20635
rect 2180 20570 2240 20605
rect 2180 20540 2195 20570
rect 2225 20540 2240 20570
rect 2180 20510 2240 20540
rect 2180 20480 2195 20510
rect 2225 20480 2240 20510
rect 2180 20445 2240 20480
rect 2180 20415 2195 20445
rect 2225 20415 2240 20445
rect 2180 20375 2240 20415
rect 2180 20345 2195 20375
rect 2225 20345 2240 20375
rect 2180 20305 2240 20345
rect 2180 20275 2195 20305
rect 2225 20275 2240 20305
rect 2180 20235 2240 20275
rect 2180 20205 2195 20235
rect 2225 20205 2240 20235
rect 2180 20170 2240 20205
rect 2180 20140 2195 20170
rect 2225 20140 2240 20170
rect 2180 20110 2240 20140
rect 2180 20080 2195 20110
rect 2225 20080 2240 20110
rect 2180 20045 2240 20080
rect 2180 20015 2195 20045
rect 2225 20015 2240 20045
rect 2180 19975 2240 20015
rect 2180 19945 2195 19975
rect 2225 19945 2240 19975
rect 2180 19905 2240 19945
rect 2180 19875 2195 19905
rect 2225 19875 2240 19905
rect 2180 19835 2240 19875
rect 2180 19805 2195 19835
rect 2225 19805 2240 19835
rect 2180 19770 2240 19805
rect 2180 19740 2195 19770
rect 2225 19740 2240 19770
rect 2180 19710 2240 19740
rect 2180 19680 2195 19710
rect 2225 19680 2240 19710
rect 2180 19645 2240 19680
rect 2180 19615 2195 19645
rect 2225 19615 2240 19645
rect 2180 19575 2240 19615
rect 2180 19545 2195 19575
rect 2225 19545 2240 19575
rect 2180 19505 2240 19545
rect 2180 19475 2195 19505
rect 2225 19475 2240 19505
rect 2180 19435 2240 19475
rect 2180 19405 2195 19435
rect 2225 19405 2240 19435
rect 2180 19370 2240 19405
rect 2180 19340 2195 19370
rect 2225 19340 2240 19370
rect 2180 19310 2240 19340
rect 2180 19280 2195 19310
rect 2225 19280 2240 19310
rect 2180 19245 2240 19280
rect 2180 19215 2195 19245
rect 2225 19215 2240 19245
rect 2180 19175 2240 19215
rect 2180 19145 2195 19175
rect 2225 19145 2240 19175
rect 2180 19105 2240 19145
rect 2180 19075 2195 19105
rect 2225 19075 2240 19105
rect 2180 19035 2240 19075
rect 2180 19005 2195 19035
rect 2225 19005 2240 19035
rect 2180 18970 2240 19005
rect 2180 18940 2195 18970
rect 2225 18940 2240 18970
rect 2180 18910 2240 18940
rect 2180 18880 2195 18910
rect 2225 18880 2240 18910
rect 2180 18845 2240 18880
rect 2180 18815 2195 18845
rect 2225 18815 2240 18845
rect 2180 18775 2240 18815
rect 2180 18745 2195 18775
rect 2225 18745 2240 18775
rect 2180 18705 2240 18745
rect 2180 18675 2195 18705
rect 2225 18675 2240 18705
rect 2180 18635 2240 18675
rect 2180 18605 2195 18635
rect 2225 18605 2240 18635
rect 2180 18570 2240 18605
rect 2180 18540 2195 18570
rect 2225 18540 2240 18570
rect 2180 18510 2240 18540
rect 2180 18480 2195 18510
rect 2225 18480 2240 18510
rect 2180 18445 2240 18480
rect 2180 18415 2195 18445
rect 2225 18415 2240 18445
rect 2180 18375 2240 18415
rect 2180 18345 2195 18375
rect 2225 18345 2240 18375
rect 2180 18305 2240 18345
rect 2180 18275 2195 18305
rect 2225 18275 2240 18305
rect 2180 18235 2240 18275
rect 2180 18205 2195 18235
rect 2225 18205 2240 18235
rect 2180 18170 2240 18205
rect 2180 18140 2195 18170
rect 2225 18140 2240 18170
rect 2180 18110 2240 18140
rect 2180 18080 2195 18110
rect 2225 18080 2240 18110
rect 2180 18045 2240 18080
rect 2180 18015 2195 18045
rect 2225 18015 2240 18045
rect 2180 17975 2240 18015
rect 2180 17945 2195 17975
rect 2225 17945 2240 17975
rect 2180 17905 2240 17945
rect 2180 17875 2195 17905
rect 2225 17875 2240 17905
rect 2180 17835 2240 17875
rect 2180 17805 2195 17835
rect 2225 17805 2240 17835
rect 2180 17770 2240 17805
rect 2180 17740 2195 17770
rect 2225 17740 2240 17770
rect 2180 17725 2240 17740
rect 6650 20910 6710 20925
rect 6650 20880 6665 20910
rect 6695 20880 6710 20910
rect 6650 20845 6710 20880
rect 6650 20815 6665 20845
rect 6695 20815 6710 20845
rect 6650 20775 6710 20815
rect 6650 20745 6665 20775
rect 6695 20745 6710 20775
rect 6650 20705 6710 20745
rect 6650 20675 6665 20705
rect 6695 20675 6710 20705
rect 6650 20635 6710 20675
rect 6650 20605 6665 20635
rect 6695 20605 6710 20635
rect 6650 20570 6710 20605
rect 6650 20540 6665 20570
rect 6695 20540 6710 20570
rect 6650 20510 6710 20540
rect 6650 20480 6665 20510
rect 6695 20480 6710 20510
rect 6650 20445 6710 20480
rect 6650 20415 6665 20445
rect 6695 20415 6710 20445
rect 6650 20375 6710 20415
rect 6650 20345 6665 20375
rect 6695 20345 6710 20375
rect 6650 20305 6710 20345
rect 6650 20275 6665 20305
rect 6695 20275 6710 20305
rect 6650 20235 6710 20275
rect 6650 20205 6665 20235
rect 6695 20205 6710 20235
rect 6650 20170 6710 20205
rect 6650 20140 6665 20170
rect 6695 20140 6710 20170
rect 6650 20110 6710 20140
rect 6650 20080 6665 20110
rect 6695 20080 6710 20110
rect 6650 20045 6710 20080
rect 6650 20015 6665 20045
rect 6695 20015 6710 20045
rect 6650 19975 6710 20015
rect 6650 19945 6665 19975
rect 6695 19945 6710 19975
rect 6650 19905 6710 19945
rect 6650 19875 6665 19905
rect 6695 19875 6710 19905
rect 6650 19835 6710 19875
rect 6650 19805 6665 19835
rect 6695 19805 6710 19835
rect 6650 19770 6710 19805
rect 6650 19740 6665 19770
rect 6695 19740 6710 19770
rect 6650 19710 6710 19740
rect 6650 19680 6665 19710
rect 6695 19680 6710 19710
rect 6650 19645 6710 19680
rect 6650 19615 6665 19645
rect 6695 19615 6710 19645
rect 6650 19575 6710 19615
rect 6650 19545 6665 19575
rect 6695 19545 6710 19575
rect 6650 19505 6710 19545
rect 6650 19475 6665 19505
rect 6695 19475 6710 19505
rect 6650 19435 6710 19475
rect 6650 19405 6665 19435
rect 6695 19405 6710 19435
rect 6650 19370 6710 19405
rect 6650 19340 6665 19370
rect 6695 19340 6710 19370
rect 6650 19310 6710 19340
rect 6650 19280 6665 19310
rect 6695 19280 6710 19310
rect 6650 19245 6710 19280
rect 6650 19215 6665 19245
rect 6695 19215 6710 19245
rect 6650 19175 6710 19215
rect 6650 19145 6665 19175
rect 6695 19145 6710 19175
rect 6650 19105 6710 19145
rect 6650 19075 6665 19105
rect 6695 19075 6710 19105
rect 6650 19035 6710 19075
rect 6650 19005 6665 19035
rect 6695 19005 6710 19035
rect 6650 18970 6710 19005
rect 6650 18940 6665 18970
rect 6695 18940 6710 18970
rect 6650 18910 6710 18940
rect 6650 18880 6665 18910
rect 6695 18880 6710 18910
rect 6650 18845 6710 18880
rect 6650 18815 6665 18845
rect 6695 18815 6710 18845
rect 6650 18775 6710 18815
rect 6650 18745 6665 18775
rect 6695 18745 6710 18775
rect 6650 18705 6710 18745
rect 6650 18675 6665 18705
rect 6695 18675 6710 18705
rect 6650 18635 6710 18675
rect 6650 18605 6665 18635
rect 6695 18605 6710 18635
rect 6650 18570 6710 18605
rect 6650 18540 6665 18570
rect 6695 18540 6710 18570
rect 6650 18510 6710 18540
rect 6650 18480 6665 18510
rect 6695 18480 6710 18510
rect 6650 18445 6710 18480
rect 6650 18415 6665 18445
rect 6695 18415 6710 18445
rect 6650 18375 6710 18415
rect 6650 18345 6665 18375
rect 6695 18345 6710 18375
rect 6650 18305 6710 18345
rect 6650 18275 6665 18305
rect 6695 18275 6710 18305
rect 6650 18235 6710 18275
rect 6650 18205 6665 18235
rect 6695 18205 6710 18235
rect 6650 18170 6710 18205
rect 6650 18140 6665 18170
rect 6695 18140 6710 18170
rect 6650 18110 6710 18140
rect 6650 18080 6665 18110
rect 6695 18080 6710 18110
rect 6650 18045 6710 18080
rect 6650 18015 6665 18045
rect 6695 18015 6710 18045
rect 6650 17975 6710 18015
rect 6650 17945 6665 17975
rect 6695 17945 6710 17975
rect 6650 17905 6710 17945
rect 6650 17875 6665 17905
rect 6695 17875 6710 17905
rect 6650 17835 6710 17875
rect 6650 17805 6665 17835
rect 6695 17805 6710 17835
rect 6650 17770 6710 17805
rect 6650 17740 6665 17770
rect 6695 17740 6710 17770
rect 6650 17725 6710 17740
rect 2285 15925 2405 15930
rect 2285 15895 2290 15925
rect 2320 15895 2330 15925
rect 2360 15895 2370 15925
rect 2400 15895 2405 15925
rect 2285 15890 2405 15895
rect 2150 15780 2270 15785
rect 2150 15750 2155 15780
rect 2185 15750 2195 15780
rect 2225 15750 2235 15780
rect 2265 15775 2270 15780
rect 2265 15750 4470 15775
rect 2150 15740 4470 15750
rect 2150 15710 2155 15740
rect 2185 15710 2195 15740
rect 2225 15710 2235 15740
rect 2265 15710 2975 15740
rect 3005 15710 3300 15740
rect 3330 15710 4470 15740
rect 2150 15700 4470 15710
rect 2150 15670 2155 15700
rect 2185 15670 2195 15700
rect 2225 15670 2235 15700
rect 2265 15670 2975 15700
rect 3005 15670 3300 15700
rect 3330 15670 4470 15700
rect 5685 15705 6740 15710
rect 5685 15675 6625 15705
rect 6655 15675 6665 15705
rect 6695 15675 6705 15705
rect 6735 15675 6740 15705
rect 5685 15670 6740 15675
rect 2150 15665 4470 15670
rect 5645 15665 6740 15670
rect 5645 15635 5650 15665
rect 5680 15635 5975 15665
rect 6005 15635 6625 15665
rect 6655 15635 6665 15665
rect 6695 15635 6705 15665
rect 6735 15635 6740 15665
rect 5645 15625 6740 15635
rect 5645 15595 5650 15625
rect 5680 15595 5975 15625
rect 6005 15595 6625 15625
rect 6655 15595 6665 15625
rect 6695 15595 6705 15625
rect 6735 15595 6740 15625
rect 5645 15590 6740 15595
rect 5690 13005 6740 13010
rect 5690 12975 6625 13005
rect 6655 12975 6665 13005
rect 6695 12975 6705 13005
rect 6735 12975 6740 13005
rect 5690 12965 6740 12975
rect 5690 12935 6625 12965
rect 6655 12935 6665 12965
rect 6695 12935 6705 12965
rect 6735 12935 6740 12965
rect 5690 12925 6740 12935
rect 5690 12895 6625 12925
rect 6655 12895 6665 12925
rect 6695 12895 6705 12925
rect 6735 12895 6740 12925
rect 5690 12890 6740 12895
rect 2150 12720 3355 12725
rect 2150 12690 2155 12720
rect 2185 12690 2195 12720
rect 2225 12690 2235 12720
rect 2265 12690 3355 12720
rect 2150 12680 3355 12690
rect 2150 12650 2155 12680
rect 2185 12650 2195 12680
rect 2225 12650 2235 12680
rect 2265 12650 3355 12680
rect 2150 12645 3355 12650
rect 2150 12560 3800 12565
rect 2150 12530 2155 12560
rect 2185 12530 2195 12560
rect 2225 12530 2235 12560
rect 2265 12530 3800 12560
rect 2150 12520 3800 12530
rect 2150 12490 2155 12520
rect 2185 12490 2195 12520
rect 2225 12490 2235 12520
rect 2265 12490 3800 12520
rect 2150 12480 3800 12490
rect 2150 12450 2155 12480
rect 2185 12450 2195 12480
rect 2225 12450 2235 12480
rect 2265 12450 3800 12480
rect 2150 12445 3800 12450
rect 5670 12160 6710 12165
rect 5670 12130 6595 12160
rect 6625 12130 6635 12160
rect 6665 12130 6675 12160
rect 6705 12130 6710 12160
rect 5670 12120 6710 12130
rect 5670 12090 6595 12120
rect 6625 12090 6635 12120
rect 6665 12090 6675 12120
rect 6705 12090 6710 12120
rect 5670 12080 6710 12090
rect 5670 12050 6595 12080
rect 6625 12050 6635 12080
rect 6665 12050 6675 12080
rect 6705 12050 6710 12080
rect 5670 12045 6710 12050
rect 5870 11205 6710 11210
rect 5870 11175 6595 11205
rect 6625 11175 6635 11205
rect 6665 11175 6675 11205
rect 6705 11175 6710 11205
rect 5870 11165 6710 11175
rect 5870 11135 6595 11165
rect 6625 11135 6635 11165
rect 6665 11135 6675 11165
rect 6705 11135 6710 11165
rect 5870 11125 6710 11135
rect 5870 11095 6595 11125
rect 6625 11095 6635 11125
rect 6665 11095 6675 11125
rect 6705 11095 6710 11125
rect 5870 11090 6710 11095
rect 5855 10500 6710 10505
rect 5855 10470 6595 10500
rect 6625 10470 6635 10500
rect 6665 10470 6675 10500
rect 6705 10470 6710 10500
rect 5855 10460 6710 10470
rect 5855 10430 6595 10460
rect 6625 10430 6635 10460
rect 6665 10430 6675 10460
rect 6705 10430 6710 10460
rect 5855 10420 6710 10430
rect 5855 10390 6595 10420
rect 6625 10390 6635 10420
rect 6665 10390 6675 10420
rect 6705 10390 6710 10420
rect 5855 10385 6710 10390
rect 5925 10035 6710 10040
rect 5925 10005 6595 10035
rect 6625 10005 6635 10035
rect 6665 10005 6675 10035
rect 6705 10005 6710 10035
rect 5925 9995 6710 10005
rect 5925 9965 6595 9995
rect 6625 9965 6635 9995
rect 6665 9965 6675 9995
rect 6705 9965 6710 9995
rect 5925 9955 6710 9965
rect 5925 9925 6595 9955
rect 6625 9925 6635 9955
rect 6665 9925 6675 9955
rect 6705 9925 6710 9955
rect 5925 9920 6710 9925
rect -90 9635 -30 9650
rect -90 9605 -75 9635
rect -45 9605 -30 9635
rect -90 9570 -30 9605
rect -90 9540 -75 9570
rect -45 9540 -30 9570
rect -90 9500 -30 9540
rect -90 9470 -75 9500
rect -45 9470 -30 9500
rect -90 9430 -30 9470
rect -90 9400 -75 9430
rect -45 9400 -30 9430
rect -90 9360 -30 9400
rect -90 9330 -75 9360
rect -45 9330 -30 9360
rect -90 9295 -30 9330
rect -90 9265 -75 9295
rect -45 9265 -30 9295
rect -90 9235 -30 9265
rect -90 9205 -75 9235
rect -45 9205 -30 9235
rect -90 9170 -30 9205
rect -90 9140 -75 9170
rect -45 9140 -30 9170
rect -90 9100 -30 9140
rect -90 9070 -75 9100
rect -45 9070 -30 9100
rect -90 9030 -30 9070
rect -90 9000 -75 9030
rect -45 9000 -30 9030
rect -90 8960 -30 9000
rect -90 8930 -75 8960
rect -45 8930 -30 8960
rect -90 8895 -30 8930
rect -90 8865 -75 8895
rect -45 8865 -30 8895
rect -90 8835 -30 8865
rect -90 8805 -75 8835
rect -45 8805 -30 8835
rect -90 8770 -30 8805
rect -90 8740 -75 8770
rect -45 8740 -30 8770
rect -90 8700 -30 8740
rect -90 8670 -75 8700
rect -45 8670 -30 8700
rect -90 8630 -30 8670
rect -90 8600 -75 8630
rect -45 8600 -30 8630
rect -90 8560 -30 8600
rect -90 8530 -75 8560
rect -45 8530 -30 8560
rect -90 8495 -30 8530
rect -90 8465 -75 8495
rect -45 8465 -30 8495
rect -90 8435 -30 8465
rect -90 8405 -75 8435
rect -45 8405 -30 8435
rect -90 8370 -30 8405
rect -90 8340 -75 8370
rect -45 8340 -30 8370
rect -90 8300 -30 8340
rect -90 8270 -75 8300
rect -45 8270 -30 8300
rect -90 8230 -30 8270
rect -90 8200 -75 8230
rect -45 8200 -30 8230
rect -90 8160 -30 8200
rect -90 8130 -75 8160
rect -45 8130 -30 8160
rect -90 8095 -30 8130
rect -90 8065 -75 8095
rect -45 8065 -30 8095
rect -90 8035 -30 8065
rect -90 8005 -75 8035
rect -45 8005 -30 8035
rect -90 7970 -30 8005
rect -90 7940 -75 7970
rect -45 7940 -30 7970
rect -90 7900 -30 7940
rect -90 7870 -75 7900
rect -45 7870 -30 7900
rect -90 7830 -30 7870
rect -90 7800 -75 7830
rect -45 7800 -30 7830
rect -90 7760 -30 7800
rect -90 7730 -75 7760
rect -45 7730 -30 7760
rect -90 7695 -30 7730
rect -90 7665 -75 7695
rect -45 7665 -30 7695
rect -90 7635 -30 7665
rect -90 7605 -75 7635
rect -45 7605 -30 7635
rect -90 7570 -30 7605
rect -90 7540 -75 7570
rect -45 7540 -30 7570
rect -90 7500 -30 7540
rect -90 7470 -75 7500
rect -45 7470 -30 7500
rect -90 7430 -30 7470
rect -90 7400 -75 7430
rect -45 7400 -30 7430
rect -90 7360 -30 7400
rect -90 7330 -75 7360
rect -45 7330 -30 7360
rect -90 7295 -30 7330
rect -90 7265 -75 7295
rect -45 7265 -30 7295
rect -90 7235 -30 7265
rect -90 7205 -75 7235
rect -45 7205 -30 7235
rect -90 7170 -30 7205
rect -90 7140 -75 7170
rect -45 7140 -30 7170
rect -90 7100 -30 7140
rect -90 7070 -75 7100
rect -45 7070 -30 7100
rect -90 7030 -30 7070
rect -90 7000 -75 7030
rect -45 7000 -30 7030
rect -90 6960 -30 7000
rect -90 6930 -75 6960
rect -45 6930 -30 6960
rect -90 6895 -30 6930
rect -90 6865 -75 6895
rect -45 6865 -30 6895
rect -90 6835 -30 6865
rect -90 6805 -75 6835
rect -45 6805 -30 6835
rect -90 6770 -30 6805
rect -90 6740 -75 6770
rect -45 6740 -30 6770
rect -90 6700 -30 6740
rect -90 6670 -75 6700
rect -45 6670 -30 6700
rect -90 6630 -30 6670
rect -90 6600 -75 6630
rect -45 6600 -30 6630
rect -90 6560 -30 6600
rect -90 6530 -75 6560
rect -45 6530 -30 6560
rect -90 6495 -30 6530
rect -90 6465 -75 6495
rect -45 6465 -30 6495
rect -90 6450 -30 6465
rect 260 9635 320 9650
rect 260 9605 275 9635
rect 305 9605 320 9635
rect 260 9570 320 9605
rect 260 9540 275 9570
rect 305 9540 320 9570
rect 260 9500 320 9540
rect 260 9470 275 9500
rect 305 9470 320 9500
rect 260 9430 320 9470
rect 260 9400 275 9430
rect 305 9400 320 9430
rect 260 9360 320 9400
rect 260 9330 275 9360
rect 305 9330 320 9360
rect 260 9295 320 9330
rect 260 9265 275 9295
rect 305 9265 320 9295
rect 260 9235 320 9265
rect 260 9205 275 9235
rect 305 9205 320 9235
rect 260 9170 320 9205
rect 260 9140 275 9170
rect 305 9140 320 9170
rect 260 9100 320 9140
rect 260 9070 275 9100
rect 305 9070 320 9100
rect 260 9030 320 9070
rect 260 9000 275 9030
rect 305 9000 320 9030
rect 260 8960 320 9000
rect 260 8930 275 8960
rect 305 8930 320 8960
rect 260 8895 320 8930
rect 260 8865 275 8895
rect 305 8865 320 8895
rect 260 8835 320 8865
rect 260 8805 275 8835
rect 305 8805 320 8835
rect 260 8770 320 8805
rect 260 8740 275 8770
rect 305 8740 320 8770
rect 260 8700 320 8740
rect 260 8670 275 8700
rect 305 8670 320 8700
rect 260 8630 320 8670
rect 260 8600 275 8630
rect 305 8600 320 8630
rect 260 8560 320 8600
rect 260 8530 275 8560
rect 305 8530 320 8560
rect 260 8495 320 8530
rect 260 8465 275 8495
rect 305 8465 320 8495
rect 260 8435 320 8465
rect 260 8405 275 8435
rect 305 8405 320 8435
rect 260 8370 320 8405
rect 260 8340 275 8370
rect 305 8340 320 8370
rect 260 8300 320 8340
rect 260 8270 275 8300
rect 305 8270 320 8300
rect 260 8230 320 8270
rect 260 8200 275 8230
rect 305 8200 320 8230
rect 260 8160 320 8200
rect 260 8130 275 8160
rect 305 8130 320 8160
rect 260 8095 320 8130
rect 260 8065 275 8095
rect 305 8065 320 8095
rect 260 8035 320 8065
rect 260 8005 275 8035
rect 305 8005 320 8035
rect 260 7970 320 8005
rect 260 7940 275 7970
rect 305 7940 320 7970
rect 260 7900 320 7940
rect 260 7870 275 7900
rect 305 7870 320 7900
rect 260 7830 320 7870
rect 260 7800 275 7830
rect 305 7800 320 7830
rect 260 7760 320 7800
rect 260 7730 275 7760
rect 305 7730 320 7760
rect 260 7695 320 7730
rect 260 7665 275 7695
rect 305 7665 320 7695
rect 260 7635 320 7665
rect 260 7605 275 7635
rect 305 7605 320 7635
rect 260 7570 320 7605
rect 260 7540 275 7570
rect 305 7540 320 7570
rect 260 7500 320 7540
rect 260 7470 275 7500
rect 305 7470 320 7500
rect 260 7430 320 7470
rect 260 7400 275 7430
rect 305 7400 320 7430
rect 260 7360 320 7400
rect 260 7330 275 7360
rect 305 7330 320 7360
rect 260 7295 320 7330
rect 260 7265 275 7295
rect 305 7265 320 7295
rect 260 7235 320 7265
rect 260 7205 275 7235
rect 305 7205 320 7235
rect 260 7170 320 7205
rect 260 7140 275 7170
rect 305 7140 320 7170
rect 260 7100 320 7140
rect 260 7070 275 7100
rect 305 7070 320 7100
rect 260 7030 320 7070
rect 260 7000 275 7030
rect 305 7000 320 7030
rect 260 6960 320 7000
rect 260 6930 275 6960
rect 305 6930 320 6960
rect 260 6895 320 6930
rect 260 6865 275 6895
rect 305 6865 320 6895
rect 260 6835 320 6865
rect 260 6805 275 6835
rect 305 6805 320 6835
rect 260 6770 320 6805
rect 260 6740 275 6770
rect 305 6740 320 6770
rect 260 6700 320 6740
rect 260 6670 275 6700
rect 305 6670 320 6700
rect 260 6630 320 6670
rect 260 6600 275 6630
rect 305 6600 320 6630
rect 260 6560 320 6600
rect 260 6530 275 6560
rect 305 6530 320 6560
rect 260 6495 320 6530
rect 260 6465 275 6495
rect 305 6465 320 6495
rect 260 6450 320 6465
rect 610 9635 670 9650
rect 610 9605 625 9635
rect 655 9605 670 9635
rect 610 9570 670 9605
rect 610 9540 625 9570
rect 655 9540 670 9570
rect 610 9500 670 9540
rect 610 9470 625 9500
rect 655 9470 670 9500
rect 610 9430 670 9470
rect 610 9400 625 9430
rect 655 9400 670 9430
rect 610 9360 670 9400
rect 610 9330 625 9360
rect 655 9330 670 9360
rect 610 9295 670 9330
rect 610 9265 625 9295
rect 655 9265 670 9295
rect 610 9235 670 9265
rect 610 9205 625 9235
rect 655 9205 670 9235
rect 610 9170 670 9205
rect 610 9140 625 9170
rect 655 9140 670 9170
rect 610 9100 670 9140
rect 610 9070 625 9100
rect 655 9070 670 9100
rect 610 9030 670 9070
rect 610 9000 625 9030
rect 655 9000 670 9030
rect 610 8960 670 9000
rect 610 8930 625 8960
rect 655 8930 670 8960
rect 610 8895 670 8930
rect 610 8865 625 8895
rect 655 8865 670 8895
rect 610 8835 670 8865
rect 610 8805 625 8835
rect 655 8805 670 8835
rect 610 8770 670 8805
rect 610 8740 625 8770
rect 655 8740 670 8770
rect 610 8700 670 8740
rect 610 8670 625 8700
rect 655 8670 670 8700
rect 610 8630 670 8670
rect 610 8600 625 8630
rect 655 8600 670 8630
rect 610 8560 670 8600
rect 610 8530 625 8560
rect 655 8530 670 8560
rect 610 8495 670 8530
rect 610 8465 625 8495
rect 655 8465 670 8495
rect 610 8435 670 8465
rect 610 8405 625 8435
rect 655 8405 670 8435
rect 610 8370 670 8405
rect 610 8340 625 8370
rect 655 8340 670 8370
rect 610 8300 670 8340
rect 610 8270 625 8300
rect 655 8270 670 8300
rect 610 8230 670 8270
rect 610 8200 625 8230
rect 655 8200 670 8230
rect 610 8160 670 8200
rect 610 8130 625 8160
rect 655 8130 670 8160
rect 610 8095 670 8130
rect 610 8065 625 8095
rect 655 8065 670 8095
rect 610 8035 670 8065
rect 610 8005 625 8035
rect 655 8005 670 8035
rect 610 7970 670 8005
rect 610 7940 625 7970
rect 655 7940 670 7970
rect 610 7900 670 7940
rect 610 7870 625 7900
rect 655 7870 670 7900
rect 610 7830 670 7870
rect 610 7800 625 7830
rect 655 7800 670 7830
rect 610 7760 670 7800
rect 610 7730 625 7760
rect 655 7730 670 7760
rect 610 7695 670 7730
rect 610 7665 625 7695
rect 655 7665 670 7695
rect 610 7635 670 7665
rect 610 7605 625 7635
rect 655 7605 670 7635
rect 610 7570 670 7605
rect 610 7540 625 7570
rect 655 7540 670 7570
rect 610 7500 670 7540
rect 610 7470 625 7500
rect 655 7470 670 7500
rect 610 7430 670 7470
rect 610 7400 625 7430
rect 655 7400 670 7430
rect 610 7360 670 7400
rect 610 7330 625 7360
rect 655 7330 670 7360
rect 610 7295 670 7330
rect 610 7265 625 7295
rect 655 7265 670 7295
rect 610 7235 670 7265
rect 610 7205 625 7235
rect 655 7205 670 7235
rect 610 7170 670 7205
rect 610 7140 625 7170
rect 655 7140 670 7170
rect 610 7100 670 7140
rect 610 7070 625 7100
rect 655 7070 670 7100
rect 610 7030 670 7070
rect 610 7000 625 7030
rect 655 7000 670 7030
rect 610 6960 670 7000
rect 610 6930 625 6960
rect 655 6930 670 6960
rect 610 6895 670 6930
rect 610 6865 625 6895
rect 655 6865 670 6895
rect 610 6835 670 6865
rect 610 6805 625 6835
rect 655 6805 670 6835
rect 610 6770 670 6805
rect 610 6740 625 6770
rect 655 6740 670 6770
rect 610 6700 670 6740
rect 610 6670 625 6700
rect 655 6670 670 6700
rect 610 6630 670 6670
rect 610 6600 625 6630
rect 655 6600 670 6630
rect 610 6560 670 6600
rect 610 6530 625 6560
rect 655 6530 670 6560
rect 610 6495 670 6530
rect 610 6465 625 6495
rect 655 6465 670 6495
rect 610 6450 670 6465
rect 960 9635 1020 9650
rect 960 9605 975 9635
rect 1005 9605 1020 9635
rect 960 9570 1020 9605
rect 960 9540 975 9570
rect 1005 9540 1020 9570
rect 960 9500 1020 9540
rect 960 9470 975 9500
rect 1005 9470 1020 9500
rect 960 9430 1020 9470
rect 960 9400 975 9430
rect 1005 9400 1020 9430
rect 960 9360 1020 9400
rect 960 9330 975 9360
rect 1005 9330 1020 9360
rect 960 9295 1020 9330
rect 960 9265 975 9295
rect 1005 9265 1020 9295
rect 960 9235 1020 9265
rect 960 9205 975 9235
rect 1005 9205 1020 9235
rect 960 9170 1020 9205
rect 960 9140 975 9170
rect 1005 9140 1020 9170
rect 960 9100 1020 9140
rect 960 9070 975 9100
rect 1005 9070 1020 9100
rect 960 9030 1020 9070
rect 960 9000 975 9030
rect 1005 9000 1020 9030
rect 960 8960 1020 9000
rect 960 8930 975 8960
rect 1005 8930 1020 8960
rect 960 8895 1020 8930
rect 960 8865 975 8895
rect 1005 8865 1020 8895
rect 960 8835 1020 8865
rect 960 8805 975 8835
rect 1005 8805 1020 8835
rect 960 8770 1020 8805
rect 960 8740 975 8770
rect 1005 8740 1020 8770
rect 960 8700 1020 8740
rect 960 8670 975 8700
rect 1005 8670 1020 8700
rect 960 8630 1020 8670
rect 960 8600 975 8630
rect 1005 8600 1020 8630
rect 960 8560 1020 8600
rect 960 8530 975 8560
rect 1005 8530 1020 8560
rect 960 8495 1020 8530
rect 960 8465 975 8495
rect 1005 8465 1020 8495
rect 960 8435 1020 8465
rect 960 8405 975 8435
rect 1005 8405 1020 8435
rect 960 8370 1020 8405
rect 960 8340 975 8370
rect 1005 8340 1020 8370
rect 960 8300 1020 8340
rect 960 8270 975 8300
rect 1005 8270 1020 8300
rect 960 8230 1020 8270
rect 960 8200 975 8230
rect 1005 8200 1020 8230
rect 960 8160 1020 8200
rect 960 8130 975 8160
rect 1005 8130 1020 8160
rect 960 8095 1020 8130
rect 960 8065 975 8095
rect 1005 8065 1020 8095
rect 960 8035 1020 8065
rect 960 8005 975 8035
rect 1005 8005 1020 8035
rect 960 7970 1020 8005
rect 960 7940 975 7970
rect 1005 7940 1020 7970
rect 960 7900 1020 7940
rect 960 7870 975 7900
rect 1005 7870 1020 7900
rect 960 7830 1020 7870
rect 960 7800 975 7830
rect 1005 7800 1020 7830
rect 960 7760 1020 7800
rect 960 7730 975 7760
rect 1005 7730 1020 7760
rect 960 7695 1020 7730
rect 960 7665 975 7695
rect 1005 7665 1020 7695
rect 960 7635 1020 7665
rect 960 7605 975 7635
rect 1005 7605 1020 7635
rect 960 7570 1020 7605
rect 960 7540 975 7570
rect 1005 7540 1020 7570
rect 960 7500 1020 7540
rect 960 7470 975 7500
rect 1005 7470 1020 7500
rect 960 7430 1020 7470
rect 960 7400 975 7430
rect 1005 7400 1020 7430
rect 960 7360 1020 7400
rect 960 7330 975 7360
rect 1005 7330 1020 7360
rect 960 7295 1020 7330
rect 960 7265 975 7295
rect 1005 7265 1020 7295
rect 960 7235 1020 7265
rect 960 7205 975 7235
rect 1005 7205 1020 7235
rect 960 7170 1020 7205
rect 960 7140 975 7170
rect 1005 7140 1020 7170
rect 960 7100 1020 7140
rect 960 7070 975 7100
rect 1005 7070 1020 7100
rect 960 7030 1020 7070
rect 960 7000 975 7030
rect 1005 7000 1020 7030
rect 960 6960 1020 7000
rect 960 6930 975 6960
rect 1005 6930 1020 6960
rect 960 6895 1020 6930
rect 960 6865 975 6895
rect 1005 6865 1020 6895
rect 960 6835 1020 6865
rect 960 6805 975 6835
rect 1005 6805 1020 6835
rect 960 6770 1020 6805
rect 960 6740 975 6770
rect 1005 6740 1020 6770
rect 960 6700 1020 6740
rect 960 6670 975 6700
rect 1005 6670 1020 6700
rect 960 6630 1020 6670
rect 960 6600 975 6630
rect 1005 6600 1020 6630
rect 960 6560 1020 6600
rect 960 6530 975 6560
rect 1005 6530 1020 6560
rect 960 6495 1020 6530
rect 960 6465 975 6495
rect 1005 6465 1020 6495
rect 960 6450 1020 6465
rect 1660 9635 1720 9650
rect 1660 9605 1675 9635
rect 1705 9605 1720 9635
rect 1660 9570 1720 9605
rect 1660 9540 1675 9570
rect 1705 9540 1720 9570
rect 1660 9500 1720 9540
rect 1660 9470 1675 9500
rect 1705 9470 1720 9500
rect 1660 9430 1720 9470
rect 1660 9400 1675 9430
rect 1705 9400 1720 9430
rect 1660 9360 1720 9400
rect 1660 9330 1675 9360
rect 1705 9330 1720 9360
rect 1660 9295 1720 9330
rect 1660 9265 1675 9295
rect 1705 9265 1720 9295
rect 1660 9235 1720 9265
rect 1660 9205 1675 9235
rect 1705 9205 1720 9235
rect 1660 9170 1720 9205
rect 1660 9140 1675 9170
rect 1705 9140 1720 9170
rect 1660 9100 1720 9140
rect 1660 9070 1675 9100
rect 1705 9070 1720 9100
rect 1660 9030 1720 9070
rect 1660 9000 1675 9030
rect 1705 9000 1720 9030
rect 1660 8960 1720 9000
rect 1660 8930 1675 8960
rect 1705 8930 1720 8960
rect 1660 8895 1720 8930
rect 1660 8865 1675 8895
rect 1705 8865 1720 8895
rect 1660 8835 1720 8865
rect 1660 8805 1675 8835
rect 1705 8805 1720 8835
rect 1660 8770 1720 8805
rect 1660 8740 1675 8770
rect 1705 8740 1720 8770
rect 1660 8700 1720 8740
rect 1660 8670 1675 8700
rect 1705 8670 1720 8700
rect 1660 8630 1720 8670
rect 1660 8600 1675 8630
rect 1705 8600 1720 8630
rect 1660 8560 1720 8600
rect 1660 8530 1675 8560
rect 1705 8530 1720 8560
rect 1660 8495 1720 8530
rect 1660 8465 1675 8495
rect 1705 8465 1720 8495
rect 1660 8435 1720 8465
rect 1660 8405 1675 8435
rect 1705 8405 1720 8435
rect 1660 8370 1720 8405
rect 1660 8340 1675 8370
rect 1705 8340 1720 8370
rect 1660 8300 1720 8340
rect 1660 8270 1675 8300
rect 1705 8270 1720 8300
rect 1660 8230 1720 8270
rect 1660 8200 1675 8230
rect 1705 8200 1720 8230
rect 1660 8160 1720 8200
rect 1660 8130 1675 8160
rect 1705 8130 1720 8160
rect 1660 8095 1720 8130
rect 1660 8065 1675 8095
rect 1705 8065 1720 8095
rect 1660 8035 1720 8065
rect 1660 8005 1675 8035
rect 1705 8005 1720 8035
rect 1660 7970 1720 8005
rect 1660 7940 1675 7970
rect 1705 7940 1720 7970
rect 1660 7900 1720 7940
rect 1660 7870 1675 7900
rect 1705 7870 1720 7900
rect 1660 7830 1720 7870
rect 1660 7800 1675 7830
rect 1705 7800 1720 7830
rect 1660 7760 1720 7800
rect 1660 7730 1675 7760
rect 1705 7730 1720 7760
rect 1660 7695 1720 7730
rect 1660 7665 1675 7695
rect 1705 7665 1720 7695
rect 1660 7635 1720 7665
rect 1660 7605 1675 7635
rect 1705 7605 1720 7635
rect 1660 7570 1720 7605
rect 1660 7540 1675 7570
rect 1705 7540 1720 7570
rect 1660 7500 1720 7540
rect 1660 7470 1675 7500
rect 1705 7470 1720 7500
rect 1660 7430 1720 7470
rect 1660 7400 1675 7430
rect 1705 7400 1720 7430
rect 1660 7360 1720 7400
rect 1660 7330 1675 7360
rect 1705 7330 1720 7360
rect 1660 7295 1720 7330
rect 1660 7265 1675 7295
rect 1705 7265 1720 7295
rect 1660 7235 1720 7265
rect 1660 7205 1675 7235
rect 1705 7205 1720 7235
rect 1660 7170 1720 7205
rect 1660 7140 1675 7170
rect 1705 7140 1720 7170
rect 1660 7100 1720 7140
rect 1660 7070 1675 7100
rect 1705 7070 1720 7100
rect 1660 7030 1720 7070
rect 1660 7000 1675 7030
rect 1705 7000 1720 7030
rect 1660 6960 1720 7000
rect 1660 6930 1675 6960
rect 1705 6930 1720 6960
rect 1660 6895 1720 6930
rect 1660 6865 1675 6895
rect 1705 6865 1720 6895
rect 1660 6835 1720 6865
rect 1660 6805 1675 6835
rect 1705 6805 1720 6835
rect 1660 6770 1720 6805
rect 1660 6740 1675 6770
rect 1705 6740 1720 6770
rect 1660 6700 1720 6740
rect 1660 6670 1675 6700
rect 1705 6670 1720 6700
rect 1660 6630 1720 6670
rect 1660 6600 1675 6630
rect 1705 6600 1720 6630
rect 1660 6560 1720 6600
rect 1660 6530 1675 6560
rect 1705 6530 1720 6560
rect 1660 6495 1720 6530
rect 1660 6465 1675 6495
rect 1705 6465 1720 6495
rect 1660 6450 1720 6465
rect 2315 9635 2375 9650
rect 2315 9605 2330 9635
rect 2360 9605 2375 9635
rect 2315 9570 2375 9605
rect 2315 9540 2330 9570
rect 2360 9540 2375 9570
rect 2315 9500 2375 9540
rect 2315 9470 2330 9500
rect 2360 9470 2375 9500
rect 2315 9430 2375 9470
rect 2315 9400 2330 9430
rect 2360 9400 2375 9430
rect 2315 9360 2375 9400
rect 2315 9330 2330 9360
rect 2360 9330 2375 9360
rect 2315 9295 2375 9330
rect 2315 9265 2330 9295
rect 2360 9265 2375 9295
rect 2315 9235 2375 9265
rect 2315 9205 2330 9235
rect 2360 9205 2375 9235
rect 2315 9170 2375 9205
rect 2315 9140 2330 9170
rect 2360 9140 2375 9170
rect 2315 9100 2375 9140
rect 2315 9070 2330 9100
rect 2360 9070 2375 9100
rect 2315 9030 2375 9070
rect 2315 9000 2330 9030
rect 2360 9000 2375 9030
rect 2315 8960 2375 9000
rect 2315 8930 2330 8960
rect 2360 8930 2375 8960
rect 2315 8895 2375 8930
rect 2315 8865 2330 8895
rect 2360 8865 2375 8895
rect 2315 8835 2375 8865
rect 2315 8805 2330 8835
rect 2360 8805 2375 8835
rect 2315 8770 2375 8805
rect 2315 8740 2330 8770
rect 2360 8740 2375 8770
rect 2315 8700 2375 8740
rect 2315 8670 2330 8700
rect 2360 8670 2375 8700
rect 2315 8630 2375 8670
rect 2315 8600 2330 8630
rect 2360 8600 2375 8630
rect 2315 8560 2375 8600
rect 2315 8530 2330 8560
rect 2360 8530 2375 8560
rect 2315 8495 2375 8530
rect 2315 8465 2330 8495
rect 2360 8465 2375 8495
rect 2315 8435 2375 8465
rect 2315 8405 2330 8435
rect 2360 8405 2375 8435
rect 2315 8370 2375 8405
rect 2315 8340 2330 8370
rect 2360 8340 2375 8370
rect 2315 8300 2375 8340
rect 2315 8270 2330 8300
rect 2360 8270 2375 8300
rect 2315 8230 2375 8270
rect 2315 8200 2330 8230
rect 2360 8200 2375 8230
rect 2315 8160 2375 8200
rect 2315 8130 2330 8160
rect 2360 8130 2375 8160
rect 2315 8095 2375 8130
rect 2315 8065 2330 8095
rect 2360 8065 2375 8095
rect 2315 8035 2375 8065
rect 2315 8005 2330 8035
rect 2360 8005 2375 8035
rect 2315 7970 2375 8005
rect 2315 7940 2330 7970
rect 2360 7940 2375 7970
rect 2315 7900 2375 7940
rect 2315 7870 2330 7900
rect 2360 7870 2375 7900
rect 2315 7830 2375 7870
rect 2315 7800 2330 7830
rect 2360 7800 2375 7830
rect 2315 7760 2375 7800
rect 2315 7730 2330 7760
rect 2360 7730 2375 7760
rect 2315 7695 2375 7730
rect 2315 7665 2330 7695
rect 2360 7665 2375 7695
rect 2315 7635 2375 7665
rect 2315 7605 2330 7635
rect 2360 7605 2375 7635
rect 2315 7570 2375 7605
rect 2315 7540 2330 7570
rect 2360 7540 2375 7570
rect 2315 7500 2375 7540
rect 2315 7470 2330 7500
rect 2360 7470 2375 7500
rect 2315 7430 2375 7470
rect 2315 7400 2330 7430
rect 2360 7400 2375 7430
rect 2315 7360 2375 7400
rect 2315 7330 2330 7360
rect 2360 7330 2375 7360
rect 2315 7295 2375 7330
rect 2315 7265 2330 7295
rect 2360 7265 2375 7295
rect 2315 7235 2375 7265
rect 2315 7205 2330 7235
rect 2360 7205 2375 7235
rect 2315 7170 2375 7205
rect 2315 7140 2330 7170
rect 2360 7140 2375 7170
rect 2315 7100 2375 7140
rect 2315 7070 2330 7100
rect 2360 7070 2375 7100
rect 2315 7030 2375 7070
rect 2315 7000 2330 7030
rect 2360 7000 2375 7030
rect 2315 6960 2375 7000
rect 2315 6930 2330 6960
rect 2360 6930 2375 6960
rect 2315 6895 2375 6930
rect 2315 6865 2330 6895
rect 2360 6865 2375 6895
rect 2315 6835 2375 6865
rect 2315 6805 2330 6835
rect 2360 6805 2375 6835
rect 2315 6770 2375 6805
rect 2315 6740 2330 6770
rect 2360 6740 2375 6770
rect 2315 6700 2375 6740
rect 2315 6670 2330 6700
rect 2360 6670 2375 6700
rect 2315 6630 2375 6670
rect 2315 6600 2330 6630
rect 2360 6600 2375 6630
rect 2315 6560 2375 6600
rect 2315 6530 2330 6560
rect 2360 6530 2375 6560
rect 2315 6495 2375 6530
rect 2315 6465 2330 6495
rect 2360 6465 2375 6495
rect 2315 6450 2375 6465
rect 3165 9635 3285 9650
rect 3165 9605 3180 9635
rect 3210 9605 3240 9635
rect 3270 9605 3285 9635
rect 3165 9570 3285 9605
rect 3165 9540 3180 9570
rect 3210 9540 3240 9570
rect 3270 9540 3285 9570
rect 3165 9500 3285 9540
rect 3165 9470 3180 9500
rect 3210 9470 3240 9500
rect 3270 9470 3285 9500
rect 3165 9430 3285 9470
rect 3165 9400 3180 9430
rect 3210 9400 3240 9430
rect 3270 9400 3285 9430
rect 3165 9360 3285 9400
rect 3165 9330 3180 9360
rect 3210 9330 3240 9360
rect 3270 9330 3285 9360
rect 3165 9295 3285 9330
rect 3165 9265 3180 9295
rect 3210 9265 3240 9295
rect 3270 9265 3285 9295
rect 3165 9235 3285 9265
rect 3165 9205 3180 9235
rect 3210 9205 3240 9235
rect 3270 9205 3285 9235
rect 3165 9170 3285 9205
rect 3165 9140 3180 9170
rect 3210 9140 3240 9170
rect 3270 9140 3285 9170
rect 3165 9100 3285 9140
rect 3165 9070 3180 9100
rect 3210 9070 3240 9100
rect 3270 9070 3285 9100
rect 3165 9030 3285 9070
rect 3165 9000 3180 9030
rect 3210 9000 3240 9030
rect 3270 9000 3285 9030
rect 3165 8960 3285 9000
rect 3165 8930 3180 8960
rect 3210 8930 3240 8960
rect 3270 8930 3285 8960
rect 3165 8895 3285 8930
rect 3165 8865 3180 8895
rect 3210 8865 3240 8895
rect 3270 8865 3285 8895
rect 3165 8835 3285 8865
rect 3165 8805 3180 8835
rect 3210 8805 3240 8835
rect 3270 8805 3285 8835
rect 3165 8770 3285 8805
rect 3165 8740 3180 8770
rect 3210 8740 3240 8770
rect 3270 8740 3285 8770
rect 3165 8700 3285 8740
rect 3165 8670 3180 8700
rect 3210 8670 3240 8700
rect 3270 8670 3285 8700
rect 3165 8630 3285 8670
rect 3165 8600 3180 8630
rect 3210 8600 3240 8630
rect 3270 8600 3285 8630
rect 3165 8560 3285 8600
rect 3165 8530 3180 8560
rect 3210 8530 3240 8560
rect 3270 8530 3285 8560
rect 3165 8495 3285 8530
rect 3165 8465 3180 8495
rect 3210 8465 3240 8495
rect 3270 8465 3285 8495
rect 3165 8435 3285 8465
rect 3165 8405 3180 8435
rect 3210 8405 3240 8435
rect 3270 8405 3285 8435
rect 3165 8370 3285 8405
rect 3165 8340 3180 8370
rect 3210 8340 3240 8370
rect 3270 8340 3285 8370
rect 3165 8300 3285 8340
rect 3165 8270 3180 8300
rect 3210 8270 3240 8300
rect 3270 8270 3285 8300
rect 3165 8230 3285 8270
rect 3165 8200 3180 8230
rect 3210 8200 3240 8230
rect 3270 8200 3285 8230
rect 3165 8160 3285 8200
rect 3165 8130 3180 8160
rect 3210 8130 3240 8160
rect 3270 8130 3285 8160
rect 3165 8095 3285 8130
rect 3165 8065 3180 8095
rect 3210 8065 3240 8095
rect 3270 8065 3285 8095
rect 3165 8035 3285 8065
rect 3165 8005 3180 8035
rect 3210 8005 3240 8035
rect 3270 8005 3285 8035
rect 3165 7970 3285 8005
rect 3165 7940 3180 7970
rect 3210 7940 3240 7970
rect 3270 7940 3285 7970
rect 3165 7900 3285 7940
rect 3165 7870 3180 7900
rect 3210 7870 3240 7900
rect 3270 7870 3285 7900
rect 3165 7830 3285 7870
rect 3165 7800 3180 7830
rect 3210 7800 3240 7830
rect 3270 7800 3285 7830
rect 3165 7760 3285 7800
rect 3165 7730 3180 7760
rect 3210 7730 3240 7760
rect 3270 7730 3285 7760
rect 3165 7695 3285 7730
rect 3165 7665 3180 7695
rect 3210 7665 3240 7695
rect 3270 7665 3285 7695
rect 3165 7635 3285 7665
rect 3165 7605 3180 7635
rect 3210 7605 3240 7635
rect 3270 7605 3285 7635
rect 3165 7570 3285 7605
rect 3165 7540 3180 7570
rect 3210 7540 3240 7570
rect 3270 7540 3285 7570
rect 3165 7500 3285 7540
rect 3165 7470 3180 7500
rect 3210 7470 3240 7500
rect 3270 7470 3285 7500
rect 3165 7430 3285 7470
rect 3165 7400 3180 7430
rect 3210 7400 3240 7430
rect 3270 7400 3285 7430
rect 3165 7360 3285 7400
rect 3165 7330 3180 7360
rect 3210 7330 3240 7360
rect 3270 7330 3285 7360
rect 3165 7295 3285 7330
rect 3165 7265 3180 7295
rect 3210 7265 3240 7295
rect 3270 7265 3285 7295
rect 3165 7235 3285 7265
rect 3165 7205 3180 7235
rect 3210 7205 3240 7235
rect 3270 7205 3285 7235
rect 3165 7170 3285 7205
rect 3165 7140 3180 7170
rect 3210 7140 3240 7170
rect 3270 7140 3285 7170
rect 3165 7100 3285 7140
rect 3165 7070 3180 7100
rect 3210 7070 3240 7100
rect 3270 7070 3285 7100
rect 3165 7030 3285 7070
rect 3165 7000 3180 7030
rect 3210 7000 3240 7030
rect 3270 7000 3285 7030
rect 3165 6960 3285 7000
rect 3165 6930 3180 6960
rect 3210 6930 3240 6960
rect 3270 6930 3285 6960
rect 3165 6895 3285 6930
rect 3165 6865 3180 6895
rect 3210 6865 3240 6895
rect 3270 6865 3285 6895
rect 3165 6835 3285 6865
rect 3165 6805 3180 6835
rect 3210 6805 3240 6835
rect 3270 6805 3285 6835
rect 3165 6770 3285 6805
rect 3165 6740 3180 6770
rect 3210 6740 3240 6770
rect 3270 6740 3285 6770
rect 3165 6700 3285 6740
rect 3165 6670 3180 6700
rect 3210 6670 3240 6700
rect 3270 6670 3285 6700
rect 3165 6630 3285 6670
rect 3165 6600 3180 6630
rect 3210 6600 3240 6630
rect 3270 6600 3285 6630
rect 3165 6560 3285 6600
rect 3165 6530 3180 6560
rect 3210 6530 3240 6560
rect 3270 6530 3285 6560
rect 3165 6495 3285 6530
rect 3165 6465 3180 6495
rect 3210 6465 3240 6495
rect 3270 6465 3285 6495
rect 3165 6450 3285 6465
rect 3335 9635 3395 9650
rect 3335 9605 3350 9635
rect 3380 9605 3395 9635
rect 3335 9570 3395 9605
rect 3335 9540 3350 9570
rect 3380 9540 3395 9570
rect 3335 9500 3395 9540
rect 3335 9470 3350 9500
rect 3380 9470 3395 9500
rect 3335 9430 3395 9470
rect 3335 9400 3350 9430
rect 3380 9400 3395 9430
rect 3335 9360 3395 9400
rect 3335 9330 3350 9360
rect 3380 9330 3395 9360
rect 3335 9295 3395 9330
rect 3335 9265 3350 9295
rect 3380 9265 3395 9295
rect 3335 9235 3395 9265
rect 3335 9205 3350 9235
rect 3380 9205 3395 9235
rect 3335 9170 3395 9205
rect 3335 9140 3350 9170
rect 3380 9140 3395 9170
rect 3335 9100 3395 9140
rect 3335 9070 3350 9100
rect 3380 9070 3395 9100
rect 3335 9030 3395 9070
rect 3335 9000 3350 9030
rect 3380 9000 3395 9030
rect 3335 8960 3395 9000
rect 3335 8930 3350 8960
rect 3380 8930 3395 8960
rect 3335 8895 3395 8930
rect 3335 8865 3350 8895
rect 3380 8865 3395 8895
rect 3335 8835 3395 8865
rect 3335 8805 3350 8835
rect 3380 8805 3395 8835
rect 3335 8770 3395 8805
rect 3335 8740 3350 8770
rect 3380 8740 3395 8770
rect 3335 8700 3395 8740
rect 3335 8670 3350 8700
rect 3380 8670 3395 8700
rect 3335 8630 3395 8670
rect 3335 8600 3350 8630
rect 3380 8600 3395 8630
rect 3335 8560 3395 8600
rect 3335 8530 3350 8560
rect 3380 8530 3395 8560
rect 3335 8495 3395 8530
rect 3335 8465 3350 8495
rect 3380 8465 3395 8495
rect 3335 8435 3395 8465
rect 3335 8405 3350 8435
rect 3380 8405 3395 8435
rect 3335 8370 3395 8405
rect 3335 8340 3350 8370
rect 3380 8340 3395 8370
rect 3335 8300 3395 8340
rect 3335 8270 3350 8300
rect 3380 8270 3395 8300
rect 3335 8230 3395 8270
rect 3335 8200 3350 8230
rect 3380 8200 3395 8230
rect 3335 8160 3395 8200
rect 3335 8130 3350 8160
rect 3380 8130 3395 8160
rect 3335 8095 3395 8130
rect 3335 8065 3350 8095
rect 3380 8065 3395 8095
rect 3335 8035 3395 8065
rect 3335 8005 3350 8035
rect 3380 8005 3395 8035
rect 3335 7970 3395 8005
rect 3335 7940 3350 7970
rect 3380 7940 3395 7970
rect 3335 7900 3395 7940
rect 3335 7870 3350 7900
rect 3380 7870 3395 7900
rect 3335 7830 3395 7870
rect 3335 7800 3350 7830
rect 3380 7800 3395 7830
rect 3335 7760 3395 7800
rect 3335 7730 3350 7760
rect 3380 7730 3395 7760
rect 3335 7695 3395 7730
rect 3335 7665 3350 7695
rect 3380 7665 3395 7695
rect 3335 7635 3395 7665
rect 3335 7605 3350 7635
rect 3380 7605 3395 7635
rect 3335 7570 3395 7605
rect 3335 7540 3350 7570
rect 3380 7540 3395 7570
rect 3335 7500 3395 7540
rect 3335 7470 3350 7500
rect 3380 7470 3395 7500
rect 3335 7430 3395 7470
rect 3335 7400 3350 7430
rect 3380 7400 3395 7430
rect 3335 7360 3395 7400
rect 3335 7330 3350 7360
rect 3380 7330 3395 7360
rect 3335 7295 3395 7330
rect 3335 7265 3350 7295
rect 3380 7265 3395 7295
rect 3335 7235 3395 7265
rect 3335 7205 3350 7235
rect 3380 7205 3395 7235
rect 3335 7170 3395 7205
rect 3335 7140 3350 7170
rect 3380 7140 3395 7170
rect 3335 7100 3395 7140
rect 3335 7070 3350 7100
rect 3380 7070 3395 7100
rect 3335 7030 3395 7070
rect 3335 7000 3350 7030
rect 3380 7000 3395 7030
rect 3335 6960 3395 7000
rect 3335 6930 3350 6960
rect 3380 6930 3395 6960
rect 3335 6895 3395 6930
rect 3335 6865 3350 6895
rect 3380 6865 3395 6895
rect 3335 6835 3395 6865
rect 3335 6805 3350 6835
rect 3380 6805 3395 6835
rect 3335 6770 3395 6805
rect 3335 6740 3350 6770
rect 3380 6740 3395 6770
rect 3335 6700 3395 6740
rect 3335 6670 3350 6700
rect 3380 6670 3395 6700
rect 3335 6630 3395 6670
rect 3335 6600 3350 6630
rect 3380 6600 3395 6630
rect 3335 6560 3395 6600
rect 3335 6530 3350 6560
rect 3380 6530 3395 6560
rect 3335 6495 3395 6530
rect 3335 6465 3350 6495
rect 3380 6465 3395 6495
rect 3335 6450 3395 6465
rect 6620 9635 6680 9650
rect 6620 9605 6635 9635
rect 6665 9605 6680 9635
rect 6620 9570 6680 9605
rect 6620 9540 6635 9570
rect 6665 9540 6680 9570
rect 6620 9500 6680 9540
rect 6620 9470 6635 9500
rect 6665 9470 6680 9500
rect 6620 9430 6680 9470
rect 6620 9400 6635 9430
rect 6665 9400 6680 9430
rect 6620 9360 6680 9400
rect 6620 9330 6635 9360
rect 6665 9330 6680 9360
rect 6620 9295 6680 9330
rect 6620 9265 6635 9295
rect 6665 9265 6680 9295
rect 6620 9235 6680 9265
rect 6620 9205 6635 9235
rect 6665 9205 6680 9235
rect 6620 9170 6680 9205
rect 6620 9140 6635 9170
rect 6665 9140 6680 9170
rect 6620 9100 6680 9140
rect 6620 9070 6635 9100
rect 6665 9070 6680 9100
rect 6620 9030 6680 9070
rect 6620 9000 6635 9030
rect 6665 9000 6680 9030
rect 6620 8960 6680 9000
rect 6620 8930 6635 8960
rect 6665 8930 6680 8960
rect 6620 8895 6680 8930
rect 6620 8865 6635 8895
rect 6665 8865 6680 8895
rect 6620 8835 6680 8865
rect 6620 8805 6635 8835
rect 6665 8805 6680 8835
rect 6620 8770 6680 8805
rect 6620 8740 6635 8770
rect 6665 8740 6680 8770
rect 6620 8700 6680 8740
rect 6620 8670 6635 8700
rect 6665 8670 6680 8700
rect 6620 8630 6680 8670
rect 6620 8600 6635 8630
rect 6665 8600 6680 8630
rect 6620 8560 6680 8600
rect 6620 8530 6635 8560
rect 6665 8530 6680 8560
rect 6620 8495 6680 8530
rect 6620 8465 6635 8495
rect 6665 8465 6680 8495
rect 6620 8435 6680 8465
rect 6620 8405 6635 8435
rect 6665 8405 6680 8435
rect 6620 8370 6680 8405
rect 6620 8340 6635 8370
rect 6665 8340 6680 8370
rect 6620 8300 6680 8340
rect 6620 8270 6635 8300
rect 6665 8270 6680 8300
rect 6620 8230 6680 8270
rect 6620 8200 6635 8230
rect 6665 8200 6680 8230
rect 6620 8160 6680 8200
rect 6620 8130 6635 8160
rect 6665 8130 6680 8160
rect 6620 8095 6680 8130
rect 6620 8065 6635 8095
rect 6665 8065 6680 8095
rect 6620 8035 6680 8065
rect 6620 8005 6635 8035
rect 6665 8005 6680 8035
rect 6620 7970 6680 8005
rect 6620 7940 6635 7970
rect 6665 7940 6680 7970
rect 6620 7900 6680 7940
rect 6620 7870 6635 7900
rect 6665 7870 6680 7900
rect 6620 7830 6680 7870
rect 6620 7800 6635 7830
rect 6665 7800 6680 7830
rect 6620 7760 6680 7800
rect 6620 7730 6635 7760
rect 6665 7730 6680 7760
rect 6620 7695 6680 7730
rect 6620 7665 6635 7695
rect 6665 7665 6680 7695
rect 6620 7635 6680 7665
rect 6620 7605 6635 7635
rect 6665 7605 6680 7635
rect 6620 7570 6680 7605
rect 6620 7540 6635 7570
rect 6665 7540 6680 7570
rect 6620 7500 6680 7540
rect 6620 7470 6635 7500
rect 6665 7470 6680 7500
rect 6620 7430 6680 7470
rect 6620 7400 6635 7430
rect 6665 7400 6680 7430
rect 6620 7360 6680 7400
rect 6620 7330 6635 7360
rect 6665 7330 6680 7360
rect 6620 7295 6680 7330
rect 6620 7265 6635 7295
rect 6665 7265 6680 7295
rect 6620 7235 6680 7265
rect 6620 7205 6635 7235
rect 6665 7205 6680 7235
rect 6620 7170 6680 7205
rect 6620 7140 6635 7170
rect 6665 7140 6680 7170
rect 6620 7100 6680 7140
rect 6620 7070 6635 7100
rect 6665 7070 6680 7100
rect 6620 7030 6680 7070
rect 6620 7000 6635 7030
rect 6665 7000 6680 7030
rect 6620 6960 6680 7000
rect 6620 6930 6635 6960
rect 6665 6930 6680 6960
rect 6620 6895 6680 6930
rect 6620 6865 6635 6895
rect 6665 6865 6680 6895
rect 6620 6835 6680 6865
rect 6620 6805 6635 6835
rect 6665 6805 6680 6835
rect 6620 6770 6680 6805
rect 6620 6740 6635 6770
rect 6665 6740 6680 6770
rect 6620 6700 6680 6740
rect 6620 6670 6635 6700
rect 6665 6670 6680 6700
rect 6620 6630 6680 6670
rect 6620 6600 6635 6630
rect 6665 6600 6680 6630
rect 6620 6560 6680 6600
rect 6620 6530 6635 6560
rect 6665 6530 6680 6560
rect 6620 6495 6680 6530
rect 6620 6465 6635 6495
rect 6665 6465 6680 6495
rect 6620 6450 6680 6465
rect 7260 9635 7320 9650
rect 7260 9605 7275 9635
rect 7305 9605 7320 9635
rect 7260 9570 7320 9605
rect 7260 9540 7275 9570
rect 7305 9540 7320 9570
rect 7260 9500 7320 9540
rect 7260 9470 7275 9500
rect 7305 9470 7320 9500
rect 7260 9430 7320 9470
rect 7260 9400 7275 9430
rect 7305 9400 7320 9430
rect 7260 9360 7320 9400
rect 7260 9330 7275 9360
rect 7305 9330 7320 9360
rect 7260 9295 7320 9330
rect 7260 9265 7275 9295
rect 7305 9265 7320 9295
rect 7260 9235 7320 9265
rect 7260 9205 7275 9235
rect 7305 9205 7320 9235
rect 7260 9170 7320 9205
rect 7260 9140 7275 9170
rect 7305 9140 7320 9170
rect 7260 9100 7320 9140
rect 7260 9070 7275 9100
rect 7305 9070 7320 9100
rect 7260 9030 7320 9070
rect 7260 9000 7275 9030
rect 7305 9000 7320 9030
rect 7260 8960 7320 9000
rect 7260 8930 7275 8960
rect 7305 8930 7320 8960
rect 7260 8895 7320 8930
rect 7260 8865 7275 8895
rect 7305 8865 7320 8895
rect 7260 8835 7320 8865
rect 7260 8805 7275 8835
rect 7305 8805 7320 8835
rect 7260 8770 7320 8805
rect 7260 8740 7275 8770
rect 7305 8740 7320 8770
rect 7260 8700 7320 8740
rect 7260 8670 7275 8700
rect 7305 8670 7320 8700
rect 7260 8630 7320 8670
rect 7260 8600 7275 8630
rect 7305 8600 7320 8630
rect 7260 8560 7320 8600
rect 7260 8530 7275 8560
rect 7305 8530 7320 8560
rect 7260 8495 7320 8530
rect 7260 8465 7275 8495
rect 7305 8465 7320 8495
rect 7260 8435 7320 8465
rect 7260 8405 7275 8435
rect 7305 8405 7320 8435
rect 7260 8370 7320 8405
rect 7260 8340 7275 8370
rect 7305 8340 7320 8370
rect 7260 8300 7320 8340
rect 7260 8270 7275 8300
rect 7305 8270 7320 8300
rect 7260 8230 7320 8270
rect 7260 8200 7275 8230
rect 7305 8200 7320 8230
rect 7260 8160 7320 8200
rect 7260 8130 7275 8160
rect 7305 8130 7320 8160
rect 7260 8095 7320 8130
rect 7260 8065 7275 8095
rect 7305 8065 7320 8095
rect 7260 8035 7320 8065
rect 7260 8005 7275 8035
rect 7305 8005 7320 8035
rect 7260 7970 7320 8005
rect 7260 7940 7275 7970
rect 7305 7940 7320 7970
rect 7260 7900 7320 7940
rect 7260 7870 7275 7900
rect 7305 7870 7320 7900
rect 7260 7830 7320 7870
rect 7260 7800 7275 7830
rect 7305 7800 7320 7830
rect 7260 7760 7320 7800
rect 7260 7730 7275 7760
rect 7305 7730 7320 7760
rect 7260 7695 7320 7730
rect 7260 7665 7275 7695
rect 7305 7665 7320 7695
rect 7260 7635 7320 7665
rect 7260 7605 7275 7635
rect 7305 7605 7320 7635
rect 7260 7570 7320 7605
rect 7260 7540 7275 7570
rect 7305 7540 7320 7570
rect 7260 7500 7320 7540
rect 7260 7470 7275 7500
rect 7305 7470 7320 7500
rect 7260 7430 7320 7470
rect 7260 7400 7275 7430
rect 7305 7400 7320 7430
rect 7260 7360 7320 7400
rect 7260 7330 7275 7360
rect 7305 7330 7320 7360
rect 7260 7295 7320 7330
rect 7260 7265 7275 7295
rect 7305 7265 7320 7295
rect 7260 7235 7320 7265
rect 7260 7205 7275 7235
rect 7305 7205 7320 7235
rect 7260 7170 7320 7205
rect 7260 7140 7275 7170
rect 7305 7140 7320 7170
rect 7260 7100 7320 7140
rect 7260 7070 7275 7100
rect 7305 7070 7320 7100
rect 7260 7030 7320 7070
rect 7260 7000 7275 7030
rect 7305 7000 7320 7030
rect 7260 6960 7320 7000
rect 7260 6930 7275 6960
rect 7305 6930 7320 6960
rect 7260 6895 7320 6930
rect 7260 6865 7275 6895
rect 7305 6865 7320 6895
rect 7260 6835 7320 6865
rect 7260 6805 7275 6835
rect 7305 6805 7320 6835
rect 7260 6770 7320 6805
rect 7260 6740 7275 6770
rect 7305 6740 7320 6770
rect 7260 6700 7320 6740
rect 7260 6670 7275 6700
rect 7305 6670 7320 6700
rect 7260 6630 7320 6670
rect 7260 6600 7275 6630
rect 7305 6600 7320 6630
rect 7260 6560 7320 6600
rect 7260 6530 7275 6560
rect 7305 6530 7320 6560
rect 7260 6495 7320 6530
rect 7260 6465 7275 6495
rect 7305 6465 7320 6495
rect 7260 6450 7320 6465
rect 7960 9635 8020 9650
rect 7960 9605 7975 9635
rect 8005 9605 8020 9635
rect 7960 9570 8020 9605
rect 7960 9540 7975 9570
rect 8005 9540 8020 9570
rect 7960 9500 8020 9540
rect 7960 9470 7975 9500
rect 8005 9470 8020 9500
rect 7960 9430 8020 9470
rect 7960 9400 7975 9430
rect 8005 9400 8020 9430
rect 7960 9360 8020 9400
rect 7960 9330 7975 9360
rect 8005 9330 8020 9360
rect 7960 9295 8020 9330
rect 7960 9265 7975 9295
rect 8005 9265 8020 9295
rect 7960 9235 8020 9265
rect 7960 9205 7975 9235
rect 8005 9205 8020 9235
rect 7960 9170 8020 9205
rect 7960 9140 7975 9170
rect 8005 9140 8020 9170
rect 7960 9100 8020 9140
rect 7960 9070 7975 9100
rect 8005 9070 8020 9100
rect 7960 9030 8020 9070
rect 7960 9000 7975 9030
rect 8005 9000 8020 9030
rect 7960 8960 8020 9000
rect 7960 8930 7975 8960
rect 8005 8930 8020 8960
rect 7960 8895 8020 8930
rect 7960 8865 7975 8895
rect 8005 8865 8020 8895
rect 7960 8835 8020 8865
rect 7960 8805 7975 8835
rect 8005 8805 8020 8835
rect 7960 8770 8020 8805
rect 7960 8740 7975 8770
rect 8005 8740 8020 8770
rect 7960 8700 8020 8740
rect 7960 8670 7975 8700
rect 8005 8670 8020 8700
rect 7960 8630 8020 8670
rect 7960 8600 7975 8630
rect 8005 8600 8020 8630
rect 7960 8560 8020 8600
rect 7960 8530 7975 8560
rect 8005 8530 8020 8560
rect 7960 8495 8020 8530
rect 7960 8465 7975 8495
rect 8005 8465 8020 8495
rect 7960 8435 8020 8465
rect 7960 8405 7975 8435
rect 8005 8405 8020 8435
rect 7960 8370 8020 8405
rect 7960 8340 7975 8370
rect 8005 8340 8020 8370
rect 7960 8300 8020 8340
rect 7960 8270 7975 8300
rect 8005 8270 8020 8300
rect 7960 8230 8020 8270
rect 7960 8200 7975 8230
rect 8005 8200 8020 8230
rect 7960 8160 8020 8200
rect 7960 8130 7975 8160
rect 8005 8130 8020 8160
rect 7960 8095 8020 8130
rect 7960 8065 7975 8095
rect 8005 8065 8020 8095
rect 7960 8035 8020 8065
rect 7960 8005 7975 8035
rect 8005 8005 8020 8035
rect 7960 7970 8020 8005
rect 7960 7940 7975 7970
rect 8005 7940 8020 7970
rect 7960 7900 8020 7940
rect 7960 7870 7975 7900
rect 8005 7870 8020 7900
rect 7960 7830 8020 7870
rect 7960 7800 7975 7830
rect 8005 7800 8020 7830
rect 7960 7760 8020 7800
rect 7960 7730 7975 7760
rect 8005 7730 8020 7760
rect 7960 7695 8020 7730
rect 7960 7665 7975 7695
rect 8005 7665 8020 7695
rect 7960 7635 8020 7665
rect 7960 7605 7975 7635
rect 8005 7605 8020 7635
rect 7960 7570 8020 7605
rect 7960 7540 7975 7570
rect 8005 7540 8020 7570
rect 7960 7500 8020 7540
rect 7960 7470 7975 7500
rect 8005 7470 8020 7500
rect 7960 7430 8020 7470
rect 7960 7400 7975 7430
rect 8005 7400 8020 7430
rect 7960 7360 8020 7400
rect 7960 7330 7975 7360
rect 8005 7330 8020 7360
rect 7960 7295 8020 7330
rect 7960 7265 7975 7295
rect 8005 7265 8020 7295
rect 7960 7235 8020 7265
rect 7960 7205 7975 7235
rect 8005 7205 8020 7235
rect 7960 7170 8020 7205
rect 7960 7140 7975 7170
rect 8005 7140 8020 7170
rect 7960 7100 8020 7140
rect 7960 7070 7975 7100
rect 8005 7070 8020 7100
rect 7960 7030 8020 7070
rect 7960 7000 7975 7030
rect 8005 7000 8020 7030
rect 7960 6960 8020 7000
rect 7960 6930 7975 6960
rect 8005 6930 8020 6960
rect 7960 6895 8020 6930
rect 7960 6865 7975 6895
rect 8005 6865 8020 6895
rect 7960 6835 8020 6865
rect 7960 6805 7975 6835
rect 8005 6805 8020 6835
rect 7960 6770 8020 6805
rect 7960 6740 7975 6770
rect 8005 6740 8020 6770
rect 7960 6700 8020 6740
rect 7960 6670 7975 6700
rect 8005 6670 8020 6700
rect 7960 6630 8020 6670
rect 7960 6600 7975 6630
rect 8005 6600 8020 6630
rect 7960 6560 8020 6600
rect 7960 6530 7975 6560
rect 8005 6530 8020 6560
rect 7960 6495 8020 6530
rect 7960 6465 7975 6495
rect 8005 6465 8020 6495
rect 7960 6450 8020 6465
rect 8310 9635 8370 9650
rect 8310 9605 8325 9635
rect 8355 9605 8370 9635
rect 8310 9570 8370 9605
rect 8310 9540 8325 9570
rect 8355 9540 8370 9570
rect 8310 9500 8370 9540
rect 8310 9470 8325 9500
rect 8355 9470 8370 9500
rect 8310 9430 8370 9470
rect 8310 9400 8325 9430
rect 8355 9400 8370 9430
rect 8310 9360 8370 9400
rect 8310 9330 8325 9360
rect 8355 9330 8370 9360
rect 8310 9295 8370 9330
rect 8310 9265 8325 9295
rect 8355 9265 8370 9295
rect 8310 9235 8370 9265
rect 8310 9205 8325 9235
rect 8355 9205 8370 9235
rect 8310 9170 8370 9205
rect 8310 9140 8325 9170
rect 8355 9140 8370 9170
rect 8310 9100 8370 9140
rect 8310 9070 8325 9100
rect 8355 9070 8370 9100
rect 8310 9030 8370 9070
rect 8310 9000 8325 9030
rect 8355 9000 8370 9030
rect 8310 8960 8370 9000
rect 8310 8930 8325 8960
rect 8355 8930 8370 8960
rect 8310 8895 8370 8930
rect 8310 8865 8325 8895
rect 8355 8865 8370 8895
rect 8310 8835 8370 8865
rect 8310 8805 8325 8835
rect 8355 8805 8370 8835
rect 8310 8770 8370 8805
rect 8310 8740 8325 8770
rect 8355 8740 8370 8770
rect 8310 8700 8370 8740
rect 8310 8670 8325 8700
rect 8355 8670 8370 8700
rect 8310 8630 8370 8670
rect 8310 8600 8325 8630
rect 8355 8600 8370 8630
rect 8310 8560 8370 8600
rect 8310 8530 8325 8560
rect 8355 8530 8370 8560
rect 8310 8495 8370 8530
rect 8310 8465 8325 8495
rect 8355 8465 8370 8495
rect 8310 8435 8370 8465
rect 8310 8405 8325 8435
rect 8355 8405 8370 8435
rect 8310 8370 8370 8405
rect 8310 8340 8325 8370
rect 8355 8340 8370 8370
rect 8310 8300 8370 8340
rect 8310 8270 8325 8300
rect 8355 8270 8370 8300
rect 8310 8230 8370 8270
rect 8310 8200 8325 8230
rect 8355 8200 8370 8230
rect 8310 8160 8370 8200
rect 8310 8130 8325 8160
rect 8355 8130 8370 8160
rect 8310 8095 8370 8130
rect 8310 8065 8325 8095
rect 8355 8065 8370 8095
rect 8310 8035 8370 8065
rect 8310 8005 8325 8035
rect 8355 8005 8370 8035
rect 8310 7970 8370 8005
rect 8310 7940 8325 7970
rect 8355 7940 8370 7970
rect 8310 7900 8370 7940
rect 8310 7870 8325 7900
rect 8355 7870 8370 7900
rect 8310 7830 8370 7870
rect 8310 7800 8325 7830
rect 8355 7800 8370 7830
rect 8310 7760 8370 7800
rect 8310 7730 8325 7760
rect 8355 7730 8370 7760
rect 8310 7695 8370 7730
rect 8310 7665 8325 7695
rect 8355 7665 8370 7695
rect 8310 7635 8370 7665
rect 8310 7605 8325 7635
rect 8355 7605 8370 7635
rect 8310 7570 8370 7605
rect 8310 7540 8325 7570
rect 8355 7540 8370 7570
rect 8310 7500 8370 7540
rect 8310 7470 8325 7500
rect 8355 7470 8370 7500
rect 8310 7430 8370 7470
rect 8310 7400 8325 7430
rect 8355 7400 8370 7430
rect 8310 7360 8370 7400
rect 8310 7330 8325 7360
rect 8355 7330 8370 7360
rect 8310 7295 8370 7330
rect 8310 7265 8325 7295
rect 8355 7265 8370 7295
rect 8310 7235 8370 7265
rect 8310 7205 8325 7235
rect 8355 7205 8370 7235
rect 8310 7170 8370 7205
rect 8310 7140 8325 7170
rect 8355 7140 8370 7170
rect 8310 7100 8370 7140
rect 8310 7070 8325 7100
rect 8355 7070 8370 7100
rect 8310 7030 8370 7070
rect 8310 7000 8325 7030
rect 8355 7000 8370 7030
rect 8310 6960 8370 7000
rect 8310 6930 8325 6960
rect 8355 6930 8370 6960
rect 8310 6895 8370 6930
rect 8310 6865 8325 6895
rect 8355 6865 8370 6895
rect 8310 6835 8370 6865
rect 8310 6805 8325 6835
rect 8355 6805 8370 6835
rect 8310 6770 8370 6805
rect 8310 6740 8325 6770
rect 8355 6740 8370 6770
rect 8310 6700 8370 6740
rect 8310 6670 8325 6700
rect 8355 6670 8370 6700
rect 8310 6630 8370 6670
rect 8310 6600 8325 6630
rect 8355 6600 8370 6630
rect 8310 6560 8370 6600
rect 8310 6530 8325 6560
rect 8355 6530 8370 6560
rect 8310 6495 8370 6530
rect 8310 6465 8325 6495
rect 8355 6465 8370 6495
rect 8310 6450 8370 6465
rect 8660 9635 8720 9650
rect 8660 9605 8675 9635
rect 8705 9605 8720 9635
rect 8660 9570 8720 9605
rect 8660 9540 8675 9570
rect 8705 9540 8720 9570
rect 8660 9500 8720 9540
rect 8660 9470 8675 9500
rect 8705 9470 8720 9500
rect 8660 9430 8720 9470
rect 8660 9400 8675 9430
rect 8705 9400 8720 9430
rect 8660 9360 8720 9400
rect 8660 9330 8675 9360
rect 8705 9330 8720 9360
rect 8660 9295 8720 9330
rect 8660 9265 8675 9295
rect 8705 9265 8720 9295
rect 8660 9235 8720 9265
rect 8660 9205 8675 9235
rect 8705 9205 8720 9235
rect 8660 9170 8720 9205
rect 8660 9140 8675 9170
rect 8705 9140 8720 9170
rect 8660 9100 8720 9140
rect 8660 9070 8675 9100
rect 8705 9070 8720 9100
rect 8660 9030 8720 9070
rect 8660 9000 8675 9030
rect 8705 9000 8720 9030
rect 8660 8960 8720 9000
rect 8660 8930 8675 8960
rect 8705 8930 8720 8960
rect 8660 8895 8720 8930
rect 8660 8865 8675 8895
rect 8705 8865 8720 8895
rect 8660 8835 8720 8865
rect 8660 8805 8675 8835
rect 8705 8805 8720 8835
rect 8660 8770 8720 8805
rect 8660 8740 8675 8770
rect 8705 8740 8720 8770
rect 8660 8700 8720 8740
rect 8660 8670 8675 8700
rect 8705 8670 8720 8700
rect 8660 8630 8720 8670
rect 8660 8600 8675 8630
rect 8705 8600 8720 8630
rect 8660 8560 8720 8600
rect 8660 8530 8675 8560
rect 8705 8530 8720 8560
rect 8660 8495 8720 8530
rect 8660 8465 8675 8495
rect 8705 8465 8720 8495
rect 8660 8435 8720 8465
rect 8660 8405 8675 8435
rect 8705 8405 8720 8435
rect 8660 8370 8720 8405
rect 8660 8340 8675 8370
rect 8705 8340 8720 8370
rect 8660 8300 8720 8340
rect 8660 8270 8675 8300
rect 8705 8270 8720 8300
rect 8660 8230 8720 8270
rect 8660 8200 8675 8230
rect 8705 8200 8720 8230
rect 8660 8160 8720 8200
rect 8660 8130 8675 8160
rect 8705 8130 8720 8160
rect 8660 8095 8720 8130
rect 8660 8065 8675 8095
rect 8705 8065 8720 8095
rect 8660 8035 8720 8065
rect 8660 8005 8675 8035
rect 8705 8005 8720 8035
rect 8660 7970 8720 8005
rect 8660 7940 8675 7970
rect 8705 7940 8720 7970
rect 8660 7900 8720 7940
rect 8660 7870 8675 7900
rect 8705 7870 8720 7900
rect 8660 7830 8720 7870
rect 8660 7800 8675 7830
rect 8705 7800 8720 7830
rect 8660 7760 8720 7800
rect 8660 7730 8675 7760
rect 8705 7730 8720 7760
rect 8660 7695 8720 7730
rect 8660 7665 8675 7695
rect 8705 7665 8720 7695
rect 8660 7635 8720 7665
rect 8660 7605 8675 7635
rect 8705 7605 8720 7635
rect 8660 7570 8720 7605
rect 8660 7540 8675 7570
rect 8705 7540 8720 7570
rect 8660 7500 8720 7540
rect 8660 7470 8675 7500
rect 8705 7470 8720 7500
rect 8660 7430 8720 7470
rect 8660 7400 8675 7430
rect 8705 7400 8720 7430
rect 8660 7360 8720 7400
rect 8660 7330 8675 7360
rect 8705 7330 8720 7360
rect 8660 7295 8720 7330
rect 8660 7265 8675 7295
rect 8705 7265 8720 7295
rect 8660 7235 8720 7265
rect 8660 7205 8675 7235
rect 8705 7205 8720 7235
rect 8660 7170 8720 7205
rect 8660 7140 8675 7170
rect 8705 7140 8720 7170
rect 8660 7100 8720 7140
rect 8660 7070 8675 7100
rect 8705 7070 8720 7100
rect 8660 7030 8720 7070
rect 8660 7000 8675 7030
rect 8705 7000 8720 7030
rect 8660 6960 8720 7000
rect 8660 6930 8675 6960
rect 8705 6930 8720 6960
rect 8660 6895 8720 6930
rect 8660 6865 8675 6895
rect 8705 6865 8720 6895
rect 8660 6835 8720 6865
rect 8660 6805 8675 6835
rect 8705 6805 8720 6835
rect 8660 6770 8720 6805
rect 8660 6740 8675 6770
rect 8705 6740 8720 6770
rect 8660 6700 8720 6740
rect 8660 6670 8675 6700
rect 8705 6670 8720 6700
rect 8660 6630 8720 6670
rect 8660 6600 8675 6630
rect 8705 6600 8720 6630
rect 8660 6560 8720 6600
rect 8660 6530 8675 6560
rect 8705 6530 8720 6560
rect 8660 6495 8720 6530
rect 8660 6465 8675 6495
rect 8705 6465 8720 6495
rect 8660 6450 8720 6465
rect 9010 9635 9070 9650
rect 9010 9605 9025 9635
rect 9055 9605 9070 9635
rect 9010 9570 9070 9605
rect 9010 9540 9025 9570
rect 9055 9540 9070 9570
rect 9010 9500 9070 9540
rect 9010 9470 9025 9500
rect 9055 9470 9070 9500
rect 9010 9430 9070 9470
rect 9010 9400 9025 9430
rect 9055 9400 9070 9430
rect 9010 9360 9070 9400
rect 9010 9330 9025 9360
rect 9055 9330 9070 9360
rect 9010 9295 9070 9330
rect 9010 9265 9025 9295
rect 9055 9265 9070 9295
rect 9010 9235 9070 9265
rect 9010 9205 9025 9235
rect 9055 9205 9070 9235
rect 9010 9170 9070 9205
rect 9010 9140 9025 9170
rect 9055 9140 9070 9170
rect 9010 9100 9070 9140
rect 9010 9070 9025 9100
rect 9055 9070 9070 9100
rect 9010 9030 9070 9070
rect 9010 9000 9025 9030
rect 9055 9000 9070 9030
rect 9010 8960 9070 9000
rect 9010 8930 9025 8960
rect 9055 8930 9070 8960
rect 9010 8895 9070 8930
rect 9010 8865 9025 8895
rect 9055 8865 9070 8895
rect 9010 8835 9070 8865
rect 9010 8805 9025 8835
rect 9055 8805 9070 8835
rect 9010 8770 9070 8805
rect 9010 8740 9025 8770
rect 9055 8740 9070 8770
rect 9010 8700 9070 8740
rect 9010 8670 9025 8700
rect 9055 8670 9070 8700
rect 9010 8630 9070 8670
rect 9010 8600 9025 8630
rect 9055 8600 9070 8630
rect 9010 8560 9070 8600
rect 9010 8530 9025 8560
rect 9055 8530 9070 8560
rect 9010 8495 9070 8530
rect 9010 8465 9025 8495
rect 9055 8465 9070 8495
rect 9010 8435 9070 8465
rect 9010 8405 9025 8435
rect 9055 8405 9070 8435
rect 9010 8370 9070 8405
rect 9010 8340 9025 8370
rect 9055 8340 9070 8370
rect 9010 8300 9070 8340
rect 9010 8270 9025 8300
rect 9055 8270 9070 8300
rect 9010 8230 9070 8270
rect 9010 8200 9025 8230
rect 9055 8200 9070 8230
rect 9010 8160 9070 8200
rect 9010 8130 9025 8160
rect 9055 8130 9070 8160
rect 9010 8095 9070 8130
rect 9010 8065 9025 8095
rect 9055 8065 9070 8095
rect 9010 8035 9070 8065
rect 9010 8005 9025 8035
rect 9055 8005 9070 8035
rect 9010 7970 9070 8005
rect 9010 7940 9025 7970
rect 9055 7940 9070 7970
rect 9010 7900 9070 7940
rect 9010 7870 9025 7900
rect 9055 7870 9070 7900
rect 9010 7830 9070 7870
rect 9010 7800 9025 7830
rect 9055 7800 9070 7830
rect 9010 7760 9070 7800
rect 9010 7730 9025 7760
rect 9055 7730 9070 7760
rect 9010 7695 9070 7730
rect 9010 7665 9025 7695
rect 9055 7665 9070 7695
rect 9010 7635 9070 7665
rect 9010 7605 9025 7635
rect 9055 7605 9070 7635
rect 9010 7570 9070 7605
rect 9010 7540 9025 7570
rect 9055 7540 9070 7570
rect 9010 7500 9070 7540
rect 9010 7470 9025 7500
rect 9055 7470 9070 7500
rect 9010 7430 9070 7470
rect 9010 7400 9025 7430
rect 9055 7400 9070 7430
rect 9010 7360 9070 7400
rect 9010 7330 9025 7360
rect 9055 7330 9070 7360
rect 9010 7295 9070 7330
rect 9010 7265 9025 7295
rect 9055 7265 9070 7295
rect 9010 7235 9070 7265
rect 9010 7205 9025 7235
rect 9055 7205 9070 7235
rect 9010 7170 9070 7205
rect 9010 7140 9025 7170
rect 9055 7140 9070 7170
rect 9010 7100 9070 7140
rect 9010 7070 9025 7100
rect 9055 7070 9070 7100
rect 9010 7030 9070 7070
rect 9010 7000 9025 7030
rect 9055 7000 9070 7030
rect 9010 6960 9070 7000
rect 9010 6930 9025 6960
rect 9055 6930 9070 6960
rect 9010 6895 9070 6930
rect 9010 6865 9025 6895
rect 9055 6865 9070 6895
rect 9010 6835 9070 6865
rect 9010 6805 9025 6835
rect 9055 6805 9070 6835
rect 9010 6770 9070 6805
rect 9010 6740 9025 6770
rect 9055 6740 9070 6770
rect 9010 6700 9070 6740
rect 9010 6670 9025 6700
rect 9055 6670 9070 6700
rect 9010 6630 9070 6670
rect 9010 6600 9025 6630
rect 9055 6600 9070 6630
rect 9010 6560 9070 6600
rect 9010 6530 9025 6560
rect 9055 6530 9070 6560
rect 9010 6495 9070 6530
rect 9010 6465 9025 6495
rect 9055 6465 9070 6495
rect 9010 6450 9070 6465
rect 2045 6430 2515 6435
rect 2045 6400 2050 6430
rect 2080 6400 2480 6430
rect 2510 6400 2515 6430
rect 2045 6395 2515 6400
rect 2845 6430 2885 6435
rect 2845 6400 2850 6430
rect 2880 6425 2885 6430
rect 3390 6430 3430 6435
rect 3390 6425 3395 6430
rect 2880 6405 3395 6425
rect 2880 6400 2885 6405
rect 2845 6395 2885 6400
rect 3390 6400 3395 6405
rect 3425 6400 3430 6430
rect 3390 6395 3430 6400
rect 5490 6430 5530 6435
rect 5490 6400 5495 6430
rect 5525 6425 5530 6430
rect 6145 6430 6185 6435
rect 6145 6425 6150 6430
rect 5525 6405 6150 6425
rect 5525 6400 5530 6405
rect 5490 6395 5530 6400
rect 6145 6400 6150 6405
rect 6180 6400 6185 6430
rect 6145 6395 6185 6400
rect 6465 6430 6935 6435
rect 6465 6400 6470 6430
rect 6500 6400 6900 6430
rect 6930 6400 6935 6430
rect 6465 6395 6935 6400
rect 2000 6375 2040 6380
rect 2000 6345 2005 6375
rect 2035 6370 2040 6375
rect 3630 6375 3670 6380
rect 3630 6370 3635 6375
rect 2035 6350 3635 6370
rect 2035 6345 2040 6350
rect 2000 6340 2040 6345
rect 3630 6345 3635 6350
rect 3665 6345 3670 6375
rect 3630 6340 3670 6345
rect 5310 6375 5350 6380
rect 5310 6345 5315 6375
rect 5345 6370 5350 6375
rect 6940 6375 6980 6380
rect 6940 6370 6945 6375
rect 5345 6350 6945 6370
rect 5345 6345 5350 6350
rect 5310 6340 5350 6345
rect 6940 6345 6945 6350
rect 6975 6345 6980 6375
rect 6940 6340 6980 6345
rect 2715 6330 2755 6335
rect 2715 6300 2720 6330
rect 2750 6325 2755 6330
rect 4850 6330 4890 6335
rect 4850 6325 4855 6330
rect 2750 6305 4855 6325
rect 2750 6300 2755 6305
rect 2715 6295 2755 6300
rect 4850 6300 4855 6305
rect 4885 6300 4890 6330
rect 4850 6295 4890 6300
rect 2990 6275 3030 6280
rect 2990 6245 2995 6275
rect 3025 6270 3030 6275
rect 5545 6275 5585 6280
rect 5545 6270 5550 6275
rect 3025 6250 5550 6270
rect 3025 6245 3030 6250
rect 2990 6240 3030 6245
rect 5545 6245 5550 6250
rect 5580 6245 5585 6275
rect 5545 6240 5585 6245
rect 1280 6205 7700 6210
rect 1280 6175 1285 6205
rect 1315 6175 1325 6205
rect 1355 6175 1365 6205
rect 1395 6175 4310 6205
rect 4340 6175 4420 6205
rect 4450 6175 4530 6205
rect 4560 6175 4640 6205
rect 4670 6175 7585 6205
rect 7615 6175 7625 6205
rect 7655 6175 7665 6205
rect 7695 6175 7700 6205
rect 1280 6165 7700 6175
rect 1280 6135 1285 6165
rect 1315 6135 1325 6165
rect 1355 6135 1365 6165
rect 1395 6135 4310 6165
rect 4340 6135 4420 6165
rect 4450 6135 4530 6165
rect 4560 6135 4640 6165
rect 4670 6135 7585 6165
rect 7615 6135 7625 6165
rect 7655 6135 7665 6165
rect 7695 6135 7700 6165
rect 1280 6125 7700 6135
rect 1280 6095 1285 6125
rect 1315 6095 1325 6125
rect 1355 6095 1365 6125
rect 1395 6095 4310 6125
rect 4340 6095 4420 6125
rect 4450 6095 4530 6125
rect 4560 6095 4640 6125
rect 4670 6095 7585 6125
rect 7615 6095 7625 6125
rect 7655 6095 7665 6125
rect 7695 6095 7700 6125
rect 1280 6090 7700 6095
rect 5870 5085 5910 5090
rect 4850 5065 4890 5070
rect 4940 5065 4980 5070
rect 4850 5035 4855 5065
rect 4885 5040 4945 5065
rect 4885 5035 4890 5040
rect 4850 5030 4890 5035
rect 4940 5035 4945 5040
rect 4975 5035 4980 5065
rect 5870 5055 5875 5085
rect 5905 5080 5910 5085
rect 6220 5085 6260 5090
rect 6220 5080 6225 5085
rect 5905 5060 6225 5080
rect 5905 5055 5910 5060
rect 5870 5050 5910 5055
rect 6220 5055 6225 5060
rect 6255 5055 6260 5085
rect 6220 5050 6260 5055
rect 4940 5030 4980 5035
rect 5870 4580 5910 4585
rect 5870 4575 5875 4580
rect 5195 4555 5875 4575
rect 5870 4550 5875 4555
rect 5905 4550 5910 4580
rect 5870 4545 5910 4550
rect 4940 4500 4980 4505
rect 4940 4470 4945 4500
rect 4975 4470 4980 4500
rect 4940 4465 4980 4470
rect 5490 3000 5530 3005
rect 5490 2995 5495 3000
rect 4720 2975 5495 2995
rect 5490 2970 5495 2975
rect 5525 2970 5530 3000
rect 5490 2965 5530 2970
rect 5320 2945 5350 2950
rect 3390 2930 3430 2935
rect 3390 2900 3395 2930
rect 3425 2925 3430 2930
rect 3425 2905 3955 2925
rect 5545 2945 5585 2950
rect 5545 2940 5550 2945
rect 5350 2920 5550 2940
rect 5320 2910 5350 2915
rect 5545 2915 5550 2920
rect 5580 2915 5585 2945
rect 5545 2910 5585 2915
rect 3425 2900 3430 2905
rect 3390 2895 3430 2900
rect 2045 2005 2085 2010
rect 2045 1975 2050 2005
rect 2080 2000 2085 2005
rect 2200 2005 2240 2010
rect 2200 2000 2205 2005
rect 2080 1980 2205 2000
rect 2080 1975 2085 1980
rect 2045 1970 2085 1975
rect 2200 1975 2205 1980
rect 2235 1975 2240 2005
rect 2200 1970 2240 1975
rect 6740 2005 6780 2010
rect 6740 1975 6745 2005
rect 6775 2000 6780 2005
rect 6895 2005 6935 2010
rect 6895 2000 6900 2005
rect 6775 1980 6900 2000
rect 6775 1975 6780 1980
rect 6740 1970 6780 1975
rect 6895 1975 6900 1980
rect 6930 1975 6935 2005
rect 6895 1970 6935 1975
rect 2000 1950 2040 1955
rect 2000 1920 2005 1950
rect 2035 1945 2040 1950
rect 2155 1950 2195 1955
rect 2155 1945 2160 1950
rect 2035 1925 2160 1945
rect 2035 1920 2040 1925
rect 2000 1915 2040 1920
rect 2155 1920 2160 1925
rect 2190 1920 2195 1950
rect 2155 1915 2195 1920
rect 6785 1950 6825 1955
rect 6785 1920 6790 1950
rect 6820 1945 6825 1950
rect 6940 1950 6980 1955
rect 6940 1945 6945 1950
rect 6820 1925 6945 1945
rect 6820 1920 6825 1925
rect 6785 1915 6825 1920
rect 6940 1920 6945 1925
rect 6975 1920 6980 1950
rect 6940 1915 6980 1920
rect 3605 1370 3625 1390
rect 5355 1370 5375 1390
rect 1280 850 7700 855
rect 1280 820 1285 850
rect 1315 820 1325 850
rect 1355 820 1365 850
rect 1395 820 4420 850
rect 4450 820 4475 850
rect 4505 820 4530 850
rect 4560 820 7585 850
rect 7615 820 7625 850
rect 7655 820 7665 850
rect 7695 820 7700 850
rect 1280 810 7700 820
rect 1280 780 1285 810
rect 1315 780 1325 810
rect 1355 780 1365 810
rect 1395 780 4420 810
rect 4450 780 4475 810
rect 4505 780 4530 810
rect 4560 780 7585 810
rect 7615 780 7625 810
rect 7655 780 7665 810
rect 7695 780 7700 810
rect 1280 770 7700 780
rect 1280 740 1285 770
rect 1315 740 1325 770
rect 1355 740 1365 770
rect 1395 740 4420 770
rect 4450 740 4475 770
rect 4505 740 4530 770
rect 4560 740 7585 770
rect 7615 740 7625 770
rect 7655 740 7665 770
rect 7695 740 7700 770
rect 1280 735 7700 740
rect 1950 455 1970 475
rect 6785 455 6805 475
rect -90 -1305 -30 -1290
rect -90 -1335 -75 -1305
rect -45 -1335 -30 -1305
rect -90 -1370 -30 -1335
rect -90 -1400 -75 -1370
rect -45 -1400 -30 -1370
rect -90 -1440 -30 -1400
rect -90 -1470 -75 -1440
rect -45 -1470 -30 -1440
rect -90 -1510 -30 -1470
rect -90 -1540 -75 -1510
rect -45 -1540 -30 -1510
rect -90 -1580 -30 -1540
rect -90 -1610 -75 -1580
rect -45 -1610 -30 -1580
rect -90 -1645 -30 -1610
rect -90 -1675 -75 -1645
rect -45 -1675 -30 -1645
rect -90 -1705 -30 -1675
rect -90 -1735 -75 -1705
rect -45 -1735 -30 -1705
rect -90 -1770 -30 -1735
rect -90 -1800 -75 -1770
rect -45 -1800 -30 -1770
rect -90 -1840 -30 -1800
rect -90 -1870 -75 -1840
rect -45 -1870 -30 -1840
rect -90 -1910 -30 -1870
rect -90 -1940 -75 -1910
rect -45 -1940 -30 -1910
rect -90 -1980 -30 -1940
rect -90 -2010 -75 -1980
rect -45 -2010 -30 -1980
rect -90 -2045 -30 -2010
rect -90 -2075 -75 -2045
rect -45 -2075 -30 -2045
rect -90 -2105 -30 -2075
rect -90 -2135 -75 -2105
rect -45 -2135 -30 -2105
rect -90 -2170 -30 -2135
rect -90 -2200 -75 -2170
rect -45 -2200 -30 -2170
rect -90 -2240 -30 -2200
rect -90 -2270 -75 -2240
rect -45 -2270 -30 -2240
rect -90 -2310 -30 -2270
rect -90 -2340 -75 -2310
rect -45 -2340 -30 -2310
rect -90 -2380 -30 -2340
rect -90 -2410 -75 -2380
rect -45 -2410 -30 -2380
rect -90 -2445 -30 -2410
rect -90 -2475 -75 -2445
rect -45 -2475 -30 -2445
rect -90 -2505 -30 -2475
rect -90 -2535 -75 -2505
rect -45 -2535 -30 -2505
rect -90 -2570 -30 -2535
rect -90 -2600 -75 -2570
rect -45 -2600 -30 -2570
rect -90 -2640 -30 -2600
rect -90 -2670 -75 -2640
rect -45 -2670 -30 -2640
rect -90 -2710 -30 -2670
rect -90 -2740 -75 -2710
rect -45 -2740 -30 -2710
rect -90 -2780 -30 -2740
rect -90 -2810 -75 -2780
rect -45 -2810 -30 -2780
rect -90 -2845 -30 -2810
rect -90 -2875 -75 -2845
rect -45 -2875 -30 -2845
rect -90 -2905 -30 -2875
rect -90 -2935 -75 -2905
rect -45 -2935 -30 -2905
rect -90 -2970 -30 -2935
rect -90 -3000 -75 -2970
rect -45 -3000 -30 -2970
rect -90 -3040 -30 -3000
rect -90 -3070 -75 -3040
rect -45 -3070 -30 -3040
rect -90 -3110 -30 -3070
rect -90 -3140 -75 -3110
rect -45 -3140 -30 -3110
rect -90 -3180 -30 -3140
rect -90 -3210 -75 -3180
rect -45 -3210 -30 -3180
rect -90 -3245 -30 -3210
rect -90 -3275 -75 -3245
rect -45 -3275 -30 -3245
rect -90 -3305 -30 -3275
rect -90 -3335 -75 -3305
rect -45 -3335 -30 -3305
rect -90 -3370 -30 -3335
rect -90 -3400 -75 -3370
rect -45 -3400 -30 -3370
rect -90 -3440 -30 -3400
rect -90 -3470 -75 -3440
rect -45 -3470 -30 -3440
rect -90 -3510 -30 -3470
rect -90 -3540 -75 -3510
rect -45 -3540 -30 -3510
rect -90 -3580 -30 -3540
rect -90 -3610 -75 -3580
rect -45 -3610 -30 -3580
rect -90 -3645 -30 -3610
rect -90 -3675 -75 -3645
rect -45 -3675 -30 -3645
rect -90 -3705 -30 -3675
rect -90 -3735 -75 -3705
rect -45 -3735 -30 -3705
rect -90 -3770 -30 -3735
rect -90 -3800 -75 -3770
rect -45 -3800 -30 -3770
rect -90 -3840 -30 -3800
rect -90 -3870 -75 -3840
rect -45 -3870 -30 -3840
rect -90 -3910 -30 -3870
rect -90 -3940 -75 -3910
rect -45 -3940 -30 -3910
rect -90 -3980 -30 -3940
rect -90 -4010 -75 -3980
rect -45 -4010 -30 -3980
rect -90 -4045 -30 -4010
rect -90 -4075 -75 -4045
rect -45 -4075 -30 -4045
rect -90 -4105 -30 -4075
rect -90 -4135 -75 -4105
rect -45 -4135 -30 -4105
rect -90 -4170 -30 -4135
rect -90 -4200 -75 -4170
rect -45 -4200 -30 -4170
rect -90 -4240 -30 -4200
rect -90 -4270 -75 -4240
rect -45 -4270 -30 -4240
rect -90 -4310 -30 -4270
rect -90 -4340 -75 -4310
rect -45 -4340 -30 -4310
rect -90 -4380 -30 -4340
rect -90 -4410 -75 -4380
rect -45 -4410 -30 -4380
rect -90 -4445 -30 -4410
rect -90 -4475 -75 -4445
rect -45 -4475 -30 -4445
rect -90 -4490 -30 -4475
rect 260 -1305 320 -1290
rect 260 -1335 275 -1305
rect 305 -1335 320 -1305
rect 260 -1370 320 -1335
rect 260 -1400 275 -1370
rect 305 -1400 320 -1370
rect 260 -1440 320 -1400
rect 260 -1470 275 -1440
rect 305 -1470 320 -1440
rect 260 -1510 320 -1470
rect 260 -1540 275 -1510
rect 305 -1540 320 -1510
rect 260 -1580 320 -1540
rect 260 -1610 275 -1580
rect 305 -1610 320 -1580
rect 260 -1645 320 -1610
rect 260 -1675 275 -1645
rect 305 -1675 320 -1645
rect 260 -1705 320 -1675
rect 260 -1735 275 -1705
rect 305 -1735 320 -1705
rect 260 -1770 320 -1735
rect 260 -1800 275 -1770
rect 305 -1800 320 -1770
rect 260 -1840 320 -1800
rect 260 -1870 275 -1840
rect 305 -1870 320 -1840
rect 260 -1910 320 -1870
rect 260 -1940 275 -1910
rect 305 -1940 320 -1910
rect 260 -1980 320 -1940
rect 260 -2010 275 -1980
rect 305 -2010 320 -1980
rect 260 -2045 320 -2010
rect 260 -2075 275 -2045
rect 305 -2075 320 -2045
rect 260 -2105 320 -2075
rect 260 -2135 275 -2105
rect 305 -2135 320 -2105
rect 260 -2170 320 -2135
rect 260 -2200 275 -2170
rect 305 -2200 320 -2170
rect 260 -2240 320 -2200
rect 260 -2270 275 -2240
rect 305 -2270 320 -2240
rect 260 -2310 320 -2270
rect 260 -2340 275 -2310
rect 305 -2340 320 -2310
rect 260 -2380 320 -2340
rect 260 -2410 275 -2380
rect 305 -2410 320 -2380
rect 260 -2445 320 -2410
rect 260 -2475 275 -2445
rect 305 -2475 320 -2445
rect 260 -2505 320 -2475
rect 260 -2535 275 -2505
rect 305 -2535 320 -2505
rect 260 -2570 320 -2535
rect 260 -2600 275 -2570
rect 305 -2600 320 -2570
rect 260 -2640 320 -2600
rect 260 -2670 275 -2640
rect 305 -2670 320 -2640
rect 260 -2710 320 -2670
rect 260 -2740 275 -2710
rect 305 -2740 320 -2710
rect 260 -2780 320 -2740
rect 260 -2810 275 -2780
rect 305 -2810 320 -2780
rect 260 -2845 320 -2810
rect 260 -2875 275 -2845
rect 305 -2875 320 -2845
rect 260 -2905 320 -2875
rect 260 -2935 275 -2905
rect 305 -2935 320 -2905
rect 260 -2970 320 -2935
rect 260 -3000 275 -2970
rect 305 -3000 320 -2970
rect 260 -3040 320 -3000
rect 260 -3070 275 -3040
rect 305 -3070 320 -3040
rect 260 -3110 320 -3070
rect 260 -3140 275 -3110
rect 305 -3140 320 -3110
rect 260 -3180 320 -3140
rect 260 -3210 275 -3180
rect 305 -3210 320 -3180
rect 260 -3245 320 -3210
rect 260 -3275 275 -3245
rect 305 -3275 320 -3245
rect 260 -3305 320 -3275
rect 260 -3335 275 -3305
rect 305 -3335 320 -3305
rect 260 -3370 320 -3335
rect 260 -3400 275 -3370
rect 305 -3400 320 -3370
rect 260 -3440 320 -3400
rect 260 -3470 275 -3440
rect 305 -3470 320 -3440
rect 260 -3510 320 -3470
rect 260 -3540 275 -3510
rect 305 -3540 320 -3510
rect 260 -3580 320 -3540
rect 260 -3610 275 -3580
rect 305 -3610 320 -3580
rect 260 -3645 320 -3610
rect 260 -3675 275 -3645
rect 305 -3675 320 -3645
rect 260 -3705 320 -3675
rect 260 -3735 275 -3705
rect 305 -3735 320 -3705
rect 260 -3770 320 -3735
rect 260 -3800 275 -3770
rect 305 -3800 320 -3770
rect 260 -3840 320 -3800
rect 260 -3870 275 -3840
rect 305 -3870 320 -3840
rect 260 -3910 320 -3870
rect 260 -3940 275 -3910
rect 305 -3940 320 -3910
rect 260 -3980 320 -3940
rect 260 -4010 275 -3980
rect 305 -4010 320 -3980
rect 260 -4045 320 -4010
rect 260 -4075 275 -4045
rect 305 -4075 320 -4045
rect 260 -4105 320 -4075
rect 260 -4135 275 -4105
rect 305 -4135 320 -4105
rect 260 -4170 320 -4135
rect 260 -4200 275 -4170
rect 305 -4200 320 -4170
rect 260 -4240 320 -4200
rect 260 -4270 275 -4240
rect 305 -4270 320 -4240
rect 260 -4310 320 -4270
rect 260 -4340 275 -4310
rect 305 -4340 320 -4310
rect 260 -4380 320 -4340
rect 260 -4410 275 -4380
rect 305 -4410 320 -4380
rect 260 -4445 320 -4410
rect 260 -4475 275 -4445
rect 305 -4475 320 -4445
rect 260 -4490 320 -4475
rect 610 -1305 670 -1290
rect 610 -1335 625 -1305
rect 655 -1335 670 -1305
rect 610 -1370 670 -1335
rect 610 -1400 625 -1370
rect 655 -1400 670 -1370
rect 610 -1440 670 -1400
rect 610 -1470 625 -1440
rect 655 -1470 670 -1440
rect 610 -1510 670 -1470
rect 610 -1540 625 -1510
rect 655 -1540 670 -1510
rect 610 -1580 670 -1540
rect 610 -1610 625 -1580
rect 655 -1610 670 -1580
rect 610 -1645 670 -1610
rect 610 -1675 625 -1645
rect 655 -1675 670 -1645
rect 610 -1705 670 -1675
rect 610 -1735 625 -1705
rect 655 -1735 670 -1705
rect 610 -1770 670 -1735
rect 610 -1800 625 -1770
rect 655 -1800 670 -1770
rect 610 -1840 670 -1800
rect 610 -1870 625 -1840
rect 655 -1870 670 -1840
rect 610 -1910 670 -1870
rect 610 -1940 625 -1910
rect 655 -1940 670 -1910
rect 610 -1980 670 -1940
rect 610 -2010 625 -1980
rect 655 -2010 670 -1980
rect 610 -2045 670 -2010
rect 610 -2075 625 -2045
rect 655 -2075 670 -2045
rect 610 -2105 670 -2075
rect 610 -2135 625 -2105
rect 655 -2135 670 -2105
rect 610 -2170 670 -2135
rect 610 -2200 625 -2170
rect 655 -2200 670 -2170
rect 610 -2240 670 -2200
rect 610 -2270 625 -2240
rect 655 -2270 670 -2240
rect 610 -2310 670 -2270
rect 610 -2340 625 -2310
rect 655 -2340 670 -2310
rect 610 -2380 670 -2340
rect 610 -2410 625 -2380
rect 655 -2410 670 -2380
rect 610 -2445 670 -2410
rect 610 -2475 625 -2445
rect 655 -2475 670 -2445
rect 610 -2505 670 -2475
rect 610 -2535 625 -2505
rect 655 -2535 670 -2505
rect 610 -2570 670 -2535
rect 610 -2600 625 -2570
rect 655 -2600 670 -2570
rect 610 -2640 670 -2600
rect 610 -2670 625 -2640
rect 655 -2670 670 -2640
rect 610 -2710 670 -2670
rect 610 -2740 625 -2710
rect 655 -2740 670 -2710
rect 610 -2780 670 -2740
rect 610 -2810 625 -2780
rect 655 -2810 670 -2780
rect 610 -2845 670 -2810
rect 610 -2875 625 -2845
rect 655 -2875 670 -2845
rect 610 -2905 670 -2875
rect 610 -2935 625 -2905
rect 655 -2935 670 -2905
rect 610 -2970 670 -2935
rect 610 -3000 625 -2970
rect 655 -3000 670 -2970
rect 610 -3040 670 -3000
rect 610 -3070 625 -3040
rect 655 -3070 670 -3040
rect 610 -3110 670 -3070
rect 610 -3140 625 -3110
rect 655 -3140 670 -3110
rect 610 -3180 670 -3140
rect 610 -3210 625 -3180
rect 655 -3210 670 -3180
rect 610 -3245 670 -3210
rect 610 -3275 625 -3245
rect 655 -3275 670 -3245
rect 610 -3305 670 -3275
rect 610 -3335 625 -3305
rect 655 -3335 670 -3305
rect 610 -3370 670 -3335
rect 610 -3400 625 -3370
rect 655 -3400 670 -3370
rect 610 -3440 670 -3400
rect 610 -3470 625 -3440
rect 655 -3470 670 -3440
rect 610 -3510 670 -3470
rect 610 -3540 625 -3510
rect 655 -3540 670 -3510
rect 610 -3580 670 -3540
rect 610 -3610 625 -3580
rect 655 -3610 670 -3580
rect 610 -3645 670 -3610
rect 610 -3675 625 -3645
rect 655 -3675 670 -3645
rect 610 -3705 670 -3675
rect 610 -3735 625 -3705
rect 655 -3735 670 -3705
rect 610 -3770 670 -3735
rect 610 -3800 625 -3770
rect 655 -3800 670 -3770
rect 610 -3840 670 -3800
rect 610 -3870 625 -3840
rect 655 -3870 670 -3840
rect 610 -3910 670 -3870
rect 610 -3940 625 -3910
rect 655 -3940 670 -3910
rect 610 -3980 670 -3940
rect 610 -4010 625 -3980
rect 655 -4010 670 -3980
rect 610 -4045 670 -4010
rect 610 -4075 625 -4045
rect 655 -4075 670 -4045
rect 610 -4105 670 -4075
rect 610 -4135 625 -4105
rect 655 -4135 670 -4105
rect 610 -4170 670 -4135
rect 610 -4200 625 -4170
rect 655 -4200 670 -4170
rect 610 -4240 670 -4200
rect 610 -4270 625 -4240
rect 655 -4270 670 -4240
rect 610 -4310 670 -4270
rect 610 -4340 625 -4310
rect 655 -4340 670 -4310
rect 610 -4380 670 -4340
rect 610 -4410 625 -4380
rect 655 -4410 670 -4380
rect 610 -4445 670 -4410
rect 610 -4475 625 -4445
rect 655 -4475 670 -4445
rect 610 -4490 670 -4475
rect 960 -1305 1020 -1290
rect 960 -1335 975 -1305
rect 1005 -1335 1020 -1305
rect 960 -1370 1020 -1335
rect 960 -1400 975 -1370
rect 1005 -1400 1020 -1370
rect 960 -1440 1020 -1400
rect 960 -1470 975 -1440
rect 1005 -1470 1020 -1440
rect 960 -1510 1020 -1470
rect 960 -1540 975 -1510
rect 1005 -1540 1020 -1510
rect 960 -1580 1020 -1540
rect 960 -1610 975 -1580
rect 1005 -1610 1020 -1580
rect 960 -1645 1020 -1610
rect 960 -1675 975 -1645
rect 1005 -1675 1020 -1645
rect 960 -1705 1020 -1675
rect 960 -1735 975 -1705
rect 1005 -1735 1020 -1705
rect 960 -1770 1020 -1735
rect 960 -1800 975 -1770
rect 1005 -1800 1020 -1770
rect 960 -1840 1020 -1800
rect 960 -1870 975 -1840
rect 1005 -1870 1020 -1840
rect 960 -1910 1020 -1870
rect 960 -1940 975 -1910
rect 1005 -1940 1020 -1910
rect 960 -1980 1020 -1940
rect 960 -2010 975 -1980
rect 1005 -2010 1020 -1980
rect 960 -2045 1020 -2010
rect 960 -2075 975 -2045
rect 1005 -2075 1020 -2045
rect 960 -2105 1020 -2075
rect 960 -2135 975 -2105
rect 1005 -2135 1020 -2105
rect 960 -2170 1020 -2135
rect 960 -2200 975 -2170
rect 1005 -2200 1020 -2170
rect 960 -2240 1020 -2200
rect 960 -2270 975 -2240
rect 1005 -2270 1020 -2240
rect 960 -2310 1020 -2270
rect 960 -2340 975 -2310
rect 1005 -2340 1020 -2310
rect 960 -2380 1020 -2340
rect 960 -2410 975 -2380
rect 1005 -2410 1020 -2380
rect 960 -2445 1020 -2410
rect 960 -2475 975 -2445
rect 1005 -2475 1020 -2445
rect 960 -2505 1020 -2475
rect 960 -2535 975 -2505
rect 1005 -2535 1020 -2505
rect 960 -2570 1020 -2535
rect 960 -2600 975 -2570
rect 1005 -2600 1020 -2570
rect 960 -2640 1020 -2600
rect 960 -2670 975 -2640
rect 1005 -2670 1020 -2640
rect 960 -2710 1020 -2670
rect 960 -2740 975 -2710
rect 1005 -2740 1020 -2710
rect 960 -2780 1020 -2740
rect 960 -2810 975 -2780
rect 1005 -2810 1020 -2780
rect 960 -2845 1020 -2810
rect 960 -2875 975 -2845
rect 1005 -2875 1020 -2845
rect 960 -2905 1020 -2875
rect 960 -2935 975 -2905
rect 1005 -2935 1020 -2905
rect 960 -2970 1020 -2935
rect 960 -3000 975 -2970
rect 1005 -3000 1020 -2970
rect 960 -3040 1020 -3000
rect 960 -3070 975 -3040
rect 1005 -3070 1020 -3040
rect 960 -3110 1020 -3070
rect 960 -3140 975 -3110
rect 1005 -3140 1020 -3110
rect 960 -3180 1020 -3140
rect 960 -3210 975 -3180
rect 1005 -3210 1020 -3180
rect 960 -3245 1020 -3210
rect 960 -3275 975 -3245
rect 1005 -3275 1020 -3245
rect 960 -3305 1020 -3275
rect 960 -3335 975 -3305
rect 1005 -3335 1020 -3305
rect 960 -3370 1020 -3335
rect 960 -3400 975 -3370
rect 1005 -3400 1020 -3370
rect 960 -3440 1020 -3400
rect 960 -3470 975 -3440
rect 1005 -3470 1020 -3440
rect 960 -3510 1020 -3470
rect 960 -3540 975 -3510
rect 1005 -3540 1020 -3510
rect 960 -3580 1020 -3540
rect 960 -3610 975 -3580
rect 1005 -3610 1020 -3580
rect 960 -3645 1020 -3610
rect 960 -3675 975 -3645
rect 1005 -3675 1020 -3645
rect 960 -3705 1020 -3675
rect 960 -3735 975 -3705
rect 1005 -3735 1020 -3705
rect 960 -3770 1020 -3735
rect 960 -3800 975 -3770
rect 1005 -3800 1020 -3770
rect 960 -3840 1020 -3800
rect 960 -3870 975 -3840
rect 1005 -3870 1020 -3840
rect 960 -3910 1020 -3870
rect 960 -3940 975 -3910
rect 1005 -3940 1020 -3910
rect 960 -3980 1020 -3940
rect 960 -4010 975 -3980
rect 1005 -4010 1020 -3980
rect 960 -4045 1020 -4010
rect 960 -4075 975 -4045
rect 1005 -4075 1020 -4045
rect 960 -4105 1020 -4075
rect 960 -4135 975 -4105
rect 1005 -4135 1020 -4105
rect 960 -4170 1020 -4135
rect 960 -4200 975 -4170
rect 1005 -4200 1020 -4170
rect 960 -4240 1020 -4200
rect 960 -4270 975 -4240
rect 1005 -4270 1020 -4240
rect 960 -4310 1020 -4270
rect 960 -4340 975 -4310
rect 1005 -4340 1020 -4310
rect 960 -4380 1020 -4340
rect 960 -4410 975 -4380
rect 1005 -4410 1020 -4380
rect 960 -4445 1020 -4410
rect 960 -4475 975 -4445
rect 1005 -4475 1020 -4445
rect 960 -4490 1020 -4475
rect 1310 -1305 1370 -1290
rect 1310 -1335 1325 -1305
rect 1355 -1335 1370 -1305
rect 1310 -1370 1370 -1335
rect 1310 -1400 1325 -1370
rect 1355 -1400 1370 -1370
rect 1310 -1440 1370 -1400
rect 1310 -1470 1325 -1440
rect 1355 -1470 1370 -1440
rect 1310 -1510 1370 -1470
rect 1310 -1540 1325 -1510
rect 1355 -1540 1370 -1510
rect 1310 -1580 1370 -1540
rect 1310 -1610 1325 -1580
rect 1355 -1610 1370 -1580
rect 1310 -1645 1370 -1610
rect 1310 -1675 1325 -1645
rect 1355 -1675 1370 -1645
rect 1310 -1705 1370 -1675
rect 1310 -1735 1325 -1705
rect 1355 -1735 1370 -1705
rect 1310 -1770 1370 -1735
rect 1310 -1800 1325 -1770
rect 1355 -1800 1370 -1770
rect 1310 -1840 1370 -1800
rect 1310 -1870 1325 -1840
rect 1355 -1870 1370 -1840
rect 1310 -1910 1370 -1870
rect 1310 -1940 1325 -1910
rect 1355 -1940 1370 -1910
rect 1310 -1980 1370 -1940
rect 1310 -2010 1325 -1980
rect 1355 -2010 1370 -1980
rect 1310 -2045 1370 -2010
rect 1310 -2075 1325 -2045
rect 1355 -2075 1370 -2045
rect 1310 -2105 1370 -2075
rect 1310 -2135 1325 -2105
rect 1355 -2135 1370 -2105
rect 1310 -2170 1370 -2135
rect 1310 -2200 1325 -2170
rect 1355 -2200 1370 -2170
rect 1310 -2240 1370 -2200
rect 1310 -2270 1325 -2240
rect 1355 -2270 1370 -2240
rect 1310 -2310 1370 -2270
rect 1310 -2340 1325 -2310
rect 1355 -2340 1370 -2310
rect 1310 -2380 1370 -2340
rect 1310 -2410 1325 -2380
rect 1355 -2410 1370 -2380
rect 1310 -2445 1370 -2410
rect 1310 -2475 1325 -2445
rect 1355 -2475 1370 -2445
rect 1310 -2505 1370 -2475
rect 1310 -2535 1325 -2505
rect 1355 -2535 1370 -2505
rect 1310 -2570 1370 -2535
rect 1310 -2600 1325 -2570
rect 1355 -2600 1370 -2570
rect 1310 -2640 1370 -2600
rect 1310 -2670 1325 -2640
rect 1355 -2670 1370 -2640
rect 1310 -2710 1370 -2670
rect 1310 -2740 1325 -2710
rect 1355 -2740 1370 -2710
rect 1310 -2780 1370 -2740
rect 1310 -2810 1325 -2780
rect 1355 -2810 1370 -2780
rect 1310 -2845 1370 -2810
rect 1310 -2875 1325 -2845
rect 1355 -2875 1370 -2845
rect 1310 -2905 1370 -2875
rect 1310 -2935 1325 -2905
rect 1355 -2935 1370 -2905
rect 1310 -2970 1370 -2935
rect 1310 -3000 1325 -2970
rect 1355 -3000 1370 -2970
rect 1310 -3040 1370 -3000
rect 1310 -3070 1325 -3040
rect 1355 -3070 1370 -3040
rect 1310 -3110 1370 -3070
rect 1310 -3140 1325 -3110
rect 1355 -3140 1370 -3110
rect 1310 -3180 1370 -3140
rect 1310 -3210 1325 -3180
rect 1355 -3210 1370 -3180
rect 1310 -3245 1370 -3210
rect 1310 -3275 1325 -3245
rect 1355 -3275 1370 -3245
rect 1310 -3305 1370 -3275
rect 1310 -3335 1325 -3305
rect 1355 -3335 1370 -3305
rect 1310 -3370 1370 -3335
rect 1310 -3400 1325 -3370
rect 1355 -3400 1370 -3370
rect 1310 -3440 1370 -3400
rect 1310 -3470 1325 -3440
rect 1355 -3470 1370 -3440
rect 1310 -3510 1370 -3470
rect 1310 -3540 1325 -3510
rect 1355 -3540 1370 -3510
rect 1310 -3580 1370 -3540
rect 1310 -3610 1325 -3580
rect 1355 -3610 1370 -3580
rect 1310 -3645 1370 -3610
rect 1310 -3675 1325 -3645
rect 1355 -3675 1370 -3645
rect 1310 -3705 1370 -3675
rect 1310 -3735 1325 -3705
rect 1355 -3735 1370 -3705
rect 1310 -3770 1370 -3735
rect 1310 -3800 1325 -3770
rect 1355 -3800 1370 -3770
rect 1310 -3840 1370 -3800
rect 1310 -3870 1325 -3840
rect 1355 -3870 1370 -3840
rect 1310 -3910 1370 -3870
rect 1310 -3940 1325 -3910
rect 1355 -3940 1370 -3910
rect 1310 -3980 1370 -3940
rect 1310 -4010 1325 -3980
rect 1355 -4010 1370 -3980
rect 1310 -4045 1370 -4010
rect 1310 -4075 1325 -4045
rect 1355 -4075 1370 -4045
rect 1310 -4105 1370 -4075
rect 1310 -4135 1325 -4105
rect 1355 -4135 1370 -4105
rect 1310 -4170 1370 -4135
rect 1310 -4200 1325 -4170
rect 1355 -4200 1370 -4170
rect 1310 -4240 1370 -4200
rect 1310 -4270 1325 -4240
rect 1355 -4270 1370 -4240
rect 1310 -4310 1370 -4270
rect 1310 -4340 1325 -4310
rect 1355 -4340 1370 -4310
rect 1310 -4380 1370 -4340
rect 1310 -4410 1325 -4380
rect 1355 -4410 1370 -4380
rect 1310 -4445 1370 -4410
rect 1310 -4475 1325 -4445
rect 1355 -4475 1370 -4445
rect 1310 -4490 1370 -4475
rect 1660 -1305 1720 -1290
rect 1660 -1335 1675 -1305
rect 1705 -1335 1720 -1305
rect 1660 -1370 1720 -1335
rect 1660 -1400 1675 -1370
rect 1705 -1400 1720 -1370
rect 1660 -1440 1720 -1400
rect 1660 -1470 1675 -1440
rect 1705 -1470 1720 -1440
rect 1660 -1510 1720 -1470
rect 1660 -1540 1675 -1510
rect 1705 -1540 1720 -1510
rect 1660 -1580 1720 -1540
rect 1660 -1610 1675 -1580
rect 1705 -1610 1720 -1580
rect 1660 -1645 1720 -1610
rect 1660 -1675 1675 -1645
rect 1705 -1675 1720 -1645
rect 1660 -1705 1720 -1675
rect 1660 -1735 1675 -1705
rect 1705 -1735 1720 -1705
rect 1660 -1770 1720 -1735
rect 1660 -1800 1675 -1770
rect 1705 -1800 1720 -1770
rect 1660 -1840 1720 -1800
rect 1660 -1870 1675 -1840
rect 1705 -1870 1720 -1840
rect 1660 -1910 1720 -1870
rect 1660 -1940 1675 -1910
rect 1705 -1940 1720 -1910
rect 1660 -1980 1720 -1940
rect 1660 -2010 1675 -1980
rect 1705 -2010 1720 -1980
rect 1660 -2045 1720 -2010
rect 1660 -2075 1675 -2045
rect 1705 -2075 1720 -2045
rect 1660 -2105 1720 -2075
rect 1660 -2135 1675 -2105
rect 1705 -2135 1720 -2105
rect 1660 -2170 1720 -2135
rect 1660 -2200 1675 -2170
rect 1705 -2200 1720 -2170
rect 1660 -2240 1720 -2200
rect 1660 -2270 1675 -2240
rect 1705 -2270 1720 -2240
rect 1660 -2310 1720 -2270
rect 1660 -2340 1675 -2310
rect 1705 -2340 1720 -2310
rect 1660 -2380 1720 -2340
rect 1660 -2410 1675 -2380
rect 1705 -2410 1720 -2380
rect 1660 -2445 1720 -2410
rect 1660 -2475 1675 -2445
rect 1705 -2475 1720 -2445
rect 1660 -2505 1720 -2475
rect 1660 -2535 1675 -2505
rect 1705 -2535 1720 -2505
rect 1660 -2570 1720 -2535
rect 1660 -2600 1675 -2570
rect 1705 -2600 1720 -2570
rect 1660 -2640 1720 -2600
rect 1660 -2670 1675 -2640
rect 1705 -2670 1720 -2640
rect 1660 -2710 1720 -2670
rect 1660 -2740 1675 -2710
rect 1705 -2740 1720 -2710
rect 1660 -2780 1720 -2740
rect 1660 -2810 1675 -2780
rect 1705 -2810 1720 -2780
rect 1660 -2845 1720 -2810
rect 1660 -2875 1675 -2845
rect 1705 -2875 1720 -2845
rect 1660 -2905 1720 -2875
rect 1660 -2935 1675 -2905
rect 1705 -2935 1720 -2905
rect 1660 -2970 1720 -2935
rect 1660 -3000 1675 -2970
rect 1705 -3000 1720 -2970
rect 1660 -3040 1720 -3000
rect 1660 -3070 1675 -3040
rect 1705 -3070 1720 -3040
rect 1660 -3110 1720 -3070
rect 1660 -3140 1675 -3110
rect 1705 -3140 1720 -3110
rect 1660 -3180 1720 -3140
rect 1660 -3210 1675 -3180
rect 1705 -3210 1720 -3180
rect 1660 -3245 1720 -3210
rect 1660 -3275 1675 -3245
rect 1705 -3275 1720 -3245
rect 1660 -3305 1720 -3275
rect 1660 -3335 1675 -3305
rect 1705 -3335 1720 -3305
rect 1660 -3370 1720 -3335
rect 1660 -3400 1675 -3370
rect 1705 -3400 1720 -3370
rect 1660 -3440 1720 -3400
rect 1660 -3470 1675 -3440
rect 1705 -3470 1720 -3440
rect 1660 -3510 1720 -3470
rect 1660 -3540 1675 -3510
rect 1705 -3540 1720 -3510
rect 1660 -3580 1720 -3540
rect 1660 -3610 1675 -3580
rect 1705 -3610 1720 -3580
rect 1660 -3645 1720 -3610
rect 1660 -3675 1675 -3645
rect 1705 -3675 1720 -3645
rect 1660 -3705 1720 -3675
rect 1660 -3735 1675 -3705
rect 1705 -3735 1720 -3705
rect 1660 -3770 1720 -3735
rect 1660 -3800 1675 -3770
rect 1705 -3800 1720 -3770
rect 1660 -3840 1720 -3800
rect 1660 -3870 1675 -3840
rect 1705 -3870 1720 -3840
rect 1660 -3910 1720 -3870
rect 1660 -3940 1675 -3910
rect 1705 -3940 1720 -3910
rect 1660 -3980 1720 -3940
rect 1660 -4010 1675 -3980
rect 1705 -4010 1720 -3980
rect 1660 -4045 1720 -4010
rect 1660 -4075 1675 -4045
rect 1705 -4075 1720 -4045
rect 1660 -4105 1720 -4075
rect 1660 -4135 1675 -4105
rect 1705 -4135 1720 -4105
rect 1660 -4170 1720 -4135
rect 1660 -4200 1675 -4170
rect 1705 -4200 1720 -4170
rect 1660 -4240 1720 -4200
rect 1660 -4270 1675 -4240
rect 1705 -4270 1720 -4240
rect 1660 -4310 1720 -4270
rect 1660 -4340 1675 -4310
rect 1705 -4340 1720 -4310
rect 1660 -4380 1720 -4340
rect 1660 -4410 1675 -4380
rect 1705 -4410 1720 -4380
rect 1660 -4445 1720 -4410
rect 1660 -4475 1675 -4445
rect 1705 -4475 1720 -4445
rect 1660 -4490 1720 -4475
rect 2010 -1305 2070 -1290
rect 2010 -1335 2025 -1305
rect 2055 -1335 2070 -1305
rect 2010 -1370 2070 -1335
rect 2010 -1400 2025 -1370
rect 2055 -1400 2070 -1370
rect 2010 -1440 2070 -1400
rect 2010 -1470 2025 -1440
rect 2055 -1470 2070 -1440
rect 2010 -1510 2070 -1470
rect 2010 -1540 2025 -1510
rect 2055 -1540 2070 -1510
rect 2010 -1580 2070 -1540
rect 2010 -1610 2025 -1580
rect 2055 -1610 2070 -1580
rect 2010 -1645 2070 -1610
rect 2010 -1675 2025 -1645
rect 2055 -1675 2070 -1645
rect 2010 -1705 2070 -1675
rect 2010 -1735 2025 -1705
rect 2055 -1735 2070 -1705
rect 2010 -1770 2070 -1735
rect 2010 -1800 2025 -1770
rect 2055 -1800 2070 -1770
rect 2010 -1840 2070 -1800
rect 2010 -1870 2025 -1840
rect 2055 -1870 2070 -1840
rect 2010 -1910 2070 -1870
rect 2010 -1940 2025 -1910
rect 2055 -1940 2070 -1910
rect 2010 -1980 2070 -1940
rect 2010 -2010 2025 -1980
rect 2055 -2010 2070 -1980
rect 2010 -2045 2070 -2010
rect 2010 -2075 2025 -2045
rect 2055 -2075 2070 -2045
rect 2010 -2105 2070 -2075
rect 2010 -2135 2025 -2105
rect 2055 -2135 2070 -2105
rect 2010 -2170 2070 -2135
rect 2010 -2200 2025 -2170
rect 2055 -2200 2070 -2170
rect 2010 -2240 2070 -2200
rect 2010 -2270 2025 -2240
rect 2055 -2270 2070 -2240
rect 2010 -2310 2070 -2270
rect 2010 -2340 2025 -2310
rect 2055 -2340 2070 -2310
rect 2010 -2380 2070 -2340
rect 2010 -2410 2025 -2380
rect 2055 -2410 2070 -2380
rect 2010 -2445 2070 -2410
rect 2010 -2475 2025 -2445
rect 2055 -2475 2070 -2445
rect 2010 -2505 2070 -2475
rect 2010 -2535 2025 -2505
rect 2055 -2535 2070 -2505
rect 2010 -2570 2070 -2535
rect 2010 -2600 2025 -2570
rect 2055 -2600 2070 -2570
rect 2010 -2640 2070 -2600
rect 2010 -2670 2025 -2640
rect 2055 -2670 2070 -2640
rect 2010 -2710 2070 -2670
rect 2010 -2740 2025 -2710
rect 2055 -2740 2070 -2710
rect 2010 -2780 2070 -2740
rect 2010 -2810 2025 -2780
rect 2055 -2810 2070 -2780
rect 2010 -2845 2070 -2810
rect 2010 -2875 2025 -2845
rect 2055 -2875 2070 -2845
rect 2010 -2905 2070 -2875
rect 2010 -2935 2025 -2905
rect 2055 -2935 2070 -2905
rect 2010 -2970 2070 -2935
rect 2010 -3000 2025 -2970
rect 2055 -3000 2070 -2970
rect 2010 -3040 2070 -3000
rect 2010 -3070 2025 -3040
rect 2055 -3070 2070 -3040
rect 2010 -3110 2070 -3070
rect 2010 -3140 2025 -3110
rect 2055 -3140 2070 -3110
rect 2010 -3180 2070 -3140
rect 2010 -3210 2025 -3180
rect 2055 -3210 2070 -3180
rect 2010 -3245 2070 -3210
rect 2010 -3275 2025 -3245
rect 2055 -3275 2070 -3245
rect 2010 -3305 2070 -3275
rect 2010 -3335 2025 -3305
rect 2055 -3335 2070 -3305
rect 2010 -3370 2070 -3335
rect 2010 -3400 2025 -3370
rect 2055 -3400 2070 -3370
rect 2010 -3440 2070 -3400
rect 2010 -3470 2025 -3440
rect 2055 -3470 2070 -3440
rect 2010 -3510 2070 -3470
rect 2010 -3540 2025 -3510
rect 2055 -3540 2070 -3510
rect 2010 -3580 2070 -3540
rect 2010 -3610 2025 -3580
rect 2055 -3610 2070 -3580
rect 2010 -3645 2070 -3610
rect 2010 -3675 2025 -3645
rect 2055 -3675 2070 -3645
rect 2010 -3705 2070 -3675
rect 2010 -3735 2025 -3705
rect 2055 -3735 2070 -3705
rect 2010 -3770 2070 -3735
rect 2010 -3800 2025 -3770
rect 2055 -3800 2070 -3770
rect 2010 -3840 2070 -3800
rect 2010 -3870 2025 -3840
rect 2055 -3870 2070 -3840
rect 2010 -3910 2070 -3870
rect 2010 -3940 2025 -3910
rect 2055 -3940 2070 -3910
rect 2010 -3980 2070 -3940
rect 2010 -4010 2025 -3980
rect 2055 -4010 2070 -3980
rect 2010 -4045 2070 -4010
rect 2010 -4075 2025 -4045
rect 2055 -4075 2070 -4045
rect 2010 -4105 2070 -4075
rect 2010 -4135 2025 -4105
rect 2055 -4135 2070 -4105
rect 2010 -4170 2070 -4135
rect 2010 -4200 2025 -4170
rect 2055 -4200 2070 -4170
rect 2010 -4240 2070 -4200
rect 2010 -4270 2025 -4240
rect 2055 -4270 2070 -4240
rect 2010 -4310 2070 -4270
rect 2010 -4340 2025 -4310
rect 2055 -4340 2070 -4310
rect 2010 -4380 2070 -4340
rect 2010 -4410 2025 -4380
rect 2055 -4410 2070 -4380
rect 2010 -4445 2070 -4410
rect 2010 -4475 2025 -4445
rect 2055 -4475 2070 -4445
rect 2010 -4490 2070 -4475
rect 2360 -1305 2420 -1290
rect 2360 -1335 2375 -1305
rect 2405 -1335 2420 -1305
rect 2360 -1370 2420 -1335
rect 2360 -1400 2375 -1370
rect 2405 -1400 2420 -1370
rect 2360 -1440 2420 -1400
rect 2360 -1470 2375 -1440
rect 2405 -1470 2420 -1440
rect 2360 -1510 2420 -1470
rect 2360 -1540 2375 -1510
rect 2405 -1540 2420 -1510
rect 2360 -1580 2420 -1540
rect 2360 -1610 2375 -1580
rect 2405 -1610 2420 -1580
rect 2360 -1645 2420 -1610
rect 2360 -1675 2375 -1645
rect 2405 -1675 2420 -1645
rect 2360 -1705 2420 -1675
rect 2360 -1735 2375 -1705
rect 2405 -1735 2420 -1705
rect 2360 -1770 2420 -1735
rect 2360 -1800 2375 -1770
rect 2405 -1800 2420 -1770
rect 2360 -1840 2420 -1800
rect 2360 -1870 2375 -1840
rect 2405 -1870 2420 -1840
rect 2360 -1910 2420 -1870
rect 2360 -1940 2375 -1910
rect 2405 -1940 2420 -1910
rect 2360 -1980 2420 -1940
rect 2360 -2010 2375 -1980
rect 2405 -2010 2420 -1980
rect 2360 -2045 2420 -2010
rect 2360 -2075 2375 -2045
rect 2405 -2075 2420 -2045
rect 2360 -2105 2420 -2075
rect 2360 -2135 2375 -2105
rect 2405 -2135 2420 -2105
rect 2360 -2170 2420 -2135
rect 2360 -2200 2375 -2170
rect 2405 -2200 2420 -2170
rect 2360 -2240 2420 -2200
rect 2360 -2270 2375 -2240
rect 2405 -2270 2420 -2240
rect 2360 -2310 2420 -2270
rect 2360 -2340 2375 -2310
rect 2405 -2340 2420 -2310
rect 2360 -2380 2420 -2340
rect 2360 -2410 2375 -2380
rect 2405 -2410 2420 -2380
rect 2360 -2445 2420 -2410
rect 2360 -2475 2375 -2445
rect 2405 -2475 2420 -2445
rect 2360 -2505 2420 -2475
rect 2360 -2535 2375 -2505
rect 2405 -2535 2420 -2505
rect 2360 -2570 2420 -2535
rect 2360 -2600 2375 -2570
rect 2405 -2600 2420 -2570
rect 2360 -2640 2420 -2600
rect 2360 -2670 2375 -2640
rect 2405 -2670 2420 -2640
rect 2360 -2710 2420 -2670
rect 2360 -2740 2375 -2710
rect 2405 -2740 2420 -2710
rect 2360 -2780 2420 -2740
rect 2360 -2810 2375 -2780
rect 2405 -2810 2420 -2780
rect 2360 -2845 2420 -2810
rect 2360 -2875 2375 -2845
rect 2405 -2875 2420 -2845
rect 2360 -2905 2420 -2875
rect 2360 -2935 2375 -2905
rect 2405 -2935 2420 -2905
rect 2360 -2970 2420 -2935
rect 2360 -3000 2375 -2970
rect 2405 -3000 2420 -2970
rect 2360 -3040 2420 -3000
rect 2360 -3070 2375 -3040
rect 2405 -3070 2420 -3040
rect 2360 -3110 2420 -3070
rect 2360 -3140 2375 -3110
rect 2405 -3140 2420 -3110
rect 2360 -3180 2420 -3140
rect 2360 -3210 2375 -3180
rect 2405 -3210 2420 -3180
rect 2360 -3245 2420 -3210
rect 2360 -3275 2375 -3245
rect 2405 -3275 2420 -3245
rect 2360 -3305 2420 -3275
rect 2360 -3335 2375 -3305
rect 2405 -3335 2420 -3305
rect 2360 -3370 2420 -3335
rect 2360 -3400 2375 -3370
rect 2405 -3400 2420 -3370
rect 2360 -3440 2420 -3400
rect 2360 -3470 2375 -3440
rect 2405 -3470 2420 -3440
rect 2360 -3510 2420 -3470
rect 2360 -3540 2375 -3510
rect 2405 -3540 2420 -3510
rect 2360 -3580 2420 -3540
rect 2360 -3610 2375 -3580
rect 2405 -3610 2420 -3580
rect 2360 -3645 2420 -3610
rect 2360 -3675 2375 -3645
rect 2405 -3675 2420 -3645
rect 2360 -3705 2420 -3675
rect 2360 -3735 2375 -3705
rect 2405 -3735 2420 -3705
rect 2360 -3770 2420 -3735
rect 2360 -3800 2375 -3770
rect 2405 -3800 2420 -3770
rect 2360 -3840 2420 -3800
rect 2360 -3870 2375 -3840
rect 2405 -3870 2420 -3840
rect 2360 -3910 2420 -3870
rect 2360 -3940 2375 -3910
rect 2405 -3940 2420 -3910
rect 2360 -3980 2420 -3940
rect 2360 -4010 2375 -3980
rect 2405 -4010 2420 -3980
rect 2360 -4045 2420 -4010
rect 2360 -4075 2375 -4045
rect 2405 -4075 2420 -4045
rect 2360 -4105 2420 -4075
rect 2360 -4135 2375 -4105
rect 2405 -4135 2420 -4105
rect 2360 -4170 2420 -4135
rect 2360 -4200 2375 -4170
rect 2405 -4200 2420 -4170
rect 2360 -4240 2420 -4200
rect 2360 -4270 2375 -4240
rect 2405 -4270 2420 -4240
rect 2360 -4310 2420 -4270
rect 2360 -4340 2375 -4310
rect 2405 -4340 2420 -4310
rect 2360 -4380 2420 -4340
rect 2360 -4410 2375 -4380
rect 2405 -4410 2420 -4380
rect 2360 -4445 2420 -4410
rect 2360 -4475 2375 -4445
rect 2405 -4475 2420 -4445
rect 2360 -4490 2420 -4475
rect 2710 -1305 2770 -1290
rect 2710 -1335 2725 -1305
rect 2755 -1335 2770 -1305
rect 2710 -1370 2770 -1335
rect 2710 -1400 2725 -1370
rect 2755 -1400 2770 -1370
rect 2710 -1440 2770 -1400
rect 2710 -1470 2725 -1440
rect 2755 -1470 2770 -1440
rect 2710 -1510 2770 -1470
rect 2710 -1540 2725 -1510
rect 2755 -1540 2770 -1510
rect 2710 -1580 2770 -1540
rect 2710 -1610 2725 -1580
rect 2755 -1610 2770 -1580
rect 2710 -1645 2770 -1610
rect 2710 -1675 2725 -1645
rect 2755 -1675 2770 -1645
rect 2710 -1705 2770 -1675
rect 2710 -1735 2725 -1705
rect 2755 -1735 2770 -1705
rect 2710 -1770 2770 -1735
rect 2710 -1800 2725 -1770
rect 2755 -1800 2770 -1770
rect 2710 -1840 2770 -1800
rect 2710 -1870 2725 -1840
rect 2755 -1870 2770 -1840
rect 2710 -1910 2770 -1870
rect 2710 -1940 2725 -1910
rect 2755 -1940 2770 -1910
rect 2710 -1980 2770 -1940
rect 2710 -2010 2725 -1980
rect 2755 -2010 2770 -1980
rect 2710 -2045 2770 -2010
rect 2710 -2075 2725 -2045
rect 2755 -2075 2770 -2045
rect 2710 -2105 2770 -2075
rect 2710 -2135 2725 -2105
rect 2755 -2135 2770 -2105
rect 2710 -2170 2770 -2135
rect 2710 -2200 2725 -2170
rect 2755 -2200 2770 -2170
rect 2710 -2240 2770 -2200
rect 2710 -2270 2725 -2240
rect 2755 -2270 2770 -2240
rect 2710 -2310 2770 -2270
rect 2710 -2340 2725 -2310
rect 2755 -2340 2770 -2310
rect 2710 -2380 2770 -2340
rect 2710 -2410 2725 -2380
rect 2755 -2410 2770 -2380
rect 2710 -2445 2770 -2410
rect 2710 -2475 2725 -2445
rect 2755 -2475 2770 -2445
rect 2710 -2505 2770 -2475
rect 2710 -2535 2725 -2505
rect 2755 -2535 2770 -2505
rect 2710 -2570 2770 -2535
rect 2710 -2600 2725 -2570
rect 2755 -2600 2770 -2570
rect 2710 -2640 2770 -2600
rect 2710 -2670 2725 -2640
rect 2755 -2670 2770 -2640
rect 2710 -2710 2770 -2670
rect 2710 -2740 2725 -2710
rect 2755 -2740 2770 -2710
rect 2710 -2780 2770 -2740
rect 2710 -2810 2725 -2780
rect 2755 -2810 2770 -2780
rect 2710 -2845 2770 -2810
rect 2710 -2875 2725 -2845
rect 2755 -2875 2770 -2845
rect 2710 -2905 2770 -2875
rect 2710 -2935 2725 -2905
rect 2755 -2935 2770 -2905
rect 2710 -2970 2770 -2935
rect 2710 -3000 2725 -2970
rect 2755 -3000 2770 -2970
rect 2710 -3040 2770 -3000
rect 2710 -3070 2725 -3040
rect 2755 -3070 2770 -3040
rect 2710 -3110 2770 -3070
rect 2710 -3140 2725 -3110
rect 2755 -3140 2770 -3110
rect 2710 -3180 2770 -3140
rect 2710 -3210 2725 -3180
rect 2755 -3210 2770 -3180
rect 2710 -3245 2770 -3210
rect 2710 -3275 2725 -3245
rect 2755 -3275 2770 -3245
rect 2710 -3305 2770 -3275
rect 2710 -3335 2725 -3305
rect 2755 -3335 2770 -3305
rect 2710 -3370 2770 -3335
rect 2710 -3400 2725 -3370
rect 2755 -3400 2770 -3370
rect 2710 -3440 2770 -3400
rect 2710 -3470 2725 -3440
rect 2755 -3470 2770 -3440
rect 2710 -3510 2770 -3470
rect 2710 -3540 2725 -3510
rect 2755 -3540 2770 -3510
rect 2710 -3580 2770 -3540
rect 2710 -3610 2725 -3580
rect 2755 -3610 2770 -3580
rect 2710 -3645 2770 -3610
rect 2710 -3675 2725 -3645
rect 2755 -3675 2770 -3645
rect 2710 -3705 2770 -3675
rect 2710 -3735 2725 -3705
rect 2755 -3735 2770 -3705
rect 2710 -3770 2770 -3735
rect 2710 -3800 2725 -3770
rect 2755 -3800 2770 -3770
rect 2710 -3840 2770 -3800
rect 2710 -3870 2725 -3840
rect 2755 -3870 2770 -3840
rect 2710 -3910 2770 -3870
rect 2710 -3940 2725 -3910
rect 2755 -3940 2770 -3910
rect 2710 -3980 2770 -3940
rect 2710 -4010 2725 -3980
rect 2755 -4010 2770 -3980
rect 2710 -4045 2770 -4010
rect 2710 -4075 2725 -4045
rect 2755 -4075 2770 -4045
rect 2710 -4105 2770 -4075
rect 2710 -4135 2725 -4105
rect 2755 -4135 2770 -4105
rect 2710 -4170 2770 -4135
rect 2710 -4200 2725 -4170
rect 2755 -4200 2770 -4170
rect 2710 -4240 2770 -4200
rect 2710 -4270 2725 -4240
rect 2755 -4270 2770 -4240
rect 2710 -4310 2770 -4270
rect 2710 -4340 2725 -4310
rect 2755 -4340 2770 -4310
rect 2710 -4380 2770 -4340
rect 2710 -4410 2725 -4380
rect 2755 -4410 2770 -4380
rect 2710 -4445 2770 -4410
rect 2710 -4475 2725 -4445
rect 2755 -4475 2770 -4445
rect 2710 -4490 2770 -4475
rect 3060 -1305 3120 -1290
rect 3060 -1335 3075 -1305
rect 3105 -1335 3120 -1305
rect 3060 -1370 3120 -1335
rect 3060 -1400 3075 -1370
rect 3105 -1400 3120 -1370
rect 3060 -1440 3120 -1400
rect 3060 -1470 3075 -1440
rect 3105 -1470 3120 -1440
rect 3060 -1510 3120 -1470
rect 3060 -1540 3075 -1510
rect 3105 -1540 3120 -1510
rect 3060 -1580 3120 -1540
rect 3060 -1610 3075 -1580
rect 3105 -1610 3120 -1580
rect 3060 -1645 3120 -1610
rect 3060 -1675 3075 -1645
rect 3105 -1675 3120 -1645
rect 3060 -1705 3120 -1675
rect 3060 -1735 3075 -1705
rect 3105 -1735 3120 -1705
rect 3060 -1770 3120 -1735
rect 3060 -1800 3075 -1770
rect 3105 -1800 3120 -1770
rect 3060 -1840 3120 -1800
rect 3060 -1870 3075 -1840
rect 3105 -1870 3120 -1840
rect 3060 -1910 3120 -1870
rect 3060 -1940 3075 -1910
rect 3105 -1940 3120 -1910
rect 3060 -1980 3120 -1940
rect 3060 -2010 3075 -1980
rect 3105 -2010 3120 -1980
rect 3060 -2045 3120 -2010
rect 3060 -2075 3075 -2045
rect 3105 -2075 3120 -2045
rect 3060 -2105 3120 -2075
rect 3060 -2135 3075 -2105
rect 3105 -2135 3120 -2105
rect 3060 -2170 3120 -2135
rect 3060 -2200 3075 -2170
rect 3105 -2200 3120 -2170
rect 3060 -2240 3120 -2200
rect 3060 -2270 3075 -2240
rect 3105 -2270 3120 -2240
rect 3060 -2310 3120 -2270
rect 3060 -2340 3075 -2310
rect 3105 -2340 3120 -2310
rect 3060 -2380 3120 -2340
rect 3060 -2410 3075 -2380
rect 3105 -2410 3120 -2380
rect 3060 -2445 3120 -2410
rect 3060 -2475 3075 -2445
rect 3105 -2475 3120 -2445
rect 3060 -2505 3120 -2475
rect 3060 -2535 3075 -2505
rect 3105 -2535 3120 -2505
rect 3060 -2570 3120 -2535
rect 3060 -2600 3075 -2570
rect 3105 -2600 3120 -2570
rect 3060 -2640 3120 -2600
rect 3060 -2670 3075 -2640
rect 3105 -2670 3120 -2640
rect 3060 -2710 3120 -2670
rect 3060 -2740 3075 -2710
rect 3105 -2740 3120 -2710
rect 3060 -2780 3120 -2740
rect 3060 -2810 3075 -2780
rect 3105 -2810 3120 -2780
rect 3060 -2845 3120 -2810
rect 3060 -2875 3075 -2845
rect 3105 -2875 3120 -2845
rect 3060 -2905 3120 -2875
rect 3060 -2935 3075 -2905
rect 3105 -2935 3120 -2905
rect 3060 -2970 3120 -2935
rect 3060 -3000 3075 -2970
rect 3105 -3000 3120 -2970
rect 3060 -3040 3120 -3000
rect 3060 -3070 3075 -3040
rect 3105 -3070 3120 -3040
rect 3060 -3110 3120 -3070
rect 3060 -3140 3075 -3110
rect 3105 -3140 3120 -3110
rect 3060 -3180 3120 -3140
rect 3060 -3210 3075 -3180
rect 3105 -3210 3120 -3180
rect 3060 -3245 3120 -3210
rect 3060 -3275 3075 -3245
rect 3105 -3275 3120 -3245
rect 3060 -3305 3120 -3275
rect 3060 -3335 3075 -3305
rect 3105 -3335 3120 -3305
rect 3060 -3370 3120 -3335
rect 3060 -3400 3075 -3370
rect 3105 -3400 3120 -3370
rect 3060 -3440 3120 -3400
rect 3060 -3470 3075 -3440
rect 3105 -3470 3120 -3440
rect 3060 -3510 3120 -3470
rect 3060 -3540 3075 -3510
rect 3105 -3540 3120 -3510
rect 3060 -3580 3120 -3540
rect 3060 -3610 3075 -3580
rect 3105 -3610 3120 -3580
rect 3060 -3645 3120 -3610
rect 3060 -3675 3075 -3645
rect 3105 -3675 3120 -3645
rect 3060 -3705 3120 -3675
rect 3060 -3735 3075 -3705
rect 3105 -3735 3120 -3705
rect 3060 -3770 3120 -3735
rect 3060 -3800 3075 -3770
rect 3105 -3800 3120 -3770
rect 3060 -3840 3120 -3800
rect 3060 -3870 3075 -3840
rect 3105 -3870 3120 -3840
rect 3060 -3910 3120 -3870
rect 3060 -3940 3075 -3910
rect 3105 -3940 3120 -3910
rect 3060 -3980 3120 -3940
rect 3060 -4010 3075 -3980
rect 3105 -4010 3120 -3980
rect 3060 -4045 3120 -4010
rect 3060 -4075 3075 -4045
rect 3105 -4075 3120 -4045
rect 3060 -4105 3120 -4075
rect 3060 -4135 3075 -4105
rect 3105 -4135 3120 -4105
rect 3060 -4170 3120 -4135
rect 3060 -4200 3075 -4170
rect 3105 -4200 3120 -4170
rect 3060 -4240 3120 -4200
rect 3060 -4270 3075 -4240
rect 3105 -4270 3120 -4240
rect 3060 -4310 3120 -4270
rect 3060 -4340 3075 -4310
rect 3105 -4340 3120 -4310
rect 3060 -4380 3120 -4340
rect 3060 -4410 3075 -4380
rect 3105 -4410 3120 -4380
rect 3060 -4445 3120 -4410
rect 3060 -4475 3075 -4445
rect 3105 -4475 3120 -4445
rect 3060 -4490 3120 -4475
rect 3410 -1305 3470 -1290
rect 3410 -1335 3425 -1305
rect 3455 -1335 3470 -1305
rect 3410 -1370 3470 -1335
rect 3410 -1400 3425 -1370
rect 3455 -1400 3470 -1370
rect 3410 -1440 3470 -1400
rect 3410 -1470 3425 -1440
rect 3455 -1470 3470 -1440
rect 3410 -1510 3470 -1470
rect 3410 -1540 3425 -1510
rect 3455 -1540 3470 -1510
rect 3410 -1580 3470 -1540
rect 3410 -1610 3425 -1580
rect 3455 -1610 3470 -1580
rect 3410 -1645 3470 -1610
rect 3410 -1675 3425 -1645
rect 3455 -1675 3470 -1645
rect 3410 -1705 3470 -1675
rect 3410 -1735 3425 -1705
rect 3455 -1735 3470 -1705
rect 3410 -1770 3470 -1735
rect 3410 -1800 3425 -1770
rect 3455 -1800 3470 -1770
rect 3410 -1840 3470 -1800
rect 3410 -1870 3425 -1840
rect 3455 -1870 3470 -1840
rect 3410 -1910 3470 -1870
rect 3410 -1940 3425 -1910
rect 3455 -1940 3470 -1910
rect 3410 -1980 3470 -1940
rect 3410 -2010 3425 -1980
rect 3455 -2010 3470 -1980
rect 3410 -2045 3470 -2010
rect 3410 -2075 3425 -2045
rect 3455 -2075 3470 -2045
rect 3410 -2105 3470 -2075
rect 3410 -2135 3425 -2105
rect 3455 -2135 3470 -2105
rect 3410 -2170 3470 -2135
rect 3410 -2200 3425 -2170
rect 3455 -2200 3470 -2170
rect 3410 -2240 3470 -2200
rect 3410 -2270 3425 -2240
rect 3455 -2270 3470 -2240
rect 3410 -2310 3470 -2270
rect 3410 -2340 3425 -2310
rect 3455 -2340 3470 -2310
rect 3410 -2380 3470 -2340
rect 3410 -2410 3425 -2380
rect 3455 -2410 3470 -2380
rect 3410 -2445 3470 -2410
rect 3410 -2475 3425 -2445
rect 3455 -2475 3470 -2445
rect 3410 -2505 3470 -2475
rect 3410 -2535 3425 -2505
rect 3455 -2535 3470 -2505
rect 3410 -2570 3470 -2535
rect 3410 -2600 3425 -2570
rect 3455 -2600 3470 -2570
rect 3410 -2640 3470 -2600
rect 3410 -2670 3425 -2640
rect 3455 -2670 3470 -2640
rect 3410 -2710 3470 -2670
rect 3410 -2740 3425 -2710
rect 3455 -2740 3470 -2710
rect 3410 -2780 3470 -2740
rect 3410 -2810 3425 -2780
rect 3455 -2810 3470 -2780
rect 3410 -2845 3470 -2810
rect 3410 -2875 3425 -2845
rect 3455 -2875 3470 -2845
rect 3410 -2905 3470 -2875
rect 3410 -2935 3425 -2905
rect 3455 -2935 3470 -2905
rect 3410 -2970 3470 -2935
rect 3410 -3000 3425 -2970
rect 3455 -3000 3470 -2970
rect 3410 -3040 3470 -3000
rect 3410 -3070 3425 -3040
rect 3455 -3070 3470 -3040
rect 3410 -3110 3470 -3070
rect 3410 -3140 3425 -3110
rect 3455 -3140 3470 -3110
rect 3410 -3180 3470 -3140
rect 3410 -3210 3425 -3180
rect 3455 -3210 3470 -3180
rect 3410 -3245 3470 -3210
rect 3410 -3275 3425 -3245
rect 3455 -3275 3470 -3245
rect 3410 -3305 3470 -3275
rect 3410 -3335 3425 -3305
rect 3455 -3335 3470 -3305
rect 3410 -3370 3470 -3335
rect 3410 -3400 3425 -3370
rect 3455 -3400 3470 -3370
rect 3410 -3440 3470 -3400
rect 3410 -3470 3425 -3440
rect 3455 -3470 3470 -3440
rect 3410 -3510 3470 -3470
rect 3410 -3540 3425 -3510
rect 3455 -3540 3470 -3510
rect 3410 -3580 3470 -3540
rect 3410 -3610 3425 -3580
rect 3455 -3610 3470 -3580
rect 3410 -3645 3470 -3610
rect 3410 -3675 3425 -3645
rect 3455 -3675 3470 -3645
rect 3410 -3705 3470 -3675
rect 3410 -3735 3425 -3705
rect 3455 -3735 3470 -3705
rect 3410 -3770 3470 -3735
rect 3410 -3800 3425 -3770
rect 3455 -3800 3470 -3770
rect 3410 -3840 3470 -3800
rect 3410 -3870 3425 -3840
rect 3455 -3870 3470 -3840
rect 3410 -3910 3470 -3870
rect 3410 -3940 3425 -3910
rect 3455 -3940 3470 -3910
rect 3410 -3980 3470 -3940
rect 3410 -4010 3425 -3980
rect 3455 -4010 3470 -3980
rect 3410 -4045 3470 -4010
rect 3410 -4075 3425 -4045
rect 3455 -4075 3470 -4045
rect 3410 -4105 3470 -4075
rect 3410 -4135 3425 -4105
rect 3455 -4135 3470 -4105
rect 3410 -4170 3470 -4135
rect 3410 -4200 3425 -4170
rect 3455 -4200 3470 -4170
rect 3410 -4240 3470 -4200
rect 3410 -4270 3425 -4240
rect 3455 -4270 3470 -4240
rect 3410 -4310 3470 -4270
rect 3410 -4340 3425 -4310
rect 3455 -4340 3470 -4310
rect 3410 -4380 3470 -4340
rect 3410 -4410 3425 -4380
rect 3455 -4410 3470 -4380
rect 3410 -4445 3470 -4410
rect 3410 -4475 3425 -4445
rect 3455 -4475 3470 -4445
rect 3410 -4490 3470 -4475
rect 3760 -1305 3820 -1290
rect 3760 -1335 3775 -1305
rect 3805 -1335 3820 -1305
rect 3760 -1370 3820 -1335
rect 3760 -1400 3775 -1370
rect 3805 -1400 3820 -1370
rect 3760 -1440 3820 -1400
rect 3760 -1470 3775 -1440
rect 3805 -1470 3820 -1440
rect 3760 -1510 3820 -1470
rect 3760 -1540 3775 -1510
rect 3805 -1540 3820 -1510
rect 3760 -1580 3820 -1540
rect 3760 -1610 3775 -1580
rect 3805 -1610 3820 -1580
rect 3760 -1645 3820 -1610
rect 3760 -1675 3775 -1645
rect 3805 -1675 3820 -1645
rect 3760 -1705 3820 -1675
rect 3760 -1735 3775 -1705
rect 3805 -1735 3820 -1705
rect 3760 -1770 3820 -1735
rect 3760 -1800 3775 -1770
rect 3805 -1800 3820 -1770
rect 3760 -1840 3820 -1800
rect 3760 -1870 3775 -1840
rect 3805 -1870 3820 -1840
rect 3760 -1910 3820 -1870
rect 3760 -1940 3775 -1910
rect 3805 -1940 3820 -1910
rect 3760 -1980 3820 -1940
rect 3760 -2010 3775 -1980
rect 3805 -2010 3820 -1980
rect 3760 -2045 3820 -2010
rect 3760 -2075 3775 -2045
rect 3805 -2075 3820 -2045
rect 3760 -2105 3820 -2075
rect 3760 -2135 3775 -2105
rect 3805 -2135 3820 -2105
rect 3760 -2170 3820 -2135
rect 3760 -2200 3775 -2170
rect 3805 -2200 3820 -2170
rect 3760 -2240 3820 -2200
rect 3760 -2270 3775 -2240
rect 3805 -2270 3820 -2240
rect 3760 -2310 3820 -2270
rect 3760 -2340 3775 -2310
rect 3805 -2340 3820 -2310
rect 3760 -2380 3820 -2340
rect 3760 -2410 3775 -2380
rect 3805 -2410 3820 -2380
rect 3760 -2445 3820 -2410
rect 3760 -2475 3775 -2445
rect 3805 -2475 3820 -2445
rect 3760 -2505 3820 -2475
rect 3760 -2535 3775 -2505
rect 3805 -2535 3820 -2505
rect 3760 -2570 3820 -2535
rect 3760 -2600 3775 -2570
rect 3805 -2600 3820 -2570
rect 3760 -2640 3820 -2600
rect 3760 -2670 3775 -2640
rect 3805 -2670 3820 -2640
rect 3760 -2710 3820 -2670
rect 3760 -2740 3775 -2710
rect 3805 -2740 3820 -2710
rect 3760 -2780 3820 -2740
rect 3760 -2810 3775 -2780
rect 3805 -2810 3820 -2780
rect 3760 -2845 3820 -2810
rect 3760 -2875 3775 -2845
rect 3805 -2875 3820 -2845
rect 3760 -2905 3820 -2875
rect 3760 -2935 3775 -2905
rect 3805 -2935 3820 -2905
rect 3760 -2970 3820 -2935
rect 3760 -3000 3775 -2970
rect 3805 -3000 3820 -2970
rect 3760 -3040 3820 -3000
rect 3760 -3070 3775 -3040
rect 3805 -3070 3820 -3040
rect 3760 -3110 3820 -3070
rect 3760 -3140 3775 -3110
rect 3805 -3140 3820 -3110
rect 3760 -3180 3820 -3140
rect 3760 -3210 3775 -3180
rect 3805 -3210 3820 -3180
rect 3760 -3245 3820 -3210
rect 3760 -3275 3775 -3245
rect 3805 -3275 3820 -3245
rect 3760 -3305 3820 -3275
rect 3760 -3335 3775 -3305
rect 3805 -3335 3820 -3305
rect 3760 -3370 3820 -3335
rect 3760 -3400 3775 -3370
rect 3805 -3400 3820 -3370
rect 3760 -3440 3820 -3400
rect 3760 -3470 3775 -3440
rect 3805 -3470 3820 -3440
rect 3760 -3510 3820 -3470
rect 3760 -3540 3775 -3510
rect 3805 -3540 3820 -3510
rect 3760 -3580 3820 -3540
rect 3760 -3610 3775 -3580
rect 3805 -3610 3820 -3580
rect 3760 -3645 3820 -3610
rect 3760 -3675 3775 -3645
rect 3805 -3675 3820 -3645
rect 3760 -3705 3820 -3675
rect 3760 -3735 3775 -3705
rect 3805 -3735 3820 -3705
rect 3760 -3770 3820 -3735
rect 3760 -3800 3775 -3770
rect 3805 -3800 3820 -3770
rect 3760 -3840 3820 -3800
rect 3760 -3870 3775 -3840
rect 3805 -3870 3820 -3840
rect 3760 -3910 3820 -3870
rect 3760 -3940 3775 -3910
rect 3805 -3940 3820 -3910
rect 3760 -3980 3820 -3940
rect 3760 -4010 3775 -3980
rect 3805 -4010 3820 -3980
rect 3760 -4045 3820 -4010
rect 3760 -4075 3775 -4045
rect 3805 -4075 3820 -4045
rect 3760 -4105 3820 -4075
rect 3760 -4135 3775 -4105
rect 3805 -4135 3820 -4105
rect 3760 -4170 3820 -4135
rect 3760 -4200 3775 -4170
rect 3805 -4200 3820 -4170
rect 3760 -4240 3820 -4200
rect 3760 -4270 3775 -4240
rect 3805 -4270 3820 -4240
rect 3760 -4310 3820 -4270
rect 3760 -4340 3775 -4310
rect 3805 -4340 3820 -4310
rect 3760 -4380 3820 -4340
rect 3760 -4410 3775 -4380
rect 3805 -4410 3820 -4380
rect 3760 -4445 3820 -4410
rect 3760 -4475 3775 -4445
rect 3805 -4475 3820 -4445
rect 3760 -4490 3820 -4475
rect 4110 -1305 4170 -1290
rect 4110 -1335 4125 -1305
rect 4155 -1335 4170 -1305
rect 4110 -1370 4170 -1335
rect 4110 -1400 4125 -1370
rect 4155 -1400 4170 -1370
rect 4110 -1440 4170 -1400
rect 4110 -1470 4125 -1440
rect 4155 -1470 4170 -1440
rect 4110 -1510 4170 -1470
rect 4110 -1540 4125 -1510
rect 4155 -1540 4170 -1510
rect 4110 -1580 4170 -1540
rect 4110 -1610 4125 -1580
rect 4155 -1610 4170 -1580
rect 4110 -1645 4170 -1610
rect 4110 -1675 4125 -1645
rect 4155 -1675 4170 -1645
rect 4110 -1705 4170 -1675
rect 4110 -1735 4125 -1705
rect 4155 -1735 4170 -1705
rect 4110 -1770 4170 -1735
rect 4110 -1800 4125 -1770
rect 4155 -1800 4170 -1770
rect 4110 -1840 4170 -1800
rect 4110 -1870 4125 -1840
rect 4155 -1870 4170 -1840
rect 4110 -1910 4170 -1870
rect 4110 -1940 4125 -1910
rect 4155 -1940 4170 -1910
rect 4110 -1980 4170 -1940
rect 4110 -2010 4125 -1980
rect 4155 -2010 4170 -1980
rect 4110 -2045 4170 -2010
rect 4110 -2075 4125 -2045
rect 4155 -2075 4170 -2045
rect 4110 -2105 4170 -2075
rect 4110 -2135 4125 -2105
rect 4155 -2135 4170 -2105
rect 4110 -2170 4170 -2135
rect 4110 -2200 4125 -2170
rect 4155 -2200 4170 -2170
rect 4110 -2240 4170 -2200
rect 4110 -2270 4125 -2240
rect 4155 -2270 4170 -2240
rect 4110 -2310 4170 -2270
rect 4110 -2340 4125 -2310
rect 4155 -2340 4170 -2310
rect 4110 -2380 4170 -2340
rect 4110 -2410 4125 -2380
rect 4155 -2410 4170 -2380
rect 4110 -2445 4170 -2410
rect 4110 -2475 4125 -2445
rect 4155 -2475 4170 -2445
rect 4110 -2505 4170 -2475
rect 4110 -2535 4125 -2505
rect 4155 -2535 4170 -2505
rect 4110 -2570 4170 -2535
rect 4110 -2600 4125 -2570
rect 4155 -2600 4170 -2570
rect 4110 -2640 4170 -2600
rect 4110 -2670 4125 -2640
rect 4155 -2670 4170 -2640
rect 4110 -2710 4170 -2670
rect 4110 -2740 4125 -2710
rect 4155 -2740 4170 -2710
rect 4110 -2780 4170 -2740
rect 4110 -2810 4125 -2780
rect 4155 -2810 4170 -2780
rect 4110 -2845 4170 -2810
rect 4110 -2875 4125 -2845
rect 4155 -2875 4170 -2845
rect 4110 -2905 4170 -2875
rect 4110 -2935 4125 -2905
rect 4155 -2935 4170 -2905
rect 4110 -2970 4170 -2935
rect 4110 -3000 4125 -2970
rect 4155 -3000 4170 -2970
rect 4110 -3040 4170 -3000
rect 4110 -3070 4125 -3040
rect 4155 -3070 4170 -3040
rect 4110 -3110 4170 -3070
rect 4110 -3140 4125 -3110
rect 4155 -3140 4170 -3110
rect 4110 -3180 4170 -3140
rect 4110 -3210 4125 -3180
rect 4155 -3210 4170 -3180
rect 4110 -3245 4170 -3210
rect 4110 -3275 4125 -3245
rect 4155 -3275 4170 -3245
rect 4110 -3305 4170 -3275
rect 4110 -3335 4125 -3305
rect 4155 -3335 4170 -3305
rect 4110 -3370 4170 -3335
rect 4110 -3400 4125 -3370
rect 4155 -3400 4170 -3370
rect 4110 -3440 4170 -3400
rect 4110 -3470 4125 -3440
rect 4155 -3470 4170 -3440
rect 4110 -3510 4170 -3470
rect 4110 -3540 4125 -3510
rect 4155 -3540 4170 -3510
rect 4110 -3580 4170 -3540
rect 4110 -3610 4125 -3580
rect 4155 -3610 4170 -3580
rect 4110 -3645 4170 -3610
rect 4110 -3675 4125 -3645
rect 4155 -3675 4170 -3645
rect 4110 -3705 4170 -3675
rect 4110 -3735 4125 -3705
rect 4155 -3735 4170 -3705
rect 4110 -3770 4170 -3735
rect 4110 -3800 4125 -3770
rect 4155 -3800 4170 -3770
rect 4110 -3840 4170 -3800
rect 4110 -3870 4125 -3840
rect 4155 -3870 4170 -3840
rect 4110 -3910 4170 -3870
rect 4110 -3940 4125 -3910
rect 4155 -3940 4170 -3910
rect 4110 -3980 4170 -3940
rect 4110 -4010 4125 -3980
rect 4155 -4010 4170 -3980
rect 4110 -4045 4170 -4010
rect 4110 -4075 4125 -4045
rect 4155 -4075 4170 -4045
rect 4110 -4105 4170 -4075
rect 4110 -4135 4125 -4105
rect 4155 -4135 4170 -4105
rect 4110 -4170 4170 -4135
rect 4110 -4200 4125 -4170
rect 4155 -4200 4170 -4170
rect 4110 -4240 4170 -4200
rect 4110 -4270 4125 -4240
rect 4155 -4270 4170 -4240
rect 4110 -4310 4170 -4270
rect 4110 -4340 4125 -4310
rect 4155 -4340 4170 -4310
rect 4110 -4380 4170 -4340
rect 4110 -4410 4125 -4380
rect 4155 -4410 4170 -4380
rect 4110 -4445 4170 -4410
rect 4110 -4475 4125 -4445
rect 4155 -4475 4170 -4445
rect 4110 -4490 4170 -4475
rect 4460 -1305 4520 -1290
rect 4460 -1335 4475 -1305
rect 4505 -1335 4520 -1305
rect 4460 -1370 4520 -1335
rect 4460 -1400 4475 -1370
rect 4505 -1400 4520 -1370
rect 4460 -1440 4520 -1400
rect 4460 -1470 4475 -1440
rect 4505 -1470 4520 -1440
rect 4460 -1510 4520 -1470
rect 4460 -1540 4475 -1510
rect 4505 -1540 4520 -1510
rect 4460 -1580 4520 -1540
rect 4460 -1610 4475 -1580
rect 4505 -1610 4520 -1580
rect 4460 -1645 4520 -1610
rect 4460 -1675 4475 -1645
rect 4505 -1675 4520 -1645
rect 4460 -1705 4520 -1675
rect 4460 -1735 4475 -1705
rect 4505 -1735 4520 -1705
rect 4460 -1770 4520 -1735
rect 4460 -1800 4475 -1770
rect 4505 -1800 4520 -1770
rect 4460 -1840 4520 -1800
rect 4460 -1870 4475 -1840
rect 4505 -1870 4520 -1840
rect 4460 -1910 4520 -1870
rect 4460 -1940 4475 -1910
rect 4505 -1940 4520 -1910
rect 4460 -1980 4520 -1940
rect 4460 -2010 4475 -1980
rect 4505 -2010 4520 -1980
rect 4460 -2045 4520 -2010
rect 4460 -2075 4475 -2045
rect 4505 -2075 4520 -2045
rect 4460 -2105 4520 -2075
rect 4460 -2135 4475 -2105
rect 4505 -2135 4520 -2105
rect 4460 -2170 4520 -2135
rect 4460 -2200 4475 -2170
rect 4505 -2200 4520 -2170
rect 4460 -2240 4520 -2200
rect 4460 -2270 4475 -2240
rect 4505 -2270 4520 -2240
rect 4460 -2310 4520 -2270
rect 4460 -2340 4475 -2310
rect 4505 -2340 4520 -2310
rect 4460 -2380 4520 -2340
rect 4460 -2410 4475 -2380
rect 4505 -2410 4520 -2380
rect 4460 -2445 4520 -2410
rect 4460 -2475 4475 -2445
rect 4505 -2475 4520 -2445
rect 4460 -2505 4520 -2475
rect 4460 -2535 4475 -2505
rect 4505 -2535 4520 -2505
rect 4460 -2570 4520 -2535
rect 4460 -2600 4475 -2570
rect 4505 -2600 4520 -2570
rect 4460 -2640 4520 -2600
rect 4460 -2670 4475 -2640
rect 4505 -2670 4520 -2640
rect 4460 -2710 4520 -2670
rect 4460 -2740 4475 -2710
rect 4505 -2740 4520 -2710
rect 4460 -2780 4520 -2740
rect 4460 -2810 4475 -2780
rect 4505 -2810 4520 -2780
rect 4460 -2845 4520 -2810
rect 4460 -2875 4475 -2845
rect 4505 -2875 4520 -2845
rect 4460 -2905 4520 -2875
rect 4460 -2935 4475 -2905
rect 4505 -2935 4520 -2905
rect 4460 -2970 4520 -2935
rect 4460 -3000 4475 -2970
rect 4505 -3000 4520 -2970
rect 4460 -3040 4520 -3000
rect 4460 -3070 4475 -3040
rect 4505 -3070 4520 -3040
rect 4460 -3110 4520 -3070
rect 4460 -3140 4475 -3110
rect 4505 -3140 4520 -3110
rect 4460 -3180 4520 -3140
rect 4460 -3210 4475 -3180
rect 4505 -3210 4520 -3180
rect 4460 -3245 4520 -3210
rect 4460 -3275 4475 -3245
rect 4505 -3275 4520 -3245
rect 4460 -3305 4520 -3275
rect 4460 -3335 4475 -3305
rect 4505 -3335 4520 -3305
rect 4460 -3370 4520 -3335
rect 4460 -3400 4475 -3370
rect 4505 -3400 4520 -3370
rect 4460 -3440 4520 -3400
rect 4460 -3470 4475 -3440
rect 4505 -3470 4520 -3440
rect 4460 -3510 4520 -3470
rect 4460 -3540 4475 -3510
rect 4505 -3540 4520 -3510
rect 4460 -3580 4520 -3540
rect 4460 -3610 4475 -3580
rect 4505 -3610 4520 -3580
rect 4460 -3645 4520 -3610
rect 4460 -3675 4475 -3645
rect 4505 -3675 4520 -3645
rect 4460 -3705 4520 -3675
rect 4460 -3735 4475 -3705
rect 4505 -3735 4520 -3705
rect 4460 -3770 4520 -3735
rect 4460 -3800 4475 -3770
rect 4505 -3800 4520 -3770
rect 4460 -3840 4520 -3800
rect 4460 -3870 4475 -3840
rect 4505 -3870 4520 -3840
rect 4460 -3910 4520 -3870
rect 4460 -3940 4475 -3910
rect 4505 -3940 4520 -3910
rect 4460 -3980 4520 -3940
rect 4460 -4010 4475 -3980
rect 4505 -4010 4520 -3980
rect 4460 -4045 4520 -4010
rect 4460 -4075 4475 -4045
rect 4505 -4075 4520 -4045
rect 4460 -4105 4520 -4075
rect 4460 -4135 4475 -4105
rect 4505 -4135 4520 -4105
rect 4460 -4170 4520 -4135
rect 4460 -4200 4475 -4170
rect 4505 -4200 4520 -4170
rect 4460 -4240 4520 -4200
rect 4460 -4270 4475 -4240
rect 4505 -4270 4520 -4240
rect 4460 -4310 4520 -4270
rect 4460 -4340 4475 -4310
rect 4505 -4340 4520 -4310
rect 4460 -4380 4520 -4340
rect 4460 -4410 4475 -4380
rect 4505 -4410 4520 -4380
rect 4460 -4445 4520 -4410
rect 4460 -4475 4475 -4445
rect 4505 -4475 4520 -4445
rect 4460 -4490 4520 -4475
rect 4810 -1305 4870 -1290
rect 4810 -1335 4825 -1305
rect 4855 -1335 4870 -1305
rect 4810 -1370 4870 -1335
rect 4810 -1400 4825 -1370
rect 4855 -1400 4870 -1370
rect 4810 -1440 4870 -1400
rect 4810 -1470 4825 -1440
rect 4855 -1470 4870 -1440
rect 4810 -1510 4870 -1470
rect 4810 -1540 4825 -1510
rect 4855 -1540 4870 -1510
rect 4810 -1580 4870 -1540
rect 4810 -1610 4825 -1580
rect 4855 -1610 4870 -1580
rect 4810 -1645 4870 -1610
rect 4810 -1675 4825 -1645
rect 4855 -1675 4870 -1645
rect 4810 -1705 4870 -1675
rect 4810 -1735 4825 -1705
rect 4855 -1735 4870 -1705
rect 4810 -1770 4870 -1735
rect 4810 -1800 4825 -1770
rect 4855 -1800 4870 -1770
rect 4810 -1840 4870 -1800
rect 4810 -1870 4825 -1840
rect 4855 -1870 4870 -1840
rect 4810 -1910 4870 -1870
rect 4810 -1940 4825 -1910
rect 4855 -1940 4870 -1910
rect 4810 -1980 4870 -1940
rect 4810 -2010 4825 -1980
rect 4855 -2010 4870 -1980
rect 4810 -2045 4870 -2010
rect 4810 -2075 4825 -2045
rect 4855 -2075 4870 -2045
rect 4810 -2105 4870 -2075
rect 4810 -2135 4825 -2105
rect 4855 -2135 4870 -2105
rect 4810 -2170 4870 -2135
rect 4810 -2200 4825 -2170
rect 4855 -2200 4870 -2170
rect 4810 -2240 4870 -2200
rect 4810 -2270 4825 -2240
rect 4855 -2270 4870 -2240
rect 4810 -2310 4870 -2270
rect 4810 -2340 4825 -2310
rect 4855 -2340 4870 -2310
rect 4810 -2380 4870 -2340
rect 4810 -2410 4825 -2380
rect 4855 -2410 4870 -2380
rect 4810 -2445 4870 -2410
rect 4810 -2475 4825 -2445
rect 4855 -2475 4870 -2445
rect 4810 -2505 4870 -2475
rect 4810 -2535 4825 -2505
rect 4855 -2535 4870 -2505
rect 4810 -2570 4870 -2535
rect 4810 -2600 4825 -2570
rect 4855 -2600 4870 -2570
rect 4810 -2640 4870 -2600
rect 4810 -2670 4825 -2640
rect 4855 -2670 4870 -2640
rect 4810 -2710 4870 -2670
rect 4810 -2740 4825 -2710
rect 4855 -2740 4870 -2710
rect 4810 -2780 4870 -2740
rect 4810 -2810 4825 -2780
rect 4855 -2810 4870 -2780
rect 4810 -2845 4870 -2810
rect 4810 -2875 4825 -2845
rect 4855 -2875 4870 -2845
rect 4810 -2905 4870 -2875
rect 4810 -2935 4825 -2905
rect 4855 -2935 4870 -2905
rect 4810 -2970 4870 -2935
rect 4810 -3000 4825 -2970
rect 4855 -3000 4870 -2970
rect 4810 -3040 4870 -3000
rect 4810 -3070 4825 -3040
rect 4855 -3070 4870 -3040
rect 4810 -3110 4870 -3070
rect 4810 -3140 4825 -3110
rect 4855 -3140 4870 -3110
rect 4810 -3180 4870 -3140
rect 4810 -3210 4825 -3180
rect 4855 -3210 4870 -3180
rect 4810 -3245 4870 -3210
rect 4810 -3275 4825 -3245
rect 4855 -3275 4870 -3245
rect 4810 -3305 4870 -3275
rect 4810 -3335 4825 -3305
rect 4855 -3335 4870 -3305
rect 4810 -3370 4870 -3335
rect 4810 -3400 4825 -3370
rect 4855 -3400 4870 -3370
rect 4810 -3440 4870 -3400
rect 4810 -3470 4825 -3440
rect 4855 -3470 4870 -3440
rect 4810 -3510 4870 -3470
rect 4810 -3540 4825 -3510
rect 4855 -3540 4870 -3510
rect 4810 -3580 4870 -3540
rect 4810 -3610 4825 -3580
rect 4855 -3610 4870 -3580
rect 4810 -3645 4870 -3610
rect 4810 -3675 4825 -3645
rect 4855 -3675 4870 -3645
rect 4810 -3705 4870 -3675
rect 4810 -3735 4825 -3705
rect 4855 -3735 4870 -3705
rect 4810 -3770 4870 -3735
rect 4810 -3800 4825 -3770
rect 4855 -3800 4870 -3770
rect 4810 -3840 4870 -3800
rect 4810 -3870 4825 -3840
rect 4855 -3870 4870 -3840
rect 4810 -3910 4870 -3870
rect 4810 -3940 4825 -3910
rect 4855 -3940 4870 -3910
rect 4810 -3980 4870 -3940
rect 4810 -4010 4825 -3980
rect 4855 -4010 4870 -3980
rect 4810 -4045 4870 -4010
rect 4810 -4075 4825 -4045
rect 4855 -4075 4870 -4045
rect 4810 -4105 4870 -4075
rect 4810 -4135 4825 -4105
rect 4855 -4135 4870 -4105
rect 4810 -4170 4870 -4135
rect 4810 -4200 4825 -4170
rect 4855 -4200 4870 -4170
rect 4810 -4240 4870 -4200
rect 4810 -4270 4825 -4240
rect 4855 -4270 4870 -4240
rect 4810 -4310 4870 -4270
rect 4810 -4340 4825 -4310
rect 4855 -4340 4870 -4310
rect 4810 -4380 4870 -4340
rect 4810 -4410 4825 -4380
rect 4855 -4410 4870 -4380
rect 4810 -4445 4870 -4410
rect 4810 -4475 4825 -4445
rect 4855 -4475 4870 -4445
rect 4810 -4490 4870 -4475
rect 5160 -1305 5220 -1290
rect 5160 -1335 5175 -1305
rect 5205 -1335 5220 -1305
rect 5160 -1370 5220 -1335
rect 5160 -1400 5175 -1370
rect 5205 -1400 5220 -1370
rect 5160 -1440 5220 -1400
rect 5160 -1470 5175 -1440
rect 5205 -1470 5220 -1440
rect 5160 -1510 5220 -1470
rect 5160 -1540 5175 -1510
rect 5205 -1540 5220 -1510
rect 5160 -1580 5220 -1540
rect 5160 -1610 5175 -1580
rect 5205 -1610 5220 -1580
rect 5160 -1645 5220 -1610
rect 5160 -1675 5175 -1645
rect 5205 -1675 5220 -1645
rect 5160 -1705 5220 -1675
rect 5160 -1735 5175 -1705
rect 5205 -1735 5220 -1705
rect 5160 -1770 5220 -1735
rect 5160 -1800 5175 -1770
rect 5205 -1800 5220 -1770
rect 5160 -1840 5220 -1800
rect 5160 -1870 5175 -1840
rect 5205 -1870 5220 -1840
rect 5160 -1910 5220 -1870
rect 5160 -1940 5175 -1910
rect 5205 -1940 5220 -1910
rect 5160 -1980 5220 -1940
rect 5160 -2010 5175 -1980
rect 5205 -2010 5220 -1980
rect 5160 -2045 5220 -2010
rect 5160 -2075 5175 -2045
rect 5205 -2075 5220 -2045
rect 5160 -2105 5220 -2075
rect 5160 -2135 5175 -2105
rect 5205 -2135 5220 -2105
rect 5160 -2170 5220 -2135
rect 5160 -2200 5175 -2170
rect 5205 -2200 5220 -2170
rect 5160 -2240 5220 -2200
rect 5160 -2270 5175 -2240
rect 5205 -2270 5220 -2240
rect 5160 -2310 5220 -2270
rect 5160 -2340 5175 -2310
rect 5205 -2340 5220 -2310
rect 5160 -2380 5220 -2340
rect 5160 -2410 5175 -2380
rect 5205 -2410 5220 -2380
rect 5160 -2445 5220 -2410
rect 5160 -2475 5175 -2445
rect 5205 -2475 5220 -2445
rect 5160 -2505 5220 -2475
rect 5160 -2535 5175 -2505
rect 5205 -2535 5220 -2505
rect 5160 -2570 5220 -2535
rect 5160 -2600 5175 -2570
rect 5205 -2600 5220 -2570
rect 5160 -2640 5220 -2600
rect 5160 -2670 5175 -2640
rect 5205 -2670 5220 -2640
rect 5160 -2710 5220 -2670
rect 5160 -2740 5175 -2710
rect 5205 -2740 5220 -2710
rect 5160 -2780 5220 -2740
rect 5160 -2810 5175 -2780
rect 5205 -2810 5220 -2780
rect 5160 -2845 5220 -2810
rect 5160 -2875 5175 -2845
rect 5205 -2875 5220 -2845
rect 5160 -2905 5220 -2875
rect 5160 -2935 5175 -2905
rect 5205 -2935 5220 -2905
rect 5160 -2970 5220 -2935
rect 5160 -3000 5175 -2970
rect 5205 -3000 5220 -2970
rect 5160 -3040 5220 -3000
rect 5160 -3070 5175 -3040
rect 5205 -3070 5220 -3040
rect 5160 -3110 5220 -3070
rect 5160 -3140 5175 -3110
rect 5205 -3140 5220 -3110
rect 5160 -3180 5220 -3140
rect 5160 -3210 5175 -3180
rect 5205 -3210 5220 -3180
rect 5160 -3245 5220 -3210
rect 5160 -3275 5175 -3245
rect 5205 -3275 5220 -3245
rect 5160 -3305 5220 -3275
rect 5160 -3335 5175 -3305
rect 5205 -3335 5220 -3305
rect 5160 -3370 5220 -3335
rect 5160 -3400 5175 -3370
rect 5205 -3400 5220 -3370
rect 5160 -3440 5220 -3400
rect 5160 -3470 5175 -3440
rect 5205 -3470 5220 -3440
rect 5160 -3510 5220 -3470
rect 5160 -3540 5175 -3510
rect 5205 -3540 5220 -3510
rect 5160 -3580 5220 -3540
rect 5160 -3610 5175 -3580
rect 5205 -3610 5220 -3580
rect 5160 -3645 5220 -3610
rect 5160 -3675 5175 -3645
rect 5205 -3675 5220 -3645
rect 5160 -3705 5220 -3675
rect 5160 -3735 5175 -3705
rect 5205 -3735 5220 -3705
rect 5160 -3770 5220 -3735
rect 5160 -3800 5175 -3770
rect 5205 -3800 5220 -3770
rect 5160 -3840 5220 -3800
rect 5160 -3870 5175 -3840
rect 5205 -3870 5220 -3840
rect 5160 -3910 5220 -3870
rect 5160 -3940 5175 -3910
rect 5205 -3940 5220 -3910
rect 5160 -3980 5220 -3940
rect 5160 -4010 5175 -3980
rect 5205 -4010 5220 -3980
rect 5160 -4045 5220 -4010
rect 5160 -4075 5175 -4045
rect 5205 -4075 5220 -4045
rect 5160 -4105 5220 -4075
rect 5160 -4135 5175 -4105
rect 5205 -4135 5220 -4105
rect 5160 -4170 5220 -4135
rect 5160 -4200 5175 -4170
rect 5205 -4200 5220 -4170
rect 5160 -4240 5220 -4200
rect 5160 -4270 5175 -4240
rect 5205 -4270 5220 -4240
rect 5160 -4310 5220 -4270
rect 5160 -4340 5175 -4310
rect 5205 -4340 5220 -4310
rect 5160 -4380 5220 -4340
rect 5160 -4410 5175 -4380
rect 5205 -4410 5220 -4380
rect 5160 -4445 5220 -4410
rect 5160 -4475 5175 -4445
rect 5205 -4475 5220 -4445
rect 5160 -4490 5220 -4475
rect 5510 -1305 5570 -1290
rect 5510 -1335 5525 -1305
rect 5555 -1335 5570 -1305
rect 5510 -1370 5570 -1335
rect 5510 -1400 5525 -1370
rect 5555 -1400 5570 -1370
rect 5510 -1440 5570 -1400
rect 5510 -1470 5525 -1440
rect 5555 -1470 5570 -1440
rect 5510 -1510 5570 -1470
rect 5510 -1540 5525 -1510
rect 5555 -1540 5570 -1510
rect 5510 -1580 5570 -1540
rect 5510 -1610 5525 -1580
rect 5555 -1610 5570 -1580
rect 5510 -1645 5570 -1610
rect 5510 -1675 5525 -1645
rect 5555 -1675 5570 -1645
rect 5510 -1705 5570 -1675
rect 5510 -1735 5525 -1705
rect 5555 -1735 5570 -1705
rect 5510 -1770 5570 -1735
rect 5510 -1800 5525 -1770
rect 5555 -1800 5570 -1770
rect 5510 -1840 5570 -1800
rect 5510 -1870 5525 -1840
rect 5555 -1870 5570 -1840
rect 5510 -1910 5570 -1870
rect 5510 -1940 5525 -1910
rect 5555 -1940 5570 -1910
rect 5510 -1980 5570 -1940
rect 5510 -2010 5525 -1980
rect 5555 -2010 5570 -1980
rect 5510 -2045 5570 -2010
rect 5510 -2075 5525 -2045
rect 5555 -2075 5570 -2045
rect 5510 -2105 5570 -2075
rect 5510 -2135 5525 -2105
rect 5555 -2135 5570 -2105
rect 5510 -2170 5570 -2135
rect 5510 -2200 5525 -2170
rect 5555 -2200 5570 -2170
rect 5510 -2240 5570 -2200
rect 5510 -2270 5525 -2240
rect 5555 -2270 5570 -2240
rect 5510 -2310 5570 -2270
rect 5510 -2340 5525 -2310
rect 5555 -2340 5570 -2310
rect 5510 -2380 5570 -2340
rect 5510 -2410 5525 -2380
rect 5555 -2410 5570 -2380
rect 5510 -2445 5570 -2410
rect 5510 -2475 5525 -2445
rect 5555 -2475 5570 -2445
rect 5510 -2505 5570 -2475
rect 5510 -2535 5525 -2505
rect 5555 -2535 5570 -2505
rect 5510 -2570 5570 -2535
rect 5510 -2600 5525 -2570
rect 5555 -2600 5570 -2570
rect 5510 -2640 5570 -2600
rect 5510 -2670 5525 -2640
rect 5555 -2670 5570 -2640
rect 5510 -2710 5570 -2670
rect 5510 -2740 5525 -2710
rect 5555 -2740 5570 -2710
rect 5510 -2780 5570 -2740
rect 5510 -2810 5525 -2780
rect 5555 -2810 5570 -2780
rect 5510 -2845 5570 -2810
rect 5510 -2875 5525 -2845
rect 5555 -2875 5570 -2845
rect 5510 -2905 5570 -2875
rect 5510 -2935 5525 -2905
rect 5555 -2935 5570 -2905
rect 5510 -2970 5570 -2935
rect 5510 -3000 5525 -2970
rect 5555 -3000 5570 -2970
rect 5510 -3040 5570 -3000
rect 5510 -3070 5525 -3040
rect 5555 -3070 5570 -3040
rect 5510 -3110 5570 -3070
rect 5510 -3140 5525 -3110
rect 5555 -3140 5570 -3110
rect 5510 -3180 5570 -3140
rect 5510 -3210 5525 -3180
rect 5555 -3210 5570 -3180
rect 5510 -3245 5570 -3210
rect 5510 -3275 5525 -3245
rect 5555 -3275 5570 -3245
rect 5510 -3305 5570 -3275
rect 5510 -3335 5525 -3305
rect 5555 -3335 5570 -3305
rect 5510 -3370 5570 -3335
rect 5510 -3400 5525 -3370
rect 5555 -3400 5570 -3370
rect 5510 -3440 5570 -3400
rect 5510 -3470 5525 -3440
rect 5555 -3470 5570 -3440
rect 5510 -3510 5570 -3470
rect 5510 -3540 5525 -3510
rect 5555 -3540 5570 -3510
rect 5510 -3580 5570 -3540
rect 5510 -3610 5525 -3580
rect 5555 -3610 5570 -3580
rect 5510 -3645 5570 -3610
rect 5510 -3675 5525 -3645
rect 5555 -3675 5570 -3645
rect 5510 -3705 5570 -3675
rect 5510 -3735 5525 -3705
rect 5555 -3735 5570 -3705
rect 5510 -3770 5570 -3735
rect 5510 -3800 5525 -3770
rect 5555 -3800 5570 -3770
rect 5510 -3840 5570 -3800
rect 5510 -3870 5525 -3840
rect 5555 -3870 5570 -3840
rect 5510 -3910 5570 -3870
rect 5510 -3940 5525 -3910
rect 5555 -3940 5570 -3910
rect 5510 -3980 5570 -3940
rect 5510 -4010 5525 -3980
rect 5555 -4010 5570 -3980
rect 5510 -4045 5570 -4010
rect 5510 -4075 5525 -4045
rect 5555 -4075 5570 -4045
rect 5510 -4105 5570 -4075
rect 5510 -4135 5525 -4105
rect 5555 -4135 5570 -4105
rect 5510 -4170 5570 -4135
rect 5510 -4200 5525 -4170
rect 5555 -4200 5570 -4170
rect 5510 -4240 5570 -4200
rect 5510 -4270 5525 -4240
rect 5555 -4270 5570 -4240
rect 5510 -4310 5570 -4270
rect 5510 -4340 5525 -4310
rect 5555 -4340 5570 -4310
rect 5510 -4380 5570 -4340
rect 5510 -4410 5525 -4380
rect 5555 -4410 5570 -4380
rect 5510 -4445 5570 -4410
rect 5510 -4475 5525 -4445
rect 5555 -4475 5570 -4445
rect 5510 -4490 5570 -4475
rect 5860 -1305 5920 -1290
rect 5860 -1335 5875 -1305
rect 5905 -1335 5920 -1305
rect 5860 -1370 5920 -1335
rect 5860 -1400 5875 -1370
rect 5905 -1400 5920 -1370
rect 5860 -1440 5920 -1400
rect 5860 -1470 5875 -1440
rect 5905 -1470 5920 -1440
rect 5860 -1510 5920 -1470
rect 5860 -1540 5875 -1510
rect 5905 -1540 5920 -1510
rect 5860 -1580 5920 -1540
rect 5860 -1610 5875 -1580
rect 5905 -1610 5920 -1580
rect 5860 -1645 5920 -1610
rect 5860 -1675 5875 -1645
rect 5905 -1675 5920 -1645
rect 5860 -1705 5920 -1675
rect 5860 -1735 5875 -1705
rect 5905 -1735 5920 -1705
rect 5860 -1770 5920 -1735
rect 5860 -1800 5875 -1770
rect 5905 -1800 5920 -1770
rect 5860 -1840 5920 -1800
rect 5860 -1870 5875 -1840
rect 5905 -1870 5920 -1840
rect 5860 -1910 5920 -1870
rect 5860 -1940 5875 -1910
rect 5905 -1940 5920 -1910
rect 5860 -1980 5920 -1940
rect 5860 -2010 5875 -1980
rect 5905 -2010 5920 -1980
rect 5860 -2045 5920 -2010
rect 5860 -2075 5875 -2045
rect 5905 -2075 5920 -2045
rect 5860 -2105 5920 -2075
rect 5860 -2135 5875 -2105
rect 5905 -2135 5920 -2105
rect 5860 -2170 5920 -2135
rect 5860 -2200 5875 -2170
rect 5905 -2200 5920 -2170
rect 5860 -2240 5920 -2200
rect 5860 -2270 5875 -2240
rect 5905 -2270 5920 -2240
rect 5860 -2310 5920 -2270
rect 5860 -2340 5875 -2310
rect 5905 -2340 5920 -2310
rect 5860 -2380 5920 -2340
rect 5860 -2410 5875 -2380
rect 5905 -2410 5920 -2380
rect 5860 -2445 5920 -2410
rect 5860 -2475 5875 -2445
rect 5905 -2475 5920 -2445
rect 5860 -2505 5920 -2475
rect 5860 -2535 5875 -2505
rect 5905 -2535 5920 -2505
rect 5860 -2570 5920 -2535
rect 5860 -2600 5875 -2570
rect 5905 -2600 5920 -2570
rect 5860 -2640 5920 -2600
rect 5860 -2670 5875 -2640
rect 5905 -2670 5920 -2640
rect 5860 -2710 5920 -2670
rect 5860 -2740 5875 -2710
rect 5905 -2740 5920 -2710
rect 5860 -2780 5920 -2740
rect 5860 -2810 5875 -2780
rect 5905 -2810 5920 -2780
rect 5860 -2845 5920 -2810
rect 5860 -2875 5875 -2845
rect 5905 -2875 5920 -2845
rect 5860 -2905 5920 -2875
rect 5860 -2935 5875 -2905
rect 5905 -2935 5920 -2905
rect 5860 -2970 5920 -2935
rect 5860 -3000 5875 -2970
rect 5905 -3000 5920 -2970
rect 5860 -3040 5920 -3000
rect 5860 -3070 5875 -3040
rect 5905 -3070 5920 -3040
rect 5860 -3110 5920 -3070
rect 5860 -3140 5875 -3110
rect 5905 -3140 5920 -3110
rect 5860 -3180 5920 -3140
rect 5860 -3210 5875 -3180
rect 5905 -3210 5920 -3180
rect 5860 -3245 5920 -3210
rect 5860 -3275 5875 -3245
rect 5905 -3275 5920 -3245
rect 5860 -3305 5920 -3275
rect 5860 -3335 5875 -3305
rect 5905 -3335 5920 -3305
rect 5860 -3370 5920 -3335
rect 5860 -3400 5875 -3370
rect 5905 -3400 5920 -3370
rect 5860 -3440 5920 -3400
rect 5860 -3470 5875 -3440
rect 5905 -3470 5920 -3440
rect 5860 -3510 5920 -3470
rect 5860 -3540 5875 -3510
rect 5905 -3540 5920 -3510
rect 5860 -3580 5920 -3540
rect 5860 -3610 5875 -3580
rect 5905 -3610 5920 -3580
rect 5860 -3645 5920 -3610
rect 5860 -3675 5875 -3645
rect 5905 -3675 5920 -3645
rect 5860 -3705 5920 -3675
rect 5860 -3735 5875 -3705
rect 5905 -3735 5920 -3705
rect 5860 -3770 5920 -3735
rect 5860 -3800 5875 -3770
rect 5905 -3800 5920 -3770
rect 5860 -3840 5920 -3800
rect 5860 -3870 5875 -3840
rect 5905 -3870 5920 -3840
rect 5860 -3910 5920 -3870
rect 5860 -3940 5875 -3910
rect 5905 -3940 5920 -3910
rect 5860 -3980 5920 -3940
rect 5860 -4010 5875 -3980
rect 5905 -4010 5920 -3980
rect 5860 -4045 5920 -4010
rect 5860 -4075 5875 -4045
rect 5905 -4075 5920 -4045
rect 5860 -4105 5920 -4075
rect 5860 -4135 5875 -4105
rect 5905 -4135 5920 -4105
rect 5860 -4170 5920 -4135
rect 5860 -4200 5875 -4170
rect 5905 -4200 5920 -4170
rect 5860 -4240 5920 -4200
rect 5860 -4270 5875 -4240
rect 5905 -4270 5920 -4240
rect 5860 -4310 5920 -4270
rect 5860 -4340 5875 -4310
rect 5905 -4340 5920 -4310
rect 5860 -4380 5920 -4340
rect 5860 -4410 5875 -4380
rect 5905 -4410 5920 -4380
rect 5860 -4445 5920 -4410
rect 5860 -4475 5875 -4445
rect 5905 -4475 5920 -4445
rect 5860 -4490 5920 -4475
rect 6210 -1305 6270 -1290
rect 6210 -1335 6225 -1305
rect 6255 -1335 6270 -1305
rect 6210 -1370 6270 -1335
rect 6210 -1400 6225 -1370
rect 6255 -1400 6270 -1370
rect 6210 -1440 6270 -1400
rect 6210 -1470 6225 -1440
rect 6255 -1470 6270 -1440
rect 6210 -1510 6270 -1470
rect 6210 -1540 6225 -1510
rect 6255 -1540 6270 -1510
rect 6210 -1580 6270 -1540
rect 6210 -1610 6225 -1580
rect 6255 -1610 6270 -1580
rect 6210 -1645 6270 -1610
rect 6210 -1675 6225 -1645
rect 6255 -1675 6270 -1645
rect 6210 -1705 6270 -1675
rect 6210 -1735 6225 -1705
rect 6255 -1735 6270 -1705
rect 6210 -1770 6270 -1735
rect 6210 -1800 6225 -1770
rect 6255 -1800 6270 -1770
rect 6210 -1840 6270 -1800
rect 6210 -1870 6225 -1840
rect 6255 -1870 6270 -1840
rect 6210 -1910 6270 -1870
rect 6210 -1940 6225 -1910
rect 6255 -1940 6270 -1910
rect 6210 -1980 6270 -1940
rect 6210 -2010 6225 -1980
rect 6255 -2010 6270 -1980
rect 6210 -2045 6270 -2010
rect 6210 -2075 6225 -2045
rect 6255 -2075 6270 -2045
rect 6210 -2105 6270 -2075
rect 6210 -2135 6225 -2105
rect 6255 -2135 6270 -2105
rect 6210 -2170 6270 -2135
rect 6210 -2200 6225 -2170
rect 6255 -2200 6270 -2170
rect 6210 -2240 6270 -2200
rect 6210 -2270 6225 -2240
rect 6255 -2270 6270 -2240
rect 6210 -2310 6270 -2270
rect 6210 -2340 6225 -2310
rect 6255 -2340 6270 -2310
rect 6210 -2380 6270 -2340
rect 6210 -2410 6225 -2380
rect 6255 -2410 6270 -2380
rect 6210 -2445 6270 -2410
rect 6210 -2475 6225 -2445
rect 6255 -2475 6270 -2445
rect 6210 -2505 6270 -2475
rect 6210 -2535 6225 -2505
rect 6255 -2535 6270 -2505
rect 6210 -2570 6270 -2535
rect 6210 -2600 6225 -2570
rect 6255 -2600 6270 -2570
rect 6210 -2640 6270 -2600
rect 6210 -2670 6225 -2640
rect 6255 -2670 6270 -2640
rect 6210 -2710 6270 -2670
rect 6210 -2740 6225 -2710
rect 6255 -2740 6270 -2710
rect 6210 -2780 6270 -2740
rect 6210 -2810 6225 -2780
rect 6255 -2810 6270 -2780
rect 6210 -2845 6270 -2810
rect 6210 -2875 6225 -2845
rect 6255 -2875 6270 -2845
rect 6210 -2905 6270 -2875
rect 6210 -2935 6225 -2905
rect 6255 -2935 6270 -2905
rect 6210 -2970 6270 -2935
rect 6210 -3000 6225 -2970
rect 6255 -3000 6270 -2970
rect 6210 -3040 6270 -3000
rect 6210 -3070 6225 -3040
rect 6255 -3070 6270 -3040
rect 6210 -3110 6270 -3070
rect 6210 -3140 6225 -3110
rect 6255 -3140 6270 -3110
rect 6210 -3180 6270 -3140
rect 6210 -3210 6225 -3180
rect 6255 -3210 6270 -3180
rect 6210 -3245 6270 -3210
rect 6210 -3275 6225 -3245
rect 6255 -3275 6270 -3245
rect 6210 -3305 6270 -3275
rect 6210 -3335 6225 -3305
rect 6255 -3335 6270 -3305
rect 6210 -3370 6270 -3335
rect 6210 -3400 6225 -3370
rect 6255 -3400 6270 -3370
rect 6210 -3440 6270 -3400
rect 6210 -3470 6225 -3440
rect 6255 -3470 6270 -3440
rect 6210 -3510 6270 -3470
rect 6210 -3540 6225 -3510
rect 6255 -3540 6270 -3510
rect 6210 -3580 6270 -3540
rect 6210 -3610 6225 -3580
rect 6255 -3610 6270 -3580
rect 6210 -3645 6270 -3610
rect 6210 -3675 6225 -3645
rect 6255 -3675 6270 -3645
rect 6210 -3705 6270 -3675
rect 6210 -3735 6225 -3705
rect 6255 -3735 6270 -3705
rect 6210 -3770 6270 -3735
rect 6210 -3800 6225 -3770
rect 6255 -3800 6270 -3770
rect 6210 -3840 6270 -3800
rect 6210 -3870 6225 -3840
rect 6255 -3870 6270 -3840
rect 6210 -3910 6270 -3870
rect 6210 -3940 6225 -3910
rect 6255 -3940 6270 -3910
rect 6210 -3980 6270 -3940
rect 6210 -4010 6225 -3980
rect 6255 -4010 6270 -3980
rect 6210 -4045 6270 -4010
rect 6210 -4075 6225 -4045
rect 6255 -4075 6270 -4045
rect 6210 -4105 6270 -4075
rect 6210 -4135 6225 -4105
rect 6255 -4135 6270 -4105
rect 6210 -4170 6270 -4135
rect 6210 -4200 6225 -4170
rect 6255 -4200 6270 -4170
rect 6210 -4240 6270 -4200
rect 6210 -4270 6225 -4240
rect 6255 -4270 6270 -4240
rect 6210 -4310 6270 -4270
rect 6210 -4340 6225 -4310
rect 6255 -4340 6270 -4310
rect 6210 -4380 6270 -4340
rect 6210 -4410 6225 -4380
rect 6255 -4410 6270 -4380
rect 6210 -4445 6270 -4410
rect 6210 -4475 6225 -4445
rect 6255 -4475 6270 -4445
rect 6210 -4490 6270 -4475
rect 6560 -1305 6620 -1290
rect 6560 -1335 6575 -1305
rect 6605 -1335 6620 -1305
rect 6560 -1370 6620 -1335
rect 6560 -1400 6575 -1370
rect 6605 -1400 6620 -1370
rect 6560 -1440 6620 -1400
rect 6560 -1470 6575 -1440
rect 6605 -1470 6620 -1440
rect 6560 -1510 6620 -1470
rect 6560 -1540 6575 -1510
rect 6605 -1540 6620 -1510
rect 6560 -1580 6620 -1540
rect 6560 -1610 6575 -1580
rect 6605 -1610 6620 -1580
rect 6560 -1645 6620 -1610
rect 6560 -1675 6575 -1645
rect 6605 -1675 6620 -1645
rect 6560 -1705 6620 -1675
rect 6560 -1735 6575 -1705
rect 6605 -1735 6620 -1705
rect 6560 -1770 6620 -1735
rect 6560 -1800 6575 -1770
rect 6605 -1800 6620 -1770
rect 6560 -1840 6620 -1800
rect 6560 -1870 6575 -1840
rect 6605 -1870 6620 -1840
rect 6560 -1910 6620 -1870
rect 6560 -1940 6575 -1910
rect 6605 -1940 6620 -1910
rect 6560 -1980 6620 -1940
rect 6560 -2010 6575 -1980
rect 6605 -2010 6620 -1980
rect 6560 -2045 6620 -2010
rect 6560 -2075 6575 -2045
rect 6605 -2075 6620 -2045
rect 6560 -2105 6620 -2075
rect 6560 -2135 6575 -2105
rect 6605 -2135 6620 -2105
rect 6560 -2170 6620 -2135
rect 6560 -2200 6575 -2170
rect 6605 -2200 6620 -2170
rect 6560 -2240 6620 -2200
rect 6560 -2270 6575 -2240
rect 6605 -2270 6620 -2240
rect 6560 -2310 6620 -2270
rect 6560 -2340 6575 -2310
rect 6605 -2340 6620 -2310
rect 6560 -2380 6620 -2340
rect 6560 -2410 6575 -2380
rect 6605 -2410 6620 -2380
rect 6560 -2445 6620 -2410
rect 6560 -2475 6575 -2445
rect 6605 -2475 6620 -2445
rect 6560 -2505 6620 -2475
rect 6560 -2535 6575 -2505
rect 6605 -2535 6620 -2505
rect 6560 -2570 6620 -2535
rect 6560 -2600 6575 -2570
rect 6605 -2600 6620 -2570
rect 6560 -2640 6620 -2600
rect 6560 -2670 6575 -2640
rect 6605 -2670 6620 -2640
rect 6560 -2710 6620 -2670
rect 6560 -2740 6575 -2710
rect 6605 -2740 6620 -2710
rect 6560 -2780 6620 -2740
rect 6560 -2810 6575 -2780
rect 6605 -2810 6620 -2780
rect 6560 -2845 6620 -2810
rect 6560 -2875 6575 -2845
rect 6605 -2875 6620 -2845
rect 6560 -2905 6620 -2875
rect 6560 -2935 6575 -2905
rect 6605 -2935 6620 -2905
rect 6560 -2970 6620 -2935
rect 6560 -3000 6575 -2970
rect 6605 -3000 6620 -2970
rect 6560 -3040 6620 -3000
rect 6560 -3070 6575 -3040
rect 6605 -3070 6620 -3040
rect 6560 -3110 6620 -3070
rect 6560 -3140 6575 -3110
rect 6605 -3140 6620 -3110
rect 6560 -3180 6620 -3140
rect 6560 -3210 6575 -3180
rect 6605 -3210 6620 -3180
rect 6560 -3245 6620 -3210
rect 6560 -3275 6575 -3245
rect 6605 -3275 6620 -3245
rect 6560 -3305 6620 -3275
rect 6560 -3335 6575 -3305
rect 6605 -3335 6620 -3305
rect 6560 -3370 6620 -3335
rect 6560 -3400 6575 -3370
rect 6605 -3400 6620 -3370
rect 6560 -3440 6620 -3400
rect 6560 -3470 6575 -3440
rect 6605 -3470 6620 -3440
rect 6560 -3510 6620 -3470
rect 6560 -3540 6575 -3510
rect 6605 -3540 6620 -3510
rect 6560 -3580 6620 -3540
rect 6560 -3610 6575 -3580
rect 6605 -3610 6620 -3580
rect 6560 -3645 6620 -3610
rect 6560 -3675 6575 -3645
rect 6605 -3675 6620 -3645
rect 6560 -3705 6620 -3675
rect 6560 -3735 6575 -3705
rect 6605 -3735 6620 -3705
rect 6560 -3770 6620 -3735
rect 6560 -3800 6575 -3770
rect 6605 -3800 6620 -3770
rect 6560 -3840 6620 -3800
rect 6560 -3870 6575 -3840
rect 6605 -3870 6620 -3840
rect 6560 -3910 6620 -3870
rect 6560 -3940 6575 -3910
rect 6605 -3940 6620 -3910
rect 6560 -3980 6620 -3940
rect 6560 -4010 6575 -3980
rect 6605 -4010 6620 -3980
rect 6560 -4045 6620 -4010
rect 6560 -4075 6575 -4045
rect 6605 -4075 6620 -4045
rect 6560 -4105 6620 -4075
rect 6560 -4135 6575 -4105
rect 6605 -4135 6620 -4105
rect 6560 -4170 6620 -4135
rect 6560 -4200 6575 -4170
rect 6605 -4200 6620 -4170
rect 6560 -4240 6620 -4200
rect 6560 -4270 6575 -4240
rect 6605 -4270 6620 -4240
rect 6560 -4310 6620 -4270
rect 6560 -4340 6575 -4310
rect 6605 -4340 6620 -4310
rect 6560 -4380 6620 -4340
rect 6560 -4410 6575 -4380
rect 6605 -4410 6620 -4380
rect 6560 -4445 6620 -4410
rect 6560 -4475 6575 -4445
rect 6605 -4475 6620 -4445
rect 6560 -4490 6620 -4475
rect 6910 -1305 6970 -1290
rect 6910 -1335 6925 -1305
rect 6955 -1335 6970 -1305
rect 6910 -1370 6970 -1335
rect 6910 -1400 6925 -1370
rect 6955 -1400 6970 -1370
rect 6910 -1440 6970 -1400
rect 6910 -1470 6925 -1440
rect 6955 -1470 6970 -1440
rect 6910 -1510 6970 -1470
rect 6910 -1540 6925 -1510
rect 6955 -1540 6970 -1510
rect 6910 -1580 6970 -1540
rect 6910 -1610 6925 -1580
rect 6955 -1610 6970 -1580
rect 6910 -1645 6970 -1610
rect 6910 -1675 6925 -1645
rect 6955 -1675 6970 -1645
rect 6910 -1705 6970 -1675
rect 6910 -1735 6925 -1705
rect 6955 -1735 6970 -1705
rect 6910 -1770 6970 -1735
rect 6910 -1800 6925 -1770
rect 6955 -1800 6970 -1770
rect 6910 -1840 6970 -1800
rect 6910 -1870 6925 -1840
rect 6955 -1870 6970 -1840
rect 6910 -1910 6970 -1870
rect 6910 -1940 6925 -1910
rect 6955 -1940 6970 -1910
rect 6910 -1980 6970 -1940
rect 6910 -2010 6925 -1980
rect 6955 -2010 6970 -1980
rect 6910 -2045 6970 -2010
rect 6910 -2075 6925 -2045
rect 6955 -2075 6970 -2045
rect 6910 -2105 6970 -2075
rect 6910 -2135 6925 -2105
rect 6955 -2135 6970 -2105
rect 6910 -2170 6970 -2135
rect 6910 -2200 6925 -2170
rect 6955 -2200 6970 -2170
rect 6910 -2240 6970 -2200
rect 6910 -2270 6925 -2240
rect 6955 -2270 6970 -2240
rect 6910 -2310 6970 -2270
rect 6910 -2340 6925 -2310
rect 6955 -2340 6970 -2310
rect 6910 -2380 6970 -2340
rect 6910 -2410 6925 -2380
rect 6955 -2410 6970 -2380
rect 6910 -2445 6970 -2410
rect 6910 -2475 6925 -2445
rect 6955 -2475 6970 -2445
rect 6910 -2505 6970 -2475
rect 6910 -2535 6925 -2505
rect 6955 -2535 6970 -2505
rect 6910 -2570 6970 -2535
rect 6910 -2600 6925 -2570
rect 6955 -2600 6970 -2570
rect 6910 -2640 6970 -2600
rect 6910 -2670 6925 -2640
rect 6955 -2670 6970 -2640
rect 6910 -2710 6970 -2670
rect 6910 -2740 6925 -2710
rect 6955 -2740 6970 -2710
rect 6910 -2780 6970 -2740
rect 6910 -2810 6925 -2780
rect 6955 -2810 6970 -2780
rect 6910 -2845 6970 -2810
rect 6910 -2875 6925 -2845
rect 6955 -2875 6970 -2845
rect 6910 -2905 6970 -2875
rect 6910 -2935 6925 -2905
rect 6955 -2935 6970 -2905
rect 6910 -2970 6970 -2935
rect 6910 -3000 6925 -2970
rect 6955 -3000 6970 -2970
rect 6910 -3040 6970 -3000
rect 6910 -3070 6925 -3040
rect 6955 -3070 6970 -3040
rect 6910 -3110 6970 -3070
rect 6910 -3140 6925 -3110
rect 6955 -3140 6970 -3110
rect 6910 -3180 6970 -3140
rect 6910 -3210 6925 -3180
rect 6955 -3210 6970 -3180
rect 6910 -3245 6970 -3210
rect 6910 -3275 6925 -3245
rect 6955 -3275 6970 -3245
rect 6910 -3305 6970 -3275
rect 6910 -3335 6925 -3305
rect 6955 -3335 6970 -3305
rect 6910 -3370 6970 -3335
rect 6910 -3400 6925 -3370
rect 6955 -3400 6970 -3370
rect 6910 -3440 6970 -3400
rect 6910 -3470 6925 -3440
rect 6955 -3470 6970 -3440
rect 6910 -3510 6970 -3470
rect 6910 -3540 6925 -3510
rect 6955 -3540 6970 -3510
rect 6910 -3580 6970 -3540
rect 6910 -3610 6925 -3580
rect 6955 -3610 6970 -3580
rect 6910 -3645 6970 -3610
rect 6910 -3675 6925 -3645
rect 6955 -3675 6970 -3645
rect 6910 -3705 6970 -3675
rect 6910 -3735 6925 -3705
rect 6955 -3735 6970 -3705
rect 6910 -3770 6970 -3735
rect 6910 -3800 6925 -3770
rect 6955 -3800 6970 -3770
rect 6910 -3840 6970 -3800
rect 6910 -3870 6925 -3840
rect 6955 -3870 6970 -3840
rect 6910 -3910 6970 -3870
rect 6910 -3940 6925 -3910
rect 6955 -3940 6970 -3910
rect 6910 -3980 6970 -3940
rect 6910 -4010 6925 -3980
rect 6955 -4010 6970 -3980
rect 6910 -4045 6970 -4010
rect 6910 -4075 6925 -4045
rect 6955 -4075 6970 -4045
rect 6910 -4105 6970 -4075
rect 6910 -4135 6925 -4105
rect 6955 -4135 6970 -4105
rect 6910 -4170 6970 -4135
rect 6910 -4200 6925 -4170
rect 6955 -4200 6970 -4170
rect 6910 -4240 6970 -4200
rect 6910 -4270 6925 -4240
rect 6955 -4270 6970 -4240
rect 6910 -4310 6970 -4270
rect 6910 -4340 6925 -4310
rect 6955 -4340 6970 -4310
rect 6910 -4380 6970 -4340
rect 6910 -4410 6925 -4380
rect 6955 -4410 6970 -4380
rect 6910 -4445 6970 -4410
rect 6910 -4475 6925 -4445
rect 6955 -4475 6970 -4445
rect 6910 -4490 6970 -4475
rect 7260 -1305 7320 -1290
rect 7260 -1335 7275 -1305
rect 7305 -1335 7320 -1305
rect 7260 -1370 7320 -1335
rect 7260 -1400 7275 -1370
rect 7305 -1400 7320 -1370
rect 7260 -1440 7320 -1400
rect 7260 -1470 7275 -1440
rect 7305 -1470 7320 -1440
rect 7260 -1510 7320 -1470
rect 7260 -1540 7275 -1510
rect 7305 -1540 7320 -1510
rect 7260 -1580 7320 -1540
rect 7260 -1610 7275 -1580
rect 7305 -1610 7320 -1580
rect 7260 -1645 7320 -1610
rect 7260 -1675 7275 -1645
rect 7305 -1675 7320 -1645
rect 7260 -1705 7320 -1675
rect 7260 -1735 7275 -1705
rect 7305 -1735 7320 -1705
rect 7260 -1770 7320 -1735
rect 7260 -1800 7275 -1770
rect 7305 -1800 7320 -1770
rect 7260 -1840 7320 -1800
rect 7260 -1870 7275 -1840
rect 7305 -1870 7320 -1840
rect 7260 -1910 7320 -1870
rect 7260 -1940 7275 -1910
rect 7305 -1940 7320 -1910
rect 7260 -1980 7320 -1940
rect 7260 -2010 7275 -1980
rect 7305 -2010 7320 -1980
rect 7260 -2045 7320 -2010
rect 7260 -2075 7275 -2045
rect 7305 -2075 7320 -2045
rect 7260 -2105 7320 -2075
rect 7260 -2135 7275 -2105
rect 7305 -2135 7320 -2105
rect 7260 -2170 7320 -2135
rect 7260 -2200 7275 -2170
rect 7305 -2200 7320 -2170
rect 7260 -2240 7320 -2200
rect 7260 -2270 7275 -2240
rect 7305 -2270 7320 -2240
rect 7260 -2310 7320 -2270
rect 7260 -2340 7275 -2310
rect 7305 -2340 7320 -2310
rect 7260 -2380 7320 -2340
rect 7260 -2410 7275 -2380
rect 7305 -2410 7320 -2380
rect 7260 -2445 7320 -2410
rect 7260 -2475 7275 -2445
rect 7305 -2475 7320 -2445
rect 7260 -2505 7320 -2475
rect 7260 -2535 7275 -2505
rect 7305 -2535 7320 -2505
rect 7260 -2570 7320 -2535
rect 7260 -2600 7275 -2570
rect 7305 -2600 7320 -2570
rect 7260 -2640 7320 -2600
rect 7260 -2670 7275 -2640
rect 7305 -2670 7320 -2640
rect 7260 -2710 7320 -2670
rect 7260 -2740 7275 -2710
rect 7305 -2740 7320 -2710
rect 7260 -2780 7320 -2740
rect 7260 -2810 7275 -2780
rect 7305 -2810 7320 -2780
rect 7260 -2845 7320 -2810
rect 7260 -2875 7275 -2845
rect 7305 -2875 7320 -2845
rect 7260 -2905 7320 -2875
rect 7260 -2935 7275 -2905
rect 7305 -2935 7320 -2905
rect 7260 -2970 7320 -2935
rect 7260 -3000 7275 -2970
rect 7305 -3000 7320 -2970
rect 7260 -3040 7320 -3000
rect 7260 -3070 7275 -3040
rect 7305 -3070 7320 -3040
rect 7260 -3110 7320 -3070
rect 7260 -3140 7275 -3110
rect 7305 -3140 7320 -3110
rect 7260 -3180 7320 -3140
rect 7260 -3210 7275 -3180
rect 7305 -3210 7320 -3180
rect 7260 -3245 7320 -3210
rect 7260 -3275 7275 -3245
rect 7305 -3275 7320 -3245
rect 7260 -3305 7320 -3275
rect 7260 -3335 7275 -3305
rect 7305 -3335 7320 -3305
rect 7260 -3370 7320 -3335
rect 7260 -3400 7275 -3370
rect 7305 -3400 7320 -3370
rect 7260 -3440 7320 -3400
rect 7260 -3470 7275 -3440
rect 7305 -3470 7320 -3440
rect 7260 -3510 7320 -3470
rect 7260 -3540 7275 -3510
rect 7305 -3540 7320 -3510
rect 7260 -3580 7320 -3540
rect 7260 -3610 7275 -3580
rect 7305 -3610 7320 -3580
rect 7260 -3645 7320 -3610
rect 7260 -3675 7275 -3645
rect 7305 -3675 7320 -3645
rect 7260 -3705 7320 -3675
rect 7260 -3735 7275 -3705
rect 7305 -3735 7320 -3705
rect 7260 -3770 7320 -3735
rect 7260 -3800 7275 -3770
rect 7305 -3800 7320 -3770
rect 7260 -3840 7320 -3800
rect 7260 -3870 7275 -3840
rect 7305 -3870 7320 -3840
rect 7260 -3910 7320 -3870
rect 7260 -3940 7275 -3910
rect 7305 -3940 7320 -3910
rect 7260 -3980 7320 -3940
rect 7260 -4010 7275 -3980
rect 7305 -4010 7320 -3980
rect 7260 -4045 7320 -4010
rect 7260 -4075 7275 -4045
rect 7305 -4075 7320 -4045
rect 7260 -4105 7320 -4075
rect 7260 -4135 7275 -4105
rect 7305 -4135 7320 -4105
rect 7260 -4170 7320 -4135
rect 7260 -4200 7275 -4170
rect 7305 -4200 7320 -4170
rect 7260 -4240 7320 -4200
rect 7260 -4270 7275 -4240
rect 7305 -4270 7320 -4240
rect 7260 -4310 7320 -4270
rect 7260 -4340 7275 -4310
rect 7305 -4340 7320 -4310
rect 7260 -4380 7320 -4340
rect 7260 -4410 7275 -4380
rect 7305 -4410 7320 -4380
rect 7260 -4445 7320 -4410
rect 7260 -4475 7275 -4445
rect 7305 -4475 7320 -4445
rect 7260 -4490 7320 -4475
rect 7610 -1305 7670 -1290
rect 7610 -1335 7625 -1305
rect 7655 -1335 7670 -1305
rect 7610 -1370 7670 -1335
rect 7610 -1400 7625 -1370
rect 7655 -1400 7670 -1370
rect 7610 -1440 7670 -1400
rect 7610 -1470 7625 -1440
rect 7655 -1470 7670 -1440
rect 7610 -1510 7670 -1470
rect 7610 -1540 7625 -1510
rect 7655 -1540 7670 -1510
rect 7610 -1580 7670 -1540
rect 7610 -1610 7625 -1580
rect 7655 -1610 7670 -1580
rect 7610 -1645 7670 -1610
rect 7610 -1675 7625 -1645
rect 7655 -1675 7670 -1645
rect 7610 -1705 7670 -1675
rect 7610 -1735 7625 -1705
rect 7655 -1735 7670 -1705
rect 7610 -1770 7670 -1735
rect 7610 -1800 7625 -1770
rect 7655 -1800 7670 -1770
rect 7610 -1840 7670 -1800
rect 7610 -1870 7625 -1840
rect 7655 -1870 7670 -1840
rect 7610 -1910 7670 -1870
rect 7610 -1940 7625 -1910
rect 7655 -1940 7670 -1910
rect 7610 -1980 7670 -1940
rect 7610 -2010 7625 -1980
rect 7655 -2010 7670 -1980
rect 7610 -2045 7670 -2010
rect 7610 -2075 7625 -2045
rect 7655 -2075 7670 -2045
rect 7610 -2105 7670 -2075
rect 7610 -2135 7625 -2105
rect 7655 -2135 7670 -2105
rect 7610 -2170 7670 -2135
rect 7610 -2200 7625 -2170
rect 7655 -2200 7670 -2170
rect 7610 -2240 7670 -2200
rect 7610 -2270 7625 -2240
rect 7655 -2270 7670 -2240
rect 7610 -2310 7670 -2270
rect 7610 -2340 7625 -2310
rect 7655 -2340 7670 -2310
rect 7610 -2380 7670 -2340
rect 7610 -2410 7625 -2380
rect 7655 -2410 7670 -2380
rect 7610 -2445 7670 -2410
rect 7610 -2475 7625 -2445
rect 7655 -2475 7670 -2445
rect 7610 -2505 7670 -2475
rect 7610 -2535 7625 -2505
rect 7655 -2535 7670 -2505
rect 7610 -2570 7670 -2535
rect 7610 -2600 7625 -2570
rect 7655 -2600 7670 -2570
rect 7610 -2640 7670 -2600
rect 7610 -2670 7625 -2640
rect 7655 -2670 7670 -2640
rect 7610 -2710 7670 -2670
rect 7610 -2740 7625 -2710
rect 7655 -2740 7670 -2710
rect 7610 -2780 7670 -2740
rect 7610 -2810 7625 -2780
rect 7655 -2810 7670 -2780
rect 7610 -2845 7670 -2810
rect 7610 -2875 7625 -2845
rect 7655 -2875 7670 -2845
rect 7610 -2905 7670 -2875
rect 7610 -2935 7625 -2905
rect 7655 -2935 7670 -2905
rect 7610 -2970 7670 -2935
rect 7610 -3000 7625 -2970
rect 7655 -3000 7670 -2970
rect 7610 -3040 7670 -3000
rect 7610 -3070 7625 -3040
rect 7655 -3070 7670 -3040
rect 7610 -3110 7670 -3070
rect 7610 -3140 7625 -3110
rect 7655 -3140 7670 -3110
rect 7610 -3180 7670 -3140
rect 7610 -3210 7625 -3180
rect 7655 -3210 7670 -3180
rect 7610 -3245 7670 -3210
rect 7610 -3275 7625 -3245
rect 7655 -3275 7670 -3245
rect 7610 -3305 7670 -3275
rect 7610 -3335 7625 -3305
rect 7655 -3335 7670 -3305
rect 7610 -3370 7670 -3335
rect 7610 -3400 7625 -3370
rect 7655 -3400 7670 -3370
rect 7610 -3440 7670 -3400
rect 7610 -3470 7625 -3440
rect 7655 -3470 7670 -3440
rect 7610 -3510 7670 -3470
rect 7610 -3540 7625 -3510
rect 7655 -3540 7670 -3510
rect 7610 -3580 7670 -3540
rect 7610 -3610 7625 -3580
rect 7655 -3610 7670 -3580
rect 7610 -3645 7670 -3610
rect 7610 -3675 7625 -3645
rect 7655 -3675 7670 -3645
rect 7610 -3705 7670 -3675
rect 7610 -3735 7625 -3705
rect 7655 -3735 7670 -3705
rect 7610 -3770 7670 -3735
rect 7610 -3800 7625 -3770
rect 7655 -3800 7670 -3770
rect 7610 -3840 7670 -3800
rect 7610 -3870 7625 -3840
rect 7655 -3870 7670 -3840
rect 7610 -3910 7670 -3870
rect 7610 -3940 7625 -3910
rect 7655 -3940 7670 -3910
rect 7610 -3980 7670 -3940
rect 7610 -4010 7625 -3980
rect 7655 -4010 7670 -3980
rect 7610 -4045 7670 -4010
rect 7610 -4075 7625 -4045
rect 7655 -4075 7670 -4045
rect 7610 -4105 7670 -4075
rect 7610 -4135 7625 -4105
rect 7655 -4135 7670 -4105
rect 7610 -4170 7670 -4135
rect 7610 -4200 7625 -4170
rect 7655 -4200 7670 -4170
rect 7610 -4240 7670 -4200
rect 7610 -4270 7625 -4240
rect 7655 -4270 7670 -4240
rect 7610 -4310 7670 -4270
rect 7610 -4340 7625 -4310
rect 7655 -4340 7670 -4310
rect 7610 -4380 7670 -4340
rect 7610 -4410 7625 -4380
rect 7655 -4410 7670 -4380
rect 7610 -4445 7670 -4410
rect 7610 -4475 7625 -4445
rect 7655 -4475 7670 -4445
rect 7610 -4490 7670 -4475
rect 7960 -1305 8020 -1290
rect 7960 -1335 7975 -1305
rect 8005 -1335 8020 -1305
rect 7960 -1370 8020 -1335
rect 7960 -1400 7975 -1370
rect 8005 -1400 8020 -1370
rect 7960 -1440 8020 -1400
rect 7960 -1470 7975 -1440
rect 8005 -1470 8020 -1440
rect 7960 -1510 8020 -1470
rect 7960 -1540 7975 -1510
rect 8005 -1540 8020 -1510
rect 7960 -1580 8020 -1540
rect 7960 -1610 7975 -1580
rect 8005 -1610 8020 -1580
rect 7960 -1645 8020 -1610
rect 7960 -1675 7975 -1645
rect 8005 -1675 8020 -1645
rect 7960 -1705 8020 -1675
rect 7960 -1735 7975 -1705
rect 8005 -1735 8020 -1705
rect 7960 -1770 8020 -1735
rect 7960 -1800 7975 -1770
rect 8005 -1800 8020 -1770
rect 7960 -1840 8020 -1800
rect 7960 -1870 7975 -1840
rect 8005 -1870 8020 -1840
rect 7960 -1910 8020 -1870
rect 7960 -1940 7975 -1910
rect 8005 -1940 8020 -1910
rect 7960 -1980 8020 -1940
rect 7960 -2010 7975 -1980
rect 8005 -2010 8020 -1980
rect 7960 -2045 8020 -2010
rect 7960 -2075 7975 -2045
rect 8005 -2075 8020 -2045
rect 7960 -2105 8020 -2075
rect 7960 -2135 7975 -2105
rect 8005 -2135 8020 -2105
rect 7960 -2170 8020 -2135
rect 7960 -2200 7975 -2170
rect 8005 -2200 8020 -2170
rect 7960 -2240 8020 -2200
rect 7960 -2270 7975 -2240
rect 8005 -2270 8020 -2240
rect 7960 -2310 8020 -2270
rect 7960 -2340 7975 -2310
rect 8005 -2340 8020 -2310
rect 7960 -2380 8020 -2340
rect 7960 -2410 7975 -2380
rect 8005 -2410 8020 -2380
rect 7960 -2445 8020 -2410
rect 7960 -2475 7975 -2445
rect 8005 -2475 8020 -2445
rect 7960 -2505 8020 -2475
rect 7960 -2535 7975 -2505
rect 8005 -2535 8020 -2505
rect 7960 -2570 8020 -2535
rect 7960 -2600 7975 -2570
rect 8005 -2600 8020 -2570
rect 7960 -2640 8020 -2600
rect 7960 -2670 7975 -2640
rect 8005 -2670 8020 -2640
rect 7960 -2710 8020 -2670
rect 7960 -2740 7975 -2710
rect 8005 -2740 8020 -2710
rect 7960 -2780 8020 -2740
rect 7960 -2810 7975 -2780
rect 8005 -2810 8020 -2780
rect 7960 -2845 8020 -2810
rect 7960 -2875 7975 -2845
rect 8005 -2875 8020 -2845
rect 7960 -2905 8020 -2875
rect 7960 -2935 7975 -2905
rect 8005 -2935 8020 -2905
rect 7960 -2970 8020 -2935
rect 7960 -3000 7975 -2970
rect 8005 -3000 8020 -2970
rect 7960 -3040 8020 -3000
rect 7960 -3070 7975 -3040
rect 8005 -3070 8020 -3040
rect 7960 -3110 8020 -3070
rect 7960 -3140 7975 -3110
rect 8005 -3140 8020 -3110
rect 7960 -3180 8020 -3140
rect 7960 -3210 7975 -3180
rect 8005 -3210 8020 -3180
rect 7960 -3245 8020 -3210
rect 7960 -3275 7975 -3245
rect 8005 -3275 8020 -3245
rect 7960 -3305 8020 -3275
rect 7960 -3335 7975 -3305
rect 8005 -3335 8020 -3305
rect 7960 -3370 8020 -3335
rect 7960 -3400 7975 -3370
rect 8005 -3400 8020 -3370
rect 7960 -3440 8020 -3400
rect 7960 -3470 7975 -3440
rect 8005 -3470 8020 -3440
rect 7960 -3510 8020 -3470
rect 7960 -3540 7975 -3510
rect 8005 -3540 8020 -3510
rect 7960 -3580 8020 -3540
rect 7960 -3610 7975 -3580
rect 8005 -3610 8020 -3580
rect 7960 -3645 8020 -3610
rect 7960 -3675 7975 -3645
rect 8005 -3675 8020 -3645
rect 7960 -3705 8020 -3675
rect 7960 -3735 7975 -3705
rect 8005 -3735 8020 -3705
rect 7960 -3770 8020 -3735
rect 7960 -3800 7975 -3770
rect 8005 -3800 8020 -3770
rect 7960 -3840 8020 -3800
rect 7960 -3870 7975 -3840
rect 8005 -3870 8020 -3840
rect 7960 -3910 8020 -3870
rect 7960 -3940 7975 -3910
rect 8005 -3940 8020 -3910
rect 7960 -3980 8020 -3940
rect 7960 -4010 7975 -3980
rect 8005 -4010 8020 -3980
rect 7960 -4045 8020 -4010
rect 7960 -4075 7975 -4045
rect 8005 -4075 8020 -4045
rect 7960 -4105 8020 -4075
rect 7960 -4135 7975 -4105
rect 8005 -4135 8020 -4105
rect 7960 -4170 8020 -4135
rect 7960 -4200 7975 -4170
rect 8005 -4200 8020 -4170
rect 7960 -4240 8020 -4200
rect 7960 -4270 7975 -4240
rect 8005 -4270 8020 -4240
rect 7960 -4310 8020 -4270
rect 7960 -4340 7975 -4310
rect 8005 -4340 8020 -4310
rect 7960 -4380 8020 -4340
rect 7960 -4410 7975 -4380
rect 8005 -4410 8020 -4380
rect 7960 -4445 8020 -4410
rect 7960 -4475 7975 -4445
rect 8005 -4475 8020 -4445
rect 7960 -4490 8020 -4475
rect 8310 -1305 8370 -1290
rect 8310 -1335 8325 -1305
rect 8355 -1335 8370 -1305
rect 8310 -1370 8370 -1335
rect 8310 -1400 8325 -1370
rect 8355 -1400 8370 -1370
rect 8310 -1440 8370 -1400
rect 8310 -1470 8325 -1440
rect 8355 -1470 8370 -1440
rect 8310 -1510 8370 -1470
rect 8310 -1540 8325 -1510
rect 8355 -1540 8370 -1510
rect 8310 -1580 8370 -1540
rect 8310 -1610 8325 -1580
rect 8355 -1610 8370 -1580
rect 8310 -1645 8370 -1610
rect 8310 -1675 8325 -1645
rect 8355 -1675 8370 -1645
rect 8310 -1705 8370 -1675
rect 8310 -1735 8325 -1705
rect 8355 -1735 8370 -1705
rect 8310 -1770 8370 -1735
rect 8310 -1800 8325 -1770
rect 8355 -1800 8370 -1770
rect 8310 -1840 8370 -1800
rect 8310 -1870 8325 -1840
rect 8355 -1870 8370 -1840
rect 8310 -1910 8370 -1870
rect 8310 -1940 8325 -1910
rect 8355 -1940 8370 -1910
rect 8310 -1980 8370 -1940
rect 8310 -2010 8325 -1980
rect 8355 -2010 8370 -1980
rect 8310 -2045 8370 -2010
rect 8310 -2075 8325 -2045
rect 8355 -2075 8370 -2045
rect 8310 -2105 8370 -2075
rect 8310 -2135 8325 -2105
rect 8355 -2135 8370 -2105
rect 8310 -2170 8370 -2135
rect 8310 -2200 8325 -2170
rect 8355 -2200 8370 -2170
rect 8310 -2240 8370 -2200
rect 8310 -2270 8325 -2240
rect 8355 -2270 8370 -2240
rect 8310 -2310 8370 -2270
rect 8310 -2340 8325 -2310
rect 8355 -2340 8370 -2310
rect 8310 -2380 8370 -2340
rect 8310 -2410 8325 -2380
rect 8355 -2410 8370 -2380
rect 8310 -2445 8370 -2410
rect 8310 -2475 8325 -2445
rect 8355 -2475 8370 -2445
rect 8310 -2505 8370 -2475
rect 8310 -2535 8325 -2505
rect 8355 -2535 8370 -2505
rect 8310 -2570 8370 -2535
rect 8310 -2600 8325 -2570
rect 8355 -2600 8370 -2570
rect 8310 -2640 8370 -2600
rect 8310 -2670 8325 -2640
rect 8355 -2670 8370 -2640
rect 8310 -2710 8370 -2670
rect 8310 -2740 8325 -2710
rect 8355 -2740 8370 -2710
rect 8310 -2780 8370 -2740
rect 8310 -2810 8325 -2780
rect 8355 -2810 8370 -2780
rect 8310 -2845 8370 -2810
rect 8310 -2875 8325 -2845
rect 8355 -2875 8370 -2845
rect 8310 -2905 8370 -2875
rect 8310 -2935 8325 -2905
rect 8355 -2935 8370 -2905
rect 8310 -2970 8370 -2935
rect 8310 -3000 8325 -2970
rect 8355 -3000 8370 -2970
rect 8310 -3040 8370 -3000
rect 8310 -3070 8325 -3040
rect 8355 -3070 8370 -3040
rect 8310 -3110 8370 -3070
rect 8310 -3140 8325 -3110
rect 8355 -3140 8370 -3110
rect 8310 -3180 8370 -3140
rect 8310 -3210 8325 -3180
rect 8355 -3210 8370 -3180
rect 8310 -3245 8370 -3210
rect 8310 -3275 8325 -3245
rect 8355 -3275 8370 -3245
rect 8310 -3305 8370 -3275
rect 8310 -3335 8325 -3305
rect 8355 -3335 8370 -3305
rect 8310 -3370 8370 -3335
rect 8310 -3400 8325 -3370
rect 8355 -3400 8370 -3370
rect 8310 -3440 8370 -3400
rect 8310 -3470 8325 -3440
rect 8355 -3470 8370 -3440
rect 8310 -3510 8370 -3470
rect 8310 -3540 8325 -3510
rect 8355 -3540 8370 -3510
rect 8310 -3580 8370 -3540
rect 8310 -3610 8325 -3580
rect 8355 -3610 8370 -3580
rect 8310 -3645 8370 -3610
rect 8310 -3675 8325 -3645
rect 8355 -3675 8370 -3645
rect 8310 -3705 8370 -3675
rect 8310 -3735 8325 -3705
rect 8355 -3735 8370 -3705
rect 8310 -3770 8370 -3735
rect 8310 -3800 8325 -3770
rect 8355 -3800 8370 -3770
rect 8310 -3840 8370 -3800
rect 8310 -3870 8325 -3840
rect 8355 -3870 8370 -3840
rect 8310 -3910 8370 -3870
rect 8310 -3940 8325 -3910
rect 8355 -3940 8370 -3910
rect 8310 -3980 8370 -3940
rect 8310 -4010 8325 -3980
rect 8355 -4010 8370 -3980
rect 8310 -4045 8370 -4010
rect 8310 -4075 8325 -4045
rect 8355 -4075 8370 -4045
rect 8310 -4105 8370 -4075
rect 8310 -4135 8325 -4105
rect 8355 -4135 8370 -4105
rect 8310 -4170 8370 -4135
rect 8310 -4200 8325 -4170
rect 8355 -4200 8370 -4170
rect 8310 -4240 8370 -4200
rect 8310 -4270 8325 -4240
rect 8355 -4270 8370 -4240
rect 8310 -4310 8370 -4270
rect 8310 -4340 8325 -4310
rect 8355 -4340 8370 -4310
rect 8310 -4380 8370 -4340
rect 8310 -4410 8325 -4380
rect 8355 -4410 8370 -4380
rect 8310 -4445 8370 -4410
rect 8310 -4475 8325 -4445
rect 8355 -4475 8370 -4445
rect 8310 -4490 8370 -4475
rect 8660 -1305 8720 -1290
rect 8660 -1335 8675 -1305
rect 8705 -1335 8720 -1305
rect 8660 -1370 8720 -1335
rect 8660 -1400 8675 -1370
rect 8705 -1400 8720 -1370
rect 8660 -1440 8720 -1400
rect 8660 -1470 8675 -1440
rect 8705 -1470 8720 -1440
rect 8660 -1510 8720 -1470
rect 8660 -1540 8675 -1510
rect 8705 -1540 8720 -1510
rect 8660 -1580 8720 -1540
rect 8660 -1610 8675 -1580
rect 8705 -1610 8720 -1580
rect 8660 -1645 8720 -1610
rect 8660 -1675 8675 -1645
rect 8705 -1675 8720 -1645
rect 8660 -1705 8720 -1675
rect 8660 -1735 8675 -1705
rect 8705 -1735 8720 -1705
rect 8660 -1770 8720 -1735
rect 8660 -1800 8675 -1770
rect 8705 -1800 8720 -1770
rect 8660 -1840 8720 -1800
rect 8660 -1870 8675 -1840
rect 8705 -1870 8720 -1840
rect 8660 -1910 8720 -1870
rect 8660 -1940 8675 -1910
rect 8705 -1940 8720 -1910
rect 8660 -1980 8720 -1940
rect 8660 -2010 8675 -1980
rect 8705 -2010 8720 -1980
rect 8660 -2045 8720 -2010
rect 8660 -2075 8675 -2045
rect 8705 -2075 8720 -2045
rect 8660 -2105 8720 -2075
rect 8660 -2135 8675 -2105
rect 8705 -2135 8720 -2105
rect 8660 -2170 8720 -2135
rect 8660 -2200 8675 -2170
rect 8705 -2200 8720 -2170
rect 8660 -2240 8720 -2200
rect 8660 -2270 8675 -2240
rect 8705 -2270 8720 -2240
rect 8660 -2310 8720 -2270
rect 8660 -2340 8675 -2310
rect 8705 -2340 8720 -2310
rect 8660 -2380 8720 -2340
rect 8660 -2410 8675 -2380
rect 8705 -2410 8720 -2380
rect 8660 -2445 8720 -2410
rect 8660 -2475 8675 -2445
rect 8705 -2475 8720 -2445
rect 8660 -2505 8720 -2475
rect 8660 -2535 8675 -2505
rect 8705 -2535 8720 -2505
rect 8660 -2570 8720 -2535
rect 8660 -2600 8675 -2570
rect 8705 -2600 8720 -2570
rect 8660 -2640 8720 -2600
rect 8660 -2670 8675 -2640
rect 8705 -2670 8720 -2640
rect 8660 -2710 8720 -2670
rect 8660 -2740 8675 -2710
rect 8705 -2740 8720 -2710
rect 8660 -2780 8720 -2740
rect 8660 -2810 8675 -2780
rect 8705 -2810 8720 -2780
rect 8660 -2845 8720 -2810
rect 8660 -2875 8675 -2845
rect 8705 -2875 8720 -2845
rect 8660 -2905 8720 -2875
rect 8660 -2935 8675 -2905
rect 8705 -2935 8720 -2905
rect 8660 -2970 8720 -2935
rect 8660 -3000 8675 -2970
rect 8705 -3000 8720 -2970
rect 8660 -3040 8720 -3000
rect 8660 -3070 8675 -3040
rect 8705 -3070 8720 -3040
rect 8660 -3110 8720 -3070
rect 8660 -3140 8675 -3110
rect 8705 -3140 8720 -3110
rect 8660 -3180 8720 -3140
rect 8660 -3210 8675 -3180
rect 8705 -3210 8720 -3180
rect 8660 -3245 8720 -3210
rect 8660 -3275 8675 -3245
rect 8705 -3275 8720 -3245
rect 8660 -3305 8720 -3275
rect 8660 -3335 8675 -3305
rect 8705 -3335 8720 -3305
rect 8660 -3370 8720 -3335
rect 8660 -3400 8675 -3370
rect 8705 -3400 8720 -3370
rect 8660 -3440 8720 -3400
rect 8660 -3470 8675 -3440
rect 8705 -3470 8720 -3440
rect 8660 -3510 8720 -3470
rect 8660 -3540 8675 -3510
rect 8705 -3540 8720 -3510
rect 8660 -3580 8720 -3540
rect 8660 -3610 8675 -3580
rect 8705 -3610 8720 -3580
rect 8660 -3645 8720 -3610
rect 8660 -3675 8675 -3645
rect 8705 -3675 8720 -3645
rect 8660 -3705 8720 -3675
rect 8660 -3735 8675 -3705
rect 8705 -3735 8720 -3705
rect 8660 -3770 8720 -3735
rect 8660 -3800 8675 -3770
rect 8705 -3800 8720 -3770
rect 8660 -3840 8720 -3800
rect 8660 -3870 8675 -3840
rect 8705 -3870 8720 -3840
rect 8660 -3910 8720 -3870
rect 8660 -3940 8675 -3910
rect 8705 -3940 8720 -3910
rect 8660 -3980 8720 -3940
rect 8660 -4010 8675 -3980
rect 8705 -4010 8720 -3980
rect 8660 -4045 8720 -4010
rect 8660 -4075 8675 -4045
rect 8705 -4075 8720 -4045
rect 8660 -4105 8720 -4075
rect 8660 -4135 8675 -4105
rect 8705 -4135 8720 -4105
rect 8660 -4170 8720 -4135
rect 8660 -4200 8675 -4170
rect 8705 -4200 8720 -4170
rect 8660 -4240 8720 -4200
rect 8660 -4270 8675 -4240
rect 8705 -4270 8720 -4240
rect 8660 -4310 8720 -4270
rect 8660 -4340 8675 -4310
rect 8705 -4340 8720 -4310
rect 8660 -4380 8720 -4340
rect 8660 -4410 8675 -4380
rect 8705 -4410 8720 -4380
rect 8660 -4445 8720 -4410
rect 8660 -4475 8675 -4445
rect 8705 -4475 8720 -4445
rect 8660 -4490 8720 -4475
rect 9010 -1305 9070 -1290
rect 9010 -1335 9025 -1305
rect 9055 -1335 9070 -1305
rect 9010 -1370 9070 -1335
rect 9010 -1400 9025 -1370
rect 9055 -1400 9070 -1370
rect 9010 -1440 9070 -1400
rect 9010 -1470 9025 -1440
rect 9055 -1470 9070 -1440
rect 9010 -1510 9070 -1470
rect 9010 -1540 9025 -1510
rect 9055 -1540 9070 -1510
rect 9010 -1580 9070 -1540
rect 9010 -1610 9025 -1580
rect 9055 -1610 9070 -1580
rect 9010 -1645 9070 -1610
rect 9010 -1675 9025 -1645
rect 9055 -1675 9070 -1645
rect 9010 -1705 9070 -1675
rect 9010 -1735 9025 -1705
rect 9055 -1735 9070 -1705
rect 9010 -1770 9070 -1735
rect 9010 -1800 9025 -1770
rect 9055 -1800 9070 -1770
rect 9010 -1840 9070 -1800
rect 9010 -1870 9025 -1840
rect 9055 -1870 9070 -1840
rect 9010 -1910 9070 -1870
rect 9010 -1940 9025 -1910
rect 9055 -1940 9070 -1910
rect 9010 -1980 9070 -1940
rect 9010 -2010 9025 -1980
rect 9055 -2010 9070 -1980
rect 9010 -2045 9070 -2010
rect 9010 -2075 9025 -2045
rect 9055 -2075 9070 -2045
rect 9010 -2105 9070 -2075
rect 9010 -2135 9025 -2105
rect 9055 -2135 9070 -2105
rect 9010 -2170 9070 -2135
rect 9010 -2200 9025 -2170
rect 9055 -2200 9070 -2170
rect 9010 -2240 9070 -2200
rect 9010 -2270 9025 -2240
rect 9055 -2270 9070 -2240
rect 9010 -2310 9070 -2270
rect 9010 -2340 9025 -2310
rect 9055 -2340 9070 -2310
rect 9010 -2380 9070 -2340
rect 9010 -2410 9025 -2380
rect 9055 -2410 9070 -2380
rect 9010 -2445 9070 -2410
rect 9010 -2475 9025 -2445
rect 9055 -2475 9070 -2445
rect 9010 -2505 9070 -2475
rect 9010 -2535 9025 -2505
rect 9055 -2535 9070 -2505
rect 9010 -2570 9070 -2535
rect 9010 -2600 9025 -2570
rect 9055 -2600 9070 -2570
rect 9010 -2640 9070 -2600
rect 9010 -2670 9025 -2640
rect 9055 -2670 9070 -2640
rect 9010 -2710 9070 -2670
rect 9010 -2740 9025 -2710
rect 9055 -2740 9070 -2710
rect 9010 -2780 9070 -2740
rect 9010 -2810 9025 -2780
rect 9055 -2810 9070 -2780
rect 9010 -2845 9070 -2810
rect 9010 -2875 9025 -2845
rect 9055 -2875 9070 -2845
rect 9010 -2905 9070 -2875
rect 9010 -2935 9025 -2905
rect 9055 -2935 9070 -2905
rect 9010 -2970 9070 -2935
rect 9010 -3000 9025 -2970
rect 9055 -3000 9070 -2970
rect 9010 -3040 9070 -3000
rect 9010 -3070 9025 -3040
rect 9055 -3070 9070 -3040
rect 9010 -3110 9070 -3070
rect 9010 -3140 9025 -3110
rect 9055 -3140 9070 -3110
rect 9010 -3180 9070 -3140
rect 9010 -3210 9025 -3180
rect 9055 -3210 9070 -3180
rect 9010 -3245 9070 -3210
rect 9010 -3275 9025 -3245
rect 9055 -3275 9070 -3245
rect 9010 -3305 9070 -3275
rect 9010 -3335 9025 -3305
rect 9055 -3335 9070 -3305
rect 9010 -3370 9070 -3335
rect 9010 -3400 9025 -3370
rect 9055 -3400 9070 -3370
rect 9010 -3440 9070 -3400
rect 9010 -3470 9025 -3440
rect 9055 -3470 9070 -3440
rect 9010 -3510 9070 -3470
rect 9010 -3540 9025 -3510
rect 9055 -3540 9070 -3510
rect 9010 -3580 9070 -3540
rect 9010 -3610 9025 -3580
rect 9055 -3610 9070 -3580
rect 9010 -3645 9070 -3610
rect 9010 -3675 9025 -3645
rect 9055 -3675 9070 -3645
rect 9010 -3705 9070 -3675
rect 9010 -3735 9025 -3705
rect 9055 -3735 9070 -3705
rect 9010 -3770 9070 -3735
rect 9010 -3800 9025 -3770
rect 9055 -3800 9070 -3770
rect 9010 -3840 9070 -3800
rect 9010 -3870 9025 -3840
rect 9055 -3870 9070 -3840
rect 9010 -3910 9070 -3870
rect 9010 -3940 9025 -3910
rect 9055 -3940 9070 -3910
rect 9010 -3980 9070 -3940
rect 9010 -4010 9025 -3980
rect 9055 -4010 9070 -3980
rect 9010 -4045 9070 -4010
rect 9010 -4075 9025 -4045
rect 9055 -4075 9070 -4045
rect 9010 -4105 9070 -4075
rect 9010 -4135 9025 -4105
rect 9055 -4135 9070 -4105
rect 9010 -4170 9070 -4135
rect 9010 -4200 9025 -4170
rect 9055 -4200 9070 -4170
rect 9010 -4240 9070 -4200
rect 9010 -4270 9025 -4240
rect 9055 -4270 9070 -4240
rect 9010 -4310 9070 -4270
rect 9010 -4340 9025 -4310
rect 9055 -4340 9070 -4310
rect 9010 -4380 9070 -4340
rect 9010 -4410 9025 -4380
rect 9055 -4410 9070 -4380
rect 9010 -4445 9070 -4410
rect 9010 -4475 9025 -4445
rect 9055 -4475 9070 -4445
rect 9010 -4490 9070 -4475
<< via2 >>
rect 2195 20880 2225 20910
rect 2195 20815 2225 20845
rect 2195 20745 2225 20775
rect 2195 20675 2225 20705
rect 2195 20605 2225 20635
rect 2195 20540 2225 20570
rect 2195 20480 2225 20510
rect 2195 20415 2225 20445
rect 2195 20345 2225 20375
rect 2195 20275 2225 20305
rect 2195 20205 2225 20235
rect 2195 20140 2225 20170
rect 2195 20080 2225 20110
rect 2195 20015 2225 20045
rect 2195 19945 2225 19975
rect 2195 19875 2225 19905
rect 2195 19805 2225 19835
rect 2195 19740 2225 19770
rect 2195 19680 2225 19710
rect 2195 19615 2225 19645
rect 2195 19545 2225 19575
rect 2195 19475 2225 19505
rect 2195 19405 2225 19435
rect 2195 19340 2225 19370
rect 2195 19280 2225 19310
rect 2195 19215 2225 19245
rect 2195 19145 2225 19175
rect 2195 19075 2225 19105
rect 2195 19005 2225 19035
rect 2195 18940 2225 18970
rect 2195 18880 2225 18910
rect 2195 18815 2225 18845
rect 2195 18745 2225 18775
rect 2195 18675 2225 18705
rect 2195 18605 2225 18635
rect 2195 18540 2225 18570
rect 2195 18480 2225 18510
rect 2195 18415 2225 18445
rect 2195 18345 2225 18375
rect 2195 18275 2225 18305
rect 2195 18205 2225 18235
rect 2195 18140 2225 18170
rect 2195 18080 2225 18110
rect 2195 18015 2225 18045
rect 2195 17945 2225 17975
rect 2195 17875 2225 17905
rect 2195 17805 2225 17835
rect 2195 17740 2225 17770
rect 6665 20880 6695 20910
rect 6665 20815 6695 20845
rect 6665 20745 6695 20775
rect 6665 20675 6695 20705
rect 6665 20605 6695 20635
rect 6665 20540 6695 20570
rect 6665 20480 6695 20510
rect 6665 20415 6695 20445
rect 6665 20345 6695 20375
rect 6665 20275 6695 20305
rect 6665 20205 6695 20235
rect 6665 20140 6695 20170
rect 6665 20080 6695 20110
rect 6665 20015 6695 20045
rect 6665 19945 6695 19975
rect 6665 19875 6695 19905
rect 6665 19805 6695 19835
rect 6665 19740 6695 19770
rect 6665 19680 6695 19710
rect 6665 19615 6695 19645
rect 6665 19545 6695 19575
rect 6665 19475 6695 19505
rect 6665 19405 6695 19435
rect 6665 19340 6695 19370
rect 6665 19280 6695 19310
rect 6665 19215 6695 19245
rect 6665 19145 6695 19175
rect 6665 19075 6695 19105
rect 6665 19005 6695 19035
rect 6665 18940 6695 18970
rect 6665 18880 6695 18910
rect 6665 18815 6695 18845
rect 6665 18745 6695 18775
rect 6665 18675 6695 18705
rect 6665 18605 6695 18635
rect 6665 18540 6695 18570
rect 6665 18480 6695 18510
rect 6665 18415 6695 18445
rect 6665 18345 6695 18375
rect 6665 18275 6695 18305
rect 6665 18205 6695 18235
rect 6665 18140 6695 18170
rect 6665 18080 6695 18110
rect 6665 18015 6695 18045
rect 6665 17945 6695 17975
rect 6665 17875 6695 17905
rect 6665 17805 6695 17835
rect 6665 17740 6695 17770
rect -75 9605 -45 9635
rect -75 9540 -45 9570
rect -75 9470 -45 9500
rect -75 9400 -45 9430
rect -75 9330 -45 9360
rect -75 9265 -45 9295
rect -75 9205 -45 9235
rect -75 9140 -45 9170
rect -75 9070 -45 9100
rect -75 9000 -45 9030
rect -75 8930 -45 8960
rect -75 8865 -45 8895
rect -75 8805 -45 8835
rect -75 8740 -45 8770
rect -75 8670 -45 8700
rect -75 8600 -45 8630
rect -75 8530 -45 8560
rect -75 8465 -45 8495
rect -75 8405 -45 8435
rect -75 8340 -45 8370
rect -75 8270 -45 8300
rect -75 8200 -45 8230
rect -75 8130 -45 8160
rect -75 8065 -45 8095
rect -75 8005 -45 8035
rect -75 7940 -45 7970
rect -75 7870 -45 7900
rect -75 7800 -45 7830
rect -75 7730 -45 7760
rect -75 7665 -45 7695
rect -75 7605 -45 7635
rect -75 7540 -45 7570
rect -75 7470 -45 7500
rect -75 7400 -45 7430
rect -75 7330 -45 7360
rect -75 7265 -45 7295
rect -75 7205 -45 7235
rect -75 7140 -45 7170
rect -75 7070 -45 7100
rect -75 7000 -45 7030
rect -75 6930 -45 6960
rect -75 6865 -45 6895
rect -75 6805 -45 6835
rect -75 6740 -45 6770
rect -75 6670 -45 6700
rect -75 6600 -45 6630
rect -75 6530 -45 6560
rect -75 6465 -45 6495
rect 275 9605 305 9635
rect 275 9540 305 9570
rect 275 9470 305 9500
rect 275 9400 305 9430
rect 275 9330 305 9360
rect 275 9265 305 9295
rect 275 9205 305 9235
rect 275 9140 305 9170
rect 275 9070 305 9100
rect 275 9000 305 9030
rect 275 8930 305 8960
rect 275 8865 305 8895
rect 275 8805 305 8835
rect 275 8740 305 8770
rect 275 8670 305 8700
rect 275 8600 305 8630
rect 275 8530 305 8560
rect 275 8465 305 8495
rect 275 8405 305 8435
rect 275 8340 305 8370
rect 275 8270 305 8300
rect 275 8200 305 8230
rect 275 8130 305 8160
rect 275 8065 305 8095
rect 275 8005 305 8035
rect 275 7940 305 7970
rect 275 7870 305 7900
rect 275 7800 305 7830
rect 275 7730 305 7760
rect 275 7665 305 7695
rect 275 7605 305 7635
rect 275 7540 305 7570
rect 275 7470 305 7500
rect 275 7400 305 7430
rect 275 7330 305 7360
rect 275 7265 305 7295
rect 275 7205 305 7235
rect 275 7140 305 7170
rect 275 7070 305 7100
rect 275 7000 305 7030
rect 275 6930 305 6960
rect 275 6865 305 6895
rect 275 6805 305 6835
rect 275 6740 305 6770
rect 275 6670 305 6700
rect 275 6600 305 6630
rect 275 6530 305 6560
rect 275 6465 305 6495
rect 625 9605 655 9635
rect 625 9540 655 9570
rect 625 9470 655 9500
rect 625 9400 655 9430
rect 625 9330 655 9360
rect 625 9265 655 9295
rect 625 9205 655 9235
rect 625 9140 655 9170
rect 625 9070 655 9100
rect 625 9000 655 9030
rect 625 8930 655 8960
rect 625 8865 655 8895
rect 625 8805 655 8835
rect 625 8740 655 8770
rect 625 8670 655 8700
rect 625 8600 655 8630
rect 625 8530 655 8560
rect 625 8465 655 8495
rect 625 8405 655 8435
rect 625 8340 655 8370
rect 625 8270 655 8300
rect 625 8200 655 8230
rect 625 8130 655 8160
rect 625 8065 655 8095
rect 625 8005 655 8035
rect 625 7940 655 7970
rect 625 7870 655 7900
rect 625 7800 655 7830
rect 625 7730 655 7760
rect 625 7665 655 7695
rect 625 7605 655 7635
rect 625 7540 655 7570
rect 625 7470 655 7500
rect 625 7400 655 7430
rect 625 7330 655 7360
rect 625 7265 655 7295
rect 625 7205 655 7235
rect 625 7140 655 7170
rect 625 7070 655 7100
rect 625 7000 655 7030
rect 625 6930 655 6960
rect 625 6865 655 6895
rect 625 6805 655 6835
rect 625 6740 655 6770
rect 625 6670 655 6700
rect 625 6600 655 6630
rect 625 6530 655 6560
rect 625 6465 655 6495
rect 975 9605 1005 9635
rect 975 9540 1005 9570
rect 975 9470 1005 9500
rect 975 9400 1005 9430
rect 975 9330 1005 9360
rect 975 9265 1005 9295
rect 975 9205 1005 9235
rect 975 9140 1005 9170
rect 975 9070 1005 9100
rect 975 9000 1005 9030
rect 975 8930 1005 8960
rect 975 8865 1005 8895
rect 975 8805 1005 8835
rect 975 8740 1005 8770
rect 975 8670 1005 8700
rect 975 8600 1005 8630
rect 975 8530 1005 8560
rect 975 8465 1005 8495
rect 975 8405 1005 8435
rect 975 8340 1005 8370
rect 975 8270 1005 8300
rect 975 8200 1005 8230
rect 975 8130 1005 8160
rect 975 8065 1005 8095
rect 975 8005 1005 8035
rect 975 7940 1005 7970
rect 975 7870 1005 7900
rect 975 7800 1005 7830
rect 975 7730 1005 7760
rect 975 7665 1005 7695
rect 975 7605 1005 7635
rect 975 7540 1005 7570
rect 975 7470 1005 7500
rect 975 7400 1005 7430
rect 975 7330 1005 7360
rect 975 7265 1005 7295
rect 975 7205 1005 7235
rect 975 7140 1005 7170
rect 975 7070 1005 7100
rect 975 7000 1005 7030
rect 975 6930 1005 6960
rect 975 6865 1005 6895
rect 975 6805 1005 6835
rect 975 6740 1005 6770
rect 975 6670 1005 6700
rect 975 6600 1005 6630
rect 975 6530 1005 6560
rect 975 6465 1005 6495
rect 1675 9605 1705 9635
rect 1675 9540 1705 9570
rect 1675 9470 1705 9500
rect 1675 9400 1705 9430
rect 1675 9330 1705 9360
rect 1675 9265 1705 9295
rect 1675 9205 1705 9235
rect 1675 9140 1705 9170
rect 1675 9070 1705 9100
rect 1675 9000 1705 9030
rect 1675 8930 1705 8960
rect 1675 8865 1705 8895
rect 1675 8805 1705 8835
rect 1675 8740 1705 8770
rect 1675 8670 1705 8700
rect 1675 8600 1705 8630
rect 1675 8530 1705 8560
rect 1675 8465 1705 8495
rect 1675 8405 1705 8435
rect 1675 8340 1705 8370
rect 1675 8270 1705 8300
rect 1675 8200 1705 8230
rect 1675 8130 1705 8160
rect 1675 8065 1705 8095
rect 1675 8005 1705 8035
rect 1675 7940 1705 7970
rect 1675 7870 1705 7900
rect 1675 7800 1705 7830
rect 1675 7730 1705 7760
rect 1675 7665 1705 7695
rect 1675 7605 1705 7635
rect 1675 7540 1705 7570
rect 1675 7470 1705 7500
rect 1675 7400 1705 7430
rect 1675 7330 1705 7360
rect 1675 7265 1705 7295
rect 1675 7205 1705 7235
rect 1675 7140 1705 7170
rect 1675 7070 1705 7100
rect 1675 7000 1705 7030
rect 1675 6930 1705 6960
rect 1675 6865 1705 6895
rect 1675 6805 1705 6835
rect 1675 6740 1705 6770
rect 1675 6670 1705 6700
rect 1675 6600 1705 6630
rect 1675 6530 1705 6560
rect 1675 6465 1705 6495
rect 2330 9605 2360 9635
rect 2330 9540 2360 9570
rect 2330 9470 2360 9500
rect 2330 9400 2360 9430
rect 2330 9330 2360 9360
rect 2330 9265 2360 9295
rect 2330 9205 2360 9235
rect 2330 9140 2360 9170
rect 2330 9070 2360 9100
rect 2330 9000 2360 9030
rect 2330 8930 2360 8960
rect 2330 8865 2360 8895
rect 2330 8805 2360 8835
rect 2330 8740 2360 8770
rect 2330 8670 2360 8700
rect 2330 8600 2360 8630
rect 2330 8530 2360 8560
rect 2330 8465 2360 8495
rect 2330 8405 2360 8435
rect 2330 8340 2360 8370
rect 2330 8270 2360 8300
rect 2330 8200 2360 8230
rect 2330 8130 2360 8160
rect 2330 8065 2360 8095
rect 2330 8005 2360 8035
rect 2330 7940 2360 7970
rect 2330 7870 2360 7900
rect 2330 7800 2360 7830
rect 2330 7730 2360 7760
rect 2330 7665 2360 7695
rect 2330 7605 2360 7635
rect 2330 7540 2360 7570
rect 2330 7470 2360 7500
rect 2330 7400 2360 7430
rect 2330 7330 2360 7360
rect 2330 7265 2360 7295
rect 2330 7205 2360 7235
rect 2330 7140 2360 7170
rect 2330 7070 2360 7100
rect 2330 7000 2360 7030
rect 2330 6930 2360 6960
rect 2330 6865 2360 6895
rect 2330 6805 2360 6835
rect 2330 6740 2360 6770
rect 2330 6670 2360 6700
rect 2330 6600 2360 6630
rect 2330 6530 2360 6560
rect 2330 6465 2360 6495
rect 3180 9605 3210 9635
rect 3240 9605 3270 9635
rect 3180 9540 3210 9570
rect 3240 9540 3270 9570
rect 3180 9470 3210 9500
rect 3240 9470 3270 9500
rect 3180 9400 3210 9430
rect 3240 9400 3270 9430
rect 3180 9330 3210 9360
rect 3240 9330 3270 9360
rect 3180 9265 3210 9295
rect 3240 9265 3270 9295
rect 3180 9205 3210 9235
rect 3240 9205 3270 9235
rect 3180 9140 3210 9170
rect 3240 9140 3270 9170
rect 3180 9070 3210 9100
rect 3240 9070 3270 9100
rect 3180 9000 3210 9030
rect 3240 9000 3270 9030
rect 3180 8930 3210 8960
rect 3240 8930 3270 8960
rect 3180 8865 3210 8895
rect 3240 8865 3270 8895
rect 3180 8805 3210 8835
rect 3240 8805 3270 8835
rect 3180 8740 3210 8770
rect 3240 8740 3270 8770
rect 3180 8670 3210 8700
rect 3240 8670 3270 8700
rect 3180 8600 3210 8630
rect 3240 8600 3270 8630
rect 3180 8530 3210 8560
rect 3240 8530 3270 8560
rect 3180 8465 3210 8495
rect 3240 8465 3270 8495
rect 3180 8405 3210 8435
rect 3240 8405 3270 8435
rect 3180 8340 3210 8370
rect 3240 8340 3270 8370
rect 3180 8270 3210 8300
rect 3240 8270 3270 8300
rect 3180 8200 3210 8230
rect 3240 8200 3270 8230
rect 3180 8130 3210 8160
rect 3240 8130 3270 8160
rect 3180 8065 3210 8095
rect 3240 8065 3270 8095
rect 3180 8005 3210 8035
rect 3240 8005 3270 8035
rect 3180 7940 3210 7970
rect 3240 7940 3270 7970
rect 3180 7870 3210 7900
rect 3240 7870 3270 7900
rect 3180 7800 3210 7830
rect 3240 7800 3270 7830
rect 3180 7730 3210 7760
rect 3240 7730 3270 7760
rect 3180 7665 3210 7695
rect 3240 7665 3270 7695
rect 3180 7605 3210 7635
rect 3240 7605 3270 7635
rect 3180 7540 3210 7570
rect 3240 7540 3270 7570
rect 3180 7470 3210 7500
rect 3240 7470 3270 7500
rect 3180 7400 3210 7430
rect 3240 7400 3270 7430
rect 3180 7330 3210 7360
rect 3240 7330 3270 7360
rect 3180 7265 3210 7295
rect 3240 7265 3270 7295
rect 3180 7205 3210 7235
rect 3240 7205 3270 7235
rect 3180 7140 3210 7170
rect 3240 7140 3270 7170
rect 3180 7070 3210 7100
rect 3240 7070 3270 7100
rect 3180 7000 3210 7030
rect 3240 7000 3270 7030
rect 3180 6930 3210 6960
rect 3240 6930 3270 6960
rect 3180 6865 3210 6895
rect 3240 6865 3270 6895
rect 3180 6805 3210 6835
rect 3240 6805 3270 6835
rect 3180 6740 3210 6770
rect 3240 6740 3270 6770
rect 3180 6670 3210 6700
rect 3240 6670 3270 6700
rect 3180 6600 3210 6630
rect 3240 6600 3270 6630
rect 3180 6530 3210 6560
rect 3240 6530 3270 6560
rect 3180 6465 3210 6495
rect 3240 6465 3270 6495
rect 3350 9605 3380 9635
rect 3350 9540 3380 9570
rect 3350 9470 3380 9500
rect 3350 9400 3380 9430
rect 3350 9330 3380 9360
rect 3350 9265 3380 9295
rect 3350 9205 3380 9235
rect 3350 9140 3380 9170
rect 3350 9070 3380 9100
rect 3350 9000 3380 9030
rect 3350 8930 3380 8960
rect 3350 8865 3380 8895
rect 3350 8805 3380 8835
rect 3350 8740 3380 8770
rect 3350 8670 3380 8700
rect 3350 8600 3380 8630
rect 3350 8530 3380 8560
rect 3350 8465 3380 8495
rect 3350 8405 3380 8435
rect 3350 8340 3380 8370
rect 3350 8270 3380 8300
rect 3350 8200 3380 8230
rect 3350 8130 3380 8160
rect 3350 8065 3380 8095
rect 3350 8005 3380 8035
rect 3350 7940 3380 7970
rect 3350 7870 3380 7900
rect 3350 7800 3380 7830
rect 3350 7730 3380 7760
rect 3350 7665 3380 7695
rect 3350 7605 3380 7635
rect 3350 7540 3380 7570
rect 3350 7470 3380 7500
rect 3350 7400 3380 7430
rect 3350 7330 3380 7360
rect 3350 7265 3380 7295
rect 3350 7205 3380 7235
rect 3350 7140 3380 7170
rect 3350 7070 3380 7100
rect 3350 7000 3380 7030
rect 3350 6930 3380 6960
rect 3350 6865 3380 6895
rect 3350 6805 3380 6835
rect 3350 6740 3380 6770
rect 3350 6670 3380 6700
rect 3350 6600 3380 6630
rect 3350 6530 3380 6560
rect 3350 6465 3380 6495
rect 6635 9605 6665 9635
rect 6635 9540 6665 9570
rect 6635 9470 6665 9500
rect 6635 9400 6665 9430
rect 6635 9330 6665 9360
rect 6635 9265 6665 9295
rect 6635 9205 6665 9235
rect 6635 9140 6665 9170
rect 6635 9070 6665 9100
rect 6635 9000 6665 9030
rect 6635 8930 6665 8960
rect 6635 8865 6665 8895
rect 6635 8805 6665 8835
rect 6635 8740 6665 8770
rect 6635 8670 6665 8700
rect 6635 8600 6665 8630
rect 6635 8530 6665 8560
rect 6635 8465 6665 8495
rect 6635 8405 6665 8435
rect 6635 8340 6665 8370
rect 6635 8270 6665 8300
rect 6635 8200 6665 8230
rect 6635 8130 6665 8160
rect 6635 8065 6665 8095
rect 6635 8005 6665 8035
rect 6635 7940 6665 7970
rect 6635 7870 6665 7900
rect 6635 7800 6665 7830
rect 6635 7730 6665 7760
rect 6635 7665 6665 7695
rect 6635 7605 6665 7635
rect 6635 7540 6665 7570
rect 6635 7470 6665 7500
rect 6635 7400 6665 7430
rect 6635 7330 6665 7360
rect 6635 7265 6665 7295
rect 6635 7205 6665 7235
rect 6635 7140 6665 7170
rect 6635 7070 6665 7100
rect 6635 7000 6665 7030
rect 6635 6930 6665 6960
rect 6635 6865 6665 6895
rect 6635 6805 6665 6835
rect 6635 6740 6665 6770
rect 6635 6670 6665 6700
rect 6635 6600 6665 6630
rect 6635 6530 6665 6560
rect 6635 6465 6665 6495
rect 7275 9605 7305 9635
rect 7275 9540 7305 9570
rect 7275 9470 7305 9500
rect 7275 9400 7305 9430
rect 7275 9330 7305 9360
rect 7275 9265 7305 9295
rect 7275 9205 7305 9235
rect 7275 9140 7305 9170
rect 7275 9070 7305 9100
rect 7275 9000 7305 9030
rect 7275 8930 7305 8960
rect 7275 8865 7305 8895
rect 7275 8805 7305 8835
rect 7275 8740 7305 8770
rect 7275 8670 7305 8700
rect 7275 8600 7305 8630
rect 7275 8530 7305 8560
rect 7275 8465 7305 8495
rect 7275 8405 7305 8435
rect 7275 8340 7305 8370
rect 7275 8270 7305 8300
rect 7275 8200 7305 8230
rect 7275 8130 7305 8160
rect 7275 8065 7305 8095
rect 7275 8005 7305 8035
rect 7275 7940 7305 7970
rect 7275 7870 7305 7900
rect 7275 7800 7305 7830
rect 7275 7730 7305 7760
rect 7275 7665 7305 7695
rect 7275 7605 7305 7635
rect 7275 7540 7305 7570
rect 7275 7470 7305 7500
rect 7275 7400 7305 7430
rect 7275 7330 7305 7360
rect 7275 7265 7305 7295
rect 7275 7205 7305 7235
rect 7275 7140 7305 7170
rect 7275 7070 7305 7100
rect 7275 7000 7305 7030
rect 7275 6930 7305 6960
rect 7275 6865 7305 6895
rect 7275 6805 7305 6835
rect 7275 6740 7305 6770
rect 7275 6670 7305 6700
rect 7275 6600 7305 6630
rect 7275 6530 7305 6560
rect 7275 6465 7305 6495
rect 7975 9605 8005 9635
rect 7975 9540 8005 9570
rect 7975 9470 8005 9500
rect 7975 9400 8005 9430
rect 7975 9330 8005 9360
rect 7975 9265 8005 9295
rect 7975 9205 8005 9235
rect 7975 9140 8005 9170
rect 7975 9070 8005 9100
rect 7975 9000 8005 9030
rect 7975 8930 8005 8960
rect 7975 8865 8005 8895
rect 7975 8805 8005 8835
rect 7975 8740 8005 8770
rect 7975 8670 8005 8700
rect 7975 8600 8005 8630
rect 7975 8530 8005 8560
rect 7975 8465 8005 8495
rect 7975 8405 8005 8435
rect 7975 8340 8005 8370
rect 7975 8270 8005 8300
rect 7975 8200 8005 8230
rect 7975 8130 8005 8160
rect 7975 8065 8005 8095
rect 7975 8005 8005 8035
rect 7975 7940 8005 7970
rect 7975 7870 8005 7900
rect 7975 7800 8005 7830
rect 7975 7730 8005 7760
rect 7975 7665 8005 7695
rect 7975 7605 8005 7635
rect 7975 7540 8005 7570
rect 7975 7470 8005 7500
rect 7975 7400 8005 7430
rect 7975 7330 8005 7360
rect 7975 7265 8005 7295
rect 7975 7205 8005 7235
rect 7975 7140 8005 7170
rect 7975 7070 8005 7100
rect 7975 7000 8005 7030
rect 7975 6930 8005 6960
rect 7975 6865 8005 6895
rect 7975 6805 8005 6835
rect 7975 6740 8005 6770
rect 7975 6670 8005 6700
rect 7975 6600 8005 6630
rect 7975 6530 8005 6560
rect 7975 6465 8005 6495
rect 8325 9605 8355 9635
rect 8325 9540 8355 9570
rect 8325 9470 8355 9500
rect 8325 9400 8355 9430
rect 8325 9330 8355 9360
rect 8325 9265 8355 9295
rect 8325 9205 8355 9235
rect 8325 9140 8355 9170
rect 8325 9070 8355 9100
rect 8325 9000 8355 9030
rect 8325 8930 8355 8960
rect 8325 8865 8355 8895
rect 8325 8805 8355 8835
rect 8325 8740 8355 8770
rect 8325 8670 8355 8700
rect 8325 8600 8355 8630
rect 8325 8530 8355 8560
rect 8325 8465 8355 8495
rect 8325 8405 8355 8435
rect 8325 8340 8355 8370
rect 8325 8270 8355 8300
rect 8325 8200 8355 8230
rect 8325 8130 8355 8160
rect 8325 8065 8355 8095
rect 8325 8005 8355 8035
rect 8325 7940 8355 7970
rect 8325 7870 8355 7900
rect 8325 7800 8355 7830
rect 8325 7730 8355 7760
rect 8325 7665 8355 7695
rect 8325 7605 8355 7635
rect 8325 7540 8355 7570
rect 8325 7470 8355 7500
rect 8325 7400 8355 7430
rect 8325 7330 8355 7360
rect 8325 7265 8355 7295
rect 8325 7205 8355 7235
rect 8325 7140 8355 7170
rect 8325 7070 8355 7100
rect 8325 7000 8355 7030
rect 8325 6930 8355 6960
rect 8325 6865 8355 6895
rect 8325 6805 8355 6835
rect 8325 6740 8355 6770
rect 8325 6670 8355 6700
rect 8325 6600 8355 6630
rect 8325 6530 8355 6560
rect 8325 6465 8355 6495
rect 8675 9605 8705 9635
rect 8675 9540 8705 9570
rect 8675 9470 8705 9500
rect 8675 9400 8705 9430
rect 8675 9330 8705 9360
rect 8675 9265 8705 9295
rect 8675 9205 8705 9235
rect 8675 9140 8705 9170
rect 8675 9070 8705 9100
rect 8675 9000 8705 9030
rect 8675 8930 8705 8960
rect 8675 8865 8705 8895
rect 8675 8805 8705 8835
rect 8675 8740 8705 8770
rect 8675 8670 8705 8700
rect 8675 8600 8705 8630
rect 8675 8530 8705 8560
rect 8675 8465 8705 8495
rect 8675 8405 8705 8435
rect 8675 8340 8705 8370
rect 8675 8270 8705 8300
rect 8675 8200 8705 8230
rect 8675 8130 8705 8160
rect 8675 8065 8705 8095
rect 8675 8005 8705 8035
rect 8675 7940 8705 7970
rect 8675 7870 8705 7900
rect 8675 7800 8705 7830
rect 8675 7730 8705 7760
rect 8675 7665 8705 7695
rect 8675 7605 8705 7635
rect 8675 7540 8705 7570
rect 8675 7470 8705 7500
rect 8675 7400 8705 7430
rect 8675 7330 8705 7360
rect 8675 7265 8705 7295
rect 8675 7205 8705 7235
rect 8675 7140 8705 7170
rect 8675 7070 8705 7100
rect 8675 7000 8705 7030
rect 8675 6930 8705 6960
rect 8675 6865 8705 6895
rect 8675 6805 8705 6835
rect 8675 6740 8705 6770
rect 8675 6670 8705 6700
rect 8675 6600 8705 6630
rect 8675 6530 8705 6560
rect 8675 6465 8705 6495
rect 9025 9605 9055 9635
rect 9025 9540 9055 9570
rect 9025 9470 9055 9500
rect 9025 9400 9055 9430
rect 9025 9330 9055 9360
rect 9025 9265 9055 9295
rect 9025 9205 9055 9235
rect 9025 9140 9055 9170
rect 9025 9070 9055 9100
rect 9025 9000 9055 9030
rect 9025 8930 9055 8960
rect 9025 8865 9055 8895
rect 9025 8805 9055 8835
rect 9025 8740 9055 8770
rect 9025 8670 9055 8700
rect 9025 8600 9055 8630
rect 9025 8530 9055 8560
rect 9025 8465 9055 8495
rect 9025 8405 9055 8435
rect 9025 8340 9055 8370
rect 9025 8270 9055 8300
rect 9025 8200 9055 8230
rect 9025 8130 9055 8160
rect 9025 8065 9055 8095
rect 9025 8005 9055 8035
rect 9025 7940 9055 7970
rect 9025 7870 9055 7900
rect 9025 7800 9055 7830
rect 9025 7730 9055 7760
rect 9025 7665 9055 7695
rect 9025 7605 9055 7635
rect 9025 7540 9055 7570
rect 9025 7470 9055 7500
rect 9025 7400 9055 7430
rect 9025 7330 9055 7360
rect 9025 7265 9055 7295
rect 9025 7205 9055 7235
rect 9025 7140 9055 7170
rect 9025 7070 9055 7100
rect 9025 7000 9055 7030
rect 9025 6930 9055 6960
rect 9025 6865 9055 6895
rect 9025 6805 9055 6835
rect 9025 6740 9055 6770
rect 9025 6670 9055 6700
rect 9025 6600 9055 6630
rect 9025 6530 9055 6560
rect 9025 6465 9055 6495
rect -75 -1335 -45 -1305
rect -75 -1400 -45 -1370
rect -75 -1470 -45 -1440
rect -75 -1540 -45 -1510
rect -75 -1610 -45 -1580
rect -75 -1675 -45 -1645
rect -75 -1735 -45 -1705
rect -75 -1800 -45 -1770
rect -75 -1870 -45 -1840
rect -75 -1940 -45 -1910
rect -75 -2010 -45 -1980
rect -75 -2075 -45 -2045
rect -75 -2135 -45 -2105
rect -75 -2200 -45 -2170
rect -75 -2270 -45 -2240
rect -75 -2340 -45 -2310
rect -75 -2410 -45 -2380
rect -75 -2475 -45 -2445
rect -75 -2535 -45 -2505
rect -75 -2600 -45 -2570
rect -75 -2670 -45 -2640
rect -75 -2740 -45 -2710
rect -75 -2810 -45 -2780
rect -75 -2875 -45 -2845
rect -75 -2935 -45 -2905
rect -75 -3000 -45 -2970
rect -75 -3070 -45 -3040
rect -75 -3140 -45 -3110
rect -75 -3210 -45 -3180
rect -75 -3275 -45 -3245
rect -75 -3335 -45 -3305
rect -75 -3400 -45 -3370
rect -75 -3470 -45 -3440
rect -75 -3540 -45 -3510
rect -75 -3610 -45 -3580
rect -75 -3675 -45 -3645
rect -75 -3735 -45 -3705
rect -75 -3800 -45 -3770
rect -75 -3870 -45 -3840
rect -75 -3940 -45 -3910
rect -75 -4010 -45 -3980
rect -75 -4075 -45 -4045
rect -75 -4135 -45 -4105
rect -75 -4200 -45 -4170
rect -75 -4270 -45 -4240
rect -75 -4340 -45 -4310
rect -75 -4410 -45 -4380
rect -75 -4475 -45 -4445
rect 275 -1335 305 -1305
rect 275 -1400 305 -1370
rect 275 -1470 305 -1440
rect 275 -1540 305 -1510
rect 275 -1610 305 -1580
rect 275 -1675 305 -1645
rect 275 -1735 305 -1705
rect 275 -1800 305 -1770
rect 275 -1870 305 -1840
rect 275 -1940 305 -1910
rect 275 -2010 305 -1980
rect 275 -2075 305 -2045
rect 275 -2135 305 -2105
rect 275 -2200 305 -2170
rect 275 -2270 305 -2240
rect 275 -2340 305 -2310
rect 275 -2410 305 -2380
rect 275 -2475 305 -2445
rect 275 -2535 305 -2505
rect 275 -2600 305 -2570
rect 275 -2670 305 -2640
rect 275 -2740 305 -2710
rect 275 -2810 305 -2780
rect 275 -2875 305 -2845
rect 275 -2935 305 -2905
rect 275 -3000 305 -2970
rect 275 -3070 305 -3040
rect 275 -3140 305 -3110
rect 275 -3210 305 -3180
rect 275 -3275 305 -3245
rect 275 -3335 305 -3305
rect 275 -3400 305 -3370
rect 275 -3470 305 -3440
rect 275 -3540 305 -3510
rect 275 -3610 305 -3580
rect 275 -3675 305 -3645
rect 275 -3735 305 -3705
rect 275 -3800 305 -3770
rect 275 -3870 305 -3840
rect 275 -3940 305 -3910
rect 275 -4010 305 -3980
rect 275 -4075 305 -4045
rect 275 -4135 305 -4105
rect 275 -4200 305 -4170
rect 275 -4270 305 -4240
rect 275 -4340 305 -4310
rect 275 -4410 305 -4380
rect 275 -4475 305 -4445
rect 625 -1335 655 -1305
rect 625 -1400 655 -1370
rect 625 -1470 655 -1440
rect 625 -1540 655 -1510
rect 625 -1610 655 -1580
rect 625 -1675 655 -1645
rect 625 -1735 655 -1705
rect 625 -1800 655 -1770
rect 625 -1870 655 -1840
rect 625 -1940 655 -1910
rect 625 -2010 655 -1980
rect 625 -2075 655 -2045
rect 625 -2135 655 -2105
rect 625 -2200 655 -2170
rect 625 -2270 655 -2240
rect 625 -2340 655 -2310
rect 625 -2410 655 -2380
rect 625 -2475 655 -2445
rect 625 -2535 655 -2505
rect 625 -2600 655 -2570
rect 625 -2670 655 -2640
rect 625 -2740 655 -2710
rect 625 -2810 655 -2780
rect 625 -2875 655 -2845
rect 625 -2935 655 -2905
rect 625 -3000 655 -2970
rect 625 -3070 655 -3040
rect 625 -3140 655 -3110
rect 625 -3210 655 -3180
rect 625 -3275 655 -3245
rect 625 -3335 655 -3305
rect 625 -3400 655 -3370
rect 625 -3470 655 -3440
rect 625 -3540 655 -3510
rect 625 -3610 655 -3580
rect 625 -3675 655 -3645
rect 625 -3735 655 -3705
rect 625 -3800 655 -3770
rect 625 -3870 655 -3840
rect 625 -3940 655 -3910
rect 625 -4010 655 -3980
rect 625 -4075 655 -4045
rect 625 -4135 655 -4105
rect 625 -4200 655 -4170
rect 625 -4270 655 -4240
rect 625 -4340 655 -4310
rect 625 -4410 655 -4380
rect 625 -4475 655 -4445
rect 975 -1335 1005 -1305
rect 975 -1400 1005 -1370
rect 975 -1470 1005 -1440
rect 975 -1540 1005 -1510
rect 975 -1610 1005 -1580
rect 975 -1675 1005 -1645
rect 975 -1735 1005 -1705
rect 975 -1800 1005 -1770
rect 975 -1870 1005 -1840
rect 975 -1940 1005 -1910
rect 975 -2010 1005 -1980
rect 975 -2075 1005 -2045
rect 975 -2135 1005 -2105
rect 975 -2200 1005 -2170
rect 975 -2270 1005 -2240
rect 975 -2340 1005 -2310
rect 975 -2410 1005 -2380
rect 975 -2475 1005 -2445
rect 975 -2535 1005 -2505
rect 975 -2600 1005 -2570
rect 975 -2670 1005 -2640
rect 975 -2740 1005 -2710
rect 975 -2810 1005 -2780
rect 975 -2875 1005 -2845
rect 975 -2935 1005 -2905
rect 975 -3000 1005 -2970
rect 975 -3070 1005 -3040
rect 975 -3140 1005 -3110
rect 975 -3210 1005 -3180
rect 975 -3275 1005 -3245
rect 975 -3335 1005 -3305
rect 975 -3400 1005 -3370
rect 975 -3470 1005 -3440
rect 975 -3540 1005 -3510
rect 975 -3610 1005 -3580
rect 975 -3675 1005 -3645
rect 975 -3735 1005 -3705
rect 975 -3800 1005 -3770
rect 975 -3870 1005 -3840
rect 975 -3940 1005 -3910
rect 975 -4010 1005 -3980
rect 975 -4075 1005 -4045
rect 975 -4135 1005 -4105
rect 975 -4200 1005 -4170
rect 975 -4270 1005 -4240
rect 975 -4340 1005 -4310
rect 975 -4410 1005 -4380
rect 975 -4475 1005 -4445
rect 1325 -1335 1355 -1305
rect 1325 -1400 1355 -1370
rect 1325 -1470 1355 -1440
rect 1325 -1540 1355 -1510
rect 1325 -1610 1355 -1580
rect 1325 -1675 1355 -1645
rect 1325 -1735 1355 -1705
rect 1325 -1800 1355 -1770
rect 1325 -1870 1355 -1840
rect 1325 -1940 1355 -1910
rect 1325 -2010 1355 -1980
rect 1325 -2075 1355 -2045
rect 1325 -2135 1355 -2105
rect 1325 -2200 1355 -2170
rect 1325 -2270 1355 -2240
rect 1325 -2340 1355 -2310
rect 1325 -2410 1355 -2380
rect 1325 -2475 1355 -2445
rect 1325 -2535 1355 -2505
rect 1325 -2600 1355 -2570
rect 1325 -2670 1355 -2640
rect 1325 -2740 1355 -2710
rect 1325 -2810 1355 -2780
rect 1325 -2875 1355 -2845
rect 1325 -2935 1355 -2905
rect 1325 -3000 1355 -2970
rect 1325 -3070 1355 -3040
rect 1325 -3140 1355 -3110
rect 1325 -3210 1355 -3180
rect 1325 -3275 1355 -3245
rect 1325 -3335 1355 -3305
rect 1325 -3400 1355 -3370
rect 1325 -3470 1355 -3440
rect 1325 -3540 1355 -3510
rect 1325 -3610 1355 -3580
rect 1325 -3675 1355 -3645
rect 1325 -3735 1355 -3705
rect 1325 -3800 1355 -3770
rect 1325 -3870 1355 -3840
rect 1325 -3940 1355 -3910
rect 1325 -4010 1355 -3980
rect 1325 -4075 1355 -4045
rect 1325 -4135 1355 -4105
rect 1325 -4200 1355 -4170
rect 1325 -4270 1355 -4240
rect 1325 -4340 1355 -4310
rect 1325 -4410 1355 -4380
rect 1325 -4475 1355 -4445
rect 1675 -1335 1705 -1305
rect 1675 -1400 1705 -1370
rect 1675 -1470 1705 -1440
rect 1675 -1540 1705 -1510
rect 1675 -1610 1705 -1580
rect 1675 -1675 1705 -1645
rect 1675 -1735 1705 -1705
rect 1675 -1800 1705 -1770
rect 1675 -1870 1705 -1840
rect 1675 -1940 1705 -1910
rect 1675 -2010 1705 -1980
rect 1675 -2075 1705 -2045
rect 1675 -2135 1705 -2105
rect 1675 -2200 1705 -2170
rect 1675 -2270 1705 -2240
rect 1675 -2340 1705 -2310
rect 1675 -2410 1705 -2380
rect 1675 -2475 1705 -2445
rect 1675 -2535 1705 -2505
rect 1675 -2600 1705 -2570
rect 1675 -2670 1705 -2640
rect 1675 -2740 1705 -2710
rect 1675 -2810 1705 -2780
rect 1675 -2875 1705 -2845
rect 1675 -2935 1705 -2905
rect 1675 -3000 1705 -2970
rect 1675 -3070 1705 -3040
rect 1675 -3140 1705 -3110
rect 1675 -3210 1705 -3180
rect 1675 -3275 1705 -3245
rect 1675 -3335 1705 -3305
rect 1675 -3400 1705 -3370
rect 1675 -3470 1705 -3440
rect 1675 -3540 1705 -3510
rect 1675 -3610 1705 -3580
rect 1675 -3675 1705 -3645
rect 1675 -3735 1705 -3705
rect 1675 -3800 1705 -3770
rect 1675 -3870 1705 -3840
rect 1675 -3940 1705 -3910
rect 1675 -4010 1705 -3980
rect 1675 -4075 1705 -4045
rect 1675 -4135 1705 -4105
rect 1675 -4200 1705 -4170
rect 1675 -4270 1705 -4240
rect 1675 -4340 1705 -4310
rect 1675 -4410 1705 -4380
rect 1675 -4475 1705 -4445
rect 2025 -1335 2055 -1305
rect 2025 -1400 2055 -1370
rect 2025 -1470 2055 -1440
rect 2025 -1540 2055 -1510
rect 2025 -1610 2055 -1580
rect 2025 -1675 2055 -1645
rect 2025 -1735 2055 -1705
rect 2025 -1800 2055 -1770
rect 2025 -1870 2055 -1840
rect 2025 -1940 2055 -1910
rect 2025 -2010 2055 -1980
rect 2025 -2075 2055 -2045
rect 2025 -2135 2055 -2105
rect 2025 -2200 2055 -2170
rect 2025 -2270 2055 -2240
rect 2025 -2340 2055 -2310
rect 2025 -2410 2055 -2380
rect 2025 -2475 2055 -2445
rect 2025 -2535 2055 -2505
rect 2025 -2600 2055 -2570
rect 2025 -2670 2055 -2640
rect 2025 -2740 2055 -2710
rect 2025 -2810 2055 -2780
rect 2025 -2875 2055 -2845
rect 2025 -2935 2055 -2905
rect 2025 -3000 2055 -2970
rect 2025 -3070 2055 -3040
rect 2025 -3140 2055 -3110
rect 2025 -3210 2055 -3180
rect 2025 -3275 2055 -3245
rect 2025 -3335 2055 -3305
rect 2025 -3400 2055 -3370
rect 2025 -3470 2055 -3440
rect 2025 -3540 2055 -3510
rect 2025 -3610 2055 -3580
rect 2025 -3675 2055 -3645
rect 2025 -3735 2055 -3705
rect 2025 -3800 2055 -3770
rect 2025 -3870 2055 -3840
rect 2025 -3940 2055 -3910
rect 2025 -4010 2055 -3980
rect 2025 -4075 2055 -4045
rect 2025 -4135 2055 -4105
rect 2025 -4200 2055 -4170
rect 2025 -4270 2055 -4240
rect 2025 -4340 2055 -4310
rect 2025 -4410 2055 -4380
rect 2025 -4475 2055 -4445
rect 2375 -1335 2405 -1305
rect 2375 -1400 2405 -1370
rect 2375 -1470 2405 -1440
rect 2375 -1540 2405 -1510
rect 2375 -1610 2405 -1580
rect 2375 -1675 2405 -1645
rect 2375 -1735 2405 -1705
rect 2375 -1800 2405 -1770
rect 2375 -1870 2405 -1840
rect 2375 -1940 2405 -1910
rect 2375 -2010 2405 -1980
rect 2375 -2075 2405 -2045
rect 2375 -2135 2405 -2105
rect 2375 -2200 2405 -2170
rect 2375 -2270 2405 -2240
rect 2375 -2340 2405 -2310
rect 2375 -2410 2405 -2380
rect 2375 -2475 2405 -2445
rect 2375 -2535 2405 -2505
rect 2375 -2600 2405 -2570
rect 2375 -2670 2405 -2640
rect 2375 -2740 2405 -2710
rect 2375 -2810 2405 -2780
rect 2375 -2875 2405 -2845
rect 2375 -2935 2405 -2905
rect 2375 -3000 2405 -2970
rect 2375 -3070 2405 -3040
rect 2375 -3140 2405 -3110
rect 2375 -3210 2405 -3180
rect 2375 -3275 2405 -3245
rect 2375 -3335 2405 -3305
rect 2375 -3400 2405 -3370
rect 2375 -3470 2405 -3440
rect 2375 -3540 2405 -3510
rect 2375 -3610 2405 -3580
rect 2375 -3675 2405 -3645
rect 2375 -3735 2405 -3705
rect 2375 -3800 2405 -3770
rect 2375 -3870 2405 -3840
rect 2375 -3940 2405 -3910
rect 2375 -4010 2405 -3980
rect 2375 -4075 2405 -4045
rect 2375 -4135 2405 -4105
rect 2375 -4200 2405 -4170
rect 2375 -4270 2405 -4240
rect 2375 -4340 2405 -4310
rect 2375 -4410 2405 -4380
rect 2375 -4475 2405 -4445
rect 2725 -1335 2755 -1305
rect 2725 -1400 2755 -1370
rect 2725 -1470 2755 -1440
rect 2725 -1540 2755 -1510
rect 2725 -1610 2755 -1580
rect 2725 -1675 2755 -1645
rect 2725 -1735 2755 -1705
rect 2725 -1800 2755 -1770
rect 2725 -1870 2755 -1840
rect 2725 -1940 2755 -1910
rect 2725 -2010 2755 -1980
rect 2725 -2075 2755 -2045
rect 2725 -2135 2755 -2105
rect 2725 -2200 2755 -2170
rect 2725 -2270 2755 -2240
rect 2725 -2340 2755 -2310
rect 2725 -2410 2755 -2380
rect 2725 -2475 2755 -2445
rect 2725 -2535 2755 -2505
rect 2725 -2600 2755 -2570
rect 2725 -2670 2755 -2640
rect 2725 -2740 2755 -2710
rect 2725 -2810 2755 -2780
rect 2725 -2875 2755 -2845
rect 2725 -2935 2755 -2905
rect 2725 -3000 2755 -2970
rect 2725 -3070 2755 -3040
rect 2725 -3140 2755 -3110
rect 2725 -3210 2755 -3180
rect 2725 -3275 2755 -3245
rect 2725 -3335 2755 -3305
rect 2725 -3400 2755 -3370
rect 2725 -3470 2755 -3440
rect 2725 -3540 2755 -3510
rect 2725 -3610 2755 -3580
rect 2725 -3675 2755 -3645
rect 2725 -3735 2755 -3705
rect 2725 -3800 2755 -3770
rect 2725 -3870 2755 -3840
rect 2725 -3940 2755 -3910
rect 2725 -4010 2755 -3980
rect 2725 -4075 2755 -4045
rect 2725 -4135 2755 -4105
rect 2725 -4200 2755 -4170
rect 2725 -4270 2755 -4240
rect 2725 -4340 2755 -4310
rect 2725 -4410 2755 -4380
rect 2725 -4475 2755 -4445
rect 3075 -1335 3105 -1305
rect 3075 -1400 3105 -1370
rect 3075 -1470 3105 -1440
rect 3075 -1540 3105 -1510
rect 3075 -1610 3105 -1580
rect 3075 -1675 3105 -1645
rect 3075 -1735 3105 -1705
rect 3075 -1800 3105 -1770
rect 3075 -1870 3105 -1840
rect 3075 -1940 3105 -1910
rect 3075 -2010 3105 -1980
rect 3075 -2075 3105 -2045
rect 3075 -2135 3105 -2105
rect 3075 -2200 3105 -2170
rect 3075 -2270 3105 -2240
rect 3075 -2340 3105 -2310
rect 3075 -2410 3105 -2380
rect 3075 -2475 3105 -2445
rect 3075 -2535 3105 -2505
rect 3075 -2600 3105 -2570
rect 3075 -2670 3105 -2640
rect 3075 -2740 3105 -2710
rect 3075 -2810 3105 -2780
rect 3075 -2875 3105 -2845
rect 3075 -2935 3105 -2905
rect 3075 -3000 3105 -2970
rect 3075 -3070 3105 -3040
rect 3075 -3140 3105 -3110
rect 3075 -3210 3105 -3180
rect 3075 -3275 3105 -3245
rect 3075 -3335 3105 -3305
rect 3075 -3400 3105 -3370
rect 3075 -3470 3105 -3440
rect 3075 -3540 3105 -3510
rect 3075 -3610 3105 -3580
rect 3075 -3675 3105 -3645
rect 3075 -3735 3105 -3705
rect 3075 -3800 3105 -3770
rect 3075 -3870 3105 -3840
rect 3075 -3940 3105 -3910
rect 3075 -4010 3105 -3980
rect 3075 -4075 3105 -4045
rect 3075 -4135 3105 -4105
rect 3075 -4200 3105 -4170
rect 3075 -4270 3105 -4240
rect 3075 -4340 3105 -4310
rect 3075 -4410 3105 -4380
rect 3075 -4475 3105 -4445
rect 3425 -1335 3455 -1305
rect 3425 -1400 3455 -1370
rect 3425 -1470 3455 -1440
rect 3425 -1540 3455 -1510
rect 3425 -1610 3455 -1580
rect 3425 -1675 3455 -1645
rect 3425 -1735 3455 -1705
rect 3425 -1800 3455 -1770
rect 3425 -1870 3455 -1840
rect 3425 -1940 3455 -1910
rect 3425 -2010 3455 -1980
rect 3425 -2075 3455 -2045
rect 3425 -2135 3455 -2105
rect 3425 -2200 3455 -2170
rect 3425 -2270 3455 -2240
rect 3425 -2340 3455 -2310
rect 3425 -2410 3455 -2380
rect 3425 -2475 3455 -2445
rect 3425 -2535 3455 -2505
rect 3425 -2600 3455 -2570
rect 3425 -2670 3455 -2640
rect 3425 -2740 3455 -2710
rect 3425 -2810 3455 -2780
rect 3425 -2875 3455 -2845
rect 3425 -2935 3455 -2905
rect 3425 -3000 3455 -2970
rect 3425 -3070 3455 -3040
rect 3425 -3140 3455 -3110
rect 3425 -3210 3455 -3180
rect 3425 -3275 3455 -3245
rect 3425 -3335 3455 -3305
rect 3425 -3400 3455 -3370
rect 3425 -3470 3455 -3440
rect 3425 -3540 3455 -3510
rect 3425 -3610 3455 -3580
rect 3425 -3675 3455 -3645
rect 3425 -3735 3455 -3705
rect 3425 -3800 3455 -3770
rect 3425 -3870 3455 -3840
rect 3425 -3940 3455 -3910
rect 3425 -4010 3455 -3980
rect 3425 -4075 3455 -4045
rect 3425 -4135 3455 -4105
rect 3425 -4200 3455 -4170
rect 3425 -4270 3455 -4240
rect 3425 -4340 3455 -4310
rect 3425 -4410 3455 -4380
rect 3425 -4475 3455 -4445
rect 3775 -1335 3805 -1305
rect 3775 -1400 3805 -1370
rect 3775 -1470 3805 -1440
rect 3775 -1540 3805 -1510
rect 3775 -1610 3805 -1580
rect 3775 -1675 3805 -1645
rect 3775 -1735 3805 -1705
rect 3775 -1800 3805 -1770
rect 3775 -1870 3805 -1840
rect 3775 -1940 3805 -1910
rect 3775 -2010 3805 -1980
rect 3775 -2075 3805 -2045
rect 3775 -2135 3805 -2105
rect 3775 -2200 3805 -2170
rect 3775 -2270 3805 -2240
rect 3775 -2340 3805 -2310
rect 3775 -2410 3805 -2380
rect 3775 -2475 3805 -2445
rect 3775 -2535 3805 -2505
rect 3775 -2600 3805 -2570
rect 3775 -2670 3805 -2640
rect 3775 -2740 3805 -2710
rect 3775 -2810 3805 -2780
rect 3775 -2875 3805 -2845
rect 3775 -2935 3805 -2905
rect 3775 -3000 3805 -2970
rect 3775 -3070 3805 -3040
rect 3775 -3140 3805 -3110
rect 3775 -3210 3805 -3180
rect 3775 -3275 3805 -3245
rect 3775 -3335 3805 -3305
rect 3775 -3400 3805 -3370
rect 3775 -3470 3805 -3440
rect 3775 -3540 3805 -3510
rect 3775 -3610 3805 -3580
rect 3775 -3675 3805 -3645
rect 3775 -3735 3805 -3705
rect 3775 -3800 3805 -3770
rect 3775 -3870 3805 -3840
rect 3775 -3940 3805 -3910
rect 3775 -4010 3805 -3980
rect 3775 -4075 3805 -4045
rect 3775 -4135 3805 -4105
rect 3775 -4200 3805 -4170
rect 3775 -4270 3805 -4240
rect 3775 -4340 3805 -4310
rect 3775 -4410 3805 -4380
rect 3775 -4475 3805 -4445
rect 4125 -1335 4155 -1305
rect 4125 -1400 4155 -1370
rect 4125 -1470 4155 -1440
rect 4125 -1540 4155 -1510
rect 4125 -1610 4155 -1580
rect 4125 -1675 4155 -1645
rect 4125 -1735 4155 -1705
rect 4125 -1800 4155 -1770
rect 4125 -1870 4155 -1840
rect 4125 -1940 4155 -1910
rect 4125 -2010 4155 -1980
rect 4125 -2075 4155 -2045
rect 4125 -2135 4155 -2105
rect 4125 -2200 4155 -2170
rect 4125 -2270 4155 -2240
rect 4125 -2340 4155 -2310
rect 4125 -2410 4155 -2380
rect 4125 -2475 4155 -2445
rect 4125 -2535 4155 -2505
rect 4125 -2600 4155 -2570
rect 4125 -2670 4155 -2640
rect 4125 -2740 4155 -2710
rect 4125 -2810 4155 -2780
rect 4125 -2875 4155 -2845
rect 4125 -2935 4155 -2905
rect 4125 -3000 4155 -2970
rect 4125 -3070 4155 -3040
rect 4125 -3140 4155 -3110
rect 4125 -3210 4155 -3180
rect 4125 -3275 4155 -3245
rect 4125 -3335 4155 -3305
rect 4125 -3400 4155 -3370
rect 4125 -3470 4155 -3440
rect 4125 -3540 4155 -3510
rect 4125 -3610 4155 -3580
rect 4125 -3675 4155 -3645
rect 4125 -3735 4155 -3705
rect 4125 -3800 4155 -3770
rect 4125 -3870 4155 -3840
rect 4125 -3940 4155 -3910
rect 4125 -4010 4155 -3980
rect 4125 -4075 4155 -4045
rect 4125 -4135 4155 -4105
rect 4125 -4200 4155 -4170
rect 4125 -4270 4155 -4240
rect 4125 -4340 4155 -4310
rect 4125 -4410 4155 -4380
rect 4125 -4475 4155 -4445
rect 4475 -1335 4505 -1305
rect 4475 -1400 4505 -1370
rect 4475 -1470 4505 -1440
rect 4475 -1540 4505 -1510
rect 4475 -1610 4505 -1580
rect 4475 -1675 4505 -1645
rect 4475 -1735 4505 -1705
rect 4475 -1800 4505 -1770
rect 4475 -1870 4505 -1840
rect 4475 -1940 4505 -1910
rect 4475 -2010 4505 -1980
rect 4475 -2075 4505 -2045
rect 4475 -2135 4505 -2105
rect 4475 -2200 4505 -2170
rect 4475 -2270 4505 -2240
rect 4475 -2340 4505 -2310
rect 4475 -2410 4505 -2380
rect 4475 -2475 4505 -2445
rect 4475 -2535 4505 -2505
rect 4475 -2600 4505 -2570
rect 4475 -2670 4505 -2640
rect 4475 -2740 4505 -2710
rect 4475 -2810 4505 -2780
rect 4475 -2875 4505 -2845
rect 4475 -2935 4505 -2905
rect 4475 -3000 4505 -2970
rect 4475 -3070 4505 -3040
rect 4475 -3140 4505 -3110
rect 4475 -3210 4505 -3180
rect 4475 -3275 4505 -3245
rect 4475 -3335 4505 -3305
rect 4475 -3400 4505 -3370
rect 4475 -3470 4505 -3440
rect 4475 -3540 4505 -3510
rect 4475 -3610 4505 -3580
rect 4475 -3675 4505 -3645
rect 4475 -3735 4505 -3705
rect 4475 -3800 4505 -3770
rect 4475 -3870 4505 -3840
rect 4475 -3940 4505 -3910
rect 4475 -4010 4505 -3980
rect 4475 -4075 4505 -4045
rect 4475 -4135 4505 -4105
rect 4475 -4200 4505 -4170
rect 4475 -4270 4505 -4240
rect 4475 -4340 4505 -4310
rect 4475 -4410 4505 -4380
rect 4475 -4475 4505 -4445
rect 4825 -1335 4855 -1305
rect 4825 -1400 4855 -1370
rect 4825 -1470 4855 -1440
rect 4825 -1540 4855 -1510
rect 4825 -1610 4855 -1580
rect 4825 -1675 4855 -1645
rect 4825 -1735 4855 -1705
rect 4825 -1800 4855 -1770
rect 4825 -1870 4855 -1840
rect 4825 -1940 4855 -1910
rect 4825 -2010 4855 -1980
rect 4825 -2075 4855 -2045
rect 4825 -2135 4855 -2105
rect 4825 -2200 4855 -2170
rect 4825 -2270 4855 -2240
rect 4825 -2340 4855 -2310
rect 4825 -2410 4855 -2380
rect 4825 -2475 4855 -2445
rect 4825 -2535 4855 -2505
rect 4825 -2600 4855 -2570
rect 4825 -2670 4855 -2640
rect 4825 -2740 4855 -2710
rect 4825 -2810 4855 -2780
rect 4825 -2875 4855 -2845
rect 4825 -2935 4855 -2905
rect 4825 -3000 4855 -2970
rect 4825 -3070 4855 -3040
rect 4825 -3140 4855 -3110
rect 4825 -3210 4855 -3180
rect 4825 -3275 4855 -3245
rect 4825 -3335 4855 -3305
rect 4825 -3400 4855 -3370
rect 4825 -3470 4855 -3440
rect 4825 -3540 4855 -3510
rect 4825 -3610 4855 -3580
rect 4825 -3675 4855 -3645
rect 4825 -3735 4855 -3705
rect 4825 -3800 4855 -3770
rect 4825 -3870 4855 -3840
rect 4825 -3940 4855 -3910
rect 4825 -4010 4855 -3980
rect 4825 -4075 4855 -4045
rect 4825 -4135 4855 -4105
rect 4825 -4200 4855 -4170
rect 4825 -4270 4855 -4240
rect 4825 -4340 4855 -4310
rect 4825 -4410 4855 -4380
rect 4825 -4475 4855 -4445
rect 5175 -1335 5205 -1305
rect 5175 -1400 5205 -1370
rect 5175 -1470 5205 -1440
rect 5175 -1540 5205 -1510
rect 5175 -1610 5205 -1580
rect 5175 -1675 5205 -1645
rect 5175 -1735 5205 -1705
rect 5175 -1800 5205 -1770
rect 5175 -1870 5205 -1840
rect 5175 -1940 5205 -1910
rect 5175 -2010 5205 -1980
rect 5175 -2075 5205 -2045
rect 5175 -2135 5205 -2105
rect 5175 -2200 5205 -2170
rect 5175 -2270 5205 -2240
rect 5175 -2340 5205 -2310
rect 5175 -2410 5205 -2380
rect 5175 -2475 5205 -2445
rect 5175 -2535 5205 -2505
rect 5175 -2600 5205 -2570
rect 5175 -2670 5205 -2640
rect 5175 -2740 5205 -2710
rect 5175 -2810 5205 -2780
rect 5175 -2875 5205 -2845
rect 5175 -2935 5205 -2905
rect 5175 -3000 5205 -2970
rect 5175 -3070 5205 -3040
rect 5175 -3140 5205 -3110
rect 5175 -3210 5205 -3180
rect 5175 -3275 5205 -3245
rect 5175 -3335 5205 -3305
rect 5175 -3400 5205 -3370
rect 5175 -3470 5205 -3440
rect 5175 -3540 5205 -3510
rect 5175 -3610 5205 -3580
rect 5175 -3675 5205 -3645
rect 5175 -3735 5205 -3705
rect 5175 -3800 5205 -3770
rect 5175 -3870 5205 -3840
rect 5175 -3940 5205 -3910
rect 5175 -4010 5205 -3980
rect 5175 -4075 5205 -4045
rect 5175 -4135 5205 -4105
rect 5175 -4200 5205 -4170
rect 5175 -4270 5205 -4240
rect 5175 -4340 5205 -4310
rect 5175 -4410 5205 -4380
rect 5175 -4475 5205 -4445
rect 5525 -1335 5555 -1305
rect 5525 -1400 5555 -1370
rect 5525 -1470 5555 -1440
rect 5525 -1540 5555 -1510
rect 5525 -1610 5555 -1580
rect 5525 -1675 5555 -1645
rect 5525 -1735 5555 -1705
rect 5525 -1800 5555 -1770
rect 5525 -1870 5555 -1840
rect 5525 -1940 5555 -1910
rect 5525 -2010 5555 -1980
rect 5525 -2075 5555 -2045
rect 5525 -2135 5555 -2105
rect 5525 -2200 5555 -2170
rect 5525 -2270 5555 -2240
rect 5525 -2340 5555 -2310
rect 5525 -2410 5555 -2380
rect 5525 -2475 5555 -2445
rect 5525 -2535 5555 -2505
rect 5525 -2600 5555 -2570
rect 5525 -2670 5555 -2640
rect 5525 -2740 5555 -2710
rect 5525 -2810 5555 -2780
rect 5525 -2875 5555 -2845
rect 5525 -2935 5555 -2905
rect 5525 -3000 5555 -2970
rect 5525 -3070 5555 -3040
rect 5525 -3140 5555 -3110
rect 5525 -3210 5555 -3180
rect 5525 -3275 5555 -3245
rect 5525 -3335 5555 -3305
rect 5525 -3400 5555 -3370
rect 5525 -3470 5555 -3440
rect 5525 -3540 5555 -3510
rect 5525 -3610 5555 -3580
rect 5525 -3675 5555 -3645
rect 5525 -3735 5555 -3705
rect 5525 -3800 5555 -3770
rect 5525 -3870 5555 -3840
rect 5525 -3940 5555 -3910
rect 5525 -4010 5555 -3980
rect 5525 -4075 5555 -4045
rect 5525 -4135 5555 -4105
rect 5525 -4200 5555 -4170
rect 5525 -4270 5555 -4240
rect 5525 -4340 5555 -4310
rect 5525 -4410 5555 -4380
rect 5525 -4475 5555 -4445
rect 5875 -1335 5905 -1305
rect 5875 -1400 5905 -1370
rect 5875 -1470 5905 -1440
rect 5875 -1540 5905 -1510
rect 5875 -1610 5905 -1580
rect 5875 -1675 5905 -1645
rect 5875 -1735 5905 -1705
rect 5875 -1800 5905 -1770
rect 5875 -1870 5905 -1840
rect 5875 -1940 5905 -1910
rect 5875 -2010 5905 -1980
rect 5875 -2075 5905 -2045
rect 5875 -2135 5905 -2105
rect 5875 -2200 5905 -2170
rect 5875 -2270 5905 -2240
rect 5875 -2340 5905 -2310
rect 5875 -2410 5905 -2380
rect 5875 -2475 5905 -2445
rect 5875 -2535 5905 -2505
rect 5875 -2600 5905 -2570
rect 5875 -2670 5905 -2640
rect 5875 -2740 5905 -2710
rect 5875 -2810 5905 -2780
rect 5875 -2875 5905 -2845
rect 5875 -2935 5905 -2905
rect 5875 -3000 5905 -2970
rect 5875 -3070 5905 -3040
rect 5875 -3140 5905 -3110
rect 5875 -3210 5905 -3180
rect 5875 -3275 5905 -3245
rect 5875 -3335 5905 -3305
rect 5875 -3400 5905 -3370
rect 5875 -3470 5905 -3440
rect 5875 -3540 5905 -3510
rect 5875 -3610 5905 -3580
rect 5875 -3675 5905 -3645
rect 5875 -3735 5905 -3705
rect 5875 -3800 5905 -3770
rect 5875 -3870 5905 -3840
rect 5875 -3940 5905 -3910
rect 5875 -4010 5905 -3980
rect 5875 -4075 5905 -4045
rect 5875 -4135 5905 -4105
rect 5875 -4200 5905 -4170
rect 5875 -4270 5905 -4240
rect 5875 -4340 5905 -4310
rect 5875 -4410 5905 -4380
rect 5875 -4475 5905 -4445
rect 6225 -1335 6255 -1305
rect 6225 -1400 6255 -1370
rect 6225 -1470 6255 -1440
rect 6225 -1540 6255 -1510
rect 6225 -1610 6255 -1580
rect 6225 -1675 6255 -1645
rect 6225 -1735 6255 -1705
rect 6225 -1800 6255 -1770
rect 6225 -1870 6255 -1840
rect 6225 -1940 6255 -1910
rect 6225 -2010 6255 -1980
rect 6225 -2075 6255 -2045
rect 6225 -2135 6255 -2105
rect 6225 -2200 6255 -2170
rect 6225 -2270 6255 -2240
rect 6225 -2340 6255 -2310
rect 6225 -2410 6255 -2380
rect 6225 -2475 6255 -2445
rect 6225 -2535 6255 -2505
rect 6225 -2600 6255 -2570
rect 6225 -2670 6255 -2640
rect 6225 -2740 6255 -2710
rect 6225 -2810 6255 -2780
rect 6225 -2875 6255 -2845
rect 6225 -2935 6255 -2905
rect 6225 -3000 6255 -2970
rect 6225 -3070 6255 -3040
rect 6225 -3140 6255 -3110
rect 6225 -3210 6255 -3180
rect 6225 -3275 6255 -3245
rect 6225 -3335 6255 -3305
rect 6225 -3400 6255 -3370
rect 6225 -3470 6255 -3440
rect 6225 -3540 6255 -3510
rect 6225 -3610 6255 -3580
rect 6225 -3675 6255 -3645
rect 6225 -3735 6255 -3705
rect 6225 -3800 6255 -3770
rect 6225 -3870 6255 -3840
rect 6225 -3940 6255 -3910
rect 6225 -4010 6255 -3980
rect 6225 -4075 6255 -4045
rect 6225 -4135 6255 -4105
rect 6225 -4200 6255 -4170
rect 6225 -4270 6255 -4240
rect 6225 -4340 6255 -4310
rect 6225 -4410 6255 -4380
rect 6225 -4475 6255 -4445
rect 6575 -1335 6605 -1305
rect 6575 -1400 6605 -1370
rect 6575 -1470 6605 -1440
rect 6575 -1540 6605 -1510
rect 6575 -1610 6605 -1580
rect 6575 -1675 6605 -1645
rect 6575 -1735 6605 -1705
rect 6575 -1800 6605 -1770
rect 6575 -1870 6605 -1840
rect 6575 -1940 6605 -1910
rect 6575 -2010 6605 -1980
rect 6575 -2075 6605 -2045
rect 6575 -2135 6605 -2105
rect 6575 -2200 6605 -2170
rect 6575 -2270 6605 -2240
rect 6575 -2340 6605 -2310
rect 6575 -2410 6605 -2380
rect 6575 -2475 6605 -2445
rect 6575 -2535 6605 -2505
rect 6575 -2600 6605 -2570
rect 6575 -2670 6605 -2640
rect 6575 -2740 6605 -2710
rect 6575 -2810 6605 -2780
rect 6575 -2875 6605 -2845
rect 6575 -2935 6605 -2905
rect 6575 -3000 6605 -2970
rect 6575 -3070 6605 -3040
rect 6575 -3140 6605 -3110
rect 6575 -3210 6605 -3180
rect 6575 -3275 6605 -3245
rect 6575 -3335 6605 -3305
rect 6575 -3400 6605 -3370
rect 6575 -3470 6605 -3440
rect 6575 -3540 6605 -3510
rect 6575 -3610 6605 -3580
rect 6575 -3675 6605 -3645
rect 6575 -3735 6605 -3705
rect 6575 -3800 6605 -3770
rect 6575 -3870 6605 -3840
rect 6575 -3940 6605 -3910
rect 6575 -4010 6605 -3980
rect 6575 -4075 6605 -4045
rect 6575 -4135 6605 -4105
rect 6575 -4200 6605 -4170
rect 6575 -4270 6605 -4240
rect 6575 -4340 6605 -4310
rect 6575 -4410 6605 -4380
rect 6575 -4475 6605 -4445
rect 6925 -1335 6955 -1305
rect 6925 -1400 6955 -1370
rect 6925 -1470 6955 -1440
rect 6925 -1540 6955 -1510
rect 6925 -1610 6955 -1580
rect 6925 -1675 6955 -1645
rect 6925 -1735 6955 -1705
rect 6925 -1800 6955 -1770
rect 6925 -1870 6955 -1840
rect 6925 -1940 6955 -1910
rect 6925 -2010 6955 -1980
rect 6925 -2075 6955 -2045
rect 6925 -2135 6955 -2105
rect 6925 -2200 6955 -2170
rect 6925 -2270 6955 -2240
rect 6925 -2340 6955 -2310
rect 6925 -2410 6955 -2380
rect 6925 -2475 6955 -2445
rect 6925 -2535 6955 -2505
rect 6925 -2600 6955 -2570
rect 6925 -2670 6955 -2640
rect 6925 -2740 6955 -2710
rect 6925 -2810 6955 -2780
rect 6925 -2875 6955 -2845
rect 6925 -2935 6955 -2905
rect 6925 -3000 6955 -2970
rect 6925 -3070 6955 -3040
rect 6925 -3140 6955 -3110
rect 6925 -3210 6955 -3180
rect 6925 -3275 6955 -3245
rect 6925 -3335 6955 -3305
rect 6925 -3400 6955 -3370
rect 6925 -3470 6955 -3440
rect 6925 -3540 6955 -3510
rect 6925 -3610 6955 -3580
rect 6925 -3675 6955 -3645
rect 6925 -3735 6955 -3705
rect 6925 -3800 6955 -3770
rect 6925 -3870 6955 -3840
rect 6925 -3940 6955 -3910
rect 6925 -4010 6955 -3980
rect 6925 -4075 6955 -4045
rect 6925 -4135 6955 -4105
rect 6925 -4200 6955 -4170
rect 6925 -4270 6955 -4240
rect 6925 -4340 6955 -4310
rect 6925 -4410 6955 -4380
rect 6925 -4475 6955 -4445
rect 7275 -1335 7305 -1305
rect 7275 -1400 7305 -1370
rect 7275 -1470 7305 -1440
rect 7275 -1540 7305 -1510
rect 7275 -1610 7305 -1580
rect 7275 -1675 7305 -1645
rect 7275 -1735 7305 -1705
rect 7275 -1800 7305 -1770
rect 7275 -1870 7305 -1840
rect 7275 -1940 7305 -1910
rect 7275 -2010 7305 -1980
rect 7275 -2075 7305 -2045
rect 7275 -2135 7305 -2105
rect 7275 -2200 7305 -2170
rect 7275 -2270 7305 -2240
rect 7275 -2340 7305 -2310
rect 7275 -2410 7305 -2380
rect 7275 -2475 7305 -2445
rect 7275 -2535 7305 -2505
rect 7275 -2600 7305 -2570
rect 7275 -2670 7305 -2640
rect 7275 -2740 7305 -2710
rect 7275 -2810 7305 -2780
rect 7275 -2875 7305 -2845
rect 7275 -2935 7305 -2905
rect 7275 -3000 7305 -2970
rect 7275 -3070 7305 -3040
rect 7275 -3140 7305 -3110
rect 7275 -3210 7305 -3180
rect 7275 -3275 7305 -3245
rect 7275 -3335 7305 -3305
rect 7275 -3400 7305 -3370
rect 7275 -3470 7305 -3440
rect 7275 -3540 7305 -3510
rect 7275 -3610 7305 -3580
rect 7275 -3675 7305 -3645
rect 7275 -3735 7305 -3705
rect 7275 -3800 7305 -3770
rect 7275 -3870 7305 -3840
rect 7275 -3940 7305 -3910
rect 7275 -4010 7305 -3980
rect 7275 -4075 7305 -4045
rect 7275 -4135 7305 -4105
rect 7275 -4200 7305 -4170
rect 7275 -4270 7305 -4240
rect 7275 -4340 7305 -4310
rect 7275 -4410 7305 -4380
rect 7275 -4475 7305 -4445
rect 7625 -1335 7655 -1305
rect 7625 -1400 7655 -1370
rect 7625 -1470 7655 -1440
rect 7625 -1540 7655 -1510
rect 7625 -1610 7655 -1580
rect 7625 -1675 7655 -1645
rect 7625 -1735 7655 -1705
rect 7625 -1800 7655 -1770
rect 7625 -1870 7655 -1840
rect 7625 -1940 7655 -1910
rect 7625 -2010 7655 -1980
rect 7625 -2075 7655 -2045
rect 7625 -2135 7655 -2105
rect 7625 -2200 7655 -2170
rect 7625 -2270 7655 -2240
rect 7625 -2340 7655 -2310
rect 7625 -2410 7655 -2380
rect 7625 -2475 7655 -2445
rect 7625 -2535 7655 -2505
rect 7625 -2600 7655 -2570
rect 7625 -2670 7655 -2640
rect 7625 -2740 7655 -2710
rect 7625 -2810 7655 -2780
rect 7625 -2875 7655 -2845
rect 7625 -2935 7655 -2905
rect 7625 -3000 7655 -2970
rect 7625 -3070 7655 -3040
rect 7625 -3140 7655 -3110
rect 7625 -3210 7655 -3180
rect 7625 -3275 7655 -3245
rect 7625 -3335 7655 -3305
rect 7625 -3400 7655 -3370
rect 7625 -3470 7655 -3440
rect 7625 -3540 7655 -3510
rect 7625 -3610 7655 -3580
rect 7625 -3675 7655 -3645
rect 7625 -3735 7655 -3705
rect 7625 -3800 7655 -3770
rect 7625 -3870 7655 -3840
rect 7625 -3940 7655 -3910
rect 7625 -4010 7655 -3980
rect 7625 -4075 7655 -4045
rect 7625 -4135 7655 -4105
rect 7625 -4200 7655 -4170
rect 7625 -4270 7655 -4240
rect 7625 -4340 7655 -4310
rect 7625 -4410 7655 -4380
rect 7625 -4475 7655 -4445
rect 7975 -1335 8005 -1305
rect 7975 -1400 8005 -1370
rect 7975 -1470 8005 -1440
rect 7975 -1540 8005 -1510
rect 7975 -1610 8005 -1580
rect 7975 -1675 8005 -1645
rect 7975 -1735 8005 -1705
rect 7975 -1800 8005 -1770
rect 7975 -1870 8005 -1840
rect 7975 -1940 8005 -1910
rect 7975 -2010 8005 -1980
rect 7975 -2075 8005 -2045
rect 7975 -2135 8005 -2105
rect 7975 -2200 8005 -2170
rect 7975 -2270 8005 -2240
rect 7975 -2340 8005 -2310
rect 7975 -2410 8005 -2380
rect 7975 -2475 8005 -2445
rect 7975 -2535 8005 -2505
rect 7975 -2600 8005 -2570
rect 7975 -2670 8005 -2640
rect 7975 -2740 8005 -2710
rect 7975 -2810 8005 -2780
rect 7975 -2875 8005 -2845
rect 7975 -2935 8005 -2905
rect 7975 -3000 8005 -2970
rect 7975 -3070 8005 -3040
rect 7975 -3140 8005 -3110
rect 7975 -3210 8005 -3180
rect 7975 -3275 8005 -3245
rect 7975 -3335 8005 -3305
rect 7975 -3400 8005 -3370
rect 7975 -3470 8005 -3440
rect 7975 -3540 8005 -3510
rect 7975 -3610 8005 -3580
rect 7975 -3675 8005 -3645
rect 7975 -3735 8005 -3705
rect 7975 -3800 8005 -3770
rect 7975 -3870 8005 -3840
rect 7975 -3940 8005 -3910
rect 7975 -4010 8005 -3980
rect 7975 -4075 8005 -4045
rect 7975 -4135 8005 -4105
rect 7975 -4200 8005 -4170
rect 7975 -4270 8005 -4240
rect 7975 -4340 8005 -4310
rect 7975 -4410 8005 -4380
rect 7975 -4475 8005 -4445
rect 8325 -1335 8355 -1305
rect 8325 -1400 8355 -1370
rect 8325 -1470 8355 -1440
rect 8325 -1540 8355 -1510
rect 8325 -1610 8355 -1580
rect 8325 -1675 8355 -1645
rect 8325 -1735 8355 -1705
rect 8325 -1800 8355 -1770
rect 8325 -1870 8355 -1840
rect 8325 -1940 8355 -1910
rect 8325 -2010 8355 -1980
rect 8325 -2075 8355 -2045
rect 8325 -2135 8355 -2105
rect 8325 -2200 8355 -2170
rect 8325 -2270 8355 -2240
rect 8325 -2340 8355 -2310
rect 8325 -2410 8355 -2380
rect 8325 -2475 8355 -2445
rect 8325 -2535 8355 -2505
rect 8325 -2600 8355 -2570
rect 8325 -2670 8355 -2640
rect 8325 -2740 8355 -2710
rect 8325 -2810 8355 -2780
rect 8325 -2875 8355 -2845
rect 8325 -2935 8355 -2905
rect 8325 -3000 8355 -2970
rect 8325 -3070 8355 -3040
rect 8325 -3140 8355 -3110
rect 8325 -3210 8355 -3180
rect 8325 -3275 8355 -3245
rect 8325 -3335 8355 -3305
rect 8325 -3400 8355 -3370
rect 8325 -3470 8355 -3440
rect 8325 -3540 8355 -3510
rect 8325 -3610 8355 -3580
rect 8325 -3675 8355 -3645
rect 8325 -3735 8355 -3705
rect 8325 -3800 8355 -3770
rect 8325 -3870 8355 -3840
rect 8325 -3940 8355 -3910
rect 8325 -4010 8355 -3980
rect 8325 -4075 8355 -4045
rect 8325 -4135 8355 -4105
rect 8325 -4200 8355 -4170
rect 8325 -4270 8355 -4240
rect 8325 -4340 8355 -4310
rect 8325 -4410 8355 -4380
rect 8325 -4475 8355 -4445
rect 8675 -1335 8705 -1305
rect 8675 -1400 8705 -1370
rect 8675 -1470 8705 -1440
rect 8675 -1540 8705 -1510
rect 8675 -1610 8705 -1580
rect 8675 -1675 8705 -1645
rect 8675 -1735 8705 -1705
rect 8675 -1800 8705 -1770
rect 8675 -1870 8705 -1840
rect 8675 -1940 8705 -1910
rect 8675 -2010 8705 -1980
rect 8675 -2075 8705 -2045
rect 8675 -2135 8705 -2105
rect 8675 -2200 8705 -2170
rect 8675 -2270 8705 -2240
rect 8675 -2340 8705 -2310
rect 8675 -2410 8705 -2380
rect 8675 -2475 8705 -2445
rect 8675 -2535 8705 -2505
rect 8675 -2600 8705 -2570
rect 8675 -2670 8705 -2640
rect 8675 -2740 8705 -2710
rect 8675 -2810 8705 -2780
rect 8675 -2875 8705 -2845
rect 8675 -2935 8705 -2905
rect 8675 -3000 8705 -2970
rect 8675 -3070 8705 -3040
rect 8675 -3140 8705 -3110
rect 8675 -3210 8705 -3180
rect 8675 -3275 8705 -3245
rect 8675 -3335 8705 -3305
rect 8675 -3400 8705 -3370
rect 8675 -3470 8705 -3440
rect 8675 -3540 8705 -3510
rect 8675 -3610 8705 -3580
rect 8675 -3675 8705 -3645
rect 8675 -3735 8705 -3705
rect 8675 -3800 8705 -3770
rect 8675 -3870 8705 -3840
rect 8675 -3940 8705 -3910
rect 8675 -4010 8705 -3980
rect 8675 -4075 8705 -4045
rect 8675 -4135 8705 -4105
rect 8675 -4200 8705 -4170
rect 8675 -4270 8705 -4240
rect 8675 -4340 8705 -4310
rect 8675 -4410 8705 -4380
rect 8675 -4475 8705 -4445
rect 9025 -1335 9055 -1305
rect 9025 -1400 9055 -1370
rect 9025 -1470 9055 -1440
rect 9025 -1540 9055 -1510
rect 9025 -1610 9055 -1580
rect 9025 -1675 9055 -1645
rect 9025 -1735 9055 -1705
rect 9025 -1800 9055 -1770
rect 9025 -1870 9055 -1840
rect 9025 -1940 9055 -1910
rect 9025 -2010 9055 -1980
rect 9025 -2075 9055 -2045
rect 9025 -2135 9055 -2105
rect 9025 -2200 9055 -2170
rect 9025 -2270 9055 -2240
rect 9025 -2340 9055 -2310
rect 9025 -2410 9055 -2380
rect 9025 -2475 9055 -2445
rect 9025 -2535 9055 -2505
rect 9025 -2600 9055 -2570
rect 9025 -2670 9055 -2640
rect 9025 -2740 9055 -2710
rect 9025 -2810 9055 -2780
rect 9025 -2875 9055 -2845
rect 9025 -2935 9055 -2905
rect 9025 -3000 9055 -2970
rect 9025 -3070 9055 -3040
rect 9025 -3140 9055 -3110
rect 9025 -3210 9055 -3180
rect 9025 -3275 9055 -3245
rect 9025 -3335 9055 -3305
rect 9025 -3400 9055 -3370
rect 9025 -3470 9055 -3440
rect 9025 -3540 9055 -3510
rect 9025 -3610 9055 -3580
rect 9025 -3675 9055 -3645
rect 9025 -3735 9055 -3705
rect 9025 -3800 9055 -3770
rect 9025 -3870 9055 -3840
rect 9025 -3940 9055 -3910
rect 9025 -4010 9055 -3980
rect 9025 -4075 9055 -4045
rect 9025 -4135 9055 -4105
rect 9025 -4200 9055 -4170
rect 9025 -4270 9055 -4240
rect 9025 -4340 9055 -4310
rect 9025 -4410 9055 -4380
rect 9025 -4475 9055 -4445
<< metal3 >>
rect 2180 20915 2240 20925
rect 2180 20875 2190 20915
rect 2230 20875 2240 20915
rect 2180 20850 2240 20875
rect 2180 20810 2190 20850
rect 2230 20810 2240 20850
rect 2180 20780 2240 20810
rect 2180 20740 2190 20780
rect 2230 20740 2240 20780
rect 2180 20710 2240 20740
rect 2180 20670 2190 20710
rect 2230 20670 2240 20710
rect 2180 20640 2240 20670
rect 2180 20600 2190 20640
rect 2230 20600 2240 20640
rect 2180 20575 2240 20600
rect 2180 20535 2190 20575
rect 2230 20535 2240 20575
rect 2180 20515 2240 20535
rect 2180 20475 2190 20515
rect 2230 20475 2240 20515
rect 2180 20450 2240 20475
rect 2180 20410 2190 20450
rect 2230 20410 2240 20450
rect 2180 20380 2240 20410
rect 2180 20340 2190 20380
rect 2230 20340 2240 20380
rect 2180 20310 2240 20340
rect 2180 20270 2190 20310
rect 2230 20270 2240 20310
rect 2180 20240 2240 20270
rect 2180 20200 2190 20240
rect 2230 20200 2240 20240
rect 2180 20175 2240 20200
rect 2180 20135 2190 20175
rect 2230 20135 2240 20175
rect 2180 20115 2240 20135
rect 2180 20075 2190 20115
rect 2230 20075 2240 20115
rect 2180 20050 2240 20075
rect 2180 20010 2190 20050
rect 2230 20010 2240 20050
rect 2180 19980 2240 20010
rect 2180 19940 2190 19980
rect 2230 19940 2240 19980
rect 2180 19910 2240 19940
rect 2180 19870 2190 19910
rect 2230 19870 2240 19910
rect 2180 19840 2240 19870
rect 2180 19800 2190 19840
rect 2230 19800 2240 19840
rect 2180 19775 2240 19800
rect 2180 19735 2190 19775
rect 2230 19735 2240 19775
rect 2180 19715 2240 19735
rect 2180 19675 2190 19715
rect 2230 19675 2240 19715
rect 2180 19650 2240 19675
rect 2180 19610 2190 19650
rect 2230 19610 2240 19650
rect 2180 19580 2240 19610
rect 2180 19540 2190 19580
rect 2230 19540 2240 19580
rect 2180 19510 2240 19540
rect 2180 19470 2190 19510
rect 2230 19470 2240 19510
rect 2180 19440 2240 19470
rect 2180 19400 2190 19440
rect 2230 19400 2240 19440
rect 2180 19375 2240 19400
rect 2180 19335 2190 19375
rect 2230 19335 2240 19375
rect 2180 19315 2240 19335
rect 2180 19275 2190 19315
rect 2230 19275 2240 19315
rect 2180 19250 2240 19275
rect 2180 19210 2190 19250
rect 2230 19210 2240 19250
rect 2180 19180 2240 19210
rect 2180 19140 2190 19180
rect 2230 19140 2240 19180
rect 2180 19110 2240 19140
rect 2180 19070 2190 19110
rect 2230 19070 2240 19110
rect 2180 19040 2240 19070
rect 2180 19000 2190 19040
rect 2230 19000 2240 19040
rect 2180 18975 2240 19000
rect 2180 18935 2190 18975
rect 2230 18935 2240 18975
rect 2180 18915 2240 18935
rect 2180 18875 2190 18915
rect 2230 18875 2240 18915
rect 2180 18850 2240 18875
rect 2180 18810 2190 18850
rect 2230 18810 2240 18850
rect 2180 18780 2240 18810
rect 2180 18740 2190 18780
rect 2230 18740 2240 18780
rect 2180 18710 2240 18740
rect 2180 18670 2190 18710
rect 2230 18670 2240 18710
rect 2180 18640 2240 18670
rect 2180 18600 2190 18640
rect 2230 18600 2240 18640
rect 2180 18575 2240 18600
rect 2180 18535 2190 18575
rect 2230 18535 2240 18575
rect 2180 18515 2240 18535
rect 2180 18475 2190 18515
rect 2230 18475 2240 18515
rect 2180 18450 2240 18475
rect 2180 18410 2190 18450
rect 2230 18410 2240 18450
rect 2180 18380 2240 18410
rect 2180 18340 2190 18380
rect 2230 18340 2240 18380
rect 2180 18310 2240 18340
rect 2180 18270 2190 18310
rect 2230 18270 2240 18310
rect 2180 18240 2240 18270
rect 2180 18200 2190 18240
rect 2230 18200 2240 18240
rect 2180 18175 2240 18200
rect 2180 18135 2190 18175
rect 2230 18135 2240 18175
rect 2180 18115 2240 18135
rect 2180 18075 2190 18115
rect 2230 18075 2240 18115
rect 2180 18050 2240 18075
rect 2180 18010 2190 18050
rect 2230 18010 2240 18050
rect 2180 17980 2240 18010
rect 2180 17940 2190 17980
rect 2230 17940 2240 17980
rect 2180 17910 2240 17940
rect 2180 17870 2190 17910
rect 2230 17870 2240 17910
rect 2180 17840 2240 17870
rect 2180 17800 2190 17840
rect 2230 17800 2240 17840
rect 2180 17775 2240 17800
rect 2180 17735 2190 17775
rect 2230 17735 2240 17775
rect 2180 17725 2240 17735
rect 6650 20915 6710 20925
rect 6650 20875 6660 20915
rect 6700 20875 6710 20915
rect 6650 20850 6710 20875
rect 6650 20810 6660 20850
rect 6700 20810 6710 20850
rect 6650 20780 6710 20810
rect 6650 20740 6660 20780
rect 6700 20740 6710 20780
rect 6650 20710 6710 20740
rect 6650 20670 6660 20710
rect 6700 20670 6710 20710
rect 6650 20640 6710 20670
rect 6650 20600 6660 20640
rect 6700 20600 6710 20640
rect 6650 20575 6710 20600
rect 6650 20535 6660 20575
rect 6700 20535 6710 20575
rect 6650 20515 6710 20535
rect 6650 20475 6660 20515
rect 6700 20475 6710 20515
rect 6650 20450 6710 20475
rect 6650 20410 6660 20450
rect 6700 20410 6710 20450
rect 6650 20380 6710 20410
rect 6650 20340 6660 20380
rect 6700 20340 6710 20380
rect 6650 20310 6710 20340
rect 6650 20270 6660 20310
rect 6700 20270 6710 20310
rect 6650 20240 6710 20270
rect 6650 20200 6660 20240
rect 6700 20200 6710 20240
rect 6650 20175 6710 20200
rect 6650 20135 6660 20175
rect 6700 20135 6710 20175
rect 6650 20115 6710 20135
rect 6650 20075 6660 20115
rect 6700 20075 6710 20115
rect 6650 20050 6710 20075
rect 6650 20010 6660 20050
rect 6700 20010 6710 20050
rect 6650 19980 6710 20010
rect 6650 19940 6660 19980
rect 6700 19940 6710 19980
rect 6650 19910 6710 19940
rect 6650 19870 6660 19910
rect 6700 19870 6710 19910
rect 6650 19840 6710 19870
rect 6650 19800 6660 19840
rect 6700 19800 6710 19840
rect 6650 19775 6710 19800
rect 6650 19735 6660 19775
rect 6700 19735 6710 19775
rect 6650 19715 6710 19735
rect 6650 19675 6660 19715
rect 6700 19675 6710 19715
rect 6650 19650 6710 19675
rect 6650 19610 6660 19650
rect 6700 19610 6710 19650
rect 6650 19580 6710 19610
rect 6650 19540 6660 19580
rect 6700 19540 6710 19580
rect 6650 19510 6710 19540
rect 6650 19470 6660 19510
rect 6700 19470 6710 19510
rect 6650 19440 6710 19470
rect 6650 19400 6660 19440
rect 6700 19400 6710 19440
rect 6650 19375 6710 19400
rect 6650 19335 6660 19375
rect 6700 19335 6710 19375
rect 6650 19315 6710 19335
rect 6650 19275 6660 19315
rect 6700 19275 6710 19315
rect 6650 19250 6710 19275
rect 6650 19210 6660 19250
rect 6700 19210 6710 19250
rect 6650 19180 6710 19210
rect 6650 19140 6660 19180
rect 6700 19140 6710 19180
rect 6650 19110 6710 19140
rect 6650 19070 6660 19110
rect 6700 19070 6710 19110
rect 6650 19040 6710 19070
rect 6650 19000 6660 19040
rect 6700 19000 6710 19040
rect 6650 18975 6710 19000
rect 6650 18935 6660 18975
rect 6700 18935 6710 18975
rect 6650 18915 6710 18935
rect 6650 18875 6660 18915
rect 6700 18875 6710 18915
rect 6650 18850 6710 18875
rect 6650 18810 6660 18850
rect 6700 18810 6710 18850
rect 6650 18780 6710 18810
rect 6650 18740 6660 18780
rect 6700 18740 6710 18780
rect 6650 18710 6710 18740
rect 6650 18670 6660 18710
rect 6700 18670 6710 18710
rect 6650 18640 6710 18670
rect 6650 18600 6660 18640
rect 6700 18600 6710 18640
rect 6650 18575 6710 18600
rect 6650 18535 6660 18575
rect 6700 18535 6710 18575
rect 6650 18515 6710 18535
rect 6650 18475 6660 18515
rect 6700 18475 6710 18515
rect 6650 18450 6710 18475
rect 6650 18410 6660 18450
rect 6700 18410 6710 18450
rect 6650 18380 6710 18410
rect 6650 18340 6660 18380
rect 6700 18340 6710 18380
rect 6650 18310 6710 18340
rect 6650 18270 6660 18310
rect 6700 18270 6710 18310
rect 6650 18240 6710 18270
rect 6650 18200 6660 18240
rect 6700 18200 6710 18240
rect 6650 18175 6710 18200
rect 6650 18135 6660 18175
rect 6700 18135 6710 18175
rect 6650 18115 6710 18135
rect 6650 18075 6660 18115
rect 6700 18075 6710 18115
rect 6650 18050 6710 18075
rect 6650 18010 6660 18050
rect 6700 18010 6710 18050
rect 6650 17980 6710 18010
rect 6650 17940 6660 17980
rect 6700 17940 6710 17980
rect 6650 17910 6710 17940
rect 6650 17870 6660 17910
rect 6700 17870 6710 17910
rect 6650 17840 6710 17870
rect 6650 17800 6660 17840
rect 6700 17800 6710 17840
rect 6650 17775 6710 17800
rect 6650 17735 6660 17775
rect 6700 17735 6710 17775
rect 6650 17725 6710 17735
rect 12890 20890 16090 20925
rect 12890 20840 12925 20890
rect 12975 20840 13020 20890
rect 13070 20840 13115 20890
rect 13165 20840 13215 20890
rect 13265 20840 13315 20890
rect 13365 20840 13415 20890
rect 13465 20840 13510 20890
rect 13560 20840 13605 20890
rect 13655 20840 13725 20890
rect 13775 20840 13820 20890
rect 13870 20840 13915 20890
rect 13965 20840 14015 20890
rect 14065 20840 14115 20890
rect 14165 20840 14215 20890
rect 14265 20840 14310 20890
rect 14360 20840 14405 20890
rect 14455 20840 14525 20890
rect 14575 20840 14620 20890
rect 14670 20840 14715 20890
rect 14765 20840 14815 20890
rect 14865 20840 14915 20890
rect 14965 20840 15015 20890
rect 15065 20840 15110 20890
rect 15160 20840 15205 20890
rect 15255 20840 15325 20890
rect 15375 20840 15420 20890
rect 15470 20840 15515 20890
rect 15565 20840 15615 20890
rect 15665 20840 15715 20890
rect 15765 20840 15815 20890
rect 15865 20840 15910 20890
rect 15960 20840 16005 20890
rect 16055 20840 16090 20890
rect 12890 20800 16090 20840
rect 12890 20750 12925 20800
rect 12975 20750 13020 20800
rect 13070 20750 13115 20800
rect 13165 20750 13215 20800
rect 13265 20750 13315 20800
rect 13365 20750 13415 20800
rect 13465 20750 13510 20800
rect 13560 20750 13605 20800
rect 13655 20750 13725 20800
rect 13775 20750 13820 20800
rect 13870 20750 13915 20800
rect 13965 20750 14015 20800
rect 14065 20750 14115 20800
rect 14165 20750 14215 20800
rect 14265 20750 14310 20800
rect 14360 20750 14405 20800
rect 14455 20750 14525 20800
rect 14575 20750 14620 20800
rect 14670 20750 14715 20800
rect 14765 20750 14815 20800
rect 14865 20750 14915 20800
rect 14965 20750 15015 20800
rect 15065 20750 15110 20800
rect 15160 20750 15205 20800
rect 15255 20750 15325 20800
rect 15375 20750 15420 20800
rect 15470 20750 15515 20800
rect 15565 20750 15615 20800
rect 15665 20750 15715 20800
rect 15765 20750 15815 20800
rect 15865 20750 15910 20800
rect 15960 20750 16005 20800
rect 16055 20750 16090 20800
rect 12890 20700 16090 20750
rect 12890 20650 12925 20700
rect 12975 20650 13020 20700
rect 13070 20650 13115 20700
rect 13165 20650 13215 20700
rect 13265 20650 13315 20700
rect 13365 20650 13415 20700
rect 13465 20650 13510 20700
rect 13560 20650 13605 20700
rect 13655 20650 13725 20700
rect 13775 20650 13820 20700
rect 13870 20650 13915 20700
rect 13965 20650 14015 20700
rect 14065 20650 14115 20700
rect 14165 20650 14215 20700
rect 14265 20650 14310 20700
rect 14360 20650 14405 20700
rect 14455 20650 14525 20700
rect 14575 20650 14620 20700
rect 14670 20650 14715 20700
rect 14765 20650 14815 20700
rect 14865 20650 14915 20700
rect 14965 20650 15015 20700
rect 15065 20650 15110 20700
rect 15160 20650 15205 20700
rect 15255 20650 15325 20700
rect 15375 20650 15420 20700
rect 15470 20650 15515 20700
rect 15565 20650 15615 20700
rect 15665 20650 15715 20700
rect 15765 20650 15815 20700
rect 15865 20650 15910 20700
rect 15960 20650 16005 20700
rect 16055 20650 16090 20700
rect 12890 20610 16090 20650
rect 12890 20560 12925 20610
rect 12975 20560 13020 20610
rect 13070 20560 13115 20610
rect 13165 20560 13215 20610
rect 13265 20560 13315 20610
rect 13365 20560 13415 20610
rect 13465 20560 13510 20610
rect 13560 20560 13605 20610
rect 13655 20560 13725 20610
rect 13775 20560 13820 20610
rect 13870 20560 13915 20610
rect 13965 20560 14015 20610
rect 14065 20560 14115 20610
rect 14165 20560 14215 20610
rect 14265 20560 14310 20610
rect 14360 20560 14405 20610
rect 14455 20560 14525 20610
rect 14575 20560 14620 20610
rect 14670 20560 14715 20610
rect 14765 20560 14815 20610
rect 14865 20560 14915 20610
rect 14965 20560 15015 20610
rect 15065 20560 15110 20610
rect 15160 20560 15205 20610
rect 15255 20560 15325 20610
rect 15375 20560 15420 20610
rect 15470 20560 15515 20610
rect 15565 20560 15615 20610
rect 15665 20560 15715 20610
rect 15765 20560 15815 20610
rect 15865 20560 15910 20610
rect 15960 20560 16005 20610
rect 16055 20560 16090 20610
rect 12890 20490 16090 20560
rect 12890 20440 12925 20490
rect 12975 20440 13020 20490
rect 13070 20440 13115 20490
rect 13165 20440 13215 20490
rect 13265 20440 13315 20490
rect 13365 20440 13415 20490
rect 13465 20440 13510 20490
rect 13560 20440 13605 20490
rect 13655 20440 13725 20490
rect 13775 20440 13820 20490
rect 13870 20440 13915 20490
rect 13965 20440 14015 20490
rect 14065 20440 14115 20490
rect 14165 20440 14215 20490
rect 14265 20440 14310 20490
rect 14360 20440 14405 20490
rect 14455 20440 14525 20490
rect 14575 20440 14620 20490
rect 14670 20440 14715 20490
rect 14765 20440 14815 20490
rect 14865 20440 14915 20490
rect 14965 20440 15015 20490
rect 15065 20440 15110 20490
rect 15160 20440 15205 20490
rect 15255 20440 15325 20490
rect 15375 20440 15420 20490
rect 15470 20440 15515 20490
rect 15565 20440 15615 20490
rect 15665 20440 15715 20490
rect 15765 20440 15815 20490
rect 15865 20440 15910 20490
rect 15960 20440 16005 20490
rect 16055 20440 16090 20490
rect 12890 20400 16090 20440
rect 12890 20350 12925 20400
rect 12975 20350 13020 20400
rect 13070 20350 13115 20400
rect 13165 20350 13215 20400
rect 13265 20350 13315 20400
rect 13365 20350 13415 20400
rect 13465 20350 13510 20400
rect 13560 20350 13605 20400
rect 13655 20350 13725 20400
rect 13775 20350 13820 20400
rect 13870 20350 13915 20400
rect 13965 20350 14015 20400
rect 14065 20350 14115 20400
rect 14165 20350 14215 20400
rect 14265 20350 14310 20400
rect 14360 20350 14405 20400
rect 14455 20350 14525 20400
rect 14575 20350 14620 20400
rect 14670 20350 14715 20400
rect 14765 20350 14815 20400
rect 14865 20350 14915 20400
rect 14965 20350 15015 20400
rect 15065 20350 15110 20400
rect 15160 20350 15205 20400
rect 15255 20350 15325 20400
rect 15375 20350 15420 20400
rect 15470 20350 15515 20400
rect 15565 20350 15615 20400
rect 15665 20350 15715 20400
rect 15765 20350 15815 20400
rect 15865 20350 15910 20400
rect 15960 20350 16005 20400
rect 16055 20350 16090 20400
rect 12890 20300 16090 20350
rect 12890 20250 12925 20300
rect 12975 20250 13020 20300
rect 13070 20250 13115 20300
rect 13165 20250 13215 20300
rect 13265 20250 13315 20300
rect 13365 20250 13415 20300
rect 13465 20250 13510 20300
rect 13560 20250 13605 20300
rect 13655 20250 13725 20300
rect 13775 20250 13820 20300
rect 13870 20250 13915 20300
rect 13965 20250 14015 20300
rect 14065 20250 14115 20300
rect 14165 20250 14215 20300
rect 14265 20250 14310 20300
rect 14360 20250 14405 20300
rect 14455 20250 14525 20300
rect 14575 20250 14620 20300
rect 14670 20250 14715 20300
rect 14765 20250 14815 20300
rect 14865 20250 14915 20300
rect 14965 20250 15015 20300
rect 15065 20250 15110 20300
rect 15160 20250 15205 20300
rect 15255 20250 15325 20300
rect 15375 20250 15420 20300
rect 15470 20250 15515 20300
rect 15565 20250 15615 20300
rect 15665 20250 15715 20300
rect 15765 20250 15815 20300
rect 15865 20250 15910 20300
rect 15960 20250 16005 20300
rect 16055 20250 16090 20300
rect 12890 20210 16090 20250
rect 12890 20160 12925 20210
rect 12975 20160 13020 20210
rect 13070 20160 13115 20210
rect 13165 20160 13215 20210
rect 13265 20160 13315 20210
rect 13365 20160 13415 20210
rect 13465 20160 13510 20210
rect 13560 20160 13605 20210
rect 13655 20160 13725 20210
rect 13775 20160 13820 20210
rect 13870 20160 13915 20210
rect 13965 20160 14015 20210
rect 14065 20160 14115 20210
rect 14165 20160 14215 20210
rect 14265 20160 14310 20210
rect 14360 20160 14405 20210
rect 14455 20160 14525 20210
rect 14575 20160 14620 20210
rect 14670 20160 14715 20210
rect 14765 20160 14815 20210
rect 14865 20160 14915 20210
rect 14965 20160 15015 20210
rect 15065 20160 15110 20210
rect 15160 20160 15205 20210
rect 15255 20160 15325 20210
rect 15375 20160 15420 20210
rect 15470 20160 15515 20210
rect 15565 20160 15615 20210
rect 15665 20160 15715 20210
rect 15765 20160 15815 20210
rect 15865 20160 15910 20210
rect 15960 20160 16005 20210
rect 16055 20160 16090 20210
rect 12890 20090 16090 20160
rect 12890 20040 12925 20090
rect 12975 20040 13020 20090
rect 13070 20040 13115 20090
rect 13165 20040 13215 20090
rect 13265 20040 13315 20090
rect 13365 20040 13415 20090
rect 13465 20040 13510 20090
rect 13560 20040 13605 20090
rect 13655 20040 13725 20090
rect 13775 20040 13820 20090
rect 13870 20040 13915 20090
rect 13965 20040 14015 20090
rect 14065 20040 14115 20090
rect 14165 20040 14215 20090
rect 14265 20040 14310 20090
rect 14360 20040 14405 20090
rect 14455 20040 14525 20090
rect 14575 20040 14620 20090
rect 14670 20040 14715 20090
rect 14765 20040 14815 20090
rect 14865 20040 14915 20090
rect 14965 20040 15015 20090
rect 15065 20040 15110 20090
rect 15160 20040 15205 20090
rect 15255 20040 15325 20090
rect 15375 20040 15420 20090
rect 15470 20040 15515 20090
rect 15565 20040 15615 20090
rect 15665 20040 15715 20090
rect 15765 20040 15815 20090
rect 15865 20040 15910 20090
rect 15960 20040 16005 20090
rect 16055 20040 16090 20090
rect 12890 20000 16090 20040
rect 12890 19950 12925 20000
rect 12975 19950 13020 20000
rect 13070 19950 13115 20000
rect 13165 19950 13215 20000
rect 13265 19950 13315 20000
rect 13365 19950 13415 20000
rect 13465 19950 13510 20000
rect 13560 19950 13605 20000
rect 13655 19950 13725 20000
rect 13775 19950 13820 20000
rect 13870 19950 13915 20000
rect 13965 19950 14015 20000
rect 14065 19950 14115 20000
rect 14165 19950 14215 20000
rect 14265 19950 14310 20000
rect 14360 19950 14405 20000
rect 14455 19950 14525 20000
rect 14575 19950 14620 20000
rect 14670 19950 14715 20000
rect 14765 19950 14815 20000
rect 14865 19950 14915 20000
rect 14965 19950 15015 20000
rect 15065 19950 15110 20000
rect 15160 19950 15205 20000
rect 15255 19950 15325 20000
rect 15375 19950 15420 20000
rect 15470 19950 15515 20000
rect 15565 19950 15615 20000
rect 15665 19950 15715 20000
rect 15765 19950 15815 20000
rect 15865 19950 15910 20000
rect 15960 19950 16005 20000
rect 16055 19950 16090 20000
rect 12890 19900 16090 19950
rect 12890 19850 12925 19900
rect 12975 19850 13020 19900
rect 13070 19850 13115 19900
rect 13165 19850 13215 19900
rect 13265 19850 13315 19900
rect 13365 19850 13415 19900
rect 13465 19850 13510 19900
rect 13560 19850 13605 19900
rect 13655 19850 13725 19900
rect 13775 19850 13820 19900
rect 13870 19850 13915 19900
rect 13965 19850 14015 19900
rect 14065 19850 14115 19900
rect 14165 19850 14215 19900
rect 14265 19850 14310 19900
rect 14360 19850 14405 19900
rect 14455 19850 14525 19900
rect 14575 19850 14620 19900
rect 14670 19850 14715 19900
rect 14765 19850 14815 19900
rect 14865 19850 14915 19900
rect 14965 19850 15015 19900
rect 15065 19850 15110 19900
rect 15160 19850 15205 19900
rect 15255 19850 15325 19900
rect 15375 19850 15420 19900
rect 15470 19850 15515 19900
rect 15565 19850 15615 19900
rect 15665 19850 15715 19900
rect 15765 19850 15815 19900
rect 15865 19850 15910 19900
rect 15960 19850 16005 19900
rect 16055 19850 16090 19900
rect 12890 19810 16090 19850
rect 12890 19760 12925 19810
rect 12975 19760 13020 19810
rect 13070 19760 13115 19810
rect 13165 19760 13215 19810
rect 13265 19760 13315 19810
rect 13365 19760 13415 19810
rect 13465 19760 13510 19810
rect 13560 19760 13605 19810
rect 13655 19760 13725 19810
rect 13775 19760 13820 19810
rect 13870 19760 13915 19810
rect 13965 19760 14015 19810
rect 14065 19760 14115 19810
rect 14165 19760 14215 19810
rect 14265 19760 14310 19810
rect 14360 19760 14405 19810
rect 14455 19760 14525 19810
rect 14575 19760 14620 19810
rect 14670 19760 14715 19810
rect 14765 19760 14815 19810
rect 14865 19760 14915 19810
rect 14965 19760 15015 19810
rect 15065 19760 15110 19810
rect 15160 19760 15205 19810
rect 15255 19760 15325 19810
rect 15375 19760 15420 19810
rect 15470 19760 15515 19810
rect 15565 19760 15615 19810
rect 15665 19760 15715 19810
rect 15765 19760 15815 19810
rect 15865 19760 15910 19810
rect 15960 19760 16005 19810
rect 16055 19760 16090 19810
rect 12890 19690 16090 19760
rect 12890 19640 12925 19690
rect 12975 19640 13020 19690
rect 13070 19640 13115 19690
rect 13165 19640 13215 19690
rect 13265 19640 13315 19690
rect 13365 19640 13415 19690
rect 13465 19640 13510 19690
rect 13560 19640 13605 19690
rect 13655 19640 13725 19690
rect 13775 19640 13820 19690
rect 13870 19640 13915 19690
rect 13965 19640 14015 19690
rect 14065 19640 14115 19690
rect 14165 19640 14215 19690
rect 14265 19640 14310 19690
rect 14360 19640 14405 19690
rect 14455 19640 14525 19690
rect 14575 19640 14620 19690
rect 14670 19640 14715 19690
rect 14765 19640 14815 19690
rect 14865 19640 14915 19690
rect 14965 19640 15015 19690
rect 15065 19640 15110 19690
rect 15160 19640 15205 19690
rect 15255 19640 15325 19690
rect 15375 19640 15420 19690
rect 15470 19640 15515 19690
rect 15565 19640 15615 19690
rect 15665 19640 15715 19690
rect 15765 19640 15815 19690
rect 15865 19640 15910 19690
rect 15960 19640 16005 19690
rect 16055 19640 16090 19690
rect 12890 19600 16090 19640
rect 12890 19550 12925 19600
rect 12975 19550 13020 19600
rect 13070 19550 13115 19600
rect 13165 19550 13215 19600
rect 13265 19550 13315 19600
rect 13365 19550 13415 19600
rect 13465 19550 13510 19600
rect 13560 19550 13605 19600
rect 13655 19550 13725 19600
rect 13775 19550 13820 19600
rect 13870 19550 13915 19600
rect 13965 19550 14015 19600
rect 14065 19550 14115 19600
rect 14165 19550 14215 19600
rect 14265 19550 14310 19600
rect 14360 19550 14405 19600
rect 14455 19550 14525 19600
rect 14575 19550 14620 19600
rect 14670 19550 14715 19600
rect 14765 19550 14815 19600
rect 14865 19550 14915 19600
rect 14965 19550 15015 19600
rect 15065 19550 15110 19600
rect 15160 19550 15205 19600
rect 15255 19550 15325 19600
rect 15375 19550 15420 19600
rect 15470 19550 15515 19600
rect 15565 19550 15615 19600
rect 15665 19550 15715 19600
rect 15765 19550 15815 19600
rect 15865 19550 15910 19600
rect 15960 19550 16005 19600
rect 16055 19550 16090 19600
rect 12890 19500 16090 19550
rect 12890 19450 12925 19500
rect 12975 19450 13020 19500
rect 13070 19450 13115 19500
rect 13165 19450 13215 19500
rect 13265 19450 13315 19500
rect 13365 19450 13415 19500
rect 13465 19450 13510 19500
rect 13560 19450 13605 19500
rect 13655 19450 13725 19500
rect 13775 19450 13820 19500
rect 13870 19450 13915 19500
rect 13965 19450 14015 19500
rect 14065 19450 14115 19500
rect 14165 19450 14215 19500
rect 14265 19450 14310 19500
rect 14360 19450 14405 19500
rect 14455 19450 14525 19500
rect 14575 19450 14620 19500
rect 14670 19450 14715 19500
rect 14765 19450 14815 19500
rect 14865 19450 14915 19500
rect 14965 19450 15015 19500
rect 15065 19450 15110 19500
rect 15160 19450 15205 19500
rect 15255 19450 15325 19500
rect 15375 19450 15420 19500
rect 15470 19450 15515 19500
rect 15565 19450 15615 19500
rect 15665 19450 15715 19500
rect 15765 19450 15815 19500
rect 15865 19450 15910 19500
rect 15960 19450 16005 19500
rect 16055 19450 16090 19500
rect 12890 19410 16090 19450
rect 12890 19360 12925 19410
rect 12975 19360 13020 19410
rect 13070 19360 13115 19410
rect 13165 19360 13215 19410
rect 13265 19360 13315 19410
rect 13365 19360 13415 19410
rect 13465 19360 13510 19410
rect 13560 19360 13605 19410
rect 13655 19360 13725 19410
rect 13775 19360 13820 19410
rect 13870 19360 13915 19410
rect 13965 19360 14015 19410
rect 14065 19360 14115 19410
rect 14165 19360 14215 19410
rect 14265 19360 14310 19410
rect 14360 19360 14405 19410
rect 14455 19360 14525 19410
rect 14575 19360 14620 19410
rect 14670 19360 14715 19410
rect 14765 19360 14815 19410
rect 14865 19360 14915 19410
rect 14965 19360 15015 19410
rect 15065 19360 15110 19410
rect 15160 19360 15205 19410
rect 15255 19360 15325 19410
rect 15375 19360 15420 19410
rect 15470 19360 15515 19410
rect 15565 19360 15615 19410
rect 15665 19360 15715 19410
rect 15765 19360 15815 19410
rect 15865 19360 15910 19410
rect 15960 19360 16005 19410
rect 16055 19360 16090 19410
rect 12890 19290 16090 19360
rect 12890 19240 12925 19290
rect 12975 19240 13020 19290
rect 13070 19240 13115 19290
rect 13165 19240 13215 19290
rect 13265 19240 13315 19290
rect 13365 19240 13415 19290
rect 13465 19240 13510 19290
rect 13560 19240 13605 19290
rect 13655 19240 13725 19290
rect 13775 19240 13820 19290
rect 13870 19240 13915 19290
rect 13965 19240 14015 19290
rect 14065 19240 14115 19290
rect 14165 19240 14215 19290
rect 14265 19240 14310 19290
rect 14360 19240 14405 19290
rect 14455 19240 14525 19290
rect 14575 19240 14620 19290
rect 14670 19240 14715 19290
rect 14765 19240 14815 19290
rect 14865 19240 14915 19290
rect 14965 19240 15015 19290
rect 15065 19240 15110 19290
rect 15160 19240 15205 19290
rect 15255 19240 15325 19290
rect 15375 19240 15420 19290
rect 15470 19240 15515 19290
rect 15565 19240 15615 19290
rect 15665 19240 15715 19290
rect 15765 19240 15815 19290
rect 15865 19240 15910 19290
rect 15960 19240 16005 19290
rect 16055 19240 16090 19290
rect 12890 19200 16090 19240
rect 12890 19150 12925 19200
rect 12975 19150 13020 19200
rect 13070 19150 13115 19200
rect 13165 19150 13215 19200
rect 13265 19150 13315 19200
rect 13365 19150 13415 19200
rect 13465 19150 13510 19200
rect 13560 19150 13605 19200
rect 13655 19150 13725 19200
rect 13775 19150 13820 19200
rect 13870 19150 13915 19200
rect 13965 19150 14015 19200
rect 14065 19150 14115 19200
rect 14165 19150 14215 19200
rect 14265 19150 14310 19200
rect 14360 19150 14405 19200
rect 14455 19150 14525 19200
rect 14575 19150 14620 19200
rect 14670 19150 14715 19200
rect 14765 19150 14815 19200
rect 14865 19150 14915 19200
rect 14965 19150 15015 19200
rect 15065 19150 15110 19200
rect 15160 19150 15205 19200
rect 15255 19150 15325 19200
rect 15375 19150 15420 19200
rect 15470 19150 15515 19200
rect 15565 19150 15615 19200
rect 15665 19150 15715 19200
rect 15765 19150 15815 19200
rect 15865 19150 15910 19200
rect 15960 19150 16005 19200
rect 16055 19150 16090 19200
rect 12890 19100 16090 19150
rect 12890 19050 12925 19100
rect 12975 19050 13020 19100
rect 13070 19050 13115 19100
rect 13165 19050 13215 19100
rect 13265 19050 13315 19100
rect 13365 19050 13415 19100
rect 13465 19050 13510 19100
rect 13560 19050 13605 19100
rect 13655 19050 13725 19100
rect 13775 19050 13820 19100
rect 13870 19050 13915 19100
rect 13965 19050 14015 19100
rect 14065 19050 14115 19100
rect 14165 19050 14215 19100
rect 14265 19050 14310 19100
rect 14360 19050 14405 19100
rect 14455 19050 14525 19100
rect 14575 19050 14620 19100
rect 14670 19050 14715 19100
rect 14765 19050 14815 19100
rect 14865 19050 14915 19100
rect 14965 19050 15015 19100
rect 15065 19050 15110 19100
rect 15160 19050 15205 19100
rect 15255 19050 15325 19100
rect 15375 19050 15420 19100
rect 15470 19050 15515 19100
rect 15565 19050 15615 19100
rect 15665 19050 15715 19100
rect 15765 19050 15815 19100
rect 15865 19050 15910 19100
rect 15960 19050 16005 19100
rect 16055 19050 16090 19100
rect 12890 19010 16090 19050
rect 12890 18960 12925 19010
rect 12975 18960 13020 19010
rect 13070 18960 13115 19010
rect 13165 18960 13215 19010
rect 13265 18960 13315 19010
rect 13365 18960 13415 19010
rect 13465 18960 13510 19010
rect 13560 18960 13605 19010
rect 13655 18960 13725 19010
rect 13775 18960 13820 19010
rect 13870 18960 13915 19010
rect 13965 18960 14015 19010
rect 14065 18960 14115 19010
rect 14165 18960 14215 19010
rect 14265 18960 14310 19010
rect 14360 18960 14405 19010
rect 14455 18960 14525 19010
rect 14575 18960 14620 19010
rect 14670 18960 14715 19010
rect 14765 18960 14815 19010
rect 14865 18960 14915 19010
rect 14965 18960 15015 19010
rect 15065 18960 15110 19010
rect 15160 18960 15205 19010
rect 15255 18960 15325 19010
rect 15375 18960 15420 19010
rect 15470 18960 15515 19010
rect 15565 18960 15615 19010
rect 15665 18960 15715 19010
rect 15765 18960 15815 19010
rect 15865 18960 15910 19010
rect 15960 18960 16005 19010
rect 16055 18960 16090 19010
rect 12890 18890 16090 18960
rect 12890 18840 12925 18890
rect 12975 18840 13020 18890
rect 13070 18840 13115 18890
rect 13165 18840 13215 18890
rect 13265 18840 13315 18890
rect 13365 18840 13415 18890
rect 13465 18840 13510 18890
rect 13560 18840 13605 18890
rect 13655 18840 13725 18890
rect 13775 18840 13820 18890
rect 13870 18840 13915 18890
rect 13965 18840 14015 18890
rect 14065 18840 14115 18890
rect 14165 18840 14215 18890
rect 14265 18840 14310 18890
rect 14360 18840 14405 18890
rect 14455 18840 14525 18890
rect 14575 18840 14620 18890
rect 14670 18840 14715 18890
rect 14765 18840 14815 18890
rect 14865 18840 14915 18890
rect 14965 18840 15015 18890
rect 15065 18840 15110 18890
rect 15160 18840 15205 18890
rect 15255 18840 15325 18890
rect 15375 18840 15420 18890
rect 15470 18840 15515 18890
rect 15565 18840 15615 18890
rect 15665 18840 15715 18890
rect 15765 18840 15815 18890
rect 15865 18840 15910 18890
rect 15960 18840 16005 18890
rect 16055 18840 16090 18890
rect 12890 18800 16090 18840
rect 12890 18750 12925 18800
rect 12975 18750 13020 18800
rect 13070 18750 13115 18800
rect 13165 18750 13215 18800
rect 13265 18750 13315 18800
rect 13365 18750 13415 18800
rect 13465 18750 13510 18800
rect 13560 18750 13605 18800
rect 13655 18750 13725 18800
rect 13775 18750 13820 18800
rect 13870 18750 13915 18800
rect 13965 18750 14015 18800
rect 14065 18750 14115 18800
rect 14165 18750 14215 18800
rect 14265 18750 14310 18800
rect 14360 18750 14405 18800
rect 14455 18750 14525 18800
rect 14575 18750 14620 18800
rect 14670 18750 14715 18800
rect 14765 18750 14815 18800
rect 14865 18750 14915 18800
rect 14965 18750 15015 18800
rect 15065 18750 15110 18800
rect 15160 18750 15205 18800
rect 15255 18750 15325 18800
rect 15375 18750 15420 18800
rect 15470 18750 15515 18800
rect 15565 18750 15615 18800
rect 15665 18750 15715 18800
rect 15765 18750 15815 18800
rect 15865 18750 15910 18800
rect 15960 18750 16005 18800
rect 16055 18750 16090 18800
rect 12890 18700 16090 18750
rect 12890 18650 12925 18700
rect 12975 18650 13020 18700
rect 13070 18650 13115 18700
rect 13165 18650 13215 18700
rect 13265 18650 13315 18700
rect 13365 18650 13415 18700
rect 13465 18650 13510 18700
rect 13560 18650 13605 18700
rect 13655 18650 13725 18700
rect 13775 18650 13820 18700
rect 13870 18650 13915 18700
rect 13965 18650 14015 18700
rect 14065 18650 14115 18700
rect 14165 18650 14215 18700
rect 14265 18650 14310 18700
rect 14360 18650 14405 18700
rect 14455 18650 14525 18700
rect 14575 18650 14620 18700
rect 14670 18650 14715 18700
rect 14765 18650 14815 18700
rect 14865 18650 14915 18700
rect 14965 18650 15015 18700
rect 15065 18650 15110 18700
rect 15160 18650 15205 18700
rect 15255 18650 15325 18700
rect 15375 18650 15420 18700
rect 15470 18650 15515 18700
rect 15565 18650 15615 18700
rect 15665 18650 15715 18700
rect 15765 18650 15815 18700
rect 15865 18650 15910 18700
rect 15960 18650 16005 18700
rect 16055 18650 16090 18700
rect 12890 18610 16090 18650
rect 12890 18560 12925 18610
rect 12975 18560 13020 18610
rect 13070 18560 13115 18610
rect 13165 18560 13215 18610
rect 13265 18560 13315 18610
rect 13365 18560 13415 18610
rect 13465 18560 13510 18610
rect 13560 18560 13605 18610
rect 13655 18560 13725 18610
rect 13775 18560 13820 18610
rect 13870 18560 13915 18610
rect 13965 18560 14015 18610
rect 14065 18560 14115 18610
rect 14165 18560 14215 18610
rect 14265 18560 14310 18610
rect 14360 18560 14405 18610
rect 14455 18560 14525 18610
rect 14575 18560 14620 18610
rect 14670 18560 14715 18610
rect 14765 18560 14815 18610
rect 14865 18560 14915 18610
rect 14965 18560 15015 18610
rect 15065 18560 15110 18610
rect 15160 18560 15205 18610
rect 15255 18560 15325 18610
rect 15375 18560 15420 18610
rect 15470 18560 15515 18610
rect 15565 18560 15615 18610
rect 15665 18560 15715 18610
rect 15765 18560 15815 18610
rect 15865 18560 15910 18610
rect 15960 18560 16005 18610
rect 16055 18560 16090 18610
rect 12890 18490 16090 18560
rect 12890 18440 12925 18490
rect 12975 18440 13020 18490
rect 13070 18440 13115 18490
rect 13165 18440 13215 18490
rect 13265 18440 13315 18490
rect 13365 18440 13415 18490
rect 13465 18440 13510 18490
rect 13560 18440 13605 18490
rect 13655 18440 13725 18490
rect 13775 18440 13820 18490
rect 13870 18440 13915 18490
rect 13965 18440 14015 18490
rect 14065 18440 14115 18490
rect 14165 18440 14215 18490
rect 14265 18440 14310 18490
rect 14360 18440 14405 18490
rect 14455 18440 14525 18490
rect 14575 18440 14620 18490
rect 14670 18440 14715 18490
rect 14765 18440 14815 18490
rect 14865 18440 14915 18490
rect 14965 18440 15015 18490
rect 15065 18440 15110 18490
rect 15160 18440 15205 18490
rect 15255 18440 15325 18490
rect 15375 18440 15420 18490
rect 15470 18440 15515 18490
rect 15565 18440 15615 18490
rect 15665 18440 15715 18490
rect 15765 18440 15815 18490
rect 15865 18440 15910 18490
rect 15960 18440 16005 18490
rect 16055 18440 16090 18490
rect 12890 18400 16090 18440
rect 12890 18350 12925 18400
rect 12975 18350 13020 18400
rect 13070 18350 13115 18400
rect 13165 18350 13215 18400
rect 13265 18350 13315 18400
rect 13365 18350 13415 18400
rect 13465 18350 13510 18400
rect 13560 18350 13605 18400
rect 13655 18350 13725 18400
rect 13775 18350 13820 18400
rect 13870 18350 13915 18400
rect 13965 18350 14015 18400
rect 14065 18350 14115 18400
rect 14165 18350 14215 18400
rect 14265 18350 14310 18400
rect 14360 18350 14405 18400
rect 14455 18350 14525 18400
rect 14575 18350 14620 18400
rect 14670 18350 14715 18400
rect 14765 18350 14815 18400
rect 14865 18350 14915 18400
rect 14965 18350 15015 18400
rect 15065 18350 15110 18400
rect 15160 18350 15205 18400
rect 15255 18350 15325 18400
rect 15375 18350 15420 18400
rect 15470 18350 15515 18400
rect 15565 18350 15615 18400
rect 15665 18350 15715 18400
rect 15765 18350 15815 18400
rect 15865 18350 15910 18400
rect 15960 18350 16005 18400
rect 16055 18350 16090 18400
rect 12890 18300 16090 18350
rect 12890 18250 12925 18300
rect 12975 18250 13020 18300
rect 13070 18250 13115 18300
rect 13165 18250 13215 18300
rect 13265 18250 13315 18300
rect 13365 18250 13415 18300
rect 13465 18250 13510 18300
rect 13560 18250 13605 18300
rect 13655 18250 13725 18300
rect 13775 18250 13820 18300
rect 13870 18250 13915 18300
rect 13965 18250 14015 18300
rect 14065 18250 14115 18300
rect 14165 18250 14215 18300
rect 14265 18250 14310 18300
rect 14360 18250 14405 18300
rect 14455 18250 14525 18300
rect 14575 18250 14620 18300
rect 14670 18250 14715 18300
rect 14765 18250 14815 18300
rect 14865 18250 14915 18300
rect 14965 18250 15015 18300
rect 15065 18250 15110 18300
rect 15160 18250 15205 18300
rect 15255 18250 15325 18300
rect 15375 18250 15420 18300
rect 15470 18250 15515 18300
rect 15565 18250 15615 18300
rect 15665 18250 15715 18300
rect 15765 18250 15815 18300
rect 15865 18250 15910 18300
rect 15960 18250 16005 18300
rect 16055 18250 16090 18300
rect 12890 18210 16090 18250
rect 12890 18160 12925 18210
rect 12975 18160 13020 18210
rect 13070 18160 13115 18210
rect 13165 18160 13215 18210
rect 13265 18160 13315 18210
rect 13365 18160 13415 18210
rect 13465 18160 13510 18210
rect 13560 18160 13605 18210
rect 13655 18160 13725 18210
rect 13775 18160 13820 18210
rect 13870 18160 13915 18210
rect 13965 18160 14015 18210
rect 14065 18160 14115 18210
rect 14165 18160 14215 18210
rect 14265 18160 14310 18210
rect 14360 18160 14405 18210
rect 14455 18160 14525 18210
rect 14575 18160 14620 18210
rect 14670 18160 14715 18210
rect 14765 18160 14815 18210
rect 14865 18160 14915 18210
rect 14965 18160 15015 18210
rect 15065 18160 15110 18210
rect 15160 18160 15205 18210
rect 15255 18160 15325 18210
rect 15375 18160 15420 18210
rect 15470 18160 15515 18210
rect 15565 18160 15615 18210
rect 15665 18160 15715 18210
rect 15765 18160 15815 18210
rect 15865 18160 15910 18210
rect 15960 18160 16005 18210
rect 16055 18160 16090 18210
rect 12890 18090 16090 18160
rect 12890 18040 12925 18090
rect 12975 18040 13020 18090
rect 13070 18040 13115 18090
rect 13165 18040 13215 18090
rect 13265 18040 13315 18090
rect 13365 18040 13415 18090
rect 13465 18040 13510 18090
rect 13560 18040 13605 18090
rect 13655 18040 13725 18090
rect 13775 18040 13820 18090
rect 13870 18040 13915 18090
rect 13965 18040 14015 18090
rect 14065 18040 14115 18090
rect 14165 18040 14215 18090
rect 14265 18040 14310 18090
rect 14360 18040 14405 18090
rect 14455 18040 14525 18090
rect 14575 18040 14620 18090
rect 14670 18040 14715 18090
rect 14765 18040 14815 18090
rect 14865 18040 14915 18090
rect 14965 18040 15015 18090
rect 15065 18040 15110 18090
rect 15160 18040 15205 18090
rect 15255 18040 15325 18090
rect 15375 18040 15420 18090
rect 15470 18040 15515 18090
rect 15565 18040 15615 18090
rect 15665 18040 15715 18090
rect 15765 18040 15815 18090
rect 15865 18040 15910 18090
rect 15960 18040 16005 18090
rect 16055 18040 16090 18090
rect 12890 18000 16090 18040
rect 12890 17950 12925 18000
rect 12975 17950 13020 18000
rect 13070 17950 13115 18000
rect 13165 17950 13215 18000
rect 13265 17950 13315 18000
rect 13365 17950 13415 18000
rect 13465 17950 13510 18000
rect 13560 17950 13605 18000
rect 13655 17950 13725 18000
rect 13775 17950 13820 18000
rect 13870 17950 13915 18000
rect 13965 17950 14015 18000
rect 14065 17950 14115 18000
rect 14165 17950 14215 18000
rect 14265 17950 14310 18000
rect 14360 17950 14405 18000
rect 14455 17950 14525 18000
rect 14575 17950 14620 18000
rect 14670 17950 14715 18000
rect 14765 17950 14815 18000
rect 14865 17950 14915 18000
rect 14965 17950 15015 18000
rect 15065 17950 15110 18000
rect 15160 17950 15205 18000
rect 15255 17950 15325 18000
rect 15375 17950 15420 18000
rect 15470 17950 15515 18000
rect 15565 17950 15615 18000
rect 15665 17950 15715 18000
rect 15765 17950 15815 18000
rect 15865 17950 15910 18000
rect 15960 17950 16005 18000
rect 16055 17950 16090 18000
rect 12890 17900 16090 17950
rect 12890 17850 12925 17900
rect 12975 17850 13020 17900
rect 13070 17850 13115 17900
rect 13165 17850 13215 17900
rect 13265 17850 13315 17900
rect 13365 17850 13415 17900
rect 13465 17850 13510 17900
rect 13560 17850 13605 17900
rect 13655 17850 13725 17900
rect 13775 17850 13820 17900
rect 13870 17850 13915 17900
rect 13965 17850 14015 17900
rect 14065 17850 14115 17900
rect 14165 17850 14215 17900
rect 14265 17850 14310 17900
rect 14360 17850 14405 17900
rect 14455 17850 14525 17900
rect 14575 17850 14620 17900
rect 14670 17850 14715 17900
rect 14765 17850 14815 17900
rect 14865 17850 14915 17900
rect 14965 17850 15015 17900
rect 15065 17850 15110 17900
rect 15160 17850 15205 17900
rect 15255 17850 15325 17900
rect 15375 17850 15420 17900
rect 15470 17850 15515 17900
rect 15565 17850 15615 17900
rect 15665 17850 15715 17900
rect 15765 17850 15815 17900
rect 15865 17850 15910 17900
rect 15960 17850 16005 17900
rect 16055 17850 16090 17900
rect 12890 17810 16090 17850
rect 12890 17760 12925 17810
rect 12975 17760 13020 17810
rect 13070 17760 13115 17810
rect 13165 17760 13215 17810
rect 13265 17760 13315 17810
rect 13365 17760 13415 17810
rect 13465 17760 13510 17810
rect 13560 17760 13605 17810
rect 13655 17760 13725 17810
rect 13775 17760 13820 17810
rect 13870 17760 13915 17810
rect 13965 17760 14015 17810
rect 14065 17760 14115 17810
rect 14165 17760 14215 17810
rect 14265 17760 14310 17810
rect 14360 17760 14405 17810
rect 14455 17760 14525 17810
rect 14575 17760 14620 17810
rect 14670 17760 14715 17810
rect 14765 17760 14815 17810
rect 14865 17760 14915 17810
rect 14965 17760 15015 17810
rect 15065 17760 15110 17810
rect 15160 17760 15205 17810
rect 15255 17760 15325 17810
rect 15375 17760 15420 17810
rect 15470 17760 15515 17810
rect 15565 17760 15615 17810
rect 15665 17760 15715 17810
rect 15765 17760 15815 17810
rect 15865 17760 15910 17810
rect 15960 17760 16005 17810
rect 16055 17760 16090 17810
rect -4840 9615 -1640 10155
rect -4840 9565 -4805 9615
rect -4755 9565 -4710 9615
rect -4660 9565 -4615 9615
rect -4565 9565 -4515 9615
rect -4465 9565 -4415 9615
rect -4365 9565 -4315 9615
rect -4265 9565 -4220 9615
rect -4170 9565 -4125 9615
rect -4075 9565 -4005 9615
rect -3955 9565 -3910 9615
rect -3860 9565 -3815 9615
rect -3765 9565 -3715 9615
rect -3665 9565 -3615 9615
rect -3565 9565 -3515 9615
rect -3465 9565 -3420 9615
rect -3370 9565 -3325 9615
rect -3275 9565 -3205 9615
rect -3155 9565 -3110 9615
rect -3060 9565 -3015 9615
rect -2965 9565 -2915 9615
rect -2865 9565 -2815 9615
rect -2765 9565 -2715 9615
rect -2665 9565 -2620 9615
rect -2570 9565 -2525 9615
rect -2475 9565 -2405 9615
rect -2355 9565 -2310 9615
rect -2260 9565 -2215 9615
rect -2165 9565 -2115 9615
rect -2065 9565 -2015 9615
rect -1965 9565 -1915 9615
rect -1865 9565 -1820 9615
rect -1770 9565 -1725 9615
rect -1675 9565 -1640 9615
rect -4840 9525 -1640 9565
rect -4840 9475 -4805 9525
rect -4755 9475 -4710 9525
rect -4660 9475 -4615 9525
rect -4565 9475 -4515 9525
rect -4465 9475 -4415 9525
rect -4365 9475 -4315 9525
rect -4265 9475 -4220 9525
rect -4170 9475 -4125 9525
rect -4075 9475 -4005 9525
rect -3955 9475 -3910 9525
rect -3860 9475 -3815 9525
rect -3765 9475 -3715 9525
rect -3665 9475 -3615 9525
rect -3565 9475 -3515 9525
rect -3465 9475 -3420 9525
rect -3370 9475 -3325 9525
rect -3275 9475 -3205 9525
rect -3155 9475 -3110 9525
rect -3060 9475 -3015 9525
rect -2965 9475 -2915 9525
rect -2865 9475 -2815 9525
rect -2765 9475 -2715 9525
rect -2665 9475 -2620 9525
rect -2570 9475 -2525 9525
rect -2475 9475 -2405 9525
rect -2355 9475 -2310 9525
rect -2260 9475 -2215 9525
rect -2165 9475 -2115 9525
rect -2065 9475 -2015 9525
rect -1965 9475 -1915 9525
rect -1865 9475 -1820 9525
rect -1770 9475 -1725 9525
rect -1675 9475 -1640 9525
rect -4840 9425 -1640 9475
rect -4840 9375 -4805 9425
rect -4755 9375 -4710 9425
rect -4660 9375 -4615 9425
rect -4565 9375 -4515 9425
rect -4465 9375 -4415 9425
rect -4365 9375 -4315 9425
rect -4265 9375 -4220 9425
rect -4170 9375 -4125 9425
rect -4075 9375 -4005 9425
rect -3955 9375 -3910 9425
rect -3860 9375 -3815 9425
rect -3765 9375 -3715 9425
rect -3665 9375 -3615 9425
rect -3565 9375 -3515 9425
rect -3465 9375 -3420 9425
rect -3370 9375 -3325 9425
rect -3275 9375 -3205 9425
rect -3155 9375 -3110 9425
rect -3060 9375 -3015 9425
rect -2965 9375 -2915 9425
rect -2865 9375 -2815 9425
rect -2765 9375 -2715 9425
rect -2665 9375 -2620 9425
rect -2570 9375 -2525 9425
rect -2475 9375 -2405 9425
rect -2355 9375 -2310 9425
rect -2260 9375 -2215 9425
rect -2165 9375 -2115 9425
rect -2065 9375 -2015 9425
rect -1965 9375 -1915 9425
rect -1865 9375 -1820 9425
rect -1770 9375 -1725 9425
rect -1675 9375 -1640 9425
rect -4840 9335 -1640 9375
rect -4840 9285 -4805 9335
rect -4755 9285 -4710 9335
rect -4660 9285 -4615 9335
rect -4565 9285 -4515 9335
rect -4465 9285 -4415 9335
rect -4365 9285 -4315 9335
rect -4265 9285 -4220 9335
rect -4170 9285 -4125 9335
rect -4075 9285 -4005 9335
rect -3955 9285 -3910 9335
rect -3860 9285 -3815 9335
rect -3765 9285 -3715 9335
rect -3665 9285 -3615 9335
rect -3565 9285 -3515 9335
rect -3465 9285 -3420 9335
rect -3370 9285 -3325 9335
rect -3275 9285 -3205 9335
rect -3155 9285 -3110 9335
rect -3060 9285 -3015 9335
rect -2965 9285 -2915 9335
rect -2865 9285 -2815 9335
rect -2765 9285 -2715 9335
rect -2665 9285 -2620 9335
rect -2570 9285 -2525 9335
rect -2475 9285 -2405 9335
rect -2355 9285 -2310 9335
rect -2260 9285 -2215 9335
rect -2165 9285 -2115 9335
rect -2065 9285 -2015 9335
rect -1965 9285 -1915 9335
rect -1865 9285 -1820 9335
rect -1770 9285 -1725 9335
rect -1675 9285 -1640 9335
rect -4840 9215 -1640 9285
rect -4840 9165 -4805 9215
rect -4755 9165 -4710 9215
rect -4660 9165 -4615 9215
rect -4565 9165 -4515 9215
rect -4465 9165 -4415 9215
rect -4365 9165 -4315 9215
rect -4265 9165 -4220 9215
rect -4170 9165 -4125 9215
rect -4075 9165 -4005 9215
rect -3955 9165 -3910 9215
rect -3860 9165 -3815 9215
rect -3765 9165 -3715 9215
rect -3665 9165 -3615 9215
rect -3565 9165 -3515 9215
rect -3465 9165 -3420 9215
rect -3370 9165 -3325 9215
rect -3275 9165 -3205 9215
rect -3155 9165 -3110 9215
rect -3060 9165 -3015 9215
rect -2965 9165 -2915 9215
rect -2865 9165 -2815 9215
rect -2765 9165 -2715 9215
rect -2665 9165 -2620 9215
rect -2570 9165 -2525 9215
rect -2475 9165 -2405 9215
rect -2355 9165 -2310 9215
rect -2260 9165 -2215 9215
rect -2165 9165 -2115 9215
rect -2065 9165 -2015 9215
rect -1965 9165 -1915 9215
rect -1865 9165 -1820 9215
rect -1770 9165 -1725 9215
rect -1675 9165 -1640 9215
rect -4840 9125 -1640 9165
rect -4840 9075 -4805 9125
rect -4755 9075 -4710 9125
rect -4660 9075 -4615 9125
rect -4565 9075 -4515 9125
rect -4465 9075 -4415 9125
rect -4365 9075 -4315 9125
rect -4265 9075 -4220 9125
rect -4170 9075 -4125 9125
rect -4075 9075 -4005 9125
rect -3955 9075 -3910 9125
rect -3860 9075 -3815 9125
rect -3765 9075 -3715 9125
rect -3665 9075 -3615 9125
rect -3565 9075 -3515 9125
rect -3465 9075 -3420 9125
rect -3370 9075 -3325 9125
rect -3275 9075 -3205 9125
rect -3155 9075 -3110 9125
rect -3060 9075 -3015 9125
rect -2965 9075 -2915 9125
rect -2865 9075 -2815 9125
rect -2765 9075 -2715 9125
rect -2665 9075 -2620 9125
rect -2570 9075 -2525 9125
rect -2475 9075 -2405 9125
rect -2355 9075 -2310 9125
rect -2260 9075 -2215 9125
rect -2165 9075 -2115 9125
rect -2065 9075 -2015 9125
rect -1965 9075 -1915 9125
rect -1865 9075 -1820 9125
rect -1770 9075 -1725 9125
rect -1675 9075 -1640 9125
rect -4840 9025 -1640 9075
rect -4840 8975 -4805 9025
rect -4755 8975 -4710 9025
rect -4660 8975 -4615 9025
rect -4565 8975 -4515 9025
rect -4465 8975 -4415 9025
rect -4365 8975 -4315 9025
rect -4265 8975 -4220 9025
rect -4170 8975 -4125 9025
rect -4075 8975 -4005 9025
rect -3955 8975 -3910 9025
rect -3860 8975 -3815 9025
rect -3765 8975 -3715 9025
rect -3665 8975 -3615 9025
rect -3565 8975 -3515 9025
rect -3465 8975 -3420 9025
rect -3370 8975 -3325 9025
rect -3275 8975 -3205 9025
rect -3155 8975 -3110 9025
rect -3060 8975 -3015 9025
rect -2965 8975 -2915 9025
rect -2865 8975 -2815 9025
rect -2765 8975 -2715 9025
rect -2665 8975 -2620 9025
rect -2570 8975 -2525 9025
rect -2475 8975 -2405 9025
rect -2355 8975 -2310 9025
rect -2260 8975 -2215 9025
rect -2165 8975 -2115 9025
rect -2065 8975 -2015 9025
rect -1965 8975 -1915 9025
rect -1865 8975 -1820 9025
rect -1770 8975 -1725 9025
rect -1675 8975 -1640 9025
rect -4840 8935 -1640 8975
rect -4840 8885 -4805 8935
rect -4755 8885 -4710 8935
rect -4660 8885 -4615 8935
rect -4565 8885 -4515 8935
rect -4465 8885 -4415 8935
rect -4365 8885 -4315 8935
rect -4265 8885 -4220 8935
rect -4170 8885 -4125 8935
rect -4075 8885 -4005 8935
rect -3955 8885 -3910 8935
rect -3860 8885 -3815 8935
rect -3765 8885 -3715 8935
rect -3665 8885 -3615 8935
rect -3565 8885 -3515 8935
rect -3465 8885 -3420 8935
rect -3370 8885 -3325 8935
rect -3275 8885 -3205 8935
rect -3155 8885 -3110 8935
rect -3060 8885 -3015 8935
rect -2965 8885 -2915 8935
rect -2865 8885 -2815 8935
rect -2765 8885 -2715 8935
rect -2665 8885 -2620 8935
rect -2570 8885 -2525 8935
rect -2475 8885 -2405 8935
rect -2355 8885 -2310 8935
rect -2260 8885 -2215 8935
rect -2165 8885 -2115 8935
rect -2065 8885 -2015 8935
rect -1965 8885 -1915 8935
rect -1865 8885 -1820 8935
rect -1770 8885 -1725 8935
rect -1675 8885 -1640 8935
rect -4840 8815 -1640 8885
rect -4840 8765 -4805 8815
rect -4755 8765 -4710 8815
rect -4660 8765 -4615 8815
rect -4565 8765 -4515 8815
rect -4465 8765 -4415 8815
rect -4365 8765 -4315 8815
rect -4265 8765 -4220 8815
rect -4170 8765 -4125 8815
rect -4075 8765 -4005 8815
rect -3955 8765 -3910 8815
rect -3860 8765 -3815 8815
rect -3765 8765 -3715 8815
rect -3665 8765 -3615 8815
rect -3565 8765 -3515 8815
rect -3465 8765 -3420 8815
rect -3370 8765 -3325 8815
rect -3275 8765 -3205 8815
rect -3155 8765 -3110 8815
rect -3060 8765 -3015 8815
rect -2965 8765 -2915 8815
rect -2865 8765 -2815 8815
rect -2765 8765 -2715 8815
rect -2665 8765 -2620 8815
rect -2570 8765 -2525 8815
rect -2475 8765 -2405 8815
rect -2355 8765 -2310 8815
rect -2260 8765 -2215 8815
rect -2165 8765 -2115 8815
rect -2065 8765 -2015 8815
rect -1965 8765 -1915 8815
rect -1865 8765 -1820 8815
rect -1770 8765 -1725 8815
rect -1675 8765 -1640 8815
rect -4840 8725 -1640 8765
rect -4840 8675 -4805 8725
rect -4755 8675 -4710 8725
rect -4660 8675 -4615 8725
rect -4565 8675 -4515 8725
rect -4465 8675 -4415 8725
rect -4365 8675 -4315 8725
rect -4265 8675 -4220 8725
rect -4170 8675 -4125 8725
rect -4075 8675 -4005 8725
rect -3955 8675 -3910 8725
rect -3860 8675 -3815 8725
rect -3765 8675 -3715 8725
rect -3665 8675 -3615 8725
rect -3565 8675 -3515 8725
rect -3465 8675 -3420 8725
rect -3370 8675 -3325 8725
rect -3275 8675 -3205 8725
rect -3155 8675 -3110 8725
rect -3060 8675 -3015 8725
rect -2965 8675 -2915 8725
rect -2865 8675 -2815 8725
rect -2765 8675 -2715 8725
rect -2665 8675 -2620 8725
rect -2570 8675 -2525 8725
rect -2475 8675 -2405 8725
rect -2355 8675 -2310 8725
rect -2260 8675 -2215 8725
rect -2165 8675 -2115 8725
rect -2065 8675 -2015 8725
rect -1965 8675 -1915 8725
rect -1865 8675 -1820 8725
rect -1770 8675 -1725 8725
rect -1675 8675 -1640 8725
rect -4840 8625 -1640 8675
rect -4840 8575 -4805 8625
rect -4755 8575 -4710 8625
rect -4660 8575 -4615 8625
rect -4565 8575 -4515 8625
rect -4465 8575 -4415 8625
rect -4365 8575 -4315 8625
rect -4265 8575 -4220 8625
rect -4170 8575 -4125 8625
rect -4075 8575 -4005 8625
rect -3955 8575 -3910 8625
rect -3860 8575 -3815 8625
rect -3765 8575 -3715 8625
rect -3665 8575 -3615 8625
rect -3565 8575 -3515 8625
rect -3465 8575 -3420 8625
rect -3370 8575 -3325 8625
rect -3275 8575 -3205 8625
rect -3155 8575 -3110 8625
rect -3060 8575 -3015 8625
rect -2965 8575 -2915 8625
rect -2865 8575 -2815 8625
rect -2765 8575 -2715 8625
rect -2665 8575 -2620 8625
rect -2570 8575 -2525 8625
rect -2475 8575 -2405 8625
rect -2355 8575 -2310 8625
rect -2260 8575 -2215 8625
rect -2165 8575 -2115 8625
rect -2065 8575 -2015 8625
rect -1965 8575 -1915 8625
rect -1865 8575 -1820 8625
rect -1770 8575 -1725 8625
rect -1675 8575 -1640 8625
rect -4840 8535 -1640 8575
rect -4840 8485 -4805 8535
rect -4755 8485 -4710 8535
rect -4660 8485 -4615 8535
rect -4565 8485 -4515 8535
rect -4465 8485 -4415 8535
rect -4365 8485 -4315 8535
rect -4265 8485 -4220 8535
rect -4170 8485 -4125 8535
rect -4075 8485 -4005 8535
rect -3955 8485 -3910 8535
rect -3860 8485 -3815 8535
rect -3765 8485 -3715 8535
rect -3665 8485 -3615 8535
rect -3565 8485 -3515 8535
rect -3465 8485 -3420 8535
rect -3370 8485 -3325 8535
rect -3275 8485 -3205 8535
rect -3155 8485 -3110 8535
rect -3060 8485 -3015 8535
rect -2965 8485 -2915 8535
rect -2865 8485 -2815 8535
rect -2765 8485 -2715 8535
rect -2665 8485 -2620 8535
rect -2570 8485 -2525 8535
rect -2475 8485 -2405 8535
rect -2355 8485 -2310 8535
rect -2260 8485 -2215 8535
rect -2165 8485 -2115 8535
rect -2065 8485 -2015 8535
rect -1965 8485 -1915 8535
rect -1865 8485 -1820 8535
rect -1770 8485 -1725 8535
rect -1675 8485 -1640 8535
rect -4840 8415 -1640 8485
rect -4840 8365 -4805 8415
rect -4755 8365 -4710 8415
rect -4660 8365 -4615 8415
rect -4565 8365 -4515 8415
rect -4465 8365 -4415 8415
rect -4365 8365 -4315 8415
rect -4265 8365 -4220 8415
rect -4170 8365 -4125 8415
rect -4075 8365 -4005 8415
rect -3955 8365 -3910 8415
rect -3860 8365 -3815 8415
rect -3765 8365 -3715 8415
rect -3665 8365 -3615 8415
rect -3565 8365 -3515 8415
rect -3465 8365 -3420 8415
rect -3370 8365 -3325 8415
rect -3275 8365 -3205 8415
rect -3155 8365 -3110 8415
rect -3060 8365 -3015 8415
rect -2965 8365 -2915 8415
rect -2865 8365 -2815 8415
rect -2765 8365 -2715 8415
rect -2665 8365 -2620 8415
rect -2570 8365 -2525 8415
rect -2475 8365 -2405 8415
rect -2355 8365 -2310 8415
rect -2260 8365 -2215 8415
rect -2165 8365 -2115 8415
rect -2065 8365 -2015 8415
rect -1965 8365 -1915 8415
rect -1865 8365 -1820 8415
rect -1770 8365 -1725 8415
rect -1675 8365 -1640 8415
rect -4840 8325 -1640 8365
rect -4840 8275 -4805 8325
rect -4755 8275 -4710 8325
rect -4660 8275 -4615 8325
rect -4565 8275 -4515 8325
rect -4465 8275 -4415 8325
rect -4365 8275 -4315 8325
rect -4265 8275 -4220 8325
rect -4170 8275 -4125 8325
rect -4075 8275 -4005 8325
rect -3955 8275 -3910 8325
rect -3860 8275 -3815 8325
rect -3765 8275 -3715 8325
rect -3665 8275 -3615 8325
rect -3565 8275 -3515 8325
rect -3465 8275 -3420 8325
rect -3370 8275 -3325 8325
rect -3275 8275 -3205 8325
rect -3155 8275 -3110 8325
rect -3060 8275 -3015 8325
rect -2965 8275 -2915 8325
rect -2865 8275 -2815 8325
rect -2765 8275 -2715 8325
rect -2665 8275 -2620 8325
rect -2570 8275 -2525 8325
rect -2475 8275 -2405 8325
rect -2355 8275 -2310 8325
rect -2260 8275 -2215 8325
rect -2165 8275 -2115 8325
rect -2065 8275 -2015 8325
rect -1965 8275 -1915 8325
rect -1865 8275 -1820 8325
rect -1770 8275 -1725 8325
rect -1675 8275 -1640 8325
rect -4840 8225 -1640 8275
rect -4840 8175 -4805 8225
rect -4755 8175 -4710 8225
rect -4660 8175 -4615 8225
rect -4565 8175 -4515 8225
rect -4465 8175 -4415 8225
rect -4365 8175 -4315 8225
rect -4265 8175 -4220 8225
rect -4170 8175 -4125 8225
rect -4075 8175 -4005 8225
rect -3955 8175 -3910 8225
rect -3860 8175 -3815 8225
rect -3765 8175 -3715 8225
rect -3665 8175 -3615 8225
rect -3565 8175 -3515 8225
rect -3465 8175 -3420 8225
rect -3370 8175 -3325 8225
rect -3275 8175 -3205 8225
rect -3155 8175 -3110 8225
rect -3060 8175 -3015 8225
rect -2965 8175 -2915 8225
rect -2865 8175 -2815 8225
rect -2765 8175 -2715 8225
rect -2665 8175 -2620 8225
rect -2570 8175 -2525 8225
rect -2475 8175 -2405 8225
rect -2355 8175 -2310 8225
rect -2260 8175 -2215 8225
rect -2165 8175 -2115 8225
rect -2065 8175 -2015 8225
rect -1965 8175 -1915 8225
rect -1865 8175 -1820 8225
rect -1770 8175 -1725 8225
rect -1675 8175 -1640 8225
rect -4840 8135 -1640 8175
rect -4840 8085 -4805 8135
rect -4755 8085 -4710 8135
rect -4660 8085 -4615 8135
rect -4565 8085 -4515 8135
rect -4465 8085 -4415 8135
rect -4365 8085 -4315 8135
rect -4265 8085 -4220 8135
rect -4170 8085 -4125 8135
rect -4075 8085 -4005 8135
rect -3955 8085 -3910 8135
rect -3860 8085 -3815 8135
rect -3765 8085 -3715 8135
rect -3665 8085 -3615 8135
rect -3565 8085 -3515 8135
rect -3465 8085 -3420 8135
rect -3370 8085 -3325 8135
rect -3275 8085 -3205 8135
rect -3155 8085 -3110 8135
rect -3060 8085 -3015 8135
rect -2965 8085 -2915 8135
rect -2865 8085 -2815 8135
rect -2765 8085 -2715 8135
rect -2665 8085 -2620 8135
rect -2570 8085 -2525 8135
rect -2475 8085 -2405 8135
rect -2355 8085 -2310 8135
rect -2260 8085 -2215 8135
rect -2165 8085 -2115 8135
rect -2065 8085 -2015 8135
rect -1965 8085 -1915 8135
rect -1865 8085 -1820 8135
rect -1770 8085 -1725 8135
rect -1675 8085 -1640 8135
rect -4840 8015 -1640 8085
rect -4840 7965 -4805 8015
rect -4755 7965 -4710 8015
rect -4660 7965 -4615 8015
rect -4565 7965 -4515 8015
rect -4465 7965 -4415 8015
rect -4365 7965 -4315 8015
rect -4265 7965 -4220 8015
rect -4170 7965 -4125 8015
rect -4075 7965 -4005 8015
rect -3955 7965 -3910 8015
rect -3860 7965 -3815 8015
rect -3765 7965 -3715 8015
rect -3665 7965 -3615 8015
rect -3565 7965 -3515 8015
rect -3465 7965 -3420 8015
rect -3370 7965 -3325 8015
rect -3275 7965 -3205 8015
rect -3155 7965 -3110 8015
rect -3060 7965 -3015 8015
rect -2965 7965 -2915 8015
rect -2865 7965 -2815 8015
rect -2765 7965 -2715 8015
rect -2665 7965 -2620 8015
rect -2570 7965 -2525 8015
rect -2475 7965 -2405 8015
rect -2355 7965 -2310 8015
rect -2260 7965 -2215 8015
rect -2165 7965 -2115 8015
rect -2065 7965 -2015 8015
rect -1965 7965 -1915 8015
rect -1865 7965 -1820 8015
rect -1770 7965 -1725 8015
rect -1675 7965 -1640 8015
rect -4840 7925 -1640 7965
rect -4840 7875 -4805 7925
rect -4755 7875 -4710 7925
rect -4660 7875 -4615 7925
rect -4565 7875 -4515 7925
rect -4465 7875 -4415 7925
rect -4365 7875 -4315 7925
rect -4265 7875 -4220 7925
rect -4170 7875 -4125 7925
rect -4075 7875 -4005 7925
rect -3955 7875 -3910 7925
rect -3860 7875 -3815 7925
rect -3765 7875 -3715 7925
rect -3665 7875 -3615 7925
rect -3565 7875 -3515 7925
rect -3465 7875 -3420 7925
rect -3370 7875 -3325 7925
rect -3275 7875 -3205 7925
rect -3155 7875 -3110 7925
rect -3060 7875 -3015 7925
rect -2965 7875 -2915 7925
rect -2865 7875 -2815 7925
rect -2765 7875 -2715 7925
rect -2665 7875 -2620 7925
rect -2570 7875 -2525 7925
rect -2475 7875 -2405 7925
rect -2355 7875 -2310 7925
rect -2260 7875 -2215 7925
rect -2165 7875 -2115 7925
rect -2065 7875 -2015 7925
rect -1965 7875 -1915 7925
rect -1865 7875 -1820 7925
rect -1770 7875 -1725 7925
rect -1675 7875 -1640 7925
rect -4840 7825 -1640 7875
rect -4840 7775 -4805 7825
rect -4755 7775 -4710 7825
rect -4660 7775 -4615 7825
rect -4565 7775 -4515 7825
rect -4465 7775 -4415 7825
rect -4365 7775 -4315 7825
rect -4265 7775 -4220 7825
rect -4170 7775 -4125 7825
rect -4075 7775 -4005 7825
rect -3955 7775 -3910 7825
rect -3860 7775 -3815 7825
rect -3765 7775 -3715 7825
rect -3665 7775 -3615 7825
rect -3565 7775 -3515 7825
rect -3465 7775 -3420 7825
rect -3370 7775 -3325 7825
rect -3275 7775 -3205 7825
rect -3155 7775 -3110 7825
rect -3060 7775 -3015 7825
rect -2965 7775 -2915 7825
rect -2865 7775 -2815 7825
rect -2765 7775 -2715 7825
rect -2665 7775 -2620 7825
rect -2570 7775 -2525 7825
rect -2475 7775 -2405 7825
rect -2355 7775 -2310 7825
rect -2260 7775 -2215 7825
rect -2165 7775 -2115 7825
rect -2065 7775 -2015 7825
rect -1965 7775 -1915 7825
rect -1865 7775 -1820 7825
rect -1770 7775 -1725 7825
rect -1675 7775 -1640 7825
rect -4840 7735 -1640 7775
rect -4840 7685 -4805 7735
rect -4755 7685 -4710 7735
rect -4660 7685 -4615 7735
rect -4565 7685 -4515 7735
rect -4465 7685 -4415 7735
rect -4365 7685 -4315 7735
rect -4265 7685 -4220 7735
rect -4170 7685 -4125 7735
rect -4075 7685 -4005 7735
rect -3955 7685 -3910 7735
rect -3860 7685 -3815 7735
rect -3765 7685 -3715 7735
rect -3665 7685 -3615 7735
rect -3565 7685 -3515 7735
rect -3465 7685 -3420 7735
rect -3370 7685 -3325 7735
rect -3275 7685 -3205 7735
rect -3155 7685 -3110 7735
rect -3060 7685 -3015 7735
rect -2965 7685 -2915 7735
rect -2865 7685 -2815 7735
rect -2765 7685 -2715 7735
rect -2665 7685 -2620 7735
rect -2570 7685 -2525 7735
rect -2475 7685 -2405 7735
rect -2355 7685 -2310 7735
rect -2260 7685 -2215 7735
rect -2165 7685 -2115 7735
rect -2065 7685 -2015 7735
rect -1965 7685 -1915 7735
rect -1865 7685 -1820 7735
rect -1770 7685 -1725 7735
rect -1675 7685 -1640 7735
rect -4840 7615 -1640 7685
rect -4840 7565 -4805 7615
rect -4755 7565 -4710 7615
rect -4660 7565 -4615 7615
rect -4565 7565 -4515 7615
rect -4465 7565 -4415 7615
rect -4365 7565 -4315 7615
rect -4265 7565 -4220 7615
rect -4170 7565 -4125 7615
rect -4075 7565 -4005 7615
rect -3955 7565 -3910 7615
rect -3860 7565 -3815 7615
rect -3765 7565 -3715 7615
rect -3665 7565 -3615 7615
rect -3565 7565 -3515 7615
rect -3465 7565 -3420 7615
rect -3370 7565 -3325 7615
rect -3275 7565 -3205 7615
rect -3155 7565 -3110 7615
rect -3060 7565 -3015 7615
rect -2965 7565 -2915 7615
rect -2865 7565 -2815 7615
rect -2765 7565 -2715 7615
rect -2665 7565 -2620 7615
rect -2570 7565 -2525 7615
rect -2475 7565 -2405 7615
rect -2355 7565 -2310 7615
rect -2260 7565 -2215 7615
rect -2165 7565 -2115 7615
rect -2065 7565 -2015 7615
rect -1965 7565 -1915 7615
rect -1865 7565 -1820 7615
rect -1770 7565 -1725 7615
rect -1675 7565 -1640 7615
rect -4840 7525 -1640 7565
rect -4840 7475 -4805 7525
rect -4755 7475 -4710 7525
rect -4660 7475 -4615 7525
rect -4565 7475 -4515 7525
rect -4465 7475 -4415 7525
rect -4365 7475 -4315 7525
rect -4265 7475 -4220 7525
rect -4170 7475 -4125 7525
rect -4075 7475 -4005 7525
rect -3955 7475 -3910 7525
rect -3860 7475 -3815 7525
rect -3765 7475 -3715 7525
rect -3665 7475 -3615 7525
rect -3565 7475 -3515 7525
rect -3465 7475 -3420 7525
rect -3370 7475 -3325 7525
rect -3275 7475 -3205 7525
rect -3155 7475 -3110 7525
rect -3060 7475 -3015 7525
rect -2965 7475 -2915 7525
rect -2865 7475 -2815 7525
rect -2765 7475 -2715 7525
rect -2665 7475 -2620 7525
rect -2570 7475 -2525 7525
rect -2475 7475 -2405 7525
rect -2355 7475 -2310 7525
rect -2260 7475 -2215 7525
rect -2165 7475 -2115 7525
rect -2065 7475 -2015 7525
rect -1965 7475 -1915 7525
rect -1865 7475 -1820 7525
rect -1770 7475 -1725 7525
rect -1675 7475 -1640 7525
rect -4840 7425 -1640 7475
rect -4840 7375 -4805 7425
rect -4755 7375 -4710 7425
rect -4660 7375 -4615 7425
rect -4565 7375 -4515 7425
rect -4465 7375 -4415 7425
rect -4365 7375 -4315 7425
rect -4265 7375 -4220 7425
rect -4170 7375 -4125 7425
rect -4075 7375 -4005 7425
rect -3955 7375 -3910 7425
rect -3860 7375 -3815 7425
rect -3765 7375 -3715 7425
rect -3665 7375 -3615 7425
rect -3565 7375 -3515 7425
rect -3465 7375 -3420 7425
rect -3370 7375 -3325 7425
rect -3275 7375 -3205 7425
rect -3155 7375 -3110 7425
rect -3060 7375 -3015 7425
rect -2965 7375 -2915 7425
rect -2865 7375 -2815 7425
rect -2765 7375 -2715 7425
rect -2665 7375 -2620 7425
rect -2570 7375 -2525 7425
rect -2475 7375 -2405 7425
rect -2355 7375 -2310 7425
rect -2260 7375 -2215 7425
rect -2165 7375 -2115 7425
rect -2065 7375 -2015 7425
rect -1965 7375 -1915 7425
rect -1865 7375 -1820 7425
rect -1770 7375 -1725 7425
rect -1675 7375 -1640 7425
rect -4840 7335 -1640 7375
rect -4840 7285 -4805 7335
rect -4755 7285 -4710 7335
rect -4660 7285 -4615 7335
rect -4565 7285 -4515 7335
rect -4465 7285 -4415 7335
rect -4365 7285 -4315 7335
rect -4265 7285 -4220 7335
rect -4170 7285 -4125 7335
rect -4075 7285 -4005 7335
rect -3955 7285 -3910 7335
rect -3860 7285 -3815 7335
rect -3765 7285 -3715 7335
rect -3665 7285 -3615 7335
rect -3565 7285 -3515 7335
rect -3465 7285 -3420 7335
rect -3370 7285 -3325 7335
rect -3275 7285 -3205 7335
rect -3155 7285 -3110 7335
rect -3060 7285 -3015 7335
rect -2965 7285 -2915 7335
rect -2865 7285 -2815 7335
rect -2765 7285 -2715 7335
rect -2665 7285 -2620 7335
rect -2570 7285 -2525 7335
rect -2475 7285 -2405 7335
rect -2355 7285 -2310 7335
rect -2260 7285 -2215 7335
rect -2165 7285 -2115 7335
rect -2065 7285 -2015 7335
rect -1965 7285 -1915 7335
rect -1865 7285 -1820 7335
rect -1770 7285 -1725 7335
rect -1675 7285 -1640 7335
rect -4840 7215 -1640 7285
rect -4840 7165 -4805 7215
rect -4755 7165 -4710 7215
rect -4660 7165 -4615 7215
rect -4565 7165 -4515 7215
rect -4465 7165 -4415 7215
rect -4365 7165 -4315 7215
rect -4265 7165 -4220 7215
rect -4170 7165 -4125 7215
rect -4075 7165 -4005 7215
rect -3955 7165 -3910 7215
rect -3860 7165 -3815 7215
rect -3765 7165 -3715 7215
rect -3665 7165 -3615 7215
rect -3565 7165 -3515 7215
rect -3465 7165 -3420 7215
rect -3370 7165 -3325 7215
rect -3275 7165 -3205 7215
rect -3155 7165 -3110 7215
rect -3060 7165 -3015 7215
rect -2965 7165 -2915 7215
rect -2865 7165 -2815 7215
rect -2765 7165 -2715 7215
rect -2665 7165 -2620 7215
rect -2570 7165 -2525 7215
rect -2475 7165 -2405 7215
rect -2355 7165 -2310 7215
rect -2260 7165 -2215 7215
rect -2165 7165 -2115 7215
rect -2065 7165 -2015 7215
rect -1965 7165 -1915 7215
rect -1865 7165 -1820 7215
rect -1770 7165 -1725 7215
rect -1675 7165 -1640 7215
rect -4840 7125 -1640 7165
rect -4840 7075 -4805 7125
rect -4755 7075 -4710 7125
rect -4660 7075 -4615 7125
rect -4565 7075 -4515 7125
rect -4465 7075 -4415 7125
rect -4365 7075 -4315 7125
rect -4265 7075 -4220 7125
rect -4170 7075 -4125 7125
rect -4075 7075 -4005 7125
rect -3955 7075 -3910 7125
rect -3860 7075 -3815 7125
rect -3765 7075 -3715 7125
rect -3665 7075 -3615 7125
rect -3565 7075 -3515 7125
rect -3465 7075 -3420 7125
rect -3370 7075 -3325 7125
rect -3275 7075 -3205 7125
rect -3155 7075 -3110 7125
rect -3060 7075 -3015 7125
rect -2965 7075 -2915 7125
rect -2865 7075 -2815 7125
rect -2765 7075 -2715 7125
rect -2665 7075 -2620 7125
rect -2570 7075 -2525 7125
rect -2475 7075 -2405 7125
rect -2355 7075 -2310 7125
rect -2260 7075 -2215 7125
rect -2165 7075 -2115 7125
rect -2065 7075 -2015 7125
rect -1965 7075 -1915 7125
rect -1865 7075 -1820 7125
rect -1770 7075 -1725 7125
rect -1675 7075 -1640 7125
rect -4840 7025 -1640 7075
rect -4840 6975 -4805 7025
rect -4755 6975 -4710 7025
rect -4660 6975 -4615 7025
rect -4565 6975 -4515 7025
rect -4465 6975 -4415 7025
rect -4365 6975 -4315 7025
rect -4265 6975 -4220 7025
rect -4170 6975 -4125 7025
rect -4075 6975 -4005 7025
rect -3955 6975 -3910 7025
rect -3860 6975 -3815 7025
rect -3765 6975 -3715 7025
rect -3665 6975 -3615 7025
rect -3565 6975 -3515 7025
rect -3465 6975 -3420 7025
rect -3370 6975 -3325 7025
rect -3275 6975 -3205 7025
rect -3155 6975 -3110 7025
rect -3060 6975 -3015 7025
rect -2965 6975 -2915 7025
rect -2865 6975 -2815 7025
rect -2765 6975 -2715 7025
rect -2665 6975 -2620 7025
rect -2570 6975 -2525 7025
rect -2475 6975 -2405 7025
rect -2355 6975 -2310 7025
rect -2260 6975 -2215 7025
rect -2165 6975 -2115 7025
rect -2065 6975 -2015 7025
rect -1965 6975 -1915 7025
rect -1865 6975 -1820 7025
rect -1770 6975 -1725 7025
rect -1675 6975 -1640 7025
rect -4840 6935 -1640 6975
rect -4840 6885 -4805 6935
rect -4755 6885 -4710 6935
rect -4660 6885 -4615 6935
rect -4565 6885 -4515 6935
rect -4465 6885 -4415 6935
rect -4365 6885 -4315 6935
rect -4265 6885 -4220 6935
rect -4170 6885 -4125 6935
rect -4075 6885 -4005 6935
rect -3955 6885 -3910 6935
rect -3860 6885 -3815 6935
rect -3765 6885 -3715 6935
rect -3665 6885 -3615 6935
rect -3565 6885 -3515 6935
rect -3465 6885 -3420 6935
rect -3370 6885 -3325 6935
rect -3275 6885 -3205 6935
rect -3155 6885 -3110 6935
rect -3060 6885 -3015 6935
rect -2965 6885 -2915 6935
rect -2865 6885 -2815 6935
rect -2765 6885 -2715 6935
rect -2665 6885 -2620 6935
rect -2570 6885 -2525 6935
rect -2475 6885 -2405 6935
rect -2355 6885 -2310 6935
rect -2260 6885 -2215 6935
rect -2165 6885 -2115 6935
rect -2065 6885 -2015 6935
rect -1965 6885 -1915 6935
rect -1865 6885 -1820 6935
rect -1770 6885 -1725 6935
rect -1675 6885 -1640 6935
rect -4840 6815 -1640 6885
rect -4840 6765 -4805 6815
rect -4755 6765 -4710 6815
rect -4660 6765 -4615 6815
rect -4565 6765 -4515 6815
rect -4465 6765 -4415 6815
rect -4365 6765 -4315 6815
rect -4265 6765 -4220 6815
rect -4170 6765 -4125 6815
rect -4075 6765 -4005 6815
rect -3955 6765 -3910 6815
rect -3860 6765 -3815 6815
rect -3765 6765 -3715 6815
rect -3665 6765 -3615 6815
rect -3565 6765 -3515 6815
rect -3465 6765 -3420 6815
rect -3370 6765 -3325 6815
rect -3275 6765 -3205 6815
rect -3155 6765 -3110 6815
rect -3060 6765 -3015 6815
rect -2965 6765 -2915 6815
rect -2865 6765 -2815 6815
rect -2765 6765 -2715 6815
rect -2665 6765 -2620 6815
rect -2570 6765 -2525 6815
rect -2475 6765 -2405 6815
rect -2355 6765 -2310 6815
rect -2260 6765 -2215 6815
rect -2165 6765 -2115 6815
rect -2065 6765 -2015 6815
rect -1965 6765 -1915 6815
rect -1865 6765 -1820 6815
rect -1770 6765 -1725 6815
rect -1675 6765 -1640 6815
rect -4840 6725 -1640 6765
rect -4840 6675 -4805 6725
rect -4755 6675 -4710 6725
rect -4660 6675 -4615 6725
rect -4565 6675 -4515 6725
rect -4465 6675 -4415 6725
rect -4365 6675 -4315 6725
rect -4265 6675 -4220 6725
rect -4170 6675 -4125 6725
rect -4075 6675 -4005 6725
rect -3955 6675 -3910 6725
rect -3860 6675 -3815 6725
rect -3765 6675 -3715 6725
rect -3665 6675 -3615 6725
rect -3565 6675 -3515 6725
rect -3465 6675 -3420 6725
rect -3370 6675 -3325 6725
rect -3275 6675 -3205 6725
rect -3155 6675 -3110 6725
rect -3060 6675 -3015 6725
rect -2965 6675 -2915 6725
rect -2865 6675 -2815 6725
rect -2765 6675 -2715 6725
rect -2665 6675 -2620 6725
rect -2570 6675 -2525 6725
rect -2475 6675 -2405 6725
rect -2355 6675 -2310 6725
rect -2260 6675 -2215 6725
rect -2165 6675 -2115 6725
rect -2065 6675 -2015 6725
rect -1965 6675 -1915 6725
rect -1865 6675 -1820 6725
rect -1770 6675 -1725 6725
rect -1675 6675 -1640 6725
rect -4840 6625 -1640 6675
rect -4840 6575 -4805 6625
rect -4755 6575 -4710 6625
rect -4660 6575 -4615 6625
rect -4565 6575 -4515 6625
rect -4465 6575 -4415 6625
rect -4365 6575 -4315 6625
rect -4265 6575 -4220 6625
rect -4170 6575 -4125 6625
rect -4075 6575 -4005 6625
rect -3955 6575 -3910 6625
rect -3860 6575 -3815 6625
rect -3765 6575 -3715 6625
rect -3665 6575 -3615 6625
rect -3565 6575 -3515 6625
rect -3465 6575 -3420 6625
rect -3370 6575 -3325 6625
rect -3275 6575 -3205 6625
rect -3155 6575 -3110 6625
rect -3060 6575 -3015 6625
rect -2965 6575 -2915 6625
rect -2865 6575 -2815 6625
rect -2765 6575 -2715 6625
rect -2665 6575 -2620 6625
rect -2570 6575 -2525 6625
rect -2475 6575 -2405 6625
rect -2355 6575 -2310 6625
rect -2260 6575 -2215 6625
rect -2165 6575 -2115 6625
rect -2065 6575 -2015 6625
rect -1965 6575 -1915 6625
rect -1865 6575 -1820 6625
rect -1770 6575 -1725 6625
rect -1675 6575 -1640 6625
rect -4840 6535 -1640 6575
rect -4840 6485 -4805 6535
rect -4755 6485 -4710 6535
rect -4660 6485 -4615 6535
rect -4565 6485 -4515 6535
rect -4465 6485 -4415 6535
rect -4365 6485 -4315 6535
rect -4265 6485 -4220 6535
rect -4170 6485 -4125 6535
rect -4075 6485 -4005 6535
rect -3955 6485 -3910 6535
rect -3860 6485 -3815 6535
rect -3765 6485 -3715 6535
rect -3665 6485 -3615 6535
rect -3565 6485 -3515 6535
rect -3465 6485 -3420 6535
rect -3370 6485 -3325 6535
rect -3275 6485 -3205 6535
rect -3155 6485 -3110 6535
rect -3060 6485 -3015 6535
rect -2965 6485 -2915 6535
rect -2865 6485 -2815 6535
rect -2765 6485 -2715 6535
rect -2665 6485 -2620 6535
rect -2570 6485 -2525 6535
rect -2475 6485 -2405 6535
rect -2355 6485 -2310 6535
rect -2260 6485 -2215 6535
rect -2165 6485 -2115 6535
rect -2065 6485 -2015 6535
rect -1965 6485 -1915 6535
rect -1865 6485 -1820 6535
rect -1770 6485 -1725 6535
rect -1675 6485 -1640 6535
rect -4840 6450 -1640 6485
rect -90 9640 -30 9650
rect -90 9600 -80 9640
rect -40 9600 -30 9640
rect -90 9575 -30 9600
rect -90 9535 -80 9575
rect -40 9535 -30 9575
rect -90 9505 -30 9535
rect -90 9465 -80 9505
rect -40 9465 -30 9505
rect -90 9435 -30 9465
rect -90 9395 -80 9435
rect -40 9395 -30 9435
rect -90 9365 -30 9395
rect -90 9325 -80 9365
rect -40 9325 -30 9365
rect -90 9300 -30 9325
rect -90 9260 -80 9300
rect -40 9260 -30 9300
rect -90 9240 -30 9260
rect -90 9200 -80 9240
rect -40 9200 -30 9240
rect -90 9175 -30 9200
rect -90 9135 -80 9175
rect -40 9135 -30 9175
rect -90 9105 -30 9135
rect -90 9065 -80 9105
rect -40 9065 -30 9105
rect -90 9035 -30 9065
rect -90 8995 -80 9035
rect -40 8995 -30 9035
rect -90 8965 -30 8995
rect -90 8925 -80 8965
rect -40 8925 -30 8965
rect -90 8900 -30 8925
rect -90 8860 -80 8900
rect -40 8860 -30 8900
rect -90 8840 -30 8860
rect -90 8800 -80 8840
rect -40 8800 -30 8840
rect -90 8775 -30 8800
rect -90 8735 -80 8775
rect -40 8735 -30 8775
rect -90 8705 -30 8735
rect -90 8665 -80 8705
rect -40 8665 -30 8705
rect -90 8635 -30 8665
rect -90 8595 -80 8635
rect -40 8595 -30 8635
rect -90 8565 -30 8595
rect -90 8525 -80 8565
rect -40 8525 -30 8565
rect -90 8500 -30 8525
rect -90 8460 -80 8500
rect -40 8460 -30 8500
rect -90 8440 -30 8460
rect -90 8400 -80 8440
rect -40 8400 -30 8440
rect -90 8375 -30 8400
rect -90 8335 -80 8375
rect -40 8335 -30 8375
rect -90 8305 -30 8335
rect -90 8265 -80 8305
rect -40 8265 -30 8305
rect -90 8235 -30 8265
rect -90 8195 -80 8235
rect -40 8195 -30 8235
rect -90 8165 -30 8195
rect -90 8125 -80 8165
rect -40 8125 -30 8165
rect -90 8100 -30 8125
rect -90 8060 -80 8100
rect -40 8060 -30 8100
rect -90 8040 -30 8060
rect -90 8000 -80 8040
rect -40 8000 -30 8040
rect -90 7975 -30 8000
rect -90 7935 -80 7975
rect -40 7935 -30 7975
rect -90 7905 -30 7935
rect -90 7865 -80 7905
rect -40 7865 -30 7905
rect -90 7835 -30 7865
rect -90 7795 -80 7835
rect -40 7795 -30 7835
rect -90 7765 -30 7795
rect -90 7725 -80 7765
rect -40 7725 -30 7765
rect -90 7700 -30 7725
rect -90 7660 -80 7700
rect -40 7660 -30 7700
rect -90 7640 -30 7660
rect -90 7600 -80 7640
rect -40 7600 -30 7640
rect -90 7575 -30 7600
rect -90 7535 -80 7575
rect -40 7535 -30 7575
rect -90 7505 -30 7535
rect -90 7465 -80 7505
rect -40 7465 -30 7505
rect -90 7435 -30 7465
rect -90 7395 -80 7435
rect -40 7395 -30 7435
rect -90 7365 -30 7395
rect -90 7325 -80 7365
rect -40 7325 -30 7365
rect -90 7300 -30 7325
rect -90 7260 -80 7300
rect -40 7260 -30 7300
rect -90 7240 -30 7260
rect -90 7200 -80 7240
rect -40 7200 -30 7240
rect -90 7175 -30 7200
rect -90 7135 -80 7175
rect -40 7135 -30 7175
rect -90 7105 -30 7135
rect -90 7065 -80 7105
rect -40 7065 -30 7105
rect -90 7035 -30 7065
rect -90 6995 -80 7035
rect -40 6995 -30 7035
rect -90 6965 -30 6995
rect -90 6925 -80 6965
rect -40 6925 -30 6965
rect -90 6900 -30 6925
rect -90 6860 -80 6900
rect -40 6860 -30 6900
rect -90 6840 -30 6860
rect -90 6800 -80 6840
rect -40 6800 -30 6840
rect -90 6775 -30 6800
rect -90 6735 -80 6775
rect -40 6735 -30 6775
rect -90 6705 -30 6735
rect -90 6665 -80 6705
rect -40 6665 -30 6705
rect -90 6635 -30 6665
rect -90 6595 -80 6635
rect -40 6595 -30 6635
rect -90 6565 -30 6595
rect -90 6525 -80 6565
rect -40 6525 -30 6565
rect -90 6500 -30 6525
rect -90 6460 -80 6500
rect -40 6460 -30 6500
rect -90 6450 -30 6460
rect 260 9640 320 9650
rect 260 9600 270 9640
rect 310 9600 320 9640
rect 260 9575 320 9600
rect 260 9535 270 9575
rect 310 9535 320 9575
rect 260 9505 320 9535
rect 260 9465 270 9505
rect 310 9465 320 9505
rect 260 9435 320 9465
rect 260 9395 270 9435
rect 310 9395 320 9435
rect 260 9365 320 9395
rect 260 9325 270 9365
rect 310 9325 320 9365
rect 260 9300 320 9325
rect 260 9260 270 9300
rect 310 9260 320 9300
rect 260 9240 320 9260
rect 260 9200 270 9240
rect 310 9200 320 9240
rect 260 9175 320 9200
rect 260 9135 270 9175
rect 310 9135 320 9175
rect 260 9105 320 9135
rect 260 9065 270 9105
rect 310 9065 320 9105
rect 260 9035 320 9065
rect 260 8995 270 9035
rect 310 8995 320 9035
rect 260 8965 320 8995
rect 260 8925 270 8965
rect 310 8925 320 8965
rect 260 8900 320 8925
rect 260 8860 270 8900
rect 310 8860 320 8900
rect 260 8840 320 8860
rect 260 8800 270 8840
rect 310 8800 320 8840
rect 260 8775 320 8800
rect 260 8735 270 8775
rect 310 8735 320 8775
rect 260 8705 320 8735
rect 260 8665 270 8705
rect 310 8665 320 8705
rect 260 8635 320 8665
rect 260 8595 270 8635
rect 310 8595 320 8635
rect 260 8565 320 8595
rect 260 8525 270 8565
rect 310 8525 320 8565
rect 260 8500 320 8525
rect 260 8460 270 8500
rect 310 8460 320 8500
rect 260 8440 320 8460
rect 260 8400 270 8440
rect 310 8400 320 8440
rect 260 8375 320 8400
rect 260 8335 270 8375
rect 310 8335 320 8375
rect 260 8305 320 8335
rect 260 8265 270 8305
rect 310 8265 320 8305
rect 260 8235 320 8265
rect 260 8195 270 8235
rect 310 8195 320 8235
rect 260 8165 320 8195
rect 260 8125 270 8165
rect 310 8125 320 8165
rect 260 8100 320 8125
rect 260 8060 270 8100
rect 310 8060 320 8100
rect 260 8040 320 8060
rect 260 8000 270 8040
rect 310 8000 320 8040
rect 260 7975 320 8000
rect 260 7935 270 7975
rect 310 7935 320 7975
rect 260 7905 320 7935
rect 260 7865 270 7905
rect 310 7865 320 7905
rect 260 7835 320 7865
rect 260 7795 270 7835
rect 310 7795 320 7835
rect 260 7765 320 7795
rect 260 7725 270 7765
rect 310 7725 320 7765
rect 260 7700 320 7725
rect 260 7660 270 7700
rect 310 7660 320 7700
rect 260 7640 320 7660
rect 260 7600 270 7640
rect 310 7600 320 7640
rect 260 7575 320 7600
rect 260 7535 270 7575
rect 310 7535 320 7575
rect 260 7505 320 7535
rect 260 7465 270 7505
rect 310 7465 320 7505
rect 260 7435 320 7465
rect 260 7395 270 7435
rect 310 7395 320 7435
rect 260 7365 320 7395
rect 260 7325 270 7365
rect 310 7325 320 7365
rect 260 7300 320 7325
rect 260 7260 270 7300
rect 310 7260 320 7300
rect 260 7240 320 7260
rect 260 7200 270 7240
rect 310 7200 320 7240
rect 260 7175 320 7200
rect 260 7135 270 7175
rect 310 7135 320 7175
rect 260 7105 320 7135
rect 260 7065 270 7105
rect 310 7065 320 7105
rect 260 7035 320 7065
rect 260 6995 270 7035
rect 310 6995 320 7035
rect 260 6965 320 6995
rect 260 6925 270 6965
rect 310 6925 320 6965
rect 260 6900 320 6925
rect 260 6860 270 6900
rect 310 6860 320 6900
rect 260 6840 320 6860
rect 260 6800 270 6840
rect 310 6800 320 6840
rect 260 6775 320 6800
rect 260 6735 270 6775
rect 310 6735 320 6775
rect 260 6705 320 6735
rect 260 6665 270 6705
rect 310 6665 320 6705
rect 260 6635 320 6665
rect 260 6595 270 6635
rect 310 6595 320 6635
rect 260 6565 320 6595
rect 260 6525 270 6565
rect 310 6525 320 6565
rect 260 6500 320 6525
rect 260 6460 270 6500
rect 310 6460 320 6500
rect 260 6450 320 6460
rect 610 9640 670 9650
rect 610 9600 620 9640
rect 660 9600 670 9640
rect 610 9575 670 9600
rect 610 9535 620 9575
rect 660 9535 670 9575
rect 610 9505 670 9535
rect 610 9465 620 9505
rect 660 9465 670 9505
rect 610 9435 670 9465
rect 610 9395 620 9435
rect 660 9395 670 9435
rect 610 9365 670 9395
rect 610 9325 620 9365
rect 660 9325 670 9365
rect 610 9300 670 9325
rect 610 9260 620 9300
rect 660 9260 670 9300
rect 610 9240 670 9260
rect 610 9200 620 9240
rect 660 9200 670 9240
rect 610 9175 670 9200
rect 610 9135 620 9175
rect 660 9135 670 9175
rect 610 9105 670 9135
rect 610 9065 620 9105
rect 660 9065 670 9105
rect 610 9035 670 9065
rect 610 8995 620 9035
rect 660 8995 670 9035
rect 610 8965 670 8995
rect 610 8925 620 8965
rect 660 8925 670 8965
rect 610 8900 670 8925
rect 610 8860 620 8900
rect 660 8860 670 8900
rect 610 8840 670 8860
rect 610 8800 620 8840
rect 660 8800 670 8840
rect 610 8775 670 8800
rect 610 8735 620 8775
rect 660 8735 670 8775
rect 610 8705 670 8735
rect 610 8665 620 8705
rect 660 8665 670 8705
rect 610 8635 670 8665
rect 610 8595 620 8635
rect 660 8595 670 8635
rect 610 8565 670 8595
rect 610 8525 620 8565
rect 660 8525 670 8565
rect 610 8500 670 8525
rect 610 8460 620 8500
rect 660 8460 670 8500
rect 610 8440 670 8460
rect 610 8400 620 8440
rect 660 8400 670 8440
rect 610 8375 670 8400
rect 610 8335 620 8375
rect 660 8335 670 8375
rect 610 8305 670 8335
rect 610 8265 620 8305
rect 660 8265 670 8305
rect 610 8235 670 8265
rect 610 8195 620 8235
rect 660 8195 670 8235
rect 610 8165 670 8195
rect 610 8125 620 8165
rect 660 8125 670 8165
rect 610 8100 670 8125
rect 610 8060 620 8100
rect 660 8060 670 8100
rect 610 8040 670 8060
rect 610 8000 620 8040
rect 660 8000 670 8040
rect 610 7975 670 8000
rect 610 7935 620 7975
rect 660 7935 670 7975
rect 610 7905 670 7935
rect 610 7865 620 7905
rect 660 7865 670 7905
rect 610 7835 670 7865
rect 610 7795 620 7835
rect 660 7795 670 7835
rect 610 7765 670 7795
rect 610 7725 620 7765
rect 660 7725 670 7765
rect 610 7700 670 7725
rect 610 7660 620 7700
rect 660 7660 670 7700
rect 610 7640 670 7660
rect 610 7600 620 7640
rect 660 7600 670 7640
rect 610 7575 670 7600
rect 610 7535 620 7575
rect 660 7535 670 7575
rect 610 7505 670 7535
rect 610 7465 620 7505
rect 660 7465 670 7505
rect 610 7435 670 7465
rect 610 7395 620 7435
rect 660 7395 670 7435
rect 610 7365 670 7395
rect 610 7325 620 7365
rect 660 7325 670 7365
rect 610 7300 670 7325
rect 610 7260 620 7300
rect 660 7260 670 7300
rect 610 7240 670 7260
rect 610 7200 620 7240
rect 660 7200 670 7240
rect 610 7175 670 7200
rect 610 7135 620 7175
rect 660 7135 670 7175
rect 610 7105 670 7135
rect 610 7065 620 7105
rect 660 7065 670 7105
rect 610 7035 670 7065
rect 610 6995 620 7035
rect 660 6995 670 7035
rect 610 6965 670 6995
rect 610 6925 620 6965
rect 660 6925 670 6965
rect 610 6900 670 6925
rect 610 6860 620 6900
rect 660 6860 670 6900
rect 610 6840 670 6860
rect 610 6800 620 6840
rect 660 6800 670 6840
rect 610 6775 670 6800
rect 610 6735 620 6775
rect 660 6735 670 6775
rect 610 6705 670 6735
rect 610 6665 620 6705
rect 660 6665 670 6705
rect 610 6635 670 6665
rect 610 6595 620 6635
rect 660 6595 670 6635
rect 610 6565 670 6595
rect 610 6525 620 6565
rect 660 6525 670 6565
rect 610 6500 670 6525
rect 610 6460 620 6500
rect 660 6460 670 6500
rect 610 6450 670 6460
rect 960 9640 1020 9650
rect 960 9600 970 9640
rect 1010 9600 1020 9640
rect 960 9575 1020 9600
rect 960 9535 970 9575
rect 1010 9535 1020 9575
rect 960 9505 1020 9535
rect 960 9465 970 9505
rect 1010 9465 1020 9505
rect 960 9435 1020 9465
rect 960 9395 970 9435
rect 1010 9395 1020 9435
rect 960 9365 1020 9395
rect 960 9325 970 9365
rect 1010 9325 1020 9365
rect 960 9300 1020 9325
rect 960 9260 970 9300
rect 1010 9260 1020 9300
rect 960 9240 1020 9260
rect 960 9200 970 9240
rect 1010 9200 1020 9240
rect 960 9175 1020 9200
rect 960 9135 970 9175
rect 1010 9135 1020 9175
rect 960 9105 1020 9135
rect 960 9065 970 9105
rect 1010 9065 1020 9105
rect 960 9035 1020 9065
rect 960 8995 970 9035
rect 1010 8995 1020 9035
rect 960 8965 1020 8995
rect 960 8925 970 8965
rect 1010 8925 1020 8965
rect 960 8900 1020 8925
rect 960 8860 970 8900
rect 1010 8860 1020 8900
rect 960 8840 1020 8860
rect 960 8800 970 8840
rect 1010 8800 1020 8840
rect 960 8775 1020 8800
rect 960 8735 970 8775
rect 1010 8735 1020 8775
rect 960 8705 1020 8735
rect 960 8665 970 8705
rect 1010 8665 1020 8705
rect 960 8635 1020 8665
rect 960 8595 970 8635
rect 1010 8595 1020 8635
rect 960 8565 1020 8595
rect 960 8525 970 8565
rect 1010 8525 1020 8565
rect 960 8500 1020 8525
rect 960 8460 970 8500
rect 1010 8460 1020 8500
rect 960 8440 1020 8460
rect 960 8400 970 8440
rect 1010 8400 1020 8440
rect 960 8375 1020 8400
rect 960 8335 970 8375
rect 1010 8335 1020 8375
rect 960 8305 1020 8335
rect 960 8265 970 8305
rect 1010 8265 1020 8305
rect 960 8235 1020 8265
rect 960 8195 970 8235
rect 1010 8195 1020 8235
rect 960 8165 1020 8195
rect 960 8125 970 8165
rect 1010 8125 1020 8165
rect 960 8100 1020 8125
rect 960 8060 970 8100
rect 1010 8060 1020 8100
rect 960 8040 1020 8060
rect 960 8000 970 8040
rect 1010 8000 1020 8040
rect 960 7975 1020 8000
rect 960 7935 970 7975
rect 1010 7935 1020 7975
rect 960 7905 1020 7935
rect 960 7865 970 7905
rect 1010 7865 1020 7905
rect 960 7835 1020 7865
rect 960 7795 970 7835
rect 1010 7795 1020 7835
rect 960 7765 1020 7795
rect 960 7725 970 7765
rect 1010 7725 1020 7765
rect 960 7700 1020 7725
rect 960 7660 970 7700
rect 1010 7660 1020 7700
rect 960 7640 1020 7660
rect 960 7600 970 7640
rect 1010 7600 1020 7640
rect 960 7575 1020 7600
rect 960 7535 970 7575
rect 1010 7535 1020 7575
rect 960 7505 1020 7535
rect 960 7465 970 7505
rect 1010 7465 1020 7505
rect 960 7435 1020 7465
rect 960 7395 970 7435
rect 1010 7395 1020 7435
rect 960 7365 1020 7395
rect 960 7325 970 7365
rect 1010 7325 1020 7365
rect 960 7300 1020 7325
rect 960 7260 970 7300
rect 1010 7260 1020 7300
rect 960 7240 1020 7260
rect 960 7200 970 7240
rect 1010 7200 1020 7240
rect 960 7175 1020 7200
rect 960 7135 970 7175
rect 1010 7135 1020 7175
rect 960 7105 1020 7135
rect 960 7065 970 7105
rect 1010 7065 1020 7105
rect 960 7035 1020 7065
rect 960 6995 970 7035
rect 1010 6995 1020 7035
rect 960 6965 1020 6995
rect 960 6925 970 6965
rect 1010 6925 1020 6965
rect 960 6900 1020 6925
rect 960 6860 970 6900
rect 1010 6860 1020 6900
rect 960 6840 1020 6860
rect 960 6800 970 6840
rect 1010 6800 1020 6840
rect 960 6775 1020 6800
rect 960 6735 970 6775
rect 1010 6735 1020 6775
rect 960 6705 1020 6735
rect 960 6665 970 6705
rect 1010 6665 1020 6705
rect 960 6635 1020 6665
rect 960 6595 970 6635
rect 1010 6595 1020 6635
rect 960 6565 1020 6595
rect 960 6525 970 6565
rect 1010 6525 1020 6565
rect 960 6500 1020 6525
rect 960 6460 970 6500
rect 1010 6460 1020 6500
rect 960 6450 1020 6460
rect 1660 9640 1720 9650
rect 1660 9600 1670 9640
rect 1710 9600 1720 9640
rect 1660 9575 1720 9600
rect 1660 9535 1670 9575
rect 1710 9535 1720 9575
rect 1660 9505 1720 9535
rect 1660 9465 1670 9505
rect 1710 9465 1720 9505
rect 1660 9435 1720 9465
rect 1660 9395 1670 9435
rect 1710 9395 1720 9435
rect 1660 9365 1720 9395
rect 1660 9325 1670 9365
rect 1710 9325 1720 9365
rect 1660 9300 1720 9325
rect 1660 9260 1670 9300
rect 1710 9260 1720 9300
rect 1660 9240 1720 9260
rect 1660 9200 1670 9240
rect 1710 9200 1720 9240
rect 1660 9175 1720 9200
rect 1660 9135 1670 9175
rect 1710 9135 1720 9175
rect 1660 9105 1720 9135
rect 1660 9065 1670 9105
rect 1710 9065 1720 9105
rect 1660 9035 1720 9065
rect 1660 8995 1670 9035
rect 1710 8995 1720 9035
rect 1660 8965 1720 8995
rect 1660 8925 1670 8965
rect 1710 8925 1720 8965
rect 1660 8900 1720 8925
rect 1660 8860 1670 8900
rect 1710 8860 1720 8900
rect 1660 8840 1720 8860
rect 1660 8800 1670 8840
rect 1710 8800 1720 8840
rect 1660 8775 1720 8800
rect 1660 8735 1670 8775
rect 1710 8735 1720 8775
rect 1660 8705 1720 8735
rect 1660 8665 1670 8705
rect 1710 8665 1720 8705
rect 1660 8635 1720 8665
rect 1660 8595 1670 8635
rect 1710 8595 1720 8635
rect 1660 8565 1720 8595
rect 1660 8525 1670 8565
rect 1710 8525 1720 8565
rect 1660 8500 1720 8525
rect 1660 8460 1670 8500
rect 1710 8460 1720 8500
rect 1660 8440 1720 8460
rect 1660 8400 1670 8440
rect 1710 8400 1720 8440
rect 1660 8375 1720 8400
rect 1660 8335 1670 8375
rect 1710 8335 1720 8375
rect 1660 8305 1720 8335
rect 1660 8265 1670 8305
rect 1710 8265 1720 8305
rect 1660 8235 1720 8265
rect 1660 8195 1670 8235
rect 1710 8195 1720 8235
rect 1660 8165 1720 8195
rect 1660 8125 1670 8165
rect 1710 8125 1720 8165
rect 1660 8100 1720 8125
rect 1660 8060 1670 8100
rect 1710 8060 1720 8100
rect 1660 8040 1720 8060
rect 1660 8000 1670 8040
rect 1710 8000 1720 8040
rect 1660 7975 1720 8000
rect 1660 7935 1670 7975
rect 1710 7935 1720 7975
rect 1660 7905 1720 7935
rect 1660 7865 1670 7905
rect 1710 7865 1720 7905
rect 1660 7835 1720 7865
rect 1660 7795 1670 7835
rect 1710 7795 1720 7835
rect 1660 7765 1720 7795
rect 1660 7725 1670 7765
rect 1710 7725 1720 7765
rect 1660 7700 1720 7725
rect 1660 7660 1670 7700
rect 1710 7660 1720 7700
rect 1660 7640 1720 7660
rect 1660 7600 1670 7640
rect 1710 7600 1720 7640
rect 1660 7575 1720 7600
rect 1660 7535 1670 7575
rect 1710 7535 1720 7575
rect 1660 7505 1720 7535
rect 1660 7465 1670 7505
rect 1710 7465 1720 7505
rect 1660 7435 1720 7465
rect 1660 7395 1670 7435
rect 1710 7395 1720 7435
rect 1660 7365 1720 7395
rect 1660 7325 1670 7365
rect 1710 7325 1720 7365
rect 1660 7300 1720 7325
rect 1660 7260 1670 7300
rect 1710 7260 1720 7300
rect 1660 7240 1720 7260
rect 1660 7200 1670 7240
rect 1710 7200 1720 7240
rect 1660 7175 1720 7200
rect 1660 7135 1670 7175
rect 1710 7135 1720 7175
rect 1660 7105 1720 7135
rect 1660 7065 1670 7105
rect 1710 7065 1720 7105
rect 1660 7035 1720 7065
rect 1660 6995 1670 7035
rect 1710 6995 1720 7035
rect 1660 6965 1720 6995
rect 1660 6925 1670 6965
rect 1710 6925 1720 6965
rect 1660 6900 1720 6925
rect 1660 6860 1670 6900
rect 1710 6860 1720 6900
rect 1660 6840 1720 6860
rect 1660 6800 1670 6840
rect 1710 6800 1720 6840
rect 1660 6775 1720 6800
rect 1660 6735 1670 6775
rect 1710 6735 1720 6775
rect 1660 6705 1720 6735
rect 1660 6665 1670 6705
rect 1710 6665 1720 6705
rect 1660 6635 1720 6665
rect 1660 6595 1670 6635
rect 1710 6595 1720 6635
rect 1660 6565 1720 6595
rect 1660 6525 1670 6565
rect 1710 6525 1720 6565
rect 1660 6500 1720 6525
rect 1660 6460 1670 6500
rect 1710 6460 1720 6500
rect 1660 6450 1720 6460
rect 2315 9640 2375 9650
rect 2315 9600 2325 9640
rect 2365 9600 2375 9640
rect 2315 9575 2375 9600
rect 2315 9535 2325 9575
rect 2365 9535 2375 9575
rect 2315 9505 2375 9535
rect 2315 9465 2325 9505
rect 2365 9465 2375 9505
rect 2315 9435 2375 9465
rect 2315 9395 2325 9435
rect 2365 9395 2375 9435
rect 2315 9365 2375 9395
rect 2315 9325 2325 9365
rect 2365 9325 2375 9365
rect 2315 9300 2375 9325
rect 2315 9260 2325 9300
rect 2365 9260 2375 9300
rect 2315 9240 2375 9260
rect 2315 9200 2325 9240
rect 2365 9200 2375 9240
rect 2315 9175 2375 9200
rect 2315 9135 2325 9175
rect 2365 9135 2375 9175
rect 2315 9105 2375 9135
rect 2315 9065 2325 9105
rect 2365 9065 2375 9105
rect 2315 9035 2375 9065
rect 2315 8995 2325 9035
rect 2365 8995 2375 9035
rect 2315 8965 2375 8995
rect 2315 8925 2325 8965
rect 2365 8925 2375 8965
rect 2315 8900 2375 8925
rect 2315 8860 2325 8900
rect 2365 8860 2375 8900
rect 2315 8840 2375 8860
rect 2315 8800 2325 8840
rect 2365 8800 2375 8840
rect 2315 8775 2375 8800
rect 2315 8735 2325 8775
rect 2365 8735 2375 8775
rect 2315 8705 2375 8735
rect 2315 8665 2325 8705
rect 2365 8665 2375 8705
rect 2315 8635 2375 8665
rect 2315 8595 2325 8635
rect 2365 8595 2375 8635
rect 2315 8565 2375 8595
rect 2315 8525 2325 8565
rect 2365 8525 2375 8565
rect 2315 8500 2375 8525
rect 2315 8460 2325 8500
rect 2365 8460 2375 8500
rect 2315 8440 2375 8460
rect 2315 8400 2325 8440
rect 2365 8400 2375 8440
rect 2315 8375 2375 8400
rect 2315 8335 2325 8375
rect 2365 8335 2375 8375
rect 2315 8305 2375 8335
rect 2315 8265 2325 8305
rect 2365 8265 2375 8305
rect 2315 8235 2375 8265
rect 2315 8195 2325 8235
rect 2365 8195 2375 8235
rect 2315 8165 2375 8195
rect 2315 8125 2325 8165
rect 2365 8125 2375 8165
rect 2315 8100 2375 8125
rect 2315 8060 2325 8100
rect 2365 8060 2375 8100
rect 2315 8040 2375 8060
rect 2315 8000 2325 8040
rect 2365 8000 2375 8040
rect 2315 7975 2375 8000
rect 2315 7935 2325 7975
rect 2365 7935 2375 7975
rect 2315 7905 2375 7935
rect 2315 7865 2325 7905
rect 2365 7865 2375 7905
rect 2315 7835 2375 7865
rect 2315 7795 2325 7835
rect 2365 7795 2375 7835
rect 2315 7765 2375 7795
rect 2315 7725 2325 7765
rect 2365 7725 2375 7765
rect 2315 7700 2375 7725
rect 2315 7660 2325 7700
rect 2365 7660 2375 7700
rect 2315 7640 2375 7660
rect 2315 7600 2325 7640
rect 2365 7600 2375 7640
rect 2315 7575 2375 7600
rect 2315 7535 2325 7575
rect 2365 7535 2375 7575
rect 2315 7505 2375 7535
rect 2315 7465 2325 7505
rect 2365 7465 2375 7505
rect 2315 7435 2375 7465
rect 2315 7395 2325 7435
rect 2365 7395 2375 7435
rect 2315 7365 2375 7395
rect 2315 7325 2325 7365
rect 2365 7325 2375 7365
rect 2315 7300 2375 7325
rect 2315 7260 2325 7300
rect 2365 7260 2375 7300
rect 2315 7240 2375 7260
rect 2315 7200 2325 7240
rect 2365 7200 2375 7240
rect 2315 7175 2375 7200
rect 2315 7135 2325 7175
rect 2365 7135 2375 7175
rect 2315 7105 2375 7135
rect 2315 7065 2325 7105
rect 2365 7065 2375 7105
rect 2315 7035 2375 7065
rect 2315 6995 2325 7035
rect 2365 6995 2375 7035
rect 2315 6965 2375 6995
rect 2315 6925 2325 6965
rect 2365 6925 2375 6965
rect 2315 6900 2375 6925
rect 2315 6860 2325 6900
rect 2365 6860 2375 6900
rect 2315 6840 2375 6860
rect 2315 6800 2325 6840
rect 2365 6800 2375 6840
rect 2315 6775 2375 6800
rect 2315 6735 2325 6775
rect 2365 6735 2375 6775
rect 2315 6705 2375 6735
rect 2315 6665 2325 6705
rect 2365 6665 2375 6705
rect 2315 6635 2375 6665
rect 2315 6595 2325 6635
rect 2365 6595 2375 6635
rect 2315 6565 2375 6595
rect 2315 6525 2325 6565
rect 2365 6525 2375 6565
rect 2315 6500 2375 6525
rect 2315 6460 2325 6500
rect 2365 6460 2375 6500
rect 2315 6450 2375 6460
rect 3165 9640 3285 9650
rect 3165 9600 3175 9640
rect 3215 9600 3235 9640
rect 3275 9600 3285 9640
rect 3165 9575 3285 9600
rect 3165 9535 3175 9575
rect 3215 9535 3235 9575
rect 3275 9535 3285 9575
rect 3165 9505 3285 9535
rect 3165 9465 3175 9505
rect 3215 9465 3235 9505
rect 3275 9465 3285 9505
rect 3165 9435 3285 9465
rect 3165 9395 3175 9435
rect 3215 9395 3235 9435
rect 3275 9395 3285 9435
rect 3165 9365 3285 9395
rect 3165 9325 3175 9365
rect 3215 9325 3235 9365
rect 3275 9325 3285 9365
rect 3165 9300 3285 9325
rect 3165 9260 3175 9300
rect 3215 9260 3235 9300
rect 3275 9260 3285 9300
rect 3165 9240 3285 9260
rect 3165 9200 3175 9240
rect 3215 9200 3235 9240
rect 3275 9200 3285 9240
rect 3165 9175 3285 9200
rect 3165 9135 3175 9175
rect 3215 9135 3235 9175
rect 3275 9135 3285 9175
rect 3165 9105 3285 9135
rect 3165 9065 3175 9105
rect 3215 9065 3235 9105
rect 3275 9065 3285 9105
rect 3165 9035 3285 9065
rect 3165 8995 3175 9035
rect 3215 8995 3235 9035
rect 3275 8995 3285 9035
rect 3165 8965 3285 8995
rect 3165 8925 3175 8965
rect 3215 8925 3235 8965
rect 3275 8925 3285 8965
rect 3165 8900 3285 8925
rect 3165 8860 3175 8900
rect 3215 8860 3235 8900
rect 3275 8860 3285 8900
rect 3165 8840 3285 8860
rect 3165 8800 3175 8840
rect 3215 8800 3235 8840
rect 3275 8800 3285 8840
rect 3165 8775 3285 8800
rect 3165 8735 3175 8775
rect 3215 8735 3235 8775
rect 3275 8735 3285 8775
rect 3165 8705 3285 8735
rect 3165 8665 3175 8705
rect 3215 8665 3235 8705
rect 3275 8665 3285 8705
rect 3165 8635 3285 8665
rect 3165 8595 3175 8635
rect 3215 8595 3235 8635
rect 3275 8595 3285 8635
rect 3165 8565 3285 8595
rect 3165 8525 3175 8565
rect 3215 8525 3235 8565
rect 3275 8525 3285 8565
rect 3165 8500 3285 8525
rect 3165 8460 3175 8500
rect 3215 8460 3235 8500
rect 3275 8460 3285 8500
rect 3165 8440 3285 8460
rect 3165 8400 3175 8440
rect 3215 8400 3235 8440
rect 3275 8400 3285 8440
rect 3165 8375 3285 8400
rect 3165 8335 3175 8375
rect 3215 8335 3235 8375
rect 3275 8335 3285 8375
rect 3165 8305 3285 8335
rect 3165 8265 3175 8305
rect 3215 8265 3235 8305
rect 3275 8265 3285 8305
rect 3165 8235 3285 8265
rect 3165 8195 3175 8235
rect 3215 8195 3235 8235
rect 3275 8195 3285 8235
rect 3165 8165 3285 8195
rect 3165 8125 3175 8165
rect 3215 8125 3235 8165
rect 3275 8125 3285 8165
rect 3165 8100 3285 8125
rect 3165 8060 3175 8100
rect 3215 8060 3235 8100
rect 3275 8060 3285 8100
rect 3165 8040 3285 8060
rect 3165 8000 3175 8040
rect 3215 8000 3235 8040
rect 3275 8000 3285 8040
rect 3165 7975 3285 8000
rect 3165 7935 3175 7975
rect 3215 7935 3235 7975
rect 3275 7935 3285 7975
rect 3165 7905 3285 7935
rect 3165 7865 3175 7905
rect 3215 7865 3235 7905
rect 3275 7865 3285 7905
rect 3165 7835 3285 7865
rect 3165 7795 3175 7835
rect 3215 7795 3235 7835
rect 3275 7795 3285 7835
rect 3165 7765 3285 7795
rect 3165 7725 3175 7765
rect 3215 7725 3235 7765
rect 3275 7725 3285 7765
rect 3165 7700 3285 7725
rect 3165 7660 3175 7700
rect 3215 7660 3235 7700
rect 3275 7660 3285 7700
rect 3165 7640 3285 7660
rect 3165 7600 3175 7640
rect 3215 7600 3235 7640
rect 3275 7600 3285 7640
rect 3165 7575 3285 7600
rect 3165 7535 3175 7575
rect 3215 7535 3235 7575
rect 3275 7535 3285 7575
rect 3165 7505 3285 7535
rect 3165 7465 3175 7505
rect 3215 7465 3235 7505
rect 3275 7465 3285 7505
rect 3165 7435 3285 7465
rect 3165 7395 3175 7435
rect 3215 7395 3235 7435
rect 3275 7395 3285 7435
rect 3165 7365 3285 7395
rect 3165 7325 3175 7365
rect 3215 7325 3235 7365
rect 3275 7325 3285 7365
rect 3165 7300 3285 7325
rect 3165 7260 3175 7300
rect 3215 7260 3235 7300
rect 3275 7260 3285 7300
rect 3165 7240 3285 7260
rect 3165 7200 3175 7240
rect 3215 7200 3235 7240
rect 3275 7200 3285 7240
rect 3165 7175 3285 7200
rect 3165 7135 3175 7175
rect 3215 7135 3235 7175
rect 3275 7135 3285 7175
rect 3165 7105 3285 7135
rect 3165 7065 3175 7105
rect 3215 7065 3235 7105
rect 3275 7065 3285 7105
rect 3165 7035 3285 7065
rect 3165 6995 3175 7035
rect 3215 6995 3235 7035
rect 3275 6995 3285 7035
rect 3165 6965 3285 6995
rect 3165 6925 3175 6965
rect 3215 6925 3235 6965
rect 3275 6925 3285 6965
rect 3165 6900 3285 6925
rect 3165 6860 3175 6900
rect 3215 6860 3235 6900
rect 3275 6860 3285 6900
rect 3165 6840 3285 6860
rect 3165 6800 3175 6840
rect 3215 6800 3235 6840
rect 3275 6800 3285 6840
rect 3165 6775 3285 6800
rect 3165 6735 3175 6775
rect 3215 6735 3235 6775
rect 3275 6735 3285 6775
rect 3165 6705 3285 6735
rect 3165 6665 3175 6705
rect 3215 6665 3235 6705
rect 3275 6665 3285 6705
rect 3165 6635 3285 6665
rect 3165 6595 3175 6635
rect 3215 6595 3235 6635
rect 3275 6595 3285 6635
rect 3165 6565 3285 6595
rect 3165 6525 3175 6565
rect 3215 6525 3235 6565
rect 3275 6525 3285 6565
rect 3165 6500 3285 6525
rect 3165 6460 3175 6500
rect 3215 6460 3235 6500
rect 3275 6460 3285 6500
rect 3165 6450 3285 6460
rect 3335 9640 3395 9650
rect 3335 9600 3345 9640
rect 3385 9600 3395 9640
rect 3335 9575 3395 9600
rect 3335 9535 3345 9575
rect 3385 9535 3395 9575
rect 3335 9505 3395 9535
rect 3335 9465 3345 9505
rect 3385 9465 3395 9505
rect 3335 9435 3395 9465
rect 3335 9395 3345 9435
rect 3385 9395 3395 9435
rect 3335 9365 3395 9395
rect 3335 9325 3345 9365
rect 3385 9325 3395 9365
rect 3335 9300 3395 9325
rect 3335 9260 3345 9300
rect 3385 9260 3395 9300
rect 3335 9240 3395 9260
rect 3335 9200 3345 9240
rect 3385 9200 3395 9240
rect 3335 9175 3395 9200
rect 3335 9135 3345 9175
rect 3385 9135 3395 9175
rect 3335 9105 3395 9135
rect 3335 9065 3345 9105
rect 3385 9065 3395 9105
rect 3335 9035 3395 9065
rect 3335 8995 3345 9035
rect 3385 8995 3395 9035
rect 3335 8965 3395 8995
rect 3335 8925 3345 8965
rect 3385 8925 3395 8965
rect 3335 8900 3395 8925
rect 3335 8860 3345 8900
rect 3385 8860 3395 8900
rect 3335 8840 3395 8860
rect 3335 8800 3345 8840
rect 3385 8800 3395 8840
rect 3335 8775 3395 8800
rect 3335 8735 3345 8775
rect 3385 8735 3395 8775
rect 3335 8705 3395 8735
rect 3335 8665 3345 8705
rect 3385 8665 3395 8705
rect 3335 8635 3395 8665
rect 3335 8595 3345 8635
rect 3385 8595 3395 8635
rect 3335 8565 3395 8595
rect 3335 8525 3345 8565
rect 3385 8525 3395 8565
rect 3335 8500 3395 8525
rect 3335 8460 3345 8500
rect 3385 8460 3395 8500
rect 3335 8440 3395 8460
rect 3335 8400 3345 8440
rect 3385 8400 3395 8440
rect 3335 8375 3395 8400
rect 3335 8335 3345 8375
rect 3385 8335 3395 8375
rect 3335 8305 3395 8335
rect 3335 8265 3345 8305
rect 3385 8265 3395 8305
rect 3335 8235 3395 8265
rect 3335 8195 3345 8235
rect 3385 8195 3395 8235
rect 3335 8165 3395 8195
rect 3335 8125 3345 8165
rect 3385 8125 3395 8165
rect 3335 8100 3395 8125
rect 3335 8060 3345 8100
rect 3385 8060 3395 8100
rect 3335 8040 3395 8060
rect 3335 8000 3345 8040
rect 3385 8000 3395 8040
rect 3335 7975 3395 8000
rect 3335 7935 3345 7975
rect 3385 7935 3395 7975
rect 3335 7905 3395 7935
rect 3335 7865 3345 7905
rect 3385 7865 3395 7905
rect 3335 7835 3395 7865
rect 3335 7795 3345 7835
rect 3385 7795 3395 7835
rect 3335 7765 3395 7795
rect 3335 7725 3345 7765
rect 3385 7725 3395 7765
rect 3335 7700 3395 7725
rect 3335 7660 3345 7700
rect 3385 7660 3395 7700
rect 3335 7640 3395 7660
rect 3335 7600 3345 7640
rect 3385 7600 3395 7640
rect 3335 7575 3395 7600
rect 3335 7535 3345 7575
rect 3385 7535 3395 7575
rect 3335 7505 3395 7535
rect 3335 7465 3345 7505
rect 3385 7465 3395 7505
rect 3335 7435 3395 7465
rect 3335 7395 3345 7435
rect 3385 7395 3395 7435
rect 3335 7365 3395 7395
rect 3335 7325 3345 7365
rect 3385 7325 3395 7365
rect 3335 7300 3395 7325
rect 3335 7260 3345 7300
rect 3385 7260 3395 7300
rect 3335 7240 3395 7260
rect 3335 7200 3345 7240
rect 3385 7200 3395 7240
rect 3335 7175 3395 7200
rect 3335 7135 3345 7175
rect 3385 7135 3395 7175
rect 3335 7105 3395 7135
rect 3335 7065 3345 7105
rect 3385 7065 3395 7105
rect 3335 7035 3395 7065
rect 3335 6995 3345 7035
rect 3385 6995 3395 7035
rect 3335 6965 3395 6995
rect 3335 6925 3345 6965
rect 3385 6925 3395 6965
rect 3335 6900 3395 6925
rect 3335 6860 3345 6900
rect 3385 6860 3395 6900
rect 3335 6840 3395 6860
rect 3335 6800 3345 6840
rect 3385 6800 3395 6840
rect 3335 6775 3395 6800
rect 3335 6735 3345 6775
rect 3385 6735 3395 6775
rect 3335 6705 3395 6735
rect 3335 6665 3345 6705
rect 3385 6665 3395 6705
rect 3335 6635 3395 6665
rect 3335 6595 3345 6635
rect 3385 6595 3395 6635
rect 3335 6565 3395 6595
rect 3335 6525 3345 6565
rect 3385 6525 3395 6565
rect 3335 6500 3395 6525
rect 3335 6460 3345 6500
rect 3385 6460 3395 6500
rect 3335 6450 3395 6460
rect 6620 9640 6680 9650
rect 6620 9600 6630 9640
rect 6670 9600 6680 9640
rect 6620 9575 6680 9600
rect 6620 9535 6630 9575
rect 6670 9535 6680 9575
rect 6620 9505 6680 9535
rect 6620 9465 6630 9505
rect 6670 9465 6680 9505
rect 6620 9435 6680 9465
rect 6620 9395 6630 9435
rect 6670 9395 6680 9435
rect 6620 9365 6680 9395
rect 6620 9325 6630 9365
rect 6670 9325 6680 9365
rect 6620 9300 6680 9325
rect 6620 9260 6630 9300
rect 6670 9260 6680 9300
rect 6620 9240 6680 9260
rect 6620 9200 6630 9240
rect 6670 9200 6680 9240
rect 6620 9175 6680 9200
rect 6620 9135 6630 9175
rect 6670 9135 6680 9175
rect 6620 9105 6680 9135
rect 6620 9065 6630 9105
rect 6670 9065 6680 9105
rect 6620 9035 6680 9065
rect 6620 8995 6630 9035
rect 6670 8995 6680 9035
rect 6620 8965 6680 8995
rect 6620 8925 6630 8965
rect 6670 8925 6680 8965
rect 6620 8900 6680 8925
rect 6620 8860 6630 8900
rect 6670 8860 6680 8900
rect 6620 8840 6680 8860
rect 6620 8800 6630 8840
rect 6670 8800 6680 8840
rect 6620 8775 6680 8800
rect 6620 8735 6630 8775
rect 6670 8735 6680 8775
rect 6620 8705 6680 8735
rect 6620 8665 6630 8705
rect 6670 8665 6680 8705
rect 6620 8635 6680 8665
rect 6620 8595 6630 8635
rect 6670 8595 6680 8635
rect 6620 8565 6680 8595
rect 6620 8525 6630 8565
rect 6670 8525 6680 8565
rect 6620 8500 6680 8525
rect 6620 8460 6630 8500
rect 6670 8460 6680 8500
rect 6620 8440 6680 8460
rect 6620 8400 6630 8440
rect 6670 8400 6680 8440
rect 6620 8375 6680 8400
rect 6620 8335 6630 8375
rect 6670 8335 6680 8375
rect 6620 8305 6680 8335
rect 6620 8265 6630 8305
rect 6670 8265 6680 8305
rect 6620 8235 6680 8265
rect 6620 8195 6630 8235
rect 6670 8195 6680 8235
rect 6620 8165 6680 8195
rect 6620 8125 6630 8165
rect 6670 8125 6680 8165
rect 6620 8100 6680 8125
rect 6620 8060 6630 8100
rect 6670 8060 6680 8100
rect 6620 8040 6680 8060
rect 6620 8000 6630 8040
rect 6670 8000 6680 8040
rect 6620 7975 6680 8000
rect 6620 7935 6630 7975
rect 6670 7935 6680 7975
rect 6620 7905 6680 7935
rect 6620 7865 6630 7905
rect 6670 7865 6680 7905
rect 6620 7835 6680 7865
rect 6620 7795 6630 7835
rect 6670 7795 6680 7835
rect 6620 7765 6680 7795
rect 6620 7725 6630 7765
rect 6670 7725 6680 7765
rect 6620 7700 6680 7725
rect 6620 7660 6630 7700
rect 6670 7660 6680 7700
rect 6620 7640 6680 7660
rect 6620 7600 6630 7640
rect 6670 7600 6680 7640
rect 6620 7575 6680 7600
rect 6620 7535 6630 7575
rect 6670 7535 6680 7575
rect 6620 7505 6680 7535
rect 6620 7465 6630 7505
rect 6670 7465 6680 7505
rect 6620 7435 6680 7465
rect 6620 7395 6630 7435
rect 6670 7395 6680 7435
rect 6620 7365 6680 7395
rect 6620 7325 6630 7365
rect 6670 7325 6680 7365
rect 6620 7300 6680 7325
rect 6620 7260 6630 7300
rect 6670 7260 6680 7300
rect 6620 7240 6680 7260
rect 6620 7200 6630 7240
rect 6670 7200 6680 7240
rect 6620 7175 6680 7200
rect 6620 7135 6630 7175
rect 6670 7135 6680 7175
rect 6620 7105 6680 7135
rect 6620 7065 6630 7105
rect 6670 7065 6680 7105
rect 6620 7035 6680 7065
rect 6620 6995 6630 7035
rect 6670 6995 6680 7035
rect 6620 6965 6680 6995
rect 6620 6925 6630 6965
rect 6670 6925 6680 6965
rect 6620 6900 6680 6925
rect 6620 6860 6630 6900
rect 6670 6860 6680 6900
rect 6620 6840 6680 6860
rect 6620 6800 6630 6840
rect 6670 6800 6680 6840
rect 6620 6775 6680 6800
rect 6620 6735 6630 6775
rect 6670 6735 6680 6775
rect 6620 6705 6680 6735
rect 6620 6665 6630 6705
rect 6670 6665 6680 6705
rect 6620 6635 6680 6665
rect 6620 6595 6630 6635
rect 6670 6595 6680 6635
rect 6620 6565 6680 6595
rect 6620 6525 6630 6565
rect 6670 6525 6680 6565
rect 6620 6500 6680 6525
rect 6620 6460 6630 6500
rect 6670 6460 6680 6500
rect 6620 6450 6680 6460
rect 7260 9640 7320 9650
rect 7260 9600 7270 9640
rect 7310 9600 7320 9640
rect 7260 9575 7320 9600
rect 7260 9535 7270 9575
rect 7310 9535 7320 9575
rect 7260 9505 7320 9535
rect 7260 9465 7270 9505
rect 7310 9465 7320 9505
rect 7260 9435 7320 9465
rect 7260 9395 7270 9435
rect 7310 9395 7320 9435
rect 7260 9365 7320 9395
rect 7260 9325 7270 9365
rect 7310 9325 7320 9365
rect 7260 9300 7320 9325
rect 7260 9260 7270 9300
rect 7310 9260 7320 9300
rect 7260 9240 7320 9260
rect 7260 9200 7270 9240
rect 7310 9200 7320 9240
rect 7260 9175 7320 9200
rect 7260 9135 7270 9175
rect 7310 9135 7320 9175
rect 7260 9105 7320 9135
rect 7260 9065 7270 9105
rect 7310 9065 7320 9105
rect 7260 9035 7320 9065
rect 7260 8995 7270 9035
rect 7310 8995 7320 9035
rect 7260 8965 7320 8995
rect 7260 8925 7270 8965
rect 7310 8925 7320 8965
rect 7260 8900 7320 8925
rect 7260 8860 7270 8900
rect 7310 8860 7320 8900
rect 7260 8840 7320 8860
rect 7260 8800 7270 8840
rect 7310 8800 7320 8840
rect 7260 8775 7320 8800
rect 7260 8735 7270 8775
rect 7310 8735 7320 8775
rect 7260 8705 7320 8735
rect 7260 8665 7270 8705
rect 7310 8665 7320 8705
rect 7260 8635 7320 8665
rect 7260 8595 7270 8635
rect 7310 8595 7320 8635
rect 7260 8565 7320 8595
rect 7260 8525 7270 8565
rect 7310 8525 7320 8565
rect 7260 8500 7320 8525
rect 7260 8460 7270 8500
rect 7310 8460 7320 8500
rect 7260 8440 7320 8460
rect 7260 8400 7270 8440
rect 7310 8400 7320 8440
rect 7260 8375 7320 8400
rect 7260 8335 7270 8375
rect 7310 8335 7320 8375
rect 7260 8305 7320 8335
rect 7260 8265 7270 8305
rect 7310 8265 7320 8305
rect 7260 8235 7320 8265
rect 7260 8195 7270 8235
rect 7310 8195 7320 8235
rect 7260 8165 7320 8195
rect 7260 8125 7270 8165
rect 7310 8125 7320 8165
rect 7260 8100 7320 8125
rect 7260 8060 7270 8100
rect 7310 8060 7320 8100
rect 7260 8040 7320 8060
rect 7260 8000 7270 8040
rect 7310 8000 7320 8040
rect 7260 7975 7320 8000
rect 7260 7935 7270 7975
rect 7310 7935 7320 7975
rect 7260 7905 7320 7935
rect 7260 7865 7270 7905
rect 7310 7865 7320 7905
rect 7260 7835 7320 7865
rect 7260 7795 7270 7835
rect 7310 7795 7320 7835
rect 7260 7765 7320 7795
rect 7260 7725 7270 7765
rect 7310 7725 7320 7765
rect 7260 7700 7320 7725
rect 7260 7660 7270 7700
rect 7310 7660 7320 7700
rect 7260 7640 7320 7660
rect 7260 7600 7270 7640
rect 7310 7600 7320 7640
rect 7260 7575 7320 7600
rect 7260 7535 7270 7575
rect 7310 7535 7320 7575
rect 7260 7505 7320 7535
rect 7260 7465 7270 7505
rect 7310 7465 7320 7505
rect 7260 7435 7320 7465
rect 7260 7395 7270 7435
rect 7310 7395 7320 7435
rect 7260 7365 7320 7395
rect 7260 7325 7270 7365
rect 7310 7325 7320 7365
rect 7260 7300 7320 7325
rect 7260 7260 7270 7300
rect 7310 7260 7320 7300
rect 7260 7240 7320 7260
rect 7260 7200 7270 7240
rect 7310 7200 7320 7240
rect 7260 7175 7320 7200
rect 7260 7135 7270 7175
rect 7310 7135 7320 7175
rect 7260 7105 7320 7135
rect 7260 7065 7270 7105
rect 7310 7065 7320 7105
rect 7260 7035 7320 7065
rect 7260 6995 7270 7035
rect 7310 6995 7320 7035
rect 7260 6965 7320 6995
rect 7260 6925 7270 6965
rect 7310 6925 7320 6965
rect 7260 6900 7320 6925
rect 7260 6860 7270 6900
rect 7310 6860 7320 6900
rect 7260 6840 7320 6860
rect 7260 6800 7270 6840
rect 7310 6800 7320 6840
rect 7260 6775 7320 6800
rect 7260 6735 7270 6775
rect 7310 6735 7320 6775
rect 7260 6705 7320 6735
rect 7260 6665 7270 6705
rect 7310 6665 7320 6705
rect 7260 6635 7320 6665
rect 7260 6595 7270 6635
rect 7310 6595 7320 6635
rect 7260 6565 7320 6595
rect 7260 6525 7270 6565
rect 7310 6525 7320 6565
rect 7260 6500 7320 6525
rect 7260 6460 7270 6500
rect 7310 6460 7320 6500
rect 7260 6450 7320 6460
rect 7960 9640 8020 9650
rect 7960 9600 7970 9640
rect 8010 9600 8020 9640
rect 7960 9575 8020 9600
rect 7960 9535 7970 9575
rect 8010 9535 8020 9575
rect 7960 9505 8020 9535
rect 7960 9465 7970 9505
rect 8010 9465 8020 9505
rect 7960 9435 8020 9465
rect 7960 9395 7970 9435
rect 8010 9395 8020 9435
rect 7960 9365 8020 9395
rect 7960 9325 7970 9365
rect 8010 9325 8020 9365
rect 7960 9300 8020 9325
rect 7960 9260 7970 9300
rect 8010 9260 8020 9300
rect 7960 9240 8020 9260
rect 7960 9200 7970 9240
rect 8010 9200 8020 9240
rect 7960 9175 8020 9200
rect 7960 9135 7970 9175
rect 8010 9135 8020 9175
rect 7960 9105 8020 9135
rect 7960 9065 7970 9105
rect 8010 9065 8020 9105
rect 7960 9035 8020 9065
rect 7960 8995 7970 9035
rect 8010 8995 8020 9035
rect 7960 8965 8020 8995
rect 7960 8925 7970 8965
rect 8010 8925 8020 8965
rect 7960 8900 8020 8925
rect 7960 8860 7970 8900
rect 8010 8860 8020 8900
rect 7960 8840 8020 8860
rect 7960 8800 7970 8840
rect 8010 8800 8020 8840
rect 7960 8775 8020 8800
rect 7960 8735 7970 8775
rect 8010 8735 8020 8775
rect 7960 8705 8020 8735
rect 7960 8665 7970 8705
rect 8010 8665 8020 8705
rect 7960 8635 8020 8665
rect 7960 8595 7970 8635
rect 8010 8595 8020 8635
rect 7960 8565 8020 8595
rect 7960 8525 7970 8565
rect 8010 8525 8020 8565
rect 7960 8500 8020 8525
rect 7960 8460 7970 8500
rect 8010 8460 8020 8500
rect 7960 8440 8020 8460
rect 7960 8400 7970 8440
rect 8010 8400 8020 8440
rect 7960 8375 8020 8400
rect 7960 8335 7970 8375
rect 8010 8335 8020 8375
rect 7960 8305 8020 8335
rect 7960 8265 7970 8305
rect 8010 8265 8020 8305
rect 7960 8235 8020 8265
rect 7960 8195 7970 8235
rect 8010 8195 8020 8235
rect 7960 8165 8020 8195
rect 7960 8125 7970 8165
rect 8010 8125 8020 8165
rect 7960 8100 8020 8125
rect 7960 8060 7970 8100
rect 8010 8060 8020 8100
rect 7960 8040 8020 8060
rect 7960 8000 7970 8040
rect 8010 8000 8020 8040
rect 7960 7975 8020 8000
rect 7960 7935 7970 7975
rect 8010 7935 8020 7975
rect 7960 7905 8020 7935
rect 7960 7865 7970 7905
rect 8010 7865 8020 7905
rect 7960 7835 8020 7865
rect 7960 7795 7970 7835
rect 8010 7795 8020 7835
rect 7960 7765 8020 7795
rect 7960 7725 7970 7765
rect 8010 7725 8020 7765
rect 7960 7700 8020 7725
rect 7960 7660 7970 7700
rect 8010 7660 8020 7700
rect 7960 7640 8020 7660
rect 7960 7600 7970 7640
rect 8010 7600 8020 7640
rect 7960 7575 8020 7600
rect 7960 7535 7970 7575
rect 8010 7535 8020 7575
rect 7960 7505 8020 7535
rect 7960 7465 7970 7505
rect 8010 7465 8020 7505
rect 7960 7435 8020 7465
rect 7960 7395 7970 7435
rect 8010 7395 8020 7435
rect 7960 7365 8020 7395
rect 7960 7325 7970 7365
rect 8010 7325 8020 7365
rect 7960 7300 8020 7325
rect 7960 7260 7970 7300
rect 8010 7260 8020 7300
rect 7960 7240 8020 7260
rect 7960 7200 7970 7240
rect 8010 7200 8020 7240
rect 7960 7175 8020 7200
rect 7960 7135 7970 7175
rect 8010 7135 8020 7175
rect 7960 7105 8020 7135
rect 7960 7065 7970 7105
rect 8010 7065 8020 7105
rect 7960 7035 8020 7065
rect 7960 6995 7970 7035
rect 8010 6995 8020 7035
rect 7960 6965 8020 6995
rect 7960 6925 7970 6965
rect 8010 6925 8020 6965
rect 7960 6900 8020 6925
rect 7960 6860 7970 6900
rect 8010 6860 8020 6900
rect 7960 6840 8020 6860
rect 7960 6800 7970 6840
rect 8010 6800 8020 6840
rect 7960 6775 8020 6800
rect 7960 6735 7970 6775
rect 8010 6735 8020 6775
rect 7960 6705 8020 6735
rect 7960 6665 7970 6705
rect 8010 6665 8020 6705
rect 7960 6635 8020 6665
rect 7960 6595 7970 6635
rect 8010 6595 8020 6635
rect 7960 6565 8020 6595
rect 7960 6525 7970 6565
rect 8010 6525 8020 6565
rect 7960 6500 8020 6525
rect 7960 6460 7970 6500
rect 8010 6460 8020 6500
rect 7960 6450 8020 6460
rect 8310 9640 8370 9650
rect 8310 9600 8320 9640
rect 8360 9600 8370 9640
rect 8310 9575 8370 9600
rect 8310 9535 8320 9575
rect 8360 9535 8370 9575
rect 8310 9505 8370 9535
rect 8310 9465 8320 9505
rect 8360 9465 8370 9505
rect 8310 9435 8370 9465
rect 8310 9395 8320 9435
rect 8360 9395 8370 9435
rect 8310 9365 8370 9395
rect 8310 9325 8320 9365
rect 8360 9325 8370 9365
rect 8310 9300 8370 9325
rect 8310 9260 8320 9300
rect 8360 9260 8370 9300
rect 8310 9240 8370 9260
rect 8310 9200 8320 9240
rect 8360 9200 8370 9240
rect 8310 9175 8370 9200
rect 8310 9135 8320 9175
rect 8360 9135 8370 9175
rect 8310 9105 8370 9135
rect 8310 9065 8320 9105
rect 8360 9065 8370 9105
rect 8310 9035 8370 9065
rect 8310 8995 8320 9035
rect 8360 8995 8370 9035
rect 8310 8965 8370 8995
rect 8310 8925 8320 8965
rect 8360 8925 8370 8965
rect 8310 8900 8370 8925
rect 8310 8860 8320 8900
rect 8360 8860 8370 8900
rect 8310 8840 8370 8860
rect 8310 8800 8320 8840
rect 8360 8800 8370 8840
rect 8310 8775 8370 8800
rect 8310 8735 8320 8775
rect 8360 8735 8370 8775
rect 8310 8705 8370 8735
rect 8310 8665 8320 8705
rect 8360 8665 8370 8705
rect 8310 8635 8370 8665
rect 8310 8595 8320 8635
rect 8360 8595 8370 8635
rect 8310 8565 8370 8595
rect 8310 8525 8320 8565
rect 8360 8525 8370 8565
rect 8310 8500 8370 8525
rect 8310 8460 8320 8500
rect 8360 8460 8370 8500
rect 8310 8440 8370 8460
rect 8310 8400 8320 8440
rect 8360 8400 8370 8440
rect 8310 8375 8370 8400
rect 8310 8335 8320 8375
rect 8360 8335 8370 8375
rect 8310 8305 8370 8335
rect 8310 8265 8320 8305
rect 8360 8265 8370 8305
rect 8310 8235 8370 8265
rect 8310 8195 8320 8235
rect 8360 8195 8370 8235
rect 8310 8165 8370 8195
rect 8310 8125 8320 8165
rect 8360 8125 8370 8165
rect 8310 8100 8370 8125
rect 8310 8060 8320 8100
rect 8360 8060 8370 8100
rect 8310 8040 8370 8060
rect 8310 8000 8320 8040
rect 8360 8000 8370 8040
rect 8310 7975 8370 8000
rect 8310 7935 8320 7975
rect 8360 7935 8370 7975
rect 8310 7905 8370 7935
rect 8310 7865 8320 7905
rect 8360 7865 8370 7905
rect 8310 7835 8370 7865
rect 8310 7795 8320 7835
rect 8360 7795 8370 7835
rect 8310 7765 8370 7795
rect 8310 7725 8320 7765
rect 8360 7725 8370 7765
rect 8310 7700 8370 7725
rect 8310 7660 8320 7700
rect 8360 7660 8370 7700
rect 8310 7640 8370 7660
rect 8310 7600 8320 7640
rect 8360 7600 8370 7640
rect 8310 7575 8370 7600
rect 8310 7535 8320 7575
rect 8360 7535 8370 7575
rect 8310 7505 8370 7535
rect 8310 7465 8320 7505
rect 8360 7465 8370 7505
rect 8310 7435 8370 7465
rect 8310 7395 8320 7435
rect 8360 7395 8370 7435
rect 8310 7365 8370 7395
rect 8310 7325 8320 7365
rect 8360 7325 8370 7365
rect 8310 7300 8370 7325
rect 8310 7260 8320 7300
rect 8360 7260 8370 7300
rect 8310 7240 8370 7260
rect 8310 7200 8320 7240
rect 8360 7200 8370 7240
rect 8310 7175 8370 7200
rect 8310 7135 8320 7175
rect 8360 7135 8370 7175
rect 8310 7105 8370 7135
rect 8310 7065 8320 7105
rect 8360 7065 8370 7105
rect 8310 7035 8370 7065
rect 8310 6995 8320 7035
rect 8360 6995 8370 7035
rect 8310 6965 8370 6995
rect 8310 6925 8320 6965
rect 8360 6925 8370 6965
rect 8310 6900 8370 6925
rect 8310 6860 8320 6900
rect 8360 6860 8370 6900
rect 8310 6840 8370 6860
rect 8310 6800 8320 6840
rect 8360 6800 8370 6840
rect 8310 6775 8370 6800
rect 8310 6735 8320 6775
rect 8360 6735 8370 6775
rect 8310 6705 8370 6735
rect 8310 6665 8320 6705
rect 8360 6665 8370 6705
rect 8310 6635 8370 6665
rect 8310 6595 8320 6635
rect 8360 6595 8370 6635
rect 8310 6565 8370 6595
rect 8310 6525 8320 6565
rect 8360 6525 8370 6565
rect 8310 6500 8370 6525
rect 8310 6460 8320 6500
rect 8360 6460 8370 6500
rect 8310 6450 8370 6460
rect 8660 9640 8720 9650
rect 8660 9600 8670 9640
rect 8710 9600 8720 9640
rect 8660 9575 8720 9600
rect 8660 9535 8670 9575
rect 8710 9535 8720 9575
rect 8660 9505 8720 9535
rect 8660 9465 8670 9505
rect 8710 9465 8720 9505
rect 8660 9435 8720 9465
rect 8660 9395 8670 9435
rect 8710 9395 8720 9435
rect 8660 9365 8720 9395
rect 8660 9325 8670 9365
rect 8710 9325 8720 9365
rect 8660 9300 8720 9325
rect 8660 9260 8670 9300
rect 8710 9260 8720 9300
rect 8660 9240 8720 9260
rect 8660 9200 8670 9240
rect 8710 9200 8720 9240
rect 8660 9175 8720 9200
rect 8660 9135 8670 9175
rect 8710 9135 8720 9175
rect 8660 9105 8720 9135
rect 8660 9065 8670 9105
rect 8710 9065 8720 9105
rect 8660 9035 8720 9065
rect 8660 8995 8670 9035
rect 8710 8995 8720 9035
rect 8660 8965 8720 8995
rect 8660 8925 8670 8965
rect 8710 8925 8720 8965
rect 8660 8900 8720 8925
rect 8660 8860 8670 8900
rect 8710 8860 8720 8900
rect 8660 8840 8720 8860
rect 8660 8800 8670 8840
rect 8710 8800 8720 8840
rect 8660 8775 8720 8800
rect 8660 8735 8670 8775
rect 8710 8735 8720 8775
rect 8660 8705 8720 8735
rect 8660 8665 8670 8705
rect 8710 8665 8720 8705
rect 8660 8635 8720 8665
rect 8660 8595 8670 8635
rect 8710 8595 8720 8635
rect 8660 8565 8720 8595
rect 8660 8525 8670 8565
rect 8710 8525 8720 8565
rect 8660 8500 8720 8525
rect 8660 8460 8670 8500
rect 8710 8460 8720 8500
rect 8660 8440 8720 8460
rect 8660 8400 8670 8440
rect 8710 8400 8720 8440
rect 8660 8375 8720 8400
rect 8660 8335 8670 8375
rect 8710 8335 8720 8375
rect 8660 8305 8720 8335
rect 8660 8265 8670 8305
rect 8710 8265 8720 8305
rect 8660 8235 8720 8265
rect 8660 8195 8670 8235
rect 8710 8195 8720 8235
rect 8660 8165 8720 8195
rect 8660 8125 8670 8165
rect 8710 8125 8720 8165
rect 8660 8100 8720 8125
rect 8660 8060 8670 8100
rect 8710 8060 8720 8100
rect 8660 8040 8720 8060
rect 8660 8000 8670 8040
rect 8710 8000 8720 8040
rect 8660 7975 8720 8000
rect 8660 7935 8670 7975
rect 8710 7935 8720 7975
rect 8660 7905 8720 7935
rect 8660 7865 8670 7905
rect 8710 7865 8720 7905
rect 8660 7835 8720 7865
rect 8660 7795 8670 7835
rect 8710 7795 8720 7835
rect 8660 7765 8720 7795
rect 8660 7725 8670 7765
rect 8710 7725 8720 7765
rect 8660 7700 8720 7725
rect 8660 7660 8670 7700
rect 8710 7660 8720 7700
rect 8660 7640 8720 7660
rect 8660 7600 8670 7640
rect 8710 7600 8720 7640
rect 8660 7575 8720 7600
rect 8660 7535 8670 7575
rect 8710 7535 8720 7575
rect 8660 7505 8720 7535
rect 8660 7465 8670 7505
rect 8710 7465 8720 7505
rect 8660 7435 8720 7465
rect 8660 7395 8670 7435
rect 8710 7395 8720 7435
rect 8660 7365 8720 7395
rect 8660 7325 8670 7365
rect 8710 7325 8720 7365
rect 8660 7300 8720 7325
rect 8660 7260 8670 7300
rect 8710 7260 8720 7300
rect 8660 7240 8720 7260
rect 8660 7200 8670 7240
rect 8710 7200 8720 7240
rect 8660 7175 8720 7200
rect 8660 7135 8670 7175
rect 8710 7135 8720 7175
rect 8660 7105 8720 7135
rect 8660 7065 8670 7105
rect 8710 7065 8720 7105
rect 8660 7035 8720 7065
rect 8660 6995 8670 7035
rect 8710 6995 8720 7035
rect 8660 6965 8720 6995
rect 8660 6925 8670 6965
rect 8710 6925 8720 6965
rect 8660 6900 8720 6925
rect 8660 6860 8670 6900
rect 8710 6860 8720 6900
rect 8660 6840 8720 6860
rect 8660 6800 8670 6840
rect 8710 6800 8720 6840
rect 8660 6775 8720 6800
rect 8660 6735 8670 6775
rect 8710 6735 8720 6775
rect 8660 6705 8720 6735
rect 8660 6665 8670 6705
rect 8710 6665 8720 6705
rect 8660 6635 8720 6665
rect 8660 6595 8670 6635
rect 8710 6595 8720 6635
rect 8660 6565 8720 6595
rect 8660 6525 8670 6565
rect 8710 6525 8720 6565
rect 8660 6500 8720 6525
rect 8660 6460 8670 6500
rect 8710 6460 8720 6500
rect 8660 6450 8720 6460
rect 9010 9640 9070 9650
rect 9010 9600 9020 9640
rect 9060 9600 9070 9640
rect 9010 9575 9070 9600
rect 9010 9535 9020 9575
rect 9060 9535 9070 9575
rect 9010 9505 9070 9535
rect 9010 9465 9020 9505
rect 9060 9465 9070 9505
rect 9010 9435 9070 9465
rect 9010 9395 9020 9435
rect 9060 9395 9070 9435
rect 9010 9365 9070 9395
rect 9010 9325 9020 9365
rect 9060 9325 9070 9365
rect 9010 9300 9070 9325
rect 9010 9260 9020 9300
rect 9060 9260 9070 9300
rect 9010 9240 9070 9260
rect 9010 9200 9020 9240
rect 9060 9200 9070 9240
rect 9010 9175 9070 9200
rect 9010 9135 9020 9175
rect 9060 9135 9070 9175
rect 9010 9105 9070 9135
rect 9010 9065 9020 9105
rect 9060 9065 9070 9105
rect 9010 9035 9070 9065
rect 9010 8995 9020 9035
rect 9060 8995 9070 9035
rect 9010 8965 9070 8995
rect 9010 8925 9020 8965
rect 9060 8925 9070 8965
rect 9010 8900 9070 8925
rect 9010 8860 9020 8900
rect 9060 8860 9070 8900
rect 9010 8840 9070 8860
rect 9010 8800 9020 8840
rect 9060 8800 9070 8840
rect 9010 8775 9070 8800
rect 9010 8735 9020 8775
rect 9060 8735 9070 8775
rect 9010 8705 9070 8735
rect 9010 8665 9020 8705
rect 9060 8665 9070 8705
rect 9010 8635 9070 8665
rect 9010 8595 9020 8635
rect 9060 8595 9070 8635
rect 9010 8565 9070 8595
rect 9010 8525 9020 8565
rect 9060 8525 9070 8565
rect 9010 8500 9070 8525
rect 9010 8460 9020 8500
rect 9060 8460 9070 8500
rect 9010 8440 9070 8460
rect 9010 8400 9020 8440
rect 9060 8400 9070 8440
rect 9010 8375 9070 8400
rect 9010 8335 9020 8375
rect 9060 8335 9070 8375
rect 9010 8305 9070 8335
rect 9010 8265 9020 8305
rect 9060 8265 9070 8305
rect 9010 8235 9070 8265
rect 9010 8195 9020 8235
rect 9060 8195 9070 8235
rect 9010 8165 9070 8195
rect 9010 8125 9020 8165
rect 9060 8125 9070 8165
rect 9010 8100 9070 8125
rect 9010 8060 9020 8100
rect 9060 8060 9070 8100
rect 9010 8040 9070 8060
rect 9010 8000 9020 8040
rect 9060 8000 9070 8040
rect 9010 7975 9070 8000
rect 9010 7935 9020 7975
rect 9060 7935 9070 7975
rect 9010 7905 9070 7935
rect 9010 7865 9020 7905
rect 9060 7865 9070 7905
rect 9010 7835 9070 7865
rect 9010 7795 9020 7835
rect 9060 7795 9070 7835
rect 9010 7765 9070 7795
rect 9010 7725 9020 7765
rect 9060 7725 9070 7765
rect 9010 7700 9070 7725
rect 9010 7660 9020 7700
rect 9060 7660 9070 7700
rect 9010 7640 9070 7660
rect 9010 7600 9020 7640
rect 9060 7600 9070 7640
rect 9010 7575 9070 7600
rect 9010 7535 9020 7575
rect 9060 7535 9070 7575
rect 9010 7505 9070 7535
rect 9010 7465 9020 7505
rect 9060 7465 9070 7505
rect 9010 7435 9070 7465
rect 9010 7395 9020 7435
rect 9060 7395 9070 7435
rect 9010 7365 9070 7395
rect 9010 7325 9020 7365
rect 9060 7325 9070 7365
rect 9010 7300 9070 7325
rect 9010 7260 9020 7300
rect 9060 7260 9070 7300
rect 9010 7240 9070 7260
rect 9010 7200 9020 7240
rect 9060 7200 9070 7240
rect 9010 7175 9070 7200
rect 9010 7135 9020 7175
rect 9060 7135 9070 7175
rect 9010 7105 9070 7135
rect 9010 7065 9020 7105
rect 9060 7065 9070 7105
rect 9010 7035 9070 7065
rect 9010 6995 9020 7035
rect 9060 6995 9070 7035
rect 9010 6965 9070 6995
rect 9010 6925 9020 6965
rect 9060 6925 9070 6965
rect 9010 6900 9070 6925
rect 9010 6860 9020 6900
rect 9060 6860 9070 6900
rect 9010 6840 9070 6860
rect 9010 6800 9020 6840
rect 9060 6800 9070 6840
rect 9010 6775 9070 6800
rect 9010 6735 9020 6775
rect 9060 6735 9070 6775
rect 9010 6705 9070 6735
rect 9010 6665 9020 6705
rect 9060 6665 9070 6705
rect 9010 6635 9070 6665
rect 9010 6595 9020 6635
rect 9060 6595 9070 6635
rect 9010 6565 9070 6595
rect 9010 6525 9020 6565
rect 9060 6525 9070 6565
rect 9010 6500 9070 6525
rect 9010 6460 9020 6500
rect 9060 6460 9070 6500
rect 9010 6450 9070 6460
rect 12890 9615 16090 17760
rect 12890 9565 12925 9615
rect 12975 9565 13020 9615
rect 13070 9565 13115 9615
rect 13165 9565 13215 9615
rect 13265 9565 13315 9615
rect 13365 9565 13415 9615
rect 13465 9565 13510 9615
rect 13560 9565 13605 9615
rect 13655 9565 13725 9615
rect 13775 9565 13820 9615
rect 13870 9565 13915 9615
rect 13965 9565 14015 9615
rect 14065 9565 14115 9615
rect 14165 9565 14215 9615
rect 14265 9565 14310 9615
rect 14360 9565 14405 9615
rect 14455 9565 14525 9615
rect 14575 9565 14620 9615
rect 14670 9565 14715 9615
rect 14765 9565 14815 9615
rect 14865 9565 14915 9615
rect 14965 9565 15015 9615
rect 15065 9565 15110 9615
rect 15160 9565 15205 9615
rect 15255 9565 15325 9615
rect 15375 9565 15420 9615
rect 15470 9565 15515 9615
rect 15565 9565 15615 9615
rect 15665 9565 15715 9615
rect 15765 9565 15815 9615
rect 15865 9565 15910 9615
rect 15960 9565 16005 9615
rect 16055 9565 16090 9615
rect 12890 9525 16090 9565
rect 12890 9475 12925 9525
rect 12975 9475 13020 9525
rect 13070 9475 13115 9525
rect 13165 9475 13215 9525
rect 13265 9475 13315 9525
rect 13365 9475 13415 9525
rect 13465 9475 13510 9525
rect 13560 9475 13605 9525
rect 13655 9475 13725 9525
rect 13775 9475 13820 9525
rect 13870 9475 13915 9525
rect 13965 9475 14015 9525
rect 14065 9475 14115 9525
rect 14165 9475 14215 9525
rect 14265 9475 14310 9525
rect 14360 9475 14405 9525
rect 14455 9475 14525 9525
rect 14575 9475 14620 9525
rect 14670 9475 14715 9525
rect 14765 9475 14815 9525
rect 14865 9475 14915 9525
rect 14965 9475 15015 9525
rect 15065 9475 15110 9525
rect 15160 9475 15205 9525
rect 15255 9475 15325 9525
rect 15375 9475 15420 9525
rect 15470 9475 15515 9525
rect 15565 9475 15615 9525
rect 15665 9475 15715 9525
rect 15765 9475 15815 9525
rect 15865 9475 15910 9525
rect 15960 9475 16005 9525
rect 16055 9475 16090 9525
rect 12890 9425 16090 9475
rect 12890 9375 12925 9425
rect 12975 9375 13020 9425
rect 13070 9375 13115 9425
rect 13165 9375 13215 9425
rect 13265 9375 13315 9425
rect 13365 9375 13415 9425
rect 13465 9375 13510 9425
rect 13560 9375 13605 9425
rect 13655 9375 13725 9425
rect 13775 9375 13820 9425
rect 13870 9375 13915 9425
rect 13965 9375 14015 9425
rect 14065 9375 14115 9425
rect 14165 9375 14215 9425
rect 14265 9375 14310 9425
rect 14360 9375 14405 9425
rect 14455 9375 14525 9425
rect 14575 9375 14620 9425
rect 14670 9375 14715 9425
rect 14765 9375 14815 9425
rect 14865 9375 14915 9425
rect 14965 9375 15015 9425
rect 15065 9375 15110 9425
rect 15160 9375 15205 9425
rect 15255 9375 15325 9425
rect 15375 9375 15420 9425
rect 15470 9375 15515 9425
rect 15565 9375 15615 9425
rect 15665 9375 15715 9425
rect 15765 9375 15815 9425
rect 15865 9375 15910 9425
rect 15960 9375 16005 9425
rect 16055 9375 16090 9425
rect 12890 9335 16090 9375
rect 12890 9285 12925 9335
rect 12975 9285 13020 9335
rect 13070 9285 13115 9335
rect 13165 9285 13215 9335
rect 13265 9285 13315 9335
rect 13365 9285 13415 9335
rect 13465 9285 13510 9335
rect 13560 9285 13605 9335
rect 13655 9285 13725 9335
rect 13775 9285 13820 9335
rect 13870 9285 13915 9335
rect 13965 9285 14015 9335
rect 14065 9285 14115 9335
rect 14165 9285 14215 9335
rect 14265 9285 14310 9335
rect 14360 9285 14405 9335
rect 14455 9285 14525 9335
rect 14575 9285 14620 9335
rect 14670 9285 14715 9335
rect 14765 9285 14815 9335
rect 14865 9285 14915 9335
rect 14965 9285 15015 9335
rect 15065 9285 15110 9335
rect 15160 9285 15205 9335
rect 15255 9285 15325 9335
rect 15375 9285 15420 9335
rect 15470 9285 15515 9335
rect 15565 9285 15615 9335
rect 15665 9285 15715 9335
rect 15765 9285 15815 9335
rect 15865 9285 15910 9335
rect 15960 9285 16005 9335
rect 16055 9285 16090 9335
rect 12890 9215 16090 9285
rect 12890 9165 12925 9215
rect 12975 9165 13020 9215
rect 13070 9165 13115 9215
rect 13165 9165 13215 9215
rect 13265 9165 13315 9215
rect 13365 9165 13415 9215
rect 13465 9165 13510 9215
rect 13560 9165 13605 9215
rect 13655 9165 13725 9215
rect 13775 9165 13820 9215
rect 13870 9165 13915 9215
rect 13965 9165 14015 9215
rect 14065 9165 14115 9215
rect 14165 9165 14215 9215
rect 14265 9165 14310 9215
rect 14360 9165 14405 9215
rect 14455 9165 14525 9215
rect 14575 9165 14620 9215
rect 14670 9165 14715 9215
rect 14765 9165 14815 9215
rect 14865 9165 14915 9215
rect 14965 9165 15015 9215
rect 15065 9165 15110 9215
rect 15160 9165 15205 9215
rect 15255 9165 15325 9215
rect 15375 9165 15420 9215
rect 15470 9165 15515 9215
rect 15565 9165 15615 9215
rect 15665 9165 15715 9215
rect 15765 9165 15815 9215
rect 15865 9165 15910 9215
rect 15960 9165 16005 9215
rect 16055 9165 16090 9215
rect 12890 9125 16090 9165
rect 12890 9075 12925 9125
rect 12975 9075 13020 9125
rect 13070 9075 13115 9125
rect 13165 9075 13215 9125
rect 13265 9075 13315 9125
rect 13365 9075 13415 9125
rect 13465 9075 13510 9125
rect 13560 9075 13605 9125
rect 13655 9075 13725 9125
rect 13775 9075 13820 9125
rect 13870 9075 13915 9125
rect 13965 9075 14015 9125
rect 14065 9075 14115 9125
rect 14165 9075 14215 9125
rect 14265 9075 14310 9125
rect 14360 9075 14405 9125
rect 14455 9075 14525 9125
rect 14575 9075 14620 9125
rect 14670 9075 14715 9125
rect 14765 9075 14815 9125
rect 14865 9075 14915 9125
rect 14965 9075 15015 9125
rect 15065 9075 15110 9125
rect 15160 9075 15205 9125
rect 15255 9075 15325 9125
rect 15375 9075 15420 9125
rect 15470 9075 15515 9125
rect 15565 9075 15615 9125
rect 15665 9075 15715 9125
rect 15765 9075 15815 9125
rect 15865 9075 15910 9125
rect 15960 9075 16005 9125
rect 16055 9075 16090 9125
rect 12890 9025 16090 9075
rect 12890 8975 12925 9025
rect 12975 8975 13020 9025
rect 13070 8975 13115 9025
rect 13165 8975 13215 9025
rect 13265 8975 13315 9025
rect 13365 8975 13415 9025
rect 13465 8975 13510 9025
rect 13560 8975 13605 9025
rect 13655 8975 13725 9025
rect 13775 8975 13820 9025
rect 13870 8975 13915 9025
rect 13965 8975 14015 9025
rect 14065 8975 14115 9025
rect 14165 8975 14215 9025
rect 14265 8975 14310 9025
rect 14360 8975 14405 9025
rect 14455 8975 14525 9025
rect 14575 8975 14620 9025
rect 14670 8975 14715 9025
rect 14765 8975 14815 9025
rect 14865 8975 14915 9025
rect 14965 8975 15015 9025
rect 15065 8975 15110 9025
rect 15160 8975 15205 9025
rect 15255 8975 15325 9025
rect 15375 8975 15420 9025
rect 15470 8975 15515 9025
rect 15565 8975 15615 9025
rect 15665 8975 15715 9025
rect 15765 8975 15815 9025
rect 15865 8975 15910 9025
rect 15960 8975 16005 9025
rect 16055 8975 16090 9025
rect 12890 8935 16090 8975
rect 12890 8885 12925 8935
rect 12975 8885 13020 8935
rect 13070 8885 13115 8935
rect 13165 8885 13215 8935
rect 13265 8885 13315 8935
rect 13365 8885 13415 8935
rect 13465 8885 13510 8935
rect 13560 8885 13605 8935
rect 13655 8885 13725 8935
rect 13775 8885 13820 8935
rect 13870 8885 13915 8935
rect 13965 8885 14015 8935
rect 14065 8885 14115 8935
rect 14165 8885 14215 8935
rect 14265 8885 14310 8935
rect 14360 8885 14405 8935
rect 14455 8885 14525 8935
rect 14575 8885 14620 8935
rect 14670 8885 14715 8935
rect 14765 8885 14815 8935
rect 14865 8885 14915 8935
rect 14965 8885 15015 8935
rect 15065 8885 15110 8935
rect 15160 8885 15205 8935
rect 15255 8885 15325 8935
rect 15375 8885 15420 8935
rect 15470 8885 15515 8935
rect 15565 8885 15615 8935
rect 15665 8885 15715 8935
rect 15765 8885 15815 8935
rect 15865 8885 15910 8935
rect 15960 8885 16005 8935
rect 16055 8885 16090 8935
rect 12890 8815 16090 8885
rect 12890 8765 12925 8815
rect 12975 8765 13020 8815
rect 13070 8765 13115 8815
rect 13165 8765 13215 8815
rect 13265 8765 13315 8815
rect 13365 8765 13415 8815
rect 13465 8765 13510 8815
rect 13560 8765 13605 8815
rect 13655 8765 13725 8815
rect 13775 8765 13820 8815
rect 13870 8765 13915 8815
rect 13965 8765 14015 8815
rect 14065 8765 14115 8815
rect 14165 8765 14215 8815
rect 14265 8765 14310 8815
rect 14360 8765 14405 8815
rect 14455 8765 14525 8815
rect 14575 8765 14620 8815
rect 14670 8765 14715 8815
rect 14765 8765 14815 8815
rect 14865 8765 14915 8815
rect 14965 8765 15015 8815
rect 15065 8765 15110 8815
rect 15160 8765 15205 8815
rect 15255 8765 15325 8815
rect 15375 8765 15420 8815
rect 15470 8765 15515 8815
rect 15565 8765 15615 8815
rect 15665 8765 15715 8815
rect 15765 8765 15815 8815
rect 15865 8765 15910 8815
rect 15960 8765 16005 8815
rect 16055 8765 16090 8815
rect 12890 8725 16090 8765
rect 12890 8675 12925 8725
rect 12975 8675 13020 8725
rect 13070 8675 13115 8725
rect 13165 8675 13215 8725
rect 13265 8675 13315 8725
rect 13365 8675 13415 8725
rect 13465 8675 13510 8725
rect 13560 8675 13605 8725
rect 13655 8675 13725 8725
rect 13775 8675 13820 8725
rect 13870 8675 13915 8725
rect 13965 8675 14015 8725
rect 14065 8675 14115 8725
rect 14165 8675 14215 8725
rect 14265 8675 14310 8725
rect 14360 8675 14405 8725
rect 14455 8675 14525 8725
rect 14575 8675 14620 8725
rect 14670 8675 14715 8725
rect 14765 8675 14815 8725
rect 14865 8675 14915 8725
rect 14965 8675 15015 8725
rect 15065 8675 15110 8725
rect 15160 8675 15205 8725
rect 15255 8675 15325 8725
rect 15375 8675 15420 8725
rect 15470 8675 15515 8725
rect 15565 8675 15615 8725
rect 15665 8675 15715 8725
rect 15765 8675 15815 8725
rect 15865 8675 15910 8725
rect 15960 8675 16005 8725
rect 16055 8675 16090 8725
rect 12890 8625 16090 8675
rect 12890 8575 12925 8625
rect 12975 8575 13020 8625
rect 13070 8575 13115 8625
rect 13165 8575 13215 8625
rect 13265 8575 13315 8625
rect 13365 8575 13415 8625
rect 13465 8575 13510 8625
rect 13560 8575 13605 8625
rect 13655 8575 13725 8625
rect 13775 8575 13820 8625
rect 13870 8575 13915 8625
rect 13965 8575 14015 8625
rect 14065 8575 14115 8625
rect 14165 8575 14215 8625
rect 14265 8575 14310 8625
rect 14360 8575 14405 8625
rect 14455 8575 14525 8625
rect 14575 8575 14620 8625
rect 14670 8575 14715 8625
rect 14765 8575 14815 8625
rect 14865 8575 14915 8625
rect 14965 8575 15015 8625
rect 15065 8575 15110 8625
rect 15160 8575 15205 8625
rect 15255 8575 15325 8625
rect 15375 8575 15420 8625
rect 15470 8575 15515 8625
rect 15565 8575 15615 8625
rect 15665 8575 15715 8625
rect 15765 8575 15815 8625
rect 15865 8575 15910 8625
rect 15960 8575 16005 8625
rect 16055 8575 16090 8625
rect 12890 8535 16090 8575
rect 12890 8485 12925 8535
rect 12975 8485 13020 8535
rect 13070 8485 13115 8535
rect 13165 8485 13215 8535
rect 13265 8485 13315 8535
rect 13365 8485 13415 8535
rect 13465 8485 13510 8535
rect 13560 8485 13605 8535
rect 13655 8485 13725 8535
rect 13775 8485 13820 8535
rect 13870 8485 13915 8535
rect 13965 8485 14015 8535
rect 14065 8485 14115 8535
rect 14165 8485 14215 8535
rect 14265 8485 14310 8535
rect 14360 8485 14405 8535
rect 14455 8485 14525 8535
rect 14575 8485 14620 8535
rect 14670 8485 14715 8535
rect 14765 8485 14815 8535
rect 14865 8485 14915 8535
rect 14965 8485 15015 8535
rect 15065 8485 15110 8535
rect 15160 8485 15205 8535
rect 15255 8485 15325 8535
rect 15375 8485 15420 8535
rect 15470 8485 15515 8535
rect 15565 8485 15615 8535
rect 15665 8485 15715 8535
rect 15765 8485 15815 8535
rect 15865 8485 15910 8535
rect 15960 8485 16005 8535
rect 16055 8485 16090 8535
rect 12890 8415 16090 8485
rect 12890 8365 12925 8415
rect 12975 8365 13020 8415
rect 13070 8365 13115 8415
rect 13165 8365 13215 8415
rect 13265 8365 13315 8415
rect 13365 8365 13415 8415
rect 13465 8365 13510 8415
rect 13560 8365 13605 8415
rect 13655 8365 13725 8415
rect 13775 8365 13820 8415
rect 13870 8365 13915 8415
rect 13965 8365 14015 8415
rect 14065 8365 14115 8415
rect 14165 8365 14215 8415
rect 14265 8365 14310 8415
rect 14360 8365 14405 8415
rect 14455 8365 14525 8415
rect 14575 8365 14620 8415
rect 14670 8365 14715 8415
rect 14765 8365 14815 8415
rect 14865 8365 14915 8415
rect 14965 8365 15015 8415
rect 15065 8365 15110 8415
rect 15160 8365 15205 8415
rect 15255 8365 15325 8415
rect 15375 8365 15420 8415
rect 15470 8365 15515 8415
rect 15565 8365 15615 8415
rect 15665 8365 15715 8415
rect 15765 8365 15815 8415
rect 15865 8365 15910 8415
rect 15960 8365 16005 8415
rect 16055 8365 16090 8415
rect 12890 8325 16090 8365
rect 12890 8275 12925 8325
rect 12975 8275 13020 8325
rect 13070 8275 13115 8325
rect 13165 8275 13215 8325
rect 13265 8275 13315 8325
rect 13365 8275 13415 8325
rect 13465 8275 13510 8325
rect 13560 8275 13605 8325
rect 13655 8275 13725 8325
rect 13775 8275 13820 8325
rect 13870 8275 13915 8325
rect 13965 8275 14015 8325
rect 14065 8275 14115 8325
rect 14165 8275 14215 8325
rect 14265 8275 14310 8325
rect 14360 8275 14405 8325
rect 14455 8275 14525 8325
rect 14575 8275 14620 8325
rect 14670 8275 14715 8325
rect 14765 8275 14815 8325
rect 14865 8275 14915 8325
rect 14965 8275 15015 8325
rect 15065 8275 15110 8325
rect 15160 8275 15205 8325
rect 15255 8275 15325 8325
rect 15375 8275 15420 8325
rect 15470 8275 15515 8325
rect 15565 8275 15615 8325
rect 15665 8275 15715 8325
rect 15765 8275 15815 8325
rect 15865 8275 15910 8325
rect 15960 8275 16005 8325
rect 16055 8275 16090 8325
rect 12890 8225 16090 8275
rect 12890 8175 12925 8225
rect 12975 8175 13020 8225
rect 13070 8175 13115 8225
rect 13165 8175 13215 8225
rect 13265 8175 13315 8225
rect 13365 8175 13415 8225
rect 13465 8175 13510 8225
rect 13560 8175 13605 8225
rect 13655 8175 13725 8225
rect 13775 8175 13820 8225
rect 13870 8175 13915 8225
rect 13965 8175 14015 8225
rect 14065 8175 14115 8225
rect 14165 8175 14215 8225
rect 14265 8175 14310 8225
rect 14360 8175 14405 8225
rect 14455 8175 14525 8225
rect 14575 8175 14620 8225
rect 14670 8175 14715 8225
rect 14765 8175 14815 8225
rect 14865 8175 14915 8225
rect 14965 8175 15015 8225
rect 15065 8175 15110 8225
rect 15160 8175 15205 8225
rect 15255 8175 15325 8225
rect 15375 8175 15420 8225
rect 15470 8175 15515 8225
rect 15565 8175 15615 8225
rect 15665 8175 15715 8225
rect 15765 8175 15815 8225
rect 15865 8175 15910 8225
rect 15960 8175 16005 8225
rect 16055 8175 16090 8225
rect 12890 8135 16090 8175
rect 12890 8085 12925 8135
rect 12975 8085 13020 8135
rect 13070 8085 13115 8135
rect 13165 8085 13215 8135
rect 13265 8085 13315 8135
rect 13365 8085 13415 8135
rect 13465 8085 13510 8135
rect 13560 8085 13605 8135
rect 13655 8085 13725 8135
rect 13775 8085 13820 8135
rect 13870 8085 13915 8135
rect 13965 8085 14015 8135
rect 14065 8085 14115 8135
rect 14165 8085 14215 8135
rect 14265 8085 14310 8135
rect 14360 8085 14405 8135
rect 14455 8085 14525 8135
rect 14575 8085 14620 8135
rect 14670 8085 14715 8135
rect 14765 8085 14815 8135
rect 14865 8085 14915 8135
rect 14965 8085 15015 8135
rect 15065 8085 15110 8135
rect 15160 8085 15205 8135
rect 15255 8085 15325 8135
rect 15375 8085 15420 8135
rect 15470 8085 15515 8135
rect 15565 8085 15615 8135
rect 15665 8085 15715 8135
rect 15765 8085 15815 8135
rect 15865 8085 15910 8135
rect 15960 8085 16005 8135
rect 16055 8085 16090 8135
rect 12890 8015 16090 8085
rect 12890 7965 12925 8015
rect 12975 7965 13020 8015
rect 13070 7965 13115 8015
rect 13165 7965 13215 8015
rect 13265 7965 13315 8015
rect 13365 7965 13415 8015
rect 13465 7965 13510 8015
rect 13560 7965 13605 8015
rect 13655 7965 13725 8015
rect 13775 7965 13820 8015
rect 13870 7965 13915 8015
rect 13965 7965 14015 8015
rect 14065 7965 14115 8015
rect 14165 7965 14215 8015
rect 14265 7965 14310 8015
rect 14360 7965 14405 8015
rect 14455 7965 14525 8015
rect 14575 7965 14620 8015
rect 14670 7965 14715 8015
rect 14765 7965 14815 8015
rect 14865 7965 14915 8015
rect 14965 7965 15015 8015
rect 15065 7965 15110 8015
rect 15160 7965 15205 8015
rect 15255 7965 15325 8015
rect 15375 7965 15420 8015
rect 15470 7965 15515 8015
rect 15565 7965 15615 8015
rect 15665 7965 15715 8015
rect 15765 7965 15815 8015
rect 15865 7965 15910 8015
rect 15960 7965 16005 8015
rect 16055 7965 16090 8015
rect 12890 7925 16090 7965
rect 12890 7875 12925 7925
rect 12975 7875 13020 7925
rect 13070 7875 13115 7925
rect 13165 7875 13215 7925
rect 13265 7875 13315 7925
rect 13365 7875 13415 7925
rect 13465 7875 13510 7925
rect 13560 7875 13605 7925
rect 13655 7875 13725 7925
rect 13775 7875 13820 7925
rect 13870 7875 13915 7925
rect 13965 7875 14015 7925
rect 14065 7875 14115 7925
rect 14165 7875 14215 7925
rect 14265 7875 14310 7925
rect 14360 7875 14405 7925
rect 14455 7875 14525 7925
rect 14575 7875 14620 7925
rect 14670 7875 14715 7925
rect 14765 7875 14815 7925
rect 14865 7875 14915 7925
rect 14965 7875 15015 7925
rect 15065 7875 15110 7925
rect 15160 7875 15205 7925
rect 15255 7875 15325 7925
rect 15375 7875 15420 7925
rect 15470 7875 15515 7925
rect 15565 7875 15615 7925
rect 15665 7875 15715 7925
rect 15765 7875 15815 7925
rect 15865 7875 15910 7925
rect 15960 7875 16005 7925
rect 16055 7875 16090 7925
rect 12890 7825 16090 7875
rect 12890 7775 12925 7825
rect 12975 7775 13020 7825
rect 13070 7775 13115 7825
rect 13165 7775 13215 7825
rect 13265 7775 13315 7825
rect 13365 7775 13415 7825
rect 13465 7775 13510 7825
rect 13560 7775 13605 7825
rect 13655 7775 13725 7825
rect 13775 7775 13820 7825
rect 13870 7775 13915 7825
rect 13965 7775 14015 7825
rect 14065 7775 14115 7825
rect 14165 7775 14215 7825
rect 14265 7775 14310 7825
rect 14360 7775 14405 7825
rect 14455 7775 14525 7825
rect 14575 7775 14620 7825
rect 14670 7775 14715 7825
rect 14765 7775 14815 7825
rect 14865 7775 14915 7825
rect 14965 7775 15015 7825
rect 15065 7775 15110 7825
rect 15160 7775 15205 7825
rect 15255 7775 15325 7825
rect 15375 7775 15420 7825
rect 15470 7775 15515 7825
rect 15565 7775 15615 7825
rect 15665 7775 15715 7825
rect 15765 7775 15815 7825
rect 15865 7775 15910 7825
rect 15960 7775 16005 7825
rect 16055 7775 16090 7825
rect 12890 7735 16090 7775
rect 12890 7685 12925 7735
rect 12975 7685 13020 7735
rect 13070 7685 13115 7735
rect 13165 7685 13215 7735
rect 13265 7685 13315 7735
rect 13365 7685 13415 7735
rect 13465 7685 13510 7735
rect 13560 7685 13605 7735
rect 13655 7685 13725 7735
rect 13775 7685 13820 7735
rect 13870 7685 13915 7735
rect 13965 7685 14015 7735
rect 14065 7685 14115 7735
rect 14165 7685 14215 7735
rect 14265 7685 14310 7735
rect 14360 7685 14405 7735
rect 14455 7685 14525 7735
rect 14575 7685 14620 7735
rect 14670 7685 14715 7735
rect 14765 7685 14815 7735
rect 14865 7685 14915 7735
rect 14965 7685 15015 7735
rect 15065 7685 15110 7735
rect 15160 7685 15205 7735
rect 15255 7685 15325 7735
rect 15375 7685 15420 7735
rect 15470 7685 15515 7735
rect 15565 7685 15615 7735
rect 15665 7685 15715 7735
rect 15765 7685 15815 7735
rect 15865 7685 15910 7735
rect 15960 7685 16005 7735
rect 16055 7685 16090 7735
rect 12890 7615 16090 7685
rect 12890 7565 12925 7615
rect 12975 7565 13020 7615
rect 13070 7565 13115 7615
rect 13165 7565 13215 7615
rect 13265 7565 13315 7615
rect 13365 7565 13415 7615
rect 13465 7565 13510 7615
rect 13560 7565 13605 7615
rect 13655 7565 13725 7615
rect 13775 7565 13820 7615
rect 13870 7565 13915 7615
rect 13965 7565 14015 7615
rect 14065 7565 14115 7615
rect 14165 7565 14215 7615
rect 14265 7565 14310 7615
rect 14360 7565 14405 7615
rect 14455 7565 14525 7615
rect 14575 7565 14620 7615
rect 14670 7565 14715 7615
rect 14765 7565 14815 7615
rect 14865 7565 14915 7615
rect 14965 7565 15015 7615
rect 15065 7565 15110 7615
rect 15160 7565 15205 7615
rect 15255 7565 15325 7615
rect 15375 7565 15420 7615
rect 15470 7565 15515 7615
rect 15565 7565 15615 7615
rect 15665 7565 15715 7615
rect 15765 7565 15815 7615
rect 15865 7565 15910 7615
rect 15960 7565 16005 7615
rect 16055 7565 16090 7615
rect 12890 7525 16090 7565
rect 12890 7475 12925 7525
rect 12975 7475 13020 7525
rect 13070 7475 13115 7525
rect 13165 7475 13215 7525
rect 13265 7475 13315 7525
rect 13365 7475 13415 7525
rect 13465 7475 13510 7525
rect 13560 7475 13605 7525
rect 13655 7475 13725 7525
rect 13775 7475 13820 7525
rect 13870 7475 13915 7525
rect 13965 7475 14015 7525
rect 14065 7475 14115 7525
rect 14165 7475 14215 7525
rect 14265 7475 14310 7525
rect 14360 7475 14405 7525
rect 14455 7475 14525 7525
rect 14575 7475 14620 7525
rect 14670 7475 14715 7525
rect 14765 7475 14815 7525
rect 14865 7475 14915 7525
rect 14965 7475 15015 7525
rect 15065 7475 15110 7525
rect 15160 7475 15205 7525
rect 15255 7475 15325 7525
rect 15375 7475 15420 7525
rect 15470 7475 15515 7525
rect 15565 7475 15615 7525
rect 15665 7475 15715 7525
rect 15765 7475 15815 7525
rect 15865 7475 15910 7525
rect 15960 7475 16005 7525
rect 16055 7475 16090 7525
rect 12890 7425 16090 7475
rect 12890 7375 12925 7425
rect 12975 7375 13020 7425
rect 13070 7375 13115 7425
rect 13165 7375 13215 7425
rect 13265 7375 13315 7425
rect 13365 7375 13415 7425
rect 13465 7375 13510 7425
rect 13560 7375 13605 7425
rect 13655 7375 13725 7425
rect 13775 7375 13820 7425
rect 13870 7375 13915 7425
rect 13965 7375 14015 7425
rect 14065 7375 14115 7425
rect 14165 7375 14215 7425
rect 14265 7375 14310 7425
rect 14360 7375 14405 7425
rect 14455 7375 14525 7425
rect 14575 7375 14620 7425
rect 14670 7375 14715 7425
rect 14765 7375 14815 7425
rect 14865 7375 14915 7425
rect 14965 7375 15015 7425
rect 15065 7375 15110 7425
rect 15160 7375 15205 7425
rect 15255 7375 15325 7425
rect 15375 7375 15420 7425
rect 15470 7375 15515 7425
rect 15565 7375 15615 7425
rect 15665 7375 15715 7425
rect 15765 7375 15815 7425
rect 15865 7375 15910 7425
rect 15960 7375 16005 7425
rect 16055 7375 16090 7425
rect 12890 7335 16090 7375
rect 12890 7285 12925 7335
rect 12975 7285 13020 7335
rect 13070 7285 13115 7335
rect 13165 7285 13215 7335
rect 13265 7285 13315 7335
rect 13365 7285 13415 7335
rect 13465 7285 13510 7335
rect 13560 7285 13605 7335
rect 13655 7285 13725 7335
rect 13775 7285 13820 7335
rect 13870 7285 13915 7335
rect 13965 7285 14015 7335
rect 14065 7285 14115 7335
rect 14165 7285 14215 7335
rect 14265 7285 14310 7335
rect 14360 7285 14405 7335
rect 14455 7285 14525 7335
rect 14575 7285 14620 7335
rect 14670 7285 14715 7335
rect 14765 7285 14815 7335
rect 14865 7285 14915 7335
rect 14965 7285 15015 7335
rect 15065 7285 15110 7335
rect 15160 7285 15205 7335
rect 15255 7285 15325 7335
rect 15375 7285 15420 7335
rect 15470 7285 15515 7335
rect 15565 7285 15615 7335
rect 15665 7285 15715 7335
rect 15765 7285 15815 7335
rect 15865 7285 15910 7335
rect 15960 7285 16005 7335
rect 16055 7285 16090 7335
rect 12890 7215 16090 7285
rect 12890 7165 12925 7215
rect 12975 7165 13020 7215
rect 13070 7165 13115 7215
rect 13165 7165 13215 7215
rect 13265 7165 13315 7215
rect 13365 7165 13415 7215
rect 13465 7165 13510 7215
rect 13560 7165 13605 7215
rect 13655 7165 13725 7215
rect 13775 7165 13820 7215
rect 13870 7165 13915 7215
rect 13965 7165 14015 7215
rect 14065 7165 14115 7215
rect 14165 7165 14215 7215
rect 14265 7165 14310 7215
rect 14360 7165 14405 7215
rect 14455 7165 14525 7215
rect 14575 7165 14620 7215
rect 14670 7165 14715 7215
rect 14765 7165 14815 7215
rect 14865 7165 14915 7215
rect 14965 7165 15015 7215
rect 15065 7165 15110 7215
rect 15160 7165 15205 7215
rect 15255 7165 15325 7215
rect 15375 7165 15420 7215
rect 15470 7165 15515 7215
rect 15565 7165 15615 7215
rect 15665 7165 15715 7215
rect 15765 7165 15815 7215
rect 15865 7165 15910 7215
rect 15960 7165 16005 7215
rect 16055 7165 16090 7215
rect 12890 7125 16090 7165
rect 12890 7075 12925 7125
rect 12975 7075 13020 7125
rect 13070 7075 13115 7125
rect 13165 7075 13215 7125
rect 13265 7075 13315 7125
rect 13365 7075 13415 7125
rect 13465 7075 13510 7125
rect 13560 7075 13605 7125
rect 13655 7075 13725 7125
rect 13775 7075 13820 7125
rect 13870 7075 13915 7125
rect 13965 7075 14015 7125
rect 14065 7075 14115 7125
rect 14165 7075 14215 7125
rect 14265 7075 14310 7125
rect 14360 7075 14405 7125
rect 14455 7075 14525 7125
rect 14575 7075 14620 7125
rect 14670 7075 14715 7125
rect 14765 7075 14815 7125
rect 14865 7075 14915 7125
rect 14965 7075 15015 7125
rect 15065 7075 15110 7125
rect 15160 7075 15205 7125
rect 15255 7075 15325 7125
rect 15375 7075 15420 7125
rect 15470 7075 15515 7125
rect 15565 7075 15615 7125
rect 15665 7075 15715 7125
rect 15765 7075 15815 7125
rect 15865 7075 15910 7125
rect 15960 7075 16005 7125
rect 16055 7075 16090 7125
rect 12890 7025 16090 7075
rect 12890 6975 12925 7025
rect 12975 6975 13020 7025
rect 13070 6975 13115 7025
rect 13165 6975 13215 7025
rect 13265 6975 13315 7025
rect 13365 6975 13415 7025
rect 13465 6975 13510 7025
rect 13560 6975 13605 7025
rect 13655 6975 13725 7025
rect 13775 6975 13820 7025
rect 13870 6975 13915 7025
rect 13965 6975 14015 7025
rect 14065 6975 14115 7025
rect 14165 6975 14215 7025
rect 14265 6975 14310 7025
rect 14360 6975 14405 7025
rect 14455 6975 14525 7025
rect 14575 6975 14620 7025
rect 14670 6975 14715 7025
rect 14765 6975 14815 7025
rect 14865 6975 14915 7025
rect 14965 6975 15015 7025
rect 15065 6975 15110 7025
rect 15160 6975 15205 7025
rect 15255 6975 15325 7025
rect 15375 6975 15420 7025
rect 15470 6975 15515 7025
rect 15565 6975 15615 7025
rect 15665 6975 15715 7025
rect 15765 6975 15815 7025
rect 15865 6975 15910 7025
rect 15960 6975 16005 7025
rect 16055 6975 16090 7025
rect 12890 6935 16090 6975
rect 12890 6885 12925 6935
rect 12975 6885 13020 6935
rect 13070 6885 13115 6935
rect 13165 6885 13215 6935
rect 13265 6885 13315 6935
rect 13365 6885 13415 6935
rect 13465 6885 13510 6935
rect 13560 6885 13605 6935
rect 13655 6885 13725 6935
rect 13775 6885 13820 6935
rect 13870 6885 13915 6935
rect 13965 6885 14015 6935
rect 14065 6885 14115 6935
rect 14165 6885 14215 6935
rect 14265 6885 14310 6935
rect 14360 6885 14405 6935
rect 14455 6885 14525 6935
rect 14575 6885 14620 6935
rect 14670 6885 14715 6935
rect 14765 6885 14815 6935
rect 14865 6885 14915 6935
rect 14965 6885 15015 6935
rect 15065 6885 15110 6935
rect 15160 6885 15205 6935
rect 15255 6885 15325 6935
rect 15375 6885 15420 6935
rect 15470 6885 15515 6935
rect 15565 6885 15615 6935
rect 15665 6885 15715 6935
rect 15765 6885 15815 6935
rect 15865 6885 15910 6935
rect 15960 6885 16005 6935
rect 16055 6885 16090 6935
rect 12890 6815 16090 6885
rect 12890 6765 12925 6815
rect 12975 6765 13020 6815
rect 13070 6765 13115 6815
rect 13165 6765 13215 6815
rect 13265 6765 13315 6815
rect 13365 6765 13415 6815
rect 13465 6765 13510 6815
rect 13560 6765 13605 6815
rect 13655 6765 13725 6815
rect 13775 6765 13820 6815
rect 13870 6765 13915 6815
rect 13965 6765 14015 6815
rect 14065 6765 14115 6815
rect 14165 6765 14215 6815
rect 14265 6765 14310 6815
rect 14360 6765 14405 6815
rect 14455 6765 14525 6815
rect 14575 6765 14620 6815
rect 14670 6765 14715 6815
rect 14765 6765 14815 6815
rect 14865 6765 14915 6815
rect 14965 6765 15015 6815
rect 15065 6765 15110 6815
rect 15160 6765 15205 6815
rect 15255 6765 15325 6815
rect 15375 6765 15420 6815
rect 15470 6765 15515 6815
rect 15565 6765 15615 6815
rect 15665 6765 15715 6815
rect 15765 6765 15815 6815
rect 15865 6765 15910 6815
rect 15960 6765 16005 6815
rect 16055 6765 16090 6815
rect 12890 6725 16090 6765
rect 12890 6675 12925 6725
rect 12975 6675 13020 6725
rect 13070 6675 13115 6725
rect 13165 6675 13215 6725
rect 13265 6675 13315 6725
rect 13365 6675 13415 6725
rect 13465 6675 13510 6725
rect 13560 6675 13605 6725
rect 13655 6675 13725 6725
rect 13775 6675 13820 6725
rect 13870 6675 13915 6725
rect 13965 6675 14015 6725
rect 14065 6675 14115 6725
rect 14165 6675 14215 6725
rect 14265 6675 14310 6725
rect 14360 6675 14405 6725
rect 14455 6675 14525 6725
rect 14575 6675 14620 6725
rect 14670 6675 14715 6725
rect 14765 6675 14815 6725
rect 14865 6675 14915 6725
rect 14965 6675 15015 6725
rect 15065 6675 15110 6725
rect 15160 6675 15205 6725
rect 15255 6675 15325 6725
rect 15375 6675 15420 6725
rect 15470 6675 15515 6725
rect 15565 6675 15615 6725
rect 15665 6675 15715 6725
rect 15765 6675 15815 6725
rect 15865 6675 15910 6725
rect 15960 6675 16005 6725
rect 16055 6675 16090 6725
rect 12890 6625 16090 6675
rect 12890 6575 12925 6625
rect 12975 6575 13020 6625
rect 13070 6575 13115 6625
rect 13165 6575 13215 6625
rect 13265 6575 13315 6625
rect 13365 6575 13415 6625
rect 13465 6575 13510 6625
rect 13560 6575 13605 6625
rect 13655 6575 13725 6625
rect 13775 6575 13820 6625
rect 13870 6575 13915 6625
rect 13965 6575 14015 6625
rect 14065 6575 14115 6625
rect 14165 6575 14215 6625
rect 14265 6575 14310 6625
rect 14360 6575 14405 6625
rect 14455 6575 14525 6625
rect 14575 6575 14620 6625
rect 14670 6575 14715 6625
rect 14765 6575 14815 6625
rect 14865 6575 14915 6625
rect 14965 6575 15015 6625
rect 15065 6575 15110 6625
rect 15160 6575 15205 6625
rect 15255 6575 15325 6625
rect 15375 6575 15420 6625
rect 15470 6575 15515 6625
rect 15565 6575 15615 6625
rect 15665 6575 15715 6625
rect 15765 6575 15815 6625
rect 15865 6575 15910 6625
rect 15960 6575 16005 6625
rect 16055 6575 16090 6625
rect 12890 6535 16090 6575
rect 12890 6485 12925 6535
rect 12975 6485 13020 6535
rect 13070 6485 13115 6535
rect 13165 6485 13215 6535
rect 13265 6485 13315 6535
rect 13365 6485 13415 6535
rect 13465 6485 13510 6535
rect 13560 6485 13605 6535
rect 13655 6485 13725 6535
rect 13775 6485 13820 6535
rect 13870 6485 13915 6535
rect 13965 6485 14015 6535
rect 14065 6485 14115 6535
rect 14165 6485 14215 6535
rect 14265 6485 14310 6535
rect 14360 6485 14405 6535
rect 14455 6485 14525 6535
rect 14575 6485 14620 6535
rect 14670 6485 14715 6535
rect 14765 6485 14815 6535
rect 14865 6485 14915 6535
rect 14965 6485 15015 6535
rect 15065 6485 15110 6535
rect 15160 6485 15205 6535
rect 15255 6485 15325 6535
rect 15375 6485 15420 6535
rect 15470 6485 15515 6535
rect 15565 6485 15615 6535
rect 15665 6485 15715 6535
rect 15765 6485 15815 6535
rect 15865 6485 15910 6535
rect 15960 6485 16005 6535
rect 16055 6485 16090 6535
rect -90 -1300 -30 -1290
rect -90 -1340 -80 -1300
rect -40 -1340 -30 -1300
rect -90 -1365 -30 -1340
rect -90 -1405 -80 -1365
rect -40 -1405 -30 -1365
rect -90 -1435 -30 -1405
rect -90 -1475 -80 -1435
rect -40 -1475 -30 -1435
rect -90 -1505 -30 -1475
rect -90 -1545 -80 -1505
rect -40 -1545 -30 -1505
rect -90 -1575 -30 -1545
rect -90 -1615 -80 -1575
rect -40 -1615 -30 -1575
rect -90 -1640 -30 -1615
rect -90 -1680 -80 -1640
rect -40 -1680 -30 -1640
rect -90 -1700 -30 -1680
rect -90 -1740 -80 -1700
rect -40 -1740 -30 -1700
rect -90 -1765 -30 -1740
rect -90 -1805 -80 -1765
rect -40 -1805 -30 -1765
rect -90 -1835 -30 -1805
rect -90 -1875 -80 -1835
rect -40 -1875 -30 -1835
rect -90 -1905 -30 -1875
rect -90 -1945 -80 -1905
rect -40 -1945 -30 -1905
rect -90 -1975 -30 -1945
rect -90 -2015 -80 -1975
rect -40 -2015 -30 -1975
rect -90 -2040 -30 -2015
rect -90 -2080 -80 -2040
rect -40 -2080 -30 -2040
rect -90 -2100 -30 -2080
rect -90 -2140 -80 -2100
rect -40 -2140 -30 -2100
rect -90 -2165 -30 -2140
rect -90 -2205 -80 -2165
rect -40 -2205 -30 -2165
rect -90 -2235 -30 -2205
rect -90 -2275 -80 -2235
rect -40 -2275 -30 -2235
rect -90 -2305 -30 -2275
rect -90 -2345 -80 -2305
rect -40 -2345 -30 -2305
rect -90 -2375 -30 -2345
rect -90 -2415 -80 -2375
rect -40 -2415 -30 -2375
rect -90 -2440 -30 -2415
rect -90 -2480 -80 -2440
rect -40 -2480 -30 -2440
rect -90 -2500 -30 -2480
rect -90 -2540 -80 -2500
rect -40 -2540 -30 -2500
rect -90 -2565 -30 -2540
rect -90 -2605 -80 -2565
rect -40 -2605 -30 -2565
rect -90 -2635 -30 -2605
rect -90 -2675 -80 -2635
rect -40 -2675 -30 -2635
rect -90 -2705 -30 -2675
rect -90 -2745 -80 -2705
rect -40 -2745 -30 -2705
rect -90 -2775 -30 -2745
rect -90 -2815 -80 -2775
rect -40 -2815 -30 -2775
rect -90 -2840 -30 -2815
rect -90 -2880 -80 -2840
rect -40 -2880 -30 -2840
rect -90 -2900 -30 -2880
rect -90 -2940 -80 -2900
rect -40 -2940 -30 -2900
rect -90 -2965 -30 -2940
rect -90 -3005 -80 -2965
rect -40 -3005 -30 -2965
rect -90 -3035 -30 -3005
rect -90 -3075 -80 -3035
rect -40 -3075 -30 -3035
rect -90 -3105 -30 -3075
rect -90 -3145 -80 -3105
rect -40 -3145 -30 -3105
rect -90 -3175 -30 -3145
rect -90 -3215 -80 -3175
rect -40 -3215 -30 -3175
rect -90 -3240 -30 -3215
rect -90 -3280 -80 -3240
rect -40 -3280 -30 -3240
rect -90 -3300 -30 -3280
rect -90 -3340 -80 -3300
rect -40 -3340 -30 -3300
rect -90 -3365 -30 -3340
rect -90 -3405 -80 -3365
rect -40 -3405 -30 -3365
rect -90 -3435 -30 -3405
rect -90 -3475 -80 -3435
rect -40 -3475 -30 -3435
rect -90 -3505 -30 -3475
rect -90 -3545 -80 -3505
rect -40 -3545 -30 -3505
rect -90 -3575 -30 -3545
rect -90 -3615 -80 -3575
rect -40 -3615 -30 -3575
rect -90 -3640 -30 -3615
rect -90 -3680 -80 -3640
rect -40 -3680 -30 -3640
rect -90 -3700 -30 -3680
rect -90 -3740 -80 -3700
rect -40 -3740 -30 -3700
rect -90 -3765 -30 -3740
rect -90 -3805 -80 -3765
rect -40 -3805 -30 -3765
rect -90 -3835 -30 -3805
rect -90 -3875 -80 -3835
rect -40 -3875 -30 -3835
rect -90 -3905 -30 -3875
rect -90 -3945 -80 -3905
rect -40 -3945 -30 -3905
rect -90 -3975 -30 -3945
rect -90 -4015 -80 -3975
rect -40 -4015 -30 -3975
rect -90 -4040 -30 -4015
rect -90 -4080 -80 -4040
rect -40 -4080 -30 -4040
rect -90 -4100 -30 -4080
rect -90 -4140 -80 -4100
rect -40 -4140 -30 -4100
rect -90 -4165 -30 -4140
rect -90 -4205 -80 -4165
rect -40 -4205 -30 -4165
rect -90 -4235 -30 -4205
rect -90 -4275 -80 -4235
rect -40 -4275 -30 -4235
rect -90 -4305 -30 -4275
rect -90 -4345 -80 -4305
rect -40 -4345 -30 -4305
rect -90 -4375 -30 -4345
rect -90 -4415 -80 -4375
rect -40 -4415 -30 -4375
rect -90 -4440 -30 -4415
rect -90 -4480 -80 -4440
rect -40 -4480 -30 -4440
rect -90 -4490 -30 -4480
rect 260 -1300 320 -1290
rect 260 -1340 270 -1300
rect 310 -1340 320 -1300
rect 260 -1365 320 -1340
rect 260 -1405 270 -1365
rect 310 -1405 320 -1365
rect 260 -1435 320 -1405
rect 260 -1475 270 -1435
rect 310 -1475 320 -1435
rect 260 -1505 320 -1475
rect 260 -1545 270 -1505
rect 310 -1545 320 -1505
rect 260 -1575 320 -1545
rect 260 -1615 270 -1575
rect 310 -1615 320 -1575
rect 260 -1640 320 -1615
rect 260 -1680 270 -1640
rect 310 -1680 320 -1640
rect 260 -1700 320 -1680
rect 260 -1740 270 -1700
rect 310 -1740 320 -1700
rect 260 -1765 320 -1740
rect 260 -1805 270 -1765
rect 310 -1805 320 -1765
rect 260 -1835 320 -1805
rect 260 -1875 270 -1835
rect 310 -1875 320 -1835
rect 260 -1905 320 -1875
rect 260 -1945 270 -1905
rect 310 -1945 320 -1905
rect 260 -1975 320 -1945
rect 260 -2015 270 -1975
rect 310 -2015 320 -1975
rect 260 -2040 320 -2015
rect 260 -2080 270 -2040
rect 310 -2080 320 -2040
rect 260 -2100 320 -2080
rect 260 -2140 270 -2100
rect 310 -2140 320 -2100
rect 260 -2165 320 -2140
rect 260 -2205 270 -2165
rect 310 -2205 320 -2165
rect 260 -2235 320 -2205
rect 260 -2275 270 -2235
rect 310 -2275 320 -2235
rect 260 -2305 320 -2275
rect 260 -2345 270 -2305
rect 310 -2345 320 -2305
rect 260 -2375 320 -2345
rect 260 -2415 270 -2375
rect 310 -2415 320 -2375
rect 260 -2440 320 -2415
rect 260 -2480 270 -2440
rect 310 -2480 320 -2440
rect 260 -2500 320 -2480
rect 260 -2540 270 -2500
rect 310 -2540 320 -2500
rect 260 -2565 320 -2540
rect 260 -2605 270 -2565
rect 310 -2605 320 -2565
rect 260 -2635 320 -2605
rect 260 -2675 270 -2635
rect 310 -2675 320 -2635
rect 260 -2705 320 -2675
rect 260 -2745 270 -2705
rect 310 -2745 320 -2705
rect 260 -2775 320 -2745
rect 260 -2815 270 -2775
rect 310 -2815 320 -2775
rect 260 -2840 320 -2815
rect 260 -2880 270 -2840
rect 310 -2880 320 -2840
rect 260 -2900 320 -2880
rect 260 -2940 270 -2900
rect 310 -2940 320 -2900
rect 260 -2965 320 -2940
rect 260 -3005 270 -2965
rect 310 -3005 320 -2965
rect 260 -3035 320 -3005
rect 260 -3075 270 -3035
rect 310 -3075 320 -3035
rect 260 -3105 320 -3075
rect 260 -3145 270 -3105
rect 310 -3145 320 -3105
rect 260 -3175 320 -3145
rect 260 -3215 270 -3175
rect 310 -3215 320 -3175
rect 260 -3240 320 -3215
rect 260 -3280 270 -3240
rect 310 -3280 320 -3240
rect 260 -3300 320 -3280
rect 260 -3340 270 -3300
rect 310 -3340 320 -3300
rect 260 -3365 320 -3340
rect 260 -3405 270 -3365
rect 310 -3405 320 -3365
rect 260 -3435 320 -3405
rect 260 -3475 270 -3435
rect 310 -3475 320 -3435
rect 260 -3505 320 -3475
rect 260 -3545 270 -3505
rect 310 -3545 320 -3505
rect 260 -3575 320 -3545
rect 260 -3615 270 -3575
rect 310 -3615 320 -3575
rect 260 -3640 320 -3615
rect 260 -3680 270 -3640
rect 310 -3680 320 -3640
rect 260 -3700 320 -3680
rect 260 -3740 270 -3700
rect 310 -3740 320 -3700
rect 260 -3765 320 -3740
rect 260 -3805 270 -3765
rect 310 -3805 320 -3765
rect 260 -3835 320 -3805
rect 260 -3875 270 -3835
rect 310 -3875 320 -3835
rect 260 -3905 320 -3875
rect 260 -3945 270 -3905
rect 310 -3945 320 -3905
rect 260 -3975 320 -3945
rect 260 -4015 270 -3975
rect 310 -4015 320 -3975
rect 260 -4040 320 -4015
rect 260 -4080 270 -4040
rect 310 -4080 320 -4040
rect 260 -4100 320 -4080
rect 260 -4140 270 -4100
rect 310 -4140 320 -4100
rect 260 -4165 320 -4140
rect 260 -4205 270 -4165
rect 310 -4205 320 -4165
rect 260 -4235 320 -4205
rect 260 -4275 270 -4235
rect 310 -4275 320 -4235
rect 260 -4305 320 -4275
rect 260 -4345 270 -4305
rect 310 -4345 320 -4305
rect 260 -4375 320 -4345
rect 260 -4415 270 -4375
rect 310 -4415 320 -4375
rect 260 -4440 320 -4415
rect 260 -4480 270 -4440
rect 310 -4480 320 -4440
rect 260 -4490 320 -4480
rect 610 -1300 670 -1290
rect 610 -1340 620 -1300
rect 660 -1340 670 -1300
rect 610 -1365 670 -1340
rect 610 -1405 620 -1365
rect 660 -1405 670 -1365
rect 610 -1435 670 -1405
rect 610 -1475 620 -1435
rect 660 -1475 670 -1435
rect 610 -1505 670 -1475
rect 610 -1545 620 -1505
rect 660 -1545 670 -1505
rect 610 -1575 670 -1545
rect 610 -1615 620 -1575
rect 660 -1615 670 -1575
rect 610 -1640 670 -1615
rect 610 -1680 620 -1640
rect 660 -1680 670 -1640
rect 610 -1700 670 -1680
rect 610 -1740 620 -1700
rect 660 -1740 670 -1700
rect 610 -1765 670 -1740
rect 610 -1805 620 -1765
rect 660 -1805 670 -1765
rect 610 -1835 670 -1805
rect 610 -1875 620 -1835
rect 660 -1875 670 -1835
rect 610 -1905 670 -1875
rect 610 -1945 620 -1905
rect 660 -1945 670 -1905
rect 610 -1975 670 -1945
rect 610 -2015 620 -1975
rect 660 -2015 670 -1975
rect 610 -2040 670 -2015
rect 610 -2080 620 -2040
rect 660 -2080 670 -2040
rect 610 -2100 670 -2080
rect 610 -2140 620 -2100
rect 660 -2140 670 -2100
rect 610 -2165 670 -2140
rect 610 -2205 620 -2165
rect 660 -2205 670 -2165
rect 610 -2235 670 -2205
rect 610 -2275 620 -2235
rect 660 -2275 670 -2235
rect 610 -2305 670 -2275
rect 610 -2345 620 -2305
rect 660 -2345 670 -2305
rect 610 -2375 670 -2345
rect 610 -2415 620 -2375
rect 660 -2415 670 -2375
rect 610 -2440 670 -2415
rect 610 -2480 620 -2440
rect 660 -2480 670 -2440
rect 610 -2500 670 -2480
rect 610 -2540 620 -2500
rect 660 -2540 670 -2500
rect 610 -2565 670 -2540
rect 610 -2605 620 -2565
rect 660 -2605 670 -2565
rect 610 -2635 670 -2605
rect 610 -2675 620 -2635
rect 660 -2675 670 -2635
rect 610 -2705 670 -2675
rect 610 -2745 620 -2705
rect 660 -2745 670 -2705
rect 610 -2775 670 -2745
rect 610 -2815 620 -2775
rect 660 -2815 670 -2775
rect 610 -2840 670 -2815
rect 610 -2880 620 -2840
rect 660 -2880 670 -2840
rect 610 -2900 670 -2880
rect 610 -2940 620 -2900
rect 660 -2940 670 -2900
rect 610 -2965 670 -2940
rect 610 -3005 620 -2965
rect 660 -3005 670 -2965
rect 610 -3035 670 -3005
rect 610 -3075 620 -3035
rect 660 -3075 670 -3035
rect 610 -3105 670 -3075
rect 610 -3145 620 -3105
rect 660 -3145 670 -3105
rect 610 -3175 670 -3145
rect 610 -3215 620 -3175
rect 660 -3215 670 -3175
rect 610 -3240 670 -3215
rect 610 -3280 620 -3240
rect 660 -3280 670 -3240
rect 610 -3300 670 -3280
rect 610 -3340 620 -3300
rect 660 -3340 670 -3300
rect 610 -3365 670 -3340
rect 610 -3405 620 -3365
rect 660 -3405 670 -3365
rect 610 -3435 670 -3405
rect 610 -3475 620 -3435
rect 660 -3475 670 -3435
rect 610 -3505 670 -3475
rect 610 -3545 620 -3505
rect 660 -3545 670 -3505
rect 610 -3575 670 -3545
rect 610 -3615 620 -3575
rect 660 -3615 670 -3575
rect 610 -3640 670 -3615
rect 610 -3680 620 -3640
rect 660 -3680 670 -3640
rect 610 -3700 670 -3680
rect 610 -3740 620 -3700
rect 660 -3740 670 -3700
rect 610 -3765 670 -3740
rect 610 -3805 620 -3765
rect 660 -3805 670 -3765
rect 610 -3835 670 -3805
rect 610 -3875 620 -3835
rect 660 -3875 670 -3835
rect 610 -3905 670 -3875
rect 610 -3945 620 -3905
rect 660 -3945 670 -3905
rect 610 -3975 670 -3945
rect 610 -4015 620 -3975
rect 660 -4015 670 -3975
rect 610 -4040 670 -4015
rect 610 -4080 620 -4040
rect 660 -4080 670 -4040
rect 610 -4100 670 -4080
rect 610 -4140 620 -4100
rect 660 -4140 670 -4100
rect 610 -4165 670 -4140
rect 610 -4205 620 -4165
rect 660 -4205 670 -4165
rect 610 -4235 670 -4205
rect 610 -4275 620 -4235
rect 660 -4275 670 -4235
rect 610 -4305 670 -4275
rect 610 -4345 620 -4305
rect 660 -4345 670 -4305
rect 610 -4375 670 -4345
rect 610 -4415 620 -4375
rect 660 -4415 670 -4375
rect 610 -4440 670 -4415
rect 610 -4480 620 -4440
rect 660 -4480 670 -4440
rect 610 -4490 670 -4480
rect 960 -1300 1020 -1290
rect 960 -1340 970 -1300
rect 1010 -1340 1020 -1300
rect 960 -1365 1020 -1340
rect 960 -1405 970 -1365
rect 1010 -1405 1020 -1365
rect 960 -1435 1020 -1405
rect 960 -1475 970 -1435
rect 1010 -1475 1020 -1435
rect 960 -1505 1020 -1475
rect 960 -1545 970 -1505
rect 1010 -1545 1020 -1505
rect 960 -1575 1020 -1545
rect 960 -1615 970 -1575
rect 1010 -1615 1020 -1575
rect 960 -1640 1020 -1615
rect 960 -1680 970 -1640
rect 1010 -1680 1020 -1640
rect 960 -1700 1020 -1680
rect 960 -1740 970 -1700
rect 1010 -1740 1020 -1700
rect 960 -1765 1020 -1740
rect 960 -1805 970 -1765
rect 1010 -1805 1020 -1765
rect 960 -1835 1020 -1805
rect 960 -1875 970 -1835
rect 1010 -1875 1020 -1835
rect 960 -1905 1020 -1875
rect 960 -1945 970 -1905
rect 1010 -1945 1020 -1905
rect 960 -1975 1020 -1945
rect 960 -2015 970 -1975
rect 1010 -2015 1020 -1975
rect 960 -2040 1020 -2015
rect 960 -2080 970 -2040
rect 1010 -2080 1020 -2040
rect 960 -2100 1020 -2080
rect 960 -2140 970 -2100
rect 1010 -2140 1020 -2100
rect 960 -2165 1020 -2140
rect 960 -2205 970 -2165
rect 1010 -2205 1020 -2165
rect 960 -2235 1020 -2205
rect 960 -2275 970 -2235
rect 1010 -2275 1020 -2235
rect 960 -2305 1020 -2275
rect 960 -2345 970 -2305
rect 1010 -2345 1020 -2305
rect 960 -2375 1020 -2345
rect 960 -2415 970 -2375
rect 1010 -2415 1020 -2375
rect 960 -2440 1020 -2415
rect 960 -2480 970 -2440
rect 1010 -2480 1020 -2440
rect 960 -2500 1020 -2480
rect 960 -2540 970 -2500
rect 1010 -2540 1020 -2500
rect 960 -2565 1020 -2540
rect 960 -2605 970 -2565
rect 1010 -2605 1020 -2565
rect 960 -2635 1020 -2605
rect 960 -2675 970 -2635
rect 1010 -2675 1020 -2635
rect 960 -2705 1020 -2675
rect 960 -2745 970 -2705
rect 1010 -2745 1020 -2705
rect 960 -2775 1020 -2745
rect 960 -2815 970 -2775
rect 1010 -2815 1020 -2775
rect 960 -2840 1020 -2815
rect 960 -2880 970 -2840
rect 1010 -2880 1020 -2840
rect 960 -2900 1020 -2880
rect 960 -2940 970 -2900
rect 1010 -2940 1020 -2900
rect 960 -2965 1020 -2940
rect 960 -3005 970 -2965
rect 1010 -3005 1020 -2965
rect 960 -3035 1020 -3005
rect 960 -3075 970 -3035
rect 1010 -3075 1020 -3035
rect 960 -3105 1020 -3075
rect 960 -3145 970 -3105
rect 1010 -3145 1020 -3105
rect 960 -3175 1020 -3145
rect 960 -3215 970 -3175
rect 1010 -3215 1020 -3175
rect 960 -3240 1020 -3215
rect 960 -3280 970 -3240
rect 1010 -3280 1020 -3240
rect 960 -3300 1020 -3280
rect 960 -3340 970 -3300
rect 1010 -3340 1020 -3300
rect 960 -3365 1020 -3340
rect 960 -3405 970 -3365
rect 1010 -3405 1020 -3365
rect 960 -3435 1020 -3405
rect 960 -3475 970 -3435
rect 1010 -3475 1020 -3435
rect 960 -3505 1020 -3475
rect 960 -3545 970 -3505
rect 1010 -3545 1020 -3505
rect 960 -3575 1020 -3545
rect 960 -3615 970 -3575
rect 1010 -3615 1020 -3575
rect 960 -3640 1020 -3615
rect 960 -3680 970 -3640
rect 1010 -3680 1020 -3640
rect 960 -3700 1020 -3680
rect 960 -3740 970 -3700
rect 1010 -3740 1020 -3700
rect 960 -3765 1020 -3740
rect 960 -3805 970 -3765
rect 1010 -3805 1020 -3765
rect 960 -3835 1020 -3805
rect 960 -3875 970 -3835
rect 1010 -3875 1020 -3835
rect 960 -3905 1020 -3875
rect 960 -3945 970 -3905
rect 1010 -3945 1020 -3905
rect 960 -3975 1020 -3945
rect 960 -4015 970 -3975
rect 1010 -4015 1020 -3975
rect 960 -4040 1020 -4015
rect 960 -4080 970 -4040
rect 1010 -4080 1020 -4040
rect 960 -4100 1020 -4080
rect 960 -4140 970 -4100
rect 1010 -4140 1020 -4100
rect 960 -4165 1020 -4140
rect 960 -4205 970 -4165
rect 1010 -4205 1020 -4165
rect 960 -4235 1020 -4205
rect 960 -4275 970 -4235
rect 1010 -4275 1020 -4235
rect 960 -4305 1020 -4275
rect 960 -4345 970 -4305
rect 1010 -4345 1020 -4305
rect 960 -4375 1020 -4345
rect 960 -4415 970 -4375
rect 1010 -4415 1020 -4375
rect 960 -4440 1020 -4415
rect 960 -4480 970 -4440
rect 1010 -4480 1020 -4440
rect 960 -4490 1020 -4480
rect 1310 -1300 1370 -1290
rect 1310 -1340 1320 -1300
rect 1360 -1340 1370 -1300
rect 1310 -1365 1370 -1340
rect 1310 -1405 1320 -1365
rect 1360 -1405 1370 -1365
rect 1310 -1435 1370 -1405
rect 1310 -1475 1320 -1435
rect 1360 -1475 1370 -1435
rect 1310 -1505 1370 -1475
rect 1310 -1545 1320 -1505
rect 1360 -1545 1370 -1505
rect 1310 -1575 1370 -1545
rect 1310 -1615 1320 -1575
rect 1360 -1615 1370 -1575
rect 1310 -1640 1370 -1615
rect 1310 -1680 1320 -1640
rect 1360 -1680 1370 -1640
rect 1310 -1700 1370 -1680
rect 1310 -1740 1320 -1700
rect 1360 -1740 1370 -1700
rect 1310 -1765 1370 -1740
rect 1310 -1805 1320 -1765
rect 1360 -1805 1370 -1765
rect 1310 -1835 1370 -1805
rect 1310 -1875 1320 -1835
rect 1360 -1875 1370 -1835
rect 1310 -1905 1370 -1875
rect 1310 -1945 1320 -1905
rect 1360 -1945 1370 -1905
rect 1310 -1975 1370 -1945
rect 1310 -2015 1320 -1975
rect 1360 -2015 1370 -1975
rect 1310 -2040 1370 -2015
rect 1310 -2080 1320 -2040
rect 1360 -2080 1370 -2040
rect 1310 -2100 1370 -2080
rect 1310 -2140 1320 -2100
rect 1360 -2140 1370 -2100
rect 1310 -2165 1370 -2140
rect 1310 -2205 1320 -2165
rect 1360 -2205 1370 -2165
rect 1310 -2235 1370 -2205
rect 1310 -2275 1320 -2235
rect 1360 -2275 1370 -2235
rect 1310 -2305 1370 -2275
rect 1310 -2345 1320 -2305
rect 1360 -2345 1370 -2305
rect 1310 -2375 1370 -2345
rect 1310 -2415 1320 -2375
rect 1360 -2415 1370 -2375
rect 1310 -2440 1370 -2415
rect 1310 -2480 1320 -2440
rect 1360 -2480 1370 -2440
rect 1310 -2500 1370 -2480
rect 1310 -2540 1320 -2500
rect 1360 -2540 1370 -2500
rect 1310 -2565 1370 -2540
rect 1310 -2605 1320 -2565
rect 1360 -2605 1370 -2565
rect 1310 -2635 1370 -2605
rect 1310 -2675 1320 -2635
rect 1360 -2675 1370 -2635
rect 1310 -2705 1370 -2675
rect 1310 -2745 1320 -2705
rect 1360 -2745 1370 -2705
rect 1310 -2775 1370 -2745
rect 1310 -2815 1320 -2775
rect 1360 -2815 1370 -2775
rect 1310 -2840 1370 -2815
rect 1310 -2880 1320 -2840
rect 1360 -2880 1370 -2840
rect 1310 -2900 1370 -2880
rect 1310 -2940 1320 -2900
rect 1360 -2940 1370 -2900
rect 1310 -2965 1370 -2940
rect 1310 -3005 1320 -2965
rect 1360 -3005 1370 -2965
rect 1310 -3035 1370 -3005
rect 1310 -3075 1320 -3035
rect 1360 -3075 1370 -3035
rect 1310 -3105 1370 -3075
rect 1310 -3145 1320 -3105
rect 1360 -3145 1370 -3105
rect 1310 -3175 1370 -3145
rect 1310 -3215 1320 -3175
rect 1360 -3215 1370 -3175
rect 1310 -3240 1370 -3215
rect 1310 -3280 1320 -3240
rect 1360 -3280 1370 -3240
rect 1310 -3300 1370 -3280
rect 1310 -3340 1320 -3300
rect 1360 -3340 1370 -3300
rect 1310 -3365 1370 -3340
rect 1310 -3405 1320 -3365
rect 1360 -3405 1370 -3365
rect 1310 -3435 1370 -3405
rect 1310 -3475 1320 -3435
rect 1360 -3475 1370 -3435
rect 1310 -3505 1370 -3475
rect 1310 -3545 1320 -3505
rect 1360 -3545 1370 -3505
rect 1310 -3575 1370 -3545
rect 1310 -3615 1320 -3575
rect 1360 -3615 1370 -3575
rect 1310 -3640 1370 -3615
rect 1310 -3680 1320 -3640
rect 1360 -3680 1370 -3640
rect 1310 -3700 1370 -3680
rect 1310 -3740 1320 -3700
rect 1360 -3740 1370 -3700
rect 1310 -3765 1370 -3740
rect 1310 -3805 1320 -3765
rect 1360 -3805 1370 -3765
rect 1310 -3835 1370 -3805
rect 1310 -3875 1320 -3835
rect 1360 -3875 1370 -3835
rect 1310 -3905 1370 -3875
rect 1310 -3945 1320 -3905
rect 1360 -3945 1370 -3905
rect 1310 -3975 1370 -3945
rect 1310 -4015 1320 -3975
rect 1360 -4015 1370 -3975
rect 1310 -4040 1370 -4015
rect 1310 -4080 1320 -4040
rect 1360 -4080 1370 -4040
rect 1310 -4100 1370 -4080
rect 1310 -4140 1320 -4100
rect 1360 -4140 1370 -4100
rect 1310 -4165 1370 -4140
rect 1310 -4205 1320 -4165
rect 1360 -4205 1370 -4165
rect 1310 -4235 1370 -4205
rect 1310 -4275 1320 -4235
rect 1360 -4275 1370 -4235
rect 1310 -4305 1370 -4275
rect 1310 -4345 1320 -4305
rect 1360 -4345 1370 -4305
rect 1310 -4375 1370 -4345
rect 1310 -4415 1320 -4375
rect 1360 -4415 1370 -4375
rect 1310 -4440 1370 -4415
rect 1310 -4480 1320 -4440
rect 1360 -4480 1370 -4440
rect 1310 -4490 1370 -4480
rect 1660 -1300 1720 -1290
rect 1660 -1340 1670 -1300
rect 1710 -1340 1720 -1300
rect 1660 -1365 1720 -1340
rect 1660 -1405 1670 -1365
rect 1710 -1405 1720 -1365
rect 1660 -1435 1720 -1405
rect 1660 -1475 1670 -1435
rect 1710 -1475 1720 -1435
rect 1660 -1505 1720 -1475
rect 1660 -1545 1670 -1505
rect 1710 -1545 1720 -1505
rect 1660 -1575 1720 -1545
rect 1660 -1615 1670 -1575
rect 1710 -1615 1720 -1575
rect 1660 -1640 1720 -1615
rect 1660 -1680 1670 -1640
rect 1710 -1680 1720 -1640
rect 1660 -1700 1720 -1680
rect 1660 -1740 1670 -1700
rect 1710 -1740 1720 -1700
rect 1660 -1765 1720 -1740
rect 1660 -1805 1670 -1765
rect 1710 -1805 1720 -1765
rect 1660 -1835 1720 -1805
rect 1660 -1875 1670 -1835
rect 1710 -1875 1720 -1835
rect 1660 -1905 1720 -1875
rect 1660 -1945 1670 -1905
rect 1710 -1945 1720 -1905
rect 1660 -1975 1720 -1945
rect 1660 -2015 1670 -1975
rect 1710 -2015 1720 -1975
rect 1660 -2040 1720 -2015
rect 1660 -2080 1670 -2040
rect 1710 -2080 1720 -2040
rect 1660 -2100 1720 -2080
rect 1660 -2140 1670 -2100
rect 1710 -2140 1720 -2100
rect 1660 -2165 1720 -2140
rect 1660 -2205 1670 -2165
rect 1710 -2205 1720 -2165
rect 1660 -2235 1720 -2205
rect 1660 -2275 1670 -2235
rect 1710 -2275 1720 -2235
rect 1660 -2305 1720 -2275
rect 1660 -2345 1670 -2305
rect 1710 -2345 1720 -2305
rect 1660 -2375 1720 -2345
rect 1660 -2415 1670 -2375
rect 1710 -2415 1720 -2375
rect 1660 -2440 1720 -2415
rect 1660 -2480 1670 -2440
rect 1710 -2480 1720 -2440
rect 1660 -2500 1720 -2480
rect 1660 -2540 1670 -2500
rect 1710 -2540 1720 -2500
rect 1660 -2565 1720 -2540
rect 1660 -2605 1670 -2565
rect 1710 -2605 1720 -2565
rect 1660 -2635 1720 -2605
rect 1660 -2675 1670 -2635
rect 1710 -2675 1720 -2635
rect 1660 -2705 1720 -2675
rect 1660 -2745 1670 -2705
rect 1710 -2745 1720 -2705
rect 1660 -2775 1720 -2745
rect 1660 -2815 1670 -2775
rect 1710 -2815 1720 -2775
rect 1660 -2840 1720 -2815
rect 1660 -2880 1670 -2840
rect 1710 -2880 1720 -2840
rect 1660 -2900 1720 -2880
rect 1660 -2940 1670 -2900
rect 1710 -2940 1720 -2900
rect 1660 -2965 1720 -2940
rect 1660 -3005 1670 -2965
rect 1710 -3005 1720 -2965
rect 1660 -3035 1720 -3005
rect 1660 -3075 1670 -3035
rect 1710 -3075 1720 -3035
rect 1660 -3105 1720 -3075
rect 1660 -3145 1670 -3105
rect 1710 -3145 1720 -3105
rect 1660 -3175 1720 -3145
rect 1660 -3215 1670 -3175
rect 1710 -3215 1720 -3175
rect 1660 -3240 1720 -3215
rect 1660 -3280 1670 -3240
rect 1710 -3280 1720 -3240
rect 1660 -3300 1720 -3280
rect 1660 -3340 1670 -3300
rect 1710 -3340 1720 -3300
rect 1660 -3365 1720 -3340
rect 1660 -3405 1670 -3365
rect 1710 -3405 1720 -3365
rect 1660 -3435 1720 -3405
rect 1660 -3475 1670 -3435
rect 1710 -3475 1720 -3435
rect 1660 -3505 1720 -3475
rect 1660 -3545 1670 -3505
rect 1710 -3545 1720 -3505
rect 1660 -3575 1720 -3545
rect 1660 -3615 1670 -3575
rect 1710 -3615 1720 -3575
rect 1660 -3640 1720 -3615
rect 1660 -3680 1670 -3640
rect 1710 -3680 1720 -3640
rect 1660 -3700 1720 -3680
rect 1660 -3740 1670 -3700
rect 1710 -3740 1720 -3700
rect 1660 -3765 1720 -3740
rect 1660 -3805 1670 -3765
rect 1710 -3805 1720 -3765
rect 1660 -3835 1720 -3805
rect 1660 -3875 1670 -3835
rect 1710 -3875 1720 -3835
rect 1660 -3905 1720 -3875
rect 1660 -3945 1670 -3905
rect 1710 -3945 1720 -3905
rect 1660 -3975 1720 -3945
rect 1660 -4015 1670 -3975
rect 1710 -4015 1720 -3975
rect 1660 -4040 1720 -4015
rect 1660 -4080 1670 -4040
rect 1710 -4080 1720 -4040
rect 1660 -4100 1720 -4080
rect 1660 -4140 1670 -4100
rect 1710 -4140 1720 -4100
rect 1660 -4165 1720 -4140
rect 1660 -4205 1670 -4165
rect 1710 -4205 1720 -4165
rect 1660 -4235 1720 -4205
rect 1660 -4275 1670 -4235
rect 1710 -4275 1720 -4235
rect 1660 -4305 1720 -4275
rect 1660 -4345 1670 -4305
rect 1710 -4345 1720 -4305
rect 1660 -4375 1720 -4345
rect 1660 -4415 1670 -4375
rect 1710 -4415 1720 -4375
rect 1660 -4440 1720 -4415
rect 1660 -4480 1670 -4440
rect 1710 -4480 1720 -4440
rect 1660 -4490 1720 -4480
rect 2010 -1300 2070 -1290
rect 2010 -1340 2020 -1300
rect 2060 -1340 2070 -1300
rect 2010 -1365 2070 -1340
rect 2010 -1405 2020 -1365
rect 2060 -1405 2070 -1365
rect 2010 -1435 2070 -1405
rect 2010 -1475 2020 -1435
rect 2060 -1475 2070 -1435
rect 2010 -1505 2070 -1475
rect 2010 -1545 2020 -1505
rect 2060 -1545 2070 -1505
rect 2010 -1575 2070 -1545
rect 2010 -1615 2020 -1575
rect 2060 -1615 2070 -1575
rect 2010 -1640 2070 -1615
rect 2010 -1680 2020 -1640
rect 2060 -1680 2070 -1640
rect 2010 -1700 2070 -1680
rect 2010 -1740 2020 -1700
rect 2060 -1740 2070 -1700
rect 2010 -1765 2070 -1740
rect 2010 -1805 2020 -1765
rect 2060 -1805 2070 -1765
rect 2010 -1835 2070 -1805
rect 2010 -1875 2020 -1835
rect 2060 -1875 2070 -1835
rect 2010 -1905 2070 -1875
rect 2010 -1945 2020 -1905
rect 2060 -1945 2070 -1905
rect 2010 -1975 2070 -1945
rect 2010 -2015 2020 -1975
rect 2060 -2015 2070 -1975
rect 2010 -2040 2070 -2015
rect 2010 -2080 2020 -2040
rect 2060 -2080 2070 -2040
rect 2010 -2100 2070 -2080
rect 2010 -2140 2020 -2100
rect 2060 -2140 2070 -2100
rect 2010 -2165 2070 -2140
rect 2010 -2205 2020 -2165
rect 2060 -2205 2070 -2165
rect 2010 -2235 2070 -2205
rect 2010 -2275 2020 -2235
rect 2060 -2275 2070 -2235
rect 2010 -2305 2070 -2275
rect 2010 -2345 2020 -2305
rect 2060 -2345 2070 -2305
rect 2010 -2375 2070 -2345
rect 2010 -2415 2020 -2375
rect 2060 -2415 2070 -2375
rect 2010 -2440 2070 -2415
rect 2010 -2480 2020 -2440
rect 2060 -2480 2070 -2440
rect 2010 -2500 2070 -2480
rect 2010 -2540 2020 -2500
rect 2060 -2540 2070 -2500
rect 2010 -2565 2070 -2540
rect 2010 -2605 2020 -2565
rect 2060 -2605 2070 -2565
rect 2010 -2635 2070 -2605
rect 2010 -2675 2020 -2635
rect 2060 -2675 2070 -2635
rect 2010 -2705 2070 -2675
rect 2010 -2745 2020 -2705
rect 2060 -2745 2070 -2705
rect 2010 -2775 2070 -2745
rect 2010 -2815 2020 -2775
rect 2060 -2815 2070 -2775
rect 2010 -2840 2070 -2815
rect 2010 -2880 2020 -2840
rect 2060 -2880 2070 -2840
rect 2010 -2900 2070 -2880
rect 2010 -2940 2020 -2900
rect 2060 -2940 2070 -2900
rect 2010 -2965 2070 -2940
rect 2010 -3005 2020 -2965
rect 2060 -3005 2070 -2965
rect 2010 -3035 2070 -3005
rect 2010 -3075 2020 -3035
rect 2060 -3075 2070 -3035
rect 2010 -3105 2070 -3075
rect 2010 -3145 2020 -3105
rect 2060 -3145 2070 -3105
rect 2010 -3175 2070 -3145
rect 2010 -3215 2020 -3175
rect 2060 -3215 2070 -3175
rect 2010 -3240 2070 -3215
rect 2010 -3280 2020 -3240
rect 2060 -3280 2070 -3240
rect 2010 -3300 2070 -3280
rect 2010 -3340 2020 -3300
rect 2060 -3340 2070 -3300
rect 2010 -3365 2070 -3340
rect 2010 -3405 2020 -3365
rect 2060 -3405 2070 -3365
rect 2010 -3435 2070 -3405
rect 2010 -3475 2020 -3435
rect 2060 -3475 2070 -3435
rect 2010 -3505 2070 -3475
rect 2010 -3545 2020 -3505
rect 2060 -3545 2070 -3505
rect 2010 -3575 2070 -3545
rect 2010 -3615 2020 -3575
rect 2060 -3615 2070 -3575
rect 2010 -3640 2070 -3615
rect 2010 -3680 2020 -3640
rect 2060 -3680 2070 -3640
rect 2010 -3700 2070 -3680
rect 2010 -3740 2020 -3700
rect 2060 -3740 2070 -3700
rect 2010 -3765 2070 -3740
rect 2010 -3805 2020 -3765
rect 2060 -3805 2070 -3765
rect 2010 -3835 2070 -3805
rect 2010 -3875 2020 -3835
rect 2060 -3875 2070 -3835
rect 2010 -3905 2070 -3875
rect 2010 -3945 2020 -3905
rect 2060 -3945 2070 -3905
rect 2010 -3975 2070 -3945
rect 2010 -4015 2020 -3975
rect 2060 -4015 2070 -3975
rect 2010 -4040 2070 -4015
rect 2010 -4080 2020 -4040
rect 2060 -4080 2070 -4040
rect 2010 -4100 2070 -4080
rect 2010 -4140 2020 -4100
rect 2060 -4140 2070 -4100
rect 2010 -4165 2070 -4140
rect 2010 -4205 2020 -4165
rect 2060 -4205 2070 -4165
rect 2010 -4235 2070 -4205
rect 2010 -4275 2020 -4235
rect 2060 -4275 2070 -4235
rect 2010 -4305 2070 -4275
rect 2010 -4345 2020 -4305
rect 2060 -4345 2070 -4305
rect 2010 -4375 2070 -4345
rect 2010 -4415 2020 -4375
rect 2060 -4415 2070 -4375
rect 2010 -4440 2070 -4415
rect 2010 -4480 2020 -4440
rect 2060 -4480 2070 -4440
rect 2010 -4490 2070 -4480
rect 2360 -1300 2420 -1290
rect 2360 -1340 2370 -1300
rect 2410 -1340 2420 -1300
rect 2360 -1365 2420 -1340
rect 2360 -1405 2370 -1365
rect 2410 -1405 2420 -1365
rect 2360 -1435 2420 -1405
rect 2360 -1475 2370 -1435
rect 2410 -1475 2420 -1435
rect 2360 -1505 2420 -1475
rect 2360 -1545 2370 -1505
rect 2410 -1545 2420 -1505
rect 2360 -1575 2420 -1545
rect 2360 -1615 2370 -1575
rect 2410 -1615 2420 -1575
rect 2360 -1640 2420 -1615
rect 2360 -1680 2370 -1640
rect 2410 -1680 2420 -1640
rect 2360 -1700 2420 -1680
rect 2360 -1740 2370 -1700
rect 2410 -1740 2420 -1700
rect 2360 -1765 2420 -1740
rect 2360 -1805 2370 -1765
rect 2410 -1805 2420 -1765
rect 2360 -1835 2420 -1805
rect 2360 -1875 2370 -1835
rect 2410 -1875 2420 -1835
rect 2360 -1905 2420 -1875
rect 2360 -1945 2370 -1905
rect 2410 -1945 2420 -1905
rect 2360 -1975 2420 -1945
rect 2360 -2015 2370 -1975
rect 2410 -2015 2420 -1975
rect 2360 -2040 2420 -2015
rect 2360 -2080 2370 -2040
rect 2410 -2080 2420 -2040
rect 2360 -2100 2420 -2080
rect 2360 -2140 2370 -2100
rect 2410 -2140 2420 -2100
rect 2360 -2165 2420 -2140
rect 2360 -2205 2370 -2165
rect 2410 -2205 2420 -2165
rect 2360 -2235 2420 -2205
rect 2360 -2275 2370 -2235
rect 2410 -2275 2420 -2235
rect 2360 -2305 2420 -2275
rect 2360 -2345 2370 -2305
rect 2410 -2345 2420 -2305
rect 2360 -2375 2420 -2345
rect 2360 -2415 2370 -2375
rect 2410 -2415 2420 -2375
rect 2360 -2440 2420 -2415
rect 2360 -2480 2370 -2440
rect 2410 -2480 2420 -2440
rect 2360 -2500 2420 -2480
rect 2360 -2540 2370 -2500
rect 2410 -2540 2420 -2500
rect 2360 -2565 2420 -2540
rect 2360 -2605 2370 -2565
rect 2410 -2605 2420 -2565
rect 2360 -2635 2420 -2605
rect 2360 -2675 2370 -2635
rect 2410 -2675 2420 -2635
rect 2360 -2705 2420 -2675
rect 2360 -2745 2370 -2705
rect 2410 -2745 2420 -2705
rect 2360 -2775 2420 -2745
rect 2360 -2815 2370 -2775
rect 2410 -2815 2420 -2775
rect 2360 -2840 2420 -2815
rect 2360 -2880 2370 -2840
rect 2410 -2880 2420 -2840
rect 2360 -2900 2420 -2880
rect 2360 -2940 2370 -2900
rect 2410 -2940 2420 -2900
rect 2360 -2965 2420 -2940
rect 2360 -3005 2370 -2965
rect 2410 -3005 2420 -2965
rect 2360 -3035 2420 -3005
rect 2360 -3075 2370 -3035
rect 2410 -3075 2420 -3035
rect 2360 -3105 2420 -3075
rect 2360 -3145 2370 -3105
rect 2410 -3145 2420 -3105
rect 2360 -3175 2420 -3145
rect 2360 -3215 2370 -3175
rect 2410 -3215 2420 -3175
rect 2360 -3240 2420 -3215
rect 2360 -3280 2370 -3240
rect 2410 -3280 2420 -3240
rect 2360 -3300 2420 -3280
rect 2360 -3340 2370 -3300
rect 2410 -3340 2420 -3300
rect 2360 -3365 2420 -3340
rect 2360 -3405 2370 -3365
rect 2410 -3405 2420 -3365
rect 2360 -3435 2420 -3405
rect 2360 -3475 2370 -3435
rect 2410 -3475 2420 -3435
rect 2360 -3505 2420 -3475
rect 2360 -3545 2370 -3505
rect 2410 -3545 2420 -3505
rect 2360 -3575 2420 -3545
rect 2360 -3615 2370 -3575
rect 2410 -3615 2420 -3575
rect 2360 -3640 2420 -3615
rect 2360 -3680 2370 -3640
rect 2410 -3680 2420 -3640
rect 2360 -3700 2420 -3680
rect 2360 -3740 2370 -3700
rect 2410 -3740 2420 -3700
rect 2360 -3765 2420 -3740
rect 2360 -3805 2370 -3765
rect 2410 -3805 2420 -3765
rect 2360 -3835 2420 -3805
rect 2360 -3875 2370 -3835
rect 2410 -3875 2420 -3835
rect 2360 -3905 2420 -3875
rect 2360 -3945 2370 -3905
rect 2410 -3945 2420 -3905
rect 2360 -3975 2420 -3945
rect 2360 -4015 2370 -3975
rect 2410 -4015 2420 -3975
rect 2360 -4040 2420 -4015
rect 2360 -4080 2370 -4040
rect 2410 -4080 2420 -4040
rect 2360 -4100 2420 -4080
rect 2360 -4140 2370 -4100
rect 2410 -4140 2420 -4100
rect 2360 -4165 2420 -4140
rect 2360 -4205 2370 -4165
rect 2410 -4205 2420 -4165
rect 2360 -4235 2420 -4205
rect 2360 -4275 2370 -4235
rect 2410 -4275 2420 -4235
rect 2360 -4305 2420 -4275
rect 2360 -4345 2370 -4305
rect 2410 -4345 2420 -4305
rect 2360 -4375 2420 -4345
rect 2360 -4415 2370 -4375
rect 2410 -4415 2420 -4375
rect 2360 -4440 2420 -4415
rect 2360 -4480 2370 -4440
rect 2410 -4480 2420 -4440
rect 2360 -4490 2420 -4480
rect 2710 -1300 2770 -1290
rect 2710 -1340 2720 -1300
rect 2760 -1340 2770 -1300
rect 2710 -1365 2770 -1340
rect 2710 -1405 2720 -1365
rect 2760 -1405 2770 -1365
rect 2710 -1435 2770 -1405
rect 2710 -1475 2720 -1435
rect 2760 -1475 2770 -1435
rect 2710 -1505 2770 -1475
rect 2710 -1545 2720 -1505
rect 2760 -1545 2770 -1505
rect 2710 -1575 2770 -1545
rect 2710 -1615 2720 -1575
rect 2760 -1615 2770 -1575
rect 2710 -1640 2770 -1615
rect 2710 -1680 2720 -1640
rect 2760 -1680 2770 -1640
rect 2710 -1700 2770 -1680
rect 2710 -1740 2720 -1700
rect 2760 -1740 2770 -1700
rect 2710 -1765 2770 -1740
rect 2710 -1805 2720 -1765
rect 2760 -1805 2770 -1765
rect 2710 -1835 2770 -1805
rect 2710 -1875 2720 -1835
rect 2760 -1875 2770 -1835
rect 2710 -1905 2770 -1875
rect 2710 -1945 2720 -1905
rect 2760 -1945 2770 -1905
rect 2710 -1975 2770 -1945
rect 2710 -2015 2720 -1975
rect 2760 -2015 2770 -1975
rect 2710 -2040 2770 -2015
rect 2710 -2080 2720 -2040
rect 2760 -2080 2770 -2040
rect 2710 -2100 2770 -2080
rect 2710 -2140 2720 -2100
rect 2760 -2140 2770 -2100
rect 2710 -2165 2770 -2140
rect 2710 -2205 2720 -2165
rect 2760 -2205 2770 -2165
rect 2710 -2235 2770 -2205
rect 2710 -2275 2720 -2235
rect 2760 -2275 2770 -2235
rect 2710 -2305 2770 -2275
rect 2710 -2345 2720 -2305
rect 2760 -2345 2770 -2305
rect 2710 -2375 2770 -2345
rect 2710 -2415 2720 -2375
rect 2760 -2415 2770 -2375
rect 2710 -2440 2770 -2415
rect 2710 -2480 2720 -2440
rect 2760 -2480 2770 -2440
rect 2710 -2500 2770 -2480
rect 2710 -2540 2720 -2500
rect 2760 -2540 2770 -2500
rect 2710 -2565 2770 -2540
rect 2710 -2605 2720 -2565
rect 2760 -2605 2770 -2565
rect 2710 -2635 2770 -2605
rect 2710 -2675 2720 -2635
rect 2760 -2675 2770 -2635
rect 2710 -2705 2770 -2675
rect 2710 -2745 2720 -2705
rect 2760 -2745 2770 -2705
rect 2710 -2775 2770 -2745
rect 2710 -2815 2720 -2775
rect 2760 -2815 2770 -2775
rect 2710 -2840 2770 -2815
rect 2710 -2880 2720 -2840
rect 2760 -2880 2770 -2840
rect 2710 -2900 2770 -2880
rect 2710 -2940 2720 -2900
rect 2760 -2940 2770 -2900
rect 2710 -2965 2770 -2940
rect 2710 -3005 2720 -2965
rect 2760 -3005 2770 -2965
rect 2710 -3035 2770 -3005
rect 2710 -3075 2720 -3035
rect 2760 -3075 2770 -3035
rect 2710 -3105 2770 -3075
rect 2710 -3145 2720 -3105
rect 2760 -3145 2770 -3105
rect 2710 -3175 2770 -3145
rect 2710 -3215 2720 -3175
rect 2760 -3215 2770 -3175
rect 2710 -3240 2770 -3215
rect 2710 -3280 2720 -3240
rect 2760 -3280 2770 -3240
rect 2710 -3300 2770 -3280
rect 2710 -3340 2720 -3300
rect 2760 -3340 2770 -3300
rect 2710 -3365 2770 -3340
rect 2710 -3405 2720 -3365
rect 2760 -3405 2770 -3365
rect 2710 -3435 2770 -3405
rect 2710 -3475 2720 -3435
rect 2760 -3475 2770 -3435
rect 2710 -3505 2770 -3475
rect 2710 -3545 2720 -3505
rect 2760 -3545 2770 -3505
rect 2710 -3575 2770 -3545
rect 2710 -3615 2720 -3575
rect 2760 -3615 2770 -3575
rect 2710 -3640 2770 -3615
rect 2710 -3680 2720 -3640
rect 2760 -3680 2770 -3640
rect 2710 -3700 2770 -3680
rect 2710 -3740 2720 -3700
rect 2760 -3740 2770 -3700
rect 2710 -3765 2770 -3740
rect 2710 -3805 2720 -3765
rect 2760 -3805 2770 -3765
rect 2710 -3835 2770 -3805
rect 2710 -3875 2720 -3835
rect 2760 -3875 2770 -3835
rect 2710 -3905 2770 -3875
rect 2710 -3945 2720 -3905
rect 2760 -3945 2770 -3905
rect 2710 -3975 2770 -3945
rect 2710 -4015 2720 -3975
rect 2760 -4015 2770 -3975
rect 2710 -4040 2770 -4015
rect 2710 -4080 2720 -4040
rect 2760 -4080 2770 -4040
rect 2710 -4100 2770 -4080
rect 2710 -4140 2720 -4100
rect 2760 -4140 2770 -4100
rect 2710 -4165 2770 -4140
rect 2710 -4205 2720 -4165
rect 2760 -4205 2770 -4165
rect 2710 -4235 2770 -4205
rect 2710 -4275 2720 -4235
rect 2760 -4275 2770 -4235
rect 2710 -4305 2770 -4275
rect 2710 -4345 2720 -4305
rect 2760 -4345 2770 -4305
rect 2710 -4375 2770 -4345
rect 2710 -4415 2720 -4375
rect 2760 -4415 2770 -4375
rect 2710 -4440 2770 -4415
rect 2710 -4480 2720 -4440
rect 2760 -4480 2770 -4440
rect 2710 -4490 2770 -4480
rect 3060 -1300 3120 -1290
rect 3060 -1340 3070 -1300
rect 3110 -1340 3120 -1300
rect 3060 -1365 3120 -1340
rect 3060 -1405 3070 -1365
rect 3110 -1405 3120 -1365
rect 3060 -1435 3120 -1405
rect 3060 -1475 3070 -1435
rect 3110 -1475 3120 -1435
rect 3060 -1505 3120 -1475
rect 3060 -1545 3070 -1505
rect 3110 -1545 3120 -1505
rect 3060 -1575 3120 -1545
rect 3060 -1615 3070 -1575
rect 3110 -1615 3120 -1575
rect 3060 -1640 3120 -1615
rect 3060 -1680 3070 -1640
rect 3110 -1680 3120 -1640
rect 3060 -1700 3120 -1680
rect 3060 -1740 3070 -1700
rect 3110 -1740 3120 -1700
rect 3060 -1765 3120 -1740
rect 3060 -1805 3070 -1765
rect 3110 -1805 3120 -1765
rect 3060 -1835 3120 -1805
rect 3060 -1875 3070 -1835
rect 3110 -1875 3120 -1835
rect 3060 -1905 3120 -1875
rect 3060 -1945 3070 -1905
rect 3110 -1945 3120 -1905
rect 3060 -1975 3120 -1945
rect 3060 -2015 3070 -1975
rect 3110 -2015 3120 -1975
rect 3060 -2040 3120 -2015
rect 3060 -2080 3070 -2040
rect 3110 -2080 3120 -2040
rect 3060 -2100 3120 -2080
rect 3060 -2140 3070 -2100
rect 3110 -2140 3120 -2100
rect 3060 -2165 3120 -2140
rect 3060 -2205 3070 -2165
rect 3110 -2205 3120 -2165
rect 3060 -2235 3120 -2205
rect 3060 -2275 3070 -2235
rect 3110 -2275 3120 -2235
rect 3060 -2305 3120 -2275
rect 3060 -2345 3070 -2305
rect 3110 -2345 3120 -2305
rect 3060 -2375 3120 -2345
rect 3060 -2415 3070 -2375
rect 3110 -2415 3120 -2375
rect 3060 -2440 3120 -2415
rect 3060 -2480 3070 -2440
rect 3110 -2480 3120 -2440
rect 3060 -2500 3120 -2480
rect 3060 -2540 3070 -2500
rect 3110 -2540 3120 -2500
rect 3060 -2565 3120 -2540
rect 3060 -2605 3070 -2565
rect 3110 -2605 3120 -2565
rect 3060 -2635 3120 -2605
rect 3060 -2675 3070 -2635
rect 3110 -2675 3120 -2635
rect 3060 -2705 3120 -2675
rect 3060 -2745 3070 -2705
rect 3110 -2745 3120 -2705
rect 3060 -2775 3120 -2745
rect 3060 -2815 3070 -2775
rect 3110 -2815 3120 -2775
rect 3060 -2840 3120 -2815
rect 3060 -2880 3070 -2840
rect 3110 -2880 3120 -2840
rect 3060 -2900 3120 -2880
rect 3060 -2940 3070 -2900
rect 3110 -2940 3120 -2900
rect 3060 -2965 3120 -2940
rect 3060 -3005 3070 -2965
rect 3110 -3005 3120 -2965
rect 3060 -3035 3120 -3005
rect 3060 -3075 3070 -3035
rect 3110 -3075 3120 -3035
rect 3060 -3105 3120 -3075
rect 3060 -3145 3070 -3105
rect 3110 -3145 3120 -3105
rect 3060 -3175 3120 -3145
rect 3060 -3215 3070 -3175
rect 3110 -3215 3120 -3175
rect 3060 -3240 3120 -3215
rect 3060 -3280 3070 -3240
rect 3110 -3280 3120 -3240
rect 3060 -3300 3120 -3280
rect 3060 -3340 3070 -3300
rect 3110 -3340 3120 -3300
rect 3060 -3365 3120 -3340
rect 3060 -3405 3070 -3365
rect 3110 -3405 3120 -3365
rect 3060 -3435 3120 -3405
rect 3060 -3475 3070 -3435
rect 3110 -3475 3120 -3435
rect 3060 -3505 3120 -3475
rect 3060 -3545 3070 -3505
rect 3110 -3545 3120 -3505
rect 3060 -3575 3120 -3545
rect 3060 -3615 3070 -3575
rect 3110 -3615 3120 -3575
rect 3060 -3640 3120 -3615
rect 3060 -3680 3070 -3640
rect 3110 -3680 3120 -3640
rect 3060 -3700 3120 -3680
rect 3060 -3740 3070 -3700
rect 3110 -3740 3120 -3700
rect 3060 -3765 3120 -3740
rect 3060 -3805 3070 -3765
rect 3110 -3805 3120 -3765
rect 3060 -3835 3120 -3805
rect 3060 -3875 3070 -3835
rect 3110 -3875 3120 -3835
rect 3060 -3905 3120 -3875
rect 3060 -3945 3070 -3905
rect 3110 -3945 3120 -3905
rect 3060 -3975 3120 -3945
rect 3060 -4015 3070 -3975
rect 3110 -4015 3120 -3975
rect 3060 -4040 3120 -4015
rect 3060 -4080 3070 -4040
rect 3110 -4080 3120 -4040
rect 3060 -4100 3120 -4080
rect 3060 -4140 3070 -4100
rect 3110 -4140 3120 -4100
rect 3060 -4165 3120 -4140
rect 3060 -4205 3070 -4165
rect 3110 -4205 3120 -4165
rect 3060 -4235 3120 -4205
rect 3060 -4275 3070 -4235
rect 3110 -4275 3120 -4235
rect 3060 -4305 3120 -4275
rect 3060 -4345 3070 -4305
rect 3110 -4345 3120 -4305
rect 3060 -4375 3120 -4345
rect 3060 -4415 3070 -4375
rect 3110 -4415 3120 -4375
rect 3060 -4440 3120 -4415
rect 3060 -4480 3070 -4440
rect 3110 -4480 3120 -4440
rect 3060 -4490 3120 -4480
rect 3410 -1300 3470 -1290
rect 3410 -1340 3420 -1300
rect 3460 -1340 3470 -1300
rect 3410 -1365 3470 -1340
rect 3410 -1405 3420 -1365
rect 3460 -1405 3470 -1365
rect 3410 -1435 3470 -1405
rect 3410 -1475 3420 -1435
rect 3460 -1475 3470 -1435
rect 3410 -1505 3470 -1475
rect 3410 -1545 3420 -1505
rect 3460 -1545 3470 -1505
rect 3410 -1575 3470 -1545
rect 3410 -1615 3420 -1575
rect 3460 -1615 3470 -1575
rect 3410 -1640 3470 -1615
rect 3410 -1680 3420 -1640
rect 3460 -1680 3470 -1640
rect 3410 -1700 3470 -1680
rect 3410 -1740 3420 -1700
rect 3460 -1740 3470 -1700
rect 3410 -1765 3470 -1740
rect 3410 -1805 3420 -1765
rect 3460 -1805 3470 -1765
rect 3410 -1835 3470 -1805
rect 3410 -1875 3420 -1835
rect 3460 -1875 3470 -1835
rect 3410 -1905 3470 -1875
rect 3410 -1945 3420 -1905
rect 3460 -1945 3470 -1905
rect 3410 -1975 3470 -1945
rect 3410 -2015 3420 -1975
rect 3460 -2015 3470 -1975
rect 3410 -2040 3470 -2015
rect 3410 -2080 3420 -2040
rect 3460 -2080 3470 -2040
rect 3410 -2100 3470 -2080
rect 3410 -2140 3420 -2100
rect 3460 -2140 3470 -2100
rect 3410 -2165 3470 -2140
rect 3410 -2205 3420 -2165
rect 3460 -2205 3470 -2165
rect 3410 -2235 3470 -2205
rect 3410 -2275 3420 -2235
rect 3460 -2275 3470 -2235
rect 3410 -2305 3470 -2275
rect 3410 -2345 3420 -2305
rect 3460 -2345 3470 -2305
rect 3410 -2375 3470 -2345
rect 3410 -2415 3420 -2375
rect 3460 -2415 3470 -2375
rect 3410 -2440 3470 -2415
rect 3410 -2480 3420 -2440
rect 3460 -2480 3470 -2440
rect 3410 -2500 3470 -2480
rect 3410 -2540 3420 -2500
rect 3460 -2540 3470 -2500
rect 3410 -2565 3470 -2540
rect 3410 -2605 3420 -2565
rect 3460 -2605 3470 -2565
rect 3410 -2635 3470 -2605
rect 3410 -2675 3420 -2635
rect 3460 -2675 3470 -2635
rect 3410 -2705 3470 -2675
rect 3410 -2745 3420 -2705
rect 3460 -2745 3470 -2705
rect 3410 -2775 3470 -2745
rect 3410 -2815 3420 -2775
rect 3460 -2815 3470 -2775
rect 3410 -2840 3470 -2815
rect 3410 -2880 3420 -2840
rect 3460 -2880 3470 -2840
rect 3410 -2900 3470 -2880
rect 3410 -2940 3420 -2900
rect 3460 -2940 3470 -2900
rect 3410 -2965 3470 -2940
rect 3410 -3005 3420 -2965
rect 3460 -3005 3470 -2965
rect 3410 -3035 3470 -3005
rect 3410 -3075 3420 -3035
rect 3460 -3075 3470 -3035
rect 3410 -3105 3470 -3075
rect 3410 -3145 3420 -3105
rect 3460 -3145 3470 -3105
rect 3410 -3175 3470 -3145
rect 3410 -3215 3420 -3175
rect 3460 -3215 3470 -3175
rect 3410 -3240 3470 -3215
rect 3410 -3280 3420 -3240
rect 3460 -3280 3470 -3240
rect 3410 -3300 3470 -3280
rect 3410 -3340 3420 -3300
rect 3460 -3340 3470 -3300
rect 3410 -3365 3470 -3340
rect 3410 -3405 3420 -3365
rect 3460 -3405 3470 -3365
rect 3410 -3435 3470 -3405
rect 3410 -3475 3420 -3435
rect 3460 -3475 3470 -3435
rect 3410 -3505 3470 -3475
rect 3410 -3545 3420 -3505
rect 3460 -3545 3470 -3505
rect 3410 -3575 3470 -3545
rect 3410 -3615 3420 -3575
rect 3460 -3615 3470 -3575
rect 3410 -3640 3470 -3615
rect 3410 -3680 3420 -3640
rect 3460 -3680 3470 -3640
rect 3410 -3700 3470 -3680
rect 3410 -3740 3420 -3700
rect 3460 -3740 3470 -3700
rect 3410 -3765 3470 -3740
rect 3410 -3805 3420 -3765
rect 3460 -3805 3470 -3765
rect 3410 -3835 3470 -3805
rect 3410 -3875 3420 -3835
rect 3460 -3875 3470 -3835
rect 3410 -3905 3470 -3875
rect 3410 -3945 3420 -3905
rect 3460 -3945 3470 -3905
rect 3410 -3975 3470 -3945
rect 3410 -4015 3420 -3975
rect 3460 -4015 3470 -3975
rect 3410 -4040 3470 -4015
rect 3410 -4080 3420 -4040
rect 3460 -4080 3470 -4040
rect 3410 -4100 3470 -4080
rect 3410 -4140 3420 -4100
rect 3460 -4140 3470 -4100
rect 3410 -4165 3470 -4140
rect 3410 -4205 3420 -4165
rect 3460 -4205 3470 -4165
rect 3410 -4235 3470 -4205
rect 3410 -4275 3420 -4235
rect 3460 -4275 3470 -4235
rect 3410 -4305 3470 -4275
rect 3410 -4345 3420 -4305
rect 3460 -4345 3470 -4305
rect 3410 -4375 3470 -4345
rect 3410 -4415 3420 -4375
rect 3460 -4415 3470 -4375
rect 3410 -4440 3470 -4415
rect 3410 -4480 3420 -4440
rect 3460 -4480 3470 -4440
rect 3410 -4490 3470 -4480
rect 3760 -1300 3820 -1290
rect 3760 -1340 3770 -1300
rect 3810 -1340 3820 -1300
rect 3760 -1365 3820 -1340
rect 3760 -1405 3770 -1365
rect 3810 -1405 3820 -1365
rect 3760 -1435 3820 -1405
rect 3760 -1475 3770 -1435
rect 3810 -1475 3820 -1435
rect 3760 -1505 3820 -1475
rect 3760 -1545 3770 -1505
rect 3810 -1545 3820 -1505
rect 3760 -1575 3820 -1545
rect 3760 -1615 3770 -1575
rect 3810 -1615 3820 -1575
rect 3760 -1640 3820 -1615
rect 3760 -1680 3770 -1640
rect 3810 -1680 3820 -1640
rect 3760 -1700 3820 -1680
rect 3760 -1740 3770 -1700
rect 3810 -1740 3820 -1700
rect 3760 -1765 3820 -1740
rect 3760 -1805 3770 -1765
rect 3810 -1805 3820 -1765
rect 3760 -1835 3820 -1805
rect 3760 -1875 3770 -1835
rect 3810 -1875 3820 -1835
rect 3760 -1905 3820 -1875
rect 3760 -1945 3770 -1905
rect 3810 -1945 3820 -1905
rect 3760 -1975 3820 -1945
rect 3760 -2015 3770 -1975
rect 3810 -2015 3820 -1975
rect 3760 -2040 3820 -2015
rect 3760 -2080 3770 -2040
rect 3810 -2080 3820 -2040
rect 3760 -2100 3820 -2080
rect 3760 -2140 3770 -2100
rect 3810 -2140 3820 -2100
rect 3760 -2165 3820 -2140
rect 3760 -2205 3770 -2165
rect 3810 -2205 3820 -2165
rect 3760 -2235 3820 -2205
rect 3760 -2275 3770 -2235
rect 3810 -2275 3820 -2235
rect 3760 -2305 3820 -2275
rect 3760 -2345 3770 -2305
rect 3810 -2345 3820 -2305
rect 3760 -2375 3820 -2345
rect 3760 -2415 3770 -2375
rect 3810 -2415 3820 -2375
rect 3760 -2440 3820 -2415
rect 3760 -2480 3770 -2440
rect 3810 -2480 3820 -2440
rect 3760 -2500 3820 -2480
rect 3760 -2540 3770 -2500
rect 3810 -2540 3820 -2500
rect 3760 -2565 3820 -2540
rect 3760 -2605 3770 -2565
rect 3810 -2605 3820 -2565
rect 3760 -2635 3820 -2605
rect 3760 -2675 3770 -2635
rect 3810 -2675 3820 -2635
rect 3760 -2705 3820 -2675
rect 3760 -2745 3770 -2705
rect 3810 -2745 3820 -2705
rect 3760 -2775 3820 -2745
rect 3760 -2815 3770 -2775
rect 3810 -2815 3820 -2775
rect 3760 -2840 3820 -2815
rect 3760 -2880 3770 -2840
rect 3810 -2880 3820 -2840
rect 3760 -2900 3820 -2880
rect 3760 -2940 3770 -2900
rect 3810 -2940 3820 -2900
rect 3760 -2965 3820 -2940
rect 3760 -3005 3770 -2965
rect 3810 -3005 3820 -2965
rect 3760 -3035 3820 -3005
rect 3760 -3075 3770 -3035
rect 3810 -3075 3820 -3035
rect 3760 -3105 3820 -3075
rect 3760 -3145 3770 -3105
rect 3810 -3145 3820 -3105
rect 3760 -3175 3820 -3145
rect 3760 -3215 3770 -3175
rect 3810 -3215 3820 -3175
rect 3760 -3240 3820 -3215
rect 3760 -3280 3770 -3240
rect 3810 -3280 3820 -3240
rect 3760 -3300 3820 -3280
rect 3760 -3340 3770 -3300
rect 3810 -3340 3820 -3300
rect 3760 -3365 3820 -3340
rect 3760 -3405 3770 -3365
rect 3810 -3405 3820 -3365
rect 3760 -3435 3820 -3405
rect 3760 -3475 3770 -3435
rect 3810 -3475 3820 -3435
rect 3760 -3505 3820 -3475
rect 3760 -3545 3770 -3505
rect 3810 -3545 3820 -3505
rect 3760 -3575 3820 -3545
rect 3760 -3615 3770 -3575
rect 3810 -3615 3820 -3575
rect 3760 -3640 3820 -3615
rect 3760 -3680 3770 -3640
rect 3810 -3680 3820 -3640
rect 3760 -3700 3820 -3680
rect 3760 -3740 3770 -3700
rect 3810 -3740 3820 -3700
rect 3760 -3765 3820 -3740
rect 3760 -3805 3770 -3765
rect 3810 -3805 3820 -3765
rect 3760 -3835 3820 -3805
rect 3760 -3875 3770 -3835
rect 3810 -3875 3820 -3835
rect 3760 -3905 3820 -3875
rect 3760 -3945 3770 -3905
rect 3810 -3945 3820 -3905
rect 3760 -3975 3820 -3945
rect 3760 -4015 3770 -3975
rect 3810 -4015 3820 -3975
rect 3760 -4040 3820 -4015
rect 3760 -4080 3770 -4040
rect 3810 -4080 3820 -4040
rect 3760 -4100 3820 -4080
rect 3760 -4140 3770 -4100
rect 3810 -4140 3820 -4100
rect 3760 -4165 3820 -4140
rect 3760 -4205 3770 -4165
rect 3810 -4205 3820 -4165
rect 3760 -4235 3820 -4205
rect 3760 -4275 3770 -4235
rect 3810 -4275 3820 -4235
rect 3760 -4305 3820 -4275
rect 3760 -4345 3770 -4305
rect 3810 -4345 3820 -4305
rect 3760 -4375 3820 -4345
rect 3760 -4415 3770 -4375
rect 3810 -4415 3820 -4375
rect 3760 -4440 3820 -4415
rect 3760 -4480 3770 -4440
rect 3810 -4480 3820 -4440
rect 3760 -4490 3820 -4480
rect 4110 -1300 4170 -1290
rect 4110 -1340 4120 -1300
rect 4160 -1340 4170 -1300
rect 4110 -1365 4170 -1340
rect 4110 -1405 4120 -1365
rect 4160 -1405 4170 -1365
rect 4110 -1435 4170 -1405
rect 4110 -1475 4120 -1435
rect 4160 -1475 4170 -1435
rect 4110 -1505 4170 -1475
rect 4110 -1545 4120 -1505
rect 4160 -1545 4170 -1505
rect 4110 -1575 4170 -1545
rect 4110 -1615 4120 -1575
rect 4160 -1615 4170 -1575
rect 4110 -1640 4170 -1615
rect 4110 -1680 4120 -1640
rect 4160 -1680 4170 -1640
rect 4110 -1700 4170 -1680
rect 4110 -1740 4120 -1700
rect 4160 -1740 4170 -1700
rect 4110 -1765 4170 -1740
rect 4110 -1805 4120 -1765
rect 4160 -1805 4170 -1765
rect 4110 -1835 4170 -1805
rect 4110 -1875 4120 -1835
rect 4160 -1875 4170 -1835
rect 4110 -1905 4170 -1875
rect 4110 -1945 4120 -1905
rect 4160 -1945 4170 -1905
rect 4110 -1975 4170 -1945
rect 4110 -2015 4120 -1975
rect 4160 -2015 4170 -1975
rect 4110 -2040 4170 -2015
rect 4110 -2080 4120 -2040
rect 4160 -2080 4170 -2040
rect 4110 -2100 4170 -2080
rect 4110 -2140 4120 -2100
rect 4160 -2140 4170 -2100
rect 4110 -2165 4170 -2140
rect 4110 -2205 4120 -2165
rect 4160 -2205 4170 -2165
rect 4110 -2235 4170 -2205
rect 4110 -2275 4120 -2235
rect 4160 -2275 4170 -2235
rect 4110 -2305 4170 -2275
rect 4110 -2345 4120 -2305
rect 4160 -2345 4170 -2305
rect 4110 -2375 4170 -2345
rect 4110 -2415 4120 -2375
rect 4160 -2415 4170 -2375
rect 4110 -2440 4170 -2415
rect 4110 -2480 4120 -2440
rect 4160 -2480 4170 -2440
rect 4110 -2500 4170 -2480
rect 4110 -2540 4120 -2500
rect 4160 -2540 4170 -2500
rect 4110 -2565 4170 -2540
rect 4110 -2605 4120 -2565
rect 4160 -2605 4170 -2565
rect 4110 -2635 4170 -2605
rect 4110 -2675 4120 -2635
rect 4160 -2675 4170 -2635
rect 4110 -2705 4170 -2675
rect 4110 -2745 4120 -2705
rect 4160 -2745 4170 -2705
rect 4110 -2775 4170 -2745
rect 4110 -2815 4120 -2775
rect 4160 -2815 4170 -2775
rect 4110 -2840 4170 -2815
rect 4110 -2880 4120 -2840
rect 4160 -2880 4170 -2840
rect 4110 -2900 4170 -2880
rect 4110 -2940 4120 -2900
rect 4160 -2940 4170 -2900
rect 4110 -2965 4170 -2940
rect 4110 -3005 4120 -2965
rect 4160 -3005 4170 -2965
rect 4110 -3035 4170 -3005
rect 4110 -3075 4120 -3035
rect 4160 -3075 4170 -3035
rect 4110 -3105 4170 -3075
rect 4110 -3145 4120 -3105
rect 4160 -3145 4170 -3105
rect 4110 -3175 4170 -3145
rect 4110 -3215 4120 -3175
rect 4160 -3215 4170 -3175
rect 4110 -3240 4170 -3215
rect 4110 -3280 4120 -3240
rect 4160 -3280 4170 -3240
rect 4110 -3300 4170 -3280
rect 4110 -3340 4120 -3300
rect 4160 -3340 4170 -3300
rect 4110 -3365 4170 -3340
rect 4110 -3405 4120 -3365
rect 4160 -3405 4170 -3365
rect 4110 -3435 4170 -3405
rect 4110 -3475 4120 -3435
rect 4160 -3475 4170 -3435
rect 4110 -3505 4170 -3475
rect 4110 -3545 4120 -3505
rect 4160 -3545 4170 -3505
rect 4110 -3575 4170 -3545
rect 4110 -3615 4120 -3575
rect 4160 -3615 4170 -3575
rect 4110 -3640 4170 -3615
rect 4110 -3680 4120 -3640
rect 4160 -3680 4170 -3640
rect 4110 -3700 4170 -3680
rect 4110 -3740 4120 -3700
rect 4160 -3740 4170 -3700
rect 4110 -3765 4170 -3740
rect 4110 -3805 4120 -3765
rect 4160 -3805 4170 -3765
rect 4110 -3835 4170 -3805
rect 4110 -3875 4120 -3835
rect 4160 -3875 4170 -3835
rect 4110 -3905 4170 -3875
rect 4110 -3945 4120 -3905
rect 4160 -3945 4170 -3905
rect 4110 -3975 4170 -3945
rect 4110 -4015 4120 -3975
rect 4160 -4015 4170 -3975
rect 4110 -4040 4170 -4015
rect 4110 -4080 4120 -4040
rect 4160 -4080 4170 -4040
rect 4110 -4100 4170 -4080
rect 4110 -4140 4120 -4100
rect 4160 -4140 4170 -4100
rect 4110 -4165 4170 -4140
rect 4110 -4205 4120 -4165
rect 4160 -4205 4170 -4165
rect 4110 -4235 4170 -4205
rect 4110 -4275 4120 -4235
rect 4160 -4275 4170 -4235
rect 4110 -4305 4170 -4275
rect 4110 -4345 4120 -4305
rect 4160 -4345 4170 -4305
rect 4110 -4375 4170 -4345
rect 4110 -4415 4120 -4375
rect 4160 -4415 4170 -4375
rect 4110 -4440 4170 -4415
rect 4110 -4480 4120 -4440
rect 4160 -4480 4170 -4440
rect 4110 -4490 4170 -4480
rect 4460 -1300 4520 -1290
rect 4460 -1340 4470 -1300
rect 4510 -1340 4520 -1300
rect 4460 -1365 4520 -1340
rect 4460 -1405 4470 -1365
rect 4510 -1405 4520 -1365
rect 4460 -1435 4520 -1405
rect 4460 -1475 4470 -1435
rect 4510 -1475 4520 -1435
rect 4460 -1505 4520 -1475
rect 4460 -1545 4470 -1505
rect 4510 -1545 4520 -1505
rect 4460 -1575 4520 -1545
rect 4460 -1615 4470 -1575
rect 4510 -1615 4520 -1575
rect 4460 -1640 4520 -1615
rect 4460 -1680 4470 -1640
rect 4510 -1680 4520 -1640
rect 4460 -1700 4520 -1680
rect 4460 -1740 4470 -1700
rect 4510 -1740 4520 -1700
rect 4460 -1765 4520 -1740
rect 4460 -1805 4470 -1765
rect 4510 -1805 4520 -1765
rect 4460 -1835 4520 -1805
rect 4460 -1875 4470 -1835
rect 4510 -1875 4520 -1835
rect 4460 -1905 4520 -1875
rect 4460 -1945 4470 -1905
rect 4510 -1945 4520 -1905
rect 4460 -1975 4520 -1945
rect 4460 -2015 4470 -1975
rect 4510 -2015 4520 -1975
rect 4460 -2040 4520 -2015
rect 4460 -2080 4470 -2040
rect 4510 -2080 4520 -2040
rect 4460 -2100 4520 -2080
rect 4460 -2140 4470 -2100
rect 4510 -2140 4520 -2100
rect 4460 -2165 4520 -2140
rect 4460 -2205 4470 -2165
rect 4510 -2205 4520 -2165
rect 4460 -2235 4520 -2205
rect 4460 -2275 4470 -2235
rect 4510 -2275 4520 -2235
rect 4460 -2305 4520 -2275
rect 4460 -2345 4470 -2305
rect 4510 -2345 4520 -2305
rect 4460 -2375 4520 -2345
rect 4460 -2415 4470 -2375
rect 4510 -2415 4520 -2375
rect 4460 -2440 4520 -2415
rect 4460 -2480 4470 -2440
rect 4510 -2480 4520 -2440
rect 4460 -2500 4520 -2480
rect 4460 -2540 4470 -2500
rect 4510 -2540 4520 -2500
rect 4460 -2565 4520 -2540
rect 4460 -2605 4470 -2565
rect 4510 -2605 4520 -2565
rect 4460 -2635 4520 -2605
rect 4460 -2675 4470 -2635
rect 4510 -2675 4520 -2635
rect 4460 -2705 4520 -2675
rect 4460 -2745 4470 -2705
rect 4510 -2745 4520 -2705
rect 4460 -2775 4520 -2745
rect 4460 -2815 4470 -2775
rect 4510 -2815 4520 -2775
rect 4460 -2840 4520 -2815
rect 4460 -2880 4470 -2840
rect 4510 -2880 4520 -2840
rect 4460 -2900 4520 -2880
rect 4460 -2940 4470 -2900
rect 4510 -2940 4520 -2900
rect 4460 -2965 4520 -2940
rect 4460 -3005 4470 -2965
rect 4510 -3005 4520 -2965
rect 4460 -3035 4520 -3005
rect 4460 -3075 4470 -3035
rect 4510 -3075 4520 -3035
rect 4460 -3105 4520 -3075
rect 4460 -3145 4470 -3105
rect 4510 -3145 4520 -3105
rect 4460 -3175 4520 -3145
rect 4460 -3215 4470 -3175
rect 4510 -3215 4520 -3175
rect 4460 -3240 4520 -3215
rect 4460 -3280 4470 -3240
rect 4510 -3280 4520 -3240
rect 4460 -3300 4520 -3280
rect 4460 -3340 4470 -3300
rect 4510 -3340 4520 -3300
rect 4460 -3365 4520 -3340
rect 4460 -3405 4470 -3365
rect 4510 -3405 4520 -3365
rect 4460 -3435 4520 -3405
rect 4460 -3475 4470 -3435
rect 4510 -3475 4520 -3435
rect 4460 -3505 4520 -3475
rect 4460 -3545 4470 -3505
rect 4510 -3545 4520 -3505
rect 4460 -3575 4520 -3545
rect 4460 -3615 4470 -3575
rect 4510 -3615 4520 -3575
rect 4460 -3640 4520 -3615
rect 4460 -3680 4470 -3640
rect 4510 -3680 4520 -3640
rect 4460 -3700 4520 -3680
rect 4460 -3740 4470 -3700
rect 4510 -3740 4520 -3700
rect 4460 -3765 4520 -3740
rect 4460 -3805 4470 -3765
rect 4510 -3805 4520 -3765
rect 4460 -3835 4520 -3805
rect 4460 -3875 4470 -3835
rect 4510 -3875 4520 -3835
rect 4460 -3905 4520 -3875
rect 4460 -3945 4470 -3905
rect 4510 -3945 4520 -3905
rect 4460 -3975 4520 -3945
rect 4460 -4015 4470 -3975
rect 4510 -4015 4520 -3975
rect 4460 -4040 4520 -4015
rect 4460 -4080 4470 -4040
rect 4510 -4080 4520 -4040
rect 4460 -4100 4520 -4080
rect 4460 -4140 4470 -4100
rect 4510 -4140 4520 -4100
rect 4460 -4165 4520 -4140
rect 4460 -4205 4470 -4165
rect 4510 -4205 4520 -4165
rect 4460 -4235 4520 -4205
rect 4460 -4275 4470 -4235
rect 4510 -4275 4520 -4235
rect 4460 -4305 4520 -4275
rect 4460 -4345 4470 -4305
rect 4510 -4345 4520 -4305
rect 4460 -4375 4520 -4345
rect 4460 -4415 4470 -4375
rect 4510 -4415 4520 -4375
rect 4460 -4440 4520 -4415
rect 4460 -4480 4470 -4440
rect 4510 -4480 4520 -4440
rect 4460 -4490 4520 -4480
rect 4810 -1300 4870 -1290
rect 4810 -1340 4820 -1300
rect 4860 -1340 4870 -1300
rect 4810 -1365 4870 -1340
rect 4810 -1405 4820 -1365
rect 4860 -1405 4870 -1365
rect 4810 -1435 4870 -1405
rect 4810 -1475 4820 -1435
rect 4860 -1475 4870 -1435
rect 4810 -1505 4870 -1475
rect 4810 -1545 4820 -1505
rect 4860 -1545 4870 -1505
rect 4810 -1575 4870 -1545
rect 4810 -1615 4820 -1575
rect 4860 -1615 4870 -1575
rect 4810 -1640 4870 -1615
rect 4810 -1680 4820 -1640
rect 4860 -1680 4870 -1640
rect 4810 -1700 4870 -1680
rect 4810 -1740 4820 -1700
rect 4860 -1740 4870 -1700
rect 4810 -1765 4870 -1740
rect 4810 -1805 4820 -1765
rect 4860 -1805 4870 -1765
rect 4810 -1835 4870 -1805
rect 4810 -1875 4820 -1835
rect 4860 -1875 4870 -1835
rect 4810 -1905 4870 -1875
rect 4810 -1945 4820 -1905
rect 4860 -1945 4870 -1905
rect 4810 -1975 4870 -1945
rect 4810 -2015 4820 -1975
rect 4860 -2015 4870 -1975
rect 4810 -2040 4870 -2015
rect 4810 -2080 4820 -2040
rect 4860 -2080 4870 -2040
rect 4810 -2100 4870 -2080
rect 4810 -2140 4820 -2100
rect 4860 -2140 4870 -2100
rect 4810 -2165 4870 -2140
rect 4810 -2205 4820 -2165
rect 4860 -2205 4870 -2165
rect 4810 -2235 4870 -2205
rect 4810 -2275 4820 -2235
rect 4860 -2275 4870 -2235
rect 4810 -2305 4870 -2275
rect 4810 -2345 4820 -2305
rect 4860 -2345 4870 -2305
rect 4810 -2375 4870 -2345
rect 4810 -2415 4820 -2375
rect 4860 -2415 4870 -2375
rect 4810 -2440 4870 -2415
rect 4810 -2480 4820 -2440
rect 4860 -2480 4870 -2440
rect 4810 -2500 4870 -2480
rect 4810 -2540 4820 -2500
rect 4860 -2540 4870 -2500
rect 4810 -2565 4870 -2540
rect 4810 -2605 4820 -2565
rect 4860 -2605 4870 -2565
rect 4810 -2635 4870 -2605
rect 4810 -2675 4820 -2635
rect 4860 -2675 4870 -2635
rect 4810 -2705 4870 -2675
rect 4810 -2745 4820 -2705
rect 4860 -2745 4870 -2705
rect 4810 -2775 4870 -2745
rect 4810 -2815 4820 -2775
rect 4860 -2815 4870 -2775
rect 4810 -2840 4870 -2815
rect 4810 -2880 4820 -2840
rect 4860 -2880 4870 -2840
rect 4810 -2900 4870 -2880
rect 4810 -2940 4820 -2900
rect 4860 -2940 4870 -2900
rect 4810 -2965 4870 -2940
rect 4810 -3005 4820 -2965
rect 4860 -3005 4870 -2965
rect 4810 -3035 4870 -3005
rect 4810 -3075 4820 -3035
rect 4860 -3075 4870 -3035
rect 4810 -3105 4870 -3075
rect 4810 -3145 4820 -3105
rect 4860 -3145 4870 -3105
rect 4810 -3175 4870 -3145
rect 4810 -3215 4820 -3175
rect 4860 -3215 4870 -3175
rect 4810 -3240 4870 -3215
rect 4810 -3280 4820 -3240
rect 4860 -3280 4870 -3240
rect 4810 -3300 4870 -3280
rect 4810 -3340 4820 -3300
rect 4860 -3340 4870 -3300
rect 4810 -3365 4870 -3340
rect 4810 -3405 4820 -3365
rect 4860 -3405 4870 -3365
rect 4810 -3435 4870 -3405
rect 4810 -3475 4820 -3435
rect 4860 -3475 4870 -3435
rect 4810 -3505 4870 -3475
rect 4810 -3545 4820 -3505
rect 4860 -3545 4870 -3505
rect 4810 -3575 4870 -3545
rect 4810 -3615 4820 -3575
rect 4860 -3615 4870 -3575
rect 4810 -3640 4870 -3615
rect 4810 -3680 4820 -3640
rect 4860 -3680 4870 -3640
rect 4810 -3700 4870 -3680
rect 4810 -3740 4820 -3700
rect 4860 -3740 4870 -3700
rect 4810 -3765 4870 -3740
rect 4810 -3805 4820 -3765
rect 4860 -3805 4870 -3765
rect 4810 -3835 4870 -3805
rect 4810 -3875 4820 -3835
rect 4860 -3875 4870 -3835
rect 4810 -3905 4870 -3875
rect 4810 -3945 4820 -3905
rect 4860 -3945 4870 -3905
rect 4810 -3975 4870 -3945
rect 4810 -4015 4820 -3975
rect 4860 -4015 4870 -3975
rect 4810 -4040 4870 -4015
rect 4810 -4080 4820 -4040
rect 4860 -4080 4870 -4040
rect 4810 -4100 4870 -4080
rect 4810 -4140 4820 -4100
rect 4860 -4140 4870 -4100
rect 4810 -4165 4870 -4140
rect 4810 -4205 4820 -4165
rect 4860 -4205 4870 -4165
rect 4810 -4235 4870 -4205
rect 4810 -4275 4820 -4235
rect 4860 -4275 4870 -4235
rect 4810 -4305 4870 -4275
rect 4810 -4345 4820 -4305
rect 4860 -4345 4870 -4305
rect 4810 -4375 4870 -4345
rect 4810 -4415 4820 -4375
rect 4860 -4415 4870 -4375
rect 4810 -4440 4870 -4415
rect 4810 -4480 4820 -4440
rect 4860 -4480 4870 -4440
rect 4810 -4490 4870 -4480
rect 5160 -1300 5220 -1290
rect 5160 -1340 5170 -1300
rect 5210 -1340 5220 -1300
rect 5160 -1365 5220 -1340
rect 5160 -1405 5170 -1365
rect 5210 -1405 5220 -1365
rect 5160 -1435 5220 -1405
rect 5160 -1475 5170 -1435
rect 5210 -1475 5220 -1435
rect 5160 -1505 5220 -1475
rect 5160 -1545 5170 -1505
rect 5210 -1545 5220 -1505
rect 5160 -1575 5220 -1545
rect 5160 -1615 5170 -1575
rect 5210 -1615 5220 -1575
rect 5160 -1640 5220 -1615
rect 5160 -1680 5170 -1640
rect 5210 -1680 5220 -1640
rect 5160 -1700 5220 -1680
rect 5160 -1740 5170 -1700
rect 5210 -1740 5220 -1700
rect 5160 -1765 5220 -1740
rect 5160 -1805 5170 -1765
rect 5210 -1805 5220 -1765
rect 5160 -1835 5220 -1805
rect 5160 -1875 5170 -1835
rect 5210 -1875 5220 -1835
rect 5160 -1905 5220 -1875
rect 5160 -1945 5170 -1905
rect 5210 -1945 5220 -1905
rect 5160 -1975 5220 -1945
rect 5160 -2015 5170 -1975
rect 5210 -2015 5220 -1975
rect 5160 -2040 5220 -2015
rect 5160 -2080 5170 -2040
rect 5210 -2080 5220 -2040
rect 5160 -2100 5220 -2080
rect 5160 -2140 5170 -2100
rect 5210 -2140 5220 -2100
rect 5160 -2165 5220 -2140
rect 5160 -2205 5170 -2165
rect 5210 -2205 5220 -2165
rect 5160 -2235 5220 -2205
rect 5160 -2275 5170 -2235
rect 5210 -2275 5220 -2235
rect 5160 -2305 5220 -2275
rect 5160 -2345 5170 -2305
rect 5210 -2345 5220 -2305
rect 5160 -2375 5220 -2345
rect 5160 -2415 5170 -2375
rect 5210 -2415 5220 -2375
rect 5160 -2440 5220 -2415
rect 5160 -2480 5170 -2440
rect 5210 -2480 5220 -2440
rect 5160 -2500 5220 -2480
rect 5160 -2540 5170 -2500
rect 5210 -2540 5220 -2500
rect 5160 -2565 5220 -2540
rect 5160 -2605 5170 -2565
rect 5210 -2605 5220 -2565
rect 5160 -2635 5220 -2605
rect 5160 -2675 5170 -2635
rect 5210 -2675 5220 -2635
rect 5160 -2705 5220 -2675
rect 5160 -2745 5170 -2705
rect 5210 -2745 5220 -2705
rect 5160 -2775 5220 -2745
rect 5160 -2815 5170 -2775
rect 5210 -2815 5220 -2775
rect 5160 -2840 5220 -2815
rect 5160 -2880 5170 -2840
rect 5210 -2880 5220 -2840
rect 5160 -2900 5220 -2880
rect 5160 -2940 5170 -2900
rect 5210 -2940 5220 -2900
rect 5160 -2965 5220 -2940
rect 5160 -3005 5170 -2965
rect 5210 -3005 5220 -2965
rect 5160 -3035 5220 -3005
rect 5160 -3075 5170 -3035
rect 5210 -3075 5220 -3035
rect 5160 -3105 5220 -3075
rect 5160 -3145 5170 -3105
rect 5210 -3145 5220 -3105
rect 5160 -3175 5220 -3145
rect 5160 -3215 5170 -3175
rect 5210 -3215 5220 -3175
rect 5160 -3240 5220 -3215
rect 5160 -3280 5170 -3240
rect 5210 -3280 5220 -3240
rect 5160 -3300 5220 -3280
rect 5160 -3340 5170 -3300
rect 5210 -3340 5220 -3300
rect 5160 -3365 5220 -3340
rect 5160 -3405 5170 -3365
rect 5210 -3405 5220 -3365
rect 5160 -3435 5220 -3405
rect 5160 -3475 5170 -3435
rect 5210 -3475 5220 -3435
rect 5160 -3505 5220 -3475
rect 5160 -3545 5170 -3505
rect 5210 -3545 5220 -3505
rect 5160 -3575 5220 -3545
rect 5160 -3615 5170 -3575
rect 5210 -3615 5220 -3575
rect 5160 -3640 5220 -3615
rect 5160 -3680 5170 -3640
rect 5210 -3680 5220 -3640
rect 5160 -3700 5220 -3680
rect 5160 -3740 5170 -3700
rect 5210 -3740 5220 -3700
rect 5160 -3765 5220 -3740
rect 5160 -3805 5170 -3765
rect 5210 -3805 5220 -3765
rect 5160 -3835 5220 -3805
rect 5160 -3875 5170 -3835
rect 5210 -3875 5220 -3835
rect 5160 -3905 5220 -3875
rect 5160 -3945 5170 -3905
rect 5210 -3945 5220 -3905
rect 5160 -3975 5220 -3945
rect 5160 -4015 5170 -3975
rect 5210 -4015 5220 -3975
rect 5160 -4040 5220 -4015
rect 5160 -4080 5170 -4040
rect 5210 -4080 5220 -4040
rect 5160 -4100 5220 -4080
rect 5160 -4140 5170 -4100
rect 5210 -4140 5220 -4100
rect 5160 -4165 5220 -4140
rect 5160 -4205 5170 -4165
rect 5210 -4205 5220 -4165
rect 5160 -4235 5220 -4205
rect 5160 -4275 5170 -4235
rect 5210 -4275 5220 -4235
rect 5160 -4305 5220 -4275
rect 5160 -4345 5170 -4305
rect 5210 -4345 5220 -4305
rect 5160 -4375 5220 -4345
rect 5160 -4415 5170 -4375
rect 5210 -4415 5220 -4375
rect 5160 -4440 5220 -4415
rect 5160 -4480 5170 -4440
rect 5210 -4480 5220 -4440
rect 5160 -4490 5220 -4480
rect 5510 -1300 5570 -1290
rect 5510 -1340 5520 -1300
rect 5560 -1340 5570 -1300
rect 5510 -1365 5570 -1340
rect 5510 -1405 5520 -1365
rect 5560 -1405 5570 -1365
rect 5510 -1435 5570 -1405
rect 5510 -1475 5520 -1435
rect 5560 -1475 5570 -1435
rect 5510 -1505 5570 -1475
rect 5510 -1545 5520 -1505
rect 5560 -1545 5570 -1505
rect 5510 -1575 5570 -1545
rect 5510 -1615 5520 -1575
rect 5560 -1615 5570 -1575
rect 5510 -1640 5570 -1615
rect 5510 -1680 5520 -1640
rect 5560 -1680 5570 -1640
rect 5510 -1700 5570 -1680
rect 5510 -1740 5520 -1700
rect 5560 -1740 5570 -1700
rect 5510 -1765 5570 -1740
rect 5510 -1805 5520 -1765
rect 5560 -1805 5570 -1765
rect 5510 -1835 5570 -1805
rect 5510 -1875 5520 -1835
rect 5560 -1875 5570 -1835
rect 5510 -1905 5570 -1875
rect 5510 -1945 5520 -1905
rect 5560 -1945 5570 -1905
rect 5510 -1975 5570 -1945
rect 5510 -2015 5520 -1975
rect 5560 -2015 5570 -1975
rect 5510 -2040 5570 -2015
rect 5510 -2080 5520 -2040
rect 5560 -2080 5570 -2040
rect 5510 -2100 5570 -2080
rect 5510 -2140 5520 -2100
rect 5560 -2140 5570 -2100
rect 5510 -2165 5570 -2140
rect 5510 -2205 5520 -2165
rect 5560 -2205 5570 -2165
rect 5510 -2235 5570 -2205
rect 5510 -2275 5520 -2235
rect 5560 -2275 5570 -2235
rect 5510 -2305 5570 -2275
rect 5510 -2345 5520 -2305
rect 5560 -2345 5570 -2305
rect 5510 -2375 5570 -2345
rect 5510 -2415 5520 -2375
rect 5560 -2415 5570 -2375
rect 5510 -2440 5570 -2415
rect 5510 -2480 5520 -2440
rect 5560 -2480 5570 -2440
rect 5510 -2500 5570 -2480
rect 5510 -2540 5520 -2500
rect 5560 -2540 5570 -2500
rect 5510 -2565 5570 -2540
rect 5510 -2605 5520 -2565
rect 5560 -2605 5570 -2565
rect 5510 -2635 5570 -2605
rect 5510 -2675 5520 -2635
rect 5560 -2675 5570 -2635
rect 5510 -2705 5570 -2675
rect 5510 -2745 5520 -2705
rect 5560 -2745 5570 -2705
rect 5510 -2775 5570 -2745
rect 5510 -2815 5520 -2775
rect 5560 -2815 5570 -2775
rect 5510 -2840 5570 -2815
rect 5510 -2880 5520 -2840
rect 5560 -2880 5570 -2840
rect 5510 -2900 5570 -2880
rect 5510 -2940 5520 -2900
rect 5560 -2940 5570 -2900
rect 5510 -2965 5570 -2940
rect 5510 -3005 5520 -2965
rect 5560 -3005 5570 -2965
rect 5510 -3035 5570 -3005
rect 5510 -3075 5520 -3035
rect 5560 -3075 5570 -3035
rect 5510 -3105 5570 -3075
rect 5510 -3145 5520 -3105
rect 5560 -3145 5570 -3105
rect 5510 -3175 5570 -3145
rect 5510 -3215 5520 -3175
rect 5560 -3215 5570 -3175
rect 5510 -3240 5570 -3215
rect 5510 -3280 5520 -3240
rect 5560 -3280 5570 -3240
rect 5510 -3300 5570 -3280
rect 5510 -3340 5520 -3300
rect 5560 -3340 5570 -3300
rect 5510 -3365 5570 -3340
rect 5510 -3405 5520 -3365
rect 5560 -3405 5570 -3365
rect 5510 -3435 5570 -3405
rect 5510 -3475 5520 -3435
rect 5560 -3475 5570 -3435
rect 5510 -3505 5570 -3475
rect 5510 -3545 5520 -3505
rect 5560 -3545 5570 -3505
rect 5510 -3575 5570 -3545
rect 5510 -3615 5520 -3575
rect 5560 -3615 5570 -3575
rect 5510 -3640 5570 -3615
rect 5510 -3680 5520 -3640
rect 5560 -3680 5570 -3640
rect 5510 -3700 5570 -3680
rect 5510 -3740 5520 -3700
rect 5560 -3740 5570 -3700
rect 5510 -3765 5570 -3740
rect 5510 -3805 5520 -3765
rect 5560 -3805 5570 -3765
rect 5510 -3835 5570 -3805
rect 5510 -3875 5520 -3835
rect 5560 -3875 5570 -3835
rect 5510 -3905 5570 -3875
rect 5510 -3945 5520 -3905
rect 5560 -3945 5570 -3905
rect 5510 -3975 5570 -3945
rect 5510 -4015 5520 -3975
rect 5560 -4015 5570 -3975
rect 5510 -4040 5570 -4015
rect 5510 -4080 5520 -4040
rect 5560 -4080 5570 -4040
rect 5510 -4100 5570 -4080
rect 5510 -4140 5520 -4100
rect 5560 -4140 5570 -4100
rect 5510 -4165 5570 -4140
rect 5510 -4205 5520 -4165
rect 5560 -4205 5570 -4165
rect 5510 -4235 5570 -4205
rect 5510 -4275 5520 -4235
rect 5560 -4275 5570 -4235
rect 5510 -4305 5570 -4275
rect 5510 -4345 5520 -4305
rect 5560 -4345 5570 -4305
rect 5510 -4375 5570 -4345
rect 5510 -4415 5520 -4375
rect 5560 -4415 5570 -4375
rect 5510 -4440 5570 -4415
rect 5510 -4480 5520 -4440
rect 5560 -4480 5570 -4440
rect 5510 -4490 5570 -4480
rect 5860 -1300 5920 -1290
rect 5860 -1340 5870 -1300
rect 5910 -1340 5920 -1300
rect 5860 -1365 5920 -1340
rect 5860 -1405 5870 -1365
rect 5910 -1405 5920 -1365
rect 5860 -1435 5920 -1405
rect 5860 -1475 5870 -1435
rect 5910 -1475 5920 -1435
rect 5860 -1505 5920 -1475
rect 5860 -1545 5870 -1505
rect 5910 -1545 5920 -1505
rect 5860 -1575 5920 -1545
rect 5860 -1615 5870 -1575
rect 5910 -1615 5920 -1575
rect 5860 -1640 5920 -1615
rect 5860 -1680 5870 -1640
rect 5910 -1680 5920 -1640
rect 5860 -1700 5920 -1680
rect 5860 -1740 5870 -1700
rect 5910 -1740 5920 -1700
rect 5860 -1765 5920 -1740
rect 5860 -1805 5870 -1765
rect 5910 -1805 5920 -1765
rect 5860 -1835 5920 -1805
rect 5860 -1875 5870 -1835
rect 5910 -1875 5920 -1835
rect 5860 -1905 5920 -1875
rect 5860 -1945 5870 -1905
rect 5910 -1945 5920 -1905
rect 5860 -1975 5920 -1945
rect 5860 -2015 5870 -1975
rect 5910 -2015 5920 -1975
rect 5860 -2040 5920 -2015
rect 5860 -2080 5870 -2040
rect 5910 -2080 5920 -2040
rect 5860 -2100 5920 -2080
rect 5860 -2140 5870 -2100
rect 5910 -2140 5920 -2100
rect 5860 -2165 5920 -2140
rect 5860 -2205 5870 -2165
rect 5910 -2205 5920 -2165
rect 5860 -2235 5920 -2205
rect 5860 -2275 5870 -2235
rect 5910 -2275 5920 -2235
rect 5860 -2305 5920 -2275
rect 5860 -2345 5870 -2305
rect 5910 -2345 5920 -2305
rect 5860 -2375 5920 -2345
rect 5860 -2415 5870 -2375
rect 5910 -2415 5920 -2375
rect 5860 -2440 5920 -2415
rect 5860 -2480 5870 -2440
rect 5910 -2480 5920 -2440
rect 5860 -2500 5920 -2480
rect 5860 -2540 5870 -2500
rect 5910 -2540 5920 -2500
rect 5860 -2565 5920 -2540
rect 5860 -2605 5870 -2565
rect 5910 -2605 5920 -2565
rect 5860 -2635 5920 -2605
rect 5860 -2675 5870 -2635
rect 5910 -2675 5920 -2635
rect 5860 -2705 5920 -2675
rect 5860 -2745 5870 -2705
rect 5910 -2745 5920 -2705
rect 5860 -2775 5920 -2745
rect 5860 -2815 5870 -2775
rect 5910 -2815 5920 -2775
rect 5860 -2840 5920 -2815
rect 5860 -2880 5870 -2840
rect 5910 -2880 5920 -2840
rect 5860 -2900 5920 -2880
rect 5860 -2940 5870 -2900
rect 5910 -2940 5920 -2900
rect 5860 -2965 5920 -2940
rect 5860 -3005 5870 -2965
rect 5910 -3005 5920 -2965
rect 5860 -3035 5920 -3005
rect 5860 -3075 5870 -3035
rect 5910 -3075 5920 -3035
rect 5860 -3105 5920 -3075
rect 5860 -3145 5870 -3105
rect 5910 -3145 5920 -3105
rect 5860 -3175 5920 -3145
rect 5860 -3215 5870 -3175
rect 5910 -3215 5920 -3175
rect 5860 -3240 5920 -3215
rect 5860 -3280 5870 -3240
rect 5910 -3280 5920 -3240
rect 5860 -3300 5920 -3280
rect 5860 -3340 5870 -3300
rect 5910 -3340 5920 -3300
rect 5860 -3365 5920 -3340
rect 5860 -3405 5870 -3365
rect 5910 -3405 5920 -3365
rect 5860 -3435 5920 -3405
rect 5860 -3475 5870 -3435
rect 5910 -3475 5920 -3435
rect 5860 -3505 5920 -3475
rect 5860 -3545 5870 -3505
rect 5910 -3545 5920 -3505
rect 5860 -3575 5920 -3545
rect 5860 -3615 5870 -3575
rect 5910 -3615 5920 -3575
rect 5860 -3640 5920 -3615
rect 5860 -3680 5870 -3640
rect 5910 -3680 5920 -3640
rect 5860 -3700 5920 -3680
rect 5860 -3740 5870 -3700
rect 5910 -3740 5920 -3700
rect 5860 -3765 5920 -3740
rect 5860 -3805 5870 -3765
rect 5910 -3805 5920 -3765
rect 5860 -3835 5920 -3805
rect 5860 -3875 5870 -3835
rect 5910 -3875 5920 -3835
rect 5860 -3905 5920 -3875
rect 5860 -3945 5870 -3905
rect 5910 -3945 5920 -3905
rect 5860 -3975 5920 -3945
rect 5860 -4015 5870 -3975
rect 5910 -4015 5920 -3975
rect 5860 -4040 5920 -4015
rect 5860 -4080 5870 -4040
rect 5910 -4080 5920 -4040
rect 5860 -4100 5920 -4080
rect 5860 -4140 5870 -4100
rect 5910 -4140 5920 -4100
rect 5860 -4165 5920 -4140
rect 5860 -4205 5870 -4165
rect 5910 -4205 5920 -4165
rect 5860 -4235 5920 -4205
rect 5860 -4275 5870 -4235
rect 5910 -4275 5920 -4235
rect 5860 -4305 5920 -4275
rect 5860 -4345 5870 -4305
rect 5910 -4345 5920 -4305
rect 5860 -4375 5920 -4345
rect 5860 -4415 5870 -4375
rect 5910 -4415 5920 -4375
rect 5860 -4440 5920 -4415
rect 5860 -4480 5870 -4440
rect 5910 -4480 5920 -4440
rect 5860 -4490 5920 -4480
rect 6210 -1300 6270 -1290
rect 6210 -1340 6220 -1300
rect 6260 -1340 6270 -1300
rect 6210 -1365 6270 -1340
rect 6210 -1405 6220 -1365
rect 6260 -1405 6270 -1365
rect 6210 -1435 6270 -1405
rect 6210 -1475 6220 -1435
rect 6260 -1475 6270 -1435
rect 6210 -1505 6270 -1475
rect 6210 -1545 6220 -1505
rect 6260 -1545 6270 -1505
rect 6210 -1575 6270 -1545
rect 6210 -1615 6220 -1575
rect 6260 -1615 6270 -1575
rect 6210 -1640 6270 -1615
rect 6210 -1680 6220 -1640
rect 6260 -1680 6270 -1640
rect 6210 -1700 6270 -1680
rect 6210 -1740 6220 -1700
rect 6260 -1740 6270 -1700
rect 6210 -1765 6270 -1740
rect 6210 -1805 6220 -1765
rect 6260 -1805 6270 -1765
rect 6210 -1835 6270 -1805
rect 6210 -1875 6220 -1835
rect 6260 -1875 6270 -1835
rect 6210 -1905 6270 -1875
rect 6210 -1945 6220 -1905
rect 6260 -1945 6270 -1905
rect 6210 -1975 6270 -1945
rect 6210 -2015 6220 -1975
rect 6260 -2015 6270 -1975
rect 6210 -2040 6270 -2015
rect 6210 -2080 6220 -2040
rect 6260 -2080 6270 -2040
rect 6210 -2100 6270 -2080
rect 6210 -2140 6220 -2100
rect 6260 -2140 6270 -2100
rect 6210 -2165 6270 -2140
rect 6210 -2205 6220 -2165
rect 6260 -2205 6270 -2165
rect 6210 -2235 6270 -2205
rect 6210 -2275 6220 -2235
rect 6260 -2275 6270 -2235
rect 6210 -2305 6270 -2275
rect 6210 -2345 6220 -2305
rect 6260 -2345 6270 -2305
rect 6210 -2375 6270 -2345
rect 6210 -2415 6220 -2375
rect 6260 -2415 6270 -2375
rect 6210 -2440 6270 -2415
rect 6210 -2480 6220 -2440
rect 6260 -2480 6270 -2440
rect 6210 -2500 6270 -2480
rect 6210 -2540 6220 -2500
rect 6260 -2540 6270 -2500
rect 6210 -2565 6270 -2540
rect 6210 -2605 6220 -2565
rect 6260 -2605 6270 -2565
rect 6210 -2635 6270 -2605
rect 6210 -2675 6220 -2635
rect 6260 -2675 6270 -2635
rect 6210 -2705 6270 -2675
rect 6210 -2745 6220 -2705
rect 6260 -2745 6270 -2705
rect 6210 -2775 6270 -2745
rect 6210 -2815 6220 -2775
rect 6260 -2815 6270 -2775
rect 6210 -2840 6270 -2815
rect 6210 -2880 6220 -2840
rect 6260 -2880 6270 -2840
rect 6210 -2900 6270 -2880
rect 6210 -2940 6220 -2900
rect 6260 -2940 6270 -2900
rect 6210 -2965 6270 -2940
rect 6210 -3005 6220 -2965
rect 6260 -3005 6270 -2965
rect 6210 -3035 6270 -3005
rect 6210 -3075 6220 -3035
rect 6260 -3075 6270 -3035
rect 6210 -3105 6270 -3075
rect 6210 -3145 6220 -3105
rect 6260 -3145 6270 -3105
rect 6210 -3175 6270 -3145
rect 6210 -3215 6220 -3175
rect 6260 -3215 6270 -3175
rect 6210 -3240 6270 -3215
rect 6210 -3280 6220 -3240
rect 6260 -3280 6270 -3240
rect 6210 -3300 6270 -3280
rect 6210 -3340 6220 -3300
rect 6260 -3340 6270 -3300
rect 6210 -3365 6270 -3340
rect 6210 -3405 6220 -3365
rect 6260 -3405 6270 -3365
rect 6210 -3435 6270 -3405
rect 6210 -3475 6220 -3435
rect 6260 -3475 6270 -3435
rect 6210 -3505 6270 -3475
rect 6210 -3545 6220 -3505
rect 6260 -3545 6270 -3505
rect 6210 -3575 6270 -3545
rect 6210 -3615 6220 -3575
rect 6260 -3615 6270 -3575
rect 6210 -3640 6270 -3615
rect 6210 -3680 6220 -3640
rect 6260 -3680 6270 -3640
rect 6210 -3700 6270 -3680
rect 6210 -3740 6220 -3700
rect 6260 -3740 6270 -3700
rect 6210 -3765 6270 -3740
rect 6210 -3805 6220 -3765
rect 6260 -3805 6270 -3765
rect 6210 -3835 6270 -3805
rect 6210 -3875 6220 -3835
rect 6260 -3875 6270 -3835
rect 6210 -3905 6270 -3875
rect 6210 -3945 6220 -3905
rect 6260 -3945 6270 -3905
rect 6210 -3975 6270 -3945
rect 6210 -4015 6220 -3975
rect 6260 -4015 6270 -3975
rect 6210 -4040 6270 -4015
rect 6210 -4080 6220 -4040
rect 6260 -4080 6270 -4040
rect 6210 -4100 6270 -4080
rect 6210 -4140 6220 -4100
rect 6260 -4140 6270 -4100
rect 6210 -4165 6270 -4140
rect 6210 -4205 6220 -4165
rect 6260 -4205 6270 -4165
rect 6210 -4235 6270 -4205
rect 6210 -4275 6220 -4235
rect 6260 -4275 6270 -4235
rect 6210 -4305 6270 -4275
rect 6210 -4345 6220 -4305
rect 6260 -4345 6270 -4305
rect 6210 -4375 6270 -4345
rect 6210 -4415 6220 -4375
rect 6260 -4415 6270 -4375
rect 6210 -4440 6270 -4415
rect 6210 -4480 6220 -4440
rect 6260 -4480 6270 -4440
rect 6210 -4490 6270 -4480
rect 6560 -1300 6620 -1290
rect 6560 -1340 6570 -1300
rect 6610 -1340 6620 -1300
rect 6560 -1365 6620 -1340
rect 6560 -1405 6570 -1365
rect 6610 -1405 6620 -1365
rect 6560 -1435 6620 -1405
rect 6560 -1475 6570 -1435
rect 6610 -1475 6620 -1435
rect 6560 -1505 6620 -1475
rect 6560 -1545 6570 -1505
rect 6610 -1545 6620 -1505
rect 6560 -1575 6620 -1545
rect 6560 -1615 6570 -1575
rect 6610 -1615 6620 -1575
rect 6560 -1640 6620 -1615
rect 6560 -1680 6570 -1640
rect 6610 -1680 6620 -1640
rect 6560 -1700 6620 -1680
rect 6560 -1740 6570 -1700
rect 6610 -1740 6620 -1700
rect 6560 -1765 6620 -1740
rect 6560 -1805 6570 -1765
rect 6610 -1805 6620 -1765
rect 6560 -1835 6620 -1805
rect 6560 -1875 6570 -1835
rect 6610 -1875 6620 -1835
rect 6560 -1905 6620 -1875
rect 6560 -1945 6570 -1905
rect 6610 -1945 6620 -1905
rect 6560 -1975 6620 -1945
rect 6560 -2015 6570 -1975
rect 6610 -2015 6620 -1975
rect 6560 -2040 6620 -2015
rect 6560 -2080 6570 -2040
rect 6610 -2080 6620 -2040
rect 6560 -2100 6620 -2080
rect 6560 -2140 6570 -2100
rect 6610 -2140 6620 -2100
rect 6560 -2165 6620 -2140
rect 6560 -2205 6570 -2165
rect 6610 -2205 6620 -2165
rect 6560 -2235 6620 -2205
rect 6560 -2275 6570 -2235
rect 6610 -2275 6620 -2235
rect 6560 -2305 6620 -2275
rect 6560 -2345 6570 -2305
rect 6610 -2345 6620 -2305
rect 6560 -2375 6620 -2345
rect 6560 -2415 6570 -2375
rect 6610 -2415 6620 -2375
rect 6560 -2440 6620 -2415
rect 6560 -2480 6570 -2440
rect 6610 -2480 6620 -2440
rect 6560 -2500 6620 -2480
rect 6560 -2540 6570 -2500
rect 6610 -2540 6620 -2500
rect 6560 -2565 6620 -2540
rect 6560 -2605 6570 -2565
rect 6610 -2605 6620 -2565
rect 6560 -2635 6620 -2605
rect 6560 -2675 6570 -2635
rect 6610 -2675 6620 -2635
rect 6560 -2705 6620 -2675
rect 6560 -2745 6570 -2705
rect 6610 -2745 6620 -2705
rect 6560 -2775 6620 -2745
rect 6560 -2815 6570 -2775
rect 6610 -2815 6620 -2775
rect 6560 -2840 6620 -2815
rect 6560 -2880 6570 -2840
rect 6610 -2880 6620 -2840
rect 6560 -2900 6620 -2880
rect 6560 -2940 6570 -2900
rect 6610 -2940 6620 -2900
rect 6560 -2965 6620 -2940
rect 6560 -3005 6570 -2965
rect 6610 -3005 6620 -2965
rect 6560 -3035 6620 -3005
rect 6560 -3075 6570 -3035
rect 6610 -3075 6620 -3035
rect 6560 -3105 6620 -3075
rect 6560 -3145 6570 -3105
rect 6610 -3145 6620 -3105
rect 6560 -3175 6620 -3145
rect 6560 -3215 6570 -3175
rect 6610 -3215 6620 -3175
rect 6560 -3240 6620 -3215
rect 6560 -3280 6570 -3240
rect 6610 -3280 6620 -3240
rect 6560 -3300 6620 -3280
rect 6560 -3340 6570 -3300
rect 6610 -3340 6620 -3300
rect 6560 -3365 6620 -3340
rect 6560 -3405 6570 -3365
rect 6610 -3405 6620 -3365
rect 6560 -3435 6620 -3405
rect 6560 -3475 6570 -3435
rect 6610 -3475 6620 -3435
rect 6560 -3505 6620 -3475
rect 6560 -3545 6570 -3505
rect 6610 -3545 6620 -3505
rect 6560 -3575 6620 -3545
rect 6560 -3615 6570 -3575
rect 6610 -3615 6620 -3575
rect 6560 -3640 6620 -3615
rect 6560 -3680 6570 -3640
rect 6610 -3680 6620 -3640
rect 6560 -3700 6620 -3680
rect 6560 -3740 6570 -3700
rect 6610 -3740 6620 -3700
rect 6560 -3765 6620 -3740
rect 6560 -3805 6570 -3765
rect 6610 -3805 6620 -3765
rect 6560 -3835 6620 -3805
rect 6560 -3875 6570 -3835
rect 6610 -3875 6620 -3835
rect 6560 -3905 6620 -3875
rect 6560 -3945 6570 -3905
rect 6610 -3945 6620 -3905
rect 6560 -3975 6620 -3945
rect 6560 -4015 6570 -3975
rect 6610 -4015 6620 -3975
rect 6560 -4040 6620 -4015
rect 6560 -4080 6570 -4040
rect 6610 -4080 6620 -4040
rect 6560 -4100 6620 -4080
rect 6560 -4140 6570 -4100
rect 6610 -4140 6620 -4100
rect 6560 -4165 6620 -4140
rect 6560 -4205 6570 -4165
rect 6610 -4205 6620 -4165
rect 6560 -4235 6620 -4205
rect 6560 -4275 6570 -4235
rect 6610 -4275 6620 -4235
rect 6560 -4305 6620 -4275
rect 6560 -4345 6570 -4305
rect 6610 -4345 6620 -4305
rect 6560 -4375 6620 -4345
rect 6560 -4415 6570 -4375
rect 6610 -4415 6620 -4375
rect 6560 -4440 6620 -4415
rect 6560 -4480 6570 -4440
rect 6610 -4480 6620 -4440
rect 6560 -4490 6620 -4480
rect 6910 -1300 6970 -1290
rect 6910 -1340 6920 -1300
rect 6960 -1340 6970 -1300
rect 6910 -1365 6970 -1340
rect 6910 -1405 6920 -1365
rect 6960 -1405 6970 -1365
rect 6910 -1435 6970 -1405
rect 6910 -1475 6920 -1435
rect 6960 -1475 6970 -1435
rect 6910 -1505 6970 -1475
rect 6910 -1545 6920 -1505
rect 6960 -1545 6970 -1505
rect 6910 -1575 6970 -1545
rect 6910 -1615 6920 -1575
rect 6960 -1615 6970 -1575
rect 6910 -1640 6970 -1615
rect 6910 -1680 6920 -1640
rect 6960 -1680 6970 -1640
rect 6910 -1700 6970 -1680
rect 6910 -1740 6920 -1700
rect 6960 -1740 6970 -1700
rect 6910 -1765 6970 -1740
rect 6910 -1805 6920 -1765
rect 6960 -1805 6970 -1765
rect 6910 -1835 6970 -1805
rect 6910 -1875 6920 -1835
rect 6960 -1875 6970 -1835
rect 6910 -1905 6970 -1875
rect 6910 -1945 6920 -1905
rect 6960 -1945 6970 -1905
rect 6910 -1975 6970 -1945
rect 6910 -2015 6920 -1975
rect 6960 -2015 6970 -1975
rect 6910 -2040 6970 -2015
rect 6910 -2080 6920 -2040
rect 6960 -2080 6970 -2040
rect 6910 -2100 6970 -2080
rect 6910 -2140 6920 -2100
rect 6960 -2140 6970 -2100
rect 6910 -2165 6970 -2140
rect 6910 -2205 6920 -2165
rect 6960 -2205 6970 -2165
rect 6910 -2235 6970 -2205
rect 6910 -2275 6920 -2235
rect 6960 -2275 6970 -2235
rect 6910 -2305 6970 -2275
rect 6910 -2345 6920 -2305
rect 6960 -2345 6970 -2305
rect 6910 -2375 6970 -2345
rect 6910 -2415 6920 -2375
rect 6960 -2415 6970 -2375
rect 6910 -2440 6970 -2415
rect 6910 -2480 6920 -2440
rect 6960 -2480 6970 -2440
rect 6910 -2500 6970 -2480
rect 6910 -2540 6920 -2500
rect 6960 -2540 6970 -2500
rect 6910 -2565 6970 -2540
rect 6910 -2605 6920 -2565
rect 6960 -2605 6970 -2565
rect 6910 -2635 6970 -2605
rect 6910 -2675 6920 -2635
rect 6960 -2675 6970 -2635
rect 6910 -2705 6970 -2675
rect 6910 -2745 6920 -2705
rect 6960 -2745 6970 -2705
rect 6910 -2775 6970 -2745
rect 6910 -2815 6920 -2775
rect 6960 -2815 6970 -2775
rect 6910 -2840 6970 -2815
rect 6910 -2880 6920 -2840
rect 6960 -2880 6970 -2840
rect 6910 -2900 6970 -2880
rect 6910 -2940 6920 -2900
rect 6960 -2940 6970 -2900
rect 6910 -2965 6970 -2940
rect 6910 -3005 6920 -2965
rect 6960 -3005 6970 -2965
rect 6910 -3035 6970 -3005
rect 6910 -3075 6920 -3035
rect 6960 -3075 6970 -3035
rect 6910 -3105 6970 -3075
rect 6910 -3145 6920 -3105
rect 6960 -3145 6970 -3105
rect 6910 -3175 6970 -3145
rect 6910 -3215 6920 -3175
rect 6960 -3215 6970 -3175
rect 6910 -3240 6970 -3215
rect 6910 -3280 6920 -3240
rect 6960 -3280 6970 -3240
rect 6910 -3300 6970 -3280
rect 6910 -3340 6920 -3300
rect 6960 -3340 6970 -3300
rect 6910 -3365 6970 -3340
rect 6910 -3405 6920 -3365
rect 6960 -3405 6970 -3365
rect 6910 -3435 6970 -3405
rect 6910 -3475 6920 -3435
rect 6960 -3475 6970 -3435
rect 6910 -3505 6970 -3475
rect 6910 -3545 6920 -3505
rect 6960 -3545 6970 -3505
rect 6910 -3575 6970 -3545
rect 6910 -3615 6920 -3575
rect 6960 -3615 6970 -3575
rect 6910 -3640 6970 -3615
rect 6910 -3680 6920 -3640
rect 6960 -3680 6970 -3640
rect 6910 -3700 6970 -3680
rect 6910 -3740 6920 -3700
rect 6960 -3740 6970 -3700
rect 6910 -3765 6970 -3740
rect 6910 -3805 6920 -3765
rect 6960 -3805 6970 -3765
rect 6910 -3835 6970 -3805
rect 6910 -3875 6920 -3835
rect 6960 -3875 6970 -3835
rect 6910 -3905 6970 -3875
rect 6910 -3945 6920 -3905
rect 6960 -3945 6970 -3905
rect 6910 -3975 6970 -3945
rect 6910 -4015 6920 -3975
rect 6960 -4015 6970 -3975
rect 6910 -4040 6970 -4015
rect 6910 -4080 6920 -4040
rect 6960 -4080 6970 -4040
rect 6910 -4100 6970 -4080
rect 6910 -4140 6920 -4100
rect 6960 -4140 6970 -4100
rect 6910 -4165 6970 -4140
rect 6910 -4205 6920 -4165
rect 6960 -4205 6970 -4165
rect 6910 -4235 6970 -4205
rect 6910 -4275 6920 -4235
rect 6960 -4275 6970 -4235
rect 6910 -4305 6970 -4275
rect 6910 -4345 6920 -4305
rect 6960 -4345 6970 -4305
rect 6910 -4375 6970 -4345
rect 6910 -4415 6920 -4375
rect 6960 -4415 6970 -4375
rect 6910 -4440 6970 -4415
rect 6910 -4480 6920 -4440
rect 6960 -4480 6970 -4440
rect 6910 -4490 6970 -4480
rect 7260 -1300 7320 -1290
rect 7260 -1340 7270 -1300
rect 7310 -1340 7320 -1300
rect 7260 -1365 7320 -1340
rect 7260 -1405 7270 -1365
rect 7310 -1405 7320 -1365
rect 7260 -1435 7320 -1405
rect 7260 -1475 7270 -1435
rect 7310 -1475 7320 -1435
rect 7260 -1505 7320 -1475
rect 7260 -1545 7270 -1505
rect 7310 -1545 7320 -1505
rect 7260 -1575 7320 -1545
rect 7260 -1615 7270 -1575
rect 7310 -1615 7320 -1575
rect 7260 -1640 7320 -1615
rect 7260 -1680 7270 -1640
rect 7310 -1680 7320 -1640
rect 7260 -1700 7320 -1680
rect 7260 -1740 7270 -1700
rect 7310 -1740 7320 -1700
rect 7260 -1765 7320 -1740
rect 7260 -1805 7270 -1765
rect 7310 -1805 7320 -1765
rect 7260 -1835 7320 -1805
rect 7260 -1875 7270 -1835
rect 7310 -1875 7320 -1835
rect 7260 -1905 7320 -1875
rect 7260 -1945 7270 -1905
rect 7310 -1945 7320 -1905
rect 7260 -1975 7320 -1945
rect 7260 -2015 7270 -1975
rect 7310 -2015 7320 -1975
rect 7260 -2040 7320 -2015
rect 7260 -2080 7270 -2040
rect 7310 -2080 7320 -2040
rect 7260 -2100 7320 -2080
rect 7260 -2140 7270 -2100
rect 7310 -2140 7320 -2100
rect 7260 -2165 7320 -2140
rect 7260 -2205 7270 -2165
rect 7310 -2205 7320 -2165
rect 7260 -2235 7320 -2205
rect 7260 -2275 7270 -2235
rect 7310 -2275 7320 -2235
rect 7260 -2305 7320 -2275
rect 7260 -2345 7270 -2305
rect 7310 -2345 7320 -2305
rect 7260 -2375 7320 -2345
rect 7260 -2415 7270 -2375
rect 7310 -2415 7320 -2375
rect 7260 -2440 7320 -2415
rect 7260 -2480 7270 -2440
rect 7310 -2480 7320 -2440
rect 7260 -2500 7320 -2480
rect 7260 -2540 7270 -2500
rect 7310 -2540 7320 -2500
rect 7260 -2565 7320 -2540
rect 7260 -2605 7270 -2565
rect 7310 -2605 7320 -2565
rect 7260 -2635 7320 -2605
rect 7260 -2675 7270 -2635
rect 7310 -2675 7320 -2635
rect 7260 -2705 7320 -2675
rect 7260 -2745 7270 -2705
rect 7310 -2745 7320 -2705
rect 7260 -2775 7320 -2745
rect 7260 -2815 7270 -2775
rect 7310 -2815 7320 -2775
rect 7260 -2840 7320 -2815
rect 7260 -2880 7270 -2840
rect 7310 -2880 7320 -2840
rect 7260 -2900 7320 -2880
rect 7260 -2940 7270 -2900
rect 7310 -2940 7320 -2900
rect 7260 -2965 7320 -2940
rect 7260 -3005 7270 -2965
rect 7310 -3005 7320 -2965
rect 7260 -3035 7320 -3005
rect 7260 -3075 7270 -3035
rect 7310 -3075 7320 -3035
rect 7260 -3105 7320 -3075
rect 7260 -3145 7270 -3105
rect 7310 -3145 7320 -3105
rect 7260 -3175 7320 -3145
rect 7260 -3215 7270 -3175
rect 7310 -3215 7320 -3175
rect 7260 -3240 7320 -3215
rect 7260 -3280 7270 -3240
rect 7310 -3280 7320 -3240
rect 7260 -3300 7320 -3280
rect 7260 -3340 7270 -3300
rect 7310 -3340 7320 -3300
rect 7260 -3365 7320 -3340
rect 7260 -3405 7270 -3365
rect 7310 -3405 7320 -3365
rect 7260 -3435 7320 -3405
rect 7260 -3475 7270 -3435
rect 7310 -3475 7320 -3435
rect 7260 -3505 7320 -3475
rect 7260 -3545 7270 -3505
rect 7310 -3545 7320 -3505
rect 7260 -3575 7320 -3545
rect 7260 -3615 7270 -3575
rect 7310 -3615 7320 -3575
rect 7260 -3640 7320 -3615
rect 7260 -3680 7270 -3640
rect 7310 -3680 7320 -3640
rect 7260 -3700 7320 -3680
rect 7260 -3740 7270 -3700
rect 7310 -3740 7320 -3700
rect 7260 -3765 7320 -3740
rect 7260 -3805 7270 -3765
rect 7310 -3805 7320 -3765
rect 7260 -3835 7320 -3805
rect 7260 -3875 7270 -3835
rect 7310 -3875 7320 -3835
rect 7260 -3905 7320 -3875
rect 7260 -3945 7270 -3905
rect 7310 -3945 7320 -3905
rect 7260 -3975 7320 -3945
rect 7260 -4015 7270 -3975
rect 7310 -4015 7320 -3975
rect 7260 -4040 7320 -4015
rect 7260 -4080 7270 -4040
rect 7310 -4080 7320 -4040
rect 7260 -4100 7320 -4080
rect 7260 -4140 7270 -4100
rect 7310 -4140 7320 -4100
rect 7260 -4165 7320 -4140
rect 7260 -4205 7270 -4165
rect 7310 -4205 7320 -4165
rect 7260 -4235 7320 -4205
rect 7260 -4275 7270 -4235
rect 7310 -4275 7320 -4235
rect 7260 -4305 7320 -4275
rect 7260 -4345 7270 -4305
rect 7310 -4345 7320 -4305
rect 7260 -4375 7320 -4345
rect 7260 -4415 7270 -4375
rect 7310 -4415 7320 -4375
rect 7260 -4440 7320 -4415
rect 7260 -4480 7270 -4440
rect 7310 -4480 7320 -4440
rect 7260 -4490 7320 -4480
rect 7610 -1300 7670 -1290
rect 7610 -1340 7620 -1300
rect 7660 -1340 7670 -1300
rect 7610 -1365 7670 -1340
rect 7610 -1405 7620 -1365
rect 7660 -1405 7670 -1365
rect 7610 -1435 7670 -1405
rect 7610 -1475 7620 -1435
rect 7660 -1475 7670 -1435
rect 7610 -1505 7670 -1475
rect 7610 -1545 7620 -1505
rect 7660 -1545 7670 -1505
rect 7610 -1575 7670 -1545
rect 7610 -1615 7620 -1575
rect 7660 -1615 7670 -1575
rect 7610 -1640 7670 -1615
rect 7610 -1680 7620 -1640
rect 7660 -1680 7670 -1640
rect 7610 -1700 7670 -1680
rect 7610 -1740 7620 -1700
rect 7660 -1740 7670 -1700
rect 7610 -1765 7670 -1740
rect 7610 -1805 7620 -1765
rect 7660 -1805 7670 -1765
rect 7610 -1835 7670 -1805
rect 7610 -1875 7620 -1835
rect 7660 -1875 7670 -1835
rect 7610 -1905 7670 -1875
rect 7610 -1945 7620 -1905
rect 7660 -1945 7670 -1905
rect 7610 -1975 7670 -1945
rect 7610 -2015 7620 -1975
rect 7660 -2015 7670 -1975
rect 7610 -2040 7670 -2015
rect 7610 -2080 7620 -2040
rect 7660 -2080 7670 -2040
rect 7610 -2100 7670 -2080
rect 7610 -2140 7620 -2100
rect 7660 -2140 7670 -2100
rect 7610 -2165 7670 -2140
rect 7610 -2205 7620 -2165
rect 7660 -2205 7670 -2165
rect 7610 -2235 7670 -2205
rect 7610 -2275 7620 -2235
rect 7660 -2275 7670 -2235
rect 7610 -2305 7670 -2275
rect 7610 -2345 7620 -2305
rect 7660 -2345 7670 -2305
rect 7610 -2375 7670 -2345
rect 7610 -2415 7620 -2375
rect 7660 -2415 7670 -2375
rect 7610 -2440 7670 -2415
rect 7610 -2480 7620 -2440
rect 7660 -2480 7670 -2440
rect 7610 -2500 7670 -2480
rect 7610 -2540 7620 -2500
rect 7660 -2540 7670 -2500
rect 7610 -2565 7670 -2540
rect 7610 -2605 7620 -2565
rect 7660 -2605 7670 -2565
rect 7610 -2635 7670 -2605
rect 7610 -2675 7620 -2635
rect 7660 -2675 7670 -2635
rect 7610 -2705 7670 -2675
rect 7610 -2745 7620 -2705
rect 7660 -2745 7670 -2705
rect 7610 -2775 7670 -2745
rect 7610 -2815 7620 -2775
rect 7660 -2815 7670 -2775
rect 7610 -2840 7670 -2815
rect 7610 -2880 7620 -2840
rect 7660 -2880 7670 -2840
rect 7610 -2900 7670 -2880
rect 7610 -2940 7620 -2900
rect 7660 -2940 7670 -2900
rect 7610 -2965 7670 -2940
rect 7610 -3005 7620 -2965
rect 7660 -3005 7670 -2965
rect 7610 -3035 7670 -3005
rect 7610 -3075 7620 -3035
rect 7660 -3075 7670 -3035
rect 7610 -3105 7670 -3075
rect 7610 -3145 7620 -3105
rect 7660 -3145 7670 -3105
rect 7610 -3175 7670 -3145
rect 7610 -3215 7620 -3175
rect 7660 -3215 7670 -3175
rect 7610 -3240 7670 -3215
rect 7610 -3280 7620 -3240
rect 7660 -3280 7670 -3240
rect 7610 -3300 7670 -3280
rect 7610 -3340 7620 -3300
rect 7660 -3340 7670 -3300
rect 7610 -3365 7670 -3340
rect 7610 -3405 7620 -3365
rect 7660 -3405 7670 -3365
rect 7610 -3435 7670 -3405
rect 7610 -3475 7620 -3435
rect 7660 -3475 7670 -3435
rect 7610 -3505 7670 -3475
rect 7610 -3545 7620 -3505
rect 7660 -3545 7670 -3505
rect 7610 -3575 7670 -3545
rect 7610 -3615 7620 -3575
rect 7660 -3615 7670 -3575
rect 7610 -3640 7670 -3615
rect 7610 -3680 7620 -3640
rect 7660 -3680 7670 -3640
rect 7610 -3700 7670 -3680
rect 7610 -3740 7620 -3700
rect 7660 -3740 7670 -3700
rect 7610 -3765 7670 -3740
rect 7610 -3805 7620 -3765
rect 7660 -3805 7670 -3765
rect 7610 -3835 7670 -3805
rect 7610 -3875 7620 -3835
rect 7660 -3875 7670 -3835
rect 7610 -3905 7670 -3875
rect 7610 -3945 7620 -3905
rect 7660 -3945 7670 -3905
rect 7610 -3975 7670 -3945
rect 7610 -4015 7620 -3975
rect 7660 -4015 7670 -3975
rect 7610 -4040 7670 -4015
rect 7610 -4080 7620 -4040
rect 7660 -4080 7670 -4040
rect 7610 -4100 7670 -4080
rect 7610 -4140 7620 -4100
rect 7660 -4140 7670 -4100
rect 7610 -4165 7670 -4140
rect 7610 -4205 7620 -4165
rect 7660 -4205 7670 -4165
rect 7610 -4235 7670 -4205
rect 7610 -4275 7620 -4235
rect 7660 -4275 7670 -4235
rect 7610 -4305 7670 -4275
rect 7610 -4345 7620 -4305
rect 7660 -4345 7670 -4305
rect 7610 -4375 7670 -4345
rect 7610 -4415 7620 -4375
rect 7660 -4415 7670 -4375
rect 7610 -4440 7670 -4415
rect 7610 -4480 7620 -4440
rect 7660 -4480 7670 -4440
rect 7610 -4490 7670 -4480
rect 7960 -1300 8020 -1290
rect 7960 -1340 7970 -1300
rect 8010 -1340 8020 -1300
rect 7960 -1365 8020 -1340
rect 7960 -1405 7970 -1365
rect 8010 -1405 8020 -1365
rect 7960 -1435 8020 -1405
rect 7960 -1475 7970 -1435
rect 8010 -1475 8020 -1435
rect 7960 -1505 8020 -1475
rect 7960 -1545 7970 -1505
rect 8010 -1545 8020 -1505
rect 7960 -1575 8020 -1545
rect 7960 -1615 7970 -1575
rect 8010 -1615 8020 -1575
rect 7960 -1640 8020 -1615
rect 7960 -1680 7970 -1640
rect 8010 -1680 8020 -1640
rect 7960 -1700 8020 -1680
rect 7960 -1740 7970 -1700
rect 8010 -1740 8020 -1700
rect 7960 -1765 8020 -1740
rect 7960 -1805 7970 -1765
rect 8010 -1805 8020 -1765
rect 7960 -1835 8020 -1805
rect 7960 -1875 7970 -1835
rect 8010 -1875 8020 -1835
rect 7960 -1905 8020 -1875
rect 7960 -1945 7970 -1905
rect 8010 -1945 8020 -1905
rect 7960 -1975 8020 -1945
rect 7960 -2015 7970 -1975
rect 8010 -2015 8020 -1975
rect 7960 -2040 8020 -2015
rect 7960 -2080 7970 -2040
rect 8010 -2080 8020 -2040
rect 7960 -2100 8020 -2080
rect 7960 -2140 7970 -2100
rect 8010 -2140 8020 -2100
rect 7960 -2165 8020 -2140
rect 7960 -2205 7970 -2165
rect 8010 -2205 8020 -2165
rect 7960 -2235 8020 -2205
rect 7960 -2275 7970 -2235
rect 8010 -2275 8020 -2235
rect 7960 -2305 8020 -2275
rect 7960 -2345 7970 -2305
rect 8010 -2345 8020 -2305
rect 7960 -2375 8020 -2345
rect 7960 -2415 7970 -2375
rect 8010 -2415 8020 -2375
rect 7960 -2440 8020 -2415
rect 7960 -2480 7970 -2440
rect 8010 -2480 8020 -2440
rect 7960 -2500 8020 -2480
rect 7960 -2540 7970 -2500
rect 8010 -2540 8020 -2500
rect 7960 -2565 8020 -2540
rect 7960 -2605 7970 -2565
rect 8010 -2605 8020 -2565
rect 7960 -2635 8020 -2605
rect 7960 -2675 7970 -2635
rect 8010 -2675 8020 -2635
rect 7960 -2705 8020 -2675
rect 7960 -2745 7970 -2705
rect 8010 -2745 8020 -2705
rect 7960 -2775 8020 -2745
rect 7960 -2815 7970 -2775
rect 8010 -2815 8020 -2775
rect 7960 -2840 8020 -2815
rect 7960 -2880 7970 -2840
rect 8010 -2880 8020 -2840
rect 7960 -2900 8020 -2880
rect 7960 -2940 7970 -2900
rect 8010 -2940 8020 -2900
rect 7960 -2965 8020 -2940
rect 7960 -3005 7970 -2965
rect 8010 -3005 8020 -2965
rect 7960 -3035 8020 -3005
rect 7960 -3075 7970 -3035
rect 8010 -3075 8020 -3035
rect 7960 -3105 8020 -3075
rect 7960 -3145 7970 -3105
rect 8010 -3145 8020 -3105
rect 7960 -3175 8020 -3145
rect 7960 -3215 7970 -3175
rect 8010 -3215 8020 -3175
rect 7960 -3240 8020 -3215
rect 7960 -3280 7970 -3240
rect 8010 -3280 8020 -3240
rect 7960 -3300 8020 -3280
rect 7960 -3340 7970 -3300
rect 8010 -3340 8020 -3300
rect 7960 -3365 8020 -3340
rect 7960 -3405 7970 -3365
rect 8010 -3405 8020 -3365
rect 7960 -3435 8020 -3405
rect 7960 -3475 7970 -3435
rect 8010 -3475 8020 -3435
rect 7960 -3505 8020 -3475
rect 7960 -3545 7970 -3505
rect 8010 -3545 8020 -3505
rect 7960 -3575 8020 -3545
rect 7960 -3615 7970 -3575
rect 8010 -3615 8020 -3575
rect 7960 -3640 8020 -3615
rect 7960 -3680 7970 -3640
rect 8010 -3680 8020 -3640
rect 7960 -3700 8020 -3680
rect 7960 -3740 7970 -3700
rect 8010 -3740 8020 -3700
rect 7960 -3765 8020 -3740
rect 7960 -3805 7970 -3765
rect 8010 -3805 8020 -3765
rect 7960 -3835 8020 -3805
rect 7960 -3875 7970 -3835
rect 8010 -3875 8020 -3835
rect 7960 -3905 8020 -3875
rect 7960 -3945 7970 -3905
rect 8010 -3945 8020 -3905
rect 7960 -3975 8020 -3945
rect 7960 -4015 7970 -3975
rect 8010 -4015 8020 -3975
rect 7960 -4040 8020 -4015
rect 7960 -4080 7970 -4040
rect 8010 -4080 8020 -4040
rect 7960 -4100 8020 -4080
rect 7960 -4140 7970 -4100
rect 8010 -4140 8020 -4100
rect 7960 -4165 8020 -4140
rect 7960 -4205 7970 -4165
rect 8010 -4205 8020 -4165
rect 7960 -4235 8020 -4205
rect 7960 -4275 7970 -4235
rect 8010 -4275 8020 -4235
rect 7960 -4305 8020 -4275
rect 7960 -4345 7970 -4305
rect 8010 -4345 8020 -4305
rect 7960 -4375 8020 -4345
rect 7960 -4415 7970 -4375
rect 8010 -4415 8020 -4375
rect 7960 -4440 8020 -4415
rect 7960 -4480 7970 -4440
rect 8010 -4480 8020 -4440
rect 7960 -4490 8020 -4480
rect 8310 -1300 8370 -1290
rect 8310 -1340 8320 -1300
rect 8360 -1340 8370 -1300
rect 8310 -1365 8370 -1340
rect 8310 -1405 8320 -1365
rect 8360 -1405 8370 -1365
rect 8310 -1435 8370 -1405
rect 8310 -1475 8320 -1435
rect 8360 -1475 8370 -1435
rect 8310 -1505 8370 -1475
rect 8310 -1545 8320 -1505
rect 8360 -1545 8370 -1505
rect 8310 -1575 8370 -1545
rect 8310 -1615 8320 -1575
rect 8360 -1615 8370 -1575
rect 8310 -1640 8370 -1615
rect 8310 -1680 8320 -1640
rect 8360 -1680 8370 -1640
rect 8310 -1700 8370 -1680
rect 8310 -1740 8320 -1700
rect 8360 -1740 8370 -1700
rect 8310 -1765 8370 -1740
rect 8310 -1805 8320 -1765
rect 8360 -1805 8370 -1765
rect 8310 -1835 8370 -1805
rect 8310 -1875 8320 -1835
rect 8360 -1875 8370 -1835
rect 8310 -1905 8370 -1875
rect 8310 -1945 8320 -1905
rect 8360 -1945 8370 -1905
rect 8310 -1975 8370 -1945
rect 8310 -2015 8320 -1975
rect 8360 -2015 8370 -1975
rect 8310 -2040 8370 -2015
rect 8310 -2080 8320 -2040
rect 8360 -2080 8370 -2040
rect 8310 -2100 8370 -2080
rect 8310 -2140 8320 -2100
rect 8360 -2140 8370 -2100
rect 8310 -2165 8370 -2140
rect 8310 -2205 8320 -2165
rect 8360 -2205 8370 -2165
rect 8310 -2235 8370 -2205
rect 8310 -2275 8320 -2235
rect 8360 -2275 8370 -2235
rect 8310 -2305 8370 -2275
rect 8310 -2345 8320 -2305
rect 8360 -2345 8370 -2305
rect 8310 -2375 8370 -2345
rect 8310 -2415 8320 -2375
rect 8360 -2415 8370 -2375
rect 8310 -2440 8370 -2415
rect 8310 -2480 8320 -2440
rect 8360 -2480 8370 -2440
rect 8310 -2500 8370 -2480
rect 8310 -2540 8320 -2500
rect 8360 -2540 8370 -2500
rect 8310 -2565 8370 -2540
rect 8310 -2605 8320 -2565
rect 8360 -2605 8370 -2565
rect 8310 -2635 8370 -2605
rect 8310 -2675 8320 -2635
rect 8360 -2675 8370 -2635
rect 8310 -2705 8370 -2675
rect 8310 -2745 8320 -2705
rect 8360 -2745 8370 -2705
rect 8310 -2775 8370 -2745
rect 8310 -2815 8320 -2775
rect 8360 -2815 8370 -2775
rect 8310 -2840 8370 -2815
rect 8310 -2880 8320 -2840
rect 8360 -2880 8370 -2840
rect 8310 -2900 8370 -2880
rect 8310 -2940 8320 -2900
rect 8360 -2940 8370 -2900
rect 8310 -2965 8370 -2940
rect 8310 -3005 8320 -2965
rect 8360 -3005 8370 -2965
rect 8310 -3035 8370 -3005
rect 8310 -3075 8320 -3035
rect 8360 -3075 8370 -3035
rect 8310 -3105 8370 -3075
rect 8310 -3145 8320 -3105
rect 8360 -3145 8370 -3105
rect 8310 -3175 8370 -3145
rect 8310 -3215 8320 -3175
rect 8360 -3215 8370 -3175
rect 8310 -3240 8370 -3215
rect 8310 -3280 8320 -3240
rect 8360 -3280 8370 -3240
rect 8310 -3300 8370 -3280
rect 8310 -3340 8320 -3300
rect 8360 -3340 8370 -3300
rect 8310 -3365 8370 -3340
rect 8310 -3405 8320 -3365
rect 8360 -3405 8370 -3365
rect 8310 -3435 8370 -3405
rect 8310 -3475 8320 -3435
rect 8360 -3475 8370 -3435
rect 8310 -3505 8370 -3475
rect 8310 -3545 8320 -3505
rect 8360 -3545 8370 -3505
rect 8310 -3575 8370 -3545
rect 8310 -3615 8320 -3575
rect 8360 -3615 8370 -3575
rect 8310 -3640 8370 -3615
rect 8310 -3680 8320 -3640
rect 8360 -3680 8370 -3640
rect 8310 -3700 8370 -3680
rect 8310 -3740 8320 -3700
rect 8360 -3740 8370 -3700
rect 8310 -3765 8370 -3740
rect 8310 -3805 8320 -3765
rect 8360 -3805 8370 -3765
rect 8310 -3835 8370 -3805
rect 8310 -3875 8320 -3835
rect 8360 -3875 8370 -3835
rect 8310 -3905 8370 -3875
rect 8310 -3945 8320 -3905
rect 8360 -3945 8370 -3905
rect 8310 -3975 8370 -3945
rect 8310 -4015 8320 -3975
rect 8360 -4015 8370 -3975
rect 8310 -4040 8370 -4015
rect 8310 -4080 8320 -4040
rect 8360 -4080 8370 -4040
rect 8310 -4100 8370 -4080
rect 8310 -4140 8320 -4100
rect 8360 -4140 8370 -4100
rect 8310 -4165 8370 -4140
rect 8310 -4205 8320 -4165
rect 8360 -4205 8370 -4165
rect 8310 -4235 8370 -4205
rect 8310 -4275 8320 -4235
rect 8360 -4275 8370 -4235
rect 8310 -4305 8370 -4275
rect 8310 -4345 8320 -4305
rect 8360 -4345 8370 -4305
rect 8310 -4375 8370 -4345
rect 8310 -4415 8320 -4375
rect 8360 -4415 8370 -4375
rect 8310 -4440 8370 -4415
rect 8310 -4480 8320 -4440
rect 8360 -4480 8370 -4440
rect 8310 -4490 8370 -4480
rect 8660 -1305 8720 -1290
rect 8660 -1335 8675 -1305
rect 8705 -1335 8720 -1305
rect 8660 -1370 8720 -1335
rect 8660 -1400 8675 -1370
rect 8705 -1400 8720 -1370
rect 8660 -1440 8720 -1400
rect 8660 -1470 8675 -1440
rect 8705 -1470 8720 -1440
rect 8660 -1510 8720 -1470
rect 8660 -1540 8675 -1510
rect 8705 -1540 8720 -1510
rect 8660 -1580 8720 -1540
rect 8660 -1610 8675 -1580
rect 8705 -1610 8720 -1580
rect 8660 -1645 8720 -1610
rect 8660 -1675 8675 -1645
rect 8705 -1675 8720 -1645
rect 8660 -1705 8720 -1675
rect 8660 -1735 8675 -1705
rect 8705 -1735 8720 -1705
rect 8660 -1770 8720 -1735
rect 8660 -1800 8675 -1770
rect 8705 -1800 8720 -1770
rect 8660 -1840 8720 -1800
rect 8660 -1870 8675 -1840
rect 8705 -1870 8720 -1840
rect 8660 -1910 8720 -1870
rect 8660 -1940 8675 -1910
rect 8705 -1940 8720 -1910
rect 8660 -1980 8720 -1940
rect 8660 -2010 8675 -1980
rect 8705 -2010 8720 -1980
rect 8660 -2045 8720 -2010
rect 8660 -2075 8675 -2045
rect 8705 -2075 8720 -2045
rect 8660 -2105 8720 -2075
rect 8660 -2135 8675 -2105
rect 8705 -2135 8720 -2105
rect 8660 -2170 8720 -2135
rect 8660 -2200 8675 -2170
rect 8705 -2200 8720 -2170
rect 8660 -2240 8720 -2200
rect 8660 -2270 8675 -2240
rect 8705 -2270 8720 -2240
rect 8660 -2310 8720 -2270
rect 8660 -2340 8675 -2310
rect 8705 -2340 8720 -2310
rect 8660 -2380 8720 -2340
rect 8660 -2410 8675 -2380
rect 8705 -2410 8720 -2380
rect 8660 -2445 8720 -2410
rect 8660 -2475 8675 -2445
rect 8705 -2475 8720 -2445
rect 8660 -2505 8720 -2475
rect 8660 -2535 8675 -2505
rect 8705 -2535 8720 -2505
rect 8660 -2570 8720 -2535
rect 8660 -2600 8675 -2570
rect 8705 -2600 8720 -2570
rect 8660 -2640 8720 -2600
rect 8660 -2670 8675 -2640
rect 8705 -2670 8720 -2640
rect 8660 -2710 8720 -2670
rect 8660 -2740 8675 -2710
rect 8705 -2740 8720 -2710
rect 8660 -2780 8720 -2740
rect 8660 -2810 8675 -2780
rect 8705 -2810 8720 -2780
rect 8660 -2845 8720 -2810
rect 8660 -2875 8675 -2845
rect 8705 -2875 8720 -2845
rect 8660 -2905 8720 -2875
rect 8660 -2935 8675 -2905
rect 8705 -2935 8720 -2905
rect 8660 -2970 8720 -2935
rect 8660 -3000 8675 -2970
rect 8705 -3000 8720 -2970
rect 8660 -3040 8720 -3000
rect 8660 -3070 8675 -3040
rect 8705 -3070 8720 -3040
rect 8660 -3110 8720 -3070
rect 8660 -3140 8675 -3110
rect 8705 -3140 8720 -3110
rect 8660 -3180 8720 -3140
rect 8660 -3210 8675 -3180
rect 8705 -3210 8720 -3180
rect 8660 -3245 8720 -3210
rect 8660 -3275 8675 -3245
rect 8705 -3275 8720 -3245
rect 8660 -3305 8720 -3275
rect 8660 -3335 8675 -3305
rect 8705 -3335 8720 -3305
rect 8660 -3370 8720 -3335
rect 8660 -3400 8675 -3370
rect 8705 -3400 8720 -3370
rect 8660 -3440 8720 -3400
rect 8660 -3470 8675 -3440
rect 8705 -3470 8720 -3440
rect 8660 -3510 8720 -3470
rect 8660 -3540 8675 -3510
rect 8705 -3540 8720 -3510
rect 8660 -3580 8720 -3540
rect 8660 -3610 8675 -3580
rect 8705 -3610 8720 -3580
rect 8660 -3645 8720 -3610
rect 8660 -3675 8675 -3645
rect 8705 -3675 8720 -3645
rect 8660 -3705 8720 -3675
rect 8660 -3735 8675 -3705
rect 8705 -3735 8720 -3705
rect 8660 -3770 8720 -3735
rect 8660 -3800 8675 -3770
rect 8705 -3800 8720 -3770
rect 8660 -3840 8720 -3800
rect 8660 -3870 8675 -3840
rect 8705 -3870 8720 -3840
rect 8660 -3910 8720 -3870
rect 8660 -3940 8675 -3910
rect 8705 -3940 8720 -3910
rect 8660 -3980 8720 -3940
rect 8660 -4010 8675 -3980
rect 8705 -4010 8720 -3980
rect 8660 -4045 8720 -4010
rect 8660 -4075 8675 -4045
rect 8705 -4075 8720 -4045
rect 8660 -4105 8720 -4075
rect 8660 -4135 8675 -4105
rect 8705 -4135 8720 -4105
rect 8660 -4170 8720 -4135
rect 8660 -4200 8675 -4170
rect 8705 -4200 8720 -4170
rect 8660 -4240 8720 -4200
rect 8660 -4270 8675 -4240
rect 8705 -4270 8720 -4240
rect 8660 -4310 8720 -4270
rect 8660 -4340 8675 -4310
rect 8705 -4340 8720 -4310
rect 8660 -4380 8720 -4340
rect 8660 -4410 8675 -4380
rect 8705 -4410 8720 -4380
rect 8660 -4445 8720 -4410
rect 8660 -4475 8675 -4445
rect 8705 -4475 8720 -4445
rect 8660 -4490 8720 -4475
rect 9010 -1305 9070 -1290
rect 9010 -1335 9025 -1305
rect 9055 -1335 9070 -1305
rect 9010 -1370 9070 -1335
rect 9010 -1400 9025 -1370
rect 9055 -1400 9070 -1370
rect 9010 -1440 9070 -1400
rect 9010 -1470 9025 -1440
rect 9055 -1470 9070 -1440
rect 9010 -1510 9070 -1470
rect 9010 -1540 9025 -1510
rect 9055 -1540 9070 -1510
rect 9010 -1580 9070 -1540
rect 9010 -1610 9025 -1580
rect 9055 -1610 9070 -1580
rect 9010 -1645 9070 -1610
rect 9010 -1675 9025 -1645
rect 9055 -1675 9070 -1645
rect 9010 -1705 9070 -1675
rect 9010 -1735 9025 -1705
rect 9055 -1735 9070 -1705
rect 9010 -1770 9070 -1735
rect 9010 -1800 9025 -1770
rect 9055 -1800 9070 -1770
rect 9010 -1840 9070 -1800
rect 9010 -1870 9025 -1840
rect 9055 -1870 9070 -1840
rect 9010 -1910 9070 -1870
rect 9010 -1940 9025 -1910
rect 9055 -1940 9070 -1910
rect 9010 -1980 9070 -1940
rect 9010 -2010 9025 -1980
rect 9055 -2010 9070 -1980
rect 9010 -2045 9070 -2010
rect 9010 -2075 9025 -2045
rect 9055 -2075 9070 -2045
rect 9010 -2105 9070 -2075
rect 9010 -2135 9025 -2105
rect 9055 -2135 9070 -2105
rect 9010 -2170 9070 -2135
rect 9010 -2200 9025 -2170
rect 9055 -2200 9070 -2170
rect 9010 -2240 9070 -2200
rect 9010 -2270 9025 -2240
rect 9055 -2270 9070 -2240
rect 9010 -2310 9070 -2270
rect 9010 -2340 9025 -2310
rect 9055 -2340 9070 -2310
rect 9010 -2380 9070 -2340
rect 9010 -2410 9025 -2380
rect 9055 -2410 9070 -2380
rect 9010 -2445 9070 -2410
rect 9010 -2475 9025 -2445
rect 9055 -2475 9070 -2445
rect 9010 -2505 9070 -2475
rect 9010 -2535 9025 -2505
rect 9055 -2535 9070 -2505
rect 9010 -2570 9070 -2535
rect 9010 -2600 9025 -2570
rect 9055 -2600 9070 -2570
rect 9010 -2640 9070 -2600
rect 9010 -2670 9025 -2640
rect 9055 -2670 9070 -2640
rect 9010 -2710 9070 -2670
rect 9010 -2740 9025 -2710
rect 9055 -2740 9070 -2710
rect 9010 -2780 9070 -2740
rect 9010 -2810 9025 -2780
rect 9055 -2810 9070 -2780
rect 9010 -2845 9070 -2810
rect 9010 -2875 9025 -2845
rect 9055 -2875 9070 -2845
rect 9010 -2905 9070 -2875
rect 9010 -2935 9025 -2905
rect 9055 -2935 9070 -2905
rect 9010 -2970 9070 -2935
rect 9010 -3000 9025 -2970
rect 9055 -3000 9070 -2970
rect 9010 -3040 9070 -3000
rect 9010 -3070 9025 -3040
rect 9055 -3070 9070 -3040
rect 9010 -3110 9070 -3070
rect 9010 -3140 9025 -3110
rect 9055 -3140 9070 -3110
rect 9010 -3180 9070 -3140
rect 9010 -3210 9025 -3180
rect 9055 -3210 9070 -3180
rect 9010 -3245 9070 -3210
rect 9010 -3275 9025 -3245
rect 9055 -3275 9070 -3245
rect 9010 -3305 9070 -3275
rect 9010 -3335 9025 -3305
rect 9055 -3335 9070 -3305
rect 9010 -3370 9070 -3335
rect 9010 -3400 9025 -3370
rect 9055 -3400 9070 -3370
rect 9010 -3440 9070 -3400
rect 9010 -3470 9025 -3440
rect 9055 -3470 9070 -3440
rect 9010 -3510 9070 -3470
rect 9010 -3540 9025 -3510
rect 9055 -3540 9070 -3510
rect 9010 -3580 9070 -3540
rect 9010 -3610 9025 -3580
rect 9055 -3610 9070 -3580
rect 9010 -3645 9070 -3610
rect 9010 -3675 9025 -3645
rect 9055 -3675 9070 -3645
rect 9010 -3705 9070 -3675
rect 9010 -3735 9025 -3705
rect 9055 -3735 9070 -3705
rect 9010 -3770 9070 -3735
rect 9010 -3800 9025 -3770
rect 9055 -3800 9070 -3770
rect 9010 -3840 9070 -3800
rect 9010 -3870 9025 -3840
rect 9055 -3870 9070 -3840
rect 9010 -3910 9070 -3870
rect 9010 -3940 9025 -3910
rect 9055 -3940 9070 -3910
rect 9010 -3980 9070 -3940
rect 9010 -4010 9025 -3980
rect 9055 -4010 9070 -3980
rect 9010 -4045 9070 -4010
rect 9010 -4075 9025 -4045
rect 9055 -4075 9070 -4045
rect 9010 -4105 9070 -4075
rect 9010 -4135 9025 -4105
rect 9055 -4135 9070 -4105
rect 9010 -4170 9070 -4135
rect 9010 -4200 9025 -4170
rect 9055 -4200 9070 -4170
rect 9010 -4240 9070 -4200
rect 9010 -4270 9025 -4240
rect 9055 -4270 9070 -4240
rect 9010 -4310 9070 -4270
rect 9010 -4340 9025 -4310
rect 9055 -4340 9070 -4310
rect 9010 -4380 9070 -4340
rect 9010 -4410 9025 -4380
rect 9055 -4410 9070 -4380
rect 9010 -4445 9070 -4410
rect 9010 -4475 9025 -4445
rect 9055 -4475 9070 -4445
rect 9010 -4490 9070 -4475
rect 12890 -1325 16090 6485
rect 12890 -1375 12925 -1325
rect 12975 -1375 13020 -1325
rect 13070 -1375 13115 -1325
rect 13165 -1375 13215 -1325
rect 13265 -1375 13315 -1325
rect 13365 -1375 13415 -1325
rect 13465 -1375 13510 -1325
rect 13560 -1375 13605 -1325
rect 13655 -1375 13725 -1325
rect 13775 -1375 13820 -1325
rect 13870 -1375 13915 -1325
rect 13965 -1375 14015 -1325
rect 14065 -1375 14115 -1325
rect 14165 -1375 14215 -1325
rect 14265 -1375 14310 -1325
rect 14360 -1375 14405 -1325
rect 14455 -1375 14525 -1325
rect 14575 -1375 14620 -1325
rect 14670 -1375 14715 -1325
rect 14765 -1375 14815 -1325
rect 14865 -1375 14915 -1325
rect 14965 -1375 15015 -1325
rect 15065 -1375 15110 -1325
rect 15160 -1375 15205 -1325
rect 15255 -1375 15325 -1325
rect 15375 -1375 15420 -1325
rect 15470 -1375 15515 -1325
rect 15565 -1375 15615 -1325
rect 15665 -1375 15715 -1325
rect 15765 -1375 15815 -1325
rect 15865 -1375 15910 -1325
rect 15960 -1375 16005 -1325
rect 16055 -1375 16090 -1325
rect 12890 -1415 16090 -1375
rect 12890 -1465 12925 -1415
rect 12975 -1465 13020 -1415
rect 13070 -1465 13115 -1415
rect 13165 -1465 13215 -1415
rect 13265 -1465 13315 -1415
rect 13365 -1465 13415 -1415
rect 13465 -1465 13510 -1415
rect 13560 -1465 13605 -1415
rect 13655 -1465 13725 -1415
rect 13775 -1465 13820 -1415
rect 13870 -1465 13915 -1415
rect 13965 -1465 14015 -1415
rect 14065 -1465 14115 -1415
rect 14165 -1465 14215 -1415
rect 14265 -1465 14310 -1415
rect 14360 -1465 14405 -1415
rect 14455 -1465 14525 -1415
rect 14575 -1465 14620 -1415
rect 14670 -1465 14715 -1415
rect 14765 -1465 14815 -1415
rect 14865 -1465 14915 -1415
rect 14965 -1465 15015 -1415
rect 15065 -1465 15110 -1415
rect 15160 -1465 15205 -1415
rect 15255 -1465 15325 -1415
rect 15375 -1465 15420 -1415
rect 15470 -1465 15515 -1415
rect 15565 -1465 15615 -1415
rect 15665 -1465 15715 -1415
rect 15765 -1465 15815 -1415
rect 15865 -1465 15910 -1415
rect 15960 -1465 16005 -1415
rect 16055 -1465 16090 -1415
rect 12890 -1515 16090 -1465
rect 12890 -1565 12925 -1515
rect 12975 -1565 13020 -1515
rect 13070 -1565 13115 -1515
rect 13165 -1565 13215 -1515
rect 13265 -1565 13315 -1515
rect 13365 -1565 13415 -1515
rect 13465 -1565 13510 -1515
rect 13560 -1565 13605 -1515
rect 13655 -1565 13725 -1515
rect 13775 -1565 13820 -1515
rect 13870 -1565 13915 -1515
rect 13965 -1565 14015 -1515
rect 14065 -1565 14115 -1515
rect 14165 -1565 14215 -1515
rect 14265 -1565 14310 -1515
rect 14360 -1565 14405 -1515
rect 14455 -1565 14525 -1515
rect 14575 -1565 14620 -1515
rect 14670 -1565 14715 -1515
rect 14765 -1565 14815 -1515
rect 14865 -1565 14915 -1515
rect 14965 -1565 15015 -1515
rect 15065 -1565 15110 -1515
rect 15160 -1565 15205 -1515
rect 15255 -1565 15325 -1515
rect 15375 -1565 15420 -1515
rect 15470 -1565 15515 -1515
rect 15565 -1565 15615 -1515
rect 15665 -1565 15715 -1515
rect 15765 -1565 15815 -1515
rect 15865 -1565 15910 -1515
rect 15960 -1565 16005 -1515
rect 16055 -1565 16090 -1515
rect 12890 -1605 16090 -1565
rect 12890 -1655 12925 -1605
rect 12975 -1655 13020 -1605
rect 13070 -1655 13115 -1605
rect 13165 -1655 13215 -1605
rect 13265 -1655 13315 -1605
rect 13365 -1655 13415 -1605
rect 13465 -1655 13510 -1605
rect 13560 -1655 13605 -1605
rect 13655 -1655 13725 -1605
rect 13775 -1655 13820 -1605
rect 13870 -1655 13915 -1605
rect 13965 -1655 14015 -1605
rect 14065 -1655 14115 -1605
rect 14165 -1655 14215 -1605
rect 14265 -1655 14310 -1605
rect 14360 -1655 14405 -1605
rect 14455 -1655 14525 -1605
rect 14575 -1655 14620 -1605
rect 14670 -1655 14715 -1605
rect 14765 -1655 14815 -1605
rect 14865 -1655 14915 -1605
rect 14965 -1655 15015 -1605
rect 15065 -1655 15110 -1605
rect 15160 -1655 15205 -1605
rect 15255 -1655 15325 -1605
rect 15375 -1655 15420 -1605
rect 15470 -1655 15515 -1605
rect 15565 -1655 15615 -1605
rect 15665 -1655 15715 -1605
rect 15765 -1655 15815 -1605
rect 15865 -1655 15910 -1605
rect 15960 -1655 16005 -1605
rect 16055 -1655 16090 -1605
rect 12890 -1725 16090 -1655
rect 12890 -1775 12925 -1725
rect 12975 -1775 13020 -1725
rect 13070 -1775 13115 -1725
rect 13165 -1775 13215 -1725
rect 13265 -1775 13315 -1725
rect 13365 -1775 13415 -1725
rect 13465 -1775 13510 -1725
rect 13560 -1775 13605 -1725
rect 13655 -1775 13725 -1725
rect 13775 -1775 13820 -1725
rect 13870 -1775 13915 -1725
rect 13965 -1775 14015 -1725
rect 14065 -1775 14115 -1725
rect 14165 -1775 14215 -1725
rect 14265 -1775 14310 -1725
rect 14360 -1775 14405 -1725
rect 14455 -1775 14525 -1725
rect 14575 -1775 14620 -1725
rect 14670 -1775 14715 -1725
rect 14765 -1775 14815 -1725
rect 14865 -1775 14915 -1725
rect 14965 -1775 15015 -1725
rect 15065 -1775 15110 -1725
rect 15160 -1775 15205 -1725
rect 15255 -1775 15325 -1725
rect 15375 -1775 15420 -1725
rect 15470 -1775 15515 -1725
rect 15565 -1775 15615 -1725
rect 15665 -1775 15715 -1725
rect 15765 -1775 15815 -1725
rect 15865 -1775 15910 -1725
rect 15960 -1775 16005 -1725
rect 16055 -1775 16090 -1725
rect 12890 -1815 16090 -1775
rect 12890 -1865 12925 -1815
rect 12975 -1865 13020 -1815
rect 13070 -1865 13115 -1815
rect 13165 -1865 13215 -1815
rect 13265 -1865 13315 -1815
rect 13365 -1865 13415 -1815
rect 13465 -1865 13510 -1815
rect 13560 -1865 13605 -1815
rect 13655 -1865 13725 -1815
rect 13775 -1865 13820 -1815
rect 13870 -1865 13915 -1815
rect 13965 -1865 14015 -1815
rect 14065 -1865 14115 -1815
rect 14165 -1865 14215 -1815
rect 14265 -1865 14310 -1815
rect 14360 -1865 14405 -1815
rect 14455 -1865 14525 -1815
rect 14575 -1865 14620 -1815
rect 14670 -1865 14715 -1815
rect 14765 -1865 14815 -1815
rect 14865 -1865 14915 -1815
rect 14965 -1865 15015 -1815
rect 15065 -1865 15110 -1815
rect 15160 -1865 15205 -1815
rect 15255 -1865 15325 -1815
rect 15375 -1865 15420 -1815
rect 15470 -1865 15515 -1815
rect 15565 -1865 15615 -1815
rect 15665 -1865 15715 -1815
rect 15765 -1865 15815 -1815
rect 15865 -1865 15910 -1815
rect 15960 -1865 16005 -1815
rect 16055 -1865 16090 -1815
rect 12890 -1915 16090 -1865
rect 12890 -1965 12925 -1915
rect 12975 -1965 13020 -1915
rect 13070 -1965 13115 -1915
rect 13165 -1965 13215 -1915
rect 13265 -1965 13315 -1915
rect 13365 -1965 13415 -1915
rect 13465 -1965 13510 -1915
rect 13560 -1965 13605 -1915
rect 13655 -1965 13725 -1915
rect 13775 -1965 13820 -1915
rect 13870 -1965 13915 -1915
rect 13965 -1965 14015 -1915
rect 14065 -1965 14115 -1915
rect 14165 -1965 14215 -1915
rect 14265 -1965 14310 -1915
rect 14360 -1965 14405 -1915
rect 14455 -1965 14525 -1915
rect 14575 -1965 14620 -1915
rect 14670 -1965 14715 -1915
rect 14765 -1965 14815 -1915
rect 14865 -1965 14915 -1915
rect 14965 -1965 15015 -1915
rect 15065 -1965 15110 -1915
rect 15160 -1965 15205 -1915
rect 15255 -1965 15325 -1915
rect 15375 -1965 15420 -1915
rect 15470 -1965 15515 -1915
rect 15565 -1965 15615 -1915
rect 15665 -1965 15715 -1915
rect 15765 -1965 15815 -1915
rect 15865 -1965 15910 -1915
rect 15960 -1965 16005 -1915
rect 16055 -1965 16090 -1915
rect 12890 -2005 16090 -1965
rect 12890 -2055 12925 -2005
rect 12975 -2055 13020 -2005
rect 13070 -2055 13115 -2005
rect 13165 -2055 13215 -2005
rect 13265 -2055 13315 -2005
rect 13365 -2055 13415 -2005
rect 13465 -2055 13510 -2005
rect 13560 -2055 13605 -2005
rect 13655 -2055 13725 -2005
rect 13775 -2055 13820 -2005
rect 13870 -2055 13915 -2005
rect 13965 -2055 14015 -2005
rect 14065 -2055 14115 -2005
rect 14165 -2055 14215 -2005
rect 14265 -2055 14310 -2005
rect 14360 -2055 14405 -2005
rect 14455 -2055 14525 -2005
rect 14575 -2055 14620 -2005
rect 14670 -2055 14715 -2005
rect 14765 -2055 14815 -2005
rect 14865 -2055 14915 -2005
rect 14965 -2055 15015 -2005
rect 15065 -2055 15110 -2005
rect 15160 -2055 15205 -2005
rect 15255 -2055 15325 -2005
rect 15375 -2055 15420 -2005
rect 15470 -2055 15515 -2005
rect 15565 -2055 15615 -2005
rect 15665 -2055 15715 -2005
rect 15765 -2055 15815 -2005
rect 15865 -2055 15910 -2005
rect 15960 -2055 16005 -2005
rect 16055 -2055 16090 -2005
rect 12890 -2125 16090 -2055
rect 12890 -2175 12925 -2125
rect 12975 -2175 13020 -2125
rect 13070 -2175 13115 -2125
rect 13165 -2175 13215 -2125
rect 13265 -2175 13315 -2125
rect 13365 -2175 13415 -2125
rect 13465 -2175 13510 -2125
rect 13560 -2175 13605 -2125
rect 13655 -2175 13725 -2125
rect 13775 -2175 13820 -2125
rect 13870 -2175 13915 -2125
rect 13965 -2175 14015 -2125
rect 14065 -2175 14115 -2125
rect 14165 -2175 14215 -2125
rect 14265 -2175 14310 -2125
rect 14360 -2175 14405 -2125
rect 14455 -2175 14525 -2125
rect 14575 -2175 14620 -2125
rect 14670 -2175 14715 -2125
rect 14765 -2175 14815 -2125
rect 14865 -2175 14915 -2125
rect 14965 -2175 15015 -2125
rect 15065 -2175 15110 -2125
rect 15160 -2175 15205 -2125
rect 15255 -2175 15325 -2125
rect 15375 -2175 15420 -2125
rect 15470 -2175 15515 -2125
rect 15565 -2175 15615 -2125
rect 15665 -2175 15715 -2125
rect 15765 -2175 15815 -2125
rect 15865 -2175 15910 -2125
rect 15960 -2175 16005 -2125
rect 16055 -2175 16090 -2125
rect 12890 -2215 16090 -2175
rect 12890 -2265 12925 -2215
rect 12975 -2265 13020 -2215
rect 13070 -2265 13115 -2215
rect 13165 -2265 13215 -2215
rect 13265 -2265 13315 -2215
rect 13365 -2265 13415 -2215
rect 13465 -2265 13510 -2215
rect 13560 -2265 13605 -2215
rect 13655 -2265 13725 -2215
rect 13775 -2265 13820 -2215
rect 13870 -2265 13915 -2215
rect 13965 -2265 14015 -2215
rect 14065 -2265 14115 -2215
rect 14165 -2265 14215 -2215
rect 14265 -2265 14310 -2215
rect 14360 -2265 14405 -2215
rect 14455 -2265 14525 -2215
rect 14575 -2265 14620 -2215
rect 14670 -2265 14715 -2215
rect 14765 -2265 14815 -2215
rect 14865 -2265 14915 -2215
rect 14965 -2265 15015 -2215
rect 15065 -2265 15110 -2215
rect 15160 -2265 15205 -2215
rect 15255 -2265 15325 -2215
rect 15375 -2265 15420 -2215
rect 15470 -2265 15515 -2215
rect 15565 -2265 15615 -2215
rect 15665 -2265 15715 -2215
rect 15765 -2265 15815 -2215
rect 15865 -2265 15910 -2215
rect 15960 -2265 16005 -2215
rect 16055 -2265 16090 -2215
rect 12890 -2315 16090 -2265
rect 12890 -2365 12925 -2315
rect 12975 -2365 13020 -2315
rect 13070 -2365 13115 -2315
rect 13165 -2365 13215 -2315
rect 13265 -2365 13315 -2315
rect 13365 -2365 13415 -2315
rect 13465 -2365 13510 -2315
rect 13560 -2365 13605 -2315
rect 13655 -2365 13725 -2315
rect 13775 -2365 13820 -2315
rect 13870 -2365 13915 -2315
rect 13965 -2365 14015 -2315
rect 14065 -2365 14115 -2315
rect 14165 -2365 14215 -2315
rect 14265 -2365 14310 -2315
rect 14360 -2365 14405 -2315
rect 14455 -2365 14525 -2315
rect 14575 -2365 14620 -2315
rect 14670 -2365 14715 -2315
rect 14765 -2365 14815 -2315
rect 14865 -2365 14915 -2315
rect 14965 -2365 15015 -2315
rect 15065 -2365 15110 -2315
rect 15160 -2365 15205 -2315
rect 15255 -2365 15325 -2315
rect 15375 -2365 15420 -2315
rect 15470 -2365 15515 -2315
rect 15565 -2365 15615 -2315
rect 15665 -2365 15715 -2315
rect 15765 -2365 15815 -2315
rect 15865 -2365 15910 -2315
rect 15960 -2365 16005 -2315
rect 16055 -2365 16090 -2315
rect 12890 -2405 16090 -2365
rect 12890 -2455 12925 -2405
rect 12975 -2455 13020 -2405
rect 13070 -2455 13115 -2405
rect 13165 -2455 13215 -2405
rect 13265 -2455 13315 -2405
rect 13365 -2455 13415 -2405
rect 13465 -2455 13510 -2405
rect 13560 -2455 13605 -2405
rect 13655 -2455 13725 -2405
rect 13775 -2455 13820 -2405
rect 13870 -2455 13915 -2405
rect 13965 -2455 14015 -2405
rect 14065 -2455 14115 -2405
rect 14165 -2455 14215 -2405
rect 14265 -2455 14310 -2405
rect 14360 -2455 14405 -2405
rect 14455 -2455 14525 -2405
rect 14575 -2455 14620 -2405
rect 14670 -2455 14715 -2405
rect 14765 -2455 14815 -2405
rect 14865 -2455 14915 -2405
rect 14965 -2455 15015 -2405
rect 15065 -2455 15110 -2405
rect 15160 -2455 15205 -2405
rect 15255 -2455 15325 -2405
rect 15375 -2455 15420 -2405
rect 15470 -2455 15515 -2405
rect 15565 -2455 15615 -2405
rect 15665 -2455 15715 -2405
rect 15765 -2455 15815 -2405
rect 15865 -2455 15910 -2405
rect 15960 -2455 16005 -2405
rect 16055 -2455 16090 -2405
rect 12890 -2525 16090 -2455
rect 12890 -2575 12925 -2525
rect 12975 -2575 13020 -2525
rect 13070 -2575 13115 -2525
rect 13165 -2575 13215 -2525
rect 13265 -2575 13315 -2525
rect 13365 -2575 13415 -2525
rect 13465 -2575 13510 -2525
rect 13560 -2575 13605 -2525
rect 13655 -2575 13725 -2525
rect 13775 -2575 13820 -2525
rect 13870 -2575 13915 -2525
rect 13965 -2575 14015 -2525
rect 14065 -2575 14115 -2525
rect 14165 -2575 14215 -2525
rect 14265 -2575 14310 -2525
rect 14360 -2575 14405 -2525
rect 14455 -2575 14525 -2525
rect 14575 -2575 14620 -2525
rect 14670 -2575 14715 -2525
rect 14765 -2575 14815 -2525
rect 14865 -2575 14915 -2525
rect 14965 -2575 15015 -2525
rect 15065 -2575 15110 -2525
rect 15160 -2575 15205 -2525
rect 15255 -2575 15325 -2525
rect 15375 -2575 15420 -2525
rect 15470 -2575 15515 -2525
rect 15565 -2575 15615 -2525
rect 15665 -2575 15715 -2525
rect 15765 -2575 15815 -2525
rect 15865 -2575 15910 -2525
rect 15960 -2575 16005 -2525
rect 16055 -2575 16090 -2525
rect 12890 -2615 16090 -2575
rect 12890 -2665 12925 -2615
rect 12975 -2665 13020 -2615
rect 13070 -2665 13115 -2615
rect 13165 -2665 13215 -2615
rect 13265 -2665 13315 -2615
rect 13365 -2665 13415 -2615
rect 13465 -2665 13510 -2615
rect 13560 -2665 13605 -2615
rect 13655 -2665 13725 -2615
rect 13775 -2665 13820 -2615
rect 13870 -2665 13915 -2615
rect 13965 -2665 14015 -2615
rect 14065 -2665 14115 -2615
rect 14165 -2665 14215 -2615
rect 14265 -2665 14310 -2615
rect 14360 -2665 14405 -2615
rect 14455 -2665 14525 -2615
rect 14575 -2665 14620 -2615
rect 14670 -2665 14715 -2615
rect 14765 -2665 14815 -2615
rect 14865 -2665 14915 -2615
rect 14965 -2665 15015 -2615
rect 15065 -2665 15110 -2615
rect 15160 -2665 15205 -2615
rect 15255 -2665 15325 -2615
rect 15375 -2665 15420 -2615
rect 15470 -2665 15515 -2615
rect 15565 -2665 15615 -2615
rect 15665 -2665 15715 -2615
rect 15765 -2665 15815 -2615
rect 15865 -2665 15910 -2615
rect 15960 -2665 16005 -2615
rect 16055 -2665 16090 -2615
rect 12890 -2715 16090 -2665
rect 12890 -2765 12925 -2715
rect 12975 -2765 13020 -2715
rect 13070 -2765 13115 -2715
rect 13165 -2765 13215 -2715
rect 13265 -2765 13315 -2715
rect 13365 -2765 13415 -2715
rect 13465 -2765 13510 -2715
rect 13560 -2765 13605 -2715
rect 13655 -2765 13725 -2715
rect 13775 -2765 13820 -2715
rect 13870 -2765 13915 -2715
rect 13965 -2765 14015 -2715
rect 14065 -2765 14115 -2715
rect 14165 -2765 14215 -2715
rect 14265 -2765 14310 -2715
rect 14360 -2765 14405 -2715
rect 14455 -2765 14525 -2715
rect 14575 -2765 14620 -2715
rect 14670 -2765 14715 -2715
rect 14765 -2765 14815 -2715
rect 14865 -2765 14915 -2715
rect 14965 -2765 15015 -2715
rect 15065 -2765 15110 -2715
rect 15160 -2765 15205 -2715
rect 15255 -2765 15325 -2715
rect 15375 -2765 15420 -2715
rect 15470 -2765 15515 -2715
rect 15565 -2765 15615 -2715
rect 15665 -2765 15715 -2715
rect 15765 -2765 15815 -2715
rect 15865 -2765 15910 -2715
rect 15960 -2765 16005 -2715
rect 16055 -2765 16090 -2715
rect 12890 -2805 16090 -2765
rect 12890 -2855 12925 -2805
rect 12975 -2855 13020 -2805
rect 13070 -2855 13115 -2805
rect 13165 -2855 13215 -2805
rect 13265 -2855 13315 -2805
rect 13365 -2855 13415 -2805
rect 13465 -2855 13510 -2805
rect 13560 -2855 13605 -2805
rect 13655 -2855 13725 -2805
rect 13775 -2855 13820 -2805
rect 13870 -2855 13915 -2805
rect 13965 -2855 14015 -2805
rect 14065 -2855 14115 -2805
rect 14165 -2855 14215 -2805
rect 14265 -2855 14310 -2805
rect 14360 -2855 14405 -2805
rect 14455 -2855 14525 -2805
rect 14575 -2855 14620 -2805
rect 14670 -2855 14715 -2805
rect 14765 -2855 14815 -2805
rect 14865 -2855 14915 -2805
rect 14965 -2855 15015 -2805
rect 15065 -2855 15110 -2805
rect 15160 -2855 15205 -2805
rect 15255 -2855 15325 -2805
rect 15375 -2855 15420 -2805
rect 15470 -2855 15515 -2805
rect 15565 -2855 15615 -2805
rect 15665 -2855 15715 -2805
rect 15765 -2855 15815 -2805
rect 15865 -2855 15910 -2805
rect 15960 -2855 16005 -2805
rect 16055 -2855 16090 -2805
rect 12890 -2925 16090 -2855
rect 12890 -2975 12925 -2925
rect 12975 -2975 13020 -2925
rect 13070 -2975 13115 -2925
rect 13165 -2975 13215 -2925
rect 13265 -2975 13315 -2925
rect 13365 -2975 13415 -2925
rect 13465 -2975 13510 -2925
rect 13560 -2975 13605 -2925
rect 13655 -2975 13725 -2925
rect 13775 -2975 13820 -2925
rect 13870 -2975 13915 -2925
rect 13965 -2975 14015 -2925
rect 14065 -2975 14115 -2925
rect 14165 -2975 14215 -2925
rect 14265 -2975 14310 -2925
rect 14360 -2975 14405 -2925
rect 14455 -2975 14525 -2925
rect 14575 -2975 14620 -2925
rect 14670 -2975 14715 -2925
rect 14765 -2975 14815 -2925
rect 14865 -2975 14915 -2925
rect 14965 -2975 15015 -2925
rect 15065 -2975 15110 -2925
rect 15160 -2975 15205 -2925
rect 15255 -2975 15325 -2925
rect 15375 -2975 15420 -2925
rect 15470 -2975 15515 -2925
rect 15565 -2975 15615 -2925
rect 15665 -2975 15715 -2925
rect 15765 -2975 15815 -2925
rect 15865 -2975 15910 -2925
rect 15960 -2975 16005 -2925
rect 16055 -2975 16090 -2925
rect 12890 -3015 16090 -2975
rect 12890 -3065 12925 -3015
rect 12975 -3065 13020 -3015
rect 13070 -3065 13115 -3015
rect 13165 -3065 13215 -3015
rect 13265 -3065 13315 -3015
rect 13365 -3065 13415 -3015
rect 13465 -3065 13510 -3015
rect 13560 -3065 13605 -3015
rect 13655 -3065 13725 -3015
rect 13775 -3065 13820 -3015
rect 13870 -3065 13915 -3015
rect 13965 -3065 14015 -3015
rect 14065 -3065 14115 -3015
rect 14165 -3065 14215 -3015
rect 14265 -3065 14310 -3015
rect 14360 -3065 14405 -3015
rect 14455 -3065 14525 -3015
rect 14575 -3065 14620 -3015
rect 14670 -3065 14715 -3015
rect 14765 -3065 14815 -3015
rect 14865 -3065 14915 -3015
rect 14965 -3065 15015 -3015
rect 15065 -3065 15110 -3015
rect 15160 -3065 15205 -3015
rect 15255 -3065 15325 -3015
rect 15375 -3065 15420 -3015
rect 15470 -3065 15515 -3015
rect 15565 -3065 15615 -3015
rect 15665 -3065 15715 -3015
rect 15765 -3065 15815 -3015
rect 15865 -3065 15910 -3015
rect 15960 -3065 16005 -3015
rect 16055 -3065 16090 -3015
rect 12890 -3115 16090 -3065
rect 12890 -3165 12925 -3115
rect 12975 -3165 13020 -3115
rect 13070 -3165 13115 -3115
rect 13165 -3165 13215 -3115
rect 13265 -3165 13315 -3115
rect 13365 -3165 13415 -3115
rect 13465 -3165 13510 -3115
rect 13560 -3165 13605 -3115
rect 13655 -3165 13725 -3115
rect 13775 -3165 13820 -3115
rect 13870 -3165 13915 -3115
rect 13965 -3165 14015 -3115
rect 14065 -3165 14115 -3115
rect 14165 -3165 14215 -3115
rect 14265 -3165 14310 -3115
rect 14360 -3165 14405 -3115
rect 14455 -3165 14525 -3115
rect 14575 -3165 14620 -3115
rect 14670 -3165 14715 -3115
rect 14765 -3165 14815 -3115
rect 14865 -3165 14915 -3115
rect 14965 -3165 15015 -3115
rect 15065 -3165 15110 -3115
rect 15160 -3165 15205 -3115
rect 15255 -3165 15325 -3115
rect 15375 -3165 15420 -3115
rect 15470 -3165 15515 -3115
rect 15565 -3165 15615 -3115
rect 15665 -3165 15715 -3115
rect 15765 -3165 15815 -3115
rect 15865 -3165 15910 -3115
rect 15960 -3165 16005 -3115
rect 16055 -3165 16090 -3115
rect 12890 -3205 16090 -3165
rect 12890 -3255 12925 -3205
rect 12975 -3255 13020 -3205
rect 13070 -3255 13115 -3205
rect 13165 -3255 13215 -3205
rect 13265 -3255 13315 -3205
rect 13365 -3255 13415 -3205
rect 13465 -3255 13510 -3205
rect 13560 -3255 13605 -3205
rect 13655 -3255 13725 -3205
rect 13775 -3255 13820 -3205
rect 13870 -3255 13915 -3205
rect 13965 -3255 14015 -3205
rect 14065 -3255 14115 -3205
rect 14165 -3255 14215 -3205
rect 14265 -3255 14310 -3205
rect 14360 -3255 14405 -3205
rect 14455 -3255 14525 -3205
rect 14575 -3255 14620 -3205
rect 14670 -3255 14715 -3205
rect 14765 -3255 14815 -3205
rect 14865 -3255 14915 -3205
rect 14965 -3255 15015 -3205
rect 15065 -3255 15110 -3205
rect 15160 -3255 15205 -3205
rect 15255 -3255 15325 -3205
rect 15375 -3255 15420 -3205
rect 15470 -3255 15515 -3205
rect 15565 -3255 15615 -3205
rect 15665 -3255 15715 -3205
rect 15765 -3255 15815 -3205
rect 15865 -3255 15910 -3205
rect 15960 -3255 16005 -3205
rect 16055 -3255 16090 -3205
rect 12890 -3325 16090 -3255
rect 12890 -3375 12925 -3325
rect 12975 -3375 13020 -3325
rect 13070 -3375 13115 -3325
rect 13165 -3375 13215 -3325
rect 13265 -3375 13315 -3325
rect 13365 -3375 13415 -3325
rect 13465 -3375 13510 -3325
rect 13560 -3375 13605 -3325
rect 13655 -3375 13725 -3325
rect 13775 -3375 13820 -3325
rect 13870 -3375 13915 -3325
rect 13965 -3375 14015 -3325
rect 14065 -3375 14115 -3325
rect 14165 -3375 14215 -3325
rect 14265 -3375 14310 -3325
rect 14360 -3375 14405 -3325
rect 14455 -3375 14525 -3325
rect 14575 -3375 14620 -3325
rect 14670 -3375 14715 -3325
rect 14765 -3375 14815 -3325
rect 14865 -3375 14915 -3325
rect 14965 -3375 15015 -3325
rect 15065 -3375 15110 -3325
rect 15160 -3375 15205 -3325
rect 15255 -3375 15325 -3325
rect 15375 -3375 15420 -3325
rect 15470 -3375 15515 -3325
rect 15565 -3375 15615 -3325
rect 15665 -3375 15715 -3325
rect 15765 -3375 15815 -3325
rect 15865 -3375 15910 -3325
rect 15960 -3375 16005 -3325
rect 16055 -3375 16090 -3325
rect 12890 -3415 16090 -3375
rect 12890 -3465 12925 -3415
rect 12975 -3465 13020 -3415
rect 13070 -3465 13115 -3415
rect 13165 -3465 13215 -3415
rect 13265 -3465 13315 -3415
rect 13365 -3465 13415 -3415
rect 13465 -3465 13510 -3415
rect 13560 -3465 13605 -3415
rect 13655 -3465 13725 -3415
rect 13775 -3465 13820 -3415
rect 13870 -3465 13915 -3415
rect 13965 -3465 14015 -3415
rect 14065 -3465 14115 -3415
rect 14165 -3465 14215 -3415
rect 14265 -3465 14310 -3415
rect 14360 -3465 14405 -3415
rect 14455 -3465 14525 -3415
rect 14575 -3465 14620 -3415
rect 14670 -3465 14715 -3415
rect 14765 -3465 14815 -3415
rect 14865 -3465 14915 -3415
rect 14965 -3465 15015 -3415
rect 15065 -3465 15110 -3415
rect 15160 -3465 15205 -3415
rect 15255 -3465 15325 -3415
rect 15375 -3465 15420 -3415
rect 15470 -3465 15515 -3415
rect 15565 -3465 15615 -3415
rect 15665 -3465 15715 -3415
rect 15765 -3465 15815 -3415
rect 15865 -3465 15910 -3415
rect 15960 -3465 16005 -3415
rect 16055 -3465 16090 -3415
rect 12890 -3515 16090 -3465
rect 12890 -3565 12925 -3515
rect 12975 -3565 13020 -3515
rect 13070 -3565 13115 -3515
rect 13165 -3565 13215 -3515
rect 13265 -3565 13315 -3515
rect 13365 -3565 13415 -3515
rect 13465 -3565 13510 -3515
rect 13560 -3565 13605 -3515
rect 13655 -3565 13725 -3515
rect 13775 -3565 13820 -3515
rect 13870 -3565 13915 -3515
rect 13965 -3565 14015 -3515
rect 14065 -3565 14115 -3515
rect 14165 -3565 14215 -3515
rect 14265 -3565 14310 -3515
rect 14360 -3565 14405 -3515
rect 14455 -3565 14525 -3515
rect 14575 -3565 14620 -3515
rect 14670 -3565 14715 -3515
rect 14765 -3565 14815 -3515
rect 14865 -3565 14915 -3515
rect 14965 -3565 15015 -3515
rect 15065 -3565 15110 -3515
rect 15160 -3565 15205 -3515
rect 15255 -3565 15325 -3515
rect 15375 -3565 15420 -3515
rect 15470 -3565 15515 -3515
rect 15565 -3565 15615 -3515
rect 15665 -3565 15715 -3515
rect 15765 -3565 15815 -3515
rect 15865 -3565 15910 -3515
rect 15960 -3565 16005 -3515
rect 16055 -3565 16090 -3515
rect 12890 -3605 16090 -3565
rect 12890 -3655 12925 -3605
rect 12975 -3655 13020 -3605
rect 13070 -3655 13115 -3605
rect 13165 -3655 13215 -3605
rect 13265 -3655 13315 -3605
rect 13365 -3655 13415 -3605
rect 13465 -3655 13510 -3605
rect 13560 -3655 13605 -3605
rect 13655 -3655 13725 -3605
rect 13775 -3655 13820 -3605
rect 13870 -3655 13915 -3605
rect 13965 -3655 14015 -3605
rect 14065 -3655 14115 -3605
rect 14165 -3655 14215 -3605
rect 14265 -3655 14310 -3605
rect 14360 -3655 14405 -3605
rect 14455 -3655 14525 -3605
rect 14575 -3655 14620 -3605
rect 14670 -3655 14715 -3605
rect 14765 -3655 14815 -3605
rect 14865 -3655 14915 -3605
rect 14965 -3655 15015 -3605
rect 15065 -3655 15110 -3605
rect 15160 -3655 15205 -3605
rect 15255 -3655 15325 -3605
rect 15375 -3655 15420 -3605
rect 15470 -3655 15515 -3605
rect 15565 -3655 15615 -3605
rect 15665 -3655 15715 -3605
rect 15765 -3655 15815 -3605
rect 15865 -3655 15910 -3605
rect 15960 -3655 16005 -3605
rect 16055 -3655 16090 -3605
rect 12890 -3725 16090 -3655
rect 12890 -3775 12925 -3725
rect 12975 -3775 13020 -3725
rect 13070 -3775 13115 -3725
rect 13165 -3775 13215 -3725
rect 13265 -3775 13315 -3725
rect 13365 -3775 13415 -3725
rect 13465 -3775 13510 -3725
rect 13560 -3775 13605 -3725
rect 13655 -3775 13725 -3725
rect 13775 -3775 13820 -3725
rect 13870 -3775 13915 -3725
rect 13965 -3775 14015 -3725
rect 14065 -3775 14115 -3725
rect 14165 -3775 14215 -3725
rect 14265 -3775 14310 -3725
rect 14360 -3775 14405 -3725
rect 14455 -3775 14525 -3725
rect 14575 -3775 14620 -3725
rect 14670 -3775 14715 -3725
rect 14765 -3775 14815 -3725
rect 14865 -3775 14915 -3725
rect 14965 -3775 15015 -3725
rect 15065 -3775 15110 -3725
rect 15160 -3775 15205 -3725
rect 15255 -3775 15325 -3725
rect 15375 -3775 15420 -3725
rect 15470 -3775 15515 -3725
rect 15565 -3775 15615 -3725
rect 15665 -3775 15715 -3725
rect 15765 -3775 15815 -3725
rect 15865 -3775 15910 -3725
rect 15960 -3775 16005 -3725
rect 16055 -3775 16090 -3725
rect 12890 -3815 16090 -3775
rect 12890 -3865 12925 -3815
rect 12975 -3865 13020 -3815
rect 13070 -3865 13115 -3815
rect 13165 -3865 13215 -3815
rect 13265 -3865 13315 -3815
rect 13365 -3865 13415 -3815
rect 13465 -3865 13510 -3815
rect 13560 -3865 13605 -3815
rect 13655 -3865 13725 -3815
rect 13775 -3865 13820 -3815
rect 13870 -3865 13915 -3815
rect 13965 -3865 14015 -3815
rect 14065 -3865 14115 -3815
rect 14165 -3865 14215 -3815
rect 14265 -3865 14310 -3815
rect 14360 -3865 14405 -3815
rect 14455 -3865 14525 -3815
rect 14575 -3865 14620 -3815
rect 14670 -3865 14715 -3815
rect 14765 -3865 14815 -3815
rect 14865 -3865 14915 -3815
rect 14965 -3865 15015 -3815
rect 15065 -3865 15110 -3815
rect 15160 -3865 15205 -3815
rect 15255 -3865 15325 -3815
rect 15375 -3865 15420 -3815
rect 15470 -3865 15515 -3815
rect 15565 -3865 15615 -3815
rect 15665 -3865 15715 -3815
rect 15765 -3865 15815 -3815
rect 15865 -3865 15910 -3815
rect 15960 -3865 16005 -3815
rect 16055 -3865 16090 -3815
rect 12890 -3915 16090 -3865
rect 12890 -3965 12925 -3915
rect 12975 -3965 13020 -3915
rect 13070 -3965 13115 -3915
rect 13165 -3965 13215 -3915
rect 13265 -3965 13315 -3915
rect 13365 -3965 13415 -3915
rect 13465 -3965 13510 -3915
rect 13560 -3965 13605 -3915
rect 13655 -3965 13725 -3915
rect 13775 -3965 13820 -3915
rect 13870 -3965 13915 -3915
rect 13965 -3965 14015 -3915
rect 14065 -3965 14115 -3915
rect 14165 -3965 14215 -3915
rect 14265 -3965 14310 -3915
rect 14360 -3965 14405 -3915
rect 14455 -3965 14525 -3915
rect 14575 -3965 14620 -3915
rect 14670 -3965 14715 -3915
rect 14765 -3965 14815 -3915
rect 14865 -3965 14915 -3915
rect 14965 -3965 15015 -3915
rect 15065 -3965 15110 -3915
rect 15160 -3965 15205 -3915
rect 15255 -3965 15325 -3915
rect 15375 -3965 15420 -3915
rect 15470 -3965 15515 -3915
rect 15565 -3965 15615 -3915
rect 15665 -3965 15715 -3915
rect 15765 -3965 15815 -3915
rect 15865 -3965 15910 -3915
rect 15960 -3965 16005 -3915
rect 16055 -3965 16090 -3915
rect 12890 -4005 16090 -3965
rect 12890 -4055 12925 -4005
rect 12975 -4055 13020 -4005
rect 13070 -4055 13115 -4005
rect 13165 -4055 13215 -4005
rect 13265 -4055 13315 -4005
rect 13365 -4055 13415 -4005
rect 13465 -4055 13510 -4005
rect 13560 -4055 13605 -4005
rect 13655 -4055 13725 -4005
rect 13775 -4055 13820 -4005
rect 13870 -4055 13915 -4005
rect 13965 -4055 14015 -4005
rect 14065 -4055 14115 -4005
rect 14165 -4055 14215 -4005
rect 14265 -4055 14310 -4005
rect 14360 -4055 14405 -4005
rect 14455 -4055 14525 -4005
rect 14575 -4055 14620 -4005
rect 14670 -4055 14715 -4005
rect 14765 -4055 14815 -4005
rect 14865 -4055 14915 -4005
rect 14965 -4055 15015 -4005
rect 15065 -4055 15110 -4005
rect 15160 -4055 15205 -4005
rect 15255 -4055 15325 -4005
rect 15375 -4055 15420 -4005
rect 15470 -4055 15515 -4005
rect 15565 -4055 15615 -4005
rect 15665 -4055 15715 -4005
rect 15765 -4055 15815 -4005
rect 15865 -4055 15910 -4005
rect 15960 -4055 16005 -4005
rect 16055 -4055 16090 -4005
rect 12890 -4125 16090 -4055
rect 12890 -4175 12925 -4125
rect 12975 -4175 13020 -4125
rect 13070 -4175 13115 -4125
rect 13165 -4175 13215 -4125
rect 13265 -4175 13315 -4125
rect 13365 -4175 13415 -4125
rect 13465 -4175 13510 -4125
rect 13560 -4175 13605 -4125
rect 13655 -4175 13725 -4125
rect 13775 -4175 13820 -4125
rect 13870 -4175 13915 -4125
rect 13965 -4175 14015 -4125
rect 14065 -4175 14115 -4125
rect 14165 -4175 14215 -4125
rect 14265 -4175 14310 -4125
rect 14360 -4175 14405 -4125
rect 14455 -4175 14525 -4125
rect 14575 -4175 14620 -4125
rect 14670 -4175 14715 -4125
rect 14765 -4175 14815 -4125
rect 14865 -4175 14915 -4125
rect 14965 -4175 15015 -4125
rect 15065 -4175 15110 -4125
rect 15160 -4175 15205 -4125
rect 15255 -4175 15325 -4125
rect 15375 -4175 15420 -4125
rect 15470 -4175 15515 -4125
rect 15565 -4175 15615 -4125
rect 15665 -4175 15715 -4125
rect 15765 -4175 15815 -4125
rect 15865 -4175 15910 -4125
rect 15960 -4175 16005 -4125
rect 16055 -4175 16090 -4125
rect 12890 -4215 16090 -4175
rect 12890 -4265 12925 -4215
rect 12975 -4265 13020 -4215
rect 13070 -4265 13115 -4215
rect 13165 -4265 13215 -4215
rect 13265 -4265 13315 -4215
rect 13365 -4265 13415 -4215
rect 13465 -4265 13510 -4215
rect 13560 -4265 13605 -4215
rect 13655 -4265 13725 -4215
rect 13775 -4265 13820 -4215
rect 13870 -4265 13915 -4215
rect 13965 -4265 14015 -4215
rect 14065 -4265 14115 -4215
rect 14165 -4265 14215 -4215
rect 14265 -4265 14310 -4215
rect 14360 -4265 14405 -4215
rect 14455 -4265 14525 -4215
rect 14575 -4265 14620 -4215
rect 14670 -4265 14715 -4215
rect 14765 -4265 14815 -4215
rect 14865 -4265 14915 -4215
rect 14965 -4265 15015 -4215
rect 15065 -4265 15110 -4215
rect 15160 -4265 15205 -4215
rect 15255 -4265 15325 -4215
rect 15375 -4265 15420 -4215
rect 15470 -4265 15515 -4215
rect 15565 -4265 15615 -4215
rect 15665 -4265 15715 -4215
rect 15765 -4265 15815 -4215
rect 15865 -4265 15910 -4215
rect 15960 -4265 16005 -4215
rect 16055 -4265 16090 -4215
rect 12890 -4315 16090 -4265
rect 12890 -4365 12925 -4315
rect 12975 -4365 13020 -4315
rect 13070 -4365 13115 -4315
rect 13165 -4365 13215 -4315
rect 13265 -4365 13315 -4315
rect 13365 -4365 13415 -4315
rect 13465 -4365 13510 -4315
rect 13560 -4365 13605 -4315
rect 13655 -4365 13725 -4315
rect 13775 -4365 13820 -4315
rect 13870 -4365 13915 -4315
rect 13965 -4365 14015 -4315
rect 14065 -4365 14115 -4315
rect 14165 -4365 14215 -4315
rect 14265 -4365 14310 -4315
rect 14360 -4365 14405 -4315
rect 14455 -4365 14525 -4315
rect 14575 -4365 14620 -4315
rect 14670 -4365 14715 -4315
rect 14765 -4365 14815 -4315
rect 14865 -4365 14915 -4315
rect 14965 -4365 15015 -4315
rect 15065 -4365 15110 -4315
rect 15160 -4365 15205 -4315
rect 15255 -4365 15325 -4315
rect 15375 -4365 15420 -4315
rect 15470 -4365 15515 -4315
rect 15565 -4365 15615 -4315
rect 15665 -4365 15715 -4315
rect 15765 -4365 15815 -4315
rect 15865 -4365 15910 -4315
rect 15960 -4365 16005 -4315
rect 16055 -4365 16090 -4315
rect 12890 -4405 16090 -4365
rect 12890 -4455 12925 -4405
rect 12975 -4455 13020 -4405
rect 13070 -4455 13115 -4405
rect 13165 -4455 13215 -4405
rect 13265 -4455 13315 -4405
rect 13365 -4455 13415 -4405
rect 13465 -4455 13510 -4405
rect 13560 -4455 13605 -4405
rect 13655 -4455 13725 -4405
rect 13775 -4455 13820 -4405
rect 13870 -4455 13915 -4405
rect 13965 -4455 14015 -4405
rect 14065 -4455 14115 -4405
rect 14165 -4455 14215 -4405
rect 14265 -4455 14310 -4405
rect 14360 -4455 14405 -4405
rect 14455 -4455 14525 -4405
rect 14575 -4455 14620 -4405
rect 14670 -4455 14715 -4405
rect 14765 -4455 14815 -4405
rect 14865 -4455 14915 -4405
rect 14965 -4455 15015 -4405
rect 15065 -4455 15110 -4405
rect 15160 -4455 15205 -4405
rect 15255 -4455 15325 -4405
rect 15375 -4455 15420 -4405
rect 15470 -4455 15515 -4405
rect 15565 -4455 15615 -4405
rect 15665 -4455 15715 -4405
rect 15765 -4455 15815 -4405
rect 15865 -4455 15910 -4405
rect 15960 -4455 16005 -4405
rect 16055 -4455 16090 -4405
rect 12890 -4490 16090 -4455
<< via3 >>
rect 2190 20910 2230 20915
rect 2190 20880 2195 20910
rect 2195 20880 2225 20910
rect 2225 20880 2230 20910
rect 2190 20875 2230 20880
rect 2190 20845 2230 20850
rect 2190 20815 2195 20845
rect 2195 20815 2225 20845
rect 2225 20815 2230 20845
rect 2190 20810 2230 20815
rect 2190 20775 2230 20780
rect 2190 20745 2195 20775
rect 2195 20745 2225 20775
rect 2225 20745 2230 20775
rect 2190 20740 2230 20745
rect 2190 20705 2230 20710
rect 2190 20675 2195 20705
rect 2195 20675 2225 20705
rect 2225 20675 2230 20705
rect 2190 20670 2230 20675
rect 2190 20635 2230 20640
rect 2190 20605 2195 20635
rect 2195 20605 2225 20635
rect 2225 20605 2230 20635
rect 2190 20600 2230 20605
rect 2190 20570 2230 20575
rect 2190 20540 2195 20570
rect 2195 20540 2225 20570
rect 2225 20540 2230 20570
rect 2190 20535 2230 20540
rect 2190 20510 2230 20515
rect 2190 20480 2195 20510
rect 2195 20480 2225 20510
rect 2225 20480 2230 20510
rect 2190 20475 2230 20480
rect 2190 20445 2230 20450
rect 2190 20415 2195 20445
rect 2195 20415 2225 20445
rect 2225 20415 2230 20445
rect 2190 20410 2230 20415
rect 2190 20375 2230 20380
rect 2190 20345 2195 20375
rect 2195 20345 2225 20375
rect 2225 20345 2230 20375
rect 2190 20340 2230 20345
rect 2190 20305 2230 20310
rect 2190 20275 2195 20305
rect 2195 20275 2225 20305
rect 2225 20275 2230 20305
rect 2190 20270 2230 20275
rect 2190 20235 2230 20240
rect 2190 20205 2195 20235
rect 2195 20205 2225 20235
rect 2225 20205 2230 20235
rect 2190 20200 2230 20205
rect 2190 20170 2230 20175
rect 2190 20140 2195 20170
rect 2195 20140 2225 20170
rect 2225 20140 2230 20170
rect 2190 20135 2230 20140
rect 2190 20110 2230 20115
rect 2190 20080 2195 20110
rect 2195 20080 2225 20110
rect 2225 20080 2230 20110
rect 2190 20075 2230 20080
rect 2190 20045 2230 20050
rect 2190 20015 2195 20045
rect 2195 20015 2225 20045
rect 2225 20015 2230 20045
rect 2190 20010 2230 20015
rect 2190 19975 2230 19980
rect 2190 19945 2195 19975
rect 2195 19945 2225 19975
rect 2225 19945 2230 19975
rect 2190 19940 2230 19945
rect 2190 19905 2230 19910
rect 2190 19875 2195 19905
rect 2195 19875 2225 19905
rect 2225 19875 2230 19905
rect 2190 19870 2230 19875
rect 2190 19835 2230 19840
rect 2190 19805 2195 19835
rect 2195 19805 2225 19835
rect 2225 19805 2230 19835
rect 2190 19800 2230 19805
rect 2190 19770 2230 19775
rect 2190 19740 2195 19770
rect 2195 19740 2225 19770
rect 2225 19740 2230 19770
rect 2190 19735 2230 19740
rect 2190 19710 2230 19715
rect 2190 19680 2195 19710
rect 2195 19680 2225 19710
rect 2225 19680 2230 19710
rect 2190 19675 2230 19680
rect 2190 19645 2230 19650
rect 2190 19615 2195 19645
rect 2195 19615 2225 19645
rect 2225 19615 2230 19645
rect 2190 19610 2230 19615
rect 2190 19575 2230 19580
rect 2190 19545 2195 19575
rect 2195 19545 2225 19575
rect 2225 19545 2230 19575
rect 2190 19540 2230 19545
rect 2190 19505 2230 19510
rect 2190 19475 2195 19505
rect 2195 19475 2225 19505
rect 2225 19475 2230 19505
rect 2190 19470 2230 19475
rect 2190 19435 2230 19440
rect 2190 19405 2195 19435
rect 2195 19405 2225 19435
rect 2225 19405 2230 19435
rect 2190 19400 2230 19405
rect 2190 19370 2230 19375
rect 2190 19340 2195 19370
rect 2195 19340 2225 19370
rect 2225 19340 2230 19370
rect 2190 19335 2230 19340
rect 2190 19310 2230 19315
rect 2190 19280 2195 19310
rect 2195 19280 2225 19310
rect 2225 19280 2230 19310
rect 2190 19275 2230 19280
rect 2190 19245 2230 19250
rect 2190 19215 2195 19245
rect 2195 19215 2225 19245
rect 2225 19215 2230 19245
rect 2190 19210 2230 19215
rect 2190 19175 2230 19180
rect 2190 19145 2195 19175
rect 2195 19145 2225 19175
rect 2225 19145 2230 19175
rect 2190 19140 2230 19145
rect 2190 19105 2230 19110
rect 2190 19075 2195 19105
rect 2195 19075 2225 19105
rect 2225 19075 2230 19105
rect 2190 19070 2230 19075
rect 2190 19035 2230 19040
rect 2190 19005 2195 19035
rect 2195 19005 2225 19035
rect 2225 19005 2230 19035
rect 2190 19000 2230 19005
rect 2190 18970 2230 18975
rect 2190 18940 2195 18970
rect 2195 18940 2225 18970
rect 2225 18940 2230 18970
rect 2190 18935 2230 18940
rect 2190 18910 2230 18915
rect 2190 18880 2195 18910
rect 2195 18880 2225 18910
rect 2225 18880 2230 18910
rect 2190 18875 2230 18880
rect 2190 18845 2230 18850
rect 2190 18815 2195 18845
rect 2195 18815 2225 18845
rect 2225 18815 2230 18845
rect 2190 18810 2230 18815
rect 2190 18775 2230 18780
rect 2190 18745 2195 18775
rect 2195 18745 2225 18775
rect 2225 18745 2230 18775
rect 2190 18740 2230 18745
rect 2190 18705 2230 18710
rect 2190 18675 2195 18705
rect 2195 18675 2225 18705
rect 2225 18675 2230 18705
rect 2190 18670 2230 18675
rect 2190 18635 2230 18640
rect 2190 18605 2195 18635
rect 2195 18605 2225 18635
rect 2225 18605 2230 18635
rect 2190 18600 2230 18605
rect 2190 18570 2230 18575
rect 2190 18540 2195 18570
rect 2195 18540 2225 18570
rect 2225 18540 2230 18570
rect 2190 18535 2230 18540
rect 2190 18510 2230 18515
rect 2190 18480 2195 18510
rect 2195 18480 2225 18510
rect 2225 18480 2230 18510
rect 2190 18475 2230 18480
rect 2190 18445 2230 18450
rect 2190 18415 2195 18445
rect 2195 18415 2225 18445
rect 2225 18415 2230 18445
rect 2190 18410 2230 18415
rect 2190 18375 2230 18380
rect 2190 18345 2195 18375
rect 2195 18345 2225 18375
rect 2225 18345 2230 18375
rect 2190 18340 2230 18345
rect 2190 18305 2230 18310
rect 2190 18275 2195 18305
rect 2195 18275 2225 18305
rect 2225 18275 2230 18305
rect 2190 18270 2230 18275
rect 2190 18235 2230 18240
rect 2190 18205 2195 18235
rect 2195 18205 2225 18235
rect 2225 18205 2230 18235
rect 2190 18200 2230 18205
rect 2190 18170 2230 18175
rect 2190 18140 2195 18170
rect 2195 18140 2225 18170
rect 2225 18140 2230 18170
rect 2190 18135 2230 18140
rect 2190 18110 2230 18115
rect 2190 18080 2195 18110
rect 2195 18080 2225 18110
rect 2225 18080 2230 18110
rect 2190 18075 2230 18080
rect 2190 18045 2230 18050
rect 2190 18015 2195 18045
rect 2195 18015 2225 18045
rect 2225 18015 2230 18045
rect 2190 18010 2230 18015
rect 2190 17975 2230 17980
rect 2190 17945 2195 17975
rect 2195 17945 2225 17975
rect 2225 17945 2230 17975
rect 2190 17940 2230 17945
rect 2190 17905 2230 17910
rect 2190 17875 2195 17905
rect 2195 17875 2225 17905
rect 2225 17875 2230 17905
rect 2190 17870 2230 17875
rect 2190 17835 2230 17840
rect 2190 17805 2195 17835
rect 2195 17805 2225 17835
rect 2225 17805 2230 17835
rect 2190 17800 2230 17805
rect 2190 17770 2230 17775
rect 2190 17740 2195 17770
rect 2195 17740 2225 17770
rect 2225 17740 2230 17770
rect 2190 17735 2230 17740
rect 6660 20910 6700 20915
rect 6660 20880 6665 20910
rect 6665 20880 6695 20910
rect 6695 20880 6700 20910
rect 6660 20875 6700 20880
rect 6660 20845 6700 20850
rect 6660 20815 6665 20845
rect 6665 20815 6695 20845
rect 6695 20815 6700 20845
rect 6660 20810 6700 20815
rect 6660 20775 6700 20780
rect 6660 20745 6665 20775
rect 6665 20745 6695 20775
rect 6695 20745 6700 20775
rect 6660 20740 6700 20745
rect 6660 20705 6700 20710
rect 6660 20675 6665 20705
rect 6665 20675 6695 20705
rect 6695 20675 6700 20705
rect 6660 20670 6700 20675
rect 6660 20635 6700 20640
rect 6660 20605 6665 20635
rect 6665 20605 6695 20635
rect 6695 20605 6700 20635
rect 6660 20600 6700 20605
rect 6660 20570 6700 20575
rect 6660 20540 6665 20570
rect 6665 20540 6695 20570
rect 6695 20540 6700 20570
rect 6660 20535 6700 20540
rect 6660 20510 6700 20515
rect 6660 20480 6665 20510
rect 6665 20480 6695 20510
rect 6695 20480 6700 20510
rect 6660 20475 6700 20480
rect 6660 20445 6700 20450
rect 6660 20415 6665 20445
rect 6665 20415 6695 20445
rect 6695 20415 6700 20445
rect 6660 20410 6700 20415
rect 6660 20375 6700 20380
rect 6660 20345 6665 20375
rect 6665 20345 6695 20375
rect 6695 20345 6700 20375
rect 6660 20340 6700 20345
rect 6660 20305 6700 20310
rect 6660 20275 6665 20305
rect 6665 20275 6695 20305
rect 6695 20275 6700 20305
rect 6660 20270 6700 20275
rect 6660 20235 6700 20240
rect 6660 20205 6665 20235
rect 6665 20205 6695 20235
rect 6695 20205 6700 20235
rect 6660 20200 6700 20205
rect 6660 20170 6700 20175
rect 6660 20140 6665 20170
rect 6665 20140 6695 20170
rect 6695 20140 6700 20170
rect 6660 20135 6700 20140
rect 6660 20110 6700 20115
rect 6660 20080 6665 20110
rect 6665 20080 6695 20110
rect 6695 20080 6700 20110
rect 6660 20075 6700 20080
rect 6660 20045 6700 20050
rect 6660 20015 6665 20045
rect 6665 20015 6695 20045
rect 6695 20015 6700 20045
rect 6660 20010 6700 20015
rect 6660 19975 6700 19980
rect 6660 19945 6665 19975
rect 6665 19945 6695 19975
rect 6695 19945 6700 19975
rect 6660 19940 6700 19945
rect 6660 19905 6700 19910
rect 6660 19875 6665 19905
rect 6665 19875 6695 19905
rect 6695 19875 6700 19905
rect 6660 19870 6700 19875
rect 6660 19835 6700 19840
rect 6660 19805 6665 19835
rect 6665 19805 6695 19835
rect 6695 19805 6700 19835
rect 6660 19800 6700 19805
rect 6660 19770 6700 19775
rect 6660 19740 6665 19770
rect 6665 19740 6695 19770
rect 6695 19740 6700 19770
rect 6660 19735 6700 19740
rect 6660 19710 6700 19715
rect 6660 19680 6665 19710
rect 6665 19680 6695 19710
rect 6695 19680 6700 19710
rect 6660 19675 6700 19680
rect 6660 19645 6700 19650
rect 6660 19615 6665 19645
rect 6665 19615 6695 19645
rect 6695 19615 6700 19645
rect 6660 19610 6700 19615
rect 6660 19575 6700 19580
rect 6660 19545 6665 19575
rect 6665 19545 6695 19575
rect 6695 19545 6700 19575
rect 6660 19540 6700 19545
rect 6660 19505 6700 19510
rect 6660 19475 6665 19505
rect 6665 19475 6695 19505
rect 6695 19475 6700 19505
rect 6660 19470 6700 19475
rect 6660 19435 6700 19440
rect 6660 19405 6665 19435
rect 6665 19405 6695 19435
rect 6695 19405 6700 19435
rect 6660 19400 6700 19405
rect 6660 19370 6700 19375
rect 6660 19340 6665 19370
rect 6665 19340 6695 19370
rect 6695 19340 6700 19370
rect 6660 19335 6700 19340
rect 6660 19310 6700 19315
rect 6660 19280 6665 19310
rect 6665 19280 6695 19310
rect 6695 19280 6700 19310
rect 6660 19275 6700 19280
rect 6660 19245 6700 19250
rect 6660 19215 6665 19245
rect 6665 19215 6695 19245
rect 6695 19215 6700 19245
rect 6660 19210 6700 19215
rect 6660 19175 6700 19180
rect 6660 19145 6665 19175
rect 6665 19145 6695 19175
rect 6695 19145 6700 19175
rect 6660 19140 6700 19145
rect 6660 19105 6700 19110
rect 6660 19075 6665 19105
rect 6665 19075 6695 19105
rect 6695 19075 6700 19105
rect 6660 19070 6700 19075
rect 6660 19035 6700 19040
rect 6660 19005 6665 19035
rect 6665 19005 6695 19035
rect 6695 19005 6700 19035
rect 6660 19000 6700 19005
rect 6660 18970 6700 18975
rect 6660 18940 6665 18970
rect 6665 18940 6695 18970
rect 6695 18940 6700 18970
rect 6660 18935 6700 18940
rect 6660 18910 6700 18915
rect 6660 18880 6665 18910
rect 6665 18880 6695 18910
rect 6695 18880 6700 18910
rect 6660 18875 6700 18880
rect 6660 18845 6700 18850
rect 6660 18815 6665 18845
rect 6665 18815 6695 18845
rect 6695 18815 6700 18845
rect 6660 18810 6700 18815
rect 6660 18775 6700 18780
rect 6660 18745 6665 18775
rect 6665 18745 6695 18775
rect 6695 18745 6700 18775
rect 6660 18740 6700 18745
rect 6660 18705 6700 18710
rect 6660 18675 6665 18705
rect 6665 18675 6695 18705
rect 6695 18675 6700 18705
rect 6660 18670 6700 18675
rect 6660 18635 6700 18640
rect 6660 18605 6665 18635
rect 6665 18605 6695 18635
rect 6695 18605 6700 18635
rect 6660 18600 6700 18605
rect 6660 18570 6700 18575
rect 6660 18540 6665 18570
rect 6665 18540 6695 18570
rect 6695 18540 6700 18570
rect 6660 18535 6700 18540
rect 6660 18510 6700 18515
rect 6660 18480 6665 18510
rect 6665 18480 6695 18510
rect 6695 18480 6700 18510
rect 6660 18475 6700 18480
rect 6660 18445 6700 18450
rect 6660 18415 6665 18445
rect 6665 18415 6695 18445
rect 6695 18415 6700 18445
rect 6660 18410 6700 18415
rect 6660 18375 6700 18380
rect 6660 18345 6665 18375
rect 6665 18345 6695 18375
rect 6695 18345 6700 18375
rect 6660 18340 6700 18345
rect 6660 18305 6700 18310
rect 6660 18275 6665 18305
rect 6665 18275 6695 18305
rect 6695 18275 6700 18305
rect 6660 18270 6700 18275
rect 6660 18235 6700 18240
rect 6660 18205 6665 18235
rect 6665 18205 6695 18235
rect 6695 18205 6700 18235
rect 6660 18200 6700 18205
rect 6660 18170 6700 18175
rect 6660 18140 6665 18170
rect 6665 18140 6695 18170
rect 6695 18140 6700 18170
rect 6660 18135 6700 18140
rect 6660 18110 6700 18115
rect 6660 18080 6665 18110
rect 6665 18080 6695 18110
rect 6695 18080 6700 18110
rect 6660 18075 6700 18080
rect 6660 18045 6700 18050
rect 6660 18015 6665 18045
rect 6665 18015 6695 18045
rect 6695 18015 6700 18045
rect 6660 18010 6700 18015
rect 6660 17975 6700 17980
rect 6660 17945 6665 17975
rect 6665 17945 6695 17975
rect 6695 17945 6700 17975
rect 6660 17940 6700 17945
rect 6660 17905 6700 17910
rect 6660 17875 6665 17905
rect 6665 17875 6695 17905
rect 6695 17875 6700 17905
rect 6660 17870 6700 17875
rect 6660 17835 6700 17840
rect 6660 17805 6665 17835
rect 6665 17805 6695 17835
rect 6695 17805 6700 17835
rect 6660 17800 6700 17805
rect 6660 17770 6700 17775
rect 6660 17740 6665 17770
rect 6665 17740 6695 17770
rect 6695 17740 6700 17770
rect 6660 17735 6700 17740
rect 12925 20840 12975 20890
rect 13020 20840 13070 20890
rect 13115 20840 13165 20890
rect 13215 20840 13265 20890
rect 13315 20840 13365 20890
rect 13415 20840 13465 20890
rect 13510 20840 13560 20890
rect 13605 20840 13655 20890
rect 13725 20840 13775 20890
rect 13820 20840 13870 20890
rect 13915 20840 13965 20890
rect 14015 20840 14065 20890
rect 14115 20840 14165 20890
rect 14215 20840 14265 20890
rect 14310 20840 14360 20890
rect 14405 20840 14455 20890
rect 14525 20840 14575 20890
rect 14620 20840 14670 20890
rect 14715 20840 14765 20890
rect 14815 20840 14865 20890
rect 14915 20840 14965 20890
rect 15015 20840 15065 20890
rect 15110 20840 15160 20890
rect 15205 20840 15255 20890
rect 15325 20840 15375 20890
rect 15420 20840 15470 20890
rect 15515 20840 15565 20890
rect 15615 20840 15665 20890
rect 15715 20840 15765 20890
rect 15815 20840 15865 20890
rect 15910 20840 15960 20890
rect 16005 20840 16055 20890
rect 12925 20750 12975 20800
rect 13020 20750 13070 20800
rect 13115 20750 13165 20800
rect 13215 20750 13265 20800
rect 13315 20750 13365 20800
rect 13415 20750 13465 20800
rect 13510 20750 13560 20800
rect 13605 20750 13655 20800
rect 13725 20750 13775 20800
rect 13820 20750 13870 20800
rect 13915 20750 13965 20800
rect 14015 20750 14065 20800
rect 14115 20750 14165 20800
rect 14215 20750 14265 20800
rect 14310 20750 14360 20800
rect 14405 20750 14455 20800
rect 14525 20750 14575 20800
rect 14620 20750 14670 20800
rect 14715 20750 14765 20800
rect 14815 20750 14865 20800
rect 14915 20750 14965 20800
rect 15015 20750 15065 20800
rect 15110 20750 15160 20800
rect 15205 20750 15255 20800
rect 15325 20750 15375 20800
rect 15420 20750 15470 20800
rect 15515 20750 15565 20800
rect 15615 20750 15665 20800
rect 15715 20750 15765 20800
rect 15815 20750 15865 20800
rect 15910 20750 15960 20800
rect 16005 20750 16055 20800
rect 12925 20650 12975 20700
rect 13020 20650 13070 20700
rect 13115 20650 13165 20700
rect 13215 20650 13265 20700
rect 13315 20650 13365 20700
rect 13415 20650 13465 20700
rect 13510 20650 13560 20700
rect 13605 20650 13655 20700
rect 13725 20650 13775 20700
rect 13820 20650 13870 20700
rect 13915 20650 13965 20700
rect 14015 20650 14065 20700
rect 14115 20650 14165 20700
rect 14215 20650 14265 20700
rect 14310 20650 14360 20700
rect 14405 20650 14455 20700
rect 14525 20650 14575 20700
rect 14620 20650 14670 20700
rect 14715 20650 14765 20700
rect 14815 20650 14865 20700
rect 14915 20650 14965 20700
rect 15015 20650 15065 20700
rect 15110 20650 15160 20700
rect 15205 20650 15255 20700
rect 15325 20650 15375 20700
rect 15420 20650 15470 20700
rect 15515 20650 15565 20700
rect 15615 20650 15665 20700
rect 15715 20650 15765 20700
rect 15815 20650 15865 20700
rect 15910 20650 15960 20700
rect 16005 20650 16055 20700
rect 12925 20560 12975 20610
rect 13020 20560 13070 20610
rect 13115 20560 13165 20610
rect 13215 20560 13265 20610
rect 13315 20560 13365 20610
rect 13415 20560 13465 20610
rect 13510 20560 13560 20610
rect 13605 20560 13655 20610
rect 13725 20560 13775 20610
rect 13820 20560 13870 20610
rect 13915 20560 13965 20610
rect 14015 20560 14065 20610
rect 14115 20560 14165 20610
rect 14215 20560 14265 20610
rect 14310 20560 14360 20610
rect 14405 20560 14455 20610
rect 14525 20560 14575 20610
rect 14620 20560 14670 20610
rect 14715 20560 14765 20610
rect 14815 20560 14865 20610
rect 14915 20560 14965 20610
rect 15015 20560 15065 20610
rect 15110 20560 15160 20610
rect 15205 20560 15255 20610
rect 15325 20560 15375 20610
rect 15420 20560 15470 20610
rect 15515 20560 15565 20610
rect 15615 20560 15665 20610
rect 15715 20560 15765 20610
rect 15815 20560 15865 20610
rect 15910 20560 15960 20610
rect 16005 20560 16055 20610
rect 12925 20440 12975 20490
rect 13020 20440 13070 20490
rect 13115 20440 13165 20490
rect 13215 20440 13265 20490
rect 13315 20440 13365 20490
rect 13415 20440 13465 20490
rect 13510 20440 13560 20490
rect 13605 20440 13655 20490
rect 13725 20440 13775 20490
rect 13820 20440 13870 20490
rect 13915 20440 13965 20490
rect 14015 20440 14065 20490
rect 14115 20440 14165 20490
rect 14215 20440 14265 20490
rect 14310 20440 14360 20490
rect 14405 20440 14455 20490
rect 14525 20440 14575 20490
rect 14620 20440 14670 20490
rect 14715 20440 14765 20490
rect 14815 20440 14865 20490
rect 14915 20440 14965 20490
rect 15015 20440 15065 20490
rect 15110 20440 15160 20490
rect 15205 20440 15255 20490
rect 15325 20440 15375 20490
rect 15420 20440 15470 20490
rect 15515 20440 15565 20490
rect 15615 20440 15665 20490
rect 15715 20440 15765 20490
rect 15815 20440 15865 20490
rect 15910 20440 15960 20490
rect 16005 20440 16055 20490
rect 12925 20350 12975 20400
rect 13020 20350 13070 20400
rect 13115 20350 13165 20400
rect 13215 20350 13265 20400
rect 13315 20350 13365 20400
rect 13415 20350 13465 20400
rect 13510 20350 13560 20400
rect 13605 20350 13655 20400
rect 13725 20350 13775 20400
rect 13820 20350 13870 20400
rect 13915 20350 13965 20400
rect 14015 20350 14065 20400
rect 14115 20350 14165 20400
rect 14215 20350 14265 20400
rect 14310 20350 14360 20400
rect 14405 20350 14455 20400
rect 14525 20350 14575 20400
rect 14620 20350 14670 20400
rect 14715 20350 14765 20400
rect 14815 20350 14865 20400
rect 14915 20350 14965 20400
rect 15015 20350 15065 20400
rect 15110 20350 15160 20400
rect 15205 20350 15255 20400
rect 15325 20350 15375 20400
rect 15420 20350 15470 20400
rect 15515 20350 15565 20400
rect 15615 20350 15665 20400
rect 15715 20350 15765 20400
rect 15815 20350 15865 20400
rect 15910 20350 15960 20400
rect 16005 20350 16055 20400
rect 12925 20250 12975 20300
rect 13020 20250 13070 20300
rect 13115 20250 13165 20300
rect 13215 20250 13265 20300
rect 13315 20250 13365 20300
rect 13415 20250 13465 20300
rect 13510 20250 13560 20300
rect 13605 20250 13655 20300
rect 13725 20250 13775 20300
rect 13820 20250 13870 20300
rect 13915 20250 13965 20300
rect 14015 20250 14065 20300
rect 14115 20250 14165 20300
rect 14215 20250 14265 20300
rect 14310 20250 14360 20300
rect 14405 20250 14455 20300
rect 14525 20250 14575 20300
rect 14620 20250 14670 20300
rect 14715 20250 14765 20300
rect 14815 20250 14865 20300
rect 14915 20250 14965 20300
rect 15015 20250 15065 20300
rect 15110 20250 15160 20300
rect 15205 20250 15255 20300
rect 15325 20250 15375 20300
rect 15420 20250 15470 20300
rect 15515 20250 15565 20300
rect 15615 20250 15665 20300
rect 15715 20250 15765 20300
rect 15815 20250 15865 20300
rect 15910 20250 15960 20300
rect 16005 20250 16055 20300
rect 12925 20160 12975 20210
rect 13020 20160 13070 20210
rect 13115 20160 13165 20210
rect 13215 20160 13265 20210
rect 13315 20160 13365 20210
rect 13415 20160 13465 20210
rect 13510 20160 13560 20210
rect 13605 20160 13655 20210
rect 13725 20160 13775 20210
rect 13820 20160 13870 20210
rect 13915 20160 13965 20210
rect 14015 20160 14065 20210
rect 14115 20160 14165 20210
rect 14215 20160 14265 20210
rect 14310 20160 14360 20210
rect 14405 20160 14455 20210
rect 14525 20160 14575 20210
rect 14620 20160 14670 20210
rect 14715 20160 14765 20210
rect 14815 20160 14865 20210
rect 14915 20160 14965 20210
rect 15015 20160 15065 20210
rect 15110 20160 15160 20210
rect 15205 20160 15255 20210
rect 15325 20160 15375 20210
rect 15420 20160 15470 20210
rect 15515 20160 15565 20210
rect 15615 20160 15665 20210
rect 15715 20160 15765 20210
rect 15815 20160 15865 20210
rect 15910 20160 15960 20210
rect 16005 20160 16055 20210
rect 12925 20040 12975 20090
rect 13020 20040 13070 20090
rect 13115 20040 13165 20090
rect 13215 20040 13265 20090
rect 13315 20040 13365 20090
rect 13415 20040 13465 20090
rect 13510 20040 13560 20090
rect 13605 20040 13655 20090
rect 13725 20040 13775 20090
rect 13820 20040 13870 20090
rect 13915 20040 13965 20090
rect 14015 20040 14065 20090
rect 14115 20040 14165 20090
rect 14215 20040 14265 20090
rect 14310 20040 14360 20090
rect 14405 20040 14455 20090
rect 14525 20040 14575 20090
rect 14620 20040 14670 20090
rect 14715 20040 14765 20090
rect 14815 20040 14865 20090
rect 14915 20040 14965 20090
rect 15015 20040 15065 20090
rect 15110 20040 15160 20090
rect 15205 20040 15255 20090
rect 15325 20040 15375 20090
rect 15420 20040 15470 20090
rect 15515 20040 15565 20090
rect 15615 20040 15665 20090
rect 15715 20040 15765 20090
rect 15815 20040 15865 20090
rect 15910 20040 15960 20090
rect 16005 20040 16055 20090
rect 12925 19950 12975 20000
rect 13020 19950 13070 20000
rect 13115 19950 13165 20000
rect 13215 19950 13265 20000
rect 13315 19950 13365 20000
rect 13415 19950 13465 20000
rect 13510 19950 13560 20000
rect 13605 19950 13655 20000
rect 13725 19950 13775 20000
rect 13820 19950 13870 20000
rect 13915 19950 13965 20000
rect 14015 19950 14065 20000
rect 14115 19950 14165 20000
rect 14215 19950 14265 20000
rect 14310 19950 14360 20000
rect 14405 19950 14455 20000
rect 14525 19950 14575 20000
rect 14620 19950 14670 20000
rect 14715 19950 14765 20000
rect 14815 19950 14865 20000
rect 14915 19950 14965 20000
rect 15015 19950 15065 20000
rect 15110 19950 15160 20000
rect 15205 19950 15255 20000
rect 15325 19950 15375 20000
rect 15420 19950 15470 20000
rect 15515 19950 15565 20000
rect 15615 19950 15665 20000
rect 15715 19950 15765 20000
rect 15815 19950 15865 20000
rect 15910 19950 15960 20000
rect 16005 19950 16055 20000
rect 12925 19850 12975 19900
rect 13020 19850 13070 19900
rect 13115 19850 13165 19900
rect 13215 19850 13265 19900
rect 13315 19850 13365 19900
rect 13415 19850 13465 19900
rect 13510 19850 13560 19900
rect 13605 19850 13655 19900
rect 13725 19850 13775 19900
rect 13820 19850 13870 19900
rect 13915 19850 13965 19900
rect 14015 19850 14065 19900
rect 14115 19850 14165 19900
rect 14215 19850 14265 19900
rect 14310 19850 14360 19900
rect 14405 19850 14455 19900
rect 14525 19850 14575 19900
rect 14620 19850 14670 19900
rect 14715 19850 14765 19900
rect 14815 19850 14865 19900
rect 14915 19850 14965 19900
rect 15015 19850 15065 19900
rect 15110 19850 15160 19900
rect 15205 19850 15255 19900
rect 15325 19850 15375 19900
rect 15420 19850 15470 19900
rect 15515 19850 15565 19900
rect 15615 19850 15665 19900
rect 15715 19850 15765 19900
rect 15815 19850 15865 19900
rect 15910 19850 15960 19900
rect 16005 19850 16055 19900
rect 12925 19760 12975 19810
rect 13020 19760 13070 19810
rect 13115 19760 13165 19810
rect 13215 19760 13265 19810
rect 13315 19760 13365 19810
rect 13415 19760 13465 19810
rect 13510 19760 13560 19810
rect 13605 19760 13655 19810
rect 13725 19760 13775 19810
rect 13820 19760 13870 19810
rect 13915 19760 13965 19810
rect 14015 19760 14065 19810
rect 14115 19760 14165 19810
rect 14215 19760 14265 19810
rect 14310 19760 14360 19810
rect 14405 19760 14455 19810
rect 14525 19760 14575 19810
rect 14620 19760 14670 19810
rect 14715 19760 14765 19810
rect 14815 19760 14865 19810
rect 14915 19760 14965 19810
rect 15015 19760 15065 19810
rect 15110 19760 15160 19810
rect 15205 19760 15255 19810
rect 15325 19760 15375 19810
rect 15420 19760 15470 19810
rect 15515 19760 15565 19810
rect 15615 19760 15665 19810
rect 15715 19760 15765 19810
rect 15815 19760 15865 19810
rect 15910 19760 15960 19810
rect 16005 19760 16055 19810
rect 12925 19640 12975 19690
rect 13020 19640 13070 19690
rect 13115 19640 13165 19690
rect 13215 19640 13265 19690
rect 13315 19640 13365 19690
rect 13415 19640 13465 19690
rect 13510 19640 13560 19690
rect 13605 19640 13655 19690
rect 13725 19640 13775 19690
rect 13820 19640 13870 19690
rect 13915 19640 13965 19690
rect 14015 19640 14065 19690
rect 14115 19640 14165 19690
rect 14215 19640 14265 19690
rect 14310 19640 14360 19690
rect 14405 19640 14455 19690
rect 14525 19640 14575 19690
rect 14620 19640 14670 19690
rect 14715 19640 14765 19690
rect 14815 19640 14865 19690
rect 14915 19640 14965 19690
rect 15015 19640 15065 19690
rect 15110 19640 15160 19690
rect 15205 19640 15255 19690
rect 15325 19640 15375 19690
rect 15420 19640 15470 19690
rect 15515 19640 15565 19690
rect 15615 19640 15665 19690
rect 15715 19640 15765 19690
rect 15815 19640 15865 19690
rect 15910 19640 15960 19690
rect 16005 19640 16055 19690
rect 12925 19550 12975 19600
rect 13020 19550 13070 19600
rect 13115 19550 13165 19600
rect 13215 19550 13265 19600
rect 13315 19550 13365 19600
rect 13415 19550 13465 19600
rect 13510 19550 13560 19600
rect 13605 19550 13655 19600
rect 13725 19550 13775 19600
rect 13820 19550 13870 19600
rect 13915 19550 13965 19600
rect 14015 19550 14065 19600
rect 14115 19550 14165 19600
rect 14215 19550 14265 19600
rect 14310 19550 14360 19600
rect 14405 19550 14455 19600
rect 14525 19550 14575 19600
rect 14620 19550 14670 19600
rect 14715 19550 14765 19600
rect 14815 19550 14865 19600
rect 14915 19550 14965 19600
rect 15015 19550 15065 19600
rect 15110 19550 15160 19600
rect 15205 19550 15255 19600
rect 15325 19550 15375 19600
rect 15420 19550 15470 19600
rect 15515 19550 15565 19600
rect 15615 19550 15665 19600
rect 15715 19550 15765 19600
rect 15815 19550 15865 19600
rect 15910 19550 15960 19600
rect 16005 19550 16055 19600
rect 12925 19450 12975 19500
rect 13020 19450 13070 19500
rect 13115 19450 13165 19500
rect 13215 19450 13265 19500
rect 13315 19450 13365 19500
rect 13415 19450 13465 19500
rect 13510 19450 13560 19500
rect 13605 19450 13655 19500
rect 13725 19450 13775 19500
rect 13820 19450 13870 19500
rect 13915 19450 13965 19500
rect 14015 19450 14065 19500
rect 14115 19450 14165 19500
rect 14215 19450 14265 19500
rect 14310 19450 14360 19500
rect 14405 19450 14455 19500
rect 14525 19450 14575 19500
rect 14620 19450 14670 19500
rect 14715 19450 14765 19500
rect 14815 19450 14865 19500
rect 14915 19450 14965 19500
rect 15015 19450 15065 19500
rect 15110 19450 15160 19500
rect 15205 19450 15255 19500
rect 15325 19450 15375 19500
rect 15420 19450 15470 19500
rect 15515 19450 15565 19500
rect 15615 19450 15665 19500
rect 15715 19450 15765 19500
rect 15815 19450 15865 19500
rect 15910 19450 15960 19500
rect 16005 19450 16055 19500
rect 12925 19360 12975 19410
rect 13020 19360 13070 19410
rect 13115 19360 13165 19410
rect 13215 19360 13265 19410
rect 13315 19360 13365 19410
rect 13415 19360 13465 19410
rect 13510 19360 13560 19410
rect 13605 19360 13655 19410
rect 13725 19360 13775 19410
rect 13820 19360 13870 19410
rect 13915 19360 13965 19410
rect 14015 19360 14065 19410
rect 14115 19360 14165 19410
rect 14215 19360 14265 19410
rect 14310 19360 14360 19410
rect 14405 19360 14455 19410
rect 14525 19360 14575 19410
rect 14620 19360 14670 19410
rect 14715 19360 14765 19410
rect 14815 19360 14865 19410
rect 14915 19360 14965 19410
rect 15015 19360 15065 19410
rect 15110 19360 15160 19410
rect 15205 19360 15255 19410
rect 15325 19360 15375 19410
rect 15420 19360 15470 19410
rect 15515 19360 15565 19410
rect 15615 19360 15665 19410
rect 15715 19360 15765 19410
rect 15815 19360 15865 19410
rect 15910 19360 15960 19410
rect 16005 19360 16055 19410
rect 12925 19240 12975 19290
rect 13020 19240 13070 19290
rect 13115 19240 13165 19290
rect 13215 19240 13265 19290
rect 13315 19240 13365 19290
rect 13415 19240 13465 19290
rect 13510 19240 13560 19290
rect 13605 19240 13655 19290
rect 13725 19240 13775 19290
rect 13820 19240 13870 19290
rect 13915 19240 13965 19290
rect 14015 19240 14065 19290
rect 14115 19240 14165 19290
rect 14215 19240 14265 19290
rect 14310 19240 14360 19290
rect 14405 19240 14455 19290
rect 14525 19240 14575 19290
rect 14620 19240 14670 19290
rect 14715 19240 14765 19290
rect 14815 19240 14865 19290
rect 14915 19240 14965 19290
rect 15015 19240 15065 19290
rect 15110 19240 15160 19290
rect 15205 19240 15255 19290
rect 15325 19240 15375 19290
rect 15420 19240 15470 19290
rect 15515 19240 15565 19290
rect 15615 19240 15665 19290
rect 15715 19240 15765 19290
rect 15815 19240 15865 19290
rect 15910 19240 15960 19290
rect 16005 19240 16055 19290
rect 12925 19150 12975 19200
rect 13020 19150 13070 19200
rect 13115 19150 13165 19200
rect 13215 19150 13265 19200
rect 13315 19150 13365 19200
rect 13415 19150 13465 19200
rect 13510 19150 13560 19200
rect 13605 19150 13655 19200
rect 13725 19150 13775 19200
rect 13820 19150 13870 19200
rect 13915 19150 13965 19200
rect 14015 19150 14065 19200
rect 14115 19150 14165 19200
rect 14215 19150 14265 19200
rect 14310 19150 14360 19200
rect 14405 19150 14455 19200
rect 14525 19150 14575 19200
rect 14620 19150 14670 19200
rect 14715 19150 14765 19200
rect 14815 19150 14865 19200
rect 14915 19150 14965 19200
rect 15015 19150 15065 19200
rect 15110 19150 15160 19200
rect 15205 19150 15255 19200
rect 15325 19150 15375 19200
rect 15420 19150 15470 19200
rect 15515 19150 15565 19200
rect 15615 19150 15665 19200
rect 15715 19150 15765 19200
rect 15815 19150 15865 19200
rect 15910 19150 15960 19200
rect 16005 19150 16055 19200
rect 12925 19050 12975 19100
rect 13020 19050 13070 19100
rect 13115 19050 13165 19100
rect 13215 19050 13265 19100
rect 13315 19050 13365 19100
rect 13415 19050 13465 19100
rect 13510 19050 13560 19100
rect 13605 19050 13655 19100
rect 13725 19050 13775 19100
rect 13820 19050 13870 19100
rect 13915 19050 13965 19100
rect 14015 19050 14065 19100
rect 14115 19050 14165 19100
rect 14215 19050 14265 19100
rect 14310 19050 14360 19100
rect 14405 19050 14455 19100
rect 14525 19050 14575 19100
rect 14620 19050 14670 19100
rect 14715 19050 14765 19100
rect 14815 19050 14865 19100
rect 14915 19050 14965 19100
rect 15015 19050 15065 19100
rect 15110 19050 15160 19100
rect 15205 19050 15255 19100
rect 15325 19050 15375 19100
rect 15420 19050 15470 19100
rect 15515 19050 15565 19100
rect 15615 19050 15665 19100
rect 15715 19050 15765 19100
rect 15815 19050 15865 19100
rect 15910 19050 15960 19100
rect 16005 19050 16055 19100
rect 12925 18960 12975 19010
rect 13020 18960 13070 19010
rect 13115 18960 13165 19010
rect 13215 18960 13265 19010
rect 13315 18960 13365 19010
rect 13415 18960 13465 19010
rect 13510 18960 13560 19010
rect 13605 18960 13655 19010
rect 13725 18960 13775 19010
rect 13820 18960 13870 19010
rect 13915 18960 13965 19010
rect 14015 18960 14065 19010
rect 14115 18960 14165 19010
rect 14215 18960 14265 19010
rect 14310 18960 14360 19010
rect 14405 18960 14455 19010
rect 14525 18960 14575 19010
rect 14620 18960 14670 19010
rect 14715 18960 14765 19010
rect 14815 18960 14865 19010
rect 14915 18960 14965 19010
rect 15015 18960 15065 19010
rect 15110 18960 15160 19010
rect 15205 18960 15255 19010
rect 15325 18960 15375 19010
rect 15420 18960 15470 19010
rect 15515 18960 15565 19010
rect 15615 18960 15665 19010
rect 15715 18960 15765 19010
rect 15815 18960 15865 19010
rect 15910 18960 15960 19010
rect 16005 18960 16055 19010
rect 12925 18840 12975 18890
rect 13020 18840 13070 18890
rect 13115 18840 13165 18890
rect 13215 18840 13265 18890
rect 13315 18840 13365 18890
rect 13415 18840 13465 18890
rect 13510 18840 13560 18890
rect 13605 18840 13655 18890
rect 13725 18840 13775 18890
rect 13820 18840 13870 18890
rect 13915 18840 13965 18890
rect 14015 18840 14065 18890
rect 14115 18840 14165 18890
rect 14215 18840 14265 18890
rect 14310 18840 14360 18890
rect 14405 18840 14455 18890
rect 14525 18840 14575 18890
rect 14620 18840 14670 18890
rect 14715 18840 14765 18890
rect 14815 18840 14865 18890
rect 14915 18840 14965 18890
rect 15015 18840 15065 18890
rect 15110 18840 15160 18890
rect 15205 18840 15255 18890
rect 15325 18840 15375 18890
rect 15420 18840 15470 18890
rect 15515 18840 15565 18890
rect 15615 18840 15665 18890
rect 15715 18840 15765 18890
rect 15815 18840 15865 18890
rect 15910 18840 15960 18890
rect 16005 18840 16055 18890
rect 12925 18750 12975 18800
rect 13020 18750 13070 18800
rect 13115 18750 13165 18800
rect 13215 18750 13265 18800
rect 13315 18750 13365 18800
rect 13415 18750 13465 18800
rect 13510 18750 13560 18800
rect 13605 18750 13655 18800
rect 13725 18750 13775 18800
rect 13820 18750 13870 18800
rect 13915 18750 13965 18800
rect 14015 18750 14065 18800
rect 14115 18750 14165 18800
rect 14215 18750 14265 18800
rect 14310 18750 14360 18800
rect 14405 18750 14455 18800
rect 14525 18750 14575 18800
rect 14620 18750 14670 18800
rect 14715 18750 14765 18800
rect 14815 18750 14865 18800
rect 14915 18750 14965 18800
rect 15015 18750 15065 18800
rect 15110 18750 15160 18800
rect 15205 18750 15255 18800
rect 15325 18750 15375 18800
rect 15420 18750 15470 18800
rect 15515 18750 15565 18800
rect 15615 18750 15665 18800
rect 15715 18750 15765 18800
rect 15815 18750 15865 18800
rect 15910 18750 15960 18800
rect 16005 18750 16055 18800
rect 12925 18650 12975 18700
rect 13020 18650 13070 18700
rect 13115 18650 13165 18700
rect 13215 18650 13265 18700
rect 13315 18650 13365 18700
rect 13415 18650 13465 18700
rect 13510 18650 13560 18700
rect 13605 18650 13655 18700
rect 13725 18650 13775 18700
rect 13820 18650 13870 18700
rect 13915 18650 13965 18700
rect 14015 18650 14065 18700
rect 14115 18650 14165 18700
rect 14215 18650 14265 18700
rect 14310 18650 14360 18700
rect 14405 18650 14455 18700
rect 14525 18650 14575 18700
rect 14620 18650 14670 18700
rect 14715 18650 14765 18700
rect 14815 18650 14865 18700
rect 14915 18650 14965 18700
rect 15015 18650 15065 18700
rect 15110 18650 15160 18700
rect 15205 18650 15255 18700
rect 15325 18650 15375 18700
rect 15420 18650 15470 18700
rect 15515 18650 15565 18700
rect 15615 18650 15665 18700
rect 15715 18650 15765 18700
rect 15815 18650 15865 18700
rect 15910 18650 15960 18700
rect 16005 18650 16055 18700
rect 12925 18560 12975 18610
rect 13020 18560 13070 18610
rect 13115 18560 13165 18610
rect 13215 18560 13265 18610
rect 13315 18560 13365 18610
rect 13415 18560 13465 18610
rect 13510 18560 13560 18610
rect 13605 18560 13655 18610
rect 13725 18560 13775 18610
rect 13820 18560 13870 18610
rect 13915 18560 13965 18610
rect 14015 18560 14065 18610
rect 14115 18560 14165 18610
rect 14215 18560 14265 18610
rect 14310 18560 14360 18610
rect 14405 18560 14455 18610
rect 14525 18560 14575 18610
rect 14620 18560 14670 18610
rect 14715 18560 14765 18610
rect 14815 18560 14865 18610
rect 14915 18560 14965 18610
rect 15015 18560 15065 18610
rect 15110 18560 15160 18610
rect 15205 18560 15255 18610
rect 15325 18560 15375 18610
rect 15420 18560 15470 18610
rect 15515 18560 15565 18610
rect 15615 18560 15665 18610
rect 15715 18560 15765 18610
rect 15815 18560 15865 18610
rect 15910 18560 15960 18610
rect 16005 18560 16055 18610
rect 12925 18440 12975 18490
rect 13020 18440 13070 18490
rect 13115 18440 13165 18490
rect 13215 18440 13265 18490
rect 13315 18440 13365 18490
rect 13415 18440 13465 18490
rect 13510 18440 13560 18490
rect 13605 18440 13655 18490
rect 13725 18440 13775 18490
rect 13820 18440 13870 18490
rect 13915 18440 13965 18490
rect 14015 18440 14065 18490
rect 14115 18440 14165 18490
rect 14215 18440 14265 18490
rect 14310 18440 14360 18490
rect 14405 18440 14455 18490
rect 14525 18440 14575 18490
rect 14620 18440 14670 18490
rect 14715 18440 14765 18490
rect 14815 18440 14865 18490
rect 14915 18440 14965 18490
rect 15015 18440 15065 18490
rect 15110 18440 15160 18490
rect 15205 18440 15255 18490
rect 15325 18440 15375 18490
rect 15420 18440 15470 18490
rect 15515 18440 15565 18490
rect 15615 18440 15665 18490
rect 15715 18440 15765 18490
rect 15815 18440 15865 18490
rect 15910 18440 15960 18490
rect 16005 18440 16055 18490
rect 12925 18350 12975 18400
rect 13020 18350 13070 18400
rect 13115 18350 13165 18400
rect 13215 18350 13265 18400
rect 13315 18350 13365 18400
rect 13415 18350 13465 18400
rect 13510 18350 13560 18400
rect 13605 18350 13655 18400
rect 13725 18350 13775 18400
rect 13820 18350 13870 18400
rect 13915 18350 13965 18400
rect 14015 18350 14065 18400
rect 14115 18350 14165 18400
rect 14215 18350 14265 18400
rect 14310 18350 14360 18400
rect 14405 18350 14455 18400
rect 14525 18350 14575 18400
rect 14620 18350 14670 18400
rect 14715 18350 14765 18400
rect 14815 18350 14865 18400
rect 14915 18350 14965 18400
rect 15015 18350 15065 18400
rect 15110 18350 15160 18400
rect 15205 18350 15255 18400
rect 15325 18350 15375 18400
rect 15420 18350 15470 18400
rect 15515 18350 15565 18400
rect 15615 18350 15665 18400
rect 15715 18350 15765 18400
rect 15815 18350 15865 18400
rect 15910 18350 15960 18400
rect 16005 18350 16055 18400
rect 12925 18250 12975 18300
rect 13020 18250 13070 18300
rect 13115 18250 13165 18300
rect 13215 18250 13265 18300
rect 13315 18250 13365 18300
rect 13415 18250 13465 18300
rect 13510 18250 13560 18300
rect 13605 18250 13655 18300
rect 13725 18250 13775 18300
rect 13820 18250 13870 18300
rect 13915 18250 13965 18300
rect 14015 18250 14065 18300
rect 14115 18250 14165 18300
rect 14215 18250 14265 18300
rect 14310 18250 14360 18300
rect 14405 18250 14455 18300
rect 14525 18250 14575 18300
rect 14620 18250 14670 18300
rect 14715 18250 14765 18300
rect 14815 18250 14865 18300
rect 14915 18250 14965 18300
rect 15015 18250 15065 18300
rect 15110 18250 15160 18300
rect 15205 18250 15255 18300
rect 15325 18250 15375 18300
rect 15420 18250 15470 18300
rect 15515 18250 15565 18300
rect 15615 18250 15665 18300
rect 15715 18250 15765 18300
rect 15815 18250 15865 18300
rect 15910 18250 15960 18300
rect 16005 18250 16055 18300
rect 12925 18160 12975 18210
rect 13020 18160 13070 18210
rect 13115 18160 13165 18210
rect 13215 18160 13265 18210
rect 13315 18160 13365 18210
rect 13415 18160 13465 18210
rect 13510 18160 13560 18210
rect 13605 18160 13655 18210
rect 13725 18160 13775 18210
rect 13820 18160 13870 18210
rect 13915 18160 13965 18210
rect 14015 18160 14065 18210
rect 14115 18160 14165 18210
rect 14215 18160 14265 18210
rect 14310 18160 14360 18210
rect 14405 18160 14455 18210
rect 14525 18160 14575 18210
rect 14620 18160 14670 18210
rect 14715 18160 14765 18210
rect 14815 18160 14865 18210
rect 14915 18160 14965 18210
rect 15015 18160 15065 18210
rect 15110 18160 15160 18210
rect 15205 18160 15255 18210
rect 15325 18160 15375 18210
rect 15420 18160 15470 18210
rect 15515 18160 15565 18210
rect 15615 18160 15665 18210
rect 15715 18160 15765 18210
rect 15815 18160 15865 18210
rect 15910 18160 15960 18210
rect 16005 18160 16055 18210
rect 12925 18040 12975 18090
rect 13020 18040 13070 18090
rect 13115 18040 13165 18090
rect 13215 18040 13265 18090
rect 13315 18040 13365 18090
rect 13415 18040 13465 18090
rect 13510 18040 13560 18090
rect 13605 18040 13655 18090
rect 13725 18040 13775 18090
rect 13820 18040 13870 18090
rect 13915 18040 13965 18090
rect 14015 18040 14065 18090
rect 14115 18040 14165 18090
rect 14215 18040 14265 18090
rect 14310 18040 14360 18090
rect 14405 18040 14455 18090
rect 14525 18040 14575 18090
rect 14620 18040 14670 18090
rect 14715 18040 14765 18090
rect 14815 18040 14865 18090
rect 14915 18040 14965 18090
rect 15015 18040 15065 18090
rect 15110 18040 15160 18090
rect 15205 18040 15255 18090
rect 15325 18040 15375 18090
rect 15420 18040 15470 18090
rect 15515 18040 15565 18090
rect 15615 18040 15665 18090
rect 15715 18040 15765 18090
rect 15815 18040 15865 18090
rect 15910 18040 15960 18090
rect 16005 18040 16055 18090
rect 12925 17950 12975 18000
rect 13020 17950 13070 18000
rect 13115 17950 13165 18000
rect 13215 17950 13265 18000
rect 13315 17950 13365 18000
rect 13415 17950 13465 18000
rect 13510 17950 13560 18000
rect 13605 17950 13655 18000
rect 13725 17950 13775 18000
rect 13820 17950 13870 18000
rect 13915 17950 13965 18000
rect 14015 17950 14065 18000
rect 14115 17950 14165 18000
rect 14215 17950 14265 18000
rect 14310 17950 14360 18000
rect 14405 17950 14455 18000
rect 14525 17950 14575 18000
rect 14620 17950 14670 18000
rect 14715 17950 14765 18000
rect 14815 17950 14865 18000
rect 14915 17950 14965 18000
rect 15015 17950 15065 18000
rect 15110 17950 15160 18000
rect 15205 17950 15255 18000
rect 15325 17950 15375 18000
rect 15420 17950 15470 18000
rect 15515 17950 15565 18000
rect 15615 17950 15665 18000
rect 15715 17950 15765 18000
rect 15815 17950 15865 18000
rect 15910 17950 15960 18000
rect 16005 17950 16055 18000
rect 12925 17850 12975 17900
rect 13020 17850 13070 17900
rect 13115 17850 13165 17900
rect 13215 17850 13265 17900
rect 13315 17850 13365 17900
rect 13415 17850 13465 17900
rect 13510 17850 13560 17900
rect 13605 17850 13655 17900
rect 13725 17850 13775 17900
rect 13820 17850 13870 17900
rect 13915 17850 13965 17900
rect 14015 17850 14065 17900
rect 14115 17850 14165 17900
rect 14215 17850 14265 17900
rect 14310 17850 14360 17900
rect 14405 17850 14455 17900
rect 14525 17850 14575 17900
rect 14620 17850 14670 17900
rect 14715 17850 14765 17900
rect 14815 17850 14865 17900
rect 14915 17850 14965 17900
rect 15015 17850 15065 17900
rect 15110 17850 15160 17900
rect 15205 17850 15255 17900
rect 15325 17850 15375 17900
rect 15420 17850 15470 17900
rect 15515 17850 15565 17900
rect 15615 17850 15665 17900
rect 15715 17850 15765 17900
rect 15815 17850 15865 17900
rect 15910 17850 15960 17900
rect 16005 17850 16055 17900
rect 12925 17760 12975 17810
rect 13020 17760 13070 17810
rect 13115 17760 13165 17810
rect 13215 17760 13265 17810
rect 13315 17760 13365 17810
rect 13415 17760 13465 17810
rect 13510 17760 13560 17810
rect 13605 17760 13655 17810
rect 13725 17760 13775 17810
rect 13820 17760 13870 17810
rect 13915 17760 13965 17810
rect 14015 17760 14065 17810
rect 14115 17760 14165 17810
rect 14215 17760 14265 17810
rect 14310 17760 14360 17810
rect 14405 17760 14455 17810
rect 14525 17760 14575 17810
rect 14620 17760 14670 17810
rect 14715 17760 14765 17810
rect 14815 17760 14865 17810
rect 14915 17760 14965 17810
rect 15015 17760 15065 17810
rect 15110 17760 15160 17810
rect 15205 17760 15255 17810
rect 15325 17760 15375 17810
rect 15420 17760 15470 17810
rect 15515 17760 15565 17810
rect 15615 17760 15665 17810
rect 15715 17760 15765 17810
rect 15815 17760 15865 17810
rect 15910 17760 15960 17810
rect 16005 17760 16055 17810
rect -4805 9565 -4755 9615
rect -4710 9565 -4660 9615
rect -4615 9565 -4565 9615
rect -4515 9565 -4465 9615
rect -4415 9565 -4365 9615
rect -4315 9565 -4265 9615
rect -4220 9565 -4170 9615
rect -4125 9565 -4075 9615
rect -4005 9565 -3955 9615
rect -3910 9565 -3860 9615
rect -3815 9565 -3765 9615
rect -3715 9565 -3665 9615
rect -3615 9565 -3565 9615
rect -3515 9565 -3465 9615
rect -3420 9565 -3370 9615
rect -3325 9565 -3275 9615
rect -3205 9565 -3155 9615
rect -3110 9565 -3060 9615
rect -3015 9565 -2965 9615
rect -2915 9565 -2865 9615
rect -2815 9565 -2765 9615
rect -2715 9565 -2665 9615
rect -2620 9565 -2570 9615
rect -2525 9565 -2475 9615
rect -2405 9565 -2355 9615
rect -2310 9565 -2260 9615
rect -2215 9565 -2165 9615
rect -2115 9565 -2065 9615
rect -2015 9565 -1965 9615
rect -1915 9565 -1865 9615
rect -1820 9565 -1770 9615
rect -1725 9565 -1675 9615
rect -4805 9475 -4755 9525
rect -4710 9475 -4660 9525
rect -4615 9475 -4565 9525
rect -4515 9475 -4465 9525
rect -4415 9475 -4365 9525
rect -4315 9475 -4265 9525
rect -4220 9475 -4170 9525
rect -4125 9475 -4075 9525
rect -4005 9475 -3955 9525
rect -3910 9475 -3860 9525
rect -3815 9475 -3765 9525
rect -3715 9475 -3665 9525
rect -3615 9475 -3565 9525
rect -3515 9475 -3465 9525
rect -3420 9475 -3370 9525
rect -3325 9475 -3275 9525
rect -3205 9475 -3155 9525
rect -3110 9475 -3060 9525
rect -3015 9475 -2965 9525
rect -2915 9475 -2865 9525
rect -2815 9475 -2765 9525
rect -2715 9475 -2665 9525
rect -2620 9475 -2570 9525
rect -2525 9475 -2475 9525
rect -2405 9475 -2355 9525
rect -2310 9475 -2260 9525
rect -2215 9475 -2165 9525
rect -2115 9475 -2065 9525
rect -2015 9475 -1965 9525
rect -1915 9475 -1865 9525
rect -1820 9475 -1770 9525
rect -1725 9475 -1675 9525
rect -4805 9375 -4755 9425
rect -4710 9375 -4660 9425
rect -4615 9375 -4565 9425
rect -4515 9375 -4465 9425
rect -4415 9375 -4365 9425
rect -4315 9375 -4265 9425
rect -4220 9375 -4170 9425
rect -4125 9375 -4075 9425
rect -4005 9375 -3955 9425
rect -3910 9375 -3860 9425
rect -3815 9375 -3765 9425
rect -3715 9375 -3665 9425
rect -3615 9375 -3565 9425
rect -3515 9375 -3465 9425
rect -3420 9375 -3370 9425
rect -3325 9375 -3275 9425
rect -3205 9375 -3155 9425
rect -3110 9375 -3060 9425
rect -3015 9375 -2965 9425
rect -2915 9375 -2865 9425
rect -2815 9375 -2765 9425
rect -2715 9375 -2665 9425
rect -2620 9375 -2570 9425
rect -2525 9375 -2475 9425
rect -2405 9375 -2355 9425
rect -2310 9375 -2260 9425
rect -2215 9375 -2165 9425
rect -2115 9375 -2065 9425
rect -2015 9375 -1965 9425
rect -1915 9375 -1865 9425
rect -1820 9375 -1770 9425
rect -1725 9375 -1675 9425
rect -4805 9285 -4755 9335
rect -4710 9285 -4660 9335
rect -4615 9285 -4565 9335
rect -4515 9285 -4465 9335
rect -4415 9285 -4365 9335
rect -4315 9285 -4265 9335
rect -4220 9285 -4170 9335
rect -4125 9285 -4075 9335
rect -4005 9285 -3955 9335
rect -3910 9285 -3860 9335
rect -3815 9285 -3765 9335
rect -3715 9285 -3665 9335
rect -3615 9285 -3565 9335
rect -3515 9285 -3465 9335
rect -3420 9285 -3370 9335
rect -3325 9285 -3275 9335
rect -3205 9285 -3155 9335
rect -3110 9285 -3060 9335
rect -3015 9285 -2965 9335
rect -2915 9285 -2865 9335
rect -2815 9285 -2765 9335
rect -2715 9285 -2665 9335
rect -2620 9285 -2570 9335
rect -2525 9285 -2475 9335
rect -2405 9285 -2355 9335
rect -2310 9285 -2260 9335
rect -2215 9285 -2165 9335
rect -2115 9285 -2065 9335
rect -2015 9285 -1965 9335
rect -1915 9285 -1865 9335
rect -1820 9285 -1770 9335
rect -1725 9285 -1675 9335
rect -4805 9165 -4755 9215
rect -4710 9165 -4660 9215
rect -4615 9165 -4565 9215
rect -4515 9165 -4465 9215
rect -4415 9165 -4365 9215
rect -4315 9165 -4265 9215
rect -4220 9165 -4170 9215
rect -4125 9165 -4075 9215
rect -4005 9165 -3955 9215
rect -3910 9165 -3860 9215
rect -3815 9165 -3765 9215
rect -3715 9165 -3665 9215
rect -3615 9165 -3565 9215
rect -3515 9165 -3465 9215
rect -3420 9165 -3370 9215
rect -3325 9165 -3275 9215
rect -3205 9165 -3155 9215
rect -3110 9165 -3060 9215
rect -3015 9165 -2965 9215
rect -2915 9165 -2865 9215
rect -2815 9165 -2765 9215
rect -2715 9165 -2665 9215
rect -2620 9165 -2570 9215
rect -2525 9165 -2475 9215
rect -2405 9165 -2355 9215
rect -2310 9165 -2260 9215
rect -2215 9165 -2165 9215
rect -2115 9165 -2065 9215
rect -2015 9165 -1965 9215
rect -1915 9165 -1865 9215
rect -1820 9165 -1770 9215
rect -1725 9165 -1675 9215
rect -4805 9075 -4755 9125
rect -4710 9075 -4660 9125
rect -4615 9075 -4565 9125
rect -4515 9075 -4465 9125
rect -4415 9075 -4365 9125
rect -4315 9075 -4265 9125
rect -4220 9075 -4170 9125
rect -4125 9075 -4075 9125
rect -4005 9075 -3955 9125
rect -3910 9075 -3860 9125
rect -3815 9075 -3765 9125
rect -3715 9075 -3665 9125
rect -3615 9075 -3565 9125
rect -3515 9075 -3465 9125
rect -3420 9075 -3370 9125
rect -3325 9075 -3275 9125
rect -3205 9075 -3155 9125
rect -3110 9075 -3060 9125
rect -3015 9075 -2965 9125
rect -2915 9075 -2865 9125
rect -2815 9075 -2765 9125
rect -2715 9075 -2665 9125
rect -2620 9075 -2570 9125
rect -2525 9075 -2475 9125
rect -2405 9075 -2355 9125
rect -2310 9075 -2260 9125
rect -2215 9075 -2165 9125
rect -2115 9075 -2065 9125
rect -2015 9075 -1965 9125
rect -1915 9075 -1865 9125
rect -1820 9075 -1770 9125
rect -1725 9075 -1675 9125
rect -4805 8975 -4755 9025
rect -4710 8975 -4660 9025
rect -4615 8975 -4565 9025
rect -4515 8975 -4465 9025
rect -4415 8975 -4365 9025
rect -4315 8975 -4265 9025
rect -4220 8975 -4170 9025
rect -4125 8975 -4075 9025
rect -4005 8975 -3955 9025
rect -3910 8975 -3860 9025
rect -3815 8975 -3765 9025
rect -3715 8975 -3665 9025
rect -3615 8975 -3565 9025
rect -3515 8975 -3465 9025
rect -3420 8975 -3370 9025
rect -3325 8975 -3275 9025
rect -3205 8975 -3155 9025
rect -3110 8975 -3060 9025
rect -3015 8975 -2965 9025
rect -2915 8975 -2865 9025
rect -2815 8975 -2765 9025
rect -2715 8975 -2665 9025
rect -2620 8975 -2570 9025
rect -2525 8975 -2475 9025
rect -2405 8975 -2355 9025
rect -2310 8975 -2260 9025
rect -2215 8975 -2165 9025
rect -2115 8975 -2065 9025
rect -2015 8975 -1965 9025
rect -1915 8975 -1865 9025
rect -1820 8975 -1770 9025
rect -1725 8975 -1675 9025
rect -4805 8885 -4755 8935
rect -4710 8885 -4660 8935
rect -4615 8885 -4565 8935
rect -4515 8885 -4465 8935
rect -4415 8885 -4365 8935
rect -4315 8885 -4265 8935
rect -4220 8885 -4170 8935
rect -4125 8885 -4075 8935
rect -4005 8885 -3955 8935
rect -3910 8885 -3860 8935
rect -3815 8885 -3765 8935
rect -3715 8885 -3665 8935
rect -3615 8885 -3565 8935
rect -3515 8885 -3465 8935
rect -3420 8885 -3370 8935
rect -3325 8885 -3275 8935
rect -3205 8885 -3155 8935
rect -3110 8885 -3060 8935
rect -3015 8885 -2965 8935
rect -2915 8885 -2865 8935
rect -2815 8885 -2765 8935
rect -2715 8885 -2665 8935
rect -2620 8885 -2570 8935
rect -2525 8885 -2475 8935
rect -2405 8885 -2355 8935
rect -2310 8885 -2260 8935
rect -2215 8885 -2165 8935
rect -2115 8885 -2065 8935
rect -2015 8885 -1965 8935
rect -1915 8885 -1865 8935
rect -1820 8885 -1770 8935
rect -1725 8885 -1675 8935
rect -4805 8765 -4755 8815
rect -4710 8765 -4660 8815
rect -4615 8765 -4565 8815
rect -4515 8765 -4465 8815
rect -4415 8765 -4365 8815
rect -4315 8765 -4265 8815
rect -4220 8765 -4170 8815
rect -4125 8765 -4075 8815
rect -4005 8765 -3955 8815
rect -3910 8765 -3860 8815
rect -3815 8765 -3765 8815
rect -3715 8765 -3665 8815
rect -3615 8765 -3565 8815
rect -3515 8765 -3465 8815
rect -3420 8765 -3370 8815
rect -3325 8765 -3275 8815
rect -3205 8765 -3155 8815
rect -3110 8765 -3060 8815
rect -3015 8765 -2965 8815
rect -2915 8765 -2865 8815
rect -2815 8765 -2765 8815
rect -2715 8765 -2665 8815
rect -2620 8765 -2570 8815
rect -2525 8765 -2475 8815
rect -2405 8765 -2355 8815
rect -2310 8765 -2260 8815
rect -2215 8765 -2165 8815
rect -2115 8765 -2065 8815
rect -2015 8765 -1965 8815
rect -1915 8765 -1865 8815
rect -1820 8765 -1770 8815
rect -1725 8765 -1675 8815
rect -4805 8675 -4755 8725
rect -4710 8675 -4660 8725
rect -4615 8675 -4565 8725
rect -4515 8675 -4465 8725
rect -4415 8675 -4365 8725
rect -4315 8675 -4265 8725
rect -4220 8675 -4170 8725
rect -4125 8675 -4075 8725
rect -4005 8675 -3955 8725
rect -3910 8675 -3860 8725
rect -3815 8675 -3765 8725
rect -3715 8675 -3665 8725
rect -3615 8675 -3565 8725
rect -3515 8675 -3465 8725
rect -3420 8675 -3370 8725
rect -3325 8675 -3275 8725
rect -3205 8675 -3155 8725
rect -3110 8675 -3060 8725
rect -3015 8675 -2965 8725
rect -2915 8675 -2865 8725
rect -2815 8675 -2765 8725
rect -2715 8675 -2665 8725
rect -2620 8675 -2570 8725
rect -2525 8675 -2475 8725
rect -2405 8675 -2355 8725
rect -2310 8675 -2260 8725
rect -2215 8675 -2165 8725
rect -2115 8675 -2065 8725
rect -2015 8675 -1965 8725
rect -1915 8675 -1865 8725
rect -1820 8675 -1770 8725
rect -1725 8675 -1675 8725
rect -4805 8575 -4755 8625
rect -4710 8575 -4660 8625
rect -4615 8575 -4565 8625
rect -4515 8575 -4465 8625
rect -4415 8575 -4365 8625
rect -4315 8575 -4265 8625
rect -4220 8575 -4170 8625
rect -4125 8575 -4075 8625
rect -4005 8575 -3955 8625
rect -3910 8575 -3860 8625
rect -3815 8575 -3765 8625
rect -3715 8575 -3665 8625
rect -3615 8575 -3565 8625
rect -3515 8575 -3465 8625
rect -3420 8575 -3370 8625
rect -3325 8575 -3275 8625
rect -3205 8575 -3155 8625
rect -3110 8575 -3060 8625
rect -3015 8575 -2965 8625
rect -2915 8575 -2865 8625
rect -2815 8575 -2765 8625
rect -2715 8575 -2665 8625
rect -2620 8575 -2570 8625
rect -2525 8575 -2475 8625
rect -2405 8575 -2355 8625
rect -2310 8575 -2260 8625
rect -2215 8575 -2165 8625
rect -2115 8575 -2065 8625
rect -2015 8575 -1965 8625
rect -1915 8575 -1865 8625
rect -1820 8575 -1770 8625
rect -1725 8575 -1675 8625
rect -4805 8485 -4755 8535
rect -4710 8485 -4660 8535
rect -4615 8485 -4565 8535
rect -4515 8485 -4465 8535
rect -4415 8485 -4365 8535
rect -4315 8485 -4265 8535
rect -4220 8485 -4170 8535
rect -4125 8485 -4075 8535
rect -4005 8485 -3955 8535
rect -3910 8485 -3860 8535
rect -3815 8485 -3765 8535
rect -3715 8485 -3665 8535
rect -3615 8485 -3565 8535
rect -3515 8485 -3465 8535
rect -3420 8485 -3370 8535
rect -3325 8485 -3275 8535
rect -3205 8485 -3155 8535
rect -3110 8485 -3060 8535
rect -3015 8485 -2965 8535
rect -2915 8485 -2865 8535
rect -2815 8485 -2765 8535
rect -2715 8485 -2665 8535
rect -2620 8485 -2570 8535
rect -2525 8485 -2475 8535
rect -2405 8485 -2355 8535
rect -2310 8485 -2260 8535
rect -2215 8485 -2165 8535
rect -2115 8485 -2065 8535
rect -2015 8485 -1965 8535
rect -1915 8485 -1865 8535
rect -1820 8485 -1770 8535
rect -1725 8485 -1675 8535
rect -4805 8365 -4755 8415
rect -4710 8365 -4660 8415
rect -4615 8365 -4565 8415
rect -4515 8365 -4465 8415
rect -4415 8365 -4365 8415
rect -4315 8365 -4265 8415
rect -4220 8365 -4170 8415
rect -4125 8365 -4075 8415
rect -4005 8365 -3955 8415
rect -3910 8365 -3860 8415
rect -3815 8365 -3765 8415
rect -3715 8365 -3665 8415
rect -3615 8365 -3565 8415
rect -3515 8365 -3465 8415
rect -3420 8365 -3370 8415
rect -3325 8365 -3275 8415
rect -3205 8365 -3155 8415
rect -3110 8365 -3060 8415
rect -3015 8365 -2965 8415
rect -2915 8365 -2865 8415
rect -2815 8365 -2765 8415
rect -2715 8365 -2665 8415
rect -2620 8365 -2570 8415
rect -2525 8365 -2475 8415
rect -2405 8365 -2355 8415
rect -2310 8365 -2260 8415
rect -2215 8365 -2165 8415
rect -2115 8365 -2065 8415
rect -2015 8365 -1965 8415
rect -1915 8365 -1865 8415
rect -1820 8365 -1770 8415
rect -1725 8365 -1675 8415
rect -4805 8275 -4755 8325
rect -4710 8275 -4660 8325
rect -4615 8275 -4565 8325
rect -4515 8275 -4465 8325
rect -4415 8275 -4365 8325
rect -4315 8275 -4265 8325
rect -4220 8275 -4170 8325
rect -4125 8275 -4075 8325
rect -4005 8275 -3955 8325
rect -3910 8275 -3860 8325
rect -3815 8275 -3765 8325
rect -3715 8275 -3665 8325
rect -3615 8275 -3565 8325
rect -3515 8275 -3465 8325
rect -3420 8275 -3370 8325
rect -3325 8275 -3275 8325
rect -3205 8275 -3155 8325
rect -3110 8275 -3060 8325
rect -3015 8275 -2965 8325
rect -2915 8275 -2865 8325
rect -2815 8275 -2765 8325
rect -2715 8275 -2665 8325
rect -2620 8275 -2570 8325
rect -2525 8275 -2475 8325
rect -2405 8275 -2355 8325
rect -2310 8275 -2260 8325
rect -2215 8275 -2165 8325
rect -2115 8275 -2065 8325
rect -2015 8275 -1965 8325
rect -1915 8275 -1865 8325
rect -1820 8275 -1770 8325
rect -1725 8275 -1675 8325
rect -4805 8175 -4755 8225
rect -4710 8175 -4660 8225
rect -4615 8175 -4565 8225
rect -4515 8175 -4465 8225
rect -4415 8175 -4365 8225
rect -4315 8175 -4265 8225
rect -4220 8175 -4170 8225
rect -4125 8175 -4075 8225
rect -4005 8175 -3955 8225
rect -3910 8175 -3860 8225
rect -3815 8175 -3765 8225
rect -3715 8175 -3665 8225
rect -3615 8175 -3565 8225
rect -3515 8175 -3465 8225
rect -3420 8175 -3370 8225
rect -3325 8175 -3275 8225
rect -3205 8175 -3155 8225
rect -3110 8175 -3060 8225
rect -3015 8175 -2965 8225
rect -2915 8175 -2865 8225
rect -2815 8175 -2765 8225
rect -2715 8175 -2665 8225
rect -2620 8175 -2570 8225
rect -2525 8175 -2475 8225
rect -2405 8175 -2355 8225
rect -2310 8175 -2260 8225
rect -2215 8175 -2165 8225
rect -2115 8175 -2065 8225
rect -2015 8175 -1965 8225
rect -1915 8175 -1865 8225
rect -1820 8175 -1770 8225
rect -1725 8175 -1675 8225
rect -4805 8085 -4755 8135
rect -4710 8085 -4660 8135
rect -4615 8085 -4565 8135
rect -4515 8085 -4465 8135
rect -4415 8085 -4365 8135
rect -4315 8085 -4265 8135
rect -4220 8085 -4170 8135
rect -4125 8085 -4075 8135
rect -4005 8085 -3955 8135
rect -3910 8085 -3860 8135
rect -3815 8085 -3765 8135
rect -3715 8085 -3665 8135
rect -3615 8085 -3565 8135
rect -3515 8085 -3465 8135
rect -3420 8085 -3370 8135
rect -3325 8085 -3275 8135
rect -3205 8085 -3155 8135
rect -3110 8085 -3060 8135
rect -3015 8085 -2965 8135
rect -2915 8085 -2865 8135
rect -2815 8085 -2765 8135
rect -2715 8085 -2665 8135
rect -2620 8085 -2570 8135
rect -2525 8085 -2475 8135
rect -2405 8085 -2355 8135
rect -2310 8085 -2260 8135
rect -2215 8085 -2165 8135
rect -2115 8085 -2065 8135
rect -2015 8085 -1965 8135
rect -1915 8085 -1865 8135
rect -1820 8085 -1770 8135
rect -1725 8085 -1675 8135
rect -4805 7965 -4755 8015
rect -4710 7965 -4660 8015
rect -4615 7965 -4565 8015
rect -4515 7965 -4465 8015
rect -4415 7965 -4365 8015
rect -4315 7965 -4265 8015
rect -4220 7965 -4170 8015
rect -4125 7965 -4075 8015
rect -4005 7965 -3955 8015
rect -3910 7965 -3860 8015
rect -3815 7965 -3765 8015
rect -3715 7965 -3665 8015
rect -3615 7965 -3565 8015
rect -3515 7965 -3465 8015
rect -3420 7965 -3370 8015
rect -3325 7965 -3275 8015
rect -3205 7965 -3155 8015
rect -3110 7965 -3060 8015
rect -3015 7965 -2965 8015
rect -2915 7965 -2865 8015
rect -2815 7965 -2765 8015
rect -2715 7965 -2665 8015
rect -2620 7965 -2570 8015
rect -2525 7965 -2475 8015
rect -2405 7965 -2355 8015
rect -2310 7965 -2260 8015
rect -2215 7965 -2165 8015
rect -2115 7965 -2065 8015
rect -2015 7965 -1965 8015
rect -1915 7965 -1865 8015
rect -1820 7965 -1770 8015
rect -1725 7965 -1675 8015
rect -4805 7875 -4755 7925
rect -4710 7875 -4660 7925
rect -4615 7875 -4565 7925
rect -4515 7875 -4465 7925
rect -4415 7875 -4365 7925
rect -4315 7875 -4265 7925
rect -4220 7875 -4170 7925
rect -4125 7875 -4075 7925
rect -4005 7875 -3955 7925
rect -3910 7875 -3860 7925
rect -3815 7875 -3765 7925
rect -3715 7875 -3665 7925
rect -3615 7875 -3565 7925
rect -3515 7875 -3465 7925
rect -3420 7875 -3370 7925
rect -3325 7875 -3275 7925
rect -3205 7875 -3155 7925
rect -3110 7875 -3060 7925
rect -3015 7875 -2965 7925
rect -2915 7875 -2865 7925
rect -2815 7875 -2765 7925
rect -2715 7875 -2665 7925
rect -2620 7875 -2570 7925
rect -2525 7875 -2475 7925
rect -2405 7875 -2355 7925
rect -2310 7875 -2260 7925
rect -2215 7875 -2165 7925
rect -2115 7875 -2065 7925
rect -2015 7875 -1965 7925
rect -1915 7875 -1865 7925
rect -1820 7875 -1770 7925
rect -1725 7875 -1675 7925
rect -4805 7775 -4755 7825
rect -4710 7775 -4660 7825
rect -4615 7775 -4565 7825
rect -4515 7775 -4465 7825
rect -4415 7775 -4365 7825
rect -4315 7775 -4265 7825
rect -4220 7775 -4170 7825
rect -4125 7775 -4075 7825
rect -4005 7775 -3955 7825
rect -3910 7775 -3860 7825
rect -3815 7775 -3765 7825
rect -3715 7775 -3665 7825
rect -3615 7775 -3565 7825
rect -3515 7775 -3465 7825
rect -3420 7775 -3370 7825
rect -3325 7775 -3275 7825
rect -3205 7775 -3155 7825
rect -3110 7775 -3060 7825
rect -3015 7775 -2965 7825
rect -2915 7775 -2865 7825
rect -2815 7775 -2765 7825
rect -2715 7775 -2665 7825
rect -2620 7775 -2570 7825
rect -2525 7775 -2475 7825
rect -2405 7775 -2355 7825
rect -2310 7775 -2260 7825
rect -2215 7775 -2165 7825
rect -2115 7775 -2065 7825
rect -2015 7775 -1965 7825
rect -1915 7775 -1865 7825
rect -1820 7775 -1770 7825
rect -1725 7775 -1675 7825
rect -4805 7685 -4755 7735
rect -4710 7685 -4660 7735
rect -4615 7685 -4565 7735
rect -4515 7685 -4465 7735
rect -4415 7685 -4365 7735
rect -4315 7685 -4265 7735
rect -4220 7685 -4170 7735
rect -4125 7685 -4075 7735
rect -4005 7685 -3955 7735
rect -3910 7685 -3860 7735
rect -3815 7685 -3765 7735
rect -3715 7685 -3665 7735
rect -3615 7685 -3565 7735
rect -3515 7685 -3465 7735
rect -3420 7685 -3370 7735
rect -3325 7685 -3275 7735
rect -3205 7685 -3155 7735
rect -3110 7685 -3060 7735
rect -3015 7685 -2965 7735
rect -2915 7685 -2865 7735
rect -2815 7685 -2765 7735
rect -2715 7685 -2665 7735
rect -2620 7685 -2570 7735
rect -2525 7685 -2475 7735
rect -2405 7685 -2355 7735
rect -2310 7685 -2260 7735
rect -2215 7685 -2165 7735
rect -2115 7685 -2065 7735
rect -2015 7685 -1965 7735
rect -1915 7685 -1865 7735
rect -1820 7685 -1770 7735
rect -1725 7685 -1675 7735
rect -4805 7565 -4755 7615
rect -4710 7565 -4660 7615
rect -4615 7565 -4565 7615
rect -4515 7565 -4465 7615
rect -4415 7565 -4365 7615
rect -4315 7565 -4265 7615
rect -4220 7565 -4170 7615
rect -4125 7565 -4075 7615
rect -4005 7565 -3955 7615
rect -3910 7565 -3860 7615
rect -3815 7565 -3765 7615
rect -3715 7565 -3665 7615
rect -3615 7565 -3565 7615
rect -3515 7565 -3465 7615
rect -3420 7565 -3370 7615
rect -3325 7565 -3275 7615
rect -3205 7565 -3155 7615
rect -3110 7565 -3060 7615
rect -3015 7565 -2965 7615
rect -2915 7565 -2865 7615
rect -2815 7565 -2765 7615
rect -2715 7565 -2665 7615
rect -2620 7565 -2570 7615
rect -2525 7565 -2475 7615
rect -2405 7565 -2355 7615
rect -2310 7565 -2260 7615
rect -2215 7565 -2165 7615
rect -2115 7565 -2065 7615
rect -2015 7565 -1965 7615
rect -1915 7565 -1865 7615
rect -1820 7565 -1770 7615
rect -1725 7565 -1675 7615
rect -4805 7475 -4755 7525
rect -4710 7475 -4660 7525
rect -4615 7475 -4565 7525
rect -4515 7475 -4465 7525
rect -4415 7475 -4365 7525
rect -4315 7475 -4265 7525
rect -4220 7475 -4170 7525
rect -4125 7475 -4075 7525
rect -4005 7475 -3955 7525
rect -3910 7475 -3860 7525
rect -3815 7475 -3765 7525
rect -3715 7475 -3665 7525
rect -3615 7475 -3565 7525
rect -3515 7475 -3465 7525
rect -3420 7475 -3370 7525
rect -3325 7475 -3275 7525
rect -3205 7475 -3155 7525
rect -3110 7475 -3060 7525
rect -3015 7475 -2965 7525
rect -2915 7475 -2865 7525
rect -2815 7475 -2765 7525
rect -2715 7475 -2665 7525
rect -2620 7475 -2570 7525
rect -2525 7475 -2475 7525
rect -2405 7475 -2355 7525
rect -2310 7475 -2260 7525
rect -2215 7475 -2165 7525
rect -2115 7475 -2065 7525
rect -2015 7475 -1965 7525
rect -1915 7475 -1865 7525
rect -1820 7475 -1770 7525
rect -1725 7475 -1675 7525
rect -4805 7375 -4755 7425
rect -4710 7375 -4660 7425
rect -4615 7375 -4565 7425
rect -4515 7375 -4465 7425
rect -4415 7375 -4365 7425
rect -4315 7375 -4265 7425
rect -4220 7375 -4170 7425
rect -4125 7375 -4075 7425
rect -4005 7375 -3955 7425
rect -3910 7375 -3860 7425
rect -3815 7375 -3765 7425
rect -3715 7375 -3665 7425
rect -3615 7375 -3565 7425
rect -3515 7375 -3465 7425
rect -3420 7375 -3370 7425
rect -3325 7375 -3275 7425
rect -3205 7375 -3155 7425
rect -3110 7375 -3060 7425
rect -3015 7375 -2965 7425
rect -2915 7375 -2865 7425
rect -2815 7375 -2765 7425
rect -2715 7375 -2665 7425
rect -2620 7375 -2570 7425
rect -2525 7375 -2475 7425
rect -2405 7375 -2355 7425
rect -2310 7375 -2260 7425
rect -2215 7375 -2165 7425
rect -2115 7375 -2065 7425
rect -2015 7375 -1965 7425
rect -1915 7375 -1865 7425
rect -1820 7375 -1770 7425
rect -1725 7375 -1675 7425
rect -4805 7285 -4755 7335
rect -4710 7285 -4660 7335
rect -4615 7285 -4565 7335
rect -4515 7285 -4465 7335
rect -4415 7285 -4365 7335
rect -4315 7285 -4265 7335
rect -4220 7285 -4170 7335
rect -4125 7285 -4075 7335
rect -4005 7285 -3955 7335
rect -3910 7285 -3860 7335
rect -3815 7285 -3765 7335
rect -3715 7285 -3665 7335
rect -3615 7285 -3565 7335
rect -3515 7285 -3465 7335
rect -3420 7285 -3370 7335
rect -3325 7285 -3275 7335
rect -3205 7285 -3155 7335
rect -3110 7285 -3060 7335
rect -3015 7285 -2965 7335
rect -2915 7285 -2865 7335
rect -2815 7285 -2765 7335
rect -2715 7285 -2665 7335
rect -2620 7285 -2570 7335
rect -2525 7285 -2475 7335
rect -2405 7285 -2355 7335
rect -2310 7285 -2260 7335
rect -2215 7285 -2165 7335
rect -2115 7285 -2065 7335
rect -2015 7285 -1965 7335
rect -1915 7285 -1865 7335
rect -1820 7285 -1770 7335
rect -1725 7285 -1675 7335
rect -4805 7165 -4755 7215
rect -4710 7165 -4660 7215
rect -4615 7165 -4565 7215
rect -4515 7165 -4465 7215
rect -4415 7165 -4365 7215
rect -4315 7165 -4265 7215
rect -4220 7165 -4170 7215
rect -4125 7165 -4075 7215
rect -4005 7165 -3955 7215
rect -3910 7165 -3860 7215
rect -3815 7165 -3765 7215
rect -3715 7165 -3665 7215
rect -3615 7165 -3565 7215
rect -3515 7165 -3465 7215
rect -3420 7165 -3370 7215
rect -3325 7165 -3275 7215
rect -3205 7165 -3155 7215
rect -3110 7165 -3060 7215
rect -3015 7165 -2965 7215
rect -2915 7165 -2865 7215
rect -2815 7165 -2765 7215
rect -2715 7165 -2665 7215
rect -2620 7165 -2570 7215
rect -2525 7165 -2475 7215
rect -2405 7165 -2355 7215
rect -2310 7165 -2260 7215
rect -2215 7165 -2165 7215
rect -2115 7165 -2065 7215
rect -2015 7165 -1965 7215
rect -1915 7165 -1865 7215
rect -1820 7165 -1770 7215
rect -1725 7165 -1675 7215
rect -4805 7075 -4755 7125
rect -4710 7075 -4660 7125
rect -4615 7075 -4565 7125
rect -4515 7075 -4465 7125
rect -4415 7075 -4365 7125
rect -4315 7075 -4265 7125
rect -4220 7075 -4170 7125
rect -4125 7075 -4075 7125
rect -4005 7075 -3955 7125
rect -3910 7075 -3860 7125
rect -3815 7075 -3765 7125
rect -3715 7075 -3665 7125
rect -3615 7075 -3565 7125
rect -3515 7075 -3465 7125
rect -3420 7075 -3370 7125
rect -3325 7075 -3275 7125
rect -3205 7075 -3155 7125
rect -3110 7075 -3060 7125
rect -3015 7075 -2965 7125
rect -2915 7075 -2865 7125
rect -2815 7075 -2765 7125
rect -2715 7075 -2665 7125
rect -2620 7075 -2570 7125
rect -2525 7075 -2475 7125
rect -2405 7075 -2355 7125
rect -2310 7075 -2260 7125
rect -2215 7075 -2165 7125
rect -2115 7075 -2065 7125
rect -2015 7075 -1965 7125
rect -1915 7075 -1865 7125
rect -1820 7075 -1770 7125
rect -1725 7075 -1675 7125
rect -4805 6975 -4755 7025
rect -4710 6975 -4660 7025
rect -4615 6975 -4565 7025
rect -4515 6975 -4465 7025
rect -4415 6975 -4365 7025
rect -4315 6975 -4265 7025
rect -4220 6975 -4170 7025
rect -4125 6975 -4075 7025
rect -4005 6975 -3955 7025
rect -3910 6975 -3860 7025
rect -3815 6975 -3765 7025
rect -3715 6975 -3665 7025
rect -3615 6975 -3565 7025
rect -3515 6975 -3465 7025
rect -3420 6975 -3370 7025
rect -3325 6975 -3275 7025
rect -3205 6975 -3155 7025
rect -3110 6975 -3060 7025
rect -3015 6975 -2965 7025
rect -2915 6975 -2865 7025
rect -2815 6975 -2765 7025
rect -2715 6975 -2665 7025
rect -2620 6975 -2570 7025
rect -2525 6975 -2475 7025
rect -2405 6975 -2355 7025
rect -2310 6975 -2260 7025
rect -2215 6975 -2165 7025
rect -2115 6975 -2065 7025
rect -2015 6975 -1965 7025
rect -1915 6975 -1865 7025
rect -1820 6975 -1770 7025
rect -1725 6975 -1675 7025
rect -4805 6885 -4755 6935
rect -4710 6885 -4660 6935
rect -4615 6885 -4565 6935
rect -4515 6885 -4465 6935
rect -4415 6885 -4365 6935
rect -4315 6885 -4265 6935
rect -4220 6885 -4170 6935
rect -4125 6885 -4075 6935
rect -4005 6885 -3955 6935
rect -3910 6885 -3860 6935
rect -3815 6885 -3765 6935
rect -3715 6885 -3665 6935
rect -3615 6885 -3565 6935
rect -3515 6885 -3465 6935
rect -3420 6885 -3370 6935
rect -3325 6885 -3275 6935
rect -3205 6885 -3155 6935
rect -3110 6885 -3060 6935
rect -3015 6885 -2965 6935
rect -2915 6885 -2865 6935
rect -2815 6885 -2765 6935
rect -2715 6885 -2665 6935
rect -2620 6885 -2570 6935
rect -2525 6885 -2475 6935
rect -2405 6885 -2355 6935
rect -2310 6885 -2260 6935
rect -2215 6885 -2165 6935
rect -2115 6885 -2065 6935
rect -2015 6885 -1965 6935
rect -1915 6885 -1865 6935
rect -1820 6885 -1770 6935
rect -1725 6885 -1675 6935
rect -4805 6765 -4755 6815
rect -4710 6765 -4660 6815
rect -4615 6765 -4565 6815
rect -4515 6765 -4465 6815
rect -4415 6765 -4365 6815
rect -4315 6765 -4265 6815
rect -4220 6765 -4170 6815
rect -4125 6765 -4075 6815
rect -4005 6765 -3955 6815
rect -3910 6765 -3860 6815
rect -3815 6765 -3765 6815
rect -3715 6765 -3665 6815
rect -3615 6765 -3565 6815
rect -3515 6765 -3465 6815
rect -3420 6765 -3370 6815
rect -3325 6765 -3275 6815
rect -3205 6765 -3155 6815
rect -3110 6765 -3060 6815
rect -3015 6765 -2965 6815
rect -2915 6765 -2865 6815
rect -2815 6765 -2765 6815
rect -2715 6765 -2665 6815
rect -2620 6765 -2570 6815
rect -2525 6765 -2475 6815
rect -2405 6765 -2355 6815
rect -2310 6765 -2260 6815
rect -2215 6765 -2165 6815
rect -2115 6765 -2065 6815
rect -2015 6765 -1965 6815
rect -1915 6765 -1865 6815
rect -1820 6765 -1770 6815
rect -1725 6765 -1675 6815
rect -4805 6675 -4755 6725
rect -4710 6675 -4660 6725
rect -4615 6675 -4565 6725
rect -4515 6675 -4465 6725
rect -4415 6675 -4365 6725
rect -4315 6675 -4265 6725
rect -4220 6675 -4170 6725
rect -4125 6675 -4075 6725
rect -4005 6675 -3955 6725
rect -3910 6675 -3860 6725
rect -3815 6675 -3765 6725
rect -3715 6675 -3665 6725
rect -3615 6675 -3565 6725
rect -3515 6675 -3465 6725
rect -3420 6675 -3370 6725
rect -3325 6675 -3275 6725
rect -3205 6675 -3155 6725
rect -3110 6675 -3060 6725
rect -3015 6675 -2965 6725
rect -2915 6675 -2865 6725
rect -2815 6675 -2765 6725
rect -2715 6675 -2665 6725
rect -2620 6675 -2570 6725
rect -2525 6675 -2475 6725
rect -2405 6675 -2355 6725
rect -2310 6675 -2260 6725
rect -2215 6675 -2165 6725
rect -2115 6675 -2065 6725
rect -2015 6675 -1965 6725
rect -1915 6675 -1865 6725
rect -1820 6675 -1770 6725
rect -1725 6675 -1675 6725
rect -4805 6575 -4755 6625
rect -4710 6575 -4660 6625
rect -4615 6575 -4565 6625
rect -4515 6575 -4465 6625
rect -4415 6575 -4365 6625
rect -4315 6575 -4265 6625
rect -4220 6575 -4170 6625
rect -4125 6575 -4075 6625
rect -4005 6575 -3955 6625
rect -3910 6575 -3860 6625
rect -3815 6575 -3765 6625
rect -3715 6575 -3665 6625
rect -3615 6575 -3565 6625
rect -3515 6575 -3465 6625
rect -3420 6575 -3370 6625
rect -3325 6575 -3275 6625
rect -3205 6575 -3155 6625
rect -3110 6575 -3060 6625
rect -3015 6575 -2965 6625
rect -2915 6575 -2865 6625
rect -2815 6575 -2765 6625
rect -2715 6575 -2665 6625
rect -2620 6575 -2570 6625
rect -2525 6575 -2475 6625
rect -2405 6575 -2355 6625
rect -2310 6575 -2260 6625
rect -2215 6575 -2165 6625
rect -2115 6575 -2065 6625
rect -2015 6575 -1965 6625
rect -1915 6575 -1865 6625
rect -1820 6575 -1770 6625
rect -1725 6575 -1675 6625
rect -4805 6485 -4755 6535
rect -4710 6485 -4660 6535
rect -4615 6485 -4565 6535
rect -4515 6485 -4465 6535
rect -4415 6485 -4365 6535
rect -4315 6485 -4265 6535
rect -4220 6485 -4170 6535
rect -4125 6485 -4075 6535
rect -4005 6485 -3955 6535
rect -3910 6485 -3860 6535
rect -3815 6485 -3765 6535
rect -3715 6485 -3665 6535
rect -3615 6485 -3565 6535
rect -3515 6485 -3465 6535
rect -3420 6485 -3370 6535
rect -3325 6485 -3275 6535
rect -3205 6485 -3155 6535
rect -3110 6485 -3060 6535
rect -3015 6485 -2965 6535
rect -2915 6485 -2865 6535
rect -2815 6485 -2765 6535
rect -2715 6485 -2665 6535
rect -2620 6485 -2570 6535
rect -2525 6485 -2475 6535
rect -2405 6485 -2355 6535
rect -2310 6485 -2260 6535
rect -2215 6485 -2165 6535
rect -2115 6485 -2065 6535
rect -2015 6485 -1965 6535
rect -1915 6485 -1865 6535
rect -1820 6485 -1770 6535
rect -1725 6485 -1675 6535
rect -80 9635 -40 9640
rect -80 9605 -75 9635
rect -75 9605 -45 9635
rect -45 9605 -40 9635
rect -80 9600 -40 9605
rect -80 9570 -40 9575
rect -80 9540 -75 9570
rect -75 9540 -45 9570
rect -45 9540 -40 9570
rect -80 9535 -40 9540
rect -80 9500 -40 9505
rect -80 9470 -75 9500
rect -75 9470 -45 9500
rect -45 9470 -40 9500
rect -80 9465 -40 9470
rect -80 9430 -40 9435
rect -80 9400 -75 9430
rect -75 9400 -45 9430
rect -45 9400 -40 9430
rect -80 9395 -40 9400
rect -80 9360 -40 9365
rect -80 9330 -75 9360
rect -75 9330 -45 9360
rect -45 9330 -40 9360
rect -80 9325 -40 9330
rect -80 9295 -40 9300
rect -80 9265 -75 9295
rect -75 9265 -45 9295
rect -45 9265 -40 9295
rect -80 9260 -40 9265
rect -80 9235 -40 9240
rect -80 9205 -75 9235
rect -75 9205 -45 9235
rect -45 9205 -40 9235
rect -80 9200 -40 9205
rect -80 9170 -40 9175
rect -80 9140 -75 9170
rect -75 9140 -45 9170
rect -45 9140 -40 9170
rect -80 9135 -40 9140
rect -80 9100 -40 9105
rect -80 9070 -75 9100
rect -75 9070 -45 9100
rect -45 9070 -40 9100
rect -80 9065 -40 9070
rect -80 9030 -40 9035
rect -80 9000 -75 9030
rect -75 9000 -45 9030
rect -45 9000 -40 9030
rect -80 8995 -40 9000
rect -80 8960 -40 8965
rect -80 8930 -75 8960
rect -75 8930 -45 8960
rect -45 8930 -40 8960
rect -80 8925 -40 8930
rect -80 8895 -40 8900
rect -80 8865 -75 8895
rect -75 8865 -45 8895
rect -45 8865 -40 8895
rect -80 8860 -40 8865
rect -80 8835 -40 8840
rect -80 8805 -75 8835
rect -75 8805 -45 8835
rect -45 8805 -40 8835
rect -80 8800 -40 8805
rect -80 8770 -40 8775
rect -80 8740 -75 8770
rect -75 8740 -45 8770
rect -45 8740 -40 8770
rect -80 8735 -40 8740
rect -80 8700 -40 8705
rect -80 8670 -75 8700
rect -75 8670 -45 8700
rect -45 8670 -40 8700
rect -80 8665 -40 8670
rect -80 8630 -40 8635
rect -80 8600 -75 8630
rect -75 8600 -45 8630
rect -45 8600 -40 8630
rect -80 8595 -40 8600
rect -80 8560 -40 8565
rect -80 8530 -75 8560
rect -75 8530 -45 8560
rect -45 8530 -40 8560
rect -80 8525 -40 8530
rect -80 8495 -40 8500
rect -80 8465 -75 8495
rect -75 8465 -45 8495
rect -45 8465 -40 8495
rect -80 8460 -40 8465
rect -80 8435 -40 8440
rect -80 8405 -75 8435
rect -75 8405 -45 8435
rect -45 8405 -40 8435
rect -80 8400 -40 8405
rect -80 8370 -40 8375
rect -80 8340 -75 8370
rect -75 8340 -45 8370
rect -45 8340 -40 8370
rect -80 8335 -40 8340
rect -80 8300 -40 8305
rect -80 8270 -75 8300
rect -75 8270 -45 8300
rect -45 8270 -40 8300
rect -80 8265 -40 8270
rect -80 8230 -40 8235
rect -80 8200 -75 8230
rect -75 8200 -45 8230
rect -45 8200 -40 8230
rect -80 8195 -40 8200
rect -80 8160 -40 8165
rect -80 8130 -75 8160
rect -75 8130 -45 8160
rect -45 8130 -40 8160
rect -80 8125 -40 8130
rect -80 8095 -40 8100
rect -80 8065 -75 8095
rect -75 8065 -45 8095
rect -45 8065 -40 8095
rect -80 8060 -40 8065
rect -80 8035 -40 8040
rect -80 8005 -75 8035
rect -75 8005 -45 8035
rect -45 8005 -40 8035
rect -80 8000 -40 8005
rect -80 7970 -40 7975
rect -80 7940 -75 7970
rect -75 7940 -45 7970
rect -45 7940 -40 7970
rect -80 7935 -40 7940
rect -80 7900 -40 7905
rect -80 7870 -75 7900
rect -75 7870 -45 7900
rect -45 7870 -40 7900
rect -80 7865 -40 7870
rect -80 7830 -40 7835
rect -80 7800 -75 7830
rect -75 7800 -45 7830
rect -45 7800 -40 7830
rect -80 7795 -40 7800
rect -80 7760 -40 7765
rect -80 7730 -75 7760
rect -75 7730 -45 7760
rect -45 7730 -40 7760
rect -80 7725 -40 7730
rect -80 7695 -40 7700
rect -80 7665 -75 7695
rect -75 7665 -45 7695
rect -45 7665 -40 7695
rect -80 7660 -40 7665
rect -80 7635 -40 7640
rect -80 7605 -75 7635
rect -75 7605 -45 7635
rect -45 7605 -40 7635
rect -80 7600 -40 7605
rect -80 7570 -40 7575
rect -80 7540 -75 7570
rect -75 7540 -45 7570
rect -45 7540 -40 7570
rect -80 7535 -40 7540
rect -80 7500 -40 7505
rect -80 7470 -75 7500
rect -75 7470 -45 7500
rect -45 7470 -40 7500
rect -80 7465 -40 7470
rect -80 7430 -40 7435
rect -80 7400 -75 7430
rect -75 7400 -45 7430
rect -45 7400 -40 7430
rect -80 7395 -40 7400
rect -80 7360 -40 7365
rect -80 7330 -75 7360
rect -75 7330 -45 7360
rect -45 7330 -40 7360
rect -80 7325 -40 7330
rect -80 7295 -40 7300
rect -80 7265 -75 7295
rect -75 7265 -45 7295
rect -45 7265 -40 7295
rect -80 7260 -40 7265
rect -80 7235 -40 7240
rect -80 7205 -75 7235
rect -75 7205 -45 7235
rect -45 7205 -40 7235
rect -80 7200 -40 7205
rect -80 7170 -40 7175
rect -80 7140 -75 7170
rect -75 7140 -45 7170
rect -45 7140 -40 7170
rect -80 7135 -40 7140
rect -80 7100 -40 7105
rect -80 7070 -75 7100
rect -75 7070 -45 7100
rect -45 7070 -40 7100
rect -80 7065 -40 7070
rect -80 7030 -40 7035
rect -80 7000 -75 7030
rect -75 7000 -45 7030
rect -45 7000 -40 7030
rect -80 6995 -40 7000
rect -80 6960 -40 6965
rect -80 6930 -75 6960
rect -75 6930 -45 6960
rect -45 6930 -40 6960
rect -80 6925 -40 6930
rect -80 6895 -40 6900
rect -80 6865 -75 6895
rect -75 6865 -45 6895
rect -45 6865 -40 6895
rect -80 6860 -40 6865
rect -80 6835 -40 6840
rect -80 6805 -75 6835
rect -75 6805 -45 6835
rect -45 6805 -40 6835
rect -80 6800 -40 6805
rect -80 6770 -40 6775
rect -80 6740 -75 6770
rect -75 6740 -45 6770
rect -45 6740 -40 6770
rect -80 6735 -40 6740
rect -80 6700 -40 6705
rect -80 6670 -75 6700
rect -75 6670 -45 6700
rect -45 6670 -40 6700
rect -80 6665 -40 6670
rect -80 6630 -40 6635
rect -80 6600 -75 6630
rect -75 6600 -45 6630
rect -45 6600 -40 6630
rect -80 6595 -40 6600
rect -80 6560 -40 6565
rect -80 6530 -75 6560
rect -75 6530 -45 6560
rect -45 6530 -40 6560
rect -80 6525 -40 6530
rect -80 6495 -40 6500
rect -80 6465 -75 6495
rect -75 6465 -45 6495
rect -45 6465 -40 6495
rect -80 6460 -40 6465
rect 270 9635 310 9640
rect 270 9605 275 9635
rect 275 9605 305 9635
rect 305 9605 310 9635
rect 270 9600 310 9605
rect 270 9570 310 9575
rect 270 9540 275 9570
rect 275 9540 305 9570
rect 305 9540 310 9570
rect 270 9535 310 9540
rect 270 9500 310 9505
rect 270 9470 275 9500
rect 275 9470 305 9500
rect 305 9470 310 9500
rect 270 9465 310 9470
rect 270 9430 310 9435
rect 270 9400 275 9430
rect 275 9400 305 9430
rect 305 9400 310 9430
rect 270 9395 310 9400
rect 270 9360 310 9365
rect 270 9330 275 9360
rect 275 9330 305 9360
rect 305 9330 310 9360
rect 270 9325 310 9330
rect 270 9295 310 9300
rect 270 9265 275 9295
rect 275 9265 305 9295
rect 305 9265 310 9295
rect 270 9260 310 9265
rect 270 9235 310 9240
rect 270 9205 275 9235
rect 275 9205 305 9235
rect 305 9205 310 9235
rect 270 9200 310 9205
rect 270 9170 310 9175
rect 270 9140 275 9170
rect 275 9140 305 9170
rect 305 9140 310 9170
rect 270 9135 310 9140
rect 270 9100 310 9105
rect 270 9070 275 9100
rect 275 9070 305 9100
rect 305 9070 310 9100
rect 270 9065 310 9070
rect 270 9030 310 9035
rect 270 9000 275 9030
rect 275 9000 305 9030
rect 305 9000 310 9030
rect 270 8995 310 9000
rect 270 8960 310 8965
rect 270 8930 275 8960
rect 275 8930 305 8960
rect 305 8930 310 8960
rect 270 8925 310 8930
rect 270 8895 310 8900
rect 270 8865 275 8895
rect 275 8865 305 8895
rect 305 8865 310 8895
rect 270 8860 310 8865
rect 270 8835 310 8840
rect 270 8805 275 8835
rect 275 8805 305 8835
rect 305 8805 310 8835
rect 270 8800 310 8805
rect 270 8770 310 8775
rect 270 8740 275 8770
rect 275 8740 305 8770
rect 305 8740 310 8770
rect 270 8735 310 8740
rect 270 8700 310 8705
rect 270 8670 275 8700
rect 275 8670 305 8700
rect 305 8670 310 8700
rect 270 8665 310 8670
rect 270 8630 310 8635
rect 270 8600 275 8630
rect 275 8600 305 8630
rect 305 8600 310 8630
rect 270 8595 310 8600
rect 270 8560 310 8565
rect 270 8530 275 8560
rect 275 8530 305 8560
rect 305 8530 310 8560
rect 270 8525 310 8530
rect 270 8495 310 8500
rect 270 8465 275 8495
rect 275 8465 305 8495
rect 305 8465 310 8495
rect 270 8460 310 8465
rect 270 8435 310 8440
rect 270 8405 275 8435
rect 275 8405 305 8435
rect 305 8405 310 8435
rect 270 8400 310 8405
rect 270 8370 310 8375
rect 270 8340 275 8370
rect 275 8340 305 8370
rect 305 8340 310 8370
rect 270 8335 310 8340
rect 270 8300 310 8305
rect 270 8270 275 8300
rect 275 8270 305 8300
rect 305 8270 310 8300
rect 270 8265 310 8270
rect 270 8230 310 8235
rect 270 8200 275 8230
rect 275 8200 305 8230
rect 305 8200 310 8230
rect 270 8195 310 8200
rect 270 8160 310 8165
rect 270 8130 275 8160
rect 275 8130 305 8160
rect 305 8130 310 8160
rect 270 8125 310 8130
rect 270 8095 310 8100
rect 270 8065 275 8095
rect 275 8065 305 8095
rect 305 8065 310 8095
rect 270 8060 310 8065
rect 270 8035 310 8040
rect 270 8005 275 8035
rect 275 8005 305 8035
rect 305 8005 310 8035
rect 270 8000 310 8005
rect 270 7970 310 7975
rect 270 7940 275 7970
rect 275 7940 305 7970
rect 305 7940 310 7970
rect 270 7935 310 7940
rect 270 7900 310 7905
rect 270 7870 275 7900
rect 275 7870 305 7900
rect 305 7870 310 7900
rect 270 7865 310 7870
rect 270 7830 310 7835
rect 270 7800 275 7830
rect 275 7800 305 7830
rect 305 7800 310 7830
rect 270 7795 310 7800
rect 270 7760 310 7765
rect 270 7730 275 7760
rect 275 7730 305 7760
rect 305 7730 310 7760
rect 270 7725 310 7730
rect 270 7695 310 7700
rect 270 7665 275 7695
rect 275 7665 305 7695
rect 305 7665 310 7695
rect 270 7660 310 7665
rect 270 7635 310 7640
rect 270 7605 275 7635
rect 275 7605 305 7635
rect 305 7605 310 7635
rect 270 7600 310 7605
rect 270 7570 310 7575
rect 270 7540 275 7570
rect 275 7540 305 7570
rect 305 7540 310 7570
rect 270 7535 310 7540
rect 270 7500 310 7505
rect 270 7470 275 7500
rect 275 7470 305 7500
rect 305 7470 310 7500
rect 270 7465 310 7470
rect 270 7430 310 7435
rect 270 7400 275 7430
rect 275 7400 305 7430
rect 305 7400 310 7430
rect 270 7395 310 7400
rect 270 7360 310 7365
rect 270 7330 275 7360
rect 275 7330 305 7360
rect 305 7330 310 7360
rect 270 7325 310 7330
rect 270 7295 310 7300
rect 270 7265 275 7295
rect 275 7265 305 7295
rect 305 7265 310 7295
rect 270 7260 310 7265
rect 270 7235 310 7240
rect 270 7205 275 7235
rect 275 7205 305 7235
rect 305 7205 310 7235
rect 270 7200 310 7205
rect 270 7170 310 7175
rect 270 7140 275 7170
rect 275 7140 305 7170
rect 305 7140 310 7170
rect 270 7135 310 7140
rect 270 7100 310 7105
rect 270 7070 275 7100
rect 275 7070 305 7100
rect 305 7070 310 7100
rect 270 7065 310 7070
rect 270 7030 310 7035
rect 270 7000 275 7030
rect 275 7000 305 7030
rect 305 7000 310 7030
rect 270 6995 310 7000
rect 270 6960 310 6965
rect 270 6930 275 6960
rect 275 6930 305 6960
rect 305 6930 310 6960
rect 270 6925 310 6930
rect 270 6895 310 6900
rect 270 6865 275 6895
rect 275 6865 305 6895
rect 305 6865 310 6895
rect 270 6860 310 6865
rect 270 6835 310 6840
rect 270 6805 275 6835
rect 275 6805 305 6835
rect 305 6805 310 6835
rect 270 6800 310 6805
rect 270 6770 310 6775
rect 270 6740 275 6770
rect 275 6740 305 6770
rect 305 6740 310 6770
rect 270 6735 310 6740
rect 270 6700 310 6705
rect 270 6670 275 6700
rect 275 6670 305 6700
rect 305 6670 310 6700
rect 270 6665 310 6670
rect 270 6630 310 6635
rect 270 6600 275 6630
rect 275 6600 305 6630
rect 305 6600 310 6630
rect 270 6595 310 6600
rect 270 6560 310 6565
rect 270 6530 275 6560
rect 275 6530 305 6560
rect 305 6530 310 6560
rect 270 6525 310 6530
rect 270 6495 310 6500
rect 270 6465 275 6495
rect 275 6465 305 6495
rect 305 6465 310 6495
rect 270 6460 310 6465
rect 620 9635 660 9640
rect 620 9605 625 9635
rect 625 9605 655 9635
rect 655 9605 660 9635
rect 620 9600 660 9605
rect 620 9570 660 9575
rect 620 9540 625 9570
rect 625 9540 655 9570
rect 655 9540 660 9570
rect 620 9535 660 9540
rect 620 9500 660 9505
rect 620 9470 625 9500
rect 625 9470 655 9500
rect 655 9470 660 9500
rect 620 9465 660 9470
rect 620 9430 660 9435
rect 620 9400 625 9430
rect 625 9400 655 9430
rect 655 9400 660 9430
rect 620 9395 660 9400
rect 620 9360 660 9365
rect 620 9330 625 9360
rect 625 9330 655 9360
rect 655 9330 660 9360
rect 620 9325 660 9330
rect 620 9295 660 9300
rect 620 9265 625 9295
rect 625 9265 655 9295
rect 655 9265 660 9295
rect 620 9260 660 9265
rect 620 9235 660 9240
rect 620 9205 625 9235
rect 625 9205 655 9235
rect 655 9205 660 9235
rect 620 9200 660 9205
rect 620 9170 660 9175
rect 620 9140 625 9170
rect 625 9140 655 9170
rect 655 9140 660 9170
rect 620 9135 660 9140
rect 620 9100 660 9105
rect 620 9070 625 9100
rect 625 9070 655 9100
rect 655 9070 660 9100
rect 620 9065 660 9070
rect 620 9030 660 9035
rect 620 9000 625 9030
rect 625 9000 655 9030
rect 655 9000 660 9030
rect 620 8995 660 9000
rect 620 8960 660 8965
rect 620 8930 625 8960
rect 625 8930 655 8960
rect 655 8930 660 8960
rect 620 8925 660 8930
rect 620 8895 660 8900
rect 620 8865 625 8895
rect 625 8865 655 8895
rect 655 8865 660 8895
rect 620 8860 660 8865
rect 620 8835 660 8840
rect 620 8805 625 8835
rect 625 8805 655 8835
rect 655 8805 660 8835
rect 620 8800 660 8805
rect 620 8770 660 8775
rect 620 8740 625 8770
rect 625 8740 655 8770
rect 655 8740 660 8770
rect 620 8735 660 8740
rect 620 8700 660 8705
rect 620 8670 625 8700
rect 625 8670 655 8700
rect 655 8670 660 8700
rect 620 8665 660 8670
rect 620 8630 660 8635
rect 620 8600 625 8630
rect 625 8600 655 8630
rect 655 8600 660 8630
rect 620 8595 660 8600
rect 620 8560 660 8565
rect 620 8530 625 8560
rect 625 8530 655 8560
rect 655 8530 660 8560
rect 620 8525 660 8530
rect 620 8495 660 8500
rect 620 8465 625 8495
rect 625 8465 655 8495
rect 655 8465 660 8495
rect 620 8460 660 8465
rect 620 8435 660 8440
rect 620 8405 625 8435
rect 625 8405 655 8435
rect 655 8405 660 8435
rect 620 8400 660 8405
rect 620 8370 660 8375
rect 620 8340 625 8370
rect 625 8340 655 8370
rect 655 8340 660 8370
rect 620 8335 660 8340
rect 620 8300 660 8305
rect 620 8270 625 8300
rect 625 8270 655 8300
rect 655 8270 660 8300
rect 620 8265 660 8270
rect 620 8230 660 8235
rect 620 8200 625 8230
rect 625 8200 655 8230
rect 655 8200 660 8230
rect 620 8195 660 8200
rect 620 8160 660 8165
rect 620 8130 625 8160
rect 625 8130 655 8160
rect 655 8130 660 8160
rect 620 8125 660 8130
rect 620 8095 660 8100
rect 620 8065 625 8095
rect 625 8065 655 8095
rect 655 8065 660 8095
rect 620 8060 660 8065
rect 620 8035 660 8040
rect 620 8005 625 8035
rect 625 8005 655 8035
rect 655 8005 660 8035
rect 620 8000 660 8005
rect 620 7970 660 7975
rect 620 7940 625 7970
rect 625 7940 655 7970
rect 655 7940 660 7970
rect 620 7935 660 7940
rect 620 7900 660 7905
rect 620 7870 625 7900
rect 625 7870 655 7900
rect 655 7870 660 7900
rect 620 7865 660 7870
rect 620 7830 660 7835
rect 620 7800 625 7830
rect 625 7800 655 7830
rect 655 7800 660 7830
rect 620 7795 660 7800
rect 620 7760 660 7765
rect 620 7730 625 7760
rect 625 7730 655 7760
rect 655 7730 660 7760
rect 620 7725 660 7730
rect 620 7695 660 7700
rect 620 7665 625 7695
rect 625 7665 655 7695
rect 655 7665 660 7695
rect 620 7660 660 7665
rect 620 7635 660 7640
rect 620 7605 625 7635
rect 625 7605 655 7635
rect 655 7605 660 7635
rect 620 7600 660 7605
rect 620 7570 660 7575
rect 620 7540 625 7570
rect 625 7540 655 7570
rect 655 7540 660 7570
rect 620 7535 660 7540
rect 620 7500 660 7505
rect 620 7470 625 7500
rect 625 7470 655 7500
rect 655 7470 660 7500
rect 620 7465 660 7470
rect 620 7430 660 7435
rect 620 7400 625 7430
rect 625 7400 655 7430
rect 655 7400 660 7430
rect 620 7395 660 7400
rect 620 7360 660 7365
rect 620 7330 625 7360
rect 625 7330 655 7360
rect 655 7330 660 7360
rect 620 7325 660 7330
rect 620 7295 660 7300
rect 620 7265 625 7295
rect 625 7265 655 7295
rect 655 7265 660 7295
rect 620 7260 660 7265
rect 620 7235 660 7240
rect 620 7205 625 7235
rect 625 7205 655 7235
rect 655 7205 660 7235
rect 620 7200 660 7205
rect 620 7170 660 7175
rect 620 7140 625 7170
rect 625 7140 655 7170
rect 655 7140 660 7170
rect 620 7135 660 7140
rect 620 7100 660 7105
rect 620 7070 625 7100
rect 625 7070 655 7100
rect 655 7070 660 7100
rect 620 7065 660 7070
rect 620 7030 660 7035
rect 620 7000 625 7030
rect 625 7000 655 7030
rect 655 7000 660 7030
rect 620 6995 660 7000
rect 620 6960 660 6965
rect 620 6930 625 6960
rect 625 6930 655 6960
rect 655 6930 660 6960
rect 620 6925 660 6930
rect 620 6895 660 6900
rect 620 6865 625 6895
rect 625 6865 655 6895
rect 655 6865 660 6895
rect 620 6860 660 6865
rect 620 6835 660 6840
rect 620 6805 625 6835
rect 625 6805 655 6835
rect 655 6805 660 6835
rect 620 6800 660 6805
rect 620 6770 660 6775
rect 620 6740 625 6770
rect 625 6740 655 6770
rect 655 6740 660 6770
rect 620 6735 660 6740
rect 620 6700 660 6705
rect 620 6670 625 6700
rect 625 6670 655 6700
rect 655 6670 660 6700
rect 620 6665 660 6670
rect 620 6630 660 6635
rect 620 6600 625 6630
rect 625 6600 655 6630
rect 655 6600 660 6630
rect 620 6595 660 6600
rect 620 6560 660 6565
rect 620 6530 625 6560
rect 625 6530 655 6560
rect 655 6530 660 6560
rect 620 6525 660 6530
rect 620 6495 660 6500
rect 620 6465 625 6495
rect 625 6465 655 6495
rect 655 6465 660 6495
rect 620 6460 660 6465
rect 970 9635 1010 9640
rect 970 9605 975 9635
rect 975 9605 1005 9635
rect 1005 9605 1010 9635
rect 970 9600 1010 9605
rect 970 9570 1010 9575
rect 970 9540 975 9570
rect 975 9540 1005 9570
rect 1005 9540 1010 9570
rect 970 9535 1010 9540
rect 970 9500 1010 9505
rect 970 9470 975 9500
rect 975 9470 1005 9500
rect 1005 9470 1010 9500
rect 970 9465 1010 9470
rect 970 9430 1010 9435
rect 970 9400 975 9430
rect 975 9400 1005 9430
rect 1005 9400 1010 9430
rect 970 9395 1010 9400
rect 970 9360 1010 9365
rect 970 9330 975 9360
rect 975 9330 1005 9360
rect 1005 9330 1010 9360
rect 970 9325 1010 9330
rect 970 9295 1010 9300
rect 970 9265 975 9295
rect 975 9265 1005 9295
rect 1005 9265 1010 9295
rect 970 9260 1010 9265
rect 970 9235 1010 9240
rect 970 9205 975 9235
rect 975 9205 1005 9235
rect 1005 9205 1010 9235
rect 970 9200 1010 9205
rect 970 9170 1010 9175
rect 970 9140 975 9170
rect 975 9140 1005 9170
rect 1005 9140 1010 9170
rect 970 9135 1010 9140
rect 970 9100 1010 9105
rect 970 9070 975 9100
rect 975 9070 1005 9100
rect 1005 9070 1010 9100
rect 970 9065 1010 9070
rect 970 9030 1010 9035
rect 970 9000 975 9030
rect 975 9000 1005 9030
rect 1005 9000 1010 9030
rect 970 8995 1010 9000
rect 970 8960 1010 8965
rect 970 8930 975 8960
rect 975 8930 1005 8960
rect 1005 8930 1010 8960
rect 970 8925 1010 8930
rect 970 8895 1010 8900
rect 970 8865 975 8895
rect 975 8865 1005 8895
rect 1005 8865 1010 8895
rect 970 8860 1010 8865
rect 970 8835 1010 8840
rect 970 8805 975 8835
rect 975 8805 1005 8835
rect 1005 8805 1010 8835
rect 970 8800 1010 8805
rect 970 8770 1010 8775
rect 970 8740 975 8770
rect 975 8740 1005 8770
rect 1005 8740 1010 8770
rect 970 8735 1010 8740
rect 970 8700 1010 8705
rect 970 8670 975 8700
rect 975 8670 1005 8700
rect 1005 8670 1010 8700
rect 970 8665 1010 8670
rect 970 8630 1010 8635
rect 970 8600 975 8630
rect 975 8600 1005 8630
rect 1005 8600 1010 8630
rect 970 8595 1010 8600
rect 970 8560 1010 8565
rect 970 8530 975 8560
rect 975 8530 1005 8560
rect 1005 8530 1010 8560
rect 970 8525 1010 8530
rect 970 8495 1010 8500
rect 970 8465 975 8495
rect 975 8465 1005 8495
rect 1005 8465 1010 8495
rect 970 8460 1010 8465
rect 970 8435 1010 8440
rect 970 8405 975 8435
rect 975 8405 1005 8435
rect 1005 8405 1010 8435
rect 970 8400 1010 8405
rect 970 8370 1010 8375
rect 970 8340 975 8370
rect 975 8340 1005 8370
rect 1005 8340 1010 8370
rect 970 8335 1010 8340
rect 970 8300 1010 8305
rect 970 8270 975 8300
rect 975 8270 1005 8300
rect 1005 8270 1010 8300
rect 970 8265 1010 8270
rect 970 8230 1010 8235
rect 970 8200 975 8230
rect 975 8200 1005 8230
rect 1005 8200 1010 8230
rect 970 8195 1010 8200
rect 970 8160 1010 8165
rect 970 8130 975 8160
rect 975 8130 1005 8160
rect 1005 8130 1010 8160
rect 970 8125 1010 8130
rect 970 8095 1010 8100
rect 970 8065 975 8095
rect 975 8065 1005 8095
rect 1005 8065 1010 8095
rect 970 8060 1010 8065
rect 970 8035 1010 8040
rect 970 8005 975 8035
rect 975 8005 1005 8035
rect 1005 8005 1010 8035
rect 970 8000 1010 8005
rect 970 7970 1010 7975
rect 970 7940 975 7970
rect 975 7940 1005 7970
rect 1005 7940 1010 7970
rect 970 7935 1010 7940
rect 970 7900 1010 7905
rect 970 7870 975 7900
rect 975 7870 1005 7900
rect 1005 7870 1010 7900
rect 970 7865 1010 7870
rect 970 7830 1010 7835
rect 970 7800 975 7830
rect 975 7800 1005 7830
rect 1005 7800 1010 7830
rect 970 7795 1010 7800
rect 970 7760 1010 7765
rect 970 7730 975 7760
rect 975 7730 1005 7760
rect 1005 7730 1010 7760
rect 970 7725 1010 7730
rect 970 7695 1010 7700
rect 970 7665 975 7695
rect 975 7665 1005 7695
rect 1005 7665 1010 7695
rect 970 7660 1010 7665
rect 970 7635 1010 7640
rect 970 7605 975 7635
rect 975 7605 1005 7635
rect 1005 7605 1010 7635
rect 970 7600 1010 7605
rect 970 7570 1010 7575
rect 970 7540 975 7570
rect 975 7540 1005 7570
rect 1005 7540 1010 7570
rect 970 7535 1010 7540
rect 970 7500 1010 7505
rect 970 7470 975 7500
rect 975 7470 1005 7500
rect 1005 7470 1010 7500
rect 970 7465 1010 7470
rect 970 7430 1010 7435
rect 970 7400 975 7430
rect 975 7400 1005 7430
rect 1005 7400 1010 7430
rect 970 7395 1010 7400
rect 970 7360 1010 7365
rect 970 7330 975 7360
rect 975 7330 1005 7360
rect 1005 7330 1010 7360
rect 970 7325 1010 7330
rect 970 7295 1010 7300
rect 970 7265 975 7295
rect 975 7265 1005 7295
rect 1005 7265 1010 7295
rect 970 7260 1010 7265
rect 970 7235 1010 7240
rect 970 7205 975 7235
rect 975 7205 1005 7235
rect 1005 7205 1010 7235
rect 970 7200 1010 7205
rect 970 7170 1010 7175
rect 970 7140 975 7170
rect 975 7140 1005 7170
rect 1005 7140 1010 7170
rect 970 7135 1010 7140
rect 970 7100 1010 7105
rect 970 7070 975 7100
rect 975 7070 1005 7100
rect 1005 7070 1010 7100
rect 970 7065 1010 7070
rect 970 7030 1010 7035
rect 970 7000 975 7030
rect 975 7000 1005 7030
rect 1005 7000 1010 7030
rect 970 6995 1010 7000
rect 970 6960 1010 6965
rect 970 6930 975 6960
rect 975 6930 1005 6960
rect 1005 6930 1010 6960
rect 970 6925 1010 6930
rect 970 6895 1010 6900
rect 970 6865 975 6895
rect 975 6865 1005 6895
rect 1005 6865 1010 6895
rect 970 6860 1010 6865
rect 970 6835 1010 6840
rect 970 6805 975 6835
rect 975 6805 1005 6835
rect 1005 6805 1010 6835
rect 970 6800 1010 6805
rect 970 6770 1010 6775
rect 970 6740 975 6770
rect 975 6740 1005 6770
rect 1005 6740 1010 6770
rect 970 6735 1010 6740
rect 970 6700 1010 6705
rect 970 6670 975 6700
rect 975 6670 1005 6700
rect 1005 6670 1010 6700
rect 970 6665 1010 6670
rect 970 6630 1010 6635
rect 970 6600 975 6630
rect 975 6600 1005 6630
rect 1005 6600 1010 6630
rect 970 6595 1010 6600
rect 970 6560 1010 6565
rect 970 6530 975 6560
rect 975 6530 1005 6560
rect 1005 6530 1010 6560
rect 970 6525 1010 6530
rect 970 6495 1010 6500
rect 970 6465 975 6495
rect 975 6465 1005 6495
rect 1005 6465 1010 6495
rect 970 6460 1010 6465
rect 1670 9635 1710 9640
rect 1670 9605 1675 9635
rect 1675 9605 1705 9635
rect 1705 9605 1710 9635
rect 1670 9600 1710 9605
rect 1670 9570 1710 9575
rect 1670 9540 1675 9570
rect 1675 9540 1705 9570
rect 1705 9540 1710 9570
rect 1670 9535 1710 9540
rect 1670 9500 1710 9505
rect 1670 9470 1675 9500
rect 1675 9470 1705 9500
rect 1705 9470 1710 9500
rect 1670 9465 1710 9470
rect 1670 9430 1710 9435
rect 1670 9400 1675 9430
rect 1675 9400 1705 9430
rect 1705 9400 1710 9430
rect 1670 9395 1710 9400
rect 1670 9360 1710 9365
rect 1670 9330 1675 9360
rect 1675 9330 1705 9360
rect 1705 9330 1710 9360
rect 1670 9325 1710 9330
rect 1670 9295 1710 9300
rect 1670 9265 1675 9295
rect 1675 9265 1705 9295
rect 1705 9265 1710 9295
rect 1670 9260 1710 9265
rect 1670 9235 1710 9240
rect 1670 9205 1675 9235
rect 1675 9205 1705 9235
rect 1705 9205 1710 9235
rect 1670 9200 1710 9205
rect 1670 9170 1710 9175
rect 1670 9140 1675 9170
rect 1675 9140 1705 9170
rect 1705 9140 1710 9170
rect 1670 9135 1710 9140
rect 1670 9100 1710 9105
rect 1670 9070 1675 9100
rect 1675 9070 1705 9100
rect 1705 9070 1710 9100
rect 1670 9065 1710 9070
rect 1670 9030 1710 9035
rect 1670 9000 1675 9030
rect 1675 9000 1705 9030
rect 1705 9000 1710 9030
rect 1670 8995 1710 9000
rect 1670 8960 1710 8965
rect 1670 8930 1675 8960
rect 1675 8930 1705 8960
rect 1705 8930 1710 8960
rect 1670 8925 1710 8930
rect 1670 8895 1710 8900
rect 1670 8865 1675 8895
rect 1675 8865 1705 8895
rect 1705 8865 1710 8895
rect 1670 8860 1710 8865
rect 1670 8835 1710 8840
rect 1670 8805 1675 8835
rect 1675 8805 1705 8835
rect 1705 8805 1710 8835
rect 1670 8800 1710 8805
rect 1670 8770 1710 8775
rect 1670 8740 1675 8770
rect 1675 8740 1705 8770
rect 1705 8740 1710 8770
rect 1670 8735 1710 8740
rect 1670 8700 1710 8705
rect 1670 8670 1675 8700
rect 1675 8670 1705 8700
rect 1705 8670 1710 8700
rect 1670 8665 1710 8670
rect 1670 8630 1710 8635
rect 1670 8600 1675 8630
rect 1675 8600 1705 8630
rect 1705 8600 1710 8630
rect 1670 8595 1710 8600
rect 1670 8560 1710 8565
rect 1670 8530 1675 8560
rect 1675 8530 1705 8560
rect 1705 8530 1710 8560
rect 1670 8525 1710 8530
rect 1670 8495 1710 8500
rect 1670 8465 1675 8495
rect 1675 8465 1705 8495
rect 1705 8465 1710 8495
rect 1670 8460 1710 8465
rect 1670 8435 1710 8440
rect 1670 8405 1675 8435
rect 1675 8405 1705 8435
rect 1705 8405 1710 8435
rect 1670 8400 1710 8405
rect 1670 8370 1710 8375
rect 1670 8340 1675 8370
rect 1675 8340 1705 8370
rect 1705 8340 1710 8370
rect 1670 8335 1710 8340
rect 1670 8300 1710 8305
rect 1670 8270 1675 8300
rect 1675 8270 1705 8300
rect 1705 8270 1710 8300
rect 1670 8265 1710 8270
rect 1670 8230 1710 8235
rect 1670 8200 1675 8230
rect 1675 8200 1705 8230
rect 1705 8200 1710 8230
rect 1670 8195 1710 8200
rect 1670 8160 1710 8165
rect 1670 8130 1675 8160
rect 1675 8130 1705 8160
rect 1705 8130 1710 8160
rect 1670 8125 1710 8130
rect 1670 8095 1710 8100
rect 1670 8065 1675 8095
rect 1675 8065 1705 8095
rect 1705 8065 1710 8095
rect 1670 8060 1710 8065
rect 1670 8035 1710 8040
rect 1670 8005 1675 8035
rect 1675 8005 1705 8035
rect 1705 8005 1710 8035
rect 1670 8000 1710 8005
rect 1670 7970 1710 7975
rect 1670 7940 1675 7970
rect 1675 7940 1705 7970
rect 1705 7940 1710 7970
rect 1670 7935 1710 7940
rect 1670 7900 1710 7905
rect 1670 7870 1675 7900
rect 1675 7870 1705 7900
rect 1705 7870 1710 7900
rect 1670 7865 1710 7870
rect 1670 7830 1710 7835
rect 1670 7800 1675 7830
rect 1675 7800 1705 7830
rect 1705 7800 1710 7830
rect 1670 7795 1710 7800
rect 1670 7760 1710 7765
rect 1670 7730 1675 7760
rect 1675 7730 1705 7760
rect 1705 7730 1710 7760
rect 1670 7725 1710 7730
rect 1670 7695 1710 7700
rect 1670 7665 1675 7695
rect 1675 7665 1705 7695
rect 1705 7665 1710 7695
rect 1670 7660 1710 7665
rect 1670 7635 1710 7640
rect 1670 7605 1675 7635
rect 1675 7605 1705 7635
rect 1705 7605 1710 7635
rect 1670 7600 1710 7605
rect 1670 7570 1710 7575
rect 1670 7540 1675 7570
rect 1675 7540 1705 7570
rect 1705 7540 1710 7570
rect 1670 7535 1710 7540
rect 1670 7500 1710 7505
rect 1670 7470 1675 7500
rect 1675 7470 1705 7500
rect 1705 7470 1710 7500
rect 1670 7465 1710 7470
rect 1670 7430 1710 7435
rect 1670 7400 1675 7430
rect 1675 7400 1705 7430
rect 1705 7400 1710 7430
rect 1670 7395 1710 7400
rect 1670 7360 1710 7365
rect 1670 7330 1675 7360
rect 1675 7330 1705 7360
rect 1705 7330 1710 7360
rect 1670 7325 1710 7330
rect 1670 7295 1710 7300
rect 1670 7265 1675 7295
rect 1675 7265 1705 7295
rect 1705 7265 1710 7295
rect 1670 7260 1710 7265
rect 1670 7235 1710 7240
rect 1670 7205 1675 7235
rect 1675 7205 1705 7235
rect 1705 7205 1710 7235
rect 1670 7200 1710 7205
rect 1670 7170 1710 7175
rect 1670 7140 1675 7170
rect 1675 7140 1705 7170
rect 1705 7140 1710 7170
rect 1670 7135 1710 7140
rect 1670 7100 1710 7105
rect 1670 7070 1675 7100
rect 1675 7070 1705 7100
rect 1705 7070 1710 7100
rect 1670 7065 1710 7070
rect 1670 7030 1710 7035
rect 1670 7000 1675 7030
rect 1675 7000 1705 7030
rect 1705 7000 1710 7030
rect 1670 6995 1710 7000
rect 1670 6960 1710 6965
rect 1670 6930 1675 6960
rect 1675 6930 1705 6960
rect 1705 6930 1710 6960
rect 1670 6925 1710 6930
rect 1670 6895 1710 6900
rect 1670 6865 1675 6895
rect 1675 6865 1705 6895
rect 1705 6865 1710 6895
rect 1670 6860 1710 6865
rect 1670 6835 1710 6840
rect 1670 6805 1675 6835
rect 1675 6805 1705 6835
rect 1705 6805 1710 6835
rect 1670 6800 1710 6805
rect 1670 6770 1710 6775
rect 1670 6740 1675 6770
rect 1675 6740 1705 6770
rect 1705 6740 1710 6770
rect 1670 6735 1710 6740
rect 1670 6700 1710 6705
rect 1670 6670 1675 6700
rect 1675 6670 1705 6700
rect 1705 6670 1710 6700
rect 1670 6665 1710 6670
rect 1670 6630 1710 6635
rect 1670 6600 1675 6630
rect 1675 6600 1705 6630
rect 1705 6600 1710 6630
rect 1670 6595 1710 6600
rect 1670 6560 1710 6565
rect 1670 6530 1675 6560
rect 1675 6530 1705 6560
rect 1705 6530 1710 6560
rect 1670 6525 1710 6530
rect 1670 6495 1710 6500
rect 1670 6465 1675 6495
rect 1675 6465 1705 6495
rect 1705 6465 1710 6495
rect 1670 6460 1710 6465
rect 2325 9635 2365 9640
rect 2325 9605 2330 9635
rect 2330 9605 2360 9635
rect 2360 9605 2365 9635
rect 2325 9600 2365 9605
rect 2325 9570 2365 9575
rect 2325 9540 2330 9570
rect 2330 9540 2360 9570
rect 2360 9540 2365 9570
rect 2325 9535 2365 9540
rect 2325 9500 2365 9505
rect 2325 9470 2330 9500
rect 2330 9470 2360 9500
rect 2360 9470 2365 9500
rect 2325 9465 2365 9470
rect 2325 9430 2365 9435
rect 2325 9400 2330 9430
rect 2330 9400 2360 9430
rect 2360 9400 2365 9430
rect 2325 9395 2365 9400
rect 2325 9360 2365 9365
rect 2325 9330 2330 9360
rect 2330 9330 2360 9360
rect 2360 9330 2365 9360
rect 2325 9325 2365 9330
rect 2325 9295 2365 9300
rect 2325 9265 2330 9295
rect 2330 9265 2360 9295
rect 2360 9265 2365 9295
rect 2325 9260 2365 9265
rect 2325 9235 2365 9240
rect 2325 9205 2330 9235
rect 2330 9205 2360 9235
rect 2360 9205 2365 9235
rect 2325 9200 2365 9205
rect 2325 9170 2365 9175
rect 2325 9140 2330 9170
rect 2330 9140 2360 9170
rect 2360 9140 2365 9170
rect 2325 9135 2365 9140
rect 2325 9100 2365 9105
rect 2325 9070 2330 9100
rect 2330 9070 2360 9100
rect 2360 9070 2365 9100
rect 2325 9065 2365 9070
rect 2325 9030 2365 9035
rect 2325 9000 2330 9030
rect 2330 9000 2360 9030
rect 2360 9000 2365 9030
rect 2325 8995 2365 9000
rect 2325 8960 2365 8965
rect 2325 8930 2330 8960
rect 2330 8930 2360 8960
rect 2360 8930 2365 8960
rect 2325 8925 2365 8930
rect 2325 8895 2365 8900
rect 2325 8865 2330 8895
rect 2330 8865 2360 8895
rect 2360 8865 2365 8895
rect 2325 8860 2365 8865
rect 2325 8835 2365 8840
rect 2325 8805 2330 8835
rect 2330 8805 2360 8835
rect 2360 8805 2365 8835
rect 2325 8800 2365 8805
rect 2325 8770 2365 8775
rect 2325 8740 2330 8770
rect 2330 8740 2360 8770
rect 2360 8740 2365 8770
rect 2325 8735 2365 8740
rect 2325 8700 2365 8705
rect 2325 8670 2330 8700
rect 2330 8670 2360 8700
rect 2360 8670 2365 8700
rect 2325 8665 2365 8670
rect 2325 8630 2365 8635
rect 2325 8600 2330 8630
rect 2330 8600 2360 8630
rect 2360 8600 2365 8630
rect 2325 8595 2365 8600
rect 2325 8560 2365 8565
rect 2325 8530 2330 8560
rect 2330 8530 2360 8560
rect 2360 8530 2365 8560
rect 2325 8525 2365 8530
rect 2325 8495 2365 8500
rect 2325 8465 2330 8495
rect 2330 8465 2360 8495
rect 2360 8465 2365 8495
rect 2325 8460 2365 8465
rect 2325 8435 2365 8440
rect 2325 8405 2330 8435
rect 2330 8405 2360 8435
rect 2360 8405 2365 8435
rect 2325 8400 2365 8405
rect 2325 8370 2365 8375
rect 2325 8340 2330 8370
rect 2330 8340 2360 8370
rect 2360 8340 2365 8370
rect 2325 8335 2365 8340
rect 2325 8300 2365 8305
rect 2325 8270 2330 8300
rect 2330 8270 2360 8300
rect 2360 8270 2365 8300
rect 2325 8265 2365 8270
rect 2325 8230 2365 8235
rect 2325 8200 2330 8230
rect 2330 8200 2360 8230
rect 2360 8200 2365 8230
rect 2325 8195 2365 8200
rect 2325 8160 2365 8165
rect 2325 8130 2330 8160
rect 2330 8130 2360 8160
rect 2360 8130 2365 8160
rect 2325 8125 2365 8130
rect 2325 8095 2365 8100
rect 2325 8065 2330 8095
rect 2330 8065 2360 8095
rect 2360 8065 2365 8095
rect 2325 8060 2365 8065
rect 2325 8035 2365 8040
rect 2325 8005 2330 8035
rect 2330 8005 2360 8035
rect 2360 8005 2365 8035
rect 2325 8000 2365 8005
rect 2325 7970 2365 7975
rect 2325 7940 2330 7970
rect 2330 7940 2360 7970
rect 2360 7940 2365 7970
rect 2325 7935 2365 7940
rect 2325 7900 2365 7905
rect 2325 7870 2330 7900
rect 2330 7870 2360 7900
rect 2360 7870 2365 7900
rect 2325 7865 2365 7870
rect 2325 7830 2365 7835
rect 2325 7800 2330 7830
rect 2330 7800 2360 7830
rect 2360 7800 2365 7830
rect 2325 7795 2365 7800
rect 2325 7760 2365 7765
rect 2325 7730 2330 7760
rect 2330 7730 2360 7760
rect 2360 7730 2365 7760
rect 2325 7725 2365 7730
rect 2325 7695 2365 7700
rect 2325 7665 2330 7695
rect 2330 7665 2360 7695
rect 2360 7665 2365 7695
rect 2325 7660 2365 7665
rect 2325 7635 2365 7640
rect 2325 7605 2330 7635
rect 2330 7605 2360 7635
rect 2360 7605 2365 7635
rect 2325 7600 2365 7605
rect 2325 7570 2365 7575
rect 2325 7540 2330 7570
rect 2330 7540 2360 7570
rect 2360 7540 2365 7570
rect 2325 7535 2365 7540
rect 2325 7500 2365 7505
rect 2325 7470 2330 7500
rect 2330 7470 2360 7500
rect 2360 7470 2365 7500
rect 2325 7465 2365 7470
rect 2325 7430 2365 7435
rect 2325 7400 2330 7430
rect 2330 7400 2360 7430
rect 2360 7400 2365 7430
rect 2325 7395 2365 7400
rect 2325 7360 2365 7365
rect 2325 7330 2330 7360
rect 2330 7330 2360 7360
rect 2360 7330 2365 7360
rect 2325 7325 2365 7330
rect 2325 7295 2365 7300
rect 2325 7265 2330 7295
rect 2330 7265 2360 7295
rect 2360 7265 2365 7295
rect 2325 7260 2365 7265
rect 2325 7235 2365 7240
rect 2325 7205 2330 7235
rect 2330 7205 2360 7235
rect 2360 7205 2365 7235
rect 2325 7200 2365 7205
rect 2325 7170 2365 7175
rect 2325 7140 2330 7170
rect 2330 7140 2360 7170
rect 2360 7140 2365 7170
rect 2325 7135 2365 7140
rect 2325 7100 2365 7105
rect 2325 7070 2330 7100
rect 2330 7070 2360 7100
rect 2360 7070 2365 7100
rect 2325 7065 2365 7070
rect 2325 7030 2365 7035
rect 2325 7000 2330 7030
rect 2330 7000 2360 7030
rect 2360 7000 2365 7030
rect 2325 6995 2365 7000
rect 2325 6960 2365 6965
rect 2325 6930 2330 6960
rect 2330 6930 2360 6960
rect 2360 6930 2365 6960
rect 2325 6925 2365 6930
rect 2325 6895 2365 6900
rect 2325 6865 2330 6895
rect 2330 6865 2360 6895
rect 2360 6865 2365 6895
rect 2325 6860 2365 6865
rect 2325 6835 2365 6840
rect 2325 6805 2330 6835
rect 2330 6805 2360 6835
rect 2360 6805 2365 6835
rect 2325 6800 2365 6805
rect 2325 6770 2365 6775
rect 2325 6740 2330 6770
rect 2330 6740 2360 6770
rect 2360 6740 2365 6770
rect 2325 6735 2365 6740
rect 2325 6700 2365 6705
rect 2325 6670 2330 6700
rect 2330 6670 2360 6700
rect 2360 6670 2365 6700
rect 2325 6665 2365 6670
rect 2325 6630 2365 6635
rect 2325 6600 2330 6630
rect 2330 6600 2360 6630
rect 2360 6600 2365 6630
rect 2325 6595 2365 6600
rect 2325 6560 2365 6565
rect 2325 6530 2330 6560
rect 2330 6530 2360 6560
rect 2360 6530 2365 6560
rect 2325 6525 2365 6530
rect 2325 6495 2365 6500
rect 2325 6465 2330 6495
rect 2330 6465 2360 6495
rect 2360 6465 2365 6495
rect 2325 6460 2365 6465
rect 3175 9635 3215 9640
rect 3175 9605 3180 9635
rect 3180 9605 3210 9635
rect 3210 9605 3215 9635
rect 3175 9600 3215 9605
rect 3235 9635 3275 9640
rect 3235 9605 3240 9635
rect 3240 9605 3270 9635
rect 3270 9605 3275 9635
rect 3235 9600 3275 9605
rect 3175 9570 3215 9575
rect 3175 9540 3180 9570
rect 3180 9540 3210 9570
rect 3210 9540 3215 9570
rect 3175 9535 3215 9540
rect 3235 9570 3275 9575
rect 3235 9540 3240 9570
rect 3240 9540 3270 9570
rect 3270 9540 3275 9570
rect 3235 9535 3275 9540
rect 3175 9500 3215 9505
rect 3175 9470 3180 9500
rect 3180 9470 3210 9500
rect 3210 9470 3215 9500
rect 3175 9465 3215 9470
rect 3235 9500 3275 9505
rect 3235 9470 3240 9500
rect 3240 9470 3270 9500
rect 3270 9470 3275 9500
rect 3235 9465 3275 9470
rect 3175 9430 3215 9435
rect 3175 9400 3180 9430
rect 3180 9400 3210 9430
rect 3210 9400 3215 9430
rect 3175 9395 3215 9400
rect 3235 9430 3275 9435
rect 3235 9400 3240 9430
rect 3240 9400 3270 9430
rect 3270 9400 3275 9430
rect 3235 9395 3275 9400
rect 3175 9360 3215 9365
rect 3175 9330 3180 9360
rect 3180 9330 3210 9360
rect 3210 9330 3215 9360
rect 3175 9325 3215 9330
rect 3235 9360 3275 9365
rect 3235 9330 3240 9360
rect 3240 9330 3270 9360
rect 3270 9330 3275 9360
rect 3235 9325 3275 9330
rect 3175 9295 3215 9300
rect 3175 9265 3180 9295
rect 3180 9265 3210 9295
rect 3210 9265 3215 9295
rect 3175 9260 3215 9265
rect 3235 9295 3275 9300
rect 3235 9265 3240 9295
rect 3240 9265 3270 9295
rect 3270 9265 3275 9295
rect 3235 9260 3275 9265
rect 3175 9235 3215 9240
rect 3175 9205 3180 9235
rect 3180 9205 3210 9235
rect 3210 9205 3215 9235
rect 3175 9200 3215 9205
rect 3235 9235 3275 9240
rect 3235 9205 3240 9235
rect 3240 9205 3270 9235
rect 3270 9205 3275 9235
rect 3235 9200 3275 9205
rect 3175 9170 3215 9175
rect 3175 9140 3180 9170
rect 3180 9140 3210 9170
rect 3210 9140 3215 9170
rect 3175 9135 3215 9140
rect 3235 9170 3275 9175
rect 3235 9140 3240 9170
rect 3240 9140 3270 9170
rect 3270 9140 3275 9170
rect 3235 9135 3275 9140
rect 3175 9100 3215 9105
rect 3175 9070 3180 9100
rect 3180 9070 3210 9100
rect 3210 9070 3215 9100
rect 3175 9065 3215 9070
rect 3235 9100 3275 9105
rect 3235 9070 3240 9100
rect 3240 9070 3270 9100
rect 3270 9070 3275 9100
rect 3235 9065 3275 9070
rect 3175 9030 3215 9035
rect 3175 9000 3180 9030
rect 3180 9000 3210 9030
rect 3210 9000 3215 9030
rect 3175 8995 3215 9000
rect 3235 9030 3275 9035
rect 3235 9000 3240 9030
rect 3240 9000 3270 9030
rect 3270 9000 3275 9030
rect 3235 8995 3275 9000
rect 3175 8960 3215 8965
rect 3175 8930 3180 8960
rect 3180 8930 3210 8960
rect 3210 8930 3215 8960
rect 3175 8925 3215 8930
rect 3235 8960 3275 8965
rect 3235 8930 3240 8960
rect 3240 8930 3270 8960
rect 3270 8930 3275 8960
rect 3235 8925 3275 8930
rect 3175 8895 3215 8900
rect 3175 8865 3180 8895
rect 3180 8865 3210 8895
rect 3210 8865 3215 8895
rect 3175 8860 3215 8865
rect 3235 8895 3275 8900
rect 3235 8865 3240 8895
rect 3240 8865 3270 8895
rect 3270 8865 3275 8895
rect 3235 8860 3275 8865
rect 3175 8835 3215 8840
rect 3175 8805 3180 8835
rect 3180 8805 3210 8835
rect 3210 8805 3215 8835
rect 3175 8800 3215 8805
rect 3235 8835 3275 8840
rect 3235 8805 3240 8835
rect 3240 8805 3270 8835
rect 3270 8805 3275 8835
rect 3235 8800 3275 8805
rect 3175 8770 3215 8775
rect 3175 8740 3180 8770
rect 3180 8740 3210 8770
rect 3210 8740 3215 8770
rect 3175 8735 3215 8740
rect 3235 8770 3275 8775
rect 3235 8740 3240 8770
rect 3240 8740 3270 8770
rect 3270 8740 3275 8770
rect 3235 8735 3275 8740
rect 3175 8700 3215 8705
rect 3175 8670 3180 8700
rect 3180 8670 3210 8700
rect 3210 8670 3215 8700
rect 3175 8665 3215 8670
rect 3235 8700 3275 8705
rect 3235 8670 3240 8700
rect 3240 8670 3270 8700
rect 3270 8670 3275 8700
rect 3235 8665 3275 8670
rect 3175 8630 3215 8635
rect 3175 8600 3180 8630
rect 3180 8600 3210 8630
rect 3210 8600 3215 8630
rect 3175 8595 3215 8600
rect 3235 8630 3275 8635
rect 3235 8600 3240 8630
rect 3240 8600 3270 8630
rect 3270 8600 3275 8630
rect 3235 8595 3275 8600
rect 3175 8560 3215 8565
rect 3175 8530 3180 8560
rect 3180 8530 3210 8560
rect 3210 8530 3215 8560
rect 3175 8525 3215 8530
rect 3235 8560 3275 8565
rect 3235 8530 3240 8560
rect 3240 8530 3270 8560
rect 3270 8530 3275 8560
rect 3235 8525 3275 8530
rect 3175 8495 3215 8500
rect 3175 8465 3180 8495
rect 3180 8465 3210 8495
rect 3210 8465 3215 8495
rect 3175 8460 3215 8465
rect 3235 8495 3275 8500
rect 3235 8465 3240 8495
rect 3240 8465 3270 8495
rect 3270 8465 3275 8495
rect 3235 8460 3275 8465
rect 3175 8435 3215 8440
rect 3175 8405 3180 8435
rect 3180 8405 3210 8435
rect 3210 8405 3215 8435
rect 3175 8400 3215 8405
rect 3235 8435 3275 8440
rect 3235 8405 3240 8435
rect 3240 8405 3270 8435
rect 3270 8405 3275 8435
rect 3235 8400 3275 8405
rect 3175 8370 3215 8375
rect 3175 8340 3180 8370
rect 3180 8340 3210 8370
rect 3210 8340 3215 8370
rect 3175 8335 3215 8340
rect 3235 8370 3275 8375
rect 3235 8340 3240 8370
rect 3240 8340 3270 8370
rect 3270 8340 3275 8370
rect 3235 8335 3275 8340
rect 3175 8300 3215 8305
rect 3175 8270 3180 8300
rect 3180 8270 3210 8300
rect 3210 8270 3215 8300
rect 3175 8265 3215 8270
rect 3235 8300 3275 8305
rect 3235 8270 3240 8300
rect 3240 8270 3270 8300
rect 3270 8270 3275 8300
rect 3235 8265 3275 8270
rect 3175 8230 3215 8235
rect 3175 8200 3180 8230
rect 3180 8200 3210 8230
rect 3210 8200 3215 8230
rect 3175 8195 3215 8200
rect 3235 8230 3275 8235
rect 3235 8200 3240 8230
rect 3240 8200 3270 8230
rect 3270 8200 3275 8230
rect 3235 8195 3275 8200
rect 3175 8160 3215 8165
rect 3175 8130 3180 8160
rect 3180 8130 3210 8160
rect 3210 8130 3215 8160
rect 3175 8125 3215 8130
rect 3235 8160 3275 8165
rect 3235 8130 3240 8160
rect 3240 8130 3270 8160
rect 3270 8130 3275 8160
rect 3235 8125 3275 8130
rect 3175 8095 3215 8100
rect 3175 8065 3180 8095
rect 3180 8065 3210 8095
rect 3210 8065 3215 8095
rect 3175 8060 3215 8065
rect 3235 8095 3275 8100
rect 3235 8065 3240 8095
rect 3240 8065 3270 8095
rect 3270 8065 3275 8095
rect 3235 8060 3275 8065
rect 3175 8035 3215 8040
rect 3175 8005 3180 8035
rect 3180 8005 3210 8035
rect 3210 8005 3215 8035
rect 3175 8000 3215 8005
rect 3235 8035 3275 8040
rect 3235 8005 3240 8035
rect 3240 8005 3270 8035
rect 3270 8005 3275 8035
rect 3235 8000 3275 8005
rect 3175 7970 3215 7975
rect 3175 7940 3180 7970
rect 3180 7940 3210 7970
rect 3210 7940 3215 7970
rect 3175 7935 3215 7940
rect 3235 7970 3275 7975
rect 3235 7940 3240 7970
rect 3240 7940 3270 7970
rect 3270 7940 3275 7970
rect 3235 7935 3275 7940
rect 3175 7900 3215 7905
rect 3175 7870 3180 7900
rect 3180 7870 3210 7900
rect 3210 7870 3215 7900
rect 3175 7865 3215 7870
rect 3235 7900 3275 7905
rect 3235 7870 3240 7900
rect 3240 7870 3270 7900
rect 3270 7870 3275 7900
rect 3235 7865 3275 7870
rect 3175 7830 3215 7835
rect 3175 7800 3180 7830
rect 3180 7800 3210 7830
rect 3210 7800 3215 7830
rect 3175 7795 3215 7800
rect 3235 7830 3275 7835
rect 3235 7800 3240 7830
rect 3240 7800 3270 7830
rect 3270 7800 3275 7830
rect 3235 7795 3275 7800
rect 3175 7760 3215 7765
rect 3175 7730 3180 7760
rect 3180 7730 3210 7760
rect 3210 7730 3215 7760
rect 3175 7725 3215 7730
rect 3235 7760 3275 7765
rect 3235 7730 3240 7760
rect 3240 7730 3270 7760
rect 3270 7730 3275 7760
rect 3235 7725 3275 7730
rect 3175 7695 3215 7700
rect 3175 7665 3180 7695
rect 3180 7665 3210 7695
rect 3210 7665 3215 7695
rect 3175 7660 3215 7665
rect 3235 7695 3275 7700
rect 3235 7665 3240 7695
rect 3240 7665 3270 7695
rect 3270 7665 3275 7695
rect 3235 7660 3275 7665
rect 3175 7635 3215 7640
rect 3175 7605 3180 7635
rect 3180 7605 3210 7635
rect 3210 7605 3215 7635
rect 3175 7600 3215 7605
rect 3235 7635 3275 7640
rect 3235 7605 3240 7635
rect 3240 7605 3270 7635
rect 3270 7605 3275 7635
rect 3235 7600 3275 7605
rect 3175 7570 3215 7575
rect 3175 7540 3180 7570
rect 3180 7540 3210 7570
rect 3210 7540 3215 7570
rect 3175 7535 3215 7540
rect 3235 7570 3275 7575
rect 3235 7540 3240 7570
rect 3240 7540 3270 7570
rect 3270 7540 3275 7570
rect 3235 7535 3275 7540
rect 3175 7500 3215 7505
rect 3175 7470 3180 7500
rect 3180 7470 3210 7500
rect 3210 7470 3215 7500
rect 3175 7465 3215 7470
rect 3235 7500 3275 7505
rect 3235 7470 3240 7500
rect 3240 7470 3270 7500
rect 3270 7470 3275 7500
rect 3235 7465 3275 7470
rect 3175 7430 3215 7435
rect 3175 7400 3180 7430
rect 3180 7400 3210 7430
rect 3210 7400 3215 7430
rect 3175 7395 3215 7400
rect 3235 7430 3275 7435
rect 3235 7400 3240 7430
rect 3240 7400 3270 7430
rect 3270 7400 3275 7430
rect 3235 7395 3275 7400
rect 3175 7360 3215 7365
rect 3175 7330 3180 7360
rect 3180 7330 3210 7360
rect 3210 7330 3215 7360
rect 3175 7325 3215 7330
rect 3235 7360 3275 7365
rect 3235 7330 3240 7360
rect 3240 7330 3270 7360
rect 3270 7330 3275 7360
rect 3235 7325 3275 7330
rect 3175 7295 3215 7300
rect 3175 7265 3180 7295
rect 3180 7265 3210 7295
rect 3210 7265 3215 7295
rect 3175 7260 3215 7265
rect 3235 7295 3275 7300
rect 3235 7265 3240 7295
rect 3240 7265 3270 7295
rect 3270 7265 3275 7295
rect 3235 7260 3275 7265
rect 3175 7235 3215 7240
rect 3175 7205 3180 7235
rect 3180 7205 3210 7235
rect 3210 7205 3215 7235
rect 3175 7200 3215 7205
rect 3235 7235 3275 7240
rect 3235 7205 3240 7235
rect 3240 7205 3270 7235
rect 3270 7205 3275 7235
rect 3235 7200 3275 7205
rect 3175 7170 3215 7175
rect 3175 7140 3180 7170
rect 3180 7140 3210 7170
rect 3210 7140 3215 7170
rect 3175 7135 3215 7140
rect 3235 7170 3275 7175
rect 3235 7140 3240 7170
rect 3240 7140 3270 7170
rect 3270 7140 3275 7170
rect 3235 7135 3275 7140
rect 3175 7100 3215 7105
rect 3175 7070 3180 7100
rect 3180 7070 3210 7100
rect 3210 7070 3215 7100
rect 3175 7065 3215 7070
rect 3235 7100 3275 7105
rect 3235 7070 3240 7100
rect 3240 7070 3270 7100
rect 3270 7070 3275 7100
rect 3235 7065 3275 7070
rect 3175 7030 3215 7035
rect 3175 7000 3180 7030
rect 3180 7000 3210 7030
rect 3210 7000 3215 7030
rect 3175 6995 3215 7000
rect 3235 7030 3275 7035
rect 3235 7000 3240 7030
rect 3240 7000 3270 7030
rect 3270 7000 3275 7030
rect 3235 6995 3275 7000
rect 3175 6960 3215 6965
rect 3175 6930 3180 6960
rect 3180 6930 3210 6960
rect 3210 6930 3215 6960
rect 3175 6925 3215 6930
rect 3235 6960 3275 6965
rect 3235 6930 3240 6960
rect 3240 6930 3270 6960
rect 3270 6930 3275 6960
rect 3235 6925 3275 6930
rect 3175 6895 3215 6900
rect 3175 6865 3180 6895
rect 3180 6865 3210 6895
rect 3210 6865 3215 6895
rect 3175 6860 3215 6865
rect 3235 6895 3275 6900
rect 3235 6865 3240 6895
rect 3240 6865 3270 6895
rect 3270 6865 3275 6895
rect 3235 6860 3275 6865
rect 3175 6835 3215 6840
rect 3175 6805 3180 6835
rect 3180 6805 3210 6835
rect 3210 6805 3215 6835
rect 3175 6800 3215 6805
rect 3235 6835 3275 6840
rect 3235 6805 3240 6835
rect 3240 6805 3270 6835
rect 3270 6805 3275 6835
rect 3235 6800 3275 6805
rect 3175 6770 3215 6775
rect 3175 6740 3180 6770
rect 3180 6740 3210 6770
rect 3210 6740 3215 6770
rect 3175 6735 3215 6740
rect 3235 6770 3275 6775
rect 3235 6740 3240 6770
rect 3240 6740 3270 6770
rect 3270 6740 3275 6770
rect 3235 6735 3275 6740
rect 3175 6700 3215 6705
rect 3175 6670 3180 6700
rect 3180 6670 3210 6700
rect 3210 6670 3215 6700
rect 3175 6665 3215 6670
rect 3235 6700 3275 6705
rect 3235 6670 3240 6700
rect 3240 6670 3270 6700
rect 3270 6670 3275 6700
rect 3235 6665 3275 6670
rect 3175 6630 3215 6635
rect 3175 6600 3180 6630
rect 3180 6600 3210 6630
rect 3210 6600 3215 6630
rect 3175 6595 3215 6600
rect 3235 6630 3275 6635
rect 3235 6600 3240 6630
rect 3240 6600 3270 6630
rect 3270 6600 3275 6630
rect 3235 6595 3275 6600
rect 3175 6560 3215 6565
rect 3175 6530 3180 6560
rect 3180 6530 3210 6560
rect 3210 6530 3215 6560
rect 3175 6525 3215 6530
rect 3235 6560 3275 6565
rect 3235 6530 3240 6560
rect 3240 6530 3270 6560
rect 3270 6530 3275 6560
rect 3235 6525 3275 6530
rect 3175 6495 3215 6500
rect 3175 6465 3180 6495
rect 3180 6465 3210 6495
rect 3210 6465 3215 6495
rect 3175 6460 3215 6465
rect 3235 6495 3275 6500
rect 3235 6465 3240 6495
rect 3240 6465 3270 6495
rect 3270 6465 3275 6495
rect 3235 6460 3275 6465
rect 3345 9635 3385 9640
rect 3345 9605 3350 9635
rect 3350 9605 3380 9635
rect 3380 9605 3385 9635
rect 3345 9600 3385 9605
rect 3345 9570 3385 9575
rect 3345 9540 3350 9570
rect 3350 9540 3380 9570
rect 3380 9540 3385 9570
rect 3345 9535 3385 9540
rect 3345 9500 3385 9505
rect 3345 9470 3350 9500
rect 3350 9470 3380 9500
rect 3380 9470 3385 9500
rect 3345 9465 3385 9470
rect 3345 9430 3385 9435
rect 3345 9400 3350 9430
rect 3350 9400 3380 9430
rect 3380 9400 3385 9430
rect 3345 9395 3385 9400
rect 3345 9360 3385 9365
rect 3345 9330 3350 9360
rect 3350 9330 3380 9360
rect 3380 9330 3385 9360
rect 3345 9325 3385 9330
rect 3345 9295 3385 9300
rect 3345 9265 3350 9295
rect 3350 9265 3380 9295
rect 3380 9265 3385 9295
rect 3345 9260 3385 9265
rect 3345 9235 3385 9240
rect 3345 9205 3350 9235
rect 3350 9205 3380 9235
rect 3380 9205 3385 9235
rect 3345 9200 3385 9205
rect 3345 9170 3385 9175
rect 3345 9140 3350 9170
rect 3350 9140 3380 9170
rect 3380 9140 3385 9170
rect 3345 9135 3385 9140
rect 3345 9100 3385 9105
rect 3345 9070 3350 9100
rect 3350 9070 3380 9100
rect 3380 9070 3385 9100
rect 3345 9065 3385 9070
rect 3345 9030 3385 9035
rect 3345 9000 3350 9030
rect 3350 9000 3380 9030
rect 3380 9000 3385 9030
rect 3345 8995 3385 9000
rect 3345 8960 3385 8965
rect 3345 8930 3350 8960
rect 3350 8930 3380 8960
rect 3380 8930 3385 8960
rect 3345 8925 3385 8930
rect 3345 8895 3385 8900
rect 3345 8865 3350 8895
rect 3350 8865 3380 8895
rect 3380 8865 3385 8895
rect 3345 8860 3385 8865
rect 3345 8835 3385 8840
rect 3345 8805 3350 8835
rect 3350 8805 3380 8835
rect 3380 8805 3385 8835
rect 3345 8800 3385 8805
rect 3345 8770 3385 8775
rect 3345 8740 3350 8770
rect 3350 8740 3380 8770
rect 3380 8740 3385 8770
rect 3345 8735 3385 8740
rect 3345 8700 3385 8705
rect 3345 8670 3350 8700
rect 3350 8670 3380 8700
rect 3380 8670 3385 8700
rect 3345 8665 3385 8670
rect 3345 8630 3385 8635
rect 3345 8600 3350 8630
rect 3350 8600 3380 8630
rect 3380 8600 3385 8630
rect 3345 8595 3385 8600
rect 3345 8560 3385 8565
rect 3345 8530 3350 8560
rect 3350 8530 3380 8560
rect 3380 8530 3385 8560
rect 3345 8525 3385 8530
rect 3345 8495 3385 8500
rect 3345 8465 3350 8495
rect 3350 8465 3380 8495
rect 3380 8465 3385 8495
rect 3345 8460 3385 8465
rect 3345 8435 3385 8440
rect 3345 8405 3350 8435
rect 3350 8405 3380 8435
rect 3380 8405 3385 8435
rect 3345 8400 3385 8405
rect 3345 8370 3385 8375
rect 3345 8340 3350 8370
rect 3350 8340 3380 8370
rect 3380 8340 3385 8370
rect 3345 8335 3385 8340
rect 3345 8300 3385 8305
rect 3345 8270 3350 8300
rect 3350 8270 3380 8300
rect 3380 8270 3385 8300
rect 3345 8265 3385 8270
rect 3345 8230 3385 8235
rect 3345 8200 3350 8230
rect 3350 8200 3380 8230
rect 3380 8200 3385 8230
rect 3345 8195 3385 8200
rect 3345 8160 3385 8165
rect 3345 8130 3350 8160
rect 3350 8130 3380 8160
rect 3380 8130 3385 8160
rect 3345 8125 3385 8130
rect 3345 8095 3385 8100
rect 3345 8065 3350 8095
rect 3350 8065 3380 8095
rect 3380 8065 3385 8095
rect 3345 8060 3385 8065
rect 3345 8035 3385 8040
rect 3345 8005 3350 8035
rect 3350 8005 3380 8035
rect 3380 8005 3385 8035
rect 3345 8000 3385 8005
rect 3345 7970 3385 7975
rect 3345 7940 3350 7970
rect 3350 7940 3380 7970
rect 3380 7940 3385 7970
rect 3345 7935 3385 7940
rect 3345 7900 3385 7905
rect 3345 7870 3350 7900
rect 3350 7870 3380 7900
rect 3380 7870 3385 7900
rect 3345 7865 3385 7870
rect 3345 7830 3385 7835
rect 3345 7800 3350 7830
rect 3350 7800 3380 7830
rect 3380 7800 3385 7830
rect 3345 7795 3385 7800
rect 3345 7760 3385 7765
rect 3345 7730 3350 7760
rect 3350 7730 3380 7760
rect 3380 7730 3385 7760
rect 3345 7725 3385 7730
rect 3345 7695 3385 7700
rect 3345 7665 3350 7695
rect 3350 7665 3380 7695
rect 3380 7665 3385 7695
rect 3345 7660 3385 7665
rect 3345 7635 3385 7640
rect 3345 7605 3350 7635
rect 3350 7605 3380 7635
rect 3380 7605 3385 7635
rect 3345 7600 3385 7605
rect 3345 7570 3385 7575
rect 3345 7540 3350 7570
rect 3350 7540 3380 7570
rect 3380 7540 3385 7570
rect 3345 7535 3385 7540
rect 3345 7500 3385 7505
rect 3345 7470 3350 7500
rect 3350 7470 3380 7500
rect 3380 7470 3385 7500
rect 3345 7465 3385 7470
rect 3345 7430 3385 7435
rect 3345 7400 3350 7430
rect 3350 7400 3380 7430
rect 3380 7400 3385 7430
rect 3345 7395 3385 7400
rect 3345 7360 3385 7365
rect 3345 7330 3350 7360
rect 3350 7330 3380 7360
rect 3380 7330 3385 7360
rect 3345 7325 3385 7330
rect 3345 7295 3385 7300
rect 3345 7265 3350 7295
rect 3350 7265 3380 7295
rect 3380 7265 3385 7295
rect 3345 7260 3385 7265
rect 3345 7235 3385 7240
rect 3345 7205 3350 7235
rect 3350 7205 3380 7235
rect 3380 7205 3385 7235
rect 3345 7200 3385 7205
rect 3345 7170 3385 7175
rect 3345 7140 3350 7170
rect 3350 7140 3380 7170
rect 3380 7140 3385 7170
rect 3345 7135 3385 7140
rect 3345 7100 3385 7105
rect 3345 7070 3350 7100
rect 3350 7070 3380 7100
rect 3380 7070 3385 7100
rect 3345 7065 3385 7070
rect 3345 7030 3385 7035
rect 3345 7000 3350 7030
rect 3350 7000 3380 7030
rect 3380 7000 3385 7030
rect 3345 6995 3385 7000
rect 3345 6960 3385 6965
rect 3345 6930 3350 6960
rect 3350 6930 3380 6960
rect 3380 6930 3385 6960
rect 3345 6925 3385 6930
rect 3345 6895 3385 6900
rect 3345 6865 3350 6895
rect 3350 6865 3380 6895
rect 3380 6865 3385 6895
rect 3345 6860 3385 6865
rect 3345 6835 3385 6840
rect 3345 6805 3350 6835
rect 3350 6805 3380 6835
rect 3380 6805 3385 6835
rect 3345 6800 3385 6805
rect 3345 6770 3385 6775
rect 3345 6740 3350 6770
rect 3350 6740 3380 6770
rect 3380 6740 3385 6770
rect 3345 6735 3385 6740
rect 3345 6700 3385 6705
rect 3345 6670 3350 6700
rect 3350 6670 3380 6700
rect 3380 6670 3385 6700
rect 3345 6665 3385 6670
rect 3345 6630 3385 6635
rect 3345 6600 3350 6630
rect 3350 6600 3380 6630
rect 3380 6600 3385 6630
rect 3345 6595 3385 6600
rect 3345 6560 3385 6565
rect 3345 6530 3350 6560
rect 3350 6530 3380 6560
rect 3380 6530 3385 6560
rect 3345 6525 3385 6530
rect 3345 6495 3385 6500
rect 3345 6465 3350 6495
rect 3350 6465 3380 6495
rect 3380 6465 3385 6495
rect 3345 6460 3385 6465
rect 6630 9635 6670 9640
rect 6630 9605 6635 9635
rect 6635 9605 6665 9635
rect 6665 9605 6670 9635
rect 6630 9600 6670 9605
rect 6630 9570 6670 9575
rect 6630 9540 6635 9570
rect 6635 9540 6665 9570
rect 6665 9540 6670 9570
rect 6630 9535 6670 9540
rect 6630 9500 6670 9505
rect 6630 9470 6635 9500
rect 6635 9470 6665 9500
rect 6665 9470 6670 9500
rect 6630 9465 6670 9470
rect 6630 9430 6670 9435
rect 6630 9400 6635 9430
rect 6635 9400 6665 9430
rect 6665 9400 6670 9430
rect 6630 9395 6670 9400
rect 6630 9360 6670 9365
rect 6630 9330 6635 9360
rect 6635 9330 6665 9360
rect 6665 9330 6670 9360
rect 6630 9325 6670 9330
rect 6630 9295 6670 9300
rect 6630 9265 6635 9295
rect 6635 9265 6665 9295
rect 6665 9265 6670 9295
rect 6630 9260 6670 9265
rect 6630 9235 6670 9240
rect 6630 9205 6635 9235
rect 6635 9205 6665 9235
rect 6665 9205 6670 9235
rect 6630 9200 6670 9205
rect 6630 9170 6670 9175
rect 6630 9140 6635 9170
rect 6635 9140 6665 9170
rect 6665 9140 6670 9170
rect 6630 9135 6670 9140
rect 6630 9100 6670 9105
rect 6630 9070 6635 9100
rect 6635 9070 6665 9100
rect 6665 9070 6670 9100
rect 6630 9065 6670 9070
rect 6630 9030 6670 9035
rect 6630 9000 6635 9030
rect 6635 9000 6665 9030
rect 6665 9000 6670 9030
rect 6630 8995 6670 9000
rect 6630 8960 6670 8965
rect 6630 8930 6635 8960
rect 6635 8930 6665 8960
rect 6665 8930 6670 8960
rect 6630 8925 6670 8930
rect 6630 8895 6670 8900
rect 6630 8865 6635 8895
rect 6635 8865 6665 8895
rect 6665 8865 6670 8895
rect 6630 8860 6670 8865
rect 6630 8835 6670 8840
rect 6630 8805 6635 8835
rect 6635 8805 6665 8835
rect 6665 8805 6670 8835
rect 6630 8800 6670 8805
rect 6630 8770 6670 8775
rect 6630 8740 6635 8770
rect 6635 8740 6665 8770
rect 6665 8740 6670 8770
rect 6630 8735 6670 8740
rect 6630 8700 6670 8705
rect 6630 8670 6635 8700
rect 6635 8670 6665 8700
rect 6665 8670 6670 8700
rect 6630 8665 6670 8670
rect 6630 8630 6670 8635
rect 6630 8600 6635 8630
rect 6635 8600 6665 8630
rect 6665 8600 6670 8630
rect 6630 8595 6670 8600
rect 6630 8560 6670 8565
rect 6630 8530 6635 8560
rect 6635 8530 6665 8560
rect 6665 8530 6670 8560
rect 6630 8525 6670 8530
rect 6630 8495 6670 8500
rect 6630 8465 6635 8495
rect 6635 8465 6665 8495
rect 6665 8465 6670 8495
rect 6630 8460 6670 8465
rect 6630 8435 6670 8440
rect 6630 8405 6635 8435
rect 6635 8405 6665 8435
rect 6665 8405 6670 8435
rect 6630 8400 6670 8405
rect 6630 8370 6670 8375
rect 6630 8340 6635 8370
rect 6635 8340 6665 8370
rect 6665 8340 6670 8370
rect 6630 8335 6670 8340
rect 6630 8300 6670 8305
rect 6630 8270 6635 8300
rect 6635 8270 6665 8300
rect 6665 8270 6670 8300
rect 6630 8265 6670 8270
rect 6630 8230 6670 8235
rect 6630 8200 6635 8230
rect 6635 8200 6665 8230
rect 6665 8200 6670 8230
rect 6630 8195 6670 8200
rect 6630 8160 6670 8165
rect 6630 8130 6635 8160
rect 6635 8130 6665 8160
rect 6665 8130 6670 8160
rect 6630 8125 6670 8130
rect 6630 8095 6670 8100
rect 6630 8065 6635 8095
rect 6635 8065 6665 8095
rect 6665 8065 6670 8095
rect 6630 8060 6670 8065
rect 6630 8035 6670 8040
rect 6630 8005 6635 8035
rect 6635 8005 6665 8035
rect 6665 8005 6670 8035
rect 6630 8000 6670 8005
rect 6630 7970 6670 7975
rect 6630 7940 6635 7970
rect 6635 7940 6665 7970
rect 6665 7940 6670 7970
rect 6630 7935 6670 7940
rect 6630 7900 6670 7905
rect 6630 7870 6635 7900
rect 6635 7870 6665 7900
rect 6665 7870 6670 7900
rect 6630 7865 6670 7870
rect 6630 7830 6670 7835
rect 6630 7800 6635 7830
rect 6635 7800 6665 7830
rect 6665 7800 6670 7830
rect 6630 7795 6670 7800
rect 6630 7760 6670 7765
rect 6630 7730 6635 7760
rect 6635 7730 6665 7760
rect 6665 7730 6670 7760
rect 6630 7725 6670 7730
rect 6630 7695 6670 7700
rect 6630 7665 6635 7695
rect 6635 7665 6665 7695
rect 6665 7665 6670 7695
rect 6630 7660 6670 7665
rect 6630 7635 6670 7640
rect 6630 7605 6635 7635
rect 6635 7605 6665 7635
rect 6665 7605 6670 7635
rect 6630 7600 6670 7605
rect 6630 7570 6670 7575
rect 6630 7540 6635 7570
rect 6635 7540 6665 7570
rect 6665 7540 6670 7570
rect 6630 7535 6670 7540
rect 6630 7500 6670 7505
rect 6630 7470 6635 7500
rect 6635 7470 6665 7500
rect 6665 7470 6670 7500
rect 6630 7465 6670 7470
rect 6630 7430 6670 7435
rect 6630 7400 6635 7430
rect 6635 7400 6665 7430
rect 6665 7400 6670 7430
rect 6630 7395 6670 7400
rect 6630 7360 6670 7365
rect 6630 7330 6635 7360
rect 6635 7330 6665 7360
rect 6665 7330 6670 7360
rect 6630 7325 6670 7330
rect 6630 7295 6670 7300
rect 6630 7265 6635 7295
rect 6635 7265 6665 7295
rect 6665 7265 6670 7295
rect 6630 7260 6670 7265
rect 6630 7235 6670 7240
rect 6630 7205 6635 7235
rect 6635 7205 6665 7235
rect 6665 7205 6670 7235
rect 6630 7200 6670 7205
rect 6630 7170 6670 7175
rect 6630 7140 6635 7170
rect 6635 7140 6665 7170
rect 6665 7140 6670 7170
rect 6630 7135 6670 7140
rect 6630 7100 6670 7105
rect 6630 7070 6635 7100
rect 6635 7070 6665 7100
rect 6665 7070 6670 7100
rect 6630 7065 6670 7070
rect 6630 7030 6670 7035
rect 6630 7000 6635 7030
rect 6635 7000 6665 7030
rect 6665 7000 6670 7030
rect 6630 6995 6670 7000
rect 6630 6960 6670 6965
rect 6630 6930 6635 6960
rect 6635 6930 6665 6960
rect 6665 6930 6670 6960
rect 6630 6925 6670 6930
rect 6630 6895 6670 6900
rect 6630 6865 6635 6895
rect 6635 6865 6665 6895
rect 6665 6865 6670 6895
rect 6630 6860 6670 6865
rect 6630 6835 6670 6840
rect 6630 6805 6635 6835
rect 6635 6805 6665 6835
rect 6665 6805 6670 6835
rect 6630 6800 6670 6805
rect 6630 6770 6670 6775
rect 6630 6740 6635 6770
rect 6635 6740 6665 6770
rect 6665 6740 6670 6770
rect 6630 6735 6670 6740
rect 6630 6700 6670 6705
rect 6630 6670 6635 6700
rect 6635 6670 6665 6700
rect 6665 6670 6670 6700
rect 6630 6665 6670 6670
rect 6630 6630 6670 6635
rect 6630 6600 6635 6630
rect 6635 6600 6665 6630
rect 6665 6600 6670 6630
rect 6630 6595 6670 6600
rect 6630 6560 6670 6565
rect 6630 6530 6635 6560
rect 6635 6530 6665 6560
rect 6665 6530 6670 6560
rect 6630 6525 6670 6530
rect 6630 6495 6670 6500
rect 6630 6465 6635 6495
rect 6635 6465 6665 6495
rect 6665 6465 6670 6495
rect 6630 6460 6670 6465
rect 7270 9635 7310 9640
rect 7270 9605 7275 9635
rect 7275 9605 7305 9635
rect 7305 9605 7310 9635
rect 7270 9600 7310 9605
rect 7270 9570 7310 9575
rect 7270 9540 7275 9570
rect 7275 9540 7305 9570
rect 7305 9540 7310 9570
rect 7270 9535 7310 9540
rect 7270 9500 7310 9505
rect 7270 9470 7275 9500
rect 7275 9470 7305 9500
rect 7305 9470 7310 9500
rect 7270 9465 7310 9470
rect 7270 9430 7310 9435
rect 7270 9400 7275 9430
rect 7275 9400 7305 9430
rect 7305 9400 7310 9430
rect 7270 9395 7310 9400
rect 7270 9360 7310 9365
rect 7270 9330 7275 9360
rect 7275 9330 7305 9360
rect 7305 9330 7310 9360
rect 7270 9325 7310 9330
rect 7270 9295 7310 9300
rect 7270 9265 7275 9295
rect 7275 9265 7305 9295
rect 7305 9265 7310 9295
rect 7270 9260 7310 9265
rect 7270 9235 7310 9240
rect 7270 9205 7275 9235
rect 7275 9205 7305 9235
rect 7305 9205 7310 9235
rect 7270 9200 7310 9205
rect 7270 9170 7310 9175
rect 7270 9140 7275 9170
rect 7275 9140 7305 9170
rect 7305 9140 7310 9170
rect 7270 9135 7310 9140
rect 7270 9100 7310 9105
rect 7270 9070 7275 9100
rect 7275 9070 7305 9100
rect 7305 9070 7310 9100
rect 7270 9065 7310 9070
rect 7270 9030 7310 9035
rect 7270 9000 7275 9030
rect 7275 9000 7305 9030
rect 7305 9000 7310 9030
rect 7270 8995 7310 9000
rect 7270 8960 7310 8965
rect 7270 8930 7275 8960
rect 7275 8930 7305 8960
rect 7305 8930 7310 8960
rect 7270 8925 7310 8930
rect 7270 8895 7310 8900
rect 7270 8865 7275 8895
rect 7275 8865 7305 8895
rect 7305 8865 7310 8895
rect 7270 8860 7310 8865
rect 7270 8835 7310 8840
rect 7270 8805 7275 8835
rect 7275 8805 7305 8835
rect 7305 8805 7310 8835
rect 7270 8800 7310 8805
rect 7270 8770 7310 8775
rect 7270 8740 7275 8770
rect 7275 8740 7305 8770
rect 7305 8740 7310 8770
rect 7270 8735 7310 8740
rect 7270 8700 7310 8705
rect 7270 8670 7275 8700
rect 7275 8670 7305 8700
rect 7305 8670 7310 8700
rect 7270 8665 7310 8670
rect 7270 8630 7310 8635
rect 7270 8600 7275 8630
rect 7275 8600 7305 8630
rect 7305 8600 7310 8630
rect 7270 8595 7310 8600
rect 7270 8560 7310 8565
rect 7270 8530 7275 8560
rect 7275 8530 7305 8560
rect 7305 8530 7310 8560
rect 7270 8525 7310 8530
rect 7270 8495 7310 8500
rect 7270 8465 7275 8495
rect 7275 8465 7305 8495
rect 7305 8465 7310 8495
rect 7270 8460 7310 8465
rect 7270 8435 7310 8440
rect 7270 8405 7275 8435
rect 7275 8405 7305 8435
rect 7305 8405 7310 8435
rect 7270 8400 7310 8405
rect 7270 8370 7310 8375
rect 7270 8340 7275 8370
rect 7275 8340 7305 8370
rect 7305 8340 7310 8370
rect 7270 8335 7310 8340
rect 7270 8300 7310 8305
rect 7270 8270 7275 8300
rect 7275 8270 7305 8300
rect 7305 8270 7310 8300
rect 7270 8265 7310 8270
rect 7270 8230 7310 8235
rect 7270 8200 7275 8230
rect 7275 8200 7305 8230
rect 7305 8200 7310 8230
rect 7270 8195 7310 8200
rect 7270 8160 7310 8165
rect 7270 8130 7275 8160
rect 7275 8130 7305 8160
rect 7305 8130 7310 8160
rect 7270 8125 7310 8130
rect 7270 8095 7310 8100
rect 7270 8065 7275 8095
rect 7275 8065 7305 8095
rect 7305 8065 7310 8095
rect 7270 8060 7310 8065
rect 7270 8035 7310 8040
rect 7270 8005 7275 8035
rect 7275 8005 7305 8035
rect 7305 8005 7310 8035
rect 7270 8000 7310 8005
rect 7270 7970 7310 7975
rect 7270 7940 7275 7970
rect 7275 7940 7305 7970
rect 7305 7940 7310 7970
rect 7270 7935 7310 7940
rect 7270 7900 7310 7905
rect 7270 7870 7275 7900
rect 7275 7870 7305 7900
rect 7305 7870 7310 7900
rect 7270 7865 7310 7870
rect 7270 7830 7310 7835
rect 7270 7800 7275 7830
rect 7275 7800 7305 7830
rect 7305 7800 7310 7830
rect 7270 7795 7310 7800
rect 7270 7760 7310 7765
rect 7270 7730 7275 7760
rect 7275 7730 7305 7760
rect 7305 7730 7310 7760
rect 7270 7725 7310 7730
rect 7270 7695 7310 7700
rect 7270 7665 7275 7695
rect 7275 7665 7305 7695
rect 7305 7665 7310 7695
rect 7270 7660 7310 7665
rect 7270 7635 7310 7640
rect 7270 7605 7275 7635
rect 7275 7605 7305 7635
rect 7305 7605 7310 7635
rect 7270 7600 7310 7605
rect 7270 7570 7310 7575
rect 7270 7540 7275 7570
rect 7275 7540 7305 7570
rect 7305 7540 7310 7570
rect 7270 7535 7310 7540
rect 7270 7500 7310 7505
rect 7270 7470 7275 7500
rect 7275 7470 7305 7500
rect 7305 7470 7310 7500
rect 7270 7465 7310 7470
rect 7270 7430 7310 7435
rect 7270 7400 7275 7430
rect 7275 7400 7305 7430
rect 7305 7400 7310 7430
rect 7270 7395 7310 7400
rect 7270 7360 7310 7365
rect 7270 7330 7275 7360
rect 7275 7330 7305 7360
rect 7305 7330 7310 7360
rect 7270 7325 7310 7330
rect 7270 7295 7310 7300
rect 7270 7265 7275 7295
rect 7275 7265 7305 7295
rect 7305 7265 7310 7295
rect 7270 7260 7310 7265
rect 7270 7235 7310 7240
rect 7270 7205 7275 7235
rect 7275 7205 7305 7235
rect 7305 7205 7310 7235
rect 7270 7200 7310 7205
rect 7270 7170 7310 7175
rect 7270 7140 7275 7170
rect 7275 7140 7305 7170
rect 7305 7140 7310 7170
rect 7270 7135 7310 7140
rect 7270 7100 7310 7105
rect 7270 7070 7275 7100
rect 7275 7070 7305 7100
rect 7305 7070 7310 7100
rect 7270 7065 7310 7070
rect 7270 7030 7310 7035
rect 7270 7000 7275 7030
rect 7275 7000 7305 7030
rect 7305 7000 7310 7030
rect 7270 6995 7310 7000
rect 7270 6960 7310 6965
rect 7270 6930 7275 6960
rect 7275 6930 7305 6960
rect 7305 6930 7310 6960
rect 7270 6925 7310 6930
rect 7270 6895 7310 6900
rect 7270 6865 7275 6895
rect 7275 6865 7305 6895
rect 7305 6865 7310 6895
rect 7270 6860 7310 6865
rect 7270 6835 7310 6840
rect 7270 6805 7275 6835
rect 7275 6805 7305 6835
rect 7305 6805 7310 6835
rect 7270 6800 7310 6805
rect 7270 6770 7310 6775
rect 7270 6740 7275 6770
rect 7275 6740 7305 6770
rect 7305 6740 7310 6770
rect 7270 6735 7310 6740
rect 7270 6700 7310 6705
rect 7270 6670 7275 6700
rect 7275 6670 7305 6700
rect 7305 6670 7310 6700
rect 7270 6665 7310 6670
rect 7270 6630 7310 6635
rect 7270 6600 7275 6630
rect 7275 6600 7305 6630
rect 7305 6600 7310 6630
rect 7270 6595 7310 6600
rect 7270 6560 7310 6565
rect 7270 6530 7275 6560
rect 7275 6530 7305 6560
rect 7305 6530 7310 6560
rect 7270 6525 7310 6530
rect 7270 6495 7310 6500
rect 7270 6465 7275 6495
rect 7275 6465 7305 6495
rect 7305 6465 7310 6495
rect 7270 6460 7310 6465
rect 7970 9635 8010 9640
rect 7970 9605 7975 9635
rect 7975 9605 8005 9635
rect 8005 9605 8010 9635
rect 7970 9600 8010 9605
rect 7970 9570 8010 9575
rect 7970 9540 7975 9570
rect 7975 9540 8005 9570
rect 8005 9540 8010 9570
rect 7970 9535 8010 9540
rect 7970 9500 8010 9505
rect 7970 9470 7975 9500
rect 7975 9470 8005 9500
rect 8005 9470 8010 9500
rect 7970 9465 8010 9470
rect 7970 9430 8010 9435
rect 7970 9400 7975 9430
rect 7975 9400 8005 9430
rect 8005 9400 8010 9430
rect 7970 9395 8010 9400
rect 7970 9360 8010 9365
rect 7970 9330 7975 9360
rect 7975 9330 8005 9360
rect 8005 9330 8010 9360
rect 7970 9325 8010 9330
rect 7970 9295 8010 9300
rect 7970 9265 7975 9295
rect 7975 9265 8005 9295
rect 8005 9265 8010 9295
rect 7970 9260 8010 9265
rect 7970 9235 8010 9240
rect 7970 9205 7975 9235
rect 7975 9205 8005 9235
rect 8005 9205 8010 9235
rect 7970 9200 8010 9205
rect 7970 9170 8010 9175
rect 7970 9140 7975 9170
rect 7975 9140 8005 9170
rect 8005 9140 8010 9170
rect 7970 9135 8010 9140
rect 7970 9100 8010 9105
rect 7970 9070 7975 9100
rect 7975 9070 8005 9100
rect 8005 9070 8010 9100
rect 7970 9065 8010 9070
rect 7970 9030 8010 9035
rect 7970 9000 7975 9030
rect 7975 9000 8005 9030
rect 8005 9000 8010 9030
rect 7970 8995 8010 9000
rect 7970 8960 8010 8965
rect 7970 8930 7975 8960
rect 7975 8930 8005 8960
rect 8005 8930 8010 8960
rect 7970 8925 8010 8930
rect 7970 8895 8010 8900
rect 7970 8865 7975 8895
rect 7975 8865 8005 8895
rect 8005 8865 8010 8895
rect 7970 8860 8010 8865
rect 7970 8835 8010 8840
rect 7970 8805 7975 8835
rect 7975 8805 8005 8835
rect 8005 8805 8010 8835
rect 7970 8800 8010 8805
rect 7970 8770 8010 8775
rect 7970 8740 7975 8770
rect 7975 8740 8005 8770
rect 8005 8740 8010 8770
rect 7970 8735 8010 8740
rect 7970 8700 8010 8705
rect 7970 8670 7975 8700
rect 7975 8670 8005 8700
rect 8005 8670 8010 8700
rect 7970 8665 8010 8670
rect 7970 8630 8010 8635
rect 7970 8600 7975 8630
rect 7975 8600 8005 8630
rect 8005 8600 8010 8630
rect 7970 8595 8010 8600
rect 7970 8560 8010 8565
rect 7970 8530 7975 8560
rect 7975 8530 8005 8560
rect 8005 8530 8010 8560
rect 7970 8525 8010 8530
rect 7970 8495 8010 8500
rect 7970 8465 7975 8495
rect 7975 8465 8005 8495
rect 8005 8465 8010 8495
rect 7970 8460 8010 8465
rect 7970 8435 8010 8440
rect 7970 8405 7975 8435
rect 7975 8405 8005 8435
rect 8005 8405 8010 8435
rect 7970 8400 8010 8405
rect 7970 8370 8010 8375
rect 7970 8340 7975 8370
rect 7975 8340 8005 8370
rect 8005 8340 8010 8370
rect 7970 8335 8010 8340
rect 7970 8300 8010 8305
rect 7970 8270 7975 8300
rect 7975 8270 8005 8300
rect 8005 8270 8010 8300
rect 7970 8265 8010 8270
rect 7970 8230 8010 8235
rect 7970 8200 7975 8230
rect 7975 8200 8005 8230
rect 8005 8200 8010 8230
rect 7970 8195 8010 8200
rect 7970 8160 8010 8165
rect 7970 8130 7975 8160
rect 7975 8130 8005 8160
rect 8005 8130 8010 8160
rect 7970 8125 8010 8130
rect 7970 8095 8010 8100
rect 7970 8065 7975 8095
rect 7975 8065 8005 8095
rect 8005 8065 8010 8095
rect 7970 8060 8010 8065
rect 7970 8035 8010 8040
rect 7970 8005 7975 8035
rect 7975 8005 8005 8035
rect 8005 8005 8010 8035
rect 7970 8000 8010 8005
rect 7970 7970 8010 7975
rect 7970 7940 7975 7970
rect 7975 7940 8005 7970
rect 8005 7940 8010 7970
rect 7970 7935 8010 7940
rect 7970 7900 8010 7905
rect 7970 7870 7975 7900
rect 7975 7870 8005 7900
rect 8005 7870 8010 7900
rect 7970 7865 8010 7870
rect 7970 7830 8010 7835
rect 7970 7800 7975 7830
rect 7975 7800 8005 7830
rect 8005 7800 8010 7830
rect 7970 7795 8010 7800
rect 7970 7760 8010 7765
rect 7970 7730 7975 7760
rect 7975 7730 8005 7760
rect 8005 7730 8010 7760
rect 7970 7725 8010 7730
rect 7970 7695 8010 7700
rect 7970 7665 7975 7695
rect 7975 7665 8005 7695
rect 8005 7665 8010 7695
rect 7970 7660 8010 7665
rect 7970 7635 8010 7640
rect 7970 7605 7975 7635
rect 7975 7605 8005 7635
rect 8005 7605 8010 7635
rect 7970 7600 8010 7605
rect 7970 7570 8010 7575
rect 7970 7540 7975 7570
rect 7975 7540 8005 7570
rect 8005 7540 8010 7570
rect 7970 7535 8010 7540
rect 7970 7500 8010 7505
rect 7970 7470 7975 7500
rect 7975 7470 8005 7500
rect 8005 7470 8010 7500
rect 7970 7465 8010 7470
rect 7970 7430 8010 7435
rect 7970 7400 7975 7430
rect 7975 7400 8005 7430
rect 8005 7400 8010 7430
rect 7970 7395 8010 7400
rect 7970 7360 8010 7365
rect 7970 7330 7975 7360
rect 7975 7330 8005 7360
rect 8005 7330 8010 7360
rect 7970 7325 8010 7330
rect 7970 7295 8010 7300
rect 7970 7265 7975 7295
rect 7975 7265 8005 7295
rect 8005 7265 8010 7295
rect 7970 7260 8010 7265
rect 7970 7235 8010 7240
rect 7970 7205 7975 7235
rect 7975 7205 8005 7235
rect 8005 7205 8010 7235
rect 7970 7200 8010 7205
rect 7970 7170 8010 7175
rect 7970 7140 7975 7170
rect 7975 7140 8005 7170
rect 8005 7140 8010 7170
rect 7970 7135 8010 7140
rect 7970 7100 8010 7105
rect 7970 7070 7975 7100
rect 7975 7070 8005 7100
rect 8005 7070 8010 7100
rect 7970 7065 8010 7070
rect 7970 7030 8010 7035
rect 7970 7000 7975 7030
rect 7975 7000 8005 7030
rect 8005 7000 8010 7030
rect 7970 6995 8010 7000
rect 7970 6960 8010 6965
rect 7970 6930 7975 6960
rect 7975 6930 8005 6960
rect 8005 6930 8010 6960
rect 7970 6925 8010 6930
rect 7970 6895 8010 6900
rect 7970 6865 7975 6895
rect 7975 6865 8005 6895
rect 8005 6865 8010 6895
rect 7970 6860 8010 6865
rect 7970 6835 8010 6840
rect 7970 6805 7975 6835
rect 7975 6805 8005 6835
rect 8005 6805 8010 6835
rect 7970 6800 8010 6805
rect 7970 6770 8010 6775
rect 7970 6740 7975 6770
rect 7975 6740 8005 6770
rect 8005 6740 8010 6770
rect 7970 6735 8010 6740
rect 7970 6700 8010 6705
rect 7970 6670 7975 6700
rect 7975 6670 8005 6700
rect 8005 6670 8010 6700
rect 7970 6665 8010 6670
rect 7970 6630 8010 6635
rect 7970 6600 7975 6630
rect 7975 6600 8005 6630
rect 8005 6600 8010 6630
rect 7970 6595 8010 6600
rect 7970 6560 8010 6565
rect 7970 6530 7975 6560
rect 7975 6530 8005 6560
rect 8005 6530 8010 6560
rect 7970 6525 8010 6530
rect 7970 6495 8010 6500
rect 7970 6465 7975 6495
rect 7975 6465 8005 6495
rect 8005 6465 8010 6495
rect 7970 6460 8010 6465
rect 8320 9635 8360 9640
rect 8320 9605 8325 9635
rect 8325 9605 8355 9635
rect 8355 9605 8360 9635
rect 8320 9600 8360 9605
rect 8320 9570 8360 9575
rect 8320 9540 8325 9570
rect 8325 9540 8355 9570
rect 8355 9540 8360 9570
rect 8320 9535 8360 9540
rect 8320 9500 8360 9505
rect 8320 9470 8325 9500
rect 8325 9470 8355 9500
rect 8355 9470 8360 9500
rect 8320 9465 8360 9470
rect 8320 9430 8360 9435
rect 8320 9400 8325 9430
rect 8325 9400 8355 9430
rect 8355 9400 8360 9430
rect 8320 9395 8360 9400
rect 8320 9360 8360 9365
rect 8320 9330 8325 9360
rect 8325 9330 8355 9360
rect 8355 9330 8360 9360
rect 8320 9325 8360 9330
rect 8320 9295 8360 9300
rect 8320 9265 8325 9295
rect 8325 9265 8355 9295
rect 8355 9265 8360 9295
rect 8320 9260 8360 9265
rect 8320 9235 8360 9240
rect 8320 9205 8325 9235
rect 8325 9205 8355 9235
rect 8355 9205 8360 9235
rect 8320 9200 8360 9205
rect 8320 9170 8360 9175
rect 8320 9140 8325 9170
rect 8325 9140 8355 9170
rect 8355 9140 8360 9170
rect 8320 9135 8360 9140
rect 8320 9100 8360 9105
rect 8320 9070 8325 9100
rect 8325 9070 8355 9100
rect 8355 9070 8360 9100
rect 8320 9065 8360 9070
rect 8320 9030 8360 9035
rect 8320 9000 8325 9030
rect 8325 9000 8355 9030
rect 8355 9000 8360 9030
rect 8320 8995 8360 9000
rect 8320 8960 8360 8965
rect 8320 8930 8325 8960
rect 8325 8930 8355 8960
rect 8355 8930 8360 8960
rect 8320 8925 8360 8930
rect 8320 8895 8360 8900
rect 8320 8865 8325 8895
rect 8325 8865 8355 8895
rect 8355 8865 8360 8895
rect 8320 8860 8360 8865
rect 8320 8835 8360 8840
rect 8320 8805 8325 8835
rect 8325 8805 8355 8835
rect 8355 8805 8360 8835
rect 8320 8800 8360 8805
rect 8320 8770 8360 8775
rect 8320 8740 8325 8770
rect 8325 8740 8355 8770
rect 8355 8740 8360 8770
rect 8320 8735 8360 8740
rect 8320 8700 8360 8705
rect 8320 8670 8325 8700
rect 8325 8670 8355 8700
rect 8355 8670 8360 8700
rect 8320 8665 8360 8670
rect 8320 8630 8360 8635
rect 8320 8600 8325 8630
rect 8325 8600 8355 8630
rect 8355 8600 8360 8630
rect 8320 8595 8360 8600
rect 8320 8560 8360 8565
rect 8320 8530 8325 8560
rect 8325 8530 8355 8560
rect 8355 8530 8360 8560
rect 8320 8525 8360 8530
rect 8320 8495 8360 8500
rect 8320 8465 8325 8495
rect 8325 8465 8355 8495
rect 8355 8465 8360 8495
rect 8320 8460 8360 8465
rect 8320 8435 8360 8440
rect 8320 8405 8325 8435
rect 8325 8405 8355 8435
rect 8355 8405 8360 8435
rect 8320 8400 8360 8405
rect 8320 8370 8360 8375
rect 8320 8340 8325 8370
rect 8325 8340 8355 8370
rect 8355 8340 8360 8370
rect 8320 8335 8360 8340
rect 8320 8300 8360 8305
rect 8320 8270 8325 8300
rect 8325 8270 8355 8300
rect 8355 8270 8360 8300
rect 8320 8265 8360 8270
rect 8320 8230 8360 8235
rect 8320 8200 8325 8230
rect 8325 8200 8355 8230
rect 8355 8200 8360 8230
rect 8320 8195 8360 8200
rect 8320 8160 8360 8165
rect 8320 8130 8325 8160
rect 8325 8130 8355 8160
rect 8355 8130 8360 8160
rect 8320 8125 8360 8130
rect 8320 8095 8360 8100
rect 8320 8065 8325 8095
rect 8325 8065 8355 8095
rect 8355 8065 8360 8095
rect 8320 8060 8360 8065
rect 8320 8035 8360 8040
rect 8320 8005 8325 8035
rect 8325 8005 8355 8035
rect 8355 8005 8360 8035
rect 8320 8000 8360 8005
rect 8320 7970 8360 7975
rect 8320 7940 8325 7970
rect 8325 7940 8355 7970
rect 8355 7940 8360 7970
rect 8320 7935 8360 7940
rect 8320 7900 8360 7905
rect 8320 7870 8325 7900
rect 8325 7870 8355 7900
rect 8355 7870 8360 7900
rect 8320 7865 8360 7870
rect 8320 7830 8360 7835
rect 8320 7800 8325 7830
rect 8325 7800 8355 7830
rect 8355 7800 8360 7830
rect 8320 7795 8360 7800
rect 8320 7760 8360 7765
rect 8320 7730 8325 7760
rect 8325 7730 8355 7760
rect 8355 7730 8360 7760
rect 8320 7725 8360 7730
rect 8320 7695 8360 7700
rect 8320 7665 8325 7695
rect 8325 7665 8355 7695
rect 8355 7665 8360 7695
rect 8320 7660 8360 7665
rect 8320 7635 8360 7640
rect 8320 7605 8325 7635
rect 8325 7605 8355 7635
rect 8355 7605 8360 7635
rect 8320 7600 8360 7605
rect 8320 7570 8360 7575
rect 8320 7540 8325 7570
rect 8325 7540 8355 7570
rect 8355 7540 8360 7570
rect 8320 7535 8360 7540
rect 8320 7500 8360 7505
rect 8320 7470 8325 7500
rect 8325 7470 8355 7500
rect 8355 7470 8360 7500
rect 8320 7465 8360 7470
rect 8320 7430 8360 7435
rect 8320 7400 8325 7430
rect 8325 7400 8355 7430
rect 8355 7400 8360 7430
rect 8320 7395 8360 7400
rect 8320 7360 8360 7365
rect 8320 7330 8325 7360
rect 8325 7330 8355 7360
rect 8355 7330 8360 7360
rect 8320 7325 8360 7330
rect 8320 7295 8360 7300
rect 8320 7265 8325 7295
rect 8325 7265 8355 7295
rect 8355 7265 8360 7295
rect 8320 7260 8360 7265
rect 8320 7235 8360 7240
rect 8320 7205 8325 7235
rect 8325 7205 8355 7235
rect 8355 7205 8360 7235
rect 8320 7200 8360 7205
rect 8320 7170 8360 7175
rect 8320 7140 8325 7170
rect 8325 7140 8355 7170
rect 8355 7140 8360 7170
rect 8320 7135 8360 7140
rect 8320 7100 8360 7105
rect 8320 7070 8325 7100
rect 8325 7070 8355 7100
rect 8355 7070 8360 7100
rect 8320 7065 8360 7070
rect 8320 7030 8360 7035
rect 8320 7000 8325 7030
rect 8325 7000 8355 7030
rect 8355 7000 8360 7030
rect 8320 6995 8360 7000
rect 8320 6960 8360 6965
rect 8320 6930 8325 6960
rect 8325 6930 8355 6960
rect 8355 6930 8360 6960
rect 8320 6925 8360 6930
rect 8320 6895 8360 6900
rect 8320 6865 8325 6895
rect 8325 6865 8355 6895
rect 8355 6865 8360 6895
rect 8320 6860 8360 6865
rect 8320 6835 8360 6840
rect 8320 6805 8325 6835
rect 8325 6805 8355 6835
rect 8355 6805 8360 6835
rect 8320 6800 8360 6805
rect 8320 6770 8360 6775
rect 8320 6740 8325 6770
rect 8325 6740 8355 6770
rect 8355 6740 8360 6770
rect 8320 6735 8360 6740
rect 8320 6700 8360 6705
rect 8320 6670 8325 6700
rect 8325 6670 8355 6700
rect 8355 6670 8360 6700
rect 8320 6665 8360 6670
rect 8320 6630 8360 6635
rect 8320 6600 8325 6630
rect 8325 6600 8355 6630
rect 8355 6600 8360 6630
rect 8320 6595 8360 6600
rect 8320 6560 8360 6565
rect 8320 6530 8325 6560
rect 8325 6530 8355 6560
rect 8355 6530 8360 6560
rect 8320 6525 8360 6530
rect 8320 6495 8360 6500
rect 8320 6465 8325 6495
rect 8325 6465 8355 6495
rect 8355 6465 8360 6495
rect 8320 6460 8360 6465
rect 8670 9635 8710 9640
rect 8670 9605 8675 9635
rect 8675 9605 8705 9635
rect 8705 9605 8710 9635
rect 8670 9600 8710 9605
rect 8670 9570 8710 9575
rect 8670 9540 8675 9570
rect 8675 9540 8705 9570
rect 8705 9540 8710 9570
rect 8670 9535 8710 9540
rect 8670 9500 8710 9505
rect 8670 9470 8675 9500
rect 8675 9470 8705 9500
rect 8705 9470 8710 9500
rect 8670 9465 8710 9470
rect 8670 9430 8710 9435
rect 8670 9400 8675 9430
rect 8675 9400 8705 9430
rect 8705 9400 8710 9430
rect 8670 9395 8710 9400
rect 8670 9360 8710 9365
rect 8670 9330 8675 9360
rect 8675 9330 8705 9360
rect 8705 9330 8710 9360
rect 8670 9325 8710 9330
rect 8670 9295 8710 9300
rect 8670 9265 8675 9295
rect 8675 9265 8705 9295
rect 8705 9265 8710 9295
rect 8670 9260 8710 9265
rect 8670 9235 8710 9240
rect 8670 9205 8675 9235
rect 8675 9205 8705 9235
rect 8705 9205 8710 9235
rect 8670 9200 8710 9205
rect 8670 9170 8710 9175
rect 8670 9140 8675 9170
rect 8675 9140 8705 9170
rect 8705 9140 8710 9170
rect 8670 9135 8710 9140
rect 8670 9100 8710 9105
rect 8670 9070 8675 9100
rect 8675 9070 8705 9100
rect 8705 9070 8710 9100
rect 8670 9065 8710 9070
rect 8670 9030 8710 9035
rect 8670 9000 8675 9030
rect 8675 9000 8705 9030
rect 8705 9000 8710 9030
rect 8670 8995 8710 9000
rect 8670 8960 8710 8965
rect 8670 8930 8675 8960
rect 8675 8930 8705 8960
rect 8705 8930 8710 8960
rect 8670 8925 8710 8930
rect 8670 8895 8710 8900
rect 8670 8865 8675 8895
rect 8675 8865 8705 8895
rect 8705 8865 8710 8895
rect 8670 8860 8710 8865
rect 8670 8835 8710 8840
rect 8670 8805 8675 8835
rect 8675 8805 8705 8835
rect 8705 8805 8710 8835
rect 8670 8800 8710 8805
rect 8670 8770 8710 8775
rect 8670 8740 8675 8770
rect 8675 8740 8705 8770
rect 8705 8740 8710 8770
rect 8670 8735 8710 8740
rect 8670 8700 8710 8705
rect 8670 8670 8675 8700
rect 8675 8670 8705 8700
rect 8705 8670 8710 8700
rect 8670 8665 8710 8670
rect 8670 8630 8710 8635
rect 8670 8600 8675 8630
rect 8675 8600 8705 8630
rect 8705 8600 8710 8630
rect 8670 8595 8710 8600
rect 8670 8560 8710 8565
rect 8670 8530 8675 8560
rect 8675 8530 8705 8560
rect 8705 8530 8710 8560
rect 8670 8525 8710 8530
rect 8670 8495 8710 8500
rect 8670 8465 8675 8495
rect 8675 8465 8705 8495
rect 8705 8465 8710 8495
rect 8670 8460 8710 8465
rect 8670 8435 8710 8440
rect 8670 8405 8675 8435
rect 8675 8405 8705 8435
rect 8705 8405 8710 8435
rect 8670 8400 8710 8405
rect 8670 8370 8710 8375
rect 8670 8340 8675 8370
rect 8675 8340 8705 8370
rect 8705 8340 8710 8370
rect 8670 8335 8710 8340
rect 8670 8300 8710 8305
rect 8670 8270 8675 8300
rect 8675 8270 8705 8300
rect 8705 8270 8710 8300
rect 8670 8265 8710 8270
rect 8670 8230 8710 8235
rect 8670 8200 8675 8230
rect 8675 8200 8705 8230
rect 8705 8200 8710 8230
rect 8670 8195 8710 8200
rect 8670 8160 8710 8165
rect 8670 8130 8675 8160
rect 8675 8130 8705 8160
rect 8705 8130 8710 8160
rect 8670 8125 8710 8130
rect 8670 8095 8710 8100
rect 8670 8065 8675 8095
rect 8675 8065 8705 8095
rect 8705 8065 8710 8095
rect 8670 8060 8710 8065
rect 8670 8035 8710 8040
rect 8670 8005 8675 8035
rect 8675 8005 8705 8035
rect 8705 8005 8710 8035
rect 8670 8000 8710 8005
rect 8670 7970 8710 7975
rect 8670 7940 8675 7970
rect 8675 7940 8705 7970
rect 8705 7940 8710 7970
rect 8670 7935 8710 7940
rect 8670 7900 8710 7905
rect 8670 7870 8675 7900
rect 8675 7870 8705 7900
rect 8705 7870 8710 7900
rect 8670 7865 8710 7870
rect 8670 7830 8710 7835
rect 8670 7800 8675 7830
rect 8675 7800 8705 7830
rect 8705 7800 8710 7830
rect 8670 7795 8710 7800
rect 8670 7760 8710 7765
rect 8670 7730 8675 7760
rect 8675 7730 8705 7760
rect 8705 7730 8710 7760
rect 8670 7725 8710 7730
rect 8670 7695 8710 7700
rect 8670 7665 8675 7695
rect 8675 7665 8705 7695
rect 8705 7665 8710 7695
rect 8670 7660 8710 7665
rect 8670 7635 8710 7640
rect 8670 7605 8675 7635
rect 8675 7605 8705 7635
rect 8705 7605 8710 7635
rect 8670 7600 8710 7605
rect 8670 7570 8710 7575
rect 8670 7540 8675 7570
rect 8675 7540 8705 7570
rect 8705 7540 8710 7570
rect 8670 7535 8710 7540
rect 8670 7500 8710 7505
rect 8670 7470 8675 7500
rect 8675 7470 8705 7500
rect 8705 7470 8710 7500
rect 8670 7465 8710 7470
rect 8670 7430 8710 7435
rect 8670 7400 8675 7430
rect 8675 7400 8705 7430
rect 8705 7400 8710 7430
rect 8670 7395 8710 7400
rect 8670 7360 8710 7365
rect 8670 7330 8675 7360
rect 8675 7330 8705 7360
rect 8705 7330 8710 7360
rect 8670 7325 8710 7330
rect 8670 7295 8710 7300
rect 8670 7265 8675 7295
rect 8675 7265 8705 7295
rect 8705 7265 8710 7295
rect 8670 7260 8710 7265
rect 8670 7235 8710 7240
rect 8670 7205 8675 7235
rect 8675 7205 8705 7235
rect 8705 7205 8710 7235
rect 8670 7200 8710 7205
rect 8670 7170 8710 7175
rect 8670 7140 8675 7170
rect 8675 7140 8705 7170
rect 8705 7140 8710 7170
rect 8670 7135 8710 7140
rect 8670 7100 8710 7105
rect 8670 7070 8675 7100
rect 8675 7070 8705 7100
rect 8705 7070 8710 7100
rect 8670 7065 8710 7070
rect 8670 7030 8710 7035
rect 8670 7000 8675 7030
rect 8675 7000 8705 7030
rect 8705 7000 8710 7030
rect 8670 6995 8710 7000
rect 8670 6960 8710 6965
rect 8670 6930 8675 6960
rect 8675 6930 8705 6960
rect 8705 6930 8710 6960
rect 8670 6925 8710 6930
rect 8670 6895 8710 6900
rect 8670 6865 8675 6895
rect 8675 6865 8705 6895
rect 8705 6865 8710 6895
rect 8670 6860 8710 6865
rect 8670 6835 8710 6840
rect 8670 6805 8675 6835
rect 8675 6805 8705 6835
rect 8705 6805 8710 6835
rect 8670 6800 8710 6805
rect 8670 6770 8710 6775
rect 8670 6740 8675 6770
rect 8675 6740 8705 6770
rect 8705 6740 8710 6770
rect 8670 6735 8710 6740
rect 8670 6700 8710 6705
rect 8670 6670 8675 6700
rect 8675 6670 8705 6700
rect 8705 6670 8710 6700
rect 8670 6665 8710 6670
rect 8670 6630 8710 6635
rect 8670 6600 8675 6630
rect 8675 6600 8705 6630
rect 8705 6600 8710 6630
rect 8670 6595 8710 6600
rect 8670 6560 8710 6565
rect 8670 6530 8675 6560
rect 8675 6530 8705 6560
rect 8705 6530 8710 6560
rect 8670 6525 8710 6530
rect 8670 6495 8710 6500
rect 8670 6465 8675 6495
rect 8675 6465 8705 6495
rect 8705 6465 8710 6495
rect 8670 6460 8710 6465
rect 9020 9635 9060 9640
rect 9020 9605 9025 9635
rect 9025 9605 9055 9635
rect 9055 9605 9060 9635
rect 9020 9600 9060 9605
rect 9020 9570 9060 9575
rect 9020 9540 9025 9570
rect 9025 9540 9055 9570
rect 9055 9540 9060 9570
rect 9020 9535 9060 9540
rect 9020 9500 9060 9505
rect 9020 9470 9025 9500
rect 9025 9470 9055 9500
rect 9055 9470 9060 9500
rect 9020 9465 9060 9470
rect 9020 9430 9060 9435
rect 9020 9400 9025 9430
rect 9025 9400 9055 9430
rect 9055 9400 9060 9430
rect 9020 9395 9060 9400
rect 9020 9360 9060 9365
rect 9020 9330 9025 9360
rect 9025 9330 9055 9360
rect 9055 9330 9060 9360
rect 9020 9325 9060 9330
rect 9020 9295 9060 9300
rect 9020 9265 9025 9295
rect 9025 9265 9055 9295
rect 9055 9265 9060 9295
rect 9020 9260 9060 9265
rect 9020 9235 9060 9240
rect 9020 9205 9025 9235
rect 9025 9205 9055 9235
rect 9055 9205 9060 9235
rect 9020 9200 9060 9205
rect 9020 9170 9060 9175
rect 9020 9140 9025 9170
rect 9025 9140 9055 9170
rect 9055 9140 9060 9170
rect 9020 9135 9060 9140
rect 9020 9100 9060 9105
rect 9020 9070 9025 9100
rect 9025 9070 9055 9100
rect 9055 9070 9060 9100
rect 9020 9065 9060 9070
rect 9020 9030 9060 9035
rect 9020 9000 9025 9030
rect 9025 9000 9055 9030
rect 9055 9000 9060 9030
rect 9020 8995 9060 9000
rect 9020 8960 9060 8965
rect 9020 8930 9025 8960
rect 9025 8930 9055 8960
rect 9055 8930 9060 8960
rect 9020 8925 9060 8930
rect 9020 8895 9060 8900
rect 9020 8865 9025 8895
rect 9025 8865 9055 8895
rect 9055 8865 9060 8895
rect 9020 8860 9060 8865
rect 9020 8835 9060 8840
rect 9020 8805 9025 8835
rect 9025 8805 9055 8835
rect 9055 8805 9060 8835
rect 9020 8800 9060 8805
rect 9020 8770 9060 8775
rect 9020 8740 9025 8770
rect 9025 8740 9055 8770
rect 9055 8740 9060 8770
rect 9020 8735 9060 8740
rect 9020 8700 9060 8705
rect 9020 8670 9025 8700
rect 9025 8670 9055 8700
rect 9055 8670 9060 8700
rect 9020 8665 9060 8670
rect 9020 8630 9060 8635
rect 9020 8600 9025 8630
rect 9025 8600 9055 8630
rect 9055 8600 9060 8630
rect 9020 8595 9060 8600
rect 9020 8560 9060 8565
rect 9020 8530 9025 8560
rect 9025 8530 9055 8560
rect 9055 8530 9060 8560
rect 9020 8525 9060 8530
rect 9020 8495 9060 8500
rect 9020 8465 9025 8495
rect 9025 8465 9055 8495
rect 9055 8465 9060 8495
rect 9020 8460 9060 8465
rect 9020 8435 9060 8440
rect 9020 8405 9025 8435
rect 9025 8405 9055 8435
rect 9055 8405 9060 8435
rect 9020 8400 9060 8405
rect 9020 8370 9060 8375
rect 9020 8340 9025 8370
rect 9025 8340 9055 8370
rect 9055 8340 9060 8370
rect 9020 8335 9060 8340
rect 9020 8300 9060 8305
rect 9020 8270 9025 8300
rect 9025 8270 9055 8300
rect 9055 8270 9060 8300
rect 9020 8265 9060 8270
rect 9020 8230 9060 8235
rect 9020 8200 9025 8230
rect 9025 8200 9055 8230
rect 9055 8200 9060 8230
rect 9020 8195 9060 8200
rect 9020 8160 9060 8165
rect 9020 8130 9025 8160
rect 9025 8130 9055 8160
rect 9055 8130 9060 8160
rect 9020 8125 9060 8130
rect 9020 8095 9060 8100
rect 9020 8065 9025 8095
rect 9025 8065 9055 8095
rect 9055 8065 9060 8095
rect 9020 8060 9060 8065
rect 9020 8035 9060 8040
rect 9020 8005 9025 8035
rect 9025 8005 9055 8035
rect 9055 8005 9060 8035
rect 9020 8000 9060 8005
rect 9020 7970 9060 7975
rect 9020 7940 9025 7970
rect 9025 7940 9055 7970
rect 9055 7940 9060 7970
rect 9020 7935 9060 7940
rect 9020 7900 9060 7905
rect 9020 7870 9025 7900
rect 9025 7870 9055 7900
rect 9055 7870 9060 7900
rect 9020 7865 9060 7870
rect 9020 7830 9060 7835
rect 9020 7800 9025 7830
rect 9025 7800 9055 7830
rect 9055 7800 9060 7830
rect 9020 7795 9060 7800
rect 9020 7760 9060 7765
rect 9020 7730 9025 7760
rect 9025 7730 9055 7760
rect 9055 7730 9060 7760
rect 9020 7725 9060 7730
rect 9020 7695 9060 7700
rect 9020 7665 9025 7695
rect 9025 7665 9055 7695
rect 9055 7665 9060 7695
rect 9020 7660 9060 7665
rect 9020 7635 9060 7640
rect 9020 7605 9025 7635
rect 9025 7605 9055 7635
rect 9055 7605 9060 7635
rect 9020 7600 9060 7605
rect 9020 7570 9060 7575
rect 9020 7540 9025 7570
rect 9025 7540 9055 7570
rect 9055 7540 9060 7570
rect 9020 7535 9060 7540
rect 9020 7500 9060 7505
rect 9020 7470 9025 7500
rect 9025 7470 9055 7500
rect 9055 7470 9060 7500
rect 9020 7465 9060 7470
rect 9020 7430 9060 7435
rect 9020 7400 9025 7430
rect 9025 7400 9055 7430
rect 9055 7400 9060 7430
rect 9020 7395 9060 7400
rect 9020 7360 9060 7365
rect 9020 7330 9025 7360
rect 9025 7330 9055 7360
rect 9055 7330 9060 7360
rect 9020 7325 9060 7330
rect 9020 7295 9060 7300
rect 9020 7265 9025 7295
rect 9025 7265 9055 7295
rect 9055 7265 9060 7295
rect 9020 7260 9060 7265
rect 9020 7235 9060 7240
rect 9020 7205 9025 7235
rect 9025 7205 9055 7235
rect 9055 7205 9060 7235
rect 9020 7200 9060 7205
rect 9020 7170 9060 7175
rect 9020 7140 9025 7170
rect 9025 7140 9055 7170
rect 9055 7140 9060 7170
rect 9020 7135 9060 7140
rect 9020 7100 9060 7105
rect 9020 7070 9025 7100
rect 9025 7070 9055 7100
rect 9055 7070 9060 7100
rect 9020 7065 9060 7070
rect 9020 7030 9060 7035
rect 9020 7000 9025 7030
rect 9025 7000 9055 7030
rect 9055 7000 9060 7030
rect 9020 6995 9060 7000
rect 9020 6960 9060 6965
rect 9020 6930 9025 6960
rect 9025 6930 9055 6960
rect 9055 6930 9060 6960
rect 9020 6925 9060 6930
rect 9020 6895 9060 6900
rect 9020 6865 9025 6895
rect 9025 6865 9055 6895
rect 9055 6865 9060 6895
rect 9020 6860 9060 6865
rect 9020 6835 9060 6840
rect 9020 6805 9025 6835
rect 9025 6805 9055 6835
rect 9055 6805 9060 6835
rect 9020 6800 9060 6805
rect 9020 6770 9060 6775
rect 9020 6740 9025 6770
rect 9025 6740 9055 6770
rect 9055 6740 9060 6770
rect 9020 6735 9060 6740
rect 9020 6700 9060 6705
rect 9020 6670 9025 6700
rect 9025 6670 9055 6700
rect 9055 6670 9060 6700
rect 9020 6665 9060 6670
rect 9020 6630 9060 6635
rect 9020 6600 9025 6630
rect 9025 6600 9055 6630
rect 9055 6600 9060 6630
rect 9020 6595 9060 6600
rect 9020 6560 9060 6565
rect 9020 6530 9025 6560
rect 9025 6530 9055 6560
rect 9055 6530 9060 6560
rect 9020 6525 9060 6530
rect 9020 6495 9060 6500
rect 9020 6465 9025 6495
rect 9025 6465 9055 6495
rect 9055 6465 9060 6495
rect 9020 6460 9060 6465
rect 12925 9565 12975 9615
rect 13020 9565 13070 9615
rect 13115 9565 13165 9615
rect 13215 9565 13265 9615
rect 13315 9565 13365 9615
rect 13415 9565 13465 9615
rect 13510 9565 13560 9615
rect 13605 9565 13655 9615
rect 13725 9565 13775 9615
rect 13820 9565 13870 9615
rect 13915 9565 13965 9615
rect 14015 9565 14065 9615
rect 14115 9565 14165 9615
rect 14215 9565 14265 9615
rect 14310 9565 14360 9615
rect 14405 9565 14455 9615
rect 14525 9565 14575 9615
rect 14620 9565 14670 9615
rect 14715 9565 14765 9615
rect 14815 9565 14865 9615
rect 14915 9565 14965 9615
rect 15015 9565 15065 9615
rect 15110 9565 15160 9615
rect 15205 9565 15255 9615
rect 15325 9565 15375 9615
rect 15420 9565 15470 9615
rect 15515 9565 15565 9615
rect 15615 9565 15665 9615
rect 15715 9565 15765 9615
rect 15815 9565 15865 9615
rect 15910 9565 15960 9615
rect 16005 9565 16055 9615
rect 12925 9475 12975 9525
rect 13020 9475 13070 9525
rect 13115 9475 13165 9525
rect 13215 9475 13265 9525
rect 13315 9475 13365 9525
rect 13415 9475 13465 9525
rect 13510 9475 13560 9525
rect 13605 9475 13655 9525
rect 13725 9475 13775 9525
rect 13820 9475 13870 9525
rect 13915 9475 13965 9525
rect 14015 9475 14065 9525
rect 14115 9475 14165 9525
rect 14215 9475 14265 9525
rect 14310 9475 14360 9525
rect 14405 9475 14455 9525
rect 14525 9475 14575 9525
rect 14620 9475 14670 9525
rect 14715 9475 14765 9525
rect 14815 9475 14865 9525
rect 14915 9475 14965 9525
rect 15015 9475 15065 9525
rect 15110 9475 15160 9525
rect 15205 9475 15255 9525
rect 15325 9475 15375 9525
rect 15420 9475 15470 9525
rect 15515 9475 15565 9525
rect 15615 9475 15665 9525
rect 15715 9475 15765 9525
rect 15815 9475 15865 9525
rect 15910 9475 15960 9525
rect 16005 9475 16055 9525
rect 12925 9375 12975 9425
rect 13020 9375 13070 9425
rect 13115 9375 13165 9425
rect 13215 9375 13265 9425
rect 13315 9375 13365 9425
rect 13415 9375 13465 9425
rect 13510 9375 13560 9425
rect 13605 9375 13655 9425
rect 13725 9375 13775 9425
rect 13820 9375 13870 9425
rect 13915 9375 13965 9425
rect 14015 9375 14065 9425
rect 14115 9375 14165 9425
rect 14215 9375 14265 9425
rect 14310 9375 14360 9425
rect 14405 9375 14455 9425
rect 14525 9375 14575 9425
rect 14620 9375 14670 9425
rect 14715 9375 14765 9425
rect 14815 9375 14865 9425
rect 14915 9375 14965 9425
rect 15015 9375 15065 9425
rect 15110 9375 15160 9425
rect 15205 9375 15255 9425
rect 15325 9375 15375 9425
rect 15420 9375 15470 9425
rect 15515 9375 15565 9425
rect 15615 9375 15665 9425
rect 15715 9375 15765 9425
rect 15815 9375 15865 9425
rect 15910 9375 15960 9425
rect 16005 9375 16055 9425
rect 12925 9285 12975 9335
rect 13020 9285 13070 9335
rect 13115 9285 13165 9335
rect 13215 9285 13265 9335
rect 13315 9285 13365 9335
rect 13415 9285 13465 9335
rect 13510 9285 13560 9335
rect 13605 9285 13655 9335
rect 13725 9285 13775 9335
rect 13820 9285 13870 9335
rect 13915 9285 13965 9335
rect 14015 9285 14065 9335
rect 14115 9285 14165 9335
rect 14215 9285 14265 9335
rect 14310 9285 14360 9335
rect 14405 9285 14455 9335
rect 14525 9285 14575 9335
rect 14620 9285 14670 9335
rect 14715 9285 14765 9335
rect 14815 9285 14865 9335
rect 14915 9285 14965 9335
rect 15015 9285 15065 9335
rect 15110 9285 15160 9335
rect 15205 9285 15255 9335
rect 15325 9285 15375 9335
rect 15420 9285 15470 9335
rect 15515 9285 15565 9335
rect 15615 9285 15665 9335
rect 15715 9285 15765 9335
rect 15815 9285 15865 9335
rect 15910 9285 15960 9335
rect 16005 9285 16055 9335
rect 12925 9165 12975 9215
rect 13020 9165 13070 9215
rect 13115 9165 13165 9215
rect 13215 9165 13265 9215
rect 13315 9165 13365 9215
rect 13415 9165 13465 9215
rect 13510 9165 13560 9215
rect 13605 9165 13655 9215
rect 13725 9165 13775 9215
rect 13820 9165 13870 9215
rect 13915 9165 13965 9215
rect 14015 9165 14065 9215
rect 14115 9165 14165 9215
rect 14215 9165 14265 9215
rect 14310 9165 14360 9215
rect 14405 9165 14455 9215
rect 14525 9165 14575 9215
rect 14620 9165 14670 9215
rect 14715 9165 14765 9215
rect 14815 9165 14865 9215
rect 14915 9165 14965 9215
rect 15015 9165 15065 9215
rect 15110 9165 15160 9215
rect 15205 9165 15255 9215
rect 15325 9165 15375 9215
rect 15420 9165 15470 9215
rect 15515 9165 15565 9215
rect 15615 9165 15665 9215
rect 15715 9165 15765 9215
rect 15815 9165 15865 9215
rect 15910 9165 15960 9215
rect 16005 9165 16055 9215
rect 12925 9075 12975 9125
rect 13020 9075 13070 9125
rect 13115 9075 13165 9125
rect 13215 9075 13265 9125
rect 13315 9075 13365 9125
rect 13415 9075 13465 9125
rect 13510 9075 13560 9125
rect 13605 9075 13655 9125
rect 13725 9075 13775 9125
rect 13820 9075 13870 9125
rect 13915 9075 13965 9125
rect 14015 9075 14065 9125
rect 14115 9075 14165 9125
rect 14215 9075 14265 9125
rect 14310 9075 14360 9125
rect 14405 9075 14455 9125
rect 14525 9075 14575 9125
rect 14620 9075 14670 9125
rect 14715 9075 14765 9125
rect 14815 9075 14865 9125
rect 14915 9075 14965 9125
rect 15015 9075 15065 9125
rect 15110 9075 15160 9125
rect 15205 9075 15255 9125
rect 15325 9075 15375 9125
rect 15420 9075 15470 9125
rect 15515 9075 15565 9125
rect 15615 9075 15665 9125
rect 15715 9075 15765 9125
rect 15815 9075 15865 9125
rect 15910 9075 15960 9125
rect 16005 9075 16055 9125
rect 12925 8975 12975 9025
rect 13020 8975 13070 9025
rect 13115 8975 13165 9025
rect 13215 8975 13265 9025
rect 13315 8975 13365 9025
rect 13415 8975 13465 9025
rect 13510 8975 13560 9025
rect 13605 8975 13655 9025
rect 13725 8975 13775 9025
rect 13820 8975 13870 9025
rect 13915 8975 13965 9025
rect 14015 8975 14065 9025
rect 14115 8975 14165 9025
rect 14215 8975 14265 9025
rect 14310 8975 14360 9025
rect 14405 8975 14455 9025
rect 14525 8975 14575 9025
rect 14620 8975 14670 9025
rect 14715 8975 14765 9025
rect 14815 8975 14865 9025
rect 14915 8975 14965 9025
rect 15015 8975 15065 9025
rect 15110 8975 15160 9025
rect 15205 8975 15255 9025
rect 15325 8975 15375 9025
rect 15420 8975 15470 9025
rect 15515 8975 15565 9025
rect 15615 8975 15665 9025
rect 15715 8975 15765 9025
rect 15815 8975 15865 9025
rect 15910 8975 15960 9025
rect 16005 8975 16055 9025
rect 12925 8885 12975 8935
rect 13020 8885 13070 8935
rect 13115 8885 13165 8935
rect 13215 8885 13265 8935
rect 13315 8885 13365 8935
rect 13415 8885 13465 8935
rect 13510 8885 13560 8935
rect 13605 8885 13655 8935
rect 13725 8885 13775 8935
rect 13820 8885 13870 8935
rect 13915 8885 13965 8935
rect 14015 8885 14065 8935
rect 14115 8885 14165 8935
rect 14215 8885 14265 8935
rect 14310 8885 14360 8935
rect 14405 8885 14455 8935
rect 14525 8885 14575 8935
rect 14620 8885 14670 8935
rect 14715 8885 14765 8935
rect 14815 8885 14865 8935
rect 14915 8885 14965 8935
rect 15015 8885 15065 8935
rect 15110 8885 15160 8935
rect 15205 8885 15255 8935
rect 15325 8885 15375 8935
rect 15420 8885 15470 8935
rect 15515 8885 15565 8935
rect 15615 8885 15665 8935
rect 15715 8885 15765 8935
rect 15815 8885 15865 8935
rect 15910 8885 15960 8935
rect 16005 8885 16055 8935
rect 12925 8765 12975 8815
rect 13020 8765 13070 8815
rect 13115 8765 13165 8815
rect 13215 8765 13265 8815
rect 13315 8765 13365 8815
rect 13415 8765 13465 8815
rect 13510 8765 13560 8815
rect 13605 8765 13655 8815
rect 13725 8765 13775 8815
rect 13820 8765 13870 8815
rect 13915 8765 13965 8815
rect 14015 8765 14065 8815
rect 14115 8765 14165 8815
rect 14215 8765 14265 8815
rect 14310 8765 14360 8815
rect 14405 8765 14455 8815
rect 14525 8765 14575 8815
rect 14620 8765 14670 8815
rect 14715 8765 14765 8815
rect 14815 8765 14865 8815
rect 14915 8765 14965 8815
rect 15015 8765 15065 8815
rect 15110 8765 15160 8815
rect 15205 8765 15255 8815
rect 15325 8765 15375 8815
rect 15420 8765 15470 8815
rect 15515 8765 15565 8815
rect 15615 8765 15665 8815
rect 15715 8765 15765 8815
rect 15815 8765 15865 8815
rect 15910 8765 15960 8815
rect 16005 8765 16055 8815
rect 12925 8675 12975 8725
rect 13020 8675 13070 8725
rect 13115 8675 13165 8725
rect 13215 8675 13265 8725
rect 13315 8675 13365 8725
rect 13415 8675 13465 8725
rect 13510 8675 13560 8725
rect 13605 8675 13655 8725
rect 13725 8675 13775 8725
rect 13820 8675 13870 8725
rect 13915 8675 13965 8725
rect 14015 8675 14065 8725
rect 14115 8675 14165 8725
rect 14215 8675 14265 8725
rect 14310 8675 14360 8725
rect 14405 8675 14455 8725
rect 14525 8675 14575 8725
rect 14620 8675 14670 8725
rect 14715 8675 14765 8725
rect 14815 8675 14865 8725
rect 14915 8675 14965 8725
rect 15015 8675 15065 8725
rect 15110 8675 15160 8725
rect 15205 8675 15255 8725
rect 15325 8675 15375 8725
rect 15420 8675 15470 8725
rect 15515 8675 15565 8725
rect 15615 8675 15665 8725
rect 15715 8675 15765 8725
rect 15815 8675 15865 8725
rect 15910 8675 15960 8725
rect 16005 8675 16055 8725
rect 12925 8575 12975 8625
rect 13020 8575 13070 8625
rect 13115 8575 13165 8625
rect 13215 8575 13265 8625
rect 13315 8575 13365 8625
rect 13415 8575 13465 8625
rect 13510 8575 13560 8625
rect 13605 8575 13655 8625
rect 13725 8575 13775 8625
rect 13820 8575 13870 8625
rect 13915 8575 13965 8625
rect 14015 8575 14065 8625
rect 14115 8575 14165 8625
rect 14215 8575 14265 8625
rect 14310 8575 14360 8625
rect 14405 8575 14455 8625
rect 14525 8575 14575 8625
rect 14620 8575 14670 8625
rect 14715 8575 14765 8625
rect 14815 8575 14865 8625
rect 14915 8575 14965 8625
rect 15015 8575 15065 8625
rect 15110 8575 15160 8625
rect 15205 8575 15255 8625
rect 15325 8575 15375 8625
rect 15420 8575 15470 8625
rect 15515 8575 15565 8625
rect 15615 8575 15665 8625
rect 15715 8575 15765 8625
rect 15815 8575 15865 8625
rect 15910 8575 15960 8625
rect 16005 8575 16055 8625
rect 12925 8485 12975 8535
rect 13020 8485 13070 8535
rect 13115 8485 13165 8535
rect 13215 8485 13265 8535
rect 13315 8485 13365 8535
rect 13415 8485 13465 8535
rect 13510 8485 13560 8535
rect 13605 8485 13655 8535
rect 13725 8485 13775 8535
rect 13820 8485 13870 8535
rect 13915 8485 13965 8535
rect 14015 8485 14065 8535
rect 14115 8485 14165 8535
rect 14215 8485 14265 8535
rect 14310 8485 14360 8535
rect 14405 8485 14455 8535
rect 14525 8485 14575 8535
rect 14620 8485 14670 8535
rect 14715 8485 14765 8535
rect 14815 8485 14865 8535
rect 14915 8485 14965 8535
rect 15015 8485 15065 8535
rect 15110 8485 15160 8535
rect 15205 8485 15255 8535
rect 15325 8485 15375 8535
rect 15420 8485 15470 8535
rect 15515 8485 15565 8535
rect 15615 8485 15665 8535
rect 15715 8485 15765 8535
rect 15815 8485 15865 8535
rect 15910 8485 15960 8535
rect 16005 8485 16055 8535
rect 12925 8365 12975 8415
rect 13020 8365 13070 8415
rect 13115 8365 13165 8415
rect 13215 8365 13265 8415
rect 13315 8365 13365 8415
rect 13415 8365 13465 8415
rect 13510 8365 13560 8415
rect 13605 8365 13655 8415
rect 13725 8365 13775 8415
rect 13820 8365 13870 8415
rect 13915 8365 13965 8415
rect 14015 8365 14065 8415
rect 14115 8365 14165 8415
rect 14215 8365 14265 8415
rect 14310 8365 14360 8415
rect 14405 8365 14455 8415
rect 14525 8365 14575 8415
rect 14620 8365 14670 8415
rect 14715 8365 14765 8415
rect 14815 8365 14865 8415
rect 14915 8365 14965 8415
rect 15015 8365 15065 8415
rect 15110 8365 15160 8415
rect 15205 8365 15255 8415
rect 15325 8365 15375 8415
rect 15420 8365 15470 8415
rect 15515 8365 15565 8415
rect 15615 8365 15665 8415
rect 15715 8365 15765 8415
rect 15815 8365 15865 8415
rect 15910 8365 15960 8415
rect 16005 8365 16055 8415
rect 12925 8275 12975 8325
rect 13020 8275 13070 8325
rect 13115 8275 13165 8325
rect 13215 8275 13265 8325
rect 13315 8275 13365 8325
rect 13415 8275 13465 8325
rect 13510 8275 13560 8325
rect 13605 8275 13655 8325
rect 13725 8275 13775 8325
rect 13820 8275 13870 8325
rect 13915 8275 13965 8325
rect 14015 8275 14065 8325
rect 14115 8275 14165 8325
rect 14215 8275 14265 8325
rect 14310 8275 14360 8325
rect 14405 8275 14455 8325
rect 14525 8275 14575 8325
rect 14620 8275 14670 8325
rect 14715 8275 14765 8325
rect 14815 8275 14865 8325
rect 14915 8275 14965 8325
rect 15015 8275 15065 8325
rect 15110 8275 15160 8325
rect 15205 8275 15255 8325
rect 15325 8275 15375 8325
rect 15420 8275 15470 8325
rect 15515 8275 15565 8325
rect 15615 8275 15665 8325
rect 15715 8275 15765 8325
rect 15815 8275 15865 8325
rect 15910 8275 15960 8325
rect 16005 8275 16055 8325
rect 12925 8175 12975 8225
rect 13020 8175 13070 8225
rect 13115 8175 13165 8225
rect 13215 8175 13265 8225
rect 13315 8175 13365 8225
rect 13415 8175 13465 8225
rect 13510 8175 13560 8225
rect 13605 8175 13655 8225
rect 13725 8175 13775 8225
rect 13820 8175 13870 8225
rect 13915 8175 13965 8225
rect 14015 8175 14065 8225
rect 14115 8175 14165 8225
rect 14215 8175 14265 8225
rect 14310 8175 14360 8225
rect 14405 8175 14455 8225
rect 14525 8175 14575 8225
rect 14620 8175 14670 8225
rect 14715 8175 14765 8225
rect 14815 8175 14865 8225
rect 14915 8175 14965 8225
rect 15015 8175 15065 8225
rect 15110 8175 15160 8225
rect 15205 8175 15255 8225
rect 15325 8175 15375 8225
rect 15420 8175 15470 8225
rect 15515 8175 15565 8225
rect 15615 8175 15665 8225
rect 15715 8175 15765 8225
rect 15815 8175 15865 8225
rect 15910 8175 15960 8225
rect 16005 8175 16055 8225
rect 12925 8085 12975 8135
rect 13020 8085 13070 8135
rect 13115 8085 13165 8135
rect 13215 8085 13265 8135
rect 13315 8085 13365 8135
rect 13415 8085 13465 8135
rect 13510 8085 13560 8135
rect 13605 8085 13655 8135
rect 13725 8085 13775 8135
rect 13820 8085 13870 8135
rect 13915 8085 13965 8135
rect 14015 8085 14065 8135
rect 14115 8085 14165 8135
rect 14215 8085 14265 8135
rect 14310 8085 14360 8135
rect 14405 8085 14455 8135
rect 14525 8085 14575 8135
rect 14620 8085 14670 8135
rect 14715 8085 14765 8135
rect 14815 8085 14865 8135
rect 14915 8085 14965 8135
rect 15015 8085 15065 8135
rect 15110 8085 15160 8135
rect 15205 8085 15255 8135
rect 15325 8085 15375 8135
rect 15420 8085 15470 8135
rect 15515 8085 15565 8135
rect 15615 8085 15665 8135
rect 15715 8085 15765 8135
rect 15815 8085 15865 8135
rect 15910 8085 15960 8135
rect 16005 8085 16055 8135
rect 12925 7965 12975 8015
rect 13020 7965 13070 8015
rect 13115 7965 13165 8015
rect 13215 7965 13265 8015
rect 13315 7965 13365 8015
rect 13415 7965 13465 8015
rect 13510 7965 13560 8015
rect 13605 7965 13655 8015
rect 13725 7965 13775 8015
rect 13820 7965 13870 8015
rect 13915 7965 13965 8015
rect 14015 7965 14065 8015
rect 14115 7965 14165 8015
rect 14215 7965 14265 8015
rect 14310 7965 14360 8015
rect 14405 7965 14455 8015
rect 14525 7965 14575 8015
rect 14620 7965 14670 8015
rect 14715 7965 14765 8015
rect 14815 7965 14865 8015
rect 14915 7965 14965 8015
rect 15015 7965 15065 8015
rect 15110 7965 15160 8015
rect 15205 7965 15255 8015
rect 15325 7965 15375 8015
rect 15420 7965 15470 8015
rect 15515 7965 15565 8015
rect 15615 7965 15665 8015
rect 15715 7965 15765 8015
rect 15815 7965 15865 8015
rect 15910 7965 15960 8015
rect 16005 7965 16055 8015
rect 12925 7875 12975 7925
rect 13020 7875 13070 7925
rect 13115 7875 13165 7925
rect 13215 7875 13265 7925
rect 13315 7875 13365 7925
rect 13415 7875 13465 7925
rect 13510 7875 13560 7925
rect 13605 7875 13655 7925
rect 13725 7875 13775 7925
rect 13820 7875 13870 7925
rect 13915 7875 13965 7925
rect 14015 7875 14065 7925
rect 14115 7875 14165 7925
rect 14215 7875 14265 7925
rect 14310 7875 14360 7925
rect 14405 7875 14455 7925
rect 14525 7875 14575 7925
rect 14620 7875 14670 7925
rect 14715 7875 14765 7925
rect 14815 7875 14865 7925
rect 14915 7875 14965 7925
rect 15015 7875 15065 7925
rect 15110 7875 15160 7925
rect 15205 7875 15255 7925
rect 15325 7875 15375 7925
rect 15420 7875 15470 7925
rect 15515 7875 15565 7925
rect 15615 7875 15665 7925
rect 15715 7875 15765 7925
rect 15815 7875 15865 7925
rect 15910 7875 15960 7925
rect 16005 7875 16055 7925
rect 12925 7775 12975 7825
rect 13020 7775 13070 7825
rect 13115 7775 13165 7825
rect 13215 7775 13265 7825
rect 13315 7775 13365 7825
rect 13415 7775 13465 7825
rect 13510 7775 13560 7825
rect 13605 7775 13655 7825
rect 13725 7775 13775 7825
rect 13820 7775 13870 7825
rect 13915 7775 13965 7825
rect 14015 7775 14065 7825
rect 14115 7775 14165 7825
rect 14215 7775 14265 7825
rect 14310 7775 14360 7825
rect 14405 7775 14455 7825
rect 14525 7775 14575 7825
rect 14620 7775 14670 7825
rect 14715 7775 14765 7825
rect 14815 7775 14865 7825
rect 14915 7775 14965 7825
rect 15015 7775 15065 7825
rect 15110 7775 15160 7825
rect 15205 7775 15255 7825
rect 15325 7775 15375 7825
rect 15420 7775 15470 7825
rect 15515 7775 15565 7825
rect 15615 7775 15665 7825
rect 15715 7775 15765 7825
rect 15815 7775 15865 7825
rect 15910 7775 15960 7825
rect 16005 7775 16055 7825
rect 12925 7685 12975 7735
rect 13020 7685 13070 7735
rect 13115 7685 13165 7735
rect 13215 7685 13265 7735
rect 13315 7685 13365 7735
rect 13415 7685 13465 7735
rect 13510 7685 13560 7735
rect 13605 7685 13655 7735
rect 13725 7685 13775 7735
rect 13820 7685 13870 7735
rect 13915 7685 13965 7735
rect 14015 7685 14065 7735
rect 14115 7685 14165 7735
rect 14215 7685 14265 7735
rect 14310 7685 14360 7735
rect 14405 7685 14455 7735
rect 14525 7685 14575 7735
rect 14620 7685 14670 7735
rect 14715 7685 14765 7735
rect 14815 7685 14865 7735
rect 14915 7685 14965 7735
rect 15015 7685 15065 7735
rect 15110 7685 15160 7735
rect 15205 7685 15255 7735
rect 15325 7685 15375 7735
rect 15420 7685 15470 7735
rect 15515 7685 15565 7735
rect 15615 7685 15665 7735
rect 15715 7685 15765 7735
rect 15815 7685 15865 7735
rect 15910 7685 15960 7735
rect 16005 7685 16055 7735
rect 12925 7565 12975 7615
rect 13020 7565 13070 7615
rect 13115 7565 13165 7615
rect 13215 7565 13265 7615
rect 13315 7565 13365 7615
rect 13415 7565 13465 7615
rect 13510 7565 13560 7615
rect 13605 7565 13655 7615
rect 13725 7565 13775 7615
rect 13820 7565 13870 7615
rect 13915 7565 13965 7615
rect 14015 7565 14065 7615
rect 14115 7565 14165 7615
rect 14215 7565 14265 7615
rect 14310 7565 14360 7615
rect 14405 7565 14455 7615
rect 14525 7565 14575 7615
rect 14620 7565 14670 7615
rect 14715 7565 14765 7615
rect 14815 7565 14865 7615
rect 14915 7565 14965 7615
rect 15015 7565 15065 7615
rect 15110 7565 15160 7615
rect 15205 7565 15255 7615
rect 15325 7565 15375 7615
rect 15420 7565 15470 7615
rect 15515 7565 15565 7615
rect 15615 7565 15665 7615
rect 15715 7565 15765 7615
rect 15815 7565 15865 7615
rect 15910 7565 15960 7615
rect 16005 7565 16055 7615
rect 12925 7475 12975 7525
rect 13020 7475 13070 7525
rect 13115 7475 13165 7525
rect 13215 7475 13265 7525
rect 13315 7475 13365 7525
rect 13415 7475 13465 7525
rect 13510 7475 13560 7525
rect 13605 7475 13655 7525
rect 13725 7475 13775 7525
rect 13820 7475 13870 7525
rect 13915 7475 13965 7525
rect 14015 7475 14065 7525
rect 14115 7475 14165 7525
rect 14215 7475 14265 7525
rect 14310 7475 14360 7525
rect 14405 7475 14455 7525
rect 14525 7475 14575 7525
rect 14620 7475 14670 7525
rect 14715 7475 14765 7525
rect 14815 7475 14865 7525
rect 14915 7475 14965 7525
rect 15015 7475 15065 7525
rect 15110 7475 15160 7525
rect 15205 7475 15255 7525
rect 15325 7475 15375 7525
rect 15420 7475 15470 7525
rect 15515 7475 15565 7525
rect 15615 7475 15665 7525
rect 15715 7475 15765 7525
rect 15815 7475 15865 7525
rect 15910 7475 15960 7525
rect 16005 7475 16055 7525
rect 12925 7375 12975 7425
rect 13020 7375 13070 7425
rect 13115 7375 13165 7425
rect 13215 7375 13265 7425
rect 13315 7375 13365 7425
rect 13415 7375 13465 7425
rect 13510 7375 13560 7425
rect 13605 7375 13655 7425
rect 13725 7375 13775 7425
rect 13820 7375 13870 7425
rect 13915 7375 13965 7425
rect 14015 7375 14065 7425
rect 14115 7375 14165 7425
rect 14215 7375 14265 7425
rect 14310 7375 14360 7425
rect 14405 7375 14455 7425
rect 14525 7375 14575 7425
rect 14620 7375 14670 7425
rect 14715 7375 14765 7425
rect 14815 7375 14865 7425
rect 14915 7375 14965 7425
rect 15015 7375 15065 7425
rect 15110 7375 15160 7425
rect 15205 7375 15255 7425
rect 15325 7375 15375 7425
rect 15420 7375 15470 7425
rect 15515 7375 15565 7425
rect 15615 7375 15665 7425
rect 15715 7375 15765 7425
rect 15815 7375 15865 7425
rect 15910 7375 15960 7425
rect 16005 7375 16055 7425
rect 12925 7285 12975 7335
rect 13020 7285 13070 7335
rect 13115 7285 13165 7335
rect 13215 7285 13265 7335
rect 13315 7285 13365 7335
rect 13415 7285 13465 7335
rect 13510 7285 13560 7335
rect 13605 7285 13655 7335
rect 13725 7285 13775 7335
rect 13820 7285 13870 7335
rect 13915 7285 13965 7335
rect 14015 7285 14065 7335
rect 14115 7285 14165 7335
rect 14215 7285 14265 7335
rect 14310 7285 14360 7335
rect 14405 7285 14455 7335
rect 14525 7285 14575 7335
rect 14620 7285 14670 7335
rect 14715 7285 14765 7335
rect 14815 7285 14865 7335
rect 14915 7285 14965 7335
rect 15015 7285 15065 7335
rect 15110 7285 15160 7335
rect 15205 7285 15255 7335
rect 15325 7285 15375 7335
rect 15420 7285 15470 7335
rect 15515 7285 15565 7335
rect 15615 7285 15665 7335
rect 15715 7285 15765 7335
rect 15815 7285 15865 7335
rect 15910 7285 15960 7335
rect 16005 7285 16055 7335
rect 12925 7165 12975 7215
rect 13020 7165 13070 7215
rect 13115 7165 13165 7215
rect 13215 7165 13265 7215
rect 13315 7165 13365 7215
rect 13415 7165 13465 7215
rect 13510 7165 13560 7215
rect 13605 7165 13655 7215
rect 13725 7165 13775 7215
rect 13820 7165 13870 7215
rect 13915 7165 13965 7215
rect 14015 7165 14065 7215
rect 14115 7165 14165 7215
rect 14215 7165 14265 7215
rect 14310 7165 14360 7215
rect 14405 7165 14455 7215
rect 14525 7165 14575 7215
rect 14620 7165 14670 7215
rect 14715 7165 14765 7215
rect 14815 7165 14865 7215
rect 14915 7165 14965 7215
rect 15015 7165 15065 7215
rect 15110 7165 15160 7215
rect 15205 7165 15255 7215
rect 15325 7165 15375 7215
rect 15420 7165 15470 7215
rect 15515 7165 15565 7215
rect 15615 7165 15665 7215
rect 15715 7165 15765 7215
rect 15815 7165 15865 7215
rect 15910 7165 15960 7215
rect 16005 7165 16055 7215
rect 12925 7075 12975 7125
rect 13020 7075 13070 7125
rect 13115 7075 13165 7125
rect 13215 7075 13265 7125
rect 13315 7075 13365 7125
rect 13415 7075 13465 7125
rect 13510 7075 13560 7125
rect 13605 7075 13655 7125
rect 13725 7075 13775 7125
rect 13820 7075 13870 7125
rect 13915 7075 13965 7125
rect 14015 7075 14065 7125
rect 14115 7075 14165 7125
rect 14215 7075 14265 7125
rect 14310 7075 14360 7125
rect 14405 7075 14455 7125
rect 14525 7075 14575 7125
rect 14620 7075 14670 7125
rect 14715 7075 14765 7125
rect 14815 7075 14865 7125
rect 14915 7075 14965 7125
rect 15015 7075 15065 7125
rect 15110 7075 15160 7125
rect 15205 7075 15255 7125
rect 15325 7075 15375 7125
rect 15420 7075 15470 7125
rect 15515 7075 15565 7125
rect 15615 7075 15665 7125
rect 15715 7075 15765 7125
rect 15815 7075 15865 7125
rect 15910 7075 15960 7125
rect 16005 7075 16055 7125
rect 12925 6975 12975 7025
rect 13020 6975 13070 7025
rect 13115 6975 13165 7025
rect 13215 6975 13265 7025
rect 13315 6975 13365 7025
rect 13415 6975 13465 7025
rect 13510 6975 13560 7025
rect 13605 6975 13655 7025
rect 13725 6975 13775 7025
rect 13820 6975 13870 7025
rect 13915 6975 13965 7025
rect 14015 6975 14065 7025
rect 14115 6975 14165 7025
rect 14215 6975 14265 7025
rect 14310 6975 14360 7025
rect 14405 6975 14455 7025
rect 14525 6975 14575 7025
rect 14620 6975 14670 7025
rect 14715 6975 14765 7025
rect 14815 6975 14865 7025
rect 14915 6975 14965 7025
rect 15015 6975 15065 7025
rect 15110 6975 15160 7025
rect 15205 6975 15255 7025
rect 15325 6975 15375 7025
rect 15420 6975 15470 7025
rect 15515 6975 15565 7025
rect 15615 6975 15665 7025
rect 15715 6975 15765 7025
rect 15815 6975 15865 7025
rect 15910 6975 15960 7025
rect 16005 6975 16055 7025
rect 12925 6885 12975 6935
rect 13020 6885 13070 6935
rect 13115 6885 13165 6935
rect 13215 6885 13265 6935
rect 13315 6885 13365 6935
rect 13415 6885 13465 6935
rect 13510 6885 13560 6935
rect 13605 6885 13655 6935
rect 13725 6885 13775 6935
rect 13820 6885 13870 6935
rect 13915 6885 13965 6935
rect 14015 6885 14065 6935
rect 14115 6885 14165 6935
rect 14215 6885 14265 6935
rect 14310 6885 14360 6935
rect 14405 6885 14455 6935
rect 14525 6885 14575 6935
rect 14620 6885 14670 6935
rect 14715 6885 14765 6935
rect 14815 6885 14865 6935
rect 14915 6885 14965 6935
rect 15015 6885 15065 6935
rect 15110 6885 15160 6935
rect 15205 6885 15255 6935
rect 15325 6885 15375 6935
rect 15420 6885 15470 6935
rect 15515 6885 15565 6935
rect 15615 6885 15665 6935
rect 15715 6885 15765 6935
rect 15815 6885 15865 6935
rect 15910 6885 15960 6935
rect 16005 6885 16055 6935
rect 12925 6765 12975 6815
rect 13020 6765 13070 6815
rect 13115 6765 13165 6815
rect 13215 6765 13265 6815
rect 13315 6765 13365 6815
rect 13415 6765 13465 6815
rect 13510 6765 13560 6815
rect 13605 6765 13655 6815
rect 13725 6765 13775 6815
rect 13820 6765 13870 6815
rect 13915 6765 13965 6815
rect 14015 6765 14065 6815
rect 14115 6765 14165 6815
rect 14215 6765 14265 6815
rect 14310 6765 14360 6815
rect 14405 6765 14455 6815
rect 14525 6765 14575 6815
rect 14620 6765 14670 6815
rect 14715 6765 14765 6815
rect 14815 6765 14865 6815
rect 14915 6765 14965 6815
rect 15015 6765 15065 6815
rect 15110 6765 15160 6815
rect 15205 6765 15255 6815
rect 15325 6765 15375 6815
rect 15420 6765 15470 6815
rect 15515 6765 15565 6815
rect 15615 6765 15665 6815
rect 15715 6765 15765 6815
rect 15815 6765 15865 6815
rect 15910 6765 15960 6815
rect 16005 6765 16055 6815
rect 12925 6675 12975 6725
rect 13020 6675 13070 6725
rect 13115 6675 13165 6725
rect 13215 6675 13265 6725
rect 13315 6675 13365 6725
rect 13415 6675 13465 6725
rect 13510 6675 13560 6725
rect 13605 6675 13655 6725
rect 13725 6675 13775 6725
rect 13820 6675 13870 6725
rect 13915 6675 13965 6725
rect 14015 6675 14065 6725
rect 14115 6675 14165 6725
rect 14215 6675 14265 6725
rect 14310 6675 14360 6725
rect 14405 6675 14455 6725
rect 14525 6675 14575 6725
rect 14620 6675 14670 6725
rect 14715 6675 14765 6725
rect 14815 6675 14865 6725
rect 14915 6675 14965 6725
rect 15015 6675 15065 6725
rect 15110 6675 15160 6725
rect 15205 6675 15255 6725
rect 15325 6675 15375 6725
rect 15420 6675 15470 6725
rect 15515 6675 15565 6725
rect 15615 6675 15665 6725
rect 15715 6675 15765 6725
rect 15815 6675 15865 6725
rect 15910 6675 15960 6725
rect 16005 6675 16055 6725
rect 12925 6575 12975 6625
rect 13020 6575 13070 6625
rect 13115 6575 13165 6625
rect 13215 6575 13265 6625
rect 13315 6575 13365 6625
rect 13415 6575 13465 6625
rect 13510 6575 13560 6625
rect 13605 6575 13655 6625
rect 13725 6575 13775 6625
rect 13820 6575 13870 6625
rect 13915 6575 13965 6625
rect 14015 6575 14065 6625
rect 14115 6575 14165 6625
rect 14215 6575 14265 6625
rect 14310 6575 14360 6625
rect 14405 6575 14455 6625
rect 14525 6575 14575 6625
rect 14620 6575 14670 6625
rect 14715 6575 14765 6625
rect 14815 6575 14865 6625
rect 14915 6575 14965 6625
rect 15015 6575 15065 6625
rect 15110 6575 15160 6625
rect 15205 6575 15255 6625
rect 15325 6575 15375 6625
rect 15420 6575 15470 6625
rect 15515 6575 15565 6625
rect 15615 6575 15665 6625
rect 15715 6575 15765 6625
rect 15815 6575 15865 6625
rect 15910 6575 15960 6625
rect 16005 6575 16055 6625
rect 12925 6485 12975 6535
rect 13020 6485 13070 6535
rect 13115 6485 13165 6535
rect 13215 6485 13265 6535
rect 13315 6485 13365 6535
rect 13415 6485 13465 6535
rect 13510 6485 13560 6535
rect 13605 6485 13655 6535
rect 13725 6485 13775 6535
rect 13820 6485 13870 6535
rect 13915 6485 13965 6535
rect 14015 6485 14065 6535
rect 14115 6485 14165 6535
rect 14215 6485 14265 6535
rect 14310 6485 14360 6535
rect 14405 6485 14455 6535
rect 14525 6485 14575 6535
rect 14620 6485 14670 6535
rect 14715 6485 14765 6535
rect 14815 6485 14865 6535
rect 14915 6485 14965 6535
rect 15015 6485 15065 6535
rect 15110 6485 15160 6535
rect 15205 6485 15255 6535
rect 15325 6485 15375 6535
rect 15420 6485 15470 6535
rect 15515 6485 15565 6535
rect 15615 6485 15665 6535
rect 15715 6485 15765 6535
rect 15815 6485 15865 6535
rect 15910 6485 15960 6535
rect 16005 6485 16055 6535
rect -80 -1305 -40 -1300
rect -80 -1335 -75 -1305
rect -75 -1335 -45 -1305
rect -45 -1335 -40 -1305
rect -80 -1340 -40 -1335
rect -80 -1370 -40 -1365
rect -80 -1400 -75 -1370
rect -75 -1400 -45 -1370
rect -45 -1400 -40 -1370
rect -80 -1405 -40 -1400
rect -80 -1440 -40 -1435
rect -80 -1470 -75 -1440
rect -75 -1470 -45 -1440
rect -45 -1470 -40 -1440
rect -80 -1475 -40 -1470
rect -80 -1510 -40 -1505
rect -80 -1540 -75 -1510
rect -75 -1540 -45 -1510
rect -45 -1540 -40 -1510
rect -80 -1545 -40 -1540
rect -80 -1580 -40 -1575
rect -80 -1610 -75 -1580
rect -75 -1610 -45 -1580
rect -45 -1610 -40 -1580
rect -80 -1615 -40 -1610
rect -80 -1645 -40 -1640
rect -80 -1675 -75 -1645
rect -75 -1675 -45 -1645
rect -45 -1675 -40 -1645
rect -80 -1680 -40 -1675
rect -80 -1705 -40 -1700
rect -80 -1735 -75 -1705
rect -75 -1735 -45 -1705
rect -45 -1735 -40 -1705
rect -80 -1740 -40 -1735
rect -80 -1770 -40 -1765
rect -80 -1800 -75 -1770
rect -75 -1800 -45 -1770
rect -45 -1800 -40 -1770
rect -80 -1805 -40 -1800
rect -80 -1840 -40 -1835
rect -80 -1870 -75 -1840
rect -75 -1870 -45 -1840
rect -45 -1870 -40 -1840
rect -80 -1875 -40 -1870
rect -80 -1910 -40 -1905
rect -80 -1940 -75 -1910
rect -75 -1940 -45 -1910
rect -45 -1940 -40 -1910
rect -80 -1945 -40 -1940
rect -80 -1980 -40 -1975
rect -80 -2010 -75 -1980
rect -75 -2010 -45 -1980
rect -45 -2010 -40 -1980
rect -80 -2015 -40 -2010
rect -80 -2045 -40 -2040
rect -80 -2075 -75 -2045
rect -75 -2075 -45 -2045
rect -45 -2075 -40 -2045
rect -80 -2080 -40 -2075
rect -80 -2105 -40 -2100
rect -80 -2135 -75 -2105
rect -75 -2135 -45 -2105
rect -45 -2135 -40 -2105
rect -80 -2140 -40 -2135
rect -80 -2170 -40 -2165
rect -80 -2200 -75 -2170
rect -75 -2200 -45 -2170
rect -45 -2200 -40 -2170
rect -80 -2205 -40 -2200
rect -80 -2240 -40 -2235
rect -80 -2270 -75 -2240
rect -75 -2270 -45 -2240
rect -45 -2270 -40 -2240
rect -80 -2275 -40 -2270
rect -80 -2310 -40 -2305
rect -80 -2340 -75 -2310
rect -75 -2340 -45 -2310
rect -45 -2340 -40 -2310
rect -80 -2345 -40 -2340
rect -80 -2380 -40 -2375
rect -80 -2410 -75 -2380
rect -75 -2410 -45 -2380
rect -45 -2410 -40 -2380
rect -80 -2415 -40 -2410
rect -80 -2445 -40 -2440
rect -80 -2475 -75 -2445
rect -75 -2475 -45 -2445
rect -45 -2475 -40 -2445
rect -80 -2480 -40 -2475
rect -80 -2505 -40 -2500
rect -80 -2535 -75 -2505
rect -75 -2535 -45 -2505
rect -45 -2535 -40 -2505
rect -80 -2540 -40 -2535
rect -80 -2570 -40 -2565
rect -80 -2600 -75 -2570
rect -75 -2600 -45 -2570
rect -45 -2600 -40 -2570
rect -80 -2605 -40 -2600
rect -80 -2640 -40 -2635
rect -80 -2670 -75 -2640
rect -75 -2670 -45 -2640
rect -45 -2670 -40 -2640
rect -80 -2675 -40 -2670
rect -80 -2710 -40 -2705
rect -80 -2740 -75 -2710
rect -75 -2740 -45 -2710
rect -45 -2740 -40 -2710
rect -80 -2745 -40 -2740
rect -80 -2780 -40 -2775
rect -80 -2810 -75 -2780
rect -75 -2810 -45 -2780
rect -45 -2810 -40 -2780
rect -80 -2815 -40 -2810
rect -80 -2845 -40 -2840
rect -80 -2875 -75 -2845
rect -75 -2875 -45 -2845
rect -45 -2875 -40 -2845
rect -80 -2880 -40 -2875
rect -80 -2905 -40 -2900
rect -80 -2935 -75 -2905
rect -75 -2935 -45 -2905
rect -45 -2935 -40 -2905
rect -80 -2940 -40 -2935
rect -80 -2970 -40 -2965
rect -80 -3000 -75 -2970
rect -75 -3000 -45 -2970
rect -45 -3000 -40 -2970
rect -80 -3005 -40 -3000
rect -80 -3040 -40 -3035
rect -80 -3070 -75 -3040
rect -75 -3070 -45 -3040
rect -45 -3070 -40 -3040
rect -80 -3075 -40 -3070
rect -80 -3110 -40 -3105
rect -80 -3140 -75 -3110
rect -75 -3140 -45 -3110
rect -45 -3140 -40 -3110
rect -80 -3145 -40 -3140
rect -80 -3180 -40 -3175
rect -80 -3210 -75 -3180
rect -75 -3210 -45 -3180
rect -45 -3210 -40 -3180
rect -80 -3215 -40 -3210
rect -80 -3245 -40 -3240
rect -80 -3275 -75 -3245
rect -75 -3275 -45 -3245
rect -45 -3275 -40 -3245
rect -80 -3280 -40 -3275
rect -80 -3305 -40 -3300
rect -80 -3335 -75 -3305
rect -75 -3335 -45 -3305
rect -45 -3335 -40 -3305
rect -80 -3340 -40 -3335
rect -80 -3370 -40 -3365
rect -80 -3400 -75 -3370
rect -75 -3400 -45 -3370
rect -45 -3400 -40 -3370
rect -80 -3405 -40 -3400
rect -80 -3440 -40 -3435
rect -80 -3470 -75 -3440
rect -75 -3470 -45 -3440
rect -45 -3470 -40 -3440
rect -80 -3475 -40 -3470
rect -80 -3510 -40 -3505
rect -80 -3540 -75 -3510
rect -75 -3540 -45 -3510
rect -45 -3540 -40 -3510
rect -80 -3545 -40 -3540
rect -80 -3580 -40 -3575
rect -80 -3610 -75 -3580
rect -75 -3610 -45 -3580
rect -45 -3610 -40 -3580
rect -80 -3615 -40 -3610
rect -80 -3645 -40 -3640
rect -80 -3675 -75 -3645
rect -75 -3675 -45 -3645
rect -45 -3675 -40 -3645
rect -80 -3680 -40 -3675
rect -80 -3705 -40 -3700
rect -80 -3735 -75 -3705
rect -75 -3735 -45 -3705
rect -45 -3735 -40 -3705
rect -80 -3740 -40 -3735
rect -80 -3770 -40 -3765
rect -80 -3800 -75 -3770
rect -75 -3800 -45 -3770
rect -45 -3800 -40 -3770
rect -80 -3805 -40 -3800
rect -80 -3840 -40 -3835
rect -80 -3870 -75 -3840
rect -75 -3870 -45 -3840
rect -45 -3870 -40 -3840
rect -80 -3875 -40 -3870
rect -80 -3910 -40 -3905
rect -80 -3940 -75 -3910
rect -75 -3940 -45 -3910
rect -45 -3940 -40 -3910
rect -80 -3945 -40 -3940
rect -80 -3980 -40 -3975
rect -80 -4010 -75 -3980
rect -75 -4010 -45 -3980
rect -45 -4010 -40 -3980
rect -80 -4015 -40 -4010
rect -80 -4045 -40 -4040
rect -80 -4075 -75 -4045
rect -75 -4075 -45 -4045
rect -45 -4075 -40 -4045
rect -80 -4080 -40 -4075
rect -80 -4105 -40 -4100
rect -80 -4135 -75 -4105
rect -75 -4135 -45 -4105
rect -45 -4135 -40 -4105
rect -80 -4140 -40 -4135
rect -80 -4170 -40 -4165
rect -80 -4200 -75 -4170
rect -75 -4200 -45 -4170
rect -45 -4200 -40 -4170
rect -80 -4205 -40 -4200
rect -80 -4240 -40 -4235
rect -80 -4270 -75 -4240
rect -75 -4270 -45 -4240
rect -45 -4270 -40 -4240
rect -80 -4275 -40 -4270
rect -80 -4310 -40 -4305
rect -80 -4340 -75 -4310
rect -75 -4340 -45 -4310
rect -45 -4340 -40 -4310
rect -80 -4345 -40 -4340
rect -80 -4380 -40 -4375
rect -80 -4410 -75 -4380
rect -75 -4410 -45 -4380
rect -45 -4410 -40 -4380
rect -80 -4415 -40 -4410
rect -80 -4445 -40 -4440
rect -80 -4475 -75 -4445
rect -75 -4475 -45 -4445
rect -45 -4475 -40 -4445
rect -80 -4480 -40 -4475
rect 270 -1305 310 -1300
rect 270 -1335 275 -1305
rect 275 -1335 305 -1305
rect 305 -1335 310 -1305
rect 270 -1340 310 -1335
rect 270 -1370 310 -1365
rect 270 -1400 275 -1370
rect 275 -1400 305 -1370
rect 305 -1400 310 -1370
rect 270 -1405 310 -1400
rect 270 -1440 310 -1435
rect 270 -1470 275 -1440
rect 275 -1470 305 -1440
rect 305 -1470 310 -1440
rect 270 -1475 310 -1470
rect 270 -1510 310 -1505
rect 270 -1540 275 -1510
rect 275 -1540 305 -1510
rect 305 -1540 310 -1510
rect 270 -1545 310 -1540
rect 270 -1580 310 -1575
rect 270 -1610 275 -1580
rect 275 -1610 305 -1580
rect 305 -1610 310 -1580
rect 270 -1615 310 -1610
rect 270 -1645 310 -1640
rect 270 -1675 275 -1645
rect 275 -1675 305 -1645
rect 305 -1675 310 -1645
rect 270 -1680 310 -1675
rect 270 -1705 310 -1700
rect 270 -1735 275 -1705
rect 275 -1735 305 -1705
rect 305 -1735 310 -1705
rect 270 -1740 310 -1735
rect 270 -1770 310 -1765
rect 270 -1800 275 -1770
rect 275 -1800 305 -1770
rect 305 -1800 310 -1770
rect 270 -1805 310 -1800
rect 270 -1840 310 -1835
rect 270 -1870 275 -1840
rect 275 -1870 305 -1840
rect 305 -1870 310 -1840
rect 270 -1875 310 -1870
rect 270 -1910 310 -1905
rect 270 -1940 275 -1910
rect 275 -1940 305 -1910
rect 305 -1940 310 -1910
rect 270 -1945 310 -1940
rect 270 -1980 310 -1975
rect 270 -2010 275 -1980
rect 275 -2010 305 -1980
rect 305 -2010 310 -1980
rect 270 -2015 310 -2010
rect 270 -2045 310 -2040
rect 270 -2075 275 -2045
rect 275 -2075 305 -2045
rect 305 -2075 310 -2045
rect 270 -2080 310 -2075
rect 270 -2105 310 -2100
rect 270 -2135 275 -2105
rect 275 -2135 305 -2105
rect 305 -2135 310 -2105
rect 270 -2140 310 -2135
rect 270 -2170 310 -2165
rect 270 -2200 275 -2170
rect 275 -2200 305 -2170
rect 305 -2200 310 -2170
rect 270 -2205 310 -2200
rect 270 -2240 310 -2235
rect 270 -2270 275 -2240
rect 275 -2270 305 -2240
rect 305 -2270 310 -2240
rect 270 -2275 310 -2270
rect 270 -2310 310 -2305
rect 270 -2340 275 -2310
rect 275 -2340 305 -2310
rect 305 -2340 310 -2310
rect 270 -2345 310 -2340
rect 270 -2380 310 -2375
rect 270 -2410 275 -2380
rect 275 -2410 305 -2380
rect 305 -2410 310 -2380
rect 270 -2415 310 -2410
rect 270 -2445 310 -2440
rect 270 -2475 275 -2445
rect 275 -2475 305 -2445
rect 305 -2475 310 -2445
rect 270 -2480 310 -2475
rect 270 -2505 310 -2500
rect 270 -2535 275 -2505
rect 275 -2535 305 -2505
rect 305 -2535 310 -2505
rect 270 -2540 310 -2535
rect 270 -2570 310 -2565
rect 270 -2600 275 -2570
rect 275 -2600 305 -2570
rect 305 -2600 310 -2570
rect 270 -2605 310 -2600
rect 270 -2640 310 -2635
rect 270 -2670 275 -2640
rect 275 -2670 305 -2640
rect 305 -2670 310 -2640
rect 270 -2675 310 -2670
rect 270 -2710 310 -2705
rect 270 -2740 275 -2710
rect 275 -2740 305 -2710
rect 305 -2740 310 -2710
rect 270 -2745 310 -2740
rect 270 -2780 310 -2775
rect 270 -2810 275 -2780
rect 275 -2810 305 -2780
rect 305 -2810 310 -2780
rect 270 -2815 310 -2810
rect 270 -2845 310 -2840
rect 270 -2875 275 -2845
rect 275 -2875 305 -2845
rect 305 -2875 310 -2845
rect 270 -2880 310 -2875
rect 270 -2905 310 -2900
rect 270 -2935 275 -2905
rect 275 -2935 305 -2905
rect 305 -2935 310 -2905
rect 270 -2940 310 -2935
rect 270 -2970 310 -2965
rect 270 -3000 275 -2970
rect 275 -3000 305 -2970
rect 305 -3000 310 -2970
rect 270 -3005 310 -3000
rect 270 -3040 310 -3035
rect 270 -3070 275 -3040
rect 275 -3070 305 -3040
rect 305 -3070 310 -3040
rect 270 -3075 310 -3070
rect 270 -3110 310 -3105
rect 270 -3140 275 -3110
rect 275 -3140 305 -3110
rect 305 -3140 310 -3110
rect 270 -3145 310 -3140
rect 270 -3180 310 -3175
rect 270 -3210 275 -3180
rect 275 -3210 305 -3180
rect 305 -3210 310 -3180
rect 270 -3215 310 -3210
rect 270 -3245 310 -3240
rect 270 -3275 275 -3245
rect 275 -3275 305 -3245
rect 305 -3275 310 -3245
rect 270 -3280 310 -3275
rect 270 -3305 310 -3300
rect 270 -3335 275 -3305
rect 275 -3335 305 -3305
rect 305 -3335 310 -3305
rect 270 -3340 310 -3335
rect 270 -3370 310 -3365
rect 270 -3400 275 -3370
rect 275 -3400 305 -3370
rect 305 -3400 310 -3370
rect 270 -3405 310 -3400
rect 270 -3440 310 -3435
rect 270 -3470 275 -3440
rect 275 -3470 305 -3440
rect 305 -3470 310 -3440
rect 270 -3475 310 -3470
rect 270 -3510 310 -3505
rect 270 -3540 275 -3510
rect 275 -3540 305 -3510
rect 305 -3540 310 -3510
rect 270 -3545 310 -3540
rect 270 -3580 310 -3575
rect 270 -3610 275 -3580
rect 275 -3610 305 -3580
rect 305 -3610 310 -3580
rect 270 -3615 310 -3610
rect 270 -3645 310 -3640
rect 270 -3675 275 -3645
rect 275 -3675 305 -3645
rect 305 -3675 310 -3645
rect 270 -3680 310 -3675
rect 270 -3705 310 -3700
rect 270 -3735 275 -3705
rect 275 -3735 305 -3705
rect 305 -3735 310 -3705
rect 270 -3740 310 -3735
rect 270 -3770 310 -3765
rect 270 -3800 275 -3770
rect 275 -3800 305 -3770
rect 305 -3800 310 -3770
rect 270 -3805 310 -3800
rect 270 -3840 310 -3835
rect 270 -3870 275 -3840
rect 275 -3870 305 -3840
rect 305 -3870 310 -3840
rect 270 -3875 310 -3870
rect 270 -3910 310 -3905
rect 270 -3940 275 -3910
rect 275 -3940 305 -3910
rect 305 -3940 310 -3910
rect 270 -3945 310 -3940
rect 270 -3980 310 -3975
rect 270 -4010 275 -3980
rect 275 -4010 305 -3980
rect 305 -4010 310 -3980
rect 270 -4015 310 -4010
rect 270 -4045 310 -4040
rect 270 -4075 275 -4045
rect 275 -4075 305 -4045
rect 305 -4075 310 -4045
rect 270 -4080 310 -4075
rect 270 -4105 310 -4100
rect 270 -4135 275 -4105
rect 275 -4135 305 -4105
rect 305 -4135 310 -4105
rect 270 -4140 310 -4135
rect 270 -4170 310 -4165
rect 270 -4200 275 -4170
rect 275 -4200 305 -4170
rect 305 -4200 310 -4170
rect 270 -4205 310 -4200
rect 270 -4240 310 -4235
rect 270 -4270 275 -4240
rect 275 -4270 305 -4240
rect 305 -4270 310 -4240
rect 270 -4275 310 -4270
rect 270 -4310 310 -4305
rect 270 -4340 275 -4310
rect 275 -4340 305 -4310
rect 305 -4340 310 -4310
rect 270 -4345 310 -4340
rect 270 -4380 310 -4375
rect 270 -4410 275 -4380
rect 275 -4410 305 -4380
rect 305 -4410 310 -4380
rect 270 -4415 310 -4410
rect 270 -4445 310 -4440
rect 270 -4475 275 -4445
rect 275 -4475 305 -4445
rect 305 -4475 310 -4445
rect 270 -4480 310 -4475
rect 620 -1305 660 -1300
rect 620 -1335 625 -1305
rect 625 -1335 655 -1305
rect 655 -1335 660 -1305
rect 620 -1340 660 -1335
rect 620 -1370 660 -1365
rect 620 -1400 625 -1370
rect 625 -1400 655 -1370
rect 655 -1400 660 -1370
rect 620 -1405 660 -1400
rect 620 -1440 660 -1435
rect 620 -1470 625 -1440
rect 625 -1470 655 -1440
rect 655 -1470 660 -1440
rect 620 -1475 660 -1470
rect 620 -1510 660 -1505
rect 620 -1540 625 -1510
rect 625 -1540 655 -1510
rect 655 -1540 660 -1510
rect 620 -1545 660 -1540
rect 620 -1580 660 -1575
rect 620 -1610 625 -1580
rect 625 -1610 655 -1580
rect 655 -1610 660 -1580
rect 620 -1615 660 -1610
rect 620 -1645 660 -1640
rect 620 -1675 625 -1645
rect 625 -1675 655 -1645
rect 655 -1675 660 -1645
rect 620 -1680 660 -1675
rect 620 -1705 660 -1700
rect 620 -1735 625 -1705
rect 625 -1735 655 -1705
rect 655 -1735 660 -1705
rect 620 -1740 660 -1735
rect 620 -1770 660 -1765
rect 620 -1800 625 -1770
rect 625 -1800 655 -1770
rect 655 -1800 660 -1770
rect 620 -1805 660 -1800
rect 620 -1840 660 -1835
rect 620 -1870 625 -1840
rect 625 -1870 655 -1840
rect 655 -1870 660 -1840
rect 620 -1875 660 -1870
rect 620 -1910 660 -1905
rect 620 -1940 625 -1910
rect 625 -1940 655 -1910
rect 655 -1940 660 -1910
rect 620 -1945 660 -1940
rect 620 -1980 660 -1975
rect 620 -2010 625 -1980
rect 625 -2010 655 -1980
rect 655 -2010 660 -1980
rect 620 -2015 660 -2010
rect 620 -2045 660 -2040
rect 620 -2075 625 -2045
rect 625 -2075 655 -2045
rect 655 -2075 660 -2045
rect 620 -2080 660 -2075
rect 620 -2105 660 -2100
rect 620 -2135 625 -2105
rect 625 -2135 655 -2105
rect 655 -2135 660 -2105
rect 620 -2140 660 -2135
rect 620 -2170 660 -2165
rect 620 -2200 625 -2170
rect 625 -2200 655 -2170
rect 655 -2200 660 -2170
rect 620 -2205 660 -2200
rect 620 -2240 660 -2235
rect 620 -2270 625 -2240
rect 625 -2270 655 -2240
rect 655 -2270 660 -2240
rect 620 -2275 660 -2270
rect 620 -2310 660 -2305
rect 620 -2340 625 -2310
rect 625 -2340 655 -2310
rect 655 -2340 660 -2310
rect 620 -2345 660 -2340
rect 620 -2380 660 -2375
rect 620 -2410 625 -2380
rect 625 -2410 655 -2380
rect 655 -2410 660 -2380
rect 620 -2415 660 -2410
rect 620 -2445 660 -2440
rect 620 -2475 625 -2445
rect 625 -2475 655 -2445
rect 655 -2475 660 -2445
rect 620 -2480 660 -2475
rect 620 -2505 660 -2500
rect 620 -2535 625 -2505
rect 625 -2535 655 -2505
rect 655 -2535 660 -2505
rect 620 -2540 660 -2535
rect 620 -2570 660 -2565
rect 620 -2600 625 -2570
rect 625 -2600 655 -2570
rect 655 -2600 660 -2570
rect 620 -2605 660 -2600
rect 620 -2640 660 -2635
rect 620 -2670 625 -2640
rect 625 -2670 655 -2640
rect 655 -2670 660 -2640
rect 620 -2675 660 -2670
rect 620 -2710 660 -2705
rect 620 -2740 625 -2710
rect 625 -2740 655 -2710
rect 655 -2740 660 -2710
rect 620 -2745 660 -2740
rect 620 -2780 660 -2775
rect 620 -2810 625 -2780
rect 625 -2810 655 -2780
rect 655 -2810 660 -2780
rect 620 -2815 660 -2810
rect 620 -2845 660 -2840
rect 620 -2875 625 -2845
rect 625 -2875 655 -2845
rect 655 -2875 660 -2845
rect 620 -2880 660 -2875
rect 620 -2905 660 -2900
rect 620 -2935 625 -2905
rect 625 -2935 655 -2905
rect 655 -2935 660 -2905
rect 620 -2940 660 -2935
rect 620 -2970 660 -2965
rect 620 -3000 625 -2970
rect 625 -3000 655 -2970
rect 655 -3000 660 -2970
rect 620 -3005 660 -3000
rect 620 -3040 660 -3035
rect 620 -3070 625 -3040
rect 625 -3070 655 -3040
rect 655 -3070 660 -3040
rect 620 -3075 660 -3070
rect 620 -3110 660 -3105
rect 620 -3140 625 -3110
rect 625 -3140 655 -3110
rect 655 -3140 660 -3110
rect 620 -3145 660 -3140
rect 620 -3180 660 -3175
rect 620 -3210 625 -3180
rect 625 -3210 655 -3180
rect 655 -3210 660 -3180
rect 620 -3215 660 -3210
rect 620 -3245 660 -3240
rect 620 -3275 625 -3245
rect 625 -3275 655 -3245
rect 655 -3275 660 -3245
rect 620 -3280 660 -3275
rect 620 -3305 660 -3300
rect 620 -3335 625 -3305
rect 625 -3335 655 -3305
rect 655 -3335 660 -3305
rect 620 -3340 660 -3335
rect 620 -3370 660 -3365
rect 620 -3400 625 -3370
rect 625 -3400 655 -3370
rect 655 -3400 660 -3370
rect 620 -3405 660 -3400
rect 620 -3440 660 -3435
rect 620 -3470 625 -3440
rect 625 -3470 655 -3440
rect 655 -3470 660 -3440
rect 620 -3475 660 -3470
rect 620 -3510 660 -3505
rect 620 -3540 625 -3510
rect 625 -3540 655 -3510
rect 655 -3540 660 -3510
rect 620 -3545 660 -3540
rect 620 -3580 660 -3575
rect 620 -3610 625 -3580
rect 625 -3610 655 -3580
rect 655 -3610 660 -3580
rect 620 -3615 660 -3610
rect 620 -3645 660 -3640
rect 620 -3675 625 -3645
rect 625 -3675 655 -3645
rect 655 -3675 660 -3645
rect 620 -3680 660 -3675
rect 620 -3705 660 -3700
rect 620 -3735 625 -3705
rect 625 -3735 655 -3705
rect 655 -3735 660 -3705
rect 620 -3740 660 -3735
rect 620 -3770 660 -3765
rect 620 -3800 625 -3770
rect 625 -3800 655 -3770
rect 655 -3800 660 -3770
rect 620 -3805 660 -3800
rect 620 -3840 660 -3835
rect 620 -3870 625 -3840
rect 625 -3870 655 -3840
rect 655 -3870 660 -3840
rect 620 -3875 660 -3870
rect 620 -3910 660 -3905
rect 620 -3940 625 -3910
rect 625 -3940 655 -3910
rect 655 -3940 660 -3910
rect 620 -3945 660 -3940
rect 620 -3980 660 -3975
rect 620 -4010 625 -3980
rect 625 -4010 655 -3980
rect 655 -4010 660 -3980
rect 620 -4015 660 -4010
rect 620 -4045 660 -4040
rect 620 -4075 625 -4045
rect 625 -4075 655 -4045
rect 655 -4075 660 -4045
rect 620 -4080 660 -4075
rect 620 -4105 660 -4100
rect 620 -4135 625 -4105
rect 625 -4135 655 -4105
rect 655 -4135 660 -4105
rect 620 -4140 660 -4135
rect 620 -4170 660 -4165
rect 620 -4200 625 -4170
rect 625 -4200 655 -4170
rect 655 -4200 660 -4170
rect 620 -4205 660 -4200
rect 620 -4240 660 -4235
rect 620 -4270 625 -4240
rect 625 -4270 655 -4240
rect 655 -4270 660 -4240
rect 620 -4275 660 -4270
rect 620 -4310 660 -4305
rect 620 -4340 625 -4310
rect 625 -4340 655 -4310
rect 655 -4340 660 -4310
rect 620 -4345 660 -4340
rect 620 -4380 660 -4375
rect 620 -4410 625 -4380
rect 625 -4410 655 -4380
rect 655 -4410 660 -4380
rect 620 -4415 660 -4410
rect 620 -4445 660 -4440
rect 620 -4475 625 -4445
rect 625 -4475 655 -4445
rect 655 -4475 660 -4445
rect 620 -4480 660 -4475
rect 970 -1305 1010 -1300
rect 970 -1335 975 -1305
rect 975 -1335 1005 -1305
rect 1005 -1335 1010 -1305
rect 970 -1340 1010 -1335
rect 970 -1370 1010 -1365
rect 970 -1400 975 -1370
rect 975 -1400 1005 -1370
rect 1005 -1400 1010 -1370
rect 970 -1405 1010 -1400
rect 970 -1440 1010 -1435
rect 970 -1470 975 -1440
rect 975 -1470 1005 -1440
rect 1005 -1470 1010 -1440
rect 970 -1475 1010 -1470
rect 970 -1510 1010 -1505
rect 970 -1540 975 -1510
rect 975 -1540 1005 -1510
rect 1005 -1540 1010 -1510
rect 970 -1545 1010 -1540
rect 970 -1580 1010 -1575
rect 970 -1610 975 -1580
rect 975 -1610 1005 -1580
rect 1005 -1610 1010 -1580
rect 970 -1615 1010 -1610
rect 970 -1645 1010 -1640
rect 970 -1675 975 -1645
rect 975 -1675 1005 -1645
rect 1005 -1675 1010 -1645
rect 970 -1680 1010 -1675
rect 970 -1705 1010 -1700
rect 970 -1735 975 -1705
rect 975 -1735 1005 -1705
rect 1005 -1735 1010 -1705
rect 970 -1740 1010 -1735
rect 970 -1770 1010 -1765
rect 970 -1800 975 -1770
rect 975 -1800 1005 -1770
rect 1005 -1800 1010 -1770
rect 970 -1805 1010 -1800
rect 970 -1840 1010 -1835
rect 970 -1870 975 -1840
rect 975 -1870 1005 -1840
rect 1005 -1870 1010 -1840
rect 970 -1875 1010 -1870
rect 970 -1910 1010 -1905
rect 970 -1940 975 -1910
rect 975 -1940 1005 -1910
rect 1005 -1940 1010 -1910
rect 970 -1945 1010 -1940
rect 970 -1980 1010 -1975
rect 970 -2010 975 -1980
rect 975 -2010 1005 -1980
rect 1005 -2010 1010 -1980
rect 970 -2015 1010 -2010
rect 970 -2045 1010 -2040
rect 970 -2075 975 -2045
rect 975 -2075 1005 -2045
rect 1005 -2075 1010 -2045
rect 970 -2080 1010 -2075
rect 970 -2105 1010 -2100
rect 970 -2135 975 -2105
rect 975 -2135 1005 -2105
rect 1005 -2135 1010 -2105
rect 970 -2140 1010 -2135
rect 970 -2170 1010 -2165
rect 970 -2200 975 -2170
rect 975 -2200 1005 -2170
rect 1005 -2200 1010 -2170
rect 970 -2205 1010 -2200
rect 970 -2240 1010 -2235
rect 970 -2270 975 -2240
rect 975 -2270 1005 -2240
rect 1005 -2270 1010 -2240
rect 970 -2275 1010 -2270
rect 970 -2310 1010 -2305
rect 970 -2340 975 -2310
rect 975 -2340 1005 -2310
rect 1005 -2340 1010 -2310
rect 970 -2345 1010 -2340
rect 970 -2380 1010 -2375
rect 970 -2410 975 -2380
rect 975 -2410 1005 -2380
rect 1005 -2410 1010 -2380
rect 970 -2415 1010 -2410
rect 970 -2445 1010 -2440
rect 970 -2475 975 -2445
rect 975 -2475 1005 -2445
rect 1005 -2475 1010 -2445
rect 970 -2480 1010 -2475
rect 970 -2505 1010 -2500
rect 970 -2535 975 -2505
rect 975 -2535 1005 -2505
rect 1005 -2535 1010 -2505
rect 970 -2540 1010 -2535
rect 970 -2570 1010 -2565
rect 970 -2600 975 -2570
rect 975 -2600 1005 -2570
rect 1005 -2600 1010 -2570
rect 970 -2605 1010 -2600
rect 970 -2640 1010 -2635
rect 970 -2670 975 -2640
rect 975 -2670 1005 -2640
rect 1005 -2670 1010 -2640
rect 970 -2675 1010 -2670
rect 970 -2710 1010 -2705
rect 970 -2740 975 -2710
rect 975 -2740 1005 -2710
rect 1005 -2740 1010 -2710
rect 970 -2745 1010 -2740
rect 970 -2780 1010 -2775
rect 970 -2810 975 -2780
rect 975 -2810 1005 -2780
rect 1005 -2810 1010 -2780
rect 970 -2815 1010 -2810
rect 970 -2845 1010 -2840
rect 970 -2875 975 -2845
rect 975 -2875 1005 -2845
rect 1005 -2875 1010 -2845
rect 970 -2880 1010 -2875
rect 970 -2905 1010 -2900
rect 970 -2935 975 -2905
rect 975 -2935 1005 -2905
rect 1005 -2935 1010 -2905
rect 970 -2940 1010 -2935
rect 970 -2970 1010 -2965
rect 970 -3000 975 -2970
rect 975 -3000 1005 -2970
rect 1005 -3000 1010 -2970
rect 970 -3005 1010 -3000
rect 970 -3040 1010 -3035
rect 970 -3070 975 -3040
rect 975 -3070 1005 -3040
rect 1005 -3070 1010 -3040
rect 970 -3075 1010 -3070
rect 970 -3110 1010 -3105
rect 970 -3140 975 -3110
rect 975 -3140 1005 -3110
rect 1005 -3140 1010 -3110
rect 970 -3145 1010 -3140
rect 970 -3180 1010 -3175
rect 970 -3210 975 -3180
rect 975 -3210 1005 -3180
rect 1005 -3210 1010 -3180
rect 970 -3215 1010 -3210
rect 970 -3245 1010 -3240
rect 970 -3275 975 -3245
rect 975 -3275 1005 -3245
rect 1005 -3275 1010 -3245
rect 970 -3280 1010 -3275
rect 970 -3305 1010 -3300
rect 970 -3335 975 -3305
rect 975 -3335 1005 -3305
rect 1005 -3335 1010 -3305
rect 970 -3340 1010 -3335
rect 970 -3370 1010 -3365
rect 970 -3400 975 -3370
rect 975 -3400 1005 -3370
rect 1005 -3400 1010 -3370
rect 970 -3405 1010 -3400
rect 970 -3440 1010 -3435
rect 970 -3470 975 -3440
rect 975 -3470 1005 -3440
rect 1005 -3470 1010 -3440
rect 970 -3475 1010 -3470
rect 970 -3510 1010 -3505
rect 970 -3540 975 -3510
rect 975 -3540 1005 -3510
rect 1005 -3540 1010 -3510
rect 970 -3545 1010 -3540
rect 970 -3580 1010 -3575
rect 970 -3610 975 -3580
rect 975 -3610 1005 -3580
rect 1005 -3610 1010 -3580
rect 970 -3615 1010 -3610
rect 970 -3645 1010 -3640
rect 970 -3675 975 -3645
rect 975 -3675 1005 -3645
rect 1005 -3675 1010 -3645
rect 970 -3680 1010 -3675
rect 970 -3705 1010 -3700
rect 970 -3735 975 -3705
rect 975 -3735 1005 -3705
rect 1005 -3735 1010 -3705
rect 970 -3740 1010 -3735
rect 970 -3770 1010 -3765
rect 970 -3800 975 -3770
rect 975 -3800 1005 -3770
rect 1005 -3800 1010 -3770
rect 970 -3805 1010 -3800
rect 970 -3840 1010 -3835
rect 970 -3870 975 -3840
rect 975 -3870 1005 -3840
rect 1005 -3870 1010 -3840
rect 970 -3875 1010 -3870
rect 970 -3910 1010 -3905
rect 970 -3940 975 -3910
rect 975 -3940 1005 -3910
rect 1005 -3940 1010 -3910
rect 970 -3945 1010 -3940
rect 970 -3980 1010 -3975
rect 970 -4010 975 -3980
rect 975 -4010 1005 -3980
rect 1005 -4010 1010 -3980
rect 970 -4015 1010 -4010
rect 970 -4045 1010 -4040
rect 970 -4075 975 -4045
rect 975 -4075 1005 -4045
rect 1005 -4075 1010 -4045
rect 970 -4080 1010 -4075
rect 970 -4105 1010 -4100
rect 970 -4135 975 -4105
rect 975 -4135 1005 -4105
rect 1005 -4135 1010 -4105
rect 970 -4140 1010 -4135
rect 970 -4170 1010 -4165
rect 970 -4200 975 -4170
rect 975 -4200 1005 -4170
rect 1005 -4200 1010 -4170
rect 970 -4205 1010 -4200
rect 970 -4240 1010 -4235
rect 970 -4270 975 -4240
rect 975 -4270 1005 -4240
rect 1005 -4270 1010 -4240
rect 970 -4275 1010 -4270
rect 970 -4310 1010 -4305
rect 970 -4340 975 -4310
rect 975 -4340 1005 -4310
rect 1005 -4340 1010 -4310
rect 970 -4345 1010 -4340
rect 970 -4380 1010 -4375
rect 970 -4410 975 -4380
rect 975 -4410 1005 -4380
rect 1005 -4410 1010 -4380
rect 970 -4415 1010 -4410
rect 970 -4445 1010 -4440
rect 970 -4475 975 -4445
rect 975 -4475 1005 -4445
rect 1005 -4475 1010 -4445
rect 970 -4480 1010 -4475
rect 1320 -1305 1360 -1300
rect 1320 -1335 1325 -1305
rect 1325 -1335 1355 -1305
rect 1355 -1335 1360 -1305
rect 1320 -1340 1360 -1335
rect 1320 -1370 1360 -1365
rect 1320 -1400 1325 -1370
rect 1325 -1400 1355 -1370
rect 1355 -1400 1360 -1370
rect 1320 -1405 1360 -1400
rect 1320 -1440 1360 -1435
rect 1320 -1470 1325 -1440
rect 1325 -1470 1355 -1440
rect 1355 -1470 1360 -1440
rect 1320 -1475 1360 -1470
rect 1320 -1510 1360 -1505
rect 1320 -1540 1325 -1510
rect 1325 -1540 1355 -1510
rect 1355 -1540 1360 -1510
rect 1320 -1545 1360 -1540
rect 1320 -1580 1360 -1575
rect 1320 -1610 1325 -1580
rect 1325 -1610 1355 -1580
rect 1355 -1610 1360 -1580
rect 1320 -1615 1360 -1610
rect 1320 -1645 1360 -1640
rect 1320 -1675 1325 -1645
rect 1325 -1675 1355 -1645
rect 1355 -1675 1360 -1645
rect 1320 -1680 1360 -1675
rect 1320 -1705 1360 -1700
rect 1320 -1735 1325 -1705
rect 1325 -1735 1355 -1705
rect 1355 -1735 1360 -1705
rect 1320 -1740 1360 -1735
rect 1320 -1770 1360 -1765
rect 1320 -1800 1325 -1770
rect 1325 -1800 1355 -1770
rect 1355 -1800 1360 -1770
rect 1320 -1805 1360 -1800
rect 1320 -1840 1360 -1835
rect 1320 -1870 1325 -1840
rect 1325 -1870 1355 -1840
rect 1355 -1870 1360 -1840
rect 1320 -1875 1360 -1870
rect 1320 -1910 1360 -1905
rect 1320 -1940 1325 -1910
rect 1325 -1940 1355 -1910
rect 1355 -1940 1360 -1910
rect 1320 -1945 1360 -1940
rect 1320 -1980 1360 -1975
rect 1320 -2010 1325 -1980
rect 1325 -2010 1355 -1980
rect 1355 -2010 1360 -1980
rect 1320 -2015 1360 -2010
rect 1320 -2045 1360 -2040
rect 1320 -2075 1325 -2045
rect 1325 -2075 1355 -2045
rect 1355 -2075 1360 -2045
rect 1320 -2080 1360 -2075
rect 1320 -2105 1360 -2100
rect 1320 -2135 1325 -2105
rect 1325 -2135 1355 -2105
rect 1355 -2135 1360 -2105
rect 1320 -2140 1360 -2135
rect 1320 -2170 1360 -2165
rect 1320 -2200 1325 -2170
rect 1325 -2200 1355 -2170
rect 1355 -2200 1360 -2170
rect 1320 -2205 1360 -2200
rect 1320 -2240 1360 -2235
rect 1320 -2270 1325 -2240
rect 1325 -2270 1355 -2240
rect 1355 -2270 1360 -2240
rect 1320 -2275 1360 -2270
rect 1320 -2310 1360 -2305
rect 1320 -2340 1325 -2310
rect 1325 -2340 1355 -2310
rect 1355 -2340 1360 -2310
rect 1320 -2345 1360 -2340
rect 1320 -2380 1360 -2375
rect 1320 -2410 1325 -2380
rect 1325 -2410 1355 -2380
rect 1355 -2410 1360 -2380
rect 1320 -2415 1360 -2410
rect 1320 -2445 1360 -2440
rect 1320 -2475 1325 -2445
rect 1325 -2475 1355 -2445
rect 1355 -2475 1360 -2445
rect 1320 -2480 1360 -2475
rect 1320 -2505 1360 -2500
rect 1320 -2535 1325 -2505
rect 1325 -2535 1355 -2505
rect 1355 -2535 1360 -2505
rect 1320 -2540 1360 -2535
rect 1320 -2570 1360 -2565
rect 1320 -2600 1325 -2570
rect 1325 -2600 1355 -2570
rect 1355 -2600 1360 -2570
rect 1320 -2605 1360 -2600
rect 1320 -2640 1360 -2635
rect 1320 -2670 1325 -2640
rect 1325 -2670 1355 -2640
rect 1355 -2670 1360 -2640
rect 1320 -2675 1360 -2670
rect 1320 -2710 1360 -2705
rect 1320 -2740 1325 -2710
rect 1325 -2740 1355 -2710
rect 1355 -2740 1360 -2710
rect 1320 -2745 1360 -2740
rect 1320 -2780 1360 -2775
rect 1320 -2810 1325 -2780
rect 1325 -2810 1355 -2780
rect 1355 -2810 1360 -2780
rect 1320 -2815 1360 -2810
rect 1320 -2845 1360 -2840
rect 1320 -2875 1325 -2845
rect 1325 -2875 1355 -2845
rect 1355 -2875 1360 -2845
rect 1320 -2880 1360 -2875
rect 1320 -2905 1360 -2900
rect 1320 -2935 1325 -2905
rect 1325 -2935 1355 -2905
rect 1355 -2935 1360 -2905
rect 1320 -2940 1360 -2935
rect 1320 -2970 1360 -2965
rect 1320 -3000 1325 -2970
rect 1325 -3000 1355 -2970
rect 1355 -3000 1360 -2970
rect 1320 -3005 1360 -3000
rect 1320 -3040 1360 -3035
rect 1320 -3070 1325 -3040
rect 1325 -3070 1355 -3040
rect 1355 -3070 1360 -3040
rect 1320 -3075 1360 -3070
rect 1320 -3110 1360 -3105
rect 1320 -3140 1325 -3110
rect 1325 -3140 1355 -3110
rect 1355 -3140 1360 -3110
rect 1320 -3145 1360 -3140
rect 1320 -3180 1360 -3175
rect 1320 -3210 1325 -3180
rect 1325 -3210 1355 -3180
rect 1355 -3210 1360 -3180
rect 1320 -3215 1360 -3210
rect 1320 -3245 1360 -3240
rect 1320 -3275 1325 -3245
rect 1325 -3275 1355 -3245
rect 1355 -3275 1360 -3245
rect 1320 -3280 1360 -3275
rect 1320 -3305 1360 -3300
rect 1320 -3335 1325 -3305
rect 1325 -3335 1355 -3305
rect 1355 -3335 1360 -3305
rect 1320 -3340 1360 -3335
rect 1320 -3370 1360 -3365
rect 1320 -3400 1325 -3370
rect 1325 -3400 1355 -3370
rect 1355 -3400 1360 -3370
rect 1320 -3405 1360 -3400
rect 1320 -3440 1360 -3435
rect 1320 -3470 1325 -3440
rect 1325 -3470 1355 -3440
rect 1355 -3470 1360 -3440
rect 1320 -3475 1360 -3470
rect 1320 -3510 1360 -3505
rect 1320 -3540 1325 -3510
rect 1325 -3540 1355 -3510
rect 1355 -3540 1360 -3510
rect 1320 -3545 1360 -3540
rect 1320 -3580 1360 -3575
rect 1320 -3610 1325 -3580
rect 1325 -3610 1355 -3580
rect 1355 -3610 1360 -3580
rect 1320 -3615 1360 -3610
rect 1320 -3645 1360 -3640
rect 1320 -3675 1325 -3645
rect 1325 -3675 1355 -3645
rect 1355 -3675 1360 -3645
rect 1320 -3680 1360 -3675
rect 1320 -3705 1360 -3700
rect 1320 -3735 1325 -3705
rect 1325 -3735 1355 -3705
rect 1355 -3735 1360 -3705
rect 1320 -3740 1360 -3735
rect 1320 -3770 1360 -3765
rect 1320 -3800 1325 -3770
rect 1325 -3800 1355 -3770
rect 1355 -3800 1360 -3770
rect 1320 -3805 1360 -3800
rect 1320 -3840 1360 -3835
rect 1320 -3870 1325 -3840
rect 1325 -3870 1355 -3840
rect 1355 -3870 1360 -3840
rect 1320 -3875 1360 -3870
rect 1320 -3910 1360 -3905
rect 1320 -3940 1325 -3910
rect 1325 -3940 1355 -3910
rect 1355 -3940 1360 -3910
rect 1320 -3945 1360 -3940
rect 1320 -3980 1360 -3975
rect 1320 -4010 1325 -3980
rect 1325 -4010 1355 -3980
rect 1355 -4010 1360 -3980
rect 1320 -4015 1360 -4010
rect 1320 -4045 1360 -4040
rect 1320 -4075 1325 -4045
rect 1325 -4075 1355 -4045
rect 1355 -4075 1360 -4045
rect 1320 -4080 1360 -4075
rect 1320 -4105 1360 -4100
rect 1320 -4135 1325 -4105
rect 1325 -4135 1355 -4105
rect 1355 -4135 1360 -4105
rect 1320 -4140 1360 -4135
rect 1320 -4170 1360 -4165
rect 1320 -4200 1325 -4170
rect 1325 -4200 1355 -4170
rect 1355 -4200 1360 -4170
rect 1320 -4205 1360 -4200
rect 1320 -4240 1360 -4235
rect 1320 -4270 1325 -4240
rect 1325 -4270 1355 -4240
rect 1355 -4270 1360 -4240
rect 1320 -4275 1360 -4270
rect 1320 -4310 1360 -4305
rect 1320 -4340 1325 -4310
rect 1325 -4340 1355 -4310
rect 1355 -4340 1360 -4310
rect 1320 -4345 1360 -4340
rect 1320 -4380 1360 -4375
rect 1320 -4410 1325 -4380
rect 1325 -4410 1355 -4380
rect 1355 -4410 1360 -4380
rect 1320 -4415 1360 -4410
rect 1320 -4445 1360 -4440
rect 1320 -4475 1325 -4445
rect 1325 -4475 1355 -4445
rect 1355 -4475 1360 -4445
rect 1320 -4480 1360 -4475
rect 1670 -1305 1710 -1300
rect 1670 -1335 1675 -1305
rect 1675 -1335 1705 -1305
rect 1705 -1335 1710 -1305
rect 1670 -1340 1710 -1335
rect 1670 -1370 1710 -1365
rect 1670 -1400 1675 -1370
rect 1675 -1400 1705 -1370
rect 1705 -1400 1710 -1370
rect 1670 -1405 1710 -1400
rect 1670 -1440 1710 -1435
rect 1670 -1470 1675 -1440
rect 1675 -1470 1705 -1440
rect 1705 -1470 1710 -1440
rect 1670 -1475 1710 -1470
rect 1670 -1510 1710 -1505
rect 1670 -1540 1675 -1510
rect 1675 -1540 1705 -1510
rect 1705 -1540 1710 -1510
rect 1670 -1545 1710 -1540
rect 1670 -1580 1710 -1575
rect 1670 -1610 1675 -1580
rect 1675 -1610 1705 -1580
rect 1705 -1610 1710 -1580
rect 1670 -1615 1710 -1610
rect 1670 -1645 1710 -1640
rect 1670 -1675 1675 -1645
rect 1675 -1675 1705 -1645
rect 1705 -1675 1710 -1645
rect 1670 -1680 1710 -1675
rect 1670 -1705 1710 -1700
rect 1670 -1735 1675 -1705
rect 1675 -1735 1705 -1705
rect 1705 -1735 1710 -1705
rect 1670 -1740 1710 -1735
rect 1670 -1770 1710 -1765
rect 1670 -1800 1675 -1770
rect 1675 -1800 1705 -1770
rect 1705 -1800 1710 -1770
rect 1670 -1805 1710 -1800
rect 1670 -1840 1710 -1835
rect 1670 -1870 1675 -1840
rect 1675 -1870 1705 -1840
rect 1705 -1870 1710 -1840
rect 1670 -1875 1710 -1870
rect 1670 -1910 1710 -1905
rect 1670 -1940 1675 -1910
rect 1675 -1940 1705 -1910
rect 1705 -1940 1710 -1910
rect 1670 -1945 1710 -1940
rect 1670 -1980 1710 -1975
rect 1670 -2010 1675 -1980
rect 1675 -2010 1705 -1980
rect 1705 -2010 1710 -1980
rect 1670 -2015 1710 -2010
rect 1670 -2045 1710 -2040
rect 1670 -2075 1675 -2045
rect 1675 -2075 1705 -2045
rect 1705 -2075 1710 -2045
rect 1670 -2080 1710 -2075
rect 1670 -2105 1710 -2100
rect 1670 -2135 1675 -2105
rect 1675 -2135 1705 -2105
rect 1705 -2135 1710 -2105
rect 1670 -2140 1710 -2135
rect 1670 -2170 1710 -2165
rect 1670 -2200 1675 -2170
rect 1675 -2200 1705 -2170
rect 1705 -2200 1710 -2170
rect 1670 -2205 1710 -2200
rect 1670 -2240 1710 -2235
rect 1670 -2270 1675 -2240
rect 1675 -2270 1705 -2240
rect 1705 -2270 1710 -2240
rect 1670 -2275 1710 -2270
rect 1670 -2310 1710 -2305
rect 1670 -2340 1675 -2310
rect 1675 -2340 1705 -2310
rect 1705 -2340 1710 -2310
rect 1670 -2345 1710 -2340
rect 1670 -2380 1710 -2375
rect 1670 -2410 1675 -2380
rect 1675 -2410 1705 -2380
rect 1705 -2410 1710 -2380
rect 1670 -2415 1710 -2410
rect 1670 -2445 1710 -2440
rect 1670 -2475 1675 -2445
rect 1675 -2475 1705 -2445
rect 1705 -2475 1710 -2445
rect 1670 -2480 1710 -2475
rect 1670 -2505 1710 -2500
rect 1670 -2535 1675 -2505
rect 1675 -2535 1705 -2505
rect 1705 -2535 1710 -2505
rect 1670 -2540 1710 -2535
rect 1670 -2570 1710 -2565
rect 1670 -2600 1675 -2570
rect 1675 -2600 1705 -2570
rect 1705 -2600 1710 -2570
rect 1670 -2605 1710 -2600
rect 1670 -2640 1710 -2635
rect 1670 -2670 1675 -2640
rect 1675 -2670 1705 -2640
rect 1705 -2670 1710 -2640
rect 1670 -2675 1710 -2670
rect 1670 -2710 1710 -2705
rect 1670 -2740 1675 -2710
rect 1675 -2740 1705 -2710
rect 1705 -2740 1710 -2710
rect 1670 -2745 1710 -2740
rect 1670 -2780 1710 -2775
rect 1670 -2810 1675 -2780
rect 1675 -2810 1705 -2780
rect 1705 -2810 1710 -2780
rect 1670 -2815 1710 -2810
rect 1670 -2845 1710 -2840
rect 1670 -2875 1675 -2845
rect 1675 -2875 1705 -2845
rect 1705 -2875 1710 -2845
rect 1670 -2880 1710 -2875
rect 1670 -2905 1710 -2900
rect 1670 -2935 1675 -2905
rect 1675 -2935 1705 -2905
rect 1705 -2935 1710 -2905
rect 1670 -2940 1710 -2935
rect 1670 -2970 1710 -2965
rect 1670 -3000 1675 -2970
rect 1675 -3000 1705 -2970
rect 1705 -3000 1710 -2970
rect 1670 -3005 1710 -3000
rect 1670 -3040 1710 -3035
rect 1670 -3070 1675 -3040
rect 1675 -3070 1705 -3040
rect 1705 -3070 1710 -3040
rect 1670 -3075 1710 -3070
rect 1670 -3110 1710 -3105
rect 1670 -3140 1675 -3110
rect 1675 -3140 1705 -3110
rect 1705 -3140 1710 -3110
rect 1670 -3145 1710 -3140
rect 1670 -3180 1710 -3175
rect 1670 -3210 1675 -3180
rect 1675 -3210 1705 -3180
rect 1705 -3210 1710 -3180
rect 1670 -3215 1710 -3210
rect 1670 -3245 1710 -3240
rect 1670 -3275 1675 -3245
rect 1675 -3275 1705 -3245
rect 1705 -3275 1710 -3245
rect 1670 -3280 1710 -3275
rect 1670 -3305 1710 -3300
rect 1670 -3335 1675 -3305
rect 1675 -3335 1705 -3305
rect 1705 -3335 1710 -3305
rect 1670 -3340 1710 -3335
rect 1670 -3370 1710 -3365
rect 1670 -3400 1675 -3370
rect 1675 -3400 1705 -3370
rect 1705 -3400 1710 -3370
rect 1670 -3405 1710 -3400
rect 1670 -3440 1710 -3435
rect 1670 -3470 1675 -3440
rect 1675 -3470 1705 -3440
rect 1705 -3470 1710 -3440
rect 1670 -3475 1710 -3470
rect 1670 -3510 1710 -3505
rect 1670 -3540 1675 -3510
rect 1675 -3540 1705 -3510
rect 1705 -3540 1710 -3510
rect 1670 -3545 1710 -3540
rect 1670 -3580 1710 -3575
rect 1670 -3610 1675 -3580
rect 1675 -3610 1705 -3580
rect 1705 -3610 1710 -3580
rect 1670 -3615 1710 -3610
rect 1670 -3645 1710 -3640
rect 1670 -3675 1675 -3645
rect 1675 -3675 1705 -3645
rect 1705 -3675 1710 -3645
rect 1670 -3680 1710 -3675
rect 1670 -3705 1710 -3700
rect 1670 -3735 1675 -3705
rect 1675 -3735 1705 -3705
rect 1705 -3735 1710 -3705
rect 1670 -3740 1710 -3735
rect 1670 -3770 1710 -3765
rect 1670 -3800 1675 -3770
rect 1675 -3800 1705 -3770
rect 1705 -3800 1710 -3770
rect 1670 -3805 1710 -3800
rect 1670 -3840 1710 -3835
rect 1670 -3870 1675 -3840
rect 1675 -3870 1705 -3840
rect 1705 -3870 1710 -3840
rect 1670 -3875 1710 -3870
rect 1670 -3910 1710 -3905
rect 1670 -3940 1675 -3910
rect 1675 -3940 1705 -3910
rect 1705 -3940 1710 -3910
rect 1670 -3945 1710 -3940
rect 1670 -3980 1710 -3975
rect 1670 -4010 1675 -3980
rect 1675 -4010 1705 -3980
rect 1705 -4010 1710 -3980
rect 1670 -4015 1710 -4010
rect 1670 -4045 1710 -4040
rect 1670 -4075 1675 -4045
rect 1675 -4075 1705 -4045
rect 1705 -4075 1710 -4045
rect 1670 -4080 1710 -4075
rect 1670 -4105 1710 -4100
rect 1670 -4135 1675 -4105
rect 1675 -4135 1705 -4105
rect 1705 -4135 1710 -4105
rect 1670 -4140 1710 -4135
rect 1670 -4170 1710 -4165
rect 1670 -4200 1675 -4170
rect 1675 -4200 1705 -4170
rect 1705 -4200 1710 -4170
rect 1670 -4205 1710 -4200
rect 1670 -4240 1710 -4235
rect 1670 -4270 1675 -4240
rect 1675 -4270 1705 -4240
rect 1705 -4270 1710 -4240
rect 1670 -4275 1710 -4270
rect 1670 -4310 1710 -4305
rect 1670 -4340 1675 -4310
rect 1675 -4340 1705 -4310
rect 1705 -4340 1710 -4310
rect 1670 -4345 1710 -4340
rect 1670 -4380 1710 -4375
rect 1670 -4410 1675 -4380
rect 1675 -4410 1705 -4380
rect 1705 -4410 1710 -4380
rect 1670 -4415 1710 -4410
rect 1670 -4445 1710 -4440
rect 1670 -4475 1675 -4445
rect 1675 -4475 1705 -4445
rect 1705 -4475 1710 -4445
rect 1670 -4480 1710 -4475
rect 2020 -1305 2060 -1300
rect 2020 -1335 2025 -1305
rect 2025 -1335 2055 -1305
rect 2055 -1335 2060 -1305
rect 2020 -1340 2060 -1335
rect 2020 -1370 2060 -1365
rect 2020 -1400 2025 -1370
rect 2025 -1400 2055 -1370
rect 2055 -1400 2060 -1370
rect 2020 -1405 2060 -1400
rect 2020 -1440 2060 -1435
rect 2020 -1470 2025 -1440
rect 2025 -1470 2055 -1440
rect 2055 -1470 2060 -1440
rect 2020 -1475 2060 -1470
rect 2020 -1510 2060 -1505
rect 2020 -1540 2025 -1510
rect 2025 -1540 2055 -1510
rect 2055 -1540 2060 -1510
rect 2020 -1545 2060 -1540
rect 2020 -1580 2060 -1575
rect 2020 -1610 2025 -1580
rect 2025 -1610 2055 -1580
rect 2055 -1610 2060 -1580
rect 2020 -1615 2060 -1610
rect 2020 -1645 2060 -1640
rect 2020 -1675 2025 -1645
rect 2025 -1675 2055 -1645
rect 2055 -1675 2060 -1645
rect 2020 -1680 2060 -1675
rect 2020 -1705 2060 -1700
rect 2020 -1735 2025 -1705
rect 2025 -1735 2055 -1705
rect 2055 -1735 2060 -1705
rect 2020 -1740 2060 -1735
rect 2020 -1770 2060 -1765
rect 2020 -1800 2025 -1770
rect 2025 -1800 2055 -1770
rect 2055 -1800 2060 -1770
rect 2020 -1805 2060 -1800
rect 2020 -1840 2060 -1835
rect 2020 -1870 2025 -1840
rect 2025 -1870 2055 -1840
rect 2055 -1870 2060 -1840
rect 2020 -1875 2060 -1870
rect 2020 -1910 2060 -1905
rect 2020 -1940 2025 -1910
rect 2025 -1940 2055 -1910
rect 2055 -1940 2060 -1910
rect 2020 -1945 2060 -1940
rect 2020 -1980 2060 -1975
rect 2020 -2010 2025 -1980
rect 2025 -2010 2055 -1980
rect 2055 -2010 2060 -1980
rect 2020 -2015 2060 -2010
rect 2020 -2045 2060 -2040
rect 2020 -2075 2025 -2045
rect 2025 -2075 2055 -2045
rect 2055 -2075 2060 -2045
rect 2020 -2080 2060 -2075
rect 2020 -2105 2060 -2100
rect 2020 -2135 2025 -2105
rect 2025 -2135 2055 -2105
rect 2055 -2135 2060 -2105
rect 2020 -2140 2060 -2135
rect 2020 -2170 2060 -2165
rect 2020 -2200 2025 -2170
rect 2025 -2200 2055 -2170
rect 2055 -2200 2060 -2170
rect 2020 -2205 2060 -2200
rect 2020 -2240 2060 -2235
rect 2020 -2270 2025 -2240
rect 2025 -2270 2055 -2240
rect 2055 -2270 2060 -2240
rect 2020 -2275 2060 -2270
rect 2020 -2310 2060 -2305
rect 2020 -2340 2025 -2310
rect 2025 -2340 2055 -2310
rect 2055 -2340 2060 -2310
rect 2020 -2345 2060 -2340
rect 2020 -2380 2060 -2375
rect 2020 -2410 2025 -2380
rect 2025 -2410 2055 -2380
rect 2055 -2410 2060 -2380
rect 2020 -2415 2060 -2410
rect 2020 -2445 2060 -2440
rect 2020 -2475 2025 -2445
rect 2025 -2475 2055 -2445
rect 2055 -2475 2060 -2445
rect 2020 -2480 2060 -2475
rect 2020 -2505 2060 -2500
rect 2020 -2535 2025 -2505
rect 2025 -2535 2055 -2505
rect 2055 -2535 2060 -2505
rect 2020 -2540 2060 -2535
rect 2020 -2570 2060 -2565
rect 2020 -2600 2025 -2570
rect 2025 -2600 2055 -2570
rect 2055 -2600 2060 -2570
rect 2020 -2605 2060 -2600
rect 2020 -2640 2060 -2635
rect 2020 -2670 2025 -2640
rect 2025 -2670 2055 -2640
rect 2055 -2670 2060 -2640
rect 2020 -2675 2060 -2670
rect 2020 -2710 2060 -2705
rect 2020 -2740 2025 -2710
rect 2025 -2740 2055 -2710
rect 2055 -2740 2060 -2710
rect 2020 -2745 2060 -2740
rect 2020 -2780 2060 -2775
rect 2020 -2810 2025 -2780
rect 2025 -2810 2055 -2780
rect 2055 -2810 2060 -2780
rect 2020 -2815 2060 -2810
rect 2020 -2845 2060 -2840
rect 2020 -2875 2025 -2845
rect 2025 -2875 2055 -2845
rect 2055 -2875 2060 -2845
rect 2020 -2880 2060 -2875
rect 2020 -2905 2060 -2900
rect 2020 -2935 2025 -2905
rect 2025 -2935 2055 -2905
rect 2055 -2935 2060 -2905
rect 2020 -2940 2060 -2935
rect 2020 -2970 2060 -2965
rect 2020 -3000 2025 -2970
rect 2025 -3000 2055 -2970
rect 2055 -3000 2060 -2970
rect 2020 -3005 2060 -3000
rect 2020 -3040 2060 -3035
rect 2020 -3070 2025 -3040
rect 2025 -3070 2055 -3040
rect 2055 -3070 2060 -3040
rect 2020 -3075 2060 -3070
rect 2020 -3110 2060 -3105
rect 2020 -3140 2025 -3110
rect 2025 -3140 2055 -3110
rect 2055 -3140 2060 -3110
rect 2020 -3145 2060 -3140
rect 2020 -3180 2060 -3175
rect 2020 -3210 2025 -3180
rect 2025 -3210 2055 -3180
rect 2055 -3210 2060 -3180
rect 2020 -3215 2060 -3210
rect 2020 -3245 2060 -3240
rect 2020 -3275 2025 -3245
rect 2025 -3275 2055 -3245
rect 2055 -3275 2060 -3245
rect 2020 -3280 2060 -3275
rect 2020 -3305 2060 -3300
rect 2020 -3335 2025 -3305
rect 2025 -3335 2055 -3305
rect 2055 -3335 2060 -3305
rect 2020 -3340 2060 -3335
rect 2020 -3370 2060 -3365
rect 2020 -3400 2025 -3370
rect 2025 -3400 2055 -3370
rect 2055 -3400 2060 -3370
rect 2020 -3405 2060 -3400
rect 2020 -3440 2060 -3435
rect 2020 -3470 2025 -3440
rect 2025 -3470 2055 -3440
rect 2055 -3470 2060 -3440
rect 2020 -3475 2060 -3470
rect 2020 -3510 2060 -3505
rect 2020 -3540 2025 -3510
rect 2025 -3540 2055 -3510
rect 2055 -3540 2060 -3510
rect 2020 -3545 2060 -3540
rect 2020 -3580 2060 -3575
rect 2020 -3610 2025 -3580
rect 2025 -3610 2055 -3580
rect 2055 -3610 2060 -3580
rect 2020 -3615 2060 -3610
rect 2020 -3645 2060 -3640
rect 2020 -3675 2025 -3645
rect 2025 -3675 2055 -3645
rect 2055 -3675 2060 -3645
rect 2020 -3680 2060 -3675
rect 2020 -3705 2060 -3700
rect 2020 -3735 2025 -3705
rect 2025 -3735 2055 -3705
rect 2055 -3735 2060 -3705
rect 2020 -3740 2060 -3735
rect 2020 -3770 2060 -3765
rect 2020 -3800 2025 -3770
rect 2025 -3800 2055 -3770
rect 2055 -3800 2060 -3770
rect 2020 -3805 2060 -3800
rect 2020 -3840 2060 -3835
rect 2020 -3870 2025 -3840
rect 2025 -3870 2055 -3840
rect 2055 -3870 2060 -3840
rect 2020 -3875 2060 -3870
rect 2020 -3910 2060 -3905
rect 2020 -3940 2025 -3910
rect 2025 -3940 2055 -3910
rect 2055 -3940 2060 -3910
rect 2020 -3945 2060 -3940
rect 2020 -3980 2060 -3975
rect 2020 -4010 2025 -3980
rect 2025 -4010 2055 -3980
rect 2055 -4010 2060 -3980
rect 2020 -4015 2060 -4010
rect 2020 -4045 2060 -4040
rect 2020 -4075 2025 -4045
rect 2025 -4075 2055 -4045
rect 2055 -4075 2060 -4045
rect 2020 -4080 2060 -4075
rect 2020 -4105 2060 -4100
rect 2020 -4135 2025 -4105
rect 2025 -4135 2055 -4105
rect 2055 -4135 2060 -4105
rect 2020 -4140 2060 -4135
rect 2020 -4170 2060 -4165
rect 2020 -4200 2025 -4170
rect 2025 -4200 2055 -4170
rect 2055 -4200 2060 -4170
rect 2020 -4205 2060 -4200
rect 2020 -4240 2060 -4235
rect 2020 -4270 2025 -4240
rect 2025 -4270 2055 -4240
rect 2055 -4270 2060 -4240
rect 2020 -4275 2060 -4270
rect 2020 -4310 2060 -4305
rect 2020 -4340 2025 -4310
rect 2025 -4340 2055 -4310
rect 2055 -4340 2060 -4310
rect 2020 -4345 2060 -4340
rect 2020 -4380 2060 -4375
rect 2020 -4410 2025 -4380
rect 2025 -4410 2055 -4380
rect 2055 -4410 2060 -4380
rect 2020 -4415 2060 -4410
rect 2020 -4445 2060 -4440
rect 2020 -4475 2025 -4445
rect 2025 -4475 2055 -4445
rect 2055 -4475 2060 -4445
rect 2020 -4480 2060 -4475
rect 2370 -1305 2410 -1300
rect 2370 -1335 2375 -1305
rect 2375 -1335 2405 -1305
rect 2405 -1335 2410 -1305
rect 2370 -1340 2410 -1335
rect 2370 -1370 2410 -1365
rect 2370 -1400 2375 -1370
rect 2375 -1400 2405 -1370
rect 2405 -1400 2410 -1370
rect 2370 -1405 2410 -1400
rect 2370 -1440 2410 -1435
rect 2370 -1470 2375 -1440
rect 2375 -1470 2405 -1440
rect 2405 -1470 2410 -1440
rect 2370 -1475 2410 -1470
rect 2370 -1510 2410 -1505
rect 2370 -1540 2375 -1510
rect 2375 -1540 2405 -1510
rect 2405 -1540 2410 -1510
rect 2370 -1545 2410 -1540
rect 2370 -1580 2410 -1575
rect 2370 -1610 2375 -1580
rect 2375 -1610 2405 -1580
rect 2405 -1610 2410 -1580
rect 2370 -1615 2410 -1610
rect 2370 -1645 2410 -1640
rect 2370 -1675 2375 -1645
rect 2375 -1675 2405 -1645
rect 2405 -1675 2410 -1645
rect 2370 -1680 2410 -1675
rect 2370 -1705 2410 -1700
rect 2370 -1735 2375 -1705
rect 2375 -1735 2405 -1705
rect 2405 -1735 2410 -1705
rect 2370 -1740 2410 -1735
rect 2370 -1770 2410 -1765
rect 2370 -1800 2375 -1770
rect 2375 -1800 2405 -1770
rect 2405 -1800 2410 -1770
rect 2370 -1805 2410 -1800
rect 2370 -1840 2410 -1835
rect 2370 -1870 2375 -1840
rect 2375 -1870 2405 -1840
rect 2405 -1870 2410 -1840
rect 2370 -1875 2410 -1870
rect 2370 -1910 2410 -1905
rect 2370 -1940 2375 -1910
rect 2375 -1940 2405 -1910
rect 2405 -1940 2410 -1910
rect 2370 -1945 2410 -1940
rect 2370 -1980 2410 -1975
rect 2370 -2010 2375 -1980
rect 2375 -2010 2405 -1980
rect 2405 -2010 2410 -1980
rect 2370 -2015 2410 -2010
rect 2370 -2045 2410 -2040
rect 2370 -2075 2375 -2045
rect 2375 -2075 2405 -2045
rect 2405 -2075 2410 -2045
rect 2370 -2080 2410 -2075
rect 2370 -2105 2410 -2100
rect 2370 -2135 2375 -2105
rect 2375 -2135 2405 -2105
rect 2405 -2135 2410 -2105
rect 2370 -2140 2410 -2135
rect 2370 -2170 2410 -2165
rect 2370 -2200 2375 -2170
rect 2375 -2200 2405 -2170
rect 2405 -2200 2410 -2170
rect 2370 -2205 2410 -2200
rect 2370 -2240 2410 -2235
rect 2370 -2270 2375 -2240
rect 2375 -2270 2405 -2240
rect 2405 -2270 2410 -2240
rect 2370 -2275 2410 -2270
rect 2370 -2310 2410 -2305
rect 2370 -2340 2375 -2310
rect 2375 -2340 2405 -2310
rect 2405 -2340 2410 -2310
rect 2370 -2345 2410 -2340
rect 2370 -2380 2410 -2375
rect 2370 -2410 2375 -2380
rect 2375 -2410 2405 -2380
rect 2405 -2410 2410 -2380
rect 2370 -2415 2410 -2410
rect 2370 -2445 2410 -2440
rect 2370 -2475 2375 -2445
rect 2375 -2475 2405 -2445
rect 2405 -2475 2410 -2445
rect 2370 -2480 2410 -2475
rect 2370 -2505 2410 -2500
rect 2370 -2535 2375 -2505
rect 2375 -2535 2405 -2505
rect 2405 -2535 2410 -2505
rect 2370 -2540 2410 -2535
rect 2370 -2570 2410 -2565
rect 2370 -2600 2375 -2570
rect 2375 -2600 2405 -2570
rect 2405 -2600 2410 -2570
rect 2370 -2605 2410 -2600
rect 2370 -2640 2410 -2635
rect 2370 -2670 2375 -2640
rect 2375 -2670 2405 -2640
rect 2405 -2670 2410 -2640
rect 2370 -2675 2410 -2670
rect 2370 -2710 2410 -2705
rect 2370 -2740 2375 -2710
rect 2375 -2740 2405 -2710
rect 2405 -2740 2410 -2710
rect 2370 -2745 2410 -2740
rect 2370 -2780 2410 -2775
rect 2370 -2810 2375 -2780
rect 2375 -2810 2405 -2780
rect 2405 -2810 2410 -2780
rect 2370 -2815 2410 -2810
rect 2370 -2845 2410 -2840
rect 2370 -2875 2375 -2845
rect 2375 -2875 2405 -2845
rect 2405 -2875 2410 -2845
rect 2370 -2880 2410 -2875
rect 2370 -2905 2410 -2900
rect 2370 -2935 2375 -2905
rect 2375 -2935 2405 -2905
rect 2405 -2935 2410 -2905
rect 2370 -2940 2410 -2935
rect 2370 -2970 2410 -2965
rect 2370 -3000 2375 -2970
rect 2375 -3000 2405 -2970
rect 2405 -3000 2410 -2970
rect 2370 -3005 2410 -3000
rect 2370 -3040 2410 -3035
rect 2370 -3070 2375 -3040
rect 2375 -3070 2405 -3040
rect 2405 -3070 2410 -3040
rect 2370 -3075 2410 -3070
rect 2370 -3110 2410 -3105
rect 2370 -3140 2375 -3110
rect 2375 -3140 2405 -3110
rect 2405 -3140 2410 -3110
rect 2370 -3145 2410 -3140
rect 2370 -3180 2410 -3175
rect 2370 -3210 2375 -3180
rect 2375 -3210 2405 -3180
rect 2405 -3210 2410 -3180
rect 2370 -3215 2410 -3210
rect 2370 -3245 2410 -3240
rect 2370 -3275 2375 -3245
rect 2375 -3275 2405 -3245
rect 2405 -3275 2410 -3245
rect 2370 -3280 2410 -3275
rect 2370 -3305 2410 -3300
rect 2370 -3335 2375 -3305
rect 2375 -3335 2405 -3305
rect 2405 -3335 2410 -3305
rect 2370 -3340 2410 -3335
rect 2370 -3370 2410 -3365
rect 2370 -3400 2375 -3370
rect 2375 -3400 2405 -3370
rect 2405 -3400 2410 -3370
rect 2370 -3405 2410 -3400
rect 2370 -3440 2410 -3435
rect 2370 -3470 2375 -3440
rect 2375 -3470 2405 -3440
rect 2405 -3470 2410 -3440
rect 2370 -3475 2410 -3470
rect 2370 -3510 2410 -3505
rect 2370 -3540 2375 -3510
rect 2375 -3540 2405 -3510
rect 2405 -3540 2410 -3510
rect 2370 -3545 2410 -3540
rect 2370 -3580 2410 -3575
rect 2370 -3610 2375 -3580
rect 2375 -3610 2405 -3580
rect 2405 -3610 2410 -3580
rect 2370 -3615 2410 -3610
rect 2370 -3645 2410 -3640
rect 2370 -3675 2375 -3645
rect 2375 -3675 2405 -3645
rect 2405 -3675 2410 -3645
rect 2370 -3680 2410 -3675
rect 2370 -3705 2410 -3700
rect 2370 -3735 2375 -3705
rect 2375 -3735 2405 -3705
rect 2405 -3735 2410 -3705
rect 2370 -3740 2410 -3735
rect 2370 -3770 2410 -3765
rect 2370 -3800 2375 -3770
rect 2375 -3800 2405 -3770
rect 2405 -3800 2410 -3770
rect 2370 -3805 2410 -3800
rect 2370 -3840 2410 -3835
rect 2370 -3870 2375 -3840
rect 2375 -3870 2405 -3840
rect 2405 -3870 2410 -3840
rect 2370 -3875 2410 -3870
rect 2370 -3910 2410 -3905
rect 2370 -3940 2375 -3910
rect 2375 -3940 2405 -3910
rect 2405 -3940 2410 -3910
rect 2370 -3945 2410 -3940
rect 2370 -3980 2410 -3975
rect 2370 -4010 2375 -3980
rect 2375 -4010 2405 -3980
rect 2405 -4010 2410 -3980
rect 2370 -4015 2410 -4010
rect 2370 -4045 2410 -4040
rect 2370 -4075 2375 -4045
rect 2375 -4075 2405 -4045
rect 2405 -4075 2410 -4045
rect 2370 -4080 2410 -4075
rect 2370 -4105 2410 -4100
rect 2370 -4135 2375 -4105
rect 2375 -4135 2405 -4105
rect 2405 -4135 2410 -4105
rect 2370 -4140 2410 -4135
rect 2370 -4170 2410 -4165
rect 2370 -4200 2375 -4170
rect 2375 -4200 2405 -4170
rect 2405 -4200 2410 -4170
rect 2370 -4205 2410 -4200
rect 2370 -4240 2410 -4235
rect 2370 -4270 2375 -4240
rect 2375 -4270 2405 -4240
rect 2405 -4270 2410 -4240
rect 2370 -4275 2410 -4270
rect 2370 -4310 2410 -4305
rect 2370 -4340 2375 -4310
rect 2375 -4340 2405 -4310
rect 2405 -4340 2410 -4310
rect 2370 -4345 2410 -4340
rect 2370 -4380 2410 -4375
rect 2370 -4410 2375 -4380
rect 2375 -4410 2405 -4380
rect 2405 -4410 2410 -4380
rect 2370 -4415 2410 -4410
rect 2370 -4445 2410 -4440
rect 2370 -4475 2375 -4445
rect 2375 -4475 2405 -4445
rect 2405 -4475 2410 -4445
rect 2370 -4480 2410 -4475
rect 2720 -1305 2760 -1300
rect 2720 -1335 2725 -1305
rect 2725 -1335 2755 -1305
rect 2755 -1335 2760 -1305
rect 2720 -1340 2760 -1335
rect 2720 -1370 2760 -1365
rect 2720 -1400 2725 -1370
rect 2725 -1400 2755 -1370
rect 2755 -1400 2760 -1370
rect 2720 -1405 2760 -1400
rect 2720 -1440 2760 -1435
rect 2720 -1470 2725 -1440
rect 2725 -1470 2755 -1440
rect 2755 -1470 2760 -1440
rect 2720 -1475 2760 -1470
rect 2720 -1510 2760 -1505
rect 2720 -1540 2725 -1510
rect 2725 -1540 2755 -1510
rect 2755 -1540 2760 -1510
rect 2720 -1545 2760 -1540
rect 2720 -1580 2760 -1575
rect 2720 -1610 2725 -1580
rect 2725 -1610 2755 -1580
rect 2755 -1610 2760 -1580
rect 2720 -1615 2760 -1610
rect 2720 -1645 2760 -1640
rect 2720 -1675 2725 -1645
rect 2725 -1675 2755 -1645
rect 2755 -1675 2760 -1645
rect 2720 -1680 2760 -1675
rect 2720 -1705 2760 -1700
rect 2720 -1735 2725 -1705
rect 2725 -1735 2755 -1705
rect 2755 -1735 2760 -1705
rect 2720 -1740 2760 -1735
rect 2720 -1770 2760 -1765
rect 2720 -1800 2725 -1770
rect 2725 -1800 2755 -1770
rect 2755 -1800 2760 -1770
rect 2720 -1805 2760 -1800
rect 2720 -1840 2760 -1835
rect 2720 -1870 2725 -1840
rect 2725 -1870 2755 -1840
rect 2755 -1870 2760 -1840
rect 2720 -1875 2760 -1870
rect 2720 -1910 2760 -1905
rect 2720 -1940 2725 -1910
rect 2725 -1940 2755 -1910
rect 2755 -1940 2760 -1910
rect 2720 -1945 2760 -1940
rect 2720 -1980 2760 -1975
rect 2720 -2010 2725 -1980
rect 2725 -2010 2755 -1980
rect 2755 -2010 2760 -1980
rect 2720 -2015 2760 -2010
rect 2720 -2045 2760 -2040
rect 2720 -2075 2725 -2045
rect 2725 -2075 2755 -2045
rect 2755 -2075 2760 -2045
rect 2720 -2080 2760 -2075
rect 2720 -2105 2760 -2100
rect 2720 -2135 2725 -2105
rect 2725 -2135 2755 -2105
rect 2755 -2135 2760 -2105
rect 2720 -2140 2760 -2135
rect 2720 -2170 2760 -2165
rect 2720 -2200 2725 -2170
rect 2725 -2200 2755 -2170
rect 2755 -2200 2760 -2170
rect 2720 -2205 2760 -2200
rect 2720 -2240 2760 -2235
rect 2720 -2270 2725 -2240
rect 2725 -2270 2755 -2240
rect 2755 -2270 2760 -2240
rect 2720 -2275 2760 -2270
rect 2720 -2310 2760 -2305
rect 2720 -2340 2725 -2310
rect 2725 -2340 2755 -2310
rect 2755 -2340 2760 -2310
rect 2720 -2345 2760 -2340
rect 2720 -2380 2760 -2375
rect 2720 -2410 2725 -2380
rect 2725 -2410 2755 -2380
rect 2755 -2410 2760 -2380
rect 2720 -2415 2760 -2410
rect 2720 -2445 2760 -2440
rect 2720 -2475 2725 -2445
rect 2725 -2475 2755 -2445
rect 2755 -2475 2760 -2445
rect 2720 -2480 2760 -2475
rect 2720 -2505 2760 -2500
rect 2720 -2535 2725 -2505
rect 2725 -2535 2755 -2505
rect 2755 -2535 2760 -2505
rect 2720 -2540 2760 -2535
rect 2720 -2570 2760 -2565
rect 2720 -2600 2725 -2570
rect 2725 -2600 2755 -2570
rect 2755 -2600 2760 -2570
rect 2720 -2605 2760 -2600
rect 2720 -2640 2760 -2635
rect 2720 -2670 2725 -2640
rect 2725 -2670 2755 -2640
rect 2755 -2670 2760 -2640
rect 2720 -2675 2760 -2670
rect 2720 -2710 2760 -2705
rect 2720 -2740 2725 -2710
rect 2725 -2740 2755 -2710
rect 2755 -2740 2760 -2710
rect 2720 -2745 2760 -2740
rect 2720 -2780 2760 -2775
rect 2720 -2810 2725 -2780
rect 2725 -2810 2755 -2780
rect 2755 -2810 2760 -2780
rect 2720 -2815 2760 -2810
rect 2720 -2845 2760 -2840
rect 2720 -2875 2725 -2845
rect 2725 -2875 2755 -2845
rect 2755 -2875 2760 -2845
rect 2720 -2880 2760 -2875
rect 2720 -2905 2760 -2900
rect 2720 -2935 2725 -2905
rect 2725 -2935 2755 -2905
rect 2755 -2935 2760 -2905
rect 2720 -2940 2760 -2935
rect 2720 -2970 2760 -2965
rect 2720 -3000 2725 -2970
rect 2725 -3000 2755 -2970
rect 2755 -3000 2760 -2970
rect 2720 -3005 2760 -3000
rect 2720 -3040 2760 -3035
rect 2720 -3070 2725 -3040
rect 2725 -3070 2755 -3040
rect 2755 -3070 2760 -3040
rect 2720 -3075 2760 -3070
rect 2720 -3110 2760 -3105
rect 2720 -3140 2725 -3110
rect 2725 -3140 2755 -3110
rect 2755 -3140 2760 -3110
rect 2720 -3145 2760 -3140
rect 2720 -3180 2760 -3175
rect 2720 -3210 2725 -3180
rect 2725 -3210 2755 -3180
rect 2755 -3210 2760 -3180
rect 2720 -3215 2760 -3210
rect 2720 -3245 2760 -3240
rect 2720 -3275 2725 -3245
rect 2725 -3275 2755 -3245
rect 2755 -3275 2760 -3245
rect 2720 -3280 2760 -3275
rect 2720 -3305 2760 -3300
rect 2720 -3335 2725 -3305
rect 2725 -3335 2755 -3305
rect 2755 -3335 2760 -3305
rect 2720 -3340 2760 -3335
rect 2720 -3370 2760 -3365
rect 2720 -3400 2725 -3370
rect 2725 -3400 2755 -3370
rect 2755 -3400 2760 -3370
rect 2720 -3405 2760 -3400
rect 2720 -3440 2760 -3435
rect 2720 -3470 2725 -3440
rect 2725 -3470 2755 -3440
rect 2755 -3470 2760 -3440
rect 2720 -3475 2760 -3470
rect 2720 -3510 2760 -3505
rect 2720 -3540 2725 -3510
rect 2725 -3540 2755 -3510
rect 2755 -3540 2760 -3510
rect 2720 -3545 2760 -3540
rect 2720 -3580 2760 -3575
rect 2720 -3610 2725 -3580
rect 2725 -3610 2755 -3580
rect 2755 -3610 2760 -3580
rect 2720 -3615 2760 -3610
rect 2720 -3645 2760 -3640
rect 2720 -3675 2725 -3645
rect 2725 -3675 2755 -3645
rect 2755 -3675 2760 -3645
rect 2720 -3680 2760 -3675
rect 2720 -3705 2760 -3700
rect 2720 -3735 2725 -3705
rect 2725 -3735 2755 -3705
rect 2755 -3735 2760 -3705
rect 2720 -3740 2760 -3735
rect 2720 -3770 2760 -3765
rect 2720 -3800 2725 -3770
rect 2725 -3800 2755 -3770
rect 2755 -3800 2760 -3770
rect 2720 -3805 2760 -3800
rect 2720 -3840 2760 -3835
rect 2720 -3870 2725 -3840
rect 2725 -3870 2755 -3840
rect 2755 -3870 2760 -3840
rect 2720 -3875 2760 -3870
rect 2720 -3910 2760 -3905
rect 2720 -3940 2725 -3910
rect 2725 -3940 2755 -3910
rect 2755 -3940 2760 -3910
rect 2720 -3945 2760 -3940
rect 2720 -3980 2760 -3975
rect 2720 -4010 2725 -3980
rect 2725 -4010 2755 -3980
rect 2755 -4010 2760 -3980
rect 2720 -4015 2760 -4010
rect 2720 -4045 2760 -4040
rect 2720 -4075 2725 -4045
rect 2725 -4075 2755 -4045
rect 2755 -4075 2760 -4045
rect 2720 -4080 2760 -4075
rect 2720 -4105 2760 -4100
rect 2720 -4135 2725 -4105
rect 2725 -4135 2755 -4105
rect 2755 -4135 2760 -4105
rect 2720 -4140 2760 -4135
rect 2720 -4170 2760 -4165
rect 2720 -4200 2725 -4170
rect 2725 -4200 2755 -4170
rect 2755 -4200 2760 -4170
rect 2720 -4205 2760 -4200
rect 2720 -4240 2760 -4235
rect 2720 -4270 2725 -4240
rect 2725 -4270 2755 -4240
rect 2755 -4270 2760 -4240
rect 2720 -4275 2760 -4270
rect 2720 -4310 2760 -4305
rect 2720 -4340 2725 -4310
rect 2725 -4340 2755 -4310
rect 2755 -4340 2760 -4310
rect 2720 -4345 2760 -4340
rect 2720 -4380 2760 -4375
rect 2720 -4410 2725 -4380
rect 2725 -4410 2755 -4380
rect 2755 -4410 2760 -4380
rect 2720 -4415 2760 -4410
rect 2720 -4445 2760 -4440
rect 2720 -4475 2725 -4445
rect 2725 -4475 2755 -4445
rect 2755 -4475 2760 -4445
rect 2720 -4480 2760 -4475
rect 3070 -1305 3110 -1300
rect 3070 -1335 3075 -1305
rect 3075 -1335 3105 -1305
rect 3105 -1335 3110 -1305
rect 3070 -1340 3110 -1335
rect 3070 -1370 3110 -1365
rect 3070 -1400 3075 -1370
rect 3075 -1400 3105 -1370
rect 3105 -1400 3110 -1370
rect 3070 -1405 3110 -1400
rect 3070 -1440 3110 -1435
rect 3070 -1470 3075 -1440
rect 3075 -1470 3105 -1440
rect 3105 -1470 3110 -1440
rect 3070 -1475 3110 -1470
rect 3070 -1510 3110 -1505
rect 3070 -1540 3075 -1510
rect 3075 -1540 3105 -1510
rect 3105 -1540 3110 -1510
rect 3070 -1545 3110 -1540
rect 3070 -1580 3110 -1575
rect 3070 -1610 3075 -1580
rect 3075 -1610 3105 -1580
rect 3105 -1610 3110 -1580
rect 3070 -1615 3110 -1610
rect 3070 -1645 3110 -1640
rect 3070 -1675 3075 -1645
rect 3075 -1675 3105 -1645
rect 3105 -1675 3110 -1645
rect 3070 -1680 3110 -1675
rect 3070 -1705 3110 -1700
rect 3070 -1735 3075 -1705
rect 3075 -1735 3105 -1705
rect 3105 -1735 3110 -1705
rect 3070 -1740 3110 -1735
rect 3070 -1770 3110 -1765
rect 3070 -1800 3075 -1770
rect 3075 -1800 3105 -1770
rect 3105 -1800 3110 -1770
rect 3070 -1805 3110 -1800
rect 3070 -1840 3110 -1835
rect 3070 -1870 3075 -1840
rect 3075 -1870 3105 -1840
rect 3105 -1870 3110 -1840
rect 3070 -1875 3110 -1870
rect 3070 -1910 3110 -1905
rect 3070 -1940 3075 -1910
rect 3075 -1940 3105 -1910
rect 3105 -1940 3110 -1910
rect 3070 -1945 3110 -1940
rect 3070 -1980 3110 -1975
rect 3070 -2010 3075 -1980
rect 3075 -2010 3105 -1980
rect 3105 -2010 3110 -1980
rect 3070 -2015 3110 -2010
rect 3070 -2045 3110 -2040
rect 3070 -2075 3075 -2045
rect 3075 -2075 3105 -2045
rect 3105 -2075 3110 -2045
rect 3070 -2080 3110 -2075
rect 3070 -2105 3110 -2100
rect 3070 -2135 3075 -2105
rect 3075 -2135 3105 -2105
rect 3105 -2135 3110 -2105
rect 3070 -2140 3110 -2135
rect 3070 -2170 3110 -2165
rect 3070 -2200 3075 -2170
rect 3075 -2200 3105 -2170
rect 3105 -2200 3110 -2170
rect 3070 -2205 3110 -2200
rect 3070 -2240 3110 -2235
rect 3070 -2270 3075 -2240
rect 3075 -2270 3105 -2240
rect 3105 -2270 3110 -2240
rect 3070 -2275 3110 -2270
rect 3070 -2310 3110 -2305
rect 3070 -2340 3075 -2310
rect 3075 -2340 3105 -2310
rect 3105 -2340 3110 -2310
rect 3070 -2345 3110 -2340
rect 3070 -2380 3110 -2375
rect 3070 -2410 3075 -2380
rect 3075 -2410 3105 -2380
rect 3105 -2410 3110 -2380
rect 3070 -2415 3110 -2410
rect 3070 -2445 3110 -2440
rect 3070 -2475 3075 -2445
rect 3075 -2475 3105 -2445
rect 3105 -2475 3110 -2445
rect 3070 -2480 3110 -2475
rect 3070 -2505 3110 -2500
rect 3070 -2535 3075 -2505
rect 3075 -2535 3105 -2505
rect 3105 -2535 3110 -2505
rect 3070 -2540 3110 -2535
rect 3070 -2570 3110 -2565
rect 3070 -2600 3075 -2570
rect 3075 -2600 3105 -2570
rect 3105 -2600 3110 -2570
rect 3070 -2605 3110 -2600
rect 3070 -2640 3110 -2635
rect 3070 -2670 3075 -2640
rect 3075 -2670 3105 -2640
rect 3105 -2670 3110 -2640
rect 3070 -2675 3110 -2670
rect 3070 -2710 3110 -2705
rect 3070 -2740 3075 -2710
rect 3075 -2740 3105 -2710
rect 3105 -2740 3110 -2710
rect 3070 -2745 3110 -2740
rect 3070 -2780 3110 -2775
rect 3070 -2810 3075 -2780
rect 3075 -2810 3105 -2780
rect 3105 -2810 3110 -2780
rect 3070 -2815 3110 -2810
rect 3070 -2845 3110 -2840
rect 3070 -2875 3075 -2845
rect 3075 -2875 3105 -2845
rect 3105 -2875 3110 -2845
rect 3070 -2880 3110 -2875
rect 3070 -2905 3110 -2900
rect 3070 -2935 3075 -2905
rect 3075 -2935 3105 -2905
rect 3105 -2935 3110 -2905
rect 3070 -2940 3110 -2935
rect 3070 -2970 3110 -2965
rect 3070 -3000 3075 -2970
rect 3075 -3000 3105 -2970
rect 3105 -3000 3110 -2970
rect 3070 -3005 3110 -3000
rect 3070 -3040 3110 -3035
rect 3070 -3070 3075 -3040
rect 3075 -3070 3105 -3040
rect 3105 -3070 3110 -3040
rect 3070 -3075 3110 -3070
rect 3070 -3110 3110 -3105
rect 3070 -3140 3075 -3110
rect 3075 -3140 3105 -3110
rect 3105 -3140 3110 -3110
rect 3070 -3145 3110 -3140
rect 3070 -3180 3110 -3175
rect 3070 -3210 3075 -3180
rect 3075 -3210 3105 -3180
rect 3105 -3210 3110 -3180
rect 3070 -3215 3110 -3210
rect 3070 -3245 3110 -3240
rect 3070 -3275 3075 -3245
rect 3075 -3275 3105 -3245
rect 3105 -3275 3110 -3245
rect 3070 -3280 3110 -3275
rect 3070 -3305 3110 -3300
rect 3070 -3335 3075 -3305
rect 3075 -3335 3105 -3305
rect 3105 -3335 3110 -3305
rect 3070 -3340 3110 -3335
rect 3070 -3370 3110 -3365
rect 3070 -3400 3075 -3370
rect 3075 -3400 3105 -3370
rect 3105 -3400 3110 -3370
rect 3070 -3405 3110 -3400
rect 3070 -3440 3110 -3435
rect 3070 -3470 3075 -3440
rect 3075 -3470 3105 -3440
rect 3105 -3470 3110 -3440
rect 3070 -3475 3110 -3470
rect 3070 -3510 3110 -3505
rect 3070 -3540 3075 -3510
rect 3075 -3540 3105 -3510
rect 3105 -3540 3110 -3510
rect 3070 -3545 3110 -3540
rect 3070 -3580 3110 -3575
rect 3070 -3610 3075 -3580
rect 3075 -3610 3105 -3580
rect 3105 -3610 3110 -3580
rect 3070 -3615 3110 -3610
rect 3070 -3645 3110 -3640
rect 3070 -3675 3075 -3645
rect 3075 -3675 3105 -3645
rect 3105 -3675 3110 -3645
rect 3070 -3680 3110 -3675
rect 3070 -3705 3110 -3700
rect 3070 -3735 3075 -3705
rect 3075 -3735 3105 -3705
rect 3105 -3735 3110 -3705
rect 3070 -3740 3110 -3735
rect 3070 -3770 3110 -3765
rect 3070 -3800 3075 -3770
rect 3075 -3800 3105 -3770
rect 3105 -3800 3110 -3770
rect 3070 -3805 3110 -3800
rect 3070 -3840 3110 -3835
rect 3070 -3870 3075 -3840
rect 3075 -3870 3105 -3840
rect 3105 -3870 3110 -3840
rect 3070 -3875 3110 -3870
rect 3070 -3910 3110 -3905
rect 3070 -3940 3075 -3910
rect 3075 -3940 3105 -3910
rect 3105 -3940 3110 -3910
rect 3070 -3945 3110 -3940
rect 3070 -3980 3110 -3975
rect 3070 -4010 3075 -3980
rect 3075 -4010 3105 -3980
rect 3105 -4010 3110 -3980
rect 3070 -4015 3110 -4010
rect 3070 -4045 3110 -4040
rect 3070 -4075 3075 -4045
rect 3075 -4075 3105 -4045
rect 3105 -4075 3110 -4045
rect 3070 -4080 3110 -4075
rect 3070 -4105 3110 -4100
rect 3070 -4135 3075 -4105
rect 3075 -4135 3105 -4105
rect 3105 -4135 3110 -4105
rect 3070 -4140 3110 -4135
rect 3070 -4170 3110 -4165
rect 3070 -4200 3075 -4170
rect 3075 -4200 3105 -4170
rect 3105 -4200 3110 -4170
rect 3070 -4205 3110 -4200
rect 3070 -4240 3110 -4235
rect 3070 -4270 3075 -4240
rect 3075 -4270 3105 -4240
rect 3105 -4270 3110 -4240
rect 3070 -4275 3110 -4270
rect 3070 -4310 3110 -4305
rect 3070 -4340 3075 -4310
rect 3075 -4340 3105 -4310
rect 3105 -4340 3110 -4310
rect 3070 -4345 3110 -4340
rect 3070 -4380 3110 -4375
rect 3070 -4410 3075 -4380
rect 3075 -4410 3105 -4380
rect 3105 -4410 3110 -4380
rect 3070 -4415 3110 -4410
rect 3070 -4445 3110 -4440
rect 3070 -4475 3075 -4445
rect 3075 -4475 3105 -4445
rect 3105 -4475 3110 -4445
rect 3070 -4480 3110 -4475
rect 3420 -1305 3460 -1300
rect 3420 -1335 3425 -1305
rect 3425 -1335 3455 -1305
rect 3455 -1335 3460 -1305
rect 3420 -1340 3460 -1335
rect 3420 -1370 3460 -1365
rect 3420 -1400 3425 -1370
rect 3425 -1400 3455 -1370
rect 3455 -1400 3460 -1370
rect 3420 -1405 3460 -1400
rect 3420 -1440 3460 -1435
rect 3420 -1470 3425 -1440
rect 3425 -1470 3455 -1440
rect 3455 -1470 3460 -1440
rect 3420 -1475 3460 -1470
rect 3420 -1510 3460 -1505
rect 3420 -1540 3425 -1510
rect 3425 -1540 3455 -1510
rect 3455 -1540 3460 -1510
rect 3420 -1545 3460 -1540
rect 3420 -1580 3460 -1575
rect 3420 -1610 3425 -1580
rect 3425 -1610 3455 -1580
rect 3455 -1610 3460 -1580
rect 3420 -1615 3460 -1610
rect 3420 -1645 3460 -1640
rect 3420 -1675 3425 -1645
rect 3425 -1675 3455 -1645
rect 3455 -1675 3460 -1645
rect 3420 -1680 3460 -1675
rect 3420 -1705 3460 -1700
rect 3420 -1735 3425 -1705
rect 3425 -1735 3455 -1705
rect 3455 -1735 3460 -1705
rect 3420 -1740 3460 -1735
rect 3420 -1770 3460 -1765
rect 3420 -1800 3425 -1770
rect 3425 -1800 3455 -1770
rect 3455 -1800 3460 -1770
rect 3420 -1805 3460 -1800
rect 3420 -1840 3460 -1835
rect 3420 -1870 3425 -1840
rect 3425 -1870 3455 -1840
rect 3455 -1870 3460 -1840
rect 3420 -1875 3460 -1870
rect 3420 -1910 3460 -1905
rect 3420 -1940 3425 -1910
rect 3425 -1940 3455 -1910
rect 3455 -1940 3460 -1910
rect 3420 -1945 3460 -1940
rect 3420 -1980 3460 -1975
rect 3420 -2010 3425 -1980
rect 3425 -2010 3455 -1980
rect 3455 -2010 3460 -1980
rect 3420 -2015 3460 -2010
rect 3420 -2045 3460 -2040
rect 3420 -2075 3425 -2045
rect 3425 -2075 3455 -2045
rect 3455 -2075 3460 -2045
rect 3420 -2080 3460 -2075
rect 3420 -2105 3460 -2100
rect 3420 -2135 3425 -2105
rect 3425 -2135 3455 -2105
rect 3455 -2135 3460 -2105
rect 3420 -2140 3460 -2135
rect 3420 -2170 3460 -2165
rect 3420 -2200 3425 -2170
rect 3425 -2200 3455 -2170
rect 3455 -2200 3460 -2170
rect 3420 -2205 3460 -2200
rect 3420 -2240 3460 -2235
rect 3420 -2270 3425 -2240
rect 3425 -2270 3455 -2240
rect 3455 -2270 3460 -2240
rect 3420 -2275 3460 -2270
rect 3420 -2310 3460 -2305
rect 3420 -2340 3425 -2310
rect 3425 -2340 3455 -2310
rect 3455 -2340 3460 -2310
rect 3420 -2345 3460 -2340
rect 3420 -2380 3460 -2375
rect 3420 -2410 3425 -2380
rect 3425 -2410 3455 -2380
rect 3455 -2410 3460 -2380
rect 3420 -2415 3460 -2410
rect 3420 -2445 3460 -2440
rect 3420 -2475 3425 -2445
rect 3425 -2475 3455 -2445
rect 3455 -2475 3460 -2445
rect 3420 -2480 3460 -2475
rect 3420 -2505 3460 -2500
rect 3420 -2535 3425 -2505
rect 3425 -2535 3455 -2505
rect 3455 -2535 3460 -2505
rect 3420 -2540 3460 -2535
rect 3420 -2570 3460 -2565
rect 3420 -2600 3425 -2570
rect 3425 -2600 3455 -2570
rect 3455 -2600 3460 -2570
rect 3420 -2605 3460 -2600
rect 3420 -2640 3460 -2635
rect 3420 -2670 3425 -2640
rect 3425 -2670 3455 -2640
rect 3455 -2670 3460 -2640
rect 3420 -2675 3460 -2670
rect 3420 -2710 3460 -2705
rect 3420 -2740 3425 -2710
rect 3425 -2740 3455 -2710
rect 3455 -2740 3460 -2710
rect 3420 -2745 3460 -2740
rect 3420 -2780 3460 -2775
rect 3420 -2810 3425 -2780
rect 3425 -2810 3455 -2780
rect 3455 -2810 3460 -2780
rect 3420 -2815 3460 -2810
rect 3420 -2845 3460 -2840
rect 3420 -2875 3425 -2845
rect 3425 -2875 3455 -2845
rect 3455 -2875 3460 -2845
rect 3420 -2880 3460 -2875
rect 3420 -2905 3460 -2900
rect 3420 -2935 3425 -2905
rect 3425 -2935 3455 -2905
rect 3455 -2935 3460 -2905
rect 3420 -2940 3460 -2935
rect 3420 -2970 3460 -2965
rect 3420 -3000 3425 -2970
rect 3425 -3000 3455 -2970
rect 3455 -3000 3460 -2970
rect 3420 -3005 3460 -3000
rect 3420 -3040 3460 -3035
rect 3420 -3070 3425 -3040
rect 3425 -3070 3455 -3040
rect 3455 -3070 3460 -3040
rect 3420 -3075 3460 -3070
rect 3420 -3110 3460 -3105
rect 3420 -3140 3425 -3110
rect 3425 -3140 3455 -3110
rect 3455 -3140 3460 -3110
rect 3420 -3145 3460 -3140
rect 3420 -3180 3460 -3175
rect 3420 -3210 3425 -3180
rect 3425 -3210 3455 -3180
rect 3455 -3210 3460 -3180
rect 3420 -3215 3460 -3210
rect 3420 -3245 3460 -3240
rect 3420 -3275 3425 -3245
rect 3425 -3275 3455 -3245
rect 3455 -3275 3460 -3245
rect 3420 -3280 3460 -3275
rect 3420 -3305 3460 -3300
rect 3420 -3335 3425 -3305
rect 3425 -3335 3455 -3305
rect 3455 -3335 3460 -3305
rect 3420 -3340 3460 -3335
rect 3420 -3370 3460 -3365
rect 3420 -3400 3425 -3370
rect 3425 -3400 3455 -3370
rect 3455 -3400 3460 -3370
rect 3420 -3405 3460 -3400
rect 3420 -3440 3460 -3435
rect 3420 -3470 3425 -3440
rect 3425 -3470 3455 -3440
rect 3455 -3470 3460 -3440
rect 3420 -3475 3460 -3470
rect 3420 -3510 3460 -3505
rect 3420 -3540 3425 -3510
rect 3425 -3540 3455 -3510
rect 3455 -3540 3460 -3510
rect 3420 -3545 3460 -3540
rect 3420 -3580 3460 -3575
rect 3420 -3610 3425 -3580
rect 3425 -3610 3455 -3580
rect 3455 -3610 3460 -3580
rect 3420 -3615 3460 -3610
rect 3420 -3645 3460 -3640
rect 3420 -3675 3425 -3645
rect 3425 -3675 3455 -3645
rect 3455 -3675 3460 -3645
rect 3420 -3680 3460 -3675
rect 3420 -3705 3460 -3700
rect 3420 -3735 3425 -3705
rect 3425 -3735 3455 -3705
rect 3455 -3735 3460 -3705
rect 3420 -3740 3460 -3735
rect 3420 -3770 3460 -3765
rect 3420 -3800 3425 -3770
rect 3425 -3800 3455 -3770
rect 3455 -3800 3460 -3770
rect 3420 -3805 3460 -3800
rect 3420 -3840 3460 -3835
rect 3420 -3870 3425 -3840
rect 3425 -3870 3455 -3840
rect 3455 -3870 3460 -3840
rect 3420 -3875 3460 -3870
rect 3420 -3910 3460 -3905
rect 3420 -3940 3425 -3910
rect 3425 -3940 3455 -3910
rect 3455 -3940 3460 -3910
rect 3420 -3945 3460 -3940
rect 3420 -3980 3460 -3975
rect 3420 -4010 3425 -3980
rect 3425 -4010 3455 -3980
rect 3455 -4010 3460 -3980
rect 3420 -4015 3460 -4010
rect 3420 -4045 3460 -4040
rect 3420 -4075 3425 -4045
rect 3425 -4075 3455 -4045
rect 3455 -4075 3460 -4045
rect 3420 -4080 3460 -4075
rect 3420 -4105 3460 -4100
rect 3420 -4135 3425 -4105
rect 3425 -4135 3455 -4105
rect 3455 -4135 3460 -4105
rect 3420 -4140 3460 -4135
rect 3420 -4170 3460 -4165
rect 3420 -4200 3425 -4170
rect 3425 -4200 3455 -4170
rect 3455 -4200 3460 -4170
rect 3420 -4205 3460 -4200
rect 3420 -4240 3460 -4235
rect 3420 -4270 3425 -4240
rect 3425 -4270 3455 -4240
rect 3455 -4270 3460 -4240
rect 3420 -4275 3460 -4270
rect 3420 -4310 3460 -4305
rect 3420 -4340 3425 -4310
rect 3425 -4340 3455 -4310
rect 3455 -4340 3460 -4310
rect 3420 -4345 3460 -4340
rect 3420 -4380 3460 -4375
rect 3420 -4410 3425 -4380
rect 3425 -4410 3455 -4380
rect 3455 -4410 3460 -4380
rect 3420 -4415 3460 -4410
rect 3420 -4445 3460 -4440
rect 3420 -4475 3425 -4445
rect 3425 -4475 3455 -4445
rect 3455 -4475 3460 -4445
rect 3420 -4480 3460 -4475
rect 3770 -1305 3810 -1300
rect 3770 -1335 3775 -1305
rect 3775 -1335 3805 -1305
rect 3805 -1335 3810 -1305
rect 3770 -1340 3810 -1335
rect 3770 -1370 3810 -1365
rect 3770 -1400 3775 -1370
rect 3775 -1400 3805 -1370
rect 3805 -1400 3810 -1370
rect 3770 -1405 3810 -1400
rect 3770 -1440 3810 -1435
rect 3770 -1470 3775 -1440
rect 3775 -1470 3805 -1440
rect 3805 -1470 3810 -1440
rect 3770 -1475 3810 -1470
rect 3770 -1510 3810 -1505
rect 3770 -1540 3775 -1510
rect 3775 -1540 3805 -1510
rect 3805 -1540 3810 -1510
rect 3770 -1545 3810 -1540
rect 3770 -1580 3810 -1575
rect 3770 -1610 3775 -1580
rect 3775 -1610 3805 -1580
rect 3805 -1610 3810 -1580
rect 3770 -1615 3810 -1610
rect 3770 -1645 3810 -1640
rect 3770 -1675 3775 -1645
rect 3775 -1675 3805 -1645
rect 3805 -1675 3810 -1645
rect 3770 -1680 3810 -1675
rect 3770 -1705 3810 -1700
rect 3770 -1735 3775 -1705
rect 3775 -1735 3805 -1705
rect 3805 -1735 3810 -1705
rect 3770 -1740 3810 -1735
rect 3770 -1770 3810 -1765
rect 3770 -1800 3775 -1770
rect 3775 -1800 3805 -1770
rect 3805 -1800 3810 -1770
rect 3770 -1805 3810 -1800
rect 3770 -1840 3810 -1835
rect 3770 -1870 3775 -1840
rect 3775 -1870 3805 -1840
rect 3805 -1870 3810 -1840
rect 3770 -1875 3810 -1870
rect 3770 -1910 3810 -1905
rect 3770 -1940 3775 -1910
rect 3775 -1940 3805 -1910
rect 3805 -1940 3810 -1910
rect 3770 -1945 3810 -1940
rect 3770 -1980 3810 -1975
rect 3770 -2010 3775 -1980
rect 3775 -2010 3805 -1980
rect 3805 -2010 3810 -1980
rect 3770 -2015 3810 -2010
rect 3770 -2045 3810 -2040
rect 3770 -2075 3775 -2045
rect 3775 -2075 3805 -2045
rect 3805 -2075 3810 -2045
rect 3770 -2080 3810 -2075
rect 3770 -2105 3810 -2100
rect 3770 -2135 3775 -2105
rect 3775 -2135 3805 -2105
rect 3805 -2135 3810 -2105
rect 3770 -2140 3810 -2135
rect 3770 -2170 3810 -2165
rect 3770 -2200 3775 -2170
rect 3775 -2200 3805 -2170
rect 3805 -2200 3810 -2170
rect 3770 -2205 3810 -2200
rect 3770 -2240 3810 -2235
rect 3770 -2270 3775 -2240
rect 3775 -2270 3805 -2240
rect 3805 -2270 3810 -2240
rect 3770 -2275 3810 -2270
rect 3770 -2310 3810 -2305
rect 3770 -2340 3775 -2310
rect 3775 -2340 3805 -2310
rect 3805 -2340 3810 -2310
rect 3770 -2345 3810 -2340
rect 3770 -2380 3810 -2375
rect 3770 -2410 3775 -2380
rect 3775 -2410 3805 -2380
rect 3805 -2410 3810 -2380
rect 3770 -2415 3810 -2410
rect 3770 -2445 3810 -2440
rect 3770 -2475 3775 -2445
rect 3775 -2475 3805 -2445
rect 3805 -2475 3810 -2445
rect 3770 -2480 3810 -2475
rect 3770 -2505 3810 -2500
rect 3770 -2535 3775 -2505
rect 3775 -2535 3805 -2505
rect 3805 -2535 3810 -2505
rect 3770 -2540 3810 -2535
rect 3770 -2570 3810 -2565
rect 3770 -2600 3775 -2570
rect 3775 -2600 3805 -2570
rect 3805 -2600 3810 -2570
rect 3770 -2605 3810 -2600
rect 3770 -2640 3810 -2635
rect 3770 -2670 3775 -2640
rect 3775 -2670 3805 -2640
rect 3805 -2670 3810 -2640
rect 3770 -2675 3810 -2670
rect 3770 -2710 3810 -2705
rect 3770 -2740 3775 -2710
rect 3775 -2740 3805 -2710
rect 3805 -2740 3810 -2710
rect 3770 -2745 3810 -2740
rect 3770 -2780 3810 -2775
rect 3770 -2810 3775 -2780
rect 3775 -2810 3805 -2780
rect 3805 -2810 3810 -2780
rect 3770 -2815 3810 -2810
rect 3770 -2845 3810 -2840
rect 3770 -2875 3775 -2845
rect 3775 -2875 3805 -2845
rect 3805 -2875 3810 -2845
rect 3770 -2880 3810 -2875
rect 3770 -2905 3810 -2900
rect 3770 -2935 3775 -2905
rect 3775 -2935 3805 -2905
rect 3805 -2935 3810 -2905
rect 3770 -2940 3810 -2935
rect 3770 -2970 3810 -2965
rect 3770 -3000 3775 -2970
rect 3775 -3000 3805 -2970
rect 3805 -3000 3810 -2970
rect 3770 -3005 3810 -3000
rect 3770 -3040 3810 -3035
rect 3770 -3070 3775 -3040
rect 3775 -3070 3805 -3040
rect 3805 -3070 3810 -3040
rect 3770 -3075 3810 -3070
rect 3770 -3110 3810 -3105
rect 3770 -3140 3775 -3110
rect 3775 -3140 3805 -3110
rect 3805 -3140 3810 -3110
rect 3770 -3145 3810 -3140
rect 3770 -3180 3810 -3175
rect 3770 -3210 3775 -3180
rect 3775 -3210 3805 -3180
rect 3805 -3210 3810 -3180
rect 3770 -3215 3810 -3210
rect 3770 -3245 3810 -3240
rect 3770 -3275 3775 -3245
rect 3775 -3275 3805 -3245
rect 3805 -3275 3810 -3245
rect 3770 -3280 3810 -3275
rect 3770 -3305 3810 -3300
rect 3770 -3335 3775 -3305
rect 3775 -3335 3805 -3305
rect 3805 -3335 3810 -3305
rect 3770 -3340 3810 -3335
rect 3770 -3370 3810 -3365
rect 3770 -3400 3775 -3370
rect 3775 -3400 3805 -3370
rect 3805 -3400 3810 -3370
rect 3770 -3405 3810 -3400
rect 3770 -3440 3810 -3435
rect 3770 -3470 3775 -3440
rect 3775 -3470 3805 -3440
rect 3805 -3470 3810 -3440
rect 3770 -3475 3810 -3470
rect 3770 -3510 3810 -3505
rect 3770 -3540 3775 -3510
rect 3775 -3540 3805 -3510
rect 3805 -3540 3810 -3510
rect 3770 -3545 3810 -3540
rect 3770 -3580 3810 -3575
rect 3770 -3610 3775 -3580
rect 3775 -3610 3805 -3580
rect 3805 -3610 3810 -3580
rect 3770 -3615 3810 -3610
rect 3770 -3645 3810 -3640
rect 3770 -3675 3775 -3645
rect 3775 -3675 3805 -3645
rect 3805 -3675 3810 -3645
rect 3770 -3680 3810 -3675
rect 3770 -3705 3810 -3700
rect 3770 -3735 3775 -3705
rect 3775 -3735 3805 -3705
rect 3805 -3735 3810 -3705
rect 3770 -3740 3810 -3735
rect 3770 -3770 3810 -3765
rect 3770 -3800 3775 -3770
rect 3775 -3800 3805 -3770
rect 3805 -3800 3810 -3770
rect 3770 -3805 3810 -3800
rect 3770 -3840 3810 -3835
rect 3770 -3870 3775 -3840
rect 3775 -3870 3805 -3840
rect 3805 -3870 3810 -3840
rect 3770 -3875 3810 -3870
rect 3770 -3910 3810 -3905
rect 3770 -3940 3775 -3910
rect 3775 -3940 3805 -3910
rect 3805 -3940 3810 -3910
rect 3770 -3945 3810 -3940
rect 3770 -3980 3810 -3975
rect 3770 -4010 3775 -3980
rect 3775 -4010 3805 -3980
rect 3805 -4010 3810 -3980
rect 3770 -4015 3810 -4010
rect 3770 -4045 3810 -4040
rect 3770 -4075 3775 -4045
rect 3775 -4075 3805 -4045
rect 3805 -4075 3810 -4045
rect 3770 -4080 3810 -4075
rect 3770 -4105 3810 -4100
rect 3770 -4135 3775 -4105
rect 3775 -4135 3805 -4105
rect 3805 -4135 3810 -4105
rect 3770 -4140 3810 -4135
rect 3770 -4170 3810 -4165
rect 3770 -4200 3775 -4170
rect 3775 -4200 3805 -4170
rect 3805 -4200 3810 -4170
rect 3770 -4205 3810 -4200
rect 3770 -4240 3810 -4235
rect 3770 -4270 3775 -4240
rect 3775 -4270 3805 -4240
rect 3805 -4270 3810 -4240
rect 3770 -4275 3810 -4270
rect 3770 -4310 3810 -4305
rect 3770 -4340 3775 -4310
rect 3775 -4340 3805 -4310
rect 3805 -4340 3810 -4310
rect 3770 -4345 3810 -4340
rect 3770 -4380 3810 -4375
rect 3770 -4410 3775 -4380
rect 3775 -4410 3805 -4380
rect 3805 -4410 3810 -4380
rect 3770 -4415 3810 -4410
rect 3770 -4445 3810 -4440
rect 3770 -4475 3775 -4445
rect 3775 -4475 3805 -4445
rect 3805 -4475 3810 -4445
rect 3770 -4480 3810 -4475
rect 4120 -1305 4160 -1300
rect 4120 -1335 4125 -1305
rect 4125 -1335 4155 -1305
rect 4155 -1335 4160 -1305
rect 4120 -1340 4160 -1335
rect 4120 -1370 4160 -1365
rect 4120 -1400 4125 -1370
rect 4125 -1400 4155 -1370
rect 4155 -1400 4160 -1370
rect 4120 -1405 4160 -1400
rect 4120 -1440 4160 -1435
rect 4120 -1470 4125 -1440
rect 4125 -1470 4155 -1440
rect 4155 -1470 4160 -1440
rect 4120 -1475 4160 -1470
rect 4120 -1510 4160 -1505
rect 4120 -1540 4125 -1510
rect 4125 -1540 4155 -1510
rect 4155 -1540 4160 -1510
rect 4120 -1545 4160 -1540
rect 4120 -1580 4160 -1575
rect 4120 -1610 4125 -1580
rect 4125 -1610 4155 -1580
rect 4155 -1610 4160 -1580
rect 4120 -1615 4160 -1610
rect 4120 -1645 4160 -1640
rect 4120 -1675 4125 -1645
rect 4125 -1675 4155 -1645
rect 4155 -1675 4160 -1645
rect 4120 -1680 4160 -1675
rect 4120 -1705 4160 -1700
rect 4120 -1735 4125 -1705
rect 4125 -1735 4155 -1705
rect 4155 -1735 4160 -1705
rect 4120 -1740 4160 -1735
rect 4120 -1770 4160 -1765
rect 4120 -1800 4125 -1770
rect 4125 -1800 4155 -1770
rect 4155 -1800 4160 -1770
rect 4120 -1805 4160 -1800
rect 4120 -1840 4160 -1835
rect 4120 -1870 4125 -1840
rect 4125 -1870 4155 -1840
rect 4155 -1870 4160 -1840
rect 4120 -1875 4160 -1870
rect 4120 -1910 4160 -1905
rect 4120 -1940 4125 -1910
rect 4125 -1940 4155 -1910
rect 4155 -1940 4160 -1910
rect 4120 -1945 4160 -1940
rect 4120 -1980 4160 -1975
rect 4120 -2010 4125 -1980
rect 4125 -2010 4155 -1980
rect 4155 -2010 4160 -1980
rect 4120 -2015 4160 -2010
rect 4120 -2045 4160 -2040
rect 4120 -2075 4125 -2045
rect 4125 -2075 4155 -2045
rect 4155 -2075 4160 -2045
rect 4120 -2080 4160 -2075
rect 4120 -2105 4160 -2100
rect 4120 -2135 4125 -2105
rect 4125 -2135 4155 -2105
rect 4155 -2135 4160 -2105
rect 4120 -2140 4160 -2135
rect 4120 -2170 4160 -2165
rect 4120 -2200 4125 -2170
rect 4125 -2200 4155 -2170
rect 4155 -2200 4160 -2170
rect 4120 -2205 4160 -2200
rect 4120 -2240 4160 -2235
rect 4120 -2270 4125 -2240
rect 4125 -2270 4155 -2240
rect 4155 -2270 4160 -2240
rect 4120 -2275 4160 -2270
rect 4120 -2310 4160 -2305
rect 4120 -2340 4125 -2310
rect 4125 -2340 4155 -2310
rect 4155 -2340 4160 -2310
rect 4120 -2345 4160 -2340
rect 4120 -2380 4160 -2375
rect 4120 -2410 4125 -2380
rect 4125 -2410 4155 -2380
rect 4155 -2410 4160 -2380
rect 4120 -2415 4160 -2410
rect 4120 -2445 4160 -2440
rect 4120 -2475 4125 -2445
rect 4125 -2475 4155 -2445
rect 4155 -2475 4160 -2445
rect 4120 -2480 4160 -2475
rect 4120 -2505 4160 -2500
rect 4120 -2535 4125 -2505
rect 4125 -2535 4155 -2505
rect 4155 -2535 4160 -2505
rect 4120 -2540 4160 -2535
rect 4120 -2570 4160 -2565
rect 4120 -2600 4125 -2570
rect 4125 -2600 4155 -2570
rect 4155 -2600 4160 -2570
rect 4120 -2605 4160 -2600
rect 4120 -2640 4160 -2635
rect 4120 -2670 4125 -2640
rect 4125 -2670 4155 -2640
rect 4155 -2670 4160 -2640
rect 4120 -2675 4160 -2670
rect 4120 -2710 4160 -2705
rect 4120 -2740 4125 -2710
rect 4125 -2740 4155 -2710
rect 4155 -2740 4160 -2710
rect 4120 -2745 4160 -2740
rect 4120 -2780 4160 -2775
rect 4120 -2810 4125 -2780
rect 4125 -2810 4155 -2780
rect 4155 -2810 4160 -2780
rect 4120 -2815 4160 -2810
rect 4120 -2845 4160 -2840
rect 4120 -2875 4125 -2845
rect 4125 -2875 4155 -2845
rect 4155 -2875 4160 -2845
rect 4120 -2880 4160 -2875
rect 4120 -2905 4160 -2900
rect 4120 -2935 4125 -2905
rect 4125 -2935 4155 -2905
rect 4155 -2935 4160 -2905
rect 4120 -2940 4160 -2935
rect 4120 -2970 4160 -2965
rect 4120 -3000 4125 -2970
rect 4125 -3000 4155 -2970
rect 4155 -3000 4160 -2970
rect 4120 -3005 4160 -3000
rect 4120 -3040 4160 -3035
rect 4120 -3070 4125 -3040
rect 4125 -3070 4155 -3040
rect 4155 -3070 4160 -3040
rect 4120 -3075 4160 -3070
rect 4120 -3110 4160 -3105
rect 4120 -3140 4125 -3110
rect 4125 -3140 4155 -3110
rect 4155 -3140 4160 -3110
rect 4120 -3145 4160 -3140
rect 4120 -3180 4160 -3175
rect 4120 -3210 4125 -3180
rect 4125 -3210 4155 -3180
rect 4155 -3210 4160 -3180
rect 4120 -3215 4160 -3210
rect 4120 -3245 4160 -3240
rect 4120 -3275 4125 -3245
rect 4125 -3275 4155 -3245
rect 4155 -3275 4160 -3245
rect 4120 -3280 4160 -3275
rect 4120 -3305 4160 -3300
rect 4120 -3335 4125 -3305
rect 4125 -3335 4155 -3305
rect 4155 -3335 4160 -3305
rect 4120 -3340 4160 -3335
rect 4120 -3370 4160 -3365
rect 4120 -3400 4125 -3370
rect 4125 -3400 4155 -3370
rect 4155 -3400 4160 -3370
rect 4120 -3405 4160 -3400
rect 4120 -3440 4160 -3435
rect 4120 -3470 4125 -3440
rect 4125 -3470 4155 -3440
rect 4155 -3470 4160 -3440
rect 4120 -3475 4160 -3470
rect 4120 -3510 4160 -3505
rect 4120 -3540 4125 -3510
rect 4125 -3540 4155 -3510
rect 4155 -3540 4160 -3510
rect 4120 -3545 4160 -3540
rect 4120 -3580 4160 -3575
rect 4120 -3610 4125 -3580
rect 4125 -3610 4155 -3580
rect 4155 -3610 4160 -3580
rect 4120 -3615 4160 -3610
rect 4120 -3645 4160 -3640
rect 4120 -3675 4125 -3645
rect 4125 -3675 4155 -3645
rect 4155 -3675 4160 -3645
rect 4120 -3680 4160 -3675
rect 4120 -3705 4160 -3700
rect 4120 -3735 4125 -3705
rect 4125 -3735 4155 -3705
rect 4155 -3735 4160 -3705
rect 4120 -3740 4160 -3735
rect 4120 -3770 4160 -3765
rect 4120 -3800 4125 -3770
rect 4125 -3800 4155 -3770
rect 4155 -3800 4160 -3770
rect 4120 -3805 4160 -3800
rect 4120 -3840 4160 -3835
rect 4120 -3870 4125 -3840
rect 4125 -3870 4155 -3840
rect 4155 -3870 4160 -3840
rect 4120 -3875 4160 -3870
rect 4120 -3910 4160 -3905
rect 4120 -3940 4125 -3910
rect 4125 -3940 4155 -3910
rect 4155 -3940 4160 -3910
rect 4120 -3945 4160 -3940
rect 4120 -3980 4160 -3975
rect 4120 -4010 4125 -3980
rect 4125 -4010 4155 -3980
rect 4155 -4010 4160 -3980
rect 4120 -4015 4160 -4010
rect 4120 -4045 4160 -4040
rect 4120 -4075 4125 -4045
rect 4125 -4075 4155 -4045
rect 4155 -4075 4160 -4045
rect 4120 -4080 4160 -4075
rect 4120 -4105 4160 -4100
rect 4120 -4135 4125 -4105
rect 4125 -4135 4155 -4105
rect 4155 -4135 4160 -4105
rect 4120 -4140 4160 -4135
rect 4120 -4170 4160 -4165
rect 4120 -4200 4125 -4170
rect 4125 -4200 4155 -4170
rect 4155 -4200 4160 -4170
rect 4120 -4205 4160 -4200
rect 4120 -4240 4160 -4235
rect 4120 -4270 4125 -4240
rect 4125 -4270 4155 -4240
rect 4155 -4270 4160 -4240
rect 4120 -4275 4160 -4270
rect 4120 -4310 4160 -4305
rect 4120 -4340 4125 -4310
rect 4125 -4340 4155 -4310
rect 4155 -4340 4160 -4310
rect 4120 -4345 4160 -4340
rect 4120 -4380 4160 -4375
rect 4120 -4410 4125 -4380
rect 4125 -4410 4155 -4380
rect 4155 -4410 4160 -4380
rect 4120 -4415 4160 -4410
rect 4120 -4445 4160 -4440
rect 4120 -4475 4125 -4445
rect 4125 -4475 4155 -4445
rect 4155 -4475 4160 -4445
rect 4120 -4480 4160 -4475
rect 4470 -1305 4510 -1300
rect 4470 -1335 4475 -1305
rect 4475 -1335 4505 -1305
rect 4505 -1335 4510 -1305
rect 4470 -1340 4510 -1335
rect 4470 -1370 4510 -1365
rect 4470 -1400 4475 -1370
rect 4475 -1400 4505 -1370
rect 4505 -1400 4510 -1370
rect 4470 -1405 4510 -1400
rect 4470 -1440 4510 -1435
rect 4470 -1470 4475 -1440
rect 4475 -1470 4505 -1440
rect 4505 -1470 4510 -1440
rect 4470 -1475 4510 -1470
rect 4470 -1510 4510 -1505
rect 4470 -1540 4475 -1510
rect 4475 -1540 4505 -1510
rect 4505 -1540 4510 -1510
rect 4470 -1545 4510 -1540
rect 4470 -1580 4510 -1575
rect 4470 -1610 4475 -1580
rect 4475 -1610 4505 -1580
rect 4505 -1610 4510 -1580
rect 4470 -1615 4510 -1610
rect 4470 -1645 4510 -1640
rect 4470 -1675 4475 -1645
rect 4475 -1675 4505 -1645
rect 4505 -1675 4510 -1645
rect 4470 -1680 4510 -1675
rect 4470 -1705 4510 -1700
rect 4470 -1735 4475 -1705
rect 4475 -1735 4505 -1705
rect 4505 -1735 4510 -1705
rect 4470 -1740 4510 -1735
rect 4470 -1770 4510 -1765
rect 4470 -1800 4475 -1770
rect 4475 -1800 4505 -1770
rect 4505 -1800 4510 -1770
rect 4470 -1805 4510 -1800
rect 4470 -1840 4510 -1835
rect 4470 -1870 4475 -1840
rect 4475 -1870 4505 -1840
rect 4505 -1870 4510 -1840
rect 4470 -1875 4510 -1870
rect 4470 -1910 4510 -1905
rect 4470 -1940 4475 -1910
rect 4475 -1940 4505 -1910
rect 4505 -1940 4510 -1910
rect 4470 -1945 4510 -1940
rect 4470 -1980 4510 -1975
rect 4470 -2010 4475 -1980
rect 4475 -2010 4505 -1980
rect 4505 -2010 4510 -1980
rect 4470 -2015 4510 -2010
rect 4470 -2045 4510 -2040
rect 4470 -2075 4475 -2045
rect 4475 -2075 4505 -2045
rect 4505 -2075 4510 -2045
rect 4470 -2080 4510 -2075
rect 4470 -2105 4510 -2100
rect 4470 -2135 4475 -2105
rect 4475 -2135 4505 -2105
rect 4505 -2135 4510 -2105
rect 4470 -2140 4510 -2135
rect 4470 -2170 4510 -2165
rect 4470 -2200 4475 -2170
rect 4475 -2200 4505 -2170
rect 4505 -2200 4510 -2170
rect 4470 -2205 4510 -2200
rect 4470 -2240 4510 -2235
rect 4470 -2270 4475 -2240
rect 4475 -2270 4505 -2240
rect 4505 -2270 4510 -2240
rect 4470 -2275 4510 -2270
rect 4470 -2310 4510 -2305
rect 4470 -2340 4475 -2310
rect 4475 -2340 4505 -2310
rect 4505 -2340 4510 -2310
rect 4470 -2345 4510 -2340
rect 4470 -2380 4510 -2375
rect 4470 -2410 4475 -2380
rect 4475 -2410 4505 -2380
rect 4505 -2410 4510 -2380
rect 4470 -2415 4510 -2410
rect 4470 -2445 4510 -2440
rect 4470 -2475 4475 -2445
rect 4475 -2475 4505 -2445
rect 4505 -2475 4510 -2445
rect 4470 -2480 4510 -2475
rect 4470 -2505 4510 -2500
rect 4470 -2535 4475 -2505
rect 4475 -2535 4505 -2505
rect 4505 -2535 4510 -2505
rect 4470 -2540 4510 -2535
rect 4470 -2570 4510 -2565
rect 4470 -2600 4475 -2570
rect 4475 -2600 4505 -2570
rect 4505 -2600 4510 -2570
rect 4470 -2605 4510 -2600
rect 4470 -2640 4510 -2635
rect 4470 -2670 4475 -2640
rect 4475 -2670 4505 -2640
rect 4505 -2670 4510 -2640
rect 4470 -2675 4510 -2670
rect 4470 -2710 4510 -2705
rect 4470 -2740 4475 -2710
rect 4475 -2740 4505 -2710
rect 4505 -2740 4510 -2710
rect 4470 -2745 4510 -2740
rect 4470 -2780 4510 -2775
rect 4470 -2810 4475 -2780
rect 4475 -2810 4505 -2780
rect 4505 -2810 4510 -2780
rect 4470 -2815 4510 -2810
rect 4470 -2845 4510 -2840
rect 4470 -2875 4475 -2845
rect 4475 -2875 4505 -2845
rect 4505 -2875 4510 -2845
rect 4470 -2880 4510 -2875
rect 4470 -2905 4510 -2900
rect 4470 -2935 4475 -2905
rect 4475 -2935 4505 -2905
rect 4505 -2935 4510 -2905
rect 4470 -2940 4510 -2935
rect 4470 -2970 4510 -2965
rect 4470 -3000 4475 -2970
rect 4475 -3000 4505 -2970
rect 4505 -3000 4510 -2970
rect 4470 -3005 4510 -3000
rect 4470 -3040 4510 -3035
rect 4470 -3070 4475 -3040
rect 4475 -3070 4505 -3040
rect 4505 -3070 4510 -3040
rect 4470 -3075 4510 -3070
rect 4470 -3110 4510 -3105
rect 4470 -3140 4475 -3110
rect 4475 -3140 4505 -3110
rect 4505 -3140 4510 -3110
rect 4470 -3145 4510 -3140
rect 4470 -3180 4510 -3175
rect 4470 -3210 4475 -3180
rect 4475 -3210 4505 -3180
rect 4505 -3210 4510 -3180
rect 4470 -3215 4510 -3210
rect 4470 -3245 4510 -3240
rect 4470 -3275 4475 -3245
rect 4475 -3275 4505 -3245
rect 4505 -3275 4510 -3245
rect 4470 -3280 4510 -3275
rect 4470 -3305 4510 -3300
rect 4470 -3335 4475 -3305
rect 4475 -3335 4505 -3305
rect 4505 -3335 4510 -3305
rect 4470 -3340 4510 -3335
rect 4470 -3370 4510 -3365
rect 4470 -3400 4475 -3370
rect 4475 -3400 4505 -3370
rect 4505 -3400 4510 -3370
rect 4470 -3405 4510 -3400
rect 4470 -3440 4510 -3435
rect 4470 -3470 4475 -3440
rect 4475 -3470 4505 -3440
rect 4505 -3470 4510 -3440
rect 4470 -3475 4510 -3470
rect 4470 -3510 4510 -3505
rect 4470 -3540 4475 -3510
rect 4475 -3540 4505 -3510
rect 4505 -3540 4510 -3510
rect 4470 -3545 4510 -3540
rect 4470 -3580 4510 -3575
rect 4470 -3610 4475 -3580
rect 4475 -3610 4505 -3580
rect 4505 -3610 4510 -3580
rect 4470 -3615 4510 -3610
rect 4470 -3645 4510 -3640
rect 4470 -3675 4475 -3645
rect 4475 -3675 4505 -3645
rect 4505 -3675 4510 -3645
rect 4470 -3680 4510 -3675
rect 4470 -3705 4510 -3700
rect 4470 -3735 4475 -3705
rect 4475 -3735 4505 -3705
rect 4505 -3735 4510 -3705
rect 4470 -3740 4510 -3735
rect 4470 -3770 4510 -3765
rect 4470 -3800 4475 -3770
rect 4475 -3800 4505 -3770
rect 4505 -3800 4510 -3770
rect 4470 -3805 4510 -3800
rect 4470 -3840 4510 -3835
rect 4470 -3870 4475 -3840
rect 4475 -3870 4505 -3840
rect 4505 -3870 4510 -3840
rect 4470 -3875 4510 -3870
rect 4470 -3910 4510 -3905
rect 4470 -3940 4475 -3910
rect 4475 -3940 4505 -3910
rect 4505 -3940 4510 -3910
rect 4470 -3945 4510 -3940
rect 4470 -3980 4510 -3975
rect 4470 -4010 4475 -3980
rect 4475 -4010 4505 -3980
rect 4505 -4010 4510 -3980
rect 4470 -4015 4510 -4010
rect 4470 -4045 4510 -4040
rect 4470 -4075 4475 -4045
rect 4475 -4075 4505 -4045
rect 4505 -4075 4510 -4045
rect 4470 -4080 4510 -4075
rect 4470 -4105 4510 -4100
rect 4470 -4135 4475 -4105
rect 4475 -4135 4505 -4105
rect 4505 -4135 4510 -4105
rect 4470 -4140 4510 -4135
rect 4470 -4170 4510 -4165
rect 4470 -4200 4475 -4170
rect 4475 -4200 4505 -4170
rect 4505 -4200 4510 -4170
rect 4470 -4205 4510 -4200
rect 4470 -4240 4510 -4235
rect 4470 -4270 4475 -4240
rect 4475 -4270 4505 -4240
rect 4505 -4270 4510 -4240
rect 4470 -4275 4510 -4270
rect 4470 -4310 4510 -4305
rect 4470 -4340 4475 -4310
rect 4475 -4340 4505 -4310
rect 4505 -4340 4510 -4310
rect 4470 -4345 4510 -4340
rect 4470 -4380 4510 -4375
rect 4470 -4410 4475 -4380
rect 4475 -4410 4505 -4380
rect 4505 -4410 4510 -4380
rect 4470 -4415 4510 -4410
rect 4470 -4445 4510 -4440
rect 4470 -4475 4475 -4445
rect 4475 -4475 4505 -4445
rect 4505 -4475 4510 -4445
rect 4470 -4480 4510 -4475
rect 4820 -1305 4860 -1300
rect 4820 -1335 4825 -1305
rect 4825 -1335 4855 -1305
rect 4855 -1335 4860 -1305
rect 4820 -1340 4860 -1335
rect 4820 -1370 4860 -1365
rect 4820 -1400 4825 -1370
rect 4825 -1400 4855 -1370
rect 4855 -1400 4860 -1370
rect 4820 -1405 4860 -1400
rect 4820 -1440 4860 -1435
rect 4820 -1470 4825 -1440
rect 4825 -1470 4855 -1440
rect 4855 -1470 4860 -1440
rect 4820 -1475 4860 -1470
rect 4820 -1510 4860 -1505
rect 4820 -1540 4825 -1510
rect 4825 -1540 4855 -1510
rect 4855 -1540 4860 -1510
rect 4820 -1545 4860 -1540
rect 4820 -1580 4860 -1575
rect 4820 -1610 4825 -1580
rect 4825 -1610 4855 -1580
rect 4855 -1610 4860 -1580
rect 4820 -1615 4860 -1610
rect 4820 -1645 4860 -1640
rect 4820 -1675 4825 -1645
rect 4825 -1675 4855 -1645
rect 4855 -1675 4860 -1645
rect 4820 -1680 4860 -1675
rect 4820 -1705 4860 -1700
rect 4820 -1735 4825 -1705
rect 4825 -1735 4855 -1705
rect 4855 -1735 4860 -1705
rect 4820 -1740 4860 -1735
rect 4820 -1770 4860 -1765
rect 4820 -1800 4825 -1770
rect 4825 -1800 4855 -1770
rect 4855 -1800 4860 -1770
rect 4820 -1805 4860 -1800
rect 4820 -1840 4860 -1835
rect 4820 -1870 4825 -1840
rect 4825 -1870 4855 -1840
rect 4855 -1870 4860 -1840
rect 4820 -1875 4860 -1870
rect 4820 -1910 4860 -1905
rect 4820 -1940 4825 -1910
rect 4825 -1940 4855 -1910
rect 4855 -1940 4860 -1910
rect 4820 -1945 4860 -1940
rect 4820 -1980 4860 -1975
rect 4820 -2010 4825 -1980
rect 4825 -2010 4855 -1980
rect 4855 -2010 4860 -1980
rect 4820 -2015 4860 -2010
rect 4820 -2045 4860 -2040
rect 4820 -2075 4825 -2045
rect 4825 -2075 4855 -2045
rect 4855 -2075 4860 -2045
rect 4820 -2080 4860 -2075
rect 4820 -2105 4860 -2100
rect 4820 -2135 4825 -2105
rect 4825 -2135 4855 -2105
rect 4855 -2135 4860 -2105
rect 4820 -2140 4860 -2135
rect 4820 -2170 4860 -2165
rect 4820 -2200 4825 -2170
rect 4825 -2200 4855 -2170
rect 4855 -2200 4860 -2170
rect 4820 -2205 4860 -2200
rect 4820 -2240 4860 -2235
rect 4820 -2270 4825 -2240
rect 4825 -2270 4855 -2240
rect 4855 -2270 4860 -2240
rect 4820 -2275 4860 -2270
rect 4820 -2310 4860 -2305
rect 4820 -2340 4825 -2310
rect 4825 -2340 4855 -2310
rect 4855 -2340 4860 -2310
rect 4820 -2345 4860 -2340
rect 4820 -2380 4860 -2375
rect 4820 -2410 4825 -2380
rect 4825 -2410 4855 -2380
rect 4855 -2410 4860 -2380
rect 4820 -2415 4860 -2410
rect 4820 -2445 4860 -2440
rect 4820 -2475 4825 -2445
rect 4825 -2475 4855 -2445
rect 4855 -2475 4860 -2445
rect 4820 -2480 4860 -2475
rect 4820 -2505 4860 -2500
rect 4820 -2535 4825 -2505
rect 4825 -2535 4855 -2505
rect 4855 -2535 4860 -2505
rect 4820 -2540 4860 -2535
rect 4820 -2570 4860 -2565
rect 4820 -2600 4825 -2570
rect 4825 -2600 4855 -2570
rect 4855 -2600 4860 -2570
rect 4820 -2605 4860 -2600
rect 4820 -2640 4860 -2635
rect 4820 -2670 4825 -2640
rect 4825 -2670 4855 -2640
rect 4855 -2670 4860 -2640
rect 4820 -2675 4860 -2670
rect 4820 -2710 4860 -2705
rect 4820 -2740 4825 -2710
rect 4825 -2740 4855 -2710
rect 4855 -2740 4860 -2710
rect 4820 -2745 4860 -2740
rect 4820 -2780 4860 -2775
rect 4820 -2810 4825 -2780
rect 4825 -2810 4855 -2780
rect 4855 -2810 4860 -2780
rect 4820 -2815 4860 -2810
rect 4820 -2845 4860 -2840
rect 4820 -2875 4825 -2845
rect 4825 -2875 4855 -2845
rect 4855 -2875 4860 -2845
rect 4820 -2880 4860 -2875
rect 4820 -2905 4860 -2900
rect 4820 -2935 4825 -2905
rect 4825 -2935 4855 -2905
rect 4855 -2935 4860 -2905
rect 4820 -2940 4860 -2935
rect 4820 -2970 4860 -2965
rect 4820 -3000 4825 -2970
rect 4825 -3000 4855 -2970
rect 4855 -3000 4860 -2970
rect 4820 -3005 4860 -3000
rect 4820 -3040 4860 -3035
rect 4820 -3070 4825 -3040
rect 4825 -3070 4855 -3040
rect 4855 -3070 4860 -3040
rect 4820 -3075 4860 -3070
rect 4820 -3110 4860 -3105
rect 4820 -3140 4825 -3110
rect 4825 -3140 4855 -3110
rect 4855 -3140 4860 -3110
rect 4820 -3145 4860 -3140
rect 4820 -3180 4860 -3175
rect 4820 -3210 4825 -3180
rect 4825 -3210 4855 -3180
rect 4855 -3210 4860 -3180
rect 4820 -3215 4860 -3210
rect 4820 -3245 4860 -3240
rect 4820 -3275 4825 -3245
rect 4825 -3275 4855 -3245
rect 4855 -3275 4860 -3245
rect 4820 -3280 4860 -3275
rect 4820 -3305 4860 -3300
rect 4820 -3335 4825 -3305
rect 4825 -3335 4855 -3305
rect 4855 -3335 4860 -3305
rect 4820 -3340 4860 -3335
rect 4820 -3370 4860 -3365
rect 4820 -3400 4825 -3370
rect 4825 -3400 4855 -3370
rect 4855 -3400 4860 -3370
rect 4820 -3405 4860 -3400
rect 4820 -3440 4860 -3435
rect 4820 -3470 4825 -3440
rect 4825 -3470 4855 -3440
rect 4855 -3470 4860 -3440
rect 4820 -3475 4860 -3470
rect 4820 -3510 4860 -3505
rect 4820 -3540 4825 -3510
rect 4825 -3540 4855 -3510
rect 4855 -3540 4860 -3510
rect 4820 -3545 4860 -3540
rect 4820 -3580 4860 -3575
rect 4820 -3610 4825 -3580
rect 4825 -3610 4855 -3580
rect 4855 -3610 4860 -3580
rect 4820 -3615 4860 -3610
rect 4820 -3645 4860 -3640
rect 4820 -3675 4825 -3645
rect 4825 -3675 4855 -3645
rect 4855 -3675 4860 -3645
rect 4820 -3680 4860 -3675
rect 4820 -3705 4860 -3700
rect 4820 -3735 4825 -3705
rect 4825 -3735 4855 -3705
rect 4855 -3735 4860 -3705
rect 4820 -3740 4860 -3735
rect 4820 -3770 4860 -3765
rect 4820 -3800 4825 -3770
rect 4825 -3800 4855 -3770
rect 4855 -3800 4860 -3770
rect 4820 -3805 4860 -3800
rect 4820 -3840 4860 -3835
rect 4820 -3870 4825 -3840
rect 4825 -3870 4855 -3840
rect 4855 -3870 4860 -3840
rect 4820 -3875 4860 -3870
rect 4820 -3910 4860 -3905
rect 4820 -3940 4825 -3910
rect 4825 -3940 4855 -3910
rect 4855 -3940 4860 -3910
rect 4820 -3945 4860 -3940
rect 4820 -3980 4860 -3975
rect 4820 -4010 4825 -3980
rect 4825 -4010 4855 -3980
rect 4855 -4010 4860 -3980
rect 4820 -4015 4860 -4010
rect 4820 -4045 4860 -4040
rect 4820 -4075 4825 -4045
rect 4825 -4075 4855 -4045
rect 4855 -4075 4860 -4045
rect 4820 -4080 4860 -4075
rect 4820 -4105 4860 -4100
rect 4820 -4135 4825 -4105
rect 4825 -4135 4855 -4105
rect 4855 -4135 4860 -4105
rect 4820 -4140 4860 -4135
rect 4820 -4170 4860 -4165
rect 4820 -4200 4825 -4170
rect 4825 -4200 4855 -4170
rect 4855 -4200 4860 -4170
rect 4820 -4205 4860 -4200
rect 4820 -4240 4860 -4235
rect 4820 -4270 4825 -4240
rect 4825 -4270 4855 -4240
rect 4855 -4270 4860 -4240
rect 4820 -4275 4860 -4270
rect 4820 -4310 4860 -4305
rect 4820 -4340 4825 -4310
rect 4825 -4340 4855 -4310
rect 4855 -4340 4860 -4310
rect 4820 -4345 4860 -4340
rect 4820 -4380 4860 -4375
rect 4820 -4410 4825 -4380
rect 4825 -4410 4855 -4380
rect 4855 -4410 4860 -4380
rect 4820 -4415 4860 -4410
rect 4820 -4445 4860 -4440
rect 4820 -4475 4825 -4445
rect 4825 -4475 4855 -4445
rect 4855 -4475 4860 -4445
rect 4820 -4480 4860 -4475
rect 5170 -1305 5210 -1300
rect 5170 -1335 5175 -1305
rect 5175 -1335 5205 -1305
rect 5205 -1335 5210 -1305
rect 5170 -1340 5210 -1335
rect 5170 -1370 5210 -1365
rect 5170 -1400 5175 -1370
rect 5175 -1400 5205 -1370
rect 5205 -1400 5210 -1370
rect 5170 -1405 5210 -1400
rect 5170 -1440 5210 -1435
rect 5170 -1470 5175 -1440
rect 5175 -1470 5205 -1440
rect 5205 -1470 5210 -1440
rect 5170 -1475 5210 -1470
rect 5170 -1510 5210 -1505
rect 5170 -1540 5175 -1510
rect 5175 -1540 5205 -1510
rect 5205 -1540 5210 -1510
rect 5170 -1545 5210 -1540
rect 5170 -1580 5210 -1575
rect 5170 -1610 5175 -1580
rect 5175 -1610 5205 -1580
rect 5205 -1610 5210 -1580
rect 5170 -1615 5210 -1610
rect 5170 -1645 5210 -1640
rect 5170 -1675 5175 -1645
rect 5175 -1675 5205 -1645
rect 5205 -1675 5210 -1645
rect 5170 -1680 5210 -1675
rect 5170 -1705 5210 -1700
rect 5170 -1735 5175 -1705
rect 5175 -1735 5205 -1705
rect 5205 -1735 5210 -1705
rect 5170 -1740 5210 -1735
rect 5170 -1770 5210 -1765
rect 5170 -1800 5175 -1770
rect 5175 -1800 5205 -1770
rect 5205 -1800 5210 -1770
rect 5170 -1805 5210 -1800
rect 5170 -1840 5210 -1835
rect 5170 -1870 5175 -1840
rect 5175 -1870 5205 -1840
rect 5205 -1870 5210 -1840
rect 5170 -1875 5210 -1870
rect 5170 -1910 5210 -1905
rect 5170 -1940 5175 -1910
rect 5175 -1940 5205 -1910
rect 5205 -1940 5210 -1910
rect 5170 -1945 5210 -1940
rect 5170 -1980 5210 -1975
rect 5170 -2010 5175 -1980
rect 5175 -2010 5205 -1980
rect 5205 -2010 5210 -1980
rect 5170 -2015 5210 -2010
rect 5170 -2045 5210 -2040
rect 5170 -2075 5175 -2045
rect 5175 -2075 5205 -2045
rect 5205 -2075 5210 -2045
rect 5170 -2080 5210 -2075
rect 5170 -2105 5210 -2100
rect 5170 -2135 5175 -2105
rect 5175 -2135 5205 -2105
rect 5205 -2135 5210 -2105
rect 5170 -2140 5210 -2135
rect 5170 -2170 5210 -2165
rect 5170 -2200 5175 -2170
rect 5175 -2200 5205 -2170
rect 5205 -2200 5210 -2170
rect 5170 -2205 5210 -2200
rect 5170 -2240 5210 -2235
rect 5170 -2270 5175 -2240
rect 5175 -2270 5205 -2240
rect 5205 -2270 5210 -2240
rect 5170 -2275 5210 -2270
rect 5170 -2310 5210 -2305
rect 5170 -2340 5175 -2310
rect 5175 -2340 5205 -2310
rect 5205 -2340 5210 -2310
rect 5170 -2345 5210 -2340
rect 5170 -2380 5210 -2375
rect 5170 -2410 5175 -2380
rect 5175 -2410 5205 -2380
rect 5205 -2410 5210 -2380
rect 5170 -2415 5210 -2410
rect 5170 -2445 5210 -2440
rect 5170 -2475 5175 -2445
rect 5175 -2475 5205 -2445
rect 5205 -2475 5210 -2445
rect 5170 -2480 5210 -2475
rect 5170 -2505 5210 -2500
rect 5170 -2535 5175 -2505
rect 5175 -2535 5205 -2505
rect 5205 -2535 5210 -2505
rect 5170 -2540 5210 -2535
rect 5170 -2570 5210 -2565
rect 5170 -2600 5175 -2570
rect 5175 -2600 5205 -2570
rect 5205 -2600 5210 -2570
rect 5170 -2605 5210 -2600
rect 5170 -2640 5210 -2635
rect 5170 -2670 5175 -2640
rect 5175 -2670 5205 -2640
rect 5205 -2670 5210 -2640
rect 5170 -2675 5210 -2670
rect 5170 -2710 5210 -2705
rect 5170 -2740 5175 -2710
rect 5175 -2740 5205 -2710
rect 5205 -2740 5210 -2710
rect 5170 -2745 5210 -2740
rect 5170 -2780 5210 -2775
rect 5170 -2810 5175 -2780
rect 5175 -2810 5205 -2780
rect 5205 -2810 5210 -2780
rect 5170 -2815 5210 -2810
rect 5170 -2845 5210 -2840
rect 5170 -2875 5175 -2845
rect 5175 -2875 5205 -2845
rect 5205 -2875 5210 -2845
rect 5170 -2880 5210 -2875
rect 5170 -2905 5210 -2900
rect 5170 -2935 5175 -2905
rect 5175 -2935 5205 -2905
rect 5205 -2935 5210 -2905
rect 5170 -2940 5210 -2935
rect 5170 -2970 5210 -2965
rect 5170 -3000 5175 -2970
rect 5175 -3000 5205 -2970
rect 5205 -3000 5210 -2970
rect 5170 -3005 5210 -3000
rect 5170 -3040 5210 -3035
rect 5170 -3070 5175 -3040
rect 5175 -3070 5205 -3040
rect 5205 -3070 5210 -3040
rect 5170 -3075 5210 -3070
rect 5170 -3110 5210 -3105
rect 5170 -3140 5175 -3110
rect 5175 -3140 5205 -3110
rect 5205 -3140 5210 -3110
rect 5170 -3145 5210 -3140
rect 5170 -3180 5210 -3175
rect 5170 -3210 5175 -3180
rect 5175 -3210 5205 -3180
rect 5205 -3210 5210 -3180
rect 5170 -3215 5210 -3210
rect 5170 -3245 5210 -3240
rect 5170 -3275 5175 -3245
rect 5175 -3275 5205 -3245
rect 5205 -3275 5210 -3245
rect 5170 -3280 5210 -3275
rect 5170 -3305 5210 -3300
rect 5170 -3335 5175 -3305
rect 5175 -3335 5205 -3305
rect 5205 -3335 5210 -3305
rect 5170 -3340 5210 -3335
rect 5170 -3370 5210 -3365
rect 5170 -3400 5175 -3370
rect 5175 -3400 5205 -3370
rect 5205 -3400 5210 -3370
rect 5170 -3405 5210 -3400
rect 5170 -3440 5210 -3435
rect 5170 -3470 5175 -3440
rect 5175 -3470 5205 -3440
rect 5205 -3470 5210 -3440
rect 5170 -3475 5210 -3470
rect 5170 -3510 5210 -3505
rect 5170 -3540 5175 -3510
rect 5175 -3540 5205 -3510
rect 5205 -3540 5210 -3510
rect 5170 -3545 5210 -3540
rect 5170 -3580 5210 -3575
rect 5170 -3610 5175 -3580
rect 5175 -3610 5205 -3580
rect 5205 -3610 5210 -3580
rect 5170 -3615 5210 -3610
rect 5170 -3645 5210 -3640
rect 5170 -3675 5175 -3645
rect 5175 -3675 5205 -3645
rect 5205 -3675 5210 -3645
rect 5170 -3680 5210 -3675
rect 5170 -3705 5210 -3700
rect 5170 -3735 5175 -3705
rect 5175 -3735 5205 -3705
rect 5205 -3735 5210 -3705
rect 5170 -3740 5210 -3735
rect 5170 -3770 5210 -3765
rect 5170 -3800 5175 -3770
rect 5175 -3800 5205 -3770
rect 5205 -3800 5210 -3770
rect 5170 -3805 5210 -3800
rect 5170 -3840 5210 -3835
rect 5170 -3870 5175 -3840
rect 5175 -3870 5205 -3840
rect 5205 -3870 5210 -3840
rect 5170 -3875 5210 -3870
rect 5170 -3910 5210 -3905
rect 5170 -3940 5175 -3910
rect 5175 -3940 5205 -3910
rect 5205 -3940 5210 -3910
rect 5170 -3945 5210 -3940
rect 5170 -3980 5210 -3975
rect 5170 -4010 5175 -3980
rect 5175 -4010 5205 -3980
rect 5205 -4010 5210 -3980
rect 5170 -4015 5210 -4010
rect 5170 -4045 5210 -4040
rect 5170 -4075 5175 -4045
rect 5175 -4075 5205 -4045
rect 5205 -4075 5210 -4045
rect 5170 -4080 5210 -4075
rect 5170 -4105 5210 -4100
rect 5170 -4135 5175 -4105
rect 5175 -4135 5205 -4105
rect 5205 -4135 5210 -4105
rect 5170 -4140 5210 -4135
rect 5170 -4170 5210 -4165
rect 5170 -4200 5175 -4170
rect 5175 -4200 5205 -4170
rect 5205 -4200 5210 -4170
rect 5170 -4205 5210 -4200
rect 5170 -4240 5210 -4235
rect 5170 -4270 5175 -4240
rect 5175 -4270 5205 -4240
rect 5205 -4270 5210 -4240
rect 5170 -4275 5210 -4270
rect 5170 -4310 5210 -4305
rect 5170 -4340 5175 -4310
rect 5175 -4340 5205 -4310
rect 5205 -4340 5210 -4310
rect 5170 -4345 5210 -4340
rect 5170 -4380 5210 -4375
rect 5170 -4410 5175 -4380
rect 5175 -4410 5205 -4380
rect 5205 -4410 5210 -4380
rect 5170 -4415 5210 -4410
rect 5170 -4445 5210 -4440
rect 5170 -4475 5175 -4445
rect 5175 -4475 5205 -4445
rect 5205 -4475 5210 -4445
rect 5170 -4480 5210 -4475
rect 5520 -1305 5560 -1300
rect 5520 -1335 5525 -1305
rect 5525 -1335 5555 -1305
rect 5555 -1335 5560 -1305
rect 5520 -1340 5560 -1335
rect 5520 -1370 5560 -1365
rect 5520 -1400 5525 -1370
rect 5525 -1400 5555 -1370
rect 5555 -1400 5560 -1370
rect 5520 -1405 5560 -1400
rect 5520 -1440 5560 -1435
rect 5520 -1470 5525 -1440
rect 5525 -1470 5555 -1440
rect 5555 -1470 5560 -1440
rect 5520 -1475 5560 -1470
rect 5520 -1510 5560 -1505
rect 5520 -1540 5525 -1510
rect 5525 -1540 5555 -1510
rect 5555 -1540 5560 -1510
rect 5520 -1545 5560 -1540
rect 5520 -1580 5560 -1575
rect 5520 -1610 5525 -1580
rect 5525 -1610 5555 -1580
rect 5555 -1610 5560 -1580
rect 5520 -1615 5560 -1610
rect 5520 -1645 5560 -1640
rect 5520 -1675 5525 -1645
rect 5525 -1675 5555 -1645
rect 5555 -1675 5560 -1645
rect 5520 -1680 5560 -1675
rect 5520 -1705 5560 -1700
rect 5520 -1735 5525 -1705
rect 5525 -1735 5555 -1705
rect 5555 -1735 5560 -1705
rect 5520 -1740 5560 -1735
rect 5520 -1770 5560 -1765
rect 5520 -1800 5525 -1770
rect 5525 -1800 5555 -1770
rect 5555 -1800 5560 -1770
rect 5520 -1805 5560 -1800
rect 5520 -1840 5560 -1835
rect 5520 -1870 5525 -1840
rect 5525 -1870 5555 -1840
rect 5555 -1870 5560 -1840
rect 5520 -1875 5560 -1870
rect 5520 -1910 5560 -1905
rect 5520 -1940 5525 -1910
rect 5525 -1940 5555 -1910
rect 5555 -1940 5560 -1910
rect 5520 -1945 5560 -1940
rect 5520 -1980 5560 -1975
rect 5520 -2010 5525 -1980
rect 5525 -2010 5555 -1980
rect 5555 -2010 5560 -1980
rect 5520 -2015 5560 -2010
rect 5520 -2045 5560 -2040
rect 5520 -2075 5525 -2045
rect 5525 -2075 5555 -2045
rect 5555 -2075 5560 -2045
rect 5520 -2080 5560 -2075
rect 5520 -2105 5560 -2100
rect 5520 -2135 5525 -2105
rect 5525 -2135 5555 -2105
rect 5555 -2135 5560 -2105
rect 5520 -2140 5560 -2135
rect 5520 -2170 5560 -2165
rect 5520 -2200 5525 -2170
rect 5525 -2200 5555 -2170
rect 5555 -2200 5560 -2170
rect 5520 -2205 5560 -2200
rect 5520 -2240 5560 -2235
rect 5520 -2270 5525 -2240
rect 5525 -2270 5555 -2240
rect 5555 -2270 5560 -2240
rect 5520 -2275 5560 -2270
rect 5520 -2310 5560 -2305
rect 5520 -2340 5525 -2310
rect 5525 -2340 5555 -2310
rect 5555 -2340 5560 -2310
rect 5520 -2345 5560 -2340
rect 5520 -2380 5560 -2375
rect 5520 -2410 5525 -2380
rect 5525 -2410 5555 -2380
rect 5555 -2410 5560 -2380
rect 5520 -2415 5560 -2410
rect 5520 -2445 5560 -2440
rect 5520 -2475 5525 -2445
rect 5525 -2475 5555 -2445
rect 5555 -2475 5560 -2445
rect 5520 -2480 5560 -2475
rect 5520 -2505 5560 -2500
rect 5520 -2535 5525 -2505
rect 5525 -2535 5555 -2505
rect 5555 -2535 5560 -2505
rect 5520 -2540 5560 -2535
rect 5520 -2570 5560 -2565
rect 5520 -2600 5525 -2570
rect 5525 -2600 5555 -2570
rect 5555 -2600 5560 -2570
rect 5520 -2605 5560 -2600
rect 5520 -2640 5560 -2635
rect 5520 -2670 5525 -2640
rect 5525 -2670 5555 -2640
rect 5555 -2670 5560 -2640
rect 5520 -2675 5560 -2670
rect 5520 -2710 5560 -2705
rect 5520 -2740 5525 -2710
rect 5525 -2740 5555 -2710
rect 5555 -2740 5560 -2710
rect 5520 -2745 5560 -2740
rect 5520 -2780 5560 -2775
rect 5520 -2810 5525 -2780
rect 5525 -2810 5555 -2780
rect 5555 -2810 5560 -2780
rect 5520 -2815 5560 -2810
rect 5520 -2845 5560 -2840
rect 5520 -2875 5525 -2845
rect 5525 -2875 5555 -2845
rect 5555 -2875 5560 -2845
rect 5520 -2880 5560 -2875
rect 5520 -2905 5560 -2900
rect 5520 -2935 5525 -2905
rect 5525 -2935 5555 -2905
rect 5555 -2935 5560 -2905
rect 5520 -2940 5560 -2935
rect 5520 -2970 5560 -2965
rect 5520 -3000 5525 -2970
rect 5525 -3000 5555 -2970
rect 5555 -3000 5560 -2970
rect 5520 -3005 5560 -3000
rect 5520 -3040 5560 -3035
rect 5520 -3070 5525 -3040
rect 5525 -3070 5555 -3040
rect 5555 -3070 5560 -3040
rect 5520 -3075 5560 -3070
rect 5520 -3110 5560 -3105
rect 5520 -3140 5525 -3110
rect 5525 -3140 5555 -3110
rect 5555 -3140 5560 -3110
rect 5520 -3145 5560 -3140
rect 5520 -3180 5560 -3175
rect 5520 -3210 5525 -3180
rect 5525 -3210 5555 -3180
rect 5555 -3210 5560 -3180
rect 5520 -3215 5560 -3210
rect 5520 -3245 5560 -3240
rect 5520 -3275 5525 -3245
rect 5525 -3275 5555 -3245
rect 5555 -3275 5560 -3245
rect 5520 -3280 5560 -3275
rect 5520 -3305 5560 -3300
rect 5520 -3335 5525 -3305
rect 5525 -3335 5555 -3305
rect 5555 -3335 5560 -3305
rect 5520 -3340 5560 -3335
rect 5520 -3370 5560 -3365
rect 5520 -3400 5525 -3370
rect 5525 -3400 5555 -3370
rect 5555 -3400 5560 -3370
rect 5520 -3405 5560 -3400
rect 5520 -3440 5560 -3435
rect 5520 -3470 5525 -3440
rect 5525 -3470 5555 -3440
rect 5555 -3470 5560 -3440
rect 5520 -3475 5560 -3470
rect 5520 -3510 5560 -3505
rect 5520 -3540 5525 -3510
rect 5525 -3540 5555 -3510
rect 5555 -3540 5560 -3510
rect 5520 -3545 5560 -3540
rect 5520 -3580 5560 -3575
rect 5520 -3610 5525 -3580
rect 5525 -3610 5555 -3580
rect 5555 -3610 5560 -3580
rect 5520 -3615 5560 -3610
rect 5520 -3645 5560 -3640
rect 5520 -3675 5525 -3645
rect 5525 -3675 5555 -3645
rect 5555 -3675 5560 -3645
rect 5520 -3680 5560 -3675
rect 5520 -3705 5560 -3700
rect 5520 -3735 5525 -3705
rect 5525 -3735 5555 -3705
rect 5555 -3735 5560 -3705
rect 5520 -3740 5560 -3735
rect 5520 -3770 5560 -3765
rect 5520 -3800 5525 -3770
rect 5525 -3800 5555 -3770
rect 5555 -3800 5560 -3770
rect 5520 -3805 5560 -3800
rect 5520 -3840 5560 -3835
rect 5520 -3870 5525 -3840
rect 5525 -3870 5555 -3840
rect 5555 -3870 5560 -3840
rect 5520 -3875 5560 -3870
rect 5520 -3910 5560 -3905
rect 5520 -3940 5525 -3910
rect 5525 -3940 5555 -3910
rect 5555 -3940 5560 -3910
rect 5520 -3945 5560 -3940
rect 5520 -3980 5560 -3975
rect 5520 -4010 5525 -3980
rect 5525 -4010 5555 -3980
rect 5555 -4010 5560 -3980
rect 5520 -4015 5560 -4010
rect 5520 -4045 5560 -4040
rect 5520 -4075 5525 -4045
rect 5525 -4075 5555 -4045
rect 5555 -4075 5560 -4045
rect 5520 -4080 5560 -4075
rect 5520 -4105 5560 -4100
rect 5520 -4135 5525 -4105
rect 5525 -4135 5555 -4105
rect 5555 -4135 5560 -4105
rect 5520 -4140 5560 -4135
rect 5520 -4170 5560 -4165
rect 5520 -4200 5525 -4170
rect 5525 -4200 5555 -4170
rect 5555 -4200 5560 -4170
rect 5520 -4205 5560 -4200
rect 5520 -4240 5560 -4235
rect 5520 -4270 5525 -4240
rect 5525 -4270 5555 -4240
rect 5555 -4270 5560 -4240
rect 5520 -4275 5560 -4270
rect 5520 -4310 5560 -4305
rect 5520 -4340 5525 -4310
rect 5525 -4340 5555 -4310
rect 5555 -4340 5560 -4310
rect 5520 -4345 5560 -4340
rect 5520 -4380 5560 -4375
rect 5520 -4410 5525 -4380
rect 5525 -4410 5555 -4380
rect 5555 -4410 5560 -4380
rect 5520 -4415 5560 -4410
rect 5520 -4445 5560 -4440
rect 5520 -4475 5525 -4445
rect 5525 -4475 5555 -4445
rect 5555 -4475 5560 -4445
rect 5520 -4480 5560 -4475
rect 5870 -1305 5910 -1300
rect 5870 -1335 5875 -1305
rect 5875 -1335 5905 -1305
rect 5905 -1335 5910 -1305
rect 5870 -1340 5910 -1335
rect 5870 -1370 5910 -1365
rect 5870 -1400 5875 -1370
rect 5875 -1400 5905 -1370
rect 5905 -1400 5910 -1370
rect 5870 -1405 5910 -1400
rect 5870 -1440 5910 -1435
rect 5870 -1470 5875 -1440
rect 5875 -1470 5905 -1440
rect 5905 -1470 5910 -1440
rect 5870 -1475 5910 -1470
rect 5870 -1510 5910 -1505
rect 5870 -1540 5875 -1510
rect 5875 -1540 5905 -1510
rect 5905 -1540 5910 -1510
rect 5870 -1545 5910 -1540
rect 5870 -1580 5910 -1575
rect 5870 -1610 5875 -1580
rect 5875 -1610 5905 -1580
rect 5905 -1610 5910 -1580
rect 5870 -1615 5910 -1610
rect 5870 -1645 5910 -1640
rect 5870 -1675 5875 -1645
rect 5875 -1675 5905 -1645
rect 5905 -1675 5910 -1645
rect 5870 -1680 5910 -1675
rect 5870 -1705 5910 -1700
rect 5870 -1735 5875 -1705
rect 5875 -1735 5905 -1705
rect 5905 -1735 5910 -1705
rect 5870 -1740 5910 -1735
rect 5870 -1770 5910 -1765
rect 5870 -1800 5875 -1770
rect 5875 -1800 5905 -1770
rect 5905 -1800 5910 -1770
rect 5870 -1805 5910 -1800
rect 5870 -1840 5910 -1835
rect 5870 -1870 5875 -1840
rect 5875 -1870 5905 -1840
rect 5905 -1870 5910 -1840
rect 5870 -1875 5910 -1870
rect 5870 -1910 5910 -1905
rect 5870 -1940 5875 -1910
rect 5875 -1940 5905 -1910
rect 5905 -1940 5910 -1910
rect 5870 -1945 5910 -1940
rect 5870 -1980 5910 -1975
rect 5870 -2010 5875 -1980
rect 5875 -2010 5905 -1980
rect 5905 -2010 5910 -1980
rect 5870 -2015 5910 -2010
rect 5870 -2045 5910 -2040
rect 5870 -2075 5875 -2045
rect 5875 -2075 5905 -2045
rect 5905 -2075 5910 -2045
rect 5870 -2080 5910 -2075
rect 5870 -2105 5910 -2100
rect 5870 -2135 5875 -2105
rect 5875 -2135 5905 -2105
rect 5905 -2135 5910 -2105
rect 5870 -2140 5910 -2135
rect 5870 -2170 5910 -2165
rect 5870 -2200 5875 -2170
rect 5875 -2200 5905 -2170
rect 5905 -2200 5910 -2170
rect 5870 -2205 5910 -2200
rect 5870 -2240 5910 -2235
rect 5870 -2270 5875 -2240
rect 5875 -2270 5905 -2240
rect 5905 -2270 5910 -2240
rect 5870 -2275 5910 -2270
rect 5870 -2310 5910 -2305
rect 5870 -2340 5875 -2310
rect 5875 -2340 5905 -2310
rect 5905 -2340 5910 -2310
rect 5870 -2345 5910 -2340
rect 5870 -2380 5910 -2375
rect 5870 -2410 5875 -2380
rect 5875 -2410 5905 -2380
rect 5905 -2410 5910 -2380
rect 5870 -2415 5910 -2410
rect 5870 -2445 5910 -2440
rect 5870 -2475 5875 -2445
rect 5875 -2475 5905 -2445
rect 5905 -2475 5910 -2445
rect 5870 -2480 5910 -2475
rect 5870 -2505 5910 -2500
rect 5870 -2535 5875 -2505
rect 5875 -2535 5905 -2505
rect 5905 -2535 5910 -2505
rect 5870 -2540 5910 -2535
rect 5870 -2570 5910 -2565
rect 5870 -2600 5875 -2570
rect 5875 -2600 5905 -2570
rect 5905 -2600 5910 -2570
rect 5870 -2605 5910 -2600
rect 5870 -2640 5910 -2635
rect 5870 -2670 5875 -2640
rect 5875 -2670 5905 -2640
rect 5905 -2670 5910 -2640
rect 5870 -2675 5910 -2670
rect 5870 -2710 5910 -2705
rect 5870 -2740 5875 -2710
rect 5875 -2740 5905 -2710
rect 5905 -2740 5910 -2710
rect 5870 -2745 5910 -2740
rect 5870 -2780 5910 -2775
rect 5870 -2810 5875 -2780
rect 5875 -2810 5905 -2780
rect 5905 -2810 5910 -2780
rect 5870 -2815 5910 -2810
rect 5870 -2845 5910 -2840
rect 5870 -2875 5875 -2845
rect 5875 -2875 5905 -2845
rect 5905 -2875 5910 -2845
rect 5870 -2880 5910 -2875
rect 5870 -2905 5910 -2900
rect 5870 -2935 5875 -2905
rect 5875 -2935 5905 -2905
rect 5905 -2935 5910 -2905
rect 5870 -2940 5910 -2935
rect 5870 -2970 5910 -2965
rect 5870 -3000 5875 -2970
rect 5875 -3000 5905 -2970
rect 5905 -3000 5910 -2970
rect 5870 -3005 5910 -3000
rect 5870 -3040 5910 -3035
rect 5870 -3070 5875 -3040
rect 5875 -3070 5905 -3040
rect 5905 -3070 5910 -3040
rect 5870 -3075 5910 -3070
rect 5870 -3110 5910 -3105
rect 5870 -3140 5875 -3110
rect 5875 -3140 5905 -3110
rect 5905 -3140 5910 -3110
rect 5870 -3145 5910 -3140
rect 5870 -3180 5910 -3175
rect 5870 -3210 5875 -3180
rect 5875 -3210 5905 -3180
rect 5905 -3210 5910 -3180
rect 5870 -3215 5910 -3210
rect 5870 -3245 5910 -3240
rect 5870 -3275 5875 -3245
rect 5875 -3275 5905 -3245
rect 5905 -3275 5910 -3245
rect 5870 -3280 5910 -3275
rect 5870 -3305 5910 -3300
rect 5870 -3335 5875 -3305
rect 5875 -3335 5905 -3305
rect 5905 -3335 5910 -3305
rect 5870 -3340 5910 -3335
rect 5870 -3370 5910 -3365
rect 5870 -3400 5875 -3370
rect 5875 -3400 5905 -3370
rect 5905 -3400 5910 -3370
rect 5870 -3405 5910 -3400
rect 5870 -3440 5910 -3435
rect 5870 -3470 5875 -3440
rect 5875 -3470 5905 -3440
rect 5905 -3470 5910 -3440
rect 5870 -3475 5910 -3470
rect 5870 -3510 5910 -3505
rect 5870 -3540 5875 -3510
rect 5875 -3540 5905 -3510
rect 5905 -3540 5910 -3510
rect 5870 -3545 5910 -3540
rect 5870 -3580 5910 -3575
rect 5870 -3610 5875 -3580
rect 5875 -3610 5905 -3580
rect 5905 -3610 5910 -3580
rect 5870 -3615 5910 -3610
rect 5870 -3645 5910 -3640
rect 5870 -3675 5875 -3645
rect 5875 -3675 5905 -3645
rect 5905 -3675 5910 -3645
rect 5870 -3680 5910 -3675
rect 5870 -3705 5910 -3700
rect 5870 -3735 5875 -3705
rect 5875 -3735 5905 -3705
rect 5905 -3735 5910 -3705
rect 5870 -3740 5910 -3735
rect 5870 -3770 5910 -3765
rect 5870 -3800 5875 -3770
rect 5875 -3800 5905 -3770
rect 5905 -3800 5910 -3770
rect 5870 -3805 5910 -3800
rect 5870 -3840 5910 -3835
rect 5870 -3870 5875 -3840
rect 5875 -3870 5905 -3840
rect 5905 -3870 5910 -3840
rect 5870 -3875 5910 -3870
rect 5870 -3910 5910 -3905
rect 5870 -3940 5875 -3910
rect 5875 -3940 5905 -3910
rect 5905 -3940 5910 -3910
rect 5870 -3945 5910 -3940
rect 5870 -3980 5910 -3975
rect 5870 -4010 5875 -3980
rect 5875 -4010 5905 -3980
rect 5905 -4010 5910 -3980
rect 5870 -4015 5910 -4010
rect 5870 -4045 5910 -4040
rect 5870 -4075 5875 -4045
rect 5875 -4075 5905 -4045
rect 5905 -4075 5910 -4045
rect 5870 -4080 5910 -4075
rect 5870 -4105 5910 -4100
rect 5870 -4135 5875 -4105
rect 5875 -4135 5905 -4105
rect 5905 -4135 5910 -4105
rect 5870 -4140 5910 -4135
rect 5870 -4170 5910 -4165
rect 5870 -4200 5875 -4170
rect 5875 -4200 5905 -4170
rect 5905 -4200 5910 -4170
rect 5870 -4205 5910 -4200
rect 5870 -4240 5910 -4235
rect 5870 -4270 5875 -4240
rect 5875 -4270 5905 -4240
rect 5905 -4270 5910 -4240
rect 5870 -4275 5910 -4270
rect 5870 -4310 5910 -4305
rect 5870 -4340 5875 -4310
rect 5875 -4340 5905 -4310
rect 5905 -4340 5910 -4310
rect 5870 -4345 5910 -4340
rect 5870 -4380 5910 -4375
rect 5870 -4410 5875 -4380
rect 5875 -4410 5905 -4380
rect 5905 -4410 5910 -4380
rect 5870 -4415 5910 -4410
rect 5870 -4445 5910 -4440
rect 5870 -4475 5875 -4445
rect 5875 -4475 5905 -4445
rect 5905 -4475 5910 -4445
rect 5870 -4480 5910 -4475
rect 6220 -1305 6260 -1300
rect 6220 -1335 6225 -1305
rect 6225 -1335 6255 -1305
rect 6255 -1335 6260 -1305
rect 6220 -1340 6260 -1335
rect 6220 -1370 6260 -1365
rect 6220 -1400 6225 -1370
rect 6225 -1400 6255 -1370
rect 6255 -1400 6260 -1370
rect 6220 -1405 6260 -1400
rect 6220 -1440 6260 -1435
rect 6220 -1470 6225 -1440
rect 6225 -1470 6255 -1440
rect 6255 -1470 6260 -1440
rect 6220 -1475 6260 -1470
rect 6220 -1510 6260 -1505
rect 6220 -1540 6225 -1510
rect 6225 -1540 6255 -1510
rect 6255 -1540 6260 -1510
rect 6220 -1545 6260 -1540
rect 6220 -1580 6260 -1575
rect 6220 -1610 6225 -1580
rect 6225 -1610 6255 -1580
rect 6255 -1610 6260 -1580
rect 6220 -1615 6260 -1610
rect 6220 -1645 6260 -1640
rect 6220 -1675 6225 -1645
rect 6225 -1675 6255 -1645
rect 6255 -1675 6260 -1645
rect 6220 -1680 6260 -1675
rect 6220 -1705 6260 -1700
rect 6220 -1735 6225 -1705
rect 6225 -1735 6255 -1705
rect 6255 -1735 6260 -1705
rect 6220 -1740 6260 -1735
rect 6220 -1770 6260 -1765
rect 6220 -1800 6225 -1770
rect 6225 -1800 6255 -1770
rect 6255 -1800 6260 -1770
rect 6220 -1805 6260 -1800
rect 6220 -1840 6260 -1835
rect 6220 -1870 6225 -1840
rect 6225 -1870 6255 -1840
rect 6255 -1870 6260 -1840
rect 6220 -1875 6260 -1870
rect 6220 -1910 6260 -1905
rect 6220 -1940 6225 -1910
rect 6225 -1940 6255 -1910
rect 6255 -1940 6260 -1910
rect 6220 -1945 6260 -1940
rect 6220 -1980 6260 -1975
rect 6220 -2010 6225 -1980
rect 6225 -2010 6255 -1980
rect 6255 -2010 6260 -1980
rect 6220 -2015 6260 -2010
rect 6220 -2045 6260 -2040
rect 6220 -2075 6225 -2045
rect 6225 -2075 6255 -2045
rect 6255 -2075 6260 -2045
rect 6220 -2080 6260 -2075
rect 6220 -2105 6260 -2100
rect 6220 -2135 6225 -2105
rect 6225 -2135 6255 -2105
rect 6255 -2135 6260 -2105
rect 6220 -2140 6260 -2135
rect 6220 -2170 6260 -2165
rect 6220 -2200 6225 -2170
rect 6225 -2200 6255 -2170
rect 6255 -2200 6260 -2170
rect 6220 -2205 6260 -2200
rect 6220 -2240 6260 -2235
rect 6220 -2270 6225 -2240
rect 6225 -2270 6255 -2240
rect 6255 -2270 6260 -2240
rect 6220 -2275 6260 -2270
rect 6220 -2310 6260 -2305
rect 6220 -2340 6225 -2310
rect 6225 -2340 6255 -2310
rect 6255 -2340 6260 -2310
rect 6220 -2345 6260 -2340
rect 6220 -2380 6260 -2375
rect 6220 -2410 6225 -2380
rect 6225 -2410 6255 -2380
rect 6255 -2410 6260 -2380
rect 6220 -2415 6260 -2410
rect 6220 -2445 6260 -2440
rect 6220 -2475 6225 -2445
rect 6225 -2475 6255 -2445
rect 6255 -2475 6260 -2445
rect 6220 -2480 6260 -2475
rect 6220 -2505 6260 -2500
rect 6220 -2535 6225 -2505
rect 6225 -2535 6255 -2505
rect 6255 -2535 6260 -2505
rect 6220 -2540 6260 -2535
rect 6220 -2570 6260 -2565
rect 6220 -2600 6225 -2570
rect 6225 -2600 6255 -2570
rect 6255 -2600 6260 -2570
rect 6220 -2605 6260 -2600
rect 6220 -2640 6260 -2635
rect 6220 -2670 6225 -2640
rect 6225 -2670 6255 -2640
rect 6255 -2670 6260 -2640
rect 6220 -2675 6260 -2670
rect 6220 -2710 6260 -2705
rect 6220 -2740 6225 -2710
rect 6225 -2740 6255 -2710
rect 6255 -2740 6260 -2710
rect 6220 -2745 6260 -2740
rect 6220 -2780 6260 -2775
rect 6220 -2810 6225 -2780
rect 6225 -2810 6255 -2780
rect 6255 -2810 6260 -2780
rect 6220 -2815 6260 -2810
rect 6220 -2845 6260 -2840
rect 6220 -2875 6225 -2845
rect 6225 -2875 6255 -2845
rect 6255 -2875 6260 -2845
rect 6220 -2880 6260 -2875
rect 6220 -2905 6260 -2900
rect 6220 -2935 6225 -2905
rect 6225 -2935 6255 -2905
rect 6255 -2935 6260 -2905
rect 6220 -2940 6260 -2935
rect 6220 -2970 6260 -2965
rect 6220 -3000 6225 -2970
rect 6225 -3000 6255 -2970
rect 6255 -3000 6260 -2970
rect 6220 -3005 6260 -3000
rect 6220 -3040 6260 -3035
rect 6220 -3070 6225 -3040
rect 6225 -3070 6255 -3040
rect 6255 -3070 6260 -3040
rect 6220 -3075 6260 -3070
rect 6220 -3110 6260 -3105
rect 6220 -3140 6225 -3110
rect 6225 -3140 6255 -3110
rect 6255 -3140 6260 -3110
rect 6220 -3145 6260 -3140
rect 6220 -3180 6260 -3175
rect 6220 -3210 6225 -3180
rect 6225 -3210 6255 -3180
rect 6255 -3210 6260 -3180
rect 6220 -3215 6260 -3210
rect 6220 -3245 6260 -3240
rect 6220 -3275 6225 -3245
rect 6225 -3275 6255 -3245
rect 6255 -3275 6260 -3245
rect 6220 -3280 6260 -3275
rect 6220 -3305 6260 -3300
rect 6220 -3335 6225 -3305
rect 6225 -3335 6255 -3305
rect 6255 -3335 6260 -3305
rect 6220 -3340 6260 -3335
rect 6220 -3370 6260 -3365
rect 6220 -3400 6225 -3370
rect 6225 -3400 6255 -3370
rect 6255 -3400 6260 -3370
rect 6220 -3405 6260 -3400
rect 6220 -3440 6260 -3435
rect 6220 -3470 6225 -3440
rect 6225 -3470 6255 -3440
rect 6255 -3470 6260 -3440
rect 6220 -3475 6260 -3470
rect 6220 -3510 6260 -3505
rect 6220 -3540 6225 -3510
rect 6225 -3540 6255 -3510
rect 6255 -3540 6260 -3510
rect 6220 -3545 6260 -3540
rect 6220 -3580 6260 -3575
rect 6220 -3610 6225 -3580
rect 6225 -3610 6255 -3580
rect 6255 -3610 6260 -3580
rect 6220 -3615 6260 -3610
rect 6220 -3645 6260 -3640
rect 6220 -3675 6225 -3645
rect 6225 -3675 6255 -3645
rect 6255 -3675 6260 -3645
rect 6220 -3680 6260 -3675
rect 6220 -3705 6260 -3700
rect 6220 -3735 6225 -3705
rect 6225 -3735 6255 -3705
rect 6255 -3735 6260 -3705
rect 6220 -3740 6260 -3735
rect 6220 -3770 6260 -3765
rect 6220 -3800 6225 -3770
rect 6225 -3800 6255 -3770
rect 6255 -3800 6260 -3770
rect 6220 -3805 6260 -3800
rect 6220 -3840 6260 -3835
rect 6220 -3870 6225 -3840
rect 6225 -3870 6255 -3840
rect 6255 -3870 6260 -3840
rect 6220 -3875 6260 -3870
rect 6220 -3910 6260 -3905
rect 6220 -3940 6225 -3910
rect 6225 -3940 6255 -3910
rect 6255 -3940 6260 -3910
rect 6220 -3945 6260 -3940
rect 6220 -3980 6260 -3975
rect 6220 -4010 6225 -3980
rect 6225 -4010 6255 -3980
rect 6255 -4010 6260 -3980
rect 6220 -4015 6260 -4010
rect 6220 -4045 6260 -4040
rect 6220 -4075 6225 -4045
rect 6225 -4075 6255 -4045
rect 6255 -4075 6260 -4045
rect 6220 -4080 6260 -4075
rect 6220 -4105 6260 -4100
rect 6220 -4135 6225 -4105
rect 6225 -4135 6255 -4105
rect 6255 -4135 6260 -4105
rect 6220 -4140 6260 -4135
rect 6220 -4170 6260 -4165
rect 6220 -4200 6225 -4170
rect 6225 -4200 6255 -4170
rect 6255 -4200 6260 -4170
rect 6220 -4205 6260 -4200
rect 6220 -4240 6260 -4235
rect 6220 -4270 6225 -4240
rect 6225 -4270 6255 -4240
rect 6255 -4270 6260 -4240
rect 6220 -4275 6260 -4270
rect 6220 -4310 6260 -4305
rect 6220 -4340 6225 -4310
rect 6225 -4340 6255 -4310
rect 6255 -4340 6260 -4310
rect 6220 -4345 6260 -4340
rect 6220 -4380 6260 -4375
rect 6220 -4410 6225 -4380
rect 6225 -4410 6255 -4380
rect 6255 -4410 6260 -4380
rect 6220 -4415 6260 -4410
rect 6220 -4445 6260 -4440
rect 6220 -4475 6225 -4445
rect 6225 -4475 6255 -4445
rect 6255 -4475 6260 -4445
rect 6220 -4480 6260 -4475
rect 6570 -1305 6610 -1300
rect 6570 -1335 6575 -1305
rect 6575 -1335 6605 -1305
rect 6605 -1335 6610 -1305
rect 6570 -1340 6610 -1335
rect 6570 -1370 6610 -1365
rect 6570 -1400 6575 -1370
rect 6575 -1400 6605 -1370
rect 6605 -1400 6610 -1370
rect 6570 -1405 6610 -1400
rect 6570 -1440 6610 -1435
rect 6570 -1470 6575 -1440
rect 6575 -1470 6605 -1440
rect 6605 -1470 6610 -1440
rect 6570 -1475 6610 -1470
rect 6570 -1510 6610 -1505
rect 6570 -1540 6575 -1510
rect 6575 -1540 6605 -1510
rect 6605 -1540 6610 -1510
rect 6570 -1545 6610 -1540
rect 6570 -1580 6610 -1575
rect 6570 -1610 6575 -1580
rect 6575 -1610 6605 -1580
rect 6605 -1610 6610 -1580
rect 6570 -1615 6610 -1610
rect 6570 -1645 6610 -1640
rect 6570 -1675 6575 -1645
rect 6575 -1675 6605 -1645
rect 6605 -1675 6610 -1645
rect 6570 -1680 6610 -1675
rect 6570 -1705 6610 -1700
rect 6570 -1735 6575 -1705
rect 6575 -1735 6605 -1705
rect 6605 -1735 6610 -1705
rect 6570 -1740 6610 -1735
rect 6570 -1770 6610 -1765
rect 6570 -1800 6575 -1770
rect 6575 -1800 6605 -1770
rect 6605 -1800 6610 -1770
rect 6570 -1805 6610 -1800
rect 6570 -1840 6610 -1835
rect 6570 -1870 6575 -1840
rect 6575 -1870 6605 -1840
rect 6605 -1870 6610 -1840
rect 6570 -1875 6610 -1870
rect 6570 -1910 6610 -1905
rect 6570 -1940 6575 -1910
rect 6575 -1940 6605 -1910
rect 6605 -1940 6610 -1910
rect 6570 -1945 6610 -1940
rect 6570 -1980 6610 -1975
rect 6570 -2010 6575 -1980
rect 6575 -2010 6605 -1980
rect 6605 -2010 6610 -1980
rect 6570 -2015 6610 -2010
rect 6570 -2045 6610 -2040
rect 6570 -2075 6575 -2045
rect 6575 -2075 6605 -2045
rect 6605 -2075 6610 -2045
rect 6570 -2080 6610 -2075
rect 6570 -2105 6610 -2100
rect 6570 -2135 6575 -2105
rect 6575 -2135 6605 -2105
rect 6605 -2135 6610 -2105
rect 6570 -2140 6610 -2135
rect 6570 -2170 6610 -2165
rect 6570 -2200 6575 -2170
rect 6575 -2200 6605 -2170
rect 6605 -2200 6610 -2170
rect 6570 -2205 6610 -2200
rect 6570 -2240 6610 -2235
rect 6570 -2270 6575 -2240
rect 6575 -2270 6605 -2240
rect 6605 -2270 6610 -2240
rect 6570 -2275 6610 -2270
rect 6570 -2310 6610 -2305
rect 6570 -2340 6575 -2310
rect 6575 -2340 6605 -2310
rect 6605 -2340 6610 -2310
rect 6570 -2345 6610 -2340
rect 6570 -2380 6610 -2375
rect 6570 -2410 6575 -2380
rect 6575 -2410 6605 -2380
rect 6605 -2410 6610 -2380
rect 6570 -2415 6610 -2410
rect 6570 -2445 6610 -2440
rect 6570 -2475 6575 -2445
rect 6575 -2475 6605 -2445
rect 6605 -2475 6610 -2445
rect 6570 -2480 6610 -2475
rect 6570 -2505 6610 -2500
rect 6570 -2535 6575 -2505
rect 6575 -2535 6605 -2505
rect 6605 -2535 6610 -2505
rect 6570 -2540 6610 -2535
rect 6570 -2570 6610 -2565
rect 6570 -2600 6575 -2570
rect 6575 -2600 6605 -2570
rect 6605 -2600 6610 -2570
rect 6570 -2605 6610 -2600
rect 6570 -2640 6610 -2635
rect 6570 -2670 6575 -2640
rect 6575 -2670 6605 -2640
rect 6605 -2670 6610 -2640
rect 6570 -2675 6610 -2670
rect 6570 -2710 6610 -2705
rect 6570 -2740 6575 -2710
rect 6575 -2740 6605 -2710
rect 6605 -2740 6610 -2710
rect 6570 -2745 6610 -2740
rect 6570 -2780 6610 -2775
rect 6570 -2810 6575 -2780
rect 6575 -2810 6605 -2780
rect 6605 -2810 6610 -2780
rect 6570 -2815 6610 -2810
rect 6570 -2845 6610 -2840
rect 6570 -2875 6575 -2845
rect 6575 -2875 6605 -2845
rect 6605 -2875 6610 -2845
rect 6570 -2880 6610 -2875
rect 6570 -2905 6610 -2900
rect 6570 -2935 6575 -2905
rect 6575 -2935 6605 -2905
rect 6605 -2935 6610 -2905
rect 6570 -2940 6610 -2935
rect 6570 -2970 6610 -2965
rect 6570 -3000 6575 -2970
rect 6575 -3000 6605 -2970
rect 6605 -3000 6610 -2970
rect 6570 -3005 6610 -3000
rect 6570 -3040 6610 -3035
rect 6570 -3070 6575 -3040
rect 6575 -3070 6605 -3040
rect 6605 -3070 6610 -3040
rect 6570 -3075 6610 -3070
rect 6570 -3110 6610 -3105
rect 6570 -3140 6575 -3110
rect 6575 -3140 6605 -3110
rect 6605 -3140 6610 -3110
rect 6570 -3145 6610 -3140
rect 6570 -3180 6610 -3175
rect 6570 -3210 6575 -3180
rect 6575 -3210 6605 -3180
rect 6605 -3210 6610 -3180
rect 6570 -3215 6610 -3210
rect 6570 -3245 6610 -3240
rect 6570 -3275 6575 -3245
rect 6575 -3275 6605 -3245
rect 6605 -3275 6610 -3245
rect 6570 -3280 6610 -3275
rect 6570 -3305 6610 -3300
rect 6570 -3335 6575 -3305
rect 6575 -3335 6605 -3305
rect 6605 -3335 6610 -3305
rect 6570 -3340 6610 -3335
rect 6570 -3370 6610 -3365
rect 6570 -3400 6575 -3370
rect 6575 -3400 6605 -3370
rect 6605 -3400 6610 -3370
rect 6570 -3405 6610 -3400
rect 6570 -3440 6610 -3435
rect 6570 -3470 6575 -3440
rect 6575 -3470 6605 -3440
rect 6605 -3470 6610 -3440
rect 6570 -3475 6610 -3470
rect 6570 -3510 6610 -3505
rect 6570 -3540 6575 -3510
rect 6575 -3540 6605 -3510
rect 6605 -3540 6610 -3510
rect 6570 -3545 6610 -3540
rect 6570 -3580 6610 -3575
rect 6570 -3610 6575 -3580
rect 6575 -3610 6605 -3580
rect 6605 -3610 6610 -3580
rect 6570 -3615 6610 -3610
rect 6570 -3645 6610 -3640
rect 6570 -3675 6575 -3645
rect 6575 -3675 6605 -3645
rect 6605 -3675 6610 -3645
rect 6570 -3680 6610 -3675
rect 6570 -3705 6610 -3700
rect 6570 -3735 6575 -3705
rect 6575 -3735 6605 -3705
rect 6605 -3735 6610 -3705
rect 6570 -3740 6610 -3735
rect 6570 -3770 6610 -3765
rect 6570 -3800 6575 -3770
rect 6575 -3800 6605 -3770
rect 6605 -3800 6610 -3770
rect 6570 -3805 6610 -3800
rect 6570 -3840 6610 -3835
rect 6570 -3870 6575 -3840
rect 6575 -3870 6605 -3840
rect 6605 -3870 6610 -3840
rect 6570 -3875 6610 -3870
rect 6570 -3910 6610 -3905
rect 6570 -3940 6575 -3910
rect 6575 -3940 6605 -3910
rect 6605 -3940 6610 -3910
rect 6570 -3945 6610 -3940
rect 6570 -3980 6610 -3975
rect 6570 -4010 6575 -3980
rect 6575 -4010 6605 -3980
rect 6605 -4010 6610 -3980
rect 6570 -4015 6610 -4010
rect 6570 -4045 6610 -4040
rect 6570 -4075 6575 -4045
rect 6575 -4075 6605 -4045
rect 6605 -4075 6610 -4045
rect 6570 -4080 6610 -4075
rect 6570 -4105 6610 -4100
rect 6570 -4135 6575 -4105
rect 6575 -4135 6605 -4105
rect 6605 -4135 6610 -4105
rect 6570 -4140 6610 -4135
rect 6570 -4170 6610 -4165
rect 6570 -4200 6575 -4170
rect 6575 -4200 6605 -4170
rect 6605 -4200 6610 -4170
rect 6570 -4205 6610 -4200
rect 6570 -4240 6610 -4235
rect 6570 -4270 6575 -4240
rect 6575 -4270 6605 -4240
rect 6605 -4270 6610 -4240
rect 6570 -4275 6610 -4270
rect 6570 -4310 6610 -4305
rect 6570 -4340 6575 -4310
rect 6575 -4340 6605 -4310
rect 6605 -4340 6610 -4310
rect 6570 -4345 6610 -4340
rect 6570 -4380 6610 -4375
rect 6570 -4410 6575 -4380
rect 6575 -4410 6605 -4380
rect 6605 -4410 6610 -4380
rect 6570 -4415 6610 -4410
rect 6570 -4445 6610 -4440
rect 6570 -4475 6575 -4445
rect 6575 -4475 6605 -4445
rect 6605 -4475 6610 -4445
rect 6570 -4480 6610 -4475
rect 6920 -1305 6960 -1300
rect 6920 -1335 6925 -1305
rect 6925 -1335 6955 -1305
rect 6955 -1335 6960 -1305
rect 6920 -1340 6960 -1335
rect 6920 -1370 6960 -1365
rect 6920 -1400 6925 -1370
rect 6925 -1400 6955 -1370
rect 6955 -1400 6960 -1370
rect 6920 -1405 6960 -1400
rect 6920 -1440 6960 -1435
rect 6920 -1470 6925 -1440
rect 6925 -1470 6955 -1440
rect 6955 -1470 6960 -1440
rect 6920 -1475 6960 -1470
rect 6920 -1510 6960 -1505
rect 6920 -1540 6925 -1510
rect 6925 -1540 6955 -1510
rect 6955 -1540 6960 -1510
rect 6920 -1545 6960 -1540
rect 6920 -1580 6960 -1575
rect 6920 -1610 6925 -1580
rect 6925 -1610 6955 -1580
rect 6955 -1610 6960 -1580
rect 6920 -1615 6960 -1610
rect 6920 -1645 6960 -1640
rect 6920 -1675 6925 -1645
rect 6925 -1675 6955 -1645
rect 6955 -1675 6960 -1645
rect 6920 -1680 6960 -1675
rect 6920 -1705 6960 -1700
rect 6920 -1735 6925 -1705
rect 6925 -1735 6955 -1705
rect 6955 -1735 6960 -1705
rect 6920 -1740 6960 -1735
rect 6920 -1770 6960 -1765
rect 6920 -1800 6925 -1770
rect 6925 -1800 6955 -1770
rect 6955 -1800 6960 -1770
rect 6920 -1805 6960 -1800
rect 6920 -1840 6960 -1835
rect 6920 -1870 6925 -1840
rect 6925 -1870 6955 -1840
rect 6955 -1870 6960 -1840
rect 6920 -1875 6960 -1870
rect 6920 -1910 6960 -1905
rect 6920 -1940 6925 -1910
rect 6925 -1940 6955 -1910
rect 6955 -1940 6960 -1910
rect 6920 -1945 6960 -1940
rect 6920 -1980 6960 -1975
rect 6920 -2010 6925 -1980
rect 6925 -2010 6955 -1980
rect 6955 -2010 6960 -1980
rect 6920 -2015 6960 -2010
rect 6920 -2045 6960 -2040
rect 6920 -2075 6925 -2045
rect 6925 -2075 6955 -2045
rect 6955 -2075 6960 -2045
rect 6920 -2080 6960 -2075
rect 6920 -2105 6960 -2100
rect 6920 -2135 6925 -2105
rect 6925 -2135 6955 -2105
rect 6955 -2135 6960 -2105
rect 6920 -2140 6960 -2135
rect 6920 -2170 6960 -2165
rect 6920 -2200 6925 -2170
rect 6925 -2200 6955 -2170
rect 6955 -2200 6960 -2170
rect 6920 -2205 6960 -2200
rect 6920 -2240 6960 -2235
rect 6920 -2270 6925 -2240
rect 6925 -2270 6955 -2240
rect 6955 -2270 6960 -2240
rect 6920 -2275 6960 -2270
rect 6920 -2310 6960 -2305
rect 6920 -2340 6925 -2310
rect 6925 -2340 6955 -2310
rect 6955 -2340 6960 -2310
rect 6920 -2345 6960 -2340
rect 6920 -2380 6960 -2375
rect 6920 -2410 6925 -2380
rect 6925 -2410 6955 -2380
rect 6955 -2410 6960 -2380
rect 6920 -2415 6960 -2410
rect 6920 -2445 6960 -2440
rect 6920 -2475 6925 -2445
rect 6925 -2475 6955 -2445
rect 6955 -2475 6960 -2445
rect 6920 -2480 6960 -2475
rect 6920 -2505 6960 -2500
rect 6920 -2535 6925 -2505
rect 6925 -2535 6955 -2505
rect 6955 -2535 6960 -2505
rect 6920 -2540 6960 -2535
rect 6920 -2570 6960 -2565
rect 6920 -2600 6925 -2570
rect 6925 -2600 6955 -2570
rect 6955 -2600 6960 -2570
rect 6920 -2605 6960 -2600
rect 6920 -2640 6960 -2635
rect 6920 -2670 6925 -2640
rect 6925 -2670 6955 -2640
rect 6955 -2670 6960 -2640
rect 6920 -2675 6960 -2670
rect 6920 -2710 6960 -2705
rect 6920 -2740 6925 -2710
rect 6925 -2740 6955 -2710
rect 6955 -2740 6960 -2710
rect 6920 -2745 6960 -2740
rect 6920 -2780 6960 -2775
rect 6920 -2810 6925 -2780
rect 6925 -2810 6955 -2780
rect 6955 -2810 6960 -2780
rect 6920 -2815 6960 -2810
rect 6920 -2845 6960 -2840
rect 6920 -2875 6925 -2845
rect 6925 -2875 6955 -2845
rect 6955 -2875 6960 -2845
rect 6920 -2880 6960 -2875
rect 6920 -2905 6960 -2900
rect 6920 -2935 6925 -2905
rect 6925 -2935 6955 -2905
rect 6955 -2935 6960 -2905
rect 6920 -2940 6960 -2935
rect 6920 -2970 6960 -2965
rect 6920 -3000 6925 -2970
rect 6925 -3000 6955 -2970
rect 6955 -3000 6960 -2970
rect 6920 -3005 6960 -3000
rect 6920 -3040 6960 -3035
rect 6920 -3070 6925 -3040
rect 6925 -3070 6955 -3040
rect 6955 -3070 6960 -3040
rect 6920 -3075 6960 -3070
rect 6920 -3110 6960 -3105
rect 6920 -3140 6925 -3110
rect 6925 -3140 6955 -3110
rect 6955 -3140 6960 -3110
rect 6920 -3145 6960 -3140
rect 6920 -3180 6960 -3175
rect 6920 -3210 6925 -3180
rect 6925 -3210 6955 -3180
rect 6955 -3210 6960 -3180
rect 6920 -3215 6960 -3210
rect 6920 -3245 6960 -3240
rect 6920 -3275 6925 -3245
rect 6925 -3275 6955 -3245
rect 6955 -3275 6960 -3245
rect 6920 -3280 6960 -3275
rect 6920 -3305 6960 -3300
rect 6920 -3335 6925 -3305
rect 6925 -3335 6955 -3305
rect 6955 -3335 6960 -3305
rect 6920 -3340 6960 -3335
rect 6920 -3370 6960 -3365
rect 6920 -3400 6925 -3370
rect 6925 -3400 6955 -3370
rect 6955 -3400 6960 -3370
rect 6920 -3405 6960 -3400
rect 6920 -3440 6960 -3435
rect 6920 -3470 6925 -3440
rect 6925 -3470 6955 -3440
rect 6955 -3470 6960 -3440
rect 6920 -3475 6960 -3470
rect 6920 -3510 6960 -3505
rect 6920 -3540 6925 -3510
rect 6925 -3540 6955 -3510
rect 6955 -3540 6960 -3510
rect 6920 -3545 6960 -3540
rect 6920 -3580 6960 -3575
rect 6920 -3610 6925 -3580
rect 6925 -3610 6955 -3580
rect 6955 -3610 6960 -3580
rect 6920 -3615 6960 -3610
rect 6920 -3645 6960 -3640
rect 6920 -3675 6925 -3645
rect 6925 -3675 6955 -3645
rect 6955 -3675 6960 -3645
rect 6920 -3680 6960 -3675
rect 6920 -3705 6960 -3700
rect 6920 -3735 6925 -3705
rect 6925 -3735 6955 -3705
rect 6955 -3735 6960 -3705
rect 6920 -3740 6960 -3735
rect 6920 -3770 6960 -3765
rect 6920 -3800 6925 -3770
rect 6925 -3800 6955 -3770
rect 6955 -3800 6960 -3770
rect 6920 -3805 6960 -3800
rect 6920 -3840 6960 -3835
rect 6920 -3870 6925 -3840
rect 6925 -3870 6955 -3840
rect 6955 -3870 6960 -3840
rect 6920 -3875 6960 -3870
rect 6920 -3910 6960 -3905
rect 6920 -3940 6925 -3910
rect 6925 -3940 6955 -3910
rect 6955 -3940 6960 -3910
rect 6920 -3945 6960 -3940
rect 6920 -3980 6960 -3975
rect 6920 -4010 6925 -3980
rect 6925 -4010 6955 -3980
rect 6955 -4010 6960 -3980
rect 6920 -4015 6960 -4010
rect 6920 -4045 6960 -4040
rect 6920 -4075 6925 -4045
rect 6925 -4075 6955 -4045
rect 6955 -4075 6960 -4045
rect 6920 -4080 6960 -4075
rect 6920 -4105 6960 -4100
rect 6920 -4135 6925 -4105
rect 6925 -4135 6955 -4105
rect 6955 -4135 6960 -4105
rect 6920 -4140 6960 -4135
rect 6920 -4170 6960 -4165
rect 6920 -4200 6925 -4170
rect 6925 -4200 6955 -4170
rect 6955 -4200 6960 -4170
rect 6920 -4205 6960 -4200
rect 6920 -4240 6960 -4235
rect 6920 -4270 6925 -4240
rect 6925 -4270 6955 -4240
rect 6955 -4270 6960 -4240
rect 6920 -4275 6960 -4270
rect 6920 -4310 6960 -4305
rect 6920 -4340 6925 -4310
rect 6925 -4340 6955 -4310
rect 6955 -4340 6960 -4310
rect 6920 -4345 6960 -4340
rect 6920 -4380 6960 -4375
rect 6920 -4410 6925 -4380
rect 6925 -4410 6955 -4380
rect 6955 -4410 6960 -4380
rect 6920 -4415 6960 -4410
rect 6920 -4445 6960 -4440
rect 6920 -4475 6925 -4445
rect 6925 -4475 6955 -4445
rect 6955 -4475 6960 -4445
rect 6920 -4480 6960 -4475
rect 7270 -1305 7310 -1300
rect 7270 -1335 7275 -1305
rect 7275 -1335 7305 -1305
rect 7305 -1335 7310 -1305
rect 7270 -1340 7310 -1335
rect 7270 -1370 7310 -1365
rect 7270 -1400 7275 -1370
rect 7275 -1400 7305 -1370
rect 7305 -1400 7310 -1370
rect 7270 -1405 7310 -1400
rect 7270 -1440 7310 -1435
rect 7270 -1470 7275 -1440
rect 7275 -1470 7305 -1440
rect 7305 -1470 7310 -1440
rect 7270 -1475 7310 -1470
rect 7270 -1510 7310 -1505
rect 7270 -1540 7275 -1510
rect 7275 -1540 7305 -1510
rect 7305 -1540 7310 -1510
rect 7270 -1545 7310 -1540
rect 7270 -1580 7310 -1575
rect 7270 -1610 7275 -1580
rect 7275 -1610 7305 -1580
rect 7305 -1610 7310 -1580
rect 7270 -1615 7310 -1610
rect 7270 -1645 7310 -1640
rect 7270 -1675 7275 -1645
rect 7275 -1675 7305 -1645
rect 7305 -1675 7310 -1645
rect 7270 -1680 7310 -1675
rect 7270 -1705 7310 -1700
rect 7270 -1735 7275 -1705
rect 7275 -1735 7305 -1705
rect 7305 -1735 7310 -1705
rect 7270 -1740 7310 -1735
rect 7270 -1770 7310 -1765
rect 7270 -1800 7275 -1770
rect 7275 -1800 7305 -1770
rect 7305 -1800 7310 -1770
rect 7270 -1805 7310 -1800
rect 7270 -1840 7310 -1835
rect 7270 -1870 7275 -1840
rect 7275 -1870 7305 -1840
rect 7305 -1870 7310 -1840
rect 7270 -1875 7310 -1870
rect 7270 -1910 7310 -1905
rect 7270 -1940 7275 -1910
rect 7275 -1940 7305 -1910
rect 7305 -1940 7310 -1910
rect 7270 -1945 7310 -1940
rect 7270 -1980 7310 -1975
rect 7270 -2010 7275 -1980
rect 7275 -2010 7305 -1980
rect 7305 -2010 7310 -1980
rect 7270 -2015 7310 -2010
rect 7270 -2045 7310 -2040
rect 7270 -2075 7275 -2045
rect 7275 -2075 7305 -2045
rect 7305 -2075 7310 -2045
rect 7270 -2080 7310 -2075
rect 7270 -2105 7310 -2100
rect 7270 -2135 7275 -2105
rect 7275 -2135 7305 -2105
rect 7305 -2135 7310 -2105
rect 7270 -2140 7310 -2135
rect 7270 -2170 7310 -2165
rect 7270 -2200 7275 -2170
rect 7275 -2200 7305 -2170
rect 7305 -2200 7310 -2170
rect 7270 -2205 7310 -2200
rect 7270 -2240 7310 -2235
rect 7270 -2270 7275 -2240
rect 7275 -2270 7305 -2240
rect 7305 -2270 7310 -2240
rect 7270 -2275 7310 -2270
rect 7270 -2310 7310 -2305
rect 7270 -2340 7275 -2310
rect 7275 -2340 7305 -2310
rect 7305 -2340 7310 -2310
rect 7270 -2345 7310 -2340
rect 7270 -2380 7310 -2375
rect 7270 -2410 7275 -2380
rect 7275 -2410 7305 -2380
rect 7305 -2410 7310 -2380
rect 7270 -2415 7310 -2410
rect 7270 -2445 7310 -2440
rect 7270 -2475 7275 -2445
rect 7275 -2475 7305 -2445
rect 7305 -2475 7310 -2445
rect 7270 -2480 7310 -2475
rect 7270 -2505 7310 -2500
rect 7270 -2535 7275 -2505
rect 7275 -2535 7305 -2505
rect 7305 -2535 7310 -2505
rect 7270 -2540 7310 -2535
rect 7270 -2570 7310 -2565
rect 7270 -2600 7275 -2570
rect 7275 -2600 7305 -2570
rect 7305 -2600 7310 -2570
rect 7270 -2605 7310 -2600
rect 7270 -2640 7310 -2635
rect 7270 -2670 7275 -2640
rect 7275 -2670 7305 -2640
rect 7305 -2670 7310 -2640
rect 7270 -2675 7310 -2670
rect 7270 -2710 7310 -2705
rect 7270 -2740 7275 -2710
rect 7275 -2740 7305 -2710
rect 7305 -2740 7310 -2710
rect 7270 -2745 7310 -2740
rect 7270 -2780 7310 -2775
rect 7270 -2810 7275 -2780
rect 7275 -2810 7305 -2780
rect 7305 -2810 7310 -2780
rect 7270 -2815 7310 -2810
rect 7270 -2845 7310 -2840
rect 7270 -2875 7275 -2845
rect 7275 -2875 7305 -2845
rect 7305 -2875 7310 -2845
rect 7270 -2880 7310 -2875
rect 7270 -2905 7310 -2900
rect 7270 -2935 7275 -2905
rect 7275 -2935 7305 -2905
rect 7305 -2935 7310 -2905
rect 7270 -2940 7310 -2935
rect 7270 -2970 7310 -2965
rect 7270 -3000 7275 -2970
rect 7275 -3000 7305 -2970
rect 7305 -3000 7310 -2970
rect 7270 -3005 7310 -3000
rect 7270 -3040 7310 -3035
rect 7270 -3070 7275 -3040
rect 7275 -3070 7305 -3040
rect 7305 -3070 7310 -3040
rect 7270 -3075 7310 -3070
rect 7270 -3110 7310 -3105
rect 7270 -3140 7275 -3110
rect 7275 -3140 7305 -3110
rect 7305 -3140 7310 -3110
rect 7270 -3145 7310 -3140
rect 7270 -3180 7310 -3175
rect 7270 -3210 7275 -3180
rect 7275 -3210 7305 -3180
rect 7305 -3210 7310 -3180
rect 7270 -3215 7310 -3210
rect 7270 -3245 7310 -3240
rect 7270 -3275 7275 -3245
rect 7275 -3275 7305 -3245
rect 7305 -3275 7310 -3245
rect 7270 -3280 7310 -3275
rect 7270 -3305 7310 -3300
rect 7270 -3335 7275 -3305
rect 7275 -3335 7305 -3305
rect 7305 -3335 7310 -3305
rect 7270 -3340 7310 -3335
rect 7270 -3370 7310 -3365
rect 7270 -3400 7275 -3370
rect 7275 -3400 7305 -3370
rect 7305 -3400 7310 -3370
rect 7270 -3405 7310 -3400
rect 7270 -3440 7310 -3435
rect 7270 -3470 7275 -3440
rect 7275 -3470 7305 -3440
rect 7305 -3470 7310 -3440
rect 7270 -3475 7310 -3470
rect 7270 -3510 7310 -3505
rect 7270 -3540 7275 -3510
rect 7275 -3540 7305 -3510
rect 7305 -3540 7310 -3510
rect 7270 -3545 7310 -3540
rect 7270 -3580 7310 -3575
rect 7270 -3610 7275 -3580
rect 7275 -3610 7305 -3580
rect 7305 -3610 7310 -3580
rect 7270 -3615 7310 -3610
rect 7270 -3645 7310 -3640
rect 7270 -3675 7275 -3645
rect 7275 -3675 7305 -3645
rect 7305 -3675 7310 -3645
rect 7270 -3680 7310 -3675
rect 7270 -3705 7310 -3700
rect 7270 -3735 7275 -3705
rect 7275 -3735 7305 -3705
rect 7305 -3735 7310 -3705
rect 7270 -3740 7310 -3735
rect 7270 -3770 7310 -3765
rect 7270 -3800 7275 -3770
rect 7275 -3800 7305 -3770
rect 7305 -3800 7310 -3770
rect 7270 -3805 7310 -3800
rect 7270 -3840 7310 -3835
rect 7270 -3870 7275 -3840
rect 7275 -3870 7305 -3840
rect 7305 -3870 7310 -3840
rect 7270 -3875 7310 -3870
rect 7270 -3910 7310 -3905
rect 7270 -3940 7275 -3910
rect 7275 -3940 7305 -3910
rect 7305 -3940 7310 -3910
rect 7270 -3945 7310 -3940
rect 7270 -3980 7310 -3975
rect 7270 -4010 7275 -3980
rect 7275 -4010 7305 -3980
rect 7305 -4010 7310 -3980
rect 7270 -4015 7310 -4010
rect 7270 -4045 7310 -4040
rect 7270 -4075 7275 -4045
rect 7275 -4075 7305 -4045
rect 7305 -4075 7310 -4045
rect 7270 -4080 7310 -4075
rect 7270 -4105 7310 -4100
rect 7270 -4135 7275 -4105
rect 7275 -4135 7305 -4105
rect 7305 -4135 7310 -4105
rect 7270 -4140 7310 -4135
rect 7270 -4170 7310 -4165
rect 7270 -4200 7275 -4170
rect 7275 -4200 7305 -4170
rect 7305 -4200 7310 -4170
rect 7270 -4205 7310 -4200
rect 7270 -4240 7310 -4235
rect 7270 -4270 7275 -4240
rect 7275 -4270 7305 -4240
rect 7305 -4270 7310 -4240
rect 7270 -4275 7310 -4270
rect 7270 -4310 7310 -4305
rect 7270 -4340 7275 -4310
rect 7275 -4340 7305 -4310
rect 7305 -4340 7310 -4310
rect 7270 -4345 7310 -4340
rect 7270 -4380 7310 -4375
rect 7270 -4410 7275 -4380
rect 7275 -4410 7305 -4380
rect 7305 -4410 7310 -4380
rect 7270 -4415 7310 -4410
rect 7270 -4445 7310 -4440
rect 7270 -4475 7275 -4445
rect 7275 -4475 7305 -4445
rect 7305 -4475 7310 -4445
rect 7270 -4480 7310 -4475
rect 7620 -1305 7660 -1300
rect 7620 -1335 7625 -1305
rect 7625 -1335 7655 -1305
rect 7655 -1335 7660 -1305
rect 7620 -1340 7660 -1335
rect 7620 -1370 7660 -1365
rect 7620 -1400 7625 -1370
rect 7625 -1400 7655 -1370
rect 7655 -1400 7660 -1370
rect 7620 -1405 7660 -1400
rect 7620 -1440 7660 -1435
rect 7620 -1470 7625 -1440
rect 7625 -1470 7655 -1440
rect 7655 -1470 7660 -1440
rect 7620 -1475 7660 -1470
rect 7620 -1510 7660 -1505
rect 7620 -1540 7625 -1510
rect 7625 -1540 7655 -1510
rect 7655 -1540 7660 -1510
rect 7620 -1545 7660 -1540
rect 7620 -1580 7660 -1575
rect 7620 -1610 7625 -1580
rect 7625 -1610 7655 -1580
rect 7655 -1610 7660 -1580
rect 7620 -1615 7660 -1610
rect 7620 -1645 7660 -1640
rect 7620 -1675 7625 -1645
rect 7625 -1675 7655 -1645
rect 7655 -1675 7660 -1645
rect 7620 -1680 7660 -1675
rect 7620 -1705 7660 -1700
rect 7620 -1735 7625 -1705
rect 7625 -1735 7655 -1705
rect 7655 -1735 7660 -1705
rect 7620 -1740 7660 -1735
rect 7620 -1770 7660 -1765
rect 7620 -1800 7625 -1770
rect 7625 -1800 7655 -1770
rect 7655 -1800 7660 -1770
rect 7620 -1805 7660 -1800
rect 7620 -1840 7660 -1835
rect 7620 -1870 7625 -1840
rect 7625 -1870 7655 -1840
rect 7655 -1870 7660 -1840
rect 7620 -1875 7660 -1870
rect 7620 -1910 7660 -1905
rect 7620 -1940 7625 -1910
rect 7625 -1940 7655 -1910
rect 7655 -1940 7660 -1910
rect 7620 -1945 7660 -1940
rect 7620 -1980 7660 -1975
rect 7620 -2010 7625 -1980
rect 7625 -2010 7655 -1980
rect 7655 -2010 7660 -1980
rect 7620 -2015 7660 -2010
rect 7620 -2045 7660 -2040
rect 7620 -2075 7625 -2045
rect 7625 -2075 7655 -2045
rect 7655 -2075 7660 -2045
rect 7620 -2080 7660 -2075
rect 7620 -2105 7660 -2100
rect 7620 -2135 7625 -2105
rect 7625 -2135 7655 -2105
rect 7655 -2135 7660 -2105
rect 7620 -2140 7660 -2135
rect 7620 -2170 7660 -2165
rect 7620 -2200 7625 -2170
rect 7625 -2200 7655 -2170
rect 7655 -2200 7660 -2170
rect 7620 -2205 7660 -2200
rect 7620 -2240 7660 -2235
rect 7620 -2270 7625 -2240
rect 7625 -2270 7655 -2240
rect 7655 -2270 7660 -2240
rect 7620 -2275 7660 -2270
rect 7620 -2310 7660 -2305
rect 7620 -2340 7625 -2310
rect 7625 -2340 7655 -2310
rect 7655 -2340 7660 -2310
rect 7620 -2345 7660 -2340
rect 7620 -2380 7660 -2375
rect 7620 -2410 7625 -2380
rect 7625 -2410 7655 -2380
rect 7655 -2410 7660 -2380
rect 7620 -2415 7660 -2410
rect 7620 -2445 7660 -2440
rect 7620 -2475 7625 -2445
rect 7625 -2475 7655 -2445
rect 7655 -2475 7660 -2445
rect 7620 -2480 7660 -2475
rect 7620 -2505 7660 -2500
rect 7620 -2535 7625 -2505
rect 7625 -2535 7655 -2505
rect 7655 -2535 7660 -2505
rect 7620 -2540 7660 -2535
rect 7620 -2570 7660 -2565
rect 7620 -2600 7625 -2570
rect 7625 -2600 7655 -2570
rect 7655 -2600 7660 -2570
rect 7620 -2605 7660 -2600
rect 7620 -2640 7660 -2635
rect 7620 -2670 7625 -2640
rect 7625 -2670 7655 -2640
rect 7655 -2670 7660 -2640
rect 7620 -2675 7660 -2670
rect 7620 -2710 7660 -2705
rect 7620 -2740 7625 -2710
rect 7625 -2740 7655 -2710
rect 7655 -2740 7660 -2710
rect 7620 -2745 7660 -2740
rect 7620 -2780 7660 -2775
rect 7620 -2810 7625 -2780
rect 7625 -2810 7655 -2780
rect 7655 -2810 7660 -2780
rect 7620 -2815 7660 -2810
rect 7620 -2845 7660 -2840
rect 7620 -2875 7625 -2845
rect 7625 -2875 7655 -2845
rect 7655 -2875 7660 -2845
rect 7620 -2880 7660 -2875
rect 7620 -2905 7660 -2900
rect 7620 -2935 7625 -2905
rect 7625 -2935 7655 -2905
rect 7655 -2935 7660 -2905
rect 7620 -2940 7660 -2935
rect 7620 -2970 7660 -2965
rect 7620 -3000 7625 -2970
rect 7625 -3000 7655 -2970
rect 7655 -3000 7660 -2970
rect 7620 -3005 7660 -3000
rect 7620 -3040 7660 -3035
rect 7620 -3070 7625 -3040
rect 7625 -3070 7655 -3040
rect 7655 -3070 7660 -3040
rect 7620 -3075 7660 -3070
rect 7620 -3110 7660 -3105
rect 7620 -3140 7625 -3110
rect 7625 -3140 7655 -3110
rect 7655 -3140 7660 -3110
rect 7620 -3145 7660 -3140
rect 7620 -3180 7660 -3175
rect 7620 -3210 7625 -3180
rect 7625 -3210 7655 -3180
rect 7655 -3210 7660 -3180
rect 7620 -3215 7660 -3210
rect 7620 -3245 7660 -3240
rect 7620 -3275 7625 -3245
rect 7625 -3275 7655 -3245
rect 7655 -3275 7660 -3245
rect 7620 -3280 7660 -3275
rect 7620 -3305 7660 -3300
rect 7620 -3335 7625 -3305
rect 7625 -3335 7655 -3305
rect 7655 -3335 7660 -3305
rect 7620 -3340 7660 -3335
rect 7620 -3370 7660 -3365
rect 7620 -3400 7625 -3370
rect 7625 -3400 7655 -3370
rect 7655 -3400 7660 -3370
rect 7620 -3405 7660 -3400
rect 7620 -3440 7660 -3435
rect 7620 -3470 7625 -3440
rect 7625 -3470 7655 -3440
rect 7655 -3470 7660 -3440
rect 7620 -3475 7660 -3470
rect 7620 -3510 7660 -3505
rect 7620 -3540 7625 -3510
rect 7625 -3540 7655 -3510
rect 7655 -3540 7660 -3510
rect 7620 -3545 7660 -3540
rect 7620 -3580 7660 -3575
rect 7620 -3610 7625 -3580
rect 7625 -3610 7655 -3580
rect 7655 -3610 7660 -3580
rect 7620 -3615 7660 -3610
rect 7620 -3645 7660 -3640
rect 7620 -3675 7625 -3645
rect 7625 -3675 7655 -3645
rect 7655 -3675 7660 -3645
rect 7620 -3680 7660 -3675
rect 7620 -3705 7660 -3700
rect 7620 -3735 7625 -3705
rect 7625 -3735 7655 -3705
rect 7655 -3735 7660 -3705
rect 7620 -3740 7660 -3735
rect 7620 -3770 7660 -3765
rect 7620 -3800 7625 -3770
rect 7625 -3800 7655 -3770
rect 7655 -3800 7660 -3770
rect 7620 -3805 7660 -3800
rect 7620 -3840 7660 -3835
rect 7620 -3870 7625 -3840
rect 7625 -3870 7655 -3840
rect 7655 -3870 7660 -3840
rect 7620 -3875 7660 -3870
rect 7620 -3910 7660 -3905
rect 7620 -3940 7625 -3910
rect 7625 -3940 7655 -3910
rect 7655 -3940 7660 -3910
rect 7620 -3945 7660 -3940
rect 7620 -3980 7660 -3975
rect 7620 -4010 7625 -3980
rect 7625 -4010 7655 -3980
rect 7655 -4010 7660 -3980
rect 7620 -4015 7660 -4010
rect 7620 -4045 7660 -4040
rect 7620 -4075 7625 -4045
rect 7625 -4075 7655 -4045
rect 7655 -4075 7660 -4045
rect 7620 -4080 7660 -4075
rect 7620 -4105 7660 -4100
rect 7620 -4135 7625 -4105
rect 7625 -4135 7655 -4105
rect 7655 -4135 7660 -4105
rect 7620 -4140 7660 -4135
rect 7620 -4170 7660 -4165
rect 7620 -4200 7625 -4170
rect 7625 -4200 7655 -4170
rect 7655 -4200 7660 -4170
rect 7620 -4205 7660 -4200
rect 7620 -4240 7660 -4235
rect 7620 -4270 7625 -4240
rect 7625 -4270 7655 -4240
rect 7655 -4270 7660 -4240
rect 7620 -4275 7660 -4270
rect 7620 -4310 7660 -4305
rect 7620 -4340 7625 -4310
rect 7625 -4340 7655 -4310
rect 7655 -4340 7660 -4310
rect 7620 -4345 7660 -4340
rect 7620 -4380 7660 -4375
rect 7620 -4410 7625 -4380
rect 7625 -4410 7655 -4380
rect 7655 -4410 7660 -4380
rect 7620 -4415 7660 -4410
rect 7620 -4445 7660 -4440
rect 7620 -4475 7625 -4445
rect 7625 -4475 7655 -4445
rect 7655 -4475 7660 -4445
rect 7620 -4480 7660 -4475
rect 7970 -1305 8010 -1300
rect 7970 -1335 7975 -1305
rect 7975 -1335 8005 -1305
rect 8005 -1335 8010 -1305
rect 7970 -1340 8010 -1335
rect 7970 -1370 8010 -1365
rect 7970 -1400 7975 -1370
rect 7975 -1400 8005 -1370
rect 8005 -1400 8010 -1370
rect 7970 -1405 8010 -1400
rect 7970 -1440 8010 -1435
rect 7970 -1470 7975 -1440
rect 7975 -1470 8005 -1440
rect 8005 -1470 8010 -1440
rect 7970 -1475 8010 -1470
rect 7970 -1510 8010 -1505
rect 7970 -1540 7975 -1510
rect 7975 -1540 8005 -1510
rect 8005 -1540 8010 -1510
rect 7970 -1545 8010 -1540
rect 7970 -1580 8010 -1575
rect 7970 -1610 7975 -1580
rect 7975 -1610 8005 -1580
rect 8005 -1610 8010 -1580
rect 7970 -1615 8010 -1610
rect 7970 -1645 8010 -1640
rect 7970 -1675 7975 -1645
rect 7975 -1675 8005 -1645
rect 8005 -1675 8010 -1645
rect 7970 -1680 8010 -1675
rect 7970 -1705 8010 -1700
rect 7970 -1735 7975 -1705
rect 7975 -1735 8005 -1705
rect 8005 -1735 8010 -1705
rect 7970 -1740 8010 -1735
rect 7970 -1770 8010 -1765
rect 7970 -1800 7975 -1770
rect 7975 -1800 8005 -1770
rect 8005 -1800 8010 -1770
rect 7970 -1805 8010 -1800
rect 7970 -1840 8010 -1835
rect 7970 -1870 7975 -1840
rect 7975 -1870 8005 -1840
rect 8005 -1870 8010 -1840
rect 7970 -1875 8010 -1870
rect 7970 -1910 8010 -1905
rect 7970 -1940 7975 -1910
rect 7975 -1940 8005 -1910
rect 8005 -1940 8010 -1910
rect 7970 -1945 8010 -1940
rect 7970 -1980 8010 -1975
rect 7970 -2010 7975 -1980
rect 7975 -2010 8005 -1980
rect 8005 -2010 8010 -1980
rect 7970 -2015 8010 -2010
rect 7970 -2045 8010 -2040
rect 7970 -2075 7975 -2045
rect 7975 -2075 8005 -2045
rect 8005 -2075 8010 -2045
rect 7970 -2080 8010 -2075
rect 7970 -2105 8010 -2100
rect 7970 -2135 7975 -2105
rect 7975 -2135 8005 -2105
rect 8005 -2135 8010 -2105
rect 7970 -2140 8010 -2135
rect 7970 -2170 8010 -2165
rect 7970 -2200 7975 -2170
rect 7975 -2200 8005 -2170
rect 8005 -2200 8010 -2170
rect 7970 -2205 8010 -2200
rect 7970 -2240 8010 -2235
rect 7970 -2270 7975 -2240
rect 7975 -2270 8005 -2240
rect 8005 -2270 8010 -2240
rect 7970 -2275 8010 -2270
rect 7970 -2310 8010 -2305
rect 7970 -2340 7975 -2310
rect 7975 -2340 8005 -2310
rect 8005 -2340 8010 -2310
rect 7970 -2345 8010 -2340
rect 7970 -2380 8010 -2375
rect 7970 -2410 7975 -2380
rect 7975 -2410 8005 -2380
rect 8005 -2410 8010 -2380
rect 7970 -2415 8010 -2410
rect 7970 -2445 8010 -2440
rect 7970 -2475 7975 -2445
rect 7975 -2475 8005 -2445
rect 8005 -2475 8010 -2445
rect 7970 -2480 8010 -2475
rect 7970 -2505 8010 -2500
rect 7970 -2535 7975 -2505
rect 7975 -2535 8005 -2505
rect 8005 -2535 8010 -2505
rect 7970 -2540 8010 -2535
rect 7970 -2570 8010 -2565
rect 7970 -2600 7975 -2570
rect 7975 -2600 8005 -2570
rect 8005 -2600 8010 -2570
rect 7970 -2605 8010 -2600
rect 7970 -2640 8010 -2635
rect 7970 -2670 7975 -2640
rect 7975 -2670 8005 -2640
rect 8005 -2670 8010 -2640
rect 7970 -2675 8010 -2670
rect 7970 -2710 8010 -2705
rect 7970 -2740 7975 -2710
rect 7975 -2740 8005 -2710
rect 8005 -2740 8010 -2710
rect 7970 -2745 8010 -2740
rect 7970 -2780 8010 -2775
rect 7970 -2810 7975 -2780
rect 7975 -2810 8005 -2780
rect 8005 -2810 8010 -2780
rect 7970 -2815 8010 -2810
rect 7970 -2845 8010 -2840
rect 7970 -2875 7975 -2845
rect 7975 -2875 8005 -2845
rect 8005 -2875 8010 -2845
rect 7970 -2880 8010 -2875
rect 7970 -2905 8010 -2900
rect 7970 -2935 7975 -2905
rect 7975 -2935 8005 -2905
rect 8005 -2935 8010 -2905
rect 7970 -2940 8010 -2935
rect 7970 -2970 8010 -2965
rect 7970 -3000 7975 -2970
rect 7975 -3000 8005 -2970
rect 8005 -3000 8010 -2970
rect 7970 -3005 8010 -3000
rect 7970 -3040 8010 -3035
rect 7970 -3070 7975 -3040
rect 7975 -3070 8005 -3040
rect 8005 -3070 8010 -3040
rect 7970 -3075 8010 -3070
rect 7970 -3110 8010 -3105
rect 7970 -3140 7975 -3110
rect 7975 -3140 8005 -3110
rect 8005 -3140 8010 -3110
rect 7970 -3145 8010 -3140
rect 7970 -3180 8010 -3175
rect 7970 -3210 7975 -3180
rect 7975 -3210 8005 -3180
rect 8005 -3210 8010 -3180
rect 7970 -3215 8010 -3210
rect 7970 -3245 8010 -3240
rect 7970 -3275 7975 -3245
rect 7975 -3275 8005 -3245
rect 8005 -3275 8010 -3245
rect 7970 -3280 8010 -3275
rect 7970 -3305 8010 -3300
rect 7970 -3335 7975 -3305
rect 7975 -3335 8005 -3305
rect 8005 -3335 8010 -3305
rect 7970 -3340 8010 -3335
rect 7970 -3370 8010 -3365
rect 7970 -3400 7975 -3370
rect 7975 -3400 8005 -3370
rect 8005 -3400 8010 -3370
rect 7970 -3405 8010 -3400
rect 7970 -3440 8010 -3435
rect 7970 -3470 7975 -3440
rect 7975 -3470 8005 -3440
rect 8005 -3470 8010 -3440
rect 7970 -3475 8010 -3470
rect 7970 -3510 8010 -3505
rect 7970 -3540 7975 -3510
rect 7975 -3540 8005 -3510
rect 8005 -3540 8010 -3510
rect 7970 -3545 8010 -3540
rect 7970 -3580 8010 -3575
rect 7970 -3610 7975 -3580
rect 7975 -3610 8005 -3580
rect 8005 -3610 8010 -3580
rect 7970 -3615 8010 -3610
rect 7970 -3645 8010 -3640
rect 7970 -3675 7975 -3645
rect 7975 -3675 8005 -3645
rect 8005 -3675 8010 -3645
rect 7970 -3680 8010 -3675
rect 7970 -3705 8010 -3700
rect 7970 -3735 7975 -3705
rect 7975 -3735 8005 -3705
rect 8005 -3735 8010 -3705
rect 7970 -3740 8010 -3735
rect 7970 -3770 8010 -3765
rect 7970 -3800 7975 -3770
rect 7975 -3800 8005 -3770
rect 8005 -3800 8010 -3770
rect 7970 -3805 8010 -3800
rect 7970 -3840 8010 -3835
rect 7970 -3870 7975 -3840
rect 7975 -3870 8005 -3840
rect 8005 -3870 8010 -3840
rect 7970 -3875 8010 -3870
rect 7970 -3910 8010 -3905
rect 7970 -3940 7975 -3910
rect 7975 -3940 8005 -3910
rect 8005 -3940 8010 -3910
rect 7970 -3945 8010 -3940
rect 7970 -3980 8010 -3975
rect 7970 -4010 7975 -3980
rect 7975 -4010 8005 -3980
rect 8005 -4010 8010 -3980
rect 7970 -4015 8010 -4010
rect 7970 -4045 8010 -4040
rect 7970 -4075 7975 -4045
rect 7975 -4075 8005 -4045
rect 8005 -4075 8010 -4045
rect 7970 -4080 8010 -4075
rect 7970 -4105 8010 -4100
rect 7970 -4135 7975 -4105
rect 7975 -4135 8005 -4105
rect 8005 -4135 8010 -4105
rect 7970 -4140 8010 -4135
rect 7970 -4170 8010 -4165
rect 7970 -4200 7975 -4170
rect 7975 -4200 8005 -4170
rect 8005 -4200 8010 -4170
rect 7970 -4205 8010 -4200
rect 7970 -4240 8010 -4235
rect 7970 -4270 7975 -4240
rect 7975 -4270 8005 -4240
rect 8005 -4270 8010 -4240
rect 7970 -4275 8010 -4270
rect 7970 -4310 8010 -4305
rect 7970 -4340 7975 -4310
rect 7975 -4340 8005 -4310
rect 8005 -4340 8010 -4310
rect 7970 -4345 8010 -4340
rect 7970 -4380 8010 -4375
rect 7970 -4410 7975 -4380
rect 7975 -4410 8005 -4380
rect 8005 -4410 8010 -4380
rect 7970 -4415 8010 -4410
rect 7970 -4445 8010 -4440
rect 7970 -4475 7975 -4445
rect 7975 -4475 8005 -4445
rect 8005 -4475 8010 -4445
rect 7970 -4480 8010 -4475
rect 8320 -1305 8360 -1300
rect 8320 -1335 8325 -1305
rect 8325 -1335 8355 -1305
rect 8355 -1335 8360 -1305
rect 8320 -1340 8360 -1335
rect 8320 -1370 8360 -1365
rect 8320 -1400 8325 -1370
rect 8325 -1400 8355 -1370
rect 8355 -1400 8360 -1370
rect 8320 -1405 8360 -1400
rect 8320 -1440 8360 -1435
rect 8320 -1470 8325 -1440
rect 8325 -1470 8355 -1440
rect 8355 -1470 8360 -1440
rect 8320 -1475 8360 -1470
rect 8320 -1510 8360 -1505
rect 8320 -1540 8325 -1510
rect 8325 -1540 8355 -1510
rect 8355 -1540 8360 -1510
rect 8320 -1545 8360 -1540
rect 8320 -1580 8360 -1575
rect 8320 -1610 8325 -1580
rect 8325 -1610 8355 -1580
rect 8355 -1610 8360 -1580
rect 8320 -1615 8360 -1610
rect 8320 -1645 8360 -1640
rect 8320 -1675 8325 -1645
rect 8325 -1675 8355 -1645
rect 8355 -1675 8360 -1645
rect 8320 -1680 8360 -1675
rect 8320 -1705 8360 -1700
rect 8320 -1735 8325 -1705
rect 8325 -1735 8355 -1705
rect 8355 -1735 8360 -1705
rect 8320 -1740 8360 -1735
rect 8320 -1770 8360 -1765
rect 8320 -1800 8325 -1770
rect 8325 -1800 8355 -1770
rect 8355 -1800 8360 -1770
rect 8320 -1805 8360 -1800
rect 8320 -1840 8360 -1835
rect 8320 -1870 8325 -1840
rect 8325 -1870 8355 -1840
rect 8355 -1870 8360 -1840
rect 8320 -1875 8360 -1870
rect 8320 -1910 8360 -1905
rect 8320 -1940 8325 -1910
rect 8325 -1940 8355 -1910
rect 8355 -1940 8360 -1910
rect 8320 -1945 8360 -1940
rect 8320 -1980 8360 -1975
rect 8320 -2010 8325 -1980
rect 8325 -2010 8355 -1980
rect 8355 -2010 8360 -1980
rect 8320 -2015 8360 -2010
rect 8320 -2045 8360 -2040
rect 8320 -2075 8325 -2045
rect 8325 -2075 8355 -2045
rect 8355 -2075 8360 -2045
rect 8320 -2080 8360 -2075
rect 8320 -2105 8360 -2100
rect 8320 -2135 8325 -2105
rect 8325 -2135 8355 -2105
rect 8355 -2135 8360 -2105
rect 8320 -2140 8360 -2135
rect 8320 -2170 8360 -2165
rect 8320 -2200 8325 -2170
rect 8325 -2200 8355 -2170
rect 8355 -2200 8360 -2170
rect 8320 -2205 8360 -2200
rect 8320 -2240 8360 -2235
rect 8320 -2270 8325 -2240
rect 8325 -2270 8355 -2240
rect 8355 -2270 8360 -2240
rect 8320 -2275 8360 -2270
rect 8320 -2310 8360 -2305
rect 8320 -2340 8325 -2310
rect 8325 -2340 8355 -2310
rect 8355 -2340 8360 -2310
rect 8320 -2345 8360 -2340
rect 8320 -2380 8360 -2375
rect 8320 -2410 8325 -2380
rect 8325 -2410 8355 -2380
rect 8355 -2410 8360 -2380
rect 8320 -2415 8360 -2410
rect 8320 -2445 8360 -2440
rect 8320 -2475 8325 -2445
rect 8325 -2475 8355 -2445
rect 8355 -2475 8360 -2445
rect 8320 -2480 8360 -2475
rect 8320 -2505 8360 -2500
rect 8320 -2535 8325 -2505
rect 8325 -2535 8355 -2505
rect 8355 -2535 8360 -2505
rect 8320 -2540 8360 -2535
rect 8320 -2570 8360 -2565
rect 8320 -2600 8325 -2570
rect 8325 -2600 8355 -2570
rect 8355 -2600 8360 -2570
rect 8320 -2605 8360 -2600
rect 8320 -2640 8360 -2635
rect 8320 -2670 8325 -2640
rect 8325 -2670 8355 -2640
rect 8355 -2670 8360 -2640
rect 8320 -2675 8360 -2670
rect 8320 -2710 8360 -2705
rect 8320 -2740 8325 -2710
rect 8325 -2740 8355 -2710
rect 8355 -2740 8360 -2710
rect 8320 -2745 8360 -2740
rect 8320 -2780 8360 -2775
rect 8320 -2810 8325 -2780
rect 8325 -2810 8355 -2780
rect 8355 -2810 8360 -2780
rect 8320 -2815 8360 -2810
rect 8320 -2845 8360 -2840
rect 8320 -2875 8325 -2845
rect 8325 -2875 8355 -2845
rect 8355 -2875 8360 -2845
rect 8320 -2880 8360 -2875
rect 8320 -2905 8360 -2900
rect 8320 -2935 8325 -2905
rect 8325 -2935 8355 -2905
rect 8355 -2935 8360 -2905
rect 8320 -2940 8360 -2935
rect 8320 -2970 8360 -2965
rect 8320 -3000 8325 -2970
rect 8325 -3000 8355 -2970
rect 8355 -3000 8360 -2970
rect 8320 -3005 8360 -3000
rect 8320 -3040 8360 -3035
rect 8320 -3070 8325 -3040
rect 8325 -3070 8355 -3040
rect 8355 -3070 8360 -3040
rect 8320 -3075 8360 -3070
rect 8320 -3110 8360 -3105
rect 8320 -3140 8325 -3110
rect 8325 -3140 8355 -3110
rect 8355 -3140 8360 -3110
rect 8320 -3145 8360 -3140
rect 8320 -3180 8360 -3175
rect 8320 -3210 8325 -3180
rect 8325 -3210 8355 -3180
rect 8355 -3210 8360 -3180
rect 8320 -3215 8360 -3210
rect 8320 -3245 8360 -3240
rect 8320 -3275 8325 -3245
rect 8325 -3275 8355 -3245
rect 8355 -3275 8360 -3245
rect 8320 -3280 8360 -3275
rect 8320 -3305 8360 -3300
rect 8320 -3335 8325 -3305
rect 8325 -3335 8355 -3305
rect 8355 -3335 8360 -3305
rect 8320 -3340 8360 -3335
rect 8320 -3370 8360 -3365
rect 8320 -3400 8325 -3370
rect 8325 -3400 8355 -3370
rect 8355 -3400 8360 -3370
rect 8320 -3405 8360 -3400
rect 8320 -3440 8360 -3435
rect 8320 -3470 8325 -3440
rect 8325 -3470 8355 -3440
rect 8355 -3470 8360 -3440
rect 8320 -3475 8360 -3470
rect 8320 -3510 8360 -3505
rect 8320 -3540 8325 -3510
rect 8325 -3540 8355 -3510
rect 8355 -3540 8360 -3510
rect 8320 -3545 8360 -3540
rect 8320 -3580 8360 -3575
rect 8320 -3610 8325 -3580
rect 8325 -3610 8355 -3580
rect 8355 -3610 8360 -3580
rect 8320 -3615 8360 -3610
rect 8320 -3645 8360 -3640
rect 8320 -3675 8325 -3645
rect 8325 -3675 8355 -3645
rect 8355 -3675 8360 -3645
rect 8320 -3680 8360 -3675
rect 8320 -3705 8360 -3700
rect 8320 -3735 8325 -3705
rect 8325 -3735 8355 -3705
rect 8355 -3735 8360 -3705
rect 8320 -3740 8360 -3735
rect 8320 -3770 8360 -3765
rect 8320 -3800 8325 -3770
rect 8325 -3800 8355 -3770
rect 8355 -3800 8360 -3770
rect 8320 -3805 8360 -3800
rect 8320 -3840 8360 -3835
rect 8320 -3870 8325 -3840
rect 8325 -3870 8355 -3840
rect 8355 -3870 8360 -3840
rect 8320 -3875 8360 -3870
rect 8320 -3910 8360 -3905
rect 8320 -3940 8325 -3910
rect 8325 -3940 8355 -3910
rect 8355 -3940 8360 -3910
rect 8320 -3945 8360 -3940
rect 8320 -3980 8360 -3975
rect 8320 -4010 8325 -3980
rect 8325 -4010 8355 -3980
rect 8355 -4010 8360 -3980
rect 8320 -4015 8360 -4010
rect 8320 -4045 8360 -4040
rect 8320 -4075 8325 -4045
rect 8325 -4075 8355 -4045
rect 8355 -4075 8360 -4045
rect 8320 -4080 8360 -4075
rect 8320 -4105 8360 -4100
rect 8320 -4135 8325 -4105
rect 8325 -4135 8355 -4105
rect 8355 -4135 8360 -4105
rect 8320 -4140 8360 -4135
rect 8320 -4170 8360 -4165
rect 8320 -4200 8325 -4170
rect 8325 -4200 8355 -4170
rect 8355 -4200 8360 -4170
rect 8320 -4205 8360 -4200
rect 8320 -4240 8360 -4235
rect 8320 -4270 8325 -4240
rect 8325 -4270 8355 -4240
rect 8355 -4270 8360 -4240
rect 8320 -4275 8360 -4270
rect 8320 -4310 8360 -4305
rect 8320 -4340 8325 -4310
rect 8325 -4340 8355 -4310
rect 8355 -4340 8360 -4310
rect 8320 -4345 8360 -4340
rect 8320 -4380 8360 -4375
rect 8320 -4410 8325 -4380
rect 8325 -4410 8355 -4380
rect 8355 -4410 8360 -4380
rect 8320 -4415 8360 -4410
rect 8320 -4445 8360 -4440
rect 8320 -4475 8325 -4445
rect 8325 -4475 8355 -4445
rect 8355 -4475 8360 -4445
rect 8320 -4480 8360 -4475
rect 12925 -1375 12975 -1325
rect 13020 -1375 13070 -1325
rect 13115 -1375 13165 -1325
rect 13215 -1375 13265 -1325
rect 13315 -1375 13365 -1325
rect 13415 -1375 13465 -1325
rect 13510 -1375 13560 -1325
rect 13605 -1375 13655 -1325
rect 13725 -1375 13775 -1325
rect 13820 -1375 13870 -1325
rect 13915 -1375 13965 -1325
rect 14015 -1375 14065 -1325
rect 14115 -1375 14165 -1325
rect 14215 -1375 14265 -1325
rect 14310 -1375 14360 -1325
rect 14405 -1375 14455 -1325
rect 14525 -1375 14575 -1325
rect 14620 -1375 14670 -1325
rect 14715 -1375 14765 -1325
rect 14815 -1375 14865 -1325
rect 14915 -1375 14965 -1325
rect 15015 -1375 15065 -1325
rect 15110 -1375 15160 -1325
rect 15205 -1375 15255 -1325
rect 15325 -1375 15375 -1325
rect 15420 -1375 15470 -1325
rect 15515 -1375 15565 -1325
rect 15615 -1375 15665 -1325
rect 15715 -1375 15765 -1325
rect 15815 -1375 15865 -1325
rect 15910 -1375 15960 -1325
rect 16005 -1375 16055 -1325
rect 12925 -1465 12975 -1415
rect 13020 -1465 13070 -1415
rect 13115 -1465 13165 -1415
rect 13215 -1465 13265 -1415
rect 13315 -1465 13365 -1415
rect 13415 -1465 13465 -1415
rect 13510 -1465 13560 -1415
rect 13605 -1465 13655 -1415
rect 13725 -1465 13775 -1415
rect 13820 -1465 13870 -1415
rect 13915 -1465 13965 -1415
rect 14015 -1465 14065 -1415
rect 14115 -1465 14165 -1415
rect 14215 -1465 14265 -1415
rect 14310 -1465 14360 -1415
rect 14405 -1465 14455 -1415
rect 14525 -1465 14575 -1415
rect 14620 -1465 14670 -1415
rect 14715 -1465 14765 -1415
rect 14815 -1465 14865 -1415
rect 14915 -1465 14965 -1415
rect 15015 -1465 15065 -1415
rect 15110 -1465 15160 -1415
rect 15205 -1465 15255 -1415
rect 15325 -1465 15375 -1415
rect 15420 -1465 15470 -1415
rect 15515 -1465 15565 -1415
rect 15615 -1465 15665 -1415
rect 15715 -1465 15765 -1415
rect 15815 -1465 15865 -1415
rect 15910 -1465 15960 -1415
rect 16005 -1465 16055 -1415
rect 12925 -1565 12975 -1515
rect 13020 -1565 13070 -1515
rect 13115 -1565 13165 -1515
rect 13215 -1565 13265 -1515
rect 13315 -1565 13365 -1515
rect 13415 -1565 13465 -1515
rect 13510 -1565 13560 -1515
rect 13605 -1565 13655 -1515
rect 13725 -1565 13775 -1515
rect 13820 -1565 13870 -1515
rect 13915 -1565 13965 -1515
rect 14015 -1565 14065 -1515
rect 14115 -1565 14165 -1515
rect 14215 -1565 14265 -1515
rect 14310 -1565 14360 -1515
rect 14405 -1565 14455 -1515
rect 14525 -1565 14575 -1515
rect 14620 -1565 14670 -1515
rect 14715 -1565 14765 -1515
rect 14815 -1565 14865 -1515
rect 14915 -1565 14965 -1515
rect 15015 -1565 15065 -1515
rect 15110 -1565 15160 -1515
rect 15205 -1565 15255 -1515
rect 15325 -1565 15375 -1515
rect 15420 -1565 15470 -1515
rect 15515 -1565 15565 -1515
rect 15615 -1565 15665 -1515
rect 15715 -1565 15765 -1515
rect 15815 -1565 15865 -1515
rect 15910 -1565 15960 -1515
rect 16005 -1565 16055 -1515
rect 12925 -1655 12975 -1605
rect 13020 -1655 13070 -1605
rect 13115 -1655 13165 -1605
rect 13215 -1655 13265 -1605
rect 13315 -1655 13365 -1605
rect 13415 -1655 13465 -1605
rect 13510 -1655 13560 -1605
rect 13605 -1655 13655 -1605
rect 13725 -1655 13775 -1605
rect 13820 -1655 13870 -1605
rect 13915 -1655 13965 -1605
rect 14015 -1655 14065 -1605
rect 14115 -1655 14165 -1605
rect 14215 -1655 14265 -1605
rect 14310 -1655 14360 -1605
rect 14405 -1655 14455 -1605
rect 14525 -1655 14575 -1605
rect 14620 -1655 14670 -1605
rect 14715 -1655 14765 -1605
rect 14815 -1655 14865 -1605
rect 14915 -1655 14965 -1605
rect 15015 -1655 15065 -1605
rect 15110 -1655 15160 -1605
rect 15205 -1655 15255 -1605
rect 15325 -1655 15375 -1605
rect 15420 -1655 15470 -1605
rect 15515 -1655 15565 -1605
rect 15615 -1655 15665 -1605
rect 15715 -1655 15765 -1605
rect 15815 -1655 15865 -1605
rect 15910 -1655 15960 -1605
rect 16005 -1655 16055 -1605
rect 12925 -1775 12975 -1725
rect 13020 -1775 13070 -1725
rect 13115 -1775 13165 -1725
rect 13215 -1775 13265 -1725
rect 13315 -1775 13365 -1725
rect 13415 -1775 13465 -1725
rect 13510 -1775 13560 -1725
rect 13605 -1775 13655 -1725
rect 13725 -1775 13775 -1725
rect 13820 -1775 13870 -1725
rect 13915 -1775 13965 -1725
rect 14015 -1775 14065 -1725
rect 14115 -1775 14165 -1725
rect 14215 -1775 14265 -1725
rect 14310 -1775 14360 -1725
rect 14405 -1775 14455 -1725
rect 14525 -1775 14575 -1725
rect 14620 -1775 14670 -1725
rect 14715 -1775 14765 -1725
rect 14815 -1775 14865 -1725
rect 14915 -1775 14965 -1725
rect 15015 -1775 15065 -1725
rect 15110 -1775 15160 -1725
rect 15205 -1775 15255 -1725
rect 15325 -1775 15375 -1725
rect 15420 -1775 15470 -1725
rect 15515 -1775 15565 -1725
rect 15615 -1775 15665 -1725
rect 15715 -1775 15765 -1725
rect 15815 -1775 15865 -1725
rect 15910 -1775 15960 -1725
rect 16005 -1775 16055 -1725
rect 12925 -1865 12975 -1815
rect 13020 -1865 13070 -1815
rect 13115 -1865 13165 -1815
rect 13215 -1865 13265 -1815
rect 13315 -1865 13365 -1815
rect 13415 -1865 13465 -1815
rect 13510 -1865 13560 -1815
rect 13605 -1865 13655 -1815
rect 13725 -1865 13775 -1815
rect 13820 -1865 13870 -1815
rect 13915 -1865 13965 -1815
rect 14015 -1865 14065 -1815
rect 14115 -1865 14165 -1815
rect 14215 -1865 14265 -1815
rect 14310 -1865 14360 -1815
rect 14405 -1865 14455 -1815
rect 14525 -1865 14575 -1815
rect 14620 -1865 14670 -1815
rect 14715 -1865 14765 -1815
rect 14815 -1865 14865 -1815
rect 14915 -1865 14965 -1815
rect 15015 -1865 15065 -1815
rect 15110 -1865 15160 -1815
rect 15205 -1865 15255 -1815
rect 15325 -1865 15375 -1815
rect 15420 -1865 15470 -1815
rect 15515 -1865 15565 -1815
rect 15615 -1865 15665 -1815
rect 15715 -1865 15765 -1815
rect 15815 -1865 15865 -1815
rect 15910 -1865 15960 -1815
rect 16005 -1865 16055 -1815
rect 12925 -1965 12975 -1915
rect 13020 -1965 13070 -1915
rect 13115 -1965 13165 -1915
rect 13215 -1965 13265 -1915
rect 13315 -1965 13365 -1915
rect 13415 -1965 13465 -1915
rect 13510 -1965 13560 -1915
rect 13605 -1965 13655 -1915
rect 13725 -1965 13775 -1915
rect 13820 -1965 13870 -1915
rect 13915 -1965 13965 -1915
rect 14015 -1965 14065 -1915
rect 14115 -1965 14165 -1915
rect 14215 -1965 14265 -1915
rect 14310 -1965 14360 -1915
rect 14405 -1965 14455 -1915
rect 14525 -1965 14575 -1915
rect 14620 -1965 14670 -1915
rect 14715 -1965 14765 -1915
rect 14815 -1965 14865 -1915
rect 14915 -1965 14965 -1915
rect 15015 -1965 15065 -1915
rect 15110 -1965 15160 -1915
rect 15205 -1965 15255 -1915
rect 15325 -1965 15375 -1915
rect 15420 -1965 15470 -1915
rect 15515 -1965 15565 -1915
rect 15615 -1965 15665 -1915
rect 15715 -1965 15765 -1915
rect 15815 -1965 15865 -1915
rect 15910 -1965 15960 -1915
rect 16005 -1965 16055 -1915
rect 12925 -2055 12975 -2005
rect 13020 -2055 13070 -2005
rect 13115 -2055 13165 -2005
rect 13215 -2055 13265 -2005
rect 13315 -2055 13365 -2005
rect 13415 -2055 13465 -2005
rect 13510 -2055 13560 -2005
rect 13605 -2055 13655 -2005
rect 13725 -2055 13775 -2005
rect 13820 -2055 13870 -2005
rect 13915 -2055 13965 -2005
rect 14015 -2055 14065 -2005
rect 14115 -2055 14165 -2005
rect 14215 -2055 14265 -2005
rect 14310 -2055 14360 -2005
rect 14405 -2055 14455 -2005
rect 14525 -2055 14575 -2005
rect 14620 -2055 14670 -2005
rect 14715 -2055 14765 -2005
rect 14815 -2055 14865 -2005
rect 14915 -2055 14965 -2005
rect 15015 -2055 15065 -2005
rect 15110 -2055 15160 -2005
rect 15205 -2055 15255 -2005
rect 15325 -2055 15375 -2005
rect 15420 -2055 15470 -2005
rect 15515 -2055 15565 -2005
rect 15615 -2055 15665 -2005
rect 15715 -2055 15765 -2005
rect 15815 -2055 15865 -2005
rect 15910 -2055 15960 -2005
rect 16005 -2055 16055 -2005
rect 12925 -2175 12975 -2125
rect 13020 -2175 13070 -2125
rect 13115 -2175 13165 -2125
rect 13215 -2175 13265 -2125
rect 13315 -2175 13365 -2125
rect 13415 -2175 13465 -2125
rect 13510 -2175 13560 -2125
rect 13605 -2175 13655 -2125
rect 13725 -2175 13775 -2125
rect 13820 -2175 13870 -2125
rect 13915 -2175 13965 -2125
rect 14015 -2175 14065 -2125
rect 14115 -2175 14165 -2125
rect 14215 -2175 14265 -2125
rect 14310 -2175 14360 -2125
rect 14405 -2175 14455 -2125
rect 14525 -2175 14575 -2125
rect 14620 -2175 14670 -2125
rect 14715 -2175 14765 -2125
rect 14815 -2175 14865 -2125
rect 14915 -2175 14965 -2125
rect 15015 -2175 15065 -2125
rect 15110 -2175 15160 -2125
rect 15205 -2175 15255 -2125
rect 15325 -2175 15375 -2125
rect 15420 -2175 15470 -2125
rect 15515 -2175 15565 -2125
rect 15615 -2175 15665 -2125
rect 15715 -2175 15765 -2125
rect 15815 -2175 15865 -2125
rect 15910 -2175 15960 -2125
rect 16005 -2175 16055 -2125
rect 12925 -2265 12975 -2215
rect 13020 -2265 13070 -2215
rect 13115 -2265 13165 -2215
rect 13215 -2265 13265 -2215
rect 13315 -2265 13365 -2215
rect 13415 -2265 13465 -2215
rect 13510 -2265 13560 -2215
rect 13605 -2265 13655 -2215
rect 13725 -2265 13775 -2215
rect 13820 -2265 13870 -2215
rect 13915 -2265 13965 -2215
rect 14015 -2265 14065 -2215
rect 14115 -2265 14165 -2215
rect 14215 -2265 14265 -2215
rect 14310 -2265 14360 -2215
rect 14405 -2265 14455 -2215
rect 14525 -2265 14575 -2215
rect 14620 -2265 14670 -2215
rect 14715 -2265 14765 -2215
rect 14815 -2265 14865 -2215
rect 14915 -2265 14965 -2215
rect 15015 -2265 15065 -2215
rect 15110 -2265 15160 -2215
rect 15205 -2265 15255 -2215
rect 15325 -2265 15375 -2215
rect 15420 -2265 15470 -2215
rect 15515 -2265 15565 -2215
rect 15615 -2265 15665 -2215
rect 15715 -2265 15765 -2215
rect 15815 -2265 15865 -2215
rect 15910 -2265 15960 -2215
rect 16005 -2265 16055 -2215
rect 12925 -2365 12975 -2315
rect 13020 -2365 13070 -2315
rect 13115 -2365 13165 -2315
rect 13215 -2365 13265 -2315
rect 13315 -2365 13365 -2315
rect 13415 -2365 13465 -2315
rect 13510 -2365 13560 -2315
rect 13605 -2365 13655 -2315
rect 13725 -2365 13775 -2315
rect 13820 -2365 13870 -2315
rect 13915 -2365 13965 -2315
rect 14015 -2365 14065 -2315
rect 14115 -2365 14165 -2315
rect 14215 -2365 14265 -2315
rect 14310 -2365 14360 -2315
rect 14405 -2365 14455 -2315
rect 14525 -2365 14575 -2315
rect 14620 -2365 14670 -2315
rect 14715 -2365 14765 -2315
rect 14815 -2365 14865 -2315
rect 14915 -2365 14965 -2315
rect 15015 -2365 15065 -2315
rect 15110 -2365 15160 -2315
rect 15205 -2365 15255 -2315
rect 15325 -2365 15375 -2315
rect 15420 -2365 15470 -2315
rect 15515 -2365 15565 -2315
rect 15615 -2365 15665 -2315
rect 15715 -2365 15765 -2315
rect 15815 -2365 15865 -2315
rect 15910 -2365 15960 -2315
rect 16005 -2365 16055 -2315
rect 12925 -2455 12975 -2405
rect 13020 -2455 13070 -2405
rect 13115 -2455 13165 -2405
rect 13215 -2455 13265 -2405
rect 13315 -2455 13365 -2405
rect 13415 -2455 13465 -2405
rect 13510 -2455 13560 -2405
rect 13605 -2455 13655 -2405
rect 13725 -2455 13775 -2405
rect 13820 -2455 13870 -2405
rect 13915 -2455 13965 -2405
rect 14015 -2455 14065 -2405
rect 14115 -2455 14165 -2405
rect 14215 -2455 14265 -2405
rect 14310 -2455 14360 -2405
rect 14405 -2455 14455 -2405
rect 14525 -2455 14575 -2405
rect 14620 -2455 14670 -2405
rect 14715 -2455 14765 -2405
rect 14815 -2455 14865 -2405
rect 14915 -2455 14965 -2405
rect 15015 -2455 15065 -2405
rect 15110 -2455 15160 -2405
rect 15205 -2455 15255 -2405
rect 15325 -2455 15375 -2405
rect 15420 -2455 15470 -2405
rect 15515 -2455 15565 -2405
rect 15615 -2455 15665 -2405
rect 15715 -2455 15765 -2405
rect 15815 -2455 15865 -2405
rect 15910 -2455 15960 -2405
rect 16005 -2455 16055 -2405
rect 12925 -2575 12975 -2525
rect 13020 -2575 13070 -2525
rect 13115 -2575 13165 -2525
rect 13215 -2575 13265 -2525
rect 13315 -2575 13365 -2525
rect 13415 -2575 13465 -2525
rect 13510 -2575 13560 -2525
rect 13605 -2575 13655 -2525
rect 13725 -2575 13775 -2525
rect 13820 -2575 13870 -2525
rect 13915 -2575 13965 -2525
rect 14015 -2575 14065 -2525
rect 14115 -2575 14165 -2525
rect 14215 -2575 14265 -2525
rect 14310 -2575 14360 -2525
rect 14405 -2575 14455 -2525
rect 14525 -2575 14575 -2525
rect 14620 -2575 14670 -2525
rect 14715 -2575 14765 -2525
rect 14815 -2575 14865 -2525
rect 14915 -2575 14965 -2525
rect 15015 -2575 15065 -2525
rect 15110 -2575 15160 -2525
rect 15205 -2575 15255 -2525
rect 15325 -2575 15375 -2525
rect 15420 -2575 15470 -2525
rect 15515 -2575 15565 -2525
rect 15615 -2575 15665 -2525
rect 15715 -2575 15765 -2525
rect 15815 -2575 15865 -2525
rect 15910 -2575 15960 -2525
rect 16005 -2575 16055 -2525
rect 12925 -2665 12975 -2615
rect 13020 -2665 13070 -2615
rect 13115 -2665 13165 -2615
rect 13215 -2665 13265 -2615
rect 13315 -2665 13365 -2615
rect 13415 -2665 13465 -2615
rect 13510 -2665 13560 -2615
rect 13605 -2665 13655 -2615
rect 13725 -2665 13775 -2615
rect 13820 -2665 13870 -2615
rect 13915 -2665 13965 -2615
rect 14015 -2665 14065 -2615
rect 14115 -2665 14165 -2615
rect 14215 -2665 14265 -2615
rect 14310 -2665 14360 -2615
rect 14405 -2665 14455 -2615
rect 14525 -2665 14575 -2615
rect 14620 -2665 14670 -2615
rect 14715 -2665 14765 -2615
rect 14815 -2665 14865 -2615
rect 14915 -2665 14965 -2615
rect 15015 -2665 15065 -2615
rect 15110 -2665 15160 -2615
rect 15205 -2665 15255 -2615
rect 15325 -2665 15375 -2615
rect 15420 -2665 15470 -2615
rect 15515 -2665 15565 -2615
rect 15615 -2665 15665 -2615
rect 15715 -2665 15765 -2615
rect 15815 -2665 15865 -2615
rect 15910 -2665 15960 -2615
rect 16005 -2665 16055 -2615
rect 12925 -2765 12975 -2715
rect 13020 -2765 13070 -2715
rect 13115 -2765 13165 -2715
rect 13215 -2765 13265 -2715
rect 13315 -2765 13365 -2715
rect 13415 -2765 13465 -2715
rect 13510 -2765 13560 -2715
rect 13605 -2765 13655 -2715
rect 13725 -2765 13775 -2715
rect 13820 -2765 13870 -2715
rect 13915 -2765 13965 -2715
rect 14015 -2765 14065 -2715
rect 14115 -2765 14165 -2715
rect 14215 -2765 14265 -2715
rect 14310 -2765 14360 -2715
rect 14405 -2765 14455 -2715
rect 14525 -2765 14575 -2715
rect 14620 -2765 14670 -2715
rect 14715 -2765 14765 -2715
rect 14815 -2765 14865 -2715
rect 14915 -2765 14965 -2715
rect 15015 -2765 15065 -2715
rect 15110 -2765 15160 -2715
rect 15205 -2765 15255 -2715
rect 15325 -2765 15375 -2715
rect 15420 -2765 15470 -2715
rect 15515 -2765 15565 -2715
rect 15615 -2765 15665 -2715
rect 15715 -2765 15765 -2715
rect 15815 -2765 15865 -2715
rect 15910 -2765 15960 -2715
rect 16005 -2765 16055 -2715
rect 12925 -2855 12975 -2805
rect 13020 -2855 13070 -2805
rect 13115 -2855 13165 -2805
rect 13215 -2855 13265 -2805
rect 13315 -2855 13365 -2805
rect 13415 -2855 13465 -2805
rect 13510 -2855 13560 -2805
rect 13605 -2855 13655 -2805
rect 13725 -2855 13775 -2805
rect 13820 -2855 13870 -2805
rect 13915 -2855 13965 -2805
rect 14015 -2855 14065 -2805
rect 14115 -2855 14165 -2805
rect 14215 -2855 14265 -2805
rect 14310 -2855 14360 -2805
rect 14405 -2855 14455 -2805
rect 14525 -2855 14575 -2805
rect 14620 -2855 14670 -2805
rect 14715 -2855 14765 -2805
rect 14815 -2855 14865 -2805
rect 14915 -2855 14965 -2805
rect 15015 -2855 15065 -2805
rect 15110 -2855 15160 -2805
rect 15205 -2855 15255 -2805
rect 15325 -2855 15375 -2805
rect 15420 -2855 15470 -2805
rect 15515 -2855 15565 -2805
rect 15615 -2855 15665 -2805
rect 15715 -2855 15765 -2805
rect 15815 -2855 15865 -2805
rect 15910 -2855 15960 -2805
rect 16005 -2855 16055 -2805
rect 12925 -2975 12975 -2925
rect 13020 -2975 13070 -2925
rect 13115 -2975 13165 -2925
rect 13215 -2975 13265 -2925
rect 13315 -2975 13365 -2925
rect 13415 -2975 13465 -2925
rect 13510 -2975 13560 -2925
rect 13605 -2975 13655 -2925
rect 13725 -2975 13775 -2925
rect 13820 -2975 13870 -2925
rect 13915 -2975 13965 -2925
rect 14015 -2975 14065 -2925
rect 14115 -2975 14165 -2925
rect 14215 -2975 14265 -2925
rect 14310 -2975 14360 -2925
rect 14405 -2975 14455 -2925
rect 14525 -2975 14575 -2925
rect 14620 -2975 14670 -2925
rect 14715 -2975 14765 -2925
rect 14815 -2975 14865 -2925
rect 14915 -2975 14965 -2925
rect 15015 -2975 15065 -2925
rect 15110 -2975 15160 -2925
rect 15205 -2975 15255 -2925
rect 15325 -2975 15375 -2925
rect 15420 -2975 15470 -2925
rect 15515 -2975 15565 -2925
rect 15615 -2975 15665 -2925
rect 15715 -2975 15765 -2925
rect 15815 -2975 15865 -2925
rect 15910 -2975 15960 -2925
rect 16005 -2975 16055 -2925
rect 12925 -3065 12975 -3015
rect 13020 -3065 13070 -3015
rect 13115 -3065 13165 -3015
rect 13215 -3065 13265 -3015
rect 13315 -3065 13365 -3015
rect 13415 -3065 13465 -3015
rect 13510 -3065 13560 -3015
rect 13605 -3065 13655 -3015
rect 13725 -3065 13775 -3015
rect 13820 -3065 13870 -3015
rect 13915 -3065 13965 -3015
rect 14015 -3065 14065 -3015
rect 14115 -3065 14165 -3015
rect 14215 -3065 14265 -3015
rect 14310 -3065 14360 -3015
rect 14405 -3065 14455 -3015
rect 14525 -3065 14575 -3015
rect 14620 -3065 14670 -3015
rect 14715 -3065 14765 -3015
rect 14815 -3065 14865 -3015
rect 14915 -3065 14965 -3015
rect 15015 -3065 15065 -3015
rect 15110 -3065 15160 -3015
rect 15205 -3065 15255 -3015
rect 15325 -3065 15375 -3015
rect 15420 -3065 15470 -3015
rect 15515 -3065 15565 -3015
rect 15615 -3065 15665 -3015
rect 15715 -3065 15765 -3015
rect 15815 -3065 15865 -3015
rect 15910 -3065 15960 -3015
rect 16005 -3065 16055 -3015
rect 12925 -3165 12975 -3115
rect 13020 -3165 13070 -3115
rect 13115 -3165 13165 -3115
rect 13215 -3165 13265 -3115
rect 13315 -3165 13365 -3115
rect 13415 -3165 13465 -3115
rect 13510 -3165 13560 -3115
rect 13605 -3165 13655 -3115
rect 13725 -3165 13775 -3115
rect 13820 -3165 13870 -3115
rect 13915 -3165 13965 -3115
rect 14015 -3165 14065 -3115
rect 14115 -3165 14165 -3115
rect 14215 -3165 14265 -3115
rect 14310 -3165 14360 -3115
rect 14405 -3165 14455 -3115
rect 14525 -3165 14575 -3115
rect 14620 -3165 14670 -3115
rect 14715 -3165 14765 -3115
rect 14815 -3165 14865 -3115
rect 14915 -3165 14965 -3115
rect 15015 -3165 15065 -3115
rect 15110 -3165 15160 -3115
rect 15205 -3165 15255 -3115
rect 15325 -3165 15375 -3115
rect 15420 -3165 15470 -3115
rect 15515 -3165 15565 -3115
rect 15615 -3165 15665 -3115
rect 15715 -3165 15765 -3115
rect 15815 -3165 15865 -3115
rect 15910 -3165 15960 -3115
rect 16005 -3165 16055 -3115
rect 12925 -3255 12975 -3205
rect 13020 -3255 13070 -3205
rect 13115 -3255 13165 -3205
rect 13215 -3255 13265 -3205
rect 13315 -3255 13365 -3205
rect 13415 -3255 13465 -3205
rect 13510 -3255 13560 -3205
rect 13605 -3255 13655 -3205
rect 13725 -3255 13775 -3205
rect 13820 -3255 13870 -3205
rect 13915 -3255 13965 -3205
rect 14015 -3255 14065 -3205
rect 14115 -3255 14165 -3205
rect 14215 -3255 14265 -3205
rect 14310 -3255 14360 -3205
rect 14405 -3255 14455 -3205
rect 14525 -3255 14575 -3205
rect 14620 -3255 14670 -3205
rect 14715 -3255 14765 -3205
rect 14815 -3255 14865 -3205
rect 14915 -3255 14965 -3205
rect 15015 -3255 15065 -3205
rect 15110 -3255 15160 -3205
rect 15205 -3255 15255 -3205
rect 15325 -3255 15375 -3205
rect 15420 -3255 15470 -3205
rect 15515 -3255 15565 -3205
rect 15615 -3255 15665 -3205
rect 15715 -3255 15765 -3205
rect 15815 -3255 15865 -3205
rect 15910 -3255 15960 -3205
rect 16005 -3255 16055 -3205
rect 12925 -3375 12975 -3325
rect 13020 -3375 13070 -3325
rect 13115 -3375 13165 -3325
rect 13215 -3375 13265 -3325
rect 13315 -3375 13365 -3325
rect 13415 -3375 13465 -3325
rect 13510 -3375 13560 -3325
rect 13605 -3375 13655 -3325
rect 13725 -3375 13775 -3325
rect 13820 -3375 13870 -3325
rect 13915 -3375 13965 -3325
rect 14015 -3375 14065 -3325
rect 14115 -3375 14165 -3325
rect 14215 -3375 14265 -3325
rect 14310 -3375 14360 -3325
rect 14405 -3375 14455 -3325
rect 14525 -3375 14575 -3325
rect 14620 -3375 14670 -3325
rect 14715 -3375 14765 -3325
rect 14815 -3375 14865 -3325
rect 14915 -3375 14965 -3325
rect 15015 -3375 15065 -3325
rect 15110 -3375 15160 -3325
rect 15205 -3375 15255 -3325
rect 15325 -3375 15375 -3325
rect 15420 -3375 15470 -3325
rect 15515 -3375 15565 -3325
rect 15615 -3375 15665 -3325
rect 15715 -3375 15765 -3325
rect 15815 -3375 15865 -3325
rect 15910 -3375 15960 -3325
rect 16005 -3375 16055 -3325
rect 12925 -3465 12975 -3415
rect 13020 -3465 13070 -3415
rect 13115 -3465 13165 -3415
rect 13215 -3465 13265 -3415
rect 13315 -3465 13365 -3415
rect 13415 -3465 13465 -3415
rect 13510 -3465 13560 -3415
rect 13605 -3465 13655 -3415
rect 13725 -3465 13775 -3415
rect 13820 -3465 13870 -3415
rect 13915 -3465 13965 -3415
rect 14015 -3465 14065 -3415
rect 14115 -3465 14165 -3415
rect 14215 -3465 14265 -3415
rect 14310 -3465 14360 -3415
rect 14405 -3465 14455 -3415
rect 14525 -3465 14575 -3415
rect 14620 -3465 14670 -3415
rect 14715 -3465 14765 -3415
rect 14815 -3465 14865 -3415
rect 14915 -3465 14965 -3415
rect 15015 -3465 15065 -3415
rect 15110 -3465 15160 -3415
rect 15205 -3465 15255 -3415
rect 15325 -3465 15375 -3415
rect 15420 -3465 15470 -3415
rect 15515 -3465 15565 -3415
rect 15615 -3465 15665 -3415
rect 15715 -3465 15765 -3415
rect 15815 -3465 15865 -3415
rect 15910 -3465 15960 -3415
rect 16005 -3465 16055 -3415
rect 12925 -3565 12975 -3515
rect 13020 -3565 13070 -3515
rect 13115 -3565 13165 -3515
rect 13215 -3565 13265 -3515
rect 13315 -3565 13365 -3515
rect 13415 -3565 13465 -3515
rect 13510 -3565 13560 -3515
rect 13605 -3565 13655 -3515
rect 13725 -3565 13775 -3515
rect 13820 -3565 13870 -3515
rect 13915 -3565 13965 -3515
rect 14015 -3565 14065 -3515
rect 14115 -3565 14165 -3515
rect 14215 -3565 14265 -3515
rect 14310 -3565 14360 -3515
rect 14405 -3565 14455 -3515
rect 14525 -3565 14575 -3515
rect 14620 -3565 14670 -3515
rect 14715 -3565 14765 -3515
rect 14815 -3565 14865 -3515
rect 14915 -3565 14965 -3515
rect 15015 -3565 15065 -3515
rect 15110 -3565 15160 -3515
rect 15205 -3565 15255 -3515
rect 15325 -3565 15375 -3515
rect 15420 -3565 15470 -3515
rect 15515 -3565 15565 -3515
rect 15615 -3565 15665 -3515
rect 15715 -3565 15765 -3515
rect 15815 -3565 15865 -3515
rect 15910 -3565 15960 -3515
rect 16005 -3565 16055 -3515
rect 12925 -3655 12975 -3605
rect 13020 -3655 13070 -3605
rect 13115 -3655 13165 -3605
rect 13215 -3655 13265 -3605
rect 13315 -3655 13365 -3605
rect 13415 -3655 13465 -3605
rect 13510 -3655 13560 -3605
rect 13605 -3655 13655 -3605
rect 13725 -3655 13775 -3605
rect 13820 -3655 13870 -3605
rect 13915 -3655 13965 -3605
rect 14015 -3655 14065 -3605
rect 14115 -3655 14165 -3605
rect 14215 -3655 14265 -3605
rect 14310 -3655 14360 -3605
rect 14405 -3655 14455 -3605
rect 14525 -3655 14575 -3605
rect 14620 -3655 14670 -3605
rect 14715 -3655 14765 -3605
rect 14815 -3655 14865 -3605
rect 14915 -3655 14965 -3605
rect 15015 -3655 15065 -3605
rect 15110 -3655 15160 -3605
rect 15205 -3655 15255 -3605
rect 15325 -3655 15375 -3605
rect 15420 -3655 15470 -3605
rect 15515 -3655 15565 -3605
rect 15615 -3655 15665 -3605
rect 15715 -3655 15765 -3605
rect 15815 -3655 15865 -3605
rect 15910 -3655 15960 -3605
rect 16005 -3655 16055 -3605
rect 12925 -3775 12975 -3725
rect 13020 -3775 13070 -3725
rect 13115 -3775 13165 -3725
rect 13215 -3775 13265 -3725
rect 13315 -3775 13365 -3725
rect 13415 -3775 13465 -3725
rect 13510 -3775 13560 -3725
rect 13605 -3775 13655 -3725
rect 13725 -3775 13775 -3725
rect 13820 -3775 13870 -3725
rect 13915 -3775 13965 -3725
rect 14015 -3775 14065 -3725
rect 14115 -3775 14165 -3725
rect 14215 -3775 14265 -3725
rect 14310 -3775 14360 -3725
rect 14405 -3775 14455 -3725
rect 14525 -3775 14575 -3725
rect 14620 -3775 14670 -3725
rect 14715 -3775 14765 -3725
rect 14815 -3775 14865 -3725
rect 14915 -3775 14965 -3725
rect 15015 -3775 15065 -3725
rect 15110 -3775 15160 -3725
rect 15205 -3775 15255 -3725
rect 15325 -3775 15375 -3725
rect 15420 -3775 15470 -3725
rect 15515 -3775 15565 -3725
rect 15615 -3775 15665 -3725
rect 15715 -3775 15765 -3725
rect 15815 -3775 15865 -3725
rect 15910 -3775 15960 -3725
rect 16005 -3775 16055 -3725
rect 12925 -3865 12975 -3815
rect 13020 -3865 13070 -3815
rect 13115 -3865 13165 -3815
rect 13215 -3865 13265 -3815
rect 13315 -3865 13365 -3815
rect 13415 -3865 13465 -3815
rect 13510 -3865 13560 -3815
rect 13605 -3865 13655 -3815
rect 13725 -3865 13775 -3815
rect 13820 -3865 13870 -3815
rect 13915 -3865 13965 -3815
rect 14015 -3865 14065 -3815
rect 14115 -3865 14165 -3815
rect 14215 -3865 14265 -3815
rect 14310 -3865 14360 -3815
rect 14405 -3865 14455 -3815
rect 14525 -3865 14575 -3815
rect 14620 -3865 14670 -3815
rect 14715 -3865 14765 -3815
rect 14815 -3865 14865 -3815
rect 14915 -3865 14965 -3815
rect 15015 -3865 15065 -3815
rect 15110 -3865 15160 -3815
rect 15205 -3865 15255 -3815
rect 15325 -3865 15375 -3815
rect 15420 -3865 15470 -3815
rect 15515 -3865 15565 -3815
rect 15615 -3865 15665 -3815
rect 15715 -3865 15765 -3815
rect 15815 -3865 15865 -3815
rect 15910 -3865 15960 -3815
rect 16005 -3865 16055 -3815
rect 12925 -3965 12975 -3915
rect 13020 -3965 13070 -3915
rect 13115 -3965 13165 -3915
rect 13215 -3965 13265 -3915
rect 13315 -3965 13365 -3915
rect 13415 -3965 13465 -3915
rect 13510 -3965 13560 -3915
rect 13605 -3965 13655 -3915
rect 13725 -3965 13775 -3915
rect 13820 -3965 13870 -3915
rect 13915 -3965 13965 -3915
rect 14015 -3965 14065 -3915
rect 14115 -3965 14165 -3915
rect 14215 -3965 14265 -3915
rect 14310 -3965 14360 -3915
rect 14405 -3965 14455 -3915
rect 14525 -3965 14575 -3915
rect 14620 -3965 14670 -3915
rect 14715 -3965 14765 -3915
rect 14815 -3965 14865 -3915
rect 14915 -3965 14965 -3915
rect 15015 -3965 15065 -3915
rect 15110 -3965 15160 -3915
rect 15205 -3965 15255 -3915
rect 15325 -3965 15375 -3915
rect 15420 -3965 15470 -3915
rect 15515 -3965 15565 -3915
rect 15615 -3965 15665 -3915
rect 15715 -3965 15765 -3915
rect 15815 -3965 15865 -3915
rect 15910 -3965 15960 -3915
rect 16005 -3965 16055 -3915
rect 12925 -4055 12975 -4005
rect 13020 -4055 13070 -4005
rect 13115 -4055 13165 -4005
rect 13215 -4055 13265 -4005
rect 13315 -4055 13365 -4005
rect 13415 -4055 13465 -4005
rect 13510 -4055 13560 -4005
rect 13605 -4055 13655 -4005
rect 13725 -4055 13775 -4005
rect 13820 -4055 13870 -4005
rect 13915 -4055 13965 -4005
rect 14015 -4055 14065 -4005
rect 14115 -4055 14165 -4005
rect 14215 -4055 14265 -4005
rect 14310 -4055 14360 -4005
rect 14405 -4055 14455 -4005
rect 14525 -4055 14575 -4005
rect 14620 -4055 14670 -4005
rect 14715 -4055 14765 -4005
rect 14815 -4055 14865 -4005
rect 14915 -4055 14965 -4005
rect 15015 -4055 15065 -4005
rect 15110 -4055 15160 -4005
rect 15205 -4055 15255 -4005
rect 15325 -4055 15375 -4005
rect 15420 -4055 15470 -4005
rect 15515 -4055 15565 -4005
rect 15615 -4055 15665 -4005
rect 15715 -4055 15765 -4005
rect 15815 -4055 15865 -4005
rect 15910 -4055 15960 -4005
rect 16005 -4055 16055 -4005
rect 12925 -4175 12975 -4125
rect 13020 -4175 13070 -4125
rect 13115 -4175 13165 -4125
rect 13215 -4175 13265 -4125
rect 13315 -4175 13365 -4125
rect 13415 -4175 13465 -4125
rect 13510 -4175 13560 -4125
rect 13605 -4175 13655 -4125
rect 13725 -4175 13775 -4125
rect 13820 -4175 13870 -4125
rect 13915 -4175 13965 -4125
rect 14015 -4175 14065 -4125
rect 14115 -4175 14165 -4125
rect 14215 -4175 14265 -4125
rect 14310 -4175 14360 -4125
rect 14405 -4175 14455 -4125
rect 14525 -4175 14575 -4125
rect 14620 -4175 14670 -4125
rect 14715 -4175 14765 -4125
rect 14815 -4175 14865 -4125
rect 14915 -4175 14965 -4125
rect 15015 -4175 15065 -4125
rect 15110 -4175 15160 -4125
rect 15205 -4175 15255 -4125
rect 15325 -4175 15375 -4125
rect 15420 -4175 15470 -4125
rect 15515 -4175 15565 -4125
rect 15615 -4175 15665 -4125
rect 15715 -4175 15765 -4125
rect 15815 -4175 15865 -4125
rect 15910 -4175 15960 -4125
rect 16005 -4175 16055 -4125
rect 12925 -4265 12975 -4215
rect 13020 -4265 13070 -4215
rect 13115 -4265 13165 -4215
rect 13215 -4265 13265 -4215
rect 13315 -4265 13365 -4215
rect 13415 -4265 13465 -4215
rect 13510 -4265 13560 -4215
rect 13605 -4265 13655 -4215
rect 13725 -4265 13775 -4215
rect 13820 -4265 13870 -4215
rect 13915 -4265 13965 -4215
rect 14015 -4265 14065 -4215
rect 14115 -4265 14165 -4215
rect 14215 -4265 14265 -4215
rect 14310 -4265 14360 -4215
rect 14405 -4265 14455 -4215
rect 14525 -4265 14575 -4215
rect 14620 -4265 14670 -4215
rect 14715 -4265 14765 -4215
rect 14815 -4265 14865 -4215
rect 14915 -4265 14965 -4215
rect 15015 -4265 15065 -4215
rect 15110 -4265 15160 -4215
rect 15205 -4265 15255 -4215
rect 15325 -4265 15375 -4215
rect 15420 -4265 15470 -4215
rect 15515 -4265 15565 -4215
rect 15615 -4265 15665 -4215
rect 15715 -4265 15765 -4215
rect 15815 -4265 15865 -4215
rect 15910 -4265 15960 -4215
rect 16005 -4265 16055 -4215
rect 12925 -4365 12975 -4315
rect 13020 -4365 13070 -4315
rect 13115 -4365 13165 -4315
rect 13215 -4365 13265 -4315
rect 13315 -4365 13365 -4315
rect 13415 -4365 13465 -4315
rect 13510 -4365 13560 -4315
rect 13605 -4365 13655 -4315
rect 13725 -4365 13775 -4315
rect 13820 -4365 13870 -4315
rect 13915 -4365 13965 -4315
rect 14015 -4365 14065 -4315
rect 14115 -4365 14165 -4315
rect 14215 -4365 14265 -4315
rect 14310 -4365 14360 -4315
rect 14405 -4365 14455 -4315
rect 14525 -4365 14575 -4315
rect 14620 -4365 14670 -4315
rect 14715 -4365 14765 -4315
rect 14815 -4365 14865 -4315
rect 14915 -4365 14965 -4315
rect 15015 -4365 15065 -4315
rect 15110 -4365 15160 -4315
rect 15205 -4365 15255 -4315
rect 15325 -4365 15375 -4315
rect 15420 -4365 15470 -4315
rect 15515 -4365 15565 -4315
rect 15615 -4365 15665 -4315
rect 15715 -4365 15765 -4315
rect 15815 -4365 15865 -4315
rect 15910 -4365 15960 -4315
rect 16005 -4365 16055 -4315
rect 12925 -4455 12975 -4405
rect 13020 -4455 13070 -4405
rect 13115 -4455 13165 -4405
rect 13215 -4455 13265 -4405
rect 13315 -4455 13365 -4405
rect 13415 -4455 13465 -4405
rect 13510 -4455 13560 -4405
rect 13605 -4455 13655 -4405
rect 13725 -4455 13775 -4405
rect 13820 -4455 13870 -4405
rect 13915 -4455 13965 -4405
rect 14015 -4455 14065 -4405
rect 14115 -4455 14165 -4405
rect 14215 -4455 14265 -4405
rect 14310 -4455 14360 -4405
rect 14405 -4455 14455 -4405
rect 14525 -4455 14575 -4405
rect 14620 -4455 14670 -4405
rect 14715 -4455 14765 -4405
rect 14815 -4455 14865 -4405
rect 14915 -4455 14965 -4405
rect 15015 -4455 15065 -4405
rect 15110 -4455 15160 -4405
rect 15205 -4455 15255 -4405
rect 15325 -4455 15375 -4405
rect 15420 -4455 15470 -4405
rect 15515 -4455 15565 -4405
rect 15615 -4455 15665 -4405
rect 15715 -4455 15765 -4405
rect 15815 -4455 15865 -4405
rect 15910 -4455 15960 -4405
rect 16005 -4455 16055 -4405
<< metal4 >>
rect 2150 20915 16090 20925
rect 2150 20875 2190 20915
rect 2230 20875 6660 20915
rect 6700 20890 16090 20915
rect 6700 20875 12925 20890
rect 2150 20850 12925 20875
rect 2150 20810 2190 20850
rect 2230 20810 6660 20850
rect 6700 20840 12925 20850
rect 12975 20840 13020 20890
rect 13070 20840 13115 20890
rect 13165 20840 13215 20890
rect 13265 20840 13315 20890
rect 13365 20840 13415 20890
rect 13465 20840 13510 20890
rect 13560 20840 13605 20890
rect 13655 20840 13725 20890
rect 13775 20840 13820 20890
rect 13870 20840 13915 20890
rect 13965 20840 14015 20890
rect 14065 20840 14115 20890
rect 14165 20840 14215 20890
rect 14265 20840 14310 20890
rect 14360 20840 14405 20890
rect 14455 20840 14525 20890
rect 14575 20840 14620 20890
rect 14670 20840 14715 20890
rect 14765 20840 14815 20890
rect 14865 20840 14915 20890
rect 14965 20840 15015 20890
rect 15065 20840 15110 20890
rect 15160 20840 15205 20890
rect 15255 20840 15325 20890
rect 15375 20840 15420 20890
rect 15470 20840 15515 20890
rect 15565 20840 15615 20890
rect 15665 20840 15715 20890
rect 15765 20840 15815 20890
rect 15865 20840 15910 20890
rect 15960 20840 16005 20890
rect 16055 20840 16090 20890
rect 6700 20810 16090 20840
rect 2150 20800 16090 20810
rect 2150 20780 12925 20800
rect 2150 20740 2190 20780
rect 2230 20740 6660 20780
rect 6700 20750 12925 20780
rect 12975 20750 13020 20800
rect 13070 20750 13115 20800
rect 13165 20750 13215 20800
rect 13265 20750 13315 20800
rect 13365 20750 13415 20800
rect 13465 20750 13510 20800
rect 13560 20750 13605 20800
rect 13655 20750 13725 20800
rect 13775 20750 13820 20800
rect 13870 20750 13915 20800
rect 13965 20750 14015 20800
rect 14065 20750 14115 20800
rect 14165 20750 14215 20800
rect 14265 20750 14310 20800
rect 14360 20750 14405 20800
rect 14455 20750 14525 20800
rect 14575 20750 14620 20800
rect 14670 20750 14715 20800
rect 14765 20750 14815 20800
rect 14865 20750 14915 20800
rect 14965 20750 15015 20800
rect 15065 20750 15110 20800
rect 15160 20750 15205 20800
rect 15255 20750 15325 20800
rect 15375 20750 15420 20800
rect 15470 20750 15515 20800
rect 15565 20750 15615 20800
rect 15665 20750 15715 20800
rect 15765 20750 15815 20800
rect 15865 20750 15910 20800
rect 15960 20750 16005 20800
rect 16055 20750 16090 20800
rect 6700 20740 16090 20750
rect 2150 20710 16090 20740
rect 2150 20670 2190 20710
rect 2230 20670 6660 20710
rect 6700 20700 16090 20710
rect 6700 20670 12925 20700
rect 2150 20650 12925 20670
rect 12975 20650 13020 20700
rect 13070 20650 13115 20700
rect 13165 20650 13215 20700
rect 13265 20650 13315 20700
rect 13365 20650 13415 20700
rect 13465 20650 13510 20700
rect 13560 20650 13605 20700
rect 13655 20650 13725 20700
rect 13775 20650 13820 20700
rect 13870 20650 13915 20700
rect 13965 20650 14015 20700
rect 14065 20650 14115 20700
rect 14165 20650 14215 20700
rect 14265 20650 14310 20700
rect 14360 20650 14405 20700
rect 14455 20650 14525 20700
rect 14575 20650 14620 20700
rect 14670 20650 14715 20700
rect 14765 20650 14815 20700
rect 14865 20650 14915 20700
rect 14965 20650 15015 20700
rect 15065 20650 15110 20700
rect 15160 20650 15205 20700
rect 15255 20650 15325 20700
rect 15375 20650 15420 20700
rect 15470 20650 15515 20700
rect 15565 20650 15615 20700
rect 15665 20650 15715 20700
rect 15765 20650 15815 20700
rect 15865 20650 15910 20700
rect 15960 20650 16005 20700
rect 16055 20650 16090 20700
rect 2150 20640 16090 20650
rect 2150 20600 2190 20640
rect 2230 20600 6660 20640
rect 6700 20610 16090 20640
rect 6700 20600 12925 20610
rect 2150 20575 12925 20600
rect 2150 20535 2190 20575
rect 2230 20535 6660 20575
rect 6700 20560 12925 20575
rect 12975 20560 13020 20610
rect 13070 20560 13115 20610
rect 13165 20560 13215 20610
rect 13265 20560 13315 20610
rect 13365 20560 13415 20610
rect 13465 20560 13510 20610
rect 13560 20560 13605 20610
rect 13655 20560 13725 20610
rect 13775 20560 13820 20610
rect 13870 20560 13915 20610
rect 13965 20560 14015 20610
rect 14065 20560 14115 20610
rect 14165 20560 14215 20610
rect 14265 20560 14310 20610
rect 14360 20560 14405 20610
rect 14455 20560 14525 20610
rect 14575 20560 14620 20610
rect 14670 20560 14715 20610
rect 14765 20560 14815 20610
rect 14865 20560 14915 20610
rect 14965 20560 15015 20610
rect 15065 20560 15110 20610
rect 15160 20560 15205 20610
rect 15255 20560 15325 20610
rect 15375 20560 15420 20610
rect 15470 20560 15515 20610
rect 15565 20560 15615 20610
rect 15665 20560 15715 20610
rect 15765 20560 15815 20610
rect 15865 20560 15910 20610
rect 15960 20560 16005 20610
rect 16055 20560 16090 20610
rect 6700 20535 16090 20560
rect 2150 20515 16090 20535
rect 2150 20475 2190 20515
rect 2230 20475 6660 20515
rect 6700 20490 16090 20515
rect 6700 20475 12925 20490
rect 2150 20450 12925 20475
rect 2150 20410 2190 20450
rect 2230 20410 6660 20450
rect 6700 20440 12925 20450
rect 12975 20440 13020 20490
rect 13070 20440 13115 20490
rect 13165 20440 13215 20490
rect 13265 20440 13315 20490
rect 13365 20440 13415 20490
rect 13465 20440 13510 20490
rect 13560 20440 13605 20490
rect 13655 20440 13725 20490
rect 13775 20440 13820 20490
rect 13870 20440 13915 20490
rect 13965 20440 14015 20490
rect 14065 20440 14115 20490
rect 14165 20440 14215 20490
rect 14265 20440 14310 20490
rect 14360 20440 14405 20490
rect 14455 20440 14525 20490
rect 14575 20440 14620 20490
rect 14670 20440 14715 20490
rect 14765 20440 14815 20490
rect 14865 20440 14915 20490
rect 14965 20440 15015 20490
rect 15065 20440 15110 20490
rect 15160 20440 15205 20490
rect 15255 20440 15325 20490
rect 15375 20440 15420 20490
rect 15470 20440 15515 20490
rect 15565 20440 15615 20490
rect 15665 20440 15715 20490
rect 15765 20440 15815 20490
rect 15865 20440 15910 20490
rect 15960 20440 16005 20490
rect 16055 20440 16090 20490
rect 6700 20410 16090 20440
rect 2150 20400 16090 20410
rect 2150 20380 12925 20400
rect 2150 20340 2190 20380
rect 2230 20340 6660 20380
rect 6700 20350 12925 20380
rect 12975 20350 13020 20400
rect 13070 20350 13115 20400
rect 13165 20350 13215 20400
rect 13265 20350 13315 20400
rect 13365 20350 13415 20400
rect 13465 20350 13510 20400
rect 13560 20350 13605 20400
rect 13655 20350 13725 20400
rect 13775 20350 13820 20400
rect 13870 20350 13915 20400
rect 13965 20350 14015 20400
rect 14065 20350 14115 20400
rect 14165 20350 14215 20400
rect 14265 20350 14310 20400
rect 14360 20350 14405 20400
rect 14455 20350 14525 20400
rect 14575 20350 14620 20400
rect 14670 20350 14715 20400
rect 14765 20350 14815 20400
rect 14865 20350 14915 20400
rect 14965 20350 15015 20400
rect 15065 20350 15110 20400
rect 15160 20350 15205 20400
rect 15255 20350 15325 20400
rect 15375 20350 15420 20400
rect 15470 20350 15515 20400
rect 15565 20350 15615 20400
rect 15665 20350 15715 20400
rect 15765 20350 15815 20400
rect 15865 20350 15910 20400
rect 15960 20350 16005 20400
rect 16055 20350 16090 20400
rect 6700 20340 16090 20350
rect 2150 20310 16090 20340
rect 2150 20270 2190 20310
rect 2230 20270 6660 20310
rect 6700 20300 16090 20310
rect 6700 20270 12925 20300
rect 2150 20250 12925 20270
rect 12975 20250 13020 20300
rect 13070 20250 13115 20300
rect 13165 20250 13215 20300
rect 13265 20250 13315 20300
rect 13365 20250 13415 20300
rect 13465 20250 13510 20300
rect 13560 20250 13605 20300
rect 13655 20250 13725 20300
rect 13775 20250 13820 20300
rect 13870 20250 13915 20300
rect 13965 20250 14015 20300
rect 14065 20250 14115 20300
rect 14165 20250 14215 20300
rect 14265 20250 14310 20300
rect 14360 20250 14405 20300
rect 14455 20250 14525 20300
rect 14575 20250 14620 20300
rect 14670 20250 14715 20300
rect 14765 20250 14815 20300
rect 14865 20250 14915 20300
rect 14965 20250 15015 20300
rect 15065 20250 15110 20300
rect 15160 20250 15205 20300
rect 15255 20250 15325 20300
rect 15375 20250 15420 20300
rect 15470 20250 15515 20300
rect 15565 20250 15615 20300
rect 15665 20250 15715 20300
rect 15765 20250 15815 20300
rect 15865 20250 15910 20300
rect 15960 20250 16005 20300
rect 16055 20250 16090 20300
rect 2150 20240 16090 20250
rect 2150 20200 2190 20240
rect 2230 20200 6660 20240
rect 6700 20210 16090 20240
rect 6700 20200 12925 20210
rect 2150 20175 12925 20200
rect 2150 20135 2190 20175
rect 2230 20135 6660 20175
rect 6700 20160 12925 20175
rect 12975 20160 13020 20210
rect 13070 20160 13115 20210
rect 13165 20160 13215 20210
rect 13265 20160 13315 20210
rect 13365 20160 13415 20210
rect 13465 20160 13510 20210
rect 13560 20160 13605 20210
rect 13655 20160 13725 20210
rect 13775 20160 13820 20210
rect 13870 20160 13915 20210
rect 13965 20160 14015 20210
rect 14065 20160 14115 20210
rect 14165 20160 14215 20210
rect 14265 20160 14310 20210
rect 14360 20160 14405 20210
rect 14455 20160 14525 20210
rect 14575 20160 14620 20210
rect 14670 20160 14715 20210
rect 14765 20160 14815 20210
rect 14865 20160 14915 20210
rect 14965 20160 15015 20210
rect 15065 20160 15110 20210
rect 15160 20160 15205 20210
rect 15255 20160 15325 20210
rect 15375 20160 15420 20210
rect 15470 20160 15515 20210
rect 15565 20160 15615 20210
rect 15665 20160 15715 20210
rect 15765 20160 15815 20210
rect 15865 20160 15910 20210
rect 15960 20160 16005 20210
rect 16055 20160 16090 20210
rect 6700 20135 16090 20160
rect 2150 20115 16090 20135
rect 2150 20075 2190 20115
rect 2230 20075 6660 20115
rect 6700 20090 16090 20115
rect 6700 20075 12925 20090
rect 2150 20050 12925 20075
rect 2150 20010 2190 20050
rect 2230 20010 6660 20050
rect 6700 20040 12925 20050
rect 12975 20040 13020 20090
rect 13070 20040 13115 20090
rect 13165 20040 13215 20090
rect 13265 20040 13315 20090
rect 13365 20040 13415 20090
rect 13465 20040 13510 20090
rect 13560 20040 13605 20090
rect 13655 20040 13725 20090
rect 13775 20040 13820 20090
rect 13870 20040 13915 20090
rect 13965 20040 14015 20090
rect 14065 20040 14115 20090
rect 14165 20040 14215 20090
rect 14265 20040 14310 20090
rect 14360 20040 14405 20090
rect 14455 20040 14525 20090
rect 14575 20040 14620 20090
rect 14670 20040 14715 20090
rect 14765 20040 14815 20090
rect 14865 20040 14915 20090
rect 14965 20040 15015 20090
rect 15065 20040 15110 20090
rect 15160 20040 15205 20090
rect 15255 20040 15325 20090
rect 15375 20040 15420 20090
rect 15470 20040 15515 20090
rect 15565 20040 15615 20090
rect 15665 20040 15715 20090
rect 15765 20040 15815 20090
rect 15865 20040 15910 20090
rect 15960 20040 16005 20090
rect 16055 20040 16090 20090
rect 6700 20010 16090 20040
rect 2150 20000 16090 20010
rect 2150 19980 12925 20000
rect 2150 19940 2190 19980
rect 2230 19940 6660 19980
rect 6700 19950 12925 19980
rect 12975 19950 13020 20000
rect 13070 19950 13115 20000
rect 13165 19950 13215 20000
rect 13265 19950 13315 20000
rect 13365 19950 13415 20000
rect 13465 19950 13510 20000
rect 13560 19950 13605 20000
rect 13655 19950 13725 20000
rect 13775 19950 13820 20000
rect 13870 19950 13915 20000
rect 13965 19950 14015 20000
rect 14065 19950 14115 20000
rect 14165 19950 14215 20000
rect 14265 19950 14310 20000
rect 14360 19950 14405 20000
rect 14455 19950 14525 20000
rect 14575 19950 14620 20000
rect 14670 19950 14715 20000
rect 14765 19950 14815 20000
rect 14865 19950 14915 20000
rect 14965 19950 15015 20000
rect 15065 19950 15110 20000
rect 15160 19950 15205 20000
rect 15255 19950 15325 20000
rect 15375 19950 15420 20000
rect 15470 19950 15515 20000
rect 15565 19950 15615 20000
rect 15665 19950 15715 20000
rect 15765 19950 15815 20000
rect 15865 19950 15910 20000
rect 15960 19950 16005 20000
rect 16055 19950 16090 20000
rect 6700 19940 16090 19950
rect 2150 19910 16090 19940
rect 2150 19870 2190 19910
rect 2230 19870 6660 19910
rect 6700 19900 16090 19910
rect 6700 19870 12925 19900
rect 2150 19850 12925 19870
rect 12975 19850 13020 19900
rect 13070 19850 13115 19900
rect 13165 19850 13215 19900
rect 13265 19850 13315 19900
rect 13365 19850 13415 19900
rect 13465 19850 13510 19900
rect 13560 19850 13605 19900
rect 13655 19850 13725 19900
rect 13775 19850 13820 19900
rect 13870 19850 13915 19900
rect 13965 19850 14015 19900
rect 14065 19850 14115 19900
rect 14165 19850 14215 19900
rect 14265 19850 14310 19900
rect 14360 19850 14405 19900
rect 14455 19850 14525 19900
rect 14575 19850 14620 19900
rect 14670 19850 14715 19900
rect 14765 19850 14815 19900
rect 14865 19850 14915 19900
rect 14965 19850 15015 19900
rect 15065 19850 15110 19900
rect 15160 19850 15205 19900
rect 15255 19850 15325 19900
rect 15375 19850 15420 19900
rect 15470 19850 15515 19900
rect 15565 19850 15615 19900
rect 15665 19850 15715 19900
rect 15765 19850 15815 19900
rect 15865 19850 15910 19900
rect 15960 19850 16005 19900
rect 16055 19850 16090 19900
rect 2150 19840 16090 19850
rect 2150 19800 2190 19840
rect 2230 19800 6660 19840
rect 6700 19810 16090 19840
rect 6700 19800 12925 19810
rect 2150 19775 12925 19800
rect 2150 19735 2190 19775
rect 2230 19735 6660 19775
rect 6700 19760 12925 19775
rect 12975 19760 13020 19810
rect 13070 19760 13115 19810
rect 13165 19760 13215 19810
rect 13265 19760 13315 19810
rect 13365 19760 13415 19810
rect 13465 19760 13510 19810
rect 13560 19760 13605 19810
rect 13655 19760 13725 19810
rect 13775 19760 13820 19810
rect 13870 19760 13915 19810
rect 13965 19760 14015 19810
rect 14065 19760 14115 19810
rect 14165 19760 14215 19810
rect 14265 19760 14310 19810
rect 14360 19760 14405 19810
rect 14455 19760 14525 19810
rect 14575 19760 14620 19810
rect 14670 19760 14715 19810
rect 14765 19760 14815 19810
rect 14865 19760 14915 19810
rect 14965 19760 15015 19810
rect 15065 19760 15110 19810
rect 15160 19760 15205 19810
rect 15255 19760 15325 19810
rect 15375 19760 15420 19810
rect 15470 19760 15515 19810
rect 15565 19760 15615 19810
rect 15665 19760 15715 19810
rect 15765 19760 15815 19810
rect 15865 19760 15910 19810
rect 15960 19760 16005 19810
rect 16055 19760 16090 19810
rect 6700 19735 16090 19760
rect 2150 19715 16090 19735
rect 2150 19675 2190 19715
rect 2230 19675 6660 19715
rect 6700 19690 16090 19715
rect 6700 19675 12925 19690
rect 2150 19650 12925 19675
rect 2150 19610 2190 19650
rect 2230 19610 6660 19650
rect 6700 19640 12925 19650
rect 12975 19640 13020 19690
rect 13070 19640 13115 19690
rect 13165 19640 13215 19690
rect 13265 19640 13315 19690
rect 13365 19640 13415 19690
rect 13465 19640 13510 19690
rect 13560 19640 13605 19690
rect 13655 19640 13725 19690
rect 13775 19640 13820 19690
rect 13870 19640 13915 19690
rect 13965 19640 14015 19690
rect 14065 19640 14115 19690
rect 14165 19640 14215 19690
rect 14265 19640 14310 19690
rect 14360 19640 14405 19690
rect 14455 19640 14525 19690
rect 14575 19640 14620 19690
rect 14670 19640 14715 19690
rect 14765 19640 14815 19690
rect 14865 19640 14915 19690
rect 14965 19640 15015 19690
rect 15065 19640 15110 19690
rect 15160 19640 15205 19690
rect 15255 19640 15325 19690
rect 15375 19640 15420 19690
rect 15470 19640 15515 19690
rect 15565 19640 15615 19690
rect 15665 19640 15715 19690
rect 15765 19640 15815 19690
rect 15865 19640 15910 19690
rect 15960 19640 16005 19690
rect 16055 19640 16090 19690
rect 6700 19610 16090 19640
rect 2150 19600 16090 19610
rect 2150 19580 12925 19600
rect 2150 19540 2190 19580
rect 2230 19540 6660 19580
rect 6700 19550 12925 19580
rect 12975 19550 13020 19600
rect 13070 19550 13115 19600
rect 13165 19550 13215 19600
rect 13265 19550 13315 19600
rect 13365 19550 13415 19600
rect 13465 19550 13510 19600
rect 13560 19550 13605 19600
rect 13655 19550 13725 19600
rect 13775 19550 13820 19600
rect 13870 19550 13915 19600
rect 13965 19550 14015 19600
rect 14065 19550 14115 19600
rect 14165 19550 14215 19600
rect 14265 19550 14310 19600
rect 14360 19550 14405 19600
rect 14455 19550 14525 19600
rect 14575 19550 14620 19600
rect 14670 19550 14715 19600
rect 14765 19550 14815 19600
rect 14865 19550 14915 19600
rect 14965 19550 15015 19600
rect 15065 19550 15110 19600
rect 15160 19550 15205 19600
rect 15255 19550 15325 19600
rect 15375 19550 15420 19600
rect 15470 19550 15515 19600
rect 15565 19550 15615 19600
rect 15665 19550 15715 19600
rect 15765 19550 15815 19600
rect 15865 19550 15910 19600
rect 15960 19550 16005 19600
rect 16055 19550 16090 19600
rect 6700 19540 16090 19550
rect 2150 19510 16090 19540
rect 2150 19470 2190 19510
rect 2230 19470 6660 19510
rect 6700 19500 16090 19510
rect 6700 19470 12925 19500
rect 2150 19450 12925 19470
rect 12975 19450 13020 19500
rect 13070 19450 13115 19500
rect 13165 19450 13215 19500
rect 13265 19450 13315 19500
rect 13365 19450 13415 19500
rect 13465 19450 13510 19500
rect 13560 19450 13605 19500
rect 13655 19450 13725 19500
rect 13775 19450 13820 19500
rect 13870 19450 13915 19500
rect 13965 19450 14015 19500
rect 14065 19450 14115 19500
rect 14165 19450 14215 19500
rect 14265 19450 14310 19500
rect 14360 19450 14405 19500
rect 14455 19450 14525 19500
rect 14575 19450 14620 19500
rect 14670 19450 14715 19500
rect 14765 19450 14815 19500
rect 14865 19450 14915 19500
rect 14965 19450 15015 19500
rect 15065 19450 15110 19500
rect 15160 19450 15205 19500
rect 15255 19450 15325 19500
rect 15375 19450 15420 19500
rect 15470 19450 15515 19500
rect 15565 19450 15615 19500
rect 15665 19450 15715 19500
rect 15765 19450 15815 19500
rect 15865 19450 15910 19500
rect 15960 19450 16005 19500
rect 16055 19450 16090 19500
rect 2150 19440 16090 19450
rect 2150 19400 2190 19440
rect 2230 19400 6660 19440
rect 6700 19410 16090 19440
rect 6700 19400 12925 19410
rect 2150 19375 12925 19400
rect 2150 19335 2190 19375
rect 2230 19335 6660 19375
rect 6700 19360 12925 19375
rect 12975 19360 13020 19410
rect 13070 19360 13115 19410
rect 13165 19360 13215 19410
rect 13265 19360 13315 19410
rect 13365 19360 13415 19410
rect 13465 19360 13510 19410
rect 13560 19360 13605 19410
rect 13655 19360 13725 19410
rect 13775 19360 13820 19410
rect 13870 19360 13915 19410
rect 13965 19360 14015 19410
rect 14065 19360 14115 19410
rect 14165 19360 14215 19410
rect 14265 19360 14310 19410
rect 14360 19360 14405 19410
rect 14455 19360 14525 19410
rect 14575 19360 14620 19410
rect 14670 19360 14715 19410
rect 14765 19360 14815 19410
rect 14865 19360 14915 19410
rect 14965 19360 15015 19410
rect 15065 19360 15110 19410
rect 15160 19360 15205 19410
rect 15255 19360 15325 19410
rect 15375 19360 15420 19410
rect 15470 19360 15515 19410
rect 15565 19360 15615 19410
rect 15665 19360 15715 19410
rect 15765 19360 15815 19410
rect 15865 19360 15910 19410
rect 15960 19360 16005 19410
rect 16055 19360 16090 19410
rect 6700 19335 16090 19360
rect 2150 19315 16090 19335
rect 2150 19275 2190 19315
rect 2230 19275 6660 19315
rect 6700 19290 16090 19315
rect 6700 19275 12925 19290
rect 2150 19250 12925 19275
rect 2150 19210 2190 19250
rect 2230 19210 6660 19250
rect 6700 19240 12925 19250
rect 12975 19240 13020 19290
rect 13070 19240 13115 19290
rect 13165 19240 13215 19290
rect 13265 19240 13315 19290
rect 13365 19240 13415 19290
rect 13465 19240 13510 19290
rect 13560 19240 13605 19290
rect 13655 19240 13725 19290
rect 13775 19240 13820 19290
rect 13870 19240 13915 19290
rect 13965 19240 14015 19290
rect 14065 19240 14115 19290
rect 14165 19240 14215 19290
rect 14265 19240 14310 19290
rect 14360 19240 14405 19290
rect 14455 19240 14525 19290
rect 14575 19240 14620 19290
rect 14670 19240 14715 19290
rect 14765 19240 14815 19290
rect 14865 19240 14915 19290
rect 14965 19240 15015 19290
rect 15065 19240 15110 19290
rect 15160 19240 15205 19290
rect 15255 19240 15325 19290
rect 15375 19240 15420 19290
rect 15470 19240 15515 19290
rect 15565 19240 15615 19290
rect 15665 19240 15715 19290
rect 15765 19240 15815 19290
rect 15865 19240 15910 19290
rect 15960 19240 16005 19290
rect 16055 19240 16090 19290
rect 6700 19210 16090 19240
rect 2150 19200 16090 19210
rect 2150 19180 12925 19200
rect 2150 19140 2190 19180
rect 2230 19140 6660 19180
rect 6700 19150 12925 19180
rect 12975 19150 13020 19200
rect 13070 19150 13115 19200
rect 13165 19150 13215 19200
rect 13265 19150 13315 19200
rect 13365 19150 13415 19200
rect 13465 19150 13510 19200
rect 13560 19150 13605 19200
rect 13655 19150 13725 19200
rect 13775 19150 13820 19200
rect 13870 19150 13915 19200
rect 13965 19150 14015 19200
rect 14065 19150 14115 19200
rect 14165 19150 14215 19200
rect 14265 19150 14310 19200
rect 14360 19150 14405 19200
rect 14455 19150 14525 19200
rect 14575 19150 14620 19200
rect 14670 19150 14715 19200
rect 14765 19150 14815 19200
rect 14865 19150 14915 19200
rect 14965 19150 15015 19200
rect 15065 19150 15110 19200
rect 15160 19150 15205 19200
rect 15255 19150 15325 19200
rect 15375 19150 15420 19200
rect 15470 19150 15515 19200
rect 15565 19150 15615 19200
rect 15665 19150 15715 19200
rect 15765 19150 15815 19200
rect 15865 19150 15910 19200
rect 15960 19150 16005 19200
rect 16055 19150 16090 19200
rect 6700 19140 16090 19150
rect 2150 19110 16090 19140
rect 2150 19070 2190 19110
rect 2230 19070 6660 19110
rect 6700 19100 16090 19110
rect 6700 19070 12925 19100
rect 2150 19050 12925 19070
rect 12975 19050 13020 19100
rect 13070 19050 13115 19100
rect 13165 19050 13215 19100
rect 13265 19050 13315 19100
rect 13365 19050 13415 19100
rect 13465 19050 13510 19100
rect 13560 19050 13605 19100
rect 13655 19050 13725 19100
rect 13775 19050 13820 19100
rect 13870 19050 13915 19100
rect 13965 19050 14015 19100
rect 14065 19050 14115 19100
rect 14165 19050 14215 19100
rect 14265 19050 14310 19100
rect 14360 19050 14405 19100
rect 14455 19050 14525 19100
rect 14575 19050 14620 19100
rect 14670 19050 14715 19100
rect 14765 19050 14815 19100
rect 14865 19050 14915 19100
rect 14965 19050 15015 19100
rect 15065 19050 15110 19100
rect 15160 19050 15205 19100
rect 15255 19050 15325 19100
rect 15375 19050 15420 19100
rect 15470 19050 15515 19100
rect 15565 19050 15615 19100
rect 15665 19050 15715 19100
rect 15765 19050 15815 19100
rect 15865 19050 15910 19100
rect 15960 19050 16005 19100
rect 16055 19050 16090 19100
rect 2150 19040 16090 19050
rect 2150 19000 2190 19040
rect 2230 19000 6660 19040
rect 6700 19010 16090 19040
rect 6700 19000 12925 19010
rect 2150 18975 12925 19000
rect 2150 18935 2190 18975
rect 2230 18935 6660 18975
rect 6700 18960 12925 18975
rect 12975 18960 13020 19010
rect 13070 18960 13115 19010
rect 13165 18960 13215 19010
rect 13265 18960 13315 19010
rect 13365 18960 13415 19010
rect 13465 18960 13510 19010
rect 13560 18960 13605 19010
rect 13655 18960 13725 19010
rect 13775 18960 13820 19010
rect 13870 18960 13915 19010
rect 13965 18960 14015 19010
rect 14065 18960 14115 19010
rect 14165 18960 14215 19010
rect 14265 18960 14310 19010
rect 14360 18960 14405 19010
rect 14455 18960 14525 19010
rect 14575 18960 14620 19010
rect 14670 18960 14715 19010
rect 14765 18960 14815 19010
rect 14865 18960 14915 19010
rect 14965 18960 15015 19010
rect 15065 18960 15110 19010
rect 15160 18960 15205 19010
rect 15255 18960 15325 19010
rect 15375 18960 15420 19010
rect 15470 18960 15515 19010
rect 15565 18960 15615 19010
rect 15665 18960 15715 19010
rect 15765 18960 15815 19010
rect 15865 18960 15910 19010
rect 15960 18960 16005 19010
rect 16055 18960 16090 19010
rect 6700 18935 16090 18960
rect 2150 18915 16090 18935
rect 2150 18875 2190 18915
rect 2230 18875 6660 18915
rect 6700 18890 16090 18915
rect 6700 18875 12925 18890
rect 2150 18850 12925 18875
rect 2150 18810 2190 18850
rect 2230 18810 6660 18850
rect 6700 18840 12925 18850
rect 12975 18840 13020 18890
rect 13070 18840 13115 18890
rect 13165 18840 13215 18890
rect 13265 18840 13315 18890
rect 13365 18840 13415 18890
rect 13465 18840 13510 18890
rect 13560 18840 13605 18890
rect 13655 18840 13725 18890
rect 13775 18840 13820 18890
rect 13870 18840 13915 18890
rect 13965 18840 14015 18890
rect 14065 18840 14115 18890
rect 14165 18840 14215 18890
rect 14265 18840 14310 18890
rect 14360 18840 14405 18890
rect 14455 18840 14525 18890
rect 14575 18840 14620 18890
rect 14670 18840 14715 18890
rect 14765 18840 14815 18890
rect 14865 18840 14915 18890
rect 14965 18840 15015 18890
rect 15065 18840 15110 18890
rect 15160 18840 15205 18890
rect 15255 18840 15325 18890
rect 15375 18840 15420 18890
rect 15470 18840 15515 18890
rect 15565 18840 15615 18890
rect 15665 18840 15715 18890
rect 15765 18840 15815 18890
rect 15865 18840 15910 18890
rect 15960 18840 16005 18890
rect 16055 18840 16090 18890
rect 6700 18810 16090 18840
rect 2150 18800 16090 18810
rect 2150 18780 12925 18800
rect 2150 18740 2190 18780
rect 2230 18740 6660 18780
rect 6700 18750 12925 18780
rect 12975 18750 13020 18800
rect 13070 18750 13115 18800
rect 13165 18750 13215 18800
rect 13265 18750 13315 18800
rect 13365 18750 13415 18800
rect 13465 18750 13510 18800
rect 13560 18750 13605 18800
rect 13655 18750 13725 18800
rect 13775 18750 13820 18800
rect 13870 18750 13915 18800
rect 13965 18750 14015 18800
rect 14065 18750 14115 18800
rect 14165 18750 14215 18800
rect 14265 18750 14310 18800
rect 14360 18750 14405 18800
rect 14455 18750 14525 18800
rect 14575 18750 14620 18800
rect 14670 18750 14715 18800
rect 14765 18750 14815 18800
rect 14865 18750 14915 18800
rect 14965 18750 15015 18800
rect 15065 18750 15110 18800
rect 15160 18750 15205 18800
rect 15255 18750 15325 18800
rect 15375 18750 15420 18800
rect 15470 18750 15515 18800
rect 15565 18750 15615 18800
rect 15665 18750 15715 18800
rect 15765 18750 15815 18800
rect 15865 18750 15910 18800
rect 15960 18750 16005 18800
rect 16055 18750 16090 18800
rect 6700 18740 16090 18750
rect 2150 18710 16090 18740
rect 2150 18670 2190 18710
rect 2230 18670 6660 18710
rect 6700 18700 16090 18710
rect 6700 18670 12925 18700
rect 2150 18650 12925 18670
rect 12975 18650 13020 18700
rect 13070 18650 13115 18700
rect 13165 18650 13215 18700
rect 13265 18650 13315 18700
rect 13365 18650 13415 18700
rect 13465 18650 13510 18700
rect 13560 18650 13605 18700
rect 13655 18650 13725 18700
rect 13775 18650 13820 18700
rect 13870 18650 13915 18700
rect 13965 18650 14015 18700
rect 14065 18650 14115 18700
rect 14165 18650 14215 18700
rect 14265 18650 14310 18700
rect 14360 18650 14405 18700
rect 14455 18650 14525 18700
rect 14575 18650 14620 18700
rect 14670 18650 14715 18700
rect 14765 18650 14815 18700
rect 14865 18650 14915 18700
rect 14965 18650 15015 18700
rect 15065 18650 15110 18700
rect 15160 18650 15205 18700
rect 15255 18650 15325 18700
rect 15375 18650 15420 18700
rect 15470 18650 15515 18700
rect 15565 18650 15615 18700
rect 15665 18650 15715 18700
rect 15765 18650 15815 18700
rect 15865 18650 15910 18700
rect 15960 18650 16005 18700
rect 16055 18650 16090 18700
rect 2150 18640 16090 18650
rect 2150 18600 2190 18640
rect 2230 18600 6660 18640
rect 6700 18610 16090 18640
rect 6700 18600 12925 18610
rect 2150 18575 12925 18600
rect 2150 18535 2190 18575
rect 2230 18535 6660 18575
rect 6700 18560 12925 18575
rect 12975 18560 13020 18610
rect 13070 18560 13115 18610
rect 13165 18560 13215 18610
rect 13265 18560 13315 18610
rect 13365 18560 13415 18610
rect 13465 18560 13510 18610
rect 13560 18560 13605 18610
rect 13655 18560 13725 18610
rect 13775 18560 13820 18610
rect 13870 18560 13915 18610
rect 13965 18560 14015 18610
rect 14065 18560 14115 18610
rect 14165 18560 14215 18610
rect 14265 18560 14310 18610
rect 14360 18560 14405 18610
rect 14455 18560 14525 18610
rect 14575 18560 14620 18610
rect 14670 18560 14715 18610
rect 14765 18560 14815 18610
rect 14865 18560 14915 18610
rect 14965 18560 15015 18610
rect 15065 18560 15110 18610
rect 15160 18560 15205 18610
rect 15255 18560 15325 18610
rect 15375 18560 15420 18610
rect 15470 18560 15515 18610
rect 15565 18560 15615 18610
rect 15665 18560 15715 18610
rect 15765 18560 15815 18610
rect 15865 18560 15910 18610
rect 15960 18560 16005 18610
rect 16055 18560 16090 18610
rect 6700 18535 16090 18560
rect 2150 18515 16090 18535
rect 2150 18475 2190 18515
rect 2230 18475 6660 18515
rect 6700 18490 16090 18515
rect 6700 18475 12925 18490
rect 2150 18450 12925 18475
rect 2150 18410 2190 18450
rect 2230 18410 6660 18450
rect 6700 18440 12925 18450
rect 12975 18440 13020 18490
rect 13070 18440 13115 18490
rect 13165 18440 13215 18490
rect 13265 18440 13315 18490
rect 13365 18440 13415 18490
rect 13465 18440 13510 18490
rect 13560 18440 13605 18490
rect 13655 18440 13725 18490
rect 13775 18440 13820 18490
rect 13870 18440 13915 18490
rect 13965 18440 14015 18490
rect 14065 18440 14115 18490
rect 14165 18440 14215 18490
rect 14265 18440 14310 18490
rect 14360 18440 14405 18490
rect 14455 18440 14525 18490
rect 14575 18440 14620 18490
rect 14670 18440 14715 18490
rect 14765 18440 14815 18490
rect 14865 18440 14915 18490
rect 14965 18440 15015 18490
rect 15065 18440 15110 18490
rect 15160 18440 15205 18490
rect 15255 18440 15325 18490
rect 15375 18440 15420 18490
rect 15470 18440 15515 18490
rect 15565 18440 15615 18490
rect 15665 18440 15715 18490
rect 15765 18440 15815 18490
rect 15865 18440 15910 18490
rect 15960 18440 16005 18490
rect 16055 18440 16090 18490
rect 6700 18410 16090 18440
rect 2150 18400 16090 18410
rect 2150 18380 12925 18400
rect 2150 18340 2190 18380
rect 2230 18340 6660 18380
rect 6700 18350 12925 18380
rect 12975 18350 13020 18400
rect 13070 18350 13115 18400
rect 13165 18350 13215 18400
rect 13265 18350 13315 18400
rect 13365 18350 13415 18400
rect 13465 18350 13510 18400
rect 13560 18350 13605 18400
rect 13655 18350 13725 18400
rect 13775 18350 13820 18400
rect 13870 18350 13915 18400
rect 13965 18350 14015 18400
rect 14065 18350 14115 18400
rect 14165 18350 14215 18400
rect 14265 18350 14310 18400
rect 14360 18350 14405 18400
rect 14455 18350 14525 18400
rect 14575 18350 14620 18400
rect 14670 18350 14715 18400
rect 14765 18350 14815 18400
rect 14865 18350 14915 18400
rect 14965 18350 15015 18400
rect 15065 18350 15110 18400
rect 15160 18350 15205 18400
rect 15255 18350 15325 18400
rect 15375 18350 15420 18400
rect 15470 18350 15515 18400
rect 15565 18350 15615 18400
rect 15665 18350 15715 18400
rect 15765 18350 15815 18400
rect 15865 18350 15910 18400
rect 15960 18350 16005 18400
rect 16055 18350 16090 18400
rect 6700 18340 16090 18350
rect 2150 18310 16090 18340
rect 2150 18270 2190 18310
rect 2230 18270 6660 18310
rect 6700 18300 16090 18310
rect 6700 18270 12925 18300
rect 2150 18250 12925 18270
rect 12975 18250 13020 18300
rect 13070 18250 13115 18300
rect 13165 18250 13215 18300
rect 13265 18250 13315 18300
rect 13365 18250 13415 18300
rect 13465 18250 13510 18300
rect 13560 18250 13605 18300
rect 13655 18250 13725 18300
rect 13775 18250 13820 18300
rect 13870 18250 13915 18300
rect 13965 18250 14015 18300
rect 14065 18250 14115 18300
rect 14165 18250 14215 18300
rect 14265 18250 14310 18300
rect 14360 18250 14405 18300
rect 14455 18250 14525 18300
rect 14575 18250 14620 18300
rect 14670 18250 14715 18300
rect 14765 18250 14815 18300
rect 14865 18250 14915 18300
rect 14965 18250 15015 18300
rect 15065 18250 15110 18300
rect 15160 18250 15205 18300
rect 15255 18250 15325 18300
rect 15375 18250 15420 18300
rect 15470 18250 15515 18300
rect 15565 18250 15615 18300
rect 15665 18250 15715 18300
rect 15765 18250 15815 18300
rect 15865 18250 15910 18300
rect 15960 18250 16005 18300
rect 16055 18250 16090 18300
rect 2150 18240 16090 18250
rect 2150 18200 2190 18240
rect 2230 18200 6660 18240
rect 6700 18210 16090 18240
rect 6700 18200 12925 18210
rect 2150 18175 12925 18200
rect 2150 18135 2190 18175
rect 2230 18135 6660 18175
rect 6700 18160 12925 18175
rect 12975 18160 13020 18210
rect 13070 18160 13115 18210
rect 13165 18160 13215 18210
rect 13265 18160 13315 18210
rect 13365 18160 13415 18210
rect 13465 18160 13510 18210
rect 13560 18160 13605 18210
rect 13655 18160 13725 18210
rect 13775 18160 13820 18210
rect 13870 18160 13915 18210
rect 13965 18160 14015 18210
rect 14065 18160 14115 18210
rect 14165 18160 14215 18210
rect 14265 18160 14310 18210
rect 14360 18160 14405 18210
rect 14455 18160 14525 18210
rect 14575 18160 14620 18210
rect 14670 18160 14715 18210
rect 14765 18160 14815 18210
rect 14865 18160 14915 18210
rect 14965 18160 15015 18210
rect 15065 18160 15110 18210
rect 15160 18160 15205 18210
rect 15255 18160 15325 18210
rect 15375 18160 15420 18210
rect 15470 18160 15515 18210
rect 15565 18160 15615 18210
rect 15665 18160 15715 18210
rect 15765 18160 15815 18210
rect 15865 18160 15910 18210
rect 15960 18160 16005 18210
rect 16055 18160 16090 18210
rect 6700 18135 16090 18160
rect 2150 18115 16090 18135
rect 2150 18075 2190 18115
rect 2230 18075 6660 18115
rect 6700 18090 16090 18115
rect 6700 18075 12925 18090
rect 2150 18050 12925 18075
rect 2150 18010 2190 18050
rect 2230 18010 6660 18050
rect 6700 18040 12925 18050
rect 12975 18040 13020 18090
rect 13070 18040 13115 18090
rect 13165 18040 13215 18090
rect 13265 18040 13315 18090
rect 13365 18040 13415 18090
rect 13465 18040 13510 18090
rect 13560 18040 13605 18090
rect 13655 18040 13725 18090
rect 13775 18040 13820 18090
rect 13870 18040 13915 18090
rect 13965 18040 14015 18090
rect 14065 18040 14115 18090
rect 14165 18040 14215 18090
rect 14265 18040 14310 18090
rect 14360 18040 14405 18090
rect 14455 18040 14525 18090
rect 14575 18040 14620 18090
rect 14670 18040 14715 18090
rect 14765 18040 14815 18090
rect 14865 18040 14915 18090
rect 14965 18040 15015 18090
rect 15065 18040 15110 18090
rect 15160 18040 15205 18090
rect 15255 18040 15325 18090
rect 15375 18040 15420 18090
rect 15470 18040 15515 18090
rect 15565 18040 15615 18090
rect 15665 18040 15715 18090
rect 15765 18040 15815 18090
rect 15865 18040 15910 18090
rect 15960 18040 16005 18090
rect 16055 18040 16090 18090
rect 6700 18010 16090 18040
rect 2150 18000 16090 18010
rect 2150 17980 12925 18000
rect 2150 17940 2190 17980
rect 2230 17940 6660 17980
rect 6700 17950 12925 17980
rect 12975 17950 13020 18000
rect 13070 17950 13115 18000
rect 13165 17950 13215 18000
rect 13265 17950 13315 18000
rect 13365 17950 13415 18000
rect 13465 17950 13510 18000
rect 13560 17950 13605 18000
rect 13655 17950 13725 18000
rect 13775 17950 13820 18000
rect 13870 17950 13915 18000
rect 13965 17950 14015 18000
rect 14065 17950 14115 18000
rect 14165 17950 14215 18000
rect 14265 17950 14310 18000
rect 14360 17950 14405 18000
rect 14455 17950 14525 18000
rect 14575 17950 14620 18000
rect 14670 17950 14715 18000
rect 14765 17950 14815 18000
rect 14865 17950 14915 18000
rect 14965 17950 15015 18000
rect 15065 17950 15110 18000
rect 15160 17950 15205 18000
rect 15255 17950 15325 18000
rect 15375 17950 15420 18000
rect 15470 17950 15515 18000
rect 15565 17950 15615 18000
rect 15665 17950 15715 18000
rect 15765 17950 15815 18000
rect 15865 17950 15910 18000
rect 15960 17950 16005 18000
rect 16055 17950 16090 18000
rect 6700 17940 16090 17950
rect 2150 17910 16090 17940
rect 2150 17870 2190 17910
rect 2230 17870 6660 17910
rect 6700 17900 16090 17910
rect 6700 17870 12925 17900
rect 2150 17850 12925 17870
rect 12975 17850 13020 17900
rect 13070 17850 13115 17900
rect 13165 17850 13215 17900
rect 13265 17850 13315 17900
rect 13365 17850 13415 17900
rect 13465 17850 13510 17900
rect 13560 17850 13605 17900
rect 13655 17850 13725 17900
rect 13775 17850 13820 17900
rect 13870 17850 13915 17900
rect 13965 17850 14015 17900
rect 14065 17850 14115 17900
rect 14165 17850 14215 17900
rect 14265 17850 14310 17900
rect 14360 17850 14405 17900
rect 14455 17850 14525 17900
rect 14575 17850 14620 17900
rect 14670 17850 14715 17900
rect 14765 17850 14815 17900
rect 14865 17850 14915 17900
rect 14965 17850 15015 17900
rect 15065 17850 15110 17900
rect 15160 17850 15205 17900
rect 15255 17850 15325 17900
rect 15375 17850 15420 17900
rect 15470 17850 15515 17900
rect 15565 17850 15615 17900
rect 15665 17850 15715 17900
rect 15765 17850 15815 17900
rect 15865 17850 15910 17900
rect 15960 17850 16005 17900
rect 16055 17850 16090 17900
rect 2150 17840 16090 17850
rect 2150 17800 2190 17840
rect 2230 17800 6660 17840
rect 6700 17810 16090 17840
rect 6700 17800 12925 17810
rect 2150 17775 12925 17800
rect 2150 17735 2190 17775
rect 2230 17735 6660 17775
rect 6700 17760 12925 17775
rect 12975 17760 13020 17810
rect 13070 17760 13115 17810
rect 13165 17760 13215 17810
rect 13265 17760 13315 17810
rect 13365 17760 13415 17810
rect 13465 17760 13510 17810
rect 13560 17760 13605 17810
rect 13655 17760 13725 17810
rect 13775 17760 13820 17810
rect 13870 17760 13915 17810
rect 13965 17760 14015 17810
rect 14065 17760 14115 17810
rect 14165 17760 14215 17810
rect 14265 17760 14310 17810
rect 14360 17760 14405 17810
rect 14455 17760 14525 17810
rect 14575 17760 14620 17810
rect 14670 17760 14715 17810
rect 14765 17760 14815 17810
rect 14865 17760 14915 17810
rect 14965 17760 15015 17810
rect 15065 17760 15110 17810
rect 15160 17760 15205 17810
rect 15255 17760 15325 17810
rect 15375 17760 15420 17810
rect 15470 17760 15515 17810
rect 15565 17760 15615 17810
rect 15665 17760 15715 17810
rect 15765 17760 15815 17810
rect 15865 17760 15910 17810
rect 15960 17760 16005 17810
rect 16055 17760 16090 17810
rect 6700 17735 16090 17760
rect 2150 17725 16090 17735
rect -4840 9640 9100 9650
rect -4840 9615 -80 9640
rect -4840 9565 -4805 9615
rect -4755 9565 -4710 9615
rect -4660 9565 -4615 9615
rect -4565 9565 -4515 9615
rect -4465 9565 -4415 9615
rect -4365 9565 -4315 9615
rect -4265 9565 -4220 9615
rect -4170 9565 -4125 9615
rect -4075 9565 -4005 9615
rect -3955 9565 -3910 9615
rect -3860 9565 -3815 9615
rect -3765 9565 -3715 9615
rect -3665 9565 -3615 9615
rect -3565 9565 -3515 9615
rect -3465 9565 -3420 9615
rect -3370 9565 -3325 9615
rect -3275 9565 -3205 9615
rect -3155 9565 -3110 9615
rect -3060 9565 -3015 9615
rect -2965 9565 -2915 9615
rect -2865 9565 -2815 9615
rect -2765 9565 -2715 9615
rect -2665 9565 -2620 9615
rect -2570 9565 -2525 9615
rect -2475 9565 -2405 9615
rect -2355 9565 -2310 9615
rect -2260 9565 -2215 9615
rect -2165 9565 -2115 9615
rect -2065 9565 -2015 9615
rect -1965 9565 -1915 9615
rect -1865 9565 -1820 9615
rect -1770 9565 -1725 9615
rect -1675 9600 -80 9615
rect -40 9600 270 9640
rect 310 9600 620 9640
rect 660 9600 970 9640
rect 1010 9600 1670 9640
rect 1710 9600 2325 9640
rect 2365 9600 3175 9640
rect 3215 9600 3235 9640
rect 3275 9600 3345 9640
rect 3385 9600 6630 9640
rect 6670 9600 7270 9640
rect 7310 9600 7970 9640
rect 8010 9600 8320 9640
rect 8360 9600 8670 9640
rect 8710 9600 9020 9640
rect 9060 9600 9100 9640
rect -1675 9575 9100 9600
rect -1675 9565 -80 9575
rect -4840 9535 -80 9565
rect -40 9535 270 9575
rect 310 9535 620 9575
rect 660 9535 970 9575
rect 1010 9535 1670 9575
rect 1710 9535 2325 9575
rect 2365 9535 3175 9575
rect 3215 9535 3235 9575
rect 3275 9535 3345 9575
rect 3385 9535 6630 9575
rect 6670 9535 7270 9575
rect 7310 9535 7970 9575
rect 8010 9535 8320 9575
rect 8360 9535 8670 9575
rect 8710 9535 9020 9575
rect 9060 9535 9100 9575
rect -4840 9525 9100 9535
rect -4840 9475 -4805 9525
rect -4755 9475 -4710 9525
rect -4660 9475 -4615 9525
rect -4565 9475 -4515 9525
rect -4465 9475 -4415 9525
rect -4365 9475 -4315 9525
rect -4265 9475 -4220 9525
rect -4170 9475 -4125 9525
rect -4075 9475 -4005 9525
rect -3955 9475 -3910 9525
rect -3860 9475 -3815 9525
rect -3765 9475 -3715 9525
rect -3665 9475 -3615 9525
rect -3565 9475 -3515 9525
rect -3465 9475 -3420 9525
rect -3370 9475 -3325 9525
rect -3275 9475 -3205 9525
rect -3155 9475 -3110 9525
rect -3060 9475 -3015 9525
rect -2965 9475 -2915 9525
rect -2865 9475 -2815 9525
rect -2765 9475 -2715 9525
rect -2665 9475 -2620 9525
rect -2570 9475 -2525 9525
rect -2475 9475 -2405 9525
rect -2355 9475 -2310 9525
rect -2260 9475 -2215 9525
rect -2165 9475 -2115 9525
rect -2065 9475 -2015 9525
rect -1965 9475 -1915 9525
rect -1865 9475 -1820 9525
rect -1770 9475 -1725 9525
rect -1675 9505 9100 9525
rect -1675 9475 -80 9505
rect -4840 9465 -80 9475
rect -40 9465 270 9505
rect 310 9465 620 9505
rect 660 9465 970 9505
rect 1010 9465 1670 9505
rect 1710 9465 2325 9505
rect 2365 9465 3175 9505
rect 3215 9465 3235 9505
rect 3275 9465 3345 9505
rect 3385 9465 6630 9505
rect 6670 9465 7270 9505
rect 7310 9465 7970 9505
rect 8010 9465 8320 9505
rect 8360 9465 8670 9505
rect 8710 9465 9020 9505
rect 9060 9465 9100 9505
rect -4840 9435 9100 9465
rect -4840 9425 -80 9435
rect -4840 9375 -4805 9425
rect -4755 9375 -4710 9425
rect -4660 9375 -4615 9425
rect -4565 9375 -4515 9425
rect -4465 9375 -4415 9425
rect -4365 9375 -4315 9425
rect -4265 9375 -4220 9425
rect -4170 9375 -4125 9425
rect -4075 9375 -4005 9425
rect -3955 9375 -3910 9425
rect -3860 9375 -3815 9425
rect -3765 9375 -3715 9425
rect -3665 9375 -3615 9425
rect -3565 9375 -3515 9425
rect -3465 9375 -3420 9425
rect -3370 9375 -3325 9425
rect -3275 9375 -3205 9425
rect -3155 9375 -3110 9425
rect -3060 9375 -3015 9425
rect -2965 9375 -2915 9425
rect -2865 9375 -2815 9425
rect -2765 9375 -2715 9425
rect -2665 9375 -2620 9425
rect -2570 9375 -2525 9425
rect -2475 9375 -2405 9425
rect -2355 9375 -2310 9425
rect -2260 9375 -2215 9425
rect -2165 9375 -2115 9425
rect -2065 9375 -2015 9425
rect -1965 9375 -1915 9425
rect -1865 9375 -1820 9425
rect -1770 9375 -1725 9425
rect -1675 9395 -80 9425
rect -40 9395 270 9435
rect 310 9395 620 9435
rect 660 9395 970 9435
rect 1010 9395 1670 9435
rect 1710 9395 2325 9435
rect 2365 9395 3175 9435
rect 3215 9395 3235 9435
rect 3275 9395 3345 9435
rect 3385 9395 6630 9435
rect 6670 9395 7270 9435
rect 7310 9395 7970 9435
rect 8010 9395 8320 9435
rect 8360 9395 8670 9435
rect 8710 9395 9020 9435
rect 9060 9395 9100 9435
rect -1675 9375 9100 9395
rect -4840 9365 9100 9375
rect -4840 9335 -80 9365
rect -4840 9285 -4805 9335
rect -4755 9285 -4710 9335
rect -4660 9285 -4615 9335
rect -4565 9285 -4515 9335
rect -4465 9285 -4415 9335
rect -4365 9285 -4315 9335
rect -4265 9285 -4220 9335
rect -4170 9285 -4125 9335
rect -4075 9285 -4005 9335
rect -3955 9285 -3910 9335
rect -3860 9285 -3815 9335
rect -3765 9285 -3715 9335
rect -3665 9285 -3615 9335
rect -3565 9285 -3515 9335
rect -3465 9285 -3420 9335
rect -3370 9285 -3325 9335
rect -3275 9285 -3205 9335
rect -3155 9285 -3110 9335
rect -3060 9285 -3015 9335
rect -2965 9285 -2915 9335
rect -2865 9285 -2815 9335
rect -2765 9285 -2715 9335
rect -2665 9285 -2620 9335
rect -2570 9285 -2525 9335
rect -2475 9285 -2405 9335
rect -2355 9285 -2310 9335
rect -2260 9285 -2215 9335
rect -2165 9285 -2115 9335
rect -2065 9285 -2015 9335
rect -1965 9285 -1915 9335
rect -1865 9285 -1820 9335
rect -1770 9285 -1725 9335
rect -1675 9325 -80 9335
rect -40 9325 270 9365
rect 310 9325 620 9365
rect 660 9325 970 9365
rect 1010 9325 1670 9365
rect 1710 9325 2325 9365
rect 2365 9325 3175 9365
rect 3215 9325 3235 9365
rect 3275 9325 3345 9365
rect 3385 9325 6630 9365
rect 6670 9325 7270 9365
rect 7310 9325 7970 9365
rect 8010 9325 8320 9365
rect 8360 9325 8670 9365
rect 8710 9325 9020 9365
rect 9060 9325 9100 9365
rect -1675 9300 9100 9325
rect -1675 9285 -80 9300
rect -4840 9260 -80 9285
rect -40 9260 270 9300
rect 310 9260 620 9300
rect 660 9260 970 9300
rect 1010 9260 1670 9300
rect 1710 9260 2325 9300
rect 2365 9260 3175 9300
rect 3215 9260 3235 9300
rect 3275 9260 3345 9300
rect 3385 9260 6630 9300
rect 6670 9260 7270 9300
rect 7310 9260 7970 9300
rect 8010 9260 8320 9300
rect 8360 9260 8670 9300
rect 8710 9260 9020 9300
rect 9060 9260 9100 9300
rect -4840 9240 9100 9260
rect -4840 9215 -80 9240
rect -4840 9165 -4805 9215
rect -4755 9165 -4710 9215
rect -4660 9165 -4615 9215
rect -4565 9165 -4515 9215
rect -4465 9165 -4415 9215
rect -4365 9165 -4315 9215
rect -4265 9165 -4220 9215
rect -4170 9165 -4125 9215
rect -4075 9165 -4005 9215
rect -3955 9165 -3910 9215
rect -3860 9165 -3815 9215
rect -3765 9165 -3715 9215
rect -3665 9165 -3615 9215
rect -3565 9165 -3515 9215
rect -3465 9165 -3420 9215
rect -3370 9165 -3325 9215
rect -3275 9165 -3205 9215
rect -3155 9165 -3110 9215
rect -3060 9165 -3015 9215
rect -2965 9165 -2915 9215
rect -2865 9165 -2815 9215
rect -2765 9165 -2715 9215
rect -2665 9165 -2620 9215
rect -2570 9165 -2525 9215
rect -2475 9165 -2405 9215
rect -2355 9165 -2310 9215
rect -2260 9165 -2215 9215
rect -2165 9165 -2115 9215
rect -2065 9165 -2015 9215
rect -1965 9165 -1915 9215
rect -1865 9165 -1820 9215
rect -1770 9165 -1725 9215
rect -1675 9200 -80 9215
rect -40 9200 270 9240
rect 310 9200 620 9240
rect 660 9200 970 9240
rect 1010 9200 1670 9240
rect 1710 9200 2325 9240
rect 2365 9200 3175 9240
rect 3215 9200 3235 9240
rect 3275 9200 3345 9240
rect 3385 9200 6630 9240
rect 6670 9200 7270 9240
rect 7310 9200 7970 9240
rect 8010 9200 8320 9240
rect 8360 9200 8670 9240
rect 8710 9200 9020 9240
rect 9060 9200 9100 9240
rect -1675 9175 9100 9200
rect -1675 9165 -80 9175
rect -4840 9135 -80 9165
rect -40 9135 270 9175
rect 310 9135 620 9175
rect 660 9135 970 9175
rect 1010 9135 1670 9175
rect 1710 9135 2325 9175
rect 2365 9135 3175 9175
rect 3215 9135 3235 9175
rect 3275 9135 3345 9175
rect 3385 9135 6630 9175
rect 6670 9135 7270 9175
rect 7310 9135 7970 9175
rect 8010 9135 8320 9175
rect 8360 9135 8670 9175
rect 8710 9135 9020 9175
rect 9060 9135 9100 9175
rect -4840 9125 9100 9135
rect -4840 9075 -4805 9125
rect -4755 9075 -4710 9125
rect -4660 9075 -4615 9125
rect -4565 9075 -4515 9125
rect -4465 9075 -4415 9125
rect -4365 9075 -4315 9125
rect -4265 9075 -4220 9125
rect -4170 9075 -4125 9125
rect -4075 9075 -4005 9125
rect -3955 9075 -3910 9125
rect -3860 9075 -3815 9125
rect -3765 9075 -3715 9125
rect -3665 9075 -3615 9125
rect -3565 9075 -3515 9125
rect -3465 9075 -3420 9125
rect -3370 9075 -3325 9125
rect -3275 9075 -3205 9125
rect -3155 9075 -3110 9125
rect -3060 9075 -3015 9125
rect -2965 9075 -2915 9125
rect -2865 9075 -2815 9125
rect -2765 9075 -2715 9125
rect -2665 9075 -2620 9125
rect -2570 9075 -2525 9125
rect -2475 9075 -2405 9125
rect -2355 9075 -2310 9125
rect -2260 9075 -2215 9125
rect -2165 9075 -2115 9125
rect -2065 9075 -2015 9125
rect -1965 9075 -1915 9125
rect -1865 9075 -1820 9125
rect -1770 9075 -1725 9125
rect -1675 9105 9100 9125
rect -1675 9075 -80 9105
rect -4840 9065 -80 9075
rect -40 9065 270 9105
rect 310 9065 620 9105
rect 660 9065 970 9105
rect 1010 9065 1670 9105
rect 1710 9065 2325 9105
rect 2365 9065 3175 9105
rect 3215 9065 3235 9105
rect 3275 9065 3345 9105
rect 3385 9065 6630 9105
rect 6670 9065 7270 9105
rect 7310 9065 7970 9105
rect 8010 9065 8320 9105
rect 8360 9065 8670 9105
rect 8710 9065 9020 9105
rect 9060 9065 9100 9105
rect -4840 9035 9100 9065
rect -4840 9025 -80 9035
rect -4840 8975 -4805 9025
rect -4755 8975 -4710 9025
rect -4660 8975 -4615 9025
rect -4565 8975 -4515 9025
rect -4465 8975 -4415 9025
rect -4365 8975 -4315 9025
rect -4265 8975 -4220 9025
rect -4170 8975 -4125 9025
rect -4075 8975 -4005 9025
rect -3955 8975 -3910 9025
rect -3860 8975 -3815 9025
rect -3765 8975 -3715 9025
rect -3665 8975 -3615 9025
rect -3565 8975 -3515 9025
rect -3465 8975 -3420 9025
rect -3370 8975 -3325 9025
rect -3275 8975 -3205 9025
rect -3155 8975 -3110 9025
rect -3060 8975 -3015 9025
rect -2965 8975 -2915 9025
rect -2865 8975 -2815 9025
rect -2765 8975 -2715 9025
rect -2665 8975 -2620 9025
rect -2570 8975 -2525 9025
rect -2475 8975 -2405 9025
rect -2355 8975 -2310 9025
rect -2260 8975 -2215 9025
rect -2165 8975 -2115 9025
rect -2065 8975 -2015 9025
rect -1965 8975 -1915 9025
rect -1865 8975 -1820 9025
rect -1770 8975 -1725 9025
rect -1675 8995 -80 9025
rect -40 8995 270 9035
rect 310 8995 620 9035
rect 660 8995 970 9035
rect 1010 8995 1670 9035
rect 1710 8995 2325 9035
rect 2365 8995 3175 9035
rect 3215 8995 3235 9035
rect 3275 8995 3345 9035
rect 3385 8995 6630 9035
rect 6670 8995 7270 9035
rect 7310 8995 7970 9035
rect 8010 8995 8320 9035
rect 8360 8995 8670 9035
rect 8710 8995 9020 9035
rect 9060 8995 9100 9035
rect -1675 8975 9100 8995
rect -4840 8965 9100 8975
rect -4840 8935 -80 8965
rect -4840 8885 -4805 8935
rect -4755 8885 -4710 8935
rect -4660 8885 -4615 8935
rect -4565 8885 -4515 8935
rect -4465 8885 -4415 8935
rect -4365 8885 -4315 8935
rect -4265 8885 -4220 8935
rect -4170 8885 -4125 8935
rect -4075 8885 -4005 8935
rect -3955 8885 -3910 8935
rect -3860 8885 -3815 8935
rect -3765 8885 -3715 8935
rect -3665 8885 -3615 8935
rect -3565 8885 -3515 8935
rect -3465 8885 -3420 8935
rect -3370 8885 -3325 8935
rect -3275 8885 -3205 8935
rect -3155 8885 -3110 8935
rect -3060 8885 -3015 8935
rect -2965 8885 -2915 8935
rect -2865 8885 -2815 8935
rect -2765 8885 -2715 8935
rect -2665 8885 -2620 8935
rect -2570 8885 -2525 8935
rect -2475 8885 -2405 8935
rect -2355 8885 -2310 8935
rect -2260 8885 -2215 8935
rect -2165 8885 -2115 8935
rect -2065 8885 -2015 8935
rect -1965 8885 -1915 8935
rect -1865 8885 -1820 8935
rect -1770 8885 -1725 8935
rect -1675 8925 -80 8935
rect -40 8925 270 8965
rect 310 8925 620 8965
rect 660 8925 970 8965
rect 1010 8925 1670 8965
rect 1710 8925 2325 8965
rect 2365 8925 3175 8965
rect 3215 8925 3235 8965
rect 3275 8925 3345 8965
rect 3385 8925 6630 8965
rect 6670 8925 7270 8965
rect 7310 8925 7970 8965
rect 8010 8925 8320 8965
rect 8360 8925 8670 8965
rect 8710 8925 9020 8965
rect 9060 8925 9100 8965
rect -1675 8900 9100 8925
rect -1675 8885 -80 8900
rect -4840 8860 -80 8885
rect -40 8860 270 8900
rect 310 8860 620 8900
rect 660 8860 970 8900
rect 1010 8860 1670 8900
rect 1710 8860 2325 8900
rect 2365 8860 3175 8900
rect 3215 8860 3235 8900
rect 3275 8860 3345 8900
rect 3385 8860 6630 8900
rect 6670 8860 7270 8900
rect 7310 8860 7970 8900
rect 8010 8860 8320 8900
rect 8360 8860 8670 8900
rect 8710 8860 9020 8900
rect 9060 8860 9100 8900
rect -4840 8840 9100 8860
rect -4840 8815 -80 8840
rect -4840 8765 -4805 8815
rect -4755 8765 -4710 8815
rect -4660 8765 -4615 8815
rect -4565 8765 -4515 8815
rect -4465 8765 -4415 8815
rect -4365 8765 -4315 8815
rect -4265 8765 -4220 8815
rect -4170 8765 -4125 8815
rect -4075 8765 -4005 8815
rect -3955 8765 -3910 8815
rect -3860 8765 -3815 8815
rect -3765 8765 -3715 8815
rect -3665 8765 -3615 8815
rect -3565 8765 -3515 8815
rect -3465 8765 -3420 8815
rect -3370 8765 -3325 8815
rect -3275 8765 -3205 8815
rect -3155 8765 -3110 8815
rect -3060 8765 -3015 8815
rect -2965 8765 -2915 8815
rect -2865 8765 -2815 8815
rect -2765 8765 -2715 8815
rect -2665 8765 -2620 8815
rect -2570 8765 -2525 8815
rect -2475 8765 -2405 8815
rect -2355 8765 -2310 8815
rect -2260 8765 -2215 8815
rect -2165 8765 -2115 8815
rect -2065 8765 -2015 8815
rect -1965 8765 -1915 8815
rect -1865 8765 -1820 8815
rect -1770 8765 -1725 8815
rect -1675 8800 -80 8815
rect -40 8800 270 8840
rect 310 8800 620 8840
rect 660 8800 970 8840
rect 1010 8800 1670 8840
rect 1710 8800 2325 8840
rect 2365 8800 3175 8840
rect 3215 8800 3235 8840
rect 3275 8800 3345 8840
rect 3385 8800 6630 8840
rect 6670 8800 7270 8840
rect 7310 8800 7970 8840
rect 8010 8800 8320 8840
rect 8360 8800 8670 8840
rect 8710 8800 9020 8840
rect 9060 8800 9100 8840
rect -1675 8775 9100 8800
rect -1675 8765 -80 8775
rect -4840 8735 -80 8765
rect -40 8735 270 8775
rect 310 8735 620 8775
rect 660 8735 970 8775
rect 1010 8735 1670 8775
rect 1710 8735 2325 8775
rect 2365 8735 3175 8775
rect 3215 8735 3235 8775
rect 3275 8735 3345 8775
rect 3385 8735 6630 8775
rect 6670 8735 7270 8775
rect 7310 8735 7970 8775
rect 8010 8735 8320 8775
rect 8360 8735 8670 8775
rect 8710 8735 9020 8775
rect 9060 8735 9100 8775
rect -4840 8725 9100 8735
rect -4840 8675 -4805 8725
rect -4755 8675 -4710 8725
rect -4660 8675 -4615 8725
rect -4565 8675 -4515 8725
rect -4465 8675 -4415 8725
rect -4365 8675 -4315 8725
rect -4265 8675 -4220 8725
rect -4170 8675 -4125 8725
rect -4075 8675 -4005 8725
rect -3955 8675 -3910 8725
rect -3860 8675 -3815 8725
rect -3765 8675 -3715 8725
rect -3665 8675 -3615 8725
rect -3565 8675 -3515 8725
rect -3465 8675 -3420 8725
rect -3370 8675 -3325 8725
rect -3275 8675 -3205 8725
rect -3155 8675 -3110 8725
rect -3060 8675 -3015 8725
rect -2965 8675 -2915 8725
rect -2865 8675 -2815 8725
rect -2765 8675 -2715 8725
rect -2665 8675 -2620 8725
rect -2570 8675 -2525 8725
rect -2475 8675 -2405 8725
rect -2355 8675 -2310 8725
rect -2260 8675 -2215 8725
rect -2165 8675 -2115 8725
rect -2065 8675 -2015 8725
rect -1965 8675 -1915 8725
rect -1865 8675 -1820 8725
rect -1770 8675 -1725 8725
rect -1675 8705 9100 8725
rect -1675 8675 -80 8705
rect -4840 8665 -80 8675
rect -40 8665 270 8705
rect 310 8665 620 8705
rect 660 8665 970 8705
rect 1010 8665 1670 8705
rect 1710 8665 2325 8705
rect 2365 8665 3175 8705
rect 3215 8665 3235 8705
rect 3275 8665 3345 8705
rect 3385 8665 6630 8705
rect 6670 8665 7270 8705
rect 7310 8665 7970 8705
rect 8010 8665 8320 8705
rect 8360 8665 8670 8705
rect 8710 8665 9020 8705
rect 9060 8665 9100 8705
rect -4840 8635 9100 8665
rect -4840 8625 -80 8635
rect -4840 8575 -4805 8625
rect -4755 8575 -4710 8625
rect -4660 8575 -4615 8625
rect -4565 8575 -4515 8625
rect -4465 8575 -4415 8625
rect -4365 8575 -4315 8625
rect -4265 8575 -4220 8625
rect -4170 8575 -4125 8625
rect -4075 8575 -4005 8625
rect -3955 8575 -3910 8625
rect -3860 8575 -3815 8625
rect -3765 8575 -3715 8625
rect -3665 8575 -3615 8625
rect -3565 8575 -3515 8625
rect -3465 8575 -3420 8625
rect -3370 8575 -3325 8625
rect -3275 8575 -3205 8625
rect -3155 8575 -3110 8625
rect -3060 8575 -3015 8625
rect -2965 8575 -2915 8625
rect -2865 8575 -2815 8625
rect -2765 8575 -2715 8625
rect -2665 8575 -2620 8625
rect -2570 8575 -2525 8625
rect -2475 8575 -2405 8625
rect -2355 8575 -2310 8625
rect -2260 8575 -2215 8625
rect -2165 8575 -2115 8625
rect -2065 8575 -2015 8625
rect -1965 8575 -1915 8625
rect -1865 8575 -1820 8625
rect -1770 8575 -1725 8625
rect -1675 8595 -80 8625
rect -40 8595 270 8635
rect 310 8595 620 8635
rect 660 8595 970 8635
rect 1010 8595 1670 8635
rect 1710 8595 2325 8635
rect 2365 8595 3175 8635
rect 3215 8595 3235 8635
rect 3275 8595 3345 8635
rect 3385 8595 6630 8635
rect 6670 8595 7270 8635
rect 7310 8595 7970 8635
rect 8010 8595 8320 8635
rect 8360 8595 8670 8635
rect 8710 8595 9020 8635
rect 9060 8595 9100 8635
rect -1675 8575 9100 8595
rect -4840 8565 9100 8575
rect -4840 8535 -80 8565
rect -4840 8485 -4805 8535
rect -4755 8485 -4710 8535
rect -4660 8485 -4615 8535
rect -4565 8485 -4515 8535
rect -4465 8485 -4415 8535
rect -4365 8485 -4315 8535
rect -4265 8485 -4220 8535
rect -4170 8485 -4125 8535
rect -4075 8485 -4005 8535
rect -3955 8485 -3910 8535
rect -3860 8485 -3815 8535
rect -3765 8485 -3715 8535
rect -3665 8485 -3615 8535
rect -3565 8485 -3515 8535
rect -3465 8485 -3420 8535
rect -3370 8485 -3325 8535
rect -3275 8485 -3205 8535
rect -3155 8485 -3110 8535
rect -3060 8485 -3015 8535
rect -2965 8485 -2915 8535
rect -2865 8485 -2815 8535
rect -2765 8485 -2715 8535
rect -2665 8485 -2620 8535
rect -2570 8485 -2525 8535
rect -2475 8485 -2405 8535
rect -2355 8485 -2310 8535
rect -2260 8485 -2215 8535
rect -2165 8485 -2115 8535
rect -2065 8485 -2015 8535
rect -1965 8485 -1915 8535
rect -1865 8485 -1820 8535
rect -1770 8485 -1725 8535
rect -1675 8525 -80 8535
rect -40 8525 270 8565
rect 310 8525 620 8565
rect 660 8525 970 8565
rect 1010 8525 1670 8565
rect 1710 8525 2325 8565
rect 2365 8525 3175 8565
rect 3215 8525 3235 8565
rect 3275 8525 3345 8565
rect 3385 8525 6630 8565
rect 6670 8525 7270 8565
rect 7310 8525 7970 8565
rect 8010 8525 8320 8565
rect 8360 8525 8670 8565
rect 8710 8525 9020 8565
rect 9060 8525 9100 8565
rect -1675 8500 9100 8525
rect -1675 8485 -80 8500
rect -4840 8460 -80 8485
rect -40 8460 270 8500
rect 310 8460 620 8500
rect 660 8460 970 8500
rect 1010 8460 1670 8500
rect 1710 8460 2325 8500
rect 2365 8460 3175 8500
rect 3215 8460 3235 8500
rect 3275 8460 3345 8500
rect 3385 8460 6630 8500
rect 6670 8460 7270 8500
rect 7310 8460 7970 8500
rect 8010 8460 8320 8500
rect 8360 8460 8670 8500
rect 8710 8460 9020 8500
rect 9060 8460 9100 8500
rect -4840 8440 9100 8460
rect -4840 8415 -80 8440
rect -4840 8365 -4805 8415
rect -4755 8365 -4710 8415
rect -4660 8365 -4615 8415
rect -4565 8365 -4515 8415
rect -4465 8365 -4415 8415
rect -4365 8365 -4315 8415
rect -4265 8365 -4220 8415
rect -4170 8365 -4125 8415
rect -4075 8365 -4005 8415
rect -3955 8365 -3910 8415
rect -3860 8365 -3815 8415
rect -3765 8365 -3715 8415
rect -3665 8365 -3615 8415
rect -3565 8365 -3515 8415
rect -3465 8365 -3420 8415
rect -3370 8365 -3325 8415
rect -3275 8365 -3205 8415
rect -3155 8365 -3110 8415
rect -3060 8365 -3015 8415
rect -2965 8365 -2915 8415
rect -2865 8365 -2815 8415
rect -2765 8365 -2715 8415
rect -2665 8365 -2620 8415
rect -2570 8365 -2525 8415
rect -2475 8365 -2405 8415
rect -2355 8365 -2310 8415
rect -2260 8365 -2215 8415
rect -2165 8365 -2115 8415
rect -2065 8365 -2015 8415
rect -1965 8365 -1915 8415
rect -1865 8365 -1820 8415
rect -1770 8365 -1725 8415
rect -1675 8400 -80 8415
rect -40 8400 270 8440
rect 310 8400 620 8440
rect 660 8400 970 8440
rect 1010 8400 1670 8440
rect 1710 8400 2325 8440
rect 2365 8400 3175 8440
rect 3215 8400 3235 8440
rect 3275 8400 3345 8440
rect 3385 8400 6630 8440
rect 6670 8400 7270 8440
rect 7310 8400 7970 8440
rect 8010 8400 8320 8440
rect 8360 8400 8670 8440
rect 8710 8400 9020 8440
rect 9060 8400 9100 8440
rect -1675 8375 9100 8400
rect -1675 8365 -80 8375
rect -4840 8335 -80 8365
rect -40 8335 270 8375
rect 310 8335 620 8375
rect 660 8335 970 8375
rect 1010 8335 1670 8375
rect 1710 8335 2325 8375
rect 2365 8335 3175 8375
rect 3215 8335 3235 8375
rect 3275 8335 3345 8375
rect 3385 8335 6630 8375
rect 6670 8335 7270 8375
rect 7310 8335 7970 8375
rect 8010 8335 8320 8375
rect 8360 8335 8670 8375
rect 8710 8335 9020 8375
rect 9060 8335 9100 8375
rect -4840 8325 9100 8335
rect -4840 8275 -4805 8325
rect -4755 8275 -4710 8325
rect -4660 8275 -4615 8325
rect -4565 8275 -4515 8325
rect -4465 8275 -4415 8325
rect -4365 8275 -4315 8325
rect -4265 8275 -4220 8325
rect -4170 8275 -4125 8325
rect -4075 8275 -4005 8325
rect -3955 8275 -3910 8325
rect -3860 8275 -3815 8325
rect -3765 8275 -3715 8325
rect -3665 8275 -3615 8325
rect -3565 8275 -3515 8325
rect -3465 8275 -3420 8325
rect -3370 8275 -3325 8325
rect -3275 8275 -3205 8325
rect -3155 8275 -3110 8325
rect -3060 8275 -3015 8325
rect -2965 8275 -2915 8325
rect -2865 8275 -2815 8325
rect -2765 8275 -2715 8325
rect -2665 8275 -2620 8325
rect -2570 8275 -2525 8325
rect -2475 8275 -2405 8325
rect -2355 8275 -2310 8325
rect -2260 8275 -2215 8325
rect -2165 8275 -2115 8325
rect -2065 8275 -2015 8325
rect -1965 8275 -1915 8325
rect -1865 8275 -1820 8325
rect -1770 8275 -1725 8325
rect -1675 8305 9100 8325
rect -1675 8275 -80 8305
rect -4840 8265 -80 8275
rect -40 8265 270 8305
rect 310 8265 620 8305
rect 660 8265 970 8305
rect 1010 8265 1670 8305
rect 1710 8265 2325 8305
rect 2365 8265 3175 8305
rect 3215 8265 3235 8305
rect 3275 8265 3345 8305
rect 3385 8265 6630 8305
rect 6670 8265 7270 8305
rect 7310 8265 7970 8305
rect 8010 8265 8320 8305
rect 8360 8265 8670 8305
rect 8710 8265 9020 8305
rect 9060 8265 9100 8305
rect -4840 8235 9100 8265
rect -4840 8225 -80 8235
rect -4840 8175 -4805 8225
rect -4755 8175 -4710 8225
rect -4660 8175 -4615 8225
rect -4565 8175 -4515 8225
rect -4465 8175 -4415 8225
rect -4365 8175 -4315 8225
rect -4265 8175 -4220 8225
rect -4170 8175 -4125 8225
rect -4075 8175 -4005 8225
rect -3955 8175 -3910 8225
rect -3860 8175 -3815 8225
rect -3765 8175 -3715 8225
rect -3665 8175 -3615 8225
rect -3565 8175 -3515 8225
rect -3465 8175 -3420 8225
rect -3370 8175 -3325 8225
rect -3275 8175 -3205 8225
rect -3155 8175 -3110 8225
rect -3060 8175 -3015 8225
rect -2965 8175 -2915 8225
rect -2865 8175 -2815 8225
rect -2765 8175 -2715 8225
rect -2665 8175 -2620 8225
rect -2570 8175 -2525 8225
rect -2475 8175 -2405 8225
rect -2355 8175 -2310 8225
rect -2260 8175 -2215 8225
rect -2165 8175 -2115 8225
rect -2065 8175 -2015 8225
rect -1965 8175 -1915 8225
rect -1865 8175 -1820 8225
rect -1770 8175 -1725 8225
rect -1675 8195 -80 8225
rect -40 8195 270 8235
rect 310 8195 620 8235
rect 660 8195 970 8235
rect 1010 8195 1670 8235
rect 1710 8195 2325 8235
rect 2365 8195 3175 8235
rect 3215 8195 3235 8235
rect 3275 8195 3345 8235
rect 3385 8195 6630 8235
rect 6670 8195 7270 8235
rect 7310 8195 7970 8235
rect 8010 8195 8320 8235
rect 8360 8195 8670 8235
rect 8710 8195 9020 8235
rect 9060 8195 9100 8235
rect -1675 8175 9100 8195
rect -4840 8165 9100 8175
rect -4840 8135 -80 8165
rect -4840 8085 -4805 8135
rect -4755 8085 -4710 8135
rect -4660 8085 -4615 8135
rect -4565 8085 -4515 8135
rect -4465 8085 -4415 8135
rect -4365 8085 -4315 8135
rect -4265 8085 -4220 8135
rect -4170 8085 -4125 8135
rect -4075 8085 -4005 8135
rect -3955 8085 -3910 8135
rect -3860 8085 -3815 8135
rect -3765 8085 -3715 8135
rect -3665 8085 -3615 8135
rect -3565 8085 -3515 8135
rect -3465 8085 -3420 8135
rect -3370 8085 -3325 8135
rect -3275 8085 -3205 8135
rect -3155 8085 -3110 8135
rect -3060 8085 -3015 8135
rect -2965 8085 -2915 8135
rect -2865 8085 -2815 8135
rect -2765 8085 -2715 8135
rect -2665 8085 -2620 8135
rect -2570 8085 -2525 8135
rect -2475 8085 -2405 8135
rect -2355 8085 -2310 8135
rect -2260 8085 -2215 8135
rect -2165 8085 -2115 8135
rect -2065 8085 -2015 8135
rect -1965 8085 -1915 8135
rect -1865 8085 -1820 8135
rect -1770 8085 -1725 8135
rect -1675 8125 -80 8135
rect -40 8125 270 8165
rect 310 8125 620 8165
rect 660 8125 970 8165
rect 1010 8125 1670 8165
rect 1710 8125 2325 8165
rect 2365 8125 3175 8165
rect 3215 8125 3235 8165
rect 3275 8125 3345 8165
rect 3385 8125 6630 8165
rect 6670 8125 7270 8165
rect 7310 8125 7970 8165
rect 8010 8125 8320 8165
rect 8360 8125 8670 8165
rect 8710 8125 9020 8165
rect 9060 8125 9100 8165
rect -1675 8100 9100 8125
rect -1675 8085 -80 8100
rect -4840 8060 -80 8085
rect -40 8060 270 8100
rect 310 8060 620 8100
rect 660 8060 970 8100
rect 1010 8060 1670 8100
rect 1710 8060 2325 8100
rect 2365 8060 3175 8100
rect 3215 8060 3235 8100
rect 3275 8060 3345 8100
rect 3385 8060 6630 8100
rect 6670 8060 7270 8100
rect 7310 8060 7970 8100
rect 8010 8060 8320 8100
rect 8360 8060 8670 8100
rect 8710 8060 9020 8100
rect 9060 8060 9100 8100
rect -4840 8040 9100 8060
rect -4840 8015 -80 8040
rect -4840 7965 -4805 8015
rect -4755 7965 -4710 8015
rect -4660 7965 -4615 8015
rect -4565 7965 -4515 8015
rect -4465 7965 -4415 8015
rect -4365 7965 -4315 8015
rect -4265 7965 -4220 8015
rect -4170 7965 -4125 8015
rect -4075 7965 -4005 8015
rect -3955 7965 -3910 8015
rect -3860 7965 -3815 8015
rect -3765 7965 -3715 8015
rect -3665 7965 -3615 8015
rect -3565 7965 -3515 8015
rect -3465 7965 -3420 8015
rect -3370 7965 -3325 8015
rect -3275 7965 -3205 8015
rect -3155 7965 -3110 8015
rect -3060 7965 -3015 8015
rect -2965 7965 -2915 8015
rect -2865 7965 -2815 8015
rect -2765 7965 -2715 8015
rect -2665 7965 -2620 8015
rect -2570 7965 -2525 8015
rect -2475 7965 -2405 8015
rect -2355 7965 -2310 8015
rect -2260 7965 -2215 8015
rect -2165 7965 -2115 8015
rect -2065 7965 -2015 8015
rect -1965 7965 -1915 8015
rect -1865 7965 -1820 8015
rect -1770 7965 -1725 8015
rect -1675 8000 -80 8015
rect -40 8000 270 8040
rect 310 8000 620 8040
rect 660 8000 970 8040
rect 1010 8000 1670 8040
rect 1710 8000 2325 8040
rect 2365 8000 3175 8040
rect 3215 8000 3235 8040
rect 3275 8000 3345 8040
rect 3385 8000 6630 8040
rect 6670 8000 7270 8040
rect 7310 8000 7970 8040
rect 8010 8000 8320 8040
rect 8360 8000 8670 8040
rect 8710 8000 9020 8040
rect 9060 8000 9100 8040
rect -1675 7975 9100 8000
rect -1675 7965 -80 7975
rect -4840 7935 -80 7965
rect -40 7935 270 7975
rect 310 7935 620 7975
rect 660 7935 970 7975
rect 1010 7935 1670 7975
rect 1710 7935 2325 7975
rect 2365 7935 3175 7975
rect 3215 7935 3235 7975
rect 3275 7935 3345 7975
rect 3385 7935 6630 7975
rect 6670 7935 7270 7975
rect 7310 7935 7970 7975
rect 8010 7935 8320 7975
rect 8360 7935 8670 7975
rect 8710 7935 9020 7975
rect 9060 7935 9100 7975
rect -4840 7925 9100 7935
rect -4840 7875 -4805 7925
rect -4755 7875 -4710 7925
rect -4660 7875 -4615 7925
rect -4565 7875 -4515 7925
rect -4465 7875 -4415 7925
rect -4365 7875 -4315 7925
rect -4265 7875 -4220 7925
rect -4170 7875 -4125 7925
rect -4075 7875 -4005 7925
rect -3955 7875 -3910 7925
rect -3860 7875 -3815 7925
rect -3765 7875 -3715 7925
rect -3665 7875 -3615 7925
rect -3565 7875 -3515 7925
rect -3465 7875 -3420 7925
rect -3370 7875 -3325 7925
rect -3275 7875 -3205 7925
rect -3155 7875 -3110 7925
rect -3060 7875 -3015 7925
rect -2965 7875 -2915 7925
rect -2865 7875 -2815 7925
rect -2765 7875 -2715 7925
rect -2665 7875 -2620 7925
rect -2570 7875 -2525 7925
rect -2475 7875 -2405 7925
rect -2355 7875 -2310 7925
rect -2260 7875 -2215 7925
rect -2165 7875 -2115 7925
rect -2065 7875 -2015 7925
rect -1965 7875 -1915 7925
rect -1865 7875 -1820 7925
rect -1770 7875 -1725 7925
rect -1675 7905 9100 7925
rect -1675 7875 -80 7905
rect -4840 7865 -80 7875
rect -40 7865 270 7905
rect 310 7865 620 7905
rect 660 7865 970 7905
rect 1010 7865 1670 7905
rect 1710 7865 2325 7905
rect 2365 7865 3175 7905
rect 3215 7865 3235 7905
rect 3275 7865 3345 7905
rect 3385 7865 6630 7905
rect 6670 7865 7270 7905
rect 7310 7865 7970 7905
rect 8010 7865 8320 7905
rect 8360 7865 8670 7905
rect 8710 7865 9020 7905
rect 9060 7865 9100 7905
rect -4840 7835 9100 7865
rect -4840 7825 -80 7835
rect -4840 7775 -4805 7825
rect -4755 7775 -4710 7825
rect -4660 7775 -4615 7825
rect -4565 7775 -4515 7825
rect -4465 7775 -4415 7825
rect -4365 7775 -4315 7825
rect -4265 7775 -4220 7825
rect -4170 7775 -4125 7825
rect -4075 7775 -4005 7825
rect -3955 7775 -3910 7825
rect -3860 7775 -3815 7825
rect -3765 7775 -3715 7825
rect -3665 7775 -3615 7825
rect -3565 7775 -3515 7825
rect -3465 7775 -3420 7825
rect -3370 7775 -3325 7825
rect -3275 7775 -3205 7825
rect -3155 7775 -3110 7825
rect -3060 7775 -3015 7825
rect -2965 7775 -2915 7825
rect -2865 7775 -2815 7825
rect -2765 7775 -2715 7825
rect -2665 7775 -2620 7825
rect -2570 7775 -2525 7825
rect -2475 7775 -2405 7825
rect -2355 7775 -2310 7825
rect -2260 7775 -2215 7825
rect -2165 7775 -2115 7825
rect -2065 7775 -2015 7825
rect -1965 7775 -1915 7825
rect -1865 7775 -1820 7825
rect -1770 7775 -1725 7825
rect -1675 7795 -80 7825
rect -40 7795 270 7835
rect 310 7795 620 7835
rect 660 7795 970 7835
rect 1010 7795 1670 7835
rect 1710 7795 2325 7835
rect 2365 7795 3175 7835
rect 3215 7795 3235 7835
rect 3275 7795 3345 7835
rect 3385 7795 6630 7835
rect 6670 7795 7270 7835
rect 7310 7795 7970 7835
rect 8010 7795 8320 7835
rect 8360 7795 8670 7835
rect 8710 7795 9020 7835
rect 9060 7795 9100 7835
rect -1675 7775 9100 7795
rect -4840 7765 9100 7775
rect -4840 7735 -80 7765
rect -4840 7685 -4805 7735
rect -4755 7685 -4710 7735
rect -4660 7685 -4615 7735
rect -4565 7685 -4515 7735
rect -4465 7685 -4415 7735
rect -4365 7685 -4315 7735
rect -4265 7685 -4220 7735
rect -4170 7685 -4125 7735
rect -4075 7685 -4005 7735
rect -3955 7685 -3910 7735
rect -3860 7685 -3815 7735
rect -3765 7685 -3715 7735
rect -3665 7685 -3615 7735
rect -3565 7685 -3515 7735
rect -3465 7685 -3420 7735
rect -3370 7685 -3325 7735
rect -3275 7685 -3205 7735
rect -3155 7685 -3110 7735
rect -3060 7685 -3015 7735
rect -2965 7685 -2915 7735
rect -2865 7685 -2815 7735
rect -2765 7685 -2715 7735
rect -2665 7685 -2620 7735
rect -2570 7685 -2525 7735
rect -2475 7685 -2405 7735
rect -2355 7685 -2310 7735
rect -2260 7685 -2215 7735
rect -2165 7685 -2115 7735
rect -2065 7685 -2015 7735
rect -1965 7685 -1915 7735
rect -1865 7685 -1820 7735
rect -1770 7685 -1725 7735
rect -1675 7725 -80 7735
rect -40 7725 270 7765
rect 310 7725 620 7765
rect 660 7725 970 7765
rect 1010 7725 1670 7765
rect 1710 7725 2325 7765
rect 2365 7725 3175 7765
rect 3215 7725 3235 7765
rect 3275 7725 3345 7765
rect 3385 7725 6630 7765
rect 6670 7725 7270 7765
rect 7310 7725 7970 7765
rect 8010 7725 8320 7765
rect 8360 7725 8670 7765
rect 8710 7725 9020 7765
rect 9060 7725 9100 7765
rect -1675 7700 9100 7725
rect -1675 7685 -80 7700
rect -4840 7660 -80 7685
rect -40 7660 270 7700
rect 310 7660 620 7700
rect 660 7660 970 7700
rect 1010 7660 1670 7700
rect 1710 7660 2325 7700
rect 2365 7660 3175 7700
rect 3215 7660 3235 7700
rect 3275 7660 3345 7700
rect 3385 7660 6630 7700
rect 6670 7660 7270 7700
rect 7310 7660 7970 7700
rect 8010 7660 8320 7700
rect 8360 7660 8670 7700
rect 8710 7660 9020 7700
rect 9060 7660 9100 7700
rect -4840 7640 9100 7660
rect -4840 7615 -80 7640
rect -4840 7565 -4805 7615
rect -4755 7565 -4710 7615
rect -4660 7565 -4615 7615
rect -4565 7565 -4515 7615
rect -4465 7565 -4415 7615
rect -4365 7565 -4315 7615
rect -4265 7565 -4220 7615
rect -4170 7565 -4125 7615
rect -4075 7565 -4005 7615
rect -3955 7565 -3910 7615
rect -3860 7565 -3815 7615
rect -3765 7565 -3715 7615
rect -3665 7565 -3615 7615
rect -3565 7565 -3515 7615
rect -3465 7565 -3420 7615
rect -3370 7565 -3325 7615
rect -3275 7565 -3205 7615
rect -3155 7565 -3110 7615
rect -3060 7565 -3015 7615
rect -2965 7565 -2915 7615
rect -2865 7565 -2815 7615
rect -2765 7565 -2715 7615
rect -2665 7565 -2620 7615
rect -2570 7565 -2525 7615
rect -2475 7565 -2405 7615
rect -2355 7565 -2310 7615
rect -2260 7565 -2215 7615
rect -2165 7565 -2115 7615
rect -2065 7565 -2015 7615
rect -1965 7565 -1915 7615
rect -1865 7565 -1820 7615
rect -1770 7565 -1725 7615
rect -1675 7600 -80 7615
rect -40 7600 270 7640
rect 310 7600 620 7640
rect 660 7600 970 7640
rect 1010 7600 1670 7640
rect 1710 7600 2325 7640
rect 2365 7600 3175 7640
rect 3215 7600 3235 7640
rect 3275 7600 3345 7640
rect 3385 7600 6630 7640
rect 6670 7600 7270 7640
rect 7310 7600 7970 7640
rect 8010 7600 8320 7640
rect 8360 7600 8670 7640
rect 8710 7600 9020 7640
rect 9060 7600 9100 7640
rect -1675 7575 9100 7600
rect -1675 7565 -80 7575
rect -4840 7535 -80 7565
rect -40 7535 270 7575
rect 310 7535 620 7575
rect 660 7535 970 7575
rect 1010 7535 1670 7575
rect 1710 7535 2325 7575
rect 2365 7535 3175 7575
rect 3215 7535 3235 7575
rect 3275 7535 3345 7575
rect 3385 7535 6630 7575
rect 6670 7535 7270 7575
rect 7310 7535 7970 7575
rect 8010 7535 8320 7575
rect 8360 7535 8670 7575
rect 8710 7535 9020 7575
rect 9060 7535 9100 7575
rect -4840 7525 9100 7535
rect -4840 7475 -4805 7525
rect -4755 7475 -4710 7525
rect -4660 7475 -4615 7525
rect -4565 7475 -4515 7525
rect -4465 7475 -4415 7525
rect -4365 7475 -4315 7525
rect -4265 7475 -4220 7525
rect -4170 7475 -4125 7525
rect -4075 7475 -4005 7525
rect -3955 7475 -3910 7525
rect -3860 7475 -3815 7525
rect -3765 7475 -3715 7525
rect -3665 7475 -3615 7525
rect -3565 7475 -3515 7525
rect -3465 7475 -3420 7525
rect -3370 7475 -3325 7525
rect -3275 7475 -3205 7525
rect -3155 7475 -3110 7525
rect -3060 7475 -3015 7525
rect -2965 7475 -2915 7525
rect -2865 7475 -2815 7525
rect -2765 7475 -2715 7525
rect -2665 7475 -2620 7525
rect -2570 7475 -2525 7525
rect -2475 7475 -2405 7525
rect -2355 7475 -2310 7525
rect -2260 7475 -2215 7525
rect -2165 7475 -2115 7525
rect -2065 7475 -2015 7525
rect -1965 7475 -1915 7525
rect -1865 7475 -1820 7525
rect -1770 7475 -1725 7525
rect -1675 7505 9100 7525
rect -1675 7475 -80 7505
rect -4840 7465 -80 7475
rect -40 7465 270 7505
rect 310 7465 620 7505
rect 660 7465 970 7505
rect 1010 7465 1670 7505
rect 1710 7465 2325 7505
rect 2365 7465 3175 7505
rect 3215 7465 3235 7505
rect 3275 7465 3345 7505
rect 3385 7465 6630 7505
rect 6670 7465 7270 7505
rect 7310 7465 7970 7505
rect 8010 7465 8320 7505
rect 8360 7465 8670 7505
rect 8710 7465 9020 7505
rect 9060 7465 9100 7505
rect -4840 7435 9100 7465
rect -4840 7425 -80 7435
rect -4840 7375 -4805 7425
rect -4755 7375 -4710 7425
rect -4660 7375 -4615 7425
rect -4565 7375 -4515 7425
rect -4465 7375 -4415 7425
rect -4365 7375 -4315 7425
rect -4265 7375 -4220 7425
rect -4170 7375 -4125 7425
rect -4075 7375 -4005 7425
rect -3955 7375 -3910 7425
rect -3860 7375 -3815 7425
rect -3765 7375 -3715 7425
rect -3665 7375 -3615 7425
rect -3565 7375 -3515 7425
rect -3465 7375 -3420 7425
rect -3370 7375 -3325 7425
rect -3275 7375 -3205 7425
rect -3155 7375 -3110 7425
rect -3060 7375 -3015 7425
rect -2965 7375 -2915 7425
rect -2865 7375 -2815 7425
rect -2765 7375 -2715 7425
rect -2665 7375 -2620 7425
rect -2570 7375 -2525 7425
rect -2475 7375 -2405 7425
rect -2355 7375 -2310 7425
rect -2260 7375 -2215 7425
rect -2165 7375 -2115 7425
rect -2065 7375 -2015 7425
rect -1965 7375 -1915 7425
rect -1865 7375 -1820 7425
rect -1770 7375 -1725 7425
rect -1675 7395 -80 7425
rect -40 7395 270 7435
rect 310 7395 620 7435
rect 660 7395 970 7435
rect 1010 7395 1670 7435
rect 1710 7395 2325 7435
rect 2365 7395 3175 7435
rect 3215 7395 3235 7435
rect 3275 7395 3345 7435
rect 3385 7395 6630 7435
rect 6670 7395 7270 7435
rect 7310 7395 7970 7435
rect 8010 7395 8320 7435
rect 8360 7395 8670 7435
rect 8710 7395 9020 7435
rect 9060 7395 9100 7435
rect -1675 7375 9100 7395
rect -4840 7365 9100 7375
rect -4840 7335 -80 7365
rect -4840 7285 -4805 7335
rect -4755 7285 -4710 7335
rect -4660 7285 -4615 7335
rect -4565 7285 -4515 7335
rect -4465 7285 -4415 7335
rect -4365 7285 -4315 7335
rect -4265 7285 -4220 7335
rect -4170 7285 -4125 7335
rect -4075 7285 -4005 7335
rect -3955 7285 -3910 7335
rect -3860 7285 -3815 7335
rect -3765 7285 -3715 7335
rect -3665 7285 -3615 7335
rect -3565 7285 -3515 7335
rect -3465 7285 -3420 7335
rect -3370 7285 -3325 7335
rect -3275 7285 -3205 7335
rect -3155 7285 -3110 7335
rect -3060 7285 -3015 7335
rect -2965 7285 -2915 7335
rect -2865 7285 -2815 7335
rect -2765 7285 -2715 7335
rect -2665 7285 -2620 7335
rect -2570 7285 -2525 7335
rect -2475 7285 -2405 7335
rect -2355 7285 -2310 7335
rect -2260 7285 -2215 7335
rect -2165 7285 -2115 7335
rect -2065 7285 -2015 7335
rect -1965 7285 -1915 7335
rect -1865 7285 -1820 7335
rect -1770 7285 -1725 7335
rect -1675 7325 -80 7335
rect -40 7325 270 7365
rect 310 7325 620 7365
rect 660 7325 970 7365
rect 1010 7325 1670 7365
rect 1710 7325 2325 7365
rect 2365 7325 3175 7365
rect 3215 7325 3235 7365
rect 3275 7325 3345 7365
rect 3385 7325 6630 7365
rect 6670 7325 7270 7365
rect 7310 7325 7970 7365
rect 8010 7325 8320 7365
rect 8360 7325 8670 7365
rect 8710 7325 9020 7365
rect 9060 7325 9100 7365
rect -1675 7300 9100 7325
rect -1675 7285 -80 7300
rect -4840 7260 -80 7285
rect -40 7260 270 7300
rect 310 7260 620 7300
rect 660 7260 970 7300
rect 1010 7260 1670 7300
rect 1710 7260 2325 7300
rect 2365 7260 3175 7300
rect 3215 7260 3235 7300
rect 3275 7260 3345 7300
rect 3385 7260 6630 7300
rect 6670 7260 7270 7300
rect 7310 7260 7970 7300
rect 8010 7260 8320 7300
rect 8360 7260 8670 7300
rect 8710 7260 9020 7300
rect 9060 7260 9100 7300
rect -4840 7240 9100 7260
rect -4840 7215 -80 7240
rect -4840 7165 -4805 7215
rect -4755 7165 -4710 7215
rect -4660 7165 -4615 7215
rect -4565 7165 -4515 7215
rect -4465 7165 -4415 7215
rect -4365 7165 -4315 7215
rect -4265 7165 -4220 7215
rect -4170 7165 -4125 7215
rect -4075 7165 -4005 7215
rect -3955 7165 -3910 7215
rect -3860 7165 -3815 7215
rect -3765 7165 -3715 7215
rect -3665 7165 -3615 7215
rect -3565 7165 -3515 7215
rect -3465 7165 -3420 7215
rect -3370 7165 -3325 7215
rect -3275 7165 -3205 7215
rect -3155 7165 -3110 7215
rect -3060 7165 -3015 7215
rect -2965 7165 -2915 7215
rect -2865 7165 -2815 7215
rect -2765 7165 -2715 7215
rect -2665 7165 -2620 7215
rect -2570 7165 -2525 7215
rect -2475 7165 -2405 7215
rect -2355 7165 -2310 7215
rect -2260 7165 -2215 7215
rect -2165 7165 -2115 7215
rect -2065 7165 -2015 7215
rect -1965 7165 -1915 7215
rect -1865 7165 -1820 7215
rect -1770 7165 -1725 7215
rect -1675 7200 -80 7215
rect -40 7200 270 7240
rect 310 7200 620 7240
rect 660 7200 970 7240
rect 1010 7200 1670 7240
rect 1710 7200 2325 7240
rect 2365 7200 3175 7240
rect 3215 7200 3235 7240
rect 3275 7200 3345 7240
rect 3385 7200 6630 7240
rect 6670 7200 7270 7240
rect 7310 7200 7970 7240
rect 8010 7200 8320 7240
rect 8360 7200 8670 7240
rect 8710 7200 9020 7240
rect 9060 7200 9100 7240
rect -1675 7175 9100 7200
rect -1675 7165 -80 7175
rect -4840 7135 -80 7165
rect -40 7135 270 7175
rect 310 7135 620 7175
rect 660 7135 970 7175
rect 1010 7135 1670 7175
rect 1710 7135 2325 7175
rect 2365 7135 3175 7175
rect 3215 7135 3235 7175
rect 3275 7135 3345 7175
rect 3385 7135 6630 7175
rect 6670 7135 7270 7175
rect 7310 7135 7970 7175
rect 8010 7135 8320 7175
rect 8360 7135 8670 7175
rect 8710 7135 9020 7175
rect 9060 7135 9100 7175
rect -4840 7125 9100 7135
rect -4840 7075 -4805 7125
rect -4755 7075 -4710 7125
rect -4660 7075 -4615 7125
rect -4565 7075 -4515 7125
rect -4465 7075 -4415 7125
rect -4365 7075 -4315 7125
rect -4265 7075 -4220 7125
rect -4170 7075 -4125 7125
rect -4075 7075 -4005 7125
rect -3955 7075 -3910 7125
rect -3860 7075 -3815 7125
rect -3765 7075 -3715 7125
rect -3665 7075 -3615 7125
rect -3565 7075 -3515 7125
rect -3465 7075 -3420 7125
rect -3370 7075 -3325 7125
rect -3275 7075 -3205 7125
rect -3155 7075 -3110 7125
rect -3060 7075 -3015 7125
rect -2965 7075 -2915 7125
rect -2865 7075 -2815 7125
rect -2765 7075 -2715 7125
rect -2665 7075 -2620 7125
rect -2570 7075 -2525 7125
rect -2475 7075 -2405 7125
rect -2355 7075 -2310 7125
rect -2260 7075 -2215 7125
rect -2165 7075 -2115 7125
rect -2065 7075 -2015 7125
rect -1965 7075 -1915 7125
rect -1865 7075 -1820 7125
rect -1770 7075 -1725 7125
rect -1675 7105 9100 7125
rect -1675 7075 -80 7105
rect -4840 7065 -80 7075
rect -40 7065 270 7105
rect 310 7065 620 7105
rect 660 7065 970 7105
rect 1010 7065 1670 7105
rect 1710 7065 2325 7105
rect 2365 7065 3175 7105
rect 3215 7065 3235 7105
rect 3275 7065 3345 7105
rect 3385 7065 6630 7105
rect 6670 7065 7270 7105
rect 7310 7065 7970 7105
rect 8010 7065 8320 7105
rect 8360 7065 8670 7105
rect 8710 7065 9020 7105
rect 9060 7065 9100 7105
rect -4840 7035 9100 7065
rect -4840 7025 -80 7035
rect -4840 6975 -4805 7025
rect -4755 6975 -4710 7025
rect -4660 6975 -4615 7025
rect -4565 6975 -4515 7025
rect -4465 6975 -4415 7025
rect -4365 6975 -4315 7025
rect -4265 6975 -4220 7025
rect -4170 6975 -4125 7025
rect -4075 6975 -4005 7025
rect -3955 6975 -3910 7025
rect -3860 6975 -3815 7025
rect -3765 6975 -3715 7025
rect -3665 6975 -3615 7025
rect -3565 6975 -3515 7025
rect -3465 6975 -3420 7025
rect -3370 6975 -3325 7025
rect -3275 6975 -3205 7025
rect -3155 6975 -3110 7025
rect -3060 6975 -3015 7025
rect -2965 6975 -2915 7025
rect -2865 6975 -2815 7025
rect -2765 6975 -2715 7025
rect -2665 6975 -2620 7025
rect -2570 6975 -2525 7025
rect -2475 6975 -2405 7025
rect -2355 6975 -2310 7025
rect -2260 6975 -2215 7025
rect -2165 6975 -2115 7025
rect -2065 6975 -2015 7025
rect -1965 6975 -1915 7025
rect -1865 6975 -1820 7025
rect -1770 6975 -1725 7025
rect -1675 6995 -80 7025
rect -40 6995 270 7035
rect 310 6995 620 7035
rect 660 6995 970 7035
rect 1010 6995 1670 7035
rect 1710 6995 2325 7035
rect 2365 6995 3175 7035
rect 3215 6995 3235 7035
rect 3275 6995 3345 7035
rect 3385 6995 6630 7035
rect 6670 6995 7270 7035
rect 7310 6995 7970 7035
rect 8010 6995 8320 7035
rect 8360 6995 8670 7035
rect 8710 6995 9020 7035
rect 9060 6995 9100 7035
rect -1675 6975 9100 6995
rect -4840 6965 9100 6975
rect -4840 6935 -80 6965
rect -4840 6885 -4805 6935
rect -4755 6885 -4710 6935
rect -4660 6885 -4615 6935
rect -4565 6885 -4515 6935
rect -4465 6885 -4415 6935
rect -4365 6885 -4315 6935
rect -4265 6885 -4220 6935
rect -4170 6885 -4125 6935
rect -4075 6885 -4005 6935
rect -3955 6885 -3910 6935
rect -3860 6885 -3815 6935
rect -3765 6885 -3715 6935
rect -3665 6885 -3615 6935
rect -3565 6885 -3515 6935
rect -3465 6885 -3420 6935
rect -3370 6885 -3325 6935
rect -3275 6885 -3205 6935
rect -3155 6885 -3110 6935
rect -3060 6885 -3015 6935
rect -2965 6885 -2915 6935
rect -2865 6885 -2815 6935
rect -2765 6885 -2715 6935
rect -2665 6885 -2620 6935
rect -2570 6885 -2525 6935
rect -2475 6885 -2405 6935
rect -2355 6885 -2310 6935
rect -2260 6885 -2215 6935
rect -2165 6885 -2115 6935
rect -2065 6885 -2015 6935
rect -1965 6885 -1915 6935
rect -1865 6885 -1820 6935
rect -1770 6885 -1725 6935
rect -1675 6925 -80 6935
rect -40 6925 270 6965
rect 310 6925 620 6965
rect 660 6925 970 6965
rect 1010 6925 1670 6965
rect 1710 6925 2325 6965
rect 2365 6925 3175 6965
rect 3215 6925 3235 6965
rect 3275 6925 3345 6965
rect 3385 6925 6630 6965
rect 6670 6925 7270 6965
rect 7310 6925 7970 6965
rect 8010 6925 8320 6965
rect 8360 6925 8670 6965
rect 8710 6925 9020 6965
rect 9060 6925 9100 6965
rect -1675 6900 9100 6925
rect -1675 6885 -80 6900
rect -4840 6860 -80 6885
rect -40 6860 270 6900
rect 310 6860 620 6900
rect 660 6860 970 6900
rect 1010 6860 1670 6900
rect 1710 6860 2325 6900
rect 2365 6860 3175 6900
rect 3215 6860 3235 6900
rect 3275 6860 3345 6900
rect 3385 6860 6630 6900
rect 6670 6860 7270 6900
rect 7310 6860 7970 6900
rect 8010 6860 8320 6900
rect 8360 6860 8670 6900
rect 8710 6860 9020 6900
rect 9060 6860 9100 6900
rect -4840 6840 9100 6860
rect -4840 6815 -80 6840
rect -4840 6765 -4805 6815
rect -4755 6765 -4710 6815
rect -4660 6765 -4615 6815
rect -4565 6765 -4515 6815
rect -4465 6765 -4415 6815
rect -4365 6765 -4315 6815
rect -4265 6765 -4220 6815
rect -4170 6765 -4125 6815
rect -4075 6765 -4005 6815
rect -3955 6765 -3910 6815
rect -3860 6765 -3815 6815
rect -3765 6765 -3715 6815
rect -3665 6765 -3615 6815
rect -3565 6765 -3515 6815
rect -3465 6765 -3420 6815
rect -3370 6765 -3325 6815
rect -3275 6765 -3205 6815
rect -3155 6765 -3110 6815
rect -3060 6765 -3015 6815
rect -2965 6765 -2915 6815
rect -2865 6765 -2815 6815
rect -2765 6765 -2715 6815
rect -2665 6765 -2620 6815
rect -2570 6765 -2525 6815
rect -2475 6765 -2405 6815
rect -2355 6765 -2310 6815
rect -2260 6765 -2215 6815
rect -2165 6765 -2115 6815
rect -2065 6765 -2015 6815
rect -1965 6765 -1915 6815
rect -1865 6765 -1820 6815
rect -1770 6765 -1725 6815
rect -1675 6800 -80 6815
rect -40 6800 270 6840
rect 310 6800 620 6840
rect 660 6800 970 6840
rect 1010 6800 1670 6840
rect 1710 6800 2325 6840
rect 2365 6800 3175 6840
rect 3215 6800 3235 6840
rect 3275 6800 3345 6840
rect 3385 6800 6630 6840
rect 6670 6800 7270 6840
rect 7310 6800 7970 6840
rect 8010 6800 8320 6840
rect 8360 6800 8670 6840
rect 8710 6800 9020 6840
rect 9060 6800 9100 6840
rect -1675 6775 9100 6800
rect -1675 6765 -80 6775
rect -4840 6735 -80 6765
rect -40 6735 270 6775
rect 310 6735 620 6775
rect 660 6735 970 6775
rect 1010 6735 1670 6775
rect 1710 6735 2325 6775
rect 2365 6735 3175 6775
rect 3215 6735 3235 6775
rect 3275 6735 3345 6775
rect 3385 6735 6630 6775
rect 6670 6735 7270 6775
rect 7310 6735 7970 6775
rect 8010 6735 8320 6775
rect 8360 6735 8670 6775
rect 8710 6735 9020 6775
rect 9060 6735 9100 6775
rect -4840 6725 9100 6735
rect -4840 6675 -4805 6725
rect -4755 6675 -4710 6725
rect -4660 6675 -4615 6725
rect -4565 6675 -4515 6725
rect -4465 6675 -4415 6725
rect -4365 6675 -4315 6725
rect -4265 6675 -4220 6725
rect -4170 6675 -4125 6725
rect -4075 6675 -4005 6725
rect -3955 6675 -3910 6725
rect -3860 6675 -3815 6725
rect -3765 6675 -3715 6725
rect -3665 6675 -3615 6725
rect -3565 6675 -3515 6725
rect -3465 6675 -3420 6725
rect -3370 6675 -3325 6725
rect -3275 6675 -3205 6725
rect -3155 6675 -3110 6725
rect -3060 6675 -3015 6725
rect -2965 6675 -2915 6725
rect -2865 6675 -2815 6725
rect -2765 6675 -2715 6725
rect -2665 6675 -2620 6725
rect -2570 6675 -2525 6725
rect -2475 6675 -2405 6725
rect -2355 6675 -2310 6725
rect -2260 6675 -2215 6725
rect -2165 6675 -2115 6725
rect -2065 6675 -2015 6725
rect -1965 6675 -1915 6725
rect -1865 6675 -1820 6725
rect -1770 6675 -1725 6725
rect -1675 6705 9100 6725
rect -1675 6675 -80 6705
rect -4840 6665 -80 6675
rect -40 6665 270 6705
rect 310 6665 620 6705
rect 660 6665 970 6705
rect 1010 6665 1670 6705
rect 1710 6665 2325 6705
rect 2365 6665 3175 6705
rect 3215 6665 3235 6705
rect 3275 6665 3345 6705
rect 3385 6665 6630 6705
rect 6670 6665 7270 6705
rect 7310 6665 7970 6705
rect 8010 6665 8320 6705
rect 8360 6665 8670 6705
rect 8710 6665 9020 6705
rect 9060 6665 9100 6705
rect -4840 6635 9100 6665
rect -4840 6625 -80 6635
rect -4840 6575 -4805 6625
rect -4755 6575 -4710 6625
rect -4660 6575 -4615 6625
rect -4565 6575 -4515 6625
rect -4465 6575 -4415 6625
rect -4365 6575 -4315 6625
rect -4265 6575 -4220 6625
rect -4170 6575 -4125 6625
rect -4075 6575 -4005 6625
rect -3955 6575 -3910 6625
rect -3860 6575 -3815 6625
rect -3765 6575 -3715 6625
rect -3665 6575 -3615 6625
rect -3565 6575 -3515 6625
rect -3465 6575 -3420 6625
rect -3370 6575 -3325 6625
rect -3275 6575 -3205 6625
rect -3155 6575 -3110 6625
rect -3060 6575 -3015 6625
rect -2965 6575 -2915 6625
rect -2865 6575 -2815 6625
rect -2765 6575 -2715 6625
rect -2665 6575 -2620 6625
rect -2570 6575 -2525 6625
rect -2475 6575 -2405 6625
rect -2355 6575 -2310 6625
rect -2260 6575 -2215 6625
rect -2165 6575 -2115 6625
rect -2065 6575 -2015 6625
rect -1965 6575 -1915 6625
rect -1865 6575 -1820 6625
rect -1770 6575 -1725 6625
rect -1675 6595 -80 6625
rect -40 6595 270 6635
rect 310 6595 620 6635
rect 660 6595 970 6635
rect 1010 6595 1670 6635
rect 1710 6595 2325 6635
rect 2365 6595 3175 6635
rect 3215 6595 3235 6635
rect 3275 6595 3345 6635
rect 3385 6595 6630 6635
rect 6670 6595 7270 6635
rect 7310 6595 7970 6635
rect 8010 6595 8320 6635
rect 8360 6595 8670 6635
rect 8710 6595 9020 6635
rect 9060 6595 9100 6635
rect -1675 6575 9100 6595
rect -4840 6565 9100 6575
rect -4840 6535 -80 6565
rect -4840 6485 -4805 6535
rect -4755 6485 -4710 6535
rect -4660 6485 -4615 6535
rect -4565 6485 -4515 6535
rect -4465 6485 -4415 6535
rect -4365 6485 -4315 6535
rect -4265 6485 -4220 6535
rect -4170 6485 -4125 6535
rect -4075 6485 -4005 6535
rect -3955 6485 -3910 6535
rect -3860 6485 -3815 6535
rect -3765 6485 -3715 6535
rect -3665 6485 -3615 6535
rect -3565 6485 -3515 6535
rect -3465 6485 -3420 6535
rect -3370 6485 -3325 6535
rect -3275 6485 -3205 6535
rect -3155 6485 -3110 6535
rect -3060 6485 -3015 6535
rect -2965 6485 -2915 6535
rect -2865 6485 -2815 6535
rect -2765 6485 -2715 6535
rect -2665 6485 -2620 6535
rect -2570 6485 -2525 6535
rect -2475 6485 -2405 6535
rect -2355 6485 -2310 6535
rect -2260 6485 -2215 6535
rect -2165 6485 -2115 6535
rect -2065 6485 -2015 6535
rect -1965 6485 -1915 6535
rect -1865 6485 -1820 6535
rect -1770 6485 -1725 6535
rect -1675 6525 -80 6535
rect -40 6525 270 6565
rect 310 6525 620 6565
rect 660 6525 970 6565
rect 1010 6525 1670 6565
rect 1710 6525 2325 6565
rect 2365 6525 3175 6565
rect 3215 6525 3235 6565
rect 3275 6525 3345 6565
rect 3385 6525 6630 6565
rect 6670 6525 7270 6565
rect 7310 6525 7970 6565
rect 8010 6525 8320 6565
rect 8360 6525 8670 6565
rect 8710 6525 9020 6565
rect 9060 6525 9100 6565
rect -1675 6500 9100 6525
rect -1675 6485 -80 6500
rect -4840 6460 -80 6485
rect -40 6460 270 6500
rect 310 6460 620 6500
rect 660 6460 970 6500
rect 1010 6460 1670 6500
rect 1710 6460 2325 6500
rect 2365 6460 3175 6500
rect 3215 6460 3235 6500
rect 3275 6460 3345 6500
rect 3385 6460 6630 6500
rect 6670 6460 7270 6500
rect 7310 6460 7970 6500
rect 8010 6460 8320 6500
rect 8360 6460 8670 6500
rect 8710 6460 9020 6500
rect 9060 6460 9100 6500
rect -4840 6450 9100 6460
rect 12890 9615 18820 9650
rect 12890 9565 12925 9615
rect 12975 9565 13020 9615
rect 13070 9565 13115 9615
rect 13165 9565 13215 9615
rect 13265 9565 13315 9615
rect 13365 9565 13415 9615
rect 13465 9565 13510 9615
rect 13560 9565 13605 9615
rect 13655 9565 13725 9615
rect 13775 9565 13820 9615
rect 13870 9565 13915 9615
rect 13965 9565 14015 9615
rect 14065 9565 14115 9615
rect 14165 9565 14215 9615
rect 14265 9565 14310 9615
rect 14360 9565 14405 9615
rect 14455 9565 14525 9615
rect 14575 9565 14620 9615
rect 14670 9565 14715 9615
rect 14765 9565 14815 9615
rect 14865 9565 14915 9615
rect 14965 9565 15015 9615
rect 15065 9565 15110 9615
rect 15160 9565 15205 9615
rect 15255 9565 15325 9615
rect 15375 9565 15420 9615
rect 15470 9565 15515 9615
rect 15565 9565 15615 9615
rect 15665 9565 15715 9615
rect 15765 9565 15815 9615
rect 15865 9565 15910 9615
rect 15960 9565 16005 9615
rect 16055 9565 18820 9615
rect 12890 9525 18820 9565
rect 12890 9475 12925 9525
rect 12975 9475 13020 9525
rect 13070 9475 13115 9525
rect 13165 9475 13215 9525
rect 13265 9475 13315 9525
rect 13365 9475 13415 9525
rect 13465 9475 13510 9525
rect 13560 9475 13605 9525
rect 13655 9475 13725 9525
rect 13775 9475 13820 9525
rect 13870 9475 13915 9525
rect 13965 9475 14015 9525
rect 14065 9475 14115 9525
rect 14165 9475 14215 9525
rect 14265 9475 14310 9525
rect 14360 9475 14405 9525
rect 14455 9475 14525 9525
rect 14575 9475 14620 9525
rect 14670 9475 14715 9525
rect 14765 9475 14815 9525
rect 14865 9475 14915 9525
rect 14965 9475 15015 9525
rect 15065 9475 15110 9525
rect 15160 9475 15205 9525
rect 15255 9475 15325 9525
rect 15375 9475 15420 9525
rect 15470 9475 15515 9525
rect 15565 9475 15615 9525
rect 15665 9475 15715 9525
rect 15765 9475 15815 9525
rect 15865 9475 15910 9525
rect 15960 9475 16005 9525
rect 16055 9475 18820 9525
rect 12890 9425 18820 9475
rect 12890 9375 12925 9425
rect 12975 9375 13020 9425
rect 13070 9375 13115 9425
rect 13165 9375 13215 9425
rect 13265 9375 13315 9425
rect 13365 9375 13415 9425
rect 13465 9375 13510 9425
rect 13560 9375 13605 9425
rect 13655 9375 13725 9425
rect 13775 9375 13820 9425
rect 13870 9375 13915 9425
rect 13965 9375 14015 9425
rect 14065 9375 14115 9425
rect 14165 9375 14215 9425
rect 14265 9375 14310 9425
rect 14360 9375 14405 9425
rect 14455 9375 14525 9425
rect 14575 9375 14620 9425
rect 14670 9375 14715 9425
rect 14765 9375 14815 9425
rect 14865 9375 14915 9425
rect 14965 9375 15015 9425
rect 15065 9375 15110 9425
rect 15160 9375 15205 9425
rect 15255 9375 15325 9425
rect 15375 9375 15420 9425
rect 15470 9375 15515 9425
rect 15565 9375 15615 9425
rect 15665 9375 15715 9425
rect 15765 9375 15815 9425
rect 15865 9375 15910 9425
rect 15960 9375 16005 9425
rect 16055 9375 18820 9425
rect 12890 9335 18820 9375
rect 12890 9285 12925 9335
rect 12975 9285 13020 9335
rect 13070 9285 13115 9335
rect 13165 9285 13215 9335
rect 13265 9285 13315 9335
rect 13365 9285 13415 9335
rect 13465 9285 13510 9335
rect 13560 9285 13605 9335
rect 13655 9285 13725 9335
rect 13775 9285 13820 9335
rect 13870 9285 13915 9335
rect 13965 9285 14015 9335
rect 14065 9285 14115 9335
rect 14165 9285 14215 9335
rect 14265 9285 14310 9335
rect 14360 9285 14405 9335
rect 14455 9285 14525 9335
rect 14575 9285 14620 9335
rect 14670 9285 14715 9335
rect 14765 9285 14815 9335
rect 14865 9285 14915 9335
rect 14965 9285 15015 9335
rect 15065 9285 15110 9335
rect 15160 9285 15205 9335
rect 15255 9285 15325 9335
rect 15375 9285 15420 9335
rect 15470 9285 15515 9335
rect 15565 9285 15615 9335
rect 15665 9285 15715 9335
rect 15765 9285 15815 9335
rect 15865 9285 15910 9335
rect 15960 9285 16005 9335
rect 16055 9285 18820 9335
rect 12890 9215 18820 9285
rect 12890 9165 12925 9215
rect 12975 9165 13020 9215
rect 13070 9165 13115 9215
rect 13165 9165 13215 9215
rect 13265 9165 13315 9215
rect 13365 9165 13415 9215
rect 13465 9165 13510 9215
rect 13560 9165 13605 9215
rect 13655 9165 13725 9215
rect 13775 9165 13820 9215
rect 13870 9165 13915 9215
rect 13965 9165 14015 9215
rect 14065 9165 14115 9215
rect 14165 9165 14215 9215
rect 14265 9165 14310 9215
rect 14360 9165 14405 9215
rect 14455 9165 14525 9215
rect 14575 9165 14620 9215
rect 14670 9165 14715 9215
rect 14765 9165 14815 9215
rect 14865 9165 14915 9215
rect 14965 9165 15015 9215
rect 15065 9165 15110 9215
rect 15160 9165 15205 9215
rect 15255 9165 15325 9215
rect 15375 9165 15420 9215
rect 15470 9165 15515 9215
rect 15565 9165 15615 9215
rect 15665 9165 15715 9215
rect 15765 9165 15815 9215
rect 15865 9165 15910 9215
rect 15960 9165 16005 9215
rect 16055 9165 18820 9215
rect 12890 9125 18820 9165
rect 12890 9075 12925 9125
rect 12975 9075 13020 9125
rect 13070 9075 13115 9125
rect 13165 9075 13215 9125
rect 13265 9075 13315 9125
rect 13365 9075 13415 9125
rect 13465 9075 13510 9125
rect 13560 9075 13605 9125
rect 13655 9075 13725 9125
rect 13775 9075 13820 9125
rect 13870 9075 13915 9125
rect 13965 9075 14015 9125
rect 14065 9075 14115 9125
rect 14165 9075 14215 9125
rect 14265 9075 14310 9125
rect 14360 9075 14405 9125
rect 14455 9075 14525 9125
rect 14575 9075 14620 9125
rect 14670 9075 14715 9125
rect 14765 9075 14815 9125
rect 14865 9075 14915 9125
rect 14965 9075 15015 9125
rect 15065 9075 15110 9125
rect 15160 9075 15205 9125
rect 15255 9075 15325 9125
rect 15375 9075 15420 9125
rect 15470 9075 15515 9125
rect 15565 9075 15615 9125
rect 15665 9075 15715 9125
rect 15765 9075 15815 9125
rect 15865 9075 15910 9125
rect 15960 9075 16005 9125
rect 16055 9075 18820 9125
rect 12890 9025 18820 9075
rect 12890 8975 12925 9025
rect 12975 8975 13020 9025
rect 13070 8975 13115 9025
rect 13165 8975 13215 9025
rect 13265 8975 13315 9025
rect 13365 8975 13415 9025
rect 13465 8975 13510 9025
rect 13560 8975 13605 9025
rect 13655 8975 13725 9025
rect 13775 8975 13820 9025
rect 13870 8975 13915 9025
rect 13965 8975 14015 9025
rect 14065 8975 14115 9025
rect 14165 8975 14215 9025
rect 14265 8975 14310 9025
rect 14360 8975 14405 9025
rect 14455 8975 14525 9025
rect 14575 8975 14620 9025
rect 14670 8975 14715 9025
rect 14765 8975 14815 9025
rect 14865 8975 14915 9025
rect 14965 8975 15015 9025
rect 15065 8975 15110 9025
rect 15160 8975 15205 9025
rect 15255 8975 15325 9025
rect 15375 8975 15420 9025
rect 15470 8975 15515 9025
rect 15565 8975 15615 9025
rect 15665 8975 15715 9025
rect 15765 8975 15815 9025
rect 15865 8975 15910 9025
rect 15960 8975 16005 9025
rect 16055 8975 18820 9025
rect 12890 8935 18820 8975
rect 12890 8885 12925 8935
rect 12975 8885 13020 8935
rect 13070 8885 13115 8935
rect 13165 8885 13215 8935
rect 13265 8885 13315 8935
rect 13365 8885 13415 8935
rect 13465 8885 13510 8935
rect 13560 8885 13605 8935
rect 13655 8885 13725 8935
rect 13775 8885 13820 8935
rect 13870 8885 13915 8935
rect 13965 8885 14015 8935
rect 14065 8885 14115 8935
rect 14165 8885 14215 8935
rect 14265 8885 14310 8935
rect 14360 8885 14405 8935
rect 14455 8885 14525 8935
rect 14575 8885 14620 8935
rect 14670 8885 14715 8935
rect 14765 8885 14815 8935
rect 14865 8885 14915 8935
rect 14965 8885 15015 8935
rect 15065 8885 15110 8935
rect 15160 8885 15205 8935
rect 15255 8885 15325 8935
rect 15375 8885 15420 8935
rect 15470 8885 15515 8935
rect 15565 8885 15615 8935
rect 15665 8885 15715 8935
rect 15765 8885 15815 8935
rect 15865 8885 15910 8935
rect 15960 8885 16005 8935
rect 16055 8885 18820 8935
rect 12890 8815 18820 8885
rect 12890 8765 12925 8815
rect 12975 8765 13020 8815
rect 13070 8765 13115 8815
rect 13165 8765 13215 8815
rect 13265 8765 13315 8815
rect 13365 8765 13415 8815
rect 13465 8765 13510 8815
rect 13560 8765 13605 8815
rect 13655 8765 13725 8815
rect 13775 8765 13820 8815
rect 13870 8765 13915 8815
rect 13965 8765 14015 8815
rect 14065 8765 14115 8815
rect 14165 8765 14215 8815
rect 14265 8765 14310 8815
rect 14360 8765 14405 8815
rect 14455 8765 14525 8815
rect 14575 8765 14620 8815
rect 14670 8765 14715 8815
rect 14765 8765 14815 8815
rect 14865 8765 14915 8815
rect 14965 8765 15015 8815
rect 15065 8765 15110 8815
rect 15160 8765 15205 8815
rect 15255 8765 15325 8815
rect 15375 8765 15420 8815
rect 15470 8765 15515 8815
rect 15565 8765 15615 8815
rect 15665 8765 15715 8815
rect 15765 8765 15815 8815
rect 15865 8765 15910 8815
rect 15960 8765 16005 8815
rect 16055 8765 18820 8815
rect 12890 8725 18820 8765
rect 12890 8675 12925 8725
rect 12975 8675 13020 8725
rect 13070 8675 13115 8725
rect 13165 8675 13215 8725
rect 13265 8675 13315 8725
rect 13365 8675 13415 8725
rect 13465 8675 13510 8725
rect 13560 8675 13605 8725
rect 13655 8675 13725 8725
rect 13775 8675 13820 8725
rect 13870 8675 13915 8725
rect 13965 8675 14015 8725
rect 14065 8675 14115 8725
rect 14165 8675 14215 8725
rect 14265 8675 14310 8725
rect 14360 8675 14405 8725
rect 14455 8675 14525 8725
rect 14575 8675 14620 8725
rect 14670 8675 14715 8725
rect 14765 8675 14815 8725
rect 14865 8675 14915 8725
rect 14965 8675 15015 8725
rect 15065 8675 15110 8725
rect 15160 8675 15205 8725
rect 15255 8675 15325 8725
rect 15375 8675 15420 8725
rect 15470 8675 15515 8725
rect 15565 8675 15615 8725
rect 15665 8675 15715 8725
rect 15765 8675 15815 8725
rect 15865 8675 15910 8725
rect 15960 8675 16005 8725
rect 16055 8675 18820 8725
rect 12890 8625 18820 8675
rect 12890 8575 12925 8625
rect 12975 8575 13020 8625
rect 13070 8575 13115 8625
rect 13165 8575 13215 8625
rect 13265 8575 13315 8625
rect 13365 8575 13415 8625
rect 13465 8575 13510 8625
rect 13560 8575 13605 8625
rect 13655 8575 13725 8625
rect 13775 8575 13820 8625
rect 13870 8575 13915 8625
rect 13965 8575 14015 8625
rect 14065 8575 14115 8625
rect 14165 8575 14215 8625
rect 14265 8575 14310 8625
rect 14360 8575 14405 8625
rect 14455 8575 14525 8625
rect 14575 8575 14620 8625
rect 14670 8575 14715 8625
rect 14765 8575 14815 8625
rect 14865 8575 14915 8625
rect 14965 8575 15015 8625
rect 15065 8575 15110 8625
rect 15160 8575 15205 8625
rect 15255 8575 15325 8625
rect 15375 8575 15420 8625
rect 15470 8575 15515 8625
rect 15565 8575 15615 8625
rect 15665 8575 15715 8625
rect 15765 8575 15815 8625
rect 15865 8575 15910 8625
rect 15960 8575 16005 8625
rect 16055 8575 18820 8625
rect 12890 8535 18820 8575
rect 12890 8485 12925 8535
rect 12975 8485 13020 8535
rect 13070 8485 13115 8535
rect 13165 8485 13215 8535
rect 13265 8485 13315 8535
rect 13365 8485 13415 8535
rect 13465 8485 13510 8535
rect 13560 8485 13605 8535
rect 13655 8485 13725 8535
rect 13775 8485 13820 8535
rect 13870 8485 13915 8535
rect 13965 8485 14015 8535
rect 14065 8485 14115 8535
rect 14165 8485 14215 8535
rect 14265 8485 14310 8535
rect 14360 8485 14405 8535
rect 14455 8485 14525 8535
rect 14575 8485 14620 8535
rect 14670 8485 14715 8535
rect 14765 8485 14815 8535
rect 14865 8485 14915 8535
rect 14965 8485 15015 8535
rect 15065 8485 15110 8535
rect 15160 8485 15205 8535
rect 15255 8485 15325 8535
rect 15375 8485 15420 8535
rect 15470 8485 15515 8535
rect 15565 8485 15615 8535
rect 15665 8485 15715 8535
rect 15765 8485 15815 8535
rect 15865 8485 15910 8535
rect 15960 8485 16005 8535
rect 16055 8485 18820 8535
rect 12890 8415 18820 8485
rect 12890 8365 12925 8415
rect 12975 8365 13020 8415
rect 13070 8365 13115 8415
rect 13165 8365 13215 8415
rect 13265 8365 13315 8415
rect 13365 8365 13415 8415
rect 13465 8365 13510 8415
rect 13560 8365 13605 8415
rect 13655 8365 13725 8415
rect 13775 8365 13820 8415
rect 13870 8365 13915 8415
rect 13965 8365 14015 8415
rect 14065 8365 14115 8415
rect 14165 8365 14215 8415
rect 14265 8365 14310 8415
rect 14360 8365 14405 8415
rect 14455 8365 14525 8415
rect 14575 8365 14620 8415
rect 14670 8365 14715 8415
rect 14765 8365 14815 8415
rect 14865 8365 14915 8415
rect 14965 8365 15015 8415
rect 15065 8365 15110 8415
rect 15160 8365 15205 8415
rect 15255 8365 15325 8415
rect 15375 8365 15420 8415
rect 15470 8365 15515 8415
rect 15565 8365 15615 8415
rect 15665 8365 15715 8415
rect 15765 8365 15815 8415
rect 15865 8365 15910 8415
rect 15960 8365 16005 8415
rect 16055 8365 18820 8415
rect 12890 8325 18820 8365
rect 12890 8275 12925 8325
rect 12975 8275 13020 8325
rect 13070 8275 13115 8325
rect 13165 8275 13215 8325
rect 13265 8275 13315 8325
rect 13365 8275 13415 8325
rect 13465 8275 13510 8325
rect 13560 8275 13605 8325
rect 13655 8275 13725 8325
rect 13775 8275 13820 8325
rect 13870 8275 13915 8325
rect 13965 8275 14015 8325
rect 14065 8275 14115 8325
rect 14165 8275 14215 8325
rect 14265 8275 14310 8325
rect 14360 8275 14405 8325
rect 14455 8275 14525 8325
rect 14575 8275 14620 8325
rect 14670 8275 14715 8325
rect 14765 8275 14815 8325
rect 14865 8275 14915 8325
rect 14965 8275 15015 8325
rect 15065 8275 15110 8325
rect 15160 8275 15205 8325
rect 15255 8275 15325 8325
rect 15375 8275 15420 8325
rect 15470 8275 15515 8325
rect 15565 8275 15615 8325
rect 15665 8275 15715 8325
rect 15765 8275 15815 8325
rect 15865 8275 15910 8325
rect 15960 8275 16005 8325
rect 16055 8275 18820 8325
rect 12890 8225 18820 8275
rect 12890 8175 12925 8225
rect 12975 8175 13020 8225
rect 13070 8175 13115 8225
rect 13165 8175 13215 8225
rect 13265 8175 13315 8225
rect 13365 8175 13415 8225
rect 13465 8175 13510 8225
rect 13560 8175 13605 8225
rect 13655 8175 13725 8225
rect 13775 8175 13820 8225
rect 13870 8175 13915 8225
rect 13965 8175 14015 8225
rect 14065 8175 14115 8225
rect 14165 8175 14215 8225
rect 14265 8175 14310 8225
rect 14360 8175 14405 8225
rect 14455 8175 14525 8225
rect 14575 8175 14620 8225
rect 14670 8175 14715 8225
rect 14765 8175 14815 8225
rect 14865 8175 14915 8225
rect 14965 8175 15015 8225
rect 15065 8175 15110 8225
rect 15160 8175 15205 8225
rect 15255 8175 15325 8225
rect 15375 8175 15420 8225
rect 15470 8175 15515 8225
rect 15565 8175 15615 8225
rect 15665 8175 15715 8225
rect 15765 8175 15815 8225
rect 15865 8175 15910 8225
rect 15960 8175 16005 8225
rect 16055 8175 18820 8225
rect 12890 8135 18820 8175
rect 12890 8085 12925 8135
rect 12975 8085 13020 8135
rect 13070 8085 13115 8135
rect 13165 8085 13215 8135
rect 13265 8085 13315 8135
rect 13365 8085 13415 8135
rect 13465 8085 13510 8135
rect 13560 8085 13605 8135
rect 13655 8085 13725 8135
rect 13775 8085 13820 8135
rect 13870 8085 13915 8135
rect 13965 8085 14015 8135
rect 14065 8085 14115 8135
rect 14165 8085 14215 8135
rect 14265 8085 14310 8135
rect 14360 8085 14405 8135
rect 14455 8085 14525 8135
rect 14575 8085 14620 8135
rect 14670 8085 14715 8135
rect 14765 8085 14815 8135
rect 14865 8085 14915 8135
rect 14965 8085 15015 8135
rect 15065 8085 15110 8135
rect 15160 8085 15205 8135
rect 15255 8085 15325 8135
rect 15375 8085 15420 8135
rect 15470 8085 15515 8135
rect 15565 8085 15615 8135
rect 15665 8085 15715 8135
rect 15765 8085 15815 8135
rect 15865 8085 15910 8135
rect 15960 8085 16005 8135
rect 16055 8085 18820 8135
rect 12890 8015 18820 8085
rect 12890 7965 12925 8015
rect 12975 7965 13020 8015
rect 13070 7965 13115 8015
rect 13165 7965 13215 8015
rect 13265 7965 13315 8015
rect 13365 7965 13415 8015
rect 13465 7965 13510 8015
rect 13560 7965 13605 8015
rect 13655 7965 13725 8015
rect 13775 7965 13820 8015
rect 13870 7965 13915 8015
rect 13965 7965 14015 8015
rect 14065 7965 14115 8015
rect 14165 7965 14215 8015
rect 14265 7965 14310 8015
rect 14360 7965 14405 8015
rect 14455 7965 14525 8015
rect 14575 7965 14620 8015
rect 14670 7965 14715 8015
rect 14765 7965 14815 8015
rect 14865 7965 14915 8015
rect 14965 7965 15015 8015
rect 15065 7965 15110 8015
rect 15160 7965 15205 8015
rect 15255 7965 15325 8015
rect 15375 7965 15420 8015
rect 15470 7965 15515 8015
rect 15565 7965 15615 8015
rect 15665 7965 15715 8015
rect 15765 7965 15815 8015
rect 15865 7965 15910 8015
rect 15960 7965 16005 8015
rect 16055 7965 18820 8015
rect 12890 7925 18820 7965
rect 12890 7875 12925 7925
rect 12975 7875 13020 7925
rect 13070 7875 13115 7925
rect 13165 7875 13215 7925
rect 13265 7875 13315 7925
rect 13365 7875 13415 7925
rect 13465 7875 13510 7925
rect 13560 7875 13605 7925
rect 13655 7875 13725 7925
rect 13775 7875 13820 7925
rect 13870 7875 13915 7925
rect 13965 7875 14015 7925
rect 14065 7875 14115 7925
rect 14165 7875 14215 7925
rect 14265 7875 14310 7925
rect 14360 7875 14405 7925
rect 14455 7875 14525 7925
rect 14575 7875 14620 7925
rect 14670 7875 14715 7925
rect 14765 7875 14815 7925
rect 14865 7875 14915 7925
rect 14965 7875 15015 7925
rect 15065 7875 15110 7925
rect 15160 7875 15205 7925
rect 15255 7875 15325 7925
rect 15375 7875 15420 7925
rect 15470 7875 15515 7925
rect 15565 7875 15615 7925
rect 15665 7875 15715 7925
rect 15765 7875 15815 7925
rect 15865 7875 15910 7925
rect 15960 7875 16005 7925
rect 16055 7875 18820 7925
rect 12890 7825 18820 7875
rect 12890 7775 12925 7825
rect 12975 7775 13020 7825
rect 13070 7775 13115 7825
rect 13165 7775 13215 7825
rect 13265 7775 13315 7825
rect 13365 7775 13415 7825
rect 13465 7775 13510 7825
rect 13560 7775 13605 7825
rect 13655 7775 13725 7825
rect 13775 7775 13820 7825
rect 13870 7775 13915 7825
rect 13965 7775 14015 7825
rect 14065 7775 14115 7825
rect 14165 7775 14215 7825
rect 14265 7775 14310 7825
rect 14360 7775 14405 7825
rect 14455 7775 14525 7825
rect 14575 7775 14620 7825
rect 14670 7775 14715 7825
rect 14765 7775 14815 7825
rect 14865 7775 14915 7825
rect 14965 7775 15015 7825
rect 15065 7775 15110 7825
rect 15160 7775 15205 7825
rect 15255 7775 15325 7825
rect 15375 7775 15420 7825
rect 15470 7775 15515 7825
rect 15565 7775 15615 7825
rect 15665 7775 15715 7825
rect 15765 7775 15815 7825
rect 15865 7775 15910 7825
rect 15960 7775 16005 7825
rect 16055 7775 18820 7825
rect 12890 7735 18820 7775
rect 12890 7685 12925 7735
rect 12975 7685 13020 7735
rect 13070 7685 13115 7735
rect 13165 7685 13215 7735
rect 13265 7685 13315 7735
rect 13365 7685 13415 7735
rect 13465 7685 13510 7735
rect 13560 7685 13605 7735
rect 13655 7685 13725 7735
rect 13775 7685 13820 7735
rect 13870 7685 13915 7735
rect 13965 7685 14015 7735
rect 14065 7685 14115 7735
rect 14165 7685 14215 7735
rect 14265 7685 14310 7735
rect 14360 7685 14405 7735
rect 14455 7685 14525 7735
rect 14575 7685 14620 7735
rect 14670 7685 14715 7735
rect 14765 7685 14815 7735
rect 14865 7685 14915 7735
rect 14965 7685 15015 7735
rect 15065 7685 15110 7735
rect 15160 7685 15205 7735
rect 15255 7685 15325 7735
rect 15375 7685 15420 7735
rect 15470 7685 15515 7735
rect 15565 7685 15615 7735
rect 15665 7685 15715 7735
rect 15765 7685 15815 7735
rect 15865 7685 15910 7735
rect 15960 7685 16005 7735
rect 16055 7685 18820 7735
rect 12890 7615 18820 7685
rect 12890 7565 12925 7615
rect 12975 7565 13020 7615
rect 13070 7565 13115 7615
rect 13165 7565 13215 7615
rect 13265 7565 13315 7615
rect 13365 7565 13415 7615
rect 13465 7565 13510 7615
rect 13560 7565 13605 7615
rect 13655 7565 13725 7615
rect 13775 7565 13820 7615
rect 13870 7565 13915 7615
rect 13965 7565 14015 7615
rect 14065 7565 14115 7615
rect 14165 7565 14215 7615
rect 14265 7565 14310 7615
rect 14360 7565 14405 7615
rect 14455 7565 14525 7615
rect 14575 7565 14620 7615
rect 14670 7565 14715 7615
rect 14765 7565 14815 7615
rect 14865 7565 14915 7615
rect 14965 7565 15015 7615
rect 15065 7565 15110 7615
rect 15160 7565 15205 7615
rect 15255 7565 15325 7615
rect 15375 7565 15420 7615
rect 15470 7565 15515 7615
rect 15565 7565 15615 7615
rect 15665 7565 15715 7615
rect 15765 7565 15815 7615
rect 15865 7565 15910 7615
rect 15960 7565 16005 7615
rect 16055 7565 18820 7615
rect 12890 7525 18820 7565
rect 12890 7475 12925 7525
rect 12975 7475 13020 7525
rect 13070 7475 13115 7525
rect 13165 7475 13215 7525
rect 13265 7475 13315 7525
rect 13365 7475 13415 7525
rect 13465 7475 13510 7525
rect 13560 7475 13605 7525
rect 13655 7475 13725 7525
rect 13775 7475 13820 7525
rect 13870 7475 13915 7525
rect 13965 7475 14015 7525
rect 14065 7475 14115 7525
rect 14165 7475 14215 7525
rect 14265 7475 14310 7525
rect 14360 7475 14405 7525
rect 14455 7475 14525 7525
rect 14575 7475 14620 7525
rect 14670 7475 14715 7525
rect 14765 7475 14815 7525
rect 14865 7475 14915 7525
rect 14965 7475 15015 7525
rect 15065 7475 15110 7525
rect 15160 7475 15205 7525
rect 15255 7475 15325 7525
rect 15375 7475 15420 7525
rect 15470 7475 15515 7525
rect 15565 7475 15615 7525
rect 15665 7475 15715 7525
rect 15765 7475 15815 7525
rect 15865 7475 15910 7525
rect 15960 7475 16005 7525
rect 16055 7475 18820 7525
rect 12890 7425 18820 7475
rect 12890 7375 12925 7425
rect 12975 7375 13020 7425
rect 13070 7375 13115 7425
rect 13165 7375 13215 7425
rect 13265 7375 13315 7425
rect 13365 7375 13415 7425
rect 13465 7375 13510 7425
rect 13560 7375 13605 7425
rect 13655 7375 13725 7425
rect 13775 7375 13820 7425
rect 13870 7375 13915 7425
rect 13965 7375 14015 7425
rect 14065 7375 14115 7425
rect 14165 7375 14215 7425
rect 14265 7375 14310 7425
rect 14360 7375 14405 7425
rect 14455 7375 14525 7425
rect 14575 7375 14620 7425
rect 14670 7375 14715 7425
rect 14765 7375 14815 7425
rect 14865 7375 14915 7425
rect 14965 7375 15015 7425
rect 15065 7375 15110 7425
rect 15160 7375 15205 7425
rect 15255 7375 15325 7425
rect 15375 7375 15420 7425
rect 15470 7375 15515 7425
rect 15565 7375 15615 7425
rect 15665 7375 15715 7425
rect 15765 7375 15815 7425
rect 15865 7375 15910 7425
rect 15960 7375 16005 7425
rect 16055 7375 18820 7425
rect 12890 7335 18820 7375
rect 12890 7285 12925 7335
rect 12975 7285 13020 7335
rect 13070 7285 13115 7335
rect 13165 7285 13215 7335
rect 13265 7285 13315 7335
rect 13365 7285 13415 7335
rect 13465 7285 13510 7335
rect 13560 7285 13605 7335
rect 13655 7285 13725 7335
rect 13775 7285 13820 7335
rect 13870 7285 13915 7335
rect 13965 7285 14015 7335
rect 14065 7285 14115 7335
rect 14165 7285 14215 7335
rect 14265 7285 14310 7335
rect 14360 7285 14405 7335
rect 14455 7285 14525 7335
rect 14575 7285 14620 7335
rect 14670 7285 14715 7335
rect 14765 7285 14815 7335
rect 14865 7285 14915 7335
rect 14965 7285 15015 7335
rect 15065 7285 15110 7335
rect 15160 7285 15205 7335
rect 15255 7285 15325 7335
rect 15375 7285 15420 7335
rect 15470 7285 15515 7335
rect 15565 7285 15615 7335
rect 15665 7285 15715 7335
rect 15765 7285 15815 7335
rect 15865 7285 15910 7335
rect 15960 7285 16005 7335
rect 16055 7285 18820 7335
rect 12890 7215 18820 7285
rect 12890 7165 12925 7215
rect 12975 7165 13020 7215
rect 13070 7165 13115 7215
rect 13165 7165 13215 7215
rect 13265 7165 13315 7215
rect 13365 7165 13415 7215
rect 13465 7165 13510 7215
rect 13560 7165 13605 7215
rect 13655 7165 13725 7215
rect 13775 7165 13820 7215
rect 13870 7165 13915 7215
rect 13965 7165 14015 7215
rect 14065 7165 14115 7215
rect 14165 7165 14215 7215
rect 14265 7165 14310 7215
rect 14360 7165 14405 7215
rect 14455 7165 14525 7215
rect 14575 7165 14620 7215
rect 14670 7165 14715 7215
rect 14765 7165 14815 7215
rect 14865 7165 14915 7215
rect 14965 7165 15015 7215
rect 15065 7165 15110 7215
rect 15160 7165 15205 7215
rect 15255 7165 15325 7215
rect 15375 7165 15420 7215
rect 15470 7165 15515 7215
rect 15565 7165 15615 7215
rect 15665 7165 15715 7215
rect 15765 7165 15815 7215
rect 15865 7165 15910 7215
rect 15960 7165 16005 7215
rect 16055 7165 18820 7215
rect 12890 7125 18820 7165
rect 12890 7075 12925 7125
rect 12975 7075 13020 7125
rect 13070 7075 13115 7125
rect 13165 7075 13215 7125
rect 13265 7075 13315 7125
rect 13365 7075 13415 7125
rect 13465 7075 13510 7125
rect 13560 7075 13605 7125
rect 13655 7075 13725 7125
rect 13775 7075 13820 7125
rect 13870 7075 13915 7125
rect 13965 7075 14015 7125
rect 14065 7075 14115 7125
rect 14165 7075 14215 7125
rect 14265 7075 14310 7125
rect 14360 7075 14405 7125
rect 14455 7075 14525 7125
rect 14575 7075 14620 7125
rect 14670 7075 14715 7125
rect 14765 7075 14815 7125
rect 14865 7075 14915 7125
rect 14965 7075 15015 7125
rect 15065 7075 15110 7125
rect 15160 7075 15205 7125
rect 15255 7075 15325 7125
rect 15375 7075 15420 7125
rect 15470 7075 15515 7125
rect 15565 7075 15615 7125
rect 15665 7075 15715 7125
rect 15765 7075 15815 7125
rect 15865 7075 15910 7125
rect 15960 7075 16005 7125
rect 16055 7075 18820 7125
rect 12890 7025 18820 7075
rect 12890 6975 12925 7025
rect 12975 6975 13020 7025
rect 13070 6975 13115 7025
rect 13165 6975 13215 7025
rect 13265 6975 13315 7025
rect 13365 6975 13415 7025
rect 13465 6975 13510 7025
rect 13560 6975 13605 7025
rect 13655 6975 13725 7025
rect 13775 6975 13820 7025
rect 13870 6975 13915 7025
rect 13965 6975 14015 7025
rect 14065 6975 14115 7025
rect 14165 6975 14215 7025
rect 14265 6975 14310 7025
rect 14360 6975 14405 7025
rect 14455 6975 14525 7025
rect 14575 6975 14620 7025
rect 14670 6975 14715 7025
rect 14765 6975 14815 7025
rect 14865 6975 14915 7025
rect 14965 6975 15015 7025
rect 15065 6975 15110 7025
rect 15160 6975 15205 7025
rect 15255 6975 15325 7025
rect 15375 6975 15420 7025
rect 15470 6975 15515 7025
rect 15565 6975 15615 7025
rect 15665 6975 15715 7025
rect 15765 6975 15815 7025
rect 15865 6975 15910 7025
rect 15960 6975 16005 7025
rect 16055 6975 18820 7025
rect 12890 6935 18820 6975
rect 12890 6885 12925 6935
rect 12975 6885 13020 6935
rect 13070 6885 13115 6935
rect 13165 6885 13215 6935
rect 13265 6885 13315 6935
rect 13365 6885 13415 6935
rect 13465 6885 13510 6935
rect 13560 6885 13605 6935
rect 13655 6885 13725 6935
rect 13775 6885 13820 6935
rect 13870 6885 13915 6935
rect 13965 6885 14015 6935
rect 14065 6885 14115 6935
rect 14165 6885 14215 6935
rect 14265 6885 14310 6935
rect 14360 6885 14405 6935
rect 14455 6885 14525 6935
rect 14575 6885 14620 6935
rect 14670 6885 14715 6935
rect 14765 6885 14815 6935
rect 14865 6885 14915 6935
rect 14965 6885 15015 6935
rect 15065 6885 15110 6935
rect 15160 6885 15205 6935
rect 15255 6885 15325 6935
rect 15375 6885 15420 6935
rect 15470 6885 15515 6935
rect 15565 6885 15615 6935
rect 15665 6885 15715 6935
rect 15765 6885 15815 6935
rect 15865 6885 15910 6935
rect 15960 6885 16005 6935
rect 16055 6885 18820 6935
rect 12890 6815 18820 6885
rect 12890 6765 12925 6815
rect 12975 6765 13020 6815
rect 13070 6765 13115 6815
rect 13165 6765 13215 6815
rect 13265 6765 13315 6815
rect 13365 6765 13415 6815
rect 13465 6765 13510 6815
rect 13560 6765 13605 6815
rect 13655 6765 13725 6815
rect 13775 6765 13820 6815
rect 13870 6765 13915 6815
rect 13965 6765 14015 6815
rect 14065 6765 14115 6815
rect 14165 6765 14215 6815
rect 14265 6765 14310 6815
rect 14360 6765 14405 6815
rect 14455 6765 14525 6815
rect 14575 6765 14620 6815
rect 14670 6765 14715 6815
rect 14765 6765 14815 6815
rect 14865 6765 14915 6815
rect 14965 6765 15015 6815
rect 15065 6765 15110 6815
rect 15160 6765 15205 6815
rect 15255 6765 15325 6815
rect 15375 6765 15420 6815
rect 15470 6765 15515 6815
rect 15565 6765 15615 6815
rect 15665 6765 15715 6815
rect 15765 6765 15815 6815
rect 15865 6765 15910 6815
rect 15960 6765 16005 6815
rect 16055 6765 18820 6815
rect 12890 6725 18820 6765
rect 12890 6675 12925 6725
rect 12975 6675 13020 6725
rect 13070 6675 13115 6725
rect 13165 6675 13215 6725
rect 13265 6675 13315 6725
rect 13365 6675 13415 6725
rect 13465 6675 13510 6725
rect 13560 6675 13605 6725
rect 13655 6675 13725 6725
rect 13775 6675 13820 6725
rect 13870 6675 13915 6725
rect 13965 6675 14015 6725
rect 14065 6675 14115 6725
rect 14165 6675 14215 6725
rect 14265 6675 14310 6725
rect 14360 6675 14405 6725
rect 14455 6675 14525 6725
rect 14575 6675 14620 6725
rect 14670 6675 14715 6725
rect 14765 6675 14815 6725
rect 14865 6675 14915 6725
rect 14965 6675 15015 6725
rect 15065 6675 15110 6725
rect 15160 6675 15205 6725
rect 15255 6675 15325 6725
rect 15375 6675 15420 6725
rect 15470 6675 15515 6725
rect 15565 6675 15615 6725
rect 15665 6675 15715 6725
rect 15765 6675 15815 6725
rect 15865 6675 15910 6725
rect 15960 6675 16005 6725
rect 16055 6675 18820 6725
rect 12890 6625 18820 6675
rect 12890 6575 12925 6625
rect 12975 6575 13020 6625
rect 13070 6575 13115 6625
rect 13165 6575 13215 6625
rect 13265 6575 13315 6625
rect 13365 6575 13415 6625
rect 13465 6575 13510 6625
rect 13560 6575 13605 6625
rect 13655 6575 13725 6625
rect 13775 6575 13820 6625
rect 13870 6575 13915 6625
rect 13965 6575 14015 6625
rect 14065 6575 14115 6625
rect 14165 6575 14215 6625
rect 14265 6575 14310 6625
rect 14360 6575 14405 6625
rect 14455 6575 14525 6625
rect 14575 6575 14620 6625
rect 14670 6575 14715 6625
rect 14765 6575 14815 6625
rect 14865 6575 14915 6625
rect 14965 6575 15015 6625
rect 15065 6575 15110 6625
rect 15160 6575 15205 6625
rect 15255 6575 15325 6625
rect 15375 6575 15420 6625
rect 15470 6575 15515 6625
rect 15565 6575 15615 6625
rect 15665 6575 15715 6625
rect 15765 6575 15815 6625
rect 15865 6575 15910 6625
rect 15960 6575 16005 6625
rect 16055 6575 18820 6625
rect 12890 6535 18820 6575
rect 12890 6485 12925 6535
rect 12975 6485 13020 6535
rect 13070 6485 13115 6535
rect 13165 6485 13215 6535
rect 13265 6485 13315 6535
rect 13365 6485 13415 6535
rect 13465 6485 13510 6535
rect 13560 6485 13605 6535
rect 13655 6485 13725 6535
rect 13775 6485 13820 6535
rect 13870 6485 13915 6535
rect 13965 6485 14015 6535
rect 14065 6485 14115 6535
rect 14165 6485 14215 6535
rect 14265 6485 14310 6535
rect 14360 6485 14405 6535
rect 14455 6485 14525 6535
rect 14575 6485 14620 6535
rect 14670 6485 14715 6535
rect 14765 6485 14815 6535
rect 14865 6485 14915 6535
rect 14965 6485 15015 6535
rect 15065 6485 15110 6535
rect 15160 6485 15205 6535
rect 15255 6485 15325 6535
rect 15375 6485 15420 6535
rect 15470 6485 15515 6535
rect 15565 6485 15615 6535
rect 15665 6485 15715 6535
rect 15765 6485 15815 6535
rect 15865 6485 15910 6535
rect 15960 6485 16005 6535
rect 16055 6485 18820 6535
rect 12890 6450 18820 6485
rect -120 -1300 16090 -1290
rect -120 -1340 -80 -1300
rect -40 -1340 270 -1300
rect 310 -1340 620 -1300
rect 660 -1340 970 -1300
rect 1010 -1340 1320 -1300
rect 1360 -1340 1670 -1300
rect 1710 -1340 2020 -1300
rect 2060 -1340 2370 -1300
rect 2410 -1340 2720 -1300
rect 2760 -1340 3070 -1300
rect 3110 -1340 3420 -1300
rect 3460 -1340 3770 -1300
rect 3810 -1340 4120 -1300
rect 4160 -1340 4470 -1300
rect 4510 -1340 4820 -1300
rect 4860 -1340 5170 -1300
rect 5210 -1340 5520 -1300
rect 5560 -1340 5870 -1300
rect 5910 -1340 6220 -1300
rect 6260 -1340 6570 -1300
rect 6610 -1340 6920 -1300
rect 6960 -1340 7270 -1300
rect 7310 -1340 7620 -1300
rect 7660 -1340 7970 -1300
rect 8010 -1340 8320 -1300
rect 8360 -1325 16090 -1300
rect 8360 -1340 12925 -1325
rect -120 -1365 12925 -1340
rect -120 -1405 -80 -1365
rect -40 -1405 270 -1365
rect 310 -1405 620 -1365
rect 660 -1405 970 -1365
rect 1010 -1405 1320 -1365
rect 1360 -1405 1670 -1365
rect 1710 -1405 2020 -1365
rect 2060 -1405 2370 -1365
rect 2410 -1405 2720 -1365
rect 2760 -1405 3070 -1365
rect 3110 -1405 3420 -1365
rect 3460 -1405 3770 -1365
rect 3810 -1405 4120 -1365
rect 4160 -1405 4470 -1365
rect 4510 -1405 4820 -1365
rect 4860 -1405 5170 -1365
rect 5210 -1405 5520 -1365
rect 5560 -1405 5870 -1365
rect 5910 -1405 6220 -1365
rect 6260 -1405 6570 -1365
rect 6610 -1405 6920 -1365
rect 6960 -1405 7270 -1365
rect 7310 -1405 7620 -1365
rect 7660 -1405 7970 -1365
rect 8010 -1405 8320 -1365
rect 8360 -1375 12925 -1365
rect 12975 -1375 13020 -1325
rect 13070 -1375 13115 -1325
rect 13165 -1375 13215 -1325
rect 13265 -1375 13315 -1325
rect 13365 -1375 13415 -1325
rect 13465 -1375 13510 -1325
rect 13560 -1375 13605 -1325
rect 13655 -1375 13725 -1325
rect 13775 -1375 13820 -1325
rect 13870 -1375 13915 -1325
rect 13965 -1375 14015 -1325
rect 14065 -1375 14115 -1325
rect 14165 -1375 14215 -1325
rect 14265 -1375 14310 -1325
rect 14360 -1375 14405 -1325
rect 14455 -1375 14525 -1325
rect 14575 -1375 14620 -1325
rect 14670 -1375 14715 -1325
rect 14765 -1375 14815 -1325
rect 14865 -1375 14915 -1325
rect 14965 -1375 15015 -1325
rect 15065 -1375 15110 -1325
rect 15160 -1375 15205 -1325
rect 15255 -1375 15325 -1325
rect 15375 -1375 15420 -1325
rect 15470 -1375 15515 -1325
rect 15565 -1375 15615 -1325
rect 15665 -1375 15715 -1325
rect 15765 -1375 15815 -1325
rect 15865 -1375 15910 -1325
rect 15960 -1375 16005 -1325
rect 16055 -1375 16090 -1325
rect 8360 -1405 16090 -1375
rect -120 -1415 16090 -1405
rect -120 -1435 12925 -1415
rect -120 -1475 -80 -1435
rect -40 -1475 270 -1435
rect 310 -1475 620 -1435
rect 660 -1475 970 -1435
rect 1010 -1475 1320 -1435
rect 1360 -1475 1670 -1435
rect 1710 -1475 2020 -1435
rect 2060 -1475 2370 -1435
rect 2410 -1475 2720 -1435
rect 2760 -1475 3070 -1435
rect 3110 -1475 3420 -1435
rect 3460 -1475 3770 -1435
rect 3810 -1475 4120 -1435
rect 4160 -1475 4470 -1435
rect 4510 -1475 4820 -1435
rect 4860 -1475 5170 -1435
rect 5210 -1475 5520 -1435
rect 5560 -1475 5870 -1435
rect 5910 -1475 6220 -1435
rect 6260 -1475 6570 -1435
rect 6610 -1475 6920 -1435
rect 6960 -1475 7270 -1435
rect 7310 -1475 7620 -1435
rect 7660 -1475 7970 -1435
rect 8010 -1475 8320 -1435
rect 8360 -1465 12925 -1435
rect 12975 -1465 13020 -1415
rect 13070 -1465 13115 -1415
rect 13165 -1465 13215 -1415
rect 13265 -1465 13315 -1415
rect 13365 -1465 13415 -1415
rect 13465 -1465 13510 -1415
rect 13560 -1465 13605 -1415
rect 13655 -1465 13725 -1415
rect 13775 -1465 13820 -1415
rect 13870 -1465 13915 -1415
rect 13965 -1465 14015 -1415
rect 14065 -1465 14115 -1415
rect 14165 -1465 14215 -1415
rect 14265 -1465 14310 -1415
rect 14360 -1465 14405 -1415
rect 14455 -1465 14525 -1415
rect 14575 -1465 14620 -1415
rect 14670 -1465 14715 -1415
rect 14765 -1465 14815 -1415
rect 14865 -1465 14915 -1415
rect 14965 -1465 15015 -1415
rect 15065 -1465 15110 -1415
rect 15160 -1465 15205 -1415
rect 15255 -1465 15325 -1415
rect 15375 -1465 15420 -1415
rect 15470 -1465 15515 -1415
rect 15565 -1465 15615 -1415
rect 15665 -1465 15715 -1415
rect 15765 -1465 15815 -1415
rect 15865 -1465 15910 -1415
rect 15960 -1465 16005 -1415
rect 16055 -1465 16090 -1415
rect 8360 -1475 16090 -1465
rect -120 -1505 16090 -1475
rect -120 -1545 -80 -1505
rect -40 -1545 270 -1505
rect 310 -1545 620 -1505
rect 660 -1545 970 -1505
rect 1010 -1545 1320 -1505
rect 1360 -1545 1670 -1505
rect 1710 -1545 2020 -1505
rect 2060 -1545 2370 -1505
rect 2410 -1545 2720 -1505
rect 2760 -1545 3070 -1505
rect 3110 -1545 3420 -1505
rect 3460 -1545 3770 -1505
rect 3810 -1545 4120 -1505
rect 4160 -1545 4470 -1505
rect 4510 -1545 4820 -1505
rect 4860 -1545 5170 -1505
rect 5210 -1545 5520 -1505
rect 5560 -1545 5870 -1505
rect 5910 -1545 6220 -1505
rect 6260 -1545 6570 -1505
rect 6610 -1545 6920 -1505
rect 6960 -1545 7270 -1505
rect 7310 -1545 7620 -1505
rect 7660 -1545 7970 -1505
rect 8010 -1545 8320 -1505
rect 8360 -1515 16090 -1505
rect 8360 -1545 12925 -1515
rect -120 -1565 12925 -1545
rect 12975 -1565 13020 -1515
rect 13070 -1565 13115 -1515
rect 13165 -1565 13215 -1515
rect 13265 -1565 13315 -1515
rect 13365 -1565 13415 -1515
rect 13465 -1565 13510 -1515
rect 13560 -1565 13605 -1515
rect 13655 -1565 13725 -1515
rect 13775 -1565 13820 -1515
rect 13870 -1565 13915 -1515
rect 13965 -1565 14015 -1515
rect 14065 -1565 14115 -1515
rect 14165 -1565 14215 -1515
rect 14265 -1565 14310 -1515
rect 14360 -1565 14405 -1515
rect 14455 -1565 14525 -1515
rect 14575 -1565 14620 -1515
rect 14670 -1565 14715 -1515
rect 14765 -1565 14815 -1515
rect 14865 -1565 14915 -1515
rect 14965 -1565 15015 -1515
rect 15065 -1565 15110 -1515
rect 15160 -1565 15205 -1515
rect 15255 -1565 15325 -1515
rect 15375 -1565 15420 -1515
rect 15470 -1565 15515 -1515
rect 15565 -1565 15615 -1515
rect 15665 -1565 15715 -1515
rect 15765 -1565 15815 -1515
rect 15865 -1565 15910 -1515
rect 15960 -1565 16005 -1515
rect 16055 -1565 16090 -1515
rect -120 -1575 16090 -1565
rect -120 -1615 -80 -1575
rect -40 -1615 270 -1575
rect 310 -1615 620 -1575
rect 660 -1615 970 -1575
rect 1010 -1615 1320 -1575
rect 1360 -1615 1670 -1575
rect 1710 -1615 2020 -1575
rect 2060 -1615 2370 -1575
rect 2410 -1615 2720 -1575
rect 2760 -1615 3070 -1575
rect 3110 -1615 3420 -1575
rect 3460 -1615 3770 -1575
rect 3810 -1615 4120 -1575
rect 4160 -1615 4470 -1575
rect 4510 -1615 4820 -1575
rect 4860 -1615 5170 -1575
rect 5210 -1615 5520 -1575
rect 5560 -1615 5870 -1575
rect 5910 -1615 6220 -1575
rect 6260 -1615 6570 -1575
rect 6610 -1615 6920 -1575
rect 6960 -1615 7270 -1575
rect 7310 -1615 7620 -1575
rect 7660 -1615 7970 -1575
rect 8010 -1615 8320 -1575
rect 8360 -1605 16090 -1575
rect 8360 -1615 12925 -1605
rect -120 -1640 12925 -1615
rect -120 -1680 -80 -1640
rect -40 -1680 270 -1640
rect 310 -1680 620 -1640
rect 660 -1680 970 -1640
rect 1010 -1680 1320 -1640
rect 1360 -1680 1670 -1640
rect 1710 -1680 2020 -1640
rect 2060 -1680 2370 -1640
rect 2410 -1680 2720 -1640
rect 2760 -1680 3070 -1640
rect 3110 -1680 3420 -1640
rect 3460 -1680 3770 -1640
rect 3810 -1680 4120 -1640
rect 4160 -1680 4470 -1640
rect 4510 -1680 4820 -1640
rect 4860 -1680 5170 -1640
rect 5210 -1680 5520 -1640
rect 5560 -1680 5870 -1640
rect 5910 -1680 6220 -1640
rect 6260 -1680 6570 -1640
rect 6610 -1680 6920 -1640
rect 6960 -1680 7270 -1640
rect 7310 -1680 7620 -1640
rect 7660 -1680 7970 -1640
rect 8010 -1680 8320 -1640
rect 8360 -1655 12925 -1640
rect 12975 -1655 13020 -1605
rect 13070 -1655 13115 -1605
rect 13165 -1655 13215 -1605
rect 13265 -1655 13315 -1605
rect 13365 -1655 13415 -1605
rect 13465 -1655 13510 -1605
rect 13560 -1655 13605 -1605
rect 13655 -1655 13725 -1605
rect 13775 -1655 13820 -1605
rect 13870 -1655 13915 -1605
rect 13965 -1655 14015 -1605
rect 14065 -1655 14115 -1605
rect 14165 -1655 14215 -1605
rect 14265 -1655 14310 -1605
rect 14360 -1655 14405 -1605
rect 14455 -1655 14525 -1605
rect 14575 -1655 14620 -1605
rect 14670 -1655 14715 -1605
rect 14765 -1655 14815 -1605
rect 14865 -1655 14915 -1605
rect 14965 -1655 15015 -1605
rect 15065 -1655 15110 -1605
rect 15160 -1655 15205 -1605
rect 15255 -1655 15325 -1605
rect 15375 -1655 15420 -1605
rect 15470 -1655 15515 -1605
rect 15565 -1655 15615 -1605
rect 15665 -1655 15715 -1605
rect 15765 -1655 15815 -1605
rect 15865 -1655 15910 -1605
rect 15960 -1655 16005 -1605
rect 16055 -1655 16090 -1605
rect 8360 -1680 16090 -1655
rect -120 -1700 16090 -1680
rect -120 -1740 -80 -1700
rect -40 -1740 270 -1700
rect 310 -1740 620 -1700
rect 660 -1740 970 -1700
rect 1010 -1740 1320 -1700
rect 1360 -1740 1670 -1700
rect 1710 -1740 2020 -1700
rect 2060 -1740 2370 -1700
rect 2410 -1740 2720 -1700
rect 2760 -1740 3070 -1700
rect 3110 -1740 3420 -1700
rect 3460 -1740 3770 -1700
rect 3810 -1740 4120 -1700
rect 4160 -1740 4470 -1700
rect 4510 -1740 4820 -1700
rect 4860 -1740 5170 -1700
rect 5210 -1740 5520 -1700
rect 5560 -1740 5870 -1700
rect 5910 -1740 6220 -1700
rect 6260 -1740 6570 -1700
rect 6610 -1740 6920 -1700
rect 6960 -1740 7270 -1700
rect 7310 -1740 7620 -1700
rect 7660 -1740 7970 -1700
rect 8010 -1740 8320 -1700
rect 8360 -1725 16090 -1700
rect 8360 -1740 12925 -1725
rect -120 -1765 12925 -1740
rect -120 -1805 -80 -1765
rect -40 -1805 270 -1765
rect 310 -1805 620 -1765
rect 660 -1805 970 -1765
rect 1010 -1805 1320 -1765
rect 1360 -1805 1670 -1765
rect 1710 -1805 2020 -1765
rect 2060 -1805 2370 -1765
rect 2410 -1805 2720 -1765
rect 2760 -1805 3070 -1765
rect 3110 -1805 3420 -1765
rect 3460 -1805 3770 -1765
rect 3810 -1805 4120 -1765
rect 4160 -1805 4470 -1765
rect 4510 -1805 4820 -1765
rect 4860 -1805 5170 -1765
rect 5210 -1805 5520 -1765
rect 5560 -1805 5870 -1765
rect 5910 -1805 6220 -1765
rect 6260 -1805 6570 -1765
rect 6610 -1805 6920 -1765
rect 6960 -1805 7270 -1765
rect 7310 -1805 7620 -1765
rect 7660 -1805 7970 -1765
rect 8010 -1805 8320 -1765
rect 8360 -1775 12925 -1765
rect 12975 -1775 13020 -1725
rect 13070 -1775 13115 -1725
rect 13165 -1775 13215 -1725
rect 13265 -1775 13315 -1725
rect 13365 -1775 13415 -1725
rect 13465 -1775 13510 -1725
rect 13560 -1775 13605 -1725
rect 13655 -1775 13725 -1725
rect 13775 -1775 13820 -1725
rect 13870 -1775 13915 -1725
rect 13965 -1775 14015 -1725
rect 14065 -1775 14115 -1725
rect 14165 -1775 14215 -1725
rect 14265 -1775 14310 -1725
rect 14360 -1775 14405 -1725
rect 14455 -1775 14525 -1725
rect 14575 -1775 14620 -1725
rect 14670 -1775 14715 -1725
rect 14765 -1775 14815 -1725
rect 14865 -1775 14915 -1725
rect 14965 -1775 15015 -1725
rect 15065 -1775 15110 -1725
rect 15160 -1775 15205 -1725
rect 15255 -1775 15325 -1725
rect 15375 -1775 15420 -1725
rect 15470 -1775 15515 -1725
rect 15565 -1775 15615 -1725
rect 15665 -1775 15715 -1725
rect 15765 -1775 15815 -1725
rect 15865 -1775 15910 -1725
rect 15960 -1775 16005 -1725
rect 16055 -1775 16090 -1725
rect 8360 -1805 16090 -1775
rect -120 -1815 16090 -1805
rect -120 -1835 12925 -1815
rect -120 -1875 -80 -1835
rect -40 -1875 270 -1835
rect 310 -1875 620 -1835
rect 660 -1875 970 -1835
rect 1010 -1875 1320 -1835
rect 1360 -1875 1670 -1835
rect 1710 -1875 2020 -1835
rect 2060 -1875 2370 -1835
rect 2410 -1875 2720 -1835
rect 2760 -1875 3070 -1835
rect 3110 -1875 3420 -1835
rect 3460 -1875 3770 -1835
rect 3810 -1875 4120 -1835
rect 4160 -1875 4470 -1835
rect 4510 -1875 4820 -1835
rect 4860 -1875 5170 -1835
rect 5210 -1875 5520 -1835
rect 5560 -1875 5870 -1835
rect 5910 -1875 6220 -1835
rect 6260 -1875 6570 -1835
rect 6610 -1875 6920 -1835
rect 6960 -1875 7270 -1835
rect 7310 -1875 7620 -1835
rect 7660 -1875 7970 -1835
rect 8010 -1875 8320 -1835
rect 8360 -1865 12925 -1835
rect 12975 -1865 13020 -1815
rect 13070 -1865 13115 -1815
rect 13165 -1865 13215 -1815
rect 13265 -1865 13315 -1815
rect 13365 -1865 13415 -1815
rect 13465 -1865 13510 -1815
rect 13560 -1865 13605 -1815
rect 13655 -1865 13725 -1815
rect 13775 -1865 13820 -1815
rect 13870 -1865 13915 -1815
rect 13965 -1865 14015 -1815
rect 14065 -1865 14115 -1815
rect 14165 -1865 14215 -1815
rect 14265 -1865 14310 -1815
rect 14360 -1865 14405 -1815
rect 14455 -1865 14525 -1815
rect 14575 -1865 14620 -1815
rect 14670 -1865 14715 -1815
rect 14765 -1865 14815 -1815
rect 14865 -1865 14915 -1815
rect 14965 -1865 15015 -1815
rect 15065 -1865 15110 -1815
rect 15160 -1865 15205 -1815
rect 15255 -1865 15325 -1815
rect 15375 -1865 15420 -1815
rect 15470 -1865 15515 -1815
rect 15565 -1865 15615 -1815
rect 15665 -1865 15715 -1815
rect 15765 -1865 15815 -1815
rect 15865 -1865 15910 -1815
rect 15960 -1865 16005 -1815
rect 16055 -1865 16090 -1815
rect 8360 -1875 16090 -1865
rect -120 -1905 16090 -1875
rect -120 -1945 -80 -1905
rect -40 -1945 270 -1905
rect 310 -1945 620 -1905
rect 660 -1945 970 -1905
rect 1010 -1945 1320 -1905
rect 1360 -1945 1670 -1905
rect 1710 -1945 2020 -1905
rect 2060 -1945 2370 -1905
rect 2410 -1945 2720 -1905
rect 2760 -1945 3070 -1905
rect 3110 -1945 3420 -1905
rect 3460 -1945 3770 -1905
rect 3810 -1945 4120 -1905
rect 4160 -1945 4470 -1905
rect 4510 -1945 4820 -1905
rect 4860 -1945 5170 -1905
rect 5210 -1945 5520 -1905
rect 5560 -1945 5870 -1905
rect 5910 -1945 6220 -1905
rect 6260 -1945 6570 -1905
rect 6610 -1945 6920 -1905
rect 6960 -1945 7270 -1905
rect 7310 -1945 7620 -1905
rect 7660 -1945 7970 -1905
rect 8010 -1945 8320 -1905
rect 8360 -1915 16090 -1905
rect 8360 -1945 12925 -1915
rect -120 -1965 12925 -1945
rect 12975 -1965 13020 -1915
rect 13070 -1965 13115 -1915
rect 13165 -1965 13215 -1915
rect 13265 -1965 13315 -1915
rect 13365 -1965 13415 -1915
rect 13465 -1965 13510 -1915
rect 13560 -1965 13605 -1915
rect 13655 -1965 13725 -1915
rect 13775 -1965 13820 -1915
rect 13870 -1965 13915 -1915
rect 13965 -1965 14015 -1915
rect 14065 -1965 14115 -1915
rect 14165 -1965 14215 -1915
rect 14265 -1965 14310 -1915
rect 14360 -1965 14405 -1915
rect 14455 -1965 14525 -1915
rect 14575 -1965 14620 -1915
rect 14670 -1965 14715 -1915
rect 14765 -1965 14815 -1915
rect 14865 -1965 14915 -1915
rect 14965 -1965 15015 -1915
rect 15065 -1965 15110 -1915
rect 15160 -1965 15205 -1915
rect 15255 -1965 15325 -1915
rect 15375 -1965 15420 -1915
rect 15470 -1965 15515 -1915
rect 15565 -1965 15615 -1915
rect 15665 -1965 15715 -1915
rect 15765 -1965 15815 -1915
rect 15865 -1965 15910 -1915
rect 15960 -1965 16005 -1915
rect 16055 -1965 16090 -1915
rect -120 -1975 16090 -1965
rect -120 -2015 -80 -1975
rect -40 -2015 270 -1975
rect 310 -2015 620 -1975
rect 660 -2015 970 -1975
rect 1010 -2015 1320 -1975
rect 1360 -2015 1670 -1975
rect 1710 -2015 2020 -1975
rect 2060 -2015 2370 -1975
rect 2410 -2015 2720 -1975
rect 2760 -2015 3070 -1975
rect 3110 -2015 3420 -1975
rect 3460 -2015 3770 -1975
rect 3810 -2015 4120 -1975
rect 4160 -2015 4470 -1975
rect 4510 -2015 4820 -1975
rect 4860 -2015 5170 -1975
rect 5210 -2015 5520 -1975
rect 5560 -2015 5870 -1975
rect 5910 -2015 6220 -1975
rect 6260 -2015 6570 -1975
rect 6610 -2015 6920 -1975
rect 6960 -2015 7270 -1975
rect 7310 -2015 7620 -1975
rect 7660 -2015 7970 -1975
rect 8010 -2015 8320 -1975
rect 8360 -2005 16090 -1975
rect 8360 -2015 12925 -2005
rect -120 -2040 12925 -2015
rect -120 -2080 -80 -2040
rect -40 -2080 270 -2040
rect 310 -2080 620 -2040
rect 660 -2080 970 -2040
rect 1010 -2080 1320 -2040
rect 1360 -2080 1670 -2040
rect 1710 -2080 2020 -2040
rect 2060 -2080 2370 -2040
rect 2410 -2080 2720 -2040
rect 2760 -2080 3070 -2040
rect 3110 -2080 3420 -2040
rect 3460 -2080 3770 -2040
rect 3810 -2080 4120 -2040
rect 4160 -2080 4470 -2040
rect 4510 -2080 4820 -2040
rect 4860 -2080 5170 -2040
rect 5210 -2080 5520 -2040
rect 5560 -2080 5870 -2040
rect 5910 -2080 6220 -2040
rect 6260 -2080 6570 -2040
rect 6610 -2080 6920 -2040
rect 6960 -2080 7270 -2040
rect 7310 -2080 7620 -2040
rect 7660 -2080 7970 -2040
rect 8010 -2080 8320 -2040
rect 8360 -2055 12925 -2040
rect 12975 -2055 13020 -2005
rect 13070 -2055 13115 -2005
rect 13165 -2055 13215 -2005
rect 13265 -2055 13315 -2005
rect 13365 -2055 13415 -2005
rect 13465 -2055 13510 -2005
rect 13560 -2055 13605 -2005
rect 13655 -2055 13725 -2005
rect 13775 -2055 13820 -2005
rect 13870 -2055 13915 -2005
rect 13965 -2055 14015 -2005
rect 14065 -2055 14115 -2005
rect 14165 -2055 14215 -2005
rect 14265 -2055 14310 -2005
rect 14360 -2055 14405 -2005
rect 14455 -2055 14525 -2005
rect 14575 -2055 14620 -2005
rect 14670 -2055 14715 -2005
rect 14765 -2055 14815 -2005
rect 14865 -2055 14915 -2005
rect 14965 -2055 15015 -2005
rect 15065 -2055 15110 -2005
rect 15160 -2055 15205 -2005
rect 15255 -2055 15325 -2005
rect 15375 -2055 15420 -2005
rect 15470 -2055 15515 -2005
rect 15565 -2055 15615 -2005
rect 15665 -2055 15715 -2005
rect 15765 -2055 15815 -2005
rect 15865 -2055 15910 -2005
rect 15960 -2055 16005 -2005
rect 16055 -2055 16090 -2005
rect 8360 -2080 16090 -2055
rect -120 -2100 16090 -2080
rect -120 -2140 -80 -2100
rect -40 -2140 270 -2100
rect 310 -2140 620 -2100
rect 660 -2140 970 -2100
rect 1010 -2140 1320 -2100
rect 1360 -2140 1670 -2100
rect 1710 -2140 2020 -2100
rect 2060 -2140 2370 -2100
rect 2410 -2140 2720 -2100
rect 2760 -2140 3070 -2100
rect 3110 -2140 3420 -2100
rect 3460 -2140 3770 -2100
rect 3810 -2140 4120 -2100
rect 4160 -2140 4470 -2100
rect 4510 -2140 4820 -2100
rect 4860 -2140 5170 -2100
rect 5210 -2140 5520 -2100
rect 5560 -2140 5870 -2100
rect 5910 -2140 6220 -2100
rect 6260 -2140 6570 -2100
rect 6610 -2140 6920 -2100
rect 6960 -2140 7270 -2100
rect 7310 -2140 7620 -2100
rect 7660 -2140 7970 -2100
rect 8010 -2140 8320 -2100
rect 8360 -2125 16090 -2100
rect 8360 -2140 12925 -2125
rect -120 -2165 12925 -2140
rect -120 -2205 -80 -2165
rect -40 -2205 270 -2165
rect 310 -2205 620 -2165
rect 660 -2205 970 -2165
rect 1010 -2205 1320 -2165
rect 1360 -2205 1670 -2165
rect 1710 -2205 2020 -2165
rect 2060 -2205 2370 -2165
rect 2410 -2205 2720 -2165
rect 2760 -2205 3070 -2165
rect 3110 -2205 3420 -2165
rect 3460 -2205 3770 -2165
rect 3810 -2205 4120 -2165
rect 4160 -2205 4470 -2165
rect 4510 -2205 4820 -2165
rect 4860 -2205 5170 -2165
rect 5210 -2205 5520 -2165
rect 5560 -2205 5870 -2165
rect 5910 -2205 6220 -2165
rect 6260 -2205 6570 -2165
rect 6610 -2205 6920 -2165
rect 6960 -2205 7270 -2165
rect 7310 -2205 7620 -2165
rect 7660 -2205 7970 -2165
rect 8010 -2205 8320 -2165
rect 8360 -2175 12925 -2165
rect 12975 -2175 13020 -2125
rect 13070 -2175 13115 -2125
rect 13165 -2175 13215 -2125
rect 13265 -2175 13315 -2125
rect 13365 -2175 13415 -2125
rect 13465 -2175 13510 -2125
rect 13560 -2175 13605 -2125
rect 13655 -2175 13725 -2125
rect 13775 -2175 13820 -2125
rect 13870 -2175 13915 -2125
rect 13965 -2175 14015 -2125
rect 14065 -2175 14115 -2125
rect 14165 -2175 14215 -2125
rect 14265 -2175 14310 -2125
rect 14360 -2175 14405 -2125
rect 14455 -2175 14525 -2125
rect 14575 -2175 14620 -2125
rect 14670 -2175 14715 -2125
rect 14765 -2175 14815 -2125
rect 14865 -2175 14915 -2125
rect 14965 -2175 15015 -2125
rect 15065 -2175 15110 -2125
rect 15160 -2175 15205 -2125
rect 15255 -2175 15325 -2125
rect 15375 -2175 15420 -2125
rect 15470 -2175 15515 -2125
rect 15565 -2175 15615 -2125
rect 15665 -2175 15715 -2125
rect 15765 -2175 15815 -2125
rect 15865 -2175 15910 -2125
rect 15960 -2175 16005 -2125
rect 16055 -2175 16090 -2125
rect 8360 -2205 16090 -2175
rect -120 -2215 16090 -2205
rect -120 -2235 12925 -2215
rect -120 -2275 -80 -2235
rect -40 -2275 270 -2235
rect 310 -2275 620 -2235
rect 660 -2275 970 -2235
rect 1010 -2275 1320 -2235
rect 1360 -2275 1670 -2235
rect 1710 -2275 2020 -2235
rect 2060 -2275 2370 -2235
rect 2410 -2275 2720 -2235
rect 2760 -2275 3070 -2235
rect 3110 -2275 3420 -2235
rect 3460 -2275 3770 -2235
rect 3810 -2275 4120 -2235
rect 4160 -2275 4470 -2235
rect 4510 -2275 4820 -2235
rect 4860 -2275 5170 -2235
rect 5210 -2275 5520 -2235
rect 5560 -2275 5870 -2235
rect 5910 -2275 6220 -2235
rect 6260 -2275 6570 -2235
rect 6610 -2275 6920 -2235
rect 6960 -2275 7270 -2235
rect 7310 -2275 7620 -2235
rect 7660 -2275 7970 -2235
rect 8010 -2275 8320 -2235
rect 8360 -2265 12925 -2235
rect 12975 -2265 13020 -2215
rect 13070 -2265 13115 -2215
rect 13165 -2265 13215 -2215
rect 13265 -2265 13315 -2215
rect 13365 -2265 13415 -2215
rect 13465 -2265 13510 -2215
rect 13560 -2265 13605 -2215
rect 13655 -2265 13725 -2215
rect 13775 -2265 13820 -2215
rect 13870 -2265 13915 -2215
rect 13965 -2265 14015 -2215
rect 14065 -2265 14115 -2215
rect 14165 -2265 14215 -2215
rect 14265 -2265 14310 -2215
rect 14360 -2265 14405 -2215
rect 14455 -2265 14525 -2215
rect 14575 -2265 14620 -2215
rect 14670 -2265 14715 -2215
rect 14765 -2265 14815 -2215
rect 14865 -2265 14915 -2215
rect 14965 -2265 15015 -2215
rect 15065 -2265 15110 -2215
rect 15160 -2265 15205 -2215
rect 15255 -2265 15325 -2215
rect 15375 -2265 15420 -2215
rect 15470 -2265 15515 -2215
rect 15565 -2265 15615 -2215
rect 15665 -2265 15715 -2215
rect 15765 -2265 15815 -2215
rect 15865 -2265 15910 -2215
rect 15960 -2265 16005 -2215
rect 16055 -2265 16090 -2215
rect 8360 -2275 16090 -2265
rect -120 -2305 16090 -2275
rect -120 -2345 -80 -2305
rect -40 -2345 270 -2305
rect 310 -2345 620 -2305
rect 660 -2345 970 -2305
rect 1010 -2345 1320 -2305
rect 1360 -2345 1670 -2305
rect 1710 -2345 2020 -2305
rect 2060 -2345 2370 -2305
rect 2410 -2345 2720 -2305
rect 2760 -2345 3070 -2305
rect 3110 -2345 3420 -2305
rect 3460 -2345 3770 -2305
rect 3810 -2345 4120 -2305
rect 4160 -2345 4470 -2305
rect 4510 -2345 4820 -2305
rect 4860 -2345 5170 -2305
rect 5210 -2345 5520 -2305
rect 5560 -2345 5870 -2305
rect 5910 -2345 6220 -2305
rect 6260 -2345 6570 -2305
rect 6610 -2345 6920 -2305
rect 6960 -2345 7270 -2305
rect 7310 -2345 7620 -2305
rect 7660 -2345 7970 -2305
rect 8010 -2345 8320 -2305
rect 8360 -2315 16090 -2305
rect 8360 -2345 12925 -2315
rect -120 -2365 12925 -2345
rect 12975 -2365 13020 -2315
rect 13070 -2365 13115 -2315
rect 13165 -2365 13215 -2315
rect 13265 -2365 13315 -2315
rect 13365 -2365 13415 -2315
rect 13465 -2365 13510 -2315
rect 13560 -2365 13605 -2315
rect 13655 -2365 13725 -2315
rect 13775 -2365 13820 -2315
rect 13870 -2365 13915 -2315
rect 13965 -2365 14015 -2315
rect 14065 -2365 14115 -2315
rect 14165 -2365 14215 -2315
rect 14265 -2365 14310 -2315
rect 14360 -2365 14405 -2315
rect 14455 -2365 14525 -2315
rect 14575 -2365 14620 -2315
rect 14670 -2365 14715 -2315
rect 14765 -2365 14815 -2315
rect 14865 -2365 14915 -2315
rect 14965 -2365 15015 -2315
rect 15065 -2365 15110 -2315
rect 15160 -2365 15205 -2315
rect 15255 -2365 15325 -2315
rect 15375 -2365 15420 -2315
rect 15470 -2365 15515 -2315
rect 15565 -2365 15615 -2315
rect 15665 -2365 15715 -2315
rect 15765 -2365 15815 -2315
rect 15865 -2365 15910 -2315
rect 15960 -2365 16005 -2315
rect 16055 -2365 16090 -2315
rect -120 -2375 16090 -2365
rect -120 -2415 -80 -2375
rect -40 -2415 270 -2375
rect 310 -2415 620 -2375
rect 660 -2415 970 -2375
rect 1010 -2415 1320 -2375
rect 1360 -2415 1670 -2375
rect 1710 -2415 2020 -2375
rect 2060 -2415 2370 -2375
rect 2410 -2415 2720 -2375
rect 2760 -2415 3070 -2375
rect 3110 -2415 3420 -2375
rect 3460 -2415 3770 -2375
rect 3810 -2415 4120 -2375
rect 4160 -2415 4470 -2375
rect 4510 -2415 4820 -2375
rect 4860 -2415 5170 -2375
rect 5210 -2415 5520 -2375
rect 5560 -2415 5870 -2375
rect 5910 -2415 6220 -2375
rect 6260 -2415 6570 -2375
rect 6610 -2415 6920 -2375
rect 6960 -2415 7270 -2375
rect 7310 -2415 7620 -2375
rect 7660 -2415 7970 -2375
rect 8010 -2415 8320 -2375
rect 8360 -2405 16090 -2375
rect 8360 -2415 12925 -2405
rect -120 -2440 12925 -2415
rect -120 -2480 -80 -2440
rect -40 -2480 270 -2440
rect 310 -2480 620 -2440
rect 660 -2480 970 -2440
rect 1010 -2480 1320 -2440
rect 1360 -2480 1670 -2440
rect 1710 -2480 2020 -2440
rect 2060 -2480 2370 -2440
rect 2410 -2480 2720 -2440
rect 2760 -2480 3070 -2440
rect 3110 -2480 3420 -2440
rect 3460 -2480 3770 -2440
rect 3810 -2480 4120 -2440
rect 4160 -2480 4470 -2440
rect 4510 -2480 4820 -2440
rect 4860 -2480 5170 -2440
rect 5210 -2480 5520 -2440
rect 5560 -2480 5870 -2440
rect 5910 -2480 6220 -2440
rect 6260 -2480 6570 -2440
rect 6610 -2480 6920 -2440
rect 6960 -2480 7270 -2440
rect 7310 -2480 7620 -2440
rect 7660 -2480 7970 -2440
rect 8010 -2480 8320 -2440
rect 8360 -2455 12925 -2440
rect 12975 -2455 13020 -2405
rect 13070 -2455 13115 -2405
rect 13165 -2455 13215 -2405
rect 13265 -2455 13315 -2405
rect 13365 -2455 13415 -2405
rect 13465 -2455 13510 -2405
rect 13560 -2455 13605 -2405
rect 13655 -2455 13725 -2405
rect 13775 -2455 13820 -2405
rect 13870 -2455 13915 -2405
rect 13965 -2455 14015 -2405
rect 14065 -2455 14115 -2405
rect 14165 -2455 14215 -2405
rect 14265 -2455 14310 -2405
rect 14360 -2455 14405 -2405
rect 14455 -2455 14525 -2405
rect 14575 -2455 14620 -2405
rect 14670 -2455 14715 -2405
rect 14765 -2455 14815 -2405
rect 14865 -2455 14915 -2405
rect 14965 -2455 15015 -2405
rect 15065 -2455 15110 -2405
rect 15160 -2455 15205 -2405
rect 15255 -2455 15325 -2405
rect 15375 -2455 15420 -2405
rect 15470 -2455 15515 -2405
rect 15565 -2455 15615 -2405
rect 15665 -2455 15715 -2405
rect 15765 -2455 15815 -2405
rect 15865 -2455 15910 -2405
rect 15960 -2455 16005 -2405
rect 16055 -2455 16090 -2405
rect 8360 -2480 16090 -2455
rect -120 -2500 16090 -2480
rect -120 -2540 -80 -2500
rect -40 -2540 270 -2500
rect 310 -2540 620 -2500
rect 660 -2540 970 -2500
rect 1010 -2540 1320 -2500
rect 1360 -2540 1670 -2500
rect 1710 -2540 2020 -2500
rect 2060 -2540 2370 -2500
rect 2410 -2540 2720 -2500
rect 2760 -2540 3070 -2500
rect 3110 -2540 3420 -2500
rect 3460 -2540 3770 -2500
rect 3810 -2540 4120 -2500
rect 4160 -2540 4470 -2500
rect 4510 -2540 4820 -2500
rect 4860 -2540 5170 -2500
rect 5210 -2540 5520 -2500
rect 5560 -2540 5870 -2500
rect 5910 -2540 6220 -2500
rect 6260 -2540 6570 -2500
rect 6610 -2540 6920 -2500
rect 6960 -2540 7270 -2500
rect 7310 -2540 7620 -2500
rect 7660 -2540 7970 -2500
rect 8010 -2540 8320 -2500
rect 8360 -2525 16090 -2500
rect 8360 -2540 12925 -2525
rect -120 -2565 12925 -2540
rect -120 -2605 -80 -2565
rect -40 -2605 270 -2565
rect 310 -2605 620 -2565
rect 660 -2605 970 -2565
rect 1010 -2605 1320 -2565
rect 1360 -2605 1670 -2565
rect 1710 -2605 2020 -2565
rect 2060 -2605 2370 -2565
rect 2410 -2605 2720 -2565
rect 2760 -2605 3070 -2565
rect 3110 -2605 3420 -2565
rect 3460 -2605 3770 -2565
rect 3810 -2605 4120 -2565
rect 4160 -2605 4470 -2565
rect 4510 -2605 4820 -2565
rect 4860 -2605 5170 -2565
rect 5210 -2605 5520 -2565
rect 5560 -2605 5870 -2565
rect 5910 -2605 6220 -2565
rect 6260 -2605 6570 -2565
rect 6610 -2605 6920 -2565
rect 6960 -2605 7270 -2565
rect 7310 -2605 7620 -2565
rect 7660 -2605 7970 -2565
rect 8010 -2605 8320 -2565
rect 8360 -2575 12925 -2565
rect 12975 -2575 13020 -2525
rect 13070 -2575 13115 -2525
rect 13165 -2575 13215 -2525
rect 13265 -2575 13315 -2525
rect 13365 -2575 13415 -2525
rect 13465 -2575 13510 -2525
rect 13560 -2575 13605 -2525
rect 13655 -2575 13725 -2525
rect 13775 -2575 13820 -2525
rect 13870 -2575 13915 -2525
rect 13965 -2575 14015 -2525
rect 14065 -2575 14115 -2525
rect 14165 -2575 14215 -2525
rect 14265 -2575 14310 -2525
rect 14360 -2575 14405 -2525
rect 14455 -2575 14525 -2525
rect 14575 -2575 14620 -2525
rect 14670 -2575 14715 -2525
rect 14765 -2575 14815 -2525
rect 14865 -2575 14915 -2525
rect 14965 -2575 15015 -2525
rect 15065 -2575 15110 -2525
rect 15160 -2575 15205 -2525
rect 15255 -2575 15325 -2525
rect 15375 -2575 15420 -2525
rect 15470 -2575 15515 -2525
rect 15565 -2575 15615 -2525
rect 15665 -2575 15715 -2525
rect 15765 -2575 15815 -2525
rect 15865 -2575 15910 -2525
rect 15960 -2575 16005 -2525
rect 16055 -2575 16090 -2525
rect 8360 -2605 16090 -2575
rect -120 -2615 16090 -2605
rect -120 -2635 12925 -2615
rect -120 -2675 -80 -2635
rect -40 -2675 270 -2635
rect 310 -2675 620 -2635
rect 660 -2675 970 -2635
rect 1010 -2675 1320 -2635
rect 1360 -2675 1670 -2635
rect 1710 -2675 2020 -2635
rect 2060 -2675 2370 -2635
rect 2410 -2675 2720 -2635
rect 2760 -2675 3070 -2635
rect 3110 -2675 3420 -2635
rect 3460 -2675 3770 -2635
rect 3810 -2675 4120 -2635
rect 4160 -2675 4470 -2635
rect 4510 -2675 4820 -2635
rect 4860 -2675 5170 -2635
rect 5210 -2675 5520 -2635
rect 5560 -2675 5870 -2635
rect 5910 -2675 6220 -2635
rect 6260 -2675 6570 -2635
rect 6610 -2675 6920 -2635
rect 6960 -2675 7270 -2635
rect 7310 -2675 7620 -2635
rect 7660 -2675 7970 -2635
rect 8010 -2675 8320 -2635
rect 8360 -2665 12925 -2635
rect 12975 -2665 13020 -2615
rect 13070 -2665 13115 -2615
rect 13165 -2665 13215 -2615
rect 13265 -2665 13315 -2615
rect 13365 -2665 13415 -2615
rect 13465 -2665 13510 -2615
rect 13560 -2665 13605 -2615
rect 13655 -2665 13725 -2615
rect 13775 -2665 13820 -2615
rect 13870 -2665 13915 -2615
rect 13965 -2665 14015 -2615
rect 14065 -2665 14115 -2615
rect 14165 -2665 14215 -2615
rect 14265 -2665 14310 -2615
rect 14360 -2665 14405 -2615
rect 14455 -2665 14525 -2615
rect 14575 -2665 14620 -2615
rect 14670 -2665 14715 -2615
rect 14765 -2665 14815 -2615
rect 14865 -2665 14915 -2615
rect 14965 -2665 15015 -2615
rect 15065 -2665 15110 -2615
rect 15160 -2665 15205 -2615
rect 15255 -2665 15325 -2615
rect 15375 -2665 15420 -2615
rect 15470 -2665 15515 -2615
rect 15565 -2665 15615 -2615
rect 15665 -2665 15715 -2615
rect 15765 -2665 15815 -2615
rect 15865 -2665 15910 -2615
rect 15960 -2665 16005 -2615
rect 16055 -2665 16090 -2615
rect 8360 -2675 16090 -2665
rect -120 -2705 16090 -2675
rect -120 -2745 -80 -2705
rect -40 -2745 270 -2705
rect 310 -2745 620 -2705
rect 660 -2745 970 -2705
rect 1010 -2745 1320 -2705
rect 1360 -2745 1670 -2705
rect 1710 -2745 2020 -2705
rect 2060 -2745 2370 -2705
rect 2410 -2745 2720 -2705
rect 2760 -2745 3070 -2705
rect 3110 -2745 3420 -2705
rect 3460 -2745 3770 -2705
rect 3810 -2745 4120 -2705
rect 4160 -2745 4470 -2705
rect 4510 -2745 4820 -2705
rect 4860 -2745 5170 -2705
rect 5210 -2745 5520 -2705
rect 5560 -2745 5870 -2705
rect 5910 -2745 6220 -2705
rect 6260 -2745 6570 -2705
rect 6610 -2745 6920 -2705
rect 6960 -2745 7270 -2705
rect 7310 -2745 7620 -2705
rect 7660 -2745 7970 -2705
rect 8010 -2745 8320 -2705
rect 8360 -2715 16090 -2705
rect 8360 -2745 12925 -2715
rect -120 -2765 12925 -2745
rect 12975 -2765 13020 -2715
rect 13070 -2765 13115 -2715
rect 13165 -2765 13215 -2715
rect 13265 -2765 13315 -2715
rect 13365 -2765 13415 -2715
rect 13465 -2765 13510 -2715
rect 13560 -2765 13605 -2715
rect 13655 -2765 13725 -2715
rect 13775 -2765 13820 -2715
rect 13870 -2765 13915 -2715
rect 13965 -2765 14015 -2715
rect 14065 -2765 14115 -2715
rect 14165 -2765 14215 -2715
rect 14265 -2765 14310 -2715
rect 14360 -2765 14405 -2715
rect 14455 -2765 14525 -2715
rect 14575 -2765 14620 -2715
rect 14670 -2765 14715 -2715
rect 14765 -2765 14815 -2715
rect 14865 -2765 14915 -2715
rect 14965 -2765 15015 -2715
rect 15065 -2765 15110 -2715
rect 15160 -2765 15205 -2715
rect 15255 -2765 15325 -2715
rect 15375 -2765 15420 -2715
rect 15470 -2765 15515 -2715
rect 15565 -2765 15615 -2715
rect 15665 -2765 15715 -2715
rect 15765 -2765 15815 -2715
rect 15865 -2765 15910 -2715
rect 15960 -2765 16005 -2715
rect 16055 -2765 16090 -2715
rect -120 -2775 16090 -2765
rect -120 -2815 -80 -2775
rect -40 -2815 270 -2775
rect 310 -2815 620 -2775
rect 660 -2815 970 -2775
rect 1010 -2815 1320 -2775
rect 1360 -2815 1670 -2775
rect 1710 -2815 2020 -2775
rect 2060 -2815 2370 -2775
rect 2410 -2815 2720 -2775
rect 2760 -2815 3070 -2775
rect 3110 -2815 3420 -2775
rect 3460 -2815 3770 -2775
rect 3810 -2815 4120 -2775
rect 4160 -2815 4470 -2775
rect 4510 -2815 4820 -2775
rect 4860 -2815 5170 -2775
rect 5210 -2815 5520 -2775
rect 5560 -2815 5870 -2775
rect 5910 -2815 6220 -2775
rect 6260 -2815 6570 -2775
rect 6610 -2815 6920 -2775
rect 6960 -2815 7270 -2775
rect 7310 -2815 7620 -2775
rect 7660 -2815 7970 -2775
rect 8010 -2815 8320 -2775
rect 8360 -2805 16090 -2775
rect 8360 -2815 12925 -2805
rect -120 -2840 12925 -2815
rect -120 -2880 -80 -2840
rect -40 -2880 270 -2840
rect 310 -2880 620 -2840
rect 660 -2880 970 -2840
rect 1010 -2880 1320 -2840
rect 1360 -2880 1670 -2840
rect 1710 -2880 2020 -2840
rect 2060 -2880 2370 -2840
rect 2410 -2880 2720 -2840
rect 2760 -2880 3070 -2840
rect 3110 -2880 3420 -2840
rect 3460 -2880 3770 -2840
rect 3810 -2880 4120 -2840
rect 4160 -2880 4470 -2840
rect 4510 -2880 4820 -2840
rect 4860 -2880 5170 -2840
rect 5210 -2880 5520 -2840
rect 5560 -2880 5870 -2840
rect 5910 -2880 6220 -2840
rect 6260 -2880 6570 -2840
rect 6610 -2880 6920 -2840
rect 6960 -2880 7270 -2840
rect 7310 -2880 7620 -2840
rect 7660 -2880 7970 -2840
rect 8010 -2880 8320 -2840
rect 8360 -2855 12925 -2840
rect 12975 -2855 13020 -2805
rect 13070 -2855 13115 -2805
rect 13165 -2855 13215 -2805
rect 13265 -2855 13315 -2805
rect 13365 -2855 13415 -2805
rect 13465 -2855 13510 -2805
rect 13560 -2855 13605 -2805
rect 13655 -2855 13725 -2805
rect 13775 -2855 13820 -2805
rect 13870 -2855 13915 -2805
rect 13965 -2855 14015 -2805
rect 14065 -2855 14115 -2805
rect 14165 -2855 14215 -2805
rect 14265 -2855 14310 -2805
rect 14360 -2855 14405 -2805
rect 14455 -2855 14525 -2805
rect 14575 -2855 14620 -2805
rect 14670 -2855 14715 -2805
rect 14765 -2855 14815 -2805
rect 14865 -2855 14915 -2805
rect 14965 -2855 15015 -2805
rect 15065 -2855 15110 -2805
rect 15160 -2855 15205 -2805
rect 15255 -2855 15325 -2805
rect 15375 -2855 15420 -2805
rect 15470 -2855 15515 -2805
rect 15565 -2855 15615 -2805
rect 15665 -2855 15715 -2805
rect 15765 -2855 15815 -2805
rect 15865 -2855 15910 -2805
rect 15960 -2855 16005 -2805
rect 16055 -2855 16090 -2805
rect 8360 -2880 16090 -2855
rect -120 -2900 16090 -2880
rect -120 -2940 -80 -2900
rect -40 -2940 270 -2900
rect 310 -2940 620 -2900
rect 660 -2940 970 -2900
rect 1010 -2940 1320 -2900
rect 1360 -2940 1670 -2900
rect 1710 -2940 2020 -2900
rect 2060 -2940 2370 -2900
rect 2410 -2940 2720 -2900
rect 2760 -2940 3070 -2900
rect 3110 -2940 3420 -2900
rect 3460 -2940 3770 -2900
rect 3810 -2940 4120 -2900
rect 4160 -2940 4470 -2900
rect 4510 -2940 4820 -2900
rect 4860 -2940 5170 -2900
rect 5210 -2940 5520 -2900
rect 5560 -2940 5870 -2900
rect 5910 -2940 6220 -2900
rect 6260 -2940 6570 -2900
rect 6610 -2940 6920 -2900
rect 6960 -2940 7270 -2900
rect 7310 -2940 7620 -2900
rect 7660 -2940 7970 -2900
rect 8010 -2940 8320 -2900
rect 8360 -2925 16090 -2900
rect 8360 -2940 12925 -2925
rect -120 -2965 12925 -2940
rect -120 -3005 -80 -2965
rect -40 -3005 270 -2965
rect 310 -3005 620 -2965
rect 660 -3005 970 -2965
rect 1010 -3005 1320 -2965
rect 1360 -3005 1670 -2965
rect 1710 -3005 2020 -2965
rect 2060 -3005 2370 -2965
rect 2410 -3005 2720 -2965
rect 2760 -3005 3070 -2965
rect 3110 -3005 3420 -2965
rect 3460 -3005 3770 -2965
rect 3810 -3005 4120 -2965
rect 4160 -3005 4470 -2965
rect 4510 -3005 4820 -2965
rect 4860 -3005 5170 -2965
rect 5210 -3005 5520 -2965
rect 5560 -3005 5870 -2965
rect 5910 -3005 6220 -2965
rect 6260 -3005 6570 -2965
rect 6610 -3005 6920 -2965
rect 6960 -3005 7270 -2965
rect 7310 -3005 7620 -2965
rect 7660 -3005 7970 -2965
rect 8010 -3005 8320 -2965
rect 8360 -2975 12925 -2965
rect 12975 -2975 13020 -2925
rect 13070 -2975 13115 -2925
rect 13165 -2975 13215 -2925
rect 13265 -2975 13315 -2925
rect 13365 -2975 13415 -2925
rect 13465 -2975 13510 -2925
rect 13560 -2975 13605 -2925
rect 13655 -2975 13725 -2925
rect 13775 -2975 13820 -2925
rect 13870 -2975 13915 -2925
rect 13965 -2975 14015 -2925
rect 14065 -2975 14115 -2925
rect 14165 -2975 14215 -2925
rect 14265 -2975 14310 -2925
rect 14360 -2975 14405 -2925
rect 14455 -2975 14525 -2925
rect 14575 -2975 14620 -2925
rect 14670 -2975 14715 -2925
rect 14765 -2975 14815 -2925
rect 14865 -2975 14915 -2925
rect 14965 -2975 15015 -2925
rect 15065 -2975 15110 -2925
rect 15160 -2975 15205 -2925
rect 15255 -2975 15325 -2925
rect 15375 -2975 15420 -2925
rect 15470 -2975 15515 -2925
rect 15565 -2975 15615 -2925
rect 15665 -2975 15715 -2925
rect 15765 -2975 15815 -2925
rect 15865 -2975 15910 -2925
rect 15960 -2975 16005 -2925
rect 16055 -2975 16090 -2925
rect 8360 -3005 16090 -2975
rect -120 -3015 16090 -3005
rect -120 -3035 12925 -3015
rect -120 -3075 -80 -3035
rect -40 -3075 270 -3035
rect 310 -3075 620 -3035
rect 660 -3075 970 -3035
rect 1010 -3075 1320 -3035
rect 1360 -3075 1670 -3035
rect 1710 -3075 2020 -3035
rect 2060 -3075 2370 -3035
rect 2410 -3075 2720 -3035
rect 2760 -3075 3070 -3035
rect 3110 -3075 3420 -3035
rect 3460 -3075 3770 -3035
rect 3810 -3075 4120 -3035
rect 4160 -3075 4470 -3035
rect 4510 -3075 4820 -3035
rect 4860 -3075 5170 -3035
rect 5210 -3075 5520 -3035
rect 5560 -3075 5870 -3035
rect 5910 -3075 6220 -3035
rect 6260 -3075 6570 -3035
rect 6610 -3075 6920 -3035
rect 6960 -3075 7270 -3035
rect 7310 -3075 7620 -3035
rect 7660 -3075 7970 -3035
rect 8010 -3075 8320 -3035
rect 8360 -3065 12925 -3035
rect 12975 -3065 13020 -3015
rect 13070 -3065 13115 -3015
rect 13165 -3065 13215 -3015
rect 13265 -3065 13315 -3015
rect 13365 -3065 13415 -3015
rect 13465 -3065 13510 -3015
rect 13560 -3065 13605 -3015
rect 13655 -3065 13725 -3015
rect 13775 -3065 13820 -3015
rect 13870 -3065 13915 -3015
rect 13965 -3065 14015 -3015
rect 14065 -3065 14115 -3015
rect 14165 -3065 14215 -3015
rect 14265 -3065 14310 -3015
rect 14360 -3065 14405 -3015
rect 14455 -3065 14525 -3015
rect 14575 -3065 14620 -3015
rect 14670 -3065 14715 -3015
rect 14765 -3065 14815 -3015
rect 14865 -3065 14915 -3015
rect 14965 -3065 15015 -3015
rect 15065 -3065 15110 -3015
rect 15160 -3065 15205 -3015
rect 15255 -3065 15325 -3015
rect 15375 -3065 15420 -3015
rect 15470 -3065 15515 -3015
rect 15565 -3065 15615 -3015
rect 15665 -3065 15715 -3015
rect 15765 -3065 15815 -3015
rect 15865 -3065 15910 -3015
rect 15960 -3065 16005 -3015
rect 16055 -3065 16090 -3015
rect 8360 -3075 16090 -3065
rect -120 -3105 16090 -3075
rect -120 -3145 -80 -3105
rect -40 -3145 270 -3105
rect 310 -3145 620 -3105
rect 660 -3145 970 -3105
rect 1010 -3145 1320 -3105
rect 1360 -3145 1670 -3105
rect 1710 -3145 2020 -3105
rect 2060 -3145 2370 -3105
rect 2410 -3145 2720 -3105
rect 2760 -3145 3070 -3105
rect 3110 -3145 3420 -3105
rect 3460 -3145 3770 -3105
rect 3810 -3145 4120 -3105
rect 4160 -3145 4470 -3105
rect 4510 -3145 4820 -3105
rect 4860 -3145 5170 -3105
rect 5210 -3145 5520 -3105
rect 5560 -3145 5870 -3105
rect 5910 -3145 6220 -3105
rect 6260 -3145 6570 -3105
rect 6610 -3145 6920 -3105
rect 6960 -3145 7270 -3105
rect 7310 -3145 7620 -3105
rect 7660 -3145 7970 -3105
rect 8010 -3145 8320 -3105
rect 8360 -3115 16090 -3105
rect 8360 -3145 12925 -3115
rect -120 -3165 12925 -3145
rect 12975 -3165 13020 -3115
rect 13070 -3165 13115 -3115
rect 13165 -3165 13215 -3115
rect 13265 -3165 13315 -3115
rect 13365 -3165 13415 -3115
rect 13465 -3165 13510 -3115
rect 13560 -3165 13605 -3115
rect 13655 -3165 13725 -3115
rect 13775 -3165 13820 -3115
rect 13870 -3165 13915 -3115
rect 13965 -3165 14015 -3115
rect 14065 -3165 14115 -3115
rect 14165 -3165 14215 -3115
rect 14265 -3165 14310 -3115
rect 14360 -3165 14405 -3115
rect 14455 -3165 14525 -3115
rect 14575 -3165 14620 -3115
rect 14670 -3165 14715 -3115
rect 14765 -3165 14815 -3115
rect 14865 -3165 14915 -3115
rect 14965 -3165 15015 -3115
rect 15065 -3165 15110 -3115
rect 15160 -3165 15205 -3115
rect 15255 -3165 15325 -3115
rect 15375 -3165 15420 -3115
rect 15470 -3165 15515 -3115
rect 15565 -3165 15615 -3115
rect 15665 -3165 15715 -3115
rect 15765 -3165 15815 -3115
rect 15865 -3165 15910 -3115
rect 15960 -3165 16005 -3115
rect 16055 -3165 16090 -3115
rect -120 -3175 16090 -3165
rect -120 -3215 -80 -3175
rect -40 -3215 270 -3175
rect 310 -3215 620 -3175
rect 660 -3215 970 -3175
rect 1010 -3215 1320 -3175
rect 1360 -3215 1670 -3175
rect 1710 -3215 2020 -3175
rect 2060 -3215 2370 -3175
rect 2410 -3215 2720 -3175
rect 2760 -3215 3070 -3175
rect 3110 -3215 3420 -3175
rect 3460 -3215 3770 -3175
rect 3810 -3215 4120 -3175
rect 4160 -3215 4470 -3175
rect 4510 -3215 4820 -3175
rect 4860 -3215 5170 -3175
rect 5210 -3215 5520 -3175
rect 5560 -3215 5870 -3175
rect 5910 -3215 6220 -3175
rect 6260 -3215 6570 -3175
rect 6610 -3215 6920 -3175
rect 6960 -3215 7270 -3175
rect 7310 -3215 7620 -3175
rect 7660 -3215 7970 -3175
rect 8010 -3215 8320 -3175
rect 8360 -3205 16090 -3175
rect 8360 -3215 12925 -3205
rect -120 -3240 12925 -3215
rect -120 -3280 -80 -3240
rect -40 -3280 270 -3240
rect 310 -3280 620 -3240
rect 660 -3280 970 -3240
rect 1010 -3280 1320 -3240
rect 1360 -3280 1670 -3240
rect 1710 -3280 2020 -3240
rect 2060 -3280 2370 -3240
rect 2410 -3280 2720 -3240
rect 2760 -3280 3070 -3240
rect 3110 -3280 3420 -3240
rect 3460 -3280 3770 -3240
rect 3810 -3280 4120 -3240
rect 4160 -3280 4470 -3240
rect 4510 -3280 4820 -3240
rect 4860 -3280 5170 -3240
rect 5210 -3280 5520 -3240
rect 5560 -3280 5870 -3240
rect 5910 -3280 6220 -3240
rect 6260 -3280 6570 -3240
rect 6610 -3280 6920 -3240
rect 6960 -3280 7270 -3240
rect 7310 -3280 7620 -3240
rect 7660 -3280 7970 -3240
rect 8010 -3280 8320 -3240
rect 8360 -3255 12925 -3240
rect 12975 -3255 13020 -3205
rect 13070 -3255 13115 -3205
rect 13165 -3255 13215 -3205
rect 13265 -3255 13315 -3205
rect 13365 -3255 13415 -3205
rect 13465 -3255 13510 -3205
rect 13560 -3255 13605 -3205
rect 13655 -3255 13725 -3205
rect 13775 -3255 13820 -3205
rect 13870 -3255 13915 -3205
rect 13965 -3255 14015 -3205
rect 14065 -3255 14115 -3205
rect 14165 -3255 14215 -3205
rect 14265 -3255 14310 -3205
rect 14360 -3255 14405 -3205
rect 14455 -3255 14525 -3205
rect 14575 -3255 14620 -3205
rect 14670 -3255 14715 -3205
rect 14765 -3255 14815 -3205
rect 14865 -3255 14915 -3205
rect 14965 -3255 15015 -3205
rect 15065 -3255 15110 -3205
rect 15160 -3255 15205 -3205
rect 15255 -3255 15325 -3205
rect 15375 -3255 15420 -3205
rect 15470 -3255 15515 -3205
rect 15565 -3255 15615 -3205
rect 15665 -3255 15715 -3205
rect 15765 -3255 15815 -3205
rect 15865 -3255 15910 -3205
rect 15960 -3255 16005 -3205
rect 16055 -3255 16090 -3205
rect 8360 -3280 16090 -3255
rect -120 -3300 16090 -3280
rect -120 -3340 -80 -3300
rect -40 -3340 270 -3300
rect 310 -3340 620 -3300
rect 660 -3340 970 -3300
rect 1010 -3340 1320 -3300
rect 1360 -3340 1670 -3300
rect 1710 -3340 2020 -3300
rect 2060 -3340 2370 -3300
rect 2410 -3340 2720 -3300
rect 2760 -3340 3070 -3300
rect 3110 -3340 3420 -3300
rect 3460 -3340 3770 -3300
rect 3810 -3340 4120 -3300
rect 4160 -3340 4470 -3300
rect 4510 -3340 4820 -3300
rect 4860 -3340 5170 -3300
rect 5210 -3340 5520 -3300
rect 5560 -3340 5870 -3300
rect 5910 -3340 6220 -3300
rect 6260 -3340 6570 -3300
rect 6610 -3340 6920 -3300
rect 6960 -3340 7270 -3300
rect 7310 -3340 7620 -3300
rect 7660 -3340 7970 -3300
rect 8010 -3340 8320 -3300
rect 8360 -3325 16090 -3300
rect 8360 -3340 12925 -3325
rect -120 -3365 12925 -3340
rect -120 -3405 -80 -3365
rect -40 -3405 270 -3365
rect 310 -3405 620 -3365
rect 660 -3405 970 -3365
rect 1010 -3405 1320 -3365
rect 1360 -3405 1670 -3365
rect 1710 -3405 2020 -3365
rect 2060 -3405 2370 -3365
rect 2410 -3405 2720 -3365
rect 2760 -3405 3070 -3365
rect 3110 -3405 3420 -3365
rect 3460 -3405 3770 -3365
rect 3810 -3405 4120 -3365
rect 4160 -3405 4470 -3365
rect 4510 -3405 4820 -3365
rect 4860 -3405 5170 -3365
rect 5210 -3405 5520 -3365
rect 5560 -3405 5870 -3365
rect 5910 -3405 6220 -3365
rect 6260 -3405 6570 -3365
rect 6610 -3405 6920 -3365
rect 6960 -3405 7270 -3365
rect 7310 -3405 7620 -3365
rect 7660 -3405 7970 -3365
rect 8010 -3405 8320 -3365
rect 8360 -3375 12925 -3365
rect 12975 -3375 13020 -3325
rect 13070 -3375 13115 -3325
rect 13165 -3375 13215 -3325
rect 13265 -3375 13315 -3325
rect 13365 -3375 13415 -3325
rect 13465 -3375 13510 -3325
rect 13560 -3375 13605 -3325
rect 13655 -3375 13725 -3325
rect 13775 -3375 13820 -3325
rect 13870 -3375 13915 -3325
rect 13965 -3375 14015 -3325
rect 14065 -3375 14115 -3325
rect 14165 -3375 14215 -3325
rect 14265 -3375 14310 -3325
rect 14360 -3375 14405 -3325
rect 14455 -3375 14525 -3325
rect 14575 -3375 14620 -3325
rect 14670 -3375 14715 -3325
rect 14765 -3375 14815 -3325
rect 14865 -3375 14915 -3325
rect 14965 -3375 15015 -3325
rect 15065 -3375 15110 -3325
rect 15160 -3375 15205 -3325
rect 15255 -3375 15325 -3325
rect 15375 -3375 15420 -3325
rect 15470 -3375 15515 -3325
rect 15565 -3375 15615 -3325
rect 15665 -3375 15715 -3325
rect 15765 -3375 15815 -3325
rect 15865 -3375 15910 -3325
rect 15960 -3375 16005 -3325
rect 16055 -3375 16090 -3325
rect 8360 -3405 16090 -3375
rect -120 -3415 16090 -3405
rect -120 -3435 12925 -3415
rect -120 -3475 -80 -3435
rect -40 -3475 270 -3435
rect 310 -3475 620 -3435
rect 660 -3475 970 -3435
rect 1010 -3475 1320 -3435
rect 1360 -3475 1670 -3435
rect 1710 -3475 2020 -3435
rect 2060 -3475 2370 -3435
rect 2410 -3475 2720 -3435
rect 2760 -3475 3070 -3435
rect 3110 -3475 3420 -3435
rect 3460 -3475 3770 -3435
rect 3810 -3475 4120 -3435
rect 4160 -3475 4470 -3435
rect 4510 -3475 4820 -3435
rect 4860 -3475 5170 -3435
rect 5210 -3475 5520 -3435
rect 5560 -3475 5870 -3435
rect 5910 -3475 6220 -3435
rect 6260 -3475 6570 -3435
rect 6610 -3475 6920 -3435
rect 6960 -3475 7270 -3435
rect 7310 -3475 7620 -3435
rect 7660 -3475 7970 -3435
rect 8010 -3475 8320 -3435
rect 8360 -3465 12925 -3435
rect 12975 -3465 13020 -3415
rect 13070 -3465 13115 -3415
rect 13165 -3465 13215 -3415
rect 13265 -3465 13315 -3415
rect 13365 -3465 13415 -3415
rect 13465 -3465 13510 -3415
rect 13560 -3465 13605 -3415
rect 13655 -3465 13725 -3415
rect 13775 -3465 13820 -3415
rect 13870 -3465 13915 -3415
rect 13965 -3465 14015 -3415
rect 14065 -3465 14115 -3415
rect 14165 -3465 14215 -3415
rect 14265 -3465 14310 -3415
rect 14360 -3465 14405 -3415
rect 14455 -3465 14525 -3415
rect 14575 -3465 14620 -3415
rect 14670 -3465 14715 -3415
rect 14765 -3465 14815 -3415
rect 14865 -3465 14915 -3415
rect 14965 -3465 15015 -3415
rect 15065 -3465 15110 -3415
rect 15160 -3465 15205 -3415
rect 15255 -3465 15325 -3415
rect 15375 -3465 15420 -3415
rect 15470 -3465 15515 -3415
rect 15565 -3465 15615 -3415
rect 15665 -3465 15715 -3415
rect 15765 -3465 15815 -3415
rect 15865 -3465 15910 -3415
rect 15960 -3465 16005 -3415
rect 16055 -3465 16090 -3415
rect 8360 -3475 16090 -3465
rect -120 -3505 16090 -3475
rect -120 -3545 -80 -3505
rect -40 -3545 270 -3505
rect 310 -3545 620 -3505
rect 660 -3545 970 -3505
rect 1010 -3545 1320 -3505
rect 1360 -3545 1670 -3505
rect 1710 -3545 2020 -3505
rect 2060 -3545 2370 -3505
rect 2410 -3545 2720 -3505
rect 2760 -3545 3070 -3505
rect 3110 -3545 3420 -3505
rect 3460 -3545 3770 -3505
rect 3810 -3545 4120 -3505
rect 4160 -3545 4470 -3505
rect 4510 -3545 4820 -3505
rect 4860 -3545 5170 -3505
rect 5210 -3545 5520 -3505
rect 5560 -3545 5870 -3505
rect 5910 -3545 6220 -3505
rect 6260 -3545 6570 -3505
rect 6610 -3545 6920 -3505
rect 6960 -3545 7270 -3505
rect 7310 -3545 7620 -3505
rect 7660 -3545 7970 -3505
rect 8010 -3545 8320 -3505
rect 8360 -3515 16090 -3505
rect 8360 -3545 12925 -3515
rect -120 -3565 12925 -3545
rect 12975 -3565 13020 -3515
rect 13070 -3565 13115 -3515
rect 13165 -3565 13215 -3515
rect 13265 -3565 13315 -3515
rect 13365 -3565 13415 -3515
rect 13465 -3565 13510 -3515
rect 13560 -3565 13605 -3515
rect 13655 -3565 13725 -3515
rect 13775 -3565 13820 -3515
rect 13870 -3565 13915 -3515
rect 13965 -3565 14015 -3515
rect 14065 -3565 14115 -3515
rect 14165 -3565 14215 -3515
rect 14265 -3565 14310 -3515
rect 14360 -3565 14405 -3515
rect 14455 -3565 14525 -3515
rect 14575 -3565 14620 -3515
rect 14670 -3565 14715 -3515
rect 14765 -3565 14815 -3515
rect 14865 -3565 14915 -3515
rect 14965 -3565 15015 -3515
rect 15065 -3565 15110 -3515
rect 15160 -3565 15205 -3515
rect 15255 -3565 15325 -3515
rect 15375 -3565 15420 -3515
rect 15470 -3565 15515 -3515
rect 15565 -3565 15615 -3515
rect 15665 -3565 15715 -3515
rect 15765 -3565 15815 -3515
rect 15865 -3565 15910 -3515
rect 15960 -3565 16005 -3515
rect 16055 -3565 16090 -3515
rect -120 -3575 16090 -3565
rect -120 -3615 -80 -3575
rect -40 -3615 270 -3575
rect 310 -3615 620 -3575
rect 660 -3615 970 -3575
rect 1010 -3615 1320 -3575
rect 1360 -3615 1670 -3575
rect 1710 -3615 2020 -3575
rect 2060 -3615 2370 -3575
rect 2410 -3615 2720 -3575
rect 2760 -3615 3070 -3575
rect 3110 -3615 3420 -3575
rect 3460 -3615 3770 -3575
rect 3810 -3615 4120 -3575
rect 4160 -3615 4470 -3575
rect 4510 -3615 4820 -3575
rect 4860 -3615 5170 -3575
rect 5210 -3615 5520 -3575
rect 5560 -3615 5870 -3575
rect 5910 -3615 6220 -3575
rect 6260 -3615 6570 -3575
rect 6610 -3615 6920 -3575
rect 6960 -3615 7270 -3575
rect 7310 -3615 7620 -3575
rect 7660 -3615 7970 -3575
rect 8010 -3615 8320 -3575
rect 8360 -3605 16090 -3575
rect 8360 -3615 12925 -3605
rect -120 -3640 12925 -3615
rect -120 -3680 -80 -3640
rect -40 -3680 270 -3640
rect 310 -3680 620 -3640
rect 660 -3680 970 -3640
rect 1010 -3680 1320 -3640
rect 1360 -3680 1670 -3640
rect 1710 -3680 2020 -3640
rect 2060 -3680 2370 -3640
rect 2410 -3680 2720 -3640
rect 2760 -3680 3070 -3640
rect 3110 -3680 3420 -3640
rect 3460 -3680 3770 -3640
rect 3810 -3680 4120 -3640
rect 4160 -3680 4470 -3640
rect 4510 -3680 4820 -3640
rect 4860 -3680 5170 -3640
rect 5210 -3680 5520 -3640
rect 5560 -3680 5870 -3640
rect 5910 -3680 6220 -3640
rect 6260 -3680 6570 -3640
rect 6610 -3680 6920 -3640
rect 6960 -3680 7270 -3640
rect 7310 -3680 7620 -3640
rect 7660 -3680 7970 -3640
rect 8010 -3680 8320 -3640
rect 8360 -3655 12925 -3640
rect 12975 -3655 13020 -3605
rect 13070 -3655 13115 -3605
rect 13165 -3655 13215 -3605
rect 13265 -3655 13315 -3605
rect 13365 -3655 13415 -3605
rect 13465 -3655 13510 -3605
rect 13560 -3655 13605 -3605
rect 13655 -3655 13725 -3605
rect 13775 -3655 13820 -3605
rect 13870 -3655 13915 -3605
rect 13965 -3655 14015 -3605
rect 14065 -3655 14115 -3605
rect 14165 -3655 14215 -3605
rect 14265 -3655 14310 -3605
rect 14360 -3655 14405 -3605
rect 14455 -3655 14525 -3605
rect 14575 -3655 14620 -3605
rect 14670 -3655 14715 -3605
rect 14765 -3655 14815 -3605
rect 14865 -3655 14915 -3605
rect 14965 -3655 15015 -3605
rect 15065 -3655 15110 -3605
rect 15160 -3655 15205 -3605
rect 15255 -3655 15325 -3605
rect 15375 -3655 15420 -3605
rect 15470 -3655 15515 -3605
rect 15565 -3655 15615 -3605
rect 15665 -3655 15715 -3605
rect 15765 -3655 15815 -3605
rect 15865 -3655 15910 -3605
rect 15960 -3655 16005 -3605
rect 16055 -3655 16090 -3605
rect 8360 -3680 16090 -3655
rect -120 -3700 16090 -3680
rect -120 -3740 -80 -3700
rect -40 -3740 270 -3700
rect 310 -3740 620 -3700
rect 660 -3740 970 -3700
rect 1010 -3740 1320 -3700
rect 1360 -3740 1670 -3700
rect 1710 -3740 2020 -3700
rect 2060 -3740 2370 -3700
rect 2410 -3740 2720 -3700
rect 2760 -3740 3070 -3700
rect 3110 -3740 3420 -3700
rect 3460 -3740 3770 -3700
rect 3810 -3740 4120 -3700
rect 4160 -3740 4470 -3700
rect 4510 -3740 4820 -3700
rect 4860 -3740 5170 -3700
rect 5210 -3740 5520 -3700
rect 5560 -3740 5870 -3700
rect 5910 -3740 6220 -3700
rect 6260 -3740 6570 -3700
rect 6610 -3740 6920 -3700
rect 6960 -3740 7270 -3700
rect 7310 -3740 7620 -3700
rect 7660 -3740 7970 -3700
rect 8010 -3740 8320 -3700
rect 8360 -3725 16090 -3700
rect 8360 -3740 12925 -3725
rect -120 -3765 12925 -3740
rect -120 -3805 -80 -3765
rect -40 -3805 270 -3765
rect 310 -3805 620 -3765
rect 660 -3805 970 -3765
rect 1010 -3805 1320 -3765
rect 1360 -3805 1670 -3765
rect 1710 -3805 2020 -3765
rect 2060 -3805 2370 -3765
rect 2410 -3805 2720 -3765
rect 2760 -3805 3070 -3765
rect 3110 -3805 3420 -3765
rect 3460 -3805 3770 -3765
rect 3810 -3805 4120 -3765
rect 4160 -3805 4470 -3765
rect 4510 -3805 4820 -3765
rect 4860 -3805 5170 -3765
rect 5210 -3805 5520 -3765
rect 5560 -3805 5870 -3765
rect 5910 -3805 6220 -3765
rect 6260 -3805 6570 -3765
rect 6610 -3805 6920 -3765
rect 6960 -3805 7270 -3765
rect 7310 -3805 7620 -3765
rect 7660 -3805 7970 -3765
rect 8010 -3805 8320 -3765
rect 8360 -3775 12925 -3765
rect 12975 -3775 13020 -3725
rect 13070 -3775 13115 -3725
rect 13165 -3775 13215 -3725
rect 13265 -3775 13315 -3725
rect 13365 -3775 13415 -3725
rect 13465 -3775 13510 -3725
rect 13560 -3775 13605 -3725
rect 13655 -3775 13725 -3725
rect 13775 -3775 13820 -3725
rect 13870 -3775 13915 -3725
rect 13965 -3775 14015 -3725
rect 14065 -3775 14115 -3725
rect 14165 -3775 14215 -3725
rect 14265 -3775 14310 -3725
rect 14360 -3775 14405 -3725
rect 14455 -3775 14525 -3725
rect 14575 -3775 14620 -3725
rect 14670 -3775 14715 -3725
rect 14765 -3775 14815 -3725
rect 14865 -3775 14915 -3725
rect 14965 -3775 15015 -3725
rect 15065 -3775 15110 -3725
rect 15160 -3775 15205 -3725
rect 15255 -3775 15325 -3725
rect 15375 -3775 15420 -3725
rect 15470 -3775 15515 -3725
rect 15565 -3775 15615 -3725
rect 15665 -3775 15715 -3725
rect 15765 -3775 15815 -3725
rect 15865 -3775 15910 -3725
rect 15960 -3775 16005 -3725
rect 16055 -3775 16090 -3725
rect 8360 -3805 16090 -3775
rect -120 -3815 16090 -3805
rect -120 -3835 12925 -3815
rect -120 -3875 -80 -3835
rect -40 -3875 270 -3835
rect 310 -3875 620 -3835
rect 660 -3875 970 -3835
rect 1010 -3875 1320 -3835
rect 1360 -3875 1670 -3835
rect 1710 -3875 2020 -3835
rect 2060 -3875 2370 -3835
rect 2410 -3875 2720 -3835
rect 2760 -3875 3070 -3835
rect 3110 -3875 3420 -3835
rect 3460 -3875 3770 -3835
rect 3810 -3875 4120 -3835
rect 4160 -3875 4470 -3835
rect 4510 -3875 4820 -3835
rect 4860 -3875 5170 -3835
rect 5210 -3875 5520 -3835
rect 5560 -3875 5870 -3835
rect 5910 -3875 6220 -3835
rect 6260 -3875 6570 -3835
rect 6610 -3875 6920 -3835
rect 6960 -3875 7270 -3835
rect 7310 -3875 7620 -3835
rect 7660 -3875 7970 -3835
rect 8010 -3875 8320 -3835
rect 8360 -3865 12925 -3835
rect 12975 -3865 13020 -3815
rect 13070 -3865 13115 -3815
rect 13165 -3865 13215 -3815
rect 13265 -3865 13315 -3815
rect 13365 -3865 13415 -3815
rect 13465 -3865 13510 -3815
rect 13560 -3865 13605 -3815
rect 13655 -3865 13725 -3815
rect 13775 -3865 13820 -3815
rect 13870 -3865 13915 -3815
rect 13965 -3865 14015 -3815
rect 14065 -3865 14115 -3815
rect 14165 -3865 14215 -3815
rect 14265 -3865 14310 -3815
rect 14360 -3865 14405 -3815
rect 14455 -3865 14525 -3815
rect 14575 -3865 14620 -3815
rect 14670 -3865 14715 -3815
rect 14765 -3865 14815 -3815
rect 14865 -3865 14915 -3815
rect 14965 -3865 15015 -3815
rect 15065 -3865 15110 -3815
rect 15160 -3865 15205 -3815
rect 15255 -3865 15325 -3815
rect 15375 -3865 15420 -3815
rect 15470 -3865 15515 -3815
rect 15565 -3865 15615 -3815
rect 15665 -3865 15715 -3815
rect 15765 -3865 15815 -3815
rect 15865 -3865 15910 -3815
rect 15960 -3865 16005 -3815
rect 16055 -3865 16090 -3815
rect 8360 -3875 16090 -3865
rect -120 -3905 16090 -3875
rect -120 -3945 -80 -3905
rect -40 -3945 270 -3905
rect 310 -3945 620 -3905
rect 660 -3945 970 -3905
rect 1010 -3945 1320 -3905
rect 1360 -3945 1670 -3905
rect 1710 -3945 2020 -3905
rect 2060 -3945 2370 -3905
rect 2410 -3945 2720 -3905
rect 2760 -3945 3070 -3905
rect 3110 -3945 3420 -3905
rect 3460 -3945 3770 -3905
rect 3810 -3945 4120 -3905
rect 4160 -3945 4470 -3905
rect 4510 -3945 4820 -3905
rect 4860 -3945 5170 -3905
rect 5210 -3945 5520 -3905
rect 5560 -3945 5870 -3905
rect 5910 -3945 6220 -3905
rect 6260 -3945 6570 -3905
rect 6610 -3945 6920 -3905
rect 6960 -3945 7270 -3905
rect 7310 -3945 7620 -3905
rect 7660 -3945 7970 -3905
rect 8010 -3945 8320 -3905
rect 8360 -3915 16090 -3905
rect 8360 -3945 12925 -3915
rect -120 -3965 12925 -3945
rect 12975 -3965 13020 -3915
rect 13070 -3965 13115 -3915
rect 13165 -3965 13215 -3915
rect 13265 -3965 13315 -3915
rect 13365 -3965 13415 -3915
rect 13465 -3965 13510 -3915
rect 13560 -3965 13605 -3915
rect 13655 -3965 13725 -3915
rect 13775 -3965 13820 -3915
rect 13870 -3965 13915 -3915
rect 13965 -3965 14015 -3915
rect 14065 -3965 14115 -3915
rect 14165 -3965 14215 -3915
rect 14265 -3965 14310 -3915
rect 14360 -3965 14405 -3915
rect 14455 -3965 14525 -3915
rect 14575 -3965 14620 -3915
rect 14670 -3965 14715 -3915
rect 14765 -3965 14815 -3915
rect 14865 -3965 14915 -3915
rect 14965 -3965 15015 -3915
rect 15065 -3965 15110 -3915
rect 15160 -3965 15205 -3915
rect 15255 -3965 15325 -3915
rect 15375 -3965 15420 -3915
rect 15470 -3965 15515 -3915
rect 15565 -3965 15615 -3915
rect 15665 -3965 15715 -3915
rect 15765 -3965 15815 -3915
rect 15865 -3965 15910 -3915
rect 15960 -3965 16005 -3915
rect 16055 -3965 16090 -3915
rect -120 -3975 16090 -3965
rect -120 -4015 -80 -3975
rect -40 -4015 270 -3975
rect 310 -4015 620 -3975
rect 660 -4015 970 -3975
rect 1010 -4015 1320 -3975
rect 1360 -4015 1670 -3975
rect 1710 -4015 2020 -3975
rect 2060 -4015 2370 -3975
rect 2410 -4015 2720 -3975
rect 2760 -4015 3070 -3975
rect 3110 -4015 3420 -3975
rect 3460 -4015 3770 -3975
rect 3810 -4015 4120 -3975
rect 4160 -4015 4470 -3975
rect 4510 -4015 4820 -3975
rect 4860 -4015 5170 -3975
rect 5210 -4015 5520 -3975
rect 5560 -4015 5870 -3975
rect 5910 -4015 6220 -3975
rect 6260 -4015 6570 -3975
rect 6610 -4015 6920 -3975
rect 6960 -4015 7270 -3975
rect 7310 -4015 7620 -3975
rect 7660 -4015 7970 -3975
rect 8010 -4015 8320 -3975
rect 8360 -4005 16090 -3975
rect 8360 -4015 12925 -4005
rect -120 -4040 12925 -4015
rect -120 -4080 -80 -4040
rect -40 -4080 270 -4040
rect 310 -4080 620 -4040
rect 660 -4080 970 -4040
rect 1010 -4080 1320 -4040
rect 1360 -4080 1670 -4040
rect 1710 -4080 2020 -4040
rect 2060 -4080 2370 -4040
rect 2410 -4080 2720 -4040
rect 2760 -4080 3070 -4040
rect 3110 -4080 3420 -4040
rect 3460 -4080 3770 -4040
rect 3810 -4080 4120 -4040
rect 4160 -4080 4470 -4040
rect 4510 -4080 4820 -4040
rect 4860 -4080 5170 -4040
rect 5210 -4080 5520 -4040
rect 5560 -4080 5870 -4040
rect 5910 -4080 6220 -4040
rect 6260 -4080 6570 -4040
rect 6610 -4080 6920 -4040
rect 6960 -4080 7270 -4040
rect 7310 -4080 7620 -4040
rect 7660 -4080 7970 -4040
rect 8010 -4080 8320 -4040
rect 8360 -4055 12925 -4040
rect 12975 -4055 13020 -4005
rect 13070 -4055 13115 -4005
rect 13165 -4055 13215 -4005
rect 13265 -4055 13315 -4005
rect 13365 -4055 13415 -4005
rect 13465 -4055 13510 -4005
rect 13560 -4055 13605 -4005
rect 13655 -4055 13725 -4005
rect 13775 -4055 13820 -4005
rect 13870 -4055 13915 -4005
rect 13965 -4055 14015 -4005
rect 14065 -4055 14115 -4005
rect 14165 -4055 14215 -4005
rect 14265 -4055 14310 -4005
rect 14360 -4055 14405 -4005
rect 14455 -4055 14525 -4005
rect 14575 -4055 14620 -4005
rect 14670 -4055 14715 -4005
rect 14765 -4055 14815 -4005
rect 14865 -4055 14915 -4005
rect 14965 -4055 15015 -4005
rect 15065 -4055 15110 -4005
rect 15160 -4055 15205 -4005
rect 15255 -4055 15325 -4005
rect 15375 -4055 15420 -4005
rect 15470 -4055 15515 -4005
rect 15565 -4055 15615 -4005
rect 15665 -4055 15715 -4005
rect 15765 -4055 15815 -4005
rect 15865 -4055 15910 -4005
rect 15960 -4055 16005 -4005
rect 16055 -4055 16090 -4005
rect 8360 -4080 16090 -4055
rect -120 -4100 16090 -4080
rect -120 -4140 -80 -4100
rect -40 -4140 270 -4100
rect 310 -4140 620 -4100
rect 660 -4140 970 -4100
rect 1010 -4140 1320 -4100
rect 1360 -4140 1670 -4100
rect 1710 -4140 2020 -4100
rect 2060 -4140 2370 -4100
rect 2410 -4140 2720 -4100
rect 2760 -4140 3070 -4100
rect 3110 -4140 3420 -4100
rect 3460 -4140 3770 -4100
rect 3810 -4140 4120 -4100
rect 4160 -4140 4470 -4100
rect 4510 -4140 4820 -4100
rect 4860 -4140 5170 -4100
rect 5210 -4140 5520 -4100
rect 5560 -4140 5870 -4100
rect 5910 -4140 6220 -4100
rect 6260 -4140 6570 -4100
rect 6610 -4140 6920 -4100
rect 6960 -4140 7270 -4100
rect 7310 -4140 7620 -4100
rect 7660 -4140 7970 -4100
rect 8010 -4140 8320 -4100
rect 8360 -4125 16090 -4100
rect 8360 -4140 12925 -4125
rect -120 -4165 12925 -4140
rect -120 -4205 -80 -4165
rect -40 -4205 270 -4165
rect 310 -4205 620 -4165
rect 660 -4205 970 -4165
rect 1010 -4205 1320 -4165
rect 1360 -4205 1670 -4165
rect 1710 -4205 2020 -4165
rect 2060 -4205 2370 -4165
rect 2410 -4205 2720 -4165
rect 2760 -4205 3070 -4165
rect 3110 -4205 3420 -4165
rect 3460 -4205 3770 -4165
rect 3810 -4205 4120 -4165
rect 4160 -4205 4470 -4165
rect 4510 -4205 4820 -4165
rect 4860 -4205 5170 -4165
rect 5210 -4205 5520 -4165
rect 5560 -4205 5870 -4165
rect 5910 -4205 6220 -4165
rect 6260 -4205 6570 -4165
rect 6610 -4205 6920 -4165
rect 6960 -4205 7270 -4165
rect 7310 -4205 7620 -4165
rect 7660 -4205 7970 -4165
rect 8010 -4205 8320 -4165
rect 8360 -4175 12925 -4165
rect 12975 -4175 13020 -4125
rect 13070 -4175 13115 -4125
rect 13165 -4175 13215 -4125
rect 13265 -4175 13315 -4125
rect 13365 -4175 13415 -4125
rect 13465 -4175 13510 -4125
rect 13560 -4175 13605 -4125
rect 13655 -4175 13725 -4125
rect 13775 -4175 13820 -4125
rect 13870 -4175 13915 -4125
rect 13965 -4175 14015 -4125
rect 14065 -4175 14115 -4125
rect 14165 -4175 14215 -4125
rect 14265 -4175 14310 -4125
rect 14360 -4175 14405 -4125
rect 14455 -4175 14525 -4125
rect 14575 -4175 14620 -4125
rect 14670 -4175 14715 -4125
rect 14765 -4175 14815 -4125
rect 14865 -4175 14915 -4125
rect 14965 -4175 15015 -4125
rect 15065 -4175 15110 -4125
rect 15160 -4175 15205 -4125
rect 15255 -4175 15325 -4125
rect 15375 -4175 15420 -4125
rect 15470 -4175 15515 -4125
rect 15565 -4175 15615 -4125
rect 15665 -4175 15715 -4125
rect 15765 -4175 15815 -4125
rect 15865 -4175 15910 -4125
rect 15960 -4175 16005 -4125
rect 16055 -4175 16090 -4125
rect 8360 -4205 16090 -4175
rect -120 -4215 16090 -4205
rect -120 -4235 12925 -4215
rect -120 -4275 -80 -4235
rect -40 -4275 270 -4235
rect 310 -4275 620 -4235
rect 660 -4275 970 -4235
rect 1010 -4275 1320 -4235
rect 1360 -4275 1670 -4235
rect 1710 -4275 2020 -4235
rect 2060 -4275 2370 -4235
rect 2410 -4275 2720 -4235
rect 2760 -4275 3070 -4235
rect 3110 -4275 3420 -4235
rect 3460 -4275 3770 -4235
rect 3810 -4275 4120 -4235
rect 4160 -4275 4470 -4235
rect 4510 -4275 4820 -4235
rect 4860 -4275 5170 -4235
rect 5210 -4275 5520 -4235
rect 5560 -4275 5870 -4235
rect 5910 -4275 6220 -4235
rect 6260 -4275 6570 -4235
rect 6610 -4275 6920 -4235
rect 6960 -4275 7270 -4235
rect 7310 -4275 7620 -4235
rect 7660 -4275 7970 -4235
rect 8010 -4275 8320 -4235
rect 8360 -4265 12925 -4235
rect 12975 -4265 13020 -4215
rect 13070 -4265 13115 -4215
rect 13165 -4265 13215 -4215
rect 13265 -4265 13315 -4215
rect 13365 -4265 13415 -4215
rect 13465 -4265 13510 -4215
rect 13560 -4265 13605 -4215
rect 13655 -4265 13725 -4215
rect 13775 -4265 13820 -4215
rect 13870 -4265 13915 -4215
rect 13965 -4265 14015 -4215
rect 14065 -4265 14115 -4215
rect 14165 -4265 14215 -4215
rect 14265 -4265 14310 -4215
rect 14360 -4265 14405 -4215
rect 14455 -4265 14525 -4215
rect 14575 -4265 14620 -4215
rect 14670 -4265 14715 -4215
rect 14765 -4265 14815 -4215
rect 14865 -4265 14915 -4215
rect 14965 -4265 15015 -4215
rect 15065 -4265 15110 -4215
rect 15160 -4265 15205 -4215
rect 15255 -4265 15325 -4215
rect 15375 -4265 15420 -4215
rect 15470 -4265 15515 -4215
rect 15565 -4265 15615 -4215
rect 15665 -4265 15715 -4215
rect 15765 -4265 15815 -4215
rect 15865 -4265 15910 -4215
rect 15960 -4265 16005 -4215
rect 16055 -4265 16090 -4215
rect 8360 -4275 16090 -4265
rect -120 -4305 16090 -4275
rect -120 -4345 -80 -4305
rect -40 -4345 270 -4305
rect 310 -4345 620 -4305
rect 660 -4345 970 -4305
rect 1010 -4345 1320 -4305
rect 1360 -4345 1670 -4305
rect 1710 -4345 2020 -4305
rect 2060 -4345 2370 -4305
rect 2410 -4345 2720 -4305
rect 2760 -4345 3070 -4305
rect 3110 -4345 3420 -4305
rect 3460 -4345 3770 -4305
rect 3810 -4345 4120 -4305
rect 4160 -4345 4470 -4305
rect 4510 -4345 4820 -4305
rect 4860 -4345 5170 -4305
rect 5210 -4345 5520 -4305
rect 5560 -4345 5870 -4305
rect 5910 -4345 6220 -4305
rect 6260 -4345 6570 -4305
rect 6610 -4345 6920 -4305
rect 6960 -4345 7270 -4305
rect 7310 -4345 7620 -4305
rect 7660 -4345 7970 -4305
rect 8010 -4345 8320 -4305
rect 8360 -4315 16090 -4305
rect 8360 -4345 12925 -4315
rect -120 -4365 12925 -4345
rect 12975 -4365 13020 -4315
rect 13070 -4365 13115 -4315
rect 13165 -4365 13215 -4315
rect 13265 -4365 13315 -4315
rect 13365 -4365 13415 -4315
rect 13465 -4365 13510 -4315
rect 13560 -4365 13605 -4315
rect 13655 -4365 13725 -4315
rect 13775 -4365 13820 -4315
rect 13870 -4365 13915 -4315
rect 13965 -4365 14015 -4315
rect 14065 -4365 14115 -4315
rect 14165 -4365 14215 -4315
rect 14265 -4365 14310 -4315
rect 14360 -4365 14405 -4315
rect 14455 -4365 14525 -4315
rect 14575 -4365 14620 -4315
rect 14670 -4365 14715 -4315
rect 14765 -4365 14815 -4315
rect 14865 -4365 14915 -4315
rect 14965 -4365 15015 -4315
rect 15065 -4365 15110 -4315
rect 15160 -4365 15205 -4315
rect 15255 -4365 15325 -4315
rect 15375 -4365 15420 -4315
rect 15470 -4365 15515 -4315
rect 15565 -4365 15615 -4315
rect 15665 -4365 15715 -4315
rect 15765 -4365 15815 -4315
rect 15865 -4365 15910 -4315
rect 15960 -4365 16005 -4315
rect 16055 -4365 16090 -4315
rect -120 -4375 16090 -4365
rect -120 -4415 -80 -4375
rect -40 -4415 270 -4375
rect 310 -4415 620 -4375
rect 660 -4415 970 -4375
rect 1010 -4415 1320 -4375
rect 1360 -4415 1670 -4375
rect 1710 -4415 2020 -4375
rect 2060 -4415 2370 -4375
rect 2410 -4415 2720 -4375
rect 2760 -4415 3070 -4375
rect 3110 -4415 3420 -4375
rect 3460 -4415 3770 -4375
rect 3810 -4415 4120 -4375
rect 4160 -4415 4470 -4375
rect 4510 -4415 4820 -4375
rect 4860 -4415 5170 -4375
rect 5210 -4415 5520 -4375
rect 5560 -4415 5870 -4375
rect 5910 -4415 6220 -4375
rect 6260 -4415 6570 -4375
rect 6610 -4415 6920 -4375
rect 6960 -4415 7270 -4375
rect 7310 -4415 7620 -4375
rect 7660 -4415 7970 -4375
rect 8010 -4415 8320 -4375
rect 8360 -4405 16090 -4375
rect 8360 -4415 12925 -4405
rect -120 -4440 12925 -4415
rect -120 -4480 -80 -4440
rect -40 -4480 270 -4440
rect 310 -4480 620 -4440
rect 660 -4480 970 -4440
rect 1010 -4480 1320 -4440
rect 1360 -4480 1670 -4440
rect 1710 -4480 2020 -4440
rect 2060 -4480 2370 -4440
rect 2410 -4480 2720 -4440
rect 2760 -4480 3070 -4440
rect 3110 -4480 3420 -4440
rect 3460 -4480 3770 -4440
rect 3810 -4480 4120 -4440
rect 4160 -4480 4470 -4440
rect 4510 -4480 4820 -4440
rect 4860 -4480 5170 -4440
rect 5210 -4480 5520 -4440
rect 5560 -4480 5870 -4440
rect 5910 -4480 6220 -4440
rect 6260 -4480 6570 -4440
rect 6610 -4480 6920 -4440
rect 6960 -4480 7270 -4440
rect 7310 -4480 7620 -4440
rect 7660 -4480 7970 -4440
rect 8010 -4480 8320 -4440
rect 8360 -4455 12925 -4440
rect 12975 -4455 13020 -4405
rect 13070 -4455 13115 -4405
rect 13165 -4455 13215 -4405
rect 13265 -4455 13315 -4405
rect 13365 -4455 13415 -4405
rect 13465 -4455 13510 -4405
rect 13560 -4455 13605 -4405
rect 13655 -4455 13725 -4405
rect 13775 -4455 13820 -4405
rect 13870 -4455 13915 -4405
rect 13965 -4455 14015 -4405
rect 14065 -4455 14115 -4405
rect 14165 -4455 14215 -4405
rect 14265 -4455 14310 -4405
rect 14360 -4455 14405 -4405
rect 14455 -4455 14525 -4405
rect 14575 -4455 14620 -4405
rect 14670 -4455 14715 -4405
rect 14765 -4455 14815 -4405
rect 14865 -4455 14915 -4405
rect 14965 -4455 15015 -4405
rect 15065 -4455 15110 -4405
rect 15160 -4455 15205 -4405
rect 15255 -4455 15325 -4405
rect 15375 -4455 15420 -4405
rect 15470 -4455 15515 -4405
rect 15565 -4455 15615 -4405
rect 15665 -4455 15715 -4405
rect 15765 -4455 15815 -4405
rect 15865 -4455 15910 -4405
rect 15960 -4455 16005 -4405
rect 16055 -4455 16090 -4405
rect 8360 -4480 16090 -4455
rect -120 -4490 16090 -4480
use bgr_11  bgr_11_0
timestamp 1754396681
transform -1 0 22290 0 -1 11485
box 15665 -6150 19905 1795
use two_stage_opamp_dummy_magic_24  two_stage_opamp_dummy_magic_24_0
timestamp 1754401177
transform 1 0 -52410 0 1 100
box 52060 -1500 61740 6110
<< labels >>
flabel metal3 -2040 10155 -2040 10155 1 FreeSans 800 0 0 320 VDDA
port 1 n
flabel metal2 5375 1380 5375 1380 3 FreeSans 400 0 160 0 VIN-
port 6 e
flabel metal2 3605 1380 3605 1380 7 FreeSans 400 0 -160 0 VIN+
port 5 w
flabel metal2 6795 455 6795 455 5 FreeSans 400 0 0 -160 VOUT-
port 4 s
flabel metal2 1960 455 1960 455 5 FreeSans 400 0 0 -160 VOUT+
port 3 s
flabel metal4 18820 6650 18820 6650 3 FreeSans 800 0 320 0 GNDA
port 2 e
<< end >>
