magic
tech sky130A
timestamp 1738585014
<< nwell >>
rect 4010 2230 5060 2750
<< nmos >>
rect 4080 1925 4095 1975
rect 4145 1925 4160 1975
rect 4210 1925 4225 1975
rect 4275 1925 4290 1975
rect 4440 1925 4455 1975
rect 4505 1925 4520 1975
rect 4570 1925 4585 1975
rect 4635 1925 4650 1975
rect 4780 1925 4795 1975
rect 4845 1925 4860 1975
rect 4910 1925 4925 1975
rect 4975 1925 4990 1975
rect 4590 1545 4640 1795
rect 4690 1545 4740 1795
rect 4790 1545 4840 1795
rect 4890 1545 4940 1795
<< pmos >>
rect 4095 2445 4145 2695
rect 4195 2445 4245 2695
rect 4295 2445 4345 2695
rect 4395 2445 4445 2695
rect 4495 2445 4545 2695
rect 4595 2445 4645 2695
rect 4695 2445 4745 2695
rect 4795 2445 4845 2695
rect 4080 2255 4095 2355
rect 4145 2255 4160 2355
rect 4210 2255 4225 2355
rect 4275 2255 4290 2355
rect 4440 2255 4455 2355
rect 4505 2255 4520 2355
rect 4570 2255 4585 2355
rect 4635 2255 4650 2355
rect 4780 2255 4795 2355
rect 4845 2255 4860 2355
rect 4910 2255 4925 2355
rect 4975 2255 4990 2355
<< ndiff >>
rect 4030 1960 4080 1975
rect 4030 1940 4045 1960
rect 4065 1940 4080 1960
rect 4030 1925 4080 1940
rect 4095 1960 4145 1975
rect 4095 1940 4110 1960
rect 4130 1940 4145 1960
rect 4095 1925 4145 1940
rect 4160 1960 4210 1975
rect 4160 1940 4175 1960
rect 4195 1940 4210 1960
rect 4160 1925 4210 1940
rect 4225 1960 4275 1975
rect 4225 1940 4240 1960
rect 4260 1940 4275 1960
rect 4225 1925 4275 1940
rect 4290 1960 4340 1975
rect 4290 1940 4305 1960
rect 4325 1940 4340 1960
rect 4290 1925 4340 1940
rect 4390 1960 4440 1975
rect 4390 1940 4405 1960
rect 4425 1940 4440 1960
rect 4390 1925 4440 1940
rect 4455 1960 4505 1975
rect 4455 1940 4470 1960
rect 4490 1940 4505 1960
rect 4455 1925 4505 1940
rect 4520 1960 4570 1975
rect 4520 1940 4535 1960
rect 4555 1940 4570 1960
rect 4520 1925 4570 1940
rect 4585 1960 4635 1975
rect 4585 1940 4600 1960
rect 4620 1940 4635 1960
rect 4585 1925 4635 1940
rect 4650 1960 4700 1975
rect 4650 1940 4665 1960
rect 4685 1940 4700 1960
rect 4650 1925 4700 1940
rect 4730 1960 4780 1975
rect 4730 1940 4745 1960
rect 4765 1940 4780 1960
rect 4730 1925 4780 1940
rect 4795 1960 4845 1975
rect 4795 1940 4810 1960
rect 4830 1940 4845 1960
rect 4795 1925 4845 1940
rect 4860 1960 4910 1975
rect 4860 1940 4875 1960
rect 4895 1940 4910 1960
rect 4860 1925 4910 1940
rect 4925 1960 4975 1975
rect 4925 1940 4940 1960
rect 4960 1940 4975 1960
rect 4925 1925 4975 1940
rect 4990 1960 5040 1975
rect 4990 1940 5005 1960
rect 5025 1940 5040 1960
rect 4990 1925 5040 1940
rect 4540 1780 4590 1795
rect 4540 1560 4555 1780
rect 4575 1560 4590 1780
rect 4540 1545 4590 1560
rect 4640 1780 4690 1795
rect 4640 1560 4655 1780
rect 4675 1560 4690 1780
rect 4640 1545 4690 1560
rect 4740 1780 4790 1795
rect 4740 1560 4755 1780
rect 4775 1560 4790 1780
rect 4740 1545 4790 1560
rect 4840 1780 4890 1795
rect 4840 1560 4855 1780
rect 4875 1560 4890 1780
rect 4840 1545 4890 1560
rect 4940 1780 4990 1795
rect 4940 1560 4955 1780
rect 4975 1560 4990 1780
rect 4940 1545 4990 1560
<< pdiff >>
rect 4045 2680 4095 2695
rect 4045 2460 4060 2680
rect 4080 2460 4095 2680
rect 4045 2445 4095 2460
rect 4145 2680 4195 2695
rect 4145 2460 4160 2680
rect 4180 2460 4195 2680
rect 4145 2445 4195 2460
rect 4245 2680 4295 2695
rect 4245 2460 4260 2680
rect 4280 2460 4295 2680
rect 4245 2445 4295 2460
rect 4345 2680 4395 2695
rect 4345 2460 4360 2680
rect 4380 2460 4395 2680
rect 4345 2445 4395 2460
rect 4445 2680 4495 2695
rect 4445 2460 4460 2680
rect 4480 2460 4495 2680
rect 4445 2445 4495 2460
rect 4545 2680 4595 2695
rect 4545 2460 4560 2680
rect 4580 2460 4595 2680
rect 4545 2445 4595 2460
rect 4645 2680 4695 2695
rect 4645 2460 4660 2680
rect 4680 2460 4695 2680
rect 4645 2445 4695 2460
rect 4745 2680 4795 2695
rect 4745 2460 4760 2680
rect 4780 2460 4795 2680
rect 4745 2445 4795 2460
rect 4845 2680 4895 2695
rect 4845 2460 4860 2680
rect 4880 2460 4895 2680
rect 4845 2445 4895 2460
rect 4030 2340 4080 2355
rect 4030 2270 4045 2340
rect 4065 2270 4080 2340
rect 4030 2255 4080 2270
rect 4095 2340 4145 2355
rect 4095 2270 4110 2340
rect 4130 2270 4145 2340
rect 4095 2255 4145 2270
rect 4160 2340 4210 2355
rect 4160 2270 4175 2340
rect 4195 2270 4210 2340
rect 4160 2255 4210 2270
rect 4225 2340 4275 2355
rect 4225 2270 4240 2340
rect 4260 2270 4275 2340
rect 4225 2255 4275 2270
rect 4290 2340 4340 2355
rect 4290 2270 4305 2340
rect 4325 2270 4340 2340
rect 4290 2255 4340 2270
rect 4390 2340 4440 2355
rect 4390 2270 4405 2340
rect 4425 2270 4440 2340
rect 4390 2255 4440 2270
rect 4455 2340 4505 2355
rect 4455 2270 4470 2340
rect 4490 2270 4505 2340
rect 4455 2255 4505 2270
rect 4520 2340 4570 2355
rect 4520 2270 4535 2340
rect 4555 2270 4570 2340
rect 4520 2255 4570 2270
rect 4585 2340 4635 2355
rect 4585 2270 4600 2340
rect 4620 2270 4635 2340
rect 4585 2255 4635 2270
rect 4650 2340 4700 2355
rect 4650 2270 4665 2340
rect 4685 2270 4700 2340
rect 4650 2255 4700 2270
rect 4730 2340 4780 2355
rect 4730 2270 4745 2340
rect 4765 2270 4780 2340
rect 4730 2255 4780 2270
rect 4795 2340 4845 2355
rect 4795 2270 4810 2340
rect 4830 2270 4845 2340
rect 4795 2255 4845 2270
rect 4860 2340 4910 2355
rect 4860 2270 4875 2340
rect 4895 2270 4910 2340
rect 4860 2255 4910 2270
rect 4925 2340 4975 2355
rect 4925 2270 4940 2340
rect 4960 2270 4975 2340
rect 4925 2255 4975 2270
rect 4990 2340 5040 2355
rect 4990 2270 5005 2340
rect 5025 2270 5040 2340
rect 4990 2255 5040 2270
<< ndiffc >>
rect 4045 1940 4065 1960
rect 4110 1940 4130 1960
rect 4175 1940 4195 1960
rect 4240 1940 4260 1960
rect 4305 1940 4325 1960
rect 4405 1940 4425 1960
rect 4470 1940 4490 1960
rect 4535 1940 4555 1960
rect 4600 1940 4620 1960
rect 4665 1940 4685 1960
rect 4745 1940 4765 1960
rect 4810 1940 4830 1960
rect 4875 1940 4895 1960
rect 4940 1940 4960 1960
rect 5005 1940 5025 1960
rect 4555 1560 4575 1780
rect 4655 1560 4675 1780
rect 4755 1560 4775 1780
rect 4855 1560 4875 1780
rect 4955 1560 4975 1780
<< pdiffc >>
rect 4060 2460 4080 2680
rect 4160 2460 4180 2680
rect 4260 2460 4280 2680
rect 4360 2460 4380 2680
rect 4460 2460 4480 2680
rect 4560 2460 4580 2680
rect 4660 2460 4680 2680
rect 4760 2460 4780 2680
rect 4860 2460 4880 2680
rect 4045 2270 4065 2340
rect 4110 2270 4130 2340
rect 4175 2270 4195 2340
rect 4240 2270 4260 2340
rect 4305 2270 4325 2340
rect 4405 2270 4425 2340
rect 4470 2270 4490 2340
rect 4535 2270 4555 2340
rect 4600 2270 4620 2340
rect 4665 2270 4685 2340
rect 4745 2270 4765 2340
rect 4810 2270 4830 2340
rect 4875 2270 4895 2340
rect 4940 2270 4960 2340
rect 5005 2270 5025 2340
<< psubdiff >>
rect 4160 1880 4210 1895
rect 4160 1860 4175 1880
rect 4195 1860 4210 1880
rect 4160 1845 4210 1860
rect 4220 1410 4270 1460
<< nsubdiff >>
rect 4940 2680 4990 2695
rect 4940 2460 4955 2680
rect 4975 2460 4990 2680
rect 4940 2445 4990 2460
<< psubdiffcont >>
rect 4175 1860 4195 1880
<< nsubdiffcont >>
rect 4955 2460 4975 2680
<< poly >>
rect 4075 2740 4115 2750
rect 4075 2720 4085 2740
rect 4105 2720 4115 2740
rect 4450 2740 4490 2750
rect 4450 2720 4460 2740
rect 4480 2720 4490 2740
rect 4830 2740 4870 2750
rect 4830 2720 4840 2740
rect 4860 2720 4870 2740
rect 4075 2710 4870 2720
rect 4095 2705 4845 2710
rect 4095 2695 4145 2705
rect 4195 2695 4245 2705
rect 4295 2695 4345 2705
rect 4395 2695 4445 2705
rect 4495 2695 4545 2705
rect 4595 2695 4645 2705
rect 4695 2695 4745 2705
rect 4795 2695 4845 2705
rect 4095 2430 4145 2445
rect 4195 2430 4245 2445
rect 4295 2430 4345 2445
rect 4395 2430 4445 2445
rect 4495 2430 4545 2445
rect 4595 2430 4645 2445
rect 4695 2430 4745 2445
rect 4795 2430 4845 2445
rect 3660 2365 4160 2380
rect 3770 2070 3785 2365
rect 4080 2355 4095 2365
rect 4145 2355 4160 2365
rect 4210 2355 4225 2370
rect 4275 2355 4290 2370
rect 4440 2355 4455 2370
rect 4505 2355 4520 2370
rect 4570 2355 4585 2370
rect 4635 2355 4650 2370
rect 4780 2355 4795 2370
rect 4845 2355 4860 2370
rect 4910 2355 4925 2370
rect 4975 2355 4990 2370
rect 4080 2240 4095 2255
rect 4145 2240 4160 2255
rect 4210 2215 4225 2255
rect 4275 2215 4290 2255
rect 4440 2245 4455 2255
rect 4505 2245 4520 2255
rect 4570 2245 4585 2255
rect 4635 2245 4650 2255
rect 4440 2240 4650 2245
rect 4780 2245 4795 2255
rect 4845 2245 4860 2255
rect 4910 2245 4925 2255
rect 4975 2245 4990 2255
rect 4410 2230 4685 2240
rect 3875 2205 4385 2215
rect 3875 2200 4355 2205
rect 4345 2185 4355 2200
rect 4375 2185 4385 2205
rect 4410 2210 4420 2230
rect 4440 2225 4655 2230
rect 4440 2210 4450 2225
rect 4410 2200 4450 2210
rect 4645 2210 4655 2225
rect 4675 2210 4685 2230
rect 4645 2200 4685 2210
rect 4780 2230 5130 2245
rect 4780 2210 4790 2230
rect 4810 2210 4820 2230
rect 4780 2200 4820 2210
rect 4345 2175 4385 2185
rect 4175 2125 4215 2135
rect 4175 2105 4185 2125
rect 4205 2110 4215 2125
rect 4205 2105 4795 2110
rect 4175 2095 4795 2105
rect 3770 2055 4520 2070
rect 4045 2020 4085 2030
rect 4045 2000 4055 2020
rect 4075 2005 4085 2020
rect 4285 2020 4325 2030
rect 4285 2005 4295 2020
rect 4075 2000 4295 2005
rect 4315 2000 4325 2020
rect 4045 1990 4325 2000
rect 4080 1985 4290 1990
rect 4080 1975 4095 1985
rect 4145 1975 4160 1985
rect 4210 1975 4225 1985
rect 4275 1975 4290 1985
rect 4440 1975 4455 2055
rect 4505 1975 4520 2055
rect 4780 2000 4795 2095
rect 4570 1975 4585 1990
rect 4635 1975 4650 1990
rect 4780 1985 5090 2000
rect 4780 1975 4795 1985
rect 4845 1975 4860 1985
rect 4910 1975 4925 1985
rect 4975 1975 4990 1985
rect 4080 1910 4095 1925
rect 4145 1910 4160 1925
rect 4210 1910 4225 1925
rect 4275 1910 4290 1925
rect 4440 1910 4455 1925
rect 4505 1910 4520 1925
rect 4335 1890 4375 1900
rect 4335 1870 4345 1890
rect 4365 1885 4375 1890
rect 4570 1885 4585 1925
rect 4635 1885 4650 1925
rect 4780 1910 4795 1925
rect 4845 1910 4860 1925
rect 4910 1910 4925 1925
rect 4975 1910 4990 1925
rect 4365 1870 4650 1885
rect 4335 1860 4375 1870
rect 4590 1795 4640 1810
rect 4690 1795 4740 1810
rect 4790 1795 4840 1810
rect 4890 1795 4940 1810
rect 4590 1535 4640 1545
rect 4690 1535 4740 1545
rect 4790 1535 4840 1545
rect 4890 1535 4940 1545
rect 4590 1525 4940 1535
rect 4590 1520 4605 1525
rect 4595 1505 4605 1520
rect 4625 1520 4905 1525
rect 4625 1505 4635 1520
rect 4595 1495 4635 1505
rect 4895 1505 4905 1520
rect 4925 1520 4940 1525
rect 4925 1505 4935 1520
rect 4895 1495 4935 1505
rect 5075 1365 5090 1985
rect 4695 1350 5090 1365
rect 4505 1255 4545 1265
rect 4505 1235 4515 1255
rect 4535 1240 4545 1255
rect 4695 1240 4710 1350
rect 5115 1325 5130 2230
rect 4940 1310 5130 1325
rect 4940 1265 4955 1310
rect 4535 1235 4710 1240
rect 4505 1225 4710 1235
rect 4935 1255 4975 1265
rect 4935 1235 4945 1255
rect 4965 1235 4975 1255
rect 4935 1225 4975 1235
<< polycont >>
rect 4085 2720 4105 2740
rect 4460 2720 4480 2740
rect 4840 2720 4860 2740
rect 4355 2185 4375 2205
rect 4420 2210 4440 2230
rect 4655 2210 4675 2230
rect 4790 2210 4810 2230
rect 4185 2105 4205 2125
rect 4055 2000 4075 2020
rect 4295 2000 4315 2020
rect 4345 1870 4365 1890
rect 4605 1505 4625 1525
rect 4905 1505 4925 1525
rect 4515 1235 4535 1255
rect 4945 1235 4965 1255
<< xpolycontact >>
rect 4010 1510 4230 1795
rect 4265 1510 4485 1795
rect 3880 1225 4100 1260
rect 4170 1225 4390 1260
rect 5025 1225 5245 1260
rect 5343 1225 5563 1260
<< xpolyres >>
rect 4230 1510 4265 1795
rect 4100 1225 4170 1260
rect 5245 1225 5343 1260
<< locali >>
rect 4075 2740 4115 2750
rect 4075 2735 4085 2740
rect 3940 2720 4085 2735
rect 4105 2735 4115 2740
rect 4450 2740 4490 2750
rect 4450 2735 4460 2740
rect 4105 2720 4460 2735
rect 4480 2735 4490 2740
rect 4830 2740 4870 2750
rect 4830 2735 4840 2740
rect 4480 2720 4840 2735
rect 4860 2735 4870 2740
rect 4860 2720 4880 2735
rect 3940 2715 4880 2720
rect 3940 1795 3960 2715
rect 4060 2710 4115 2715
rect 4450 2710 4490 2715
rect 4830 2710 4880 2715
rect 4060 2690 4080 2710
rect 4460 2690 4480 2710
rect 4860 2690 4880 2710
rect 4045 2680 4090 2690
rect 4045 2460 4060 2680
rect 4080 2460 4090 2680
rect 4045 2450 4090 2460
rect 4150 2680 4190 2690
rect 4150 2460 4160 2680
rect 4180 2460 4190 2680
rect 4150 2450 4190 2460
rect 4250 2680 4290 2690
rect 4250 2460 4260 2680
rect 4280 2460 4290 2680
rect 4250 2450 4290 2460
rect 4350 2680 4390 2690
rect 4350 2460 4360 2680
rect 4380 2460 4390 2680
rect 4350 2450 4390 2460
rect 4450 2680 4490 2690
rect 4450 2460 4460 2680
rect 4480 2460 4490 2680
rect 4450 2450 4490 2460
rect 4550 2680 4590 2690
rect 4550 2460 4560 2680
rect 4580 2460 4590 2680
rect 4550 2450 4590 2460
rect 4650 2680 4690 2690
rect 4650 2460 4660 2680
rect 4680 2460 4690 2680
rect 4650 2450 4690 2460
rect 4750 2680 4790 2690
rect 4750 2460 4760 2680
rect 4780 2460 4790 2680
rect 4750 2450 4790 2460
rect 4850 2680 4890 2690
rect 4850 2460 4860 2680
rect 4880 2460 4890 2680
rect 4850 2450 4890 2460
rect 4945 2680 4985 2690
rect 4945 2460 4955 2680
rect 4975 2460 4985 2680
rect 4945 2450 4985 2460
rect 4260 2430 4280 2450
rect 4660 2430 4680 2450
rect 4125 2410 4680 2430
rect 4125 2390 4145 2410
rect 4045 2370 4325 2390
rect 4045 2350 4065 2370
rect 4175 2350 4195 2370
rect 4305 2350 4325 2370
rect 4745 2370 5025 2390
rect 4745 2350 4765 2370
rect 4875 2350 4895 2370
rect 5005 2350 5025 2370
rect 4035 2340 4075 2350
rect 4035 2270 4045 2340
rect 4065 2270 4075 2340
rect 4035 2260 4075 2270
rect 4100 2340 4140 2350
rect 4100 2270 4110 2340
rect 4130 2270 4140 2340
rect 4100 2260 4140 2270
rect 4165 2340 4205 2350
rect 4165 2270 4175 2340
rect 4195 2270 4205 2340
rect 4165 2260 4205 2270
rect 4230 2340 4270 2350
rect 4230 2270 4240 2340
rect 4260 2270 4270 2340
rect 4230 2260 4270 2270
rect 4295 2340 4340 2350
rect 4295 2270 4305 2340
rect 4325 2270 4340 2340
rect 4295 2260 4340 2270
rect 4395 2340 4435 2350
rect 4395 2270 4405 2340
rect 4425 2270 4435 2340
rect 4395 2260 4435 2270
rect 4460 2340 4500 2350
rect 4460 2270 4470 2340
rect 4490 2270 4500 2340
rect 4460 2260 4500 2270
rect 4525 2340 4565 2350
rect 4525 2270 4535 2340
rect 4555 2270 4565 2340
rect 4525 2260 4565 2270
rect 4590 2340 4635 2350
rect 4590 2270 4600 2340
rect 4620 2270 4635 2340
rect 4590 2260 4635 2270
rect 4655 2340 4695 2350
rect 4655 2270 4665 2340
rect 4685 2270 4695 2340
rect 4655 2260 4695 2270
rect 4735 2340 4775 2350
rect 4735 2270 4745 2340
rect 4765 2270 4775 2340
rect 4735 2260 4775 2270
rect 4800 2340 4840 2350
rect 4800 2270 4810 2340
rect 4830 2270 4840 2340
rect 4800 2260 4840 2270
rect 4865 2340 4905 2350
rect 4865 2270 4875 2340
rect 4895 2270 4905 2340
rect 4865 2260 4905 2270
rect 4930 2340 4970 2350
rect 4930 2270 4940 2340
rect 4960 2270 4970 2340
rect 4930 2260 4970 2270
rect 4995 2340 5035 2350
rect 4995 2270 5005 2340
rect 5025 2270 5035 2340
rect 4995 2260 5035 2270
rect 4110 2175 4130 2260
rect 4240 2175 4260 2260
rect 4405 2240 4430 2260
rect 4410 2230 4450 2240
rect 4345 2205 4385 2215
rect 4345 2185 4355 2205
rect 4375 2185 4385 2205
rect 4410 2210 4420 2230
rect 4440 2210 4450 2230
rect 4410 2200 4450 2210
rect 4345 2175 4385 2185
rect 4415 2175 4435 2200
rect 4055 2150 4130 2175
rect 4185 2155 4260 2175
rect 4055 2030 4075 2150
rect 4185 2135 4205 2155
rect 4175 2125 4215 2135
rect 4175 2105 4185 2125
rect 4205 2105 4215 2125
rect 4175 2095 4215 2105
rect 4045 2020 4085 2030
rect 4045 2000 4055 2020
rect 4075 2000 4085 2020
rect 4045 1990 4085 2000
rect 4045 1970 4065 1990
rect 4175 1970 4195 2095
rect 4285 2020 4325 2030
rect 4285 2000 4295 2020
rect 4315 2000 4325 2020
rect 4285 1990 4325 2000
rect 4305 1970 4325 1990
rect 4035 1960 4075 1970
rect 4035 1940 4045 1960
rect 4065 1940 4075 1960
rect 4035 1930 4075 1940
rect 4100 1960 4140 1970
rect 4100 1940 4110 1960
rect 4130 1940 4140 1960
rect 4100 1930 4140 1940
rect 4165 1960 4205 1970
rect 4165 1940 4175 1960
rect 4195 1940 4205 1960
rect 4165 1930 4205 1940
rect 4230 1960 4270 1970
rect 4230 1940 4240 1960
rect 4260 1940 4270 1960
rect 4230 1930 4270 1940
rect 4295 1960 4335 1970
rect 4295 1940 4305 1960
rect 4325 1940 4335 1960
rect 4295 1930 4335 1940
rect 4110 1880 4130 1930
rect 4165 1880 4205 1890
rect 4240 1880 4260 1930
rect 4355 1900 4375 2175
rect 4415 2155 4490 2175
rect 4470 1970 4490 2155
rect 4535 2165 4555 2260
rect 4665 2240 4685 2260
rect 5005 2240 5025 2260
rect 4645 2230 4685 2240
rect 4645 2210 4655 2230
rect 4675 2210 4685 2230
rect 4645 2200 4685 2210
rect 4780 2230 4820 2240
rect 4780 2210 4790 2230
rect 4810 2210 4820 2230
rect 5005 2220 5140 2240
rect 4780 2200 4820 2210
rect 4780 2165 4800 2200
rect 4535 2145 4800 2165
rect 4600 1970 4620 2145
rect 4395 1960 4435 1970
rect 4395 1940 4405 1960
rect 4425 1940 4435 1960
rect 4395 1930 4435 1940
rect 4460 1960 4500 1970
rect 4460 1940 4470 1960
rect 4490 1940 4500 1960
rect 4460 1930 4500 1940
rect 4525 1960 4565 1970
rect 4525 1940 4535 1960
rect 4555 1940 4565 1960
rect 4525 1930 4565 1940
rect 4590 1960 4630 1970
rect 4590 1940 4600 1960
rect 4620 1940 4630 1960
rect 4590 1930 4630 1940
rect 4655 1960 4695 1970
rect 4655 1940 4665 1960
rect 4685 1940 4695 1960
rect 4655 1930 4695 1940
rect 4735 1960 4775 1970
rect 4735 1940 4745 1960
rect 4765 1940 4775 1960
rect 4735 1930 4775 1940
rect 4800 1960 4840 1970
rect 4800 1940 4810 1960
rect 4830 1940 4840 1960
rect 4800 1930 4840 1940
rect 4865 1960 4905 1970
rect 4865 1940 4875 1960
rect 4895 1940 4905 1960
rect 4865 1930 4905 1940
rect 4930 1960 4970 1970
rect 4930 1940 4940 1960
rect 4960 1940 4970 1960
rect 4930 1930 4970 1940
rect 4995 1960 5035 1970
rect 4995 1940 5005 1960
rect 5025 1940 5035 1960
rect 4995 1930 5035 1940
rect 4110 1860 4175 1880
rect 4195 1860 4260 1880
rect 4335 1890 4375 1900
rect 4405 1910 4425 1930
rect 4535 1910 4555 1930
rect 4665 1910 4685 1930
rect 4405 1890 4685 1910
rect 4745 1910 4765 1930
rect 4875 1910 4895 1930
rect 5005 1910 5025 1930
rect 4745 1905 5025 1910
rect 4335 1870 4345 1890
rect 4365 1870 4375 1890
rect 4335 1860 4375 1870
rect 4165 1850 4205 1860
rect 4535 1830 4555 1890
rect 4745 1885 5100 1905
rect 4535 1810 4775 1830
rect 3940 1775 4010 1795
rect 4755 1790 4775 1810
rect 4545 1780 4585 1790
rect 4545 1560 4555 1780
rect 4575 1560 4585 1780
rect 4545 1550 4585 1560
rect 4645 1780 4685 1790
rect 4645 1560 4655 1780
rect 4675 1560 4685 1780
rect 4645 1550 4685 1560
rect 4745 1780 4785 1790
rect 4745 1560 4755 1780
rect 4775 1560 4785 1780
rect 4745 1550 4785 1560
rect 4845 1780 4885 1790
rect 4845 1560 4855 1780
rect 4875 1560 4885 1780
rect 4845 1550 4885 1560
rect 4945 1780 4985 1790
rect 4945 1560 4955 1780
rect 4975 1560 4985 1780
rect 4945 1550 4985 1560
rect 4555 1530 4575 1550
rect 4595 1530 4635 1535
rect 4895 1530 4935 1535
rect 4955 1530 4975 1550
rect 4485 1525 4975 1530
rect 4485 1510 4605 1525
rect 4595 1505 4605 1510
rect 4625 1510 4905 1525
rect 4625 1505 4635 1510
rect 4595 1495 4635 1505
rect 4895 1505 4905 1510
rect 4925 1510 4975 1525
rect 4925 1505 4935 1510
rect 4895 1495 4935 1505
rect 4225 1445 4265 1455
rect 4225 1425 4235 1445
rect 4255 1425 4265 1445
rect 4225 1415 4265 1425
rect 5080 1345 5100 1885
rect 4740 1325 5100 1345
rect 3685 1225 3880 1245
rect 4505 1255 4545 1265
rect 4505 1245 4515 1255
rect 4390 1235 4515 1245
rect 4535 1235 4545 1255
rect 4390 1225 4545 1235
rect 3685 1205 3705 1225
rect 4740 1205 4760 1325
rect 5120 1305 5140 2220
rect 3665 1195 3715 1205
rect 3665 1165 3675 1195
rect 3705 1165 3715 1195
rect 3665 1155 3715 1165
rect 4630 1195 4760 1205
rect 4630 1160 4640 1195
rect 4675 1185 4760 1195
rect 4675 1160 4685 1185
rect 4630 1150 4685 1160
rect 4740 1120 4760 1185
rect 4820 1285 5140 1305
rect 4820 1205 4840 1285
rect 4935 1260 4975 1265
rect 4935 1255 5025 1260
rect 4935 1235 4945 1255
rect 4965 1240 5025 1255
rect 4965 1235 4975 1240
rect 4935 1225 4975 1235
rect 5563 1225 5880 1245
rect 5860 1205 5880 1225
rect 4820 1195 4935 1205
rect 4820 1185 4890 1195
rect 4820 1120 4840 1185
rect 4880 1160 4890 1185
rect 4925 1160 4935 1195
rect 4880 1150 4935 1160
rect 5850 1195 5900 1205
rect 5850 1165 5860 1195
rect 5890 1165 5900 1195
rect 5850 1155 5900 1165
rect 4740 1101 4840 1120
rect 4740 1100 4805 1101
<< viali >>
rect 4160 2460 4180 2680
rect 4360 2460 4380 2680
rect 4560 2460 4580 2680
rect 4760 2460 4780 2680
rect 4955 2460 4975 2680
rect 4470 2270 4490 2340
rect 4600 2270 4620 2340
rect 4810 2270 4830 2340
rect 4940 2270 4960 2340
rect 4110 1940 4130 1960
rect 4240 1940 4260 1960
rect 4810 1940 4830 1960
rect 4940 1940 4960 1960
rect 4175 1860 4195 1880
rect 4655 1560 4675 1780
rect 4855 1560 4875 1780
rect 4235 1425 4255 1445
rect 3675 1165 3705 1195
rect 4640 1160 4675 1195
rect 4890 1160 4925 1195
rect 5860 1165 5890 1195
<< metal1 >>
rect 3990 2680 5060 2750
rect 3990 2460 4160 2680
rect 4180 2460 4360 2680
rect 4380 2460 4560 2680
rect 4580 2460 4760 2680
rect 4780 2460 4955 2680
rect 4975 2460 5060 2680
rect 3990 2340 5060 2460
rect 3990 2270 4470 2340
rect 4490 2270 4600 2340
rect 4620 2270 4810 2340
rect 4830 2270 4940 2340
rect 4960 2270 5060 2340
rect 3990 2230 5060 2270
rect 3990 1960 5060 2015
rect 3990 1940 4110 1960
rect 4130 1940 4240 1960
rect 4260 1940 4810 1960
rect 4830 1940 4940 1960
rect 4960 1940 5060 1960
rect 3990 1880 5060 1940
rect 3990 1860 4175 1880
rect 4195 1860 5060 1880
rect 3990 1780 5060 1860
rect 3990 1560 4655 1780
rect 4675 1560 4855 1780
rect 4875 1560 5060 1780
rect 3990 1445 5060 1560
rect 3990 1425 4235 1445
rect 4255 1425 5060 1445
rect 3990 1385 5060 1425
rect 3665 1195 3715 1205
rect 3665 1165 3675 1195
rect 3705 1165 3715 1195
rect 3665 1155 3715 1165
rect 4630 1195 4685 1205
rect 4630 1160 4640 1195
rect 4675 1160 4685 1195
rect 4630 1150 4685 1160
rect 4880 1195 4935 1205
rect 4880 1160 4890 1195
rect 4925 1160 4935 1195
rect 4880 1150 4935 1160
rect 5850 1195 5900 1205
rect 5850 1165 5860 1195
rect 5890 1165 5900 1195
rect 5850 1155 5900 1165
<< via1 >>
rect 3675 1165 3705 1195
rect 4640 1160 4675 1195
rect 4890 1160 4925 1195
rect 5860 1165 5890 1195
<< metal2 >>
rect 3665 1195 3715 1205
rect 3665 1165 3675 1195
rect 3705 1165 3715 1195
rect 3665 1155 3715 1165
rect 4630 1195 4685 1205
rect 4630 1160 4640 1195
rect 4675 1160 4685 1195
rect 4630 1150 4685 1160
rect 4880 1195 4935 1205
rect 4880 1160 4890 1195
rect 4925 1160 4935 1195
rect 4880 1150 4935 1160
rect 5850 1195 5900 1205
rect 5850 1165 5860 1195
rect 5890 1165 5900 1195
rect 5850 1155 5900 1165
<< via2 >>
rect 3675 1165 3705 1195
rect 4640 1160 4675 1195
rect 4890 1160 4925 1195
rect 5860 1165 5890 1195
<< metal3 >>
rect 3665 1195 3715 1205
rect 3665 1165 3675 1195
rect 3705 1165 3715 1195
rect 3665 1155 3715 1165
rect 3670 1030 3715 1155
rect 4630 1195 4685 1205
rect 4630 1160 4640 1195
rect 4675 1160 4685 1195
rect 4630 1150 4685 1160
rect 4880 1195 4935 1205
rect 4880 1160 4890 1195
rect 4925 1160 4935 1195
rect 4880 1150 4935 1160
rect 5850 1195 5900 1205
rect 5850 1165 5860 1195
rect 5890 1165 5900 1195
rect 5850 1155 5900 1165
rect 5850 1030 5895 1155
rect 3670 0 4700 1030
rect 4865 0 5895 1030
<< via3 >>
rect 4640 1160 4675 1195
rect 4890 1160 4925 1195
<< mimcap >>
rect 3685 1005 4685 1015
rect 3685 970 4640 1005
rect 4675 970 4685 1005
rect 3685 15 4685 970
rect 4880 1005 5880 1015
rect 4880 970 4890 1005
rect 4925 970 5880 1005
rect 4880 15 5880 970
<< mimcapcontact >>
rect 4640 970 4675 1005
rect 4890 970 4925 1005
<< metal4 >>
rect 4630 1195 4685 1205
rect 4630 1160 4640 1195
rect 4675 1160 4685 1195
rect 4630 1005 4685 1160
rect 4630 970 4640 1005
rect 4675 970 4685 1005
rect 4630 965 4685 970
rect 4880 1195 4935 1205
rect 4880 1160 4890 1195
rect 4925 1160 4935 1195
rect 4880 1005 4935 1160
rect 4880 970 4890 1005
rect 4925 970 4935 1005
rect 4880 965 4935 970
<< labels >>
flabel locali 4775 1830 4775 1830 2 FreeSans 400 0 0 0 v_common_n
flabel locali 4680 2410 4680 2410 4 FreeSans 400 0 0 0 v_common_p
flabel locali 4490 2130 4490 2130 3 FreeSans 160 0 80 0 n_left
flabel locali 4620 2130 4620 2130 3 FreeSans 160 0 80 0 n_right
flabel locali 4260 2155 4260 2155 3 FreeSans 160 0 80 0 p_right
flabel locali 4055 2150 4055 2150 7 FreeSans 160 0 -80 0 p_left
flabel locali 4535 1510 4535 1510 5 FreeSans 160 0 0 -80 n_bias
flabel locali 3940 2610 3940 2610 7 FreeSans 160 0 -80 0 p_bias
<< end >>
