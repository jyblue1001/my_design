magic
tech sky130A
timestamp 1755893231
<< nwell >>
rect 16315 1155 16695 1295
rect 16825 1155 17315 1295
rect 17445 1155 18155 1295
rect 18285 1155 18775 1295
rect 16375 695 16760 835
rect 16910 595 18690 935
rect 18845 695 19170 935
rect 16360 15 17725 155
rect 17875 15 19240 155
<< pwell >>
rect 17780 -4320 17820 -4120
<< nmos >>
rect 17000 -480 17020 -230
rect 17060 -480 17080 -230
rect 18520 -480 18540 -230
rect 18580 -480 18600 -230
rect 16570 -1045 17070 -795
rect 17190 -1045 17690 -795
rect 17910 -1045 18410 -795
rect 18530 -1045 19030 -795
rect 16780 -1350 17780 -1250
rect 17820 -1350 18820 -1250
rect 16640 -1670 16655 -1570
rect 16695 -1670 16710 -1570
rect 16750 -1670 16765 -1570
rect 16805 -1670 16820 -1570
rect 16860 -1670 16875 -1570
rect 17065 -1670 17080 -1570
rect 17120 -1670 17135 -1570
rect 17175 -1670 17190 -1570
rect 17230 -1670 17245 -1570
rect 17285 -1670 17300 -1570
rect 17340 -1670 17355 -1570
rect 17395 -1670 17410 -1570
rect 17450 -1670 17465 -1570
rect 17655 -1670 17670 -1570
rect 17710 -1670 17725 -1570
rect 17765 -1670 17780 -1570
rect 17820 -1670 17835 -1570
rect 17875 -1670 17890 -1570
rect 17930 -1670 17945 -1570
rect 17985 -1670 18000 -1570
rect 18190 -1670 18205 -1570
rect 18245 -1670 18260 -1570
rect 18300 -1670 18315 -1570
rect 18355 -1670 18370 -1570
rect 18410 -1670 18425 -1570
rect 18465 -1670 18480 -1570
rect 18520 -1670 18535 -1570
rect 18575 -1670 18590 -1570
<< pmos >>
rect 16415 1175 16430 1275
rect 16470 1175 16485 1275
rect 16525 1175 16540 1275
rect 16580 1175 16595 1275
rect 16925 1175 16940 1275
rect 16980 1175 16995 1275
rect 17035 1175 17050 1275
rect 17090 1175 17105 1275
rect 17145 1175 17160 1275
rect 17200 1175 17215 1275
rect 17545 1175 17560 1275
rect 17600 1175 17615 1275
rect 17655 1175 17670 1275
rect 17710 1175 17725 1275
rect 17765 1175 17780 1275
rect 17820 1175 17835 1275
rect 17875 1175 17890 1275
rect 17930 1175 17945 1275
rect 17985 1175 18000 1275
rect 18040 1175 18055 1275
rect 18385 1175 18400 1275
rect 18440 1175 18455 1275
rect 18495 1175 18510 1275
rect 18550 1175 18565 1275
rect 18605 1175 18620 1275
rect 18660 1175 18675 1275
rect 16475 715 16490 815
rect 16530 715 16545 815
rect 16585 715 16600 815
rect 16640 715 16655 815
rect 17010 615 17060 915
rect 17100 615 17150 915
rect 17190 615 17240 915
rect 17280 615 17330 915
rect 17370 615 17420 915
rect 17460 615 17510 915
rect 17550 615 17600 915
rect 17640 615 17690 915
rect 17730 615 17780 915
rect 17820 615 17870 915
rect 17910 615 17960 915
rect 18000 615 18050 915
rect 18090 615 18140 915
rect 18180 615 18230 915
rect 18270 615 18320 915
rect 18360 615 18410 915
rect 18450 615 18500 915
rect 18540 615 18590 915
rect 18945 715 18960 915
rect 19000 715 19015 915
rect 19055 715 19070 915
rect 16460 35 16480 135
rect 16520 35 16540 135
rect 16580 35 16600 135
rect 16640 35 16660 135
rect 16700 35 16720 135
rect 16760 35 16780 135
rect 16820 35 16840 135
rect 16880 35 16900 135
rect 16940 35 16960 135
rect 17000 35 17020 135
rect 17060 35 17080 135
rect 17120 35 17140 135
rect 17180 35 17200 135
rect 17240 35 17260 135
rect 17300 35 17320 135
rect 17360 35 17380 135
rect 17420 35 17440 135
rect 17480 35 17500 135
rect 17540 35 17560 135
rect 17600 35 17620 135
rect 17980 35 18000 135
rect 18040 35 18060 135
rect 18100 35 18120 135
rect 18160 35 18180 135
rect 18220 35 18240 135
rect 18280 35 18300 135
rect 18340 35 18360 135
rect 18400 35 18420 135
rect 18460 35 18480 135
rect 18520 35 18540 135
rect 18580 35 18600 135
rect 18640 35 18660 135
rect 18700 35 18720 135
rect 18760 35 18780 135
rect 18820 35 18840 135
rect 18880 35 18900 135
rect 18940 35 18960 135
rect 19000 35 19020 135
rect 19060 35 19080 135
rect 19120 35 19140 135
<< ndiff >>
rect 16960 -245 17000 -230
rect 16960 -265 16970 -245
rect 16990 -265 17000 -245
rect 16960 -295 17000 -265
rect 16960 -315 16970 -295
rect 16990 -315 17000 -295
rect 16960 -345 17000 -315
rect 16960 -365 16970 -345
rect 16990 -365 17000 -345
rect 16960 -395 17000 -365
rect 16960 -415 16970 -395
rect 16990 -415 17000 -395
rect 16960 -445 17000 -415
rect 16960 -465 16970 -445
rect 16990 -465 17000 -445
rect 16960 -480 17000 -465
rect 17020 -245 17060 -230
rect 17020 -265 17030 -245
rect 17050 -265 17060 -245
rect 17020 -295 17060 -265
rect 17020 -315 17030 -295
rect 17050 -315 17060 -295
rect 17020 -345 17060 -315
rect 17020 -365 17030 -345
rect 17050 -365 17060 -345
rect 17020 -395 17060 -365
rect 17020 -415 17030 -395
rect 17050 -415 17060 -395
rect 17020 -445 17060 -415
rect 17020 -465 17030 -445
rect 17050 -465 17060 -445
rect 17020 -480 17060 -465
rect 17080 -245 17120 -230
rect 17080 -265 17090 -245
rect 17110 -265 17120 -245
rect 17080 -295 17120 -265
rect 17080 -315 17090 -295
rect 17110 -315 17120 -295
rect 17080 -345 17120 -315
rect 17080 -365 17090 -345
rect 17110 -365 17120 -345
rect 18480 -245 18520 -230
rect 18480 -265 18490 -245
rect 18510 -265 18520 -245
rect 18480 -295 18520 -265
rect 18480 -315 18490 -295
rect 18510 -315 18520 -295
rect 18480 -345 18520 -315
rect 17080 -395 17120 -365
rect 17080 -415 17090 -395
rect 17110 -415 17120 -395
rect 17080 -445 17120 -415
rect 17080 -465 17090 -445
rect 17110 -465 17120 -445
rect 17080 -480 17120 -465
rect 18480 -365 18490 -345
rect 18510 -365 18520 -345
rect 18480 -395 18520 -365
rect 18480 -415 18490 -395
rect 18510 -415 18520 -395
rect 18480 -445 18520 -415
rect 18480 -465 18490 -445
rect 18510 -465 18520 -445
rect 18480 -480 18520 -465
rect 18540 -245 18580 -230
rect 18540 -265 18550 -245
rect 18570 -265 18580 -245
rect 18540 -295 18580 -265
rect 18540 -315 18550 -295
rect 18570 -315 18580 -295
rect 18540 -345 18580 -315
rect 18540 -365 18550 -345
rect 18570 -365 18580 -345
rect 18540 -395 18580 -365
rect 18540 -415 18550 -395
rect 18570 -415 18580 -395
rect 18540 -445 18580 -415
rect 18540 -465 18550 -445
rect 18570 -465 18580 -445
rect 18540 -480 18580 -465
rect 18600 -245 18640 -230
rect 18600 -265 18610 -245
rect 18630 -265 18640 -245
rect 18600 -295 18640 -265
rect 18600 -315 18610 -295
rect 18630 -315 18640 -295
rect 18600 -345 18640 -315
rect 18600 -365 18610 -345
rect 18630 -365 18640 -345
rect 18600 -395 18640 -365
rect 18600 -415 18610 -395
rect 18630 -415 18640 -395
rect 18600 -445 18640 -415
rect 18600 -465 18610 -445
rect 18630 -465 18640 -445
rect 18600 -480 18640 -465
rect 16530 -810 16570 -795
rect 16530 -830 16540 -810
rect 16560 -830 16570 -810
rect 16530 -860 16570 -830
rect 16530 -880 16540 -860
rect 16560 -880 16570 -860
rect 16530 -910 16570 -880
rect 16530 -930 16540 -910
rect 16560 -930 16570 -910
rect 16530 -960 16570 -930
rect 16530 -980 16540 -960
rect 16560 -980 16570 -960
rect 16530 -1010 16570 -980
rect 16530 -1030 16540 -1010
rect 16560 -1030 16570 -1010
rect 16530 -1045 16570 -1030
rect 17070 -810 17110 -795
rect 17150 -810 17190 -795
rect 17070 -830 17080 -810
rect 17100 -830 17110 -810
rect 17150 -830 17160 -810
rect 17180 -830 17190 -810
rect 17070 -860 17110 -830
rect 17150 -860 17190 -830
rect 17070 -880 17080 -860
rect 17100 -880 17110 -860
rect 17150 -880 17160 -860
rect 17180 -880 17190 -860
rect 17070 -910 17110 -880
rect 17150 -910 17190 -880
rect 17070 -930 17080 -910
rect 17100 -930 17110 -910
rect 17150 -930 17160 -910
rect 17180 -930 17190 -910
rect 17070 -960 17110 -930
rect 17150 -960 17190 -930
rect 17070 -980 17080 -960
rect 17100 -980 17110 -960
rect 17150 -980 17160 -960
rect 17180 -980 17190 -960
rect 17070 -1010 17110 -980
rect 17150 -1010 17190 -980
rect 17070 -1030 17080 -1010
rect 17100 -1030 17110 -1010
rect 17150 -1030 17160 -1010
rect 17180 -1030 17190 -1010
rect 17070 -1040 17110 -1030
rect 17150 -1040 17190 -1030
rect 17070 -1045 17190 -1040
rect 17690 -810 17730 -795
rect 17690 -830 17700 -810
rect 17720 -830 17730 -810
rect 17690 -860 17730 -830
rect 17690 -880 17700 -860
rect 17720 -880 17730 -860
rect 17690 -910 17730 -880
rect 17690 -930 17700 -910
rect 17720 -930 17730 -910
rect 17690 -960 17730 -930
rect 17690 -980 17700 -960
rect 17720 -980 17730 -960
rect 17690 -1010 17730 -980
rect 17690 -1030 17700 -1010
rect 17720 -1030 17730 -1010
rect 17690 -1045 17730 -1030
rect 17870 -810 17910 -795
rect 17870 -830 17880 -810
rect 17900 -830 17910 -810
rect 17870 -860 17910 -830
rect 17870 -880 17880 -860
rect 17900 -880 17910 -860
rect 17870 -910 17910 -880
rect 17870 -930 17880 -910
rect 17900 -930 17910 -910
rect 17870 -960 17910 -930
rect 17870 -980 17880 -960
rect 17900 -980 17910 -960
rect 17870 -1010 17910 -980
rect 17870 -1030 17880 -1010
rect 17900 -1030 17910 -1010
rect 17870 -1045 17910 -1030
rect 18410 -810 18450 -795
rect 18490 -810 18530 -795
rect 18410 -830 18420 -810
rect 18440 -830 18450 -810
rect 18490 -830 18500 -810
rect 18520 -830 18530 -810
rect 18410 -860 18450 -830
rect 18490 -860 18530 -830
rect 18410 -880 18420 -860
rect 18440 -880 18450 -860
rect 18490 -880 18500 -860
rect 18520 -880 18530 -860
rect 18410 -910 18450 -880
rect 18490 -910 18530 -880
rect 18410 -930 18420 -910
rect 18440 -930 18450 -910
rect 18490 -930 18500 -910
rect 18520 -930 18530 -910
rect 18410 -960 18450 -930
rect 18490 -960 18530 -930
rect 18410 -980 18420 -960
rect 18440 -980 18450 -960
rect 18490 -980 18500 -960
rect 18520 -980 18530 -960
rect 18410 -1010 18450 -980
rect 18490 -1010 18530 -980
rect 18410 -1030 18420 -1010
rect 18440 -1030 18450 -1010
rect 18490 -1030 18500 -1010
rect 18520 -1030 18530 -1010
rect 18410 -1045 18450 -1030
rect 18490 -1045 18530 -1030
rect 19030 -810 19070 -795
rect 19030 -830 19040 -810
rect 19060 -830 19070 -810
rect 19030 -860 19070 -830
rect 19030 -880 19040 -860
rect 19060 -880 19070 -860
rect 19030 -910 19070 -880
rect 19030 -930 19040 -910
rect 19060 -930 19070 -910
rect 19030 -960 19070 -930
rect 19030 -980 19040 -960
rect 19060 -980 19070 -960
rect 19030 -1010 19070 -980
rect 19030 -1030 19040 -1010
rect 19060 -1030 19070 -1010
rect 19030 -1045 19070 -1030
rect 16740 -1265 16780 -1250
rect 16740 -1285 16750 -1265
rect 16770 -1285 16780 -1265
rect 16740 -1315 16780 -1285
rect 16740 -1335 16750 -1315
rect 16770 -1335 16780 -1315
rect 16740 -1350 16780 -1335
rect 17780 -1265 17820 -1250
rect 17780 -1285 17790 -1265
rect 17810 -1285 17820 -1265
rect 17780 -1315 17820 -1285
rect 17780 -1335 17790 -1315
rect 17810 -1335 17820 -1315
rect 17780 -1350 17820 -1335
rect 18820 -1265 18860 -1250
rect 18820 -1285 18830 -1265
rect 18850 -1285 18860 -1265
rect 18820 -1315 18860 -1285
rect 18820 -1335 18830 -1315
rect 18850 -1335 18860 -1315
rect 18820 -1350 18860 -1335
rect 16600 -1585 16640 -1570
rect 16600 -1605 16610 -1585
rect 16630 -1605 16640 -1585
rect 16600 -1635 16640 -1605
rect 16600 -1655 16610 -1635
rect 16630 -1655 16640 -1635
rect 16600 -1670 16640 -1655
rect 16655 -1585 16695 -1570
rect 16655 -1605 16665 -1585
rect 16685 -1605 16695 -1585
rect 16655 -1635 16695 -1605
rect 16655 -1655 16665 -1635
rect 16685 -1655 16695 -1635
rect 16655 -1670 16695 -1655
rect 16710 -1585 16750 -1570
rect 16710 -1605 16720 -1585
rect 16740 -1605 16750 -1585
rect 16710 -1635 16750 -1605
rect 16710 -1655 16720 -1635
rect 16740 -1655 16750 -1635
rect 16710 -1670 16750 -1655
rect 16765 -1585 16805 -1570
rect 16765 -1605 16775 -1585
rect 16795 -1605 16805 -1585
rect 16765 -1635 16805 -1605
rect 16765 -1655 16775 -1635
rect 16795 -1655 16805 -1635
rect 16765 -1670 16805 -1655
rect 16820 -1585 16860 -1570
rect 16820 -1605 16830 -1585
rect 16850 -1605 16860 -1585
rect 16820 -1635 16860 -1605
rect 16820 -1655 16830 -1635
rect 16850 -1655 16860 -1635
rect 16820 -1670 16860 -1655
rect 16875 -1585 16915 -1570
rect 16875 -1605 16885 -1585
rect 16905 -1605 16915 -1585
rect 16875 -1635 16915 -1605
rect 16875 -1655 16885 -1635
rect 16905 -1655 16915 -1635
rect 16875 -1670 16915 -1655
rect 17025 -1585 17065 -1570
rect 17025 -1605 17035 -1585
rect 17055 -1605 17065 -1585
rect 17025 -1635 17065 -1605
rect 17025 -1655 17035 -1635
rect 17055 -1655 17065 -1635
rect 17025 -1670 17065 -1655
rect 17080 -1585 17120 -1570
rect 17080 -1605 17090 -1585
rect 17110 -1605 17120 -1585
rect 17080 -1635 17120 -1605
rect 17080 -1655 17090 -1635
rect 17110 -1655 17120 -1635
rect 17080 -1670 17120 -1655
rect 17135 -1585 17175 -1570
rect 17135 -1605 17145 -1585
rect 17165 -1605 17175 -1585
rect 17135 -1635 17175 -1605
rect 17135 -1655 17145 -1635
rect 17165 -1655 17175 -1635
rect 17135 -1670 17175 -1655
rect 17190 -1585 17230 -1570
rect 17190 -1605 17200 -1585
rect 17220 -1605 17230 -1585
rect 17190 -1635 17230 -1605
rect 17190 -1655 17200 -1635
rect 17220 -1655 17230 -1635
rect 17190 -1670 17230 -1655
rect 17245 -1585 17285 -1570
rect 17245 -1605 17255 -1585
rect 17275 -1605 17285 -1585
rect 17245 -1635 17285 -1605
rect 17245 -1655 17255 -1635
rect 17275 -1655 17285 -1635
rect 17245 -1670 17285 -1655
rect 17300 -1585 17340 -1570
rect 17300 -1605 17310 -1585
rect 17330 -1605 17340 -1585
rect 17300 -1635 17340 -1605
rect 17300 -1655 17310 -1635
rect 17330 -1655 17340 -1635
rect 17300 -1670 17340 -1655
rect 17355 -1585 17395 -1570
rect 17355 -1605 17365 -1585
rect 17385 -1605 17395 -1585
rect 17355 -1635 17395 -1605
rect 17355 -1655 17365 -1635
rect 17385 -1655 17395 -1635
rect 17355 -1670 17395 -1655
rect 17410 -1585 17450 -1570
rect 17410 -1605 17420 -1585
rect 17440 -1605 17450 -1585
rect 17410 -1635 17450 -1605
rect 17410 -1655 17420 -1635
rect 17440 -1655 17450 -1635
rect 17410 -1670 17450 -1655
rect 17465 -1585 17505 -1570
rect 17465 -1605 17475 -1585
rect 17495 -1605 17505 -1585
rect 17465 -1635 17505 -1605
rect 17465 -1655 17475 -1635
rect 17495 -1655 17505 -1635
rect 17465 -1670 17505 -1655
rect 17615 -1585 17655 -1570
rect 17615 -1605 17625 -1585
rect 17645 -1605 17655 -1585
rect 17615 -1635 17655 -1605
rect 17615 -1655 17625 -1635
rect 17645 -1655 17655 -1635
rect 17615 -1670 17655 -1655
rect 17670 -1585 17710 -1570
rect 17670 -1605 17680 -1585
rect 17700 -1605 17710 -1585
rect 17670 -1635 17710 -1605
rect 17670 -1655 17680 -1635
rect 17700 -1655 17710 -1635
rect 17670 -1670 17710 -1655
rect 17725 -1585 17765 -1570
rect 17725 -1605 17735 -1585
rect 17755 -1605 17765 -1585
rect 17725 -1635 17765 -1605
rect 17725 -1655 17735 -1635
rect 17755 -1655 17765 -1635
rect 17725 -1670 17765 -1655
rect 17780 -1585 17820 -1570
rect 17780 -1605 17790 -1585
rect 17810 -1605 17820 -1585
rect 17780 -1635 17820 -1605
rect 17780 -1655 17790 -1635
rect 17810 -1655 17820 -1635
rect 17780 -1670 17820 -1655
rect 17835 -1585 17875 -1570
rect 17835 -1605 17845 -1585
rect 17865 -1605 17875 -1585
rect 17835 -1635 17875 -1605
rect 17835 -1655 17845 -1635
rect 17865 -1655 17875 -1635
rect 17835 -1670 17875 -1655
rect 17890 -1585 17930 -1570
rect 17890 -1605 17900 -1585
rect 17920 -1605 17930 -1585
rect 17890 -1635 17930 -1605
rect 17890 -1655 17900 -1635
rect 17920 -1655 17930 -1635
rect 17890 -1670 17930 -1655
rect 17945 -1585 17985 -1570
rect 17945 -1605 17955 -1585
rect 17975 -1605 17985 -1585
rect 17945 -1635 17985 -1605
rect 17945 -1655 17955 -1635
rect 17975 -1655 17985 -1635
rect 17945 -1670 17985 -1655
rect 18000 -1585 18040 -1570
rect 18000 -1605 18010 -1585
rect 18030 -1605 18040 -1585
rect 18000 -1635 18040 -1605
rect 18000 -1655 18010 -1635
rect 18030 -1655 18040 -1635
rect 18000 -1670 18040 -1655
rect 18150 -1585 18190 -1570
rect 18150 -1605 18160 -1585
rect 18180 -1605 18190 -1585
rect 18150 -1635 18190 -1605
rect 18150 -1655 18160 -1635
rect 18180 -1655 18190 -1635
rect 18150 -1670 18190 -1655
rect 18205 -1585 18245 -1570
rect 18205 -1605 18215 -1585
rect 18235 -1605 18245 -1585
rect 18205 -1635 18245 -1605
rect 18205 -1655 18215 -1635
rect 18235 -1655 18245 -1635
rect 18205 -1670 18245 -1655
rect 18260 -1585 18300 -1570
rect 18260 -1605 18270 -1585
rect 18290 -1605 18300 -1585
rect 18260 -1635 18300 -1605
rect 18260 -1655 18270 -1635
rect 18290 -1655 18300 -1635
rect 18260 -1670 18300 -1655
rect 18315 -1585 18355 -1570
rect 18315 -1605 18325 -1585
rect 18345 -1605 18355 -1585
rect 18315 -1635 18355 -1605
rect 18315 -1655 18325 -1635
rect 18345 -1655 18355 -1635
rect 18315 -1670 18355 -1655
rect 18370 -1585 18410 -1570
rect 18370 -1605 18380 -1585
rect 18400 -1605 18410 -1585
rect 18370 -1635 18410 -1605
rect 18370 -1655 18380 -1635
rect 18400 -1655 18410 -1635
rect 18370 -1670 18410 -1655
rect 18425 -1585 18465 -1570
rect 18425 -1605 18435 -1585
rect 18455 -1605 18465 -1585
rect 18425 -1635 18465 -1605
rect 18425 -1655 18435 -1635
rect 18455 -1655 18465 -1635
rect 18425 -1670 18465 -1655
rect 18480 -1585 18520 -1570
rect 18480 -1605 18490 -1585
rect 18510 -1605 18520 -1585
rect 18480 -1635 18520 -1605
rect 18480 -1655 18490 -1635
rect 18510 -1655 18520 -1635
rect 18480 -1670 18520 -1655
rect 18535 -1585 18575 -1570
rect 18535 -1605 18545 -1585
rect 18565 -1605 18575 -1585
rect 18535 -1635 18575 -1605
rect 18535 -1655 18545 -1635
rect 18565 -1655 18575 -1635
rect 18535 -1670 18575 -1655
rect 18590 -1585 18630 -1570
rect 18590 -1605 18600 -1585
rect 18620 -1605 18630 -1585
rect 18590 -1635 18630 -1605
rect 18590 -1655 18600 -1635
rect 18620 -1655 18630 -1635
rect 18590 -1670 18630 -1655
<< pdiff >>
rect 16375 1260 16415 1275
rect 16375 1240 16385 1260
rect 16405 1240 16415 1260
rect 16375 1210 16415 1240
rect 16375 1190 16385 1210
rect 16405 1190 16415 1210
rect 16375 1175 16415 1190
rect 16430 1260 16470 1275
rect 16430 1240 16440 1260
rect 16460 1240 16470 1260
rect 16430 1210 16470 1240
rect 16430 1190 16440 1210
rect 16460 1190 16470 1210
rect 16430 1175 16470 1190
rect 16485 1260 16525 1275
rect 16485 1240 16495 1260
rect 16515 1240 16525 1260
rect 16485 1210 16525 1240
rect 16485 1190 16495 1210
rect 16515 1190 16525 1210
rect 16485 1175 16525 1190
rect 16540 1260 16580 1275
rect 16540 1240 16550 1260
rect 16570 1240 16580 1260
rect 16540 1210 16580 1240
rect 16540 1190 16550 1210
rect 16570 1190 16580 1210
rect 16540 1175 16580 1190
rect 16595 1260 16635 1275
rect 16595 1240 16605 1260
rect 16625 1240 16635 1260
rect 16595 1210 16635 1240
rect 16595 1190 16605 1210
rect 16625 1190 16635 1210
rect 16595 1175 16635 1190
rect 16885 1260 16925 1275
rect 16885 1188 16895 1260
rect 16915 1188 16925 1260
rect 16885 1175 16925 1188
rect 16940 1260 16980 1275
rect 16940 1188 16950 1260
rect 16970 1188 16980 1260
rect 16940 1175 16980 1188
rect 16995 1260 17035 1275
rect 16995 1188 17005 1260
rect 17025 1188 17035 1260
rect 16995 1175 17035 1188
rect 17050 1260 17090 1275
rect 17050 1188 17060 1260
rect 17080 1188 17090 1260
rect 17050 1175 17090 1188
rect 17105 1260 17145 1275
rect 17105 1188 17115 1260
rect 17135 1188 17145 1260
rect 17105 1175 17145 1188
rect 17160 1260 17200 1275
rect 17160 1188 17170 1260
rect 17190 1188 17200 1260
rect 17160 1175 17200 1188
rect 17215 1260 17255 1275
rect 17215 1188 17225 1260
rect 17245 1188 17255 1260
rect 17215 1175 17255 1188
rect 17505 1260 17545 1275
rect 17505 1240 17515 1260
rect 17535 1240 17545 1260
rect 17505 1210 17545 1240
rect 17505 1190 17515 1210
rect 17535 1190 17545 1210
rect 17505 1175 17545 1190
rect 17560 1260 17600 1275
rect 17560 1240 17570 1260
rect 17590 1240 17600 1260
rect 17560 1210 17600 1240
rect 17560 1190 17570 1210
rect 17590 1190 17600 1210
rect 17560 1175 17600 1190
rect 17615 1260 17655 1275
rect 17615 1240 17625 1260
rect 17645 1240 17655 1260
rect 17615 1210 17655 1240
rect 17615 1190 17625 1210
rect 17645 1190 17655 1210
rect 17615 1175 17655 1190
rect 17670 1260 17710 1275
rect 17670 1240 17680 1260
rect 17700 1240 17710 1260
rect 17670 1210 17710 1240
rect 17670 1190 17680 1210
rect 17700 1190 17710 1210
rect 17670 1175 17710 1190
rect 17725 1260 17765 1275
rect 17725 1240 17735 1260
rect 17755 1240 17765 1260
rect 17725 1210 17765 1240
rect 17725 1190 17735 1210
rect 17755 1190 17765 1210
rect 17725 1175 17765 1190
rect 17780 1260 17820 1275
rect 17780 1240 17790 1260
rect 17810 1240 17820 1260
rect 17780 1210 17820 1240
rect 17780 1190 17790 1210
rect 17810 1190 17820 1210
rect 17780 1175 17820 1190
rect 17835 1260 17875 1275
rect 17835 1240 17845 1260
rect 17865 1240 17875 1260
rect 17835 1210 17875 1240
rect 17835 1190 17845 1210
rect 17865 1190 17875 1210
rect 17835 1175 17875 1190
rect 17890 1260 17930 1275
rect 17890 1240 17900 1260
rect 17920 1240 17930 1260
rect 17890 1210 17930 1240
rect 17890 1190 17900 1210
rect 17920 1190 17930 1210
rect 17890 1175 17930 1190
rect 17945 1260 17985 1275
rect 17945 1240 17955 1260
rect 17975 1240 17985 1260
rect 17945 1210 17985 1240
rect 17945 1190 17955 1210
rect 17975 1190 17985 1210
rect 17945 1175 17985 1190
rect 18000 1260 18040 1275
rect 18000 1240 18010 1260
rect 18030 1240 18040 1260
rect 18000 1210 18040 1240
rect 18000 1190 18010 1210
rect 18030 1190 18040 1210
rect 18000 1175 18040 1190
rect 18055 1260 18095 1275
rect 18055 1240 18065 1260
rect 18085 1240 18095 1260
rect 18055 1210 18095 1240
rect 18055 1190 18065 1210
rect 18085 1190 18095 1210
rect 18055 1175 18095 1190
rect 18345 1260 18385 1275
rect 18345 1190 18355 1260
rect 18375 1190 18385 1260
rect 18345 1175 18385 1190
rect 18400 1260 18440 1275
rect 18400 1190 18410 1260
rect 18430 1190 18440 1260
rect 18400 1175 18440 1190
rect 18455 1260 18495 1275
rect 18455 1190 18465 1260
rect 18485 1190 18495 1260
rect 18455 1175 18495 1190
rect 18510 1260 18550 1275
rect 18510 1190 18520 1260
rect 18540 1190 18550 1260
rect 18510 1175 18550 1190
rect 18565 1260 18605 1275
rect 18565 1190 18575 1260
rect 18595 1190 18605 1260
rect 18565 1175 18605 1190
rect 18620 1260 18660 1275
rect 18620 1190 18630 1260
rect 18650 1190 18660 1260
rect 18620 1175 18660 1190
rect 18675 1260 18715 1275
rect 18675 1190 18685 1260
rect 18705 1190 18715 1260
rect 18675 1175 18715 1190
rect 16970 900 17010 915
rect 16970 880 16980 900
rect 17000 880 17010 900
rect 16970 850 17010 880
rect 16970 830 16980 850
rect 17000 830 17010 850
rect 16435 800 16475 815
rect 16435 780 16445 800
rect 16465 780 16475 800
rect 16435 750 16475 780
rect 16435 730 16445 750
rect 16465 730 16475 750
rect 16435 715 16475 730
rect 16490 800 16530 815
rect 16490 780 16500 800
rect 16520 780 16530 800
rect 16490 750 16530 780
rect 16490 730 16500 750
rect 16520 730 16530 750
rect 16490 715 16530 730
rect 16545 800 16585 815
rect 16545 780 16555 800
rect 16575 780 16585 800
rect 16545 750 16585 780
rect 16545 730 16555 750
rect 16575 730 16585 750
rect 16545 715 16585 730
rect 16600 800 16640 815
rect 16600 780 16610 800
rect 16630 780 16640 800
rect 16600 750 16640 780
rect 16600 730 16610 750
rect 16630 730 16640 750
rect 16600 715 16640 730
rect 16655 800 16700 815
rect 16655 780 16665 800
rect 16685 780 16700 800
rect 16655 750 16700 780
rect 16655 730 16665 750
rect 16685 730 16700 750
rect 16655 715 16700 730
rect 16970 800 17010 830
rect 16970 780 16980 800
rect 17000 780 17010 800
rect 16970 750 17010 780
rect 16970 730 16980 750
rect 17000 730 17010 750
rect 16970 700 17010 730
rect 16970 680 16980 700
rect 17000 680 17010 700
rect 16970 650 17010 680
rect 16970 630 16980 650
rect 17000 630 17010 650
rect 16970 615 17010 630
rect 17060 900 17100 915
rect 17060 880 17070 900
rect 17090 880 17100 900
rect 17060 850 17100 880
rect 17060 830 17070 850
rect 17090 830 17100 850
rect 17060 800 17100 830
rect 17060 780 17070 800
rect 17090 780 17100 800
rect 17060 750 17100 780
rect 17060 730 17070 750
rect 17090 730 17100 750
rect 17060 700 17100 730
rect 17060 680 17070 700
rect 17090 680 17100 700
rect 17060 650 17100 680
rect 17060 630 17070 650
rect 17090 630 17100 650
rect 17060 615 17100 630
rect 17150 900 17190 915
rect 17150 880 17160 900
rect 17180 880 17190 900
rect 17150 850 17190 880
rect 17150 830 17160 850
rect 17180 830 17190 850
rect 17150 800 17190 830
rect 17150 780 17160 800
rect 17180 780 17190 800
rect 17150 750 17190 780
rect 17150 730 17160 750
rect 17180 730 17190 750
rect 17150 700 17190 730
rect 17150 680 17160 700
rect 17180 680 17190 700
rect 17150 650 17190 680
rect 17150 630 17160 650
rect 17180 630 17190 650
rect 17150 615 17190 630
rect 17240 900 17280 915
rect 17240 880 17250 900
rect 17270 880 17280 900
rect 17240 850 17280 880
rect 17240 830 17250 850
rect 17270 830 17280 850
rect 17240 800 17280 830
rect 17240 780 17250 800
rect 17270 780 17280 800
rect 17240 750 17280 780
rect 17240 730 17250 750
rect 17270 730 17280 750
rect 17240 700 17280 730
rect 17240 680 17250 700
rect 17270 680 17280 700
rect 17240 650 17280 680
rect 17240 630 17250 650
rect 17270 630 17280 650
rect 17240 615 17280 630
rect 17330 900 17370 915
rect 17330 880 17340 900
rect 17360 880 17370 900
rect 17330 850 17370 880
rect 17330 830 17340 850
rect 17360 830 17370 850
rect 17330 800 17370 830
rect 17330 780 17340 800
rect 17360 780 17370 800
rect 17330 750 17370 780
rect 17330 730 17340 750
rect 17360 730 17370 750
rect 17330 700 17370 730
rect 17330 680 17340 700
rect 17360 680 17370 700
rect 17330 650 17370 680
rect 17330 630 17340 650
rect 17360 630 17370 650
rect 17330 615 17370 630
rect 17420 900 17460 915
rect 17420 880 17430 900
rect 17450 880 17460 900
rect 17420 850 17460 880
rect 17420 830 17430 850
rect 17450 830 17460 850
rect 17420 800 17460 830
rect 17420 780 17430 800
rect 17450 780 17460 800
rect 17420 750 17460 780
rect 17420 730 17430 750
rect 17450 730 17460 750
rect 17420 700 17460 730
rect 17420 680 17430 700
rect 17450 680 17460 700
rect 17420 650 17460 680
rect 17420 630 17430 650
rect 17450 630 17460 650
rect 17420 615 17460 630
rect 17510 900 17550 915
rect 17510 880 17520 900
rect 17540 880 17550 900
rect 17510 850 17550 880
rect 17510 830 17520 850
rect 17540 830 17550 850
rect 17510 800 17550 830
rect 17510 780 17520 800
rect 17540 780 17550 800
rect 17510 750 17550 780
rect 17510 730 17520 750
rect 17540 730 17550 750
rect 17510 700 17550 730
rect 17510 680 17520 700
rect 17540 680 17550 700
rect 17510 650 17550 680
rect 17510 630 17520 650
rect 17540 630 17550 650
rect 17510 615 17550 630
rect 17600 900 17640 915
rect 17600 880 17610 900
rect 17630 880 17640 900
rect 17600 850 17640 880
rect 17600 830 17610 850
rect 17630 830 17640 850
rect 17600 800 17640 830
rect 17600 780 17610 800
rect 17630 780 17640 800
rect 17600 750 17640 780
rect 17600 730 17610 750
rect 17630 730 17640 750
rect 17600 700 17640 730
rect 17600 680 17610 700
rect 17630 680 17640 700
rect 17600 650 17640 680
rect 17600 630 17610 650
rect 17630 630 17640 650
rect 17600 615 17640 630
rect 17690 900 17730 915
rect 17690 880 17700 900
rect 17720 880 17730 900
rect 17690 850 17730 880
rect 17690 830 17700 850
rect 17720 830 17730 850
rect 17690 800 17730 830
rect 17690 780 17700 800
rect 17720 780 17730 800
rect 17690 750 17730 780
rect 17690 730 17700 750
rect 17720 730 17730 750
rect 17690 700 17730 730
rect 17690 680 17700 700
rect 17720 680 17730 700
rect 17690 650 17730 680
rect 17690 630 17700 650
rect 17720 630 17730 650
rect 17690 615 17730 630
rect 17780 900 17820 915
rect 17780 880 17790 900
rect 17810 880 17820 900
rect 17780 850 17820 880
rect 17780 830 17790 850
rect 17810 830 17820 850
rect 17780 800 17820 830
rect 17780 780 17790 800
rect 17810 780 17820 800
rect 17780 750 17820 780
rect 17780 730 17790 750
rect 17810 730 17820 750
rect 17780 700 17820 730
rect 17780 680 17790 700
rect 17810 680 17820 700
rect 17780 650 17820 680
rect 17780 630 17790 650
rect 17810 630 17820 650
rect 17780 615 17820 630
rect 17870 900 17910 915
rect 17870 880 17880 900
rect 17900 880 17910 900
rect 17870 850 17910 880
rect 17870 830 17880 850
rect 17900 830 17910 850
rect 17870 800 17910 830
rect 17870 780 17880 800
rect 17900 780 17910 800
rect 17870 750 17910 780
rect 17870 730 17880 750
rect 17900 730 17910 750
rect 17870 700 17910 730
rect 17870 680 17880 700
rect 17900 680 17910 700
rect 17870 650 17910 680
rect 17870 630 17880 650
rect 17900 630 17910 650
rect 17870 615 17910 630
rect 17960 900 18000 915
rect 17960 880 17970 900
rect 17990 880 18000 900
rect 17960 850 18000 880
rect 17960 830 17970 850
rect 17990 830 18000 850
rect 17960 800 18000 830
rect 17960 780 17970 800
rect 17990 780 18000 800
rect 17960 750 18000 780
rect 17960 730 17970 750
rect 17990 730 18000 750
rect 17960 700 18000 730
rect 17960 680 17970 700
rect 17990 680 18000 700
rect 17960 650 18000 680
rect 17960 630 17970 650
rect 17990 630 18000 650
rect 17960 615 18000 630
rect 18050 900 18090 915
rect 18050 880 18060 900
rect 18080 880 18090 900
rect 18050 850 18090 880
rect 18050 830 18060 850
rect 18080 830 18090 850
rect 18050 800 18090 830
rect 18050 780 18060 800
rect 18080 780 18090 800
rect 18050 750 18090 780
rect 18050 730 18060 750
rect 18080 730 18090 750
rect 18050 700 18090 730
rect 18050 680 18060 700
rect 18080 680 18090 700
rect 18050 650 18090 680
rect 18050 630 18060 650
rect 18080 630 18090 650
rect 18050 615 18090 630
rect 18140 900 18180 915
rect 18140 880 18150 900
rect 18170 880 18180 900
rect 18140 850 18180 880
rect 18140 830 18150 850
rect 18170 830 18180 850
rect 18140 800 18180 830
rect 18140 780 18150 800
rect 18170 780 18180 800
rect 18140 750 18180 780
rect 18140 730 18150 750
rect 18170 730 18180 750
rect 18140 700 18180 730
rect 18140 680 18150 700
rect 18170 680 18180 700
rect 18140 650 18180 680
rect 18140 630 18150 650
rect 18170 630 18180 650
rect 18140 615 18180 630
rect 18230 900 18270 915
rect 18230 880 18240 900
rect 18260 880 18270 900
rect 18230 850 18270 880
rect 18230 830 18240 850
rect 18260 830 18270 850
rect 18230 800 18270 830
rect 18230 780 18240 800
rect 18260 780 18270 800
rect 18230 750 18270 780
rect 18230 730 18240 750
rect 18260 730 18270 750
rect 18230 700 18270 730
rect 18230 680 18240 700
rect 18260 680 18270 700
rect 18230 650 18270 680
rect 18230 630 18240 650
rect 18260 630 18270 650
rect 18230 615 18270 630
rect 18320 900 18360 915
rect 18320 880 18330 900
rect 18350 880 18360 900
rect 18320 850 18360 880
rect 18320 830 18330 850
rect 18350 830 18360 850
rect 18320 800 18360 830
rect 18320 780 18330 800
rect 18350 780 18360 800
rect 18320 750 18360 780
rect 18320 730 18330 750
rect 18350 730 18360 750
rect 18320 700 18360 730
rect 18320 680 18330 700
rect 18350 680 18360 700
rect 18320 650 18360 680
rect 18320 630 18330 650
rect 18350 630 18360 650
rect 18320 615 18360 630
rect 18410 900 18450 915
rect 18410 880 18420 900
rect 18440 880 18450 900
rect 18410 850 18450 880
rect 18410 830 18420 850
rect 18440 830 18450 850
rect 18410 800 18450 830
rect 18410 780 18420 800
rect 18440 780 18450 800
rect 18410 750 18450 780
rect 18410 730 18420 750
rect 18440 730 18450 750
rect 18410 700 18450 730
rect 18410 680 18420 700
rect 18440 680 18450 700
rect 18410 650 18450 680
rect 18410 630 18420 650
rect 18440 630 18450 650
rect 18410 615 18450 630
rect 18500 900 18540 915
rect 18500 880 18510 900
rect 18530 880 18540 900
rect 18500 850 18540 880
rect 18500 830 18510 850
rect 18530 830 18540 850
rect 18500 800 18540 830
rect 18500 780 18510 800
rect 18530 780 18540 800
rect 18500 750 18540 780
rect 18500 730 18510 750
rect 18530 730 18540 750
rect 18500 700 18540 730
rect 18500 680 18510 700
rect 18530 680 18540 700
rect 18500 650 18540 680
rect 18500 630 18510 650
rect 18530 630 18540 650
rect 18500 615 18540 630
rect 18590 900 18630 915
rect 18590 880 18600 900
rect 18620 880 18630 900
rect 18590 850 18630 880
rect 18590 830 18600 850
rect 18620 830 18630 850
rect 18590 800 18630 830
rect 18590 780 18600 800
rect 18620 780 18630 800
rect 18590 750 18630 780
rect 18590 730 18600 750
rect 18620 730 18630 750
rect 18590 700 18630 730
rect 18905 900 18945 915
rect 18905 880 18915 900
rect 18935 880 18945 900
rect 18905 850 18945 880
rect 18905 830 18915 850
rect 18935 830 18945 850
rect 18905 800 18945 830
rect 18905 780 18915 800
rect 18935 780 18945 800
rect 18905 750 18945 780
rect 18905 730 18915 750
rect 18935 730 18945 750
rect 18905 715 18945 730
rect 18960 900 19000 915
rect 18960 880 18970 900
rect 18990 880 19000 900
rect 18960 850 19000 880
rect 18960 830 18970 850
rect 18990 830 19000 850
rect 18960 800 19000 830
rect 18960 780 18970 800
rect 18990 780 19000 800
rect 18960 750 19000 780
rect 18960 730 18970 750
rect 18990 730 19000 750
rect 18960 715 19000 730
rect 19015 900 19055 915
rect 19015 880 19025 900
rect 19045 880 19055 900
rect 19015 850 19055 880
rect 19015 830 19025 850
rect 19045 830 19055 850
rect 19015 800 19055 830
rect 19015 780 19025 800
rect 19045 780 19055 800
rect 19015 750 19055 780
rect 19015 730 19025 750
rect 19045 730 19055 750
rect 19015 715 19055 730
rect 19070 900 19110 915
rect 19070 880 19080 900
rect 19100 880 19110 900
rect 19070 850 19110 880
rect 19070 830 19080 850
rect 19100 830 19110 850
rect 19070 800 19110 830
rect 19070 780 19080 800
rect 19100 780 19110 800
rect 19070 750 19110 780
rect 19070 730 19080 750
rect 19100 730 19110 750
rect 19070 715 19110 730
rect 18590 680 18600 700
rect 18620 680 18630 700
rect 18590 650 18630 680
rect 18590 630 18600 650
rect 18620 630 18630 650
rect 18590 615 18630 630
rect 16420 120 16460 135
rect 16420 100 16430 120
rect 16450 100 16460 120
rect 16420 70 16460 100
rect 16420 50 16430 70
rect 16450 50 16460 70
rect 16420 35 16460 50
rect 16480 120 16520 135
rect 16480 100 16490 120
rect 16510 100 16520 120
rect 16480 70 16520 100
rect 16480 50 16490 70
rect 16510 50 16520 70
rect 16480 35 16520 50
rect 16540 120 16580 135
rect 16540 100 16550 120
rect 16570 100 16580 120
rect 16540 70 16580 100
rect 16540 50 16550 70
rect 16570 50 16580 70
rect 16540 35 16580 50
rect 16600 120 16640 135
rect 16600 100 16610 120
rect 16630 100 16640 120
rect 16600 70 16640 100
rect 16600 50 16610 70
rect 16630 50 16640 70
rect 16600 35 16640 50
rect 16660 120 16700 135
rect 16660 100 16670 120
rect 16690 100 16700 120
rect 16660 70 16700 100
rect 16660 50 16670 70
rect 16690 50 16700 70
rect 16660 35 16700 50
rect 16720 120 16760 135
rect 16720 100 16730 120
rect 16750 100 16760 120
rect 16720 70 16760 100
rect 16720 50 16730 70
rect 16750 50 16760 70
rect 16720 35 16760 50
rect 16780 120 16820 135
rect 16780 100 16790 120
rect 16810 100 16820 120
rect 16780 70 16820 100
rect 16780 50 16790 70
rect 16810 50 16820 70
rect 16780 35 16820 50
rect 16840 120 16880 135
rect 16840 100 16850 120
rect 16870 100 16880 120
rect 16840 70 16880 100
rect 16840 50 16850 70
rect 16870 50 16880 70
rect 16840 35 16880 50
rect 16900 120 16940 135
rect 16900 100 16910 120
rect 16930 100 16940 120
rect 16900 70 16940 100
rect 16900 50 16910 70
rect 16930 50 16940 70
rect 16900 35 16940 50
rect 16960 120 17000 135
rect 16960 100 16970 120
rect 16990 100 17000 120
rect 16960 70 17000 100
rect 16960 50 16970 70
rect 16990 50 17000 70
rect 16960 35 17000 50
rect 17020 120 17060 135
rect 17020 100 17030 120
rect 17050 100 17060 120
rect 17020 70 17060 100
rect 17020 50 17030 70
rect 17050 50 17060 70
rect 17020 35 17060 50
rect 17080 120 17120 135
rect 17080 100 17090 120
rect 17110 100 17120 120
rect 17080 70 17120 100
rect 17080 50 17090 70
rect 17110 50 17120 70
rect 17080 35 17120 50
rect 17140 120 17180 135
rect 17140 100 17150 120
rect 17170 100 17180 120
rect 17140 70 17180 100
rect 17140 50 17150 70
rect 17170 50 17180 70
rect 17140 35 17180 50
rect 17200 120 17240 135
rect 17200 100 17210 120
rect 17230 100 17240 120
rect 17200 70 17240 100
rect 17200 50 17210 70
rect 17230 50 17240 70
rect 17200 35 17240 50
rect 17260 120 17300 135
rect 17260 100 17270 120
rect 17290 100 17300 120
rect 17260 70 17300 100
rect 17260 50 17270 70
rect 17290 50 17300 70
rect 17260 35 17300 50
rect 17320 120 17360 135
rect 17320 100 17330 120
rect 17350 100 17360 120
rect 17320 70 17360 100
rect 17320 50 17330 70
rect 17350 50 17360 70
rect 17320 35 17360 50
rect 17380 120 17420 135
rect 17380 100 17390 120
rect 17410 100 17420 120
rect 17380 70 17420 100
rect 17380 50 17390 70
rect 17410 50 17420 70
rect 17380 35 17420 50
rect 17440 120 17480 135
rect 17440 100 17450 120
rect 17470 100 17480 120
rect 17440 70 17480 100
rect 17440 50 17450 70
rect 17470 50 17480 70
rect 17440 35 17480 50
rect 17500 120 17540 135
rect 17500 100 17510 120
rect 17530 100 17540 120
rect 17500 70 17540 100
rect 17500 50 17510 70
rect 17530 50 17540 70
rect 17500 35 17540 50
rect 17560 120 17600 135
rect 17560 100 17570 120
rect 17590 100 17600 120
rect 17560 70 17600 100
rect 17560 50 17570 70
rect 17590 50 17600 70
rect 17560 35 17600 50
rect 17620 120 17660 135
rect 17620 100 17630 120
rect 17650 100 17660 120
rect 17620 70 17660 100
rect 17620 50 17630 70
rect 17650 50 17660 70
rect 17620 35 17660 50
rect 17940 120 17980 135
rect 17940 100 17950 120
rect 17970 100 17980 120
rect 17940 70 17980 100
rect 17940 50 17950 70
rect 17970 50 17980 70
rect 17940 35 17980 50
rect 18000 120 18040 135
rect 18000 100 18010 120
rect 18030 100 18040 120
rect 18000 70 18040 100
rect 18000 50 18010 70
rect 18030 50 18040 70
rect 18000 35 18040 50
rect 18060 120 18100 135
rect 18060 100 18070 120
rect 18090 100 18100 120
rect 18060 70 18100 100
rect 18060 50 18070 70
rect 18090 50 18100 70
rect 18060 35 18100 50
rect 18120 120 18160 135
rect 18120 100 18130 120
rect 18150 100 18160 120
rect 18120 70 18160 100
rect 18120 50 18130 70
rect 18150 50 18160 70
rect 18120 35 18160 50
rect 18180 120 18220 135
rect 18180 100 18190 120
rect 18210 100 18220 120
rect 18180 70 18220 100
rect 18180 50 18190 70
rect 18210 50 18220 70
rect 18180 35 18220 50
rect 18240 120 18280 135
rect 18240 100 18250 120
rect 18270 100 18280 120
rect 18240 70 18280 100
rect 18240 50 18250 70
rect 18270 50 18280 70
rect 18240 35 18280 50
rect 18300 120 18340 135
rect 18300 100 18310 120
rect 18330 100 18340 120
rect 18300 70 18340 100
rect 18300 50 18310 70
rect 18330 50 18340 70
rect 18300 35 18340 50
rect 18360 120 18400 135
rect 18360 100 18370 120
rect 18390 100 18400 120
rect 18360 70 18400 100
rect 18360 50 18370 70
rect 18390 50 18400 70
rect 18360 35 18400 50
rect 18420 120 18460 135
rect 18420 100 18430 120
rect 18450 100 18460 120
rect 18420 70 18460 100
rect 18420 50 18430 70
rect 18450 50 18460 70
rect 18420 35 18460 50
rect 18480 120 18520 135
rect 18480 100 18490 120
rect 18510 100 18520 120
rect 18480 70 18520 100
rect 18480 50 18490 70
rect 18510 50 18520 70
rect 18480 35 18520 50
rect 18540 120 18580 135
rect 18540 100 18550 120
rect 18570 100 18580 120
rect 18540 70 18580 100
rect 18540 50 18550 70
rect 18570 50 18580 70
rect 18540 35 18580 50
rect 18600 120 18640 135
rect 18600 100 18610 120
rect 18630 100 18640 120
rect 18600 70 18640 100
rect 18600 50 18610 70
rect 18630 50 18640 70
rect 18600 35 18640 50
rect 18660 120 18700 135
rect 18660 100 18670 120
rect 18690 100 18700 120
rect 18660 70 18700 100
rect 18660 50 18670 70
rect 18690 50 18700 70
rect 18660 35 18700 50
rect 18720 120 18760 135
rect 18720 100 18730 120
rect 18750 100 18760 120
rect 18720 70 18760 100
rect 18720 50 18730 70
rect 18750 50 18760 70
rect 18720 35 18760 50
rect 18780 120 18820 135
rect 18780 100 18790 120
rect 18810 100 18820 120
rect 18780 70 18820 100
rect 18780 50 18790 70
rect 18810 50 18820 70
rect 18780 35 18820 50
rect 18840 120 18880 135
rect 18840 100 18850 120
rect 18870 100 18880 120
rect 18840 70 18880 100
rect 18840 50 18850 70
rect 18870 50 18880 70
rect 18840 35 18880 50
rect 18900 120 18940 135
rect 18900 100 18910 120
rect 18930 100 18940 120
rect 18900 70 18940 100
rect 18900 50 18910 70
rect 18930 50 18940 70
rect 18900 35 18940 50
rect 18960 120 19000 135
rect 18960 100 18970 120
rect 18990 100 19000 120
rect 18960 70 19000 100
rect 18960 50 18970 70
rect 18990 50 19000 70
rect 18960 35 19000 50
rect 19020 120 19060 135
rect 19020 100 19030 120
rect 19050 100 19060 120
rect 19020 70 19060 100
rect 19020 50 19030 70
rect 19050 50 19060 70
rect 19020 35 19060 50
rect 19080 120 19120 135
rect 19080 100 19090 120
rect 19110 100 19120 120
rect 19080 70 19120 100
rect 19080 50 19090 70
rect 19110 50 19120 70
rect 19080 35 19120 50
rect 19140 120 19180 135
rect 19140 100 19150 120
rect 19170 100 19180 120
rect 19140 70 19180 100
rect 19140 50 19150 70
rect 19170 50 19180 70
rect 19140 35 19180 50
<< ndiffc >>
rect 16970 -265 16990 -245
rect 16970 -315 16990 -295
rect 16970 -365 16990 -345
rect 16970 -415 16990 -395
rect 16970 -465 16990 -445
rect 17030 -265 17050 -245
rect 17030 -315 17050 -295
rect 17030 -365 17050 -345
rect 17030 -415 17050 -395
rect 17030 -465 17050 -445
rect 17090 -265 17110 -245
rect 17090 -315 17110 -295
rect 17090 -365 17110 -345
rect 18490 -265 18510 -245
rect 18490 -315 18510 -295
rect 17090 -415 17110 -395
rect 17090 -465 17110 -445
rect 18490 -365 18510 -345
rect 18490 -415 18510 -395
rect 18490 -465 18510 -445
rect 18550 -265 18570 -245
rect 18550 -315 18570 -295
rect 18550 -365 18570 -345
rect 18550 -415 18570 -395
rect 18550 -465 18570 -445
rect 18610 -265 18630 -245
rect 18610 -315 18630 -295
rect 18610 -365 18630 -345
rect 18610 -415 18630 -395
rect 18610 -465 18630 -445
rect 16540 -830 16560 -810
rect 16540 -880 16560 -860
rect 16540 -930 16560 -910
rect 16540 -980 16560 -960
rect 16540 -1030 16560 -1010
rect 17080 -830 17100 -810
rect 17160 -830 17180 -810
rect 17080 -880 17100 -860
rect 17160 -880 17180 -860
rect 17080 -930 17100 -910
rect 17160 -930 17180 -910
rect 17080 -980 17100 -960
rect 17160 -980 17180 -960
rect 17080 -1030 17100 -1010
rect 17160 -1030 17180 -1010
rect 17700 -830 17720 -810
rect 17700 -880 17720 -860
rect 17700 -930 17720 -910
rect 17700 -980 17720 -960
rect 17700 -1030 17720 -1010
rect 17880 -830 17900 -810
rect 17880 -880 17900 -860
rect 17880 -930 17900 -910
rect 17880 -980 17900 -960
rect 17880 -1030 17900 -1010
rect 18420 -830 18440 -810
rect 18500 -830 18520 -810
rect 18420 -880 18440 -860
rect 18500 -880 18520 -860
rect 18420 -930 18440 -910
rect 18500 -930 18520 -910
rect 18420 -980 18440 -960
rect 18500 -980 18520 -960
rect 18420 -1030 18440 -1010
rect 18500 -1030 18520 -1010
rect 19040 -830 19060 -810
rect 19040 -880 19060 -860
rect 19040 -930 19060 -910
rect 19040 -980 19060 -960
rect 19040 -1030 19060 -1010
rect 16750 -1285 16770 -1265
rect 16750 -1335 16770 -1315
rect 17790 -1285 17810 -1265
rect 17790 -1335 17810 -1315
rect 18830 -1285 18850 -1265
rect 18830 -1335 18850 -1315
rect 16610 -1605 16630 -1585
rect 16610 -1655 16630 -1635
rect 16665 -1605 16685 -1585
rect 16665 -1655 16685 -1635
rect 16720 -1605 16740 -1585
rect 16720 -1655 16740 -1635
rect 16775 -1605 16795 -1585
rect 16775 -1655 16795 -1635
rect 16830 -1605 16850 -1585
rect 16830 -1655 16850 -1635
rect 16885 -1605 16905 -1585
rect 16885 -1655 16905 -1635
rect 17035 -1605 17055 -1585
rect 17035 -1655 17055 -1635
rect 17090 -1605 17110 -1585
rect 17090 -1655 17110 -1635
rect 17145 -1605 17165 -1585
rect 17145 -1655 17165 -1635
rect 17200 -1605 17220 -1585
rect 17200 -1655 17220 -1635
rect 17255 -1605 17275 -1585
rect 17255 -1655 17275 -1635
rect 17310 -1605 17330 -1585
rect 17310 -1655 17330 -1635
rect 17365 -1605 17385 -1585
rect 17365 -1655 17385 -1635
rect 17420 -1605 17440 -1585
rect 17420 -1655 17440 -1635
rect 17475 -1605 17495 -1585
rect 17475 -1655 17495 -1635
rect 17625 -1605 17645 -1585
rect 17625 -1655 17645 -1635
rect 17680 -1605 17700 -1585
rect 17680 -1655 17700 -1635
rect 17735 -1605 17755 -1585
rect 17735 -1655 17755 -1635
rect 17790 -1605 17810 -1585
rect 17790 -1655 17810 -1635
rect 17845 -1605 17865 -1585
rect 17845 -1655 17865 -1635
rect 17900 -1605 17920 -1585
rect 17900 -1655 17920 -1635
rect 17955 -1605 17975 -1585
rect 17955 -1655 17975 -1635
rect 18010 -1605 18030 -1585
rect 18010 -1655 18030 -1635
rect 18160 -1605 18180 -1585
rect 18160 -1655 18180 -1635
rect 18215 -1605 18235 -1585
rect 18215 -1655 18235 -1635
rect 18270 -1605 18290 -1585
rect 18270 -1655 18290 -1635
rect 18325 -1605 18345 -1585
rect 18325 -1655 18345 -1635
rect 18380 -1605 18400 -1585
rect 18380 -1655 18400 -1635
rect 18435 -1605 18455 -1585
rect 18435 -1655 18455 -1635
rect 18490 -1605 18510 -1585
rect 18490 -1655 18510 -1635
rect 18545 -1605 18565 -1585
rect 18545 -1655 18565 -1635
rect 18600 -1605 18620 -1585
rect 18600 -1655 18620 -1635
<< pdiffc >>
rect 16385 1240 16405 1260
rect 16385 1190 16405 1210
rect 16440 1240 16460 1260
rect 16440 1190 16460 1210
rect 16495 1240 16515 1260
rect 16495 1190 16515 1210
rect 16550 1240 16570 1260
rect 16550 1190 16570 1210
rect 16605 1240 16625 1260
rect 16605 1190 16625 1210
rect 16895 1188 16915 1260
rect 16950 1188 16970 1260
rect 17005 1188 17025 1260
rect 17060 1188 17080 1260
rect 17115 1188 17135 1260
rect 17170 1188 17190 1260
rect 17225 1188 17245 1260
rect 17515 1240 17535 1260
rect 17515 1190 17535 1210
rect 17570 1240 17590 1260
rect 17570 1190 17590 1210
rect 17625 1240 17645 1260
rect 17625 1190 17645 1210
rect 17680 1240 17700 1260
rect 17680 1190 17700 1210
rect 17735 1240 17755 1260
rect 17735 1190 17755 1210
rect 17790 1240 17810 1260
rect 17790 1190 17810 1210
rect 17845 1240 17865 1260
rect 17845 1190 17865 1210
rect 17900 1240 17920 1260
rect 17900 1190 17920 1210
rect 17955 1240 17975 1260
rect 17955 1190 17975 1210
rect 18010 1240 18030 1260
rect 18010 1190 18030 1210
rect 18065 1240 18085 1260
rect 18065 1190 18085 1210
rect 18355 1190 18375 1260
rect 18410 1190 18430 1260
rect 18465 1190 18485 1260
rect 18520 1190 18540 1260
rect 18575 1190 18595 1260
rect 18630 1190 18650 1260
rect 18685 1190 18705 1260
rect 16980 880 17000 900
rect 16980 830 17000 850
rect 16445 780 16465 800
rect 16445 730 16465 750
rect 16500 780 16520 800
rect 16500 730 16520 750
rect 16555 780 16575 800
rect 16555 730 16575 750
rect 16610 780 16630 800
rect 16610 730 16630 750
rect 16665 780 16685 800
rect 16665 730 16685 750
rect 16980 780 17000 800
rect 16980 730 17000 750
rect 16980 680 17000 700
rect 16980 630 17000 650
rect 17070 880 17090 900
rect 17070 830 17090 850
rect 17070 780 17090 800
rect 17070 730 17090 750
rect 17070 680 17090 700
rect 17070 630 17090 650
rect 17160 880 17180 900
rect 17160 830 17180 850
rect 17160 780 17180 800
rect 17160 730 17180 750
rect 17160 680 17180 700
rect 17160 630 17180 650
rect 17250 880 17270 900
rect 17250 830 17270 850
rect 17250 780 17270 800
rect 17250 730 17270 750
rect 17250 680 17270 700
rect 17250 630 17270 650
rect 17340 880 17360 900
rect 17340 830 17360 850
rect 17340 780 17360 800
rect 17340 730 17360 750
rect 17340 680 17360 700
rect 17340 630 17360 650
rect 17430 880 17450 900
rect 17430 830 17450 850
rect 17430 780 17450 800
rect 17430 730 17450 750
rect 17430 680 17450 700
rect 17430 630 17450 650
rect 17520 880 17540 900
rect 17520 830 17540 850
rect 17520 780 17540 800
rect 17520 730 17540 750
rect 17520 680 17540 700
rect 17520 630 17540 650
rect 17610 880 17630 900
rect 17610 830 17630 850
rect 17610 780 17630 800
rect 17610 730 17630 750
rect 17610 680 17630 700
rect 17610 630 17630 650
rect 17700 880 17720 900
rect 17700 830 17720 850
rect 17700 780 17720 800
rect 17700 730 17720 750
rect 17700 680 17720 700
rect 17700 630 17720 650
rect 17790 880 17810 900
rect 17790 830 17810 850
rect 17790 780 17810 800
rect 17790 730 17810 750
rect 17790 680 17810 700
rect 17790 630 17810 650
rect 17880 880 17900 900
rect 17880 830 17900 850
rect 17880 780 17900 800
rect 17880 730 17900 750
rect 17880 680 17900 700
rect 17880 630 17900 650
rect 17970 880 17990 900
rect 17970 830 17990 850
rect 17970 780 17990 800
rect 17970 730 17990 750
rect 17970 680 17990 700
rect 17970 630 17990 650
rect 18060 880 18080 900
rect 18060 830 18080 850
rect 18060 780 18080 800
rect 18060 730 18080 750
rect 18060 680 18080 700
rect 18060 630 18080 650
rect 18150 880 18170 900
rect 18150 830 18170 850
rect 18150 780 18170 800
rect 18150 730 18170 750
rect 18150 680 18170 700
rect 18150 630 18170 650
rect 18240 880 18260 900
rect 18240 830 18260 850
rect 18240 780 18260 800
rect 18240 730 18260 750
rect 18240 680 18260 700
rect 18240 630 18260 650
rect 18330 880 18350 900
rect 18330 830 18350 850
rect 18330 780 18350 800
rect 18330 730 18350 750
rect 18330 680 18350 700
rect 18330 630 18350 650
rect 18420 880 18440 900
rect 18420 830 18440 850
rect 18420 780 18440 800
rect 18420 730 18440 750
rect 18420 680 18440 700
rect 18420 630 18440 650
rect 18510 880 18530 900
rect 18510 830 18530 850
rect 18510 780 18530 800
rect 18510 730 18530 750
rect 18510 680 18530 700
rect 18510 630 18530 650
rect 18600 880 18620 900
rect 18600 830 18620 850
rect 18600 780 18620 800
rect 18600 730 18620 750
rect 18915 880 18935 900
rect 18915 830 18935 850
rect 18915 780 18935 800
rect 18915 730 18935 750
rect 18970 880 18990 900
rect 18970 830 18990 850
rect 18970 780 18990 800
rect 18970 730 18990 750
rect 19025 880 19045 900
rect 19025 830 19045 850
rect 19025 780 19045 800
rect 19025 730 19045 750
rect 19080 880 19100 900
rect 19080 830 19100 850
rect 19080 780 19100 800
rect 19080 730 19100 750
rect 18600 680 18620 700
rect 18600 630 18620 650
rect 16430 100 16450 120
rect 16430 50 16450 70
rect 16490 100 16510 120
rect 16490 50 16510 70
rect 16550 100 16570 120
rect 16550 50 16570 70
rect 16610 100 16630 120
rect 16610 50 16630 70
rect 16670 100 16690 120
rect 16670 50 16690 70
rect 16730 100 16750 120
rect 16730 50 16750 70
rect 16790 100 16810 120
rect 16790 50 16810 70
rect 16850 100 16870 120
rect 16850 50 16870 70
rect 16910 100 16930 120
rect 16910 50 16930 70
rect 16970 100 16990 120
rect 16970 50 16990 70
rect 17030 100 17050 120
rect 17030 50 17050 70
rect 17090 100 17110 120
rect 17090 50 17110 70
rect 17150 100 17170 120
rect 17150 50 17170 70
rect 17210 100 17230 120
rect 17210 50 17230 70
rect 17270 100 17290 120
rect 17270 50 17290 70
rect 17330 100 17350 120
rect 17330 50 17350 70
rect 17390 100 17410 120
rect 17390 50 17410 70
rect 17450 100 17470 120
rect 17450 50 17470 70
rect 17510 100 17530 120
rect 17510 50 17530 70
rect 17570 100 17590 120
rect 17570 50 17590 70
rect 17630 100 17650 120
rect 17630 50 17650 70
rect 17950 100 17970 120
rect 17950 50 17970 70
rect 18010 100 18030 120
rect 18010 50 18030 70
rect 18070 100 18090 120
rect 18070 50 18090 70
rect 18130 100 18150 120
rect 18130 50 18150 70
rect 18190 100 18210 120
rect 18190 50 18210 70
rect 18250 100 18270 120
rect 18250 50 18270 70
rect 18310 100 18330 120
rect 18310 50 18330 70
rect 18370 100 18390 120
rect 18370 50 18390 70
rect 18430 100 18450 120
rect 18430 50 18450 70
rect 18490 100 18510 120
rect 18490 50 18510 70
rect 18550 100 18570 120
rect 18550 50 18570 70
rect 18610 100 18630 120
rect 18610 50 18630 70
rect 18670 100 18690 120
rect 18670 50 18690 70
rect 18730 100 18750 120
rect 18730 50 18750 70
rect 18790 100 18810 120
rect 18790 50 18810 70
rect 18850 100 18870 120
rect 18850 50 18870 70
rect 18910 100 18930 120
rect 18910 50 18930 70
rect 18970 100 18990 120
rect 18970 50 18990 70
rect 19030 100 19050 120
rect 19030 50 19050 70
rect 19090 100 19110 120
rect 19090 50 19110 70
rect 19150 100 19170 120
rect 19150 50 19170 70
<< psubdiff >>
rect 17560 -245 17600 -230
rect 17560 -265 17570 -245
rect 17590 -265 17600 -245
rect 17560 -285 17600 -265
rect 17560 -305 17570 -285
rect 17590 -305 17600 -285
rect 17560 -325 17600 -305
rect 17560 -345 17570 -325
rect 17590 -345 17600 -325
rect 17560 -360 17600 -345
rect 18000 -245 18040 -230
rect 18000 -265 18010 -245
rect 18030 -265 18040 -245
rect 18000 -285 18040 -265
rect 18000 -305 18010 -285
rect 18030 -305 18040 -285
rect 18000 -325 18040 -305
rect 18000 -345 18010 -325
rect 18030 -345 18040 -325
rect 18000 -360 18040 -345
rect 17110 -810 17150 -795
rect 17110 -830 17120 -810
rect 17140 -830 17150 -810
rect 17110 -860 17150 -830
rect 17110 -880 17120 -860
rect 17140 -880 17150 -860
rect 17110 -910 17150 -880
rect 17110 -930 17120 -910
rect 17140 -930 17150 -910
rect 17110 -960 17150 -930
rect 17110 -980 17120 -960
rect 17140 -980 17150 -960
rect 17110 -1010 17150 -980
rect 17110 -1030 17120 -1010
rect 17140 -1030 17150 -1010
rect 17110 -1040 17150 -1030
rect 18450 -810 18490 -795
rect 18450 -830 18460 -810
rect 18480 -830 18490 -810
rect 18450 -860 18490 -830
rect 18450 -880 18460 -860
rect 18480 -880 18490 -860
rect 18450 -910 18490 -880
rect 18450 -930 18460 -910
rect 18480 -930 18490 -910
rect 18450 -960 18490 -930
rect 18450 -980 18460 -960
rect 18480 -980 18490 -960
rect 18450 -1010 18490 -980
rect 18450 -1030 18460 -1010
rect 18480 -1030 18490 -1010
rect 18450 -1045 18490 -1030
rect 18860 -1265 18900 -1250
rect 18860 -1285 18870 -1265
rect 18890 -1285 18900 -1265
rect 18860 -1315 18900 -1285
rect 18860 -1335 18870 -1315
rect 18890 -1335 18900 -1315
rect 18860 -1350 18900 -1335
rect 16560 -1585 16600 -1570
rect 16560 -1605 16570 -1585
rect 16590 -1605 16600 -1585
rect 16560 -1635 16600 -1605
rect 16560 -1655 16570 -1635
rect 16590 -1655 16600 -1635
rect 16560 -1670 16600 -1655
rect 16915 -1585 16955 -1570
rect 16915 -1605 16925 -1585
rect 16945 -1605 16955 -1585
rect 16915 -1635 16955 -1605
rect 16915 -1655 16925 -1635
rect 16945 -1655 16955 -1635
rect 16915 -1670 16955 -1655
rect 16985 -1585 17025 -1570
rect 16985 -1605 16995 -1585
rect 17015 -1605 17025 -1585
rect 16985 -1635 17025 -1605
rect 16985 -1655 16995 -1635
rect 17015 -1655 17025 -1635
rect 16985 -1670 17025 -1655
rect 17505 -1585 17545 -1570
rect 17505 -1605 17515 -1585
rect 17535 -1605 17545 -1585
rect 17505 -1635 17545 -1605
rect 17505 -1655 17515 -1635
rect 17535 -1655 17545 -1635
rect 17505 -1670 17545 -1655
rect 17575 -1585 17615 -1570
rect 17575 -1605 17585 -1585
rect 17605 -1605 17615 -1585
rect 17575 -1635 17615 -1605
rect 17575 -1655 17585 -1635
rect 17605 -1655 17615 -1635
rect 17575 -1670 17615 -1655
rect 18040 -1585 18080 -1570
rect 18040 -1605 18050 -1585
rect 18070 -1605 18080 -1585
rect 18040 -1635 18080 -1605
rect 18040 -1655 18050 -1635
rect 18070 -1655 18080 -1635
rect 18040 -1670 18080 -1655
rect 18110 -1585 18150 -1570
rect 18110 -1605 18120 -1585
rect 18140 -1605 18150 -1585
rect 18110 -1635 18150 -1605
rect 18110 -1655 18120 -1635
rect 18140 -1655 18150 -1635
rect 18110 -1670 18150 -1655
rect 18630 -1585 18670 -1570
rect 18630 -1605 18640 -1585
rect 18660 -1605 18670 -1585
rect 18630 -1635 18670 -1605
rect 18630 -1655 18640 -1635
rect 18660 -1655 18670 -1635
rect 18630 -1670 18670 -1655
rect 17775 -4210 17825 -4195
rect 17775 -4230 17790 -4210
rect 17810 -4230 17825 -4210
rect 17775 -4250 17825 -4230
rect 17775 -4270 17790 -4250
rect 17810 -4270 17825 -4250
rect 17775 -4290 17825 -4270
rect 17775 -4310 17790 -4290
rect 17810 -4310 17825 -4290
rect 17775 -4325 17825 -4310
<< nsubdiff >>
rect 16335 1262 16375 1275
rect 16335 1240 16345 1262
rect 16365 1240 16375 1262
rect 16335 1210 16375 1240
rect 16335 1190 16345 1210
rect 16365 1190 16375 1210
rect 16335 1175 16375 1190
rect 16635 1262 16675 1275
rect 16635 1240 16645 1262
rect 16665 1240 16675 1262
rect 16635 1210 16675 1240
rect 16635 1190 16645 1210
rect 16665 1190 16675 1210
rect 16635 1175 16675 1190
rect 16845 1262 16885 1275
rect 16845 1190 16855 1262
rect 16875 1190 16885 1262
rect 16845 1175 16885 1190
rect 17255 1262 17295 1275
rect 17255 1190 17265 1262
rect 17285 1190 17295 1262
rect 17255 1175 17295 1190
rect 17465 1262 17505 1275
rect 17465 1240 17475 1262
rect 17495 1240 17505 1262
rect 17465 1210 17505 1240
rect 17465 1190 17475 1210
rect 17495 1190 17505 1210
rect 17465 1175 17505 1190
rect 18095 1262 18135 1275
rect 18095 1240 18105 1262
rect 18125 1240 18135 1262
rect 18095 1210 18135 1240
rect 18095 1190 18105 1210
rect 18125 1190 18135 1210
rect 18095 1175 18135 1190
rect 18305 1262 18345 1275
rect 18305 1190 18315 1262
rect 18335 1190 18345 1262
rect 18305 1175 18345 1190
rect 18715 1262 18755 1275
rect 18715 1190 18725 1262
rect 18745 1190 18755 1262
rect 18715 1175 18755 1190
rect 16930 900 16970 915
rect 16930 880 16940 900
rect 16960 880 16970 900
rect 16930 850 16970 880
rect 16930 830 16940 850
rect 16960 830 16970 850
rect 16395 800 16435 815
rect 16395 780 16405 800
rect 16425 780 16435 800
rect 16395 750 16435 780
rect 16395 730 16405 750
rect 16425 730 16435 750
rect 16395 715 16435 730
rect 16700 800 16740 815
rect 16700 780 16710 800
rect 16730 780 16740 800
rect 16700 750 16740 780
rect 16700 730 16710 750
rect 16730 730 16740 750
rect 16700 715 16740 730
rect 16930 800 16970 830
rect 16930 780 16940 800
rect 16960 780 16970 800
rect 16930 750 16970 780
rect 16930 730 16940 750
rect 16960 730 16970 750
rect 16930 700 16970 730
rect 16930 680 16940 700
rect 16960 680 16970 700
rect 16930 650 16970 680
rect 16930 630 16940 650
rect 16960 630 16970 650
rect 16930 615 16970 630
rect 18630 900 18670 915
rect 18630 880 18640 900
rect 18660 880 18670 900
rect 18630 850 18670 880
rect 18630 830 18640 850
rect 18660 830 18670 850
rect 18630 800 18670 830
rect 18630 780 18640 800
rect 18660 780 18670 800
rect 18630 750 18670 780
rect 18630 730 18640 750
rect 18660 730 18670 750
rect 18630 700 18670 730
rect 18865 900 18905 915
rect 18865 880 18875 900
rect 18895 880 18905 900
rect 18865 850 18905 880
rect 18865 830 18875 850
rect 18895 830 18905 850
rect 18865 800 18905 830
rect 18865 780 18875 800
rect 18895 780 18905 800
rect 18865 750 18905 780
rect 18865 730 18875 750
rect 18895 730 18905 750
rect 18865 715 18905 730
rect 19110 900 19150 915
rect 19110 880 19120 900
rect 19140 880 19150 900
rect 19110 850 19150 880
rect 19110 830 19120 850
rect 19140 830 19150 850
rect 19110 800 19150 830
rect 19110 780 19120 800
rect 19140 780 19150 800
rect 19110 750 19150 780
rect 19110 730 19120 750
rect 19140 730 19150 750
rect 19110 715 19150 730
rect 18630 680 18640 700
rect 18660 680 18670 700
rect 18630 650 18670 680
rect 18630 630 18640 650
rect 18660 630 18670 650
rect 18630 615 18670 630
rect 16380 120 16420 135
rect 16380 100 16390 120
rect 16410 100 16420 120
rect 16380 70 16420 100
rect 16380 50 16390 70
rect 16410 50 16420 70
rect 16380 35 16420 50
rect 17660 120 17700 135
rect 17660 100 17670 120
rect 17690 100 17700 120
rect 17660 70 17700 100
rect 17660 50 17670 70
rect 17690 50 17700 70
rect 17660 35 17700 50
rect 17900 120 17940 135
rect 17900 100 17910 120
rect 17930 100 17940 120
rect 17900 70 17940 100
rect 17900 50 17910 70
rect 17930 50 17940 70
rect 17900 35 17940 50
rect 19180 120 19220 135
rect 19180 100 19190 120
rect 19210 100 19220 120
rect 19180 70 19220 100
rect 19180 50 19190 70
rect 19210 50 19220 70
rect 19180 35 19220 50
<< psubdiffcont >>
rect 17570 -265 17590 -245
rect 17570 -305 17590 -285
rect 17570 -345 17590 -325
rect 18010 -265 18030 -245
rect 18010 -305 18030 -285
rect 18010 -345 18030 -325
rect 17120 -830 17140 -810
rect 17120 -880 17140 -860
rect 17120 -930 17140 -910
rect 17120 -980 17140 -960
rect 17120 -1030 17140 -1010
rect 18460 -830 18480 -810
rect 18460 -880 18480 -860
rect 18460 -930 18480 -910
rect 18460 -980 18480 -960
rect 18460 -1030 18480 -1010
rect 18870 -1285 18890 -1265
rect 18870 -1335 18890 -1315
rect 16570 -1605 16590 -1585
rect 16570 -1655 16590 -1635
rect 16925 -1605 16945 -1585
rect 16925 -1655 16945 -1635
rect 16995 -1605 17015 -1585
rect 16995 -1655 17015 -1635
rect 17515 -1605 17535 -1585
rect 17515 -1655 17535 -1635
rect 17585 -1605 17605 -1585
rect 17585 -1655 17605 -1635
rect 18050 -1605 18070 -1585
rect 18050 -1655 18070 -1635
rect 18120 -1605 18140 -1585
rect 18120 -1655 18140 -1635
rect 18640 -1605 18660 -1585
rect 18640 -1655 18660 -1635
rect 17790 -4230 17810 -4210
rect 17790 -4270 17810 -4250
rect 17790 -4310 17810 -4290
<< nsubdiffcont >>
rect 16345 1240 16365 1262
rect 16345 1190 16365 1210
rect 16645 1240 16665 1262
rect 16645 1190 16665 1210
rect 16855 1190 16875 1262
rect 17265 1190 17285 1262
rect 17475 1240 17495 1262
rect 17475 1190 17495 1210
rect 18105 1240 18125 1262
rect 18105 1190 18125 1210
rect 18315 1190 18335 1262
rect 18725 1190 18745 1262
rect 16940 880 16960 900
rect 16940 830 16960 850
rect 16405 780 16425 800
rect 16405 730 16425 750
rect 16710 780 16730 800
rect 16710 730 16730 750
rect 16940 780 16960 800
rect 16940 730 16960 750
rect 16940 680 16960 700
rect 16940 630 16960 650
rect 18640 880 18660 900
rect 18640 830 18660 850
rect 18640 780 18660 800
rect 18640 730 18660 750
rect 18875 880 18895 900
rect 18875 830 18895 850
rect 18875 780 18895 800
rect 18875 730 18895 750
rect 19120 880 19140 900
rect 19120 830 19140 850
rect 19120 780 19140 800
rect 19120 730 19140 750
rect 18640 680 18660 700
rect 18640 630 18660 650
rect 16390 100 16410 120
rect 16390 50 16410 70
rect 17670 100 17690 120
rect 17670 50 17690 70
rect 17910 100 17930 120
rect 17910 50 17930 70
rect 19190 100 19210 120
rect 19190 50 19210 70
<< poly >>
rect 16485 1455 16525 1465
rect 16485 1435 16495 1455
rect 16515 1435 16525 1455
rect 16485 1425 16525 1435
rect 17780 1455 17820 1465
rect 17780 1435 17790 1455
rect 17810 1435 17820 1455
rect 17780 1425 17820 1435
rect 16365 1320 16405 1330
rect 16365 1300 16375 1320
rect 16395 1305 16405 1320
rect 16395 1300 16430 1305
rect 16495 1300 16515 1425
rect 16605 1320 16645 1330
rect 16605 1305 16615 1320
rect 16580 1300 16615 1305
rect 16635 1300 16645 1320
rect 16365 1290 16430 1300
rect 16415 1275 16430 1290
rect 16470 1285 16540 1300
rect 16470 1275 16485 1285
rect 16525 1275 16540 1285
rect 16580 1290 16645 1300
rect 16885 1320 16925 1330
rect 16885 1300 16895 1320
rect 16915 1300 16925 1320
rect 17055 1320 17085 1330
rect 17055 1300 17060 1320
rect 17080 1300 17085 1320
rect 17215 1320 17255 1330
rect 17215 1300 17225 1320
rect 17245 1300 17255 1320
rect 16580 1275 16595 1290
rect 16885 1285 16940 1300
rect 16925 1275 16940 1285
rect 16980 1285 17160 1300
rect 16980 1275 16995 1285
rect 17035 1275 17050 1285
rect 17090 1275 17105 1285
rect 17145 1275 17160 1285
rect 17200 1285 17255 1300
rect 17495 1320 17535 1330
rect 17495 1300 17505 1320
rect 17525 1305 17535 1320
rect 17525 1300 17560 1305
rect 17790 1300 17810 1425
rect 18065 1320 18105 1330
rect 18065 1305 18075 1320
rect 18040 1300 18075 1305
rect 18095 1300 18105 1320
rect 17495 1290 17560 1300
rect 17200 1275 17215 1285
rect 17545 1275 17560 1290
rect 17600 1285 18000 1300
rect 17600 1275 17615 1285
rect 17655 1275 17670 1285
rect 17710 1275 17725 1285
rect 17765 1275 17780 1285
rect 17820 1275 17835 1285
rect 17875 1275 17890 1285
rect 17930 1275 17945 1285
rect 17985 1275 18000 1285
rect 18040 1290 18105 1300
rect 18345 1320 18385 1330
rect 18345 1300 18355 1320
rect 18375 1305 18385 1320
rect 18515 1320 18545 1330
rect 18375 1300 18400 1305
rect 18515 1300 18520 1320
rect 18540 1300 18545 1320
rect 18675 1320 18715 1330
rect 18675 1305 18685 1320
rect 18660 1300 18685 1305
rect 18705 1300 18715 1320
rect 18345 1290 18400 1300
rect 18040 1275 18055 1290
rect 18385 1275 18400 1290
rect 18440 1285 18620 1300
rect 18440 1275 18455 1285
rect 18495 1275 18510 1285
rect 18550 1275 18565 1285
rect 18605 1275 18620 1285
rect 18660 1290 18715 1300
rect 18660 1275 18675 1290
rect 16415 1160 16430 1175
rect 16470 1160 16485 1175
rect 16525 1160 16540 1175
rect 16580 1160 16595 1175
rect 16925 1160 16940 1175
rect 16980 1160 16995 1175
rect 17035 1160 17050 1175
rect 17090 1160 17105 1175
rect 17145 1160 17160 1175
rect 17200 1160 17215 1175
rect 17545 1160 17560 1175
rect 17600 1160 17615 1175
rect 17655 1160 17670 1175
rect 17710 1160 17725 1175
rect 17765 1160 17780 1175
rect 17820 1160 17835 1175
rect 17875 1160 17890 1175
rect 17930 1160 17945 1175
rect 17985 1160 18000 1175
rect 18040 1160 18055 1175
rect 18385 1160 18400 1175
rect 18440 1160 18455 1175
rect 18495 1160 18510 1175
rect 18550 1160 18565 1175
rect 18605 1160 18620 1175
rect 18660 1160 18675 1175
rect 16970 960 17010 970
rect 16970 940 16980 960
rect 17000 945 17010 960
rect 18590 960 18630 970
rect 18590 945 18600 960
rect 17000 940 17060 945
rect 16970 930 17060 940
rect 18540 940 18600 945
rect 18620 940 18630 960
rect 18540 930 18630 940
rect 18910 960 18940 970
rect 18910 940 18915 960
rect 18935 945 18940 960
rect 19080 960 19110 970
rect 19080 945 19085 960
rect 18935 940 18960 945
rect 18910 930 18960 940
rect 19055 940 19085 945
rect 19105 940 19110 960
rect 19055 930 19110 940
rect 17010 915 17060 930
rect 17100 915 17150 930
rect 17190 915 17240 930
rect 17280 915 17330 930
rect 17370 915 17420 930
rect 17460 915 17510 930
rect 17550 915 17600 930
rect 17640 915 17690 930
rect 17730 915 17780 930
rect 17820 915 17870 930
rect 17910 915 17960 930
rect 18000 915 18050 930
rect 18090 915 18140 930
rect 18180 915 18230 930
rect 18270 915 18320 930
rect 18360 915 18410 930
rect 18450 915 18500 930
rect 18540 915 18590 930
rect 18945 915 18960 930
rect 19000 915 19015 930
rect 19055 915 19070 930
rect 16440 860 16470 870
rect 16440 840 16445 860
rect 16465 840 16470 860
rect 16660 860 16690 870
rect 16660 840 16665 860
rect 16685 840 16690 860
rect 16440 825 16490 840
rect 16475 815 16490 825
rect 16530 815 16545 830
rect 16585 815 16600 830
rect 16640 825 16690 840
rect 16640 815 16655 825
rect 16475 700 16490 715
rect 16530 705 16545 715
rect 16585 705 16600 715
rect 16530 690 16600 705
rect 16640 700 16655 715
rect 16545 670 16555 690
rect 16575 670 16585 690
rect 16545 660 16585 670
rect 18945 700 18960 715
rect 19000 640 19015 715
rect 19055 700 19070 715
rect 19000 630 19040 640
rect 17010 600 17060 615
rect 17100 595 17150 615
rect 17190 600 17240 615
rect 17280 600 17330 615
rect 17370 600 17420 615
rect 17460 600 17510 615
rect 17550 600 17600 615
rect 17640 600 17690 615
rect 17730 600 17780 615
rect 17820 600 17870 615
rect 17910 600 17960 615
rect 18000 600 18050 615
rect 18090 600 18140 615
rect 18180 600 18230 615
rect 18270 600 18320 615
rect 18360 600 18410 615
rect 18450 600 18500 615
rect 18540 600 18590 615
rect 19000 610 19010 630
rect 19030 610 19040 630
rect 19000 600 19040 610
rect 17110 590 17145 595
rect 17110 570 17115 590
rect 17135 570 17145 590
rect 17110 560 17145 570
rect 17195 590 17235 600
rect 17195 570 17205 590
rect 17225 570 17235 590
rect 17195 560 17235 570
rect 17285 590 17325 600
rect 17285 570 17295 590
rect 17315 570 17325 590
rect 17285 560 17325 570
rect 17375 590 17415 600
rect 17375 570 17385 590
rect 17405 570 17415 590
rect 17375 560 17415 570
rect 17465 590 17505 600
rect 17465 570 17475 590
rect 17495 570 17505 590
rect 17465 560 17505 570
rect 17555 590 17595 600
rect 17555 570 17565 590
rect 17585 570 17595 590
rect 17555 560 17595 570
rect 17645 590 17685 600
rect 17645 570 17655 590
rect 17675 570 17685 590
rect 17645 560 17685 570
rect 17735 590 17770 600
rect 17735 570 17745 590
rect 17765 570 17770 590
rect 17735 560 17770 570
rect 17830 590 17865 600
rect 17830 570 17835 590
rect 17855 570 17865 590
rect 17830 560 17865 570
rect 17915 590 17955 600
rect 17915 570 17925 590
rect 17945 570 17955 590
rect 17915 560 17955 570
rect 18005 590 18045 600
rect 18005 570 18015 590
rect 18035 570 18045 590
rect 18005 560 18045 570
rect 18095 590 18135 600
rect 18095 570 18105 590
rect 18125 570 18135 590
rect 18095 560 18135 570
rect 18185 590 18225 600
rect 18185 570 18195 590
rect 18215 570 18225 590
rect 18185 560 18225 570
rect 18275 590 18315 600
rect 18275 570 18285 590
rect 18305 570 18315 590
rect 18275 560 18315 570
rect 18365 590 18405 600
rect 18365 570 18375 590
rect 18395 570 18405 590
rect 18365 560 18405 570
rect 18455 590 18490 600
rect 18455 570 18465 590
rect 18485 570 18490 590
rect 18455 560 18490 570
rect 16425 180 16455 190
rect 16425 160 16430 180
rect 16450 165 16455 180
rect 17625 180 17655 190
rect 17625 165 17630 180
rect 16450 160 16480 165
rect 16425 150 16480 160
rect 17600 160 17630 165
rect 17650 160 17655 180
rect 17600 150 17655 160
rect 17945 180 17975 190
rect 17945 160 17950 180
rect 17970 165 17975 180
rect 19145 180 19175 190
rect 19145 165 19150 180
rect 17970 160 18000 165
rect 17945 150 18000 160
rect 19120 160 19150 165
rect 19170 160 19175 180
rect 19120 150 19175 160
rect 16460 135 16480 150
rect 16520 135 16540 150
rect 16580 135 16600 150
rect 16640 135 16660 150
rect 16700 135 16720 150
rect 16760 135 16780 150
rect 16820 135 16840 150
rect 16880 135 16900 150
rect 16940 135 16960 150
rect 17000 135 17020 150
rect 17060 135 17080 150
rect 17120 135 17140 150
rect 17180 135 17200 150
rect 17240 135 17260 150
rect 17300 135 17320 150
rect 17360 135 17380 150
rect 17420 135 17440 150
rect 17480 135 17500 150
rect 17540 135 17560 150
rect 17600 135 17620 150
rect 17980 135 18000 150
rect 18040 135 18060 150
rect 18100 135 18120 150
rect 18160 135 18180 150
rect 18220 135 18240 150
rect 18280 135 18300 150
rect 18340 135 18360 150
rect 18400 135 18420 150
rect 18460 135 18480 150
rect 18520 135 18540 150
rect 18580 135 18600 150
rect 18640 135 18660 150
rect 18700 135 18720 150
rect 18760 135 18780 150
rect 18820 135 18840 150
rect 18880 135 18900 150
rect 18940 135 18960 150
rect 19000 135 19020 150
rect 19060 135 19080 150
rect 19120 135 19140 150
rect 16460 20 16480 35
rect 16520 15 16540 35
rect 16580 25 16600 35
rect 16640 25 16660 35
rect 16700 25 16720 35
rect 16760 25 16780 35
rect 16515 5 16545 15
rect 16580 10 16780 25
rect 16820 25 16840 35
rect 16880 25 16900 35
rect 16820 10 16900 25
rect 16940 25 16960 35
rect 17000 25 17020 35
rect 17060 25 17080 35
rect 17120 25 17140 35
rect 16940 10 17140 25
rect 17180 25 17200 35
rect 17240 25 17260 35
rect 17180 10 17260 25
rect 17300 25 17320 35
rect 17360 25 17380 35
rect 17420 25 17440 35
rect 17480 25 17500 35
rect 17300 10 17500 25
rect 17540 20 17560 35
rect 17600 20 17620 35
rect 17980 20 18000 35
rect 18040 20 18060 35
rect 18100 25 18120 35
rect 18160 25 18180 35
rect 18220 25 18240 35
rect 18280 25 18300 35
rect 17535 10 17565 20
rect 16515 -15 16520 5
rect 16540 -15 16545 5
rect 16515 -25 16545 -15
rect 16600 -10 16610 10
rect 16630 -10 16640 10
rect 16600 -20 16640 -10
rect 16845 -10 16850 10
rect 16870 -10 16875 10
rect 16845 -20 16875 -10
rect 16960 -10 16970 10
rect 16990 -10 17000 10
rect 16960 -20 17000 -10
rect 17205 -10 17210 10
rect 17230 -10 17235 10
rect 17205 -20 17235 -10
rect 17320 -10 17330 10
rect 17350 -10 17360 10
rect 17320 -20 17360 -10
rect 17535 -10 17540 10
rect 17560 -10 17565 10
rect 17535 -20 17565 -10
rect 18035 10 18065 20
rect 18100 10 18300 25
rect 18340 25 18360 35
rect 18400 25 18420 35
rect 18340 10 18420 25
rect 18460 25 18480 35
rect 18520 25 18540 35
rect 18580 25 18600 35
rect 18640 25 18660 35
rect 18460 10 18660 25
rect 18700 25 18720 35
rect 18760 25 18780 35
rect 18700 10 18780 25
rect 18820 25 18840 35
rect 18880 25 18900 35
rect 18940 25 18960 35
rect 19000 25 19020 35
rect 18820 10 19020 25
rect 19060 15 19080 35
rect 19120 20 19140 35
rect 18035 -10 18040 10
rect 18060 -10 18065 10
rect 18035 -20 18065 -10
rect 18240 -10 18250 10
rect 18270 -10 18280 10
rect 18240 -20 18280 -10
rect 18365 -10 18370 10
rect 18390 -10 18395 10
rect 18365 -20 18395 -10
rect 18600 -10 18610 10
rect 18630 -10 18640 10
rect 18600 -20 18640 -10
rect 18725 -10 18730 10
rect 18750 -10 18755 10
rect 18725 -20 18755 -10
rect 18960 -10 18970 10
rect 18990 -10 19000 10
rect 18960 -20 19000 -10
rect 19055 5 19085 15
rect 19055 -15 19060 5
rect 19080 -15 19085 5
rect 19055 -25 19085 -15
rect 17007 -185 17037 -175
rect 17007 -200 17012 -185
rect 17000 -205 17012 -200
rect 17032 -205 17037 -185
rect 17000 -215 17037 -205
rect 18563 -185 18593 -175
rect 18563 -205 18568 -185
rect 18588 -200 18593 -185
rect 18588 -205 18600 -200
rect 18563 -215 18600 -205
rect 17000 -230 17020 -215
rect 17060 -230 17080 -215
rect 18520 -230 18540 -215
rect 18580 -230 18600 -215
rect 17000 -495 17020 -480
rect 17060 -495 17080 -480
rect 18520 -495 18540 -480
rect 18580 -495 18600 -480
rect 17060 -505 17105 -495
rect 17060 -525 17080 -505
rect 17100 -525 17105 -505
rect 17060 -535 17105 -525
rect 18440 -505 18540 -495
rect 18440 -525 18445 -505
rect 18465 -510 18540 -505
rect 18465 -525 18470 -510
rect 18440 -535 18470 -525
rect 16620 -750 16660 -740
rect 16620 -770 16630 -750
rect 16650 -770 16660 -750
rect 16620 -780 16660 -770
rect 16740 -750 16780 -740
rect 16740 -770 16750 -750
rect 16770 -770 16780 -750
rect 16740 -780 16780 -770
rect 16860 -750 16900 -740
rect 16860 -770 16870 -750
rect 16890 -770 16900 -750
rect 16860 -780 16900 -770
rect 16980 -750 17020 -740
rect 16980 -770 16990 -750
rect 17010 -770 17020 -750
rect 16980 -780 17020 -770
rect 17300 -750 17340 -740
rect 17300 -770 17310 -750
rect 17330 -770 17340 -750
rect 17300 -780 17340 -770
rect 17420 -750 17460 -740
rect 17420 -770 17430 -750
rect 17450 -770 17460 -750
rect 17420 -780 17460 -770
rect 17540 -750 17580 -740
rect 17540 -770 17550 -750
rect 17570 -770 17580 -750
rect 17540 -780 17580 -770
rect 18020 -750 18060 -740
rect 18020 -770 18030 -750
rect 18050 -770 18060 -750
rect 18020 -780 18060 -770
rect 18140 -750 18180 -740
rect 18140 -770 18150 -750
rect 18170 -770 18180 -750
rect 18140 -780 18180 -770
rect 18260 -750 18300 -740
rect 18260 -770 18270 -750
rect 18290 -770 18300 -750
rect 18260 -780 18300 -770
rect 18580 -750 18620 -740
rect 18580 -770 18590 -750
rect 18610 -770 18620 -750
rect 18580 -780 18620 -770
rect 18700 -750 18740 -740
rect 18700 -770 18710 -750
rect 18730 -770 18740 -750
rect 18700 -780 18740 -770
rect 18820 -750 18860 -740
rect 18820 -770 18830 -750
rect 18850 -770 18860 -750
rect 18820 -780 18860 -770
rect 18940 -750 18980 -740
rect 18940 -770 18950 -750
rect 18970 -770 18980 -750
rect 18940 -780 18980 -770
rect 16570 -795 17070 -780
rect 17190 -795 17690 -780
rect 17910 -795 18410 -780
rect 18530 -795 19030 -780
rect 16570 -1060 17070 -1045
rect 17190 -1060 17690 -1045
rect 17910 -1060 18410 -1045
rect 18530 -1060 19030 -1045
rect 16820 -1205 16860 -1195
rect 16820 -1225 16830 -1205
rect 16850 -1225 16860 -1205
rect 16820 -1235 16860 -1225
rect 16900 -1205 16940 -1195
rect 16900 -1225 16910 -1205
rect 16930 -1225 16940 -1205
rect 16900 -1235 16940 -1225
rect 16980 -1205 17020 -1195
rect 16980 -1225 16990 -1205
rect 17010 -1225 17020 -1205
rect 16980 -1235 17020 -1225
rect 17060 -1205 17100 -1195
rect 17060 -1225 17070 -1205
rect 17090 -1225 17100 -1205
rect 17060 -1235 17100 -1225
rect 17140 -1205 17180 -1195
rect 17140 -1225 17150 -1205
rect 17170 -1225 17180 -1205
rect 17140 -1235 17180 -1225
rect 17220 -1205 17260 -1195
rect 17220 -1225 17230 -1205
rect 17250 -1225 17260 -1205
rect 17220 -1235 17260 -1225
rect 17300 -1205 17340 -1195
rect 17300 -1225 17310 -1205
rect 17330 -1225 17340 -1205
rect 17300 -1235 17340 -1225
rect 17380 -1205 17420 -1195
rect 17380 -1225 17390 -1205
rect 17410 -1225 17420 -1205
rect 17380 -1235 17420 -1225
rect 17460 -1205 17500 -1195
rect 17460 -1225 17470 -1205
rect 17490 -1225 17500 -1205
rect 17460 -1235 17500 -1225
rect 17540 -1205 17580 -1195
rect 17540 -1225 17550 -1205
rect 17570 -1225 17580 -1205
rect 17540 -1235 17580 -1225
rect 17620 -1205 17660 -1195
rect 17620 -1225 17630 -1205
rect 17650 -1225 17660 -1205
rect 17620 -1235 17660 -1225
rect 17700 -1205 17740 -1195
rect 17700 -1225 17710 -1205
rect 17730 -1225 17740 -1205
rect 17700 -1235 17740 -1225
rect 17860 -1205 17900 -1195
rect 17860 -1225 17870 -1205
rect 17890 -1225 17900 -1205
rect 17860 -1235 17900 -1225
rect 17940 -1205 17980 -1195
rect 17940 -1225 17950 -1205
rect 17970 -1225 17980 -1205
rect 17940 -1235 17980 -1225
rect 18020 -1205 18060 -1195
rect 18020 -1225 18030 -1205
rect 18050 -1225 18060 -1205
rect 18020 -1235 18060 -1225
rect 18100 -1205 18140 -1195
rect 18100 -1225 18110 -1205
rect 18130 -1225 18140 -1205
rect 18100 -1235 18140 -1225
rect 18180 -1205 18220 -1195
rect 18180 -1225 18190 -1205
rect 18210 -1225 18220 -1205
rect 18180 -1235 18220 -1225
rect 18260 -1205 18300 -1195
rect 18260 -1225 18270 -1205
rect 18290 -1225 18300 -1205
rect 18260 -1235 18300 -1225
rect 18340 -1205 18380 -1195
rect 18340 -1225 18350 -1205
rect 18370 -1225 18380 -1205
rect 18340 -1235 18380 -1225
rect 18420 -1205 18460 -1195
rect 18420 -1225 18430 -1205
rect 18450 -1225 18460 -1205
rect 18420 -1235 18460 -1225
rect 18500 -1205 18540 -1195
rect 18500 -1225 18510 -1205
rect 18530 -1225 18540 -1205
rect 18500 -1235 18540 -1225
rect 18580 -1205 18620 -1195
rect 18580 -1225 18590 -1205
rect 18610 -1225 18620 -1205
rect 18580 -1235 18620 -1225
rect 18660 -1205 18700 -1195
rect 18660 -1225 18670 -1205
rect 18690 -1225 18700 -1205
rect 18660 -1235 18700 -1225
rect 18740 -1205 18780 -1195
rect 18740 -1225 18750 -1205
rect 18770 -1225 18780 -1205
rect 18740 -1235 18780 -1225
rect 16780 -1250 17780 -1235
rect 17820 -1250 18820 -1235
rect 16780 -1365 17780 -1350
rect 17820 -1365 18820 -1350
rect 16600 -1525 16640 -1515
rect 16600 -1545 16610 -1525
rect 16630 -1540 16640 -1525
rect 16770 -1525 16800 -1515
rect 16630 -1545 16655 -1540
rect 16770 -1545 16775 -1525
rect 16795 -1545 16800 -1525
rect 16880 -1525 16920 -1515
rect 16880 -1540 16890 -1525
rect 16860 -1545 16890 -1540
rect 16910 -1545 16920 -1525
rect 16600 -1555 16655 -1545
rect 16640 -1570 16655 -1555
rect 16695 -1560 16820 -1545
rect 16695 -1570 16710 -1560
rect 16750 -1570 16765 -1560
rect 16805 -1570 16820 -1560
rect 16860 -1555 16920 -1545
rect 17025 -1525 17065 -1515
rect 17025 -1545 17035 -1525
rect 17055 -1540 17065 -1525
rect 17305 -1525 17335 -1515
rect 17055 -1545 17080 -1540
rect 17305 -1545 17310 -1525
rect 17330 -1545 17335 -1525
rect 17465 -1525 17505 -1515
rect 17465 -1540 17475 -1525
rect 17450 -1545 17475 -1540
rect 17495 -1545 17505 -1525
rect 17025 -1555 17080 -1545
rect 16860 -1570 16875 -1555
rect 17065 -1570 17080 -1555
rect 17120 -1560 17410 -1545
rect 17120 -1570 17135 -1560
rect 17175 -1570 17190 -1560
rect 17230 -1570 17245 -1560
rect 17285 -1570 17300 -1560
rect 17340 -1570 17355 -1560
rect 17395 -1570 17410 -1560
rect 17450 -1555 17505 -1545
rect 17615 -1525 17655 -1515
rect 17615 -1545 17625 -1525
rect 17645 -1540 17655 -1525
rect 17785 -1525 17815 -1515
rect 17645 -1545 17670 -1540
rect 17785 -1545 17790 -1525
rect 17810 -1545 17815 -1525
rect 18005 -1525 18045 -1515
rect 18005 -1540 18015 -1525
rect 17985 -1545 18015 -1540
rect 18035 -1545 18045 -1525
rect 17615 -1555 17670 -1545
rect 17450 -1570 17465 -1555
rect 17655 -1570 17670 -1555
rect 17710 -1560 17945 -1545
rect 17710 -1570 17725 -1560
rect 17765 -1570 17780 -1560
rect 17820 -1570 17835 -1560
rect 17875 -1570 17890 -1560
rect 17930 -1570 17945 -1560
rect 17985 -1555 18045 -1545
rect 18150 -1525 18190 -1515
rect 18150 -1545 18160 -1525
rect 18180 -1540 18190 -1525
rect 18320 -1525 18350 -1515
rect 18180 -1545 18205 -1540
rect 18320 -1545 18325 -1525
rect 18345 -1545 18350 -1525
rect 18590 -1525 18630 -1515
rect 18590 -1540 18600 -1525
rect 18575 -1545 18600 -1540
rect 18620 -1545 18630 -1525
rect 18150 -1555 18205 -1545
rect 17985 -1570 18000 -1555
rect 18190 -1570 18205 -1555
rect 18245 -1560 18535 -1545
rect 18245 -1570 18260 -1560
rect 18300 -1570 18315 -1560
rect 18355 -1570 18370 -1560
rect 18410 -1570 18425 -1560
rect 18465 -1570 18480 -1560
rect 18520 -1570 18535 -1560
rect 18575 -1555 18630 -1545
rect 18575 -1570 18590 -1555
rect 16640 -1685 16655 -1670
rect 16695 -1685 16710 -1670
rect 16750 -1685 16765 -1670
rect 16805 -1685 16820 -1670
rect 16860 -1685 16875 -1670
rect 17065 -1685 17080 -1670
rect 17120 -1685 17135 -1670
rect 17175 -1685 17190 -1670
rect 17230 -1685 17245 -1670
rect 17285 -1685 17300 -1670
rect 17340 -1685 17355 -1670
rect 17395 -1685 17410 -1670
rect 17450 -1685 17465 -1670
rect 17655 -1685 17670 -1670
rect 17710 -1685 17725 -1670
rect 17765 -1685 17780 -1670
rect 17820 -1685 17835 -1670
rect 17875 -1685 17890 -1670
rect 17930 -1685 17945 -1670
rect 17985 -1685 18000 -1670
rect 18190 -1685 18205 -1670
rect 18245 -1685 18260 -1670
rect 18300 -1685 18315 -1670
rect 18355 -1685 18370 -1670
rect 18410 -1685 18425 -1670
rect 18465 -1685 18480 -1670
rect 18520 -1685 18535 -1670
rect 18575 -1685 18590 -1670
<< polycont >>
rect 16495 1435 16515 1455
rect 17790 1435 17810 1455
rect 16375 1300 16395 1320
rect 16615 1300 16635 1320
rect 16895 1300 16915 1320
rect 17060 1300 17080 1320
rect 17225 1300 17245 1320
rect 17505 1300 17525 1320
rect 18075 1300 18095 1320
rect 18355 1300 18375 1320
rect 18520 1300 18540 1320
rect 18685 1300 18705 1320
rect 16980 940 17000 960
rect 18600 940 18620 960
rect 18915 940 18935 960
rect 19085 940 19105 960
rect 16445 840 16465 860
rect 16665 840 16685 860
rect 16555 670 16575 690
rect 19010 610 19030 630
rect 17115 570 17135 590
rect 17205 570 17225 590
rect 17295 570 17315 590
rect 17385 570 17405 590
rect 17475 570 17495 590
rect 17565 570 17585 590
rect 17655 570 17675 590
rect 17745 570 17765 590
rect 17835 570 17855 590
rect 17925 570 17945 590
rect 18015 570 18035 590
rect 18105 570 18125 590
rect 18195 570 18215 590
rect 18285 570 18305 590
rect 18375 570 18395 590
rect 18465 570 18485 590
rect 16430 160 16450 180
rect 17630 160 17650 180
rect 17950 160 17970 180
rect 19150 160 19170 180
rect 16520 -15 16540 5
rect 16610 -10 16630 10
rect 16850 -10 16870 10
rect 16970 -10 16990 10
rect 17210 -10 17230 10
rect 17330 -10 17350 10
rect 17540 -10 17560 10
rect 18040 -10 18060 10
rect 18250 -10 18270 10
rect 18370 -10 18390 10
rect 18610 -10 18630 10
rect 18730 -10 18750 10
rect 18970 -10 18990 10
rect 19060 -15 19080 5
rect 17012 -205 17032 -185
rect 18568 -205 18588 -185
rect 17080 -525 17100 -505
rect 18445 -525 18465 -505
rect 16630 -770 16650 -750
rect 16750 -770 16770 -750
rect 16870 -770 16890 -750
rect 16990 -770 17010 -750
rect 17310 -770 17330 -750
rect 17430 -770 17450 -750
rect 17550 -770 17570 -750
rect 18030 -770 18050 -750
rect 18150 -770 18170 -750
rect 18270 -770 18290 -750
rect 18590 -770 18610 -750
rect 18710 -770 18730 -750
rect 18830 -770 18850 -750
rect 18950 -770 18970 -750
rect 16830 -1225 16850 -1205
rect 16910 -1225 16930 -1205
rect 16990 -1225 17010 -1205
rect 17070 -1225 17090 -1205
rect 17150 -1225 17170 -1205
rect 17230 -1225 17250 -1205
rect 17310 -1225 17330 -1205
rect 17390 -1225 17410 -1205
rect 17470 -1225 17490 -1205
rect 17550 -1225 17570 -1205
rect 17630 -1225 17650 -1205
rect 17710 -1225 17730 -1205
rect 17870 -1225 17890 -1205
rect 17950 -1225 17970 -1205
rect 18030 -1225 18050 -1205
rect 18110 -1225 18130 -1205
rect 18190 -1225 18210 -1205
rect 18270 -1225 18290 -1205
rect 18350 -1225 18370 -1205
rect 18430 -1225 18450 -1205
rect 18510 -1225 18530 -1205
rect 18590 -1225 18610 -1205
rect 18670 -1225 18690 -1205
rect 18750 -1225 18770 -1205
rect 16610 -1545 16630 -1525
rect 16775 -1545 16795 -1525
rect 16890 -1545 16910 -1525
rect 17035 -1545 17055 -1525
rect 17310 -1545 17330 -1525
rect 17475 -1545 17495 -1525
rect 17625 -1545 17645 -1525
rect 17790 -1545 17810 -1525
rect 18015 -1545 18035 -1525
rect 18160 -1545 18180 -1525
rect 18325 -1545 18345 -1525
rect 18600 -1545 18620 -1525
<< xpolycontact >>
rect 17470 -2035 17690 -2000
rect 17904 -2035 18124 -2000
rect 15950 -3376 15985 -3156
rect 15950 -3784 15985 -3565
rect 16160 -3285 16195 -3065
rect 16160 -3889 16195 -3669
rect 16220 -3285 16255 -3065
rect 16220 -3889 16255 -3669
rect 16280 -3285 16315 -3065
rect 16280 -3889 16315 -3669
rect 16485 -3160 16520 -2940
rect 16485 -3964 16520 -3744
rect 16545 -3160 16580 -2940
rect 16545 -3964 16580 -3744
rect 16605 -3160 16640 -2940
rect 16605 -3964 16640 -3744
rect 18960 -3160 18995 -2940
rect 18960 -3964 18995 -3744
rect 19020 -3160 19055 -2940
rect 19020 -3964 19055 -3744
rect 19080 -3160 19115 -2940
rect 19080 -3964 19115 -3744
rect 19285 -3257 19320 -3037
rect 19285 -3889 19320 -3669
rect 19345 -3257 19380 -3037
rect 19345 -3889 19380 -3669
rect 19405 -3257 19440 -3037
rect 19405 -3889 19440 -3669
rect 19610 -3376 19645 -3156
rect 19610 -3784 19645 -3565
<< ppolyres >>
rect 15950 -3565 15985 -3376
rect 19610 -3565 19645 -3376
<< xpolyres >>
rect 17690 -2035 17904 -2000
rect 16160 -3669 16195 -3285
rect 16220 -3669 16255 -3285
rect 16280 -3669 16315 -3285
rect 16485 -3744 16520 -3160
rect 16545 -3744 16580 -3160
rect 16605 -3744 16640 -3160
rect 18960 -3744 18995 -3160
rect 19020 -3744 19055 -3160
rect 19080 -3744 19115 -3160
rect 19285 -3669 19320 -3257
rect 19345 -3669 19380 -3257
rect 19405 -3669 19440 -3257
<< locali >>
rect 16485 1455 16525 1465
rect 16485 1435 16495 1455
rect 16515 1435 16525 1455
rect 16485 1425 16525 1435
rect 17780 1455 17820 1465
rect 17780 1435 17790 1455
rect 17810 1435 17820 1455
rect 17780 1425 17820 1435
rect 16365 1320 16405 1330
rect 16365 1300 16375 1320
rect 16395 1300 16405 1320
rect 16365 1290 16405 1300
rect 16485 1320 16525 1330
rect 16485 1300 16495 1320
rect 16515 1300 16525 1320
rect 16485 1290 16525 1300
rect 16605 1320 16645 1330
rect 16605 1300 16615 1320
rect 16635 1300 16645 1320
rect 16605 1290 16645 1300
rect 16885 1320 16925 1330
rect 16885 1300 16895 1320
rect 16915 1300 16925 1320
rect 16885 1290 16925 1300
rect 16945 1320 16975 1330
rect 16945 1300 16950 1320
rect 16970 1300 16975 1320
rect 16945 1290 16975 1300
rect 16995 1320 17035 1330
rect 16995 1300 17005 1320
rect 17025 1300 17035 1320
rect 16995 1290 17035 1300
rect 17055 1320 17085 1330
rect 17055 1300 17060 1320
rect 17080 1300 17085 1320
rect 17055 1290 17085 1300
rect 17105 1320 17145 1330
rect 17105 1300 17115 1320
rect 17135 1300 17145 1320
rect 17105 1290 17145 1300
rect 17215 1320 17255 1330
rect 17215 1300 17225 1320
rect 17245 1300 17255 1320
rect 17215 1290 17255 1300
rect 17495 1320 17535 1330
rect 17495 1300 17505 1320
rect 17525 1300 17535 1320
rect 17495 1290 17535 1300
rect 17560 1320 17600 1330
rect 17560 1300 17570 1320
rect 17590 1300 17600 1320
rect 17560 1290 17600 1300
rect 17620 1320 17650 1330
rect 17620 1300 17625 1320
rect 17645 1300 17650 1320
rect 16385 1270 16405 1290
rect 16495 1270 16515 1290
rect 16605 1270 16625 1290
rect 16895 1270 16915 1290
rect 16950 1270 16970 1290
rect 17005 1270 17025 1290
rect 17115 1270 17135 1290
rect 17225 1270 17245 1290
rect 17515 1270 17535 1290
rect 17570 1270 17590 1290
rect 16340 1262 16410 1270
rect 16340 1240 16345 1262
rect 16365 1260 16410 1262
rect 16365 1240 16385 1260
rect 16405 1240 16410 1260
rect 16340 1210 16410 1240
rect 16340 1190 16345 1210
rect 16365 1190 16385 1210
rect 16405 1190 16410 1210
rect 16340 1180 16410 1190
rect 16435 1260 16465 1270
rect 16435 1240 16440 1260
rect 16460 1240 16465 1260
rect 16435 1210 16465 1240
rect 16435 1190 16440 1210
rect 16460 1190 16465 1210
rect 16435 1180 16465 1190
rect 16490 1260 16520 1270
rect 16490 1240 16495 1260
rect 16515 1240 16520 1260
rect 16490 1210 16520 1240
rect 16490 1190 16495 1210
rect 16515 1190 16520 1210
rect 16490 1180 16520 1190
rect 16545 1260 16575 1270
rect 16545 1240 16550 1260
rect 16570 1240 16575 1260
rect 16545 1210 16575 1240
rect 16545 1190 16550 1210
rect 16570 1190 16575 1210
rect 16545 1180 16575 1190
rect 16600 1262 16670 1270
rect 16600 1260 16645 1262
rect 16600 1240 16605 1260
rect 16625 1240 16645 1260
rect 16665 1240 16670 1262
rect 16600 1210 16670 1240
rect 16600 1190 16605 1210
rect 16625 1190 16645 1210
rect 16665 1190 16670 1210
rect 16600 1180 16670 1190
rect 16850 1262 16920 1270
rect 16850 1190 16855 1262
rect 16875 1260 16920 1262
rect 16875 1190 16895 1260
rect 16850 1188 16895 1190
rect 16915 1188 16920 1260
rect 16850 1180 16920 1188
rect 16945 1260 16975 1270
rect 16945 1188 16950 1260
rect 16970 1188 16975 1260
rect 16945 1180 16975 1188
rect 17000 1260 17030 1270
rect 17000 1188 17005 1260
rect 17025 1188 17030 1260
rect 17000 1180 17030 1188
rect 17055 1260 17085 1270
rect 17055 1188 17060 1260
rect 17080 1188 17085 1260
rect 17055 1180 17085 1188
rect 17110 1260 17140 1270
rect 17110 1188 17115 1260
rect 17135 1188 17140 1260
rect 17110 1180 17140 1188
rect 17165 1260 17195 1270
rect 17165 1188 17170 1260
rect 17190 1188 17195 1260
rect 17165 1180 17195 1188
rect 17220 1262 17290 1270
rect 17220 1260 17265 1262
rect 17220 1188 17225 1260
rect 17245 1190 17265 1260
rect 17285 1190 17290 1262
rect 17245 1188 17290 1190
rect 17220 1180 17290 1188
rect 17470 1262 17540 1270
rect 17470 1240 17475 1262
rect 17495 1260 17540 1262
rect 17495 1240 17515 1260
rect 17535 1240 17540 1260
rect 17470 1210 17540 1240
rect 17470 1190 17475 1210
rect 17495 1190 17515 1210
rect 17535 1190 17540 1210
rect 17470 1180 17540 1190
rect 17565 1260 17595 1270
rect 17565 1240 17570 1260
rect 17590 1240 17595 1260
rect 17565 1210 17595 1240
rect 17565 1190 17570 1210
rect 17590 1190 17595 1210
rect 17565 1180 17595 1190
rect 17620 1260 17650 1300
rect 17670 1320 17710 1330
rect 17670 1300 17680 1320
rect 17700 1300 17710 1320
rect 17670 1290 17710 1300
rect 17730 1320 17760 1330
rect 17730 1300 17735 1320
rect 17755 1300 17760 1320
rect 17680 1270 17700 1290
rect 17620 1240 17625 1260
rect 17645 1240 17650 1260
rect 17620 1210 17650 1240
rect 17620 1190 17625 1210
rect 17645 1190 17650 1210
rect 17620 1180 17650 1190
rect 17675 1260 17705 1270
rect 17675 1240 17680 1260
rect 17700 1240 17705 1260
rect 17675 1210 17705 1240
rect 17675 1190 17680 1210
rect 17700 1190 17705 1210
rect 17675 1180 17705 1190
rect 17730 1260 17760 1300
rect 17780 1320 17820 1330
rect 17780 1300 17790 1320
rect 17810 1300 17820 1320
rect 17780 1290 17820 1300
rect 17840 1320 17870 1330
rect 17840 1300 17845 1320
rect 17865 1300 17870 1320
rect 17790 1270 17810 1290
rect 17730 1240 17735 1260
rect 17755 1240 17760 1260
rect 17730 1210 17760 1240
rect 17730 1190 17735 1210
rect 17755 1190 17760 1210
rect 17730 1180 17760 1190
rect 17785 1260 17815 1270
rect 17785 1240 17790 1260
rect 17810 1240 17815 1260
rect 17785 1210 17815 1240
rect 17785 1190 17790 1210
rect 17810 1190 17815 1210
rect 17785 1180 17815 1190
rect 17840 1260 17870 1300
rect 17890 1320 17930 1330
rect 17890 1300 17900 1320
rect 17920 1300 17930 1320
rect 17890 1290 17930 1300
rect 17950 1320 17980 1330
rect 17950 1300 17955 1320
rect 17975 1300 17980 1320
rect 17900 1270 17920 1290
rect 17840 1240 17845 1260
rect 17865 1240 17870 1260
rect 17840 1210 17870 1240
rect 17840 1190 17845 1210
rect 17865 1190 17870 1210
rect 17840 1180 17870 1190
rect 17895 1260 17925 1270
rect 17895 1240 17900 1260
rect 17920 1240 17925 1260
rect 17895 1210 17925 1240
rect 17895 1190 17900 1210
rect 17920 1190 17925 1210
rect 17895 1180 17925 1190
rect 17950 1260 17980 1300
rect 18000 1320 18040 1330
rect 18000 1300 18010 1320
rect 18030 1300 18040 1320
rect 18000 1290 18040 1300
rect 18065 1320 18105 1330
rect 18065 1300 18075 1320
rect 18095 1300 18105 1320
rect 18065 1290 18105 1300
rect 18345 1320 18385 1330
rect 18345 1300 18355 1320
rect 18375 1300 18385 1320
rect 18345 1290 18385 1300
rect 18455 1320 18495 1330
rect 18455 1300 18465 1320
rect 18485 1300 18495 1320
rect 18455 1290 18495 1300
rect 18515 1320 18545 1330
rect 18515 1300 18520 1320
rect 18540 1300 18545 1320
rect 18515 1290 18545 1300
rect 18565 1320 18605 1330
rect 18565 1300 18575 1320
rect 18595 1300 18605 1320
rect 18565 1290 18605 1300
rect 18625 1320 18655 1330
rect 18625 1300 18630 1320
rect 18650 1300 18655 1320
rect 18625 1290 18655 1300
rect 18675 1320 18715 1330
rect 18675 1300 18685 1320
rect 18705 1300 18715 1320
rect 18675 1290 18715 1300
rect 18010 1270 18030 1290
rect 18065 1270 18085 1290
rect 18355 1270 18375 1290
rect 18465 1270 18485 1290
rect 18575 1270 18595 1290
rect 18630 1270 18650 1290
rect 18685 1270 18705 1290
rect 17950 1240 17955 1260
rect 17975 1240 17980 1260
rect 17950 1210 17980 1240
rect 17950 1190 17955 1210
rect 17975 1190 17980 1210
rect 17950 1180 17980 1190
rect 18005 1260 18035 1270
rect 18005 1240 18010 1260
rect 18030 1240 18035 1260
rect 18005 1210 18035 1240
rect 18005 1190 18010 1210
rect 18030 1190 18035 1210
rect 18005 1180 18035 1190
rect 18060 1262 18130 1270
rect 18060 1260 18105 1262
rect 18060 1240 18065 1260
rect 18085 1240 18105 1260
rect 18125 1240 18130 1262
rect 18060 1210 18130 1240
rect 18060 1190 18065 1210
rect 18085 1190 18105 1210
rect 18125 1190 18130 1210
rect 18060 1180 18130 1190
rect 18310 1262 18380 1270
rect 18310 1190 18315 1262
rect 18335 1260 18380 1262
rect 18335 1190 18355 1260
rect 18375 1190 18380 1260
rect 18310 1180 18380 1190
rect 18405 1260 18435 1270
rect 18405 1190 18410 1260
rect 18430 1190 18435 1260
rect 18405 1180 18435 1190
rect 18460 1260 18490 1270
rect 18460 1190 18465 1260
rect 18485 1190 18490 1260
rect 18460 1180 18490 1190
rect 18515 1260 18545 1270
rect 18515 1190 18520 1260
rect 18540 1190 18545 1260
rect 18515 1180 18545 1190
rect 18570 1260 18600 1270
rect 18570 1190 18575 1260
rect 18595 1190 18600 1260
rect 18570 1180 18600 1190
rect 18625 1260 18655 1270
rect 18625 1190 18630 1260
rect 18650 1190 18655 1260
rect 18625 1180 18655 1190
rect 18680 1262 18750 1270
rect 18680 1260 18725 1262
rect 18680 1190 18685 1260
rect 18705 1190 18725 1260
rect 18745 1190 18750 1262
rect 18680 1180 18750 1190
rect 16440 1160 16460 1180
rect 16550 1160 16570 1180
rect 16950 1160 16970 1180
rect 17060 1160 17080 1180
rect 17170 1160 17190 1180
rect 17625 1160 17645 1180
rect 17735 1160 17755 1180
rect 17845 1160 17865 1180
rect 17955 1160 17975 1180
rect 18410 1160 18430 1180
rect 18520 1160 18540 1180
rect 18630 1160 18650 1180
rect 16430 1150 16470 1160
rect 16430 1130 16440 1150
rect 16460 1130 16470 1150
rect 16430 1120 16470 1130
rect 16540 1150 16580 1160
rect 16540 1130 16550 1150
rect 16570 1130 16580 1150
rect 16540 1120 16580 1130
rect 16940 1150 16980 1160
rect 16940 1130 16950 1150
rect 16970 1130 16980 1150
rect 16940 1120 16980 1130
rect 17050 1150 17090 1160
rect 17050 1130 17060 1150
rect 17080 1130 17090 1150
rect 17050 1120 17090 1130
rect 17160 1150 17200 1160
rect 17160 1130 17170 1150
rect 17190 1130 17200 1150
rect 17160 1120 17200 1130
rect 17615 1150 17655 1160
rect 17615 1130 17625 1150
rect 17645 1130 17655 1150
rect 17615 1120 17655 1130
rect 17725 1150 17765 1160
rect 17725 1130 17735 1150
rect 17755 1130 17765 1150
rect 17725 1120 17765 1130
rect 17835 1150 17875 1160
rect 17835 1130 17845 1150
rect 17865 1130 17875 1150
rect 17835 1120 17875 1130
rect 17945 1150 17985 1160
rect 17945 1130 17955 1150
rect 17975 1130 17985 1150
rect 17945 1120 17985 1130
rect 18400 1150 18440 1160
rect 18400 1130 18410 1150
rect 18430 1130 18440 1150
rect 18400 1120 18440 1130
rect 18510 1150 18550 1160
rect 18510 1130 18520 1150
rect 18540 1130 18550 1150
rect 18510 1120 18550 1130
rect 18620 1150 18660 1160
rect 18620 1130 18630 1150
rect 18650 1130 18660 1150
rect 18620 1120 18660 1130
rect 16970 960 17010 970
rect 16970 940 16980 960
rect 17000 940 17010 960
rect 16970 930 17010 940
rect 17150 960 17190 970
rect 17150 940 17160 960
rect 17180 940 17190 960
rect 17150 930 17190 940
rect 17330 960 17370 970
rect 17330 940 17340 960
rect 17360 940 17370 960
rect 17330 930 17370 940
rect 17510 960 17550 970
rect 17510 940 17520 960
rect 17540 940 17550 960
rect 17510 930 17550 940
rect 17690 960 17730 970
rect 17690 940 17700 960
rect 17720 940 17730 960
rect 17690 930 17730 940
rect 17870 960 17910 970
rect 17870 940 17880 960
rect 17900 940 17910 960
rect 17870 930 17910 940
rect 18050 960 18090 970
rect 18050 940 18060 960
rect 18080 940 18090 960
rect 18050 930 18090 940
rect 18230 960 18270 970
rect 18230 940 18240 960
rect 18260 940 18270 960
rect 18230 930 18270 940
rect 18410 960 18450 970
rect 18410 940 18420 960
rect 18440 940 18450 960
rect 18410 930 18450 940
rect 18590 960 18630 970
rect 18590 940 18600 960
rect 18620 940 18630 960
rect 18590 930 18630 940
rect 18905 960 18945 970
rect 18905 940 18915 960
rect 18935 940 18945 960
rect 18905 930 18945 940
rect 19015 960 19055 970
rect 19015 940 19025 960
rect 19045 940 19055 960
rect 19015 930 19055 940
rect 19075 960 19115 970
rect 19075 940 19085 960
rect 19105 940 19115 960
rect 19075 930 19115 940
rect 16980 910 17000 930
rect 17160 910 17180 930
rect 17340 910 17360 930
rect 17520 910 17540 930
rect 17700 910 17720 930
rect 17880 910 17900 930
rect 18060 910 18080 930
rect 18240 910 18260 930
rect 18420 910 18440 930
rect 18600 910 18620 930
rect 16935 900 17005 910
rect 16935 880 16940 900
rect 16960 880 16980 900
rect 17000 880 17005 900
rect 16440 860 16470 870
rect 16440 840 16445 860
rect 16465 840 16470 860
rect 16440 810 16470 840
rect 16545 860 16585 870
rect 16545 840 16555 860
rect 16575 840 16585 860
rect 16545 830 16585 840
rect 16655 860 16695 870
rect 16655 840 16665 860
rect 16685 840 16695 860
rect 16655 830 16695 840
rect 16935 850 17005 880
rect 16935 830 16940 850
rect 16960 830 16980 850
rect 17000 830 17005 850
rect 16555 810 16575 830
rect 16660 810 16690 830
rect 16400 800 16470 810
rect 16400 780 16405 800
rect 16425 780 16445 800
rect 16465 780 16470 800
rect 16400 750 16470 780
rect 16400 730 16405 750
rect 16425 730 16445 750
rect 16465 730 16470 750
rect 16400 720 16470 730
rect 16495 800 16525 810
rect 16495 780 16500 800
rect 16520 780 16525 800
rect 16495 750 16525 780
rect 16495 730 16500 750
rect 16520 730 16525 750
rect 16495 720 16525 730
rect 16550 800 16580 810
rect 16550 780 16555 800
rect 16575 780 16580 800
rect 16550 750 16580 780
rect 16550 730 16555 750
rect 16575 730 16580 750
rect 16550 720 16580 730
rect 16605 800 16635 810
rect 16605 780 16610 800
rect 16630 780 16635 800
rect 16605 750 16635 780
rect 16605 730 16610 750
rect 16630 730 16635 750
rect 16605 720 16635 730
rect 16660 800 16735 810
rect 16660 780 16665 800
rect 16685 780 16710 800
rect 16730 780 16735 800
rect 16660 750 16735 780
rect 16660 730 16665 750
rect 16685 730 16710 750
rect 16730 730 16735 750
rect 16660 720 16735 730
rect 16935 800 17005 830
rect 16935 780 16940 800
rect 16960 780 16980 800
rect 17000 780 17005 800
rect 16935 750 17005 780
rect 16935 730 16940 750
rect 16960 730 16980 750
rect 17000 730 17005 750
rect 16500 700 16520 720
rect 16610 700 16630 720
rect 16935 700 17005 730
rect 16480 690 16520 700
rect 16480 670 16490 690
rect 16510 670 16520 690
rect 16480 660 16520 670
rect 16545 690 16585 700
rect 16545 670 16555 690
rect 16575 670 16585 690
rect 16545 660 16585 670
rect 16610 690 16650 700
rect 16610 670 16620 690
rect 16640 670 16650 690
rect 16610 660 16650 670
rect 16935 680 16940 700
rect 16960 680 16980 700
rect 17000 680 17005 700
rect 16935 650 17005 680
rect 16935 630 16940 650
rect 16960 630 16980 650
rect 17000 630 17005 650
rect 16935 620 17005 630
rect 17065 900 17095 910
rect 17065 880 17070 900
rect 17090 880 17095 900
rect 17065 850 17095 880
rect 17065 830 17070 850
rect 17090 830 17095 850
rect 17065 800 17095 830
rect 17065 780 17070 800
rect 17090 780 17095 800
rect 17065 750 17095 780
rect 17065 730 17070 750
rect 17090 730 17095 750
rect 17065 700 17095 730
rect 17065 680 17070 700
rect 17090 680 17095 700
rect 17065 650 17095 680
rect 17065 630 17070 650
rect 17090 630 17095 650
rect 17065 620 17095 630
rect 17155 900 17185 910
rect 17155 880 17160 900
rect 17180 880 17185 900
rect 17155 850 17185 880
rect 17155 830 17160 850
rect 17180 830 17185 850
rect 17155 800 17185 830
rect 17155 780 17160 800
rect 17180 780 17185 800
rect 17155 750 17185 780
rect 17155 730 17160 750
rect 17180 730 17185 750
rect 17155 700 17185 730
rect 17155 680 17160 700
rect 17180 680 17185 700
rect 17155 650 17185 680
rect 17155 630 17160 650
rect 17180 630 17185 650
rect 17155 620 17185 630
rect 17245 900 17275 910
rect 17245 880 17250 900
rect 17270 880 17275 900
rect 17245 850 17275 880
rect 17245 830 17250 850
rect 17270 830 17275 850
rect 17245 800 17275 830
rect 17245 780 17250 800
rect 17270 780 17275 800
rect 17245 750 17275 780
rect 17245 730 17250 750
rect 17270 730 17275 750
rect 17245 700 17275 730
rect 17245 680 17250 700
rect 17270 680 17275 700
rect 17245 650 17275 680
rect 17245 630 17250 650
rect 17270 630 17275 650
rect 17245 620 17275 630
rect 17335 900 17365 910
rect 17335 880 17340 900
rect 17360 880 17365 900
rect 17335 850 17365 880
rect 17335 830 17340 850
rect 17360 830 17365 850
rect 17335 800 17365 830
rect 17335 780 17340 800
rect 17360 780 17365 800
rect 17335 750 17365 780
rect 17335 730 17340 750
rect 17360 730 17365 750
rect 17335 700 17365 730
rect 17335 680 17340 700
rect 17360 680 17365 700
rect 17335 650 17365 680
rect 17335 630 17340 650
rect 17360 630 17365 650
rect 17335 620 17365 630
rect 17425 900 17455 910
rect 17425 880 17430 900
rect 17450 880 17455 900
rect 17425 850 17455 880
rect 17425 830 17430 850
rect 17450 830 17455 850
rect 17425 800 17455 830
rect 17425 780 17430 800
rect 17450 780 17455 800
rect 17425 750 17455 780
rect 17425 730 17430 750
rect 17450 730 17455 750
rect 17425 700 17455 730
rect 17425 680 17430 700
rect 17450 680 17455 700
rect 17425 650 17455 680
rect 17425 630 17430 650
rect 17450 630 17455 650
rect 17425 620 17455 630
rect 17515 900 17545 910
rect 17515 880 17520 900
rect 17540 880 17545 900
rect 17515 850 17545 880
rect 17515 830 17520 850
rect 17540 830 17545 850
rect 17515 800 17545 830
rect 17515 780 17520 800
rect 17540 780 17545 800
rect 17515 750 17545 780
rect 17515 730 17520 750
rect 17540 730 17545 750
rect 17515 700 17545 730
rect 17515 680 17520 700
rect 17540 680 17545 700
rect 17515 650 17545 680
rect 17515 630 17520 650
rect 17540 630 17545 650
rect 17515 620 17545 630
rect 17605 900 17635 910
rect 17605 880 17610 900
rect 17630 880 17635 900
rect 17605 850 17635 880
rect 17605 830 17610 850
rect 17630 830 17635 850
rect 17605 800 17635 830
rect 17605 780 17610 800
rect 17630 780 17635 800
rect 17605 750 17635 780
rect 17605 730 17610 750
rect 17630 730 17635 750
rect 17605 700 17635 730
rect 17605 680 17610 700
rect 17630 680 17635 700
rect 17605 650 17635 680
rect 17605 630 17610 650
rect 17630 630 17635 650
rect 17605 620 17635 630
rect 17695 900 17725 910
rect 17695 880 17700 900
rect 17720 880 17725 900
rect 17695 850 17725 880
rect 17695 830 17700 850
rect 17720 830 17725 850
rect 17695 800 17725 830
rect 17695 780 17700 800
rect 17720 780 17725 800
rect 17695 750 17725 780
rect 17695 730 17700 750
rect 17720 730 17725 750
rect 17695 700 17725 730
rect 17695 680 17700 700
rect 17720 680 17725 700
rect 17695 650 17725 680
rect 17695 630 17700 650
rect 17720 630 17725 650
rect 17695 620 17725 630
rect 17785 900 17815 910
rect 17785 880 17790 900
rect 17810 880 17815 900
rect 17785 850 17815 880
rect 17785 830 17790 850
rect 17810 830 17815 850
rect 17785 800 17815 830
rect 17785 780 17790 800
rect 17810 780 17815 800
rect 17785 750 17815 780
rect 17785 730 17790 750
rect 17810 730 17815 750
rect 17785 700 17815 730
rect 17785 680 17790 700
rect 17810 680 17815 700
rect 17785 650 17815 680
rect 17785 630 17790 650
rect 17810 630 17815 650
rect 17785 620 17815 630
rect 17875 900 17905 910
rect 17875 880 17880 900
rect 17900 880 17905 900
rect 17875 850 17905 880
rect 17875 830 17880 850
rect 17900 830 17905 850
rect 17875 800 17905 830
rect 17875 780 17880 800
rect 17900 780 17905 800
rect 17875 750 17905 780
rect 17875 730 17880 750
rect 17900 730 17905 750
rect 17875 700 17905 730
rect 17875 680 17880 700
rect 17900 680 17905 700
rect 17875 650 17905 680
rect 17875 630 17880 650
rect 17900 630 17905 650
rect 17875 620 17905 630
rect 17965 900 17995 910
rect 17965 880 17970 900
rect 17990 880 17995 900
rect 17965 850 17995 880
rect 17965 830 17970 850
rect 17990 830 17995 850
rect 17965 800 17995 830
rect 17965 780 17970 800
rect 17990 780 17995 800
rect 17965 750 17995 780
rect 17965 730 17970 750
rect 17990 730 17995 750
rect 17965 700 17995 730
rect 17965 680 17970 700
rect 17990 680 17995 700
rect 17965 650 17995 680
rect 17965 630 17970 650
rect 17990 630 17995 650
rect 17965 620 17995 630
rect 18055 900 18085 910
rect 18055 880 18060 900
rect 18080 880 18085 900
rect 18055 850 18085 880
rect 18055 830 18060 850
rect 18080 830 18085 850
rect 18055 800 18085 830
rect 18055 780 18060 800
rect 18080 780 18085 800
rect 18055 750 18085 780
rect 18055 730 18060 750
rect 18080 730 18085 750
rect 18055 700 18085 730
rect 18055 680 18060 700
rect 18080 680 18085 700
rect 18055 650 18085 680
rect 18055 630 18060 650
rect 18080 630 18085 650
rect 18055 620 18085 630
rect 18145 900 18175 910
rect 18145 880 18150 900
rect 18170 880 18175 900
rect 18145 850 18175 880
rect 18145 830 18150 850
rect 18170 830 18175 850
rect 18145 800 18175 830
rect 18145 780 18150 800
rect 18170 780 18175 800
rect 18145 750 18175 780
rect 18145 730 18150 750
rect 18170 730 18175 750
rect 18145 700 18175 730
rect 18145 680 18150 700
rect 18170 680 18175 700
rect 18145 650 18175 680
rect 18145 630 18150 650
rect 18170 630 18175 650
rect 18145 620 18175 630
rect 18235 900 18265 910
rect 18235 880 18240 900
rect 18260 880 18265 900
rect 18235 850 18265 880
rect 18235 830 18240 850
rect 18260 830 18265 850
rect 18235 800 18265 830
rect 18235 780 18240 800
rect 18260 780 18265 800
rect 18235 750 18265 780
rect 18235 730 18240 750
rect 18260 730 18265 750
rect 18235 700 18265 730
rect 18235 680 18240 700
rect 18260 680 18265 700
rect 18235 650 18265 680
rect 18235 630 18240 650
rect 18260 630 18265 650
rect 18235 620 18265 630
rect 18325 900 18355 910
rect 18325 880 18330 900
rect 18350 880 18355 900
rect 18325 850 18355 880
rect 18325 830 18330 850
rect 18350 830 18355 850
rect 18325 800 18355 830
rect 18325 780 18330 800
rect 18350 780 18355 800
rect 18325 750 18355 780
rect 18325 730 18330 750
rect 18350 730 18355 750
rect 18325 700 18355 730
rect 18325 680 18330 700
rect 18350 680 18355 700
rect 18325 650 18355 680
rect 18325 630 18330 650
rect 18350 630 18355 650
rect 18325 620 18355 630
rect 18415 900 18445 910
rect 18415 880 18420 900
rect 18440 880 18445 900
rect 18415 850 18445 880
rect 18415 830 18420 850
rect 18440 830 18445 850
rect 18415 800 18445 830
rect 18415 780 18420 800
rect 18440 780 18445 800
rect 18415 750 18445 780
rect 18415 730 18420 750
rect 18440 730 18445 750
rect 18415 700 18445 730
rect 18415 680 18420 700
rect 18440 680 18445 700
rect 18415 650 18445 680
rect 18415 630 18420 650
rect 18440 630 18445 650
rect 18415 620 18445 630
rect 18505 900 18535 910
rect 18505 880 18510 900
rect 18530 880 18535 900
rect 18505 850 18535 880
rect 18505 830 18510 850
rect 18530 830 18535 850
rect 18505 800 18535 830
rect 18505 780 18510 800
rect 18530 780 18535 800
rect 18505 750 18535 780
rect 18505 730 18510 750
rect 18530 730 18535 750
rect 18505 700 18535 730
rect 18505 680 18510 700
rect 18530 680 18535 700
rect 18505 650 18535 680
rect 18505 630 18510 650
rect 18530 630 18535 650
rect 18505 620 18535 630
rect 18595 900 18665 910
rect 18595 880 18600 900
rect 18620 880 18640 900
rect 18660 880 18665 900
rect 18595 850 18665 880
rect 18595 830 18600 850
rect 18620 830 18640 850
rect 18660 830 18665 850
rect 18595 800 18665 830
rect 18595 780 18600 800
rect 18620 780 18640 800
rect 18660 780 18665 800
rect 18595 750 18665 780
rect 18595 730 18600 750
rect 18620 730 18640 750
rect 18660 730 18665 750
rect 18595 700 18665 730
rect 18870 900 18940 910
rect 18870 880 18875 900
rect 18895 880 18915 900
rect 18935 880 18940 900
rect 18870 850 18940 880
rect 18870 830 18875 850
rect 18895 830 18915 850
rect 18935 830 18940 850
rect 18870 800 18940 830
rect 18870 780 18875 800
rect 18895 780 18915 800
rect 18935 780 18940 800
rect 18870 750 18940 780
rect 18870 730 18875 750
rect 18895 730 18915 750
rect 18935 730 18940 750
rect 18870 720 18940 730
rect 18965 900 18995 910
rect 18965 880 18970 900
rect 18990 880 18995 900
rect 18965 850 18995 880
rect 18965 830 18970 850
rect 18990 830 18995 850
rect 18965 800 18995 830
rect 18965 780 18970 800
rect 18990 780 18995 800
rect 18965 750 18995 780
rect 18965 730 18970 750
rect 18990 730 18995 750
rect 18965 720 18995 730
rect 19020 900 19050 910
rect 19020 880 19025 900
rect 19045 880 19050 900
rect 19020 850 19050 880
rect 19020 830 19025 850
rect 19045 830 19050 850
rect 19020 800 19050 830
rect 19020 780 19025 800
rect 19045 780 19050 800
rect 19020 750 19050 780
rect 19020 730 19025 750
rect 19045 730 19050 750
rect 19020 720 19050 730
rect 19075 900 19145 910
rect 19075 880 19080 900
rect 19100 880 19120 900
rect 19140 880 19145 900
rect 19075 850 19145 880
rect 19075 830 19080 850
rect 19100 830 19120 850
rect 19140 830 19145 850
rect 19075 800 19145 830
rect 19075 780 19080 800
rect 19100 780 19120 800
rect 19140 780 19145 800
rect 19075 750 19145 780
rect 19075 730 19080 750
rect 19100 730 19120 750
rect 19140 730 19145 750
rect 19075 720 19145 730
rect 18595 680 18600 700
rect 18620 680 18640 700
rect 18660 680 18665 700
rect 18595 650 18665 680
rect 18595 630 18600 650
rect 18620 630 18640 650
rect 18660 630 18665 650
rect 18595 620 18665 630
rect 19000 630 19040 640
rect 19000 610 19010 630
rect 19030 610 19040 630
rect 19000 600 19040 610
rect 17110 590 17145 600
rect 17110 570 17115 590
rect 17135 570 17145 590
rect 17110 560 17145 570
rect 17195 590 17235 600
rect 17195 570 17205 590
rect 17225 570 17235 590
rect 17195 560 17235 570
rect 17285 590 17325 600
rect 17285 570 17295 590
rect 17315 570 17325 590
rect 17285 560 17325 570
rect 17375 590 17415 600
rect 17375 570 17385 590
rect 17405 570 17415 590
rect 17375 560 17415 570
rect 17465 590 17505 600
rect 17465 570 17475 590
rect 17495 570 17505 590
rect 17465 560 17505 570
rect 17555 590 17595 600
rect 17555 570 17565 590
rect 17585 570 17595 590
rect 17555 560 17595 570
rect 17645 590 17685 600
rect 17645 570 17655 590
rect 17675 570 17685 590
rect 17645 560 17685 570
rect 17735 590 17770 600
rect 17735 570 17745 590
rect 17765 570 17770 590
rect 17735 560 17770 570
rect 17830 590 17865 600
rect 17830 570 17835 590
rect 17855 570 17865 590
rect 17830 560 17865 570
rect 17915 590 17955 600
rect 17915 570 17925 590
rect 17945 570 17955 590
rect 17915 560 17955 570
rect 18005 590 18045 600
rect 18005 570 18015 590
rect 18035 570 18045 590
rect 18005 560 18045 570
rect 18095 590 18135 600
rect 18095 570 18105 590
rect 18125 570 18135 590
rect 18095 560 18135 570
rect 18185 590 18225 600
rect 18185 570 18195 590
rect 18215 570 18225 590
rect 18185 560 18225 570
rect 18275 590 18315 600
rect 18275 570 18285 590
rect 18305 570 18315 590
rect 18275 560 18315 570
rect 18365 590 18405 600
rect 18365 570 18375 590
rect 18395 570 18405 590
rect 18365 560 18405 570
rect 18455 590 18490 600
rect 18455 570 18465 590
rect 18485 570 18490 590
rect 18455 560 18490 570
rect 16425 180 16455 190
rect 16425 160 16430 180
rect 16450 160 16455 180
rect 16425 150 16455 160
rect 17625 180 17655 190
rect 17625 160 17630 180
rect 17650 160 17655 180
rect 17625 150 17655 160
rect 17945 180 17975 190
rect 17945 160 17950 180
rect 17970 160 17975 180
rect 17945 150 17975 160
rect 19145 180 19175 190
rect 19145 160 19150 180
rect 19170 160 19175 180
rect 19145 150 19175 160
rect 16385 120 16455 130
rect 16385 100 16390 120
rect 16410 100 16430 120
rect 16450 100 16455 120
rect 16385 70 16455 100
rect 16385 50 16390 70
rect 16410 50 16430 70
rect 16450 50 16455 70
rect 16385 40 16455 50
rect 16485 120 16515 130
rect 16485 100 16490 120
rect 16510 100 16515 120
rect 16485 70 16515 100
rect 16485 50 16490 70
rect 16510 50 16515 70
rect 16485 40 16515 50
rect 16545 120 16575 130
rect 16545 100 16550 120
rect 16570 100 16575 120
rect 16545 70 16575 100
rect 16545 50 16550 70
rect 16570 50 16575 70
rect 16545 40 16575 50
rect 16605 120 16635 130
rect 16605 100 16610 120
rect 16630 100 16635 120
rect 16605 70 16635 100
rect 16605 50 16610 70
rect 16630 50 16635 70
rect 16605 40 16635 50
rect 16665 120 16695 130
rect 16665 100 16670 120
rect 16690 100 16695 120
rect 16665 70 16695 100
rect 16665 50 16670 70
rect 16690 50 16695 70
rect 16665 40 16695 50
rect 16725 120 16755 130
rect 16725 100 16730 120
rect 16750 100 16755 120
rect 16725 70 16755 100
rect 16725 50 16730 70
rect 16750 50 16755 70
rect 16725 40 16755 50
rect 16785 120 16815 130
rect 16785 100 16790 120
rect 16810 100 16815 120
rect 16785 70 16815 100
rect 16785 50 16790 70
rect 16810 50 16815 70
rect 16785 40 16815 50
rect 16845 120 16875 130
rect 16845 100 16850 120
rect 16870 100 16875 120
rect 16845 70 16875 100
rect 16845 50 16850 70
rect 16870 50 16875 70
rect 16845 40 16875 50
rect 16905 120 16935 130
rect 16905 100 16910 120
rect 16930 100 16935 120
rect 16905 70 16935 100
rect 16905 50 16910 70
rect 16930 50 16935 70
rect 16905 40 16935 50
rect 16965 120 16995 130
rect 16965 100 16970 120
rect 16990 100 16995 120
rect 16965 70 16995 100
rect 16965 50 16970 70
rect 16990 50 16995 70
rect 16965 40 16995 50
rect 17025 120 17055 130
rect 17025 100 17030 120
rect 17050 100 17055 120
rect 17025 70 17055 100
rect 17025 50 17030 70
rect 17050 50 17055 70
rect 17025 40 17055 50
rect 17085 120 17115 130
rect 17085 100 17090 120
rect 17110 100 17115 120
rect 17085 70 17115 100
rect 17085 50 17090 70
rect 17110 50 17115 70
rect 17085 40 17115 50
rect 17145 120 17175 130
rect 17145 100 17150 120
rect 17170 100 17175 120
rect 17145 70 17175 100
rect 17145 50 17150 70
rect 17170 50 17175 70
rect 17145 40 17175 50
rect 17205 120 17235 130
rect 17205 100 17210 120
rect 17230 100 17235 120
rect 17205 70 17235 100
rect 17205 50 17210 70
rect 17230 50 17235 70
rect 17205 40 17235 50
rect 17265 120 17295 130
rect 17265 100 17270 120
rect 17290 100 17295 120
rect 17265 70 17295 100
rect 17265 50 17270 70
rect 17290 50 17295 70
rect 17265 40 17295 50
rect 17325 120 17355 130
rect 17325 100 17330 120
rect 17350 100 17355 120
rect 17325 70 17355 100
rect 17325 50 17330 70
rect 17350 50 17355 70
rect 17325 40 17355 50
rect 17385 120 17415 130
rect 17385 100 17390 120
rect 17410 100 17415 120
rect 17385 70 17415 100
rect 17385 50 17390 70
rect 17410 50 17415 70
rect 17385 40 17415 50
rect 17445 120 17475 130
rect 17445 100 17450 120
rect 17470 100 17475 120
rect 17445 70 17475 100
rect 17445 50 17450 70
rect 17470 50 17475 70
rect 17445 40 17475 50
rect 17505 120 17535 130
rect 17505 100 17510 120
rect 17530 100 17535 120
rect 17505 70 17535 100
rect 17505 50 17510 70
rect 17530 50 17535 70
rect 17505 40 17535 50
rect 17565 120 17595 130
rect 17565 100 17570 120
rect 17590 100 17595 120
rect 17565 70 17595 100
rect 17565 50 17570 70
rect 17590 50 17595 70
rect 17565 40 17595 50
rect 17625 120 17695 130
rect 17625 100 17630 120
rect 17650 100 17670 120
rect 17690 100 17695 120
rect 17625 70 17695 100
rect 17625 50 17630 70
rect 17650 50 17670 70
rect 17690 50 17695 70
rect 17625 40 17695 50
rect 17905 120 17975 130
rect 17905 100 17910 120
rect 17930 100 17950 120
rect 17970 100 17975 120
rect 17905 70 17975 100
rect 17905 50 17910 70
rect 17930 50 17950 70
rect 17970 50 17975 70
rect 17905 40 17975 50
rect 18005 120 18035 130
rect 18005 100 18010 120
rect 18030 100 18035 120
rect 18005 70 18035 100
rect 18005 50 18010 70
rect 18030 50 18035 70
rect 18005 40 18035 50
rect 18065 120 18095 130
rect 18065 100 18070 120
rect 18090 100 18095 120
rect 18065 70 18095 100
rect 18065 50 18070 70
rect 18090 50 18095 70
rect 18065 40 18095 50
rect 18125 120 18155 130
rect 18125 100 18130 120
rect 18150 100 18155 120
rect 18125 70 18155 100
rect 18125 50 18130 70
rect 18150 50 18155 70
rect 18125 40 18155 50
rect 18185 120 18215 130
rect 18185 100 18190 120
rect 18210 100 18215 120
rect 18185 70 18215 100
rect 18185 50 18190 70
rect 18210 50 18215 70
rect 18185 40 18215 50
rect 18245 120 18275 130
rect 18245 100 18250 120
rect 18270 100 18275 120
rect 18245 70 18275 100
rect 18245 50 18250 70
rect 18270 50 18275 70
rect 18245 40 18275 50
rect 18305 120 18335 130
rect 18305 100 18310 120
rect 18330 100 18335 120
rect 18305 70 18335 100
rect 18305 50 18310 70
rect 18330 50 18335 70
rect 18305 40 18335 50
rect 18365 120 18395 130
rect 18365 100 18370 120
rect 18390 100 18395 120
rect 18365 70 18395 100
rect 18365 50 18370 70
rect 18390 50 18395 70
rect 18365 40 18395 50
rect 18425 120 18455 130
rect 18425 100 18430 120
rect 18450 100 18455 120
rect 18425 70 18455 100
rect 18425 50 18430 70
rect 18450 50 18455 70
rect 18425 40 18455 50
rect 18485 120 18515 130
rect 18485 100 18490 120
rect 18510 100 18515 120
rect 18485 70 18515 100
rect 18485 50 18490 70
rect 18510 50 18515 70
rect 18485 40 18515 50
rect 18545 120 18575 130
rect 18545 100 18550 120
rect 18570 100 18575 120
rect 18545 70 18575 100
rect 18545 50 18550 70
rect 18570 50 18575 70
rect 18545 40 18575 50
rect 18605 120 18635 130
rect 18605 100 18610 120
rect 18630 100 18635 120
rect 18605 70 18635 100
rect 18605 50 18610 70
rect 18630 50 18635 70
rect 18605 40 18635 50
rect 18665 120 18695 130
rect 18665 100 18670 120
rect 18690 100 18695 120
rect 18665 70 18695 100
rect 18665 50 18670 70
rect 18690 50 18695 70
rect 18665 40 18695 50
rect 18725 120 18755 130
rect 18725 100 18730 120
rect 18750 100 18755 120
rect 18725 70 18755 100
rect 18725 50 18730 70
rect 18750 50 18755 70
rect 18725 40 18755 50
rect 18785 120 18815 130
rect 18785 100 18790 120
rect 18810 100 18815 120
rect 18785 70 18815 100
rect 18785 50 18790 70
rect 18810 50 18815 70
rect 18785 40 18815 50
rect 18845 120 18875 130
rect 18845 100 18850 120
rect 18870 100 18875 120
rect 18845 70 18875 100
rect 18845 50 18850 70
rect 18870 50 18875 70
rect 18845 40 18875 50
rect 18905 120 18935 130
rect 18905 100 18910 120
rect 18930 100 18935 120
rect 18905 70 18935 100
rect 18905 50 18910 70
rect 18930 50 18935 70
rect 18905 40 18935 50
rect 18965 120 18995 130
rect 18965 100 18970 120
rect 18990 100 18995 120
rect 18965 70 18995 100
rect 18965 50 18970 70
rect 18990 50 18995 70
rect 18965 40 18995 50
rect 19025 120 19055 130
rect 19025 100 19030 120
rect 19050 100 19055 120
rect 19025 70 19055 100
rect 19025 50 19030 70
rect 19050 50 19055 70
rect 19025 40 19055 50
rect 19085 120 19115 130
rect 19085 100 19090 120
rect 19110 100 19115 120
rect 19085 70 19115 100
rect 19085 50 19090 70
rect 19110 50 19115 70
rect 19085 40 19115 50
rect 19145 120 19215 130
rect 19145 100 19150 120
rect 19170 100 19190 120
rect 19210 100 19215 120
rect 19145 70 19215 100
rect 19145 50 19150 70
rect 19170 50 19190 70
rect 19210 50 19215 70
rect 19145 40 19215 50
rect 16515 5 16545 15
rect 16515 -15 16520 5
rect 16540 -15 16545 5
rect 16515 -25 16545 -15
rect 16600 10 16640 20
rect 16600 -10 16610 10
rect 16630 -10 16640 10
rect 16600 -20 16640 -10
rect 16845 10 16875 20
rect 16845 -10 16850 10
rect 16870 -10 16875 10
rect 16845 -20 16875 -10
rect 16960 10 17000 20
rect 16960 -10 16970 10
rect 16990 -10 17000 10
rect 16960 -20 17000 -10
rect 17205 10 17235 20
rect 17205 -10 17210 10
rect 17230 -10 17235 10
rect 17205 -20 17235 -10
rect 17320 10 17360 20
rect 17320 -10 17330 10
rect 17350 -10 17360 10
rect 17320 -20 17360 -10
rect 17535 10 17565 20
rect 17535 -10 17540 10
rect 17560 -10 17565 10
rect 17535 -20 17565 -10
rect 18035 10 18065 20
rect 18035 -10 18040 10
rect 18060 -10 18065 10
rect 18035 -20 18065 -10
rect 18240 10 18280 20
rect 18240 -10 18250 10
rect 18270 -10 18280 10
rect 18240 -20 18280 -10
rect 18365 10 18395 20
rect 18365 -10 18370 10
rect 18390 -10 18395 10
rect 18365 -20 18395 -10
rect 18600 10 18640 20
rect 18600 -10 18610 10
rect 18630 -10 18640 10
rect 18600 -20 18640 -10
rect 18725 10 18755 20
rect 18725 -10 18730 10
rect 18750 -10 18755 10
rect 18725 -20 18755 -10
rect 18960 10 19000 20
rect 18960 -10 18970 10
rect 18990 -10 19000 10
rect 18960 -20 19000 -10
rect 19055 5 19085 15
rect 19055 -15 19060 5
rect 19080 -15 19085 5
rect 19055 -25 19085 -15
rect 17007 -185 17037 -175
rect 17007 -205 17012 -185
rect 17032 -205 17037 -185
rect 17007 -215 17037 -205
rect 18563 -185 18593 -175
rect 18563 -205 18568 -185
rect 18588 -205 18593 -185
rect 18563 -215 18593 -205
rect 16965 -245 16995 -235
rect 16965 -265 16970 -245
rect 16990 -265 16995 -245
rect 16965 -295 16995 -265
rect 16965 -315 16970 -295
rect 16990 -315 16995 -295
rect 16965 -345 16995 -315
rect 16965 -365 16970 -345
rect 16990 -365 16995 -345
rect 16965 -395 16995 -365
rect 16965 -415 16970 -395
rect 16990 -415 16995 -395
rect 16965 -445 16995 -415
rect 16965 -465 16970 -445
rect 16990 -465 16995 -445
rect 16965 -475 16995 -465
rect 17025 -245 17055 -235
rect 17025 -265 17030 -245
rect 17050 -265 17055 -245
rect 17025 -295 17055 -265
rect 17025 -315 17030 -295
rect 17050 -315 17055 -295
rect 17025 -345 17055 -315
rect 17025 -365 17030 -345
rect 17050 -365 17055 -345
rect 17025 -395 17055 -365
rect 17025 -415 17030 -395
rect 17050 -415 17055 -395
rect 17025 -445 17055 -415
rect 17025 -465 17030 -445
rect 17050 -465 17055 -445
rect 17025 -475 17055 -465
rect 17085 -245 17115 -235
rect 17085 -265 17090 -245
rect 17110 -265 17115 -245
rect 17085 -295 17115 -265
rect 17085 -315 17090 -295
rect 17110 -315 17115 -295
rect 17085 -345 17115 -315
rect 17085 -365 17090 -345
rect 17110 -365 17115 -345
rect 17560 -245 17600 -235
rect 17560 -265 17570 -245
rect 17590 -265 17600 -245
rect 17560 -285 17600 -265
rect 17560 -305 17570 -285
rect 17590 -305 17600 -285
rect 17560 -325 17600 -305
rect 17560 -345 17570 -325
rect 17590 -345 17600 -325
rect 17560 -355 17600 -345
rect 18000 -245 18040 -235
rect 18000 -265 18010 -245
rect 18030 -265 18040 -245
rect 18000 -285 18040 -265
rect 18000 -305 18010 -285
rect 18030 -305 18040 -285
rect 18000 -325 18040 -305
rect 18000 -345 18010 -325
rect 18030 -345 18040 -325
rect 18000 -355 18040 -345
rect 18485 -245 18515 -235
rect 18485 -265 18490 -245
rect 18510 -265 18515 -245
rect 18485 -295 18515 -265
rect 18485 -315 18490 -295
rect 18510 -315 18515 -295
rect 18485 -345 18515 -315
rect 17085 -395 17115 -365
rect 17085 -415 17090 -395
rect 17110 -415 17115 -395
rect 17085 -445 17115 -415
rect 17085 -465 17090 -445
rect 17110 -465 17115 -445
rect 17085 -475 17115 -465
rect 18485 -365 18490 -345
rect 18510 -365 18515 -345
rect 18485 -395 18515 -365
rect 18485 -415 18490 -395
rect 18510 -415 18515 -395
rect 18485 -445 18515 -415
rect 18485 -465 18490 -445
rect 18510 -465 18515 -445
rect 18485 -475 18515 -465
rect 18545 -245 18575 -235
rect 18545 -265 18550 -245
rect 18570 -265 18575 -245
rect 18545 -295 18575 -265
rect 18545 -315 18550 -295
rect 18570 -315 18575 -295
rect 18545 -345 18575 -315
rect 18545 -365 18550 -345
rect 18570 -365 18575 -345
rect 18545 -395 18575 -365
rect 18545 -415 18550 -395
rect 18570 -415 18575 -395
rect 18545 -445 18575 -415
rect 18545 -465 18550 -445
rect 18570 -465 18575 -445
rect 18545 -475 18575 -465
rect 18605 -245 18635 -235
rect 18605 -265 18610 -245
rect 18630 -265 18635 -245
rect 18605 -295 18635 -265
rect 18605 -315 18610 -295
rect 18630 -315 18635 -295
rect 18605 -345 18635 -315
rect 18605 -365 18610 -345
rect 18630 -365 18635 -345
rect 18605 -395 18635 -365
rect 18605 -415 18610 -395
rect 18630 -415 18635 -395
rect 18605 -445 18635 -415
rect 18605 -465 18610 -445
rect 18630 -465 18635 -445
rect 18605 -475 18635 -465
rect 17075 -505 17105 -495
rect 17075 -525 17080 -505
rect 17100 -525 17105 -505
rect 17075 -535 17105 -525
rect 18440 -505 18470 -495
rect 18440 -525 18445 -505
rect 18465 -525 18470 -505
rect 18440 -535 18470 -525
rect 16620 -750 16660 -740
rect 16620 -770 16630 -750
rect 16650 -770 16660 -750
rect 16620 -780 16660 -770
rect 16740 -750 16780 -740
rect 16740 -770 16750 -750
rect 16770 -770 16780 -750
rect 16740 -780 16780 -770
rect 16860 -750 16900 -740
rect 16860 -770 16870 -750
rect 16890 -770 16900 -750
rect 16860 -780 16900 -770
rect 16980 -750 17020 -740
rect 16980 -770 16990 -750
rect 17010 -770 17020 -750
rect 16980 -780 17020 -770
rect 17300 -750 17340 -740
rect 17300 -770 17310 -750
rect 17330 -770 17340 -750
rect 17300 -780 17340 -770
rect 17420 -750 17460 -740
rect 17420 -770 17430 -750
rect 17450 -770 17460 -750
rect 17420 -780 17460 -770
rect 17540 -750 17580 -740
rect 17540 -770 17550 -750
rect 17570 -770 17580 -750
rect 18020 -750 18060 -740
rect 17540 -780 17580 -770
rect 17695 -765 17725 -755
rect 17695 -785 17700 -765
rect 17720 -785 17725 -765
rect 16535 -810 16565 -800
rect 16535 -830 16540 -810
rect 16560 -830 16565 -810
rect 16535 -860 16565 -830
rect 16535 -880 16540 -860
rect 16560 -880 16565 -860
rect 16535 -910 16565 -880
rect 16535 -930 16540 -910
rect 16560 -930 16565 -910
rect 16535 -960 16565 -930
rect 16535 -980 16540 -960
rect 16560 -980 16565 -960
rect 16535 -1010 16565 -980
rect 16535 -1030 16540 -1010
rect 16560 -1030 16565 -1010
rect 16535 -1040 16565 -1030
rect 17075 -810 17185 -800
rect 17075 -830 17080 -810
rect 17100 -830 17120 -810
rect 17140 -830 17160 -810
rect 17180 -830 17185 -810
rect 17075 -860 17185 -830
rect 17075 -880 17080 -860
rect 17100 -880 17120 -860
rect 17140 -880 17160 -860
rect 17180 -880 17185 -860
rect 17075 -910 17185 -880
rect 17075 -930 17080 -910
rect 17100 -930 17120 -910
rect 17140 -930 17160 -910
rect 17180 -930 17185 -910
rect 17075 -960 17185 -930
rect 17075 -980 17080 -960
rect 17100 -980 17120 -960
rect 17140 -980 17160 -960
rect 17180 -980 17185 -960
rect 17075 -1010 17185 -980
rect 17075 -1030 17080 -1010
rect 17100 -1030 17120 -1010
rect 17140 -1030 17160 -1010
rect 17180 -1030 17185 -1010
rect 17075 -1040 17185 -1030
rect 17695 -810 17725 -785
rect 17695 -830 17700 -810
rect 17720 -830 17725 -810
rect 17695 -860 17725 -830
rect 17695 -880 17700 -860
rect 17720 -880 17725 -860
rect 17695 -910 17725 -880
rect 17695 -930 17700 -910
rect 17720 -930 17725 -910
rect 17695 -960 17725 -930
rect 17695 -980 17700 -960
rect 17720 -980 17725 -960
rect 17695 -1010 17725 -980
rect 17695 -1030 17700 -1010
rect 17720 -1030 17725 -1010
rect 17695 -1040 17725 -1030
rect 17875 -765 17905 -755
rect 17875 -785 17880 -765
rect 17900 -785 17905 -765
rect 18020 -770 18030 -750
rect 18050 -770 18060 -750
rect 18020 -780 18060 -770
rect 18140 -750 18180 -740
rect 18140 -770 18150 -750
rect 18170 -770 18180 -750
rect 18140 -780 18180 -770
rect 18260 -750 18300 -740
rect 18260 -770 18270 -750
rect 18290 -770 18300 -750
rect 18260 -780 18300 -770
rect 18580 -750 18620 -740
rect 18580 -770 18590 -750
rect 18610 -770 18620 -750
rect 18580 -780 18620 -770
rect 18700 -750 18740 -740
rect 18700 -770 18710 -750
rect 18730 -770 18740 -750
rect 18700 -780 18740 -770
rect 18820 -750 18860 -740
rect 18820 -770 18830 -750
rect 18850 -770 18860 -750
rect 18820 -780 18860 -770
rect 18940 -750 18980 -740
rect 18940 -770 18950 -750
rect 18970 -770 18980 -750
rect 18940 -780 18980 -770
rect 19030 -770 19070 -760
rect 17875 -810 17905 -785
rect 19030 -790 19040 -770
rect 19060 -790 19070 -770
rect 19030 -800 19070 -790
rect 17875 -830 17880 -810
rect 17900 -830 17905 -810
rect 17875 -860 17905 -830
rect 17875 -880 17880 -860
rect 17900 -880 17905 -860
rect 17875 -910 17905 -880
rect 17875 -930 17880 -910
rect 17900 -930 17905 -910
rect 17875 -960 17905 -930
rect 17875 -980 17880 -960
rect 17900 -980 17905 -960
rect 17875 -1010 17905 -980
rect 17875 -1030 17880 -1010
rect 17900 -1030 17905 -1010
rect 17875 -1040 17905 -1030
rect 18415 -810 18525 -800
rect 18415 -830 18420 -810
rect 18440 -830 18460 -810
rect 18480 -830 18500 -810
rect 18520 -830 18525 -810
rect 18415 -860 18525 -830
rect 18415 -880 18420 -860
rect 18440 -880 18460 -860
rect 18480 -880 18500 -860
rect 18520 -880 18525 -860
rect 18415 -910 18525 -880
rect 18415 -930 18420 -910
rect 18440 -930 18460 -910
rect 18480 -930 18500 -910
rect 18520 -930 18525 -910
rect 18415 -960 18525 -930
rect 18415 -980 18420 -960
rect 18440 -980 18460 -960
rect 18480 -980 18500 -960
rect 18520 -980 18525 -960
rect 18415 -1010 18525 -980
rect 18415 -1030 18420 -1010
rect 18440 -1030 18460 -1010
rect 18480 -1030 18500 -1010
rect 18520 -1030 18525 -1010
rect 18415 -1040 18525 -1030
rect 19035 -810 19065 -800
rect 19035 -830 19040 -810
rect 19060 -830 19065 -810
rect 19035 -860 19065 -830
rect 19035 -880 19040 -860
rect 19060 -880 19065 -860
rect 19035 -910 19065 -880
rect 19035 -930 19040 -910
rect 19060 -930 19065 -910
rect 19035 -960 19065 -930
rect 19035 -980 19040 -960
rect 19060 -980 19065 -960
rect 19035 -1010 19065 -980
rect 19035 -1030 19040 -1010
rect 19060 -1030 19065 -1010
rect 19035 -1040 19065 -1030
rect 17120 -1060 17140 -1040
rect 18460 -1060 18480 -1040
rect 17110 -1070 17150 -1060
rect 17110 -1090 17120 -1070
rect 17140 -1090 17150 -1070
rect 17110 -1100 17150 -1090
rect 18450 -1070 18490 -1060
rect 18450 -1090 18460 -1070
rect 18480 -1090 18490 -1070
rect 18450 -1100 18490 -1090
rect 16740 -1205 16780 -1195
rect 16740 -1225 16750 -1205
rect 16770 -1225 16780 -1205
rect 16740 -1235 16780 -1225
rect 16820 -1205 16860 -1195
rect 16820 -1225 16830 -1205
rect 16850 -1225 16860 -1205
rect 16820 -1235 16860 -1225
rect 16900 -1205 16940 -1195
rect 16900 -1225 16910 -1205
rect 16930 -1225 16940 -1205
rect 16900 -1235 16940 -1225
rect 16980 -1205 17020 -1195
rect 16980 -1225 16990 -1205
rect 17010 -1225 17020 -1205
rect 16980 -1235 17020 -1225
rect 17060 -1205 17100 -1195
rect 17060 -1225 17070 -1205
rect 17090 -1225 17100 -1205
rect 17060 -1235 17100 -1225
rect 17140 -1205 17180 -1195
rect 17140 -1225 17150 -1205
rect 17170 -1225 17180 -1205
rect 17140 -1235 17180 -1225
rect 17220 -1205 17260 -1195
rect 17220 -1225 17230 -1205
rect 17250 -1225 17260 -1205
rect 17220 -1235 17260 -1225
rect 17300 -1205 17340 -1195
rect 17300 -1225 17310 -1205
rect 17330 -1225 17340 -1205
rect 17300 -1235 17340 -1225
rect 17380 -1205 17420 -1195
rect 17380 -1225 17390 -1205
rect 17410 -1225 17420 -1205
rect 17380 -1235 17420 -1225
rect 17460 -1205 17500 -1195
rect 17460 -1225 17470 -1205
rect 17490 -1225 17500 -1205
rect 17460 -1235 17500 -1225
rect 17540 -1205 17580 -1195
rect 17540 -1225 17550 -1205
rect 17570 -1225 17580 -1205
rect 17540 -1235 17580 -1225
rect 17620 -1205 17660 -1195
rect 17620 -1225 17630 -1205
rect 17650 -1225 17660 -1205
rect 17620 -1235 17660 -1225
rect 17700 -1205 17740 -1195
rect 17700 -1225 17710 -1205
rect 17730 -1225 17740 -1205
rect 17700 -1235 17740 -1225
rect 17780 -1205 17820 -1195
rect 17780 -1225 17790 -1205
rect 17810 -1225 17820 -1205
rect 17780 -1235 17820 -1225
rect 17860 -1205 17900 -1195
rect 17860 -1225 17870 -1205
rect 17890 -1225 17900 -1205
rect 17860 -1235 17900 -1225
rect 17940 -1205 17980 -1195
rect 17940 -1225 17950 -1205
rect 17970 -1225 17980 -1205
rect 17940 -1235 17980 -1225
rect 18020 -1205 18060 -1195
rect 18020 -1225 18030 -1205
rect 18050 -1225 18060 -1205
rect 18020 -1235 18060 -1225
rect 18100 -1205 18140 -1195
rect 18100 -1225 18110 -1205
rect 18130 -1225 18140 -1205
rect 18100 -1235 18140 -1225
rect 18180 -1205 18220 -1195
rect 18180 -1225 18190 -1205
rect 18210 -1225 18220 -1205
rect 18180 -1235 18220 -1225
rect 18260 -1205 18300 -1195
rect 18260 -1225 18270 -1205
rect 18290 -1225 18300 -1205
rect 18260 -1235 18300 -1225
rect 18340 -1205 18380 -1195
rect 18340 -1225 18350 -1205
rect 18370 -1225 18380 -1205
rect 18340 -1235 18380 -1225
rect 18420 -1205 18460 -1195
rect 18420 -1225 18430 -1205
rect 18450 -1225 18460 -1205
rect 18420 -1235 18460 -1225
rect 18500 -1205 18540 -1195
rect 18500 -1225 18510 -1205
rect 18530 -1225 18540 -1205
rect 18500 -1235 18540 -1225
rect 18580 -1205 18620 -1195
rect 18580 -1225 18590 -1205
rect 18610 -1225 18620 -1205
rect 18580 -1235 18620 -1225
rect 18660 -1205 18700 -1195
rect 18660 -1225 18670 -1205
rect 18690 -1225 18700 -1205
rect 18660 -1235 18700 -1225
rect 18740 -1205 18780 -1195
rect 18740 -1225 18750 -1205
rect 18770 -1225 18780 -1205
rect 18740 -1235 18780 -1225
rect 16750 -1255 16770 -1235
rect 17790 -1255 17810 -1235
rect 16745 -1265 16775 -1255
rect 16745 -1280 16750 -1265
rect 16700 -1285 16750 -1280
rect 16770 -1285 16775 -1265
rect 16700 -1290 16775 -1285
rect 16700 -1310 16710 -1290
rect 16730 -1310 16775 -1290
rect 16700 -1315 16775 -1310
rect 16700 -1320 16750 -1315
rect 16745 -1335 16750 -1320
rect 16770 -1335 16775 -1315
rect 16745 -1345 16775 -1335
rect 17785 -1265 17815 -1255
rect 17785 -1285 17790 -1265
rect 17810 -1285 17815 -1265
rect 17785 -1315 17815 -1285
rect 17785 -1335 17790 -1315
rect 17810 -1335 17815 -1315
rect 17785 -1345 17815 -1335
rect 18825 -1260 18895 -1255
rect 18825 -1265 18935 -1260
rect 18825 -1285 18830 -1265
rect 18850 -1285 18870 -1265
rect 18890 -1270 18935 -1265
rect 18890 -1285 18905 -1270
rect 18825 -1290 18905 -1285
rect 18925 -1290 18935 -1270
rect 18825 -1310 18935 -1290
rect 18825 -1315 18905 -1310
rect 18825 -1335 18830 -1315
rect 18850 -1335 18870 -1315
rect 18890 -1330 18905 -1315
rect 18925 -1330 18935 -1310
rect 18890 -1335 18935 -1330
rect 18825 -1340 18935 -1335
rect 18825 -1345 18895 -1340
rect 16600 -1525 16640 -1515
rect 16600 -1545 16610 -1525
rect 16630 -1545 16640 -1525
rect 16600 -1555 16640 -1545
rect 16660 -1525 16690 -1515
rect 16660 -1545 16665 -1525
rect 16685 -1545 16690 -1525
rect 16660 -1555 16690 -1545
rect 16710 -1525 16750 -1515
rect 16710 -1545 16720 -1525
rect 16740 -1545 16750 -1525
rect 16710 -1555 16750 -1545
rect 16770 -1525 16800 -1515
rect 16770 -1545 16775 -1525
rect 16795 -1545 16800 -1525
rect 16770 -1555 16800 -1545
rect 16820 -1525 16860 -1515
rect 16820 -1545 16830 -1525
rect 16850 -1545 16860 -1525
rect 16820 -1555 16860 -1545
rect 16880 -1525 16920 -1515
rect 16880 -1545 16890 -1525
rect 16910 -1545 16920 -1525
rect 16880 -1555 16920 -1545
rect 17025 -1525 17065 -1515
rect 17025 -1545 17035 -1525
rect 17055 -1545 17065 -1525
rect 17025 -1555 17065 -1545
rect 17135 -1525 17175 -1515
rect 17135 -1545 17145 -1525
rect 17165 -1545 17175 -1525
rect 17135 -1555 17175 -1545
rect 17245 -1525 17285 -1515
rect 17245 -1545 17255 -1525
rect 17275 -1545 17285 -1525
rect 17245 -1555 17285 -1545
rect 17305 -1525 17335 -1515
rect 17305 -1545 17310 -1525
rect 17330 -1545 17335 -1525
rect 17305 -1555 17335 -1545
rect 17355 -1525 17395 -1515
rect 17355 -1545 17365 -1525
rect 17385 -1545 17395 -1525
rect 17355 -1555 17395 -1545
rect 17465 -1525 17505 -1515
rect 17465 -1545 17475 -1525
rect 17495 -1545 17505 -1525
rect 17465 -1555 17505 -1545
rect 17615 -1525 17655 -1515
rect 17615 -1545 17625 -1525
rect 17645 -1545 17655 -1525
rect 17615 -1555 17655 -1545
rect 17725 -1525 17765 -1515
rect 17725 -1545 17735 -1525
rect 17755 -1545 17765 -1525
rect 17725 -1555 17765 -1545
rect 17785 -1525 17815 -1515
rect 17785 -1545 17790 -1525
rect 17810 -1545 17815 -1525
rect 17785 -1555 17815 -1545
rect 17835 -1525 17875 -1515
rect 17835 -1545 17845 -1525
rect 17865 -1545 17875 -1525
rect 17835 -1555 17875 -1545
rect 17945 -1525 17985 -1515
rect 17945 -1545 17955 -1525
rect 17975 -1545 17985 -1525
rect 17945 -1555 17985 -1545
rect 18005 -1525 18045 -1515
rect 18005 -1545 18015 -1525
rect 18035 -1545 18045 -1525
rect 18005 -1555 18045 -1545
rect 18150 -1525 18190 -1515
rect 18150 -1545 18160 -1525
rect 18180 -1545 18190 -1525
rect 18150 -1555 18190 -1545
rect 18260 -1525 18300 -1515
rect 18260 -1545 18270 -1525
rect 18290 -1545 18300 -1525
rect 18260 -1555 18300 -1545
rect 18320 -1525 18350 -1515
rect 18320 -1545 18325 -1525
rect 18345 -1545 18350 -1525
rect 18320 -1555 18350 -1545
rect 18370 -1525 18410 -1515
rect 18370 -1545 18380 -1525
rect 18400 -1545 18410 -1525
rect 18370 -1555 18410 -1545
rect 18480 -1525 18520 -1515
rect 18480 -1545 18490 -1525
rect 18510 -1545 18520 -1525
rect 18480 -1555 18520 -1545
rect 18590 -1525 18630 -1515
rect 18590 -1545 18600 -1525
rect 18620 -1545 18630 -1525
rect 18590 -1555 18630 -1545
rect 16605 -1575 16635 -1555
rect 16665 -1575 16685 -1555
rect 16720 -1575 16740 -1555
rect 16830 -1575 16850 -1555
rect 16880 -1575 16910 -1555
rect 17030 -1575 17060 -1555
rect 17145 -1575 17165 -1555
rect 17255 -1575 17275 -1555
rect 17365 -1575 17385 -1555
rect 17470 -1575 17500 -1555
rect 17620 -1575 17650 -1555
rect 17735 -1575 17755 -1555
rect 17845 -1575 17865 -1555
rect 17955 -1575 17975 -1555
rect 18010 -1575 18035 -1555
rect 18155 -1575 18185 -1555
rect 18270 -1575 18290 -1555
rect 18380 -1575 18400 -1555
rect 18490 -1575 18510 -1555
rect 18595 -1575 18625 -1555
rect 16565 -1585 16635 -1575
rect 16565 -1605 16570 -1585
rect 16590 -1605 16610 -1585
rect 16630 -1605 16635 -1585
rect 16565 -1635 16635 -1605
rect 16565 -1655 16570 -1635
rect 16590 -1655 16610 -1635
rect 16630 -1655 16635 -1635
rect 16565 -1665 16635 -1655
rect 16660 -1585 16690 -1575
rect 16660 -1605 16665 -1585
rect 16685 -1605 16690 -1585
rect 16660 -1635 16690 -1605
rect 16660 -1655 16665 -1635
rect 16685 -1655 16690 -1635
rect 16660 -1665 16690 -1655
rect 16715 -1585 16745 -1575
rect 16715 -1605 16720 -1585
rect 16740 -1605 16745 -1585
rect 16715 -1635 16745 -1605
rect 16715 -1655 16720 -1635
rect 16740 -1655 16745 -1635
rect 16715 -1665 16745 -1655
rect 16770 -1585 16800 -1575
rect 16770 -1605 16775 -1585
rect 16795 -1605 16800 -1585
rect 16770 -1635 16800 -1605
rect 16770 -1655 16775 -1635
rect 16795 -1655 16800 -1635
rect 16770 -1665 16800 -1655
rect 16825 -1585 16855 -1575
rect 16825 -1605 16830 -1585
rect 16850 -1605 16855 -1585
rect 16825 -1635 16855 -1605
rect 16825 -1655 16830 -1635
rect 16850 -1655 16855 -1635
rect 16825 -1665 16855 -1655
rect 16880 -1585 16950 -1575
rect 16880 -1605 16885 -1585
rect 16905 -1605 16925 -1585
rect 16945 -1605 16950 -1585
rect 16880 -1635 16950 -1605
rect 16880 -1655 16885 -1635
rect 16905 -1655 16925 -1635
rect 16945 -1655 16950 -1635
rect 16880 -1665 16950 -1655
rect 16990 -1585 17060 -1575
rect 16990 -1605 16995 -1585
rect 17015 -1605 17035 -1585
rect 17055 -1605 17060 -1585
rect 16990 -1635 17060 -1605
rect 16990 -1655 16995 -1635
rect 17015 -1655 17035 -1635
rect 17055 -1655 17060 -1635
rect 16990 -1665 17060 -1655
rect 17085 -1585 17115 -1575
rect 17085 -1605 17090 -1585
rect 17110 -1605 17115 -1585
rect 17085 -1635 17115 -1605
rect 17085 -1655 17090 -1635
rect 17110 -1655 17115 -1635
rect 17085 -1665 17115 -1655
rect 17140 -1585 17170 -1575
rect 17140 -1605 17145 -1585
rect 17165 -1605 17170 -1585
rect 17140 -1635 17170 -1605
rect 17140 -1655 17145 -1635
rect 17165 -1655 17170 -1635
rect 17140 -1665 17170 -1655
rect 17195 -1585 17225 -1575
rect 17195 -1605 17200 -1585
rect 17220 -1605 17225 -1585
rect 17195 -1635 17225 -1605
rect 17195 -1655 17200 -1635
rect 17220 -1655 17225 -1635
rect 17195 -1665 17225 -1655
rect 17250 -1585 17280 -1575
rect 17250 -1605 17255 -1585
rect 17275 -1605 17280 -1585
rect 17250 -1635 17280 -1605
rect 17250 -1655 17255 -1635
rect 17275 -1655 17280 -1635
rect 17250 -1665 17280 -1655
rect 17305 -1585 17335 -1575
rect 17305 -1605 17310 -1585
rect 17330 -1605 17335 -1585
rect 17305 -1635 17335 -1605
rect 17305 -1655 17310 -1635
rect 17330 -1655 17335 -1635
rect 17305 -1665 17335 -1655
rect 17360 -1585 17390 -1575
rect 17360 -1605 17365 -1585
rect 17385 -1605 17390 -1585
rect 17360 -1635 17390 -1605
rect 17360 -1655 17365 -1635
rect 17385 -1655 17390 -1635
rect 17360 -1665 17390 -1655
rect 17415 -1585 17445 -1575
rect 17415 -1605 17420 -1585
rect 17440 -1605 17445 -1585
rect 17415 -1635 17445 -1605
rect 17415 -1655 17420 -1635
rect 17440 -1655 17445 -1635
rect 17415 -1665 17445 -1655
rect 17470 -1585 17540 -1575
rect 17470 -1605 17475 -1585
rect 17495 -1605 17515 -1585
rect 17535 -1605 17540 -1585
rect 17470 -1635 17540 -1605
rect 17470 -1655 17475 -1635
rect 17495 -1655 17515 -1635
rect 17535 -1655 17540 -1635
rect 17470 -1665 17540 -1655
rect 17580 -1585 17650 -1575
rect 17580 -1605 17585 -1585
rect 17605 -1605 17625 -1585
rect 17645 -1605 17650 -1585
rect 17580 -1635 17650 -1605
rect 17580 -1655 17585 -1635
rect 17605 -1655 17625 -1635
rect 17645 -1655 17650 -1635
rect 17580 -1665 17650 -1655
rect 17675 -1585 17705 -1575
rect 17675 -1605 17680 -1585
rect 17700 -1605 17705 -1585
rect 17675 -1635 17705 -1605
rect 17675 -1655 17680 -1635
rect 17700 -1655 17705 -1635
rect 17675 -1665 17705 -1655
rect 17730 -1585 17760 -1575
rect 17730 -1605 17735 -1585
rect 17755 -1605 17760 -1585
rect 17730 -1635 17760 -1605
rect 17730 -1655 17735 -1635
rect 17755 -1655 17760 -1635
rect 17730 -1665 17760 -1655
rect 17785 -1585 17815 -1575
rect 17785 -1605 17790 -1585
rect 17810 -1605 17815 -1585
rect 17785 -1635 17815 -1605
rect 17785 -1655 17790 -1635
rect 17810 -1655 17815 -1635
rect 17785 -1665 17815 -1655
rect 17840 -1585 17870 -1575
rect 17840 -1605 17845 -1585
rect 17865 -1605 17870 -1585
rect 17840 -1635 17870 -1605
rect 17840 -1655 17845 -1635
rect 17865 -1655 17870 -1635
rect 17840 -1665 17870 -1655
rect 17895 -1585 17925 -1575
rect 17895 -1605 17900 -1585
rect 17920 -1605 17925 -1585
rect 17895 -1635 17925 -1605
rect 17895 -1655 17900 -1635
rect 17920 -1655 17925 -1635
rect 17895 -1665 17925 -1655
rect 17950 -1585 17980 -1575
rect 17950 -1605 17955 -1585
rect 17975 -1605 17980 -1585
rect 17950 -1635 17980 -1605
rect 17950 -1655 17955 -1635
rect 17975 -1655 17980 -1635
rect 17950 -1665 17980 -1655
rect 18005 -1585 18075 -1575
rect 18005 -1605 18010 -1585
rect 18030 -1605 18050 -1585
rect 18070 -1605 18075 -1585
rect 18005 -1635 18075 -1605
rect 18005 -1655 18010 -1635
rect 18030 -1655 18050 -1635
rect 18070 -1655 18075 -1635
rect 18005 -1665 18075 -1655
rect 18115 -1585 18185 -1575
rect 18115 -1605 18120 -1585
rect 18140 -1605 18160 -1585
rect 18180 -1605 18185 -1585
rect 18115 -1635 18185 -1605
rect 18115 -1655 18120 -1635
rect 18140 -1655 18160 -1635
rect 18180 -1655 18185 -1635
rect 18115 -1665 18185 -1655
rect 18210 -1585 18240 -1575
rect 18210 -1605 18215 -1585
rect 18235 -1605 18240 -1585
rect 18210 -1635 18240 -1605
rect 18210 -1655 18215 -1635
rect 18235 -1655 18240 -1635
rect 18210 -1665 18240 -1655
rect 18265 -1585 18295 -1575
rect 18265 -1605 18270 -1585
rect 18290 -1605 18295 -1585
rect 18265 -1635 18295 -1605
rect 18265 -1655 18270 -1635
rect 18290 -1655 18295 -1635
rect 18265 -1665 18295 -1655
rect 18320 -1585 18350 -1575
rect 18320 -1605 18325 -1585
rect 18345 -1605 18350 -1585
rect 18320 -1635 18350 -1605
rect 18320 -1655 18325 -1635
rect 18345 -1655 18350 -1635
rect 18320 -1665 18350 -1655
rect 18375 -1585 18405 -1575
rect 18375 -1605 18380 -1585
rect 18400 -1605 18405 -1585
rect 18375 -1635 18405 -1605
rect 18375 -1655 18380 -1635
rect 18400 -1655 18405 -1635
rect 18375 -1665 18405 -1655
rect 18430 -1585 18460 -1575
rect 18430 -1605 18435 -1585
rect 18455 -1605 18460 -1585
rect 18430 -1635 18460 -1605
rect 18430 -1655 18435 -1635
rect 18455 -1655 18460 -1635
rect 18430 -1665 18460 -1655
rect 18485 -1585 18515 -1575
rect 18485 -1605 18490 -1585
rect 18510 -1605 18515 -1585
rect 18485 -1635 18515 -1605
rect 18485 -1655 18490 -1635
rect 18510 -1655 18515 -1635
rect 18485 -1665 18515 -1655
rect 18540 -1585 18570 -1575
rect 18540 -1605 18545 -1585
rect 18565 -1605 18570 -1585
rect 18540 -1635 18570 -1605
rect 18540 -1655 18545 -1635
rect 18565 -1655 18570 -1635
rect 18540 -1665 18570 -1655
rect 18595 -1585 18665 -1575
rect 18595 -1605 18600 -1585
rect 18620 -1605 18640 -1585
rect 18660 -1605 18665 -1585
rect 18595 -1635 18665 -1605
rect 18595 -1655 18600 -1635
rect 18620 -1655 18640 -1635
rect 18660 -1655 18665 -1635
rect 18595 -1665 18665 -1655
rect 16775 -1685 16795 -1665
rect 17090 -1685 17110 -1665
rect 17310 -1685 17330 -1665
rect 17680 -1685 17700 -1665
rect 17790 -1685 17810 -1665
rect 17900 -1685 17920 -1665
rect 18325 -1685 18345 -1665
rect 18545 -1685 18565 -1665
rect 16765 -1695 16805 -1685
rect 16765 -1715 16775 -1695
rect 16795 -1715 16805 -1695
rect 16765 -1725 16805 -1715
rect 17080 -1695 17120 -1685
rect 17080 -1715 17090 -1695
rect 17110 -1715 17120 -1695
rect 17080 -1725 17120 -1715
rect 17190 -1695 17230 -1685
rect 17190 -1715 17200 -1695
rect 17220 -1715 17230 -1695
rect 17190 -1725 17230 -1715
rect 17300 -1695 17340 -1685
rect 17300 -1715 17310 -1695
rect 17330 -1715 17340 -1695
rect 17300 -1725 17340 -1715
rect 17410 -1695 17450 -1685
rect 17410 -1715 17420 -1695
rect 17440 -1715 17450 -1695
rect 17410 -1725 17450 -1715
rect 17670 -1695 17710 -1685
rect 17670 -1715 17680 -1695
rect 17700 -1715 17710 -1695
rect 17670 -1725 17710 -1715
rect 17780 -1695 17820 -1685
rect 17780 -1715 17790 -1695
rect 17810 -1715 17820 -1695
rect 17780 -1725 17820 -1715
rect 17890 -1695 17930 -1685
rect 17890 -1715 17900 -1695
rect 17920 -1715 17930 -1695
rect 17890 -1725 17930 -1715
rect 18205 -1695 18245 -1685
rect 18205 -1715 18215 -1695
rect 18235 -1715 18245 -1695
rect 18205 -1725 18245 -1715
rect 18315 -1695 18355 -1685
rect 18315 -1715 18325 -1695
rect 18345 -1715 18355 -1695
rect 18315 -1725 18355 -1715
rect 18425 -1695 18465 -1685
rect 18425 -1715 18435 -1695
rect 18455 -1715 18465 -1695
rect 18425 -1725 18465 -1715
rect 18535 -1695 18575 -1685
rect 18535 -1715 18545 -1695
rect 18565 -1715 18575 -1695
rect 18535 -1725 18575 -1715
rect 17425 -2005 17470 -2000
rect 17425 -2030 17435 -2005
rect 17460 -2030 17470 -2005
rect 17425 -2035 17470 -2030
rect 18124 -2005 18169 -2000
rect 18124 -2030 18134 -2005
rect 18159 -2030 18169 -2005
rect 18124 -2035 18169 -2030
rect 16795 -2240 18805 -2115
rect 17440 -2795 17480 -2240
rect 18120 -2795 18160 -2240
rect 16485 -2905 16520 -2895
rect 16485 -2930 16490 -2905
rect 16515 -2930 16520 -2905
rect 16795 -2920 18805 -2795
rect 19080 -2905 19115 -2895
rect 16485 -2940 16520 -2930
rect 16160 -3030 16195 -3020
rect 16160 -3055 16165 -3030
rect 16190 -3055 16195 -3030
rect 16160 -3065 16195 -3055
rect 15950 -3121 15985 -3110
rect 15950 -3146 15955 -3121
rect 15980 -3146 15985 -3121
rect 15950 -3156 15985 -3146
rect 16255 -3100 16280 -3065
rect 16580 -2975 16605 -2940
rect 17440 -3475 17480 -2920
rect 18120 -3475 18160 -2920
rect 19080 -2930 19085 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2940 19115 -2930
rect 18995 -2975 19020 -2940
rect 19405 -3002 19440 -2992
rect 19405 -3027 19410 -3002
rect 19435 -3027 19440 -3002
rect 19405 -3037 19440 -3027
rect 19320 -3072 19345 -3037
rect 19610 -3120 19645 -3110
rect 19610 -3145 19615 -3120
rect 19640 -3145 19645 -3120
rect 19610 -3156 19645 -3145
rect 16795 -3600 18805 -3475
rect 15950 -3794 15985 -3784
rect 15950 -3819 15955 -3794
rect 15980 -3819 15985 -3794
rect 15950 -3829 15985 -3819
rect 16195 -3889 16220 -3854
rect 16280 -3899 16315 -3889
rect 16280 -3924 16285 -3899
rect 16310 -3924 16315 -3899
rect 16280 -3934 16315 -3924
rect 16520 -3964 16545 -3929
rect 16605 -3974 16640 -3964
rect 16605 -3999 16610 -3974
rect 16635 -3999 16640 -3974
rect 16605 -4009 16640 -3999
rect 17440 -4125 17480 -3600
rect 17780 -4210 17820 -4120
rect 18120 -4125 18160 -3600
rect 19055 -3964 19080 -3929
rect 19380 -3889 19405 -3854
rect 19610 -3794 19645 -3784
rect 19610 -3819 19615 -3794
rect 19640 -3819 19645 -3794
rect 19610 -3829 19645 -3819
rect 19285 -3899 19320 -3889
rect 19285 -3924 19290 -3899
rect 19315 -3924 19320 -3899
rect 19285 -3934 19320 -3924
rect 18960 -3974 18995 -3964
rect 18960 -3999 18965 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4009 18995 -3999
rect 17780 -4230 17790 -4210
rect 17810 -4230 17820 -4210
rect 17780 -4250 17820 -4230
rect 17780 -4270 17790 -4250
rect 17810 -4270 17820 -4250
rect 17780 -4290 17820 -4270
rect 17780 -4310 17790 -4290
rect 17810 -4310 17820 -4290
rect 17780 -4320 17820 -4310
<< viali >>
rect 16495 1435 16515 1455
rect 17790 1435 17810 1455
rect 16375 1300 16395 1320
rect 16495 1300 16515 1320
rect 16615 1300 16635 1320
rect 16895 1300 16915 1320
rect 16950 1300 16970 1320
rect 17005 1300 17025 1320
rect 17060 1300 17080 1320
rect 17115 1300 17135 1320
rect 17225 1300 17245 1320
rect 17505 1300 17525 1320
rect 17570 1300 17590 1320
rect 17625 1300 17645 1320
rect 17680 1300 17700 1320
rect 17735 1300 17755 1320
rect 17790 1300 17810 1320
rect 17845 1300 17865 1320
rect 17900 1300 17920 1320
rect 17955 1300 17975 1320
rect 18010 1300 18030 1320
rect 18075 1300 18095 1320
rect 18355 1300 18375 1320
rect 18465 1300 18485 1320
rect 18520 1300 18540 1320
rect 18575 1300 18595 1320
rect 18630 1300 18650 1320
rect 18685 1300 18705 1320
rect 16440 1130 16460 1150
rect 16550 1130 16570 1150
rect 16950 1130 16970 1150
rect 17060 1130 17080 1150
rect 17170 1130 17190 1150
rect 17625 1130 17645 1150
rect 17735 1130 17755 1150
rect 17845 1130 17865 1150
rect 17955 1130 17975 1150
rect 18410 1130 18430 1150
rect 18520 1130 18540 1150
rect 18630 1130 18650 1150
rect 16980 940 17000 960
rect 17160 940 17180 960
rect 17340 940 17360 960
rect 17520 940 17540 960
rect 17700 940 17720 960
rect 17880 940 17900 960
rect 18060 940 18080 960
rect 18240 940 18260 960
rect 18420 940 18440 960
rect 18600 940 18620 960
rect 18915 940 18935 960
rect 19025 940 19045 960
rect 19085 940 19105 960
rect 16980 880 17000 900
rect 16445 840 16465 860
rect 16555 840 16575 860
rect 16665 840 16685 860
rect 16980 830 17000 850
rect 16980 780 17000 800
rect 16980 730 17000 750
rect 16490 670 16510 690
rect 16555 670 16575 690
rect 16620 670 16640 690
rect 16980 680 17000 700
rect 16980 630 17000 650
rect 17070 880 17090 900
rect 17070 830 17090 850
rect 17070 780 17090 800
rect 17070 730 17090 750
rect 17070 680 17090 700
rect 17070 630 17090 650
rect 17160 880 17180 900
rect 17160 830 17180 850
rect 17160 780 17180 800
rect 17160 730 17180 750
rect 17160 680 17180 700
rect 17160 630 17180 650
rect 17250 880 17270 900
rect 17250 830 17270 850
rect 17250 780 17270 800
rect 17250 730 17270 750
rect 17250 680 17270 700
rect 17250 630 17270 650
rect 17340 880 17360 900
rect 17340 830 17360 850
rect 17340 780 17360 800
rect 17340 730 17360 750
rect 17340 680 17360 700
rect 17340 630 17360 650
rect 17430 880 17450 900
rect 17430 830 17450 850
rect 17430 780 17450 800
rect 17430 730 17450 750
rect 17430 680 17450 700
rect 17430 630 17450 650
rect 17520 880 17540 900
rect 17520 830 17540 850
rect 17520 780 17540 800
rect 17520 730 17540 750
rect 17520 680 17540 700
rect 17520 630 17540 650
rect 17610 880 17630 900
rect 17610 830 17630 850
rect 17610 780 17630 800
rect 17610 730 17630 750
rect 17610 680 17630 700
rect 17610 630 17630 650
rect 17700 880 17720 900
rect 17700 830 17720 850
rect 17700 780 17720 800
rect 17700 730 17720 750
rect 17700 680 17720 700
rect 17700 630 17720 650
rect 17790 880 17810 900
rect 17790 830 17810 850
rect 17790 780 17810 800
rect 17790 730 17810 750
rect 17790 680 17810 700
rect 17790 630 17810 650
rect 17880 880 17900 900
rect 17880 830 17900 850
rect 17880 780 17900 800
rect 17880 730 17900 750
rect 17880 680 17900 700
rect 17880 630 17900 650
rect 17970 880 17990 900
rect 17970 830 17990 850
rect 17970 780 17990 800
rect 17970 730 17990 750
rect 17970 680 17990 700
rect 17970 630 17990 650
rect 18060 880 18080 900
rect 18060 830 18080 850
rect 18060 780 18080 800
rect 18060 730 18080 750
rect 18060 680 18080 700
rect 18060 630 18080 650
rect 18150 880 18170 900
rect 18150 830 18170 850
rect 18150 780 18170 800
rect 18150 730 18170 750
rect 18150 680 18170 700
rect 18150 630 18170 650
rect 18240 880 18260 900
rect 18240 830 18260 850
rect 18240 780 18260 800
rect 18240 730 18260 750
rect 18240 680 18260 700
rect 18240 630 18260 650
rect 18330 880 18350 900
rect 18330 830 18350 850
rect 18330 780 18350 800
rect 18330 730 18350 750
rect 18330 680 18350 700
rect 18330 630 18350 650
rect 18420 880 18440 900
rect 18420 830 18440 850
rect 18420 780 18440 800
rect 18420 730 18440 750
rect 18420 680 18440 700
rect 18420 630 18440 650
rect 18510 880 18530 900
rect 18510 830 18530 850
rect 18510 780 18530 800
rect 18510 730 18530 750
rect 18510 680 18530 700
rect 18510 630 18530 650
rect 18600 880 18620 900
rect 18600 830 18620 850
rect 18600 780 18620 800
rect 18600 730 18620 750
rect 18915 880 18935 900
rect 18915 830 18935 850
rect 18915 780 18935 800
rect 18915 730 18935 750
rect 18970 880 18990 900
rect 18970 830 18990 850
rect 18970 780 18990 800
rect 18970 730 18990 750
rect 19025 880 19045 900
rect 19025 830 19045 850
rect 19025 780 19045 800
rect 19025 730 19045 750
rect 19080 880 19100 900
rect 19080 830 19100 850
rect 19080 780 19100 800
rect 19080 730 19100 750
rect 18600 680 18620 700
rect 18600 630 18620 650
rect 19010 610 19030 630
rect 17115 570 17135 590
rect 17205 570 17225 590
rect 17295 570 17315 590
rect 17385 570 17405 590
rect 17475 570 17495 590
rect 17565 570 17585 590
rect 17655 570 17675 590
rect 17745 570 17765 590
rect 17835 570 17855 590
rect 17925 570 17945 590
rect 18015 570 18035 590
rect 18105 570 18125 590
rect 18195 570 18215 590
rect 18285 570 18305 590
rect 18375 570 18395 590
rect 18465 570 18485 590
rect 16430 160 16450 180
rect 17630 160 17650 180
rect 17950 160 17970 180
rect 19150 160 19170 180
rect 16430 100 16450 120
rect 16430 50 16450 70
rect 16490 100 16510 120
rect 16490 50 16510 70
rect 16550 100 16570 120
rect 16550 50 16570 70
rect 16610 100 16630 120
rect 16610 50 16630 70
rect 16670 100 16690 120
rect 16670 50 16690 70
rect 16730 100 16750 120
rect 16730 50 16750 70
rect 16790 100 16810 120
rect 16790 50 16810 70
rect 16850 100 16870 120
rect 16850 50 16870 70
rect 16910 100 16930 120
rect 16910 50 16930 70
rect 16970 100 16990 120
rect 16970 50 16990 70
rect 17030 100 17050 120
rect 17030 50 17050 70
rect 17090 100 17110 120
rect 17090 50 17110 70
rect 17150 100 17170 120
rect 17150 50 17170 70
rect 17210 100 17230 120
rect 17210 50 17230 70
rect 17270 100 17290 120
rect 17270 50 17290 70
rect 17330 100 17350 120
rect 17330 50 17350 70
rect 17390 100 17410 120
rect 17390 50 17410 70
rect 17450 100 17470 120
rect 17450 50 17470 70
rect 17510 100 17530 120
rect 17510 50 17530 70
rect 17570 100 17590 120
rect 17570 50 17590 70
rect 17630 100 17650 120
rect 17630 50 17650 70
rect 17950 100 17970 120
rect 17950 50 17970 70
rect 18010 100 18030 120
rect 18010 50 18030 70
rect 18070 100 18090 120
rect 18070 50 18090 70
rect 18130 100 18150 120
rect 18130 50 18150 70
rect 18190 100 18210 120
rect 18190 50 18210 70
rect 18250 100 18270 120
rect 18250 50 18270 70
rect 18310 100 18330 120
rect 18310 50 18330 70
rect 18370 100 18390 120
rect 18370 50 18390 70
rect 18430 100 18450 120
rect 18430 50 18450 70
rect 18490 100 18510 120
rect 18490 50 18510 70
rect 18550 100 18570 120
rect 18550 50 18570 70
rect 18610 100 18630 120
rect 18610 50 18630 70
rect 18670 100 18690 120
rect 18670 50 18690 70
rect 18730 100 18750 120
rect 18730 50 18750 70
rect 18790 100 18810 120
rect 18790 50 18810 70
rect 18850 100 18870 120
rect 18850 50 18870 70
rect 18910 100 18930 120
rect 18910 50 18930 70
rect 18970 100 18990 120
rect 18970 50 18990 70
rect 19030 100 19050 120
rect 19030 50 19050 70
rect 19090 100 19110 120
rect 19090 50 19110 70
rect 19150 100 19170 120
rect 19150 50 19170 70
rect 16520 -15 16540 5
rect 16610 -10 16630 10
rect 16850 -10 16870 10
rect 16970 -10 16990 10
rect 17210 -10 17230 10
rect 17330 -10 17350 10
rect 17540 -10 17560 10
rect 18040 -10 18060 10
rect 18250 -10 18270 10
rect 18370 -10 18390 10
rect 18610 -10 18630 10
rect 18730 -10 18750 10
rect 18970 -10 18990 10
rect 19060 -15 19080 5
rect 17012 -205 17032 -185
rect 18568 -205 18588 -185
rect 16970 -265 16990 -245
rect 16970 -315 16990 -295
rect 16970 -365 16990 -345
rect 16970 -415 16990 -395
rect 16970 -465 16990 -445
rect 17030 -265 17050 -245
rect 17030 -315 17050 -295
rect 17030 -365 17050 -345
rect 17030 -415 17050 -395
rect 17030 -465 17050 -445
rect 17090 -265 17110 -245
rect 17090 -315 17110 -295
rect 17090 -365 17110 -345
rect 17570 -265 17590 -245
rect 17570 -305 17590 -285
rect 17570 -345 17590 -325
rect 18010 -265 18030 -245
rect 18010 -305 18030 -285
rect 18010 -345 18030 -325
rect 18490 -265 18510 -245
rect 18490 -315 18510 -295
rect 17090 -415 17110 -395
rect 17090 -465 17110 -445
rect 18490 -365 18510 -345
rect 18490 -415 18510 -395
rect 18490 -465 18510 -445
rect 18550 -265 18570 -245
rect 18550 -315 18570 -295
rect 18550 -365 18570 -345
rect 18550 -415 18570 -395
rect 18550 -465 18570 -445
rect 18610 -265 18630 -245
rect 18610 -315 18630 -295
rect 18610 -365 18630 -345
rect 18610 -415 18630 -395
rect 18610 -465 18630 -445
rect 17080 -525 17100 -505
rect 18445 -525 18465 -505
rect 16630 -770 16650 -750
rect 16750 -770 16770 -750
rect 16870 -770 16890 -750
rect 16990 -770 17010 -750
rect 17310 -770 17330 -750
rect 17430 -770 17450 -750
rect 17550 -770 17570 -750
rect 17700 -785 17720 -765
rect 16540 -830 16560 -810
rect 16540 -880 16560 -860
rect 16540 -930 16560 -910
rect 16540 -980 16560 -960
rect 16540 -1030 16560 -1010
rect 17880 -785 17900 -765
rect 18030 -770 18050 -750
rect 18150 -770 18170 -750
rect 18270 -770 18290 -750
rect 18590 -770 18610 -750
rect 18710 -770 18730 -750
rect 18830 -770 18850 -750
rect 18950 -770 18970 -750
rect 19040 -790 19060 -770
rect 17120 -1090 17140 -1070
rect 18460 -1090 18480 -1070
rect 16750 -1225 16770 -1205
rect 16830 -1225 16850 -1205
rect 16910 -1225 16930 -1205
rect 16990 -1225 17010 -1205
rect 17070 -1225 17090 -1205
rect 17150 -1225 17170 -1205
rect 17230 -1225 17250 -1205
rect 17310 -1225 17330 -1205
rect 17390 -1225 17410 -1205
rect 17470 -1225 17490 -1205
rect 17550 -1225 17570 -1205
rect 17630 -1225 17650 -1205
rect 17710 -1225 17730 -1205
rect 17790 -1225 17810 -1205
rect 17870 -1225 17890 -1205
rect 17950 -1225 17970 -1205
rect 18030 -1225 18050 -1205
rect 18110 -1225 18130 -1205
rect 18190 -1225 18210 -1205
rect 18270 -1225 18290 -1205
rect 18350 -1225 18370 -1205
rect 18430 -1225 18450 -1205
rect 18510 -1225 18530 -1205
rect 18590 -1225 18610 -1205
rect 18670 -1225 18690 -1205
rect 18750 -1225 18770 -1205
rect 16710 -1310 16730 -1290
rect 18905 -1290 18925 -1270
rect 18905 -1330 18925 -1310
rect 16610 -1545 16630 -1525
rect 16665 -1545 16685 -1525
rect 16720 -1545 16740 -1525
rect 16775 -1545 16795 -1525
rect 16830 -1545 16850 -1525
rect 16890 -1545 16910 -1525
rect 17035 -1545 17055 -1525
rect 17145 -1545 17165 -1525
rect 17255 -1545 17275 -1525
rect 17310 -1545 17330 -1525
rect 17365 -1545 17385 -1525
rect 17475 -1545 17495 -1525
rect 17625 -1545 17645 -1525
rect 17735 -1545 17755 -1525
rect 17790 -1545 17810 -1525
rect 17845 -1545 17865 -1525
rect 17955 -1545 17975 -1525
rect 18015 -1545 18035 -1525
rect 18160 -1545 18180 -1525
rect 18270 -1545 18290 -1525
rect 18325 -1545 18345 -1525
rect 18380 -1545 18400 -1525
rect 18490 -1545 18510 -1525
rect 18600 -1545 18620 -1525
rect 17200 -1605 17220 -1585
rect 17200 -1655 17220 -1635
rect 17420 -1605 17440 -1585
rect 17420 -1655 17440 -1635
rect 18215 -1605 18235 -1585
rect 18215 -1655 18235 -1635
rect 18435 -1605 18455 -1585
rect 18435 -1655 18455 -1635
rect 16775 -1715 16795 -1695
rect 17090 -1715 17110 -1695
rect 17200 -1715 17220 -1695
rect 17310 -1715 17330 -1695
rect 17420 -1715 17440 -1695
rect 17680 -1715 17700 -1695
rect 17790 -1715 17810 -1695
rect 17900 -1715 17920 -1695
rect 18215 -1715 18235 -1695
rect 18325 -1715 18345 -1695
rect 18435 -1715 18455 -1695
rect 18545 -1715 18565 -1695
rect 17435 -2030 17460 -2005
rect 18134 -2030 18159 -2005
rect 16490 -2930 16515 -2905
rect 16165 -3055 16190 -3030
rect 15955 -3146 15980 -3121
rect 19085 -2930 19110 -2905
rect 19410 -3027 19435 -3002
rect 19615 -3145 19640 -3120
rect 15955 -3819 15980 -3794
rect 16285 -3924 16310 -3899
rect 16610 -3999 16635 -3974
rect 19615 -3819 19640 -3794
rect 19290 -3924 19315 -3899
rect 18965 -3999 18990 -3974
rect 17790 -4230 17810 -4210
rect 17790 -4270 17810 -4250
rect 17790 -4310 17810 -4290
<< metal1 >>
rect 15645 -45 15765 -40
rect 15645 -75 15650 -45
rect 15680 -75 15690 -45
rect 15720 -75 15730 -45
rect 15760 -75 15765 -45
rect 15645 -85 15765 -75
rect 15645 -115 15650 -85
rect 15680 -115 15690 -85
rect 15720 -115 15730 -85
rect 15760 -115 15765 -85
rect 15645 -125 15765 -115
rect 15645 -155 15650 -125
rect 15680 -155 15690 -125
rect 15720 -155 15730 -125
rect 15760 -155 15765 -125
rect 15645 -4345 15765 -155
rect 15790 -1795 15815 1640
rect 15890 1155 15930 1160
rect 15890 1125 15895 1155
rect 15925 1125 15930 1155
rect 15890 -1385 15930 1125
rect 15890 -1415 15895 -1385
rect 15925 -1415 15930 -1385
rect 15890 -1420 15930 -1415
rect 15945 185 15985 190
rect 15945 155 15950 185
rect 15980 155 15985 185
rect 15785 -1800 15825 -1795
rect 15785 -1830 15790 -1800
rect 15820 -1830 15825 -1800
rect 15785 -1835 15825 -1830
rect 15945 -3110 15985 155
rect 16040 -1740 16060 1640
rect 16030 -1745 16070 -1740
rect 16030 -1775 16035 -1745
rect 16065 -1775 16070 -1745
rect 16030 -1780 16070 -1775
rect 16115 -1850 16135 1640
rect 16485 1460 16525 1465
rect 16485 1430 16490 1460
rect 16520 1430 16525 1460
rect 16485 1425 16525 1430
rect 16365 1405 16405 1410
rect 16365 1375 16370 1405
rect 16400 1375 16405 1405
rect 16365 1365 16405 1375
rect 16365 1335 16370 1365
rect 16400 1335 16405 1365
rect 16365 1325 16405 1335
rect 16365 1295 16370 1325
rect 16400 1295 16405 1325
rect 16365 1290 16405 1295
rect 16485 1405 16525 1410
rect 16485 1375 16490 1405
rect 16520 1375 16525 1405
rect 16485 1365 16525 1375
rect 16485 1335 16490 1365
rect 16520 1335 16525 1365
rect 16485 1325 16525 1335
rect 16485 1295 16490 1325
rect 16520 1295 16525 1325
rect 16485 1290 16525 1295
rect 16605 1405 16645 1410
rect 16605 1375 16610 1405
rect 16640 1375 16645 1405
rect 16605 1365 16645 1375
rect 16605 1335 16610 1365
rect 16640 1335 16645 1365
rect 16605 1325 16645 1335
rect 16605 1295 16610 1325
rect 16640 1295 16645 1325
rect 16605 1290 16645 1295
rect 16885 1405 16925 1410
rect 16885 1375 16890 1405
rect 16920 1375 16925 1405
rect 16885 1365 16925 1375
rect 16885 1335 16890 1365
rect 16920 1335 16925 1365
rect 16885 1325 16925 1335
rect 16950 1330 16970 1640
rect 17050 1460 17090 1465
rect 17050 1430 17055 1460
rect 17085 1430 17090 1460
rect 17050 1425 17090 1430
rect 16995 1405 17035 1410
rect 16995 1375 17000 1405
rect 17030 1375 17035 1405
rect 16995 1365 17035 1375
rect 16995 1335 17000 1365
rect 17030 1335 17035 1365
rect 16885 1295 16890 1325
rect 16920 1295 16925 1325
rect 16885 1290 16925 1295
rect 16945 1320 16975 1330
rect 16945 1300 16950 1320
rect 16970 1300 16975 1320
rect 16945 1290 16975 1300
rect 16995 1325 17035 1335
rect 16995 1295 17000 1325
rect 17030 1295 17035 1325
rect 16995 1290 17035 1295
rect 17055 1320 17085 1425
rect 17055 1300 17060 1320
rect 17080 1300 17085 1320
rect 17055 1290 17085 1300
rect 17105 1405 17145 1410
rect 17105 1375 17110 1405
rect 17140 1375 17145 1405
rect 17105 1365 17145 1375
rect 17105 1335 17110 1365
rect 17140 1335 17145 1365
rect 17105 1325 17145 1335
rect 17105 1295 17110 1325
rect 17140 1295 17145 1325
rect 17105 1290 17145 1295
rect 17215 1405 17255 1410
rect 17215 1375 17220 1405
rect 17250 1375 17255 1405
rect 17215 1365 17255 1375
rect 17215 1335 17220 1365
rect 17250 1335 17255 1365
rect 17215 1325 17255 1335
rect 17215 1295 17220 1325
rect 17250 1295 17255 1325
rect 17215 1290 17255 1295
rect 17495 1405 17535 1410
rect 17495 1375 17500 1405
rect 17530 1375 17535 1405
rect 17495 1365 17535 1375
rect 17495 1335 17500 1365
rect 17530 1335 17535 1365
rect 17495 1325 17535 1335
rect 17495 1295 17500 1325
rect 17530 1295 17535 1325
rect 17495 1290 17535 1295
rect 17560 1405 17600 1410
rect 17560 1375 17565 1405
rect 17595 1375 17600 1405
rect 17560 1365 17600 1375
rect 17560 1335 17565 1365
rect 17595 1335 17600 1365
rect 17560 1325 17600 1335
rect 17560 1295 17565 1325
rect 17595 1295 17600 1325
rect 17560 1290 17600 1295
rect 17620 1320 17650 1640
rect 17620 1300 17625 1320
rect 17645 1300 17650 1320
rect 17620 1290 17650 1300
rect 17670 1405 17710 1410
rect 17670 1375 17675 1405
rect 17705 1375 17710 1405
rect 17670 1365 17710 1375
rect 17670 1335 17675 1365
rect 17705 1335 17710 1365
rect 17670 1325 17710 1335
rect 17670 1295 17675 1325
rect 17705 1295 17710 1325
rect 17670 1290 17710 1295
rect 17730 1320 17760 1640
rect 17780 1460 17820 1465
rect 17780 1430 17785 1460
rect 17815 1430 17820 1460
rect 17780 1425 17820 1430
rect 17730 1300 17735 1320
rect 17755 1300 17760 1320
rect 17730 1290 17760 1300
rect 17780 1405 17820 1410
rect 17780 1375 17785 1405
rect 17815 1375 17820 1405
rect 17780 1365 17820 1375
rect 17780 1335 17785 1365
rect 17815 1335 17820 1365
rect 17780 1325 17820 1335
rect 17780 1295 17785 1325
rect 17815 1295 17820 1325
rect 17780 1290 17820 1295
rect 17840 1320 17870 1640
rect 17840 1300 17845 1320
rect 17865 1300 17870 1320
rect 17840 1290 17870 1300
rect 17890 1405 17930 1410
rect 17890 1375 17895 1405
rect 17925 1375 17930 1405
rect 17890 1365 17930 1375
rect 17890 1335 17895 1365
rect 17925 1335 17930 1365
rect 17890 1325 17930 1335
rect 17890 1295 17895 1325
rect 17925 1295 17930 1325
rect 17890 1290 17930 1295
rect 17950 1320 17980 1640
rect 18510 1430 18515 1460
rect 18545 1430 18550 1460
rect 18510 1425 18550 1430
rect 17950 1300 17955 1320
rect 17975 1300 17980 1320
rect 17950 1290 17980 1300
rect 18000 1405 18040 1410
rect 18000 1375 18005 1405
rect 18035 1375 18040 1405
rect 18000 1365 18040 1375
rect 18000 1335 18005 1365
rect 18035 1335 18040 1365
rect 18000 1325 18040 1335
rect 18000 1295 18005 1325
rect 18035 1295 18040 1325
rect 18000 1290 18040 1295
rect 18065 1405 18105 1410
rect 18065 1375 18070 1405
rect 18100 1375 18105 1405
rect 18065 1365 18105 1375
rect 18065 1335 18070 1365
rect 18100 1335 18105 1365
rect 18065 1325 18105 1335
rect 18065 1295 18070 1325
rect 18100 1295 18105 1325
rect 18065 1290 18105 1295
rect 18345 1405 18385 1410
rect 18345 1375 18350 1405
rect 18380 1375 18385 1405
rect 18345 1365 18385 1375
rect 18345 1335 18350 1365
rect 18380 1335 18385 1365
rect 18345 1325 18385 1335
rect 18345 1295 18350 1325
rect 18380 1295 18385 1325
rect 18345 1290 18385 1295
rect 18455 1405 18495 1410
rect 18455 1375 18460 1405
rect 18490 1375 18495 1405
rect 18455 1365 18495 1375
rect 18455 1335 18460 1365
rect 18490 1335 18495 1365
rect 18455 1325 18495 1335
rect 18520 1330 18540 1425
rect 18565 1405 18605 1410
rect 18565 1375 18570 1405
rect 18600 1375 18605 1405
rect 18565 1365 18605 1375
rect 18565 1335 18570 1365
rect 18600 1335 18605 1365
rect 18455 1295 18460 1325
rect 18490 1295 18495 1325
rect 18455 1290 18495 1295
rect 18515 1320 18545 1330
rect 18515 1300 18520 1320
rect 18540 1300 18545 1320
rect 18515 1290 18545 1300
rect 18565 1325 18605 1335
rect 18630 1330 18650 1640
rect 18675 1405 18715 1410
rect 18675 1375 18680 1405
rect 18710 1375 18715 1405
rect 18675 1365 18715 1375
rect 18675 1335 18680 1365
rect 18710 1335 18715 1365
rect 18565 1295 18570 1325
rect 18600 1295 18605 1325
rect 18565 1290 18605 1295
rect 18625 1320 18655 1330
rect 18625 1300 18630 1320
rect 18650 1300 18655 1320
rect 18625 1290 18655 1300
rect 18675 1325 18715 1335
rect 18675 1295 18680 1325
rect 18710 1295 18715 1325
rect 18675 1290 18715 1295
rect 16430 1155 16470 1160
rect 16430 1125 16435 1155
rect 16465 1125 16470 1155
rect 16430 1120 16470 1125
rect 16540 1155 16580 1160
rect 16540 1125 16545 1155
rect 16575 1125 16580 1155
rect 16540 1100 16580 1125
rect 16940 1155 16980 1160
rect 16940 1125 16945 1155
rect 16975 1125 16980 1155
rect 16940 1120 16980 1125
rect 17050 1155 17090 1160
rect 17050 1125 17055 1155
rect 17085 1125 17090 1155
rect 17050 1120 17090 1125
rect 17160 1155 17200 1160
rect 17160 1125 17165 1155
rect 17195 1125 17200 1155
rect 17160 1120 17200 1125
rect 17615 1155 17655 1160
rect 17615 1125 17620 1155
rect 17650 1125 17655 1155
rect 17615 1120 17655 1125
rect 17725 1155 17765 1160
rect 17725 1125 17730 1155
rect 17760 1125 17765 1155
rect 17725 1120 17765 1125
rect 17835 1155 17875 1160
rect 17835 1125 17840 1155
rect 17870 1125 17875 1155
rect 17835 1120 17875 1125
rect 17945 1155 17985 1160
rect 17945 1125 17950 1155
rect 17980 1125 17985 1155
rect 17945 1120 17985 1125
rect 18400 1155 18440 1160
rect 18400 1125 18405 1155
rect 18435 1125 18440 1155
rect 18400 1120 18440 1125
rect 18510 1155 18550 1160
rect 18510 1125 18515 1155
rect 18545 1125 18550 1155
rect 18510 1120 18550 1125
rect 18620 1155 18660 1160
rect 18620 1125 18625 1155
rect 18655 1125 18660 1155
rect 18620 1120 18660 1125
rect 16540 1070 16545 1100
rect 16575 1070 16580 1100
rect 16540 1065 16580 1070
rect 16435 1045 16475 1050
rect 16435 1015 16440 1045
rect 16470 1015 16475 1045
rect 16435 1005 16475 1015
rect 16435 975 16440 1005
rect 16470 975 16475 1005
rect 16435 965 16475 975
rect 16435 935 16440 965
rect 16470 935 16475 965
rect 16435 930 16475 935
rect 16655 1045 16695 1050
rect 16655 1015 16660 1045
rect 16690 1015 16695 1045
rect 16655 1005 16695 1015
rect 16655 975 16660 1005
rect 16690 975 16695 1005
rect 16655 965 16695 975
rect 16655 935 16660 965
rect 16690 935 16695 965
rect 16655 930 16695 935
rect 16970 1045 17010 1050
rect 16970 1015 16975 1045
rect 17005 1015 17010 1045
rect 16970 1005 17010 1015
rect 16970 975 16975 1005
rect 17005 975 17010 1005
rect 16970 965 17010 975
rect 16970 935 16975 965
rect 17005 935 17010 965
rect 16970 930 17010 935
rect 17150 1045 17190 1050
rect 17150 1015 17155 1045
rect 17185 1015 17190 1045
rect 17150 1005 17190 1015
rect 17150 975 17155 1005
rect 17185 975 17190 1005
rect 17150 965 17190 975
rect 17150 935 17155 965
rect 17185 935 17190 965
rect 17150 930 17190 935
rect 17330 1045 17370 1050
rect 17330 1015 17335 1045
rect 17365 1015 17370 1045
rect 17330 1005 17370 1015
rect 17330 975 17335 1005
rect 17365 975 17370 1005
rect 17330 965 17370 975
rect 17330 935 17335 965
rect 17365 935 17370 965
rect 17330 930 17370 935
rect 17510 1045 17550 1050
rect 17510 1015 17515 1045
rect 17545 1015 17550 1045
rect 17510 1005 17550 1015
rect 17510 975 17515 1005
rect 17545 975 17550 1005
rect 17510 965 17550 975
rect 17510 935 17515 965
rect 17545 935 17550 965
rect 17510 930 17550 935
rect 17690 1045 17730 1050
rect 17690 1015 17695 1045
rect 17725 1015 17730 1045
rect 17690 1005 17730 1015
rect 17690 975 17695 1005
rect 17725 975 17730 1005
rect 17690 965 17730 975
rect 17690 935 17695 965
rect 17725 935 17730 965
rect 17690 930 17730 935
rect 17870 1045 17910 1050
rect 17870 1015 17875 1045
rect 17905 1015 17910 1045
rect 17870 1005 17910 1015
rect 17870 975 17875 1005
rect 17905 975 17910 1005
rect 17870 965 17910 975
rect 17870 935 17875 965
rect 17905 935 17910 965
rect 17870 930 17910 935
rect 18050 1045 18090 1050
rect 18050 1015 18055 1045
rect 18085 1015 18090 1045
rect 18050 1005 18090 1015
rect 18050 975 18055 1005
rect 18085 975 18090 1005
rect 18050 965 18090 975
rect 18050 935 18055 965
rect 18085 935 18090 965
rect 18050 930 18090 935
rect 18230 1045 18270 1050
rect 18230 1015 18235 1045
rect 18265 1015 18270 1045
rect 18230 1005 18270 1015
rect 18230 975 18235 1005
rect 18265 975 18270 1005
rect 18230 965 18270 975
rect 18230 935 18235 965
rect 18265 935 18270 965
rect 18230 930 18270 935
rect 18410 1045 18450 1050
rect 18410 1015 18415 1045
rect 18445 1015 18450 1045
rect 18410 1005 18450 1015
rect 18410 975 18415 1005
rect 18445 975 18450 1005
rect 18410 965 18450 975
rect 18410 935 18415 965
rect 18445 935 18450 965
rect 18410 930 18450 935
rect 18590 1045 18630 1050
rect 18590 1015 18595 1045
rect 18625 1015 18630 1045
rect 18590 1005 18630 1015
rect 18590 975 18595 1005
rect 18625 975 18630 1005
rect 18590 965 18630 975
rect 18590 935 18595 965
rect 18625 935 18630 965
rect 18590 930 18630 935
rect 18905 1045 18945 1050
rect 18905 1015 18910 1045
rect 18940 1015 18945 1045
rect 18905 1005 18945 1015
rect 18905 975 18910 1005
rect 18940 975 18945 1005
rect 18905 965 18945 975
rect 18905 935 18910 965
rect 18940 935 18945 965
rect 18905 930 18945 935
rect 16445 870 16465 930
rect 16665 870 16685 930
rect 16975 900 17005 910
rect 16975 880 16980 900
rect 17000 880 17005 900
rect 16435 860 16475 870
rect 16435 840 16445 860
rect 16465 840 16475 860
rect 16435 830 16475 840
rect 16545 865 16585 870
rect 16545 835 16550 865
rect 16580 835 16585 865
rect 16545 830 16585 835
rect 16655 860 16695 870
rect 16655 840 16665 860
rect 16685 840 16695 860
rect 16655 830 16695 840
rect 16780 865 16820 870
rect 16780 835 16785 865
rect 16815 835 16820 865
rect 16780 830 16820 835
rect 16975 850 17005 880
rect 16975 830 16980 850
rect 17000 830 17005 850
rect 16480 695 16520 700
rect 16480 665 16485 695
rect 16515 665 16520 695
rect 16315 540 16355 545
rect 16315 510 16320 540
rect 16350 510 16355 540
rect 16315 505 16355 510
rect 16260 485 16300 490
rect 16260 455 16265 485
rect 16295 455 16300 485
rect 16260 450 16300 455
rect 16205 430 16245 435
rect 16205 400 16210 430
rect 16240 400 16245 430
rect 16205 395 16245 400
rect 16215 -1280 16235 395
rect 16270 -175 16290 450
rect 16260 -180 16300 -175
rect 16260 -210 16265 -180
rect 16295 -210 16300 -180
rect 16260 -215 16300 -210
rect 16205 -1285 16245 -1280
rect 16205 -1315 16210 -1285
rect 16240 -1315 16245 -1285
rect 16205 -1320 16245 -1315
rect 16105 -1855 16145 -1850
rect 16105 -1885 16110 -1855
rect 16140 -1885 16145 -1855
rect 16105 -1890 16145 -1885
rect 16155 -1945 16195 -1940
rect 16155 -1975 16160 -1945
rect 16190 -1975 16195 -1945
rect 16155 -3020 16195 -1975
rect 16270 -2095 16290 -215
rect 16325 -495 16345 505
rect 16420 320 16460 325
rect 16420 290 16425 320
rect 16455 290 16460 320
rect 16420 280 16460 290
rect 16420 250 16425 280
rect 16455 250 16460 280
rect 16420 240 16460 250
rect 16420 210 16425 240
rect 16455 210 16460 240
rect 16420 205 16460 210
rect 16425 180 16455 205
rect 16425 160 16430 180
rect 16450 160 16455 180
rect 16425 120 16455 160
rect 16480 185 16520 665
rect 16545 690 16585 700
rect 16545 670 16555 690
rect 16575 670 16585 690
rect 16545 660 16585 670
rect 16610 695 16650 700
rect 16610 665 16615 695
rect 16645 665 16650 695
rect 16610 660 16650 665
rect 16555 435 16575 660
rect 16790 490 16810 830
rect 16975 800 17005 830
rect 16975 780 16980 800
rect 17000 780 17005 800
rect 16975 750 17005 780
rect 16975 730 16980 750
rect 17000 730 17005 750
rect 16975 700 17005 730
rect 16975 680 16980 700
rect 17000 680 17005 700
rect 16975 650 17005 680
rect 16975 630 16980 650
rect 17000 630 17005 650
rect 16975 620 17005 630
rect 17065 900 17095 910
rect 17065 880 17070 900
rect 17090 880 17095 900
rect 17065 850 17095 880
rect 17065 830 17070 850
rect 17090 830 17095 850
rect 17065 800 17095 830
rect 17065 780 17070 800
rect 17090 780 17095 800
rect 17065 750 17095 780
rect 17065 730 17070 750
rect 17090 730 17095 750
rect 17065 700 17095 730
rect 17065 680 17070 700
rect 17090 680 17095 700
rect 17065 650 17095 680
rect 17065 630 17070 650
rect 17090 630 17095 650
rect 16780 485 16820 490
rect 16780 455 16785 485
rect 16815 455 16820 485
rect 16780 450 16820 455
rect 16545 430 16585 435
rect 16545 400 16550 430
rect 16580 400 16585 430
rect 16545 395 16585 400
rect 17065 380 17095 630
rect 17155 900 17185 910
rect 17155 880 17160 900
rect 17180 880 17185 900
rect 17155 850 17185 880
rect 17155 830 17160 850
rect 17180 830 17185 850
rect 17155 800 17185 830
rect 17155 780 17160 800
rect 17180 780 17185 800
rect 17155 750 17185 780
rect 17155 730 17160 750
rect 17180 730 17185 750
rect 17155 700 17185 730
rect 17155 680 17160 700
rect 17180 680 17185 700
rect 17155 650 17185 680
rect 17155 630 17160 650
rect 17180 630 17185 650
rect 17155 620 17185 630
rect 17245 900 17275 910
rect 17245 880 17250 900
rect 17270 880 17275 900
rect 17245 850 17275 880
rect 17245 830 17250 850
rect 17270 830 17275 850
rect 17245 800 17275 830
rect 17245 780 17250 800
rect 17270 780 17275 800
rect 17245 750 17275 780
rect 17245 730 17250 750
rect 17270 730 17275 750
rect 17245 700 17275 730
rect 17245 680 17250 700
rect 17270 680 17275 700
rect 17245 650 17275 680
rect 17245 630 17250 650
rect 17270 630 17275 650
rect 17245 620 17275 630
rect 17335 900 17365 910
rect 17335 880 17340 900
rect 17360 880 17365 900
rect 17335 850 17365 880
rect 17335 830 17340 850
rect 17360 830 17365 850
rect 17335 800 17365 830
rect 17335 780 17340 800
rect 17360 780 17365 800
rect 17335 750 17365 780
rect 17335 730 17340 750
rect 17360 730 17365 750
rect 17335 700 17365 730
rect 17335 680 17340 700
rect 17360 680 17365 700
rect 17335 650 17365 680
rect 17335 630 17340 650
rect 17360 630 17365 650
rect 17335 620 17365 630
rect 17425 900 17455 910
rect 17425 880 17430 900
rect 17450 880 17455 900
rect 17425 850 17455 880
rect 17425 830 17430 850
rect 17450 830 17455 850
rect 17425 800 17455 830
rect 17425 780 17430 800
rect 17450 780 17455 800
rect 17425 750 17455 780
rect 17425 730 17430 750
rect 17450 730 17455 750
rect 17425 700 17455 730
rect 17425 680 17430 700
rect 17450 680 17455 700
rect 17425 650 17455 680
rect 17425 630 17430 650
rect 17450 630 17455 650
rect 17425 620 17455 630
rect 17515 900 17545 910
rect 17515 880 17520 900
rect 17540 880 17545 900
rect 17515 850 17545 880
rect 17515 830 17520 850
rect 17540 830 17545 850
rect 17515 800 17545 830
rect 17515 780 17520 800
rect 17540 780 17545 800
rect 17515 750 17545 780
rect 17515 730 17520 750
rect 17540 730 17545 750
rect 17515 700 17545 730
rect 17515 680 17520 700
rect 17540 680 17545 700
rect 17515 650 17545 680
rect 17515 630 17520 650
rect 17540 630 17545 650
rect 17515 620 17545 630
rect 17605 900 17635 910
rect 17605 880 17610 900
rect 17630 880 17635 900
rect 17605 850 17635 880
rect 17605 830 17610 850
rect 17630 830 17635 850
rect 17605 800 17635 830
rect 17605 780 17610 800
rect 17630 780 17635 800
rect 17605 750 17635 780
rect 17605 730 17610 750
rect 17630 730 17635 750
rect 17605 700 17635 730
rect 17605 680 17610 700
rect 17630 680 17635 700
rect 17605 650 17635 680
rect 17605 630 17610 650
rect 17630 630 17635 650
rect 17605 620 17635 630
rect 17695 900 17725 910
rect 17695 880 17700 900
rect 17720 880 17725 900
rect 17695 850 17725 880
rect 17695 830 17700 850
rect 17720 830 17725 850
rect 17695 800 17725 830
rect 17695 780 17700 800
rect 17720 780 17725 800
rect 17695 750 17725 780
rect 17695 730 17700 750
rect 17720 730 17725 750
rect 17695 700 17725 730
rect 17695 680 17700 700
rect 17720 680 17725 700
rect 17695 650 17725 680
rect 17695 630 17700 650
rect 17720 630 17725 650
rect 17695 620 17725 630
rect 17785 900 17815 910
rect 17785 880 17790 900
rect 17810 880 17815 900
rect 17785 850 17815 880
rect 17785 830 17790 850
rect 17810 830 17815 850
rect 17785 800 17815 830
rect 17785 780 17790 800
rect 17810 780 17815 800
rect 17785 750 17815 780
rect 17785 730 17790 750
rect 17810 730 17815 750
rect 17785 700 17815 730
rect 17785 680 17790 700
rect 17810 680 17815 700
rect 17785 650 17815 680
rect 17785 630 17790 650
rect 17810 630 17815 650
rect 17110 595 17145 600
rect 17140 565 17145 595
rect 17110 560 17145 565
rect 17195 595 17235 600
rect 17195 565 17200 595
rect 17230 565 17235 595
rect 17195 560 17235 565
rect 17250 435 17270 620
rect 17285 595 17325 600
rect 17285 565 17290 595
rect 17320 565 17325 595
rect 17285 560 17325 565
rect 17375 595 17415 600
rect 17375 565 17380 595
rect 17410 565 17415 595
rect 17375 560 17415 565
rect 17430 490 17450 620
rect 17465 595 17505 600
rect 17465 565 17470 595
rect 17500 565 17505 595
rect 17465 560 17505 565
rect 17555 595 17595 600
rect 17555 565 17560 595
rect 17590 565 17595 595
rect 17555 560 17595 565
rect 17610 545 17630 620
rect 17645 595 17770 600
rect 17645 565 17650 595
rect 17680 565 17695 595
rect 17725 565 17740 595
rect 17645 560 17770 565
rect 17600 540 17640 545
rect 17600 510 17605 540
rect 17635 510 17640 540
rect 17600 505 17640 510
rect 17420 485 17460 490
rect 17420 455 17425 485
rect 17455 455 17460 485
rect 17420 450 17460 455
rect 17240 430 17280 435
rect 17240 400 17245 430
rect 17275 400 17280 430
rect 17240 395 17280 400
rect 17060 375 17100 380
rect 17060 345 17065 375
rect 17095 345 17100 375
rect 17060 340 17100 345
rect 16540 320 16580 325
rect 16540 290 16545 320
rect 16575 290 16580 320
rect 16540 280 16580 290
rect 16540 250 16545 280
rect 16575 250 16580 280
rect 16540 240 16580 250
rect 16540 210 16545 240
rect 16575 210 16580 240
rect 16540 205 16580 210
rect 16660 320 16700 325
rect 16660 290 16665 320
rect 16695 290 16700 320
rect 16660 280 16700 290
rect 16660 250 16665 280
rect 16695 250 16700 280
rect 16660 240 16700 250
rect 16660 210 16665 240
rect 16695 210 16700 240
rect 16660 205 16700 210
rect 16780 320 16820 325
rect 16780 290 16785 320
rect 16815 290 16820 320
rect 16780 280 16820 290
rect 16780 250 16785 280
rect 16815 250 16820 280
rect 16780 240 16820 250
rect 16780 210 16785 240
rect 16815 210 16820 240
rect 16780 205 16820 210
rect 16900 320 16940 325
rect 16900 290 16905 320
rect 16935 290 16940 320
rect 16900 280 16940 290
rect 16900 250 16905 280
rect 16935 250 16940 280
rect 16900 240 16940 250
rect 16900 210 16905 240
rect 16935 210 16940 240
rect 16900 205 16940 210
rect 17020 320 17060 325
rect 17020 290 17025 320
rect 17055 290 17060 320
rect 17020 280 17060 290
rect 17020 250 17025 280
rect 17055 250 17060 280
rect 17020 240 17060 250
rect 17020 210 17025 240
rect 17055 210 17060 240
rect 17020 205 17060 210
rect 17140 320 17180 325
rect 17140 290 17145 320
rect 17175 290 17180 320
rect 17140 280 17180 290
rect 17140 250 17145 280
rect 17175 250 17180 280
rect 17140 240 17180 250
rect 17140 210 17145 240
rect 17175 210 17180 240
rect 17140 205 17180 210
rect 17260 320 17300 325
rect 17260 290 17265 320
rect 17295 290 17300 320
rect 17260 280 17300 290
rect 17260 250 17265 280
rect 17295 250 17300 280
rect 17260 240 17300 250
rect 17260 210 17265 240
rect 17295 210 17300 240
rect 17260 205 17300 210
rect 17380 320 17420 325
rect 17380 290 17385 320
rect 17415 290 17420 320
rect 17380 280 17420 290
rect 17380 250 17385 280
rect 17415 250 17420 280
rect 17380 240 17420 250
rect 17380 210 17385 240
rect 17415 210 17420 240
rect 17380 205 17420 210
rect 17500 320 17540 325
rect 17500 290 17505 320
rect 17535 290 17540 320
rect 17500 280 17540 290
rect 17500 250 17505 280
rect 17535 250 17540 280
rect 17500 240 17540 250
rect 17500 210 17505 240
rect 17535 210 17540 240
rect 17500 205 17540 210
rect 17620 320 17660 325
rect 17620 290 17625 320
rect 17655 290 17660 320
rect 17620 280 17660 290
rect 17620 250 17625 280
rect 17655 250 17660 280
rect 17620 240 17660 250
rect 17620 210 17625 240
rect 17655 210 17660 240
rect 17620 205 17660 210
rect 16480 155 16485 185
rect 16515 155 16520 185
rect 16480 150 16520 155
rect 16425 100 16430 120
rect 16450 100 16455 120
rect 16425 70 16455 100
rect 16425 50 16430 70
rect 16450 50 16455 70
rect 16425 40 16455 50
rect 16485 120 16515 150
rect 16485 100 16490 120
rect 16510 100 16515 120
rect 16485 70 16515 100
rect 16485 50 16490 70
rect 16510 50 16515 70
rect 16485 40 16515 50
rect 16545 120 16575 205
rect 16545 100 16550 120
rect 16570 100 16575 120
rect 16545 70 16575 100
rect 16545 50 16550 70
rect 16570 50 16575 70
rect 16545 40 16575 50
rect 16605 120 16635 130
rect 16605 100 16610 120
rect 16630 100 16635 120
rect 16605 70 16635 100
rect 16605 50 16610 70
rect 16630 50 16635 70
rect 16605 20 16635 50
rect 16665 120 16695 205
rect 16665 100 16670 120
rect 16690 100 16695 120
rect 16665 70 16695 100
rect 16665 50 16670 70
rect 16690 50 16695 70
rect 16665 40 16695 50
rect 16725 120 16755 130
rect 16725 100 16730 120
rect 16750 100 16755 120
rect 16725 70 16755 100
rect 16725 50 16730 70
rect 16750 50 16755 70
rect 16600 15 16640 20
rect 16515 5 16545 15
rect 16515 -15 16520 5
rect 16540 -15 16545 5
rect 16515 -40 16545 -15
rect 16600 -15 16605 15
rect 16635 -15 16640 15
rect 16600 -20 16640 -15
rect 16725 -40 16755 50
rect 16785 120 16815 205
rect 16840 185 16880 190
rect 16840 155 16845 185
rect 16875 155 16880 185
rect 16840 150 16880 155
rect 16785 100 16790 120
rect 16810 100 16815 120
rect 16785 70 16815 100
rect 16785 50 16790 70
rect 16810 50 16815 70
rect 16785 40 16815 50
rect 16845 120 16875 150
rect 16845 100 16850 120
rect 16870 100 16875 120
rect 16845 70 16875 100
rect 16845 50 16850 70
rect 16870 50 16875 70
rect 16845 40 16875 50
rect 16905 120 16935 205
rect 16905 100 16910 120
rect 16930 100 16935 120
rect 16905 70 16935 100
rect 16905 50 16910 70
rect 16930 50 16935 70
rect 16905 40 16935 50
rect 16965 120 16995 130
rect 16965 100 16970 120
rect 16990 100 16995 120
rect 16965 70 16995 100
rect 16965 50 16970 70
rect 16990 50 16995 70
rect 16965 20 16995 50
rect 17025 120 17055 205
rect 17025 100 17030 120
rect 17050 100 17055 120
rect 17025 70 17055 100
rect 17025 50 17030 70
rect 17050 50 17055 70
rect 17025 40 17055 50
rect 17085 120 17115 130
rect 17085 100 17090 120
rect 17110 100 17115 120
rect 17085 70 17115 100
rect 17085 50 17090 70
rect 17110 50 17115 70
rect 16845 10 16875 20
rect 16845 -10 16850 10
rect 16870 -10 16875 10
rect 16845 -40 16875 -10
rect 16960 15 17000 20
rect 16960 -15 16965 15
rect 16995 -15 17000 15
rect 16960 -20 17000 -15
rect 16510 -45 16550 -40
rect 16510 -75 16515 -45
rect 16545 -75 16550 -45
rect 16510 -85 16550 -75
rect 16510 -115 16515 -85
rect 16545 -115 16550 -85
rect 16510 -125 16550 -115
rect 16510 -155 16515 -125
rect 16545 -155 16550 -125
rect 16510 -160 16550 -155
rect 16720 -45 16760 -40
rect 16720 -75 16725 -45
rect 16755 -75 16760 -45
rect 16720 -85 16760 -75
rect 16720 -115 16725 -85
rect 16755 -115 16760 -85
rect 16720 -125 16760 -115
rect 16720 -155 16725 -125
rect 16755 -155 16760 -125
rect 16720 -160 16760 -155
rect 16840 -45 16880 -40
rect 16840 -75 16845 -45
rect 16875 -75 16880 -45
rect 16840 -85 16880 -75
rect 16840 -115 16845 -85
rect 16875 -115 16880 -85
rect 16840 -125 16880 -115
rect 16840 -155 16845 -125
rect 16875 -155 16880 -125
rect 16840 -160 16880 -155
rect 16970 -235 16990 -20
rect 17085 -40 17115 50
rect 17145 120 17175 205
rect 17200 185 17240 190
rect 17200 155 17205 185
rect 17235 155 17240 185
rect 17200 150 17240 155
rect 17145 100 17150 120
rect 17170 100 17175 120
rect 17145 70 17175 100
rect 17145 50 17150 70
rect 17170 50 17175 70
rect 17145 40 17175 50
rect 17205 120 17235 150
rect 17205 100 17210 120
rect 17230 100 17235 120
rect 17205 70 17235 100
rect 17205 50 17210 70
rect 17230 50 17235 70
rect 17205 40 17235 50
rect 17265 120 17295 205
rect 17265 100 17270 120
rect 17290 100 17295 120
rect 17265 70 17295 100
rect 17265 50 17270 70
rect 17290 50 17295 70
rect 17265 40 17295 50
rect 17325 120 17355 130
rect 17325 100 17330 120
rect 17350 100 17355 120
rect 17325 70 17355 100
rect 17325 50 17330 70
rect 17350 50 17355 70
rect 17325 20 17355 50
rect 17385 120 17415 205
rect 17385 100 17390 120
rect 17410 100 17415 120
rect 17385 70 17415 100
rect 17385 50 17390 70
rect 17410 50 17415 70
rect 17385 40 17415 50
rect 17445 120 17475 130
rect 17445 100 17450 120
rect 17470 100 17475 120
rect 17445 70 17475 100
rect 17445 50 17450 70
rect 17470 50 17475 70
rect 17205 10 17235 20
rect 17205 -10 17210 10
rect 17230 -10 17235 10
rect 17205 -40 17235 -10
rect 17320 15 17360 20
rect 17320 -15 17325 15
rect 17355 -15 17360 15
rect 17320 -20 17360 -15
rect 17445 -40 17475 50
rect 17505 120 17535 205
rect 17560 185 17600 190
rect 17560 155 17565 185
rect 17595 155 17600 185
rect 17560 150 17600 155
rect 17625 180 17655 205
rect 17625 160 17630 180
rect 17650 160 17655 180
rect 17505 100 17510 120
rect 17530 100 17535 120
rect 17505 70 17535 100
rect 17505 50 17510 70
rect 17530 50 17535 70
rect 17505 40 17535 50
rect 17565 120 17595 150
rect 17565 100 17570 120
rect 17590 100 17595 120
rect 17565 70 17595 100
rect 17565 50 17570 70
rect 17590 50 17595 70
rect 17565 40 17595 50
rect 17625 120 17655 160
rect 17690 185 17730 560
rect 17785 380 17815 630
rect 17875 900 17905 910
rect 17875 880 17880 900
rect 17900 880 17905 900
rect 17875 850 17905 880
rect 17875 830 17880 850
rect 17900 830 17905 850
rect 17875 800 17905 830
rect 17875 780 17880 800
rect 17900 780 17905 800
rect 17875 750 17905 780
rect 17875 730 17880 750
rect 17900 730 17905 750
rect 17875 700 17905 730
rect 17875 680 17880 700
rect 17900 680 17905 700
rect 17875 650 17905 680
rect 17875 630 17880 650
rect 17900 630 17905 650
rect 17875 620 17905 630
rect 17965 900 17995 910
rect 17965 880 17970 900
rect 17990 880 17995 900
rect 17965 850 17995 880
rect 17965 830 17970 850
rect 17990 830 17995 850
rect 17965 800 17995 830
rect 17965 780 17970 800
rect 17990 780 17995 800
rect 17965 750 17995 780
rect 17965 730 17970 750
rect 17990 730 17995 750
rect 17965 700 17995 730
rect 17965 680 17970 700
rect 17990 680 17995 700
rect 17965 650 17995 680
rect 17965 630 17970 650
rect 17990 630 17995 650
rect 17965 620 17995 630
rect 18055 900 18085 910
rect 18055 880 18060 900
rect 18080 880 18085 900
rect 18055 850 18085 880
rect 18055 830 18060 850
rect 18080 830 18085 850
rect 18055 800 18085 830
rect 18055 780 18060 800
rect 18080 780 18085 800
rect 18055 750 18085 780
rect 18055 730 18060 750
rect 18080 730 18085 750
rect 18055 700 18085 730
rect 18055 680 18060 700
rect 18080 680 18085 700
rect 18055 650 18085 680
rect 18055 630 18060 650
rect 18080 630 18085 650
rect 18055 620 18085 630
rect 18145 900 18175 910
rect 18145 880 18150 900
rect 18170 880 18175 900
rect 18145 850 18175 880
rect 18145 830 18150 850
rect 18170 830 18175 850
rect 18145 800 18175 830
rect 18145 780 18150 800
rect 18170 780 18175 800
rect 18145 750 18175 780
rect 18145 730 18150 750
rect 18170 730 18175 750
rect 18145 700 18175 730
rect 18145 680 18150 700
rect 18170 680 18175 700
rect 18145 650 18175 680
rect 18145 630 18150 650
rect 18170 630 18175 650
rect 18145 620 18175 630
rect 18235 900 18265 910
rect 18235 880 18240 900
rect 18260 880 18265 900
rect 18235 850 18265 880
rect 18235 830 18240 850
rect 18260 830 18265 850
rect 18235 800 18265 830
rect 18235 780 18240 800
rect 18260 780 18265 800
rect 18235 750 18265 780
rect 18235 730 18240 750
rect 18260 730 18265 750
rect 18235 700 18265 730
rect 18235 680 18240 700
rect 18260 680 18265 700
rect 18235 650 18265 680
rect 18235 630 18240 650
rect 18260 630 18265 650
rect 18235 620 18265 630
rect 18325 900 18355 910
rect 18325 880 18330 900
rect 18350 880 18355 900
rect 18325 850 18355 880
rect 18325 830 18330 850
rect 18350 830 18355 850
rect 18325 800 18355 830
rect 18325 780 18330 800
rect 18350 780 18355 800
rect 18325 750 18355 780
rect 18325 730 18330 750
rect 18350 730 18355 750
rect 18325 700 18355 730
rect 18325 680 18330 700
rect 18350 680 18355 700
rect 18325 650 18355 680
rect 18325 630 18330 650
rect 18350 630 18355 650
rect 18325 620 18355 630
rect 18415 900 18445 910
rect 18415 880 18420 900
rect 18440 880 18445 900
rect 18415 850 18445 880
rect 18415 830 18420 850
rect 18440 830 18445 850
rect 18415 800 18445 830
rect 18415 780 18420 800
rect 18440 780 18445 800
rect 18415 750 18445 780
rect 18415 730 18420 750
rect 18440 730 18445 750
rect 18415 700 18445 730
rect 18415 680 18420 700
rect 18440 680 18445 700
rect 18415 650 18445 680
rect 18415 630 18420 650
rect 18440 630 18445 650
rect 18415 620 18445 630
rect 18505 900 18535 910
rect 18505 880 18510 900
rect 18530 880 18535 900
rect 18505 850 18535 880
rect 18505 830 18510 850
rect 18530 830 18535 850
rect 18505 800 18535 830
rect 18505 780 18510 800
rect 18530 780 18535 800
rect 18505 750 18535 780
rect 18505 730 18510 750
rect 18530 730 18535 750
rect 18505 700 18535 730
rect 18505 680 18510 700
rect 18530 680 18535 700
rect 18505 650 18535 680
rect 18505 630 18510 650
rect 18530 630 18535 650
rect 17830 595 17865 600
rect 17860 565 17865 595
rect 17830 560 17865 565
rect 17915 595 17955 600
rect 17915 565 17920 595
rect 17950 565 17955 595
rect 17915 560 17955 565
rect 17970 545 17990 620
rect 18005 595 18045 600
rect 18005 565 18010 595
rect 18040 565 18045 595
rect 18005 560 18045 565
rect 18095 595 18135 600
rect 18095 565 18100 595
rect 18130 565 18135 595
rect 18095 560 18135 565
rect 17960 540 18000 545
rect 17960 510 17965 540
rect 17995 510 18000 540
rect 17960 505 18000 510
rect 18150 490 18170 620
rect 18185 595 18225 600
rect 18185 565 18190 595
rect 18220 565 18225 595
rect 18185 560 18225 565
rect 18275 595 18315 600
rect 18275 565 18280 595
rect 18310 565 18315 595
rect 18275 560 18315 565
rect 18140 485 18180 490
rect 18140 455 18145 485
rect 18175 455 18180 485
rect 18140 450 18180 455
rect 18330 435 18350 620
rect 18365 595 18405 600
rect 18365 565 18370 595
rect 18400 565 18405 595
rect 18365 560 18405 565
rect 18455 595 18490 600
rect 18455 565 18460 595
rect 18455 560 18490 565
rect 18320 430 18360 435
rect 18320 400 18325 430
rect 18355 400 18360 430
rect 18320 395 18360 400
rect 18505 380 18535 630
rect 18595 900 18625 910
rect 18595 880 18600 900
rect 18620 880 18625 900
rect 18595 850 18625 880
rect 18595 830 18600 850
rect 18620 830 18625 850
rect 18595 800 18625 830
rect 18595 780 18600 800
rect 18620 780 18625 800
rect 18595 750 18625 780
rect 18595 730 18600 750
rect 18620 730 18625 750
rect 18595 700 18625 730
rect 18910 900 18940 930
rect 18910 880 18915 900
rect 18935 880 18940 900
rect 18910 850 18940 880
rect 18910 830 18915 850
rect 18935 830 18940 850
rect 18910 800 18940 830
rect 18910 780 18915 800
rect 18935 780 18940 800
rect 18910 750 18940 780
rect 18910 730 18915 750
rect 18935 730 18940 750
rect 18910 720 18940 730
rect 18965 900 18995 1640
rect 19325 1100 19365 1105
rect 19325 1070 19330 1100
rect 19360 1070 19365 1100
rect 19015 1045 19055 1050
rect 19015 1015 19020 1045
rect 19050 1015 19055 1045
rect 19015 1005 19055 1015
rect 19015 975 19020 1005
rect 19050 975 19055 1005
rect 19015 965 19055 975
rect 19015 935 19020 965
rect 19050 935 19055 965
rect 19015 930 19055 935
rect 19075 1045 19115 1050
rect 19075 1015 19080 1045
rect 19110 1015 19115 1045
rect 19075 1005 19115 1015
rect 19075 975 19080 1005
rect 19110 975 19115 1005
rect 19075 965 19115 975
rect 19075 935 19080 965
rect 19110 935 19115 965
rect 19075 930 19115 935
rect 18965 880 18970 900
rect 18990 880 18995 900
rect 18965 850 18995 880
rect 18965 830 18970 850
rect 18990 830 18995 850
rect 18965 800 18995 830
rect 18965 780 18970 800
rect 18990 780 18995 800
rect 18965 750 18995 780
rect 18965 730 18970 750
rect 18990 730 18995 750
rect 18965 720 18995 730
rect 19020 900 19050 930
rect 19020 880 19025 900
rect 19045 880 19050 900
rect 19020 850 19050 880
rect 19020 830 19025 850
rect 19045 830 19050 850
rect 19020 800 19050 830
rect 19020 780 19025 800
rect 19045 780 19050 800
rect 19020 750 19050 780
rect 19020 730 19025 750
rect 19045 730 19050 750
rect 19020 720 19050 730
rect 19075 900 19105 930
rect 19075 880 19080 900
rect 19100 880 19105 900
rect 19075 850 19105 880
rect 19075 830 19080 850
rect 19100 830 19105 850
rect 19075 800 19105 830
rect 19075 780 19080 800
rect 19100 780 19105 800
rect 19075 750 19105 780
rect 19075 730 19080 750
rect 19100 730 19105 750
rect 19075 720 19105 730
rect 18595 680 18600 700
rect 18620 680 18625 700
rect 18595 650 18625 680
rect 18595 630 18600 650
rect 18620 630 18625 650
rect 18595 620 18625 630
rect 19000 635 19040 640
rect 19000 605 19005 635
rect 19035 605 19040 635
rect 19000 600 19040 605
rect 17780 375 17820 380
rect 17780 345 17785 375
rect 17815 345 17820 375
rect 17780 340 17820 345
rect 18500 375 18540 380
rect 18500 345 18505 375
rect 18535 345 18540 375
rect 18500 340 18540 345
rect 17940 320 17980 325
rect 17940 290 17945 320
rect 17975 290 17980 320
rect 17940 280 17980 290
rect 17940 250 17945 280
rect 17975 250 17980 280
rect 17940 240 17980 250
rect 17940 210 17945 240
rect 17975 210 17980 240
rect 17940 205 17980 210
rect 18060 320 18100 325
rect 18060 290 18065 320
rect 18095 290 18100 320
rect 18060 280 18100 290
rect 18060 250 18065 280
rect 18095 250 18100 280
rect 18060 240 18100 250
rect 18060 210 18065 240
rect 18095 210 18100 240
rect 18060 205 18100 210
rect 18180 320 18220 325
rect 18180 290 18185 320
rect 18215 290 18220 320
rect 18180 280 18220 290
rect 18180 250 18185 280
rect 18215 250 18220 280
rect 18180 240 18220 250
rect 18180 210 18185 240
rect 18215 210 18220 240
rect 18180 205 18220 210
rect 18300 320 18340 325
rect 18300 290 18305 320
rect 18335 290 18340 320
rect 18300 280 18340 290
rect 18300 250 18305 280
rect 18335 250 18340 280
rect 18300 240 18340 250
rect 18300 210 18305 240
rect 18335 210 18340 240
rect 18300 205 18340 210
rect 18420 320 18460 325
rect 18420 290 18425 320
rect 18455 290 18460 320
rect 18420 280 18460 290
rect 18420 250 18425 280
rect 18455 250 18460 280
rect 18420 240 18460 250
rect 18420 210 18425 240
rect 18455 210 18460 240
rect 18420 205 18460 210
rect 18540 320 18580 325
rect 18540 290 18545 320
rect 18575 290 18580 320
rect 18540 280 18580 290
rect 18540 250 18545 280
rect 18575 250 18580 280
rect 18540 240 18580 250
rect 18540 210 18545 240
rect 18575 210 18580 240
rect 18540 205 18580 210
rect 18660 320 18700 325
rect 18660 290 18665 320
rect 18695 290 18700 320
rect 18660 280 18700 290
rect 18660 250 18665 280
rect 18695 250 18700 280
rect 18660 240 18700 250
rect 18660 210 18665 240
rect 18695 210 18700 240
rect 18660 205 18700 210
rect 18780 320 18820 325
rect 18780 290 18785 320
rect 18815 290 18820 320
rect 18780 280 18820 290
rect 18780 250 18785 280
rect 18815 250 18820 280
rect 18780 240 18820 250
rect 18780 210 18785 240
rect 18815 210 18820 240
rect 18780 205 18820 210
rect 18900 320 18940 325
rect 18900 290 18905 320
rect 18935 290 18940 320
rect 18900 280 18940 290
rect 18900 250 18905 280
rect 18935 250 18940 280
rect 18900 240 18940 250
rect 18900 210 18905 240
rect 18935 210 18940 240
rect 18900 205 18940 210
rect 19020 320 19060 325
rect 19020 290 19025 320
rect 19055 290 19060 320
rect 19020 280 19060 290
rect 19020 250 19025 280
rect 19055 250 19060 280
rect 19020 240 19060 250
rect 19020 210 19025 240
rect 19055 210 19060 240
rect 19020 205 19060 210
rect 19140 320 19180 325
rect 19140 290 19145 320
rect 19175 290 19180 320
rect 19140 280 19180 290
rect 19140 250 19145 280
rect 19175 250 19180 280
rect 19140 240 19180 250
rect 19140 210 19145 240
rect 19175 210 19180 240
rect 19140 205 19180 210
rect 17690 155 17695 185
rect 17725 155 17730 185
rect 17690 150 17730 155
rect 17870 185 17910 190
rect 17870 155 17875 185
rect 17905 155 17910 185
rect 17870 150 17910 155
rect 17945 180 17975 205
rect 17945 160 17950 180
rect 17970 160 17975 180
rect 17625 100 17630 120
rect 17650 100 17655 120
rect 17625 70 17655 100
rect 17625 50 17630 70
rect 17650 50 17655 70
rect 17625 40 17655 50
rect 17535 10 17565 20
rect 17535 -10 17540 10
rect 17560 -10 17565 10
rect 17535 -40 17565 -10
rect 17080 -45 17120 -40
rect 17080 -75 17085 -45
rect 17115 -75 17120 -45
rect 17080 -85 17120 -75
rect 17080 -115 17085 -85
rect 17115 -115 17120 -85
rect 17080 -125 17120 -115
rect 17080 -155 17085 -125
rect 17115 -155 17120 -125
rect 17080 -160 17120 -155
rect 17200 -45 17240 -40
rect 17200 -75 17205 -45
rect 17235 -75 17240 -45
rect 17200 -85 17240 -75
rect 17200 -115 17205 -85
rect 17235 -115 17240 -85
rect 17200 -125 17240 -115
rect 17200 -155 17205 -125
rect 17235 -155 17240 -125
rect 17200 -160 17240 -155
rect 17440 -45 17480 -40
rect 17440 -75 17445 -45
rect 17475 -75 17480 -45
rect 17440 -85 17480 -75
rect 17440 -115 17445 -85
rect 17475 -115 17480 -85
rect 17440 -125 17480 -115
rect 17440 -155 17445 -125
rect 17475 -155 17480 -125
rect 17440 -160 17480 -155
rect 17530 -45 17570 -40
rect 17530 -75 17535 -45
rect 17565 -75 17570 -45
rect 17530 -85 17570 -75
rect 17530 -115 17535 -85
rect 17565 -115 17570 -85
rect 17530 -125 17570 -115
rect 17530 -155 17535 -125
rect 17565 -155 17570 -125
rect 17530 -160 17570 -155
rect 17007 -180 17037 -175
rect 17007 -215 17037 -210
rect 17090 -235 17110 -160
rect 16965 -245 16995 -235
rect 16965 -265 16970 -245
rect 16990 -265 16995 -245
rect 16965 -295 16995 -265
rect 16965 -315 16970 -295
rect 16990 -315 16995 -295
rect 16965 -345 16995 -315
rect 16965 -365 16970 -345
rect 16990 -365 16995 -345
rect 16965 -395 16995 -365
rect 16965 -415 16970 -395
rect 16990 -415 16995 -395
rect 16965 -445 16995 -415
rect 16965 -465 16970 -445
rect 16990 -465 16995 -445
rect 16965 -475 16995 -465
rect 17025 -245 17055 -235
rect 17025 -265 17030 -245
rect 17050 -265 17055 -245
rect 17025 -295 17055 -265
rect 17025 -315 17030 -295
rect 17050 -315 17055 -295
rect 17025 -345 17055 -315
rect 17025 -365 17030 -345
rect 17050 -365 17055 -345
rect 17025 -395 17055 -365
rect 17025 -415 17030 -395
rect 17050 -415 17055 -395
rect 17025 -445 17055 -415
rect 17025 -465 17030 -445
rect 17050 -465 17055 -445
rect 16315 -500 16355 -495
rect 16315 -530 16320 -500
rect 16350 -530 16355 -500
rect 16315 -535 16355 -530
rect 16325 -1995 16345 -535
rect 17025 -605 17055 -465
rect 17085 -245 17115 -235
rect 17085 -265 17090 -245
rect 17110 -265 17115 -245
rect 17085 -295 17115 -265
rect 17085 -315 17090 -295
rect 17110 -315 17115 -295
rect 17085 -345 17115 -315
rect 17085 -365 17090 -345
rect 17110 -365 17115 -345
rect 17560 -240 17600 -235
rect 17560 -270 17565 -240
rect 17595 -270 17600 -240
rect 17560 -280 17600 -270
rect 17560 -310 17565 -280
rect 17595 -310 17600 -280
rect 17560 -320 17600 -310
rect 17560 -350 17565 -320
rect 17595 -350 17600 -320
rect 17560 -355 17600 -350
rect 17085 -395 17115 -365
rect 17085 -415 17090 -395
rect 17110 -415 17115 -395
rect 17085 -445 17115 -415
rect 17085 -465 17090 -445
rect 17110 -465 17115 -445
rect 17085 -475 17115 -465
rect 17075 -500 17105 -495
rect 17075 -535 17105 -530
rect 16530 -610 16570 -605
rect 16530 -640 16535 -610
rect 16565 -640 16570 -610
rect 16530 -645 16570 -640
rect 17020 -610 17060 -605
rect 17020 -640 17025 -610
rect 17055 -640 17060 -610
rect 17020 -645 17060 -640
rect 16535 -810 16565 -645
rect 16620 -665 16660 -660
rect 16620 -695 16625 -665
rect 16655 -695 16660 -665
rect 16620 -705 16660 -695
rect 16620 -735 16625 -705
rect 16655 -735 16660 -705
rect 16620 -745 16660 -735
rect 16620 -775 16625 -745
rect 16655 -775 16660 -745
rect 16620 -780 16660 -775
rect 16740 -665 16780 -660
rect 16740 -695 16745 -665
rect 16775 -695 16780 -665
rect 16740 -705 16780 -695
rect 16740 -735 16745 -705
rect 16775 -735 16780 -705
rect 16740 -745 16780 -735
rect 16740 -775 16745 -745
rect 16775 -775 16780 -745
rect 16740 -780 16780 -775
rect 16860 -665 16900 -660
rect 16860 -695 16865 -665
rect 16895 -695 16900 -665
rect 16860 -705 16900 -695
rect 16860 -735 16865 -705
rect 16895 -735 16900 -705
rect 16860 -745 16900 -735
rect 16860 -775 16865 -745
rect 16895 -775 16900 -745
rect 16860 -780 16900 -775
rect 16980 -665 17020 -660
rect 16980 -695 16985 -665
rect 17015 -695 17020 -665
rect 16980 -705 17020 -695
rect 16980 -735 16985 -705
rect 17015 -735 17020 -705
rect 16980 -745 17020 -735
rect 16980 -775 16985 -745
rect 17015 -775 17020 -745
rect 16980 -780 17020 -775
rect 17300 -665 17340 -660
rect 17300 -695 17305 -665
rect 17335 -695 17340 -665
rect 17300 -705 17340 -695
rect 17300 -735 17305 -705
rect 17335 -735 17340 -705
rect 17300 -745 17340 -735
rect 17300 -775 17305 -745
rect 17335 -775 17340 -745
rect 17300 -780 17340 -775
rect 17420 -665 17460 -660
rect 17420 -695 17425 -665
rect 17455 -695 17460 -665
rect 17420 -705 17460 -695
rect 17420 -735 17425 -705
rect 17455 -735 17460 -705
rect 17420 -745 17460 -735
rect 17420 -775 17425 -745
rect 17455 -775 17460 -745
rect 17420 -780 17460 -775
rect 17540 -665 17580 -660
rect 17540 -695 17545 -665
rect 17575 -695 17580 -665
rect 17540 -705 17580 -695
rect 17540 -735 17545 -705
rect 17575 -735 17580 -705
rect 17540 -745 17580 -735
rect 17540 -775 17545 -745
rect 17575 -775 17580 -745
rect 17540 -780 17580 -775
rect 17695 -765 17725 150
rect 17695 -785 17700 -765
rect 17720 -785 17725 -765
rect 17695 -795 17725 -785
rect 17740 -240 17860 -235
rect 17740 -270 17745 -240
rect 17775 -270 17785 -240
rect 17815 -270 17825 -240
rect 17855 -270 17860 -240
rect 17740 -280 17860 -270
rect 17740 -310 17745 -280
rect 17775 -310 17785 -280
rect 17815 -310 17825 -280
rect 17855 -310 17860 -280
rect 17740 -320 17860 -310
rect 17740 -350 17745 -320
rect 17775 -350 17785 -320
rect 17815 -350 17825 -320
rect 17855 -350 17860 -320
rect 16535 -830 16540 -810
rect 16560 -830 16565 -810
rect 16535 -860 16565 -830
rect 16535 -880 16540 -860
rect 16560 -880 16565 -860
rect 16535 -910 16565 -880
rect 16535 -930 16540 -910
rect 16560 -930 16565 -910
rect 16535 -960 16565 -930
rect 16535 -980 16540 -960
rect 16560 -980 16565 -960
rect 16535 -1010 16565 -980
rect 16535 -1030 16540 -1010
rect 16560 -1030 16565 -1010
rect 16535 -1040 16565 -1030
rect 17110 -1065 17150 -1060
rect 17110 -1095 17115 -1065
rect 17145 -1095 17150 -1065
rect 17110 -1105 17150 -1095
rect 17110 -1135 17115 -1105
rect 17145 -1135 17150 -1105
rect 17110 -1145 17150 -1135
rect 17110 -1175 17115 -1145
rect 17145 -1175 17150 -1145
rect 17110 -1180 17150 -1175
rect 17740 -1065 17860 -350
rect 17875 -765 17905 150
rect 17945 120 17975 160
rect 18000 185 18040 190
rect 18000 155 18005 185
rect 18035 155 18040 185
rect 18000 150 18040 155
rect 17945 100 17950 120
rect 17970 100 17975 120
rect 17945 70 17975 100
rect 17945 50 17950 70
rect 17970 50 17975 70
rect 17945 40 17975 50
rect 18005 120 18035 150
rect 18005 100 18010 120
rect 18030 100 18035 120
rect 18005 70 18035 100
rect 18005 50 18010 70
rect 18030 50 18035 70
rect 18005 40 18035 50
rect 18065 120 18095 205
rect 18065 100 18070 120
rect 18090 100 18095 120
rect 18065 70 18095 100
rect 18065 50 18070 70
rect 18090 50 18095 70
rect 18065 40 18095 50
rect 18125 120 18155 130
rect 18125 100 18130 120
rect 18150 100 18155 120
rect 18125 70 18155 100
rect 18125 50 18130 70
rect 18150 50 18155 70
rect 18035 10 18065 20
rect 18035 -10 18040 10
rect 18060 -10 18065 10
rect 18035 -40 18065 -10
rect 18125 -40 18155 50
rect 18185 120 18215 205
rect 18185 100 18190 120
rect 18210 100 18215 120
rect 18185 70 18215 100
rect 18185 50 18190 70
rect 18210 50 18215 70
rect 18185 40 18215 50
rect 18245 120 18275 130
rect 18245 100 18250 120
rect 18270 100 18275 120
rect 18245 70 18275 100
rect 18245 50 18250 70
rect 18270 50 18275 70
rect 18245 20 18275 50
rect 18305 120 18335 205
rect 18360 185 18400 190
rect 18360 155 18365 185
rect 18395 155 18400 185
rect 18360 150 18400 155
rect 18305 100 18310 120
rect 18330 100 18335 120
rect 18305 70 18335 100
rect 18305 50 18310 70
rect 18330 50 18335 70
rect 18305 40 18335 50
rect 18365 120 18395 150
rect 18365 100 18370 120
rect 18390 100 18395 120
rect 18365 70 18395 100
rect 18365 50 18370 70
rect 18390 50 18395 70
rect 18365 40 18395 50
rect 18425 120 18455 205
rect 18425 100 18430 120
rect 18450 100 18455 120
rect 18425 70 18455 100
rect 18425 50 18430 70
rect 18450 50 18455 70
rect 18425 40 18455 50
rect 18485 120 18515 130
rect 18485 100 18490 120
rect 18510 100 18515 120
rect 18485 70 18515 100
rect 18485 50 18490 70
rect 18510 50 18515 70
rect 18240 15 18280 20
rect 18240 -15 18245 15
rect 18275 -15 18280 15
rect 18240 -20 18280 -15
rect 18365 10 18395 20
rect 18365 -10 18370 10
rect 18390 -10 18395 10
rect 18365 -40 18395 -10
rect 18485 -40 18515 50
rect 18545 120 18575 205
rect 18545 100 18550 120
rect 18570 100 18575 120
rect 18545 70 18575 100
rect 18545 50 18550 70
rect 18570 50 18575 70
rect 18545 40 18575 50
rect 18605 120 18635 130
rect 18605 100 18610 120
rect 18630 100 18635 120
rect 18605 70 18635 100
rect 18605 50 18610 70
rect 18630 50 18635 70
rect 18605 20 18635 50
rect 18665 120 18695 205
rect 18720 185 18760 190
rect 18720 155 18725 185
rect 18755 155 18760 185
rect 18720 150 18760 155
rect 18665 100 18670 120
rect 18690 100 18695 120
rect 18665 70 18695 100
rect 18665 50 18670 70
rect 18690 50 18695 70
rect 18665 40 18695 50
rect 18725 120 18755 150
rect 18725 100 18730 120
rect 18750 100 18755 120
rect 18725 70 18755 100
rect 18725 50 18730 70
rect 18750 50 18755 70
rect 18725 40 18755 50
rect 18785 120 18815 205
rect 18785 100 18790 120
rect 18810 100 18815 120
rect 18785 70 18815 100
rect 18785 50 18790 70
rect 18810 50 18815 70
rect 18785 40 18815 50
rect 18845 120 18875 130
rect 18845 100 18850 120
rect 18870 100 18875 120
rect 18845 70 18875 100
rect 18845 50 18850 70
rect 18870 50 18875 70
rect 18600 15 18640 20
rect 18600 -15 18605 15
rect 18635 -15 18640 15
rect 18600 -20 18640 -15
rect 18725 10 18755 20
rect 18725 -10 18730 10
rect 18750 -10 18755 10
rect 18030 -45 18070 -40
rect 18030 -75 18035 -45
rect 18065 -75 18070 -45
rect 18030 -80 18070 -75
rect 18120 -45 18160 -40
rect 18120 -75 18125 -45
rect 18155 -75 18160 -45
rect 18120 -80 18160 -75
rect 18360 -45 18400 -40
rect 18360 -75 18365 -45
rect 18395 -75 18400 -45
rect 18360 -80 18400 -75
rect 18480 -45 18520 -40
rect 18480 -75 18485 -45
rect 18515 -75 18520 -45
rect 18480 -80 18520 -75
rect 18000 -240 18040 -235
rect 18000 -270 18005 -240
rect 18035 -270 18040 -240
rect 18000 -280 18040 -270
rect 18000 -310 18005 -280
rect 18035 -310 18040 -280
rect 18000 -320 18040 -310
rect 18000 -350 18005 -320
rect 18035 -350 18040 -320
rect 18000 -355 18040 -350
rect 18485 -245 18515 -80
rect 18563 -180 18593 -175
rect 18563 -215 18593 -210
rect 18610 -235 18630 -20
rect 18725 -40 18755 -10
rect 18845 -40 18875 50
rect 18905 120 18935 205
rect 18905 100 18910 120
rect 18930 100 18935 120
rect 18905 70 18935 100
rect 18905 50 18910 70
rect 18930 50 18935 70
rect 18905 40 18935 50
rect 18965 120 18995 130
rect 18965 100 18970 120
rect 18990 100 18995 120
rect 18965 70 18995 100
rect 18965 50 18970 70
rect 18990 50 18995 70
rect 18965 20 18995 50
rect 19025 120 19055 205
rect 19080 185 19120 190
rect 19080 155 19085 185
rect 19115 155 19120 185
rect 19080 150 19120 155
rect 19145 180 19175 205
rect 19145 160 19150 180
rect 19170 160 19175 180
rect 19025 100 19030 120
rect 19050 100 19055 120
rect 19025 70 19055 100
rect 19025 50 19030 70
rect 19050 50 19055 70
rect 19025 40 19055 50
rect 19085 120 19115 150
rect 19085 100 19090 120
rect 19110 100 19115 120
rect 19085 70 19115 100
rect 19085 50 19090 70
rect 19110 50 19115 70
rect 19085 40 19115 50
rect 19145 120 19175 160
rect 19145 100 19150 120
rect 19170 100 19175 120
rect 19145 70 19175 100
rect 19145 50 19150 70
rect 19170 50 19175 70
rect 19145 40 19175 50
rect 18960 15 19000 20
rect 18960 -15 18965 15
rect 18995 -15 19000 15
rect 18960 -20 19000 -15
rect 19055 5 19085 15
rect 19055 -15 19060 5
rect 19080 -15 19085 5
rect 19055 -40 19085 -15
rect 18720 -45 18760 -40
rect 18720 -75 18725 -45
rect 18755 -75 18760 -45
rect 18720 -80 18760 -75
rect 18840 -45 18880 -40
rect 18840 -75 18845 -45
rect 18875 -75 18880 -45
rect 18840 -80 18880 -75
rect 19050 -45 19130 -40
rect 19050 -75 19055 -45
rect 19085 -75 19095 -45
rect 19125 -75 19130 -45
rect 19050 -80 19130 -75
rect 18485 -265 18490 -245
rect 18510 -265 18515 -245
rect 18485 -295 18515 -265
rect 18485 -315 18490 -295
rect 18510 -315 18515 -295
rect 18485 -345 18515 -315
rect 18485 -365 18490 -345
rect 18510 -365 18515 -345
rect 18485 -395 18515 -365
rect 18485 -415 18490 -395
rect 18510 -415 18515 -395
rect 18485 -445 18515 -415
rect 18485 -465 18490 -445
rect 18510 -465 18515 -445
rect 18485 -475 18515 -465
rect 18545 -245 18575 -235
rect 18545 -265 18550 -245
rect 18570 -265 18575 -245
rect 18545 -295 18575 -265
rect 18545 -315 18550 -295
rect 18570 -315 18575 -295
rect 18545 -345 18575 -315
rect 18545 -365 18550 -345
rect 18570 -365 18575 -345
rect 18545 -395 18575 -365
rect 18545 -415 18550 -395
rect 18570 -415 18575 -395
rect 18545 -445 18575 -415
rect 18545 -465 18550 -445
rect 18570 -465 18575 -445
rect 18440 -500 18470 -495
rect 18440 -535 18470 -530
rect 18545 -605 18575 -465
rect 18605 -245 18635 -235
rect 18605 -265 18610 -245
rect 18630 -265 18635 -245
rect 18605 -295 18635 -265
rect 18605 -315 18610 -295
rect 18630 -315 18635 -295
rect 18605 -345 18635 -315
rect 18605 -365 18610 -345
rect 18630 -365 18635 -345
rect 18605 -395 18635 -365
rect 18605 -415 18610 -395
rect 18630 -415 18635 -395
rect 18605 -445 18635 -415
rect 18605 -465 18610 -445
rect 18630 -465 18635 -445
rect 18605 -475 18635 -465
rect 18540 -610 18580 -605
rect 18540 -640 18545 -610
rect 18575 -640 18580 -610
rect 18540 -645 18580 -640
rect 19030 -610 19070 -605
rect 19030 -640 19035 -610
rect 19065 -640 19070 -610
rect 19030 -645 19070 -640
rect 17875 -785 17880 -765
rect 17900 -785 17905 -765
rect 18020 -665 18060 -660
rect 18020 -695 18025 -665
rect 18055 -695 18060 -665
rect 18020 -705 18060 -695
rect 18020 -735 18025 -705
rect 18055 -735 18060 -705
rect 18020 -745 18060 -735
rect 18020 -775 18025 -745
rect 18055 -775 18060 -745
rect 18020 -780 18060 -775
rect 18140 -665 18180 -660
rect 18140 -695 18145 -665
rect 18175 -695 18180 -665
rect 18140 -705 18180 -695
rect 18140 -735 18145 -705
rect 18175 -735 18180 -705
rect 18140 -745 18180 -735
rect 18140 -775 18145 -745
rect 18175 -775 18180 -745
rect 18140 -780 18180 -775
rect 18260 -665 18300 -660
rect 18260 -695 18265 -665
rect 18295 -695 18300 -665
rect 18260 -705 18300 -695
rect 18260 -735 18265 -705
rect 18295 -735 18300 -705
rect 18260 -745 18300 -735
rect 18260 -775 18265 -745
rect 18295 -775 18300 -745
rect 18260 -780 18300 -775
rect 18580 -665 18620 -660
rect 18580 -695 18585 -665
rect 18615 -695 18620 -665
rect 18580 -705 18620 -695
rect 18580 -735 18585 -705
rect 18615 -735 18620 -705
rect 18580 -745 18620 -735
rect 18580 -775 18585 -745
rect 18615 -775 18620 -745
rect 18580 -780 18620 -775
rect 18700 -665 18740 -660
rect 18700 -695 18705 -665
rect 18735 -695 18740 -665
rect 18700 -705 18740 -695
rect 18700 -735 18705 -705
rect 18735 -735 18740 -705
rect 18700 -745 18740 -735
rect 18700 -775 18705 -745
rect 18735 -775 18740 -745
rect 18700 -780 18740 -775
rect 18820 -665 18860 -660
rect 18820 -695 18825 -665
rect 18855 -695 18860 -665
rect 18820 -705 18860 -695
rect 18820 -735 18825 -705
rect 18855 -735 18860 -705
rect 18820 -745 18860 -735
rect 18820 -775 18825 -745
rect 18855 -775 18860 -745
rect 18820 -780 18860 -775
rect 18940 -665 18980 -660
rect 18940 -695 18945 -665
rect 18975 -695 18980 -665
rect 18940 -705 18980 -695
rect 18940 -735 18945 -705
rect 18975 -735 18980 -705
rect 18940 -745 18980 -735
rect 18940 -775 18945 -745
rect 18975 -775 18980 -745
rect 19040 -760 19060 -645
rect 18940 -780 18980 -775
rect 19030 -770 19070 -760
rect 17875 -795 17905 -785
rect 19030 -790 19040 -770
rect 19060 -790 19070 -770
rect 19030 -800 19070 -790
rect 17740 -1095 17745 -1065
rect 17775 -1095 17785 -1065
rect 17815 -1095 17825 -1065
rect 17855 -1095 17860 -1065
rect 17740 -1105 17860 -1095
rect 17740 -1135 17745 -1105
rect 17775 -1135 17785 -1105
rect 17815 -1135 17825 -1105
rect 17855 -1135 17860 -1105
rect 17740 -1145 17860 -1135
rect 17740 -1175 17745 -1145
rect 17775 -1175 17785 -1145
rect 17815 -1175 17825 -1145
rect 17855 -1175 17860 -1145
rect 17740 -1180 17860 -1175
rect 18450 -1065 18490 -1060
rect 18450 -1095 18455 -1065
rect 18485 -1095 18490 -1065
rect 18450 -1105 18490 -1095
rect 18450 -1135 18455 -1105
rect 18485 -1135 18490 -1105
rect 18450 -1145 18490 -1135
rect 18450 -1175 18455 -1145
rect 18485 -1175 18490 -1145
rect 18450 -1180 18490 -1175
rect 16740 -1200 16780 -1195
rect 16740 -1230 16745 -1200
rect 16775 -1230 16780 -1200
rect 16740 -1235 16780 -1230
rect 16820 -1200 16860 -1195
rect 16820 -1230 16825 -1200
rect 16855 -1230 16860 -1200
rect 16820 -1235 16860 -1230
rect 16900 -1200 16940 -1195
rect 16900 -1230 16905 -1200
rect 16935 -1230 16940 -1200
rect 16900 -1235 16940 -1230
rect 16980 -1200 17020 -1195
rect 16980 -1230 16985 -1200
rect 17015 -1230 17020 -1200
rect 16980 -1235 17020 -1230
rect 17060 -1200 17100 -1195
rect 17060 -1230 17065 -1200
rect 17095 -1230 17100 -1200
rect 17060 -1235 17100 -1230
rect 17140 -1200 17180 -1195
rect 17140 -1230 17145 -1200
rect 17175 -1230 17180 -1200
rect 17140 -1235 17180 -1230
rect 17220 -1200 17260 -1195
rect 17220 -1230 17225 -1200
rect 17255 -1230 17260 -1200
rect 17220 -1235 17260 -1230
rect 17300 -1200 17340 -1195
rect 17300 -1230 17305 -1200
rect 17335 -1230 17340 -1200
rect 17300 -1235 17340 -1230
rect 17380 -1200 17420 -1195
rect 17380 -1230 17385 -1200
rect 17415 -1230 17420 -1200
rect 17380 -1235 17420 -1230
rect 17460 -1200 17500 -1195
rect 17460 -1230 17465 -1200
rect 17495 -1230 17500 -1200
rect 17460 -1235 17500 -1230
rect 17540 -1200 17580 -1195
rect 17540 -1230 17545 -1200
rect 17575 -1230 17580 -1200
rect 17540 -1235 17580 -1230
rect 17620 -1200 17660 -1195
rect 17620 -1230 17625 -1200
rect 17655 -1230 17660 -1200
rect 17620 -1235 17660 -1230
rect 17700 -1200 17740 -1195
rect 17700 -1230 17705 -1200
rect 17735 -1230 17740 -1200
rect 17700 -1235 17740 -1230
rect 17780 -1200 17820 -1195
rect 17780 -1230 17785 -1200
rect 17815 -1230 17820 -1200
rect 17780 -1235 17820 -1230
rect 17860 -1200 17900 -1195
rect 17860 -1230 17865 -1200
rect 17895 -1230 17900 -1200
rect 17860 -1235 17900 -1230
rect 17940 -1200 17980 -1195
rect 17940 -1230 17945 -1200
rect 17975 -1230 17980 -1200
rect 17940 -1235 17980 -1230
rect 18020 -1200 18060 -1195
rect 18020 -1230 18025 -1200
rect 18055 -1230 18060 -1200
rect 18020 -1235 18060 -1230
rect 18100 -1200 18140 -1195
rect 18100 -1230 18105 -1200
rect 18135 -1230 18140 -1200
rect 18100 -1235 18140 -1230
rect 18180 -1200 18220 -1195
rect 18180 -1230 18185 -1200
rect 18215 -1230 18220 -1200
rect 18180 -1235 18220 -1230
rect 18260 -1200 18300 -1195
rect 18260 -1230 18265 -1200
rect 18295 -1230 18300 -1200
rect 18260 -1235 18300 -1230
rect 18340 -1200 18380 -1195
rect 18340 -1230 18345 -1200
rect 18375 -1230 18380 -1200
rect 18340 -1235 18380 -1230
rect 18420 -1200 18460 -1195
rect 18420 -1230 18425 -1200
rect 18455 -1230 18460 -1200
rect 18420 -1235 18460 -1230
rect 18500 -1200 18540 -1195
rect 18500 -1230 18505 -1200
rect 18535 -1230 18540 -1200
rect 18500 -1235 18540 -1230
rect 18580 -1200 18620 -1195
rect 18580 -1230 18585 -1200
rect 18615 -1230 18620 -1200
rect 18580 -1235 18620 -1230
rect 18660 -1200 18700 -1195
rect 18660 -1230 18665 -1200
rect 18695 -1230 18700 -1200
rect 18660 -1235 18700 -1230
rect 18740 -1200 18780 -1195
rect 18740 -1230 18745 -1200
rect 18775 -1230 18780 -1200
rect 18740 -1235 18780 -1230
rect 18895 -1265 18935 -1260
rect 16700 -1285 16740 -1280
rect 16700 -1315 16705 -1285
rect 16735 -1315 16740 -1285
rect 16700 -1320 16740 -1315
rect 18895 -1295 18900 -1265
rect 18930 -1295 18935 -1265
rect 18895 -1305 18935 -1295
rect 18895 -1335 18900 -1305
rect 18930 -1335 18935 -1305
rect 18895 -1340 18935 -1335
rect 16655 -1385 16695 -1380
rect 16655 -1415 16660 -1385
rect 16690 -1415 16695 -1385
rect 16655 -1420 16695 -1415
rect 16765 -1385 16805 -1380
rect 16765 -1415 16770 -1385
rect 16800 -1415 16805 -1385
rect 16765 -1420 16805 -1415
rect 17300 -1385 17340 -1380
rect 17300 -1415 17305 -1385
rect 17335 -1415 17340 -1385
rect 17300 -1420 17340 -1415
rect 17780 -1385 17820 -1380
rect 17780 -1415 17785 -1385
rect 17815 -1415 17820 -1385
rect 17780 -1420 17820 -1415
rect 18315 -1385 18355 -1380
rect 18315 -1415 18320 -1385
rect 18350 -1415 18355 -1385
rect 18315 -1420 18355 -1415
rect 16600 -1440 16640 -1435
rect 16600 -1470 16605 -1440
rect 16635 -1470 16640 -1440
rect 16600 -1480 16640 -1470
rect 16600 -1510 16605 -1480
rect 16635 -1510 16640 -1480
rect 16600 -1520 16640 -1510
rect 16600 -1550 16605 -1520
rect 16635 -1550 16640 -1520
rect 16600 -1555 16640 -1550
rect 16660 -1525 16690 -1420
rect 16660 -1545 16665 -1525
rect 16685 -1545 16690 -1525
rect 16660 -1555 16690 -1545
rect 16710 -1440 16750 -1435
rect 16710 -1470 16715 -1440
rect 16745 -1470 16750 -1440
rect 16710 -1480 16750 -1470
rect 16710 -1510 16715 -1480
rect 16745 -1510 16750 -1480
rect 16710 -1520 16750 -1510
rect 16710 -1550 16715 -1520
rect 16745 -1550 16750 -1520
rect 16710 -1555 16750 -1550
rect 16770 -1525 16800 -1420
rect 16770 -1545 16775 -1525
rect 16795 -1545 16800 -1525
rect 16770 -1555 16800 -1545
rect 16820 -1440 16860 -1435
rect 16820 -1470 16825 -1440
rect 16855 -1470 16860 -1440
rect 16820 -1480 16860 -1470
rect 16820 -1510 16825 -1480
rect 16855 -1510 16860 -1480
rect 16820 -1520 16860 -1510
rect 16820 -1550 16825 -1520
rect 16855 -1550 16860 -1520
rect 16820 -1555 16860 -1550
rect 16880 -1440 16920 -1435
rect 16880 -1470 16885 -1440
rect 16915 -1470 16920 -1440
rect 16880 -1480 16920 -1470
rect 16880 -1510 16885 -1480
rect 16915 -1510 16920 -1480
rect 16880 -1520 16920 -1510
rect 16880 -1550 16885 -1520
rect 16915 -1550 16920 -1520
rect 16880 -1555 16920 -1550
rect 17025 -1440 17065 -1435
rect 17025 -1470 17030 -1440
rect 17060 -1470 17065 -1440
rect 17025 -1480 17065 -1470
rect 17025 -1510 17030 -1480
rect 17060 -1510 17065 -1480
rect 17025 -1520 17065 -1510
rect 17025 -1550 17030 -1520
rect 17060 -1550 17065 -1520
rect 17025 -1555 17065 -1550
rect 17135 -1440 17175 -1435
rect 17135 -1470 17140 -1440
rect 17170 -1470 17175 -1440
rect 17135 -1480 17175 -1470
rect 17135 -1510 17140 -1480
rect 17170 -1510 17175 -1480
rect 17135 -1520 17175 -1510
rect 17135 -1550 17140 -1520
rect 17170 -1550 17175 -1520
rect 17135 -1555 17175 -1550
rect 17245 -1440 17285 -1435
rect 17245 -1470 17250 -1440
rect 17280 -1470 17285 -1440
rect 17245 -1480 17285 -1470
rect 17245 -1510 17250 -1480
rect 17280 -1510 17285 -1480
rect 17245 -1520 17285 -1510
rect 17245 -1550 17250 -1520
rect 17280 -1550 17285 -1520
rect 17245 -1555 17285 -1550
rect 17305 -1525 17335 -1420
rect 17305 -1545 17310 -1525
rect 17330 -1545 17335 -1525
rect 17305 -1555 17335 -1545
rect 17355 -1440 17395 -1435
rect 17355 -1470 17360 -1440
rect 17390 -1470 17395 -1440
rect 17355 -1480 17395 -1470
rect 17355 -1510 17360 -1480
rect 17390 -1510 17395 -1480
rect 17355 -1520 17395 -1510
rect 17355 -1550 17360 -1520
rect 17390 -1550 17395 -1520
rect 17355 -1555 17395 -1550
rect 17465 -1440 17505 -1435
rect 17465 -1470 17470 -1440
rect 17500 -1470 17505 -1440
rect 17465 -1480 17505 -1470
rect 17465 -1510 17470 -1480
rect 17500 -1510 17505 -1480
rect 17465 -1520 17505 -1510
rect 17465 -1550 17470 -1520
rect 17500 -1550 17505 -1520
rect 17465 -1555 17505 -1550
rect 17615 -1440 17655 -1435
rect 17615 -1470 17620 -1440
rect 17650 -1470 17655 -1440
rect 17615 -1480 17655 -1470
rect 17615 -1510 17620 -1480
rect 17650 -1510 17655 -1480
rect 17615 -1520 17655 -1510
rect 17615 -1550 17620 -1520
rect 17650 -1550 17655 -1520
rect 17615 -1555 17655 -1550
rect 17725 -1440 17765 -1435
rect 17725 -1470 17730 -1440
rect 17760 -1470 17765 -1440
rect 17725 -1480 17765 -1470
rect 17725 -1510 17730 -1480
rect 17760 -1510 17765 -1480
rect 17725 -1520 17765 -1510
rect 17725 -1550 17730 -1520
rect 17760 -1550 17765 -1520
rect 17725 -1555 17765 -1550
rect 17785 -1525 17815 -1420
rect 17785 -1545 17790 -1525
rect 17810 -1545 17815 -1525
rect 17785 -1555 17815 -1545
rect 17835 -1440 17875 -1435
rect 17835 -1470 17840 -1440
rect 17870 -1470 17875 -1440
rect 17835 -1480 17875 -1470
rect 17835 -1510 17840 -1480
rect 17870 -1510 17875 -1480
rect 17835 -1520 17875 -1510
rect 17835 -1550 17840 -1520
rect 17870 -1550 17875 -1520
rect 17835 -1555 17875 -1550
rect 17945 -1440 17985 -1435
rect 17945 -1470 17950 -1440
rect 17980 -1470 17985 -1440
rect 17945 -1480 17985 -1470
rect 17945 -1510 17950 -1480
rect 17980 -1510 17985 -1480
rect 17945 -1520 17985 -1510
rect 17945 -1550 17950 -1520
rect 17980 -1550 17985 -1520
rect 17945 -1555 17985 -1550
rect 18005 -1440 18045 -1435
rect 18005 -1470 18010 -1440
rect 18040 -1470 18045 -1440
rect 18005 -1480 18045 -1470
rect 18005 -1510 18010 -1480
rect 18040 -1510 18045 -1480
rect 18005 -1520 18045 -1510
rect 18005 -1550 18010 -1520
rect 18040 -1550 18045 -1520
rect 18005 -1555 18045 -1550
rect 18150 -1440 18190 -1435
rect 18150 -1470 18155 -1440
rect 18185 -1470 18190 -1440
rect 18150 -1480 18190 -1470
rect 18150 -1510 18155 -1480
rect 18185 -1510 18190 -1480
rect 18150 -1520 18190 -1510
rect 18150 -1550 18155 -1520
rect 18185 -1550 18190 -1520
rect 18150 -1555 18190 -1550
rect 18260 -1440 18300 -1435
rect 18260 -1470 18265 -1440
rect 18295 -1470 18300 -1440
rect 18260 -1480 18300 -1470
rect 18260 -1510 18265 -1480
rect 18295 -1510 18300 -1480
rect 18260 -1520 18300 -1510
rect 18260 -1550 18265 -1520
rect 18295 -1550 18300 -1520
rect 18260 -1555 18300 -1550
rect 18320 -1525 18350 -1420
rect 18320 -1545 18325 -1525
rect 18345 -1545 18350 -1525
rect 18320 -1555 18350 -1545
rect 18370 -1440 18410 -1435
rect 18370 -1470 18375 -1440
rect 18405 -1470 18410 -1440
rect 18370 -1480 18410 -1470
rect 18370 -1510 18375 -1480
rect 18405 -1510 18410 -1480
rect 18370 -1520 18410 -1510
rect 18370 -1550 18375 -1520
rect 18405 -1550 18410 -1520
rect 18370 -1555 18410 -1550
rect 18480 -1440 18520 -1435
rect 18480 -1470 18485 -1440
rect 18515 -1470 18520 -1440
rect 18480 -1480 18520 -1470
rect 18480 -1510 18485 -1480
rect 18515 -1510 18520 -1480
rect 18480 -1520 18520 -1510
rect 18480 -1550 18485 -1520
rect 18515 -1550 18520 -1520
rect 18480 -1555 18520 -1550
rect 18590 -1440 18630 -1435
rect 18590 -1470 18595 -1440
rect 18625 -1470 18630 -1440
rect 18590 -1480 18630 -1470
rect 18590 -1510 18595 -1480
rect 18625 -1510 18630 -1480
rect 18590 -1520 18630 -1510
rect 18590 -1550 18595 -1520
rect 18625 -1550 18630 -1520
rect 18590 -1555 18630 -1550
rect 17195 -1585 17225 -1575
rect 17195 -1605 17200 -1585
rect 17220 -1605 17225 -1585
rect 17195 -1635 17225 -1605
rect 17195 -1655 17200 -1635
rect 17220 -1655 17225 -1635
rect 17195 -1685 17225 -1655
rect 17415 -1585 17445 -1575
rect 17415 -1605 17420 -1585
rect 17440 -1605 17445 -1585
rect 17415 -1635 17445 -1605
rect 17415 -1655 17420 -1635
rect 17440 -1655 17445 -1635
rect 17415 -1685 17445 -1655
rect 18210 -1585 18240 -1575
rect 18210 -1605 18215 -1585
rect 18235 -1605 18240 -1585
rect 18210 -1635 18240 -1605
rect 18210 -1655 18215 -1635
rect 18235 -1655 18240 -1635
rect 18210 -1685 18240 -1655
rect 18430 -1585 18460 -1575
rect 18430 -1605 18435 -1585
rect 18455 -1605 18460 -1585
rect 18430 -1635 18460 -1605
rect 18430 -1655 18435 -1635
rect 18455 -1655 18460 -1635
rect 18430 -1685 18460 -1655
rect 16765 -1695 16805 -1685
rect 16765 -1715 16775 -1695
rect 16795 -1715 16805 -1695
rect 16765 -1725 16805 -1715
rect 17080 -1695 17120 -1685
rect 17080 -1715 17090 -1695
rect 17110 -1715 17120 -1695
rect 17080 -1725 17120 -1715
rect 17190 -1690 17230 -1685
rect 17190 -1720 17195 -1690
rect 17225 -1720 17230 -1690
rect 16775 -1850 16795 -1725
rect 17090 -1740 17110 -1725
rect 17080 -1745 17120 -1740
rect 17080 -1775 17085 -1745
rect 17115 -1775 17120 -1745
rect 17080 -1780 17120 -1775
rect 17190 -1800 17230 -1720
rect 17300 -1695 17340 -1685
rect 17300 -1715 17310 -1695
rect 17330 -1715 17340 -1695
rect 17300 -1725 17340 -1715
rect 17410 -1690 17450 -1685
rect 17410 -1720 17415 -1690
rect 17445 -1720 17450 -1690
rect 17410 -1725 17450 -1720
rect 17670 -1690 17710 -1685
rect 17670 -1720 17675 -1690
rect 17705 -1720 17710 -1690
rect 17670 -1725 17710 -1720
rect 17780 -1690 17820 -1685
rect 17780 -1720 17785 -1690
rect 17815 -1720 17820 -1690
rect 17780 -1725 17820 -1720
rect 17890 -1690 17930 -1685
rect 17890 -1720 17895 -1690
rect 17925 -1720 17930 -1690
rect 17890 -1725 17930 -1720
rect 18205 -1690 18245 -1685
rect 18205 -1720 18210 -1690
rect 18240 -1720 18245 -1690
rect 18205 -1725 18245 -1720
rect 18315 -1695 18355 -1685
rect 18315 -1715 18325 -1695
rect 18345 -1715 18355 -1695
rect 18315 -1725 18355 -1715
rect 18425 -1690 18465 -1685
rect 18425 -1720 18430 -1690
rect 18460 -1720 18465 -1690
rect 18425 -1725 18465 -1720
rect 18535 -1695 18575 -1685
rect 18535 -1715 18545 -1695
rect 18565 -1715 18575 -1695
rect 18535 -1725 18575 -1715
rect 17310 -1740 17330 -1725
rect 17300 -1745 17340 -1740
rect 17300 -1775 17305 -1745
rect 17335 -1775 17340 -1745
rect 17300 -1780 17340 -1775
rect 17190 -1830 17195 -1800
rect 17225 -1830 17230 -1800
rect 17190 -1835 17230 -1830
rect 16765 -1855 16805 -1850
rect 16765 -1885 16770 -1855
rect 16800 -1885 16805 -1855
rect 17790 -1885 17810 -1725
rect 18325 -1740 18345 -1725
rect 18315 -1745 18355 -1740
rect 18315 -1775 18320 -1745
rect 18350 -1775 18355 -1745
rect 18315 -1780 18355 -1775
rect 18435 -1795 18455 -1725
rect 18545 -1740 18565 -1725
rect 18535 -1745 18575 -1740
rect 18535 -1775 18540 -1745
rect 18570 -1775 18575 -1745
rect 18535 -1780 18575 -1775
rect 18885 -1750 18925 -1745
rect 18885 -1780 18890 -1750
rect 18920 -1780 18925 -1750
rect 18425 -1800 18465 -1795
rect 18425 -1830 18430 -1800
rect 18460 -1830 18465 -1800
rect 18425 -1835 18465 -1830
rect 16765 -1890 16805 -1885
rect 17780 -1890 17820 -1885
rect 17780 -1920 17785 -1890
rect 17815 -1920 17820 -1890
rect 17780 -1925 17820 -1920
rect 16315 -2000 16355 -1995
rect 16315 -2030 16320 -2000
rect 16350 -2030 16355 -2000
rect 16315 -2035 16355 -2030
rect 17425 -2035 17430 -2000
rect 17465 -2035 17470 -2000
rect 18124 -2035 18129 -2000
rect 18164 -2035 18169 -2000
rect 18830 -2005 18870 -2000
rect 18830 -2035 18835 -2005
rect 18865 -2035 18870 -2005
rect 17425 -2060 17465 -2035
rect 17425 -2090 17430 -2060
rect 17460 -2090 17465 -2060
rect 17425 -2095 17465 -2090
rect 16260 -2100 16300 -2095
rect 16260 -2130 16265 -2100
rect 16295 -2130 16300 -2100
rect 16260 -2135 16300 -2130
rect 16480 -2100 16520 -2095
rect 16480 -2130 16485 -2100
rect 16515 -2130 16520 -2100
rect 16480 -2135 16520 -2130
rect 16730 -2100 16770 -2095
rect 16730 -2130 16735 -2100
rect 16765 -2130 16770 -2100
rect 16730 -2135 16770 -2130
rect 16490 -2895 16510 -2135
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 16160 -3025 16195 -3020
rect 16160 -3065 16195 -3060
rect 16740 -3100 16760 -2135
rect 16945 -2615 18655 -2265
rect 15820 -3115 15860 -3110
rect 15820 -3145 15825 -3115
rect 15855 -3145 15860 -3115
rect 15820 -4255 15860 -3145
rect 15950 -3116 15985 -3110
rect 16730 -3105 16770 -3100
rect 16730 -3135 16735 -3105
rect 16765 -3135 16770 -3105
rect 16730 -3140 16770 -3135
rect 15950 -3156 15985 -3151
rect 16945 -3625 17295 -2615
rect 17625 -3105 17975 -2945
rect 17625 -3135 17785 -3105
rect 17815 -3135 17975 -3105
rect 17625 -3295 17975 -3135
rect 18305 -3105 18655 -2615
rect 18305 -3135 18620 -3105
rect 18650 -3135 18655 -3105
rect 18305 -3625 18655 -3135
rect 18830 -3105 18870 -2035
rect 18830 -3135 18835 -3105
rect 18865 -3135 18870 -3105
rect 18830 -3140 18870 -3135
rect 15950 -3789 15985 -3784
rect 15950 -3829 15985 -3824
rect 15820 -4285 15825 -4255
rect 15855 -4285 15860 -4255
rect 15820 -4290 15860 -4285
rect 15645 -4375 15650 -4345
rect 15680 -4375 15690 -4345
rect 15720 -4375 15730 -4345
rect 15760 -4375 15765 -4345
rect 15645 -4385 15765 -4375
rect 15645 -4415 15650 -4385
rect 15680 -4415 15690 -4385
rect 15720 -4415 15730 -4385
rect 15760 -4415 15765 -4385
rect 15645 -4425 15765 -4415
rect 15645 -4455 15650 -4425
rect 15680 -4455 15690 -4425
rect 15720 -4455 15730 -4425
rect 15760 -4455 15765 -4425
rect 15645 -4460 15765 -4455
rect 15960 -4475 15980 -3829
rect 16280 -3894 16315 -3889
rect 16280 -3934 16315 -3929
rect 16290 -4105 16310 -3934
rect 16605 -3969 16640 -3964
rect 16945 -3975 18655 -3625
rect 16605 -4009 16640 -4004
rect 16615 -4105 16635 -4009
rect 16280 -4110 16320 -4105
rect 16280 -4140 16285 -4110
rect 16315 -4140 16320 -4110
rect 16280 -4150 16320 -4140
rect 16280 -4180 16285 -4150
rect 16315 -4180 16320 -4150
rect 16280 -4190 16320 -4180
rect 16280 -4220 16285 -4190
rect 16315 -4220 16320 -4190
rect 16280 -4225 16320 -4220
rect 16605 -4110 16645 -4105
rect 16605 -4140 16610 -4110
rect 16640 -4140 16645 -4110
rect 16605 -4150 16645 -4140
rect 16605 -4180 16610 -4150
rect 16640 -4180 16645 -4150
rect 16605 -4190 16645 -4180
rect 16605 -4220 16610 -4190
rect 16640 -4220 16645 -4190
rect 16605 -4225 16645 -4220
rect 17780 -4205 17820 -4200
rect 17780 -4235 17785 -4205
rect 17815 -4235 17820 -4205
rect 17780 -4245 17820 -4235
rect 17250 -4255 17300 -4245
rect 17250 -4285 17260 -4255
rect 17290 -4285 17300 -4255
rect 17250 -4295 17300 -4285
rect 17780 -4275 17785 -4245
rect 17815 -4275 17820 -4245
rect 17780 -4285 17820 -4275
rect 17780 -4315 17785 -4285
rect 17815 -4315 17820 -4285
rect 17780 -4320 17820 -4315
rect 16900 -4335 16950 -4325
rect 16900 -4365 16910 -4335
rect 16940 -4365 16950 -4335
rect 16900 -4385 16950 -4365
rect 16900 -4415 16910 -4385
rect 16940 -4415 16950 -4385
rect 16900 -4435 16950 -4415
rect 16900 -4465 16910 -4435
rect 16940 -4465 16950 -4435
rect 16900 -4475 16950 -4465
rect 18650 -4470 18700 -4460
rect 15950 -4480 15990 -4475
rect 15950 -4510 15955 -4480
rect 15985 -4510 15990 -4480
rect 15950 -4515 15990 -4510
rect 16205 -4480 16245 -4475
rect 16205 -4510 16210 -4480
rect 16240 -4510 16245 -4480
rect 18650 -4500 18660 -4470
rect 18690 -4500 18700 -4470
rect 18650 -4510 18700 -4500
rect 18885 -4470 18925 -1780
rect 19090 -1750 19130 -80
rect 19090 -1780 19095 -1750
rect 19125 -1780 19130 -1750
rect 19090 -1785 19130 -1780
rect 19325 -500 19365 1070
rect 19325 -530 19330 -500
rect 19360 -530 19365 -500
rect 19325 -1945 19365 -530
rect 19325 -1975 19330 -1945
rect 19360 -1975 19365 -1945
rect 19325 -1980 19365 -1975
rect 19405 375 19445 1640
rect 19405 345 19410 375
rect 19440 345 19445 375
rect 19405 -180 19445 345
rect 19405 -210 19410 -180
rect 19440 -210 19445 -180
rect 19080 -2060 19120 -2055
rect 19080 -2090 19085 -2060
rect 19115 -2090 19120 -2060
rect 19080 -2895 19120 -2090
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19405 -2995 19445 -210
rect 19545 -1885 19565 1640
rect 19610 1460 19650 1465
rect 19610 1430 19615 1460
rect 19645 1430 19650 1460
rect 19610 635 19650 1430
rect 19610 605 19615 635
rect 19645 605 19650 635
rect 19610 185 19650 605
rect 19610 155 19615 185
rect 19645 155 19650 185
rect 19535 -1890 19575 -1885
rect 19535 -1920 19540 -1890
rect 19570 -1920 19575 -1890
rect 19535 -1925 19575 -1920
rect 19405 -2997 19440 -2995
rect 19405 -3037 19440 -3032
rect 19610 -3115 19650 155
rect 19785 -1795 19805 1640
rect 19775 -1800 19815 -1795
rect 19775 -1830 19780 -1800
rect 19810 -1830 19815 -1800
rect 19775 -1835 19815 -1830
rect 19610 -3160 19645 -3150
rect 19610 -3789 19645 -3784
rect 19610 -3829 19645 -3824
rect 19285 -3894 19320 -3889
rect 19285 -3934 19320 -3929
rect 18960 -3969 18995 -3964
rect 18960 -4009 18995 -4004
rect 18965 -4200 18985 -4009
rect 19290 -4200 19310 -3934
rect 18955 -4205 18995 -4200
rect 18955 -4235 18960 -4205
rect 18990 -4235 18995 -4205
rect 18955 -4245 18995 -4235
rect 18955 -4275 18960 -4245
rect 18990 -4275 18995 -4245
rect 18955 -4285 18995 -4275
rect 18955 -4315 18960 -4285
rect 18990 -4315 18995 -4285
rect 18955 -4320 18995 -4315
rect 19280 -4205 19320 -4200
rect 19280 -4235 19285 -4205
rect 19315 -4235 19320 -4205
rect 19280 -4245 19320 -4235
rect 19280 -4275 19285 -4245
rect 19315 -4275 19320 -4245
rect 19280 -4285 19320 -4275
rect 19280 -4315 19285 -4285
rect 19315 -4315 19320 -4285
rect 19280 -4320 19320 -4315
rect 19620 -4465 19640 -3829
rect 18885 -4500 18890 -4470
rect 18920 -4500 18925 -4470
rect 18885 -4505 18925 -4500
rect 19355 -4470 19395 -4465
rect 19355 -4500 19360 -4470
rect 19390 -4500 19395 -4470
rect 19355 -4505 19395 -4500
rect 19610 -4470 19650 -4465
rect 19610 -4500 19615 -4470
rect 19645 -4500 19650 -4470
rect 19610 -4505 19650 -4500
rect 16205 -4515 16245 -4510
rect 17955 -4520 17995 -4515
rect 17955 -4550 17960 -4520
rect 17990 -4550 17995 -4520
rect 17955 -4555 17995 -4550
<< via1 >>
rect 15650 -75 15680 -45
rect 15690 -75 15720 -45
rect 15730 -75 15760 -45
rect 15650 -115 15680 -85
rect 15690 -115 15720 -85
rect 15730 -115 15760 -85
rect 15650 -155 15680 -125
rect 15690 -155 15720 -125
rect 15730 -155 15760 -125
rect 15895 1125 15925 1155
rect 15895 -1415 15925 -1385
rect 15950 155 15980 185
rect 15790 -1830 15820 -1800
rect 16035 -1775 16065 -1745
rect 16490 1455 16520 1460
rect 16490 1435 16495 1455
rect 16495 1435 16515 1455
rect 16515 1435 16520 1455
rect 16490 1430 16520 1435
rect 16370 1375 16400 1405
rect 16370 1335 16400 1365
rect 16370 1320 16400 1325
rect 16370 1300 16375 1320
rect 16375 1300 16395 1320
rect 16395 1300 16400 1320
rect 16370 1295 16400 1300
rect 16490 1375 16520 1405
rect 16490 1335 16520 1365
rect 16490 1320 16520 1325
rect 16490 1300 16495 1320
rect 16495 1300 16515 1320
rect 16515 1300 16520 1320
rect 16490 1295 16520 1300
rect 16610 1375 16640 1405
rect 16610 1335 16640 1365
rect 16610 1320 16640 1325
rect 16610 1300 16615 1320
rect 16615 1300 16635 1320
rect 16635 1300 16640 1320
rect 16610 1295 16640 1300
rect 16890 1375 16920 1405
rect 16890 1335 16920 1365
rect 17055 1430 17085 1460
rect 17000 1375 17030 1405
rect 17000 1335 17030 1365
rect 16890 1320 16920 1325
rect 16890 1300 16895 1320
rect 16895 1300 16915 1320
rect 16915 1300 16920 1320
rect 16890 1295 16920 1300
rect 17000 1320 17030 1325
rect 17000 1300 17005 1320
rect 17005 1300 17025 1320
rect 17025 1300 17030 1320
rect 17000 1295 17030 1300
rect 17110 1375 17140 1405
rect 17110 1335 17140 1365
rect 17110 1320 17140 1325
rect 17110 1300 17115 1320
rect 17115 1300 17135 1320
rect 17135 1300 17140 1320
rect 17110 1295 17140 1300
rect 17220 1375 17250 1405
rect 17220 1335 17250 1365
rect 17220 1320 17250 1325
rect 17220 1300 17225 1320
rect 17225 1300 17245 1320
rect 17245 1300 17250 1320
rect 17220 1295 17250 1300
rect 17500 1375 17530 1405
rect 17500 1335 17530 1365
rect 17500 1320 17530 1325
rect 17500 1300 17505 1320
rect 17505 1300 17525 1320
rect 17525 1300 17530 1320
rect 17500 1295 17530 1300
rect 17565 1375 17595 1405
rect 17565 1335 17595 1365
rect 17565 1320 17595 1325
rect 17565 1300 17570 1320
rect 17570 1300 17590 1320
rect 17590 1300 17595 1320
rect 17565 1295 17595 1300
rect 17675 1375 17705 1405
rect 17675 1335 17705 1365
rect 17675 1320 17705 1325
rect 17675 1300 17680 1320
rect 17680 1300 17700 1320
rect 17700 1300 17705 1320
rect 17675 1295 17705 1300
rect 17785 1455 17815 1460
rect 17785 1435 17790 1455
rect 17790 1435 17810 1455
rect 17810 1435 17815 1455
rect 17785 1430 17815 1435
rect 17785 1375 17815 1405
rect 17785 1335 17815 1365
rect 17785 1320 17815 1325
rect 17785 1300 17790 1320
rect 17790 1300 17810 1320
rect 17810 1300 17815 1320
rect 17785 1295 17815 1300
rect 17895 1375 17925 1405
rect 17895 1335 17925 1365
rect 17895 1320 17925 1325
rect 17895 1300 17900 1320
rect 17900 1300 17920 1320
rect 17920 1300 17925 1320
rect 17895 1295 17925 1300
rect 18515 1430 18545 1460
rect 18005 1375 18035 1405
rect 18005 1335 18035 1365
rect 18005 1320 18035 1325
rect 18005 1300 18010 1320
rect 18010 1300 18030 1320
rect 18030 1300 18035 1320
rect 18005 1295 18035 1300
rect 18070 1375 18100 1405
rect 18070 1335 18100 1365
rect 18070 1320 18100 1325
rect 18070 1300 18075 1320
rect 18075 1300 18095 1320
rect 18095 1300 18100 1320
rect 18070 1295 18100 1300
rect 18350 1375 18380 1405
rect 18350 1335 18380 1365
rect 18350 1320 18380 1325
rect 18350 1300 18355 1320
rect 18355 1300 18375 1320
rect 18375 1300 18380 1320
rect 18350 1295 18380 1300
rect 18460 1375 18490 1405
rect 18460 1335 18490 1365
rect 18570 1375 18600 1405
rect 18570 1335 18600 1365
rect 18460 1320 18490 1325
rect 18460 1300 18465 1320
rect 18465 1300 18485 1320
rect 18485 1300 18490 1320
rect 18460 1295 18490 1300
rect 18680 1375 18710 1405
rect 18680 1335 18710 1365
rect 18570 1320 18600 1325
rect 18570 1300 18575 1320
rect 18575 1300 18595 1320
rect 18595 1300 18600 1320
rect 18570 1295 18600 1300
rect 18680 1320 18710 1325
rect 18680 1300 18685 1320
rect 18685 1300 18705 1320
rect 18705 1300 18710 1320
rect 18680 1295 18710 1300
rect 16435 1150 16465 1155
rect 16435 1130 16440 1150
rect 16440 1130 16460 1150
rect 16460 1130 16465 1150
rect 16435 1125 16465 1130
rect 16545 1150 16575 1155
rect 16545 1130 16550 1150
rect 16550 1130 16570 1150
rect 16570 1130 16575 1150
rect 16545 1125 16575 1130
rect 16945 1150 16975 1155
rect 16945 1130 16950 1150
rect 16950 1130 16970 1150
rect 16970 1130 16975 1150
rect 16945 1125 16975 1130
rect 17055 1150 17085 1155
rect 17055 1130 17060 1150
rect 17060 1130 17080 1150
rect 17080 1130 17085 1150
rect 17055 1125 17085 1130
rect 17165 1150 17195 1155
rect 17165 1130 17170 1150
rect 17170 1130 17190 1150
rect 17190 1130 17195 1150
rect 17165 1125 17195 1130
rect 17620 1150 17650 1155
rect 17620 1130 17625 1150
rect 17625 1130 17645 1150
rect 17645 1130 17650 1150
rect 17620 1125 17650 1130
rect 17730 1150 17760 1155
rect 17730 1130 17735 1150
rect 17735 1130 17755 1150
rect 17755 1130 17760 1150
rect 17730 1125 17760 1130
rect 17840 1150 17870 1155
rect 17840 1130 17845 1150
rect 17845 1130 17865 1150
rect 17865 1130 17870 1150
rect 17840 1125 17870 1130
rect 17950 1150 17980 1155
rect 17950 1130 17955 1150
rect 17955 1130 17975 1150
rect 17975 1130 17980 1150
rect 17950 1125 17980 1130
rect 18405 1150 18435 1155
rect 18405 1130 18410 1150
rect 18410 1130 18430 1150
rect 18430 1130 18435 1150
rect 18405 1125 18435 1130
rect 18515 1150 18545 1155
rect 18515 1130 18520 1150
rect 18520 1130 18540 1150
rect 18540 1130 18545 1150
rect 18515 1125 18545 1130
rect 18625 1150 18655 1155
rect 18625 1130 18630 1150
rect 18630 1130 18650 1150
rect 18650 1130 18655 1150
rect 18625 1125 18655 1130
rect 16545 1070 16575 1100
rect 16440 1015 16470 1045
rect 16440 975 16470 1005
rect 16440 935 16470 965
rect 16660 1015 16690 1045
rect 16660 975 16690 1005
rect 16660 935 16690 965
rect 16975 1015 17005 1045
rect 16975 975 17005 1005
rect 16975 960 17005 965
rect 16975 940 16980 960
rect 16980 940 17000 960
rect 17000 940 17005 960
rect 16975 935 17005 940
rect 17155 1015 17185 1045
rect 17155 975 17185 1005
rect 17155 960 17185 965
rect 17155 940 17160 960
rect 17160 940 17180 960
rect 17180 940 17185 960
rect 17155 935 17185 940
rect 17335 1015 17365 1045
rect 17335 975 17365 1005
rect 17335 960 17365 965
rect 17335 940 17340 960
rect 17340 940 17360 960
rect 17360 940 17365 960
rect 17335 935 17365 940
rect 17515 1015 17545 1045
rect 17515 975 17545 1005
rect 17515 960 17545 965
rect 17515 940 17520 960
rect 17520 940 17540 960
rect 17540 940 17545 960
rect 17515 935 17545 940
rect 17695 1015 17725 1045
rect 17695 975 17725 1005
rect 17695 960 17725 965
rect 17695 940 17700 960
rect 17700 940 17720 960
rect 17720 940 17725 960
rect 17695 935 17725 940
rect 17875 1015 17905 1045
rect 17875 975 17905 1005
rect 17875 960 17905 965
rect 17875 940 17880 960
rect 17880 940 17900 960
rect 17900 940 17905 960
rect 17875 935 17905 940
rect 18055 1015 18085 1045
rect 18055 975 18085 1005
rect 18055 960 18085 965
rect 18055 940 18060 960
rect 18060 940 18080 960
rect 18080 940 18085 960
rect 18055 935 18085 940
rect 18235 1015 18265 1045
rect 18235 975 18265 1005
rect 18235 960 18265 965
rect 18235 940 18240 960
rect 18240 940 18260 960
rect 18260 940 18265 960
rect 18235 935 18265 940
rect 18415 1015 18445 1045
rect 18415 975 18445 1005
rect 18415 960 18445 965
rect 18415 940 18420 960
rect 18420 940 18440 960
rect 18440 940 18445 960
rect 18415 935 18445 940
rect 18595 1015 18625 1045
rect 18595 975 18625 1005
rect 18595 960 18625 965
rect 18595 940 18600 960
rect 18600 940 18620 960
rect 18620 940 18625 960
rect 18595 935 18625 940
rect 18910 1015 18940 1045
rect 18910 975 18940 1005
rect 18910 960 18940 965
rect 18910 940 18915 960
rect 18915 940 18935 960
rect 18935 940 18940 960
rect 18910 935 18940 940
rect 16550 860 16580 865
rect 16550 840 16555 860
rect 16555 840 16575 860
rect 16575 840 16580 860
rect 16550 835 16580 840
rect 16785 835 16815 865
rect 16485 690 16515 695
rect 16485 670 16490 690
rect 16490 670 16510 690
rect 16510 670 16515 690
rect 16485 665 16515 670
rect 16320 510 16350 540
rect 16265 455 16295 485
rect 16210 400 16240 430
rect 16265 -210 16295 -180
rect 16210 -1315 16240 -1285
rect 16110 -1885 16140 -1855
rect 16160 -1975 16190 -1945
rect 16425 290 16455 320
rect 16425 250 16455 280
rect 16425 210 16455 240
rect 16615 690 16645 695
rect 16615 670 16620 690
rect 16620 670 16640 690
rect 16640 670 16645 690
rect 16615 665 16645 670
rect 16785 455 16815 485
rect 16550 400 16580 430
rect 17110 590 17140 595
rect 17110 570 17115 590
rect 17115 570 17135 590
rect 17135 570 17140 590
rect 17110 565 17140 570
rect 17200 590 17230 595
rect 17200 570 17205 590
rect 17205 570 17225 590
rect 17225 570 17230 590
rect 17200 565 17230 570
rect 17290 590 17320 595
rect 17290 570 17295 590
rect 17295 570 17315 590
rect 17315 570 17320 590
rect 17290 565 17320 570
rect 17380 590 17410 595
rect 17380 570 17385 590
rect 17385 570 17405 590
rect 17405 570 17410 590
rect 17380 565 17410 570
rect 17470 590 17500 595
rect 17470 570 17475 590
rect 17475 570 17495 590
rect 17495 570 17500 590
rect 17470 565 17500 570
rect 17560 590 17590 595
rect 17560 570 17565 590
rect 17565 570 17585 590
rect 17585 570 17590 590
rect 17560 565 17590 570
rect 17650 590 17680 595
rect 17650 570 17655 590
rect 17655 570 17675 590
rect 17675 570 17680 590
rect 17650 565 17680 570
rect 17695 565 17725 595
rect 17740 590 17770 595
rect 17740 570 17745 590
rect 17745 570 17765 590
rect 17765 570 17770 590
rect 17740 565 17770 570
rect 17605 510 17635 540
rect 17425 455 17455 485
rect 17245 400 17275 430
rect 17065 345 17095 375
rect 16545 290 16575 320
rect 16545 250 16575 280
rect 16545 210 16575 240
rect 16665 290 16695 320
rect 16665 250 16695 280
rect 16665 210 16695 240
rect 16785 290 16815 320
rect 16785 250 16815 280
rect 16785 210 16815 240
rect 16905 290 16935 320
rect 16905 250 16935 280
rect 16905 210 16935 240
rect 17025 290 17055 320
rect 17025 250 17055 280
rect 17025 210 17055 240
rect 17145 290 17175 320
rect 17145 250 17175 280
rect 17145 210 17175 240
rect 17265 290 17295 320
rect 17265 250 17295 280
rect 17265 210 17295 240
rect 17385 290 17415 320
rect 17385 250 17415 280
rect 17385 210 17415 240
rect 17505 290 17535 320
rect 17505 250 17535 280
rect 17505 210 17535 240
rect 17625 290 17655 320
rect 17625 250 17655 280
rect 17625 210 17655 240
rect 16485 155 16515 185
rect 16605 10 16635 15
rect 16605 -10 16610 10
rect 16610 -10 16630 10
rect 16630 -10 16635 10
rect 16605 -15 16635 -10
rect 16845 155 16875 185
rect 16965 10 16995 15
rect 16965 -10 16970 10
rect 16970 -10 16990 10
rect 16990 -10 16995 10
rect 16965 -15 16995 -10
rect 16515 -75 16545 -45
rect 16515 -115 16545 -85
rect 16515 -155 16545 -125
rect 16725 -75 16755 -45
rect 16725 -115 16755 -85
rect 16725 -155 16755 -125
rect 16845 -75 16875 -45
rect 16845 -115 16875 -85
rect 16845 -155 16875 -125
rect 17205 155 17235 185
rect 17325 10 17355 15
rect 17325 -10 17330 10
rect 17330 -10 17350 10
rect 17350 -10 17355 10
rect 17325 -15 17355 -10
rect 17565 155 17595 185
rect 17830 590 17860 595
rect 17830 570 17835 590
rect 17835 570 17855 590
rect 17855 570 17860 590
rect 17830 565 17860 570
rect 17920 590 17950 595
rect 17920 570 17925 590
rect 17925 570 17945 590
rect 17945 570 17950 590
rect 17920 565 17950 570
rect 18010 590 18040 595
rect 18010 570 18015 590
rect 18015 570 18035 590
rect 18035 570 18040 590
rect 18010 565 18040 570
rect 18100 590 18130 595
rect 18100 570 18105 590
rect 18105 570 18125 590
rect 18125 570 18130 590
rect 18100 565 18130 570
rect 17965 510 17995 540
rect 18190 590 18220 595
rect 18190 570 18195 590
rect 18195 570 18215 590
rect 18215 570 18220 590
rect 18190 565 18220 570
rect 18280 590 18310 595
rect 18280 570 18285 590
rect 18285 570 18305 590
rect 18305 570 18310 590
rect 18280 565 18310 570
rect 18145 455 18175 485
rect 18370 590 18400 595
rect 18370 570 18375 590
rect 18375 570 18395 590
rect 18395 570 18400 590
rect 18370 565 18400 570
rect 18460 590 18490 595
rect 18460 570 18465 590
rect 18465 570 18485 590
rect 18485 570 18490 590
rect 18460 565 18490 570
rect 18325 400 18355 430
rect 19330 1070 19360 1100
rect 19020 1015 19050 1045
rect 19020 975 19050 1005
rect 19020 960 19050 965
rect 19020 940 19025 960
rect 19025 940 19045 960
rect 19045 940 19050 960
rect 19020 935 19050 940
rect 19080 1015 19110 1045
rect 19080 975 19110 1005
rect 19080 960 19110 965
rect 19080 940 19085 960
rect 19085 940 19105 960
rect 19105 940 19110 960
rect 19080 935 19110 940
rect 19005 630 19035 635
rect 19005 610 19010 630
rect 19010 610 19030 630
rect 19030 610 19035 630
rect 19005 605 19035 610
rect 17785 345 17815 375
rect 18505 345 18535 375
rect 17945 290 17975 320
rect 17945 250 17975 280
rect 17945 210 17975 240
rect 18065 290 18095 320
rect 18065 250 18095 280
rect 18065 210 18095 240
rect 18185 290 18215 320
rect 18185 250 18215 280
rect 18185 210 18215 240
rect 18305 290 18335 320
rect 18305 250 18335 280
rect 18305 210 18335 240
rect 18425 290 18455 320
rect 18425 250 18455 280
rect 18425 210 18455 240
rect 18545 290 18575 320
rect 18545 250 18575 280
rect 18545 210 18575 240
rect 18665 290 18695 320
rect 18665 250 18695 280
rect 18665 210 18695 240
rect 18785 290 18815 320
rect 18785 250 18815 280
rect 18785 210 18815 240
rect 18905 290 18935 320
rect 18905 250 18935 280
rect 18905 210 18935 240
rect 19025 290 19055 320
rect 19025 250 19055 280
rect 19025 210 19055 240
rect 19145 290 19175 320
rect 19145 250 19175 280
rect 19145 210 19175 240
rect 17695 155 17725 185
rect 17875 155 17905 185
rect 17085 -75 17115 -45
rect 17085 -115 17115 -85
rect 17085 -155 17115 -125
rect 17205 -75 17235 -45
rect 17205 -115 17235 -85
rect 17205 -155 17235 -125
rect 17445 -75 17475 -45
rect 17445 -115 17475 -85
rect 17445 -155 17475 -125
rect 17535 -75 17565 -45
rect 17535 -115 17565 -85
rect 17535 -155 17565 -125
rect 17007 -185 17037 -180
rect 17007 -205 17012 -185
rect 17012 -205 17032 -185
rect 17032 -205 17037 -185
rect 17007 -210 17037 -205
rect 16320 -530 16350 -500
rect 17565 -245 17595 -240
rect 17565 -265 17570 -245
rect 17570 -265 17590 -245
rect 17590 -265 17595 -245
rect 17565 -270 17595 -265
rect 17565 -285 17595 -280
rect 17565 -305 17570 -285
rect 17570 -305 17590 -285
rect 17590 -305 17595 -285
rect 17565 -310 17595 -305
rect 17565 -325 17595 -320
rect 17565 -345 17570 -325
rect 17570 -345 17590 -325
rect 17590 -345 17595 -325
rect 17565 -350 17595 -345
rect 17075 -505 17105 -500
rect 17075 -525 17080 -505
rect 17080 -525 17100 -505
rect 17100 -525 17105 -505
rect 17075 -530 17105 -525
rect 16535 -640 16565 -610
rect 17025 -640 17055 -610
rect 16625 -695 16655 -665
rect 16625 -735 16655 -705
rect 16625 -750 16655 -745
rect 16625 -770 16630 -750
rect 16630 -770 16650 -750
rect 16650 -770 16655 -750
rect 16625 -775 16655 -770
rect 16745 -695 16775 -665
rect 16745 -735 16775 -705
rect 16745 -750 16775 -745
rect 16745 -770 16750 -750
rect 16750 -770 16770 -750
rect 16770 -770 16775 -750
rect 16745 -775 16775 -770
rect 16865 -695 16895 -665
rect 16865 -735 16895 -705
rect 16865 -750 16895 -745
rect 16865 -770 16870 -750
rect 16870 -770 16890 -750
rect 16890 -770 16895 -750
rect 16865 -775 16895 -770
rect 16985 -695 17015 -665
rect 16985 -735 17015 -705
rect 16985 -750 17015 -745
rect 16985 -770 16990 -750
rect 16990 -770 17010 -750
rect 17010 -770 17015 -750
rect 16985 -775 17015 -770
rect 17305 -695 17335 -665
rect 17305 -735 17335 -705
rect 17305 -750 17335 -745
rect 17305 -770 17310 -750
rect 17310 -770 17330 -750
rect 17330 -770 17335 -750
rect 17305 -775 17335 -770
rect 17425 -695 17455 -665
rect 17425 -735 17455 -705
rect 17425 -750 17455 -745
rect 17425 -770 17430 -750
rect 17430 -770 17450 -750
rect 17450 -770 17455 -750
rect 17425 -775 17455 -770
rect 17545 -695 17575 -665
rect 17545 -735 17575 -705
rect 17545 -750 17575 -745
rect 17545 -770 17550 -750
rect 17550 -770 17570 -750
rect 17570 -770 17575 -750
rect 17545 -775 17575 -770
rect 17745 -270 17775 -240
rect 17785 -270 17815 -240
rect 17825 -270 17855 -240
rect 17745 -310 17775 -280
rect 17785 -310 17815 -280
rect 17825 -310 17855 -280
rect 17745 -350 17775 -320
rect 17785 -350 17815 -320
rect 17825 -350 17855 -320
rect 17115 -1070 17145 -1065
rect 17115 -1090 17120 -1070
rect 17120 -1090 17140 -1070
rect 17140 -1090 17145 -1070
rect 17115 -1095 17145 -1090
rect 17115 -1135 17145 -1105
rect 17115 -1175 17145 -1145
rect 18005 155 18035 185
rect 18365 155 18395 185
rect 18245 10 18275 15
rect 18245 -10 18250 10
rect 18250 -10 18270 10
rect 18270 -10 18275 10
rect 18245 -15 18275 -10
rect 18725 155 18755 185
rect 18605 10 18635 15
rect 18605 -10 18610 10
rect 18610 -10 18630 10
rect 18630 -10 18635 10
rect 18605 -15 18635 -10
rect 18035 -75 18065 -45
rect 18125 -75 18155 -45
rect 18365 -75 18395 -45
rect 18485 -75 18515 -45
rect 18005 -245 18035 -240
rect 18005 -265 18010 -245
rect 18010 -265 18030 -245
rect 18030 -265 18035 -245
rect 18005 -270 18035 -265
rect 18005 -285 18035 -280
rect 18005 -305 18010 -285
rect 18010 -305 18030 -285
rect 18030 -305 18035 -285
rect 18005 -310 18035 -305
rect 18005 -325 18035 -320
rect 18005 -345 18010 -325
rect 18010 -345 18030 -325
rect 18030 -345 18035 -325
rect 18005 -350 18035 -345
rect 18563 -185 18593 -180
rect 18563 -205 18568 -185
rect 18568 -205 18588 -185
rect 18588 -205 18593 -185
rect 18563 -210 18593 -205
rect 19085 155 19115 185
rect 18965 10 18995 15
rect 18965 -10 18970 10
rect 18970 -10 18990 10
rect 18990 -10 18995 10
rect 18965 -15 18995 -10
rect 18725 -75 18755 -45
rect 18845 -75 18875 -45
rect 19055 -75 19085 -45
rect 19095 -75 19125 -45
rect 18440 -505 18470 -500
rect 18440 -525 18445 -505
rect 18445 -525 18465 -505
rect 18465 -525 18470 -505
rect 18440 -530 18470 -525
rect 18545 -640 18575 -610
rect 19035 -640 19065 -610
rect 18025 -695 18055 -665
rect 18025 -735 18055 -705
rect 18025 -750 18055 -745
rect 18025 -770 18030 -750
rect 18030 -770 18050 -750
rect 18050 -770 18055 -750
rect 18025 -775 18055 -770
rect 18145 -695 18175 -665
rect 18145 -735 18175 -705
rect 18145 -750 18175 -745
rect 18145 -770 18150 -750
rect 18150 -770 18170 -750
rect 18170 -770 18175 -750
rect 18145 -775 18175 -770
rect 18265 -695 18295 -665
rect 18265 -735 18295 -705
rect 18265 -750 18295 -745
rect 18265 -770 18270 -750
rect 18270 -770 18290 -750
rect 18290 -770 18295 -750
rect 18265 -775 18295 -770
rect 18585 -695 18615 -665
rect 18585 -735 18615 -705
rect 18585 -750 18615 -745
rect 18585 -770 18590 -750
rect 18590 -770 18610 -750
rect 18610 -770 18615 -750
rect 18585 -775 18615 -770
rect 18705 -695 18735 -665
rect 18705 -735 18735 -705
rect 18705 -750 18735 -745
rect 18705 -770 18710 -750
rect 18710 -770 18730 -750
rect 18730 -770 18735 -750
rect 18705 -775 18735 -770
rect 18825 -695 18855 -665
rect 18825 -735 18855 -705
rect 18825 -750 18855 -745
rect 18825 -770 18830 -750
rect 18830 -770 18850 -750
rect 18850 -770 18855 -750
rect 18825 -775 18855 -770
rect 18945 -695 18975 -665
rect 18945 -735 18975 -705
rect 18945 -750 18975 -745
rect 18945 -770 18950 -750
rect 18950 -770 18970 -750
rect 18970 -770 18975 -750
rect 18945 -775 18975 -770
rect 17745 -1095 17775 -1065
rect 17785 -1095 17815 -1065
rect 17825 -1095 17855 -1065
rect 17745 -1135 17775 -1105
rect 17785 -1135 17815 -1105
rect 17825 -1135 17855 -1105
rect 17745 -1175 17775 -1145
rect 17785 -1175 17815 -1145
rect 17825 -1175 17855 -1145
rect 18455 -1070 18485 -1065
rect 18455 -1090 18460 -1070
rect 18460 -1090 18480 -1070
rect 18480 -1090 18485 -1070
rect 18455 -1095 18485 -1090
rect 18455 -1135 18485 -1105
rect 18455 -1175 18485 -1145
rect 16745 -1205 16775 -1200
rect 16745 -1225 16750 -1205
rect 16750 -1225 16770 -1205
rect 16770 -1225 16775 -1205
rect 16745 -1230 16775 -1225
rect 16825 -1205 16855 -1200
rect 16825 -1225 16830 -1205
rect 16830 -1225 16850 -1205
rect 16850 -1225 16855 -1205
rect 16825 -1230 16855 -1225
rect 16905 -1205 16935 -1200
rect 16905 -1225 16910 -1205
rect 16910 -1225 16930 -1205
rect 16930 -1225 16935 -1205
rect 16905 -1230 16935 -1225
rect 16985 -1205 17015 -1200
rect 16985 -1225 16990 -1205
rect 16990 -1225 17010 -1205
rect 17010 -1225 17015 -1205
rect 16985 -1230 17015 -1225
rect 17065 -1205 17095 -1200
rect 17065 -1225 17070 -1205
rect 17070 -1225 17090 -1205
rect 17090 -1225 17095 -1205
rect 17065 -1230 17095 -1225
rect 17145 -1205 17175 -1200
rect 17145 -1225 17150 -1205
rect 17150 -1225 17170 -1205
rect 17170 -1225 17175 -1205
rect 17145 -1230 17175 -1225
rect 17225 -1205 17255 -1200
rect 17225 -1225 17230 -1205
rect 17230 -1225 17250 -1205
rect 17250 -1225 17255 -1205
rect 17225 -1230 17255 -1225
rect 17305 -1205 17335 -1200
rect 17305 -1225 17310 -1205
rect 17310 -1225 17330 -1205
rect 17330 -1225 17335 -1205
rect 17305 -1230 17335 -1225
rect 17385 -1205 17415 -1200
rect 17385 -1225 17390 -1205
rect 17390 -1225 17410 -1205
rect 17410 -1225 17415 -1205
rect 17385 -1230 17415 -1225
rect 17465 -1205 17495 -1200
rect 17465 -1225 17470 -1205
rect 17470 -1225 17490 -1205
rect 17490 -1225 17495 -1205
rect 17465 -1230 17495 -1225
rect 17545 -1205 17575 -1200
rect 17545 -1225 17550 -1205
rect 17550 -1225 17570 -1205
rect 17570 -1225 17575 -1205
rect 17545 -1230 17575 -1225
rect 17625 -1205 17655 -1200
rect 17625 -1225 17630 -1205
rect 17630 -1225 17650 -1205
rect 17650 -1225 17655 -1205
rect 17625 -1230 17655 -1225
rect 17705 -1205 17735 -1200
rect 17705 -1225 17710 -1205
rect 17710 -1225 17730 -1205
rect 17730 -1225 17735 -1205
rect 17705 -1230 17735 -1225
rect 17785 -1205 17815 -1200
rect 17785 -1225 17790 -1205
rect 17790 -1225 17810 -1205
rect 17810 -1225 17815 -1205
rect 17785 -1230 17815 -1225
rect 17865 -1205 17895 -1200
rect 17865 -1225 17870 -1205
rect 17870 -1225 17890 -1205
rect 17890 -1225 17895 -1205
rect 17865 -1230 17895 -1225
rect 17945 -1205 17975 -1200
rect 17945 -1225 17950 -1205
rect 17950 -1225 17970 -1205
rect 17970 -1225 17975 -1205
rect 17945 -1230 17975 -1225
rect 18025 -1205 18055 -1200
rect 18025 -1225 18030 -1205
rect 18030 -1225 18050 -1205
rect 18050 -1225 18055 -1205
rect 18025 -1230 18055 -1225
rect 18105 -1205 18135 -1200
rect 18105 -1225 18110 -1205
rect 18110 -1225 18130 -1205
rect 18130 -1225 18135 -1205
rect 18105 -1230 18135 -1225
rect 18185 -1205 18215 -1200
rect 18185 -1225 18190 -1205
rect 18190 -1225 18210 -1205
rect 18210 -1225 18215 -1205
rect 18185 -1230 18215 -1225
rect 18265 -1205 18295 -1200
rect 18265 -1225 18270 -1205
rect 18270 -1225 18290 -1205
rect 18290 -1225 18295 -1205
rect 18265 -1230 18295 -1225
rect 18345 -1205 18375 -1200
rect 18345 -1225 18350 -1205
rect 18350 -1225 18370 -1205
rect 18370 -1225 18375 -1205
rect 18345 -1230 18375 -1225
rect 18425 -1205 18455 -1200
rect 18425 -1225 18430 -1205
rect 18430 -1225 18450 -1205
rect 18450 -1225 18455 -1205
rect 18425 -1230 18455 -1225
rect 18505 -1205 18535 -1200
rect 18505 -1225 18510 -1205
rect 18510 -1225 18530 -1205
rect 18530 -1225 18535 -1205
rect 18505 -1230 18535 -1225
rect 18585 -1205 18615 -1200
rect 18585 -1225 18590 -1205
rect 18590 -1225 18610 -1205
rect 18610 -1225 18615 -1205
rect 18585 -1230 18615 -1225
rect 18665 -1205 18695 -1200
rect 18665 -1225 18670 -1205
rect 18670 -1225 18690 -1205
rect 18690 -1225 18695 -1205
rect 18665 -1230 18695 -1225
rect 18745 -1205 18775 -1200
rect 18745 -1225 18750 -1205
rect 18750 -1225 18770 -1205
rect 18770 -1225 18775 -1205
rect 18745 -1230 18775 -1225
rect 16705 -1290 16735 -1285
rect 16705 -1310 16710 -1290
rect 16710 -1310 16730 -1290
rect 16730 -1310 16735 -1290
rect 16705 -1315 16735 -1310
rect 18900 -1270 18930 -1265
rect 18900 -1290 18905 -1270
rect 18905 -1290 18925 -1270
rect 18925 -1290 18930 -1270
rect 18900 -1295 18930 -1290
rect 18900 -1310 18930 -1305
rect 18900 -1330 18905 -1310
rect 18905 -1330 18925 -1310
rect 18925 -1330 18930 -1310
rect 18900 -1335 18930 -1330
rect 16660 -1415 16690 -1385
rect 16770 -1415 16800 -1385
rect 17305 -1415 17335 -1385
rect 17785 -1415 17815 -1385
rect 18320 -1415 18350 -1385
rect 16605 -1470 16635 -1440
rect 16605 -1510 16635 -1480
rect 16605 -1525 16635 -1520
rect 16605 -1545 16610 -1525
rect 16610 -1545 16630 -1525
rect 16630 -1545 16635 -1525
rect 16605 -1550 16635 -1545
rect 16715 -1470 16745 -1440
rect 16715 -1510 16745 -1480
rect 16715 -1525 16745 -1520
rect 16715 -1545 16720 -1525
rect 16720 -1545 16740 -1525
rect 16740 -1545 16745 -1525
rect 16715 -1550 16745 -1545
rect 16825 -1470 16855 -1440
rect 16825 -1510 16855 -1480
rect 16825 -1525 16855 -1520
rect 16825 -1545 16830 -1525
rect 16830 -1545 16850 -1525
rect 16850 -1545 16855 -1525
rect 16825 -1550 16855 -1545
rect 16885 -1470 16915 -1440
rect 16885 -1510 16915 -1480
rect 16885 -1525 16915 -1520
rect 16885 -1545 16890 -1525
rect 16890 -1545 16910 -1525
rect 16910 -1545 16915 -1525
rect 16885 -1550 16915 -1545
rect 17030 -1470 17060 -1440
rect 17030 -1510 17060 -1480
rect 17030 -1525 17060 -1520
rect 17030 -1545 17035 -1525
rect 17035 -1545 17055 -1525
rect 17055 -1545 17060 -1525
rect 17030 -1550 17060 -1545
rect 17140 -1470 17170 -1440
rect 17140 -1510 17170 -1480
rect 17140 -1525 17170 -1520
rect 17140 -1545 17145 -1525
rect 17145 -1545 17165 -1525
rect 17165 -1545 17170 -1525
rect 17140 -1550 17170 -1545
rect 17250 -1470 17280 -1440
rect 17250 -1510 17280 -1480
rect 17250 -1525 17280 -1520
rect 17250 -1545 17255 -1525
rect 17255 -1545 17275 -1525
rect 17275 -1545 17280 -1525
rect 17250 -1550 17280 -1545
rect 17360 -1470 17390 -1440
rect 17360 -1510 17390 -1480
rect 17360 -1525 17390 -1520
rect 17360 -1545 17365 -1525
rect 17365 -1545 17385 -1525
rect 17385 -1545 17390 -1525
rect 17360 -1550 17390 -1545
rect 17470 -1470 17500 -1440
rect 17470 -1510 17500 -1480
rect 17470 -1525 17500 -1520
rect 17470 -1545 17475 -1525
rect 17475 -1545 17495 -1525
rect 17495 -1545 17500 -1525
rect 17470 -1550 17500 -1545
rect 17620 -1470 17650 -1440
rect 17620 -1510 17650 -1480
rect 17620 -1525 17650 -1520
rect 17620 -1545 17625 -1525
rect 17625 -1545 17645 -1525
rect 17645 -1545 17650 -1525
rect 17620 -1550 17650 -1545
rect 17730 -1470 17760 -1440
rect 17730 -1510 17760 -1480
rect 17730 -1525 17760 -1520
rect 17730 -1545 17735 -1525
rect 17735 -1545 17755 -1525
rect 17755 -1545 17760 -1525
rect 17730 -1550 17760 -1545
rect 17840 -1470 17870 -1440
rect 17840 -1510 17870 -1480
rect 17840 -1525 17870 -1520
rect 17840 -1545 17845 -1525
rect 17845 -1545 17865 -1525
rect 17865 -1545 17870 -1525
rect 17840 -1550 17870 -1545
rect 17950 -1470 17980 -1440
rect 17950 -1510 17980 -1480
rect 17950 -1525 17980 -1520
rect 17950 -1545 17955 -1525
rect 17955 -1545 17975 -1525
rect 17975 -1545 17980 -1525
rect 17950 -1550 17980 -1545
rect 18010 -1470 18040 -1440
rect 18010 -1510 18040 -1480
rect 18010 -1525 18040 -1520
rect 18010 -1545 18015 -1525
rect 18015 -1545 18035 -1525
rect 18035 -1545 18040 -1525
rect 18010 -1550 18040 -1545
rect 18155 -1470 18185 -1440
rect 18155 -1510 18185 -1480
rect 18155 -1525 18185 -1520
rect 18155 -1545 18160 -1525
rect 18160 -1545 18180 -1525
rect 18180 -1545 18185 -1525
rect 18155 -1550 18185 -1545
rect 18265 -1470 18295 -1440
rect 18265 -1510 18295 -1480
rect 18265 -1525 18295 -1520
rect 18265 -1545 18270 -1525
rect 18270 -1545 18290 -1525
rect 18290 -1545 18295 -1525
rect 18265 -1550 18295 -1545
rect 18375 -1470 18405 -1440
rect 18375 -1510 18405 -1480
rect 18375 -1525 18405 -1520
rect 18375 -1545 18380 -1525
rect 18380 -1545 18400 -1525
rect 18400 -1545 18405 -1525
rect 18375 -1550 18405 -1545
rect 18485 -1470 18515 -1440
rect 18485 -1510 18515 -1480
rect 18485 -1525 18515 -1520
rect 18485 -1545 18490 -1525
rect 18490 -1545 18510 -1525
rect 18510 -1545 18515 -1525
rect 18485 -1550 18515 -1545
rect 18595 -1470 18625 -1440
rect 18595 -1510 18625 -1480
rect 18595 -1525 18625 -1520
rect 18595 -1545 18600 -1525
rect 18600 -1545 18620 -1525
rect 18620 -1545 18625 -1525
rect 18595 -1550 18625 -1545
rect 17195 -1695 17225 -1690
rect 17195 -1715 17200 -1695
rect 17200 -1715 17220 -1695
rect 17220 -1715 17225 -1695
rect 17195 -1720 17225 -1715
rect 17085 -1775 17115 -1745
rect 17415 -1695 17445 -1690
rect 17415 -1715 17420 -1695
rect 17420 -1715 17440 -1695
rect 17440 -1715 17445 -1695
rect 17415 -1720 17445 -1715
rect 17675 -1695 17705 -1690
rect 17675 -1715 17680 -1695
rect 17680 -1715 17700 -1695
rect 17700 -1715 17705 -1695
rect 17675 -1720 17705 -1715
rect 17785 -1695 17815 -1690
rect 17785 -1715 17790 -1695
rect 17790 -1715 17810 -1695
rect 17810 -1715 17815 -1695
rect 17785 -1720 17815 -1715
rect 17895 -1695 17925 -1690
rect 17895 -1715 17900 -1695
rect 17900 -1715 17920 -1695
rect 17920 -1715 17925 -1695
rect 17895 -1720 17925 -1715
rect 18210 -1695 18240 -1690
rect 18210 -1715 18215 -1695
rect 18215 -1715 18235 -1695
rect 18235 -1715 18240 -1695
rect 18210 -1720 18240 -1715
rect 18430 -1695 18460 -1690
rect 18430 -1715 18435 -1695
rect 18435 -1715 18455 -1695
rect 18455 -1715 18460 -1695
rect 18430 -1720 18460 -1715
rect 17305 -1775 17335 -1745
rect 17195 -1830 17225 -1800
rect 16770 -1885 16800 -1855
rect 18320 -1775 18350 -1745
rect 18540 -1775 18570 -1745
rect 18890 -1780 18920 -1750
rect 18430 -1830 18460 -1800
rect 17785 -1920 17815 -1890
rect 16320 -2030 16350 -2000
rect 17430 -2005 17465 -2000
rect 17430 -2030 17435 -2005
rect 17435 -2030 17460 -2005
rect 17460 -2030 17465 -2005
rect 17430 -2035 17465 -2030
rect 18129 -2005 18164 -2000
rect 18129 -2030 18134 -2005
rect 18134 -2030 18159 -2005
rect 18159 -2030 18164 -2005
rect 18129 -2035 18164 -2030
rect 18835 -2035 18865 -2005
rect 17430 -2090 17460 -2060
rect 16265 -2130 16295 -2100
rect 16485 -2130 16515 -2100
rect 16735 -2130 16765 -2100
rect 16485 -2905 16520 -2900
rect 16485 -2930 16490 -2905
rect 16490 -2930 16515 -2905
rect 16515 -2930 16520 -2905
rect 16485 -2935 16520 -2930
rect 16160 -3030 16195 -3025
rect 16160 -3055 16165 -3030
rect 16165 -3055 16190 -3030
rect 16190 -3055 16195 -3030
rect 16160 -3060 16195 -3055
rect 15825 -3145 15855 -3115
rect 15950 -3121 15985 -3116
rect 15950 -3146 15955 -3121
rect 15955 -3146 15980 -3121
rect 15980 -3146 15985 -3121
rect 16735 -3135 16765 -3105
rect 15950 -3151 15985 -3146
rect 17785 -3135 17815 -3105
rect 18620 -3135 18650 -3105
rect 18835 -3135 18865 -3105
rect 15950 -3794 15985 -3789
rect 15950 -3819 15955 -3794
rect 15955 -3819 15980 -3794
rect 15980 -3819 15985 -3794
rect 15950 -3824 15985 -3819
rect 15825 -4285 15855 -4255
rect 15650 -4375 15680 -4345
rect 15690 -4375 15720 -4345
rect 15730 -4375 15760 -4345
rect 15650 -4415 15680 -4385
rect 15690 -4415 15720 -4385
rect 15730 -4415 15760 -4385
rect 15650 -4455 15680 -4425
rect 15690 -4455 15720 -4425
rect 15730 -4455 15760 -4425
rect 16280 -3899 16315 -3894
rect 16280 -3924 16285 -3899
rect 16285 -3924 16310 -3899
rect 16310 -3924 16315 -3899
rect 16280 -3929 16315 -3924
rect 16605 -3974 16640 -3969
rect 16605 -3999 16610 -3974
rect 16610 -3999 16635 -3974
rect 16635 -3999 16640 -3974
rect 16605 -4004 16640 -3999
rect 16285 -4140 16315 -4110
rect 16285 -4180 16315 -4150
rect 16285 -4220 16315 -4190
rect 16610 -4140 16640 -4110
rect 16610 -4180 16640 -4150
rect 16610 -4220 16640 -4190
rect 17785 -4210 17815 -4205
rect 17785 -4230 17790 -4210
rect 17790 -4230 17810 -4210
rect 17810 -4230 17815 -4210
rect 17785 -4235 17815 -4230
rect 17260 -4285 17290 -4255
rect 17785 -4250 17815 -4245
rect 17785 -4270 17790 -4250
rect 17790 -4270 17810 -4250
rect 17810 -4270 17815 -4250
rect 17785 -4275 17815 -4270
rect 17785 -4290 17815 -4285
rect 17785 -4310 17790 -4290
rect 17790 -4310 17810 -4290
rect 17810 -4310 17815 -4290
rect 17785 -4315 17815 -4310
rect 16910 -4365 16940 -4335
rect 16910 -4415 16940 -4385
rect 16910 -4465 16940 -4435
rect 15955 -4510 15985 -4480
rect 16210 -4510 16240 -4480
rect 18660 -4500 18690 -4470
rect 19095 -1780 19125 -1750
rect 19330 -530 19360 -500
rect 19330 -1975 19360 -1945
rect 19410 345 19440 375
rect 19410 -210 19440 -180
rect 19085 -2090 19115 -2060
rect 19080 -2905 19115 -2900
rect 19080 -2930 19085 -2905
rect 19085 -2930 19110 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2935 19115 -2930
rect 19615 1430 19645 1460
rect 19615 605 19645 635
rect 19615 155 19645 185
rect 19540 -1920 19570 -1890
rect 19405 -3002 19440 -2997
rect 19405 -3027 19410 -3002
rect 19410 -3027 19435 -3002
rect 19435 -3027 19440 -3002
rect 19405 -3032 19440 -3027
rect 19780 -1830 19810 -1800
rect 19610 -3120 19645 -3115
rect 19610 -3145 19615 -3120
rect 19615 -3145 19640 -3120
rect 19640 -3145 19645 -3120
rect 19610 -3150 19645 -3145
rect 19610 -3794 19645 -3789
rect 19610 -3819 19615 -3794
rect 19615 -3819 19640 -3794
rect 19640 -3819 19645 -3794
rect 19610 -3824 19645 -3819
rect 19285 -3899 19320 -3894
rect 19285 -3924 19290 -3899
rect 19290 -3924 19315 -3899
rect 19315 -3924 19320 -3899
rect 19285 -3929 19320 -3924
rect 18960 -3974 18995 -3969
rect 18960 -3999 18965 -3974
rect 18965 -3999 18990 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4004 18995 -3999
rect 18960 -4235 18990 -4205
rect 18960 -4275 18990 -4245
rect 18960 -4315 18990 -4285
rect 19285 -4235 19315 -4205
rect 19285 -4275 19315 -4245
rect 19285 -4315 19315 -4285
rect 18890 -4500 18920 -4470
rect 19360 -4500 19390 -4470
rect 19615 -4500 19645 -4470
rect 17960 -4550 17990 -4520
<< metal2 >>
rect 16485 1460 18500 1465
rect 18590 1460 19650 1465
rect 16485 1430 16490 1460
rect 16520 1430 17055 1460
rect 17085 1430 17785 1460
rect 17815 1430 18515 1460
rect 18545 1430 19615 1460
rect 19645 1430 19650 1460
rect 16485 1425 19650 1430
rect 16365 1405 18715 1410
rect 16365 1375 16370 1405
rect 16400 1375 16490 1405
rect 16520 1375 16610 1405
rect 16640 1375 16890 1405
rect 16920 1375 17000 1405
rect 17030 1375 17110 1405
rect 17140 1375 17220 1405
rect 17250 1375 17500 1405
rect 17530 1375 17565 1405
rect 17595 1375 17675 1405
rect 17705 1375 17785 1405
rect 17815 1375 17895 1405
rect 17925 1375 18005 1405
rect 18035 1375 18070 1405
rect 18100 1375 18350 1405
rect 18380 1375 18460 1405
rect 18490 1375 18570 1405
rect 18600 1375 18680 1405
rect 18710 1375 18715 1405
rect 16365 1365 18715 1375
rect 16365 1335 16370 1365
rect 16400 1335 16490 1365
rect 16520 1335 16610 1365
rect 16640 1335 16890 1365
rect 16920 1335 17000 1365
rect 17030 1335 17110 1365
rect 17140 1335 17220 1365
rect 17250 1335 17500 1365
rect 17530 1335 17565 1365
rect 17595 1335 17675 1365
rect 17705 1335 17785 1365
rect 17815 1335 17895 1365
rect 17925 1335 18005 1365
rect 18035 1335 18070 1365
rect 18100 1335 18350 1365
rect 18380 1335 18460 1365
rect 18490 1335 18570 1365
rect 18600 1335 18680 1365
rect 18710 1335 18715 1365
rect 16365 1325 18715 1335
rect 16365 1295 16370 1325
rect 16400 1295 16490 1325
rect 16520 1295 16610 1325
rect 16640 1295 16890 1325
rect 16920 1295 17000 1325
rect 17030 1295 17110 1325
rect 17140 1295 17220 1325
rect 17250 1295 17500 1325
rect 17530 1295 17565 1325
rect 17595 1295 17675 1325
rect 17705 1295 17785 1325
rect 17815 1295 17895 1325
rect 17925 1295 18005 1325
rect 18035 1295 18070 1325
rect 18100 1295 18350 1325
rect 18380 1295 18460 1325
rect 18490 1295 18570 1325
rect 18600 1295 18680 1325
rect 18710 1295 18715 1325
rect 16365 1290 18715 1295
rect 15890 1155 16470 1160
rect 15890 1125 15895 1155
rect 15925 1125 16435 1155
rect 16465 1125 16470 1155
rect 15890 1120 16470 1125
rect 16540 1155 16580 1160
rect 16540 1125 16545 1155
rect 16575 1125 16580 1155
rect 16540 1120 16580 1125
rect 16940 1155 16980 1160
rect 16940 1125 16945 1155
rect 16975 1150 16980 1155
rect 17050 1155 17090 1160
rect 17050 1150 17055 1155
rect 16975 1130 17055 1150
rect 16975 1125 16980 1130
rect 16940 1120 16980 1125
rect 17050 1125 17055 1130
rect 17085 1150 17090 1155
rect 17160 1155 17200 1160
rect 17160 1150 17165 1155
rect 17085 1130 17165 1150
rect 17085 1125 17090 1130
rect 17050 1120 17090 1125
rect 17160 1125 17165 1130
rect 17195 1125 17200 1155
rect 17160 1120 17200 1125
rect 17615 1155 17655 1160
rect 17615 1125 17620 1155
rect 17650 1150 17655 1155
rect 17725 1155 17765 1160
rect 17725 1150 17730 1155
rect 17650 1130 17730 1150
rect 17650 1125 17655 1130
rect 17615 1120 17655 1125
rect 17725 1125 17730 1130
rect 17760 1150 17765 1155
rect 17835 1155 17875 1160
rect 17835 1150 17840 1155
rect 17760 1130 17840 1150
rect 17760 1125 17765 1130
rect 17725 1120 17765 1125
rect 17835 1125 17840 1130
rect 17870 1150 17875 1155
rect 17945 1155 17985 1160
rect 17945 1150 17950 1155
rect 17870 1130 17950 1150
rect 17870 1125 17875 1130
rect 17835 1120 17875 1125
rect 17945 1125 17950 1130
rect 17980 1125 17985 1155
rect 17945 1120 17985 1125
rect 18400 1155 18440 1160
rect 18400 1125 18405 1155
rect 18435 1150 18440 1155
rect 18510 1155 18550 1160
rect 18510 1150 18515 1155
rect 18435 1130 18515 1150
rect 18435 1125 18440 1130
rect 18400 1120 18440 1125
rect 18510 1125 18515 1130
rect 18545 1150 18550 1155
rect 18620 1155 18660 1160
rect 18620 1150 18625 1155
rect 18545 1130 18625 1150
rect 18545 1125 18550 1130
rect 18510 1120 18550 1125
rect 18620 1125 18625 1130
rect 18655 1125 18660 1155
rect 18620 1120 18660 1125
rect 16540 1100 19365 1105
rect 16540 1070 16545 1100
rect 16575 1070 19330 1100
rect 19360 1070 19365 1100
rect 16540 1065 19365 1070
rect 16435 1045 18630 1050
rect 16435 1015 16440 1045
rect 16470 1015 16660 1045
rect 16690 1015 16975 1045
rect 17005 1015 17155 1045
rect 17185 1015 17335 1045
rect 17365 1015 17515 1045
rect 17545 1015 17695 1045
rect 17725 1015 17875 1045
rect 17905 1015 18055 1045
rect 18085 1015 18235 1045
rect 18265 1015 18415 1045
rect 18445 1015 18595 1045
rect 18625 1015 18630 1045
rect 16435 1005 18630 1015
rect 16435 975 16440 1005
rect 16470 975 16660 1005
rect 16690 975 16975 1005
rect 17005 975 17155 1005
rect 17185 975 17335 1005
rect 17365 975 17515 1005
rect 17545 975 17695 1005
rect 17725 975 17875 1005
rect 17905 975 18055 1005
rect 18085 975 18235 1005
rect 18265 975 18415 1005
rect 18445 975 18595 1005
rect 18625 975 18630 1005
rect 16435 965 18630 975
rect 16435 935 16440 965
rect 16470 935 16660 965
rect 16690 935 16975 965
rect 17005 935 17155 965
rect 17185 935 17335 965
rect 17365 935 17515 965
rect 17545 935 17695 965
rect 17725 935 17875 965
rect 17905 935 18055 965
rect 18085 935 18235 965
rect 18265 935 18415 965
rect 18445 935 18595 965
rect 18625 935 18630 965
rect 16435 930 18630 935
rect 18905 1045 19115 1050
rect 18905 1015 18910 1045
rect 18940 1015 19020 1045
rect 19050 1015 19080 1045
rect 19110 1015 19115 1045
rect 18905 1005 19115 1015
rect 18905 975 18910 1005
rect 18940 975 19020 1005
rect 19050 975 19080 1005
rect 19110 975 19115 1005
rect 18905 965 19115 975
rect 18905 935 18910 965
rect 18940 935 19020 965
rect 19050 935 19080 965
rect 19110 935 19115 965
rect 18905 930 19115 935
rect 16545 865 16585 870
rect 16545 835 16550 865
rect 16580 860 16585 865
rect 16780 865 16820 870
rect 16780 860 16785 865
rect 16580 840 16785 860
rect 16580 835 16585 840
rect 16545 830 16585 835
rect 16780 835 16785 840
rect 16815 835 16820 865
rect 16780 830 16820 835
rect 16480 695 16650 700
rect 16480 665 16485 695
rect 16515 665 16615 695
rect 16645 665 16650 695
rect 16480 660 16650 665
rect 19000 635 19650 640
rect 19000 605 19005 635
rect 19035 605 19615 635
rect 19645 605 19650 635
rect 19000 600 19650 605
rect 17110 595 18490 600
rect 17140 565 17200 595
rect 17230 565 17290 595
rect 17320 565 17380 595
rect 17410 565 17470 595
rect 17500 565 17560 595
rect 17590 565 17650 595
rect 17680 565 17695 595
rect 17725 565 17740 595
rect 17770 565 17830 595
rect 17860 565 17920 595
rect 17950 565 18010 595
rect 18040 565 18100 595
rect 18130 565 18190 595
rect 18220 565 18280 595
rect 18310 565 18370 595
rect 18400 565 18460 595
rect 17110 560 18490 565
rect 16315 540 16355 545
rect 16315 510 16320 540
rect 16350 535 16355 540
rect 17600 540 17640 545
rect 17600 535 17605 540
rect 16350 515 17605 535
rect 16350 510 16355 515
rect 16315 505 16355 510
rect 17600 510 17605 515
rect 17635 535 17640 540
rect 17960 540 18000 545
rect 17960 535 17965 540
rect 17635 515 17965 535
rect 17635 510 17640 515
rect 17600 505 17640 510
rect 17960 510 17965 515
rect 17995 510 18000 540
rect 17960 505 18000 510
rect 16260 485 16300 490
rect 16260 455 16265 485
rect 16295 480 16300 485
rect 16780 485 16820 490
rect 16780 480 16785 485
rect 16295 460 16785 480
rect 16295 455 16300 460
rect 16260 450 16300 455
rect 16780 455 16785 460
rect 16815 480 16820 485
rect 17420 485 17460 490
rect 17420 480 17425 485
rect 16815 460 17425 480
rect 16815 455 16820 460
rect 16780 450 16820 455
rect 17420 455 17425 460
rect 17455 480 17460 485
rect 18140 485 18180 490
rect 18140 480 18145 485
rect 17455 460 18145 480
rect 17455 455 17460 460
rect 17420 450 17460 455
rect 18140 455 18145 460
rect 18175 455 18180 485
rect 18140 450 18180 455
rect 16205 430 16245 435
rect 16205 400 16210 430
rect 16240 425 16245 430
rect 16545 430 16585 435
rect 16545 425 16550 430
rect 16240 405 16550 425
rect 16240 400 16245 405
rect 16205 395 16245 400
rect 16545 400 16550 405
rect 16580 425 16585 430
rect 17240 430 17280 435
rect 17240 425 17245 430
rect 16580 405 17245 425
rect 16580 400 16585 405
rect 16545 395 16585 400
rect 17240 400 17245 405
rect 17275 425 17280 430
rect 18320 430 18360 435
rect 18320 425 18325 430
rect 17275 405 18325 425
rect 17275 400 17280 405
rect 17240 395 17280 400
rect 18320 400 18325 405
rect 18355 400 18360 430
rect 18320 395 18360 400
rect 17060 375 19445 380
rect 17060 345 17065 375
rect 17095 345 17785 375
rect 17815 345 18505 375
rect 18535 345 19410 375
rect 19440 345 19445 375
rect 17060 340 19445 345
rect 16420 320 19180 325
rect 16420 290 16425 320
rect 16455 290 16545 320
rect 16575 290 16665 320
rect 16695 290 16785 320
rect 16815 290 16905 320
rect 16935 290 17025 320
rect 17055 290 17145 320
rect 17175 290 17265 320
rect 17295 290 17385 320
rect 17415 290 17505 320
rect 17535 290 17625 320
rect 17655 290 17945 320
rect 17975 290 18065 320
rect 18095 290 18185 320
rect 18215 290 18305 320
rect 18335 290 18425 320
rect 18455 290 18545 320
rect 18575 290 18665 320
rect 18695 290 18785 320
rect 18815 290 18905 320
rect 18935 290 19025 320
rect 19055 290 19145 320
rect 19175 290 19180 320
rect 16420 280 19180 290
rect 16420 250 16425 280
rect 16455 250 16545 280
rect 16575 250 16665 280
rect 16695 250 16785 280
rect 16815 250 16905 280
rect 16935 250 17025 280
rect 17055 250 17145 280
rect 17175 250 17265 280
rect 17295 250 17385 280
rect 17415 250 17505 280
rect 17535 250 17625 280
rect 17655 250 17945 280
rect 17975 250 18065 280
rect 18095 250 18185 280
rect 18215 250 18305 280
rect 18335 250 18425 280
rect 18455 250 18545 280
rect 18575 250 18665 280
rect 18695 250 18785 280
rect 18815 250 18905 280
rect 18935 250 19025 280
rect 19055 250 19145 280
rect 19175 250 19180 280
rect 16420 240 19180 250
rect 16420 210 16425 240
rect 16455 210 16545 240
rect 16575 210 16665 240
rect 16695 210 16785 240
rect 16815 210 16905 240
rect 16935 210 17025 240
rect 17055 210 17145 240
rect 17175 210 17265 240
rect 17295 210 17385 240
rect 17415 210 17505 240
rect 17535 210 17625 240
rect 17655 210 17945 240
rect 17975 210 18065 240
rect 18095 210 18185 240
rect 18215 210 18305 240
rect 18335 210 18425 240
rect 18455 210 18545 240
rect 18575 210 18665 240
rect 18695 210 18785 240
rect 18815 210 18905 240
rect 18935 210 19025 240
rect 19055 210 19145 240
rect 19175 210 19180 240
rect 16420 205 19180 210
rect 15945 185 17730 190
rect 15945 155 15950 185
rect 15980 155 16485 185
rect 16515 155 16845 185
rect 16875 155 17205 185
rect 17235 155 17565 185
rect 17595 155 17695 185
rect 17725 155 17730 185
rect 15945 150 17730 155
rect 17870 185 19650 190
rect 17870 155 17875 185
rect 17905 155 18005 185
rect 18035 155 18365 185
rect 18395 155 18725 185
rect 18755 155 19085 185
rect 19115 155 19615 185
rect 19645 155 19650 185
rect 17870 150 19650 155
rect 16845 130 16875 150
rect 18725 135 18755 150
rect 16600 15 16640 20
rect 16600 -15 16605 15
rect 16635 10 16640 15
rect 16960 15 17000 20
rect 16960 10 16965 15
rect 16635 -10 16965 10
rect 16635 -15 16640 -10
rect 16600 -20 16640 -15
rect 16960 -15 16965 -10
rect 16995 10 17000 15
rect 17320 15 17360 20
rect 17320 10 17325 15
rect 16995 -10 17325 10
rect 16995 -15 17000 -10
rect 16960 -20 17000 -15
rect 17320 -15 17325 -10
rect 17355 -15 17360 15
rect 17320 -20 17360 -15
rect 18240 15 18280 20
rect 18240 -15 18245 15
rect 18275 10 18280 15
rect 18600 15 18640 20
rect 18600 10 18605 15
rect 18275 -10 18605 10
rect 18275 -15 18280 -10
rect 18240 -20 18280 -15
rect 18600 -15 18605 -10
rect 18635 10 18640 15
rect 18960 15 19000 20
rect 18960 10 18965 15
rect 18635 -10 18965 10
rect 18635 -15 18640 -10
rect 18600 -20 18640 -15
rect 18960 -15 18965 -10
rect 18995 -15 19000 15
rect 18960 -20 19000 -15
rect 15645 -45 17570 -40
rect 15645 -75 15650 -45
rect 15680 -75 15690 -45
rect 15720 -75 15730 -45
rect 15760 -75 16515 -45
rect 16545 -75 16725 -45
rect 16755 -75 16845 -45
rect 16875 -75 17085 -45
rect 17115 -75 17205 -45
rect 17235 -75 17445 -45
rect 17475 -75 17535 -45
rect 17565 -75 17570 -45
rect 15645 -85 17570 -75
rect 18030 -45 19130 -40
rect 18030 -75 18035 -45
rect 18065 -75 18125 -45
rect 18155 -75 18365 -45
rect 18395 -75 18485 -45
rect 18515 -75 18725 -45
rect 18755 -75 18845 -45
rect 18875 -75 19055 -45
rect 19085 -75 19095 -45
rect 19125 -75 19130 -45
rect 18030 -80 19130 -75
rect 15645 -115 15650 -85
rect 15680 -115 15690 -85
rect 15720 -115 15730 -85
rect 15760 -115 16515 -85
rect 16545 -115 16725 -85
rect 16755 -115 16845 -85
rect 16875 -115 17085 -85
rect 17115 -115 17205 -85
rect 17235 -115 17445 -85
rect 17475 -115 17535 -85
rect 17565 -115 17570 -85
rect 15645 -125 17570 -115
rect 15645 -155 15650 -125
rect 15680 -155 15690 -125
rect 15720 -155 15730 -125
rect 15760 -155 16515 -125
rect 16545 -155 16725 -125
rect 16755 -155 16845 -125
rect 16875 -155 17085 -125
rect 17115 -155 17205 -125
rect 17235 -155 17445 -125
rect 17475 -155 17535 -125
rect 17565 -155 17570 -125
rect 15645 -160 17570 -155
rect 16260 -180 16300 -175
rect 16260 -210 16265 -180
rect 16295 -185 16300 -180
rect 17005 -180 17037 -175
rect 17005 -185 17007 -180
rect 16295 -205 17007 -185
rect 16295 -210 16300 -205
rect 16260 -215 16300 -210
rect 17005 -210 17007 -205
rect 18563 -180 19445 -175
rect 18562 -205 18563 -185
rect 17005 -215 17037 -210
rect 18593 -210 19410 -180
rect 19440 -210 19445 -180
rect 18563 -215 19445 -210
rect 17560 -240 18040 -235
rect 17560 -270 17565 -240
rect 17595 -270 17745 -240
rect 17775 -270 17785 -240
rect 17815 -270 17825 -240
rect 17855 -270 18005 -240
rect 18035 -270 18040 -240
rect 17560 -280 18040 -270
rect 17560 -310 17565 -280
rect 17595 -310 17745 -280
rect 17775 -310 17785 -280
rect 17815 -310 17825 -280
rect 17855 -310 18005 -280
rect 18035 -310 18040 -280
rect 17560 -320 18040 -310
rect 17560 -350 17565 -320
rect 17595 -350 17745 -320
rect 17775 -350 17785 -320
rect 17815 -350 17825 -320
rect 17855 -350 18005 -320
rect 18035 -350 18040 -320
rect 17560 -355 18040 -350
rect 16315 -500 16355 -495
rect 16315 -530 16320 -500
rect 16350 -505 16355 -500
rect 17075 -500 17105 -495
rect 16350 -525 17075 -505
rect 16350 -530 16355 -525
rect 16315 -535 16355 -530
rect 17075 -535 17105 -530
rect 18440 -500 19365 -495
rect 18470 -530 19330 -500
rect 19360 -530 19365 -500
rect 18440 -535 19365 -530
rect 16530 -610 17060 -605
rect 16530 -640 16535 -610
rect 16565 -640 17025 -610
rect 17055 -640 17060 -610
rect 16530 -645 17060 -640
rect 18540 -610 19070 -605
rect 18540 -640 18545 -610
rect 18575 -640 19035 -610
rect 19065 -640 19070 -610
rect 18540 -645 19070 -640
rect 16620 -665 18980 -660
rect 16620 -695 16625 -665
rect 16655 -695 16745 -665
rect 16775 -695 16865 -665
rect 16895 -695 16985 -665
rect 17015 -695 17305 -665
rect 17335 -695 17425 -665
rect 17455 -695 17545 -665
rect 17575 -695 18025 -665
rect 18055 -695 18145 -665
rect 18175 -695 18265 -665
rect 18295 -695 18585 -665
rect 18615 -695 18705 -665
rect 18735 -695 18825 -665
rect 18855 -695 18945 -665
rect 18975 -695 18980 -665
rect 16620 -705 18980 -695
rect 16620 -735 16625 -705
rect 16655 -735 16745 -705
rect 16775 -735 16865 -705
rect 16895 -735 16985 -705
rect 17015 -735 17305 -705
rect 17335 -735 17425 -705
rect 17455 -735 17545 -705
rect 17575 -735 18025 -705
rect 18055 -735 18145 -705
rect 18175 -735 18265 -705
rect 18295 -735 18585 -705
rect 18615 -735 18705 -705
rect 18735 -735 18825 -705
rect 18855 -735 18945 -705
rect 18975 -735 18980 -705
rect 16620 -745 18980 -735
rect 16620 -775 16625 -745
rect 16655 -775 16745 -745
rect 16775 -775 16865 -745
rect 16895 -775 16985 -745
rect 17015 -775 17305 -745
rect 17335 -775 17425 -745
rect 17455 -775 17545 -745
rect 17575 -775 18025 -745
rect 18055 -775 18145 -745
rect 18175 -775 18265 -745
rect 18295 -775 18585 -745
rect 18615 -775 18705 -745
rect 18735 -775 18825 -745
rect 18855 -775 18945 -745
rect 18975 -775 18980 -745
rect 16620 -780 18980 -775
rect 17110 -1065 18490 -1060
rect 17110 -1095 17115 -1065
rect 17145 -1095 17745 -1065
rect 17775 -1095 17785 -1065
rect 17815 -1095 17825 -1065
rect 17855 -1095 18455 -1065
rect 18485 -1095 18490 -1065
rect 17110 -1105 18490 -1095
rect 17110 -1135 17115 -1105
rect 17145 -1135 17745 -1105
rect 17775 -1135 17785 -1105
rect 17815 -1135 17825 -1105
rect 17855 -1135 18455 -1105
rect 18485 -1135 18490 -1105
rect 17110 -1145 18490 -1135
rect 17110 -1175 17115 -1145
rect 17145 -1175 17745 -1145
rect 17775 -1175 17785 -1145
rect 17815 -1175 17825 -1145
rect 17855 -1175 18455 -1145
rect 18485 -1175 18490 -1145
rect 17110 -1180 18490 -1175
rect 16740 -1200 16780 -1195
rect 16740 -1230 16745 -1200
rect 16775 -1205 16780 -1200
rect 16820 -1200 16860 -1195
rect 16820 -1205 16825 -1200
rect 16775 -1225 16825 -1205
rect 16775 -1230 16780 -1225
rect 16740 -1235 16780 -1230
rect 16820 -1230 16825 -1225
rect 16855 -1205 16860 -1200
rect 16900 -1200 16940 -1195
rect 16900 -1205 16905 -1200
rect 16855 -1225 16905 -1205
rect 16855 -1230 16860 -1225
rect 16820 -1235 16860 -1230
rect 16900 -1230 16905 -1225
rect 16935 -1205 16940 -1200
rect 16980 -1200 17020 -1195
rect 16980 -1205 16985 -1200
rect 16935 -1225 16985 -1205
rect 16935 -1230 16940 -1225
rect 16900 -1235 16940 -1230
rect 16980 -1230 16985 -1225
rect 17015 -1205 17020 -1200
rect 17060 -1200 17100 -1195
rect 17060 -1205 17065 -1200
rect 17015 -1225 17065 -1205
rect 17015 -1230 17020 -1225
rect 16980 -1235 17020 -1230
rect 17060 -1230 17065 -1225
rect 17095 -1205 17100 -1200
rect 17140 -1200 17180 -1195
rect 17140 -1205 17145 -1200
rect 17095 -1225 17145 -1205
rect 17095 -1230 17100 -1225
rect 17060 -1235 17100 -1230
rect 17140 -1230 17145 -1225
rect 17175 -1205 17180 -1200
rect 17220 -1200 17260 -1195
rect 17220 -1205 17225 -1200
rect 17175 -1225 17225 -1205
rect 17175 -1230 17180 -1225
rect 17140 -1235 17180 -1230
rect 17220 -1230 17225 -1225
rect 17255 -1205 17260 -1200
rect 17300 -1200 17340 -1195
rect 17300 -1205 17305 -1200
rect 17255 -1225 17305 -1205
rect 17255 -1230 17260 -1225
rect 17220 -1235 17260 -1230
rect 17300 -1230 17305 -1225
rect 17335 -1205 17340 -1200
rect 17380 -1200 17420 -1195
rect 17380 -1205 17385 -1200
rect 17335 -1225 17385 -1205
rect 17335 -1230 17340 -1225
rect 17300 -1235 17340 -1230
rect 17380 -1230 17385 -1225
rect 17415 -1205 17420 -1200
rect 17460 -1200 17500 -1195
rect 17460 -1205 17465 -1200
rect 17415 -1225 17465 -1205
rect 17415 -1230 17420 -1225
rect 17380 -1235 17420 -1230
rect 17460 -1230 17465 -1225
rect 17495 -1205 17500 -1200
rect 17540 -1200 17580 -1195
rect 17540 -1205 17545 -1200
rect 17495 -1225 17545 -1205
rect 17495 -1230 17500 -1225
rect 17460 -1235 17500 -1230
rect 17540 -1230 17545 -1225
rect 17575 -1205 17580 -1200
rect 17620 -1200 17660 -1195
rect 17620 -1205 17625 -1200
rect 17575 -1225 17625 -1205
rect 17575 -1230 17580 -1225
rect 17540 -1235 17580 -1230
rect 17620 -1230 17625 -1225
rect 17655 -1205 17660 -1200
rect 17700 -1200 17740 -1195
rect 17700 -1205 17705 -1200
rect 17655 -1225 17705 -1205
rect 17655 -1230 17660 -1225
rect 17620 -1235 17660 -1230
rect 17700 -1230 17705 -1225
rect 17735 -1230 17740 -1200
rect 17700 -1235 17740 -1230
rect 17780 -1200 17820 -1195
rect 17780 -1230 17785 -1200
rect 17815 -1205 17820 -1200
rect 17860 -1200 17900 -1195
rect 17860 -1205 17865 -1200
rect 17815 -1225 17865 -1205
rect 17815 -1230 17820 -1225
rect 17780 -1235 17820 -1230
rect 17860 -1230 17865 -1225
rect 17895 -1205 17900 -1200
rect 17940 -1200 17980 -1195
rect 17940 -1205 17945 -1200
rect 17895 -1225 17945 -1205
rect 17895 -1230 17900 -1225
rect 17860 -1235 17900 -1230
rect 17940 -1230 17945 -1225
rect 17975 -1205 17980 -1200
rect 18020 -1200 18060 -1195
rect 18020 -1205 18025 -1200
rect 17975 -1225 18025 -1205
rect 17975 -1230 17980 -1225
rect 17940 -1235 17980 -1230
rect 18020 -1230 18025 -1225
rect 18055 -1205 18060 -1200
rect 18100 -1200 18140 -1195
rect 18100 -1205 18105 -1200
rect 18055 -1225 18105 -1205
rect 18055 -1230 18060 -1225
rect 18020 -1235 18060 -1230
rect 18100 -1230 18105 -1225
rect 18135 -1205 18140 -1200
rect 18180 -1200 18220 -1195
rect 18180 -1205 18185 -1200
rect 18135 -1225 18185 -1205
rect 18135 -1230 18140 -1225
rect 18100 -1235 18140 -1230
rect 18180 -1230 18185 -1225
rect 18215 -1205 18220 -1200
rect 18260 -1200 18300 -1195
rect 18260 -1205 18265 -1200
rect 18215 -1225 18265 -1205
rect 18215 -1230 18220 -1225
rect 18180 -1235 18220 -1230
rect 18260 -1230 18265 -1225
rect 18295 -1205 18300 -1200
rect 18340 -1200 18380 -1195
rect 18340 -1205 18345 -1200
rect 18295 -1225 18345 -1205
rect 18295 -1230 18300 -1225
rect 18260 -1235 18300 -1230
rect 18340 -1230 18345 -1225
rect 18375 -1205 18380 -1200
rect 18420 -1200 18460 -1195
rect 18420 -1205 18425 -1200
rect 18375 -1225 18425 -1205
rect 18375 -1230 18380 -1225
rect 18340 -1235 18380 -1230
rect 18420 -1230 18425 -1225
rect 18455 -1205 18460 -1200
rect 18500 -1200 18540 -1195
rect 18500 -1205 18505 -1200
rect 18455 -1225 18505 -1205
rect 18455 -1230 18460 -1225
rect 18420 -1235 18460 -1230
rect 18500 -1230 18505 -1225
rect 18535 -1205 18540 -1200
rect 18580 -1200 18620 -1195
rect 18580 -1205 18585 -1200
rect 18535 -1225 18585 -1205
rect 18535 -1230 18540 -1225
rect 18500 -1235 18540 -1230
rect 18580 -1230 18585 -1225
rect 18615 -1205 18620 -1200
rect 18660 -1200 18700 -1195
rect 18660 -1205 18665 -1200
rect 18615 -1225 18665 -1205
rect 18615 -1230 18620 -1225
rect 18580 -1235 18620 -1230
rect 18660 -1230 18665 -1225
rect 18695 -1205 18700 -1200
rect 18740 -1200 18780 -1195
rect 18740 -1205 18745 -1200
rect 18695 -1225 18745 -1205
rect 18695 -1230 18700 -1225
rect 18660 -1235 18700 -1230
rect 18740 -1230 18745 -1225
rect 18775 -1230 18780 -1200
rect 18740 -1235 18780 -1230
rect 18895 -1265 18935 -1260
rect 16205 -1285 16245 -1280
rect 16205 -1315 16210 -1285
rect 16240 -1290 16245 -1285
rect 16700 -1285 16740 -1280
rect 16700 -1290 16705 -1285
rect 16240 -1310 16705 -1290
rect 16240 -1315 16245 -1310
rect 16205 -1320 16245 -1315
rect 16700 -1315 16705 -1310
rect 16735 -1315 16740 -1285
rect 16700 -1320 16740 -1315
rect 18895 -1295 18900 -1265
rect 18930 -1295 18935 -1265
rect 18895 -1305 18935 -1295
rect 18895 -1335 18900 -1305
rect 18930 -1335 18935 -1305
rect 18895 -1340 18935 -1335
rect 15890 -1385 18355 -1380
rect 15890 -1415 15895 -1385
rect 15925 -1415 16660 -1385
rect 16690 -1415 16770 -1385
rect 16800 -1415 17305 -1385
rect 17335 -1415 17785 -1385
rect 17815 -1415 18320 -1385
rect 18350 -1415 18355 -1385
rect 15890 -1420 18355 -1415
rect 16600 -1440 18630 -1435
rect 16600 -1470 16605 -1440
rect 16635 -1470 16715 -1440
rect 16745 -1470 16825 -1440
rect 16855 -1470 16885 -1440
rect 16915 -1470 17030 -1440
rect 17060 -1470 17140 -1440
rect 17170 -1470 17250 -1440
rect 17280 -1470 17360 -1440
rect 17390 -1470 17470 -1440
rect 17500 -1470 17620 -1440
rect 17650 -1470 17730 -1440
rect 17760 -1470 17840 -1440
rect 17870 -1470 17950 -1440
rect 17980 -1470 18010 -1440
rect 18040 -1470 18155 -1440
rect 18185 -1470 18265 -1440
rect 18295 -1470 18375 -1440
rect 18405 -1470 18485 -1440
rect 18515 -1470 18595 -1440
rect 18625 -1470 18630 -1440
rect 16600 -1480 18630 -1470
rect 16600 -1510 16605 -1480
rect 16635 -1510 16715 -1480
rect 16745 -1510 16825 -1480
rect 16855 -1510 16885 -1480
rect 16915 -1510 17030 -1480
rect 17060 -1510 17140 -1480
rect 17170 -1510 17250 -1480
rect 17280 -1510 17360 -1480
rect 17390 -1510 17470 -1480
rect 17500 -1510 17620 -1480
rect 17650 -1510 17730 -1480
rect 17760 -1510 17840 -1480
rect 17870 -1510 17950 -1480
rect 17980 -1510 18010 -1480
rect 18040 -1510 18155 -1480
rect 18185 -1510 18265 -1480
rect 18295 -1510 18375 -1480
rect 18405 -1510 18485 -1480
rect 18515 -1510 18595 -1480
rect 18625 -1510 18630 -1480
rect 16600 -1520 18630 -1510
rect 16600 -1550 16605 -1520
rect 16635 -1550 16715 -1520
rect 16745 -1550 16825 -1520
rect 16855 -1550 16885 -1520
rect 16915 -1550 17030 -1520
rect 17060 -1550 17140 -1520
rect 17170 -1550 17250 -1520
rect 17280 -1550 17360 -1520
rect 17390 -1550 17470 -1520
rect 17500 -1550 17620 -1520
rect 17650 -1550 17730 -1520
rect 17760 -1550 17840 -1520
rect 17870 -1550 17950 -1520
rect 17980 -1550 18010 -1520
rect 18040 -1550 18155 -1520
rect 18185 -1550 18265 -1520
rect 18295 -1550 18375 -1520
rect 18405 -1550 18485 -1520
rect 18515 -1550 18595 -1520
rect 18625 -1550 18630 -1520
rect 16600 -1555 18630 -1550
rect 17190 -1690 17450 -1685
rect 17190 -1720 17195 -1690
rect 17225 -1720 17415 -1690
rect 17445 -1720 17450 -1690
rect 17190 -1725 17450 -1720
rect 17670 -1690 17710 -1685
rect 17670 -1720 17675 -1690
rect 17705 -1695 17710 -1690
rect 17780 -1690 17820 -1685
rect 17780 -1695 17785 -1690
rect 17705 -1715 17785 -1695
rect 17705 -1720 17710 -1715
rect 17670 -1725 17710 -1720
rect 17780 -1720 17785 -1715
rect 17815 -1695 17820 -1690
rect 17890 -1690 17930 -1685
rect 17890 -1695 17895 -1690
rect 17815 -1715 17895 -1695
rect 17815 -1720 17820 -1715
rect 17780 -1725 17820 -1720
rect 17890 -1720 17895 -1715
rect 17925 -1720 17930 -1690
rect 17890 -1725 17930 -1720
rect 18205 -1690 18465 -1685
rect 18205 -1720 18210 -1690
rect 18240 -1720 18430 -1690
rect 18460 -1720 18465 -1690
rect 18205 -1725 18465 -1720
rect 16030 -1745 16070 -1740
rect 16030 -1775 16035 -1745
rect 16065 -1750 16070 -1745
rect 17080 -1745 17120 -1740
rect 17080 -1750 17085 -1745
rect 16065 -1770 17085 -1750
rect 16065 -1775 16070 -1770
rect 16030 -1780 16070 -1775
rect 17080 -1775 17085 -1770
rect 17115 -1750 17120 -1745
rect 17300 -1745 17340 -1740
rect 17300 -1750 17305 -1745
rect 17115 -1770 17305 -1750
rect 17115 -1775 17120 -1770
rect 17080 -1780 17120 -1775
rect 17300 -1775 17305 -1770
rect 17335 -1750 17340 -1745
rect 18315 -1745 18355 -1740
rect 18315 -1750 18320 -1745
rect 17335 -1770 18320 -1750
rect 17335 -1775 17340 -1770
rect 17300 -1780 17340 -1775
rect 18315 -1775 18320 -1770
rect 18350 -1750 18355 -1745
rect 18535 -1745 18575 -1740
rect 18535 -1750 18540 -1745
rect 18350 -1770 18540 -1750
rect 18350 -1775 18355 -1770
rect 18315 -1780 18355 -1775
rect 18535 -1775 18540 -1770
rect 18570 -1775 18575 -1745
rect 18535 -1780 18575 -1775
rect 18885 -1750 19130 -1745
rect 18885 -1780 18890 -1750
rect 18920 -1780 19095 -1750
rect 19125 -1780 19130 -1750
rect 18885 -1785 19130 -1780
rect 15785 -1800 17230 -1795
rect 15785 -1830 15790 -1800
rect 15820 -1830 17195 -1800
rect 17225 -1830 17230 -1800
rect 15785 -1835 17230 -1830
rect 18425 -1800 18465 -1795
rect 18425 -1830 18430 -1800
rect 18460 -1805 18465 -1800
rect 19775 -1800 19815 -1795
rect 19775 -1805 19780 -1800
rect 18460 -1825 19780 -1805
rect 18460 -1830 18465 -1825
rect 18425 -1835 18465 -1830
rect 19775 -1830 19780 -1825
rect 19810 -1830 19815 -1800
rect 19775 -1835 19815 -1830
rect 16105 -1855 16145 -1850
rect 16105 -1885 16110 -1855
rect 16140 -1860 16145 -1855
rect 16765 -1855 16805 -1850
rect 16765 -1860 16770 -1855
rect 16140 -1880 16770 -1860
rect 16140 -1885 16145 -1880
rect 16105 -1890 16145 -1885
rect 16765 -1885 16770 -1880
rect 16800 -1885 16805 -1855
rect 16765 -1890 16805 -1885
rect 17780 -1890 17820 -1885
rect 17780 -1920 17785 -1890
rect 17815 -1895 17820 -1890
rect 19535 -1890 19575 -1885
rect 19535 -1895 19540 -1890
rect 17815 -1915 19540 -1895
rect 17815 -1920 17820 -1915
rect 17780 -1925 17820 -1920
rect 19535 -1920 19540 -1915
rect 19570 -1920 19575 -1890
rect 19535 -1925 19575 -1920
rect 16155 -1945 19365 -1940
rect 16155 -1975 16160 -1945
rect 16190 -1975 19330 -1945
rect 19360 -1975 19365 -1945
rect 16155 -1980 19365 -1975
rect 16315 -2000 16355 -1995
rect 16315 -2030 16320 -2000
rect 16350 -2005 16355 -2000
rect 17425 -2005 17430 -2000
rect 16350 -2025 17430 -2005
rect 16350 -2030 16355 -2025
rect 16315 -2035 16355 -2030
rect 17425 -2035 17430 -2025
rect 17465 -2035 17470 -2000
rect 18124 -2035 18129 -2000
rect 18164 -2005 18870 -2000
rect 18164 -2035 18835 -2005
rect 18865 -2035 18870 -2005
rect 18165 -2040 18870 -2035
rect 17425 -2060 19120 -2055
rect 17425 -2090 17430 -2060
rect 17460 -2090 19085 -2060
rect 19115 -2090 19120 -2060
rect 17425 -2095 19120 -2090
rect 16260 -2100 16300 -2095
rect 16260 -2130 16265 -2100
rect 16295 -2105 16300 -2100
rect 16480 -2100 16520 -2095
rect 16480 -2105 16485 -2100
rect 16295 -2125 16485 -2105
rect 16295 -2130 16300 -2125
rect 16260 -2135 16300 -2130
rect 16480 -2130 16485 -2125
rect 16515 -2105 16520 -2100
rect 16730 -2100 16770 -2095
rect 16730 -2105 16735 -2100
rect 16515 -2125 16735 -2105
rect 16515 -2130 16520 -2125
rect 16480 -2135 16520 -2130
rect 16730 -2130 16735 -2125
rect 16765 -2130 16770 -2100
rect 16730 -2135 16770 -2130
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19405 -2997 19440 -2992
rect 16160 -3025 16195 -3020
rect 19405 -3037 19440 -3032
rect 16160 -3065 16195 -3060
rect 16730 -3105 17820 -3100
rect 15820 -3115 15985 -3110
rect 15820 -3145 15825 -3115
rect 15855 -3116 15985 -3115
rect 15855 -3145 15950 -3116
rect 15820 -3150 15950 -3145
rect 16730 -3135 16735 -3105
rect 16765 -3135 17785 -3105
rect 17815 -3135 17820 -3105
rect 16730 -3140 17820 -3135
rect 18615 -3105 18870 -3100
rect 18615 -3135 18620 -3105
rect 18650 -3135 18835 -3105
rect 18865 -3135 18870 -3105
rect 18615 -3140 18870 -3135
rect 19610 -3115 19645 -3110
rect 15950 -3156 15985 -3151
rect 19610 -3160 19645 -3150
rect 15950 -3789 15985 -3784
rect 15950 -3829 15985 -3824
rect 19610 -3789 19645 -3784
rect 19610 -3829 19645 -3824
rect 15960 -3830 15980 -3829
rect 19620 -3830 19640 -3829
rect 16280 -3894 16315 -3889
rect 16280 -3934 16315 -3929
rect 19285 -3894 19320 -3889
rect 19285 -3934 19320 -3929
rect 16290 -3935 16310 -3934
rect 19290 -3935 19310 -3934
rect 16605 -3969 16640 -3964
rect 16605 -4009 16640 -4004
rect 18960 -3969 18995 -3964
rect 18960 -4009 18995 -4004
rect 16615 -4010 16635 -4009
rect 18965 -4010 18985 -4009
rect 15640 -4110 16645 -4105
rect 15640 -4140 16285 -4110
rect 16315 -4140 16610 -4110
rect 16640 -4140 16645 -4110
rect 15640 -4150 16645 -4140
rect 15640 -4180 16285 -4150
rect 16315 -4180 16610 -4150
rect 16640 -4180 16645 -4150
rect 15640 -4190 16645 -4180
rect 15640 -4220 16285 -4190
rect 16315 -4220 16610 -4190
rect 16640 -4220 16645 -4190
rect 15640 -4225 16645 -4220
rect 17780 -4205 19320 -4200
rect 17780 -4235 17785 -4205
rect 17815 -4235 18960 -4205
rect 18990 -4235 19285 -4205
rect 19315 -4235 19320 -4205
rect 17780 -4245 19320 -4235
rect 17250 -4250 17300 -4245
rect 15820 -4255 17300 -4250
rect 15820 -4285 15825 -4255
rect 15855 -4285 17260 -4255
rect 17290 -4285 17300 -4255
rect 15820 -4290 17300 -4285
rect 17250 -4295 17300 -4290
rect 17780 -4275 17785 -4245
rect 17815 -4275 18960 -4245
rect 18990 -4275 19285 -4245
rect 19315 -4275 19320 -4245
rect 17780 -4285 19320 -4275
rect 17780 -4315 17785 -4285
rect 17815 -4315 18960 -4285
rect 18990 -4315 19285 -4285
rect 19315 -4315 19320 -4285
rect 17780 -4320 19320 -4315
rect 16900 -4335 16950 -4325
rect 16900 -4340 16910 -4335
rect 15645 -4345 16910 -4340
rect 15645 -4375 15650 -4345
rect 15680 -4375 15690 -4345
rect 15720 -4375 15730 -4345
rect 15760 -4365 16910 -4345
rect 16940 -4365 16950 -4335
rect 15760 -4375 16950 -4365
rect 15645 -4385 16950 -4375
rect 15645 -4415 15650 -4385
rect 15680 -4415 15690 -4385
rect 15720 -4415 15730 -4385
rect 15760 -4415 16910 -4385
rect 16940 -4415 16950 -4385
rect 15645 -4425 16950 -4415
rect 15645 -4455 15650 -4425
rect 15680 -4455 15690 -4425
rect 15720 -4455 15730 -4425
rect 15760 -4435 16950 -4425
rect 15760 -4455 16910 -4435
rect 15645 -4460 16910 -4455
rect 16900 -4465 16910 -4460
rect 16940 -4465 16950 -4435
rect 16900 -4475 16950 -4465
rect 18650 -4465 18700 -4460
rect 18650 -4470 18925 -4465
rect 15950 -4480 15990 -4475
rect 15950 -4510 15955 -4480
rect 15985 -4485 15990 -4480
rect 16205 -4480 16245 -4475
rect 16205 -4485 16210 -4480
rect 15985 -4505 16210 -4485
rect 15985 -4510 15990 -4505
rect 15950 -4515 15990 -4510
rect 16205 -4510 16210 -4505
rect 16240 -4510 16245 -4480
rect 18650 -4500 18660 -4470
rect 18690 -4500 18890 -4470
rect 18920 -4500 18925 -4470
rect 18650 -4505 18925 -4500
rect 19355 -4470 19395 -4465
rect 19355 -4500 19360 -4470
rect 19390 -4475 19395 -4470
rect 19610 -4470 19650 -4465
rect 19610 -4475 19615 -4470
rect 19390 -4495 19615 -4475
rect 19390 -4500 19395 -4495
rect 19355 -4505 19395 -4500
rect 19610 -4500 19615 -4495
rect 19645 -4500 19650 -4470
rect 19610 -4505 19650 -4500
rect 18650 -4510 18700 -4505
rect 16205 -4515 16245 -4510
rect 17955 -4520 17995 -4515
rect 17955 -4550 17960 -4520
rect 17990 -4525 17995 -4520
rect 17990 -4545 19905 -4525
rect 17990 -4550 17995 -4545
rect 17955 -4555 17995 -4550
<< via2 >>
rect 17260 -4285 17290 -4255
rect 16910 -4365 16940 -4335
rect 16910 -4415 16940 -4385
rect 16910 -4465 16940 -4435
rect 16210 -4510 16240 -4480
rect 18660 -4500 18690 -4470
rect 19360 -4500 19390 -4470
rect 17960 -4550 17990 -4520
<< metal3 >>
rect 17250 -4250 17300 -4245
rect 17250 -4290 17255 -4250
rect 17295 -4290 17300 -4250
rect 17250 -4295 17300 -4290
rect 16900 -4330 16950 -4325
rect 16900 -4370 16905 -4330
rect 16945 -4370 16950 -4330
rect 16900 -4380 16950 -4370
rect 16900 -4420 16905 -4380
rect 16945 -4420 16950 -4380
rect 16900 -4430 16950 -4420
rect 16900 -4470 16905 -4430
rect 16945 -4470 16950 -4430
rect 16900 -4475 16950 -4470
rect 18650 -4465 18700 -4460
rect 16205 -4480 16245 -4475
rect 16205 -4510 16210 -4480
rect 16240 -4510 16245 -4480
rect 18650 -4505 18655 -4465
rect 18695 -4505 18700 -4465
rect 18650 -4510 18700 -4505
rect 19355 -4470 19395 -4465
rect 19355 -4500 19360 -4470
rect 19390 -4500 19395 -4470
rect 16205 -4630 16245 -4510
rect 17955 -4520 17995 -4515
rect 17955 -4550 17960 -4520
rect 17990 -4550 17995 -4520
rect 17955 -4630 17995 -4550
rect 19355 -4630 19395 -4500
rect 15760 -4725 15990 -4630
rect 16110 -4725 16340 -4630
rect 16460 -4725 16690 -4630
rect 16810 -4725 17040 -4630
rect 15760 -4775 17040 -4725
rect 15760 -4860 15990 -4775
rect 16110 -4860 16340 -4775
rect 16460 -4860 16690 -4775
rect 16810 -4860 17040 -4775
rect 17160 -4725 17390 -4630
rect 17510 -4725 17740 -4630
rect 17860 -4725 18090 -4630
rect 18210 -4725 18440 -4630
rect 17160 -4775 18440 -4725
rect 17160 -4860 17390 -4775
rect 17510 -4860 17740 -4775
rect 17860 -4860 18090 -4775
rect 18210 -4860 18440 -4775
rect 18560 -4725 18790 -4630
rect 18910 -4725 19140 -4630
rect 19260 -4725 19490 -4630
rect 19610 -4725 19840 -4630
rect 18560 -4775 19840 -4725
rect 18560 -4860 18790 -4775
rect 18910 -4860 19140 -4775
rect 19260 -4860 19490 -4775
rect 19610 -4860 19840 -4775
rect 16200 -4980 16250 -4860
rect 17950 -4980 18000 -4860
rect 19350 -4980 19400 -4860
rect 15760 -5075 15990 -4980
rect 16110 -5075 16340 -4980
rect 16460 -5075 16690 -4980
rect 16810 -5075 17040 -4980
rect 15760 -5125 17040 -5075
rect 15760 -5210 15990 -5125
rect 16110 -5210 16340 -5125
rect 16460 -5210 16690 -5125
rect 16810 -5210 17040 -5125
rect 17160 -5075 17390 -4980
rect 17510 -5075 17740 -4980
rect 17860 -5075 18090 -4980
rect 18210 -5075 18440 -4980
rect 17160 -5125 18440 -5075
rect 17160 -5210 17390 -5125
rect 17510 -5210 17740 -5125
rect 17860 -5210 18090 -5125
rect 18210 -5210 18440 -5125
rect 18560 -5075 18790 -4980
rect 18910 -5075 19140 -4980
rect 19260 -5075 19490 -4980
rect 19610 -5075 19840 -4980
rect 18560 -5125 19840 -5075
rect 18560 -5210 18790 -5125
rect 18910 -5210 19140 -5125
rect 19260 -5210 19490 -5125
rect 19610 -5210 19840 -5125
rect 16200 -5330 16250 -5210
rect 17950 -5330 18000 -5210
rect 19350 -5330 19400 -5210
rect 15760 -5425 15990 -5330
rect 16110 -5425 16340 -5330
rect 16460 -5425 16690 -5330
rect 16810 -5425 17040 -5330
rect 15760 -5475 17040 -5425
rect 15760 -5560 15990 -5475
rect 16110 -5560 16340 -5475
rect 16460 -5560 16690 -5475
rect 16810 -5560 17040 -5475
rect 17160 -5425 17390 -5330
rect 17510 -5425 17740 -5330
rect 17860 -5425 18090 -5330
rect 18210 -5425 18440 -5330
rect 17160 -5475 18440 -5425
rect 17160 -5560 17390 -5475
rect 17510 -5560 17740 -5475
rect 17860 -5560 18090 -5475
rect 18210 -5560 18440 -5475
rect 18560 -5425 18790 -5330
rect 18910 -5425 19140 -5330
rect 19260 -5425 19490 -5330
rect 19610 -5425 19840 -5330
rect 18560 -5475 19840 -5425
rect 18560 -5560 18790 -5475
rect 18910 -5560 19140 -5475
rect 19260 -5560 19490 -5475
rect 19610 -5560 19840 -5475
rect 16200 -5680 16250 -5560
rect 17950 -5680 18000 -5560
rect 19350 -5680 19400 -5560
rect 15760 -5775 15990 -5680
rect 16110 -5775 16340 -5680
rect 16460 -5775 16690 -5680
rect 16810 -5775 17040 -5680
rect 15760 -5825 17040 -5775
rect 15760 -5910 15990 -5825
rect 16110 -5910 16340 -5825
rect 16460 -5910 16690 -5825
rect 16810 -5910 17040 -5825
rect 17160 -5775 17390 -5680
rect 17510 -5775 17740 -5680
rect 17860 -5775 18090 -5680
rect 18210 -5775 18440 -5680
rect 17160 -5825 18440 -5775
rect 17160 -5910 17390 -5825
rect 17510 -5910 17740 -5825
rect 17860 -5910 18090 -5825
rect 18210 -5910 18440 -5825
rect 18560 -5775 18790 -5680
rect 18910 -5775 19140 -5680
rect 19260 -5775 19490 -5680
rect 19610 -5775 19840 -5680
rect 18560 -5825 19840 -5775
rect 18560 -5910 18790 -5825
rect 18910 -5910 19140 -5825
rect 19260 -5910 19490 -5825
rect 19610 -5910 19840 -5825
rect 16200 -6030 16250 -5910
rect 17950 -6030 18000 -5910
rect 19350 -6030 19400 -5910
rect 15760 -6125 15990 -6030
rect 16110 -6125 16340 -6030
rect 16460 -6125 16690 -6030
rect 16810 -6125 17040 -6030
rect 15760 -6175 17040 -6125
rect 15760 -6260 15990 -6175
rect 16110 -6260 16340 -6175
rect 16460 -6260 16690 -6175
rect 16810 -6260 17040 -6175
rect 17160 -6125 17390 -6030
rect 17510 -6125 17740 -6030
rect 17860 -6125 18090 -6030
rect 18210 -6125 18440 -6030
rect 17160 -6175 18440 -6125
rect 17160 -6260 17390 -6175
rect 17510 -6260 17740 -6175
rect 17860 -6260 18090 -6175
rect 18210 -6260 18440 -6175
rect 18560 -6125 18790 -6030
rect 18910 -6125 19140 -6030
rect 19260 -6125 19490 -6030
rect 19610 -6125 19840 -6030
rect 18560 -6175 19840 -6125
rect 18560 -6260 18790 -6175
rect 18910 -6260 19140 -6175
rect 19260 -6260 19490 -6175
rect 19610 -6260 19840 -6175
<< via3 >>
rect 17255 -4255 17295 -4250
rect 17255 -4285 17260 -4255
rect 17260 -4285 17290 -4255
rect 17290 -4285 17295 -4255
rect 17255 -4290 17295 -4285
rect 16905 -4335 16945 -4330
rect 16905 -4365 16910 -4335
rect 16910 -4365 16940 -4335
rect 16940 -4365 16945 -4335
rect 16905 -4370 16945 -4365
rect 16905 -4385 16945 -4380
rect 16905 -4415 16910 -4385
rect 16910 -4415 16940 -4385
rect 16940 -4415 16945 -4385
rect 16905 -4420 16945 -4415
rect 16905 -4435 16945 -4430
rect 16905 -4465 16910 -4435
rect 16910 -4465 16940 -4435
rect 16940 -4465 16945 -4435
rect 16905 -4470 16945 -4465
rect 18655 -4470 18695 -4465
rect 18655 -4500 18660 -4470
rect 18660 -4500 18690 -4470
rect 18690 -4500 18695 -4470
rect 18655 -4505 18695 -4500
<< mimcap >>
rect 15775 -4730 15975 -4645
rect 15775 -4770 15855 -4730
rect 15895 -4770 15975 -4730
rect 15775 -4845 15975 -4770
rect 16125 -4730 16325 -4645
rect 16125 -4770 16205 -4730
rect 16245 -4770 16325 -4730
rect 16125 -4845 16325 -4770
rect 16475 -4730 16675 -4645
rect 16475 -4770 16555 -4730
rect 16595 -4770 16675 -4730
rect 16475 -4845 16675 -4770
rect 16825 -4730 17025 -4645
rect 16825 -4770 16905 -4730
rect 16945 -4770 17025 -4730
rect 16825 -4845 17025 -4770
rect 17175 -4730 17375 -4645
rect 17175 -4770 17255 -4730
rect 17295 -4770 17375 -4730
rect 17175 -4845 17375 -4770
rect 17525 -4730 17725 -4645
rect 17525 -4770 17605 -4730
rect 17645 -4770 17725 -4730
rect 17525 -4845 17725 -4770
rect 17875 -4730 18075 -4645
rect 17875 -4770 17955 -4730
rect 17995 -4770 18075 -4730
rect 17875 -4845 18075 -4770
rect 18225 -4730 18425 -4645
rect 18225 -4770 18305 -4730
rect 18345 -4770 18425 -4730
rect 18225 -4845 18425 -4770
rect 18575 -4730 18775 -4645
rect 18575 -4770 18655 -4730
rect 18695 -4770 18775 -4730
rect 18575 -4845 18775 -4770
rect 18925 -4730 19125 -4645
rect 18925 -4770 19005 -4730
rect 19045 -4770 19125 -4730
rect 18925 -4845 19125 -4770
rect 19275 -4730 19475 -4645
rect 19275 -4770 19355 -4730
rect 19395 -4770 19475 -4730
rect 19275 -4845 19475 -4770
rect 19625 -4730 19825 -4645
rect 19625 -4770 19705 -4730
rect 19745 -4770 19825 -4730
rect 19625 -4845 19825 -4770
rect 15775 -5080 15975 -4995
rect 15775 -5120 15855 -5080
rect 15895 -5120 15975 -5080
rect 15775 -5195 15975 -5120
rect 16125 -5080 16325 -4995
rect 16125 -5120 16205 -5080
rect 16245 -5120 16325 -5080
rect 16125 -5195 16325 -5120
rect 16475 -5080 16675 -4995
rect 16475 -5120 16555 -5080
rect 16595 -5120 16675 -5080
rect 16475 -5195 16675 -5120
rect 16825 -5080 17025 -4995
rect 16825 -5120 16905 -5080
rect 16945 -5120 17025 -5080
rect 16825 -5195 17025 -5120
rect 17175 -5080 17375 -4995
rect 17175 -5120 17255 -5080
rect 17295 -5120 17375 -5080
rect 17175 -5195 17375 -5120
rect 17525 -5080 17725 -4995
rect 17525 -5120 17605 -5080
rect 17645 -5120 17725 -5080
rect 17525 -5195 17725 -5120
rect 17875 -5080 18075 -4995
rect 17875 -5120 17955 -5080
rect 17995 -5120 18075 -5080
rect 17875 -5195 18075 -5120
rect 18225 -5080 18425 -4995
rect 18225 -5120 18305 -5080
rect 18345 -5120 18425 -5080
rect 18225 -5195 18425 -5120
rect 18575 -5080 18775 -4995
rect 18575 -5120 18655 -5080
rect 18695 -5120 18775 -5080
rect 18575 -5195 18775 -5120
rect 18925 -5080 19125 -4995
rect 18925 -5120 19005 -5080
rect 19045 -5120 19125 -5080
rect 18925 -5195 19125 -5120
rect 19275 -5080 19475 -4995
rect 19275 -5120 19355 -5080
rect 19395 -5120 19475 -5080
rect 19275 -5195 19475 -5120
rect 19625 -5080 19825 -4995
rect 19625 -5120 19705 -5080
rect 19745 -5120 19825 -5080
rect 19625 -5195 19825 -5120
rect 15775 -5430 15975 -5345
rect 15775 -5470 15855 -5430
rect 15895 -5470 15975 -5430
rect 15775 -5545 15975 -5470
rect 16125 -5430 16325 -5345
rect 16125 -5470 16205 -5430
rect 16245 -5470 16325 -5430
rect 16125 -5545 16325 -5470
rect 16475 -5430 16675 -5345
rect 16475 -5470 16555 -5430
rect 16595 -5470 16675 -5430
rect 16475 -5545 16675 -5470
rect 16825 -5430 17025 -5345
rect 16825 -5470 16905 -5430
rect 16945 -5470 17025 -5430
rect 16825 -5545 17025 -5470
rect 17175 -5430 17375 -5345
rect 17175 -5470 17255 -5430
rect 17295 -5470 17375 -5430
rect 17175 -5545 17375 -5470
rect 17525 -5430 17725 -5345
rect 17525 -5470 17605 -5430
rect 17645 -5470 17725 -5430
rect 17525 -5545 17725 -5470
rect 17875 -5430 18075 -5345
rect 17875 -5470 17955 -5430
rect 17995 -5470 18075 -5430
rect 17875 -5545 18075 -5470
rect 18225 -5430 18425 -5345
rect 18225 -5470 18305 -5430
rect 18345 -5470 18425 -5430
rect 18225 -5545 18425 -5470
rect 18575 -5430 18775 -5345
rect 18575 -5470 18655 -5430
rect 18695 -5470 18775 -5430
rect 18575 -5545 18775 -5470
rect 18925 -5430 19125 -5345
rect 18925 -5470 19005 -5430
rect 19045 -5470 19125 -5430
rect 18925 -5545 19125 -5470
rect 19275 -5430 19475 -5345
rect 19275 -5470 19355 -5430
rect 19395 -5470 19475 -5430
rect 19275 -5545 19475 -5470
rect 19625 -5430 19825 -5345
rect 19625 -5470 19705 -5430
rect 19745 -5470 19825 -5430
rect 19625 -5545 19825 -5470
rect 15775 -5780 15975 -5695
rect 15775 -5820 15855 -5780
rect 15895 -5820 15975 -5780
rect 15775 -5895 15975 -5820
rect 16125 -5780 16325 -5695
rect 16125 -5820 16205 -5780
rect 16245 -5820 16325 -5780
rect 16125 -5895 16325 -5820
rect 16475 -5780 16675 -5695
rect 16475 -5820 16555 -5780
rect 16595 -5820 16675 -5780
rect 16475 -5895 16675 -5820
rect 16825 -5780 17025 -5695
rect 16825 -5820 16905 -5780
rect 16945 -5820 17025 -5780
rect 16825 -5895 17025 -5820
rect 17175 -5780 17375 -5695
rect 17175 -5820 17255 -5780
rect 17295 -5820 17375 -5780
rect 17175 -5895 17375 -5820
rect 17525 -5780 17725 -5695
rect 17525 -5820 17605 -5780
rect 17645 -5820 17725 -5780
rect 17525 -5895 17725 -5820
rect 17875 -5780 18075 -5695
rect 17875 -5820 17955 -5780
rect 17995 -5820 18075 -5780
rect 17875 -5895 18075 -5820
rect 18225 -5780 18425 -5695
rect 18225 -5820 18305 -5780
rect 18345 -5820 18425 -5780
rect 18225 -5895 18425 -5820
rect 18575 -5780 18775 -5695
rect 18575 -5820 18655 -5780
rect 18695 -5820 18775 -5780
rect 18575 -5895 18775 -5820
rect 18925 -5780 19125 -5695
rect 18925 -5820 19005 -5780
rect 19045 -5820 19125 -5780
rect 18925 -5895 19125 -5820
rect 19275 -5780 19475 -5695
rect 19275 -5820 19355 -5780
rect 19395 -5820 19475 -5780
rect 19275 -5895 19475 -5820
rect 19625 -5780 19825 -5695
rect 19625 -5820 19705 -5780
rect 19745 -5820 19825 -5780
rect 19625 -5895 19825 -5820
rect 15775 -6130 15975 -6045
rect 15775 -6170 15855 -6130
rect 15895 -6170 15975 -6130
rect 15775 -6245 15975 -6170
rect 16125 -6130 16325 -6045
rect 16125 -6170 16205 -6130
rect 16245 -6170 16325 -6130
rect 16125 -6245 16325 -6170
rect 16475 -6130 16675 -6045
rect 16475 -6170 16555 -6130
rect 16595 -6170 16675 -6130
rect 16475 -6245 16675 -6170
rect 16825 -6130 17025 -6045
rect 16825 -6170 16905 -6130
rect 16945 -6170 17025 -6130
rect 16825 -6245 17025 -6170
rect 17175 -6130 17375 -6045
rect 17175 -6170 17255 -6130
rect 17295 -6170 17375 -6130
rect 17175 -6245 17375 -6170
rect 17525 -6130 17725 -6045
rect 17525 -6170 17605 -6130
rect 17645 -6170 17725 -6130
rect 17525 -6245 17725 -6170
rect 17875 -6130 18075 -6045
rect 17875 -6170 17955 -6130
rect 17995 -6170 18075 -6130
rect 17875 -6245 18075 -6170
rect 18225 -6130 18425 -6045
rect 18225 -6170 18305 -6130
rect 18345 -6170 18425 -6130
rect 18225 -6245 18425 -6170
rect 18575 -6130 18775 -6045
rect 18575 -6170 18655 -6130
rect 18695 -6170 18775 -6130
rect 18575 -6245 18775 -6170
rect 18925 -6130 19125 -6045
rect 18925 -6170 19005 -6130
rect 19045 -6170 19125 -6130
rect 18925 -6245 19125 -6170
rect 19275 -6130 19475 -6045
rect 19275 -6170 19355 -6130
rect 19395 -6170 19475 -6130
rect 19275 -6245 19475 -6170
rect 19625 -6130 19825 -6045
rect 19625 -6170 19705 -6130
rect 19745 -6170 19825 -6130
rect 19625 -6245 19825 -6170
<< mimcapcontact >>
rect 15855 -4770 15895 -4730
rect 16205 -4770 16245 -4730
rect 16555 -4770 16595 -4730
rect 16905 -4770 16945 -4730
rect 17255 -4770 17295 -4730
rect 17605 -4770 17645 -4730
rect 17955 -4770 17995 -4730
rect 18305 -4770 18345 -4730
rect 18655 -4770 18695 -4730
rect 19005 -4770 19045 -4730
rect 19355 -4770 19395 -4730
rect 19705 -4770 19745 -4730
rect 15855 -5120 15895 -5080
rect 16205 -5120 16245 -5080
rect 16555 -5120 16595 -5080
rect 16905 -5120 16945 -5080
rect 17255 -5120 17295 -5080
rect 17605 -5120 17645 -5080
rect 17955 -5120 17995 -5080
rect 18305 -5120 18345 -5080
rect 18655 -5120 18695 -5080
rect 19005 -5120 19045 -5080
rect 19355 -5120 19395 -5080
rect 19705 -5120 19745 -5080
rect 15855 -5470 15895 -5430
rect 16205 -5470 16245 -5430
rect 16555 -5470 16595 -5430
rect 16905 -5470 16945 -5430
rect 17255 -5470 17295 -5430
rect 17605 -5470 17645 -5430
rect 17955 -5470 17995 -5430
rect 18305 -5470 18345 -5430
rect 18655 -5470 18695 -5430
rect 19005 -5470 19045 -5430
rect 19355 -5470 19395 -5430
rect 19705 -5470 19745 -5430
rect 15855 -5820 15895 -5780
rect 16205 -5820 16245 -5780
rect 16555 -5820 16595 -5780
rect 16905 -5820 16945 -5780
rect 17255 -5820 17295 -5780
rect 17605 -5820 17645 -5780
rect 17955 -5820 17995 -5780
rect 18305 -5820 18345 -5780
rect 18655 -5820 18695 -5780
rect 19005 -5820 19045 -5780
rect 19355 -5820 19395 -5780
rect 19705 -5820 19745 -5780
rect 15855 -6170 15895 -6130
rect 16205 -6170 16245 -6130
rect 16555 -6170 16595 -6130
rect 16905 -6170 16945 -6130
rect 17255 -6170 17295 -6130
rect 17605 -6170 17645 -6130
rect 17955 -6170 17995 -6130
rect 18305 -6170 18345 -6130
rect 18655 -6170 18695 -6130
rect 19005 -6170 19045 -6130
rect 19355 -6170 19395 -6130
rect 19705 -6170 19745 -6130
<< metal4 >>
rect 17250 -4250 17300 -4245
rect 17250 -4290 17255 -4250
rect 17295 -4290 17300 -4250
rect 16900 -4330 16950 -4325
rect 16900 -4370 16905 -4330
rect 16945 -4370 16950 -4330
rect 16900 -4380 16950 -4370
rect 16900 -4420 16905 -4380
rect 16945 -4420 16950 -4380
rect 16900 -4430 16950 -4420
rect 16900 -4470 16905 -4430
rect 16945 -4470 16950 -4430
rect 16900 -4725 16950 -4470
rect 15850 -4730 16950 -4725
rect 15850 -4770 15855 -4730
rect 15895 -4770 16205 -4730
rect 16245 -4770 16555 -4730
rect 16595 -4770 16905 -4730
rect 16945 -4770 16950 -4730
rect 15850 -4775 16950 -4770
rect 17250 -4725 17300 -4290
rect 18650 -4465 18700 -4460
rect 18650 -4505 18655 -4465
rect 18695 -4505 18700 -4465
rect 18650 -4725 18700 -4505
rect 17250 -4730 18350 -4725
rect 17250 -4770 17255 -4730
rect 17295 -4770 17605 -4730
rect 17645 -4770 17955 -4730
rect 17995 -4770 18305 -4730
rect 18345 -4770 18350 -4730
rect 17250 -4775 18350 -4770
rect 18650 -4730 19750 -4725
rect 18650 -4770 18655 -4730
rect 18695 -4770 19005 -4730
rect 19045 -4770 19355 -4730
rect 19395 -4770 19705 -4730
rect 19745 -4770 19750 -4730
rect 18650 -4775 19750 -4770
rect 16200 -5075 16250 -4775
rect 17950 -5075 18000 -4775
rect 19350 -5075 19400 -4775
rect 15850 -5080 16950 -5075
rect 15850 -5120 15855 -5080
rect 15895 -5120 16205 -5080
rect 16245 -5120 16555 -5080
rect 16595 -5120 16905 -5080
rect 16945 -5120 16950 -5080
rect 15850 -5125 16950 -5120
rect 17250 -5080 18350 -5075
rect 17250 -5120 17255 -5080
rect 17295 -5120 17605 -5080
rect 17645 -5120 17955 -5080
rect 17995 -5120 18305 -5080
rect 18345 -5120 18350 -5080
rect 17250 -5125 18350 -5120
rect 18650 -5080 19750 -5075
rect 18650 -5120 18655 -5080
rect 18695 -5120 19005 -5080
rect 19045 -5120 19355 -5080
rect 19395 -5120 19705 -5080
rect 19745 -5120 19750 -5080
rect 18650 -5125 19750 -5120
rect 16200 -5425 16250 -5125
rect 17950 -5425 18000 -5125
rect 19350 -5425 19400 -5125
rect 15850 -5430 16950 -5425
rect 15850 -5470 15855 -5430
rect 15895 -5470 16205 -5430
rect 16245 -5470 16555 -5430
rect 16595 -5470 16905 -5430
rect 16945 -5470 16950 -5430
rect 15850 -5475 16950 -5470
rect 17250 -5430 18350 -5425
rect 17250 -5470 17255 -5430
rect 17295 -5470 17605 -5430
rect 17645 -5470 17955 -5430
rect 17995 -5470 18305 -5430
rect 18345 -5470 18350 -5430
rect 17250 -5475 18350 -5470
rect 18650 -5430 19750 -5425
rect 18650 -5470 18655 -5430
rect 18695 -5470 19005 -5430
rect 19045 -5470 19355 -5430
rect 19395 -5470 19705 -5430
rect 19745 -5470 19750 -5430
rect 18650 -5475 19750 -5470
rect 16200 -5775 16250 -5475
rect 17950 -5775 18000 -5475
rect 19350 -5775 19400 -5475
rect 15850 -5780 16950 -5775
rect 15850 -5820 15855 -5780
rect 15895 -5820 16205 -5780
rect 16245 -5820 16555 -5780
rect 16595 -5820 16905 -5780
rect 16945 -5820 16950 -5780
rect 15850 -5825 16950 -5820
rect 17250 -5780 18350 -5775
rect 17250 -5820 17255 -5780
rect 17295 -5820 17605 -5780
rect 17645 -5820 17955 -5780
rect 17995 -5820 18305 -5780
rect 18345 -5820 18350 -5780
rect 17250 -5825 18350 -5820
rect 18650 -5780 19750 -5775
rect 18650 -5820 18655 -5780
rect 18695 -5820 19005 -5780
rect 19045 -5820 19355 -5780
rect 19395 -5820 19705 -5780
rect 19745 -5820 19750 -5780
rect 18650 -5825 19750 -5820
rect 16200 -6125 16250 -5825
rect 17950 -6125 18000 -5825
rect 19350 -6125 19400 -5825
rect 15850 -6130 16950 -6125
rect 15850 -6170 15855 -6130
rect 15895 -6170 16205 -6130
rect 16245 -6170 16555 -6130
rect 16595 -6170 16905 -6130
rect 16945 -6170 16950 -6130
rect 15850 -6175 16950 -6170
rect 17250 -6130 18350 -6125
rect 17250 -6170 17255 -6130
rect 17295 -6170 17605 -6130
rect 17645 -6170 17955 -6130
rect 17995 -6170 18305 -6130
rect 18345 -6170 18350 -6130
rect 17250 -6175 18350 -6170
rect 18650 -6130 19750 -6125
rect 18650 -6170 18655 -6130
rect 18695 -6170 19005 -6130
rect 19045 -6170 19355 -6130
rect 19395 -6170 19705 -6130
rect 19745 -6170 19750 -6130
rect 18650 -6175 19750 -6170
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 18145 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_18
timestamp 1723858470
transform 1 0 16785 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_19
timestamp 1723858470
transform 1 0 17465 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_20
timestamp 1723858470
transform 1 0 18145 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_21
timestamp 1723858470
transform 1 0 18145 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_22
timestamp 1723858470
transform 1 0 17465 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23
timestamp 1723858470
transform 1 0 17465 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_24
timestamp 1723858470
transform 1 0 16785 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25
timestamp 1723858470
transform 1 0 16785 0 1 -3455
box 0 0 670 670
<< labels >>
flabel metal3 19355 -4485 19355 -4485 7 FreeSans 400 180 -40 0 cap_res2
flabel metal2 15995 -4505 15995 -4505 5 FreeSans 400 0 0 -40 cap_res1
flabel metal1 18780 -1215 18780 -1215 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal1 16235 -1015 16235 -1015 3 FreeSans 400 0 200 0 START_UP
flabel metal2 17060 -645 17060 -645 3 FreeSans 400 0 200 0 V_p_1
flabel metal1 15890 -1330 15890 -1330 7 FreeSans 400 0 -200 0 NFET_GATE_10uA
flabel metal2 18580 -645 18580 -645 3 FreeSans 400 180 200 0 V_p_2
flabel metal2 16670 -510 16670 -510 1 FreeSans 400 0 0 80 Vin+
flabel metal2 16665 -205 16665 -205 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 18930 -505 18930 -505 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal2 18030 -60 18030 -60 7 FreeSans 240 0 -120 0 1st_Vout_2
flabel metal2 16620 -20 16620 -20 5 FreeSans 400 0 0 -40 V_mir1
flabel metal2 17570 -60 17570 -60 3 FreeSans 240 0 120 0 1st_Vout_1
flabel via1 17800 1455 17800 1455 1 FreeSans 400 0 0 200 PFET_GATE_10uA
flabel metal1 19795 1640 19795 1640 1 FreeSans 240 0 0 80 V_CMFB_S4
port 9 n
flabel metal1 16960 1640 16960 1640 1 FreeSans 240 0 0 80 V_CMFB_S1
port 6 n
flabel metal1 18640 1640 18640 1640 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal1 16125 1640 16125 1640 1 FreeSans 240 0 0 80 ERR_AMP_CUR_BIAS
port 7 n
flabel metal1 17750 1640 17750 1640 1 FreeSans 240 0 0 80 TAIL_CUR_MIR_BIAS
port 5 n
flabel metal1 15805 1640 15805 1640 1 FreeSans 240 0 0 80 V_CMFB_S2
port 10 n
flabel metal1 19415 1635 19415 1635 7 FreeSans 240 0 -160 0 ERR_AMP_REF
port 2 w
flabel metal1 16040 1630 16040 1630 7 FreeSans 240 0 -160 0 VB2_CUR_BIAS
port 11 w
flabel metal1 19560 1635 19560 1635 3 FreeSans 240 0 160 0 VB3_CUR_BIAS
port 8 e
flabel metal2 18430 590 18430 590 5 FreeSans 400 0 0 -40 V_TOP
flabel metal1 18980 1635 18980 1635 1 FreeSans 240 0 0 80 VB1_CUR_BIAS
port 4 n
<< end >>
