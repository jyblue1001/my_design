magic
tech sky130A
timestamp 1751507027
<< metal1 >>
rect 2945 3045 2965 4295
rect 2980 3355 3020 3360
rect 2980 3325 2985 3355
rect 3015 3325 3020 3355
rect 2980 3320 3020 3325
rect 2990 2855 3010 3320
rect 4085 2410 4105 4295
rect 7075 3355 7115 3360
rect 7075 3325 7080 3355
rect 7110 3325 7115 3355
rect 7075 3320 7115 3325
rect 7085 2855 7105 3320
rect 7130 3045 7150 4185
rect 4075 2405 4115 2410
rect 4075 2375 4080 2405
rect 4110 2375 4115 2405
rect 4075 2370 4115 2375
rect 2460 2225 2500 2265
rect 7590 2225 7630 2265
<< via1 >>
rect 2985 3325 3015 3355
rect 7080 3325 7110 3355
rect 4080 2375 4110 2405
<< metal2 >>
rect 2980 3355 3020 3360
rect 2980 3350 2985 3355
rect 2935 3330 2985 3350
rect 2980 3325 2985 3330
rect 3015 3325 3020 3355
rect 2980 3320 3020 3325
rect 7075 3355 7115 3360
rect 7075 3325 7080 3355
rect 7110 3350 7115 3355
rect 7110 3330 7160 3350
rect 7110 3325 7115 3330
rect 7075 3320 7115 3325
rect 4075 2405 4115 2410
rect 4075 2375 4080 2405
rect 4110 2400 4115 2405
rect 4110 2380 4965 2400
rect 4110 2375 4115 2380
rect 4075 2370 4115 2375
rect 4065 2290 4080 2310
rect 2460 2225 2500 2265
rect 7590 2225 7630 2265
rect 4065 2070 4080 2090
<< metal4 >>
rect 940 6700 990 6750
rect 975 0 1025 50
use bgr  bgr_0
timestamp 1751468312
transform -1 0 8031 0 -1 12099
box -200 535 6100 5350
use two_stage_opamp_dummy_magic  two_stage_opamp_dummy_magic_0
timestamp 1751484366
transform 1 0 -26855 0 1 555
box 26855 -555 36545 6195
<< labels >>
flabel metal4 965 6750 965 6750 1 FreeSans 800 0 0 400 VDDA
port 1 n
flabel metal2 7610 2225 7610 2225 5 FreeSans 400 0 0 -200 VOUT+
port 3 s
flabel metal2 4065 2080 4065 2080 7 FreeSans 400 0 -200 0 VIN+
port 5 w
flabel metal2 4065 2300 4065 2300 7 FreeSans 400 0 -200 0 VIN-
port 6 w
flabel metal2 2480 2225 2480 2225 5 FreeSans 400 0 0 -200 VOUT-
port 4 s
flabel metal4 1000 0 1000 0 5 FreeSans 800 0 0 -400 GNDA
port 2 s
<< end >>
