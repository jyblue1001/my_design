magic
tech sky130A
timestamp 1738312014
<< nwell >>
rect 605 105 1335 210
<< nmos >>
rect 665 -35 680 15
rect 845 -35 860 15
rect 900 -35 915 15
rect 1025 -35 1040 15
rect 1080 -35 1095 15
rect 1135 -35 1150 15
rect 1260 -35 1275 15
<< pmos >>
rect 665 125 680 175
rect 720 125 735 175
rect 845 125 860 175
rect 900 125 915 175
rect 1260 125 1275 175
<< ndiff >>
rect 625 0 665 15
rect 625 -20 635 0
rect 655 -20 665 0
rect 625 -35 665 -20
rect 680 0 720 15
rect 680 -20 690 0
rect 710 -20 720 0
rect 680 -35 720 -20
rect 805 0 845 15
rect 805 -20 815 0
rect 835 -20 845 0
rect 805 -35 845 -20
rect 860 0 900 15
rect 860 -20 870 0
rect 890 -20 900 0
rect 860 -35 900 -20
rect 915 0 955 15
rect 915 -20 925 0
rect 945 -20 955 0
rect 915 -35 955 -20
rect 985 0 1025 15
rect 985 -20 995 0
rect 1015 -20 1025 0
rect 985 -35 1025 -20
rect 1040 0 1080 15
rect 1040 -20 1050 0
rect 1070 -20 1080 0
rect 1040 -35 1080 -20
rect 1095 0 1135 15
rect 1095 -20 1105 0
rect 1125 -20 1135 0
rect 1095 -35 1135 -20
rect 1150 0 1190 15
rect 1150 -20 1160 0
rect 1180 -20 1190 0
rect 1150 -35 1190 -20
rect 1220 0 1260 15
rect 1220 -20 1230 0
rect 1250 -20 1260 0
rect 1220 -35 1260 -20
rect 1275 0 1315 15
rect 1275 -20 1285 0
rect 1305 -20 1315 0
rect 1275 -35 1315 -20
<< pdiff >>
rect 625 160 665 175
rect 625 140 635 160
rect 655 140 665 160
rect 625 125 665 140
rect 680 160 720 175
rect 680 140 690 160
rect 710 140 720 160
rect 680 125 720 140
rect 735 160 775 175
rect 735 140 745 160
rect 765 140 775 160
rect 735 125 775 140
rect 805 160 845 175
rect 805 140 815 160
rect 835 140 845 160
rect 805 125 845 140
rect 860 160 900 175
rect 860 140 870 160
rect 890 140 900 160
rect 860 125 900 140
rect 915 160 955 175
rect 915 140 925 160
rect 945 140 955 160
rect 915 125 955 140
rect 1220 160 1260 175
rect 1220 140 1230 160
rect 1250 140 1260 160
rect 1220 125 1260 140
rect 1275 160 1315 175
rect 1275 140 1285 160
rect 1305 140 1315 160
rect 1275 125 1315 140
<< ndiffc >>
rect 635 -20 655 0
rect 690 -20 710 0
rect 815 -20 835 0
rect 870 -20 890 0
rect 925 -20 945 0
rect 995 -20 1015 0
rect 1050 -20 1070 0
rect 1105 -20 1125 0
rect 1160 -20 1180 0
rect 1230 -20 1250 0
rect 1285 -20 1305 0
<< pdiffc >>
rect 635 140 655 160
rect 690 140 710 160
rect 745 140 765 160
rect 815 140 835 160
rect 870 140 890 160
rect 925 140 945 160
rect 1230 140 1250 160
rect 1285 140 1305 160
<< psubdiff >>
rect 765 0 805 15
rect 765 -20 775 0
rect 795 -20 805 0
rect 765 -35 805 -20
<< nsubdiff >>
rect 1180 160 1220 175
rect 1180 140 1190 160
rect 1210 140 1220 160
rect 1180 125 1220 140
<< psubdiffcont >>
rect 775 -20 795 0
<< nsubdiffcont >>
rect 1190 140 1210 160
<< poly >>
rect 820 220 860 230
rect 820 200 830 220
rect 850 200 860 220
rect 665 185 735 200
rect 820 190 860 200
rect 665 175 680 185
rect 720 175 735 185
rect 845 175 860 190
rect 900 175 915 190
rect 1260 175 1275 190
rect 665 70 680 125
rect 720 110 735 125
rect 605 55 680 70
rect 665 15 680 55
rect 705 60 745 70
rect 705 40 715 60
rect 735 40 745 60
rect 705 30 745 40
rect 845 15 860 125
rect 900 110 915 125
rect 1260 110 1275 125
rect 900 100 990 110
rect 900 95 960 100
rect 950 80 960 95
rect 980 80 990 100
rect 950 70 990 80
rect 1135 95 1275 110
rect 885 60 925 70
rect 885 40 895 60
rect 915 40 925 60
rect 1135 40 1150 95
rect 885 30 1150 40
rect 1175 60 1215 70
rect 1175 40 1185 60
rect 1205 45 1215 60
rect 1205 40 1275 45
rect 1175 30 1275 40
rect 900 25 1150 30
rect 900 15 915 25
rect 1025 15 1040 25
rect 1080 15 1095 25
rect 1135 15 1150 25
rect 1260 15 1275 30
rect 665 -50 680 -35
rect 845 -50 860 -35
rect 900 -50 915 -35
rect 1025 -50 1040 -35
rect 1080 -50 1095 -35
rect 1135 -50 1150 -35
rect 1260 -50 1275 -35
<< polycont >>
rect 830 200 850 220
rect 715 40 735 60
rect 960 80 980 100
rect 895 40 915 60
rect 1185 40 1205 60
<< locali >>
rect 820 220 860 230
rect 820 200 830 220
rect 850 210 860 220
rect 850 200 1305 210
rect 820 190 1305 200
rect 1285 170 1305 190
rect 630 160 660 170
rect 630 140 635 160
rect 655 140 660 160
rect 630 130 660 140
rect 685 160 715 170
rect 685 140 690 160
rect 710 140 715 160
rect 685 130 715 140
rect 740 160 770 170
rect 740 140 745 160
rect 765 140 770 160
rect 740 130 770 140
rect 810 160 840 170
rect 810 140 815 160
rect 835 140 840 160
rect 810 130 840 140
rect 865 160 895 170
rect 865 140 870 160
rect 890 140 895 160
rect 865 130 895 140
rect 920 160 1030 170
rect 920 140 925 160
rect 945 150 1030 160
rect 945 140 950 150
rect 920 130 950 140
rect 695 70 715 130
rect 815 110 835 130
rect 815 100 990 110
rect 815 90 960 100
rect 950 80 960 90
rect 980 80 990 100
rect 950 70 990 80
rect 695 60 745 70
rect 695 40 715 60
rect 735 50 745 60
rect 885 60 925 70
rect 885 50 895 60
rect 735 40 895 50
rect 915 40 925 60
rect 695 30 925 40
rect 695 10 715 30
rect 950 10 970 70
rect 1010 50 1030 150
rect 1185 160 1255 170
rect 1185 140 1190 160
rect 1210 140 1230 160
rect 1250 140 1255 160
rect 1185 130 1255 140
rect 1280 160 1310 170
rect 1280 140 1285 160
rect 1305 140 1310 160
rect 1280 130 1310 140
rect 1285 75 1305 130
rect 1175 60 1215 70
rect 1175 50 1185 60
rect 995 40 1185 50
rect 1205 40 1215 60
rect 995 30 1215 40
rect 1285 55 1345 75
rect 995 10 1015 30
rect 1105 10 1125 30
rect 1285 10 1305 55
rect 630 0 660 10
rect 630 -20 635 0
rect 655 -20 660 0
rect 630 -30 660 -20
rect 685 0 715 10
rect 685 -20 690 0
rect 710 -20 715 0
rect 685 -30 715 -20
rect 770 0 840 10
rect 770 -20 775 0
rect 795 -20 815 0
rect 835 -20 840 0
rect 770 -30 840 -20
rect 865 0 895 10
rect 865 -20 870 0
rect 890 -20 895 0
rect 865 -30 895 -20
rect 920 0 970 10
rect 920 -20 925 0
rect 945 -10 970 0
rect 990 0 1020 10
rect 945 -20 950 -10
rect 920 -30 950 -20
rect 990 -20 995 0
rect 1015 -20 1020 0
rect 990 -30 1020 -20
rect 1045 0 1075 10
rect 1045 -20 1050 0
rect 1070 -20 1075 0
rect 1045 -30 1075 -20
rect 1100 0 1130 10
rect 1100 -20 1105 0
rect 1125 -20 1130 0
rect 1100 -30 1130 -20
rect 1155 0 1185 10
rect 1155 -20 1160 0
rect 1180 -20 1185 0
rect 1155 -30 1185 -20
rect 1225 0 1255 10
rect 1225 -20 1230 0
rect 1250 -20 1255 0
rect 1225 -30 1255 -20
rect 1280 0 1310 10
rect 1280 -20 1285 0
rect 1305 -20 1310 0
rect 1280 -30 1310 -20
<< viali >>
rect 635 140 655 160
rect 745 140 765 160
rect 870 140 890 160
rect 1190 140 1210 160
rect 1230 140 1250 160
rect 635 -20 655 0
rect 775 -20 795 0
rect 815 -20 835 0
rect 1050 -20 1070 0
rect 1160 -20 1180 0
rect 1230 -20 1250 0
<< metal1 >>
rect 605 160 1335 175
rect 605 140 635 160
rect 655 140 745 160
rect 765 140 870 160
rect 890 140 1190 160
rect 1210 140 1230 160
rect 1250 140 1335 160
rect 605 125 1335 140
rect 605 0 1335 15
rect 605 -20 635 0
rect 655 -20 775 0
rect 795 -20 815 0
rect 835 -20 1050 0
rect 1070 -20 1160 0
rect 1180 -20 1230 0
rect 1250 -20 1335 0
rect 605 -35 1335 -20
<< labels >>
flabel metal1 605 150 605 150 7 FreeSans 160 0 -80 0 VDDA
flabel metal1 605 -10 605 -10 7 FreeSans 160 0 -80 0 GNDA
flabel poly 605 60 605 60 7 FreeSans 160 0 -80 0 VIN
flabel locali 1345 65 1345 65 3 FreeSans 160 0 80 0 VOUT
flabel locali 1030 80 1030 80 3 FreeSans 160 0 80 0 C
flabel locali 760 50 760 50 1 FreeSans 160 0 0 80 CLK
flabel locali 815 90 815 90 5 FreeSans 160 0 0 0 A
<< end >>
