* NGSPICE file created from pfd.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends


* Top level circuit pfd

Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_0/A sky130_fd_sc_hd__nor2_1_0/B
+ sky130_fd_sc_hd__nor2_1_0/VGND VSUBS sky130_fd_sc_hd__nor2_1_0/VPB sky130_fd_sc_hd__nor2_1_0/VPWR
+ sky130_fd_sc_hd__nor2_1_0/Y sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_1/A sky130_fd_sc_hd__nor2_1_1/B
+ sky130_fd_sc_hd__nor2_1_1/VGND VSUBS sky130_fd_sc_hd__nor2_1_1/VPB sky130_fd_sc_hd__nor2_1_1/VPWR
+ sky130_fd_sc_hd__nor2_1_1/Y sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_2 sky130_fd_sc_hd__nor2_1_2/A sky130_fd_sc_hd__nor2_1_2/B
+ sky130_fd_sc_hd__nor2_1_2/VGND VSUBS sky130_fd_sc_hd__nor2_1_2/VPB sky130_fd_sc_hd__nor2_1_2/VPWR
+ sky130_fd_sc_hd__nor2_1_2/Y sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_3 sky130_fd_sc_hd__nor2_1_3/A sky130_fd_sc_hd__nor2_1_3/B
+ sky130_fd_sc_hd__nor2_1_3/VGND VSUBS sky130_fd_sc_hd__nor2_1_3/VPB sky130_fd_sc_hd__nor2_1_3/VPWR
+ sky130_fd_sc_hd__nor2_1_3/Y sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_4 sky130_fd_sc_hd__nor2_1_4/A sky130_fd_sc_hd__nor2_1_4/B
+ sky130_fd_sc_hd__nor2_1_4/VGND VSUBS sky130_fd_sc_hd__nor2_1_4/VPB sky130_fd_sc_hd__nor2_1_4/VPWR
+ sky130_fd_sc_hd__nor2_1_4/Y sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_5 sky130_fd_sc_hd__nor2_1_5/A sky130_fd_sc_hd__nor2_1_5/B
+ sky130_fd_sc_hd__nor2_1_5/VGND VSUBS sky130_fd_sc_hd__nor2_1_5/VPB sky130_fd_sc_hd__nor2_1_5/VPWR
+ sky130_fd_sc_hd__nor2_1_5/Y sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_6 sky130_fd_sc_hd__nor2_1_6/A sky130_fd_sc_hd__nor2_1_6/B
+ sky130_fd_sc_hd__nor2_1_6/VGND VSUBS sky130_fd_sc_hd__nor2_1_6/VPB sky130_fd_sc_hd__nor2_1_6/VPWR
+ sky130_fd_sc_hd__nor2_1_6/Y sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_7 sky130_fd_sc_hd__nor2_1_7/A sky130_fd_sc_hd__nor2_1_7/B
+ sky130_fd_sc_hd__nor2_1_7/VGND VSUBS sky130_fd_sc_hd__nor2_1_7/VPB sky130_fd_sc_hd__nor2_1_7/VPWR
+ sky130_fd_sc_hd__nor2_1_7/Y sky130_fd_sc_hd__nor2_1
.end

