** sch_path: /foss/designs/my_design/projects/ASU/EEE572/schematic/tb_boost_converter.sch
**.subckt tb_boost_converter
V1 net1 net2 12
V2 V_CTRL_VTC GND pulse(0 1.8 1000ns 200ns 200ns 4800ns 10us)
L46 net4 net1 100u m=1
D1 V_DIODE V_OUT D1N914 area=1
C3 V_CAP net2 100u m=1
R15 net6 net2 2 m=1
R16 V_OUT net5 0.05 m=1
Vmeas net4 V_DIODE 0
.save i(vmeas)
Vmeas1 V_DIODE net3 0
.save i(vmeas1)
Vmeas2 net5 V_CAP 0
.save i(vmeas2)
Vmeas3 V_OUT net6 0
.save i(vmeas3)
M1 net3 V_CTRL_VTC net2 net7 nmos w=5u l=0.18u m=1
**** begin user architecture code
.lib /foss/pdks/sky130A/libs.tech/combined/sky130.lib.spice tt



.options method=gear
.options wnflag=1
.options savecurrents

.include /foss/pdks/volare/gf180mcu/versions/0fe599b2afb6708d281543108caf8310912f54af/gf180mcuD/libs.tech/ngspice/.spiceinit

.control
  save all
  * dc V1 0.0 2.0 0.005
  tran 10ns 200us
  remzerovec
  write tb_boost_converter.raw
  set appendwrite

.endc




**** end user architecture code
**.ends
.GLOBAL GND
.end
