magic
tech sky130A
timestamp 1738239501
<< nwell >>
rect 120 -4500 2050 -3915
<< pwell >>
rect 800 -4600 815 -4595
rect 295 -4730 1610 -4605
rect 860 -4735 1610 -4730
rect 860 -4740 1225 -4735
rect 860 -4800 1025 -4740
rect 1140 -4775 1225 -4740
rect 1140 -4790 1190 -4775
rect 1210 -4790 1225 -4775
rect 1140 -4800 1225 -4790
rect 1170 -4805 1210 -4800
rect 1220 -4830 1260 -4805
<< nmos >>
rect 365 -4710 380 -4610
rect 510 -4710 525 -4610
rect 655 -4710 670 -4610
rect 800 -4710 815 -4610
rect 945 -4710 960 -4610
rect 1090 -4710 1105 -4610
rect 1235 -4710 1250 -4610
rect 1380 -4710 1395 -4610
rect 1525 -4710 1540 -4610
rect 210 -4965 270 -4865
rect 320 -4965 380 -4865
rect 430 -4965 490 -4865
rect 540 -4965 600 -4865
rect 870 -4965 930 -4865
rect 980 -4965 1040 -4865
rect 1090 -4965 1150 -4865
rect 1200 -4965 1260 -4865
rect 1590 -4965 1650 -4865
rect 1700 -4965 1760 -4865
rect 1810 -4965 1870 -4865
rect 1920 -4965 1980 -4865
<< pmos >>
rect 190 -4035 250 -3935
rect 300 -4035 360 -3935
rect 410 -4035 470 -3935
rect 520 -4035 580 -3935
rect 630 -4035 690 -3935
rect 740 -4035 800 -3935
rect 850 -4035 910 -3935
rect 960 -4035 1020 -3935
rect 1150 -4035 1210 -3935
rect 1260 -4035 1320 -3935
rect 1370 -4035 1430 -3935
rect 1480 -4035 1540 -3935
rect 1590 -4035 1650 -3935
rect 1700 -4035 1760 -3935
rect 1810 -4035 1870 -3935
rect 1920 -4035 1980 -3935
rect 365 -4480 380 -4280
rect 510 -4480 525 -4280
rect 655 -4480 670 -4280
rect 800 -4480 815 -4280
rect 945 -4480 960 -4280
rect 1090 -4480 1105 -4280
rect 1235 -4480 1250 -4280
rect 1380 -4480 1395 -4280
rect 1525 -4480 1540 -4280
<< ndiff >>
rect 315 -4625 365 -4610
rect 315 -4695 330 -4625
rect 350 -4695 365 -4625
rect 315 -4710 365 -4695
rect 380 -4625 430 -4610
rect 380 -4695 395 -4625
rect 415 -4695 430 -4625
rect 380 -4710 430 -4695
rect 460 -4625 510 -4610
rect 460 -4695 475 -4625
rect 495 -4695 510 -4625
rect 460 -4710 510 -4695
rect 525 -4625 575 -4610
rect 525 -4695 540 -4625
rect 560 -4695 575 -4625
rect 525 -4710 575 -4695
rect 605 -4625 655 -4610
rect 605 -4695 620 -4625
rect 640 -4695 655 -4625
rect 605 -4710 655 -4695
rect 670 -4625 720 -4610
rect 670 -4695 685 -4625
rect 705 -4695 720 -4625
rect 670 -4710 720 -4695
rect 750 -4625 800 -4610
rect 750 -4695 765 -4625
rect 785 -4695 800 -4625
rect 750 -4710 800 -4695
rect 815 -4625 865 -4610
rect 815 -4695 830 -4625
rect 850 -4695 865 -4625
rect 815 -4710 865 -4695
rect 895 -4625 945 -4610
rect 895 -4695 910 -4625
rect 930 -4695 945 -4625
rect 895 -4710 945 -4695
rect 960 -4625 1010 -4610
rect 960 -4695 975 -4625
rect 995 -4695 1010 -4625
rect 960 -4710 1010 -4695
rect 1040 -4625 1090 -4610
rect 1040 -4695 1055 -4625
rect 1075 -4695 1090 -4625
rect 1040 -4710 1090 -4695
rect 1105 -4625 1155 -4610
rect 1105 -4695 1120 -4625
rect 1140 -4695 1155 -4625
rect 1105 -4710 1155 -4695
rect 1185 -4625 1235 -4610
rect 1185 -4695 1200 -4625
rect 1220 -4695 1235 -4625
rect 1185 -4710 1235 -4695
rect 1250 -4625 1300 -4610
rect 1250 -4695 1265 -4625
rect 1285 -4695 1300 -4625
rect 1250 -4710 1300 -4695
rect 1330 -4625 1380 -4610
rect 1330 -4695 1345 -4625
rect 1365 -4695 1380 -4625
rect 1330 -4710 1380 -4695
rect 1395 -4625 1445 -4610
rect 1395 -4695 1410 -4625
rect 1430 -4695 1445 -4625
rect 1395 -4710 1445 -4695
rect 1475 -4625 1525 -4610
rect 1475 -4695 1490 -4625
rect 1510 -4695 1525 -4625
rect 1475 -4710 1525 -4695
rect 1540 -4625 1590 -4610
rect 1540 -4695 1555 -4625
rect 1575 -4695 1590 -4625
rect 1540 -4710 1590 -4695
rect 160 -4880 210 -4865
rect 160 -4950 175 -4880
rect 195 -4950 210 -4880
rect 160 -4965 210 -4950
rect 270 -4880 320 -4865
rect 270 -4950 285 -4880
rect 305 -4950 320 -4880
rect 270 -4965 320 -4950
rect 380 -4880 430 -4865
rect 380 -4950 395 -4880
rect 415 -4950 430 -4880
rect 380 -4965 430 -4950
rect 490 -4880 540 -4865
rect 490 -4950 505 -4880
rect 525 -4950 540 -4880
rect 490 -4965 540 -4950
rect 600 -4880 650 -4865
rect 600 -4950 615 -4880
rect 635 -4950 650 -4880
rect 600 -4965 650 -4950
rect 820 -4880 870 -4865
rect 820 -4950 835 -4880
rect 855 -4950 870 -4880
rect 820 -4965 870 -4950
rect 930 -4880 980 -4865
rect 930 -4950 945 -4880
rect 965 -4950 980 -4880
rect 930 -4965 980 -4950
rect 1040 -4880 1090 -4865
rect 1040 -4950 1055 -4880
rect 1075 -4950 1090 -4880
rect 1040 -4965 1090 -4950
rect 1150 -4880 1200 -4865
rect 1150 -4950 1165 -4880
rect 1185 -4950 1200 -4880
rect 1150 -4965 1200 -4950
rect 1260 -4880 1310 -4865
rect 1260 -4950 1275 -4880
rect 1295 -4950 1310 -4880
rect 1260 -4965 1310 -4950
rect 1540 -4880 1590 -4865
rect 1540 -4950 1555 -4880
rect 1575 -4950 1590 -4880
rect 1540 -4965 1590 -4950
rect 1650 -4880 1700 -4865
rect 1650 -4950 1665 -4880
rect 1685 -4950 1700 -4880
rect 1650 -4965 1700 -4950
rect 1760 -4880 1810 -4865
rect 1760 -4950 1775 -4880
rect 1795 -4950 1810 -4880
rect 1760 -4965 1810 -4950
rect 1870 -4880 1920 -4865
rect 1870 -4950 1885 -4880
rect 1905 -4950 1920 -4880
rect 1870 -4965 1920 -4950
rect 1980 -4880 2030 -4865
rect 1980 -4950 1995 -4880
rect 2015 -4950 2030 -4880
rect 1980 -4965 2030 -4950
<< pdiff >>
rect 140 -3950 190 -3935
rect 140 -4020 155 -3950
rect 175 -4020 190 -3950
rect 140 -4035 190 -4020
rect 250 -3950 300 -3935
rect 250 -4020 265 -3950
rect 285 -4020 300 -3950
rect 250 -4035 300 -4020
rect 360 -3950 410 -3935
rect 360 -4020 375 -3950
rect 395 -4020 410 -3950
rect 360 -4035 410 -4020
rect 470 -3950 520 -3935
rect 470 -4020 485 -3950
rect 505 -4020 520 -3950
rect 470 -4035 520 -4020
rect 580 -3950 630 -3935
rect 580 -4020 595 -3950
rect 615 -4020 630 -3950
rect 580 -4035 630 -4020
rect 690 -3950 740 -3935
rect 690 -4020 705 -3950
rect 725 -4020 740 -3950
rect 690 -4035 740 -4020
rect 800 -3950 850 -3935
rect 800 -4020 815 -3950
rect 835 -4020 850 -3950
rect 800 -4035 850 -4020
rect 910 -3950 960 -3935
rect 910 -4020 925 -3950
rect 945 -4020 960 -3950
rect 910 -4035 960 -4020
rect 1020 -3950 1070 -3935
rect 1020 -4020 1035 -3950
rect 1055 -4020 1070 -3950
rect 1020 -4035 1070 -4020
rect 1100 -3950 1150 -3935
rect 1100 -4020 1115 -3950
rect 1135 -4020 1150 -3950
rect 1100 -4035 1150 -4020
rect 1210 -3950 1260 -3935
rect 1210 -4020 1225 -3950
rect 1245 -4020 1260 -3950
rect 1210 -4035 1260 -4020
rect 1320 -3950 1370 -3935
rect 1320 -4020 1335 -3950
rect 1355 -4020 1370 -3950
rect 1320 -4035 1370 -4020
rect 1430 -3950 1480 -3935
rect 1430 -4020 1445 -3950
rect 1465 -4020 1480 -3950
rect 1430 -4035 1480 -4020
rect 1540 -3950 1590 -3935
rect 1540 -4020 1555 -3950
rect 1575 -4020 1590 -3950
rect 1540 -4035 1590 -4020
rect 1650 -3950 1700 -3935
rect 1650 -4020 1665 -3950
rect 1685 -4020 1700 -3950
rect 1650 -4035 1700 -4020
rect 1760 -3950 1810 -3935
rect 1760 -4020 1775 -3950
rect 1795 -4020 1810 -3950
rect 1760 -4035 1810 -4020
rect 1870 -3950 1920 -3935
rect 1870 -4020 1885 -3950
rect 1905 -4020 1920 -3950
rect 1870 -4035 1920 -4020
rect 1980 -3950 2030 -3935
rect 1980 -4020 1995 -3950
rect 2015 -4020 2030 -3950
rect 1980 -4035 2030 -4020
rect 315 -4295 365 -4280
rect 315 -4465 330 -4295
rect 350 -4465 365 -4295
rect 315 -4480 365 -4465
rect 380 -4295 430 -4280
rect 380 -4465 395 -4295
rect 415 -4465 430 -4295
rect 380 -4480 430 -4465
rect 460 -4295 510 -4280
rect 460 -4465 475 -4295
rect 495 -4465 510 -4295
rect 460 -4480 510 -4465
rect 525 -4295 575 -4280
rect 525 -4465 540 -4295
rect 560 -4465 575 -4295
rect 525 -4480 575 -4465
rect 605 -4295 655 -4280
rect 605 -4465 620 -4295
rect 640 -4465 655 -4295
rect 605 -4480 655 -4465
rect 670 -4295 720 -4280
rect 670 -4465 685 -4295
rect 705 -4465 720 -4295
rect 670 -4480 720 -4465
rect 750 -4295 800 -4280
rect 750 -4465 765 -4295
rect 785 -4465 800 -4295
rect 750 -4480 800 -4465
rect 815 -4295 865 -4280
rect 815 -4465 830 -4295
rect 850 -4465 865 -4295
rect 815 -4480 865 -4465
rect 895 -4295 945 -4280
rect 895 -4465 910 -4295
rect 930 -4465 945 -4295
rect 895 -4480 945 -4465
rect 960 -4295 1010 -4280
rect 960 -4465 975 -4295
rect 995 -4465 1010 -4295
rect 960 -4480 1010 -4465
rect 1040 -4295 1090 -4280
rect 1040 -4465 1055 -4295
rect 1075 -4465 1090 -4295
rect 1040 -4480 1090 -4465
rect 1105 -4295 1155 -4280
rect 1105 -4465 1120 -4295
rect 1140 -4465 1155 -4295
rect 1105 -4480 1155 -4465
rect 1185 -4295 1235 -4280
rect 1185 -4465 1200 -4295
rect 1220 -4465 1235 -4295
rect 1185 -4480 1235 -4465
rect 1250 -4295 1300 -4280
rect 1250 -4465 1265 -4295
rect 1285 -4465 1300 -4295
rect 1250 -4480 1300 -4465
rect 1330 -4295 1380 -4280
rect 1330 -4465 1345 -4295
rect 1365 -4465 1380 -4295
rect 1330 -4480 1380 -4465
rect 1395 -4295 1445 -4280
rect 1395 -4465 1410 -4295
rect 1430 -4465 1445 -4295
rect 1395 -4480 1445 -4465
rect 1475 -4295 1525 -4280
rect 1475 -4465 1490 -4295
rect 1510 -4465 1525 -4295
rect 1475 -4480 1525 -4465
rect 1540 -4295 1590 -4280
rect 1540 -4465 1555 -4295
rect 1575 -4465 1590 -4295
rect 1540 -4480 1590 -4465
<< ndiffc >>
rect 330 -4695 350 -4625
rect 395 -4695 415 -4625
rect 475 -4695 495 -4625
rect 540 -4695 560 -4625
rect 620 -4695 640 -4625
rect 685 -4695 705 -4625
rect 765 -4695 785 -4625
rect 830 -4695 850 -4625
rect 910 -4695 930 -4625
rect 975 -4695 995 -4625
rect 1055 -4695 1075 -4625
rect 1120 -4695 1140 -4625
rect 1200 -4695 1220 -4625
rect 1265 -4695 1285 -4625
rect 1345 -4695 1365 -4625
rect 1410 -4695 1430 -4625
rect 1490 -4695 1510 -4625
rect 1555 -4695 1575 -4625
rect 175 -4950 195 -4880
rect 285 -4950 305 -4880
rect 395 -4950 415 -4880
rect 505 -4950 525 -4880
rect 615 -4950 635 -4880
rect 835 -4950 855 -4880
rect 945 -4950 965 -4880
rect 1055 -4950 1075 -4880
rect 1165 -4950 1185 -4880
rect 1275 -4950 1295 -4880
rect 1555 -4950 1575 -4880
rect 1665 -4950 1685 -4880
rect 1775 -4950 1795 -4880
rect 1885 -4950 1905 -4880
rect 1995 -4950 2015 -4880
<< pdiffc >>
rect 155 -4020 175 -3950
rect 265 -4020 285 -3950
rect 375 -4020 395 -3950
rect 485 -4020 505 -3950
rect 595 -4020 615 -3950
rect 705 -4020 725 -3950
rect 815 -4020 835 -3950
rect 925 -4020 945 -3950
rect 1035 -4020 1055 -3950
rect 1115 -4020 1135 -3950
rect 1225 -4020 1245 -3950
rect 1335 -4020 1355 -3950
rect 1445 -4020 1465 -3950
rect 1555 -4020 1575 -3950
rect 1665 -4020 1685 -3950
rect 1775 -4020 1795 -3950
rect 1885 -4020 1905 -3950
rect 1995 -4020 2015 -3950
rect 330 -4465 350 -4295
rect 395 -4465 415 -4295
rect 475 -4465 495 -4295
rect 540 -4465 560 -4295
rect 620 -4465 640 -4295
rect 685 -4465 705 -4295
rect 765 -4465 785 -4295
rect 830 -4465 850 -4295
rect 910 -4465 930 -4295
rect 975 -4465 995 -4295
rect 1055 -4465 1075 -4295
rect 1120 -4465 1140 -4295
rect 1200 -4465 1220 -4295
rect 1265 -4465 1285 -4295
rect 1345 -4465 1365 -4295
rect 1410 -4465 1430 -4295
rect 1490 -4465 1510 -4295
rect 1555 -4465 1575 -4295
<< psubdiff >>
rect 1620 -4625 1670 -4610
rect 1620 -4695 1635 -4625
rect 1655 -4695 1670 -4625
rect 1620 -4710 1670 -4695
<< nsubdiff >>
rect 1620 -4295 1670 -4280
rect 1620 -4465 1635 -4295
rect 1655 -4465 1670 -4295
rect 1620 -4480 1670 -4465
<< psubdiffcont >>
rect 1635 -4695 1655 -4625
<< nsubdiffcont >>
rect 1635 -4465 1655 -4295
<< poly >>
rect -40 -3690 2255 -3675
rect -40 -4150 -25 -3690
rect 190 -3935 250 -3920
rect 300 -3935 360 -3920
rect 410 -3935 470 -3920
rect 520 -3935 580 -3920
rect 630 -3935 690 -3920
rect 740 -3935 800 -3920
rect 850 -3935 910 -3920
rect 960 -3935 1020 -3920
rect 1150 -3935 1210 -3920
rect 1260 -3935 1320 -3920
rect 1370 -3935 1430 -3920
rect 1480 -3935 1540 -3920
rect 1590 -3935 1650 -3920
rect 1700 -3935 1760 -3920
rect 1810 -3935 1870 -3920
rect 1920 -3935 1980 -3920
rect 190 -4045 250 -4035
rect 300 -4045 360 -4035
rect 410 -4045 470 -4035
rect 520 -4045 580 -4035
rect 630 -4045 690 -4035
rect 740 -4045 800 -4035
rect 850 -4045 910 -4035
rect 960 -4045 1020 -4035
rect 190 -4065 1020 -4045
rect 1150 -4045 1210 -4035
rect 1260 -4045 1320 -4035
rect 1370 -4045 1430 -4035
rect 1480 -4045 1540 -4035
rect 1590 -4045 1650 -4035
rect 1700 -4045 1760 -4035
rect 1810 -4045 1870 -4035
rect 1920 -4045 1980 -4035
rect 1150 -4060 1980 -4045
rect 2005 -4060 2045 -4050
rect 0 -4135 40 -4125
rect 0 -4150 10 -4135
rect -40 -4155 10 -4150
rect 30 -4155 40 -4135
rect 770 -4150 785 -4065
rect -40 -4165 40 -4155
rect 755 -4160 795 -4150
rect 755 -4180 765 -4160
rect 785 -4180 795 -4160
rect 755 -4190 795 -4180
rect 655 -4230 1540 -4215
rect 1715 -4225 1730 -4060
rect 2005 -4080 2015 -4060
rect 2035 -4080 2045 -4060
rect 2005 -4090 2045 -4080
rect 365 -4280 380 -4265
rect 510 -4280 525 -4265
rect 655 -4280 670 -4230
rect 800 -4280 815 -4265
rect 945 -4280 960 -4265
rect 1090 -4280 1105 -4265
rect 1235 -4280 1250 -4265
rect 1380 -4280 1395 -4265
rect 1525 -4280 1540 -4230
rect 1700 -4235 1740 -4225
rect 1700 -4255 1710 -4235
rect 1730 -4255 1740 -4235
rect 1700 -4265 1740 -4255
rect 2005 -4455 2020 -4090
rect 2060 -4170 2255 -4160
rect 2060 -4190 2070 -4170
rect 2090 -4175 2255 -4170
rect 2090 -4190 2100 -4175
rect 2060 -4200 2100 -4190
rect 2005 -4470 2255 -4455
rect 365 -4535 380 -4480
rect 510 -4520 525 -4480
rect 655 -4520 670 -4480
rect 800 -4495 815 -4480
rect 0 -4550 380 -4535
rect 365 -4610 380 -4550
rect 485 -4530 525 -4520
rect 485 -4550 495 -4530
rect 515 -4550 525 -4530
rect 485 -4560 525 -4550
rect 630 -4530 670 -4520
rect 630 -4550 640 -4530
rect 660 -4550 670 -4530
rect 695 -4505 815 -4495
rect 695 -4525 705 -4505
rect 725 -4510 815 -4505
rect 725 -4525 735 -4510
rect 695 -4535 735 -4525
rect 630 -4560 670 -4550
rect 510 -4610 525 -4560
rect 655 -4585 670 -4560
rect 655 -4600 815 -4585
rect 655 -4610 670 -4600
rect 800 -4610 815 -4600
rect 945 -4610 960 -4480
rect 1090 -4490 1105 -4480
rect 1010 -4505 1105 -4490
rect 1130 -4505 1170 -4495
rect 1235 -4505 1250 -4480
rect 1380 -4505 1395 -4480
rect 1525 -4495 1540 -4480
rect 1010 -4555 1025 -4505
rect 1130 -4525 1140 -4505
rect 1160 -4520 1505 -4505
rect 1160 -4525 1170 -4520
rect 1130 -4530 1170 -4525
rect 985 -4565 1025 -4555
rect 1170 -4560 1210 -4555
rect 985 -4585 995 -4565
rect 1015 -4585 1025 -4565
rect 985 -4595 1025 -4585
rect 1090 -4565 1210 -4560
rect 1090 -4575 1180 -4565
rect 1090 -4610 1105 -4575
rect 1170 -4585 1180 -4575
rect 1200 -4585 1210 -4565
rect 1170 -4595 1210 -4585
rect 1235 -4610 1250 -4520
rect 1490 -4540 1505 -4520
rect 1490 -4555 1540 -4540
rect 1275 -4570 1315 -4560
rect 1275 -4590 1285 -4570
rect 1305 -4585 1315 -4570
rect 1305 -4590 1395 -4585
rect 1275 -4600 1395 -4590
rect 1380 -4610 1395 -4600
rect 1525 -4610 1540 -4555
rect 1715 -4565 1755 -4555
rect 1715 -4585 1725 -4565
rect 1745 -4585 1755 -4565
rect 1715 -4595 1755 -4585
rect 365 -4725 380 -4710
rect 510 -4725 525 -4710
rect 655 -4725 670 -4710
rect 800 -4725 815 -4710
rect 945 -4750 960 -4710
rect 1090 -4725 1105 -4710
rect 0 -4765 960 -4750
rect 1235 -4790 1250 -4710
rect 1380 -4725 1395 -4710
rect 1380 -4735 1435 -4725
rect 1380 -4755 1405 -4735
rect 1425 -4755 1435 -4735
rect 1380 -4765 1435 -4755
rect 1525 -4790 1540 -4710
rect 1170 -4800 1210 -4790
rect 165 -4820 205 -4810
rect 165 -4840 175 -4820
rect 195 -4830 205 -4820
rect 385 -4820 425 -4810
rect 385 -4830 395 -4820
rect 195 -4840 395 -4830
rect 415 -4830 425 -4820
rect 605 -4820 645 -4810
rect 605 -4830 615 -4820
rect 415 -4840 615 -4830
rect 635 -4830 645 -4820
rect 1170 -4820 1180 -4800
rect 1200 -4820 1210 -4800
rect 1235 -4805 1540 -4790
rect 1170 -4830 1210 -4820
rect 635 -4840 1260 -4830
rect 1740 -4840 1755 -4595
rect 2005 -4815 2020 -4470
rect 2005 -4825 2045 -4815
rect 165 -4855 1260 -4840
rect 210 -4865 270 -4855
rect 320 -4865 380 -4855
rect 430 -4865 490 -4855
rect 540 -4865 600 -4855
rect 870 -4865 930 -4855
rect 980 -4865 1040 -4855
rect 1090 -4865 1150 -4855
rect 1200 -4865 1260 -4855
rect 1590 -4855 1980 -4840
rect 2005 -4845 2015 -4825
rect 2035 -4845 2045 -4825
rect 2005 -4855 2045 -4845
rect 1590 -4865 1650 -4855
rect 1700 -4865 1760 -4855
rect 1810 -4865 1870 -4855
rect 1920 -4865 1980 -4855
rect 210 -4980 270 -4965
rect 320 -4980 380 -4965
rect 430 -4980 490 -4965
rect 540 -4980 600 -4965
rect 870 -4980 930 -4965
rect 980 -4980 1040 -4965
rect 1090 -4980 1150 -4965
rect 1200 -4980 1260 -4965
rect 1590 -4980 1650 -4965
rect 1700 -4980 1760 -4965
rect 1810 -4980 1870 -4965
rect 1920 -4980 1980 -4965
<< polycont >>
rect 10 -4155 30 -4135
rect 765 -4180 785 -4160
rect 2015 -4080 2035 -4060
rect 1710 -4255 1730 -4235
rect 2070 -4190 2090 -4170
rect 495 -4550 515 -4530
rect 640 -4550 660 -4530
rect 705 -4525 725 -4505
rect 1140 -4525 1160 -4505
rect 995 -4585 1015 -4565
rect 1180 -4585 1200 -4565
rect 1285 -4590 1305 -4570
rect 1725 -4585 1745 -4565
rect 1405 -4755 1425 -4735
rect 175 -4840 195 -4820
rect 395 -4840 415 -4820
rect 615 -4840 635 -4820
rect 1180 -4820 1200 -4800
rect 2015 -4845 2035 -4825
<< locali >>
rect 155 -3920 1055 -3900
rect 155 -3940 175 -3920
rect 375 -3940 395 -3920
rect 595 -3940 615 -3920
rect 815 -3940 835 -3920
rect 1035 -3940 1055 -3920
rect 1115 -3920 2015 -3900
rect 1115 -3940 1135 -3920
rect 1335 -3940 1355 -3920
rect 1555 -3940 1575 -3920
rect 1775 -3940 1795 -3920
rect 1995 -3940 2015 -3920
rect 145 -3950 185 -3940
rect 145 -4020 155 -3950
rect 175 -4020 185 -3950
rect 145 -4030 185 -4020
rect 255 -3950 295 -3940
rect 255 -4020 265 -3950
rect 285 -4020 295 -3950
rect 255 -4030 295 -4020
rect 365 -3950 405 -3940
rect 365 -4020 375 -3950
rect 395 -4020 405 -3950
rect 365 -4030 405 -4020
rect 475 -3950 515 -3940
rect 475 -4020 485 -3950
rect 505 -4020 515 -3950
rect 475 -4030 515 -4020
rect 585 -3950 625 -3940
rect 585 -4020 595 -3950
rect 615 -4020 625 -3950
rect 585 -4030 625 -4020
rect 695 -3950 735 -3940
rect 695 -4020 705 -3950
rect 725 -4020 735 -3950
rect 695 -4030 735 -4020
rect 805 -3950 845 -3940
rect 805 -4020 815 -3950
rect 835 -4020 845 -3950
rect 805 -4030 845 -4020
rect 915 -3950 955 -3940
rect 915 -4020 925 -3950
rect 945 -4020 955 -3950
rect 915 -4030 955 -4020
rect 1025 -3950 1065 -3940
rect 1025 -4020 1035 -3950
rect 1055 -4020 1065 -3950
rect 1025 -4030 1065 -4020
rect 1105 -3950 1145 -3940
rect 1105 -4020 1115 -3950
rect 1135 -4020 1145 -3950
rect 1105 -4030 1145 -4020
rect 1215 -3950 1255 -3940
rect 1215 -4020 1225 -3950
rect 1245 -4020 1255 -3950
rect 1215 -4030 1255 -4020
rect 1325 -3950 1365 -3940
rect 1325 -4020 1335 -3950
rect 1355 -4020 1365 -3950
rect 1325 -4030 1365 -4020
rect 1435 -3950 1475 -3940
rect 1435 -4020 1445 -3950
rect 1465 -4020 1475 -3950
rect 1435 -4030 1475 -4020
rect 1545 -3950 1585 -3940
rect 1545 -4020 1555 -3950
rect 1575 -4020 1585 -3950
rect 1545 -4030 1585 -4020
rect 1655 -3950 1695 -3940
rect 1655 -4020 1665 -3950
rect 1685 -4020 1695 -3950
rect 1655 -4030 1695 -4020
rect 1765 -3950 1805 -3940
rect 1765 -4020 1775 -3950
rect 1795 -4020 1805 -3950
rect 1765 -4030 1805 -4020
rect 1875 -3950 1915 -3940
rect 1875 -4020 1885 -3950
rect 1905 -4020 1915 -3950
rect 1875 -4030 1915 -4020
rect 1985 -3950 2025 -3940
rect 1985 -4020 1995 -3950
rect 2015 -4020 2025 -3950
rect 1985 -4030 2025 -4020
rect 155 -4050 175 -4030
rect 1035 -4035 1055 -4030
rect 100 -4070 175 -4050
rect 2005 -4050 2025 -4030
rect 2005 -4060 2045 -4050
rect 0 -4135 40 -4125
rect 0 -4155 10 -4135
rect 30 -4145 40 -4135
rect 100 -4145 120 -4070
rect 2005 -4080 2015 -4060
rect 2035 -4080 2045 -4060
rect 2005 -4090 2045 -4080
rect 30 -4155 120 -4145
rect 0 -4165 120 -4155
rect 100 -4725 120 -4165
rect 685 -4130 2205 -4110
rect 685 -4285 705 -4130
rect 755 -4160 795 -4150
rect 755 -4180 765 -4160
rect 785 -4170 2100 -4160
rect 785 -4180 2070 -4170
rect 755 -4190 795 -4180
rect 2060 -4190 2070 -4180
rect 2090 -4190 2100 -4170
rect 765 -4285 785 -4190
rect 2060 -4200 2100 -4190
rect 1700 -4235 1740 -4225
rect 1700 -4245 1710 -4235
rect 830 -4255 1710 -4245
rect 1730 -4245 1740 -4235
rect 1730 -4255 2165 -4245
rect 830 -4265 2165 -4255
rect 830 -4285 850 -4265
rect 1555 -4285 1575 -4265
rect 320 -4295 360 -4285
rect 320 -4465 330 -4295
rect 350 -4465 360 -4295
rect 320 -4475 360 -4465
rect 385 -4295 425 -4285
rect 385 -4465 395 -4295
rect 415 -4465 425 -4295
rect 385 -4475 425 -4465
rect 465 -4295 505 -4285
rect 465 -4465 475 -4295
rect 495 -4465 505 -4295
rect 465 -4475 505 -4465
rect 530 -4295 570 -4285
rect 530 -4465 540 -4295
rect 560 -4465 570 -4295
rect 530 -4475 570 -4465
rect 610 -4295 650 -4285
rect 610 -4465 620 -4295
rect 640 -4465 650 -4295
rect 610 -4475 650 -4465
rect 675 -4295 715 -4285
rect 675 -4465 685 -4295
rect 705 -4465 715 -4295
rect 675 -4475 715 -4465
rect 755 -4295 795 -4285
rect 755 -4465 765 -4295
rect 785 -4465 795 -4295
rect 755 -4475 795 -4465
rect 820 -4295 860 -4285
rect 820 -4465 830 -4295
rect 850 -4465 860 -4295
rect 820 -4475 860 -4465
rect 900 -4295 940 -4285
rect 900 -4465 910 -4295
rect 930 -4465 940 -4295
rect 900 -4475 940 -4465
rect 965 -4295 1005 -4285
rect 965 -4465 975 -4295
rect 995 -4445 1005 -4295
rect 1045 -4295 1085 -4285
rect 995 -4465 1010 -4445
rect 965 -4475 1010 -4465
rect 1045 -4465 1055 -4295
rect 1075 -4465 1085 -4295
rect 1045 -4475 1085 -4465
rect 1110 -4295 1150 -4285
rect 1110 -4465 1120 -4295
rect 1140 -4465 1150 -4295
rect 1110 -4475 1150 -4465
rect 1190 -4295 1230 -4285
rect 1190 -4465 1200 -4295
rect 1220 -4465 1230 -4295
rect 1190 -4475 1230 -4465
rect 1255 -4295 1295 -4285
rect 1255 -4465 1265 -4295
rect 1285 -4465 1295 -4295
rect 1255 -4475 1295 -4465
rect 1335 -4295 1375 -4285
rect 1335 -4465 1345 -4295
rect 1365 -4465 1375 -4295
rect 1335 -4475 1375 -4465
rect 1400 -4295 1440 -4285
rect 1400 -4465 1410 -4295
rect 1430 -4465 1440 -4295
rect 1400 -4475 1440 -4465
rect 1480 -4295 1520 -4285
rect 1480 -4465 1490 -4295
rect 1510 -4465 1520 -4295
rect 1480 -4475 1520 -4465
rect 1545 -4295 1585 -4285
rect 1545 -4465 1555 -4295
rect 1575 -4465 1585 -4295
rect 1545 -4475 1585 -4465
rect 1625 -4295 1665 -4285
rect 1625 -4465 1635 -4295
rect 1655 -4465 1665 -4295
rect 1625 -4475 1665 -4465
rect 405 -4530 425 -4475
rect 485 -4530 525 -4520
rect 405 -4550 495 -4530
rect 515 -4550 525 -4530
rect 405 -4615 425 -4550
rect 485 -4560 525 -4550
rect 550 -4530 570 -4475
rect 695 -4495 715 -4475
rect 695 -4505 735 -4495
rect 630 -4530 670 -4520
rect 550 -4550 640 -4530
rect 660 -4550 670 -4530
rect 550 -4615 570 -4550
rect 630 -4560 670 -4550
rect 695 -4525 705 -4505
rect 725 -4525 735 -4505
rect 695 -4535 735 -4525
rect 695 -4615 715 -4535
rect 765 -4615 785 -4475
rect 820 -4615 840 -4475
rect 920 -4495 940 -4475
rect 1055 -4495 1075 -4475
rect 920 -4515 1075 -4495
rect 920 -4615 940 -4515
rect 985 -4565 1025 -4555
rect 985 -4585 995 -4565
rect 1015 -4585 1025 -4565
rect 985 -4595 1025 -4585
rect 985 -4615 1005 -4595
rect 1055 -4615 1075 -4515
rect 1120 -4495 1140 -4475
rect 1120 -4505 1170 -4495
rect 1120 -4525 1140 -4505
rect 1160 -4525 1170 -4505
rect 1120 -4530 1170 -4525
rect 1120 -4615 1140 -4530
rect 1195 -4555 1215 -4475
rect 1170 -4565 1215 -4555
rect 1170 -4585 1180 -4565
rect 1200 -4585 1215 -4565
rect 1170 -4595 1215 -4585
rect 1275 -4560 1295 -4475
rect 1275 -4570 1315 -4560
rect 1275 -4590 1285 -4570
rect 1305 -4590 1315 -4570
rect 1275 -4600 1315 -4590
rect 1275 -4615 1295 -4600
rect 1345 -4615 1365 -4475
rect 1410 -4555 1430 -4475
rect 1410 -4565 2125 -4555
rect 1410 -4575 1725 -4565
rect 1410 -4615 1430 -4575
rect 1555 -4615 1575 -4575
rect 1715 -4585 1725 -4575
rect 1745 -4575 2125 -4565
rect 1745 -4585 1755 -4575
rect 1715 -4595 1755 -4585
rect 320 -4625 360 -4615
rect 320 -4695 330 -4625
rect 350 -4695 360 -4625
rect 320 -4705 360 -4695
rect 385 -4625 425 -4615
rect 385 -4695 395 -4625
rect 415 -4695 425 -4625
rect 385 -4705 425 -4695
rect 465 -4625 505 -4615
rect 465 -4695 475 -4625
rect 495 -4695 505 -4625
rect 465 -4705 505 -4695
rect 530 -4625 570 -4615
rect 530 -4695 540 -4625
rect 560 -4695 570 -4625
rect 530 -4705 570 -4695
rect 610 -4625 650 -4615
rect 610 -4695 620 -4625
rect 640 -4695 650 -4625
rect 610 -4705 650 -4695
rect 675 -4625 715 -4615
rect 675 -4695 685 -4625
rect 705 -4695 715 -4625
rect 675 -4705 715 -4695
rect 755 -4625 795 -4615
rect 755 -4695 765 -4625
rect 785 -4695 795 -4625
rect 755 -4705 795 -4695
rect 820 -4625 860 -4615
rect 820 -4695 830 -4625
rect 850 -4695 860 -4625
rect 820 -4705 860 -4695
rect 900 -4625 940 -4615
rect 900 -4695 910 -4625
rect 930 -4695 940 -4625
rect 900 -4705 940 -4695
rect 965 -4625 1005 -4615
rect 965 -4695 975 -4625
rect 995 -4695 1005 -4625
rect 965 -4705 1005 -4695
rect 1045 -4625 1085 -4615
rect 1045 -4695 1055 -4625
rect 1075 -4695 1085 -4625
rect 1045 -4705 1085 -4695
rect 1110 -4625 1150 -4615
rect 1110 -4695 1120 -4625
rect 1140 -4695 1150 -4625
rect 1110 -4705 1150 -4695
rect 1190 -4625 1230 -4615
rect 1190 -4695 1200 -4625
rect 1220 -4695 1230 -4625
rect 1190 -4705 1230 -4695
rect 1255 -4625 1295 -4615
rect 1255 -4695 1265 -4625
rect 1285 -4695 1295 -4625
rect 1255 -4705 1295 -4695
rect 1335 -4625 1375 -4615
rect 1335 -4695 1345 -4625
rect 1365 -4695 1375 -4625
rect 1335 -4705 1375 -4695
rect 1400 -4625 1445 -4615
rect 1400 -4695 1410 -4625
rect 1430 -4695 1445 -4625
rect 1400 -4705 1445 -4695
rect 1480 -4625 1520 -4615
rect 1480 -4695 1490 -4625
rect 1510 -4695 1520 -4625
rect 1480 -4705 1520 -4695
rect 1545 -4625 1585 -4615
rect 1545 -4695 1555 -4625
rect 1575 -4695 1585 -4625
rect 1545 -4705 1585 -4695
rect 1625 -4625 1665 -4615
rect 1625 -4695 1635 -4625
rect 1655 -4695 1665 -4625
rect 1625 -4705 1665 -4695
rect 100 -4745 855 -4725
rect 1345 -4740 1365 -4705
rect 165 -4820 205 -4810
rect 165 -4840 175 -4820
rect 195 -4840 205 -4820
rect 165 -4850 205 -4840
rect 385 -4820 425 -4810
rect 385 -4840 395 -4820
rect 415 -4840 425 -4820
rect 385 -4850 425 -4840
rect 605 -4820 645 -4810
rect 605 -4840 615 -4820
rect 635 -4840 645 -4820
rect 605 -4850 645 -4840
rect 175 -4870 195 -4850
rect 395 -4870 415 -4850
rect 615 -4870 635 -4850
rect 835 -4870 855 -4745
rect 1190 -4760 1365 -4740
rect 1395 -4735 1435 -4725
rect 1395 -4755 1405 -4735
rect 1425 -4745 1435 -4735
rect 1425 -4755 2085 -4745
rect 1190 -4790 1210 -4760
rect 1395 -4765 2085 -4755
rect 1170 -4800 1210 -4790
rect 1170 -4820 1180 -4800
rect 1200 -4820 1210 -4800
rect 1170 -4830 1210 -4820
rect 2005 -4825 2045 -4815
rect 2005 -4845 2015 -4825
rect 2035 -4845 2045 -4825
rect 2005 -4855 2045 -4845
rect 1055 -4870 1075 -4865
rect 2005 -4870 2025 -4855
rect 165 -4880 205 -4870
rect 165 -4950 175 -4880
rect 195 -4950 205 -4880
rect 165 -4960 205 -4950
rect 275 -4880 315 -4870
rect 275 -4950 285 -4880
rect 305 -4950 315 -4880
rect 275 -4960 315 -4950
rect 385 -4880 425 -4870
rect 385 -4950 395 -4880
rect 415 -4950 425 -4880
rect 385 -4960 425 -4950
rect 495 -4880 535 -4870
rect 495 -4950 505 -4880
rect 525 -4950 535 -4880
rect 495 -4960 535 -4950
rect 605 -4880 645 -4870
rect 605 -4950 615 -4880
rect 635 -4950 645 -4880
rect 605 -4960 645 -4950
rect 825 -4880 865 -4870
rect 825 -4950 835 -4880
rect 855 -4950 865 -4880
rect 825 -4960 865 -4950
rect 935 -4880 975 -4870
rect 935 -4950 945 -4880
rect 965 -4950 975 -4880
rect 935 -4960 975 -4950
rect 1045 -4880 1085 -4870
rect 1045 -4950 1055 -4880
rect 1075 -4950 1085 -4880
rect 1045 -4960 1085 -4950
rect 1155 -4880 1195 -4870
rect 1155 -4950 1165 -4880
rect 1185 -4950 1195 -4880
rect 1155 -4960 1195 -4950
rect 1265 -4880 1305 -4870
rect 1265 -4950 1275 -4880
rect 1295 -4950 1305 -4880
rect 1265 -4960 1305 -4950
rect 1545 -4880 1585 -4870
rect 1545 -4950 1555 -4880
rect 1575 -4950 1585 -4880
rect 1545 -4960 1585 -4950
rect 1655 -4880 1695 -4870
rect 1655 -4950 1665 -4880
rect 1685 -4950 1695 -4880
rect 1655 -4960 1695 -4950
rect 1765 -4880 1805 -4870
rect 1765 -4950 1775 -4880
rect 1795 -4950 1805 -4880
rect 1765 -4960 1805 -4950
rect 1875 -4880 1915 -4870
rect 1875 -4950 1885 -4880
rect 1905 -4950 1915 -4880
rect 1875 -4960 1915 -4950
rect 1985 -4880 2025 -4870
rect 1985 -4950 1995 -4880
rect 2015 -4950 2025 -4880
rect 1985 -4960 2025 -4950
rect 175 -4980 195 -4960
rect 395 -4980 415 -4960
rect 615 -4980 635 -4960
rect 25 -5000 635 -4980
rect 835 -4980 855 -4960
rect 1055 -4980 1075 -4960
rect 1275 -4980 1295 -4960
rect 835 -5000 1295 -4980
rect 1555 -4980 1575 -4960
rect 1775 -4980 1795 -4960
rect 1995 -4980 2015 -4960
rect 1555 -5000 2015 -4980
rect 2065 -5340 2085 -4765
rect 835 -5360 2085 -5340
rect 835 -5500 860 -5360
rect 2105 -5380 2125 -4575
rect 805 -5510 860 -5500
rect 805 -5545 815 -5510
rect 850 -5545 860 -5510
rect 805 -5555 860 -5545
rect 1025 -5400 2125 -5380
rect 1025 -5500 1045 -5400
rect 2145 -5420 2165 -4265
rect 1335 -5440 2165 -5420
rect 1335 -5500 1355 -5440
rect 2185 -5460 2205 -4130
rect 1025 -5510 1080 -5500
rect 1025 -5545 1035 -5510
rect 1070 -5545 1080 -5510
rect 1025 -5555 1080 -5545
rect 1230 -5510 1355 -5500
rect 1230 -5545 1240 -5510
rect 1275 -5520 1355 -5510
rect 1470 -5480 2205 -5460
rect 1470 -5500 1490 -5480
rect 1470 -5510 1665 -5500
rect 1470 -5520 1620 -5510
rect 1275 -5545 1285 -5520
rect 1230 -5555 1285 -5545
rect 1610 -5545 1620 -5520
rect 1655 -5545 1665 -5510
rect 1610 -5555 1665 -5545
<< viali >>
rect 265 -4020 285 -3950
rect 485 -4020 505 -3950
rect 705 -4020 725 -3950
rect 925 -4020 945 -3950
rect 1225 -4020 1245 -3950
rect 1445 -4020 1465 -3950
rect 1665 -4020 1685 -3950
rect 1885 -4020 1905 -3950
rect 330 -4465 350 -4295
rect 475 -4465 495 -4295
rect 620 -4465 640 -4295
rect 975 -4465 995 -4295
rect 1200 -4465 1220 -4295
rect 1490 -4465 1510 -4295
rect 1635 -4465 1655 -4295
rect 330 -4695 350 -4625
rect 475 -4695 495 -4625
rect 620 -4695 640 -4625
rect 975 -4695 995 -4625
rect 1200 -4695 1220 -4625
rect 1490 -4695 1510 -4625
rect 1635 -4695 1655 -4625
rect 285 -4950 305 -4880
rect 505 -4950 525 -4880
rect 945 -4950 965 -4880
rect 1165 -4950 1185 -4880
rect 1665 -4950 1685 -4880
rect 1885 -4950 1905 -4880
rect 815 -5545 850 -5510
rect 1035 -5545 1070 -5510
rect 1240 -5545 1275 -5510
rect 1620 -5545 1655 -5510
<< metal1 >>
rect 145 -3950 2255 -3845
rect 145 -4020 265 -3950
rect 285 -4020 485 -3950
rect 505 -4020 705 -3950
rect 725 -4020 925 -3950
rect 945 -4020 1225 -3950
rect 1245 -4020 1445 -3950
rect 1465 -4020 1665 -3950
rect 1685 -4020 1885 -3950
rect 1905 -4020 2255 -3950
rect 145 -4295 2255 -4020
rect 145 -4465 330 -4295
rect 350 -4465 475 -4295
rect 495 -4465 620 -4295
rect 640 -4465 975 -4295
rect 995 -4465 1200 -4295
rect 1220 -4465 1490 -4295
rect 1510 -4465 1635 -4295
rect 1655 -4465 2255 -4295
rect 145 -4480 2255 -4465
rect 145 -4625 2255 -4610
rect 145 -4695 330 -4625
rect 350 -4695 475 -4625
rect 495 -4695 620 -4625
rect 640 -4695 975 -4625
rect 995 -4695 1200 -4625
rect 1220 -4695 1490 -4625
rect 1510 -4695 1635 -4625
rect 1655 -4695 2255 -4625
rect 145 -4880 2255 -4695
rect 145 -4950 285 -4880
rect 305 -4950 505 -4880
rect 525 -4950 945 -4880
rect 965 -4950 1165 -4880
rect 1185 -4950 1665 -4880
rect 1685 -4950 1885 -4880
rect 1905 -4950 2255 -4880
rect 145 -4965 2255 -4950
rect 805 -5510 860 -5500
rect 805 -5545 815 -5510
rect 850 -5545 860 -5510
rect 805 -5555 860 -5545
rect 1025 -5510 1080 -5500
rect 1025 -5545 1035 -5510
rect 1070 -5545 1080 -5510
rect 1025 -5555 1080 -5545
rect 1230 -5510 1285 -5500
rect 1230 -5545 1240 -5510
rect 1275 -5545 1285 -5510
rect 1230 -5555 1285 -5545
rect 1610 -5510 1665 -5500
rect 1610 -5545 1620 -5510
rect 1655 -5545 1665 -5510
rect 1610 -5555 1665 -5545
<< via1 >>
rect 815 -5545 850 -5510
rect 1035 -5545 1070 -5510
rect 1240 -5545 1275 -5510
rect 1620 -5545 1655 -5510
<< metal2 >>
rect 805 -5510 860 -5500
rect 805 -5545 815 -5510
rect 850 -5545 860 -5510
rect 805 -5555 860 -5545
rect 1025 -5510 1080 -5500
rect 1025 -5545 1035 -5510
rect 1070 -5545 1080 -5510
rect 1025 -5555 1080 -5545
rect 1230 -5510 1285 -5500
rect 1230 -5545 1240 -5510
rect 1275 -5545 1285 -5510
rect 1230 -5555 1285 -5545
rect 1610 -5510 1665 -5500
rect 1610 -5545 1620 -5510
rect 1655 -5545 1665 -5510
rect 1610 -5555 1665 -5545
<< via2 >>
rect 815 -5545 850 -5510
rect 1035 -5545 1070 -5510
rect 1240 -5545 1275 -5510
rect 1620 -5545 1655 -5510
<< metal3 >>
rect 805 -5510 860 -5500
rect 805 -5545 815 -5510
rect 850 -5545 860 -5510
rect 805 -5675 860 -5545
rect 1025 -5510 1080 -5500
rect 1025 -5545 1035 -5510
rect 1070 -5545 1080 -5510
rect 1025 -5555 1080 -5545
rect 1230 -5510 1285 -5500
rect 1230 -5545 1240 -5510
rect 1275 -5545 1285 -5510
rect 1230 -5555 1285 -5545
rect 1610 -5510 1665 -5500
rect 1610 -5545 1620 -5510
rect 1655 -5545 1665 -5510
rect 1610 -5675 1665 -5545
rect 805 -5965 1095 -5675
rect 1215 -6305 1665 -5675
<< via3 >>
rect 1035 -5545 1070 -5510
rect 1240 -5545 1275 -5510
<< mimcap >>
rect 820 -5700 1080 -5690
rect 820 -5735 1035 -5700
rect 1070 -5735 1080 -5700
rect 820 -5950 1080 -5735
rect 1230 -5700 1650 -5690
rect 1230 -5735 1240 -5700
rect 1275 -5735 1650 -5700
rect 1230 -6290 1650 -5735
<< mimcapcontact >>
rect 1035 -5735 1070 -5700
rect 1240 -5735 1275 -5700
<< metal4 >>
rect 1025 -5510 1080 -5500
rect 1025 -5545 1035 -5510
rect 1070 -5545 1080 -5510
rect 1025 -5700 1080 -5545
rect 1025 -5735 1035 -5700
rect 1070 -5735 1080 -5700
rect 1025 -5745 1080 -5735
rect 1230 -5510 1285 -5500
rect 1230 -5545 1240 -5510
rect 1275 -5545 1285 -5510
rect 1230 -5700 1285 -5545
rect 1230 -5735 1240 -5700
rect 1275 -5735 1285 -5700
rect 1230 -5745 1285 -5735
<< labels >>
flabel poly 0 -4540 0 -4540 7 FreeSans 400 0 -200 0 UP_PFD
flabel poly 0 -4760 0 -4760 7 FreeSans 400 0 -200 0 DOWN_PFD
flabel locali 25 -4990 25 -4990 7 FreeSans 400 0 -200 0 I_IN
<< end >>
