* PEX produced on Mon Feb 17 07:07:27 AM CET 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from opamp_cell_4.ext - technology: sky130A

.subckt rail_to_rail_opamp_magic VDDA VIN+ VIN- VOUT GNDA
X0 VDDA.t34 n_left.t4 n_left.t5 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X1 a_7050_3820.t3 a_7050_3820.t2 GNDA.t15 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X2 GNDA.t6 a_7340_3850.t5 VOUT.t7 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X3 VDDA.t15 p_bias.t7 p_bias.t8 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X4 a_7170_3160.t1 VIN-.t0 n_left.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X5 p_bias.t0 a_7070_3110.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_5p73 l=1
X6 VDDA.t24 p_bias.t9 a_6820_4420.t7 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X7 a_6820_4420.t12 a_6820_4420.t11 a_6820_4420.t12 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X8 a_6820_4420.t6 p_bias.t10 VDDA.t6 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X9 GNDA.t9 a_7070_3110.t7 a_7070_3110.t8 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X10 p_bias.t6 p_bias.t5 VDDA.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X11 p_bias.t4 p_bias.t3 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X12 GNDA.t30 GNDA.t29 GNDA.t30 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X13 GNDA.t5 a_7070_3110.t9 a_7170_3160.t2 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X14 a_6820_4420.t2 VIN+.t0 a_7340_3850.t0 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X15 a_7170_3160.t3 a_7070_3110.t10 GNDA.t10 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X16 VDDA.t55 VDDA.t52 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X17 a_7070_3110.t6 a_7070_3110.t5 GNDA.t33 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X18 VDDA.t51 VDDA.t49 VDDA.t51 VDDA.t50 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X19 VOUT.t2 n_right.t5 VDDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X20 GNDA.t14 a_7050_3820.t6 a_7340_3850.t4 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X21 a_7070_3110.t4 a_7070_3110.t3 GNDA.t35 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X22 a_7340_3850.t2 VIN+.t1 a_6820_4420.t3 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X23 n_left.t3 n_left.t2 VDDA.t32 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X24 a_7340_3850.t1 a_10210_2370.t0 GNDA.t7 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X25 a_7170_3160.t12 a_7170_3160.t11 a_7170_3160.t12 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X26 VOUT.t6 a_7340_3850.t6 GNDA.t34 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X27 GNDA.t28 GNDA.t26 GNDA.t27 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X28 VOUT.t8 a_10210_2370.t1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X29 VDDA.t4 n_right.t6 VOUT.t0 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X30 a_7340_3850.t3 a_7050_3820.t7 GNDA.t13 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X31 n_left.t1 VIN-.t1 a_7170_3160.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X32 VOUT.t9 a_10210_5296.t1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X33 VDDA.t48 VDDA.t45 VDDA.t47 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X34 GNDA.t32 a_7340_3850.t7 VOUT.t5 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X35 a_6820_4420.t5 p_bias.t11 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X36 VDDA.t44 VDDA.t42 VDDA.t44 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X37 VOUT.t1 n_right.t7 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X38 a_7170_3160.t10 a_7170_3160.t8 a_7170_3160.t9 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X39 VDDA.t13 p_bias.t12 a_6820_4420.t4 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X40 VDDA.t17 p_bias.t1 p_bias.t2 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X41 VOUT.t4 a_7340_3850.t8 GNDA.t2 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X42 a_7170_3160.t7 a_7070_3110.t11 GNDA.t31 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X43 GNDA.t25 GNDA.t24 GNDA.t25 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X44 a_10210_5296.t0 n_right.t0 GNDA.t1 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X45 a_6820_4420.t10 a_6820_4420.t8 a_6820_4420.t9 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X46 VDDA.t30 n_left.t6 n_right.t4 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X47 VDDA.t41 VDDA.t38 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X48 GNDA.t11 a_7070_3110.t12 a_7170_3160.t6 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X49 a_6820_4420.t1 VIN-.t2 a_7050_3820.t1 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X50 VDDA.t37 VDDA.t35 VDDA.t37 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X51 GNDA.t23 GNDA.t21 GNDA.t22 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X52 a_7170_3160.t4 VIN+.t2 n_right.t2 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X53 GNDA.t8 a_7070_3110.t1 a_7070_3110.t2 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X54 GNDA.t20 GNDA.t18 GNDA.t19 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X55 n_right.t3 n_left.t7 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X56 GNDA.t12 a_7050_3820.t4 a_7050_3820.t5 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X57 GNDA.t17 GNDA.t16 GNDA.t17 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X58 a_7050_3820.t0 VIN-.t3 a_6820_4420.t0 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X59 VDDA.t57 n_right.t8 VOUT.t3 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X60 n_right.t1 VIN+.t3 a_7170_3160.t5 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
R0 n_left.n1 n_left.t6 401.668
R1 n_left.n5 n_left.n4 325.248
R2 n_left.n4 n_left.n0 313
R3 n_left.n3 n_left.t2 252.248
R4 n_left.n2 n_left.n1 208.868
R5 n_left.n1 n_left.t7 192.8
R6 n_left.n2 n_left.t4 192.8
R7 n_left.n4 n_left.n3 152
R8 n_left.n0 n_left.t0 60.0005
R9 n_left.n0 n_left.t1 60.0005
R10 n_left.n3 n_left.n2 59.4472
R11 n_left.t5 n_left.n5 49.2505
R12 n_left.n5 n_left.t3 49.2505
R13 VDDA.n98 VDDA.n3 585
R14 VDDA.n76 VDDA.n68 585
R15 VDDA.n16 VDDA.t35 384.967
R16 VDDA.n81 VDDA.t49 384.967
R17 VDDA.n85 VDDA.t45 384.967
R18 VDDA.n20 VDDA.t38 384.967
R19 VDDA.n69 VDDA.t42 374.878
R20 VDDA.n99 VDDA.t52 352.834
R21 VDDA.n86 VDDA.t48 341.752
R22 VDDA.n80 VDDA.t51 341.752
R23 VDDA.n19 VDDA.t41 341.752
R24 VDDA.n15 VDDA.t37 341.75
R25 VDDA.n22 VDDA.n13 315.647
R26 VDDA.n83 VDDA.n7 315.647
R27 VDDA.n84 VDDA.n5 315.647
R28 VDDA.n82 VDDA.n8 315.647
R29 VDDA.n21 VDDA.n18 315.647
R30 VDDA.n17 VDDA.n14 315.647
R31 VDDA.n15 VDDA.t36 304.659
R32 VDDA.n92 VDDA.n3 290.733
R33 VDDA.n90 VDDA.n3 290.733
R34 VDDA.n74 VDDA.n68 290.733
R35 VDDA.n70 VDDA.n68 290.733
R36 VDDA.n90 VDDA.n88 233.841
R37 VDDA.n77 VDDA.n76 230.308
R38 VDDA.n69 VDDA.n10 230.308
R39 VDDA.n19 VDDA.n9 185.001
R40 VDDA.n80 VDDA.n79 185.001
R41 VDDA.n87 VDDA.n86 185.001
R42 VDDA.n75 VDDA.n12 185
R43 VDDA.n73 VDDA.n11 185
R44 VDDA.n78 VDDA.n11 185
R45 VDDA.n72 VDDA.n71 185
R46 VDDA.n91 VDDA.n89 185
R47 VDDA.n94 VDDA.n93 185
R48 VDDA.n4 VDDA.n2 185
R49 VDDA.n98 VDDA.n97 185
R50 VDDA.n97 VDDA.n96 185
R51 VDDA.t7 VDDA.t16 145.038
R52 VDDA.n94 VDDA.n89 120.001
R53 VDDA.n97 VDDA.n4 120.001
R54 VDDA.n12 VDDA.n11 120.001
R55 VDDA.n71 VDDA.n11 120.001
R56 VDDA.n67 VDDA.n66 119.737
R57 VDDA.n26 VDDA.n25 119.737
R58 VDDA.n31 VDDA.n30 119.737
R59 VDDA.n35 VDDA.n34 119.737
R60 VDDA.n38 VDDA.n37 119.737
R61 VDDA.t39 VDDA.n9 119.656
R62 VDDA.n79 VDDA.n78 108.779
R63 VDDA.t36 VDDA.t56 94.2753
R64 VDDA.t56 VDDA.t21 94.2753
R65 VDDA.t21 VDDA.t3 94.2753
R66 VDDA.t3 VDDA.t18 94.2753
R67 VDDA.t18 VDDA.t39 94.2753
R68 VDDA.t29 VDDA.t27 94.2753
R69 VDDA.t31 VDDA.t46 94.2753
R70 VDDA.n87 VDDA.t0 94.2753
R71 VDDA.t11 VDDA.t26 94.2753
R72 VDDA.t2 VDDA.t20 94.2753
R73 VDDA.t43 VDDA.t50 83.3974
R74 VDDA.t25 VDDA.t12 83.3974
R75 VDDA.n83 VDDA.n82 83.2005
R76 VDDA.n84 VDDA.n83 83.2005
R77 VDDA.n22 VDDA.n17 83.2005
R78 VDDA.n22 VDDA.n21 83.2005
R79 VDDA.t9 VDDA.t33 76.1455
R80 VDDA.t58 VDDA.t53 76.1455
R81 VDDA.n78 VDDA.n77 69.8479
R82 VDDA.n78 VDDA.n10 69.8479
R83 VDDA.n96 VDDA.n88 69.8479
R84 VDDA.n96 VDDA.n95 69.8479
R85 VDDA.n23 VDDA.n22 69.3203
R86 VDDA.t33 VDDA.t14 68.8936
R87 VDDA.n96 VDDA.t58 68.8936
R88 VDDA.t50 VDDA.t23 61.6417
R89 VDDA.t5 VDDA.t25 61.6417
R90 VDDA.t16 VDDA.n87 50.7639
R91 VDDA.n13 VDDA.t22 49.2505
R92 VDDA.n13 VDDA.t4 49.2505
R93 VDDA.n7 VDDA.t28 49.2505
R94 VDDA.n7 VDDA.t34 49.2505
R95 VDDA.n5 VDDA.t32 49.2505
R96 VDDA.n5 VDDA.t47 49.2505
R97 VDDA.t51 VDDA.n8 49.2505
R98 VDDA.n8 VDDA.t30 49.2505
R99 VDDA.n18 VDDA.t19 49.2505
R100 VDDA.n18 VDDA.t40 49.2505
R101 VDDA.t37 VDDA.n14 49.2505
R102 VDDA.n14 VDDA.t57 49.2505
R103 VDDA.n89 VDDA.n88 45.3071
R104 VDDA.n95 VDDA.n94 45.3071
R105 VDDA.n71 VDDA.n10 45.3071
R106 VDDA.n77 VDDA.n12 45.3071
R107 VDDA.n95 VDDA.n4 45.3071
R108 VDDA.n83 VDDA.n6 41.6005
R109 VDDA.t26 VDDA.t7 39.886
R110 VDDA.n64 VDDA.n23 39.4988
R111 VDDA.n101 VDDA.n0 39.4379
R112 VDDA.n79 VDDA.t43 36.26
R113 VDDA VDDA.n101 33.434
R114 VDDA.t23 VDDA.t29 32.6341
R115 VDDA.t20 VDDA.t5 32.6341
R116 VDDA.n64 VDDA.n63 32.0005
R117 VDDA.n63 VDDA.n62 32.0005
R118 VDDA.n59 VDDA.n58 32.0005
R119 VDDA.n58 VDDA.n27 32.0005
R120 VDDA.n54 VDDA.n27 32.0005
R121 VDDA.n54 VDDA.n53 32.0005
R122 VDDA.n53 VDDA.n52 32.0005
R123 VDDA.n52 VDDA.n29 32.0005
R124 VDDA.n48 VDDA.n29 32.0005
R125 VDDA.n48 VDDA.n47 32.0005
R126 VDDA.n47 VDDA.n46 32.0005
R127 VDDA.n46 VDDA.n33 32.0005
R128 VDDA.n42 VDDA.n33 32.0005
R129 VDDA.n42 VDDA.n41 32.0005
R130 VDDA.n41 VDDA.n40 32.0005
R131 VDDA.n40 VDDA.n0 32.0005
R132 VDDA.n86 VDDA.n85 30.754
R133 VDDA.n20 VDDA.n19 30.754
R134 VDDA.n16 VDDA.n15 30.186
R135 VDDA.n81 VDDA.n80 30.186
R136 VDDA.n62 VDDA.n6 25.6005
R137 VDDA.t14 VDDA.t31 25.3822
R138 VDDA.t46 VDDA.t0 25.3822
R139 VDDA.n99 VDDA.n98 22.0449
R140 VDDA.n3 VDDA.t55 19.7005
R141 VDDA.t44 VDDA.n67 19.7005
R142 VDDA.n67 VDDA.t24 19.7005
R143 VDDA.n25 VDDA.t10 19.7005
R144 VDDA.n25 VDDA.t15 19.7005
R145 VDDA.n30 VDDA.t1 19.7005
R146 VDDA.n30 VDDA.t17 19.7005
R147 VDDA.n34 VDDA.t8 19.7005
R148 VDDA.n34 VDDA.t13 19.7005
R149 VDDA.n37 VDDA.t6 19.7005
R150 VDDA.n37 VDDA.t54 19.7005
R151 VDDA.n68 VDDA.t44 19.7005
R152 VDDA.t27 VDDA.t9 18.1303
R153 VDDA.t53 VDDA.t2 18.1303
R154 VDDA.n85 VDDA.n84 16.0005
R155 VDDA.n82 VDDA.n81 16.0005
R156 VDDA.n21 VDDA.n20 16.0005
R157 VDDA.n17 VDDA.n16 16.0005
R158 VDDA.t12 VDDA.t11 10.8784
R159 VDDA.n100 VDDA.n99 9.613
R160 VDDA.n65 VDDA.n64 9.3005
R161 VDDA.n63 VDDA.n24 9.3005
R162 VDDA.n62 VDDA.n61 9.3005
R163 VDDA.n60 VDDA.n59 9.3005
R164 VDDA.n58 VDDA.n57 9.3005
R165 VDDA.n56 VDDA.n27 9.3005
R166 VDDA.n55 VDDA.n54 9.3005
R167 VDDA.n53 VDDA.n28 9.3005
R168 VDDA.n52 VDDA.n51 9.3005
R169 VDDA.n50 VDDA.n29 9.3005
R170 VDDA.n49 VDDA.n48 9.3005
R171 VDDA.n47 VDDA.n32 9.3005
R172 VDDA.n46 VDDA.n45 9.3005
R173 VDDA.n44 VDDA.n33 9.3005
R174 VDDA.n43 VDDA.n42 9.3005
R175 VDDA.n41 VDDA.n36 9.3005
R176 VDDA.n40 VDDA.n39 9.3005
R177 VDDA.n1 VDDA.n0 9.3005
R178 VDDA.n78 VDDA.n9 7.25241
R179 VDDA.n93 VDDA.n91 7.11161
R180 VDDA.n98 VDDA.n2 7.11161
R181 VDDA.n76 VDDA.n75 7.11161
R182 VDDA.n73 VDDA.n72 7.11161
R183 VDDA.n59 VDDA.n6 6.4005
R184 VDDA.n93 VDDA.n92 3.53508
R185 VDDA.n91 VDDA.n90 3.53508
R186 VDDA.n92 VDDA.n2 3.53508
R187 VDDA.n75 VDDA.n74 3.53508
R188 VDDA.n72 VDDA.n70 3.53508
R189 VDDA.n74 VDDA.n73 3.53508
R190 VDDA.n70 VDDA.n69 3.53508
R191 VDDA.n101 VDDA.n100 0.1925
R192 VDDA.n65 VDDA.n24 0.15675
R193 VDDA.n61 VDDA.n24 0.15675
R194 VDDA.n61 VDDA.n60 0.15675
R195 VDDA.n57 VDDA.n56 0.15675
R196 VDDA.n56 VDDA.n55 0.15675
R197 VDDA.n55 VDDA.n28 0.15675
R198 VDDA.n51 VDDA.n50 0.15675
R199 VDDA.n50 VDDA.n49 0.15675
R200 VDDA.n49 VDDA.n32 0.15675
R201 VDDA.n45 VDDA.n44 0.15675
R202 VDDA.n44 VDDA.n43 0.15675
R203 VDDA.n43 VDDA.n36 0.15675
R204 VDDA.n39 VDDA.n1 0.15675
R205 VDDA.n66 VDDA.n23 0.100307
R206 VDDA.n66 VDDA.n65 0.09425
R207 VDDA.n57 VDDA.n26 0.09425
R208 VDDA.n51 VDDA.n31 0.09425
R209 VDDA.n45 VDDA.n35 0.09425
R210 VDDA.n39 VDDA.n38 0.09425
R211 VDDA.n60 VDDA.n26 0.063
R212 VDDA.n31 VDDA.n28 0.063
R213 VDDA.n35 VDDA.n32 0.063
R214 VDDA.n38 VDDA.n36 0.063
R215 VDDA.n100 VDDA.n1 0.063
R216 a_7050_3820.n5 a_7050_3820.n4 427.647
R217 a_7050_3820.n1 a_7050_3820.t6 321.334
R218 a_7050_3820.n4 a_7050_3820.n0 210.601
R219 a_7050_3820.n2 a_7050_3820.n1 208.868
R220 a_7050_3820.n3 a_7050_3820.t2 174.056
R221 a_7050_3820.n4 a_7050_3820.n3 152
R222 a_7050_3820.n2 a_7050_3820.t4 112.468
R223 a_7050_3820.n1 a_7050_3820.t7 112.468
R224 a_7050_3820.n3 a_7050_3820.n2 61.5894
R225 a_7050_3820.n0 a_7050_3820.t5 60.0005
R226 a_7050_3820.n0 a_7050_3820.t3 60.0005
R227 a_7050_3820.n5 a_7050_3820.t1 49.2505
R228 a_7050_3820.t0 a_7050_3820.n5 49.2505
R229 GNDA.t0 GNDA.t1 36609.1
R230 GNDA.n16 GNDA.t1 3567.2
R231 GNDA.n73 GNDA.t0 1186
R232 GNDA.t0 GNDA.n11 1186
R233 GNDA.t0 GNDA.n10 1186
R234 GNDA.t0 GNDA.n72 1186
R235 GNDA.n16 GNDA.t3 806.668
R236 GNDA.t0 GNDA.n69 614.872
R237 GNDA.n66 GNDA.n18 589.889
R238 GNDA.n15 GNDA.n14 589.889
R239 GNDA.n68 GNDA.n67 585
R240 GNDA.n69 GNDA.n68 585
R241 GNDA.n18 GNDA.n17 585
R242 GNDA.n13 GNDA.n12 585
R243 GNDA.n69 GNDA.n12 585
R244 GNDA.n17 GNDA.n15 585
R245 GNDA.n16 GNDA.t7 340.536
R246 GNDA.n71 GNDA.t29 304.634
R247 GNDA.n74 GNDA.t21 304.634
R248 GNDA.n24 GNDA.t16 304.634
R249 GNDA.n27 GNDA.t18 304.634
R250 GNDA.n19 GNDA.t24 292.584
R251 GNDA.n1 GNDA.t26 292.584
R252 GNDA.n15 GNDA.n12 275.8
R253 GNDA.n68 GNDA.n18 275.8
R254 GNDA.n72 GNDA.t30 245
R255 GNDA.n73 GNDA.t23 245
R256 GNDA.t17 GNDA.n10 245
R257 GNDA.n11 GNDA.t20 245
R258 GNDA.n76 GNDA.n7 204.201
R259 GNDA.n25 GNDA.n23 204.201
R260 GNDA.n29 GNDA.n22 204.201
R261 GNDA.n28 GNDA.n26 204.201
R262 GNDA.n70 GNDA.n8 204.201
R263 GNDA.n75 GNDA.n9 204.201
R264 GNDA.n17 GNDA.n16 150.052
R265 GNDA.n66 GNDA.t25 132.058
R266 GNDA.n14 GNDA.t28 132.058
R267 GNDA.n3 GNDA.n2 97.8707
R268 GNDA.n43 GNDA.n42 97.8707
R269 GNDA.n50 GNDA.n39 97.8707
R270 GNDA.n57 GNDA.n36 97.8707
R271 GNDA.n65 GNDA.n64 97.8707
R272 GNDA.n76 GNDA.n8 83.2005
R273 GNDA.n76 GNDA.n75 83.2005
R274 GNDA.n69 GNDA.t4 78.9749
R275 GNDA.n17 GNDA.t4 78.9749
R276 GNDA.n29 GNDA.n25 66.5605
R277 GNDA.n29 GNDA.n28 66.5605
R278 GNDA.n30 GNDA.n29 65.9634
R279 GNDA.n7 GNDA.t13 60.0005
R280 GNDA.n7 GNDA.t12 60.0005
R281 GNDA.n23 GNDA.t17 60.0005
R282 GNDA.n23 GNDA.t6 60.0005
R283 GNDA.n22 GNDA.t34 60.0005
R284 GNDA.n22 GNDA.t32 60.0005
R285 GNDA.n26 GNDA.t2 60.0005
R286 GNDA.n26 GNDA.t19 60.0005
R287 GNDA.t30 GNDA.n70 60.0005
R288 GNDA.n70 GNDA.t14 60.0005
R289 GNDA.n9 GNDA.t15 60.0005
R290 GNDA.n9 GNDA.t22 60.0005
R291 GNDA.n77 GNDA.n76 41.6005
R292 GNDA.n33 GNDA.n30 39.4985
R293 GNDA.n87 GNDA.n0 39.1796
R294 GNDA GNDA.n87 33.0217
R295 GNDA.n34 GNDA.n33 32.0005
R296 GNDA.n62 GNDA.n34 32.0005
R297 GNDA.n62 GNDA.n61 32.0005
R298 GNDA.n61 GNDA.n60 32.0005
R299 GNDA.n60 GNDA.n35 32.0005
R300 GNDA.n55 GNDA.n35 32.0005
R301 GNDA.n55 GNDA.n54 32.0005
R302 GNDA.n54 GNDA.n53 32.0005
R303 GNDA.n53 GNDA.n38 32.0005
R304 GNDA.n48 GNDA.n38 32.0005
R305 GNDA.n48 GNDA.n47 32.0005
R306 GNDA.n47 GNDA.n46 32.0005
R307 GNDA.n46 GNDA.n41 32.0005
R308 GNDA.n41 GNDA.n6 32.0005
R309 GNDA.n78 GNDA.n6 32.0005
R310 GNDA.n82 GNDA.n4 32.0005
R311 GNDA.n83 GNDA.n82 32.0005
R312 GNDA.n83 GNDA.n0 32.0005
R313 GNDA.n27 GNDA.n11 27.2005
R314 GNDA.n24 GNDA.n10 27.2005
R315 GNDA.n74 GNDA.n73 25.6005
R316 GNDA.n72 GNDA.n71 25.6005
R317 GNDA.n77 GNDA.n4 25.6005
R318 GNDA.n2 GNDA.t10 24.0005
R319 GNDA.n2 GNDA.t27 24.0005
R320 GNDA.n42 GNDA.t33 24.0005
R321 GNDA.n42 GNDA.t11 24.0005
R322 GNDA.n39 GNDA.t35 24.0005
R323 GNDA.n39 GNDA.t8 24.0005
R324 GNDA.n36 GNDA.t31 24.0005
R325 GNDA.n36 GNDA.t9 24.0005
R326 GNDA.t25 GNDA.n65 24.0005
R327 GNDA.n65 GNDA.t5 24.0005
R328 GNDA.n13 GNDA.n1 22.4005
R329 GNDA.n67 GNDA.n19 22.4005
R330 GNDA.n28 GNDA.n27 14.0805
R331 GNDA.n25 GNDA.n24 14.0805
R332 GNDA.n75 GNDA.n74 12.8005
R333 GNDA.n71 GNDA.n8 12.8005
R334 GNDA.n86 GNDA.n1 9.58175
R335 GNDA.n31 GNDA.n19 9.58175
R336 GNDA.n85 GNDA.n0 9.3005
R337 GNDA.n84 GNDA.n83 9.3005
R338 GNDA.n82 GNDA.n81 9.3005
R339 GNDA.n80 GNDA.n4 9.3005
R340 GNDA.n33 GNDA.n32 9.3005
R341 GNDA.n34 GNDA.n20 9.3005
R342 GNDA.n63 GNDA.n62 9.3005
R343 GNDA.n61 GNDA.n21 9.3005
R344 GNDA.n60 GNDA.n59 9.3005
R345 GNDA.n58 GNDA.n35 9.3005
R346 GNDA.n56 GNDA.n55 9.3005
R347 GNDA.n54 GNDA.n37 9.3005
R348 GNDA.n53 GNDA.n52 9.3005
R349 GNDA.n51 GNDA.n38 9.3005
R350 GNDA.n49 GNDA.n48 9.3005
R351 GNDA.n47 GNDA.n40 9.3005
R352 GNDA.n46 GNDA.n45 9.3005
R353 GNDA.n44 GNDA.n41 9.3005
R354 GNDA.n6 GNDA.n5 9.3005
R355 GNDA.n79 GNDA.n78 9.3005
R356 GNDA.n78 GNDA.n77 6.4005
R357 GNDA.n14 GNDA.n13 4.88834
R358 GNDA.n67 GNDA.n66 4.88834
R359 GNDA.n87 GNDA.n86 0.421712
R360 GNDA.n32 GNDA.n20 0.15675
R361 GNDA.n63 GNDA.n21 0.15675
R362 GNDA.n59 GNDA.n21 0.15675
R363 GNDA.n59 GNDA.n58 0.15675
R364 GNDA.n56 GNDA.n37 0.15675
R365 GNDA.n52 GNDA.n37 0.15675
R366 GNDA.n52 GNDA.n51 0.15675
R367 GNDA.n49 GNDA.n40 0.15675
R368 GNDA.n45 GNDA.n40 0.15675
R369 GNDA.n45 GNDA.n44 0.15675
R370 GNDA.n79 GNDA.n5 0.15675
R371 GNDA.n80 GNDA.n79 0.15675
R372 GNDA.n81 GNDA.n80 0.15675
R373 GNDA.n85 GNDA.n84 0.15675
R374 GNDA.n31 GNDA.n30 0.131895
R375 GNDA.n64 GNDA.n20 0.09425
R376 GNDA.n58 GNDA.n57 0.09425
R377 GNDA.n51 GNDA.n50 0.09425
R378 GNDA.n44 GNDA.n43 0.09425
R379 GNDA.n81 GNDA.n3 0.09425
R380 GNDA.n86 GNDA.n85 0.09425
R381 GNDA.n32 GNDA.n31 0.063
R382 GNDA.n64 GNDA.n63 0.063
R383 GNDA.n57 GNDA.n56 0.063
R384 GNDA.n50 GNDA.n49 0.063
R385 GNDA.n43 GNDA.n5 0.063
R386 GNDA.n84 GNDA.n3 0.063
R387 a_7340_3850.t1 a_7340_3850.n6 1112.76
R388 a_7340_3850.n3 a_7340_3850.n2 416.863
R389 a_7340_3850.n2 a_7340_3850.n0 366.848
R390 a_7340_3850.n2 a_7340_3850.n1 271.401
R391 a_7340_3850.n3 a_7340_3850.t8 208.868
R392 a_7340_3850.n4 a_7340_3850.t7 208.868
R393 a_7340_3850.n5 a_7340_3850.t6 208.868
R394 a_7340_3850.n6 a_7340_3850.t5 208.868
R395 a_7340_3850.n6 a_7340_3850.n5 208.868
R396 a_7340_3850.n5 a_7340_3850.n4 208.868
R397 a_7340_3850.n4 a_7340_3850.n3 193.804
R398 a_7340_3850.n1 a_7340_3850.t4 60.0005
R399 a_7340_3850.n1 a_7340_3850.t3 60.0005
R400 a_7340_3850.n0 a_7340_3850.t0 49.2505
R401 a_7340_3850.n0 a_7340_3850.t2 49.2505
R402 VOUT.n2 VOUT.n1 424.447
R403 VOUT.n2 VOUT.n0 354.046
R404 VOUT.n7 VOUT.n6 313
R405 VOUT.n7 VOUT.n5 242.601
R406 VOUT.n3 VOUT.n2 220.8
R407 VOUT.n8 VOUT.n7 220.8
R408 VOUT VOUT.n3 70.4005
R409 VOUT.n8 VOUT.t8 70.0829
R410 VOUT.n3 VOUT.t9 63.6829
R411 VOUT.n6 VOUT.t5 60.0005
R412 VOUT.n6 VOUT.t4 60.0005
R413 VOUT.n5 VOUT.t7 60.0005
R414 VOUT.n5 VOUT.t6 60.0005
R415 VOUT.n9 VOUT.n8 54.4005
R416 VOUT.n0 VOUT.t3 49.2505
R417 VOUT.n0 VOUT.t2 49.2505
R418 VOUT.n1 VOUT.t0 49.2505
R419 VOUT.n1 VOUT.t1 49.2505
R420 VOUT VOUT.n9 12.8005
R421 VOUT.n9 VOUT.n4 6.4005
R422 p_bias p_bias.t0 918.318
R423 p_bias p_bias.n11 540.801
R424 p_bias.n8 p_bias.t10 377.567
R425 p_bias.n3 p_bias.t9 377.567
R426 p_bias.n9 p_bias.n8 257.067
R427 p_bias.n7 p_bias.n6 257.067
R428 p_bias.n4 p_bias.n3 257.067
R429 p_bias.n11 p_bias.n0 154.321
R430 p_bias.n2 p_bias.n1 154.321
R431 p_bias.n5 p_bias.n2 152
R432 p_bias.n11 p_bias.n10 152
R433 p_bias.n8 p_bias.t12 120.501
R434 p_bias.n9 p_bias.t5 120.501
R435 p_bias.n7 p_bias.t1 120.501
R436 p_bias.n6 p_bias.t3 120.501
R437 p_bias.n3 p_bias.t11 120.501
R438 p_bias.n4 p_bias.t7 120.501
R439 p_bias.n11 p_bias.n2 115.201
R440 p_bias.n10 p_bias.n9 85.6894
R441 p_bias.n10 p_bias.n7 85.6894
R442 p_bias.n6 p_bias.n5 85.6894
R443 p_bias.n5 p_bias.n4 85.6894
R444 p_bias.n0 p_bias.t2 19.7005
R445 p_bias.n0 p_bias.t6 19.7005
R446 p_bias.n1 p_bias.t8 19.7005
R447 p_bias.n1 p_bias.t4 19.7005
R448 VIN-.n2 VIN-.n1 2008.33
R449 VIN- VIN-.n2 618.567
R450 VIN-.n0 VIN-.t2 401.668
R451 VIN-.n2 VIN-.n0 369.534
R452 VIN-.n1 VIN-.t0 321.334
R453 VIN-.n0 VIN-.t3 192.8
R454 VIN-.n1 VIN-.t1 112.468
R455 a_7170_3160.n7 a_7170_3160.n5 482.582
R456 a_7170_3160.n3 a_7170_3160.t8 304.634
R457 a_7170_3160.n0 a_7170_3160.t11 304.634
R458 a_7170_3160.n3 a_7170_3160.t10 277.914
R459 a_7170_3160.t12 a_7170_3160.n0 276.289
R460 a_7170_3160.n8 a_7170_3160.n1 204.201
R461 a_7170_3160.n4 a_7170_3160.n2 204.201
R462 a_7170_3160.n10 a_7170_3160.n9 204.201
R463 a_7170_3160.n7 a_7170_3160.n6 120.981
R464 a_7170_3160.n8 a_7170_3160.n4 74.6672
R465 a_7170_3160.n9 a_7170_3160.n8 74.6672
R466 a_7170_3160.n1 a_7170_3160.t5 60.0005
R467 a_7170_3160.n1 a_7170_3160.t1 60.0005
R468 a_7170_3160.n2 a_7170_3160.t0 60.0005
R469 a_7170_3160.n2 a_7170_3160.t9 60.0005
R470 a_7170_3160.t12 a_7170_3160.n10 60.0005
R471 a_7170_3160.n10 a_7170_3160.t4 60.0005
R472 a_7170_3160.n8 a_7170_3160.n7 37.763
R473 a_7170_3160.n5 a_7170_3160.t6 24.0005
R474 a_7170_3160.n5 a_7170_3160.t3 24.0005
R475 a_7170_3160.n6 a_7170_3160.t2 24.0005
R476 a_7170_3160.n6 a_7170_3160.t7 24.0005
R477 a_7170_3160.n4 a_7170_3160.n3 16.0005
R478 a_7170_3160.n9 a_7170_3160.n0 16.0005
R479 a_7070_3110.n4 a_7070_3110.t10 317.317
R480 a_7070_3110.n2 a_7070_3110.t9 317.317
R481 a_7070_3110.n5 a_7070_3110.n4 257.067
R482 a_7070_3110.n3 a_7070_3110.n2 257.067
R483 a_7070_3110.n10 a_7070_3110.n9 257.067
R484 a_7070_3110.t0 a_7070_3110.n12 194.478
R485 a_7070_3110.n8 a_7070_3110.n7 152
R486 a_7070_3110.n12 a_7070_3110.n11 152
R487 a_7070_3110.n1 a_7070_3110.n0 120.981
R488 a_7070_3110.n7 a_7070_3110.n6 117.781
R489 a_7070_3110.n7 a_7070_3110.n1 108.8
R490 a_7070_3110.n8 a_7070_3110.n5 85.6894
R491 a_7070_3110.n11 a_7070_3110.n3 85.6894
R492 a_7070_3110.n11 a_7070_3110.n10 85.6894
R493 a_7070_3110.n9 a_7070_3110.n8 85.6894
R494 a_7070_3110.n4 a_7070_3110.t12 60.2505
R495 a_7070_3110.n5 a_7070_3110.t5 60.2505
R496 a_7070_3110.n2 a_7070_3110.t11 60.2505
R497 a_7070_3110.n3 a_7070_3110.t7 60.2505
R498 a_7070_3110.n10 a_7070_3110.t3 60.2505
R499 a_7070_3110.n9 a_7070_3110.t1 60.2505
R500 a_7070_3110.n6 a_7070_3110.t2 24.0005
R501 a_7070_3110.n6 a_7070_3110.t6 24.0005
R502 a_7070_3110.n0 a_7070_3110.t8 24.0005
R503 a_7070_3110.n0 a_7070_3110.t4 24.0005
R504 a_7070_3110.n12 a_7070_3110.n1 3.2005
R505 a_6820_4420.n8 a_6820_4420.n6 522.322
R506 a_6820_4420.n3 a_6820_4420.t8 384.967
R507 a_6820_4420.n0 a_6820_4420.t11 384.967
R508 a_6820_4420.n3 a_6820_4420.t10 379.166
R509 a_6820_4420.t12 a_6820_4420.n0 376.56
R510 a_6820_4420.n4 a_6820_4420.n2 315.647
R511 a_6820_4420.n5 a_6820_4420.n1 315.647
R512 a_6820_4420.n11 a_6820_4420.n10 314.503
R513 a_6820_4420.n8 a_6820_4420.n7 160.721
R514 a_6820_4420.n5 a_6820_4420.n4 83.2005
R515 a_6820_4420.n2 a_6820_4420.t0 49.2505
R516 a_6820_4420.n2 a_6820_4420.t9 49.2505
R517 a_6820_4420.n1 a_6820_4420.t3 49.2505
R518 a_6820_4420.n1 a_6820_4420.t1 49.2505
R519 a_6820_4420.t12 a_6820_4420.n11 49.2505
R520 a_6820_4420.n11 a_6820_4420.t2 49.2505
R521 a_6820_4420.n10 a_6820_4420.n9 42.6672
R522 a_6820_4420.n9 a_6820_4420.n8 37.763
R523 a_6820_4420.n9 a_6820_4420.n5 23.4672
R524 a_6820_4420.n6 a_6820_4420.t7 19.7005
R525 a_6820_4420.n6 a_6820_4420.t5 19.7005
R526 a_6820_4420.n7 a_6820_4420.t4 19.7005
R527 a_6820_4420.n7 a_6820_4420.t6 19.7005
R528 a_6820_4420.n4 a_6820_4420.n3 16.0005
R529 a_6820_4420.n10 a_6820_4420.n0 16.0005
R530 VIN+.n0 VIN+.t1 377.567
R531 VIN+.n1 VIN+.t2 297.233
R532 VIN+.n2 VIN+.n1 243.44
R533 VIN+.n2 VIN+.n0 224.496
R534 VIN+.n0 VIN+.t0 216.9
R535 VIN+.n1 VIN+.t3 136.567
R536 VIN+ VIN+.n2 3.438
R537 n_right.t0 n_right.n6 1010.36
R538 n_right.n3 n_right.n2 416.101
R539 n_right.n2 n_right.n0 354.046
R540 n_right.n6 n_right.t8 289.2
R541 n_right.n5 n_right.t5 289.2
R542 n_right.n4 n_right.t6 289.2
R543 n_right.n3 n_right.t7 289.2
R544 n_right.n2 n_right.n1 284.2
R545 n_right.n6 n_right.n5 208.868
R546 n_right.n5 n_right.n4 208.868
R547 n_right.n4 n_right.n3 208.868
R548 n_right.n1 n_right.t2 60.0005
R549 n_right.n1 n_right.t1 60.0005
R550 n_right.n0 n_right.t4 49.2505
R551 n_right.n0 n_right.t3 49.2505
R552 a_10210_2370.t0 a_10210_2370.t1 245.883
R553 a_10210_5296.t0 a_10210_5296.t1 323.964
C0 VIN+ VIN- 0.126393f
C1 VIN+ VDDA 0.256632f
C2 VOUT VDDA 0.469696f
C3 VIN- VDDA 0.171402f
C4 VIN- p_bias 0.010861f
C5 p_bias VDDA 2.78755f
C6 VOUT GNDA 1.46613f
C7 VIN+ GNDA 0.962537f
C8 VIN- GNDA 1.24201f
C9 VDDA GNDA 13.276419f
C10 p_bias GNDA 3.947242f
C11 a_6820_4420.t11 GNDA 0.030769f
C12 a_6820_4420.n0 GNDA 0.124795f
C13 a_6820_4420.t3 GNDA 0.020325f
C14 a_6820_4420.t1 GNDA 0.020325f
C15 a_6820_4420.n1 GNDA 0.044943f
C16 a_6820_4420.t0 GNDA 0.020325f
C17 a_6820_4420.t9 GNDA 0.020325f
C18 a_6820_4420.n2 GNDA 0.044943f
C19 a_6820_4420.t10 GNDA 0.077457f
C20 a_6820_4420.t8 GNDA 0.030769f
C21 a_6820_4420.n3 GNDA 0.097952f
C22 a_6820_4420.n4 GNDA 0.087903f
C23 a_6820_4420.n5 GNDA 0.089425f
C24 a_6820_4420.t7 GNDA 0.050813f
C25 a_6820_4420.t5 GNDA 0.050813f
C26 a_6820_4420.n6 GNDA 0.295523f
C27 a_6820_4420.t4 GNDA 0.050813f
C28 a_6820_4420.t6 GNDA 0.050813f
C29 a_6820_4420.n7 GNDA 0.144587f
C30 a_6820_4420.n8 GNDA 0.360746f
C31 a_6820_4420.n9 GNDA 0.13437f
C32 a_6820_4420.n10 GNDA 0.085474f
C33 a_6820_4420.t2 GNDA 0.020325f
C34 a_6820_4420.n11 GNDA 0.045257f
C35 a_6820_4420.t12 GNDA 0.100208f
C36 p_bias.t2 GNDA 0.019014f
C37 p_bias.t6 GNDA 0.019014f
C38 p_bias.n0 GNDA 0.052203f
C39 p_bias.t8 GNDA 0.019014f
C40 p_bias.t4 GNDA 0.019014f
C41 p_bias.n1 GNDA 0.052203f
C42 p_bias.n2 GNDA 0.06614f
C43 p_bias.t1 GNDA 0.052478f
C44 p_bias.t3 GNDA 0.052478f
C45 p_bias.t7 GNDA 0.052478f
C46 p_bias.t11 GNDA 0.052478f
C47 p_bias.t9 GNDA 0.072156f
C48 p_bias.n3 GNDA 0.040407f
C49 p_bias.n4 GNDA 0.028673f
C50 p_bias.n5 GNDA 0.012321f
C51 p_bias.n6 GNDA 0.028673f
C52 p_bias.n7 GNDA 0.028673f
C53 p_bias.t5 GNDA 0.052478f
C54 p_bias.t12 GNDA 0.052478f
C55 p_bias.t10 GNDA 0.072156f
C56 p_bias.n8 GNDA 0.040407f
C57 p_bias.n9 GNDA 0.028673f
C58 p_bias.n10 GNDA 0.012321f
C59 p_bias.n11 GNDA 0.116466f
C60 p_bias.t0 GNDA 1.60533f
C61 VDDA.n2 GNDA 0.013168f
C62 VDDA.n3 GNDA 0.027433f
C63 VDDA.t0 GNDA 0.079061f
C64 VDDA.n9 GNDA 0.091281f
C65 VDDA.t37 GNDA 0.016775f
C66 VDDA.t39 GNDA 0.141352f
C67 VDDA.t18 GNDA 0.124581f
C68 VDDA.t3 GNDA 0.124581f
C69 VDDA.t21 GNDA 0.124581f
C70 VDDA.t56 GNDA 0.124581f
C71 VDDA.t36 GNDA 0.246253f
C72 VDDA.n15 GNDA 0.100543f
C73 VDDA.n16 GNDA 0.010064f
C74 VDDA.n17 GNDA 0.015819f
C75 VDDA.t41 GNDA 0.01311f
C76 VDDA.n19 GNDA 0.027517f
C77 VDDA.n21 GNDA 0.015819f
C78 VDDA.n22 GNDA 0.022642f
C79 VDDA.n23 GNDA 0.065783f
C80 VDDA.n25 GNDA 0.01915f
C81 VDDA.n26 GNDA 0.064099f
C82 VDDA.n30 GNDA 0.01915f
C83 VDDA.n31 GNDA 0.064099f
C84 VDDA.n34 GNDA 0.01915f
C85 VDDA.n35 GNDA 0.064099f
C86 VDDA.n37 GNDA 0.01915f
C87 VDDA.n38 GNDA 0.064099f
C88 VDDA.n66 GNDA 0.066097f
C89 VDDA.n67 GNDA 0.01915f
C90 VDDA.t44 GNDA 0.018289f
C91 VDDA.n68 GNDA 0.027433f
C92 VDDA.t42 GNDA 0.036978f
C93 VDDA.n69 GNDA 0.025838f
C94 VDDA.n72 GNDA 0.013168f
C95 VDDA.n73 GNDA 0.013168f
C96 VDDA.n75 GNDA 0.013168f
C97 VDDA.n76 GNDA 0.01329f
C98 VDDA.n78 GNDA 0.076665f
C99 VDDA.t46 GNDA 0.079061f
C100 VDDA.t31 GNDA 0.079061f
C101 VDDA.t14 GNDA 0.062291f
C102 VDDA.t33 GNDA 0.095832f
C103 VDDA.t9 GNDA 0.062291f
C104 VDDA.t27 GNDA 0.07427f
C105 VDDA.t29 GNDA 0.083853f
C106 VDDA.t23 GNDA 0.062291f
C107 VDDA.t50 GNDA 0.095832f
C108 VDDA.t43 GNDA 0.079061f
C109 VDDA.n79 GNDA 0.103272f
C110 VDDA.t51 GNDA 0.016775f
C111 VDDA.n80 GNDA 0.032694f
C112 VDDA.n81 GNDA 0.010064f
C113 VDDA.n82 GNDA 0.015819f
C114 VDDA.n83 GNDA 0.020442f
C115 VDDA.n84 GNDA 0.015819f
C116 VDDA.t48 GNDA 0.01311f
C117 VDDA.n86 GNDA 0.027517f
C118 VDDA.n87 GNDA 0.10326f
C119 VDDA.t16 GNDA 0.129373f
C120 VDDA.t7 GNDA 0.122185f
C121 VDDA.t26 GNDA 0.088644f
C122 VDDA.t11 GNDA 0.069478f
C123 VDDA.t12 GNDA 0.062291f
C124 VDDA.t25 GNDA 0.095832f
C125 VDDA.t5 GNDA 0.062291f
C126 VDDA.t20 GNDA 0.083853f
C127 VDDA.t2 GNDA 0.07427f
C128 VDDA.t53 GNDA 0.062291f
C129 VDDA.t58 GNDA 0.095832f
C130 VDDA.n90 GNDA 0.013089f
C131 VDDA.n91 GNDA 0.013168f
C132 VDDA.n93 GNDA 0.013168f
C133 VDDA.n96 GNDA 0.198851f
C134 VDDA.n98 GNDA 0.012531f
C135 VDDA.t52 GNDA 0.036236f
C136 VDDA.n99 GNDA 0.012784f
C137 VDDA.n100 GNDA 0.018616f
C138 VDDA.n101 GNDA 0.024948f
.ends

