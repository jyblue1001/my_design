magic
tech sky130A
timestamp 1739812747
<< psubdiff >>
rect 2605 195 2655 210
rect 2605 175 2620 195
rect 2640 175 2655 195
rect 2605 160 2655 175
<< psubdiffcont >>
rect 2620 175 2640 195
<< xpolycontact >>
rect 5520 295 5740 330
rect 6476 295 6696 330
<< xpolyres >>
rect 5740 295 6476 330
<< locali >>
rect 1135 320 1185 330
rect 1135 290 1145 320
rect 1175 290 1185 320
rect 5480 325 5520 330
rect 5480 300 5485 325
rect 5510 300 5520 325
rect 5480 295 5520 300
rect 6696 325 6736 330
rect 6696 300 6706 325
rect 6731 300 6736 325
rect 6696 295 6736 300
rect 1135 280 1185 290
rect 2475 220 2780 230
rect 2475 185 2485 220
rect 2520 210 2735 220
rect 2520 185 2530 210
rect 2475 175 2530 185
rect 2605 195 2655 210
rect 2605 175 2620 195
rect 2640 175 2655 195
rect 2725 185 2735 210
rect 2770 185 2780 220
rect 2725 175 2780 185
rect 2605 160 2655 175
<< viali >>
rect 1145 290 1175 320
rect 5485 300 5510 325
rect 6706 300 6731 325
rect 2485 185 2520 220
rect 2735 185 2770 220
<< metal1 >>
rect 1135 325 5520 330
rect 1135 320 5485 325
rect 1135 290 1145 320
rect 1175 300 5485 320
rect 5510 300 5520 325
rect 1175 295 5520 300
rect 6695 325 9720 330
rect 6695 300 6706 325
rect 6731 320 9720 325
rect 6731 300 9680 320
rect 6695 295 9680 300
rect 1175 290 1185 295
rect 1135 280 1185 290
rect 9670 290 9680 295
rect 9710 290 9720 320
rect 9670 280 9720 290
rect 2475 220 2530 230
rect 2475 185 2485 220
rect 2520 185 2530 220
rect 2475 175 2530 185
rect 2725 220 2780 230
rect 2725 185 2735 220
rect 2770 185 2780 220
rect 2725 175 2780 185
<< via1 >>
rect 1145 290 1175 320
rect 9680 290 9710 320
rect 2485 185 2520 220
rect 2735 185 2770 220
<< metal2 >>
rect 1135 320 1185 330
rect 1135 290 1145 320
rect 1175 290 1185 320
rect 1135 280 1185 290
rect 9670 320 9720 330
rect 9670 290 9680 320
rect 9710 290 9720 320
rect 9670 280 9720 290
rect 2475 220 2530 230
rect 2475 185 2485 220
rect 2520 185 2530 220
rect 2475 175 2530 185
rect 2725 220 2780 230
rect 2725 185 2735 220
rect 2770 185 2780 220
rect 2725 175 2780 185
<< via2 >>
rect 1145 290 1175 320
rect 9680 290 9710 320
rect 2485 185 2520 220
rect 2735 185 2770 220
<< metal3 >>
rect 1135 320 1185 330
rect 1135 290 1145 320
rect 1175 290 1185 320
rect 1135 55 1185 290
rect 9670 320 9720 330
rect 9670 290 9680 320
rect 9710 290 9720 320
rect 2475 220 2530 230
rect 2475 185 2485 220
rect 2520 185 2530 220
rect 2475 175 2530 185
rect 2725 220 2780 230
rect 2725 185 2735 220
rect 2770 185 2780 220
rect 2725 175 2780 185
rect 9670 55 9720 290
rect 1135 -5975 2545 55
rect 2710 -5975 9720 55
<< via3 >>
rect 2485 185 2520 220
rect 2735 185 2770 220
<< mimcap >>
rect 1150 30 2530 40
rect 1150 -5 2485 30
rect 2520 -5 2530 30
rect 1150 -5960 2530 -5
rect 2725 30 9705 40
rect 2725 -5 2735 30
rect 2770 -5 9705 30
rect 2725 -5960 9705 -5
<< mimcapcontact >>
rect 2485 -5 2520 30
rect 2735 -5 2770 30
<< metal4 >>
rect 2475 220 2530 230
rect 2475 185 2485 220
rect 2520 185 2530 220
rect 2475 30 2530 185
rect 2475 -5 2485 30
rect 2520 -5 2530 30
rect 2475 -10 2530 -5
rect 2725 220 2780 230
rect 2725 185 2735 220
rect 2770 185 2780 220
rect 2725 30 2780 185
rect 2725 -5 2735 30
rect 2770 -5 2780 30
rect 2725 -10 2780 -5
<< labels >>
flabel metal1 1485 330 1485 330 1 FreeSans 800 0 0 400 V_OUT
port 1 n
flabel metal1 8230 330 8230 330 1 FreeSans 800 0 0 400 R1_C1
flabel locali 2630 160 2630 160 5 FreeSans 800 0 0 -400 GNDA
<< end >>
