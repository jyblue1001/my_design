* PEX produced on Sat Jul  5 05:14:37 PM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 VDDA.t315 bgr_0.V_TOP.t14 bgr_0.Vin-.t4 VDDA.t314 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X1 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 GNDA.t216 GNDA.t215 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X2 bgr_0.1st_Vout_1.t11 bgr_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X3 bgr_0.V_TOP.t15 VDDA.t313 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X4 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA.t314 GNDA.t316 GNDA.t315 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X5 two_stage_opamp_dummy_magic_0.VOUT+.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X6 GNDA.t248 GNDA.t313 bgr_0.Vbe2.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 two_stage_opamp_dummy_magic_0.Y.t25 GNDA.t47 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X8 two_stage_opamp_dummy_magic_0.VOUT+.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 two_stage_opamp_dummy_magic_0.VOUT+.t21 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 bgr_0.NFET_GATE_10uA.t1 bgr_0.NFET_GATE_10uA.t0 GNDA.t44 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X11 bgr_0.1st_Vout_1.t12 bgr_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 bgr_0.V_TOP.t16 VDDA.t312 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X13 VDDA.t202 bgr_0.V_mir2.t10 bgr_0.V_mir2.t11 VDDA.t201 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X14 two_stage_opamp_dummy_magic_0.V_err_gate.t6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 VDDA.t262 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X15 two_stage_opamp_dummy_magic_0.VOUT+.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X16 two_stage_opamp_dummy_magic_0.VOUT+.t23 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 two_stage_opamp_dummy_magic_0.Y.t8 two_stage_opamp_dummy_magic_0.Vb2.t11 two_stage_opamp_dummy_magic_0.VD4.t20 two_stage_opamp_dummy_magic_0.VD4.t19 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X18 VDDA.t47 two_stage_opamp_dummy_magic_0.X.t25 two_stage_opamp_dummy_magic_0.VOUT-.t13 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X19 two_stage_opamp_dummy_magic_0.Y.t11 two_stage_opamp_dummy_magic_0.Vb1.t6 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA.t126 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X20 two_stage_opamp_dummy_magic_0.VOUT+.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X21 two_stage_opamp_dummy_magic_0.VOUT+.t25 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 VDDA.t42 two_stage_opamp_dummy_magic_0.X.t26 two_stage_opamp_dummy_magic_0.VOUT-.t12 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X23 VDDA.t145 bgr_0.PFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X24 two_stage_opamp_dummy_magic_0.VOUT+.t26 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X25 two_stage_opamp_dummy_magic_0.VOUT-.t18 GNDA.t310 GNDA.t312 GNDA.t311 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X26 a_14520_5068.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA.t91 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X27 bgr_0.V_TOP.t17 VDDA.t311 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X28 VDDA.t65 two_stage_opamp_dummy_magic_0.V_err_gate.t14 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X29 VDDA.t29 bgr_0.V_mir1.t17 bgr_0.1st_Vout_1.t4 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X30 two_stage_opamp_dummy_magic_0.VOUT-.t19 two_stage_opamp_dummy_magic_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X31 bgr_0.START_UP_NFET1.t0 bgr_0.START_UP_NFET1 GNDA.t8 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X32 two_stage_opamp_dummy_magic_0.VOUT-.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X33 two_stage_opamp_dummy_magic_0.VOUT-.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 two_stage_opamp_dummy_magic_0.VOUT+.t27 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 two_stage_opamp_dummy_magic_0.VOUT+.t28 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 two_stage_opamp_dummy_magic_0.VOUT+.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 two_stage_opamp_dummy_magic_0.VOUT-.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 bgr_0.1st_Vout_1.t13 bgr_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 two_stage_opamp_dummy_magic_0.V_p_mir.t3 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 GNDA.t18 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X40 two_stage_opamp_dummy_magic_0.VOUT+.t16 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA.t322 GNDA.t321 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X41 VDDA.t14 two_stage_opamp_dummy_magic_0.Y.t26 two_stage_opamp_dummy_magic_0.VOUT+.t1 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X42 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 two_stage_opamp_dummy_magic_0.X.t27 VDDA.t130 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X43 two_stage_opamp_dummy_magic_0.VOUT+.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 bgr_0.V_mir2.t16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 bgr_0.V_p_2.t5 GNDA.t182 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X45 bgr_0.Vin-.t6 bgr_0.V_TOP.t18 VDDA.t310 VDDA.t309 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X46 VDDA.t430 VDDA.t428 two_stage_opamp_dummy_magic_0.V_err_gate.t12 VDDA.t429 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X47 GNDA.t176 bgr_0.NFET_GATE_10uA.t5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA.t175 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X48 GNDA.t38 bgr_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X49 two_stage_opamp_dummy_magic_0.V_err_p.t19 two_stage_opamp_dummy_magic_0.V_err_gate.t15 VDDA.t67 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X50 two_stage_opamp_dummy_magic_0.VOUT+.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 two_stage_opamp_dummy_magic_0.VOUT-.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X52 two_stage_opamp_dummy_magic_0.Y.t2 two_stage_opamp_dummy_magic_0.Vb2.t12 two_stage_opamp_dummy_magic_0.VD4.t18 two_stage_opamp_dummy_magic_0.VD4.t17 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X53 two_stage_opamp_dummy_magic_0.V_err_p.t0 two_stage_opamp_dummy_magic_0.V_tot.t4 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X54 two_stage_opamp_dummy_magic_0.X.t11 two_stage_opamp_dummy_magic_0.Vb1.t7 two_stage_opamp_dummy_magic_0.VD1.t20 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X55 two_stage_opamp_dummy_magic_0.VOUT-.t24 two_stage_opamp_dummy_magic_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 two_stage_opamp_dummy_magic_0.X.t28 GNDA.t21 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X57 bgr_0.1st_Vout_1.t3 bgr_0.Vin+.t6 bgr_0.V_p_1.t4 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X58 two_stage_opamp_dummy_magic_0.VOUT-.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 bgr_0.1st_Vout_2.t11 bgr_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X60 GNDA.t327 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_0.V_source.t38 GNDA.t326 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X61 VDDA.t427 VDDA.t425 bgr_0.V_TOP.t2 VDDA.t426 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X62 GNDA.t158 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 two_stage_opamp_dummy_magic_0.V_source.t37 GNDA.t157 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X63 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 two_stage_opamp_dummy_magic_0.Y.t27 VDDA.t15 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X64 two_stage_opamp_dummy_magic_0.VD1.t3 VIN-.t0 two_stage_opamp_dummy_magic_0.V_source.t8 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X65 two_stage_opamp_dummy_magic_0.V_err_p.t18 two_stage_opamp_dummy_magic_0.V_err_gate.t16 VDDA.t23 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X66 two_stage_opamp_dummy_magic_0.VOUT-.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X67 GNDA.t40 bgr_0.NFET_GATE_10uA.t7 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X68 GNDA.t309 GNDA.t307 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA.t308 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X69 VDDA.t179 bgr_0.V_mir1.t18 bgr_0.1st_Vout_1.t8 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X70 two_stage_opamp_dummy_magic_0.VOUT+.t32 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X71 two_stage_opamp_dummy_magic_0.VOUT-.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 two_stage_opamp_dummy_magic_0.err_amp_out.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 GNDA.t214 GNDA.t213 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X73 two_stage_opamp_dummy_magic_0.VOUT-.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X74 two_stage_opamp_dummy_magic_0.VOUT-.t29 two_stage_opamp_dummy_magic_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X75 two_stage_opamp_dummy_magic_0.VOUT+.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 two_stage_opamp_dummy_magic_0.VD1.t0 VIN-.t1 two_stage_opamp_dummy_magic_0.V_source.t2 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X77 two_stage_opamp_dummy_magic_0.VOUT-.t30 two_stage_opamp_dummy_magic_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X78 bgr_0.NFET_GATE_10uA.t4 bgr_0.PFET_GATE_10uA.t11 VDDA.t448 VDDA.t447 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X79 two_stage_opamp_dummy_magic_0.err_amp_out.t9 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 GNDA.t212 GNDA.t211 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X80 bgr_0.1st_Vout_2.t12 bgr_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 VDDA.t31 bgr_0.PFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 VDDA.t30 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X82 GNDA.t306 GNDA.t304 two_stage_opamp_dummy_magic_0.X.t20 GNDA.t305 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X83 two_stage_opamp_dummy_magic_0.VOUT+.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VDDA.t424 VDDA.t422 bgr_0.NFET_GATE_10uA.t2 VDDA.t423 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X85 two_stage_opamp_dummy_magic_0.Y.t20 GNDA.t301 GNDA.t303 GNDA.t302 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X86 VDDA.t115 two_stage_opamp_dummy_magic_0.X.t29 two_stage_opamp_dummy_magic_0.VOUT-.t11 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X87 VDDA.t442 bgr_0.1st_Vout_1.t14 bgr_0.V_TOP.t11 VDDA.t441 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X88 GNDA.t300 GNDA.t298 two_stage_opamp_dummy_magic_0.VD1.t8 GNDA.t299 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X89 two_stage_opamp_dummy_magic_0.VOUT-.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 two_stage_opamp_dummy_magic_0.VD3.t36 VDDA.t419 VDDA.t421 VDDA.t420 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X91 two_stage_opamp_dummy_magic_0.VOUT-.t32 two_stage_opamp_dummy_magic_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X92 two_stage_opamp_dummy_magic_0.VOUT-.t0 a_14240_2076.t0 GNDA.t6 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X93 two_stage_opamp_dummy_magic_0.VOUT+.t35 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 two_stage_opamp_dummy_magic_0.VOUT-.t33 two_stage_opamp_dummy_magic_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 VDDA.t462 bgr_0.V_mir2.t8 bgr_0.V_mir2.t9 VDDA.t461 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X96 two_stage_opamp_dummy_magic_0.VD3.t30 two_stage_opamp_dummy_magic_0.VD3.t28 two_stage_opamp_dummy_magic_0.X.t18 two_stage_opamp_dummy_magic_0.VD3.t29 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X97 GNDA.t122 bgr_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X98 VDDA.t25 two_stage_opamp_dummy_magic_0.V_err_gate.t17 two_stage_opamp_dummy_magic_0.V_err_p.t17 VDDA.t24 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X99 two_stage_opamp_dummy_magic_0.VOUT+.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 two_stage_opamp_dummy_magic_0.Vb3.t4 bgr_0.NFET_GATE_10uA.t9 GNDA.t124 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X101 GNDA.t297 GNDA.t295 two_stage_opamp_dummy_magic_0.VD1.t7 GNDA.t296 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X102 VDDA.t440 bgr_0.1st_Vout_1.t15 bgr_0.V_TOP.t10 VDDA.t439 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X103 two_stage_opamp_dummy_magic_0.VOUT-.t34 two_stage_opamp_dummy_magic_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 bgr_0.V_TOP.t3 bgr_0.cap_res1.t0 GNDA.t96 sky130_fd_pr__res_high_po_0p35 l=2.05
X105 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 two_stage_opamp_dummy_magic_0.X.t30 VDDA.t102 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X106 two_stage_opamp_dummy_magic_0.V_source.t36 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA.t220 GNDA.t219 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X107 a_11220_17410.t0 GNDA.t90 GNDA.t23 sky130_fd_pr__res_xhigh_po_0p35 l=6
X108 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 two_stage_opamp_dummy_magic_0.X.t31 VDDA.t58 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X109 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 two_stage_opamp_dummy_magic_0.V_err_gate.t18 VDDA.t93 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X110 two_stage_opamp_dummy_magic_0.VOUT+.t37 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 two_stage_opamp_dummy_magic_0.Vb1.t0 bgr_0.PFET_GATE_10uA.t13 VDDA.t72 VDDA.t71 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X112 two_stage_opamp_dummy_magic_0.VOUT-.t35 two_stage_opamp_dummy_magic_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 bgr_0.PFET_GATE_10uA.t9 bgr_0.1st_Vout_2.t13 VDDA.t466 VDDA.t465 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X114 two_stage_opamp_dummy_magic_0.VOUT-.t36 two_stage_opamp_dummy_magic_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 GNDA.t138 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_0.V_source.t35 GNDA.t137 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X116 two_stage_opamp_dummy_magic_0.VD3.t37 two_stage_opamp_dummy_magic_0.Vb3.t8 VDDA.t450 VDDA.t449 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X117 two_stage_opamp_dummy_magic_0.VOUT-.t37 two_stage_opamp_dummy_magic_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X118 two_stage_opamp_dummy_magic_0.VOUT-.t38 two_stage_opamp_dummy_magic_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X119 two_stage_opamp_dummy_magic_0.VOUT-.t39 two_stage_opamp_dummy_magic_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 two_stage_opamp_dummy_magic_0.VOUT+.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 two_stage_opamp_dummy_magic_0.VOUT+.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X122 VDDA.t218 bgr_0.V_mir1.t10 bgr_0.V_mir1.t11 VDDA.t217 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X123 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 two_stage_opamp_dummy_magic_0.Y.t28 VDDA.t254 GNDA.t177 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X124 two_stage_opamp_dummy_magic_0.VOUT+.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 two_stage_opamp_dummy_magic_0.VOUT+.t41 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 GNDA.t210 GNDA.t209 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X127 GNDA.t93 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 two_stage_opamp_dummy_magic_0.VOUT+.t4 GNDA.t92 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X128 two_stage_opamp_dummy_magic_0.VOUT+.t42 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X129 bgr_0.1st_Vout_1.t16 bgr_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X130 VDDA.t61 bgr_0.1st_Vout_2.t14 bgr_0.PFET_GATE_10uA.t2 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X131 two_stage_opamp_dummy_magic_0.VD4.t28 two_stage_opamp_dummy_magic_0.Vb3.t9 VDDA.t261 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X132 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 two_stage_opamp_dummy_magic_0.Y.t29 GNDA.t178 VDDA.t255 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X133 bgr_0.V_TOP.t19 VDDA.t308 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 two_stage_opamp_dummy_magic_0.VD4.t16 two_stage_opamp_dummy_magic_0.Vb2.t13 two_stage_opamp_dummy_magic_0.Y.t3 two_stage_opamp_dummy_magic_0.VD4.t15 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X135 two_stage_opamp_dummy_magic_0.VOUT-.t40 two_stage_opamp_dummy_magic_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 bgr_0.1st_Vout_1.t17 bgr_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X137 two_stage_opamp_dummy_magic_0.VD1.t19 two_stage_opamp_dummy_magic_0.Vb1.t8 two_stage_opamp_dummy_magic_0.X.t17 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X138 two_stage_opamp_dummy_magic_0.VOUT-.t41 two_stage_opamp_dummy_magic_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X139 a_14640_5068.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 GNDA.t70 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X140 two_stage_opamp_dummy_magic_0.Y.t15 two_stage_opamp_dummy_magic_0.Vb1.t9 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X141 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA.t292 GNDA.t294 GNDA.t293 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X142 two_stage_opamp_dummy_magic_0.VOUT-.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 two_stage_opamp_dummy_magic_0.VOUT+.t43 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X144 two_stage_opamp_dummy_magic_0.V_source.t6 VIN+.t0 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X145 two_stage_opamp_dummy_magic_0.VOUT-.t43 two_stage_opamp_dummy_magic_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X146 VDDA.t132 bgr_0.V_mir2.t17 bgr_0.1st_Vout_2.t6 VDDA.t131 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X147 two_stage_opamp_dummy_magic_0.VOUT+.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X148 two_stage_opamp_dummy_magic_0.VOUT+.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 bgr_0.1st_Vout_1.t18 bgr_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 a_13730_17020.t1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X151 GNDA.t104 two_stage_opamp_dummy_magic_0.Y.t30 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X152 two_stage_opamp_dummy_magic_0.V_source.t0 VIN+.t1 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X153 two_stage_opamp_dummy_magic_0.VOUT-.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 bgr_0.V_CUR_REF_REG.t2 VDDA.t416 VDDA.t418 VDDA.t417 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X155 a_11220_17410.t1 a_12828_17530.t1 GNDA.t23 sky130_fd_pr__res_xhigh_po_0p35 l=6
X156 two_stage_opamp_dummy_magic_0.VOUT-.t45 two_stage_opamp_dummy_magic_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 VDDA.t127 two_stage_opamp_dummy_magic_0.Y.t31 two_stage_opamp_dummy_magic_0.VOUT+.t8 VDDA.t126 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X158 two_stage_opamp_dummy_magic_0.VOUT+.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 bgr_0.PFET_GATE_10uA.t14 VDDA.t177 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X160 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 two_stage_opamp_dummy_magic_0.X.t32 VDDA.t83 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X161 two_stage_opamp_dummy_magic_0.VOUT-.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X162 two_stage_opamp_dummy_magic_0.VOUT-.t47 two_stage_opamp_dummy_magic_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 two_stage_opamp_dummy_magic_0.V_source.t39 two_stage_opamp_dummy_magic_0.Vb1.t3 two_stage_opamp_dummy_magic_0.Vb1.t4 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=3.1
X164 two_stage_opamp_dummy_magic_0.V_source.t34 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA.t77 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X165 VDDA.t216 bgr_0.PFET_GATE_10uA.t15 bgr_0.V_CUR_REF_REG.t1 VDDA.t215 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X166 two_stage_opamp_dummy_magic_0.VD3.t20 two_stage_opamp_dummy_magic_0.Vb3.t10 VDDA.t33 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X167 two_stage_opamp_dummy_magic_0.VOUT-.t48 two_stage_opamp_dummy_magic_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 bgr_0.PFET_GATE_10uA.t3 bgr_0.cap_res2.t20 GNDA.t96 sky130_fd_pr__res_high_po_0p35 l=2.05
X169 two_stage_opamp_dummy_magic_0.VD4.t14 two_stage_opamp_dummy_magic_0.Vb2.t14 two_stage_opamp_dummy_magic_0.Y.t4 two_stage_opamp_dummy_magic_0.VD4.t13 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X170 bgr_0.V_p_1.t9 bgr_0.Vin-.t8 bgr_0.V_mir1.t16 GNDA.t187 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X171 VDDA.t80 bgr_0.V_mir1.t8 bgr_0.V_mir1.t9 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X172 two_stage_opamp_dummy_magic_0.VOUT-.t49 two_stage_opamp_dummy_magic_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X173 two_stage_opamp_dummy_magic_0.VOUT-.t50 two_stage_opamp_dummy_magic_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X174 GNDA.t291 GNDA.t289 two_stage_opamp_dummy_magic_0.Y.t19 GNDA.t290 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X175 bgr_0.1st_Vout_2.t15 bgr_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 two_stage_opamp_dummy_magic_0.VOUT+.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 two_stage_opamp_dummy_magic_0.VOUT+.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X178 VDDA.t438 bgr_0.1st_Vout_1.t19 bgr_0.V_TOP.t9 VDDA.t437 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X179 VDDA.t307 bgr_0.V_TOP.t20 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 VDDA.t306 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X180 two_stage_opamp_dummy_magic_0.VOUT+.t49 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X181 GNDA.t218 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_0.V_source.t33 GNDA.t217 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X182 two_stage_opamp_dummy_magic_0.VOUT+.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 bgr_0.V_p_2.t10 bgr_0.V_CUR_REF_REG.t3 bgr_0.1st_Vout_2.t10 GNDA.t320 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X184 two_stage_opamp_dummy_magic_0.VOUT+.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X185 two_stage_opamp_dummy_magic_0.VOUT-.t51 two_stage_opamp_dummy_magic_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X186 two_stage_opamp_dummy_magic_0.VOUT+.t2 two_stage_opamp_dummy_magic_0.Y.t32 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X187 two_stage_opamp_dummy_magic_0.VOUT-.t52 two_stage_opamp_dummy_magic_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 bgr_0.V_p_1.t8 bgr_0.Vin-.t9 bgr_0.V_mir1.t15 GNDA.t186 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X189 bgr_0.1st_Vout_2.t16 bgr_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X190 GNDA.t32 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_0.V_source.t32 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X191 bgr_0.V_TOP.t4 VDDA.t413 VDDA.t415 VDDA.t414 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X192 two_stage_opamp_dummy_magic_0.VOUT+.t52 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X193 bgr_0.Vin-.t7 bgr_0.START_UP.t6 bgr_0.V_TOP.t13 VDDA.t455 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X194 VDDA.t412 VDDA.t410 two_stage_opamp_dummy_magic_0.V_err_p.t21 VDDA.t411 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X195 two_stage_opamp_dummy_magic_0.VD1.t18 two_stage_opamp_dummy_magic_0.Vb1.t10 two_stage_opamp_dummy_magic_0.X.t10 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X196 two_stage_opamp_dummy_magic_0.VOUT+.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 two_stage_opamp_dummy_magic_0.VOUT-.t53 two_stage_opamp_dummy_magic_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X198 bgr_0.1st_Vout_1.t20 bgr_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X199 bgr_0.V_TOP.t21 VDDA.t297 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 two_stage_opamp_dummy_magic_0.err_amp_out.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_0.V_err_p.t9 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X201 two_stage_opamp_dummy_magic_0.VOUT+.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 two_stage_opamp_dummy_magic_0.VOUT+.t55 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 a_14240_2076.t1 GNDA.t154 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X204 VDDA.t70 two_stage_opamp_dummy_magic_0.Vb3.t11 two_stage_opamp_dummy_magic_0.VD3.t21 VDDA.t69 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X205 GNDA.t127 two_stage_opamp_dummy_magic_0.X.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X206 two_stage_opamp_dummy_magic_0.VOUT+.t56 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X207 two_stage_opamp_dummy_magic_0.V_source.t31 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA.t82 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X208 a_13730_17020.t0 GNDA.t4 GNDA.t3 sky130_fd_pr__res_xhigh_po_0p35 l=6.3
X209 bgr_0.1st_Vout_1.t21 bgr_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X210 bgr_0.V_TOP.t22 VDDA.t296 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 two_stage_opamp_dummy_magic_0.VD4.t37 two_stage_opamp_dummy_magic_0.VD4.t35 two_stage_opamp_dummy_magic_0.Y.t7 two_stage_opamp_dummy_magic_0.VD4.t36 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X212 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 VDDA.t407 VDDA.t409 VDDA.t408 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X213 a_11220_17290.t1 a_12828_17650.t1 GNDA.t23 sky130_fd_pr__res_xhigh_po_0p35 l=6
X214 VDDA.t229 two_stage_opamp_dummy_magic_0.Vb3.t12 two_stage_opamp_dummy_magic_0.VD4.t25 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X215 two_stage_opamp_dummy_magic_0.VOUT-.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X216 two_stage_opamp_dummy_magic_0.VOUT-.t55 two_stage_opamp_dummy_magic_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 two_stage_opamp_dummy_magic_0.VOUT-.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X218 two_stage_opamp_dummy_magic_0.VOUT+.t57 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 bgr_0.V_p_2.t9 bgr_0.V_CUR_REF_REG.t4 bgr_0.1st_Vout_2.t9 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X220 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 bgr_0.PFET_GATE_10uA.t16 VDDA.t200 VDDA.t199 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X221 two_stage_opamp_dummy_magic_0.VOUT-.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VDDA.t214 bgr_0.PFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 VDDA.t213 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X223 two_stage_opamp_dummy_magic_0.V_source.t12 VIN+.t2 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA.t147 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X224 two_stage_opamp_dummy_magic_0.VOUT+.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X225 GNDA.t20 two_stage_opamp_dummy_magic_0.Y.t33 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X226 a_11220_17290.t0 GNDA.t24 GNDA.t23 sky130_fd_pr__res_xhigh_po_0p35 l=6
X227 two_stage_opamp_dummy_magic_0.V_source.t13 VIN-.t2 two_stage_opamp_dummy_magic_0.VD1.t5 GNDA.t180 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X228 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA.t287 GNDA.t288 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X229 bgr_0.1st_Vout_1.t22 bgr_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 two_stage_opamp_dummy_magic_0.VOUT+.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 two_stage_opamp_dummy_magic_0.VOUT+.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 bgr_0.START_UP.t3 bgr_0.V_TOP.t23 VDDA.t305 VDDA.t304 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X233 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t5 VDDA.t252 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X234 two_stage_opamp_dummy_magic_0.V_source.t30 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA.t75 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X235 bgr_0.1st_Vout_2.t5 bgr_0.V_mir2.t18 VDDA.t134 VDDA.t133 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X236 bgr_0.V_TOP.t24 VDDA.t303 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X237 two_stage_opamp_dummy_magic_0.VOUT+.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 two_stage_opamp_dummy_magic_0.VOUT+.t62 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X239 two_stage_opamp_dummy_magic_0.VOUT-.t58 two_stage_opamp_dummy_magic_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 two_stage_opamp_dummy_magic_0.VOUT-.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 VDDA.t111 two_stage_opamp_dummy_magic_0.Vb3.t13 two_stage_opamp_dummy_magic_0.VD3.t22 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X242 VDDA.t181 bgr_0.V_mir1.t19 bgr_0.1st_Vout_1.t9 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X243 two_stage_opamp_dummy_magic_0.VOUT-.t10 two_stage_opamp_dummy_magic_0.X.t34 VDDA.t171 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X244 two_stage_opamp_dummy_magic_0.VD2.t1 two_stage_opamp_dummy_magic_0.Vb1.t11 two_stage_opamp_dummy_magic_0.Y.t1 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X245 two_stage_opamp_dummy_magic_0.VOUT+.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X246 two_stage_opamp_dummy_magic_0.VOUT+.t64 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X247 bgr_0.1st_Vout_1.t23 bgr_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 GNDA.t88 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 two_stage_opamp_dummy_magic_0.V_source.t29 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X249 bgr_0.V_p_2.t0 bgr_0.V_CUR_REF_REG.t5 bgr_0.1st_Vout_2.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X250 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 two_stage_opamp_dummy_magic_0.Y.t34 VDDA.t137 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X251 two_stage_opamp_dummy_magic_0.V_err_p.t20 VDDA.t404 VDDA.t406 VDDA.t405 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X252 two_stage_opamp_dummy_magic_0.VOUT-.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X253 two_stage_opamp_dummy_magic_0.VOUT-.t61 two_stage_opamp_dummy_magic_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 VDDA.t9 two_stage_opamp_dummy_magic_0.Vb3.t14 two_stage_opamp_dummy_magic_0.VD4.t21 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X255 two_stage_opamp_dummy_magic_0.VOUT+.t65 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 two_stage_opamp_dummy_magic_0.VOUT+.t66 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X257 two_stage_opamp_dummy_magic_0.VOUT-.t62 two_stage_opamp_dummy_magic_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X258 bgr_0.V_TOP.t25 VDDA.t302 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 GNDA.t229 GNDA.t279 bgr_0.Vbe2.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X260 two_stage_opamp_dummy_magic_0.VOUT-.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X261 two_stage_opamp_dummy_magic_0.VOUT+.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 two_stage_opamp_dummy_magic_0.VOUT+.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X263 VDDA.t259 two_stage_opamp_dummy_magic_0.Vb3.t15 two_stage_opamp_dummy_magic_0.VD3.t34 VDDA.t258 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X264 two_stage_opamp_dummy_magic_0.VOUT+.t9 two_stage_opamp_dummy_magic_0.Y.t35 VDDA.t139 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X265 two_stage_opamp_dummy_magic_0.Y.t13 two_stage_opamp_dummy_magic_0.Vb2.t15 two_stage_opamp_dummy_magic_0.VD4.t12 two_stage_opamp_dummy_magic_0.VD4.t11 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X266 two_stage_opamp_dummy_magic_0.VOUT-.t64 two_stage_opamp_dummy_magic_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X267 bgr_0.1st_Vout_2.t17 bgr_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 GNDA.t34 bgr_0.NFET_GATE_10uA.t10 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X269 two_stage_opamp_dummy_magic_0.VOUT+.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X270 VDDA.t95 two_stage_opamp_dummy_magic_0.V_err_gate.t19 two_stage_opamp_dummy_magic_0.V_err_p.t16 VDDA.t94 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X271 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0 ps=0 w=3.6 l=0.2
X272 two_stage_opamp_dummy_magic_0.VOUT-.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X273 a_14640_5068.t1 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA.t338 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X274 VDDA.t166 two_stage_opamp_dummy_magic_0.V_err_gate.t20 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X275 two_stage_opamp_dummy_magic_0.VD1.t17 two_stage_opamp_dummy_magic_0.Vb1.t12 two_stage_opamp_dummy_magic_0.X.t16 GNDA.t140 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X276 two_stage_opamp_dummy_magic_0.VOUT+.t70 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 two_stage_opamp_dummy_magic_0.V_tot.t5 two_stage_opamp_dummy_magic_0.V_err_p.t3 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X278 bgr_0.V_mir2.t7 bgr_0.V_mir2.t6 VDDA.t105 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X279 VDDA.t301 bgr_0.V_TOP.t26 bgr_0.Vin-.t3 VDDA.t300 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X280 GNDA.t148 two_stage_opamp_dummy_magic_0.X.t35 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 VDDA.t221 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X281 VDDA.t403 VDDA.t401 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 VDDA.t402 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X282 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 bgr_0.PFET_GATE_10uA.t18 VDDA.t198 VDDA.t197 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X283 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 VIN+.t3 two_stage_opamp_dummy_magic_0.V_p_mir.t0 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X284 two_stage_opamp_dummy_magic_0.V_source.t14 VIN-.t3 two_stage_opamp_dummy_magic_0.VD1.t6 GNDA.t181 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X285 two_stage_opamp_dummy_magic_0.VOUT-.t66 two_stage_opamp_dummy_magic_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X286 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 VDDA.t398 VDDA.t400 VDDA.t399 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=1.28 ps=7.2 w=3.2 l=0.2
X287 VDDA.t53 two_stage_opamp_dummy_magic_0.Y.t36 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X288 two_stage_opamp_dummy_magic_0.VOUT+.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X289 two_stage_opamp_dummy_magic_0.VOUT-.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 bgr_0.Vin-.t1 a_12828_17650.t0 GNDA.t23 sky130_fd_pr__res_xhigh_po_0p35 l=6
X291 two_stage_opamp_dummy_magic_0.VOUT-.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X292 two_stage_opamp_dummy_magic_0.VOUT+.t72 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X293 two_stage_opamp_dummy_magic_0.VOUT+.t73 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X294 GNDA.t231 GNDA.t283 bgr_0.Vbe2.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X295 two_stage_opamp_dummy_magic_0.V_source.t20 VIN-.t4 two_stage_opamp_dummy_magic_0.VD1.t10 GNDA.t331 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X296 two_stage_opamp_dummy_magic_0.Y.t17 two_stage_opamp_dummy_magic_0.Vb2.t16 two_stage_opamp_dummy_magic_0.VD4.t10 two_stage_opamp_dummy_magic_0.VD4.t9 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X297 VDDA.t136 two_stage_opamp_dummy_magic_0.Vb3.t16 two_stage_opamp_dummy_magic_0.VD3.t23 VDDA.t135 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X298 GNDA.t46 two_stage_opamp_dummy_magic_0.Y.t37 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X299 two_stage_opamp_dummy_magic_0.VD4.t30 VDDA.t395 VDDA.t397 VDDA.t396 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X300 GNDA.t13 two_stage_opamp_dummy_magic_0.Y.t38 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X301 two_stage_opamp_dummy_magic_0.VOUT+.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X302 two_stage_opamp_dummy_magic_0.VOUT-.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X303 two_stage_opamp_dummy_magic_0.VOUT-.t70 two_stage_opamp_dummy_magic_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 bgr_0.1st_Vout_2.t18 bgr_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 GNDA.t36 bgr_0.NFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X306 bgr_0.PFET_GATE_10uA.t0 bgr_0.1st_Vout_2.t19 VDDA.t7 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X307 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 two_stage_opamp_dummy_magic_0.V_tot.t6 two_stage_opamp_dummy_magic_0.V_err_gate.t1 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X308 two_stage_opamp_dummy_magic_0.VOUT+.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 two_stage_opamp_dummy_magic_0.VOUT+.t76 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA.t284 GNDA.t286 GNDA.t285 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X311 GNDA.t282 GNDA.t280 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA.t281 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X312 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_tot.t7 two_stage_opamp_dummy_magic_0.V_err_gate.t0 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X313 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 bgr_0.NFET_GATE_10uA.t12 GNDA.t118 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X314 bgr_0.START_UP.t5 bgr_0.START_UP.t4 bgr_0.START_UP_NFET1.t0 GNDA.t161 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X315 two_stage_opamp_dummy_magic_0.VOUT-.t2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA.t65 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X316 two_stage_opamp_dummy_magic_0.VOUT-.t9 two_stage_opamp_dummy_magic_0.X.t36 VDDA.t223 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X317 two_stage_opamp_dummy_magic_0.VOUT+.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X318 two_stage_opamp_dummy_magic_0.VOUT-.t71 two_stage_opamp_dummy_magic_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 two_stage_opamp_dummy_magic_0.VOUT-.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X320 two_stage_opamp_dummy_magic_0.VOUT-.t73 two_stage_opamp_dummy_magic_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X321 two_stage_opamp_dummy_magic_0.VOUT-.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 two_stage_opamp_dummy_magic_0.VOUT+.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X323 two_stage_opamp_dummy_magic_0.VOUT+.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 two_stage_opamp_dummy_magic_0.VOUT+.t80 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 GNDA.t120 bgr_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA.t119 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X326 bgr_0.V_p_1.t3 bgr_0.Vin+.t7 bgr_0.1st_Vout_1.t5 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X327 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 two_stage_opamp_dummy_magic_0.V_err_gate.t21 VDDA.t168 VDDA.t167 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X328 two_stage_opamp_dummy_magic_0.Vb2.t5 bgr_0.NFET_GATE_10uA.t14 GNDA.t57 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X329 two_stage_opamp_dummy_magic_0.Vb2.t4 bgr_0.NFET_GATE_10uA.t15 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X330 two_stage_opamp_dummy_magic_0.VOUT+.t81 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 two_stage_opamp_dummy_magic_0.VD3.t19 two_stage_opamp_dummy_magic_0.Vb2.t17 two_stage_opamp_dummy_magic_0.X.t3 two_stage_opamp_dummy_magic_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X332 bgr_0.1st_Vout_2.t20 bgr_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X333 two_stage_opamp_dummy_magic_0.VOUT+.t0 two_stage_opamp_dummy_magic_0.Y.t39 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X334 two_stage_opamp_dummy_magic_0.VOUT+.t7 two_stage_opamp_dummy_magic_0.Y.t40 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X335 VDDA.t183 two_stage_opamp_dummy_magic_0.X.t37 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X336 bgr_0.Vin+.t4 bgr_0.V_TOP.t27 VDDA.t299 VDDA.t298 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X337 two_stage_opamp_dummy_magic_0.VOUT-.t75 two_stage_opamp_dummy_magic_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 two_stage_opamp_dummy_magic_0.VOUT-.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X339 two_stage_opamp_dummy_magic_0.VOUT-.t14 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA.t150 GNDA.t149 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X340 two_stage_opamp_dummy_magic_0.VOUT+.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X341 VDDA.t156 two_stage_opamp_dummy_magic_0.V_err_gate.t22 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 VDDA.t155 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X342 two_stage_opamp_dummy_magic_0.VD3.t32 two_stage_opamp_dummy_magic_0.Vb3.t17 VDDA.t208 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X343 VDDA.t468 bgr_0.PFET_GATE_10uA.t19 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 VDDA.t467 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X344 two_stage_opamp_dummy_magic_0.VOUT-.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 bgr_0.PFET_GATE_10uA.t20 VDDA.t454 VDDA.t453 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X346 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 two_stage_opamp_dummy_magic_0.V_tot.t8 two_stage_opamp_dummy_magic_0.V_err_p.t1 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X347 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 GNDA.t208 GNDA.t207 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X348 two_stage_opamp_dummy_magic_0.VD1.t16 two_stage_opamp_dummy_magic_0.Vb1.t13 two_stage_opamp_dummy_magic_0.X.t21 GNDA.t330 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X349 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 two_stage_opamp_dummy_magic_0.Y.t0 GNDA.t2 sky130_fd_pr__res_high_po_1p41 l=1.41
X350 two_stage_opamp_dummy_magic_0.err_amp_out.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 two_stage_opamp_dummy_magic_0.V_err_p.t6 VDDA.t253 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X351 two_stage_opamp_dummy_magic_0.VOUT-.t78 two_stage_opamp_dummy_magic_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 GNDA.t100 two_stage_opamp_dummy_magic_0.X.t38 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X353 two_stage_opamp_dummy_magic_0.VOUT-.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 two_stage_opamp_dummy_magic_0.VOUT+.t83 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X355 two_stage_opamp_dummy_magic_0.VOUT+.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 bgr_0.V_TOP.t28 VDDA.t295 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X357 bgr_0.Vin+.t0 a_12828_17530.t0 GNDA.t23 sky130_fd_pr__res_xhigh_po_0p35 l=6
X358 two_stage_opamp_dummy_magic_0.V_source.t10 VIN+.t4 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X359 two_stage_opamp_dummy_magic_0.VOUT+.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 two_stage_opamp_dummy_magic_0.VD4.t22 two_stage_opamp_dummy_magic_0.Vb3.t18 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X361 VDDA.t124 two_stage_opamp_dummy_magic_0.Y.t41 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X362 two_stage_opamp_dummy_magic_0.VOUT-.t80 two_stage_opamp_dummy_magic_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 bgr_0.1st_Vout_1.t24 bgr_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X364 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA.t276 GNDA.t278 GNDA.t277 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X365 GNDA.t275 GNDA.t273 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 GNDA.t274 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X366 two_stage_opamp_dummy_magic_0.Vb3.t3 bgr_0.NFET_GATE_10uA.t16 GNDA.t53 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X367 GNDA.t55 bgr_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X368 two_stage_opamp_dummy_magic_0.V_source.t11 VIN+.t5 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X369 bgr_0.V_mir1.t7 bgr_0.V_mir1.t6 VDDA.t107 VDDA.t106 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X370 GNDA.t102 two_stage_opamp_dummy_magic_0.Y.t42 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X371 a_5230_5068.t1 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA.t114 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X372 two_stage_opamp_dummy_magic_0.VOUT-.t81 two_stage_opamp_dummy_magic_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X373 two_stage_opamp_dummy_magic_0.VOUT-.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X374 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 two_stage_opamp_dummy_magic_0.V_err_gate.t4 VDDA.t251 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X375 two_stage_opamp_dummy_magic_0.VOUT-.t83 two_stage_opamp_dummy_magic_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X376 bgr_0.V_p_2.t4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 bgr_0.V_mir2.t15 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X377 two_stage_opamp_dummy_magic_0.VOUT-.t84 two_stage_opamp_dummy_magic_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 VDDA.t464 bgr_0.PFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_0.Vb1.t5 VDDA.t463 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X379 two_stage_opamp_dummy_magic_0.VD2.t5 two_stage_opamp_dummy_magic_0.Vb1.t14 two_stage_opamp_dummy_magic_0.Y.t6 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X380 two_stage_opamp_dummy_magic_0.VOUT+.t86 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X381 two_stage_opamp_dummy_magic_0.VOUT-.t85 two_stage_opamp_dummy_magic_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 two_stage_opamp_dummy_magic_0.VOUT-.t8 two_stage_opamp_dummy_magic_0.X.t39 VDDA.t129 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X383 two_stage_opamp_dummy_magic_0.VOUT+.t87 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 two_stage_opamp_dummy_magic_0.VD4.t26 two_stage_opamp_dummy_magic_0.Vb3.t19 VDDA.t231 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X385 bgr_0.V_p_1.t2 bgr_0.Vin+.t8 bgr_0.1st_Vout_1.t10 GNDA.t162 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X386 two_stage_opamp_dummy_magic_0.VOUT-.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 VDDA.t294 bgr_0.V_TOP.t29 bgr_0.START_UP.t2 VDDA.t293 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X388 two_stage_opamp_dummy_magic_0.V_err_p.t15 two_stage_opamp_dummy_magic_0.V_err_gate.t23 VDDA.t158 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X389 two_stage_opamp_dummy_magic_0.VD4.t8 two_stage_opamp_dummy_magic_0.Vb2.t18 two_stage_opamp_dummy_magic_0.Y.t23 two_stage_opamp_dummy_magic_0.VD4.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X390 two_stage_opamp_dummy_magic_0.VOUT-.t87 two_stage_opamp_dummy_magic_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 bgr_0.1st_Vout_2.t21 bgr_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X392 bgr_0.V_mir1.t5 bgr_0.V_mir1.t4 VDDA.t82 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X393 two_stage_opamp_dummy_magic_0.VOUT+.t88 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X394 two_stage_opamp_dummy_magic_0.VOUT-.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X395 two_stage_opamp_dummy_magic_0.Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2.t19 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4 as=0.72 ps=4 w=3.6 l=0.2
X396 a_14520_5068.t1 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA.t143 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X397 bgr_0.V_p_2.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 bgr_0.V_mir2.t14 GNDA.t173 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X398 two_stage_opamp_dummy_magic_0.VOUT+.t6 two_stage_opamp_dummy_magic_0.Y.t43 VDDA.t121 VDDA.t120 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X399 two_stage_opamp_dummy_magic_0.VOUT+.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VDDA.t169 two_stage_opamp_dummy_magic_0.X.t40 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X401 two_stage_opamp_dummy_magic_0.VOUT-.t89 two_stage_opamp_dummy_magic_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 bgr_0.1st_Vout_2.t22 bgr_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X403 VDDA.t97 two_stage_opamp_dummy_magic_0.V_err_gate.t24 two_stage_opamp_dummy_magic_0.V_err_p.t14 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X404 two_stage_opamp_dummy_magic_0.err_amp_out.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 two_stage_opamp_dummy_magic_0.V_err_p.t7 VDDA.t250 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X405 two_stage_opamp_dummy_magic_0.err_amp_out.t11 GNDA.t270 GNDA.t272 GNDA.t271 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X406 two_stage_opamp_dummy_magic_0.VD1.t15 two_stage_opamp_dummy_magic_0.Vb1.t15 two_stage_opamp_dummy_magic_0.X.t15 GNDA.t130 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X407 GNDA.t156 two_stage_opamp_dummy_magic_0.X.t41 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 VDDA.t233 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X408 two_stage_opamp_dummy_magic_0.VOUT+.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X409 two_stage_opamp_dummy_magic_0.VOUT+.t91 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X410 VDDA.t241 two_stage_opamp_dummy_magic_0.Vb3.t20 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=0.64 ps=3.6 w=3.2 l=0.2
X411 GNDA.t129 two_stage_opamp_dummy_magic_0.X.t42 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 VDDA.t184 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X412 two_stage_opamp_dummy_magic_0.VOUT+.t92 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X413 two_stage_opamp_dummy_magic_0.V_source.t5 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X414 VDDA.t190 two_stage_opamp_dummy_magic_0.Y.t44 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA.t134 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X415 two_stage_opamp_dummy_magic_0.V_source.t40 VIN-.t5 two_stage_opamp_dummy_magic_0.VD1.t21 GNDA.t341 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X416 bgr_0.1st_Vout_1.t0 bgr_0.V_mir1.t20 VDDA.t3 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X417 VDDA.t99 two_stage_opamp_dummy_magic_0.V_err_gate.t25 two_stage_opamp_dummy_magic_0.V_err_p.t13 VDDA.t98 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X418 VDDA.t191 two_stage_opamp_dummy_magic_0.Y.t45 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X419 GNDA.t345 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 two_stage_opamp_dummy_magic_0.VOUT+.t18 GNDA.t344 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X420 GNDA.t196 VDDA.t469 bgr_0.V_TOP.t12 GNDA.t185 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X421 two_stage_opamp_dummy_magic_0.VD3.t33 two_stage_opamp_dummy_magic_0.Vb3.t21 VDDA.t237 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X422 two_stage_opamp_dummy_magic_0.VOUT-.t90 two_stage_opamp_dummy_magic_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 two_stage_opamp_dummy_magic_0.X.t24 two_stage_opamp_dummy_magic_0.VD3.t25 two_stage_opamp_dummy_magic_0.VD3.t27 two_stage_opamp_dummy_magic_0.VD3.t26 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X424 GNDA.t206 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 two_stage_opamp_dummy_magic_0.err_amp_out.t8 GNDA.t205 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X425 two_stage_opamp_dummy_magic_0.VOUT-.t91 two_stage_opamp_dummy_magic_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X426 two_stage_opamp_dummy_magic_0.VOUT-.t92 two_stage_opamp_dummy_magic_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X427 bgr_0.1st_Vout_2.t4 bgr_0.V_mir2.t19 VDDA.t225 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X428 two_stage_opamp_dummy_magic_0.VOUT-.t93 two_stage_opamp_dummy_magic_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X429 two_stage_opamp_dummy_magic_0.VOUT-.t94 two_stage_opamp_dummy_magic_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X430 bgr_0.1st_Vout_2.t23 bgr_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X431 two_stage_opamp_dummy_magic_0.VOUT-.t95 two_stage_opamp_dummy_magic_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X432 GNDA.t29 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 two_stage_opamp_dummy_magic_0.VOUT-.t1 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X433 two_stage_opamp_dummy_magic_0.VOUT+.t93 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X434 bgr_0.1st_Vout_2.t24 bgr_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X435 VDDA.t175 bgr_0.PFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X436 two_stage_opamp_dummy_magic_0.VOUT+.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X437 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 two_stage_opamp_dummy_magic_0.V_err_gate.t26 VDDA.t162 VDDA.t161 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X438 bgr_0.1st_Vout_1.t25 bgr_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 two_stage_opamp_dummy_magic_0.VOUT-.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 bgr_0.V_TOP.t30 VDDA.t292 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 two_stage_opamp_dummy_magic_0.V_tot.t9 two_stage_opamp_dummy_magic_0.V_err_gate.t13 VDDA.t443 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X442 two_stage_opamp_dummy_magic_0.VOUT+.t95 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 bgr_0.START_UP.t1 bgr_0.V_TOP.t31 VDDA.t291 VDDA.t290 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X444 two_stage_opamp_dummy_magic_0.VOUT+.t96 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X445 two_stage_opamp_dummy_magic_0.VOUT-.t97 two_stage_opamp_dummy_magic_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X446 two_stage_opamp_dummy_magic_0.VOUT-.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X447 GNDA.t269 GNDA.t267 two_stage_opamp_dummy_magic_0.VOUT+.t15 GNDA.t268 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X448 two_stage_opamp_dummy_magic_0.VD2.t14 two_stage_opamp_dummy_magic_0.Vb1.t16 two_stage_opamp_dummy_magic_0.Y.t18 GNDA.t153 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X449 two_stage_opamp_dummy_magic_0.VOUT-.t7 two_stage_opamp_dummy_magic_0.X.t43 VDDA.t85 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X450 two_stage_opamp_dummy_magic_0.VOUT-.t6 two_stage_opamp_dummy_magic_0.X.t44 VDDA.t17 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X451 bgr_0.1st_Vout_1.t26 bgr_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 bgr_0.V_mir2.t5 bgr_0.V_mir2.t4 VDDA.t247 VDDA.t246 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X453 two_stage_opamp_dummy_magic_0.VOUT-.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X454 two_stage_opamp_dummy_magic_0.VOUT-.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 two_stage_opamp_dummy_magic_0.X.t4 two_stage_opamp_dummy_magic_0.Vb2.t20 two_stage_opamp_dummy_magic_0.VD3.t17 two_stage_opamp_dummy_magic_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X456 bgr_0.1st_Vout_2.t25 bgr_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 two_stage_opamp_dummy_magic_0.V_err_gate.t27 VDDA.t164 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X458 two_stage_opamp_dummy_magic_0.VOUT-.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 bgr_0.V_TOP.t8 bgr_0.1st_Vout_1.t27 VDDA.t436 VDDA.t435 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X460 two_stage_opamp_dummy_magic_0.VOUT+.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X461 two_stage_opamp_dummy_magic_0.VOUT+.t98 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 two_stage_opamp_dummy_magic_0.VOUT+.t99 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 bgr_0.1st_Vout_1.t28 bgr_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X464 GNDA.t266 GNDA.t263 GNDA.t265 GNDA.t264 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X465 GNDA.t248 GNDA.t261 bgr_0.Vbe2.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X466 bgr_0.V_mir2.t3 bgr_0.V_mir2.t2 VDDA.t245 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X467 VDDA.t289 bgr_0.V_TOP.t32 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 VDDA.t288 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X468 GNDA.t42 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 two_stage_opamp_dummy_magic_0.V_source.t28 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X469 VDDA.t18 two_stage_opamp_dummy_magic_0.X.t45 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X470 two_stage_opamp_dummy_magic_0.VOUT+.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X471 two_stage_opamp_dummy_magic_0.VOUT+.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 VDDA.t394 VDDA.t392 bgr_0.V_TOP.t1 VDDA.t393 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X473 two_stage_opamp_dummy_magic_0.V_err_gate.t3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 VDDA.t249 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X474 two_stage_opamp_dummy_magic_0.VOUT-.t102 two_stage_opamp_dummy_magic_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 VDDA.t152 two_stage_opamp_dummy_magic_0.V_err_gate.t28 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 VDDA.t151 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X476 two_stage_opamp_dummy_magic_0.VOUT+.t102 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 bgr_0.V_TOP.t33 VDDA.t287 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X478 VDDA.t78 two_stage_opamp_dummy_magic_0.Vb3.t22 two_stage_opamp_dummy_magic_0.VD4.t23 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X479 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 VDDA.t389 VDDA.t391 VDDA.t390 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X480 GNDA.t195 VDDA.t386 VDDA.t388 VDDA.t387 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X481 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 a_5750_2076.t0 GNDA.t142 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X482 two_stage_opamp_dummy_magic_0.V_source.t27 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA.t343 GNDA.t342 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X483 two_stage_opamp_dummy_magic_0.VOUT-.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X484 two_stage_opamp_dummy_magic_0.VOUT-.t104 two_stage_opamp_dummy_magic_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 two_stage_opamp_dummy_magic_0.VOUT-.t105 two_stage_opamp_dummy_magic_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X486 GNDA.t229 GNDA.t260 bgr_0.Vbe2.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X487 bgr_0.1st_Vout_1.t29 bgr_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X488 two_stage_opamp_dummy_magic_0.V_source.t7 VIN+.t6 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X489 bgr_0.V_TOP.t34 VDDA.t286 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X490 VDDA.t188 two_stage_opamp_dummy_magic_0.Y.t46 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X491 two_stage_opamp_dummy_magic_0.VOUT-.t106 two_stage_opamp_dummy_magic_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X492 two_stage_opamp_dummy_magic_0.VOUT+.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 bgr_0.PFET_GATE_10uA.t1 bgr_0.1st_Vout_2.t26 VDDA.t38 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X494 a_13790_17550.t0 bgr_0.V_CUR_REF_REG.t0 GNDA.t60 sky130_fd_pr__res_xhigh_po_0p35 l=6
X495 GNDA.t204 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X496 two_stage_opamp_dummy_magic_0.VOUT+.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X497 VDDA.t196 bgr_0.PFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 VDDA.t195 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X498 VDDA.t285 bgr_0.V_TOP.t35 bgr_0.Vin+.t3 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X499 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 VDDA.t383 VDDA.t385 VDDA.t384 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X500 a_5350_5068.t0 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA.t12 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X501 bgr_0.1st_Vout_2.t27 bgr_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X502 two_stage_opamp_dummy_magic_0.VOUT+.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X503 GNDA.t194 VDDA.t470 bgr_0.V_p_2.t6 GNDA.t193 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=5
X504 two_stage_opamp_dummy_magic_0.VOUT+.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X505 GNDA.t202 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 GNDA.t201 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X506 two_stage_opamp_dummy_magic_0.X.t22 two_stage_opamp_dummy_magic_0.Vb1.t17 two_stage_opamp_dummy_magic_0.VD1.t14 GNDA.t333 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X507 bgr_0.V_p_1.t7 bgr_0.Vin-.t10 bgr_0.V_mir1.t14 GNDA.t185 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X508 VDDA.t1 two_stage_opamp_dummy_magic_0.Vb3.t23 two_stage_opamp_dummy_magic_0.VD4.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X509 two_stage_opamp_dummy_magic_0.X.t7 two_stage_opamp_dummy_magic_0.Vb2.t21 two_stage_opamp_dummy_magic_0.VD3.t15 two_stage_opamp_dummy_magic_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X510 two_stage_opamp_dummy_magic_0.VOUT+.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X511 two_stage_opamp_dummy_magic_0.VOUT-.t107 two_stage_opamp_dummy_magic_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X512 bgr_0.V_TOP.t6 bgr_0.1st_Vout_1.t30 VDDA.t432 VDDA.t431 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X513 two_stage_opamp_dummy_magic_0.VOUT-.t16 VDDA.t380 VDDA.t382 VDDA.t381 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X514 two_stage_opamp_dummy_magic_0.VD2.t21 two_stage_opamp_dummy_magic_0.Vb1.t18 two_stage_opamp_dummy_magic_0.Y.t24 GNDA.t340 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X515 two_stage_opamp_dummy_magic_0.VOUT-.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X516 bgr_0.V_TOP.t36 VDDA.t283 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X517 two_stage_opamp_dummy_magic_0.VOUT-.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 two_stage_opamp_dummy_magic_0.VOUT+.t14 GNDA.t257 GNDA.t259 GNDA.t258 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X519 GNDA.t231 GNDA.t262 bgr_0.Vbe2.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X520 two_stage_opamp_dummy_magic_0.VD1.t4 VIN-.t6 two_stage_opamp_dummy_magic_0.V_source.t9 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X521 bgr_0.1st_Vout_1.t1 bgr_0.V_mir1.t21 VDDA.t5 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X522 two_stage_opamp_dummy_magic_0.VOUT+.t108 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 two_stage_opamp_dummy_magic_0.VOUT+.t109 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X524 two_stage_opamp_dummy_magic_0.VOUT-.t110 two_stage_opamp_dummy_magic_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 two_stage_opamp_dummy_magic_0.VOUT+.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X526 two_stage_opamp_dummy_magic_0.VOUT+.t111 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X527 two_stage_opamp_dummy_magic_0.VOUT+.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 two_stage_opamp_dummy_magic_0.VOUT+.t113 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 bgr_0.Vin+.t2 bgr_0.V_TOP.t37 VDDA.t282 VDDA.t281 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X530 bgr_0.V_mir2.t13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 bgr_0.V_p_2.t2 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X531 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_0.Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 sky130_fd_pr__pfet_01v8 ad=1.44 pd=8 as=0.72 ps=4 w=3.6 l=0.2
X532 bgr_0.1st_Vout_2.t28 bgr_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X533 bgr_0.PFET_GATE_10uA.t7 VDDA.t471 GNDA.t192 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X534 two_stage_opamp_dummy_magic_0.VD1.t2 VIN-.t7 two_stage_opamp_dummy_magic_0.V_source.t4 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X535 two_stage_opamp_dummy_magic_0.VOUT-.t111 two_stage_opamp_dummy_magic_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 bgr_0.1st_Vout_2.t29 bgr_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X537 two_stage_opamp_dummy_magic_0.VOUT+.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X538 two_stage_opamp_dummy_magic_0.VOUT+.t115 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X539 VDDA.t192 two_stage_opamp_dummy_magic_0.X.t46 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X540 two_stage_opamp_dummy_magic_0.VOUT-.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X541 GNDA.t256 GNDA.t254 bgr_0.NFET_GATE_10uA.t3 GNDA.t255 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X542 two_stage_opamp_dummy_magic_0.VOUT-.t113 two_stage_opamp_dummy_magic_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X543 GNDA.t152 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 two_stage_opamp_dummy_magic_0.V_source.t26 GNDA.t151 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X544 two_stage_opamp_dummy_magic_0.V_err_gate.t7 bgr_0.NFET_GATE_10uA.t18 GNDA.t164 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X545 bgr_0.1st_Vout_1.t2 bgr_0.Vin+.t9 bgr_0.V_p_1.t1 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X546 VDDA.t256 two_stage_opamp_dummy_magic_0.X.t47 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA.t179 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X547 two_stage_opamp_dummy_magic_0.VOUT+.t3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA.t84 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X548 VDDA.t379 VDDA.t377 VDDA.t379 VDDA.t378 sky130_fd_pr__pfet_01v8 ad=0.64 pd=3.6 as=0 ps=0 w=3.2 l=0.2
X549 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.X.t12 GNDA.t63 sky130_fd_pr__res_high_po_1p41 l=1.41
X550 bgr_0.V_TOP.t7 bgr_0.1st_Vout_1.t31 VDDA.t434 VDDA.t433 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X551 two_stage_opamp_dummy_magic_0.VOUT+.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X552 two_stage_opamp_dummy_magic_0.VOUT-.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 bgr_0.PFET_GATE_10uA.t24 VDDA.t76 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X554 two_stage_opamp_dummy_magic_0.VOUT+.t117 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X555 two_stage_opamp_dummy_magic_0.VOUT+.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X556 bgr_0.Vin-.t5 bgr_0.V_TOP.t38 VDDA.t280 VDDA.t279 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X557 VDDA.t160 bgr_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 VDDA.t159 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X558 VDDA.t376 VDDA.t374 two_stage_opamp_dummy_magic_0.VD3.t35 VDDA.t375 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X559 two_stage_opamp_dummy_magic_0.VOUT-.t115 two_stage_opamp_dummy_magic_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X560 two_stage_opamp_dummy_magic_0.V_source.t25 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA.t67 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X561 two_stage_opamp_dummy_magic_0.VD3.t13 two_stage_opamp_dummy_magic_0.Vb2.t22 two_stage_opamp_dummy_magic_0.X.t6 two_stage_opamp_dummy_magic_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X562 two_stage_opamp_dummy_magic_0.VOUT+.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X563 a_13790_17550.t1 GNDA.t89 GNDA.t60 sky130_fd_pr__res_xhigh_po_0p35 l=6
X564 two_stage_opamp_dummy_magic_0.VOUT-.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 two_stage_opamp_dummy_magic_0.VOUT-.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X566 bgr_0.V_TOP.t5 VDDA.t371 VDDA.t373 VDDA.t372 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X567 GNDA.t200 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t7 GNDA.t199 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X568 VDDA.t370 VDDA.t368 two_stage_opamp_dummy_magic_0.VD4.t29 VDDA.t369 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X569 two_stage_opamp_dummy_magic_0.VOUT-.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 two_stage_opamp_dummy_magic_0.VOUT-.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X571 two_stage_opamp_dummy_magic_0.VOUT+.t120 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 GNDA.t191 VDDA.t365 VDDA.t367 VDDA.t366 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X573 bgr_0.V_TOP.t39 VDDA.t278 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 two_stage_opamp_dummy_magic_0.VOUT-.t120 two_stage_opamp_dummy_magic_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X575 two_stage_opamp_dummy_magic_0.VOUT+.t121 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X576 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 bgr_0.NFET_GATE_10uA.t19 GNDA.t166 GNDA.t165 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X577 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 bgr_0.NFET_GATE_10uA.t20 GNDA.t168 GNDA.t167 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X578 two_stage_opamp_dummy_magic_0.VOUT+.t122 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X579 two_stage_opamp_dummy_magic_0.VOUT-.t121 two_stage_opamp_dummy_magic_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 bgr_0.1st_Vout_1.t32 bgr_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X581 VDDA.t227 bgr_0.V_mir2.t20 bgr_0.1st_Vout_2.t3 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X582 VDDA.t364 VDDA.t362 two_stage_opamp_dummy_magic_0.err_amp_out.t5 VDDA.t363 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X583 two_stage_opamp_dummy_magic_0.X.t14 two_stage_opamp_dummy_magic_0.Vb1.t19 two_stage_opamp_dummy_magic_0.VD1.t13 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X584 two_stage_opamp_dummy_magic_0.VOUT+.t123 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X585 bgr_0.V_TOP.t40 VDDA.t277 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X586 VDDA.t276 bgr_0.V_TOP.t41 bgr_0.Vin+.t1 VDDA.t275 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X587 VDDA.t361 VDDA.t359 GNDA.t190 VDDA.t360 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X588 two_stage_opamp_dummy_magic_0.VOUT+.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X589 two_stage_opamp_dummy_magic_0.VD2.t10 two_stage_opamp_dummy_magic_0.Vb1.t20 two_stage_opamp_dummy_magic_0.Y.t14 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X590 two_stage_opamp_dummy_magic_0.VD3.t11 two_stage_opamp_dummy_magic_0.Vb2.t23 two_stage_opamp_dummy_magic_0.X.t5 two_stage_opamp_dummy_magic_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X591 bgr_0.V_mir1.t3 bgr_0.V_mir1.t2 VDDA.t109 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X592 two_stage_opamp_dummy_magic_0.VOUT+.t125 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X593 two_stage_opamp_dummy_magic_0.Vb2.t3 bgr_0.NFET_GATE_10uA.t21 GNDA.t170 GNDA.t169 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X594 two_stage_opamp_dummy_magic_0.Y.t21 two_stage_opamp_dummy_magic_0.Vb2.t24 two_stage_opamp_dummy_magic_0.VD4.t6 two_stage_opamp_dummy_magic_0.VD4.t5 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X595 GNDA.t229 GNDA.t228 bgr_0.Vbe2.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X596 bgr_0.V_mir2.t12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 bgr_0.V_p_2.t1 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X597 bgr_0.PFET_GATE_10uA.t6 VDDA.t356 VDDA.t358 VDDA.t357 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X598 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 two_stage_opamp_dummy_magic_0.Y.t47 GNDA.t133 VDDA.t189 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X599 two_stage_opamp_dummy_magic_0.VD2.t15 VIN+.t7 two_stage_opamp_dummy_magic_0.V_source.t15 GNDA.t221 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X600 two_stage_opamp_dummy_magic_0.VOUT-.t122 two_stage_opamp_dummy_magic_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X601 two_stage_opamp_dummy_magic_0.VOUT+.t13 VDDA.t353 VDDA.t355 VDDA.t354 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X602 VDDA.t112 GNDA.t251 GNDA.t253 GNDA.t252 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X603 two_stage_opamp_dummy_magic_0.VOUT+.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 GNDA.t325 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 two_stage_opamp_dummy_magic_0.V_source.t24 GNDA.t324 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X605 two_stage_opamp_dummy_magic_0.V_err_gate.t10 two_stage_opamp_dummy_magic_0.V_tot.t10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 VDDA.t257 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X606 two_stage_opamp_dummy_magic_0.VOUT-.t123 two_stage_opamp_dummy_magic_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 VDDA.t352 VDDA.t350 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 VDDA.t351 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X608 two_stage_opamp_dummy_magic_0.VD4.t24 two_stage_opamp_dummy_magic_0.Vb3.t24 VDDA.t204 VDDA.t203 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X609 two_stage_opamp_dummy_magic_0.VD3.t9 two_stage_opamp_dummy_magic_0.Vb2.t25 two_stage_opamp_dummy_magic_0.X.t8 two_stage_opamp_dummy_magic_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X610 two_stage_opamp_dummy_magic_0.VOUT+.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X611 bgr_0.V_TOP.t42 VDDA.t274 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X612 two_stage_opamp_dummy_magic_0.VOUT+.t17 a_5750_2076.t1 GNDA.t337 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X613 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 bgr_0.PFET_GATE_10uA.t26 VDDA.t452 VDDA.t451 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X614 two_stage_opamp_dummy_magic_0.VOUT-.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X615 two_stage_opamp_dummy_magic_0.VOUT-.t125 two_stage_opamp_dummy_magic_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X616 two_stage_opamp_dummy_magic_0.Y.t5 two_stage_opamp_dummy_magic_0.Vb1.t21 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X617 VDDA.t349 VDDA.t347 two_stage_opamp_dummy_magic_0.VOUT-.t15 VDDA.t348 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X618 two_stage_opamp_dummy_magic_0.VOUT+.t128 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X619 bgr_0.1st_Vout_2.t2 bgr_0.V_mir2.t21 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X620 two_stage_opamp_dummy_magic_0.V_source.t23 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 GNDA.t72 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X621 VDDA.t346 VDDA.t343 VDDA.t345 VDDA.t344 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0 ps=0 w=0.63 l=0.2
X622 bgr_0.1st_Vout_2.t30 bgr_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X623 a_5350_5068.t1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA.t336 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X624 GNDA.t231 GNDA.t230 bgr_0.Vin-.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X625 two_stage_opamp_dummy_magic_0.VOUT-.t126 two_stage_opamp_dummy_magic_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 GNDA.t108 bgr_0.NFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X627 two_stage_opamp_dummy_magic_0.VOUT-.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X628 two_stage_opamp_dummy_magic_0.VOUT-.t128 two_stage_opamp_dummy_magic_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X629 VDDA.t186 two_stage_opamp_dummy_magic_0.Y.t48 two_stage_opamp_dummy_magic_0.VOUT+.t10 VDDA.t185 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X630 two_stage_opamp_dummy_magic_0.VOUT+.t129 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X631 two_stage_opamp_dummy_magic_0.VOUT-.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X632 two_stage_opamp_dummy_magic_0.V_source.t22 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA.t10 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X633 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 bgr_0.V_TOP.t43 VDDA.t273 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X634 bgr_0.1st_Vout_2.t31 bgr_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 VDDA.t340 VDDA.t342 VDDA.t341 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X636 two_stage_opamp_dummy_magic_0.VD3.t7 two_stage_opamp_dummy_magic_0.Vb2.t26 two_stage_opamp_dummy_magic_0.X.t0 two_stage_opamp_dummy_magic_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X637 two_stage_opamp_dummy_magic_0.VD4.t27 two_stage_opamp_dummy_magic_0.Vb3.t25 VDDA.t235 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X638 two_stage_opamp_dummy_magic_0.V_err_p.t12 two_stage_opamp_dummy_magic_0.V_err_gate.t29 VDDA.t154 VDDA.t153 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X639 two_stage_opamp_dummy_magic_0.VOUT+.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X640 two_stage_opamp_dummy_magic_0.VOUT+.t131 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 two_stage_opamp_dummy_magic_0.X.t13 two_stage_opamp_dummy_magic_0.Vb1.t22 two_stage_opamp_dummy_magic_0.VD1.t12 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X642 VDDA.t239 bgr_0.1st_Vout_2.t32 bgr_0.PFET_GATE_10uA.t4 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X643 VDDA.t339 VDDA.t337 two_stage_opamp_dummy_magic_0.Vb1.t2 VDDA.t338 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X644 two_stage_opamp_dummy_magic_0.VOUT-.t130 two_stage_opamp_dummy_magic_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 two_stage_opamp_dummy_magic_0.Vb1.t1 VDDA.t334 VDDA.t336 VDDA.t335 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X646 two_stage_opamp_dummy_magic_0.V_err_p.t2 two_stage_opamp_dummy_magic_0.V_tot.t11 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 VDDA.t48 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X647 two_stage_opamp_dummy_magic_0.VOUT-.t131 two_stage_opamp_dummy_magic_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_0.X.t48 GNDA.t329 VDDA.t444 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X649 two_stage_opamp_dummy_magic_0.VD2.t2 VIN+.t8 two_stage_opamp_dummy_magic_0.V_source.t1 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X650 GNDA.t250 GNDA.t249 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X651 bgr_0.1st_Vout_2.t33 bgr_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X652 two_stage_opamp_dummy_magic_0.VOUT-.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 two_stage_opamp_dummy_magic_0.VOUT-.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X654 bgr_0.1st_Vout_2.t34 bgr_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 two_stage_opamp_dummy_magic_0.VOUT-.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 two_stage_opamp_dummy_magic_0.VOUT+.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X657 bgr_0.V_mir1.t13 bgr_0.Vin-.t11 bgr_0.V_p_1.t6 GNDA.t184 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X658 two_stage_opamp_dummy_magic_0.VOUT-.t135 two_stage_opamp_dummy_magic_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 two_stage_opamp_dummy_magic_0.VOUT-.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X660 two_stage_opamp_dummy_magic_0.VD2.t19 VIN+.t9 two_stage_opamp_dummy_magic_0.V_source.t19 GNDA.t328 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X661 two_stage_opamp_dummy_magic_0.VD3.t31 two_stage_opamp_dummy_magic_0.Vb3.t26 VDDA.t206 VDDA.t205 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X662 two_stage_opamp_dummy_magic_0.VOUT+.t133 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X663 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 two_stage_opamp_dummy_magic_0.Y.t49 GNDA.t131 VDDA.t187 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X664 VDDA.t333 VDDA.t331 GNDA.t189 VDDA.t332 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X665 bgr_0.1st_Vout_1.t33 bgr_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X666 GNDA.t347 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 two_stage_opamp_dummy_magic_0.V_p_mir.t2 GNDA.t346 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X667 two_stage_opamp_dummy_magic_0.V_err_gate.t2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X668 VDDA.t330 VDDA.t328 two_stage_opamp_dummy_magic_0.Vb2.t8 VDDA.t329 sky130_fd_pr__pfet_01v8 ad=0.252 pd=2.06 as=0.126 ps=1.03 w=0.63 l=0.2
X669 two_stage_opamp_dummy_magic_0.X.t9 two_stage_opamp_dummy_magic_0.Vb2.t27 two_stage_opamp_dummy_magic_0.VD3.t5 two_stage_opamp_dummy_magic_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X670 two_stage_opamp_dummy_magic_0.Y.t22 two_stage_opamp_dummy_magic_0.Vb1.t23 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA.t332 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X671 VDDA.t74 two_stage_opamp_dummy_magic_0.X.t49 two_stage_opamp_dummy_magic_0.VOUT-.t5 VDDA.t73 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X672 GNDA.t110 bgr_0.NFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X673 VDDA.t271 bgr_0.V_TOP.t44 bgr_0.START_UP.t0 VDDA.t270 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X674 two_stage_opamp_dummy_magic_0.VOUT-.t137 two_stage_opamp_dummy_magic_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X675 two_stage_opamp_dummy_magic_0.VD4.t4 two_stage_opamp_dummy_magic_0.Vb2.t28 two_stage_opamp_dummy_magic_0.Y.t10 two_stage_opamp_dummy_magic_0.VD4.t3 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X676 two_stage_opamp_dummy_magic_0.VOUT-.t138 two_stage_opamp_dummy_magic_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X677 two_stage_opamp_dummy_magic_0.V_source.t21 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA.t160 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X678 VDDA.t34 GNDA.t241 GNDA.t243 GNDA.t242 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X679 two_stage_opamp_dummy_magic_0.VOUT-.t139 two_stage_opamp_dummy_magic_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X680 VDDA.t147 two_stage_opamp_dummy_magic_0.V_err_gate.t30 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 VDDA.t146 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X681 two_stage_opamp_dummy_magic_0.VOUT+.t134 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X682 GNDA.t248 GNDA.t247 bgr_0.Vbe2.t0 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X683 two_stage_opamp_dummy_magic_0.VOUT+.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X684 two_stage_opamp_dummy_magic_0.VOUT+.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X685 VDDA.t117 two_stage_opamp_dummy_magic_0.Y.t50 two_stage_opamp_dummy_magic_0.VOUT+.t5 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X686 VDDA.t327 VDDA.t325 two_stage_opamp_dummy_magic_0.VOUT+.t12 VDDA.t326 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X687 VDDA.t243 bgr_0.V_mir2.t0 bgr_0.V_mir2.t1 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X688 VDDA.t458 bgr_0.PFET_GATE_10uA.t27 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 VDDA.t457 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X689 two_stage_opamp_dummy_magic_0.VOUT-.t140 two_stage_opamp_dummy_magic_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X690 bgr_0.1st_Vout_1.t34 bgr_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X691 GNDA.t246 GNDA.t244 VDDA.t35 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X692 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 bgr_0.PFET_GATE_10uA.t28 VDDA.t141 VDDA.t140 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X693 two_stage_opamp_dummy_magic_0.VOUT+.t137 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 bgr_0.V_TOP.t45 VDDA.t269 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 two_stage_opamp_dummy_magic_0.V_err_p.t11 two_stage_opamp_dummy_magic_0.V_err_gate.t31 VDDA.t149 VDDA.t148 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X696 bgr_0.1st_Vout_1.t6 bgr_0.V_mir1.t22 VDDA.t101 VDDA.t100 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X697 two_stage_opamp_dummy_magic_0.X.t23 two_stage_opamp_dummy_magic_0.Vb1.t24 two_stage_opamp_dummy_magic_0.VD1.t11 GNDA.t339 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X698 two_stage_opamp_dummy_magic_0.VOUT+.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X699 two_stage_opamp_dummy_magic_0.V_err_p.t4 two_stage_opamp_dummy_magic_0.V_tot.t12 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X700 two_stage_opamp_dummy_magic_0.V_err_p.t8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 two_stage_opamp_dummy_magic_0.err_amp_out.t1 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X701 two_stage_opamp_dummy_magic_0.VOUT-.t141 two_stage_opamp_dummy_magic_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_0.X.t50 GNDA.t334 VDDA.t456 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X703 bgr_0.1st_Vout_1.t35 bgr_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X704 bgr_0.1st_Vout_2.t8 bgr_0.V_CUR_REF_REG.t6 bgr_0.V_p_2.t8 GNDA.t319 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X705 bgr_0.V_TOP.t46 VDDA.t268 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X706 two_stage_opamp_dummy_magic_0.VD4.t2 two_stage_opamp_dummy_magic_0.Vb2.t29 two_stage_opamp_dummy_magic_0.Y.t16 two_stage_opamp_dummy_magic_0.VD4.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X707 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 two_stage_opamp_dummy_magic_0.Y.t51 VDDA.t118 GNDA.t101 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X708 two_stage_opamp_dummy_magic_0.V_p_mir.t1 VIN-.t8 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA.t159 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X709 two_stage_opamp_dummy_magic_0.VD1.t9 VIN-.t9 two_stage_opamp_dummy_magic_0.V_source.t18 GNDA.t323 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X710 two_stage_opamp_dummy_magic_0.VOUT-.t142 two_stage_opamp_dummy_magic_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X711 two_stage_opamp_dummy_magic_0.VOUT+.t139 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X712 two_stage_opamp_dummy_magic_0.VOUT+.t140 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 two_stage_opamp_dummy_magic_0.VOUT+.t141 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X714 bgr_0.V_p_1.t10 VDDA.t472 GNDA.t188 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=5
X715 GNDA.t113 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 two_stage_opamp_dummy_magic_0.VOUT-.t3 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X716 bgr_0.1st_Vout_2.t35 bgr_0.cap_res2.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X717 bgr_0.V_mir1.t12 bgr_0.Vin-.t12 bgr_0.V_p_1.t5 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X718 VDDA.t324 VDDA.t322 bgr_0.PFET_GATE_10uA.t5 VDDA.t323 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X719 two_stage_opamp_dummy_magic_0.VOUT+.t142 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 two_stage_opamp_dummy_magic_0.VOUT+.t143 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X721 two_stage_opamp_dummy_magic_0.VOUT-.t143 two_stage_opamp_dummy_magic_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X722 two_stage_opamp_dummy_magic_0.VD1.t1 VIN-.t10 two_stage_opamp_dummy_magic_0.V_source.t3 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X723 two_stage_opamp_dummy_magic_0.X.t2 two_stage_opamp_dummy_magic_0.Vb2.t30 two_stage_opamp_dummy_magic_0.VD3.t3 two_stage_opamp_dummy_magic_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X724 bgr_0.V_TOP.t47 VDDA.t267 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X725 VDDA.t446 two_stage_opamp_dummy_magic_0.Vb3.t27 two_stage_opamp_dummy_magic_0.VD4.t31 VDDA.t445 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X726 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 two_stage_opamp_dummy_magic_0.Y.t52 GNDA.t145 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X727 VDDA.t220 bgr_0.V_mir1.t0 bgr_0.V_mir1.t1 VDDA.t219 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X728 two_stage_opamp_dummy_magic_0.VOUT-.t144 two_stage_opamp_dummy_magic_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X729 two_stage_opamp_dummy_magic_0.VOUT-.t145 two_stage_opamp_dummy_magic_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X730 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 bgr_0.V_TOP.t48 VDDA.t266 VDDA.t265 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X731 bgr_0.V_TOP.t0 bgr_0.START_UP.t7 bgr_0.Vin-.t0 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X732 two_stage_opamp_dummy_magic_0.V_err_gate.t11 VDDA.t319 VDDA.t321 VDDA.t320 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X733 two_stage_opamp_dummy_magic_0.VOUT+.t144 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 bgr_0.1st_Vout_2.t7 bgr_0.V_CUR_REF_REG.t7 bgr_0.V_p_2.t7 GNDA.t318 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X735 two_stage_opamp_dummy_magic_0.V_err_gate.t9 two_stage_opamp_dummy_magic_0.V_tot.t13 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X736 two_stage_opamp_dummy_magic_0.VOUT-.t146 two_stage_opamp_dummy_magic_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 VDDA.t460 bgr_0.1st_Vout_2.t36 bgr_0.PFET_GATE_10uA.t8 VDDA.t459 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X738 bgr_0.1st_Vout_1.t36 bgr_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X739 two_stage_opamp_dummy_magic_0.Y.t9 two_stage_opamp_dummy_magic_0.Vb1.t25 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X740 two_stage_opamp_dummy_magic_0.Vb2.t1 two_stage_opamp_dummy_magic_0.Vb2.t0 VDDA.t63 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.126 pd=1.03 as=0.126 ps=1.03 w=0.63 l=0.2
X741 GNDA.t227 GNDA.t225 two_stage_opamp_dummy_magic_0.VOUT-.t17 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X742 VDDA.t194 two_stage_opamp_dummy_magic_0.X.t51 two_stage_opamp_dummy_magic_0.VOUT-.t4 VDDA.t193 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X743 two_stage_opamp_dummy_magic_0.VOUT-.t147 two_stage_opamp_dummy_magic_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 a_5230_5068.t0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA.t78 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X745 two_stage_opamp_dummy_magic_0.VOUT+.t145 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X746 two_stage_opamp_dummy_magic_0.VOUT+.t146 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 two_stage_opamp_dummy_magic_0.VOUT+.t147 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X748 two_stage_opamp_dummy_magic_0.VOUT-.t148 two_stage_opamp_dummy_magic_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 two_stage_opamp_dummy_magic_0.VOUT-.t149 two_stage_opamp_dummy_magic_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X750 two_stage_opamp_dummy_magic_0.VOUT+.t148 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 VDDA.t89 two_stage_opamp_dummy_magic_0.V_err_gate.t32 two_stage_opamp_dummy_magic_0.V_err_p.t10 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X752 two_stage_opamp_dummy_magic_0.Y.t12 two_stage_opamp_dummy_magic_0.VD4.t32 two_stage_opamp_dummy_magic_0.VD4.t34 two_stage_opamp_dummy_magic_0.VD4.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X753 two_stage_opamp_dummy_magic_0.VOUT+.t149 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X754 two_stage_opamp_dummy_magic_0.VOUT-.t150 two_stage_opamp_dummy_magic_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 VDDA.t318 VDDA.t316 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 VDDA.t317 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X756 two_stage_opamp_dummy_magic_0.VOUT+.t150 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X757 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 bgr_0.PFET_GATE_10uA.t29 VDDA.t143 VDDA.t142 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X758 two_stage_opamp_dummy_magic_0.X.t1 two_stage_opamp_dummy_magic_0.Vb2.t31 two_stage_opamp_dummy_magic_0.VD3.t1 two_stage_opamp_dummy_magic_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X759 two_stage_opamp_dummy_magic_0.VOUT-.t151 two_stage_opamp_dummy_magic_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X760 VDDA.t52 bgr_0.V_mir2.t22 bgr_0.1st_Vout_2.t1 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X761 VDDA.t211 two_stage_opamp_dummy_magic_0.Y.t53 two_stage_opamp_dummy_magic_0.VOUT+.t11 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X762 two_stage_opamp_dummy_magic_0.VOUT+.t151 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X763 two_stage_opamp_dummy_magic_0.VOUT-.t152 two_stage_opamp_dummy_magic_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X764 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 two_stage_opamp_dummy_magic_0.X.t52 VDDA.t44 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X765 two_stage_opamp_dummy_magic_0.VOUT-.t153 two_stage_opamp_dummy_magic_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X766 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 two_stage_opamp_dummy_magic_0.V_err_gate.t33 VDDA.t91 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X767 two_stage_opamp_dummy_magic_0.VOUT+.t152 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X768 two_stage_opamp_dummy_magic_0.X.t19 GNDA.t238 GNDA.t240 GNDA.t239 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X769 two_stage_opamp_dummy_magic_0.V_err_p.t5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t0 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X770 GNDA.t198 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 two_stage_opamp_dummy_magic_0.err_amp_out.t6 GNDA.t197 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X771 two_stage_opamp_dummy_magic_0.VOUT+.t153 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X772 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 two_stage_opamp_dummy_magic_0.X.t53 GNDA.t48 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X773 two_stage_opamp_dummy_magic_0.VOUT+.t154 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X774 two_stage_opamp_dummy_magic_0.VOUT-.t154 two_stage_opamp_dummy_magic_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X775 two_stage_opamp_dummy_magic_0.VOUT-.t155 two_stage_opamp_dummy_magic_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X776 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 two_stage_opamp_dummy_magic_0.X.t54 GNDA.t49 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X777 two_stage_opamp_dummy_magic_0.VOUT+.t155 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X778 bgr_0.V_TOP.t49 VDDA.t264 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X779 bgr_0.1st_Vout_1.t7 bgr_0.Vin+.t10 bgr_0.V_p_1.t0 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X780 GNDA.t237 GNDA.t235 two_stage_opamp_dummy_magic_0.V_source.t16 GNDA.t236 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X781 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA.t232 GNDA.t234 GNDA.t233 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X782 two_stage_opamp_dummy_magic_0.VOUT+.t156 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X783 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 two_stage_opamp_dummy_magic_0.Y.t54 VDDA.t212 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X784 GNDA.t224 GNDA.t222 VDDA.t232 GNDA.t223 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X785 two_stage_opamp_dummy_magic_0.VD2.t18 VIN+.t10 two_stage_opamp_dummy_magic_0.V_source.t17 GNDA.t317 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X786 bgr_0.Vin+.t5 bgr_0.Vbe2.t8 GNDA.t335 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X787 VDDA.t173 two_stage_opamp_dummy_magic_0.Vb3.t28 two_stage_opamp_dummy_magic_0.VD3.t24 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X788 two_stage_opamp_dummy_magic_0.VOUT-.t156 two_stage_opamp_dummy_magic_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_0.V_TOP.n0 bgr_0.V_TOP.t43 369.534
R1 bgr_0.V_TOP.n11 bgr_0.V_TOP.n9 339.961
R2 bgr_0.V_TOP.n11 bgr_0.V_TOP.n10 339.272
R3 bgr_0.V_TOP.n7 bgr_0.V_TOP.n6 339.272
R4 bgr_0.V_TOP.n15 bgr_0.V_TOP.n14 339.272
R5 bgr_0.V_TOP.n17 bgr_0.V_TOP.n16 339.272
R6 bgr_0.V_TOP.n12 bgr_0.V_TOP.n8 334.772
R7 bgr_0.V_TOP.n27 bgr_0.V_TOP.n26 224.934
R8 bgr_0.V_TOP.n26 bgr_0.V_TOP.n25 224.934
R9 bgr_0.V_TOP.n25 bgr_0.V_TOP.n24 224.934
R10 bgr_0.V_TOP.n24 bgr_0.V_TOP.n23 224.934
R11 bgr_0.V_TOP.n23 bgr_0.V_TOP.n22 224.934
R12 bgr_0.V_TOP.n22 bgr_0.V_TOP.n21 224.934
R13 bgr_0.V_TOP.n21 bgr_0.V_TOP.n20 224.934
R14 bgr_0.V_TOP.n1 bgr_0.V_TOP.n0 224.934
R15 bgr_0.V_TOP.n2 bgr_0.V_TOP.n1 224.934
R16 bgr_0.V_TOP.n3 bgr_0.V_TOP.n2 224.934
R17 bgr_0.V_TOP.n4 bgr_0.V_TOP.n3 224.934
R18 bgr_0.V_TOP.n5 bgr_0.V_TOP.n4 224.934
R19 bgr_0.V_TOP bgr_0.V_TOP.t32 214.222
R20 bgr_0.V_TOP bgr_0.V_TOP.n40 205.502
R21 bgr_0.V_TOP.n7 bgr_0.V_TOP.t3 176.114
R22 bgr_0.V_TOP.n19 bgr_0.V_TOP.n18 163.175
R23 bgr_0.V_TOP.n27 bgr_0.V_TOP.t31 144.601
R24 bgr_0.V_TOP.n26 bgr_0.V_TOP.t44 144.601
R25 bgr_0.V_TOP.n25 bgr_0.V_TOP.t18 144.601
R26 bgr_0.V_TOP.n24 bgr_0.V_TOP.t26 144.601
R27 bgr_0.V_TOP.n23 bgr_0.V_TOP.t37 144.601
R28 bgr_0.V_TOP.n22 bgr_0.V_TOP.t35 144.601
R29 bgr_0.V_TOP.n21 bgr_0.V_TOP.t48 144.601
R30 bgr_0.V_TOP.n20 bgr_0.V_TOP.t20 144.601
R31 bgr_0.V_TOP.n0 bgr_0.V_TOP.t29 144.601
R32 bgr_0.V_TOP.n1 bgr_0.V_TOP.t23 144.601
R33 bgr_0.V_TOP.n2 bgr_0.V_TOP.t14 144.601
R34 bgr_0.V_TOP.n3 bgr_0.V_TOP.t38 144.601
R35 bgr_0.V_TOP.n4 bgr_0.V_TOP.t41 144.601
R36 bgr_0.V_TOP.n5 bgr_0.V_TOP.t27 144.601
R37 bgr_0.V_TOP.n18 bgr_0.V_TOP.t12 95.4466
R38 bgr_0.V_TOP bgr_0.V_TOP.n27 69.6227
R39 bgr_0.V_TOP.n20 bgr_0.V_TOP.n19 69.6227
R40 bgr_0.V_TOP.n19 bgr_0.V_TOP.n5 69.6227
R41 bgr_0.V_TOP.n6 bgr_0.V_TOP.t2 39.4005
R42 bgr_0.V_TOP.n6 bgr_0.V_TOP.t6 39.4005
R43 bgr_0.V_TOP.n8 bgr_0.V_TOP.t11 39.4005
R44 bgr_0.V_TOP.n8 bgr_0.V_TOP.t7 39.4005
R45 bgr_0.V_TOP.n10 bgr_0.V_TOP.t13 39.4005
R46 bgr_0.V_TOP.n10 bgr_0.V_TOP.t4 39.4005
R47 bgr_0.V_TOP.n9 bgr_0.V_TOP.t1 39.4005
R48 bgr_0.V_TOP.n9 bgr_0.V_TOP.t0 39.4005
R49 bgr_0.V_TOP.n14 bgr_0.V_TOP.t9 39.4005
R50 bgr_0.V_TOP.n14 bgr_0.V_TOP.t8 39.4005
R51 bgr_0.V_TOP.n16 bgr_0.V_TOP.t10 39.4005
R52 bgr_0.V_TOP.n16 bgr_0.V_TOP.t5 39.4005
R53 bgr_0.V_TOP.n12 bgr_0.V_TOP.n11 8.313
R54 bgr_0.V_TOP.n18 bgr_0.V_TOP.n17 5.188
R55 bgr_0.V_TOP.n28 bgr_0.V_TOP.t49 4.8295
R56 bgr_0.V_TOP.n29 bgr_0.V_TOP.t25 4.8295
R57 bgr_0.V_TOP.n31 bgr_0.V_TOP.t21 4.8295
R58 bgr_0.V_TOP.n32 bgr_0.V_TOP.t34 4.8295
R59 bgr_0.V_TOP.n34 bgr_0.V_TOP.t30 4.8295
R60 bgr_0.V_TOP.n35 bgr_0.V_TOP.t46 4.8295
R61 bgr_0.V_TOP.n37 bgr_0.V_TOP.t24 4.8295
R62 bgr_0.V_TOP.n28 bgr_0.V_TOP.t39 4.5005
R63 bgr_0.V_TOP.n30 bgr_0.V_TOP.t28 4.5005
R64 bgr_0.V_TOP.n29 bgr_0.V_TOP.t33 4.5005
R65 bgr_0.V_TOP.n31 bgr_0.V_TOP.t15 4.5005
R66 bgr_0.V_TOP.n33 bgr_0.V_TOP.t40 4.5005
R67 bgr_0.V_TOP.n32 bgr_0.V_TOP.t45 4.5005
R68 bgr_0.V_TOP.n34 bgr_0.V_TOP.t22 4.5005
R69 bgr_0.V_TOP.n36 bgr_0.V_TOP.t16 4.5005
R70 bgr_0.V_TOP.n35 bgr_0.V_TOP.t19 4.5005
R71 bgr_0.V_TOP.n37 bgr_0.V_TOP.t17 4.5005
R72 bgr_0.V_TOP.n38 bgr_0.V_TOP.t42 4.5005
R73 bgr_0.V_TOP.n39 bgr_0.V_TOP.t47 4.5005
R74 bgr_0.V_TOP.n40 bgr_0.V_TOP.t36 4.5005
R75 bgr_0.V_TOP.n13 bgr_0.V_TOP.n12 4.5005
R76 bgr_0.V_TOP.n17 bgr_0.V_TOP.n15 2.1255
R77 bgr_0.V_TOP.n15 bgr_0.V_TOP.n13 2.1255
R78 bgr_0.V_TOP.n13 bgr_0.V_TOP.n7 2.1255
R79 bgr_0.V_TOP.n30 bgr_0.V_TOP.n28 0.3295
R80 bgr_0.V_TOP.n30 bgr_0.V_TOP.n29 0.3295
R81 bgr_0.V_TOP.n33 bgr_0.V_TOP.n31 0.3295
R82 bgr_0.V_TOP.n33 bgr_0.V_TOP.n32 0.3295
R83 bgr_0.V_TOP.n36 bgr_0.V_TOP.n34 0.3295
R84 bgr_0.V_TOP.n36 bgr_0.V_TOP.n35 0.3295
R85 bgr_0.V_TOP.n38 bgr_0.V_TOP.n37 0.3295
R86 bgr_0.V_TOP.n39 bgr_0.V_TOP.n38 0.3295
R87 bgr_0.V_TOP.n40 bgr_0.V_TOP.n39 0.3295
R88 bgr_0.V_TOP.n33 bgr_0.V_TOP.n30 0.2825
R89 bgr_0.V_TOP.n36 bgr_0.V_TOP.n33 0.2825
R90 bgr_0.V_TOP.n38 bgr_0.V_TOP.n36 0.2825
R91 bgr_0.Vin-.n14 bgr_0.Vin-.t10 688.859
R92 bgr_0.Vin-.n16 bgr_0.Vin-.n15 514.134
R93 bgr_0.Vin-.n12 bgr_0.Vin-.n11 345.115
R94 bgr_0.Vin-.n18 bgr_0.Vin-.n17 214.713
R95 bgr_0.Vin-.n14 bgr_0.Vin-.t12 174.726
R96 bgr_0.Vin-.n15 bgr_0.Vin-.t8 174.726
R97 bgr_0.Vin-.n16 bgr_0.Vin-.t11 174.726
R98 bgr_0.Vin-.n17 bgr_0.Vin-.t9 174.726
R99 bgr_0.Vin-.n10 bgr_0.Vin-.n8 173.029
R100 bgr_0.Vin-.n10 bgr_0.Vin-.n9 168.654
R101 bgr_0.Vin-.n12 bgr_0.Vin-.t1 162.921
R102 bgr_0.Vin-.n15 bgr_0.Vin-.n14 128.534
R103 bgr_0.Vin-.n17 bgr_0.Vin-.n16 128.534
R104 bgr_0.Vin-.n5 bgr_0.Vin-.n4 83.5719
R105 bgr_0.Vin-.n3 bgr_0.Vin-.n0 83.5719
R106 bgr_0.Vin-.n3 bgr_0.Vin-.n1 73.3165
R107 bgr_0.Vin-.t2 bgr_0.Vin-.n2 65.0341
R108 bgr_0.Vin-.n11 bgr_0.Vin-.t0 39.4005
R109 bgr_0.Vin-.n11 bgr_0.Vin-.t7 39.4005
R110 bgr_0.Vin-.n4 bgr_0.Vin-.n3 26.074
R111 bgr_0.Vin-.n19 bgr_0.Vin-.n18 17.526
R112 bgr_0.Vin-.n9 bgr_0.Vin-.t4 13.1338
R113 bgr_0.Vin-.n9 bgr_0.Vin-.t5 13.1338
R114 bgr_0.Vin-.n8 bgr_0.Vin-.t3 13.1338
R115 bgr_0.Vin-.n8 bgr_0.Vin-.t6 13.1338
R116 bgr_0.Vin-.n18 bgr_0.Vin-.n13 12.5317
R117 bgr_0.Vin-.n13 bgr_0.Vin-.n12 6.40675
R118 bgr_0.Vin-.n13 bgr_0.Vin-.n10 3.8755
R119 bgr_0.Vin-.n19 bgr_0.Vin-.n1 2.19742
R120 bgr_0.Vin-.n5 bgr_0.Vin-.n2 1.56483
R121 bgr_0.Vin-.n21 bgr_0.Vin-.n20 1.5505
R122 bgr_0.Vin-.n7 bgr_0.Vin-.n6 1.5505
R123 bgr_0.Vin-.n21 bgr_0.Vin-.n1 1.19225
R124 bgr_0.Vin-.n6 bgr_0.Vin-.n0 0.885803
R125 bgr_0.Vin-.n6 bgr_0.Vin-.n5 0.77514
R126 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n0 0.756696
R127 bgr_0.Vin-.n7 bgr_0.Vin-.n2 0.539177
R128 bgr_0.Vin-.n4 bgr_0.Vin-.t2 0.290206
R129 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter bgr_0.Vin-.n21 0.203382
R130 bgr_0.Vin-.n20 bgr_0.Vin-.n7 0.0183571
R131 bgr_0.Vin-.n20 bgr_0.Vin-.n19 0.0183571
R132 VDDA.n376 VDDA.n343 6600
R133 VDDA.n378 VDDA.n343 6600
R134 VDDA.n378 VDDA.n344 6570
R135 VDDA.n376 VDDA.n344 6570
R136 VDDA.n331 VDDA.n266 4710
R137 VDDA.n331 VDDA.n267 4710
R138 VDDA.n333 VDDA.n266 4710
R139 VDDA.n333 VDDA.n267 4710
R140 VDDA.n289 VDDA.n288 4710
R141 VDDA.n291 VDDA.n288 4710
R142 VDDA.n289 VDDA.n282 4710
R143 VDDA.n291 VDDA.n282 4710
R144 VDDA.n143 VDDA.n129 4605
R145 VDDA.n145 VDDA.n129 4605
R146 VDDA.n69 VDDA.n65 4605
R147 VDDA.n69 VDDA.n66 4605
R148 VDDA.n179 VDDA.n175 4590
R149 VDDA.n179 VDDA.n176 4590
R150 VDDA.n181 VDDA.n176 4590
R151 VDDA.n181 VDDA.n175 4590
R152 VDDA.n143 VDDA.n130 4575
R153 VDDA.n145 VDDA.n130 4575
R154 VDDA.n71 VDDA.n65 4575
R155 VDDA.n71 VDDA.n66 4575
R156 VDDA.n205 VDDA.n198 4020
R157 VDDA.n207 VDDA.n198 4020
R158 VDDA.n205 VDDA.n204 4020
R159 VDDA.n207 VDDA.n204 4020
R160 VDDA.n93 VDDA.n86 4020
R161 VDDA.n95 VDDA.n86 4020
R162 VDDA.n93 VDDA.n92 4020
R163 VDDA.n95 VDDA.n92 4020
R164 VDDA.n442 VDDA.n410 3420
R165 VDDA.n444 VDDA.n410 3420
R166 VDDA.n444 VDDA.n411 3420
R167 VDDA.n442 VDDA.n411 3420
R168 VDDA.n122 VDDA.n115 3390
R169 VDDA.n124 VDDA.n115 3390
R170 VDDA.n122 VDDA.n121 3390
R171 VDDA.n124 VDDA.n121 3390
R172 VDDA.n49 VDDA.n42 3390
R173 VDDA.n51 VDDA.n42 3390
R174 VDDA.n49 VDDA.n48 3390
R175 VDDA.n51 VDDA.n48 3390
R176 VDDA.n23 VDDA.n17 2940
R177 VDDA.n25 VDDA.n17 2940
R178 VDDA.n25 VDDA.n22 2940
R179 VDDA.n23 VDDA.n22 2940
R180 VDDA.n31 VDDA.n12 2940
R181 VDDA.n33 VDDA.n12 2940
R182 VDDA.n33 VDDA.n30 2940
R183 VDDA.n31 VDDA.n30 2940
R184 VDDA.n235 VDDA.n224 2415
R185 VDDA.n232 VDDA.n225 2400
R186 VDDA.n235 VDDA.n225 2370
R187 VDDA.n458 VDDA.n404 2145
R188 VDDA.n232 VDDA.n224 2115
R189 VDDA.n458 VDDA.n405 2100
R190 VDDA.n455 VDDA.n405 2100
R191 VDDA.n423 VDDA.n416 2100
R192 VDDA.n425 VDDA.n416 2100
R193 VDDA.n425 VDDA.n417 2100
R194 VDDA.n423 VDDA.n417 2100
R195 VDDA.n455 VDDA.n404 2055
R196 VDDA.n391 VDDA.n389 1770
R197 VDDA.n393 VDDA.n389 1770
R198 VDDA.n391 VDDA.n386 1770
R199 VDDA.n393 VDDA.n386 1770
R200 VDDA.n352 VDDA.n350 1770
R201 VDDA.n354 VDDA.n350 1770
R202 VDDA.n352 VDDA.n347 1770
R203 VDDA.n354 VDDA.n347 1770
R204 VDDA.n247 VDDA.n220 1575
R205 VDDA.n246 VDDA.n220 1575
R206 VDDA.n246 VDDA.n219 1545
R207 VDDA.n247 VDDA.n219 1545
R208 VDDA.n140 VDDA.t347 1216.42
R209 VDDA.n148 VDDA.t380 1216.42
R210 VDDA.n63 VDDA.t353 1216.42
R211 VDDA.n74 VDDA.t325 1216.42
R212 VDDA.n375 VDDA.n342 704
R213 VDDA.n379 VDDA.n342 704
R214 VDDA.n19 VDDA.t364 689.4
R215 VDDA.n18 VDDA.t391 689.4
R216 VDDA.n14 VDDA.t430 689.4
R217 VDDA.n13 VDDA.t321 689.4
R218 VDDA.n172 VDDA.t406 663.801
R219 VDDA.n185 VDDA.t412 663.801
R220 VDDA.n201 VDDA.t368 660.109
R221 VDDA.n199 VDDA.t395 660.109
R222 VDDA.n89 VDDA.t374 660.109
R223 VDDA.n87 VDDA.t419 660.109
R224 VDDA.n444 VDDA.t417 652.576
R225 VDDA.n242 VDDA.t330 647.54
R226 VDDA.n251 VDDA.t346 647.54
R227 VDDA.n216 VDDA.n215 631.654
R228 VDDA.n152 VDDA.n151 626.534
R229 VDDA.n155 VDDA.n154 626.534
R230 VDDA.n157 VDDA.n156 626.534
R231 VDDA.n159 VDDA.n158 626.534
R232 VDDA.n161 VDDA.n160 626.534
R233 VDDA.n163 VDDA.n162 626.534
R234 VDDA.n165 VDDA.n164 626.534
R235 VDDA.n167 VDDA.n166 626.534
R236 VDDA.n169 VDDA.n168 626.534
R237 VDDA.n171 VDDA.n170 626.534
R238 VDDA.n229 VDDA.t377 623.958
R239 VDDA.n238 VDDA.t398 623.958
R240 VDDA.t377 VDDA.n228 615.926
R241 VDDA.n118 VDDA.t359 573.75
R242 VDDA.n116 VDDA.t386 573.75
R243 VDDA.n45 VDDA.t331 573.75
R244 VDDA.n43 VDDA.t365 573.75
R245 VDDA.n374 VDDA.n341 518.4
R246 VDDA.n380 VDDA.n341 518.4
R247 VDDA.n293 VDDA.n292 496
R248 VDDA.n293 VDDA.n281 496
R249 VDDA.n146 VDDA.n128 491.2
R250 VDDA.n142 VDDA.n128 491.2
R251 VDDA.n68 VDDA.n40 491.2
R252 VDDA.n68 VDDA.n67 491.2
R253 VDDA.n178 VDDA.n153 489.601
R254 VDDA.n178 VDDA.n177 489.601
R255 VDDA.n209 VDDA.n208 428.8
R256 VDDA.n209 VDDA.n197 428.8
R257 VDDA.n97 VDDA.n96 428.8
R258 VDDA.n97 VDDA.n85 428.8
R259 VDDA.n387 VDDA.t334 419.108
R260 VDDA.n384 VDDA.t337 419.108
R261 VDDA.n348 VDDA.t413 413.084
R262 VDDA.n345 VDDA.t392 413.084
R263 VDDA.n452 VDDA.t401 409.067
R264 VDDA.n461 VDDA.t340 409.067
R265 VDDA.n439 VDDA.t422 409.067
R266 VDDA.n447 VDDA.t416 409.067
R267 VDDA.n420 VDDA.t316 409.067
R268 VDDA.n428 VDDA.t383 390.322
R269 VDDA.t411 VDDA.n175 389.375
R270 VDDA.t405 VDDA.n176 389.375
R271 VDDA.t429 VDDA.n30 389.375
R272 VDDA.t320 VDDA.n12 389.375
R273 VDDA.n387 VDDA.t336 389.185
R274 VDDA.n384 VDDA.t339 389.185
R275 VDDA.n183 VDDA.n182 387.2
R276 VDDA.n182 VDDA.n174 387.2
R277 VDDA.n439 VDDA.t424 387.051
R278 VDDA.n447 VDDA.t418 387.051
R279 VDDA.n264 VDDA.t358 384.918
R280 VDDA.n268 VDDA.t324 384.918
R281 VDDA.n283 VDDA.t373 384.918
R282 VDDA.n285 VDDA.t427 384.918
R283 VDDA.n348 VDDA.t415 384.918
R284 VDDA.n345 VDDA.t394 384.918
R285 VDDA.t363 VDDA.n22 384.168
R286 VDDA.t390 VDDA.n17 384.168
R287 VDDA.n270 VDDA.n269 384
R288 VDDA.n269 VDDA.n265 384
R289 VDDA.n287 VDDA.n286 384
R290 VDDA.n287 VDDA.n284 384
R291 VDDA.n420 VDDA.t318 370.728
R292 VDDA.n428 VDDA.t385 370.728
R293 VDDA.n452 VDDA.t403 370.3
R294 VDDA.n461 VDDA.t342 370.3
R295 VDDA.n441 VDDA.n409 364.8
R296 VDDA.n445 VDDA.n409 364.8
R297 VDDA.n373 VDDA.t350 360.868
R298 VDDA.n381 VDDA.t407 360.868
R299 VDDA.n264 VDDA.t356 358.858
R300 VDDA.n268 VDDA.t322 358.858
R301 VDDA.n283 VDDA.t371 358.858
R302 VDDA.n285 VDDA.t425 358.858
R303 VDDA.n126 VDDA.n125 355.2
R304 VDDA.n126 VDDA.n114 355.2
R305 VDDA.n53 VDDA.n52 355.2
R306 VDDA.n53 VDDA.n41 355.2
R307 VDDA.t323 VDDA.n331 351.591
R308 VDDA.n333 VDDA.t357 351.591
R309 VDDA.t426 VDDA.n289 351.591
R310 VDDA.n291 VDDA.t372 351.591
R311 VDDA.t329 VDDA.n246 346.668
R312 VDDA.n247 VDDA.t344 346.668
R313 VDDA.n413 VDDA.n412 345.127
R314 VDDA.n419 VDDA.n418 345.127
R315 VDDA.n401 VDDA.n400 344.7
R316 VDDA.n450 VDDA.n449 344.7
R317 VDDA.t338 VDDA.n391 344.394
R318 VDDA.n393 VDDA.t335 344.394
R319 VDDA.t393 VDDA.n352 344.394
R320 VDDA.n354 VDDA.t414 344.394
R321 VDDA.t402 VDDA.n455 344.394
R322 VDDA.n458 VDDA.t341 344.394
R323 VDDA.n275 VDDA.n273 342.3
R324 VDDA.n303 VDDA.n302 341.675
R325 VDDA.n301 VDDA.n300 341.675
R326 VDDA.n299 VDDA.n298 341.675
R327 VDDA.n297 VDDA.n296 341.675
R328 VDDA.n279 VDDA.n278 341.675
R329 VDDA.n277 VDDA.n276 341.675
R330 VDDA.n275 VDDA.n274 341.675
R331 VDDA.t423 VDDA.n442 340.635
R332 VDDA.t317 VDDA.n423 340.635
R333 VDDA.n425 VDDA.t384 340.635
R334 VDDA.n407 VDDA.n406 339.272
R335 VDDA.n431 VDDA.n430 339.272
R336 VDDA.n433 VDDA.n432 339.272
R337 VDDA.n435 VDDA.n434 339.272
R338 VDDA.n437 VDDA.n436 339.272
R339 VDDA.n336 VDDA.n260 337.175
R340 VDDA.n262 VDDA.n261 337.175
R341 VDDA.n312 VDDA.n311 337.175
R342 VDDA.n315 VDDA.n309 337.175
R343 VDDA.n307 VDDA.n306 337.175
R344 VDDA.n319 VDDA.n318 337.175
R345 VDDA.n322 VDDA.n305 337.175
R346 VDDA.n325 VDDA.n324 337.175
R347 VDDA.n328 VDDA.n272 337.175
R348 VDDA.n294 VDDA.n280 337.175
R349 VDDA.n397 VDDA.n383 335.022
R350 VDDA.n173 VDDA.t404 332.75
R351 VDDA.n184 VDDA.t410 332.75
R352 VDDA.n19 VDDA.t362 332.75
R353 VDDA.n18 VDDA.t389 332.75
R354 VDDA.n14 VDDA.t428 332.75
R355 VDDA.n13 VDDA.t319 332.75
R356 VDDA.n243 VDDA.t328 314.274
R357 VDDA.n250 VDDA.t343 314.274
R358 VDDA.n21 VDDA.n16 313.601
R359 VDDA.n28 VDDA.n16 307.2
R360 VDDA.n36 VDDA.n11 307.2
R361 VDDA.n29 VDDA.n11 307.2
R362 VDDA.t360 VDDA.n122 285.815
R363 VDDA.n124 VDDA.t387 285.815
R364 VDDA.t332 VDDA.n49 285.815
R365 VDDA.n51 VDDA.t366 285.815
R366 VDDA.t351 VDDA.n376 278.95
R367 VDDA.n378 VDDA.t408 278.95
R368 VDDA.n118 VDDA.t361 277.916
R369 VDDA.n116 VDDA.t388 277.916
R370 VDDA.n45 VDDA.t333 277.916
R371 VDDA.n43 VDDA.t367 277.916
R372 VDDA.n147 VDDA.n146 276.8
R373 VDDA.n142 VDDA.n141 276.8
R374 VDDA.n73 VDDA.n40 276.8
R375 VDDA.n67 VDDA.n64 276.8
R376 VDDA.n373 VDDA.t352 270.705
R377 VDDA.n381 VDDA.t409 270.705
R378 VDDA.n236 VDDA.n223 257.601
R379 VDDA.n440 VDDA.n408 246.4
R380 VDDA.t369 VDDA.n205 239.915
R381 VDDA.n207 VDDA.t396 239.915
R382 VDDA.t375 VDDA.n93 239.915
R383 VDDA.n95 VDDA.t420 239.915
R384 VDDA.n203 VDDA.n202 230.4
R385 VDDA.n203 VDDA.n200 230.4
R386 VDDA.n91 VDDA.n90 230.4
R387 VDDA.n91 VDDA.n88 230.4
R388 VDDA.n459 VDDA.n403 228.8
R389 VDDA.n231 VDDA.n223 225.601
R390 VDDA.n422 VDDA.n415 224
R391 VDDA.n426 VDDA.n415 224
R392 VDDA.n454 VDDA.n403 219.201
R393 VDDA.n120 VDDA.n119 211.201
R394 VDDA.n120 VDDA.n117 211.201
R395 VDDA.n47 VDDA.n46 211.201
R396 VDDA.n47 VDDA.n44 211.201
R397 VDDA.n26 VDDA.n20 211.201
R398 VDDA.n27 VDDA.n26 211.201
R399 VDDA.n35 VDDA.n34 211.201
R400 VDDA.n231 VDDA.n230 204.8
R401 VDDA.n141 VDDA.n127 204.8
R402 VDDA.n147 VDDA.n127 204.8
R403 VDDA.n73 VDDA.n72 204.8
R404 VDDA.n72 VDDA.n64 204.8
R405 VDDA.n34 VDDA.n15 202.971
R406 VDDA.n208 VDDA.n200 198.4
R407 VDDA.n202 VDDA.n197 198.4
R408 VDDA.n96 VDDA.n88 198.4
R409 VDDA.n90 VDDA.n85 198.4
R410 VDDA.t62 VDDA.t329 190
R411 VDDA.t344 VDDA.t62 190
R412 VDDA.n237 VDDA.n236 188.8
R413 VDDA.n335 VDDA.n334 188.8
R414 VDDA.n330 VDDA.n329 188.8
R415 VDDA.n394 VDDA.n388 188.8
R416 VDDA.n390 VDDA.n388 188.8
R417 VDDA.n355 VDDA.n349 188.8
R418 VDDA.n351 VDDA.n349 188.8
R419 VDDA.n446 VDDA.n445 188.8
R420 VDDA.t153 VDDA.t411 186.607
R421 VDDA.t165 VDDA.t153 186.607
R422 VDDA.t161 VDDA.t165 186.607
R423 VDDA.t94 VDDA.t161 186.607
R424 VDDA.t148 VDDA.t94 186.607
R425 VDDA.t155 VDDA.t148 186.607
R426 VDDA.t90 VDDA.t155 186.607
R427 VDDA.t96 VDDA.t90 186.607
R428 VDDA.t66 VDDA.t96 186.607
R429 VDDA.t151 VDDA.t66 186.607
R430 VDDA.t92 VDDA.t98 186.607
R431 VDDA.t98 VDDA.t22 186.607
R432 VDDA.t22 VDDA.t146 186.607
R433 VDDA.t146 VDDA.t167 186.607
R434 VDDA.t167 VDDA.t88 186.607
R435 VDDA.t88 VDDA.t157 186.607
R436 VDDA.t157 VDDA.t64 186.607
R437 VDDA.t64 VDDA.t163 186.607
R438 VDDA.t163 VDDA.t24 186.607
R439 VDDA.t24 VDDA.t405 186.607
R440 VDDA.t249 VDDA.t429 186.607
R441 VDDA.t27 VDDA.t249 186.607
R442 VDDA.t150 VDDA.t27 186.607
R443 VDDA.t251 VDDA.t150 186.607
R444 VDDA.t262 VDDA.t251 186.607
R445 VDDA.t443 VDDA.t257 186.607
R446 VDDA.t257 VDDA.t252 186.607
R447 VDDA.t252 VDDA.t248 186.607
R448 VDDA.t248 VDDA.t103 186.607
R449 VDDA.t103 VDDA.t320 186.607
R450 VDDA.t263 VDDA.t363 183.333
R451 VDDA.t48 VDDA.t263 183.333
R452 VDDA.t59 VDDA.t48 183.333
R453 VDDA.t86 VDDA.t59 183.333
R454 VDDA.t253 VDDA.t86 183.333
R455 VDDA.t68 VDDA.t45 183.333
R456 VDDA.t45 VDDA.t87 183.333
R457 VDDA.t87 VDDA.t250 183.333
R458 VDDA.t250 VDDA.t43 183.333
R459 VDDA.t43 VDDA.t390 183.333
R460 VDDA.n375 VDDA.n374 182.4
R461 VDDA.n380 VDDA.n379 182.4
R462 VDDA.n139 VDDA.t349 178.124
R463 VDDA.n149 VDDA.t382 178.124
R464 VDDA.n62 VDDA.t355 178.124
R465 VDDA.n75 VDDA.t327 178.124
R466 VDDA.n446 VDDA.n408 176
R467 VDDA.n226 VDDA.n221 174.393
R468 VDDA.t465 VDDA.t323 172.727
R469 VDDA.t226 VDDA.t465 172.727
R470 VDDA.t133 VDDA.t226 172.727
R471 VDDA.t242 VDDA.t133 172.727
R472 VDDA.t246 VDDA.t242 172.727
R473 VDDA.t238 VDDA.t246 172.727
R474 VDDA.t6 VDDA.t238 172.727
R475 VDDA.t51 VDDA.t6 172.727
R476 VDDA.t224 VDDA.t51 172.727
R477 VDDA.t104 VDDA.t461 172.727
R478 VDDA.t459 VDDA.t104 172.727
R479 VDDA.t37 VDDA.t459 172.727
R480 VDDA.t131 VDDA.t37 172.727
R481 VDDA.t49 VDDA.t131 172.727
R482 VDDA.t201 VDDA.t49 172.727
R483 VDDA.t244 VDDA.t201 172.727
R484 VDDA.t60 VDDA.t244 172.727
R485 VDDA.t357 VDDA.t60 172.727
R486 VDDA.t431 VDDA.t426 172.727
R487 VDDA.t79 VDDA.t431 172.727
R488 VDDA.t106 VDDA.t79 172.727
R489 VDDA.t28 VDDA.t106 172.727
R490 VDDA.t2 VDDA.t28 172.727
R491 VDDA.t441 VDDA.t2 172.727
R492 VDDA.t433 VDDA.t441 172.727
R493 VDDA.t219 VDDA.t433 172.727
R494 VDDA.t81 VDDA.t219 172.727
R495 VDDA.t4 VDDA.t178 172.727
R496 VDDA.t437 VDDA.t4 172.727
R497 VDDA.t435 VDDA.t437 172.727
R498 VDDA.t217 VDDA.t435 172.727
R499 VDDA.t108 VDDA.t217 172.727
R500 VDDA.t180 VDDA.t108 172.727
R501 VDDA.t100 VDDA.t180 172.727
R502 VDDA.t439 VDDA.t100 172.727
R503 VDDA.t372 VDDA.t439 172.727
R504 VDDA.n235 VDDA.t399 172.554
R505 VDDA.t378 VDDA.n232 170.873
R506 VDDA.n340 VDDA.n339 168.435
R507 VDDA.n359 VDDA.n358 168.435
R508 VDDA.n361 VDDA.n360 168.435
R509 VDDA.n363 VDDA.n362 168.435
R510 VDDA.n365 VDDA.n364 168.435
R511 VDDA.n367 VDDA.n366 168.435
R512 VDDA.n369 VDDA.n368 168.435
R513 VDDA.n371 VDDA.n370 168.435
R514 VDDA.n245 VDDA.n218 164.8
R515 VDDA.n248 VDDA.n218 164.8
R516 VDDA.t348 VDDA.n143 161.817
R517 VDDA.n145 VDDA.t381 161.817
R518 VDDA.t326 VDDA.n65 161.817
R519 VDDA.t354 VDDA.n66 161.817
R520 VDDA.n195 VDDA.n193 160.428
R521 VDDA.n192 VDDA.n190 160.428
R522 VDDA.n83 VDDA.n81 160.428
R523 VDDA.n80 VDDA.n78 160.428
R524 VDDA.t272 VDDA.t351 159.814
R525 VDDA.t293 VDDA.t272 159.814
R526 VDDA.t304 VDDA.t293 159.814
R527 VDDA.t314 VDDA.t304 159.814
R528 VDDA.t279 VDDA.t314 159.814
R529 VDDA.t275 VDDA.t279 159.814
R530 VDDA.t298 VDDA.t275 159.814
R531 VDDA.t306 VDDA.t298 159.814
R532 VDDA.t284 VDDA.t265 159.814
R533 VDDA.t281 VDDA.t284 159.814
R534 VDDA.t300 VDDA.t281 159.814
R535 VDDA.t309 VDDA.t300 159.814
R536 VDDA.t270 VDDA.t309 159.814
R537 VDDA.t290 VDDA.t270 159.814
R538 VDDA.t288 VDDA.t290 159.814
R539 VDDA.t408 VDDA.t288 159.814
R540 VDDA.n195 VDDA.n194 159.803
R541 VDDA.n192 VDDA.n191 159.803
R542 VDDA.n83 VDDA.n82 159.803
R543 VDDA.n80 VDDA.n79 159.803
R544 VDDA.t71 VDDA.t338 158.333
R545 VDDA.t335 VDDA.t463 158.333
R546 VDDA.t36 VDDA.t393 158.333
R547 VDDA.t414 VDDA.t455 158.333
R548 VDDA.t75 VDDA.t402 158.333
R549 VDDA.t144 VDDA.t75 158.333
R550 VDDA.t159 VDDA.t197 158.333
R551 VDDA.t341 VDDA.t159 158.333
R552 VDDA.t447 VDDA.t423 155.97
R553 VDDA.t467 VDDA.t447 155.97
R554 VDDA.t451 VDDA.t467 155.97
R555 VDDA.t30 VDDA.t451 155.97
R556 VDDA.t453 VDDA.t30 155.97
R557 VDDA.t457 VDDA.t453 155.97
R558 VDDA.t174 VDDA.t176 155.97
R559 VDDA.t140 VDDA.t174 155.97
R560 VDDA.t215 VDDA.t140 155.97
R561 VDDA.t417 VDDA.t215 155.97
R562 VDDA.t199 VDDA.t317 155.97
R563 VDDA.t195 VDDA.t199 155.97
R564 VDDA.t213 VDDA.t142 155.97
R565 VDDA.t384 VDDA.t213 155.97
R566 VDDA.n201 VDDA.t370 155.125
R567 VDDA.n199 VDDA.t397 155.125
R568 VDDA.n89 VDDA.t376 155.125
R569 VDDA.n87 VDDA.t421 155.125
R570 VDDA.n139 VDDA.n138 151.882
R571 VDDA.n62 VDDA.n61 151.882
R572 VDDA.n150 VDDA.n149 151.321
R573 VDDA.n76 VDDA.n75 151.321
R574 VDDA.n125 VDDA.n117 150.4
R575 VDDA.n119 VDDA.n114 150.4
R576 VDDA.n52 VDDA.n44 150.4
R577 VDDA.n46 VDDA.n41 150.4
R578 VDDA.n211 VDDA.n210 146.002
R579 VDDA.n99 VDDA.n98 146.002
R580 VDDA.n113 VDDA.n112 145.429
R581 VDDA.n132 VDDA.n131 145.429
R582 VDDA.n134 VDDA.n133 145.429
R583 VDDA.n136 VDDA.n135 145.429
R584 VDDA.n138 VDDA.n137 145.429
R585 VDDA.n39 VDDA.n38 145.429
R586 VDDA.n55 VDDA.n54 145.429
R587 VDDA.n57 VDDA.n56 145.429
R588 VDDA.n59 VDDA.n58 145.429
R589 VDDA.n61 VDDA.n60 145.429
R590 VDDA.n149 VDDA.n148 135.387
R591 VDDA.n140 VDDA.n139 135.387
R592 VDDA.n75 VDDA.n74 135.387
R593 VDDA.n63 VDDA.n62 135.387
R594 VDDA.t182 VDDA.t360 121.513
R595 VDDA.t444 VDDA.t182 121.513
R596 VDDA.t221 VDDA.t444 121.513
R597 VDDA.t456 VDDA.t221 121.513
R598 VDDA.t113 VDDA.t456 121.513
R599 VDDA.t184 VDDA.t57 121.513
R600 VDDA.t56 VDDA.t184 121.513
R601 VDDA.t233 VDDA.t56 121.513
R602 VDDA.t26 VDDA.t233 121.513
R603 VDDA.t387 VDDA.t26 121.513
R604 VDDA.t10 VDDA.t332 121.513
R605 VDDA.t209 VDDA.t10 121.513
R606 VDDA.t119 VDDA.t209 121.513
R607 VDDA.t55 VDDA.t119 121.513
R608 VDDA.t125 VDDA.t55 121.513
R609 VDDA.t21 VDDA.t189 121.513
R610 VDDA.t187 VDDA.t21 121.513
R611 VDDA.t54 VDDA.t187 121.513
R612 VDDA.t255 VDDA.t54 121.513
R613 VDDA.t366 VDDA.t255 121.513
R614 VDDA.n334 VDDA.n265 118.4
R615 VDDA.n330 VDDA.n270 118.4
R616 VDDA.n292 VDDA.n284 118.4
R617 VDDA.n286 VDDA.n281 118.4
R618 VDDA.n395 VDDA.n394 118.4
R619 VDDA.n390 VDDA.n385 118.4
R620 VDDA.n356 VDDA.n355 118.4
R621 VDDA.n351 VDDA.n346 118.4
R622 VDDA.n454 VDDA.n453 118.4
R623 VDDA.n460 VDDA.n459 118.4
R624 VDDA.n441 VDDA.n440 118.4
R625 VDDA.n422 VDDA.n421 118.4
R626 VDDA.n427 VDDA.n426 118.4
R627 VDDA.n245 VDDA.n244 110.4
R628 VDDA.n249 VDDA.n248 110.4
R629 VDDA.n453 VDDA.n402 105.6
R630 VDDA.n460 VDDA.n402 105.6
R631 VDDA.n421 VDDA.n414 105.6
R632 VDDA.n427 VDDA.n414 105.6
R633 VDDA.t399 VDDA.t240 102.704
R634 VDDA.n183 VDDA.n153 102.4
R635 VDDA.n177 VDDA.n174 102.4
R636 VDDA.n21 VDDA.n20 102.4
R637 VDDA.n240 VDDA.n239 101.267
R638 VDDA.t234 VDDA.t369 98.2764
R639 VDDA.t0 VDDA.t234 98.2764
R640 VDDA.t230 VDDA.t0 98.2764
R641 VDDA.t8 VDDA.t230 98.2764
R642 VDDA.t260 VDDA.t8 98.2764
R643 VDDA.t203 VDDA.t445 98.2764
R644 VDDA.t77 VDDA.t203 98.2764
R645 VDDA.t39 VDDA.t77 98.2764
R646 VDDA.t228 VDDA.t39 98.2764
R647 VDDA.t396 VDDA.t228 98.2764
R648 VDDA.t236 VDDA.t375 98.2764
R649 VDDA.t135 VDDA.t236 98.2764
R650 VDDA.t32 VDDA.t135 98.2764
R651 VDDA.t110 VDDA.t32 98.2764
R652 VDDA.t449 VDDA.t110 98.2764
R653 VDDA.t205 VDDA.t172 98.2764
R654 VDDA.t258 VDDA.t205 98.2764
R655 VDDA.t207 VDDA.t258 98.2764
R656 VDDA.t69 VDDA.t207 98.2764
R657 VDDA.t420 VDDA.t69 98.2764
R658 VDDA.n103 VDDA.n101 97.4034
R659 VDDA.n2 VDDA.n0 97.4034
R660 VDDA.n111 VDDA.n110 96.8409
R661 VDDA.n109 VDDA.n108 96.8409
R662 VDDA.n107 VDDA.n106 96.8409
R663 VDDA.n105 VDDA.n104 96.8409
R664 VDDA.n103 VDDA.n102 96.8409
R665 VDDA.n10 VDDA.n9 96.8409
R666 VDDA.n8 VDDA.n7 96.8409
R667 VDDA.n6 VDDA.n5 96.8409
R668 VDDA.n4 VDDA.n3 96.8409
R669 VDDA.n2 VDDA.n1 96.8409
R670 VDDA.n28 VDDA.n27 96.0005
R671 VDDA.n29 VDDA.n15 96.0005
R672 VDDA.n36 VDDA.n35 96.0005
R673 VDDA.n180 VDDA.t151 93.3041
R674 VDDA.n180 VDDA.t92 93.3041
R675 VDDA.n32 VDDA.t262 93.3041
R676 VDDA.n32 VDDA.t443 93.3041
R677 VDDA.n219 VDDA.n218 92.5005
R678 VDDA.t62 VDDA.n219 92.5005
R679 VDDA.n220 VDDA.n217 92.5005
R680 VDDA.t62 VDDA.n220 92.5005
R681 VDDA.n224 VDDA.n223 92.5005
R682 VDDA.n233 VDDA.n224 92.5005
R683 VDDA.n225 VDDA.n222 92.5005
R684 VDDA.n234 VDDA.n225 92.5005
R685 VDDA.n208 VDDA.n207 92.5005
R686 VDDA.n204 VDDA.n203 92.5005
R687 VDDA.n206 VDDA.n204 92.5005
R688 VDDA.n205 VDDA.n197 92.5005
R689 VDDA.n209 VDDA.n198 92.5005
R690 VDDA.n206 VDDA.n198 92.5005
R691 VDDA.n175 VDDA.n153 92.5005
R692 VDDA.n179 VDDA.n178 92.5005
R693 VDDA.n180 VDDA.n179 92.5005
R694 VDDA.n177 VDDA.n176 92.5005
R695 VDDA.n182 VDDA.n181 92.5005
R696 VDDA.n181 VDDA.n180 92.5005
R697 VDDA.n125 VDDA.n124 92.5005
R698 VDDA.n121 VDDA.n120 92.5005
R699 VDDA.n123 VDDA.n121 92.5005
R700 VDDA.n122 VDDA.n114 92.5005
R701 VDDA.n126 VDDA.n115 92.5005
R702 VDDA.n123 VDDA.n115 92.5005
R703 VDDA.n130 VDDA.n127 92.5005
R704 VDDA.n144 VDDA.n130 92.5005
R705 VDDA.n129 VDDA.n128 92.5005
R706 VDDA.n144 VDDA.n129 92.5005
R707 VDDA.n96 VDDA.n95 92.5005
R708 VDDA.n92 VDDA.n91 92.5005
R709 VDDA.n94 VDDA.n92 92.5005
R710 VDDA.n93 VDDA.n85 92.5005
R711 VDDA.n97 VDDA.n86 92.5005
R712 VDDA.n94 VDDA.n86 92.5005
R713 VDDA.n52 VDDA.n51 92.5005
R714 VDDA.n48 VDDA.n47 92.5005
R715 VDDA.n50 VDDA.n48 92.5005
R716 VDDA.n49 VDDA.n41 92.5005
R717 VDDA.n53 VDDA.n42 92.5005
R718 VDDA.n50 VDDA.n42 92.5005
R719 VDDA.n72 VDDA.n71 92.5005
R720 VDDA.n71 VDDA.n70 92.5005
R721 VDDA.n69 VDDA.n68 92.5005
R722 VDDA.n70 VDDA.n69 92.5005
R723 VDDA.n23 VDDA.n16 92.5005
R724 VDDA.n24 VDDA.n23 92.5005
R725 VDDA.n22 VDDA.n21 92.5005
R726 VDDA.n26 VDDA.n25 92.5005
R727 VDDA.n25 VDDA.n24 92.5005
R728 VDDA.n28 VDDA.n17 92.5005
R729 VDDA.n31 VDDA.n11 92.5005
R730 VDDA.n32 VDDA.n31 92.5005
R731 VDDA.n30 VDDA.n29 92.5005
R732 VDDA.n34 VDDA.n33 92.5005
R733 VDDA.n33 VDDA.n32 92.5005
R734 VDDA.n36 VDDA.n12 92.5005
R735 VDDA.n317 VDDA.n267 92.5005
R736 VDDA.n332 VDDA.n267 92.5005
R737 VDDA.n334 VDDA.n333 92.5005
R738 VDDA.n269 VDDA.n266 92.5005
R739 VDDA.n332 VDDA.n266 92.5005
R740 VDDA.n331 VDDA.n330 92.5005
R741 VDDA.n292 VDDA.n291 92.5005
R742 VDDA.n288 VDDA.n287 92.5005
R743 VDDA.n290 VDDA.n288 92.5005
R744 VDDA.n289 VDDA.n281 92.5005
R745 VDDA.n293 VDDA.n282 92.5005
R746 VDDA.n290 VDDA.n282 92.5005
R747 VDDA.n394 VDDA.n393 92.5005
R748 VDDA.n389 VDDA.n388 92.5005
R749 VDDA.n392 VDDA.n389 92.5005
R750 VDDA.n391 VDDA.n390 92.5005
R751 VDDA.n396 VDDA.n386 92.5005
R752 VDDA.n392 VDDA.n386 92.5005
R753 VDDA.n376 VDDA.n375 92.5005
R754 VDDA.n343 VDDA.n342 92.5005
R755 VDDA.n377 VDDA.n343 92.5005
R756 VDDA.n379 VDDA.n378 92.5005
R757 VDDA.n344 VDDA.n341 92.5005
R758 VDDA.n377 VDDA.n344 92.5005
R759 VDDA.n355 VDDA.n354 92.5005
R760 VDDA.n350 VDDA.n349 92.5005
R761 VDDA.n353 VDDA.n350 92.5005
R762 VDDA.n352 VDDA.n351 92.5005
R763 VDDA.n357 VDDA.n347 92.5005
R764 VDDA.n353 VDDA.n347 92.5005
R765 VDDA.n455 VDDA.n454 92.5005
R766 VDDA.n404 VDDA.n403 92.5005
R767 VDDA.n456 VDDA.n404 92.5005
R768 VDDA.n459 VDDA.n458 92.5005
R769 VDDA.n405 VDDA.n402 92.5005
R770 VDDA.n457 VDDA.n405 92.5005
R771 VDDA.n442 VDDA.n441 92.5005
R772 VDDA.n410 VDDA.n409 92.5005
R773 VDDA.n443 VDDA.n410 92.5005
R774 VDDA.n445 VDDA.n444 92.5005
R775 VDDA.n411 VDDA.n408 92.5005
R776 VDDA.n443 VDDA.n411 92.5005
R777 VDDA.n423 VDDA.n422 92.5005
R778 VDDA.n416 VDDA.n415 92.5005
R779 VDDA.n424 VDDA.n416 92.5005
R780 VDDA.n426 VDDA.n425 92.5005
R781 VDDA.n417 VDDA.n414 92.5005
R782 VDDA.n424 VDDA.n417 92.5005
R783 VDDA.n24 VDDA.t253 91.6672
R784 VDDA.n24 VDDA.t68 91.6672
R785 VDDA.n228 VDDA.n227 87.4672
R786 VDDA.n332 VDDA.t224 86.3641
R787 VDDA.t461 VDDA.n332 86.3641
R788 VDDA.n290 VDDA.t81 86.3641
R789 VDDA.t178 VDDA.n290 86.3641
R790 VDDA.n227 VDDA.t379 85.438
R791 VDDA.n239 VDDA.t400 85.438
R792 VDDA.n233 VDDA.t378 81.3068
R793 VDDA.n239 VDDA.n238 81.0672
R794 VDDA.n229 VDDA.n227 81.0672
R795 VDDA.n377 VDDA.t306 79.907
R796 VDDA.t265 VDDA.n377 79.907
R797 VDDA.n392 VDDA.t71 79.1672
R798 VDDA.t463 VDDA.n392 79.1672
R799 VDDA.n353 VDDA.t36 79.1672
R800 VDDA.t455 VDDA.n353 79.1672
R801 VDDA.t197 VDDA.n457 79.1672
R802 VDDA.n151 VDDA.t154 78.8005
R803 VDDA.n151 VDDA.t166 78.8005
R804 VDDA.n154 VDDA.t162 78.8005
R805 VDDA.n154 VDDA.t95 78.8005
R806 VDDA.n156 VDDA.t149 78.8005
R807 VDDA.n156 VDDA.t156 78.8005
R808 VDDA.n158 VDDA.t91 78.8005
R809 VDDA.n158 VDDA.t97 78.8005
R810 VDDA.n160 VDDA.t67 78.8005
R811 VDDA.n160 VDDA.t152 78.8005
R812 VDDA.n162 VDDA.t93 78.8005
R813 VDDA.n162 VDDA.t99 78.8005
R814 VDDA.n164 VDDA.t23 78.8005
R815 VDDA.n164 VDDA.t147 78.8005
R816 VDDA.n166 VDDA.t168 78.8005
R817 VDDA.n166 VDDA.t89 78.8005
R818 VDDA.n168 VDDA.t158 78.8005
R819 VDDA.n168 VDDA.t65 78.8005
R820 VDDA.n170 VDDA.t164 78.8005
R821 VDDA.n170 VDDA.t25 78.8005
R822 VDDA.n443 VDDA.t457 77.9856
R823 VDDA.t176 VDDA.n443 77.9856
R824 VDDA.n424 VDDA.t195 77.9856
R825 VDDA.t142 VDDA.n424 77.9856
R826 VDDA.n237 VDDA.n222 64.0005
R827 VDDA.n329 VDDA.n271 64.0005
R828 VDDA.n321 VDDA.n271 64.0005
R829 VDDA.n321 VDDA.n320 64.0005
R830 VDDA.n320 VDDA.n317 64.0005
R831 VDDA.n317 VDDA.n316 64.0005
R832 VDDA.n316 VDDA.n308 64.0005
R833 VDDA.n308 VDDA.n263 64.0005
R834 VDDA.n335 VDDA.n263 64.0005
R835 VDDA.n357 VDDA.n356 64.0005
R836 VDDA.n357 VDDA.n346 64.0005
R837 VDDA.t170 VDDA.t348 62.9523
R838 VDDA.t73 VDDA.t170 62.9523
R839 VDDA.t222 VDDA.t73 62.9523
R840 VDDA.t193 VDDA.t222 62.9523
R841 VDDA.t128 VDDA.t193 62.9523
R842 VDDA.t16 VDDA.t41 62.9523
R843 VDDA.t46 VDDA.t16 62.9523
R844 VDDA.t84 VDDA.t46 62.9523
R845 VDDA.t114 VDDA.t84 62.9523
R846 VDDA.t381 VDDA.t114 62.9523
R847 VDDA.t122 VDDA.t326 62.9523
R848 VDDA.t210 VDDA.t122 62.9523
R849 VDDA.t120 VDDA.t210 62.9523
R850 VDDA.t13 VDDA.t120 62.9523
R851 VDDA.t19 VDDA.t13 62.9523
R852 VDDA.t185 VDDA.t138 62.9523
R853 VDDA.t138 VDDA.t116 62.9523
R854 VDDA.t116 VDDA.t11 62.9523
R855 VDDA.t11 VDDA.t126 62.9523
R856 VDDA.t126 VDDA.t354 62.9523
R857 VDDA.n396 VDDA.n395 62.7205
R858 VDDA.n396 VDDA.n385 62.7205
R859 VDDA.n215 VDDA.t63 62.5402
R860 VDDA.n215 VDDA.t345 62.5402
R861 VDDA.n246 VDDA.n245 61.6672
R862 VDDA.n248 VDDA.n247 61.6672
R863 VDDA.n146 VDDA.n145 61.6672
R864 VDDA.n143 VDDA.n142 61.6672
R865 VDDA.n65 VDDA.n40 61.6672
R866 VDDA.n67 VDDA.n66 61.6672
R867 VDDA.n123 VDDA.t113 60.7563
R868 VDDA.t57 VDDA.n123 60.7563
R869 VDDA.n50 VDDA.t125 60.7563
R870 VDDA.t189 VDDA.n50 60.7563
R871 VDDA.n256 VDDA.t471 59.5681
R872 VDDA.n255 VDDA.t469 59.5681
R873 VDDA.n244 VDDA.n217 57.6005
R874 VDDA.n249 VDDA.n217 57.6005
R875 VDDA.n456 VDDA.t144 57.5763
R876 VDDA.n255 VDDA.t472 51.8888
R877 VDDA.n230 VDDA.n222 51.2005
R878 VDDA.n206 VDDA.t260 49.1384
R879 VDDA.t445 VDDA.n206 49.1384
R880 VDDA.n94 VDDA.t449 49.1384
R881 VDDA.t172 VDDA.n94 49.1384
R882 VDDA.n257 VDDA.t470 48.9557
R883 VDDA.n252 VDDA.n251 46.6538
R884 VDDA.n242 VDDA.n241 42.1538
R885 VDDA.n172 VDDA.n171 42.0963
R886 VDDA.n186 VDDA.n185 41.5338
R887 VDDA.n260 VDDA.t245 39.4005
R888 VDDA.n260 VDDA.t61 39.4005
R889 VDDA.n261 VDDA.t50 39.4005
R890 VDDA.n261 VDDA.t202 39.4005
R891 VDDA.n311 VDDA.t38 39.4005
R892 VDDA.n311 VDDA.t132 39.4005
R893 VDDA.n309 VDDA.t105 39.4005
R894 VDDA.n309 VDDA.t460 39.4005
R895 VDDA.n306 VDDA.t225 39.4005
R896 VDDA.n306 VDDA.t462 39.4005
R897 VDDA.n318 VDDA.t7 39.4005
R898 VDDA.n318 VDDA.t52 39.4005
R899 VDDA.n305 VDDA.t247 39.4005
R900 VDDA.n305 VDDA.t239 39.4005
R901 VDDA.n324 VDDA.t134 39.4005
R902 VDDA.n324 VDDA.t243 39.4005
R903 VDDA.n272 VDDA.t466 39.4005
R904 VDDA.n272 VDDA.t227 39.4005
R905 VDDA.n302 VDDA.t101 39.4005
R906 VDDA.n302 VDDA.t440 39.4005
R907 VDDA.n300 VDDA.t109 39.4005
R908 VDDA.n300 VDDA.t181 39.4005
R909 VDDA.n298 VDDA.t436 39.4005
R910 VDDA.n298 VDDA.t218 39.4005
R911 VDDA.n296 VDDA.t5 39.4005
R912 VDDA.n296 VDDA.t438 39.4005
R913 VDDA.n280 VDDA.t82 39.4005
R914 VDDA.n280 VDDA.t179 39.4005
R915 VDDA.n278 VDDA.t434 39.4005
R916 VDDA.n278 VDDA.t220 39.4005
R917 VDDA.n276 VDDA.t3 39.4005
R918 VDDA.n276 VDDA.t442 39.4005
R919 VDDA.n274 VDDA.t107 39.4005
R920 VDDA.n274 VDDA.t29 39.4005
R921 VDDA.n273 VDDA.t432 39.4005
R922 VDDA.n273 VDDA.t80 39.4005
R923 VDDA.n383 VDDA.t72 39.4005
R924 VDDA.n383 VDDA.t464 39.4005
R925 VDDA.n400 VDDA.t198 39.4005
R926 VDDA.n400 VDDA.t160 39.4005
R927 VDDA.n449 VDDA.t76 39.4005
R928 VDDA.n449 VDDA.t145 39.4005
R929 VDDA.n406 VDDA.t141 39.4005
R930 VDDA.n406 VDDA.t216 39.4005
R931 VDDA.n430 VDDA.t177 39.4005
R932 VDDA.n430 VDDA.t175 39.4005
R933 VDDA.n432 VDDA.t454 39.4005
R934 VDDA.n432 VDDA.t458 39.4005
R935 VDDA.n434 VDDA.t452 39.4005
R936 VDDA.n434 VDDA.t31 39.4005
R937 VDDA.n436 VDDA.t448 39.4005
R938 VDDA.n436 VDDA.t468 39.4005
R939 VDDA.n412 VDDA.t143 39.4005
R940 VDDA.n412 VDDA.t214 39.4005
R941 VDDA.n418 VDDA.t200 39.4005
R942 VDDA.n418 VDDA.t196 39.4005
R943 VDDA.n144 VDDA.t128 31.4764
R944 VDDA.t41 VDDA.n144 31.4764
R945 VDDA.n70 VDDA.t19 31.4764
R946 VDDA.n70 VDDA.t185 31.4764
R947 VDDA.n29 VDDA.n28 28.663
R948 VDDA.n251 VDDA.n250 27.3072
R949 VDDA.n243 VDDA.n242 27.3072
R950 VDDA.n185 VDDA.n184 25.6005
R951 VDDA.n173 VDDA.n172 25.6005
R952 VDDA.n258 VDDA.n254 24.7453
R953 VDDA.n250 VDDA.n249 24.5338
R954 VDDA.n244 VDDA.n243 24.5338
R955 VDDA.n238 VDDA.n237 24.5338
R956 VDDA.n230 VDDA.n229 24.5338
R957 VDDA.n457 VDDA.n456 21.5914
R958 VDDA.n254 VDDA.n253 21.5392
R959 VDDA.n202 VDDA.n201 21.3338
R960 VDDA.n200 VDDA.n199 21.3338
R961 VDDA.n184 VDDA.n183 21.3338
R962 VDDA.n174 VDDA.n173 21.3338
R963 VDDA.n119 VDDA.n118 21.3338
R964 VDDA.n117 VDDA.n116 21.3338
R965 VDDA.n148 VDDA.n147 21.3338
R966 VDDA.n141 VDDA.n140 21.3338
R967 VDDA.n90 VDDA.n89 21.3338
R968 VDDA.n88 VDDA.n87 21.3338
R969 VDDA.n46 VDDA.n45 21.3338
R970 VDDA.n44 VDDA.n43 21.3338
R971 VDDA.n74 VDDA.n73 21.3338
R972 VDDA.n64 VDDA.n63 21.3338
R973 VDDA.n20 VDDA.n19 21.3338
R974 VDDA.n27 VDDA.n18 21.3338
R975 VDDA.n15 VDDA.n14 21.3338
R976 VDDA.n35 VDDA.n13 21.3338
R977 VDDA.n265 VDDA.n264 21.3338
R978 VDDA.n270 VDDA.n268 21.3338
R979 VDDA.n284 VDDA.n283 21.3338
R980 VDDA.n286 VDDA.n285 21.3338
R981 VDDA.n395 VDDA.n387 21.3338
R982 VDDA.n385 VDDA.n384 21.3338
R983 VDDA.n356 VDDA.n348 21.3338
R984 VDDA.n346 VDDA.n345 21.3338
R985 VDDA.n37 VDDA.n36 19.5505
R986 VDDA.n127 VDDA.n126 19.538
R987 VDDA.n72 VDDA.n53 19.538
R988 VDDA.n211 VDDA.n209 19.2005
R989 VDDA.n99 VDDA.n97 19.2005
R990 VDDA.n381 VDDA.n380 19.2005
R991 VDDA.n374 VDDA.n373 19.2005
R992 VDDA.n461 VDDA.n460 19.2005
R993 VDDA.n453 VDDA.n452 19.2005
R994 VDDA.n447 VDDA.n446 19.2005
R995 VDDA.n440 VDDA.n439 19.2005
R996 VDDA.n428 VDDA.n427 19.2005
R997 VDDA.n421 VDDA.n420 19.2005
R998 VDDA.n236 VDDA.n235 18.5005
R999 VDDA.t240 VDDA.n234 17.1176
R1000 VDDA.n188 VDDA.n111 16.8443
R1001 VDDA.n232 VDDA.n231 16.8187
R1002 VDDA.n372 VDDA.n357 16.363
R1003 VDDA.n468 VDDA.t274 15.0181
R1004 VDDA.n420 VDDA.n419 14.363
R1005 VDDA.n228 VDDA.n221 14.0505
R1006 VDDA.n373 VDDA.n372 13.8005
R1007 VDDA.n382 VDDA.n381 13.8005
R1008 VDDA.n452 VDDA.n451 13.8005
R1009 VDDA.n439 VDDA.n438 13.8005
R1010 VDDA.n429 VDDA.n428 13.8005
R1011 VDDA.n448 VDDA.n447 13.8005
R1012 VDDA.n462 VDDA.n461 13.8005
R1013 VDDA.n37 VDDA.n10 13.6255
R1014 VDDA.n213 VDDA.n189 13.563
R1015 VDDA.n339 VDDA.t291 13.1338
R1016 VDDA.n339 VDDA.t289 13.1338
R1017 VDDA.n358 VDDA.t310 13.1338
R1018 VDDA.n358 VDDA.t271 13.1338
R1019 VDDA.n360 VDDA.t282 13.1338
R1020 VDDA.n360 VDDA.t301 13.1338
R1021 VDDA.n362 VDDA.t266 13.1338
R1022 VDDA.n362 VDDA.t285 13.1338
R1023 VDDA.n364 VDDA.t299 13.1338
R1024 VDDA.n364 VDDA.t307 13.1338
R1025 VDDA.n366 VDDA.t280 13.1338
R1026 VDDA.n366 VDDA.t276 13.1338
R1027 VDDA.n368 VDDA.t305 13.1338
R1028 VDDA.n368 VDDA.t315 13.1338
R1029 VDDA.n370 VDDA.t273 13.1338
R1030 VDDA.n370 VDDA.t294 13.1338
R1031 VDDA.t379 VDDA.n226 12.313
R1032 VDDA.n226 VDDA.t241 12.313
R1033 VDDA.n210 VDDA.t261 11.2576
R1034 VDDA.n210 VDDA.t446 11.2576
R1035 VDDA.n194 VDDA.t204 11.2576
R1036 VDDA.n194 VDDA.t78 11.2576
R1037 VDDA.n193 VDDA.t40 11.2576
R1038 VDDA.n193 VDDA.t229 11.2576
R1039 VDDA.n191 VDDA.t231 11.2576
R1040 VDDA.n191 VDDA.t9 11.2576
R1041 VDDA.n190 VDDA.t235 11.2576
R1042 VDDA.n190 VDDA.t1 11.2576
R1043 VDDA.n98 VDDA.t450 11.2576
R1044 VDDA.n98 VDDA.t173 11.2576
R1045 VDDA.n82 VDDA.t206 11.2576
R1046 VDDA.n82 VDDA.t259 11.2576
R1047 VDDA.n81 VDDA.t208 11.2576
R1048 VDDA.n81 VDDA.t70 11.2576
R1049 VDDA.n79 VDDA.t33 11.2576
R1050 VDDA.n79 VDDA.t111 11.2576
R1051 VDDA.n78 VDDA.t237 11.2576
R1052 VDDA.n78 VDDA.t136 11.2576
R1053 VDDA.n189 VDDA.n188 9.5005
R1054 VDDA.n212 VDDA.n211 9.3005
R1055 VDDA.n100 VDDA.n99 9.3005
R1056 VDDA.n325 VDDA.n271 9.3005
R1057 VDDA.n322 VDDA.n321 9.3005
R1058 VDDA.n320 VDDA.n319 9.3005
R1059 VDDA.n317 VDDA.n307 9.3005
R1060 VDDA.n316 VDDA.n315 9.3005
R1061 VDDA.n312 VDDA.n308 9.3005
R1062 VDDA.n263 VDDA.n262 9.3005
R1063 VDDA.n336 VDDA.n335 9.3005
R1064 VDDA.n329 VDDA.n328 9.3005
R1065 VDDA.n294 VDDA.n293 9.3005
R1066 VDDA.n397 VDDA.n396 9.3005
R1067 VDDA.n241 VDDA.n240 8.938
R1068 VDDA.n258 VDDA.n257 8.03219
R1069 VDDA.n110 VDDA.t83 8.0005
R1070 VDDA.n110 VDDA.t112 8.0005
R1071 VDDA.n108 VDDA.t102 8.0005
R1072 VDDA.n108 VDDA.t192 8.0005
R1073 VDDA.n106 VDDA.t58 8.0005
R1074 VDDA.n106 VDDA.t256 8.0005
R1075 VDDA.n104 VDDA.t130 8.0005
R1076 VDDA.n104 VDDA.t18 8.0005
R1077 VDDA.n102 VDDA.t44 8.0005
R1078 VDDA.n102 VDDA.t169 8.0005
R1079 VDDA.n101 VDDA.t35 8.0005
R1080 VDDA.n101 VDDA.t183 8.0005
R1081 VDDA.n9 VDDA.t232 8.0005
R1082 VDDA.n9 VDDA.t191 8.0005
R1083 VDDA.n7 VDDA.t15 8.0005
R1084 VDDA.n7 VDDA.t188 8.0005
R1085 VDDA.n5 VDDA.t254 8.0005
R1086 VDDA.n5 VDDA.t53 8.0005
R1087 VDDA.n3 VDDA.t118 8.0005
R1088 VDDA.n3 VDDA.t124 8.0005
R1089 VDDA.n1 VDDA.t212 8.0005
R1090 VDDA.n1 VDDA.t190 8.0005
R1091 VDDA.n0 VDDA.t137 8.0005
R1092 VDDA.n0 VDDA.t34 8.0005
R1093 VDDA.n213 VDDA.n212 7.8755
R1094 VDDA.n189 VDDA.n100 7.8755
R1095 VDDA.n463 VDDA.n462 7.44175
R1096 VDDA.n253 VDDA.n252 6.6255
R1097 VDDA.n112 VDDA.t85 6.56717
R1098 VDDA.n112 VDDA.t115 6.56717
R1099 VDDA.n131 VDDA.t17 6.56717
R1100 VDDA.n131 VDDA.t47 6.56717
R1101 VDDA.n133 VDDA.t129 6.56717
R1102 VDDA.n133 VDDA.t42 6.56717
R1103 VDDA.n135 VDDA.t223 6.56717
R1104 VDDA.n135 VDDA.t194 6.56717
R1105 VDDA.n137 VDDA.t171 6.56717
R1106 VDDA.n137 VDDA.t74 6.56717
R1107 VDDA.n38 VDDA.t123 6.56717
R1108 VDDA.n38 VDDA.t211 6.56717
R1109 VDDA.n54 VDDA.t121 6.56717
R1110 VDDA.n54 VDDA.t14 6.56717
R1111 VDDA.n56 VDDA.t20 6.56717
R1112 VDDA.n56 VDDA.t186 6.56717
R1113 VDDA.n58 VDDA.t139 6.56717
R1114 VDDA.n58 VDDA.t117 6.56717
R1115 VDDA.n60 VDDA.t12 6.56717
R1116 VDDA.n60 VDDA.t127 6.56717
R1117 VDDA.n399 VDDA.n398 6.13371
R1118 VDDA.n338 VDDA.n337 6.098
R1119 VDDA.n77 VDDA.n76 5.438
R1120 VDDA.n241 VDDA.n216 5.1255
R1121 VDDA.n214 VDDA.n77 5.0005
R1122 VDDA.n212 VDDA.n196 4.5005
R1123 VDDA.n188 VDDA.n187 4.5005
R1124 VDDA.n100 VDDA.n84 4.5005
R1125 VDDA.n214 VDDA.n213 4.5005
R1126 VDDA.n295 VDDA.n294 4.5005
R1127 VDDA.n328 VDDA.n327 4.5005
R1128 VDDA.n326 VDDA.n325 4.5005
R1129 VDDA.n323 VDDA.n322 4.5005
R1130 VDDA.n319 VDDA.n304 4.5005
R1131 VDDA.n310 VDDA.n307 4.5005
R1132 VDDA.n315 VDDA.n314 4.5005
R1133 VDDA.n313 VDDA.n312 4.5005
R1134 VDDA.n262 VDDA.n259 4.5005
R1135 VDDA.n337 VDDA.n336 4.5005
R1136 VDDA.n398 VDDA.n397 4.5005
R1137 VDDA.n234 VDDA.n233 4.27978
R1138 VDDA.n256 VDDA.n255 4.12334
R1139 VDDA.n469 VDDA 4.08025
R1140 VDDA.n327 VDDA.n303 3.3755
R1141 VDDA.n77 VDDA.n37 3.09425
R1142 VDDA.n187 VDDA.n186 2.938
R1143 VDDA.n257 VDDA.n256 2.93377
R1144 VDDA.n451 VDDA.n448 2.5005
R1145 VDDA.n398 VDDA.n382 2.47371
R1146 VDDA.n253 VDDA.n214 1.938
R1147 VDDA.n438 VDDA.n429 1.813
R1148 VDDA VDDA.n469 1.20605
R1149 VDDA VDDA.n468 1.0815
R1150 VDDA.n372 VDDA.n371 1.0005
R1151 VDDA.n371 VDDA.n369 1.0005
R1152 VDDA.n369 VDDA.n367 1.0005
R1153 VDDA.n367 VDDA.n365 1.0005
R1154 VDDA.n365 VDDA.n363 1.0005
R1155 VDDA.n363 VDDA.n361 1.0005
R1156 VDDA.n361 VDDA.n359 1.0005
R1157 VDDA.n359 VDDA.n340 1.0005
R1158 VDDA.n382 VDDA.n340 1.0005
R1159 VDDA.n187 VDDA.n150 0.938
R1160 VDDA.n338 VDDA.n258 0.840625
R1161 VDDA.n469 VDDA.n254 0.7948
R1162 VDDA.n399 VDDA.n338 0.74075
R1163 VDDA.n240 VDDA.n221 0.6255
R1164 VDDA.n196 VDDA.n195 0.6255
R1165 VDDA.n196 VDDA.n192 0.6255
R1166 VDDA.n84 VDDA.n83 0.6255
R1167 VDDA.n84 VDDA.n80 0.6255
R1168 VDDA.n277 VDDA.n275 0.6255
R1169 VDDA.n279 VDDA.n277 0.6255
R1170 VDDA.n295 VDDA.n279 0.6255
R1171 VDDA.n297 VDDA.n295 0.6255
R1172 VDDA.n299 VDDA.n297 0.6255
R1173 VDDA.n301 VDDA.n299 0.6255
R1174 VDDA.n303 VDDA.n301 0.6255
R1175 VDDA.n327 VDDA.n326 0.6255
R1176 VDDA.n326 VDDA.n323 0.6255
R1177 VDDA.n323 VDDA.n304 0.6255
R1178 VDDA.n310 VDDA.n304 0.6255
R1179 VDDA.n314 VDDA.n310 0.6255
R1180 VDDA.n314 VDDA.n313 0.6255
R1181 VDDA.n313 VDDA.n259 0.6255
R1182 VDDA.n337 VDDA.n259 0.6255
R1183 VDDA.n171 VDDA.n169 0.563
R1184 VDDA.n169 VDDA.n167 0.563
R1185 VDDA.n167 VDDA.n165 0.563
R1186 VDDA.n165 VDDA.n163 0.563
R1187 VDDA.n163 VDDA.n161 0.563
R1188 VDDA.n161 VDDA.n159 0.563
R1189 VDDA.n159 VDDA.n157 0.563
R1190 VDDA.n157 VDDA.n155 0.563
R1191 VDDA.n155 VDDA.n152 0.563
R1192 VDDA.n186 VDDA.n152 0.563
R1193 VDDA.n138 VDDA.n136 0.563
R1194 VDDA.n136 VDDA.n134 0.563
R1195 VDDA.n134 VDDA.n132 0.563
R1196 VDDA.n132 VDDA.n113 0.563
R1197 VDDA.n150 VDDA.n113 0.563
R1198 VDDA.n105 VDDA.n103 0.563
R1199 VDDA.n107 VDDA.n105 0.563
R1200 VDDA.n109 VDDA.n107 0.563
R1201 VDDA.n111 VDDA.n109 0.563
R1202 VDDA.n61 VDDA.n59 0.563
R1203 VDDA.n59 VDDA.n57 0.563
R1204 VDDA.n57 VDDA.n55 0.563
R1205 VDDA.n55 VDDA.n39 0.563
R1206 VDDA.n76 VDDA.n39 0.563
R1207 VDDA.n4 VDDA.n2 0.563
R1208 VDDA.n6 VDDA.n4 0.563
R1209 VDDA.n8 VDDA.n6 0.563
R1210 VDDA.n10 VDDA.n8 0.563
R1211 VDDA.n419 VDDA.n413 0.563
R1212 VDDA.n429 VDDA.n413 0.563
R1213 VDDA.n438 VDDA.n437 0.563
R1214 VDDA.n437 VDDA.n435 0.563
R1215 VDDA.n435 VDDA.n433 0.563
R1216 VDDA.n433 VDDA.n431 0.563
R1217 VDDA.n431 VDDA.n407 0.563
R1218 VDDA.n448 VDDA.n407 0.563
R1219 VDDA.n451 VDDA.n450 0.563
R1220 VDDA.n450 VDDA.n401 0.563
R1221 VDDA.n462 VDDA.n401 0.563
R1222 VDDA.n463 VDDA.n399 0.546875
R1223 VDDA.n468 VDDA.n463 0.370625
R1224 VDDA.n252 VDDA.n216 0.2505
R1225 VDDA.t267 VDDA.t283 0.1603
R1226 VDDA.t311 VDDA.t303 0.1603
R1227 VDDA.t308 VDDA.t268 0.1603
R1228 VDDA.t296 VDDA.t292 0.1603
R1229 VDDA.t269 VDDA.t286 0.1603
R1230 VDDA.t313 VDDA.t297 0.1603
R1231 VDDA.t287 VDDA.t302 0.1603
R1232 VDDA.t278 VDDA.t264 0.1603
R1233 VDDA.n465 VDDA.t295 0.159278
R1234 VDDA.n466 VDDA.t277 0.159278
R1235 VDDA.n467 VDDA.t312 0.159278
R1236 VDDA.n467 VDDA.t267 0.1368
R1237 VDDA.n467 VDDA.t311 0.1368
R1238 VDDA.n466 VDDA.t308 0.1368
R1239 VDDA.n466 VDDA.t296 0.1368
R1240 VDDA.n465 VDDA.t269 0.1368
R1241 VDDA.n465 VDDA.t313 0.1368
R1242 VDDA.n464 VDDA.t287 0.1368
R1243 VDDA.n464 VDDA.t278 0.1368
R1244 VDDA.t295 VDDA.n464 0.00152174
R1245 VDDA.t277 VDDA.n465 0.00152174
R1246 VDDA.t312 VDDA.n466 0.00152174
R1247 VDDA.t274 VDDA.n467 0.00152174
R1248 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 628.034
R1249 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 626.784
R1250 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 622.284
R1251 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t21 289.2
R1252 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.t7 289.2
R1253 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 227.252
R1254 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 212.733
R1255 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 212.733
R1256 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 176.733
R1257 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 176.733
R1258 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 176.733
R1259 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 176.733
R1260 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 176.733
R1261 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 152
R1262 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 152
R1263 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 two_stage_opamp_dummy_magic_0.err_amp_mir.t11 112.468
R1264 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 two_stage_opamp_dummy_magic_0.err_amp_mir.t15 112.468
R1265 two_stage_opamp_dummy_magic_0.err_amp_mir.n5 two_stage_opamp_dummy_magic_0.err_amp_mir.t17 112.468
R1266 two_stage_opamp_dummy_magic_0.err_amp_mir.n4 two_stage_opamp_dummy_magic_0.err_amp_mir.t19 112.468
R1267 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.t13 112.468
R1268 two_stage_opamp_dummy_magic_0.err_amp_mir.n10 two_stage_opamp_dummy_magic_0.err_amp_mir.t18 112.468
R1269 two_stage_opamp_dummy_magic_0.err_amp_mir.n11 two_stage_opamp_dummy_magic_0.err_amp_mir.t20 112.468
R1270 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 two_stage_opamp_dummy_magic_0.err_amp_mir.t9 112.468
R1271 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t5 78.8005
R1272 two_stage_opamp_dummy_magic_0.err_amp_mir.n17 two_stage_opamp_dummy_magic_0.err_amp_mir.t2 78.8005
R1273 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t3 78.8005
R1274 two_stage_opamp_dummy_magic_0.err_amp_mir.n16 two_stage_opamp_dummy_magic_0.err_amp_mir.t4 78.8005
R1275 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t1 78.8005
R1276 two_stage_opamp_dummy_magic_0.err_amp_mir.n15 two_stage_opamp_dummy_magic_0.err_amp_mir.t6 78.8005
R1277 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t16 48.0005
R1278 two_stage_opamp_dummy_magic_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_0.err_amp_mir.t10 48.0005
R1279 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t14 48.0005
R1280 two_stage_opamp_dummy_magic_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_0.err_amp_mir.t12 48.0005
R1281 two_stage_opamp_dummy_magic_0.err_amp_mir.t0 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 48.0005
R1282 two_stage_opamp_dummy_magic_0.err_amp_mir.n20 two_stage_opamp_dummy_magic_0.err_amp_mir.t8 48.0005
R1283 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 two_stage_opamp_dummy_magic_0.err_amp_mir.n7 45.5227
R1284 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n6 45.5227
R1285 two_stage_opamp_dummy_magic_0.err_amp_mir.n13 two_stage_opamp_dummy_magic_0.err_amp_mir.n12 45.5227
R1286 two_stage_opamp_dummy_magic_0.err_amp_mir.n9 two_stage_opamp_dummy_magic_0.err_amp_mir.n8 45.5227
R1287 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n2 15.488
R1288 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n14 14.238
R1289 two_stage_opamp_dummy_magic_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 6.1255
R1290 two_stage_opamp_dummy_magic_0.err_amp_mir.n19 two_stage_opamp_dummy_magic_0.err_amp_mir.n18 5.7505
R1291 GNDA.n404 GNDA.n30 227083
R1292 GNDA.n1688 GNDA.n1687 40282.1
R1293 GNDA.n2471 GNDA.n57 30529.2
R1294 GNDA.n407 GNDA.n403 29344.6
R1295 GNDA.n1619 GNDA.n84 28608.1
R1296 GNDA.n2471 GNDA.n56 28430.8
R1297 GNDA.n405 GNDA.n403 28430.8
R1298 GNDA.n406 GNDA.n404 26656.2
R1299 GNDA.n1686 GNDA.n1619 26648.4
R1300 GNDA.n405 GNDA.n80 23523.1
R1301 GNDA.n80 GNDA.n56 23523.1
R1302 GNDA.n1687 GNDA.n83 21442.2
R1303 GNDA.n2452 GNDA.n2451 21037.5
R1304 GNDA.n1687 GNDA.n84 19885.8
R1305 GNDA.n2454 GNDA.n80 19630.8
R1306 GNDA.n2453 GNDA.n81 19055.4
R1307 GNDA.n405 GNDA.n81 17609.2
R1308 GNDA.n2456 GNDA.n56 17609.2
R1309 GNDA.n1690 GNDA.n1686 17265.8
R1310 GNDA.n2454 GNDA.n2453 15992.3
R1311 GNDA.n1688 GNDA.n1686 15892.5
R1312 GNDA.n1692 GNDA.n1621 12361.8
R1313 GNDA.n1696 GNDA.n1621 12312.5
R1314 GNDA.n404 GNDA.n56 11934.7
R1315 GNDA.n1692 GNDA.n1622 11918.5
R1316 GNDA.n1696 GNDA.n1622 11869.2
R1317 GNDA.n496 GNDA.n81 10910.2
R1318 GNDA.n2455 GNDA.n2454 10879.5
R1319 GNDA.n481 GNDA.n336 10441
R1320 GNDA.n477 GNDA.n336 10441
R1321 GNDA.n481 GNDA.n337 10441
R1322 GNDA.n477 GNDA.n337 10441
R1323 GNDA.n1736 GNDA.n1619 10371.4
R1324 GNDA.n2490 GNDA.n31 9259
R1325 GNDA.n1699 GNDA.n1648 9062
R1326 GNDA.n2490 GNDA.n32 8914.25
R1327 GNDA.n107 GNDA.n103 8175.5
R1328 GNDA.n2436 GNDA.n103 8126.25
R1329 GNDA.n1703 GNDA.n1643 7880
R1330 GNDA.n1703 GNDA.n1644 7880
R1331 GNDA.n1742 GNDA.n1616 7880
R1332 GNDA.n1738 GNDA.n1616 7880
R1333 GNDA.n1646 GNDA.n1643 7830.75
R1334 GNDA.n1646 GNDA.n1644 7830.75
R1335 GNDA.n1742 GNDA.n1617 7830.75
R1336 GNDA.n1738 GNDA.n1617 7830.75
R1337 GNDA.n107 GNDA.n101 7732.25
R1338 GNDA.n2478 GNDA.n40 7732.25
R1339 GNDA.n2478 GNDA.n41 7732.25
R1340 GNDA.n2480 GNDA.n40 7732.25
R1341 GNDA.n2480 GNDA.n41 7732.25
R1342 GNDA.n485 GNDA.n333 7732.25
R1343 GNDA.n485 GNDA.n334 7732.25
R1344 GNDA.n335 GNDA.n333 7732.25
R1345 GNDA.n335 GNDA.n334 7732.25
R1346 GNDA.n2436 GNDA.n101 7683
R1347 GNDA.n2183 GNDA.n314 6845.75
R1348 GNDA.n2187 GNDA.n314 6845.75
R1349 GNDA.n2183 GNDA.n313 6796.5
R1350 GNDA.n2187 GNDA.n313 6796.5
R1351 GNDA.n2181 GNDA.n498 6698
R1352 GNDA.n2176 GNDA.n498 6698
R1353 GNDA.n2181 GNDA.n497 6648.75
R1354 GNDA.n2176 GNDA.n497 6648.75
R1355 GNDA.n395 GNDA.n318 6008.5
R1356 GNDA.n74 GNDA.n71 5860.75
R1357 GNDA.n2458 GNDA.n71 5811.5
R1358 GNDA.n494 GNDA.n318 5762.25
R1359 GNDA.n407 GNDA.n406 5446.53
R1360 GNDA.n395 GNDA.n319 5319
R1361 GNDA.n465 GNDA.n462 5319
R1362 GNDA.n443 GNDA.n442 5319
R1363 GNDA.n75 GNDA.n74 5319
R1364 GNDA.n494 GNDA.n319 5269.75
R1365 GNDA.n2458 GNDA.n75 5269.75
R1366 GNDA.n402 GNDA.n371 5171.25
R1367 GNDA.n408 GNDA.n31 5171.25
R1368 GNDA.n411 GNDA.n32 5171.25
R1369 GNDA.n2470 GNDA.n58 5171.25
R1370 GNDA.n2453 GNDA.n2452 5144.1
R1371 GNDA.n398 GNDA.n371 5122
R1372 GNDA.n2466 GNDA.n58 5122
R1373 GNDA.n1701 GNDA.n1648 4974.25
R1374 GNDA.n1720 GNDA.n1634 4974.25
R1375 GNDA.n1724 GNDA.n1634 4974.25
R1376 GNDA.n402 GNDA.n372 4944.7
R1377 GNDA.n2470 GNDA.n59 4944.7
R1378 GNDA.n459 GNDA.n449 4925
R1379 GNDA.n459 GNDA.n450 4925
R1380 GNDA.n398 GNDA.n372 4895.45
R1381 GNDA.n2466 GNDA.n59 4895.45
R1382 GNDA.n449 GNDA.n360 4728
R1383 GNDA.n450 GNDA.n360 4728
R1384 GNDA.n2440 GNDA.n96 4678.75
R1385 GNDA.n2440 GNDA.n95 4629.5
R1386 GNDA.n167 GNDA.n96 4629.5
R1387 GNDA.n2450 GNDA.n84 4598.65
R1388 GNDA.n2162 GNDA.n512 4580.25
R1389 GNDA.n2162 GNDA.n513 4580.25
R1390 GNDA.n167 GNDA.n95 4580.25
R1391 GNDA.n2158 GNDA.n511 4580.25
R1392 GNDA.n521 GNDA.n511 4580.25
R1393 GNDA.n1735 GNDA.n1623 4531
R1394 GNDA.n1735 GNDA.n1624 4531
R1395 GNDA.n1623 GNDA.n1620 4531
R1396 GNDA.n1624 GNDA.n1620 4531
R1397 GNDA.n1720 GNDA.n1633 4531
R1398 GNDA.n1724 GNDA.n1633 4531
R1399 GNDA.n2129 GNDA.n512 4481.75
R1400 GNDA.n2129 GNDA.n513 4481.75
R1401 GNDA.n2158 GNDA.n518 4481.75
R1402 GNDA.n521 GNDA.n518 4481.75
R1403 GNDA.n496 GNDA.n495 4275.41
R1404 GNDA.n2451 GNDA.n2450 4159.38
R1405 GNDA.n1689 GNDA.n1688 4073.68
R1406 GNDA.n406 GNDA.n405 3964.58
R1407 GNDA.n54 GNDA.n50 3619.88
R1408 GNDA.n368 GNDA.n366 3619.88
R1409 GNDA.n438 GNDA.n408 3595.25
R1410 GNDA.n2493 GNDA.n27 3447.5
R1411 GNDA.n446 GNDA.n27 3398.25
R1412 GNDA.n2493 GNDA.n28 3349
R1413 GNDA.n446 GNDA.n28 3299.75
R1414 GNDA.n1691 GNDA.n1690 3287.9
R1415 GNDA.n438 GNDA.n411 3250.5
R1416 GNDA.n50 GNDA.n48 2437.88
R1417 GNDA.n366 GNDA.n326 2437.88
R1418 GNDA.n386 GNDA.n383 2326.02
R1419 GNDA.n393 GNDA.n383 2326.02
R1420 GNDA.n66 GNDA.n63 2326.02
R1421 GNDA.n77 GNDA.n63 2326.02
R1422 GNDA.n1684 GNDA.n1654 2142.38
R1423 GNDA.n1717 GNDA.n1632 2142.38
R1424 GNDA.n1654 GNDA.n1653 1846.88
R1425 GNDA.n1728 GNDA.n1632 1846.88
R1426 GNDA.n1689 GNDA.n79 1749.05
R1427 GNDA.n1853 GNDA.n608 1672.5
R1428 GNDA.n2473 GNDA.n50 1456.78
R1429 GNDA.n366 GNDA.n325 1456.78
R1430 GNDA.n1690 GNDA.n1689 1226.55
R1431 GNDA.n441 GNDA.n407 1184.62
R1432 GNDA.n2455 GNDA.n79 1163.28
R1433 GNDA.n390 GNDA.n383 1114.8
R1434 GNDA.n2463 GNDA.n63 1114.8
R1435 GNDA.n752 GNDA.n625 1064.42
R1436 GNDA.n1450 GNDA.n598 1064.42
R1437 GNDA.n1432 GNDA.n625 1041.66
R1438 GNDA.n1877 GNDA.n598 1041.66
R1439 GNDA.n1681 GNDA.n1654 991.841
R1440 GNDA.n1712 GNDA.n1632 991.841
R1441 GNDA.n2182 GNDA.n317 991.54
R1442 GNDA.n2457 GNDA.n2456 971.551
R1443 GNDA.n2456 GNDA.n2455 890.324
R1444 GNDA.n83 GNDA.n79 831.111
R1445 GNDA.n1693 GNDA.n1637 803.201
R1446 GNDA.n1695 GNDA.n1637 800
R1447 GNDA.n1694 GNDA.n1693 774.4
R1448 GNDA.n1695 GNDA.n1694 771.201
R1449 GNDA.n327 GNDA.t251 734.418
R1450 GNDA.n323 GNDA.t244 734.418
R1451 GNDA.n51 GNDA.t241 734.418
R1452 GNDA.n46 GNDA.t222 734.418
R1453 GNDA.n467 GNDA.n466 691.201
R1454 GNDA.n365 GNDA.n357 691.201
R1455 GNDA.n2487 GNDA.t263 682.201
R1456 GNDA.n479 GNDA.n478 678.4
R1457 GNDA.n480 GNDA.n479 672
R1458 GNDA.n2081 GNDA.n554 669.307
R1459 GNDA.n434 GNDA.t235 666.134
R1460 GNDA.n2067 GNDA.n2066 662.155
R1461 GNDA.n2340 GNDA.n145 662.155
R1462 GNDA.n392 GNDA.n384 617.601
R1463 GNDA.n68 GNDA.n67 617.601
R1464 GNDA.n2489 GNDA.n33 601.601
R1465 GNDA.n441 GNDA.t305 592.308
R1466 GNDA.t302 GNDA.n57 592.308
R1467 GNDA.n2082 GNDA.n555 585
R1468 GNDA.n2084 GNDA.n2083 585
R1469 GNDA.n2085 GNDA.n2084 585
R1470 GNDA.n567 GNDA.n566 585
R1471 GNDA.n2068 GNDA.n567 585
R1472 GNDA.n2071 GNDA.n2070 585
R1473 GNDA.n2070 GNDA.n2069 585
R1474 GNDA.n2072 GNDA.n565 585
R1475 GNDA.n565 GNDA.n564 585
R1476 GNDA.n2074 GNDA.n2073 585
R1477 GNDA.n2075 GNDA.n2074 585
R1478 GNDA.n563 GNDA.n562 585
R1479 GNDA.n2076 GNDA.n563 585
R1480 GNDA.n2079 GNDA.n2078 585
R1481 GNDA.n2078 GNDA.n2077 585
R1482 GNDA.n553 GNDA.n552 585
R1483 GNDA.n2086 GNDA.n553 585
R1484 GNDA.n2089 GNDA.n2088 585
R1485 GNDA.n2088 GNDA.n2087 585
R1486 GNDA.n2090 GNDA.n551 585
R1487 GNDA.n551 GNDA.n550 585
R1488 GNDA.n2093 GNDA.n2092 585
R1489 GNDA.n2094 GNDA.n2093 585
R1490 GNDA.n2091 GNDA.n547 585
R1491 GNDA.n2095 GNDA.n547 585
R1492 GNDA.n2097 GNDA.n549 585
R1493 GNDA.n2097 GNDA.n2096 585
R1494 GNDA.n904 GNDA.n741 585
R1495 GNDA.n741 GNDA.n740 585
R1496 GNDA.n906 GNDA.n905 585
R1497 GNDA.n907 GNDA.n906 585
R1498 GNDA.n739 GNDA.n738 585
R1499 GNDA.n908 GNDA.n739 585
R1500 GNDA.n912 GNDA.n911 585
R1501 GNDA.n911 GNDA.n910 585
R1502 GNDA.n913 GNDA.n737 585
R1503 GNDA.n909 GNDA.n737 585
R1504 GNDA.n915 GNDA.n914 585
R1505 GNDA.n915 GNDA.n621 585
R1506 GNDA.n916 GNDA.n736 585
R1507 GNDA.n916 GNDA.n622 585
R1508 GNDA.n919 GNDA.n918 585
R1509 GNDA.n918 GNDA.n917 585
R1510 GNDA.n920 GNDA.n735 585
R1511 GNDA.n735 GNDA.n734 585
R1512 GNDA.n923 GNDA.n922 585
R1513 GNDA.n924 GNDA.n923 585
R1514 GNDA.n921 GNDA.n731 585
R1515 GNDA.n925 GNDA.n731 585
R1516 GNDA.n927 GNDA.n733 585
R1517 GNDA.n927 GNDA.n926 585
R1518 GNDA.n928 GNDA.n730 585
R1519 GNDA.n928 GNDA.n568 585
R1520 GNDA.n751 GNDA.n750 585
R1521 GNDA.n884 GNDA.n751 585
R1522 GNDA.n887 GNDA.n886 585
R1523 GNDA.n886 GNDA.n885 585
R1524 GNDA.n888 GNDA.n749 585
R1525 GNDA.n749 GNDA.n748 585
R1526 GNDA.n890 GNDA.n889 585
R1527 GNDA.n891 GNDA.n890 585
R1528 GNDA.n747 GNDA.n746 585
R1529 GNDA.n892 GNDA.n747 585
R1530 GNDA.n895 GNDA.n894 585
R1531 GNDA.n894 GNDA.n893 585
R1532 GNDA.n896 GNDA.n745 585
R1533 GNDA.n745 GNDA.n744 585
R1534 GNDA.n898 GNDA.n897 585
R1535 GNDA.n899 GNDA.n898 585
R1536 GNDA.n743 GNDA.n742 585
R1537 GNDA.n900 GNDA.n743 585
R1538 GNDA.n903 GNDA.n902 585
R1539 GNDA.n902 GNDA.n901 585
R1540 GNDA.n1423 GNDA.n1422 585
R1541 GNDA.n1449 GNDA.n1423 585
R1542 GNDA.n1447 GNDA.n1446 585
R1543 GNDA.n1448 GNDA.n1447 585
R1544 GNDA.n1445 GNDA.n1425 585
R1545 GNDA.n1425 GNDA.n1424 585
R1546 GNDA.n1444 GNDA.n1443 585
R1547 GNDA.n1443 GNDA.n1442 585
R1548 GNDA.n1427 GNDA.n1426 585
R1549 GNDA.n1441 GNDA.n1427 585
R1550 GNDA.n1439 GNDA.n1438 585
R1551 GNDA.n1440 GNDA.n1439 585
R1552 GNDA.n1437 GNDA.n1429 585
R1553 GNDA.n1429 GNDA.n1428 585
R1554 GNDA.n1436 GNDA.n1435 585
R1555 GNDA.n1435 GNDA.n1434 585
R1556 GNDA.n1431 GNDA.n1430 585
R1557 GNDA.n1433 GNDA.n1431 585
R1558 GNDA.n633 GNDA.n632 585
R1559 GNDA.n1432 GNDA.n632 585
R1560 GNDA.n1878 GNDA.n596 585
R1561 GNDA.n1878 GNDA.n1877 585
R1562 GNDA.n601 GNDA.n597 585
R1563 GNDA.n1876 GNDA.n597 585
R1564 GNDA.n1874 GNDA.n1873 585
R1565 GNDA.n1875 GNDA.n1874 585
R1566 GNDA.n1872 GNDA.n600 585
R1567 GNDA.n600 GNDA.n599 585
R1568 GNDA.n1871 GNDA.n1870 585
R1569 GNDA.n1870 GNDA.n1869 585
R1570 GNDA.n603 GNDA.n602 585
R1571 GNDA.n1868 GNDA.n603 585
R1572 GNDA.n1866 GNDA.n1865 585
R1573 GNDA.n1867 GNDA.n1866 585
R1574 GNDA.n1864 GNDA.n605 585
R1575 GNDA.n605 GNDA.n604 585
R1576 GNDA.n1863 GNDA.n1862 585
R1577 GNDA.n1862 GNDA.n1861 585
R1578 GNDA.n607 GNDA.n606 585
R1579 GNDA.n1860 GNDA.n607 585
R1580 GNDA.n1859 GNDA.n1858 585
R1581 GNDA.n609 GNDA.n608 585
R1582 GNDA.n1881 GNDA.n1880 585
R1583 GNDA.n1882 GNDA.n595 585
R1584 GNDA.n1884 GNDA.n1883 585
R1585 GNDA.n1886 GNDA.n594 585
R1586 GNDA.n1889 GNDA.n1888 585
R1587 GNDA.n1890 GNDA.n593 585
R1588 GNDA.n1892 GNDA.n1891 585
R1589 GNDA.n1894 GNDA.n592 585
R1590 GNDA.n1897 GNDA.n1896 585
R1591 GNDA.n1898 GNDA.n591 585
R1592 GNDA.n1900 GNDA.n1899 585
R1593 GNDA.n1902 GNDA.n589 585
R1594 GNDA.n1602 GNDA.n1601 585
R1595 GNDA.n1600 GNDA.n631 585
R1596 GNDA.n1599 GNDA.n1598 585
R1597 GNDA.n1597 GNDA.n1596 585
R1598 GNDA.n1595 GNDA.n1594 585
R1599 GNDA.n1593 GNDA.n1592 585
R1600 GNDA.n1591 GNDA.n1590 585
R1601 GNDA.n1589 GNDA.n1588 585
R1602 GNDA.n1587 GNDA.n1586 585
R1603 GNDA.n1585 GNDA.n1584 585
R1604 GNDA.n1583 GNDA.n1582 585
R1605 GNDA.n1581 GNDA.n1580 585
R1606 GNDA.n959 GNDA.n958 585
R1607 GNDA.n947 GNDA.n720 585
R1608 GNDA.n948 GNDA.n723 585
R1609 GNDA.n951 GNDA.n950 585
R1610 GNDA.n946 GNDA.n725 585
R1611 GNDA.n944 GNDA.n943 585
R1612 GNDA.n727 GNDA.n726 585
R1613 GNDA.n937 GNDA.n936 585
R1614 GNDA.n934 GNDA.n729 585
R1615 GNDA.n932 GNDA.n931 585
R1616 GNDA.n1561 GNDA.n655 585
R1617 GNDA.n1562 GNDA.n653 585
R1618 GNDA.n1563 GNDA.n652 585
R1619 GNDA.n650 GNDA.n648 585
R1620 GNDA.n1569 GNDA.n647 585
R1621 GNDA.n1570 GNDA.n645 585
R1622 GNDA.n1571 GNDA.n644 585
R1623 GNDA.n642 GNDA.n640 585
R1624 GNDA.n1576 GNDA.n639 585
R1625 GNDA.n1577 GNDA.n637 585
R1626 GNDA.n573 GNDA.n570 585
R1627 GNDA.n1933 GNDA.n1932 585
R1628 GNDA.n577 GNDA.n576 585
R1629 GNDA.n1923 GNDA.n579 585
R1630 GNDA.n1925 GNDA.n1924 585
R1631 GNDA.n1920 GNDA.n581 585
R1632 GNDA.n1919 GNDA.n1918 585
R1633 GNDA.n1910 GNDA.n583 585
R1634 GNDA.n1912 GNDA.n1911 585
R1635 GNDA.n1908 GNDA.n585 585
R1636 GNDA.n1907 GNDA.n1906 585
R1637 GNDA.n1907 GNDA.n570 585
R1638 GNDA.n931 GNDA.n930 585
R1639 GNDA.n729 GNDA.n728 585
R1640 GNDA.n938 GNDA.n937 585
R1641 GNDA.n940 GNDA.n727 585
R1642 GNDA.n943 GNDA.n942 585
R1643 GNDA.n725 GNDA.n724 585
R1644 GNDA.n952 GNDA.n951 585
R1645 GNDA.n954 GNDA.n723 585
R1646 GNDA.n955 GNDA.n720 585
R1647 GNDA.n958 GNDA.n957 585
R1648 GNDA.n1579 GNDA.n635 585
R1649 GNDA.n1579 GNDA.n588 585
R1650 GNDA.n1578 GNDA.n1577 585
R1651 GNDA.n1576 GNDA.n1575 585
R1652 GNDA.n1574 GNDA.n640 585
R1653 GNDA.n1572 GNDA.n1571 585
R1654 GNDA.n1570 GNDA.n641 585
R1655 GNDA.n1569 GNDA.n1568 585
R1656 GNDA.n1566 GNDA.n648 585
R1657 GNDA.n1564 GNDA.n1563 585
R1658 GNDA.n1562 GNDA.n649 585
R1659 GNDA.n1561 GNDA.n1560 585
R1660 GNDA.n1903 GNDA.n587 585
R1661 GNDA.n1903 GNDA.n588 585
R1662 GNDA.n1906 GNDA.n1905 585
R1663 GNDA.n585 GNDA.n584 585
R1664 GNDA.n1913 GNDA.n1912 585
R1665 GNDA.n1915 GNDA.n583 585
R1666 GNDA.n1918 GNDA.n1917 585
R1667 GNDA.n581 GNDA.n580 585
R1668 GNDA.n1926 GNDA.n1925 585
R1669 GNDA.n1928 GNDA.n579 585
R1670 GNDA.n1929 GNDA.n577 585
R1671 GNDA.n1932 GNDA.n1931 585
R1672 GNDA.n578 GNDA.n569 585
R1673 GNDA.n1820 GNDA.n569 585
R1674 GNDA.n1221 GNDA.n586 585
R1675 GNDA.n1272 GNDA.n1271 585
R1676 GNDA.n1270 GNDA.n1220 585
R1677 GNDA.n1269 GNDA.n1268 585
R1678 GNDA.n1267 GNDA.n1266 585
R1679 GNDA.n1265 GNDA.n1264 585
R1680 GNDA.n1263 GNDA.n1262 585
R1681 GNDA.n1261 GNDA.n1260 585
R1682 GNDA.n1259 GNDA.n1258 585
R1683 GNDA.n1257 GNDA.n1256 585
R1684 GNDA.n1255 GNDA.n1254 585
R1685 GNDA.n1253 GNDA.n1252 585
R1686 GNDA.n689 GNDA.n688 585
R1687 GNDA.n687 GNDA.n666 585
R1688 GNDA.n686 GNDA.n685 585
R1689 GNDA.n684 GNDA.n683 585
R1690 GNDA.n682 GNDA.n681 585
R1691 GNDA.n680 GNDA.n679 585
R1692 GNDA.n678 GNDA.n677 585
R1693 GNDA.n676 GNDA.n675 585
R1694 GNDA.n674 GNDA.n673 585
R1695 GNDA.n672 GNDA.n671 585
R1696 GNDA.n670 GNDA.n669 585
R1697 GNDA.n668 GNDA.n667 585
R1698 GNDA.n2333 GNDA.n146 585
R1699 GNDA.n1232 GNDA.n148 585
R1700 GNDA.n1233 GNDA.n1230 585
R1701 GNDA.n1236 GNDA.n1229 585
R1702 GNDA.n1237 GNDA.n1228 585
R1703 GNDA.n1240 GNDA.n1227 585
R1704 GNDA.n1241 GNDA.n1226 585
R1705 GNDA.n1244 GNDA.n1225 585
R1706 GNDA.n1245 GNDA.n1224 585
R1707 GNDA.n1248 GNDA.n1223 585
R1708 GNDA.n1249 GNDA.n161 585
R1709 GNDA.n2333 GNDA.n161 585
R1710 GNDA.n1251 GNDA.n1222 585
R1711 GNDA.n1251 GNDA.n187 585
R1712 GNDA.n1250 GNDA.n1249 585
R1713 GNDA.n1248 GNDA.n1247 585
R1714 GNDA.n1246 GNDA.n1245 585
R1715 GNDA.n1244 GNDA.n1243 585
R1716 GNDA.n1242 GNDA.n1241 585
R1717 GNDA.n1240 GNDA.n1239 585
R1718 GNDA.n1238 GNDA.n1237 585
R1719 GNDA.n1236 GNDA.n1235 585
R1720 GNDA.n1234 GNDA.n1233 585
R1721 GNDA.n1232 GNDA.n1231 585
R1722 GNDA.n2302 GNDA.n199 585
R1723 GNDA.n2302 GNDA.n205 585
R1724 GNDA.n1205 GNDA.n1081 585
R1725 GNDA.n1079 GNDA.n1076 585
R1726 GNDA.n1075 GNDA.n1074 585
R1727 GNDA.n1073 GNDA.n1070 585
R1728 GNDA.n1069 GNDA.n1068 585
R1729 GNDA.n1067 GNDA.n1064 585
R1730 GNDA.n1063 GNDA.n1062 585
R1731 GNDA.n1061 GNDA.n1058 585
R1732 GNDA.n1057 GNDA.n545 585
R1733 GNDA.n2101 GNDA.n2100 585
R1734 GNDA.n2098 GNDA.n544 585
R1735 GNDA.n2098 GNDA.n546 585
R1736 GNDA.n2100 GNDA.n2099 585
R1737 GNDA.n1059 GNDA.n545 585
R1738 GNDA.n1061 GNDA.n1060 585
R1739 GNDA.n1065 GNDA.n1062 585
R1740 GNDA.n1067 GNDA.n1066 585
R1741 GNDA.n1071 GNDA.n1068 585
R1742 GNDA.n1073 GNDA.n1072 585
R1743 GNDA.n1077 GNDA.n1074 585
R1744 GNDA.n1079 GNDA.n1078 585
R1745 GNDA.n1081 GNDA.n1080 585
R1746 GNDA.n2102 GNDA.n543 585
R1747 GNDA.n2103 GNDA.n2102 585
R1748 GNDA.n2106 GNDA.n2105 585
R1749 GNDA.n2105 GNDA.n2104 585
R1750 GNDA.n2107 GNDA.n542 585
R1751 GNDA.n542 GNDA.n541 585
R1752 GNDA.n2109 GNDA.n2108 585
R1753 GNDA.n2110 GNDA.n2109 585
R1754 GNDA.n540 GNDA.n539 585
R1755 GNDA.n2111 GNDA.n540 585
R1756 GNDA.n2114 GNDA.n2113 585
R1757 GNDA.n2113 GNDA.n2112 585
R1758 GNDA.n2115 GNDA.n538 585
R1759 GNDA.n538 GNDA.n537 585
R1760 GNDA.n2117 GNDA.n2116 585
R1761 GNDA.n2118 GNDA.n2117 585
R1762 GNDA.n536 GNDA.n535 585
R1763 GNDA.n2119 GNDA.n536 585
R1764 GNDA.n2123 GNDA.n2122 585
R1765 GNDA.n2122 GNDA.n2121 585
R1766 GNDA.n2124 GNDA.n534 585
R1767 GNDA.n2120 GNDA.n534 585
R1768 GNDA.n2126 GNDA.n2125 585
R1769 GNDA.n2126 GNDA.n317 585
R1770 GNDA.n1207 GNDA.n1082 585
R1771 GNDA.n1207 GNDA.n1206 585
R1772 GNDA.n1108 GNDA.n1107 585
R1773 GNDA.n1103 GNDA.n1102 585
R1774 GNDA.n1179 GNDA.n1178 585
R1775 GNDA.n1182 GNDA.n1181 585
R1776 GNDA.n1101 GNDA.n1098 585
R1777 GNDA.n1094 GNDA.n1093 585
R1778 GNDA.n1190 GNDA.n1189 585
R1779 GNDA.n1193 GNDA.n1192 585
R1780 GNDA.n1092 GNDA.n1089 585
R1781 GNDA.n1085 GNDA.n1084 585
R1782 GNDA.n1201 GNDA.n1200 585
R1783 GNDA.n1204 GNDA.n1203 585
R1784 GNDA.n962 GNDA.n570 585
R1785 GNDA.n960 GNDA.n570 585
R1786 GNDA.n1212 GNDA.n1211 585
R1787 GNDA.n1054 GNDA.n697 585
R1788 GNDA.n701 GNDA.n700 585
R1789 GNDA.n978 GNDA.n977 585
R1790 GNDA.n980 GNDA.n979 585
R1791 GNDA.n984 GNDA.n983 585
R1792 GNDA.n982 GNDA.n968 585
R1793 GNDA.n991 GNDA.n990 585
R1794 GNDA.n993 GNDA.n992 585
R1795 GNDA.n997 GNDA.n996 585
R1796 GNDA.n995 GNDA.n966 585
R1797 GNDA.n964 GNDA.n963 585
R1798 GNDA.n1210 GNDA.n698 585
R1799 GNDA.n698 GNDA.n187 585
R1800 GNDA.n2302 GNDA.n193 585
R1801 GNDA.n2302 GNDA.n206 585
R1802 GNDA.n880 GNDA.n752 585
R1803 GNDA.n883 GNDA.n882 585
R1804 GNDA.n784 GNDA.n783 585
R1805 GNDA.n775 GNDA.n774 585
R1806 GNDA.n855 GNDA.n854 585
R1807 GNDA.n858 GNDA.n857 585
R1808 GNDA.n773 GNDA.n770 585
R1809 GNDA.n766 GNDA.n765 585
R1810 GNDA.n866 GNDA.n865 585
R1811 GNDA.n869 GNDA.n868 585
R1812 GNDA.n764 GNDA.n761 585
R1813 GNDA.n757 GNDA.n755 585
R1814 GNDA.n877 GNDA.n876 585
R1815 GNDA.n879 GNDA.n754 585
R1816 GNDA.n782 GNDA.n777 585
R1817 GNDA.n782 GNDA.n588 585
R1818 GNDA.n722 GNDA.n569 585
R1819 GNDA.n781 GNDA.n569 585
R1820 GNDA.n2295 GNDA.n281 585
R1821 GNDA.n279 GNDA.n276 585
R1822 GNDA.n275 GNDA.n274 585
R1823 GNDA.n273 GNDA.n270 585
R1824 GNDA.n269 GNDA.n268 585
R1825 GNDA.n267 GNDA.n264 585
R1826 GNDA.n263 GNDA.n262 585
R1827 GNDA.n261 GNDA.n259 585
R1828 GNDA.n258 GNDA.n184 585
R1829 GNDA.n2306 GNDA.n2305 585
R1830 GNDA.n185 GNDA.n183 585
R1831 GNDA.n187 GNDA.n185 585
R1832 GNDA.n2305 GNDA.n2304 585
R1833 GNDA.n186 GNDA.n184 585
R1834 GNDA.n261 GNDA.n260 585
R1835 GNDA.n265 GNDA.n262 585
R1836 GNDA.n267 GNDA.n266 585
R1837 GNDA.n271 GNDA.n268 585
R1838 GNDA.n273 GNDA.n272 585
R1839 GNDA.n277 GNDA.n274 585
R1840 GNDA.n279 GNDA.n278 585
R1841 GNDA.n281 GNDA.n280 585
R1842 GNDA.n2309 GNDA.n2308 585
R1843 GNDA.n2310 GNDA.n181 585
R1844 GNDA.n2312 GNDA.n2311 585
R1845 GNDA.n2314 GNDA.n180 585
R1846 GNDA.n2317 GNDA.n2316 585
R1847 GNDA.n2318 GNDA.n179 585
R1848 GNDA.n2320 GNDA.n2319 585
R1849 GNDA.n2322 GNDA.n178 585
R1850 GNDA.n2325 GNDA.n2324 585
R1851 GNDA.n2326 GNDA.n177 585
R1852 GNDA.n2328 GNDA.n2327 585
R1853 GNDA.n2330 GNDA.n176 585
R1854 GNDA.n2297 GNDA.n282 585
R1855 GNDA.n2297 GNDA.n2296 585
R1856 GNDA.n660 GNDA.n570 585
R1857 GNDA.n657 GNDA.n570 585
R1858 GNDA.n1299 GNDA.n1298 585
R1859 GNDA.n1295 GNDA.n1294 585
R1860 GNDA.n1370 GNDA.n1369 585
R1861 GNDA.n1373 GNDA.n1372 585
R1862 GNDA.n1293 GNDA.n1290 585
R1863 GNDA.n1286 GNDA.n1285 585
R1864 GNDA.n1381 GNDA.n1380 585
R1865 GNDA.n1384 GNDA.n1383 585
R1866 GNDA.n1284 GNDA.n1281 585
R1867 GNDA.n1277 GNDA.n1276 585
R1868 GNDA.n1392 GNDA.n1391 585
R1869 GNDA.n1395 GNDA.n1394 585
R1870 GNDA.n208 GNDA.n207 585
R1871 GNDA.n207 GNDA.n187 585
R1872 GNDA.n2302 GNDA.n188 585
R1873 GNDA.n2302 GNDA.n2301 585
R1874 GNDA.n1450 GNDA.n1421 585
R1875 GNDA.n1452 GNDA.n1451 585
R1876 GNDA.n1553 GNDA.n1399 585
R1877 GNDA.n1551 GNDA.n1550 585
R1878 GNDA.n1472 GNDA.n1400 585
R1879 GNDA.n1470 GNDA.n1469 585
R1880 GNDA.n1479 GNDA.n1478 585
R1881 GNDA.n1482 GNDA.n1481 585
R1882 GNDA.n1467 GNDA.n1464 585
R1883 GNDA.n1460 GNDA.n1459 585
R1884 GNDA.n1490 GNDA.n1489 585
R1885 GNDA.n1493 GNDA.n1492 585
R1886 GNDA.n1458 GNDA.n1419 585
R1887 GNDA.n1456 GNDA.n1455 585
R1888 GNDA.n1555 GNDA.n1554 585
R1889 GNDA.n1554 GNDA.n588 585
R1890 GNDA.n1558 GNDA.n569 585
R1891 GNDA.n1398 GNDA.n569 585
R1892 GNDA.n2198 GNDA.n2197 585
R1893 GNDA.n303 GNDA.n302 585
R1894 GNDA.n2269 GNDA.n2268 585
R1895 GNDA.n2272 GNDA.n2271 585
R1896 GNDA.n301 GNDA.n298 585
R1897 GNDA.n294 GNDA.n293 585
R1898 GNDA.n2280 GNDA.n2279 585
R1899 GNDA.n2283 GNDA.n2282 585
R1900 GNDA.n292 GNDA.n289 585
R1901 GNDA.n285 GNDA.n284 585
R1902 GNDA.n2291 GNDA.n2290 585
R1903 GNDA.n2294 GNDA.n2293 585
R1904 GNDA.n256 GNDA.n255 585
R1905 GNDA.n253 GNDA.n209 585
R1906 GNDA.n252 GNDA.n251 585
R1907 GNDA.n250 GNDA.n249 585
R1908 GNDA.n248 GNDA.n211 585
R1909 GNDA.n246 GNDA.n245 585
R1910 GNDA.n244 GNDA.n212 585
R1911 GNDA.n243 GNDA.n242 585
R1912 GNDA.n240 GNDA.n213 585
R1913 GNDA.n238 GNDA.n237 585
R1914 GNDA.n236 GNDA.n214 585
R1915 GNDA.n235 GNDA.n234 585
R1916 GNDA.n489 GNDA.n325 585
R1917 GNDA.n370 GNDA.n325 585
R1918 GNDA.n2474 GNDA.n2473 585
R1919 GNDA.n2473 GNDA.n2472 585
R1920 GNDA.n1105 GNDA.n525 585
R1921 GNDA.n1105 GNDA.n172 585
R1922 GNDA.n2127 GNDA.n533 585
R1923 GNDA.n2128 GNDA.n2127 585
R1924 GNDA.n2133 GNDA.n2132 585
R1925 GNDA.n2132 GNDA.n2131 585
R1926 GNDA.n2134 GNDA.n532 585
R1927 GNDA.n532 GNDA.n531 585
R1928 GNDA.n2136 GNDA.n2135 585
R1929 GNDA.n2137 GNDA.n2136 585
R1930 GNDA.n530 GNDA.n529 585
R1931 GNDA.n2138 GNDA.n530 585
R1932 GNDA.n2142 GNDA.n2141 585
R1933 GNDA.n2141 GNDA.n2140 585
R1934 GNDA.n2143 GNDA.n528 585
R1935 GNDA.n2139 GNDA.n528 585
R1936 GNDA.n2145 GNDA.n2144 585
R1937 GNDA.n2146 GNDA.n2145 585
R1938 GNDA.n527 GNDA.n526 585
R1939 GNDA.n2147 GNDA.n527 585
R1940 GNDA.n2150 GNDA.n2149 585
R1941 GNDA.n2149 GNDA.n2148 585
R1942 GNDA.n2151 GNDA.n523 585
R1943 GNDA.n523 GNDA.n519 585
R1944 GNDA.n2155 GNDA.n2154 585
R1945 GNDA.n524 GNDA.n522 585
R1946 GNDA.n2196 GNDA.n305 585
R1947 GNDA.n2196 GNDA.n169 585
R1948 GNDA.n2331 GNDA.n174 585
R1949 GNDA.n2332 GNDA.n2331 585
R1950 GNDA.n506 GNDA.n175 585
R1951 GNDA.n175 GNDA.n173 585
R1952 GNDA.n507 GNDA.n505 585
R1953 GNDA.n505 GNDA.n504 585
R1954 GNDA.n509 GNDA.n508 585
R1955 GNDA.n510 GNDA.n509 585
R1956 GNDA.n503 GNDA.n502 585
R1957 GNDA.n2164 GNDA.n503 585
R1958 GNDA.n2168 GNDA.n2167 585
R1959 GNDA.n2167 GNDA.n2166 585
R1960 GNDA.n2169 GNDA.n500 585
R1961 GNDA.n2165 GNDA.n500 585
R1962 GNDA.n2173 GNDA.n2172 585
R1963 GNDA.n2174 GNDA.n2173 585
R1964 GNDA.n2171 GNDA.n501 585
R1965 GNDA.n501 GNDA.n312 585
R1966 GNDA.n2170 GNDA.n309 585
R1967 GNDA.n2189 GNDA.n309 585
R1968 GNDA.n2191 GNDA.n311 585
R1969 GNDA.n2191 GNDA.n2190 585
R1970 GNDA.n2193 GNDA.n2192 585
R1971 GNDA.n2195 GNDA.n2194 585
R1972 GNDA.n2444 GNDA.n2443 585
R1973 GNDA.n2443 GNDA.n2442 585
R1974 GNDA.n232 GNDA.n215 585
R1975 GNDA.n232 GNDA.n216 585
R1976 GNDA.n231 GNDA.n218 585
R1977 GNDA.n231 GNDA.n230 585
R1978 GNDA.n221 GNDA.n217 585
R1979 GNDA.n229 GNDA.n217 585
R1980 GNDA.n227 GNDA.n226 585
R1981 GNDA.n228 GNDA.n227 585
R1982 GNDA.n225 GNDA.n220 585
R1983 GNDA.n220 GNDA.n219 585
R1984 GNDA.n224 GNDA.n223 585
R1985 GNDA.n223 GNDA.n222 585
R1986 GNDA.n115 GNDA.n114 585
R1987 GNDA.n117 GNDA.n115 585
R1988 GNDA.n2429 GNDA.n2428 585
R1989 GNDA.n2428 GNDA.n2427 585
R1990 GNDA.n2430 GNDA.n109 585
R1991 GNDA.n109 GNDA.n104 585
R1992 GNDA.n2433 GNDA.n2432 585
R1993 GNDA.n2434 GNDA.n2433 585
R1994 GNDA.n2431 GNDA.n113 585
R1995 GNDA.n113 GNDA.n108 585
R1996 GNDA.n112 GNDA.n111 585
R1997 GNDA.n93 GNDA.n92 585
R1998 GNDA.n2445 GNDA.n88 585
R1999 GNDA.n88 GNDA.n86 585
R2000 GNDA.n2448 GNDA.n2447 585
R2001 GNDA.n2449 GNDA.n2448 585
R2002 GNDA.n2414 GNDA.n87 585
R2003 GNDA.n87 GNDA.n85 585
R2004 GNDA.n2418 GNDA.n2417 585
R2005 GNDA.n2417 GNDA.n2416 585
R2006 GNDA.n124 GNDA.n122 585
R2007 GNDA.n122 GNDA.n120 585
R2008 GNDA.n2425 GNDA.n2424 585
R2009 GNDA.n2426 GNDA.n2425 585
R2010 GNDA.n2344 GNDA.n121 585
R2011 GNDA.n121 GNDA.n119 585
R2012 GNDA.n2351 GNDA.n2350 585
R2013 GNDA.n2352 GNDA.n2351 585
R2014 GNDA.n2342 GNDA.n144 585
R2015 GNDA.n2353 GNDA.n144 585
R2016 GNDA.n2356 GNDA.n2355 585
R2017 GNDA.n2355 GNDA.n2354 585
R2018 GNDA.n143 GNDA.n141 585
R2019 GNDA.n2341 GNDA.n143 585
R2020 GNDA.n2339 GNDA.n2338 585
R2021 GNDA.n2340 GNDA.n2339 585
R2022 GNDA.n2032 GNDA.n1957 585
R2023 GNDA.n1957 GNDA.n1956 585
R2024 GNDA.n2035 GNDA.n2034 585
R2025 GNDA.n2036 GNDA.n2035 585
R2026 GNDA.n1958 GNDA.n1953 585
R2027 GNDA.n2037 GNDA.n1953 585
R2028 GNDA.n2040 GNDA.n2039 585
R2029 GNDA.n2039 GNDA.n2038 585
R2030 GNDA.n1952 GNDA.n1950 585
R2031 GNDA.n1955 GNDA.n1952 585
R2032 GNDA.n1946 GNDA.n1945 585
R2033 GNDA.n1954 GNDA.n1945 585
R2034 GNDA.n2048 GNDA.n2047 585
R2035 GNDA.n2052 GNDA.n2048 585
R2036 GNDA.n2055 GNDA.n2054 585
R2037 GNDA.n2054 GNDA.n2053 585
R2038 GNDA.n1944 GNDA.n1942 585
R2039 GNDA.n2051 GNDA.n1944 585
R2040 GNDA.n2049 GNDA.n1938 585
R2041 GNDA.n2050 GNDA.n2049 585
R2042 GNDA.n2062 GNDA.n574 585
R2043 GNDA.n574 GNDA.n572 585
R2044 GNDA.n2065 GNDA.n2064 585
R2045 GNDA.n2066 GNDA.n2065 585
R2046 GNDA.n2031 GNDA.n2030 585
R2047 GNDA.n2030 GNDA.n2029 585
R2048 GNDA.n1823 GNDA.n1746 585
R2049 GNDA.n1746 GNDA.n1745 585
R2050 GNDA.n1826 GNDA.n1825 585
R2051 GNDA.n1827 GNDA.n1826 585
R2052 GNDA.n1747 GNDA.n1614 585
R2053 GNDA.n1828 GNDA.n1614 585
R2054 GNDA.n1831 GNDA.n1830 585
R2055 GNDA.n1830 GNDA.n1829 585
R2056 GNDA.n1609 GNDA.n1606 585
R2057 GNDA.n1606 GNDA.n1605 585
R2058 GNDA.n1838 GNDA.n1837 585
R2059 GNDA.n1839 GNDA.n1838 585
R2060 GNDA.n1607 GNDA.n620 585
R2061 GNDA.n1840 GNDA.n620 585
R2062 GNDA.n1843 GNDA.n1842 585
R2063 GNDA.n1842 GNDA.n1841 585
R2064 GNDA.n616 GNDA.n613 585
R2065 GNDA.n613 GNDA.n612 585
R2066 GNDA.n1850 GNDA.n1849 585
R2067 GNDA.n1851 GNDA.n1850 585
R2068 GNDA.n614 GNDA.n611 585
R2069 GNDA.n1852 GNDA.n611 585
R2070 GNDA.n1855 GNDA.n1854 585
R2071 GNDA.n1854 GNDA.n1853 585
R2072 GNDA.n1822 GNDA.n1821 585
R2073 GNDA.n1821 GNDA.n571 585
R2074 GNDA.n488 GNDA.n328 569.601
R2075 GNDA.n2475 GNDA.n47 569.601
R2076 GNDA.n1744 GNDA.n1743 556.322
R2077 GNDA.n331 GNDA.t310 535.191
R2078 GNDA.n329 GNDA.t225 535.191
R2079 GNDA.n44 GNDA.t257 535.191
R2080 GNDA.n42 GNDA.t267 535.191
R2081 GNDA.n901 GNDA.n740 534.218
R2082 GNDA.n106 GNDA.n100 531.201
R2083 GNDA.n2437 GNDA.n100 528
R2084 GNDA.n901 GNDA.n900 512.29
R2085 GNDA.n900 GNDA.n899 512.29
R2086 GNDA.n899 GNDA.n744 512.29
R2087 GNDA.n893 GNDA.n744 512.29
R2088 GNDA.n893 GNDA.n892 512.29
R2089 GNDA.n891 GNDA.n748 512.29
R2090 GNDA.n885 GNDA.n748 512.29
R2091 GNDA.n885 GNDA.n884 512.29
R2092 GNDA.n884 GNDA.n883 512.29
R2093 GNDA.n883 GNDA.n752 512.29
R2094 GNDA.n1433 GNDA.n1432 512.29
R2095 GNDA.n1434 GNDA.n1433 512.29
R2096 GNDA.n1434 GNDA.n1428 512.29
R2097 GNDA.n1440 GNDA.n1428 512.29
R2098 GNDA.n1441 GNDA.n1440 512.29
R2099 GNDA.n1442 GNDA.n1424 512.29
R2100 GNDA.n1448 GNDA.n1424 512.29
R2101 GNDA.n1449 GNDA.n1448 512.29
R2102 GNDA.n1451 GNDA.n1449 512.29
R2103 GNDA.n1451 GNDA.n1450 512.29
R2104 GNDA.n1877 GNDA.n1876 512.29
R2105 GNDA.n1876 GNDA.n1875 512.29
R2106 GNDA.n1875 GNDA.n599 512.29
R2107 GNDA.n1869 GNDA.n599 512.29
R2108 GNDA.n1869 GNDA.n1868 512.29
R2109 GNDA.n1867 GNDA.n604 512.29
R2110 GNDA.n1861 GNDA.n604 512.29
R2111 GNDA.n1861 GNDA.n1860 512.29
R2112 GNDA.n1860 GNDA.n1859 512.29
R2113 GNDA.n1859 GNDA.n608 512.29
R2114 GNDA.n1704 GNDA.n1641 512
R2115 GNDA.n1704 GNDA.n1642 512
R2116 GNDA.n1739 GNDA.n1618 512
R2117 GNDA.n1741 GNDA.n1618 512
R2118 GNDA.n1645 GNDA.n1641 508.8
R2119 GNDA.n1645 GNDA.n1642 508.8
R2120 GNDA.n1740 GNDA.n1739 508.8
R2121 GNDA.n1741 GNDA.n1740 508.8
R2122 GNDA.n106 GNDA.n105 499.2
R2123 GNDA.t248 GNDA.n118 496.098
R2124 GNDA.n378 GNDA.n373 496
R2125 GNDA.n2481 GNDA.n38 496
R2126 GNDA.n343 GNDA.t249 493.418
R2127 GNDA.n344 GNDA.t232 493.418
R2128 GNDA.n338 GNDA.t298 493.418
R2129 GNDA.n340 GNDA.t314 493.418
R2130 GNDA.n341 GNDA.t295 493.418
R2131 GNDA.n342 GNDA.t287 493.418
R2132 GNDA.n463 GNDA.t301 493.418
R2133 GNDA.n358 GNDA.t289 493.418
R2134 GNDA.n362 GNDA.t238 493.418
R2135 GNDA.n361 GNDA.t304 493.418
R2136 GNDA.n379 GNDA.n378 489.601
R2137 GNDA.n2481 GNDA.n39 489.601
R2138 GNDA.n2452 GNDA.n82 488.889
R2139 GNDA.n2437 GNDA.n99 486.401
R2140 GNDA.n483 GNDA.n482 463.603
R2141 GNDA.n476 GNDA.n475 463.603
R2142 GNDA.n2185 GNDA.n2184 444.8
R2143 GNDA.n2186 GNDA.n2185 444.8
R2144 GNDA.n2186 GNDA.n315 441.601
R2145 GNDA.n2184 GNDA.n316 438.401
R2146 GNDA.n2180 GNDA.n2179 435.2
R2147 GNDA.n2067 GNDA.n571 434.906
R2148 GNDA.n2029 GNDA.n145 434.906
R2149 GNDA.n2488 GNDA.n34 428.8
R2150 GNDA.n2180 GNDA.n499 425.601
R2151 GNDA.n2178 GNDA.n2177 422.401
R2152 GNDA.n473 GNDA.n472 422.401
R2153 GNDA.n345 GNDA.n339 422.401
R2154 GNDA.n464 GNDA.n359 422.401
R2155 GNDA.n364 GNDA.n363 422.401
R2156 GNDA.n2177 GNDA.n499 419.2
R2157 GNDA.n1655 GNDA.t284 413.084
R2158 GNDA.n1656 GNDA.t280 413.084
R2159 GNDA.n1627 GNDA.t276 413.084
R2160 GNDA.n1625 GNDA.t254 413.084
R2161 GNDA.n1629 GNDA.t292 413.084
R2162 GNDA.n1714 GNDA.t307 413.084
R2163 GNDA.n322 GNDA.n321 390.401
R2164 GNDA.n1700 GNDA.n1699 383.118
R2165 GNDA.n73 GNDA.n69 380.8
R2166 GNDA.t333 GNDA.t155 372.308
R2167 GNDA.t130 GNDA.t125 372.308
R2168 GNDA.t62 GNDA.t130 372.308
R2169 GNDA.t62 GNDA.t26 372.308
R2170 GNDA.t26 GNDA.t115 372.308
R2171 GNDA.t203 GNDA.t209 372.308
R2172 GNDA.t199 GNDA.t211 372.308
R2173 GNDA.t340 GNDA.t141 372.308
R2174 GNDA.t141 GNDA.t139 372.308
R2175 GNDA.t111 GNDA.t79 372.308
R2176 GNDA.t79 GNDA.t126 372.308
R2177 GNDA.t126 GNDA.t153 372.308
R2178 GNDA.n598 GNDA.n590 370.214
R2179 GNDA.n1604 GNDA.n625 370.214
R2180 GNDA.n623 GNDA.n598 365.957
R2181 GNDA.n625 GNDA.n624 365.957
R2182 GNDA.n493 GNDA.n320 361.601
R2183 GNDA.n448 GNDA.t140 355.385
R2184 GNDA.t213 GNDA.n444 355.385
R2185 GNDA.n461 GNDA.t201 355.385
R2186 GNDA.t332 GNDA.n29 355.385
R2187 GNDA.t139 GNDA.n30 355.385
R2188 GNDA.n1719 GNDA.n1615 354.024
R2189 GNDA.n1853 GNDA.n1852 352.627
R2190 GNDA.n1852 GNDA.n1851 352.627
R2191 GNDA.n1851 GNDA.n612 352.627
R2192 GNDA.n1841 GNDA.n612 352.627
R2193 GNDA.n1841 GNDA.n1840 352.627
R2194 GNDA.n1839 GNDA.n1605 352.627
R2195 GNDA.n1829 GNDA.n1605 352.627
R2196 GNDA.n1829 GNDA.n1828 352.627
R2197 GNDA.n1828 GNDA.n1827 352.627
R2198 GNDA.n1745 GNDA.n571 352.627
R2199 GNDA.n2066 GNDA.n572 352.627
R2200 GNDA.n2050 GNDA.n572 352.627
R2201 GNDA.n2051 GNDA.n2050 352.627
R2202 GNDA.n2053 GNDA.n2051 352.627
R2203 GNDA.n2053 GNDA.n2052 352.627
R2204 GNDA.n1955 GNDA.n1954 352.627
R2205 GNDA.n2038 GNDA.n1955 352.627
R2206 GNDA.n2038 GNDA.n2037 352.627
R2207 GNDA.n2037 GNDA.n2036 352.627
R2208 GNDA.n2036 GNDA.n1956 352.627
R2209 GNDA.n2029 GNDA.n1956 352.627
R2210 GNDA.n2341 GNDA.n2340 352.627
R2211 GNDA.n2354 GNDA.n2341 352.627
R2212 GNDA.n2354 GNDA.n2353 352.627
R2213 GNDA.n2353 GNDA.n2352 352.627
R2214 GNDA.n2352 GNDA.n119 352.627
R2215 GNDA.n2426 GNDA.n120 352.627
R2216 GNDA.n2460 GNDA.n2459 352
R2217 GNDA.n2416 GNDA.n85 343.452
R2218 GNDA.n2449 GNDA.n86 343.452
R2219 GNDA.n493 GNDA.n492 342.401
R2220 GNDA.n2459 GNDA.n70 342.401
R2221 GNDA.n1698 GNDA.n1697 341.38
R2222 GNDA.n412 GNDA.n33 336
R2223 GNDA.n435 GNDA.n34 336
R2224 GNDA.n399 GNDA.n381 332.8
R2225 GNDA.n2467 GNDA.n61 332.8
R2226 GNDA.n453 GNDA.t270 332.75
R2227 GNDA.n451 GNDA.t273 332.75
R2228 GNDA.t248 GNDA.n166 172.876
R2229 GNDA.t229 GNDA.n623 327.661
R2230 GNDA.t229 GNDA.n624 327.661
R2231 GNDA.n1275 GNDA.t231 172.876
R2232 GNDA.n1214 GNDA.t231 172.876
R2233 GNDA.t248 GNDA.n170 172.876
R2234 GNDA.t248 GNDA.n171 172.615
R2235 GNDA.t229 GNDA.n590 323.404
R2236 GNDA.t229 GNDA.n1604 323.404
R2237 GNDA.n1274 GNDA.t231 172.615
R2238 GNDA.n691 GNDA.t231 172.615
R2239 GNDA.t248 GNDA.n116 172.615
R2240 GNDA.n1722 GNDA.n1721 323.2
R2241 GNDA.n1701 GNDA.n1700 322.861
R2242 GNDA.n401 GNDA.n400 321.281
R2243 GNDA.n2469 GNDA.n2468 321.281
R2244 GNDA.n400 GNDA.n399 318.08
R2245 GNDA.n2468 GNDA.n2467 318.08
R2246 GNDA.n1723 GNDA.n1722 316.8
R2247 GNDA.n489 GNDA.n488 310.401
R2248 GNDA.n373 GNDA.n332 310.401
R2249 GNDA.n2475 GNDA.n2474 310.401
R2250 GNDA.n43 GNDA.n38 310.401
R2251 GNDA.n2439 GNDA.n2438 304
R2252 GNDA.n379 GNDA.n330 304
R2253 GNDA.n45 GNDA.n39 304
R2254 GNDA.n2416 GNDA.n118 301.474
R2255 GNDA.n2438 GNDA.n98 300.8
R2256 GNDA.n2439 GNDA.n97 300.8
R2257 GNDA.n456 GNDA.n455 300.8
R2258 GNDA.n455 GNDA.n454 300.8
R2259 GNDA.n381 GNDA.n380 300.8
R2260 GNDA.n61 GNDA.n60 300.8
R2261 GNDA.n2161 GNDA.n514 297.601
R2262 GNDA.n2161 GNDA.n2160 297.601
R2263 GNDA.n98 GNDA.n97 297.601
R2264 GNDA.n2159 GNDA.n517 297.601
R2265 GNDA.n520 GNDA.n517 297.601
R2266 GNDA.n392 GNDA.n391 296
R2267 GNDA.n2462 GNDA.n67 296
R2268 GNDA.n1732 GNDA.n1731 294.401
R2269 GNDA.n1731 GNDA.n1730 294.401
R2270 GNDA.n1721 GNDA.n1635 294.401
R2271 GNDA.n2467 GNDA.n2466 292.5
R2272 GNDA.n2466 GNDA.n2465 292.5
R2273 GNDA.n2468 GNDA.n59 292.5
R2274 GNDA.n64 GNDA.n59 292.5
R2275 GNDA.n61 GNDA.n58 292.5
R2276 GNDA.n64 GNDA.n58 292.5
R2277 GNDA.n2459 GNDA.n2458 292.5
R2278 GNDA.n2458 GNDA.n2457 292.5
R2279 GNDA.n75 GNDA.n70 292.5
R2280 GNDA.n76 GNDA.n75 292.5
R2281 GNDA.n74 GNDA.n73 292.5
R2282 GNDA.n74 GNDA.n62 292.5
R2283 GNDA.n71 GNDA.n69 292.5
R2284 GNDA.n76 GNDA.n71 292.5
R2285 GNDA.n2463 GNDA.n2462 292.5
R2286 GNDA.n2464 GNDA.n2463 292.5
R2287 GNDA.n443 GNDA.n357 292.5
R2288 GNDA.n444 GNDA.n443 292.5
R2289 GNDA.n442 GNDA.n365 292.5
R2290 GNDA.n442 GNDA.n441 292.5
R2291 GNDA.n466 GNDA.n465 292.5
R2292 GNDA.n465 GNDA.n57 292.5
R2293 GNDA.n467 GNDA.n462 292.5
R2294 GNDA.n462 GNDA.n461 292.5
R2295 GNDA.n456 GNDA.n450 292.5
R2296 GNDA.n450 GNDA.n29 292.5
R2297 GNDA.n455 GNDA.n360 292.5
R2298 GNDA.n460 GNDA.n360 292.5
R2299 GNDA.n454 GNDA.n449 292.5
R2300 GNDA.n449 GNDA.n448 292.5
R2301 GNDA.n459 GNDA.n458 292.5
R2302 GNDA.n460 GNDA.n459 292.5
R2303 GNDA.n2494 GNDA.n2493 292.5
R2304 GNDA.n2493 GNDA.n2492 292.5
R2305 GNDA.n28 GNDA.n25 292.5
R2306 GNDA.n460 GNDA.n28 292.5
R2307 GNDA.n446 GNDA.n445 292.5
R2308 GNDA.n447 GNDA.n446 292.5
R2309 GNDA.n27 GNDA.n26 292.5
R2310 GNDA.n460 GNDA.n27 292.5
R2311 GNDA.n373 GNDA.n334 292.5
R2312 GNDA.n483 GNDA.n334 292.5
R2313 GNDA.n378 GNDA.n335 292.5
R2314 GNDA.n484 GNDA.n335 292.5
R2315 GNDA.n379 GNDA.n333 292.5
R2316 GNDA.n369 GNDA.n333 292.5
R2317 GNDA.n486 GNDA.n485 292.5
R2318 GNDA.n485 GNDA.n484 292.5
R2319 GNDA.n2490 GNDA.n2489 292.5
R2320 GNDA.n2491 GNDA.n2490 292.5
R2321 GNDA.n34 GNDA.n32 292.5
R2322 GNDA.n460 GNDA.n32 292.5
R2323 GNDA.n435 GNDA.n411 292.5
R2324 GNDA.n411 GNDA.n410 292.5
R2325 GNDA.n438 GNDA.n437 292.5
R2326 GNDA.n439 GNDA.n438 292.5
R2327 GNDA.n412 GNDA.n408 292.5
R2328 GNDA.n410 GNDA.n408 292.5
R2329 GNDA.n33 GNDA.n31 292.5
R2330 GNDA.n460 GNDA.n31 292.5
R2331 GNDA.n2470 GNDA.n2469 292.5
R2332 GNDA.n2471 GNDA.n2470 292.5
R2333 GNDA.n41 GNDA.n39 292.5
R2334 GNDA.n55 GNDA.n41 292.5
R2335 GNDA.n2481 GNDA.n2480 292.5
R2336 GNDA.n2480 GNDA.n2479 292.5
R2337 GNDA.n40 GNDA.n38 292.5
R2338 GNDA.n475 GNDA.n40 292.5
R2339 GNDA.n2478 GNDA.n2477 292.5
R2340 GNDA.n2479 GNDA.n2478 292.5
R2341 GNDA.n478 GNDA.n477 292.5
R2342 GNDA.n477 GNDA.n476 292.5
R2343 GNDA.n479 GNDA.n337 292.5
R2344 GNDA.n460 GNDA.n337 292.5
R2345 GNDA.n481 GNDA.n480 292.5
R2346 GNDA.n482 GNDA.n481 292.5
R2347 GNDA.n470 GNDA.n336 292.5
R2348 GNDA.n460 GNDA.n336 292.5
R2349 GNDA.n488 GNDA.n326 292.5
R2350 GNDA.t112 GNDA.n326 292.5
R2351 GNDA.n368 GNDA.n367 292.5
R2352 GNDA.t112 GNDA.n368 292.5
R2353 GNDA.n2475 GNDA.n48 292.5
R2354 GNDA.t83 GNDA.n48 292.5
R2355 GNDA.n54 GNDA.n53 292.5
R2356 GNDA.t83 GNDA.n54 292.5
R2357 GNDA.n402 GNDA.n401 292.5
R2358 GNDA.n403 GNDA.n402 292.5
R2359 GNDA.n400 GNDA.n372 292.5
R2360 GNDA.n382 GNDA.n372 292.5
R2361 GNDA.n399 GNDA.n398 292.5
R2362 GNDA.n398 GNDA.n397 292.5
R2363 GNDA.n381 GNDA.n371 292.5
R2364 GNDA.n382 GNDA.n371 292.5
R2365 GNDA.n321 GNDA.n318 292.5
R2366 GNDA.n388 GNDA.n318 292.5
R2367 GNDA.n395 GNDA.n322 292.5
R2368 GNDA.n396 GNDA.n395 292.5
R2369 GNDA.n492 GNDA.n319 292.5
R2370 GNDA.n388 GNDA.n319 292.5
R2371 GNDA.n494 GNDA.n493 292.5
R2372 GNDA.n495 GNDA.n494 292.5
R2373 GNDA.n391 GNDA.n390 292.5
R2374 GNDA.n390 GNDA.n389 292.5
R2375 GNDA.n2187 GNDA.n2186 292.5
R2376 GNDA.n2188 GNDA.n2187 292.5
R2377 GNDA.n2185 GNDA.n314 292.5
R2378 GNDA.n2156 GNDA.n314 292.5
R2379 GNDA.n2184 GNDA.n2183 292.5
R2380 GNDA.n2183 GNDA.n2182 292.5
R2381 GNDA.n315 GNDA.n313 292.5
R2382 GNDA.n2156 GNDA.n313 292.5
R2383 GNDA.n2177 GNDA.n2176 292.5
R2384 GNDA.n2176 GNDA.n2175 292.5
R2385 GNDA.n2179 GNDA.n498 292.5
R2386 GNDA.n2157 GNDA.n498 292.5
R2387 GNDA.n2181 GNDA.n2180 292.5
R2388 GNDA.n2182 GNDA.n2181 292.5
R2389 GNDA.n499 GNDA.n497 292.5
R2390 GNDA.n2157 GNDA.n497 292.5
R2391 GNDA.n103 GNDA.n100 292.5
R2392 GNDA.n103 GNDA.n102 292.5
R2393 GNDA.n107 GNDA.n106 292.5
R2394 GNDA.n2435 GNDA.n107 292.5
R2395 GNDA.n105 GNDA.n101 292.5
R2396 GNDA.n308 GNDA.n101 292.5
R2397 GNDA.n2437 GNDA.n2436 292.5
R2398 GNDA.n2436 GNDA.n2435 292.5
R2399 GNDA.n517 GNDA.n511 292.5
R2400 GNDA.n2163 GNDA.n511 292.5
R2401 GNDA.n521 GNDA.n520 292.5
R2402 GNDA.n2157 GNDA.n521 292.5
R2403 GNDA.n518 GNDA.n516 292.5
R2404 GNDA.n2130 GNDA.n518 292.5
R2405 GNDA.n2159 GNDA.n2158 292.5
R2406 GNDA.n2158 GNDA.n2157 292.5
R2407 GNDA.n2440 GNDA.n2439 292.5
R2408 GNDA.n2441 GNDA.n2440 292.5
R2409 GNDA.n2438 GNDA.n96 292.5
R2410 GNDA.n2435 GNDA.n96 292.5
R2411 GNDA.n167 GNDA.n98 292.5
R2412 GNDA.n168 GNDA.n167 292.5
R2413 GNDA.n97 GNDA.n95 292.5
R2414 GNDA.n2435 GNDA.n95 292.5
R2415 GNDA.n2162 GNDA.n2161 292.5
R2416 GNDA.n2163 GNDA.n2162 292.5
R2417 GNDA.n2160 GNDA.n513 292.5
R2418 GNDA.n2157 GNDA.n513 292.5
R2419 GNDA.n2129 GNDA.n515 292.5
R2420 GNDA.n2130 GNDA.n2129 292.5
R2421 GNDA.n514 GNDA.n512 292.5
R2422 GNDA.n2157 GNDA.n512 292.5
R2423 GNDA.n1724 GNDA.n1723 292.5
R2424 GNDA.n1725 GNDA.n1724 292.5
R2425 GNDA.n1722 GNDA.n1634 292.5
R2426 GNDA.n1711 GNDA.n1634 292.5
R2427 GNDA.n1721 GNDA.n1720 292.5
R2428 GNDA.n1720 GNDA.n1719 292.5
R2429 GNDA.n1635 GNDA.n1633 292.5
R2430 GNDA.n1711 GNDA.n1633 292.5
R2431 GNDA.n1699 GNDA.n1698 292.5
R2432 GNDA.n1702 GNDA.n1701 292.5
R2433 GNDA.n1648 GNDA.n1636 292.5
R2434 GNDA.n1650 GNDA.n1648 292.5
R2435 GNDA.n1644 GNDA.n1642 292.5
R2436 GNDA.n1691 GNDA.n1644 292.5
R2437 GNDA.n1646 GNDA.n1645 292.5
R2438 GNDA.n1702 GNDA.n1646 292.5
R2439 GNDA.n1643 GNDA.n1641 292.5
R2440 GNDA.n1649 GNDA.n1643 292.5
R2441 GNDA.n1704 GNDA.n1703 292.5
R2442 GNDA.n1703 GNDA.n1702 292.5
R2443 GNDA.n1696 GNDA.n1695 292.5
R2444 GNDA.n1697 GNDA.n1696 292.5
R2445 GNDA.n1637 GNDA.n1621 292.5
R2446 GNDA.n1736 GNDA.n1621 292.5
R2447 GNDA.n1693 GNDA.n1692 292.5
R2448 GNDA.n1692 GNDA.n1615 292.5
R2449 GNDA.n1694 GNDA.n1622 292.5
R2450 GNDA.n1736 GNDA.n1622 292.5
R2451 GNDA.n1729 GNDA.n1728 292.5
R2452 GNDA.n1728 GNDA.n1727 292.5
R2453 GNDA.n1712 GNDA.n1631 292.5
R2454 GNDA.n1713 GNDA.n1712 292.5
R2455 GNDA.n1717 GNDA.n1716 292.5
R2456 GNDA.n1718 GNDA.n1717 292.5
R2457 GNDA.n1732 GNDA.n1624 292.5
R2458 GNDA.n1651 GNDA.n1624 292.5
R2459 GNDA.n1731 GNDA.n1620 292.5
R2460 GNDA.n1736 GNDA.n1620 292.5
R2461 GNDA.n1730 GNDA.n1623 292.5
R2462 GNDA.n1726 GNDA.n1623 292.5
R2463 GNDA.n1735 GNDA.n1734 292.5
R2464 GNDA.n1736 GNDA.n1735 292.5
R2465 GNDA.n1684 GNDA.n1683 292.5
R2466 GNDA.n1685 GNDA.n1684 292.5
R2467 GNDA.n1682 GNDA.n1681 292.5
R2468 GNDA.n1681 GNDA.n1647 292.5
R2469 GNDA.n1653 GNDA.n1628 292.5
R2470 GNDA.n1653 GNDA.n1652 292.5
R2471 GNDA.n1739 GNDA.n1738 292.5
R2472 GNDA.n1738 GNDA.n1737 292.5
R2473 GNDA.n1740 GNDA.n1617 292.5
R2474 GNDA.n1711 GNDA.n1617 292.5
R2475 GNDA.n1742 GNDA.n1741 292.5
R2476 GNDA.n1743 GNDA.n1742 292.5
R2477 GNDA.n1618 GNDA.n1616 292.5
R2478 GNDA.n1711 GNDA.n1616 292.5
R2479 GNDA.n515 GNDA.n514 291.2
R2480 GNDA.n2160 GNDA.n515 291.2
R2481 GNDA.n2159 GNDA.n516 291.2
R2482 GNDA.n520 GNDA.n516 291.2
R2483 GNDA.n1723 GNDA.n1635 288
R2484 GNDA.n1658 GNDA.n1657 281.601
R2485 GNDA.n1715 GNDA.n1630 281.601
R2486 GNDA.n1683 GNDA.n1682 278.401
R2487 GNDA.n1716 GNDA.n1631 278.401
R2488 GNDA.n892 GNDA.t229 267.529
R2489 GNDA.t229 GNDA.n1441 267.529
R2490 GNDA.n1868 GNDA.t229 267.529
R2491 GNDA.n1697 GNDA.n1691 265.517
R2492 GNDA.n2293 GNDA.n282 259.416
R2493 GNDA.n2339 GNDA.n146 259.416
R2494 GNDA.n2065 GNDA.n573 259.416
R2495 GNDA.n1394 GNDA.n660 259.416
R2496 GNDA.n1854 GNDA.n609 259.416
R2497 GNDA.n1456 GNDA.n1421 259.416
R2498 GNDA.n880 GNDA.n879 259.416
R2499 GNDA.n963 GNDA.n962 259.416
R2500 GNDA.n1203 GNDA.n1082 259.416
R2501 GNDA.n453 GNDA.t272 258.601
R2502 GNDA.n451 GNDA.t275 258.601
R2503 GNDA.n1857 GNDA.n1856 254.494
R2504 GNDA.n881 GNDA.n753 254.392
R2505 GNDA.n1454 GNDA.n1453 254.392
R2506 GNDA.n1879 GNDA.n590 254.34
R2507 GNDA.n1885 GNDA.n590 254.34
R2508 GNDA.n1887 GNDA.n590 254.34
R2509 GNDA.n1893 GNDA.n590 254.34
R2510 GNDA.n1895 GNDA.n590 254.34
R2511 GNDA.n1901 GNDA.n590 254.34
R2512 GNDA.n1604 GNDA.n1603 254.34
R2513 GNDA.n1604 GNDA.n630 254.34
R2514 GNDA.n1604 GNDA.n629 254.34
R2515 GNDA.n1604 GNDA.n628 254.34
R2516 GNDA.n1604 GNDA.n627 254.34
R2517 GNDA.n1604 GNDA.n626 254.34
R2518 GNDA.n719 GNDA.n570 254.34
R2519 GNDA.n949 GNDA.n570 254.34
R2520 GNDA.n945 GNDA.n570 254.34
R2521 GNDA.n935 GNDA.n570 254.34
R2522 GNDA.n933 GNDA.n570 254.34
R2523 GNDA.n654 GNDA.n570 254.34
R2524 GNDA.n651 GNDA.n570 254.34
R2525 GNDA.n646 GNDA.n570 254.34
R2526 GNDA.n643 GNDA.n570 254.34
R2527 GNDA.n638 GNDA.n570 254.34
R2528 GNDA.n1936 GNDA.n1935 254.34
R2529 GNDA.n1934 GNDA.n570 254.34
R2530 GNDA.n1922 GNDA.n570 254.34
R2531 GNDA.n1921 GNDA.n570 254.34
R2532 GNDA.n582 GNDA.n570 254.34
R2533 GNDA.n1909 GNDA.n570 254.34
R2534 GNDA.n929 GNDA.n569 254.34
R2535 GNDA.n939 GNDA.n569 254.34
R2536 GNDA.n941 GNDA.n569 254.34
R2537 GNDA.n953 GNDA.n569 254.34
R2538 GNDA.n956 GNDA.n569 254.34
R2539 GNDA.n636 GNDA.n569 254.34
R2540 GNDA.n1573 GNDA.n569 254.34
R2541 GNDA.n1567 GNDA.n569 254.34
R2542 GNDA.n1565 GNDA.n569 254.34
R2543 GNDA.n1559 GNDA.n569 254.34
R2544 GNDA.n1904 GNDA.n569 254.34
R2545 GNDA.n1914 GNDA.n569 254.34
R2546 GNDA.n1916 GNDA.n569 254.34
R2547 GNDA.n1927 GNDA.n569 254.34
R2548 GNDA.n1930 GNDA.n569 254.34
R2549 GNDA.n1819 GNDA.n1818 254.34
R2550 GNDA.n1274 GNDA.n1273 254.34
R2551 GNDA.n1274 GNDA.n1219 254.34
R2552 GNDA.n1274 GNDA.n1218 254.34
R2553 GNDA.n1274 GNDA.n1217 254.34
R2554 GNDA.n1274 GNDA.n1216 254.34
R2555 GNDA.n1274 GNDA.n1215 254.34
R2556 GNDA.n691 GNDA.n690 254.34
R2557 GNDA.n691 GNDA.n665 254.34
R2558 GNDA.n691 GNDA.n664 254.34
R2559 GNDA.n691 GNDA.n663 254.34
R2560 GNDA.n691 GNDA.n662 254.34
R2561 GNDA.n691 GNDA.n661 254.34
R2562 GNDA.n2336 GNDA.n2335 254.34
R2563 GNDA.n2334 GNDA.n2333 254.34
R2564 GNDA.n2333 GNDA.n165 254.34
R2565 GNDA.n2333 GNDA.n164 254.34
R2566 GNDA.n2333 GNDA.n163 254.34
R2567 GNDA.n2333 GNDA.n162 254.34
R2568 GNDA.n2302 GNDA.n204 254.34
R2569 GNDA.n2302 GNDA.n203 254.34
R2570 GNDA.n2302 GNDA.n202 254.34
R2571 GNDA.n2302 GNDA.n201 254.34
R2572 GNDA.n2302 GNDA.n200 254.34
R2573 GNDA.n2028 GNDA.n2027 254.34
R2574 GNDA.n2333 GNDA.n160 254.34
R2575 GNDA.n2333 GNDA.n159 254.34
R2576 GNDA.n2333 GNDA.n158 254.34
R2577 GNDA.n2333 GNDA.n157 254.34
R2578 GNDA.n2333 GNDA.n156 254.34
R2579 GNDA.n2302 GNDA.n198 254.34
R2580 GNDA.n2302 GNDA.n197 254.34
R2581 GNDA.n2302 GNDA.n196 254.34
R2582 GNDA.n2302 GNDA.n195 254.34
R2583 GNDA.n2302 GNDA.n194 254.34
R2584 GNDA.n2333 GNDA.n155 254.34
R2585 GNDA.n1106 GNDA.n166 254.34
R2586 GNDA.n1180 GNDA.n166 254.34
R2587 GNDA.n1100 GNDA.n166 254.34
R2588 GNDA.n1191 GNDA.n166 254.34
R2589 GNDA.n1091 GNDA.n166 254.34
R2590 GNDA.n1202 GNDA.n166 254.34
R2591 GNDA.n961 GNDA.n718 254.34
R2592 GNDA.n1214 GNDA.n1213 254.34
R2593 GNDA.n1214 GNDA.n696 254.34
R2594 GNDA.n1214 GNDA.n695 254.34
R2595 GNDA.n1214 GNDA.n694 254.34
R2596 GNDA.n1214 GNDA.n693 254.34
R2597 GNDA.n1214 GNDA.n692 254.34
R2598 GNDA.n1209 GNDA.n1056 254.34
R2599 GNDA.n778 GNDA.n624 254.34
R2600 GNDA.n856 GNDA.n624 254.34
R2601 GNDA.n772 GNDA.n624 254.34
R2602 GNDA.n867 GNDA.n624 254.34
R2603 GNDA.n763 GNDA.n624 254.34
R2604 GNDA.n878 GNDA.n624 254.34
R2605 GNDA.n780 GNDA.n779 254.34
R2606 GNDA.n2333 GNDA.n154 254.34
R2607 GNDA.n2333 GNDA.n153 254.34
R2608 GNDA.n2333 GNDA.n152 254.34
R2609 GNDA.n2333 GNDA.n151 254.34
R2610 GNDA.n2333 GNDA.n150 254.34
R2611 GNDA.n2303 GNDA.n2302 254.34
R2612 GNDA.n2302 GNDA.n192 254.34
R2613 GNDA.n2302 GNDA.n191 254.34
R2614 GNDA.n2302 GNDA.n190 254.34
R2615 GNDA.n2302 GNDA.n189 254.34
R2616 GNDA.n2307 GNDA.n171 254.34
R2617 GNDA.n2313 GNDA.n171 254.34
R2618 GNDA.n2315 GNDA.n171 254.34
R2619 GNDA.n2321 GNDA.n171 254.34
R2620 GNDA.n2323 GNDA.n171 254.34
R2621 GNDA.n2329 GNDA.n171 254.34
R2622 GNDA.n2333 GNDA.n149 254.34
R2623 GNDA.n1396 GNDA.n658 254.34
R2624 GNDA.n1297 GNDA.n1275 254.34
R2625 GNDA.n1371 GNDA.n1275 254.34
R2626 GNDA.n1292 GNDA.n1275 254.34
R2627 GNDA.n1382 GNDA.n1275 254.34
R2628 GNDA.n1283 GNDA.n1275 254.34
R2629 GNDA.n1393 GNDA.n1275 254.34
R2630 GNDA.n2300 GNDA.n2299 254.34
R2631 GNDA.n1552 GNDA.n623 254.34
R2632 GNDA.n1468 GNDA.n623 254.34
R2633 GNDA.n1480 GNDA.n623 254.34
R2634 GNDA.n1466 GNDA.n623 254.34
R2635 GNDA.n1491 GNDA.n623 254.34
R2636 GNDA.n1457 GNDA.n623 254.34
R2637 GNDA.n1557 GNDA.n1556 254.34
R2638 GNDA.n306 GNDA.n170 254.34
R2639 GNDA.n2270 GNDA.n170 254.34
R2640 GNDA.n300 GNDA.n170 254.34
R2641 GNDA.n2281 GNDA.n170 254.34
R2642 GNDA.n291 GNDA.n170 254.34
R2643 GNDA.n2292 GNDA.n170 254.34
R2644 GNDA.n254 GNDA.n116 254.34
R2645 GNDA.n210 GNDA.n116 254.34
R2646 GNDA.n247 GNDA.n116 254.34
R2647 GNDA.n241 GNDA.n116 254.34
R2648 GNDA.n239 GNDA.n116 254.34
R2649 GNDA.n233 GNDA.n116 254.34
R2650 GNDA.n2153 GNDA.n2152 254.34
R2651 GNDA.n310 GNDA.n307 254.34
R2652 GNDA.n110 GNDA.n91 254.34
R2653 GNDA.n1743 GNDA.n1615 252.875
R2654 GNDA.n2085 GNDA.n554 250.349
R2655 GNDA.n2308 GNDA.n2306 249.663
R2656 GNDA.n255 GNDA.n161 249.663
R2657 GNDA.n1907 GNDA.n586 249.663
R2658 GNDA.n689 GNDA.n637 249.663
R2659 GNDA.n1880 GNDA.n1878 249.663
R2660 GNDA.n1602 GNDA.n632 249.663
R2661 GNDA.n902 GNDA.n741 249.663
R2662 GNDA.n932 GNDA.n567 249.663
R2663 GNDA.n2102 GNDA.n2101 249.663
R2664 GNDA.n2450 GNDA.n2449 248.049
R2665 GNDA.t229 GNDA.n891 244.762
R2666 GNDA.n1442 GNDA.t229 244.762
R2667 GNDA.t229 GNDA.n1867 244.762
R2668 GNDA.n2451 GNDA.n83 241.291
R2669 GNDA.n1682 GNDA.n1628 240
R2670 GNDA.n1729 GNDA.n1631 240
R2671 GNDA.n490 GNDA.n324 240
R2672 GNDA.n52 GNDA.n49 240
R2673 GNDA.n1840 GNDA.t229 239.004
R2674 GNDA.n1827 GNDA.n1744 239.004
R2675 GNDA.n2052 GNDA.t231 239.004
R2676 GNDA.t248 GNDA.n119 239.004
R2677 GNDA.n385 GNDA.n384 238.4
R2678 GNDA.n2461 GNDA.n68 238.4
R2679 GNDA.t140 GNDA.t274 236.923
R2680 GNDA.t339 GNDA.t215 236.923
R2681 GNDA.t330 GNDA.t205 236.923
R2682 GNDA.t239 GNDA.t213 236.923
R2683 GNDA.t201 GNDA.t290 236.923
R2684 GNDA.t207 GNDA.t25 236.923
R2685 GNDA.t5 GNDA.t197 236.923
R2686 GNDA.t332 GNDA.t271 236.923
R2687 GNDA.n437 GNDA.n412 233.601
R2688 GNDA.n352 GNDA.n350 227.096
R2689 GNDA.n349 GNDA.n347 227.096
R2690 GNDA.n352 GNDA.n351 226.534
R2691 GNDA.n349 GNDA.n348 226.534
R2692 GNDA.n331 GNDA.t312 224.525
R2693 GNDA.n329 GNDA.t227 224.525
R2694 GNDA.n44 GNDA.t259 224.525
R2695 GNDA.n42 GNDA.t269 224.525
R2696 GNDA.n2494 GNDA.n26 224
R2697 GNDA.n355 GNDA.n354 222.034
R2698 GNDA.n1533 GNDA.n1408 221.667
R2699 GNDA.n1350 GNDA.n1349 221.667
R2700 GNDA.n2249 GNDA.n2248 221.667
R2701 GNDA.n835 GNDA.n834 221.667
R2702 GNDA.n1035 GNDA.n1034 221.667
R2703 GNDA.n1159 GNDA.n1158 221.667
R2704 GNDA.n1802 GNDA.n1756 221.667
R2705 GNDA.n2011 GNDA.n1967 221.667
R2706 GNDA.n2394 GNDA.n2393 221.667
R2707 GNDA.n445 GNDA.n26 220.8
R2708 GNDA.n458 GNDA.n452 211.201
R2709 GNDA.n458 GNDA.n457 211.201
R2710 GNDA.n367 GNDA.n324 211.201
R2711 GNDA.n367 GNDA.n328 211.201
R2712 GNDA.n53 GNDA.n47 211.201
R2713 GNDA.n53 GNDA.n52 211.201
R2714 GNDA.n445 GNDA.n25 209.601
R2715 GNDA.n2495 GNDA.n2494 208
R2716 GNDA.n15 GNDA.n13 206.052
R2717 GNDA.n4 GNDA.n2 206.052
R2718 GNDA.n23 GNDA.n22 205.488
R2719 GNDA.n21 GNDA.n20 205.488
R2720 GNDA.n19 GNDA.n18 205.488
R2721 GNDA.n17 GNDA.n16 205.488
R2722 GNDA.n15 GNDA.n14 205.488
R2723 GNDA.n12 GNDA.n11 205.488
R2724 GNDA.n10 GNDA.n9 205.488
R2725 GNDA.n8 GNDA.n7 205.488
R2726 GNDA.n6 GNDA.n5 205.488
R2727 GNDA.n4 GNDA.n3 205.488
R2728 GNDA.n2442 GNDA.n2441 200.225
R2729 GNDA.n2196 GNDA.n2195 197
R2730 GNDA.n2443 GNDA.n92 197
R2731 GNDA.n2030 GNDA.n205 197
R2732 GNDA.n2301 GNDA.n207 197
R2733 GNDA.n1821 GNDA.n1820 197
R2734 GNDA.n1554 GNDA.n1398 197
R2735 GNDA.n782 GNDA.n781 197
R2736 GNDA.n698 GNDA.n206 197
R2737 GNDA.n2084 GNDA.n555 197
R2738 GNDA.n1105 GNDA.n524 197
R2739 GNDA.n77 GNDA.n68 195
R2740 GNDA.n78 GNDA.n77 195
R2741 GNDA.n67 GNDA.n66 195
R2742 GNDA.n66 GNDA.n65 195
R2743 GNDA.n393 GNDA.n392 195
R2744 GNDA.n394 GNDA.n393 195
R2745 GNDA.n386 GNDA.n384 195
R2746 GNDA.n387 GNDA.n386 195
R2747 GNDA.n486 GNDA.n332 192
R2748 GNDA.n2477 GNDA.n43 192
R2749 GNDA.n2331 GNDA.n175 187.249
R2750 GNDA.n232 GNDA.n231 187.249
R2751 GNDA.n1251 GNDA.n1250 187.249
R2752 GNDA.n2304 GNDA.n185 187.249
R2753 GNDA.n1905 GNDA.n1903 187.249
R2754 GNDA.n1579 GNDA.n1578 187.249
R2755 GNDA.n930 GNDA.n928 187.249
R2756 GNDA.n2099 GNDA.n2098 187.249
R2757 GNDA.n2132 GNDA.n2127 187.249
R2758 GNDA.n460 GNDA.t209 186.155
R2759 GNDA.n460 GNDA.t199 186.155
R2760 GNDA.n1498 GNDA.n1497 185
R2761 GNDA.n1499 GNDA.n1416 185
R2762 GNDA.n1416 GNDA.t228 185
R2763 GNDA.n1501 GNDA.n1500 185
R2764 GNDA.n1503 GNDA.n1415 185
R2765 GNDA.n1506 GNDA.n1505 185
R2766 GNDA.n1507 GNDA.n1414 185
R2767 GNDA.n1509 GNDA.n1508 185
R2768 GNDA.n1511 GNDA.n1413 185
R2769 GNDA.n1514 GNDA.n1513 185
R2770 GNDA.n1515 GNDA.n1412 185
R2771 GNDA.n1517 GNDA.n1516 185
R2772 GNDA.n1519 GNDA.n1411 185
R2773 GNDA.n1522 GNDA.n1521 185
R2774 GNDA.n1523 GNDA.n1410 185
R2775 GNDA.n1525 GNDA.n1524 185
R2776 GNDA.n1527 GNDA.n1409 185
R2777 GNDA.n1530 GNDA.n1529 185
R2778 GNDA.n1531 GNDA.n1408 185
R2779 GNDA.n1548 GNDA.n1547 185
R2780 GNDA.n1545 GNDA.n1402 185
R2781 GNDA.n1544 GNDA.n1404 185
R2782 GNDA.n1542 GNDA.n1541 185
R2783 GNDA.n1540 GNDA.n1405 185
R2784 GNDA.n1539 GNDA.n1538 185
R2785 GNDA.n1536 GNDA.n1406 185
R2786 GNDA.n1536 GNDA.t228 185
R2787 GNDA.n1535 GNDA.n1407 185
R2788 GNDA.n1533 GNDA.n1532 185
R2789 GNDA.n1316 GNDA.n1315 185
R2790 GNDA.n1317 GNDA.n1314 185
R2791 GNDA.n1317 GNDA.t230 185
R2792 GNDA.n1320 GNDA.n1319 185
R2793 GNDA.n1321 GNDA.n1313 185
R2794 GNDA.n1323 GNDA.n1322 185
R2795 GNDA.n1325 GNDA.n1312 185
R2796 GNDA.n1328 GNDA.n1327 185
R2797 GNDA.n1329 GNDA.n1311 185
R2798 GNDA.n1331 GNDA.n1330 185
R2799 GNDA.n1333 GNDA.n1310 185
R2800 GNDA.n1336 GNDA.n1335 185
R2801 GNDA.n1337 GNDA.n1309 185
R2802 GNDA.n1339 GNDA.n1338 185
R2803 GNDA.n1341 GNDA.n1308 185
R2804 GNDA.n1344 GNDA.n1343 185
R2805 GNDA.n1345 GNDA.n1307 185
R2806 GNDA.n1347 GNDA.n1346 185
R2807 GNDA.n1349 GNDA.n1306 185
R2808 GNDA.n1366 GNDA.n1301 185
R2809 GNDA.n1364 GNDA.n1363 185
R2810 GNDA.n1362 GNDA.n1302 185
R2811 GNDA.n1361 GNDA.n1360 185
R2812 GNDA.n1358 GNDA.n1303 185
R2813 GNDA.n1356 GNDA.n1355 185
R2814 GNDA.n1354 GNDA.n1304 185
R2815 GNDA.n1304 GNDA.t230 185
R2816 GNDA.n1353 GNDA.n1352 185
R2817 GNDA.n1350 GNDA.n1305 185
R2818 GNDA.n2215 GNDA.n2214 185
R2819 GNDA.n2216 GNDA.n2213 185
R2820 GNDA.n2216 GNDA.t313 185
R2821 GNDA.n2219 GNDA.n2218 185
R2822 GNDA.n2220 GNDA.n2212 185
R2823 GNDA.n2222 GNDA.n2221 185
R2824 GNDA.n2224 GNDA.n2211 185
R2825 GNDA.n2227 GNDA.n2226 185
R2826 GNDA.n2228 GNDA.n2210 185
R2827 GNDA.n2230 GNDA.n2229 185
R2828 GNDA.n2232 GNDA.n2209 185
R2829 GNDA.n2235 GNDA.n2234 185
R2830 GNDA.n2236 GNDA.n2208 185
R2831 GNDA.n2238 GNDA.n2237 185
R2832 GNDA.n2240 GNDA.n2207 185
R2833 GNDA.n2243 GNDA.n2242 185
R2834 GNDA.n2244 GNDA.n2206 185
R2835 GNDA.n2246 GNDA.n2245 185
R2836 GNDA.n2248 GNDA.n2205 185
R2837 GNDA.n2265 GNDA.n2200 185
R2838 GNDA.n2263 GNDA.n2262 185
R2839 GNDA.n2261 GNDA.n2201 185
R2840 GNDA.n2260 GNDA.n2259 185
R2841 GNDA.n2257 GNDA.n2202 185
R2842 GNDA.n2255 GNDA.n2254 185
R2843 GNDA.n2253 GNDA.n2203 185
R2844 GNDA.n2203 GNDA.t313 185
R2845 GNDA.n2252 GNDA.n2251 185
R2846 GNDA.n2249 GNDA.n2204 185
R2847 GNDA.n801 GNDA.n800 185
R2848 GNDA.n802 GNDA.n799 185
R2849 GNDA.n802 GNDA.t279 185
R2850 GNDA.n805 GNDA.n804 185
R2851 GNDA.n806 GNDA.n798 185
R2852 GNDA.n808 GNDA.n807 185
R2853 GNDA.n810 GNDA.n797 185
R2854 GNDA.n813 GNDA.n812 185
R2855 GNDA.n814 GNDA.n796 185
R2856 GNDA.n816 GNDA.n815 185
R2857 GNDA.n818 GNDA.n795 185
R2858 GNDA.n821 GNDA.n820 185
R2859 GNDA.n822 GNDA.n794 185
R2860 GNDA.n824 GNDA.n823 185
R2861 GNDA.n826 GNDA.n793 185
R2862 GNDA.n829 GNDA.n828 185
R2863 GNDA.n830 GNDA.n792 185
R2864 GNDA.n832 GNDA.n831 185
R2865 GNDA.n834 GNDA.n791 185
R2866 GNDA.n851 GNDA.n786 185
R2867 GNDA.n849 GNDA.n848 185
R2868 GNDA.n847 GNDA.n787 185
R2869 GNDA.n846 GNDA.n845 185
R2870 GNDA.n843 GNDA.n788 185
R2871 GNDA.n841 GNDA.n840 185
R2872 GNDA.n839 GNDA.n789 185
R2873 GNDA.n789 GNDA.t279 185
R2874 GNDA.n838 GNDA.n837 185
R2875 GNDA.n835 GNDA.n790 185
R2876 GNDA.n1001 GNDA.n716 185
R2877 GNDA.n1002 GNDA.n715 185
R2878 GNDA.n1002 GNDA.t283 185
R2879 GNDA.n1005 GNDA.n1004 185
R2880 GNDA.n1006 GNDA.n714 185
R2881 GNDA.n1008 GNDA.n1007 185
R2882 GNDA.n1010 GNDA.n713 185
R2883 GNDA.n1013 GNDA.n1012 185
R2884 GNDA.n1014 GNDA.n712 185
R2885 GNDA.n1016 GNDA.n1015 185
R2886 GNDA.n1018 GNDA.n711 185
R2887 GNDA.n1021 GNDA.n1020 185
R2888 GNDA.n1022 GNDA.n710 185
R2889 GNDA.n1024 GNDA.n1023 185
R2890 GNDA.n1026 GNDA.n709 185
R2891 GNDA.n1029 GNDA.n1028 185
R2892 GNDA.n1030 GNDA.n708 185
R2893 GNDA.n1032 GNDA.n1031 185
R2894 GNDA.n1034 GNDA.n707 185
R2895 GNDA.n1051 GNDA.n699 185
R2896 GNDA.n1049 GNDA.n1048 185
R2897 GNDA.n1047 GNDA.n703 185
R2898 GNDA.n1046 GNDA.n1045 185
R2899 GNDA.n1043 GNDA.n704 185
R2900 GNDA.n1041 GNDA.n1040 185
R2901 GNDA.n1039 GNDA.n705 185
R2902 GNDA.n705 GNDA.t283 185
R2903 GNDA.n1038 GNDA.n1037 185
R2904 GNDA.n1035 GNDA.n706 185
R2905 GNDA.n1125 GNDA.n1124 185
R2906 GNDA.n1126 GNDA.n1123 185
R2907 GNDA.n1126 GNDA.t261 185
R2908 GNDA.n1129 GNDA.n1128 185
R2909 GNDA.n1130 GNDA.n1122 185
R2910 GNDA.n1132 GNDA.n1131 185
R2911 GNDA.n1134 GNDA.n1121 185
R2912 GNDA.n1137 GNDA.n1136 185
R2913 GNDA.n1138 GNDA.n1120 185
R2914 GNDA.n1140 GNDA.n1139 185
R2915 GNDA.n1142 GNDA.n1119 185
R2916 GNDA.n1145 GNDA.n1144 185
R2917 GNDA.n1146 GNDA.n1118 185
R2918 GNDA.n1148 GNDA.n1147 185
R2919 GNDA.n1150 GNDA.n1117 185
R2920 GNDA.n1153 GNDA.n1152 185
R2921 GNDA.n1154 GNDA.n1116 185
R2922 GNDA.n1156 GNDA.n1155 185
R2923 GNDA.n1158 GNDA.n1115 185
R2924 GNDA.n1175 GNDA.n1110 185
R2925 GNDA.n1173 GNDA.n1172 185
R2926 GNDA.n1171 GNDA.n1111 185
R2927 GNDA.n1170 GNDA.n1169 185
R2928 GNDA.n1167 GNDA.n1112 185
R2929 GNDA.n1165 GNDA.n1164 185
R2930 GNDA.n1163 GNDA.n1113 185
R2931 GNDA.n1113 GNDA.t261 185
R2932 GNDA.n1162 GNDA.n1161 185
R2933 GNDA.n1159 GNDA.n1114 185
R2934 GNDA.n1767 GNDA.n1766 185
R2935 GNDA.n1768 GNDA.n1764 185
R2936 GNDA.n1764 GNDA.t260 185
R2937 GNDA.n1770 GNDA.n1769 185
R2938 GNDA.n1772 GNDA.n1763 185
R2939 GNDA.n1775 GNDA.n1774 185
R2940 GNDA.n1776 GNDA.n1762 185
R2941 GNDA.n1778 GNDA.n1777 185
R2942 GNDA.n1780 GNDA.n1761 185
R2943 GNDA.n1783 GNDA.n1782 185
R2944 GNDA.n1784 GNDA.n1760 185
R2945 GNDA.n1786 GNDA.n1785 185
R2946 GNDA.n1788 GNDA.n1759 185
R2947 GNDA.n1791 GNDA.n1790 185
R2948 GNDA.n1792 GNDA.n1758 185
R2949 GNDA.n1794 GNDA.n1793 185
R2950 GNDA.n1796 GNDA.n1757 185
R2951 GNDA.n1799 GNDA.n1798 185
R2952 GNDA.n1800 GNDA.n1756 185
R2953 GNDA.n1817 GNDA.n1816 185
R2954 GNDA.n1814 GNDA.n1749 185
R2955 GNDA.n1813 GNDA.n1752 185
R2956 GNDA.n1811 GNDA.n1810 185
R2957 GNDA.n1809 GNDA.n1753 185
R2958 GNDA.n1808 GNDA.n1807 185
R2959 GNDA.n1805 GNDA.n1754 185
R2960 GNDA.n1805 GNDA.t260 185
R2961 GNDA.n1804 GNDA.n1755 185
R2962 GNDA.n1802 GNDA.n1801 185
R2963 GNDA.n1975 GNDA.n1937 185
R2964 GNDA.n1977 GNDA.n1976 185
R2965 GNDA.n1976 GNDA.t262 185
R2966 GNDA.n1979 GNDA.n1978 185
R2967 GNDA.n1981 GNDA.n1974 185
R2968 GNDA.n1984 GNDA.n1983 185
R2969 GNDA.n1985 GNDA.n1973 185
R2970 GNDA.n1987 GNDA.n1986 185
R2971 GNDA.n1989 GNDA.n1972 185
R2972 GNDA.n1992 GNDA.n1991 185
R2973 GNDA.n1993 GNDA.n1971 185
R2974 GNDA.n1995 GNDA.n1994 185
R2975 GNDA.n1997 GNDA.n1970 185
R2976 GNDA.n2000 GNDA.n1999 185
R2977 GNDA.n2001 GNDA.n1969 185
R2978 GNDA.n2003 GNDA.n2002 185
R2979 GNDA.n2005 GNDA.n1968 185
R2980 GNDA.n2008 GNDA.n2007 185
R2981 GNDA.n2009 GNDA.n1967 185
R2982 GNDA.n2026 GNDA.n2025 185
R2983 GNDA.n2023 GNDA.n1960 185
R2984 GNDA.n2022 GNDA.n1963 185
R2985 GNDA.n2020 GNDA.n2019 185
R2986 GNDA.n2018 GNDA.n1964 185
R2987 GNDA.n2017 GNDA.n2016 185
R2988 GNDA.n2014 GNDA.n1965 185
R2989 GNDA.n2014 GNDA.t262 185
R2990 GNDA.n2013 GNDA.n1966 185
R2991 GNDA.n2011 GNDA.n2010 185
R2992 GNDA.n2360 GNDA.n139 185
R2993 GNDA.n2361 GNDA.n138 185
R2994 GNDA.n2361 GNDA.t247 185
R2995 GNDA.n2364 GNDA.n2363 185
R2996 GNDA.n2365 GNDA.n137 185
R2997 GNDA.n2367 GNDA.n2366 185
R2998 GNDA.n2369 GNDA.n136 185
R2999 GNDA.n2372 GNDA.n2371 185
R3000 GNDA.n2373 GNDA.n135 185
R3001 GNDA.n2375 GNDA.n2374 185
R3002 GNDA.n2377 GNDA.n134 185
R3003 GNDA.n2380 GNDA.n2379 185
R3004 GNDA.n2381 GNDA.n133 185
R3005 GNDA.n2383 GNDA.n2382 185
R3006 GNDA.n2385 GNDA.n132 185
R3007 GNDA.n2388 GNDA.n2387 185
R3008 GNDA.n2389 GNDA.n131 185
R3009 GNDA.n2391 GNDA.n2390 185
R3010 GNDA.n2393 GNDA.n130 185
R3011 GNDA.n2410 GNDA.n90 185
R3012 GNDA.n2408 GNDA.n2407 185
R3013 GNDA.n2406 GNDA.n126 185
R3014 GNDA.n2405 GNDA.n2404 185
R3015 GNDA.n2402 GNDA.n127 185
R3016 GNDA.n2400 GNDA.n2399 185
R3017 GNDA.n2398 GNDA.n128 185
R3018 GNDA.n128 GNDA.t247 185
R3019 GNDA.n2397 GNDA.n2396 185
R3020 GNDA.n2394 GNDA.n129 185
R3021 GNDA.n2411 GNDA.n89 185
R3022 GNDA.n2415 GNDA.n2413 185
R3023 GNDA.n2420 GNDA.n2419 185
R3024 GNDA.n2423 GNDA.n2422 185
R3025 GNDA.n125 GNDA.n123 185
R3026 GNDA.n2349 GNDA.n2348 185
R3027 GNDA.n2346 GNDA.n2343 185
R3028 GNDA.n142 GNDA.n140 185
R3029 GNDA.n2358 GNDA.n2357 185
R3030 GNDA.n1962 GNDA.n1959 185
R3031 GNDA.n1951 GNDA.n1949 185
R3032 GNDA.n2042 GNDA.n2041 185
R3033 GNDA.n2044 GNDA.n1948 185
R3034 GNDA.n2046 GNDA.n2045 185
R3035 GNDA.n1943 GNDA.n1941 185
R3036 GNDA.n2057 GNDA.n2056 185
R3037 GNDA.n2059 GNDA.n1940 185
R3038 GNDA.n2061 GNDA.n2060 185
R3039 GNDA.n1751 GNDA.n1748 185
R3040 GNDA.n1613 GNDA.n1612 185
R3041 GNDA.n1833 GNDA.n1832 185
R3042 GNDA.n1836 GNDA.n1835 185
R3043 GNDA.n1611 GNDA.n1608 185
R3044 GNDA.n619 GNDA.n618 185
R3045 GNDA.n1845 GNDA.n1844 185
R3046 GNDA.n1848 GNDA.n1847 185
R3047 GNDA.n617 GNDA.n615 185
R3048 GNDA.n1177 GNDA.n1176 185
R3049 GNDA.n1099 GNDA.n1097 185
R3050 GNDA.n1184 GNDA.n1183 185
R3051 GNDA.n1186 GNDA.n1096 185
R3052 GNDA.n1188 GNDA.n1187 185
R3053 GNDA.n1090 GNDA.n1088 185
R3054 GNDA.n1195 GNDA.n1194 185
R3055 GNDA.n1197 GNDA.n1087 185
R3056 GNDA.n1199 GNDA.n1198 185
R3057 GNDA.n1053 GNDA.n1052 185
R3058 GNDA.n976 GNDA.n975 185
R3059 GNDA.n974 GNDA.n972 185
R3060 GNDA.n981 GNDA.n971 185
R3061 GNDA.n986 GNDA.n985 185
R3062 GNDA.n989 GNDA.n988 185
R3063 GNDA.n970 GNDA.n967 185
R3064 GNDA.n994 GNDA.n717 185
R3065 GNDA.n999 GNDA.n998 185
R3066 GNDA.n853 GNDA.n852 185
R3067 GNDA.n771 GNDA.n769 185
R3068 GNDA.n860 GNDA.n859 185
R3069 GNDA.n862 GNDA.n768 185
R3070 GNDA.n864 GNDA.n863 185
R3071 GNDA.n762 GNDA.n760 185
R3072 GNDA.n871 GNDA.n870 185
R3073 GNDA.n873 GNDA.n759 185
R3074 GNDA.n875 GNDA.n874 185
R3075 GNDA.n2267 GNDA.n2266 185
R3076 GNDA.n299 GNDA.n297 185
R3077 GNDA.n2274 GNDA.n2273 185
R3078 GNDA.n2276 GNDA.n296 185
R3079 GNDA.n2278 GNDA.n2277 185
R3080 GNDA.n290 GNDA.n288 185
R3081 GNDA.n2285 GNDA.n2284 185
R3082 GNDA.n2287 GNDA.n287 185
R3083 GNDA.n2289 GNDA.n2288 185
R3084 GNDA.n1368 GNDA.n1367 185
R3085 GNDA.n1291 GNDA.n1289 185
R3086 GNDA.n1375 GNDA.n1374 185
R3087 GNDA.n1377 GNDA.n1288 185
R3088 GNDA.n1379 GNDA.n1378 185
R3089 GNDA.n1282 GNDA.n1280 185
R3090 GNDA.n1386 GNDA.n1385 185
R3091 GNDA.n1388 GNDA.n1279 185
R3092 GNDA.n1390 GNDA.n1389 185
R3093 GNDA.n1403 GNDA.n1401 185
R3094 GNDA.n1475 GNDA.n1473 185
R3095 GNDA.n1477 GNDA.n1476 185
R3096 GNDA.n1465 GNDA.n1463 185
R3097 GNDA.n1484 GNDA.n1483 185
R3098 GNDA.n1486 GNDA.n1462 185
R3099 GNDA.n1488 GNDA.n1487 185
R3100 GNDA.n1420 GNDA.n1418 185
R3101 GNDA.n1495 GNDA.n1494 185
R3102 GNDA.n492 GNDA.n491 182.4
R3103 GNDA.n72 GNDA.n70 182.4
R3104 GNDA.n2068 GNDA.n2067 181.233
R3105 GNDA.n2103 GNDA.n145 181.233
R3106 GNDA.t252 GNDA.n483 181.226
R3107 GNDA.n475 GNDA.t223 181.226
R3108 GNDA.n1700 GNDA.n1636 179.917
R3109 GNDA.n1734 GNDA.n1626 176
R3110 GNDA.n1734 GNDA.n1733 176
R3111 GNDA.n2291 GNDA.n284 175.546
R3112 GNDA.n2282 GNDA.n292 175.546
R3113 GNDA.n2280 GNDA.n293 175.546
R3114 GNDA.n2271 GNDA.n301 175.546
R3115 GNDA.n2269 GNDA.n302 175.546
R3116 GNDA.n505 GNDA.n175 175.546
R3117 GNDA.n509 GNDA.n505 175.546
R3118 GNDA.n509 GNDA.n503 175.546
R3119 GNDA.n2167 GNDA.n503 175.546
R3120 GNDA.n2167 GNDA.n500 175.546
R3121 GNDA.n2173 GNDA.n500 175.546
R3122 GNDA.n2173 GNDA.n501 175.546
R3123 GNDA.n501 GNDA.n309 175.546
R3124 GNDA.n2191 GNDA.n309 175.546
R3125 GNDA.n2192 GNDA.n2191 175.546
R3126 GNDA.n2312 GNDA.n181 175.546
R3127 GNDA.n2316 GNDA.n2314 175.546
R3128 GNDA.n2320 GNDA.n179 175.546
R3129 GNDA.n2324 GNDA.n2322 175.546
R3130 GNDA.n2328 GNDA.n177 175.546
R3131 GNDA.n259 GNDA.n258 175.546
R3132 GNDA.n264 GNDA.n263 175.546
R3133 GNDA.n270 GNDA.n269 175.546
R3134 GNDA.n276 GNDA.n275 175.546
R3135 GNDA.n2296 GNDA.n2295 175.546
R3136 GNDA.n2339 GNDA.n143 175.546
R3137 GNDA.n2355 GNDA.n143 175.546
R3138 GNDA.n2355 GNDA.n144 175.546
R3139 GNDA.n2351 GNDA.n144 175.546
R3140 GNDA.n2351 GNDA.n121 175.546
R3141 GNDA.n2425 GNDA.n121 175.546
R3142 GNDA.n2425 GNDA.n122 175.546
R3143 GNDA.n2417 GNDA.n122 175.546
R3144 GNDA.n2417 GNDA.n87 175.546
R3145 GNDA.n2448 GNDA.n87 175.546
R3146 GNDA.n2448 GNDA.n88 175.546
R3147 GNDA.n231 GNDA.n217 175.546
R3148 GNDA.n227 GNDA.n217 175.546
R3149 GNDA.n227 GNDA.n220 175.546
R3150 GNDA.n223 GNDA.n220 175.546
R3151 GNDA.n223 GNDA.n115 175.546
R3152 GNDA.n2428 GNDA.n115 175.546
R3153 GNDA.n2428 GNDA.n109 175.546
R3154 GNDA.n2433 GNDA.n109 175.546
R3155 GNDA.n2433 GNDA.n113 175.546
R3156 GNDA.n113 GNDA.n112 175.546
R3157 GNDA.n253 GNDA.n252 175.546
R3158 GNDA.n249 GNDA.n248 175.546
R3159 GNDA.n246 GNDA.n212 175.546
R3160 GNDA.n242 GNDA.n240 175.546
R3161 GNDA.n238 GNDA.n214 175.546
R3162 GNDA.n1223 GNDA.n161 175.546
R3163 GNDA.n1225 GNDA.n1224 175.546
R3164 GNDA.n1227 GNDA.n1226 175.546
R3165 GNDA.n1229 GNDA.n1228 175.546
R3166 GNDA.n1230 GNDA.n148 175.546
R3167 GNDA.n2065 GNDA.n574 175.546
R3168 GNDA.n2049 GNDA.n574 175.546
R3169 GNDA.n2049 GNDA.n1944 175.546
R3170 GNDA.n2054 GNDA.n1944 175.546
R3171 GNDA.n2054 GNDA.n2048 175.546
R3172 GNDA.n2048 GNDA.n1945 175.546
R3173 GNDA.n1952 GNDA.n1945 175.546
R3174 GNDA.n2039 GNDA.n1952 175.546
R3175 GNDA.n2039 GNDA.n1953 175.546
R3176 GNDA.n2035 GNDA.n1953 175.546
R3177 GNDA.n2035 GNDA.n1957 175.546
R3178 GNDA.n1247 GNDA.n1246 175.546
R3179 GNDA.n1243 GNDA.n1242 175.546
R3180 GNDA.n1239 GNDA.n1238 175.546
R3181 GNDA.n1235 GNDA.n1234 175.546
R3182 GNDA.n1231 GNDA.n199 175.546
R3183 GNDA.n1272 GNDA.n1220 175.546
R3184 GNDA.n1268 GNDA.n1267 175.546
R3185 GNDA.n1264 GNDA.n1263 175.546
R3186 GNDA.n1260 GNDA.n1259 175.546
R3187 GNDA.n1256 GNDA.n1255 175.546
R3188 GNDA.n1908 GNDA.n1907 175.546
R3189 GNDA.n1911 GNDA.n1910 175.546
R3190 GNDA.n1920 GNDA.n1919 175.546
R3191 GNDA.n1924 GNDA.n1923 175.546
R3192 GNDA.n1933 GNDA.n576 175.546
R3193 GNDA.n1392 GNDA.n1276 175.546
R3194 GNDA.n1383 GNDA.n1284 175.546
R3195 GNDA.n1381 GNDA.n1285 175.546
R3196 GNDA.n1372 GNDA.n1293 175.546
R3197 GNDA.n1370 GNDA.n1294 175.546
R3198 GNDA.n260 GNDA.n186 175.546
R3199 GNDA.n266 GNDA.n265 175.546
R3200 GNDA.n272 GNDA.n271 175.546
R3201 GNDA.n278 GNDA.n277 175.546
R3202 GNDA.n280 GNDA.n188 175.546
R3203 GNDA.n685 GNDA.n666 175.546
R3204 GNDA.n683 GNDA.n682 175.546
R3205 GNDA.n679 GNDA.n678 175.546
R3206 GNDA.n675 GNDA.n674 175.546
R3207 GNDA.n671 GNDA.n670 175.546
R3208 GNDA.n642 GNDA.n639 175.546
R3209 GNDA.n645 GNDA.n644 175.546
R3210 GNDA.n650 GNDA.n647 175.546
R3211 GNDA.n653 GNDA.n652 175.546
R3212 GNDA.n657 GNDA.n655 175.546
R3213 GNDA.n1854 GNDA.n611 175.546
R3214 GNDA.n1850 GNDA.n611 175.546
R3215 GNDA.n1850 GNDA.n613 175.546
R3216 GNDA.n1842 GNDA.n613 175.546
R3217 GNDA.n1842 GNDA.n620 175.546
R3218 GNDA.n1838 GNDA.n620 175.546
R3219 GNDA.n1838 GNDA.n1606 175.546
R3220 GNDA.n1830 GNDA.n1606 175.546
R3221 GNDA.n1830 GNDA.n1614 175.546
R3222 GNDA.n1826 GNDA.n1614 175.546
R3223 GNDA.n1826 GNDA.n1746 175.546
R3224 GNDA.n1913 GNDA.n584 175.546
R3225 GNDA.n1917 GNDA.n1915 175.546
R3226 GNDA.n1926 GNDA.n580 175.546
R3227 GNDA.n1929 GNDA.n1928 175.546
R3228 GNDA.n1931 GNDA.n578 175.546
R3229 GNDA.n1884 GNDA.n595 175.546
R3230 GNDA.n1888 GNDA.n1886 175.546
R3231 GNDA.n1892 GNDA.n593 175.546
R3232 GNDA.n1896 GNDA.n1894 175.546
R3233 GNDA.n1900 GNDA.n591 175.546
R3234 GNDA.n1878 GNDA.n597 175.546
R3235 GNDA.n1874 GNDA.n597 175.546
R3236 GNDA.n1874 GNDA.n600 175.546
R3237 GNDA.n1870 GNDA.n600 175.546
R3238 GNDA.n1870 GNDA.n603 175.546
R3239 GNDA.n1866 GNDA.n603 175.546
R3240 GNDA.n1866 GNDA.n605 175.546
R3241 GNDA.n1862 GNDA.n605 175.546
R3242 GNDA.n1862 GNDA.n607 175.546
R3243 GNDA.n1858 GNDA.n607 175.546
R3244 GNDA.n1492 GNDA.n1458 175.546
R3245 GNDA.n1490 GNDA.n1459 175.546
R3246 GNDA.n1481 GNDA.n1467 175.546
R3247 GNDA.n1479 GNDA.n1469 175.546
R3248 GNDA.n1551 GNDA.n1400 175.546
R3249 GNDA.n1575 GNDA.n1574 175.546
R3250 GNDA.n1572 GNDA.n641 175.546
R3251 GNDA.n1568 GNDA.n1566 175.546
R3252 GNDA.n1564 GNDA.n649 175.546
R3253 GNDA.n1560 GNDA.n1558 175.546
R3254 GNDA.n1598 GNDA.n631 175.546
R3255 GNDA.n1596 GNDA.n1595 175.546
R3256 GNDA.n1592 GNDA.n1591 175.546
R3257 GNDA.n1588 GNDA.n1587 175.546
R3258 GNDA.n1584 GNDA.n1583 175.546
R3259 GNDA.n1431 GNDA.n632 175.546
R3260 GNDA.n1435 GNDA.n1431 175.546
R3261 GNDA.n1435 GNDA.n1429 175.546
R3262 GNDA.n1439 GNDA.n1429 175.546
R3263 GNDA.n1439 GNDA.n1427 175.546
R3264 GNDA.n1443 GNDA.n1427 175.546
R3265 GNDA.n1443 GNDA.n1425 175.546
R3266 GNDA.n1447 GNDA.n1425 175.546
R3267 GNDA.n1447 GNDA.n1423 175.546
R3268 GNDA.n1452 GNDA.n1423 175.546
R3269 GNDA.n877 GNDA.n755 175.546
R3270 GNDA.n868 GNDA.n764 175.546
R3271 GNDA.n866 GNDA.n765 175.546
R3272 GNDA.n857 GNDA.n773 175.546
R3273 GNDA.n855 GNDA.n774 175.546
R3274 GNDA.n902 GNDA.n743 175.546
R3275 GNDA.n898 GNDA.n743 175.546
R3276 GNDA.n898 GNDA.n745 175.546
R3277 GNDA.n894 GNDA.n745 175.546
R3278 GNDA.n894 GNDA.n747 175.546
R3279 GNDA.n890 GNDA.n747 175.546
R3280 GNDA.n890 GNDA.n749 175.546
R3281 GNDA.n886 GNDA.n749 175.546
R3282 GNDA.n886 GNDA.n751 175.546
R3283 GNDA.n882 GNDA.n751 175.546
R3284 GNDA.n938 GNDA.n728 175.546
R3285 GNDA.n942 GNDA.n940 175.546
R3286 GNDA.n952 GNDA.n724 175.546
R3287 GNDA.n955 GNDA.n954 175.546
R3288 GNDA.n957 GNDA.n722 175.546
R3289 GNDA.n906 GNDA.n741 175.546
R3290 GNDA.n906 GNDA.n739 175.546
R3291 GNDA.n911 GNDA.n739 175.546
R3292 GNDA.n911 GNDA.n737 175.546
R3293 GNDA.n915 GNDA.n737 175.546
R3294 GNDA.n916 GNDA.n915 175.546
R3295 GNDA.n918 GNDA.n916 175.546
R3296 GNDA.n918 GNDA.n735 175.546
R3297 GNDA.n923 GNDA.n735 175.546
R3298 GNDA.n923 GNDA.n731 175.546
R3299 GNDA.n927 GNDA.n731 175.546
R3300 GNDA.n996 GNDA.n995 175.546
R3301 GNDA.n992 GNDA.n991 175.546
R3302 GNDA.n983 GNDA.n982 175.546
R3303 GNDA.n979 GNDA.n978 175.546
R3304 GNDA.n700 GNDA.n697 175.546
R3305 GNDA.n936 GNDA.n934 175.546
R3306 GNDA.n944 GNDA.n726 175.546
R3307 GNDA.n950 GNDA.n946 175.546
R3308 GNDA.n948 GNDA.n947 175.546
R3309 GNDA.n960 GNDA.n959 175.546
R3310 GNDA.n1060 GNDA.n1059 175.546
R3311 GNDA.n1066 GNDA.n1065 175.546
R3312 GNDA.n1072 GNDA.n1071 175.546
R3313 GNDA.n1078 GNDA.n1077 175.546
R3314 GNDA.n1080 GNDA.n193 175.546
R3315 GNDA.n2070 GNDA.n567 175.546
R3316 GNDA.n2070 GNDA.n565 175.546
R3317 GNDA.n2074 GNDA.n565 175.546
R3318 GNDA.n2074 GNDA.n563 175.546
R3319 GNDA.n2078 GNDA.n563 175.546
R3320 GNDA.n2078 GNDA.n553 175.546
R3321 GNDA.n2088 GNDA.n553 175.546
R3322 GNDA.n2088 GNDA.n551 175.546
R3323 GNDA.n2093 GNDA.n551 175.546
R3324 GNDA.n2093 GNDA.n547 175.546
R3325 GNDA.n2097 GNDA.n547 175.546
R3326 GNDA.n1201 GNDA.n1084 175.546
R3327 GNDA.n1192 GNDA.n1092 175.546
R3328 GNDA.n1190 GNDA.n1093 175.546
R3329 GNDA.n1181 GNDA.n1101 175.546
R3330 GNDA.n1179 GNDA.n1102 175.546
R3331 GNDA.n2132 GNDA.n532 175.546
R3332 GNDA.n2136 GNDA.n532 175.546
R3333 GNDA.n2136 GNDA.n530 175.546
R3334 GNDA.n2141 GNDA.n530 175.546
R3335 GNDA.n2141 GNDA.n528 175.546
R3336 GNDA.n2145 GNDA.n528 175.546
R3337 GNDA.n2145 GNDA.n527 175.546
R3338 GNDA.n2149 GNDA.n527 175.546
R3339 GNDA.n2149 GNDA.n523 175.546
R3340 GNDA.n2154 GNDA.n523 175.546
R3341 GNDA.n2105 GNDA.n2102 175.546
R3342 GNDA.n2105 GNDA.n542 175.546
R3343 GNDA.n2109 GNDA.n542 175.546
R3344 GNDA.n2109 GNDA.n540 175.546
R3345 GNDA.n2113 GNDA.n540 175.546
R3346 GNDA.n2113 GNDA.n538 175.546
R3347 GNDA.n2117 GNDA.n538 175.546
R3348 GNDA.n2117 GNDA.n536 175.546
R3349 GNDA.n2122 GNDA.n536 175.546
R3350 GNDA.n2122 GNDA.n534 175.546
R3351 GNDA.n2126 GNDA.n534 175.546
R3352 GNDA.n1058 GNDA.n1057 175.546
R3353 GNDA.n1064 GNDA.n1063 175.546
R3354 GNDA.n1070 GNDA.n1069 175.546
R3355 GNDA.n1076 GNDA.n1075 175.546
R3356 GNDA.n1206 GNDA.n1205 175.546
R3357 GNDA.n1726 GNDA.n1725 164.369
R3358 GNDA.n1651 GNDA.n1650 164.369
R3359 GNDA.n1547 GNDA.n1403 163.333
R3360 GNDA.n1367 GNDA.n1366 163.333
R3361 GNDA.n2266 GNDA.n2265 163.333
R3362 GNDA.n852 GNDA.n851 163.333
R3363 GNDA.n1052 GNDA.n1051 163.333
R3364 GNDA.n1176 GNDA.n1175 163.333
R3365 GNDA.n1816 GNDA.n1751 163.333
R3366 GNDA.n2025 GNDA.n1962 163.333
R3367 GNDA.n2411 GNDA.n2410 163.333
R3368 GNDA.n1655 GNDA.t286 160.725
R3369 GNDA.n1656 GNDA.t282 160.725
R3370 GNDA.n1627 GNDA.t278 160.725
R3371 GNDA.n1625 GNDA.t256 160.725
R3372 GNDA.n1629 GNDA.t294 160.725
R3373 GNDA.n1714 GNDA.t309 160.725
R3374 GNDA.n559 GNDA.t89 157.555
R3375 GNDA.n558 GNDA.t4 157.555
R3376 GNDA.n437 GNDA.n436 156.8
R3377 GNDA.n487 GNDA.n330 153.601
R3378 GNDA.n2476 GNDA.n45 153.601
R3379 GNDA.n1659 GNDA.t8 153.294
R3380 GNDA.n327 GNDA.t253 152.994
R3381 GNDA.n323 GNDA.t246 152.994
R3382 GNDA.n51 GNDA.t243 152.994
R3383 GNDA.n46 GNDA.t224 152.994
R3384 GNDA.n2335 GNDA.n2334 152.643
R3385 GNDA.n1935 GNDA.n1934 152.643
R3386 GNDA.n102 GNDA.n94 150.988
R3387 GNDA.n491 GNDA.n322 150.4
R3388 GNDA.n2489 GNDA.n2488 150.4
R3389 GNDA.n73 GNDA.n72 150.4
R3390 GNDA.n1495 GNDA.n1418 150
R3391 GNDA.n1487 GNDA.n1486 150
R3392 GNDA.n1484 GNDA.n1463 150
R3393 GNDA.n1476 GNDA.n1475 150
R3394 GNDA.n1536 GNDA.n1535 150
R3395 GNDA.n1538 GNDA.n1536 150
R3396 GNDA.n1542 GNDA.n1405 150
R3397 GNDA.n1545 GNDA.n1544 150
R3398 GNDA.n1517 GNDA.n1412 150
R3399 GNDA.n1521 GNDA.n1519 150
R3400 GNDA.n1525 GNDA.n1410 150
R3401 GNDA.n1529 GNDA.n1527 150
R3402 GNDA.n1513 GNDA.n1511 150
R3403 GNDA.n1509 GNDA.n1414 150
R3404 GNDA.n1505 GNDA.n1503 150
R3405 GNDA.n1501 GNDA.n1416 150
R3406 GNDA.n1497 GNDA.n1416 150
R3407 GNDA.n1389 GNDA.n1388 150
R3408 GNDA.n1386 GNDA.n1280 150
R3409 GNDA.n1378 GNDA.n1377 150
R3410 GNDA.n1375 GNDA.n1289 150
R3411 GNDA.n1352 GNDA.n1304 150
R3412 GNDA.n1356 GNDA.n1304 150
R3413 GNDA.n1360 GNDA.n1358 150
R3414 GNDA.n1364 GNDA.n1302 150
R3415 GNDA.n1335 GNDA.n1333 150
R3416 GNDA.n1339 GNDA.n1309 150
R3417 GNDA.n1343 GNDA.n1341 150
R3418 GNDA.n1347 GNDA.n1307 150
R3419 GNDA.n1331 GNDA.n1311 150
R3420 GNDA.n1327 GNDA.n1325 150
R3421 GNDA.n1323 GNDA.n1313 150
R3422 GNDA.n1319 GNDA.n1317 150
R3423 GNDA.n1317 GNDA.n1316 150
R3424 GNDA.n2288 GNDA.n2287 150
R3425 GNDA.n2285 GNDA.n288 150
R3426 GNDA.n2277 GNDA.n2276 150
R3427 GNDA.n2274 GNDA.n297 150
R3428 GNDA.n2251 GNDA.n2203 150
R3429 GNDA.n2255 GNDA.n2203 150
R3430 GNDA.n2259 GNDA.n2257 150
R3431 GNDA.n2263 GNDA.n2201 150
R3432 GNDA.n2234 GNDA.n2232 150
R3433 GNDA.n2238 GNDA.n2208 150
R3434 GNDA.n2242 GNDA.n2240 150
R3435 GNDA.n2246 GNDA.n2206 150
R3436 GNDA.n2230 GNDA.n2210 150
R3437 GNDA.n2226 GNDA.n2224 150
R3438 GNDA.n2222 GNDA.n2212 150
R3439 GNDA.n2218 GNDA.n2216 150
R3440 GNDA.n2216 GNDA.n2215 150
R3441 GNDA.n874 GNDA.n873 150
R3442 GNDA.n871 GNDA.n760 150
R3443 GNDA.n863 GNDA.n862 150
R3444 GNDA.n860 GNDA.n769 150
R3445 GNDA.n837 GNDA.n789 150
R3446 GNDA.n841 GNDA.n789 150
R3447 GNDA.n845 GNDA.n843 150
R3448 GNDA.n849 GNDA.n787 150
R3449 GNDA.n820 GNDA.n818 150
R3450 GNDA.n824 GNDA.n794 150
R3451 GNDA.n828 GNDA.n826 150
R3452 GNDA.n832 GNDA.n792 150
R3453 GNDA.n816 GNDA.n796 150
R3454 GNDA.n812 GNDA.n810 150
R3455 GNDA.n808 GNDA.n798 150
R3456 GNDA.n804 GNDA.n802 150
R3457 GNDA.n802 GNDA.n801 150
R3458 GNDA.n999 GNDA.n717 150
R3459 GNDA.n988 GNDA.n970 150
R3460 GNDA.n986 GNDA.n971 150
R3461 GNDA.n975 GNDA.n974 150
R3462 GNDA.n1037 GNDA.n705 150
R3463 GNDA.n1041 GNDA.n705 150
R3464 GNDA.n1045 GNDA.n1043 150
R3465 GNDA.n1049 GNDA.n703 150
R3466 GNDA.n1020 GNDA.n1018 150
R3467 GNDA.n1024 GNDA.n710 150
R3468 GNDA.n1028 GNDA.n1026 150
R3469 GNDA.n1032 GNDA.n708 150
R3470 GNDA.n1016 GNDA.n712 150
R3471 GNDA.n1012 GNDA.n1010 150
R3472 GNDA.n1008 GNDA.n714 150
R3473 GNDA.n1004 GNDA.n1002 150
R3474 GNDA.n1002 GNDA.n1001 150
R3475 GNDA.n1198 GNDA.n1197 150
R3476 GNDA.n1195 GNDA.n1088 150
R3477 GNDA.n1187 GNDA.n1186 150
R3478 GNDA.n1184 GNDA.n1097 150
R3479 GNDA.n1161 GNDA.n1113 150
R3480 GNDA.n1165 GNDA.n1113 150
R3481 GNDA.n1169 GNDA.n1167 150
R3482 GNDA.n1173 GNDA.n1111 150
R3483 GNDA.n1144 GNDA.n1142 150
R3484 GNDA.n1148 GNDA.n1118 150
R3485 GNDA.n1152 GNDA.n1150 150
R3486 GNDA.n1156 GNDA.n1116 150
R3487 GNDA.n1140 GNDA.n1120 150
R3488 GNDA.n1136 GNDA.n1134 150
R3489 GNDA.n1132 GNDA.n1122 150
R3490 GNDA.n1128 GNDA.n1126 150
R3491 GNDA.n1126 GNDA.n1125 150
R3492 GNDA.n1847 GNDA.n617 150
R3493 GNDA.n1845 GNDA.n618 150
R3494 GNDA.n1835 GNDA.n1611 150
R3495 GNDA.n1833 GNDA.n1612 150
R3496 GNDA.n1805 GNDA.n1804 150
R3497 GNDA.n1807 GNDA.n1805 150
R3498 GNDA.n1811 GNDA.n1753 150
R3499 GNDA.n1814 GNDA.n1813 150
R3500 GNDA.n1786 GNDA.n1760 150
R3501 GNDA.n1790 GNDA.n1788 150
R3502 GNDA.n1794 GNDA.n1758 150
R3503 GNDA.n1798 GNDA.n1796 150
R3504 GNDA.n1782 GNDA.n1780 150
R3505 GNDA.n1778 GNDA.n1762 150
R3506 GNDA.n1774 GNDA.n1772 150
R3507 GNDA.n1770 GNDA.n1764 150
R3508 GNDA.n1766 GNDA.n1764 150
R3509 GNDA.n2060 GNDA.n2059 150
R3510 GNDA.n2057 GNDA.n1941 150
R3511 GNDA.n2045 GNDA.n2044 150
R3512 GNDA.n2042 GNDA.n1949 150
R3513 GNDA.n2014 GNDA.n2013 150
R3514 GNDA.n2016 GNDA.n2014 150
R3515 GNDA.n2020 GNDA.n1964 150
R3516 GNDA.n2023 GNDA.n2022 150
R3517 GNDA.n1995 GNDA.n1971 150
R3518 GNDA.n1999 GNDA.n1997 150
R3519 GNDA.n2003 GNDA.n1969 150
R3520 GNDA.n2007 GNDA.n2005 150
R3521 GNDA.n1991 GNDA.n1989 150
R3522 GNDA.n1987 GNDA.n1973 150
R3523 GNDA.n1983 GNDA.n1981 150
R3524 GNDA.n1979 GNDA.n1976 150
R3525 GNDA.n1976 GNDA.n1975 150
R3526 GNDA.n2358 GNDA.n140 150
R3527 GNDA.n2348 GNDA.n2346 150
R3528 GNDA.n2422 GNDA.n125 150
R3529 GNDA.n2420 GNDA.n2413 150
R3530 GNDA.n2396 GNDA.n128 150
R3531 GNDA.n2400 GNDA.n128 150
R3532 GNDA.n2404 GNDA.n2402 150
R3533 GNDA.n2408 GNDA.n126 150
R3534 GNDA.n2379 GNDA.n2377 150
R3535 GNDA.n2383 GNDA.n133 150
R3536 GNDA.n2387 GNDA.n2385 150
R3537 GNDA.n2391 GNDA.n131 150
R3538 GNDA.n2375 GNDA.n135 150
R3539 GNDA.n2371 GNDA.n2369 150
R3540 GNDA.n2367 GNDA.n137 150
R3541 GNDA.n2363 GNDA.n2361 150
R3542 GNDA.n2361 GNDA.n2360 150
R3543 GNDA.n556 GNDA.t90 148.906
R3544 GNDA.n556 GNDA.t24 148.653
R3545 GNDA.n482 GNDA.t299 147.511
R3546 GNDA.n476 GNDA.t315 147.511
R3547 GNDA.t293 GNDA.t22 145.403
R3548 GNDA.t320 GNDA.t281 145.403
R3549 GNDA.n94 GNDA.n86 145.013
R3550 GNDA.n1662 GNDA.n1660 139.638
R3551 GNDA.t255 GNDA.t43 139.081
R3552 GNDA.t43 GNDA.t33 139.081
R3553 GNDA.t33 GNDA.t163 139.081
R3554 GNDA.t123 GNDA.t107 139.081
R3555 GNDA.t54 GNDA.t123 139.081
R3556 GNDA.t277 GNDA.t54 139.081
R3557 GNDA.n1678 GNDA.n1677 139.077
R3558 GNDA.n1676 GNDA.n1675 139.077
R3559 GNDA.n1674 GNDA.n1673 139.077
R3560 GNDA.n1672 GNDA.n1671 139.077
R3561 GNDA.n1670 GNDA.n1669 139.077
R3562 GNDA.n1668 GNDA.n1667 139.077
R3563 GNDA.n1666 GNDA.n1665 139.077
R3564 GNDA.n1664 GNDA.n1663 139.077
R3565 GNDA.n1662 GNDA.n1661 139.077
R3566 GNDA.t339 GNDA.t274 135.386
R3567 GNDA.t330 GNDA.t215 135.386
R3568 GNDA.t239 GNDA.t205 135.386
R3569 GNDA.t290 GNDA.t207 135.386
R3570 GNDA.t197 GNDA.t25 135.386
R3571 GNDA.t5 GNDA.t271 135.386
R3572 GNDA.n370 GNDA.n369 134.867
R3573 GNDA.n2472 GNDA.n55 134.867
R3574 GNDA.n478 GNDA.n473 134.4
R3575 GNDA.n467 GNDA.n359 134.4
R3576 GNDA.n466 GNDA.n464 134.4
R3577 GNDA.n365 GNDA.n364 134.4
R3578 GNDA.n363 GNDA.n357 134.4
R3579 GNDA.n1737 GNDA.t163 132.76
R3580 GNDA.t107 GNDA.n1649 132.76
R3581 GNDA.n480 GNDA.n339 128
R3582 GNDA.n1718 GNDA.t15 126.438
R3583 GNDA.n1685 GNDA.t193 126.438
R3584 GNDA.n2197 GNDA.n2196 124.832
R3585 GNDA.n2331 GNDA.n2330 124.832
R3586 GNDA.n2443 GNDA.n88 124.832
R3587 GNDA.n234 GNDA.n232 124.832
R3588 GNDA.n2030 GNDA.n1957 124.832
R3589 GNDA.n1252 GNDA.n1251 124.832
R3590 GNDA.n1298 GNDA.n207 124.832
R3591 GNDA.n667 GNDA.n185 124.832
R3592 GNDA.n1821 GNDA.n1746 124.832
R3593 GNDA.n1903 GNDA.n1902 124.832
R3594 GNDA.n1554 GNDA.n1553 124.832
R3595 GNDA.n1580 GNDA.n1579 124.832
R3596 GNDA.n783 GNDA.n782 124.832
R3597 GNDA.n928 GNDA.n927 124.832
R3598 GNDA.n1212 GNDA.n698 124.832
R3599 GNDA.n2098 GNDA.n2097 124.832
R3600 GNDA.n1107 GNDA.n1105 124.832
R3601 GNDA.n2127 GNDA.n2126 124.832
R3602 GNDA.t56 GNDA.t183 120.115
R3603 GNDA.t173 GNDA.t37 120.115
R3604 GNDA.n2067 GNDA.n568 119.035
R3605 GNDA.n546 GNDA.n145 119.035
R3606 GNDA.n1657 GNDA.n1628 118.4
R3607 GNDA.n1683 GNDA.n1658 118.4
R3608 GNDA.n1730 GNDA.n1626 118.4
R3609 GNDA.n1733 GNDA.n1732 118.4
R3610 GNDA.n1716 GNDA.n1715 118.4
R3611 GNDA.n1729 GNDA.n1630 118.4
R3612 GNDA.n343 GNDA.t250 113.974
R3613 GNDA.n344 GNDA.t234 113.974
R3614 GNDA.n338 GNDA.t300 113.974
R3615 GNDA.n340 GNDA.t316 113.974
R3616 GNDA.n341 GNDA.t297 113.974
R3617 GNDA.n342 GNDA.t288 113.974
R3618 GNDA.n463 GNDA.t303 113.974
R3619 GNDA.n358 GNDA.t291 113.974
R3620 GNDA.n362 GNDA.t240 113.974
R3621 GNDA.n361 GNDA.t306 113.974
R3622 GNDA.t229 GNDA.n1839 113.624
R3623 GNDA.n1745 GNDA.n1744 113.624
R3624 GNDA.n1954 GNDA.t231 113.624
R3625 GNDA.t248 GNDA.n2426 113.624
R3626 GNDA.n457 GNDA.n456 108.8
R3627 GNDA.n454 GNDA.n452 108.8
R3628 GNDA.n2067 GNDA.n569 103.144
R3629 GNDA.n2302 GNDA.n145 103.144
R3630 GNDA.n1719 GNDA.n1718 101.15
R3631 GNDA.t161 GNDA.t162 101.15
R3632 GNDA.t318 GNDA.t7 101.15
R3633 GNDA.n1698 GNDA.n1685 101.15
R3634 GNDA.n2067 GNDA.n570 99.6276
R3635 GNDA.n2333 GNDA.n145 99.6276
R3636 GNDA.n432 GNDA.n431 99.0842
R3637 GNDA.n430 GNDA.n429 99.0842
R3638 GNDA.n428 GNDA.n427 99.0842
R3639 GNDA.n426 GNDA.n425 99.0842
R3640 GNDA.n424 GNDA.n423 99.0842
R3641 GNDA.n422 GNDA.n421 99.0842
R3642 GNDA.n420 GNDA.n419 99.0842
R3643 GNDA.n418 GNDA.n417 99.0842
R3644 GNDA.n416 GNDA.n415 99.0842
R3645 GNDA.n414 GNDA.n413 99.0842
R3646 GNDA.n36 GNDA.n35 99.0842
R3647 GNDA.n2450 GNDA.n82 98.4712
R3648 GNDA.n907 GNDA.n740 96.5152
R3649 GNDA.n908 GNDA.n907 96.5152
R3650 GNDA.n910 GNDA.n908 96.5152
R3651 GNDA.n910 GNDA.n909 96.5152
R3652 GNDA.n909 GNDA.n621 96.5152
R3653 GNDA.n917 GNDA.n622 96.5152
R3654 GNDA.n917 GNDA.n734 96.5152
R3655 GNDA.n924 GNDA.n734 96.5152
R3656 GNDA.n925 GNDA.n924 96.5152
R3657 GNDA.n926 GNDA.n925 96.5152
R3658 GNDA.n926 GNDA.n568 96.5152
R3659 GNDA.n2069 GNDA.n2068 96.5152
R3660 GNDA.n2069 GNDA.n564 96.5152
R3661 GNDA.n2075 GNDA.n564 96.5152
R3662 GNDA.n2076 GNDA.n2075 96.5152
R3663 GNDA.n2077 GNDA.n2076 96.5152
R3664 GNDA.n2087 GNDA.n2086 96.5152
R3665 GNDA.n2087 GNDA.n550 96.5152
R3666 GNDA.n2094 GNDA.n550 96.5152
R3667 GNDA.n2095 GNDA.n2094 96.5152
R3668 GNDA.n2096 GNDA.n2095 96.5152
R3669 GNDA.n2096 GNDA.n546 96.5152
R3670 GNDA.n2104 GNDA.n2103 96.5152
R3671 GNDA.n2104 GNDA.n541 96.5152
R3672 GNDA.n2110 GNDA.n541 96.5152
R3673 GNDA.n2111 GNDA.n2110 96.5152
R3674 GNDA.n2112 GNDA.n2111 96.5152
R3675 GNDA.n2118 GNDA.n537 96.5152
R3676 GNDA.n2119 GNDA.n2118 96.5152
R3677 GNDA.n2121 GNDA.n2119 96.5152
R3678 GNDA.n2121 GNDA.n2120 96.5152
R3679 GNDA.n2120 GNDA.n317 96.5152
R3680 GNDA.n2182 GNDA.n496 95.7359
R3681 GNDA.n2450 GNDA.n85 95.4038
R3682 GNDA.n2482 GNDA.n37 95.101
R3683 GNDA.n377 GNDA.n374 95.101
R3684 GNDA.n2487 GNDA.t266 94.8842
R3685 GNDA.n434 GNDA.t237 94.8842
R3686 GNDA.t15 GNDA.t308 94.8281
R3687 GNDA.t169 GNDA.t99 94.8281
R3688 GNDA.t35 GNDA.t0 94.8281
R3689 GNDA.t193 GNDA.t285 94.8281
R3690 GNDA.n2484 GNDA.n2483 94.601
R3691 GNDA.n376 GNDA.n375 94.601
R3692 GNDA.t245 GNDA.t128 92.7208
R3693 GNDA.t30 GNDA.t116 92.7208
R3694 GNDA.t105 GNDA.t16 92.7208
R3695 GNDA.t86 GNDA.t136 92.7208
R3696 GNDA.t217 GNDA.t71 92.7208
R3697 GNDA.t71 GNDA.t87 92.7208
R3698 GNDA.t31 GNDA.t159 92.7208
R3699 GNDA.t9 GNDA.t31 92.7208
R3700 GNDA.t14 GNDA.t132 92.7208
R3701 GNDA.t103 GNDA.t101 92.7208
R3702 GNDA.t134 GNDA.t146 92.7208
R3703 GNDA.t242 GNDA.t106 92.7208
R3704 GNDA.t231 GNDA.n570 91.423
R3705 GNDA.n2333 GNDA.t248 91.423
R3706 GNDA.t80 GNDA.t311 88.5063
R3707 GNDA.t268 GNDA.t135 88.5063
R3708 GNDA.n1706 GNDA.n1705 85.2845
R3709 GNDA.n1639 GNDA.n1638 85.2845
R3710 GNDA.n555 GNDA.n554 84.306
R3711 GNDA.t186 GNDA.t58 82.1844
R3712 GNDA.t119 GNDA.t61 82.1844
R3713 GNDA.t165 GNDA.t319 82.1844
R3714 GNDA.t182 GNDA.t175 82.1844
R3715 GNDA.t128 GNDA.t226 80.0771
R3716 GNDA.t28 GNDA.t80 80.0771
R3717 GNDA.t135 GNDA.t321 80.0771
R3718 GNDA.t106 GNDA.t258 80.0771
R3719 GNDA.n2292 GNDA.n2291 76.3222
R3720 GNDA.n292 GNDA.n291 76.3222
R3721 GNDA.n2281 GNDA.n2280 76.3222
R3722 GNDA.n301 GNDA.n300 76.3222
R3723 GNDA.n2270 GNDA.n2269 76.3222
R3724 GNDA.n2197 GNDA.n306 76.3222
R3725 GNDA.n2192 GNDA.n307 76.3222
R3726 GNDA.n2308 GNDA.n2307 76.3222
R3727 GNDA.n2313 GNDA.n2312 76.3222
R3728 GNDA.n2316 GNDA.n2315 76.3222
R3729 GNDA.n2321 GNDA.n2320 76.3222
R3730 GNDA.n2324 GNDA.n2323 76.3222
R3731 GNDA.n2329 GNDA.n2328 76.3222
R3732 GNDA.n2306 GNDA.n150 76.3222
R3733 GNDA.n259 GNDA.n151 76.3222
R3734 GNDA.n264 GNDA.n152 76.3222
R3735 GNDA.n270 GNDA.n153 76.3222
R3736 GNDA.n2295 GNDA.n154 76.3222
R3737 GNDA.n2296 GNDA.n149 76.3222
R3738 GNDA.n112 GNDA.n110 76.3222
R3739 GNDA.n255 GNDA.n254 76.3222
R3740 GNDA.n252 GNDA.n210 76.3222
R3741 GNDA.n248 GNDA.n247 76.3222
R3742 GNDA.n241 GNDA.n212 76.3222
R3743 GNDA.n240 GNDA.n239 76.3222
R3744 GNDA.n233 GNDA.n214 76.3222
R3745 GNDA.n1224 GNDA.n162 76.3222
R3746 GNDA.n1226 GNDA.n163 76.3222
R3747 GNDA.n1228 GNDA.n164 76.3222
R3748 GNDA.n1230 GNDA.n165 76.3222
R3749 GNDA.n2335 GNDA.n146 76.3222
R3750 GNDA.n1250 GNDA.n204 76.3222
R3751 GNDA.n1246 GNDA.n203 76.3222
R3752 GNDA.n1242 GNDA.n202 76.3222
R3753 GNDA.n1238 GNDA.n201 76.3222
R3754 GNDA.n1234 GNDA.n200 76.3222
R3755 GNDA.n2027 GNDA.n199 76.3222
R3756 GNDA.n1273 GNDA.n586 76.3222
R3757 GNDA.n1220 GNDA.n1219 76.3222
R3758 GNDA.n1267 GNDA.n1218 76.3222
R3759 GNDA.n1263 GNDA.n1217 76.3222
R3760 GNDA.n1259 GNDA.n1216 76.3222
R3761 GNDA.n1255 GNDA.n1215 76.3222
R3762 GNDA.n1911 GNDA.n1909 76.3222
R3763 GNDA.n1919 GNDA.n582 76.3222
R3764 GNDA.n1924 GNDA.n1921 76.3222
R3765 GNDA.n1922 GNDA.n576 76.3222
R3766 GNDA.n1935 GNDA.n573 76.3222
R3767 GNDA.n1393 GNDA.n1392 76.3222
R3768 GNDA.n1284 GNDA.n1283 76.3222
R3769 GNDA.n1382 GNDA.n1381 76.3222
R3770 GNDA.n1293 GNDA.n1292 76.3222
R3771 GNDA.n1371 GNDA.n1370 76.3222
R3772 GNDA.n1298 GNDA.n1297 76.3222
R3773 GNDA.n2304 GNDA.n2303 76.3222
R3774 GNDA.n260 GNDA.n192 76.3222
R3775 GNDA.n266 GNDA.n191 76.3222
R3776 GNDA.n272 GNDA.n190 76.3222
R3777 GNDA.n278 GNDA.n189 76.3222
R3778 GNDA.n2300 GNDA.n188 76.3222
R3779 GNDA.n690 GNDA.n689 76.3222
R3780 GNDA.n685 GNDA.n665 76.3222
R3781 GNDA.n682 GNDA.n664 76.3222
R3782 GNDA.n678 GNDA.n663 76.3222
R3783 GNDA.n674 GNDA.n662 76.3222
R3784 GNDA.n670 GNDA.n661 76.3222
R3785 GNDA.n639 GNDA.n638 76.3222
R3786 GNDA.n644 GNDA.n643 76.3222
R3787 GNDA.n647 GNDA.n646 76.3222
R3788 GNDA.n652 GNDA.n651 76.3222
R3789 GNDA.n655 GNDA.n654 76.3222
R3790 GNDA.n660 GNDA.n658 76.3222
R3791 GNDA.n1905 GNDA.n1904 76.3222
R3792 GNDA.n1914 GNDA.n1913 76.3222
R3793 GNDA.n1917 GNDA.n1916 76.3222
R3794 GNDA.n1927 GNDA.n1926 76.3222
R3795 GNDA.n1930 GNDA.n1929 76.3222
R3796 GNDA.n1819 GNDA.n578 76.3222
R3797 GNDA.n1880 GNDA.n1879 76.3222
R3798 GNDA.n1885 GNDA.n1884 76.3222
R3799 GNDA.n1888 GNDA.n1887 76.3222
R3800 GNDA.n1893 GNDA.n1892 76.3222
R3801 GNDA.n1896 GNDA.n1895 76.3222
R3802 GNDA.n1901 GNDA.n1900 76.3222
R3803 GNDA.n1858 GNDA.n1857 76.3222
R3804 GNDA.n1458 GNDA.n1457 76.3222
R3805 GNDA.n1491 GNDA.n1490 76.3222
R3806 GNDA.n1467 GNDA.n1466 76.3222
R3807 GNDA.n1480 GNDA.n1479 76.3222
R3808 GNDA.n1468 GNDA.n1400 76.3222
R3809 GNDA.n1553 GNDA.n1552 76.3222
R3810 GNDA.n1578 GNDA.n636 76.3222
R3811 GNDA.n1574 GNDA.n1573 76.3222
R3812 GNDA.n1567 GNDA.n641 76.3222
R3813 GNDA.n1566 GNDA.n1565 76.3222
R3814 GNDA.n1559 GNDA.n649 76.3222
R3815 GNDA.n1558 GNDA.n1557 76.3222
R3816 GNDA.n1603 GNDA.n1602 76.3222
R3817 GNDA.n1598 GNDA.n630 76.3222
R3818 GNDA.n1595 GNDA.n629 76.3222
R3819 GNDA.n1591 GNDA.n628 76.3222
R3820 GNDA.n1587 GNDA.n627 76.3222
R3821 GNDA.n1583 GNDA.n626 76.3222
R3822 GNDA.n1453 GNDA.n1421 76.3222
R3823 GNDA.n878 GNDA.n877 76.3222
R3824 GNDA.n764 GNDA.n763 76.3222
R3825 GNDA.n867 GNDA.n866 76.3222
R3826 GNDA.n773 GNDA.n772 76.3222
R3827 GNDA.n856 GNDA.n855 76.3222
R3828 GNDA.n783 GNDA.n778 76.3222
R3829 GNDA.n881 GNDA.n880 76.3222
R3830 GNDA.n930 GNDA.n929 76.3222
R3831 GNDA.n939 GNDA.n938 76.3222
R3832 GNDA.n942 GNDA.n941 76.3222
R3833 GNDA.n953 GNDA.n952 76.3222
R3834 GNDA.n956 GNDA.n955 76.3222
R3835 GNDA.n780 GNDA.n722 76.3222
R3836 GNDA.n995 GNDA.n692 76.3222
R3837 GNDA.n992 GNDA.n693 76.3222
R3838 GNDA.n982 GNDA.n694 76.3222
R3839 GNDA.n979 GNDA.n695 76.3222
R3840 GNDA.n700 GNDA.n696 76.3222
R3841 GNDA.n1213 GNDA.n1212 76.3222
R3842 GNDA.n934 GNDA.n933 76.3222
R3843 GNDA.n935 GNDA.n726 76.3222
R3844 GNDA.n946 GNDA.n945 76.3222
R3845 GNDA.n949 GNDA.n948 76.3222
R3846 GNDA.n959 GNDA.n719 76.3222
R3847 GNDA.n962 GNDA.n961 76.3222
R3848 GNDA.n2099 GNDA.n198 76.3222
R3849 GNDA.n1060 GNDA.n197 76.3222
R3850 GNDA.n1066 GNDA.n196 76.3222
R3851 GNDA.n1072 GNDA.n195 76.3222
R3852 GNDA.n1078 GNDA.n194 76.3222
R3853 GNDA.n1056 GNDA.n193 76.3222
R3854 GNDA.n1857 GNDA.n609 76.3222
R3855 GNDA.n1879 GNDA.n595 76.3222
R3856 GNDA.n1886 GNDA.n1885 76.3222
R3857 GNDA.n1887 GNDA.n593 76.3222
R3858 GNDA.n1894 GNDA.n1893 76.3222
R3859 GNDA.n1895 GNDA.n591 76.3222
R3860 GNDA.n1902 GNDA.n1901 76.3222
R3861 GNDA.n1603 GNDA.n631 76.3222
R3862 GNDA.n1596 GNDA.n630 76.3222
R3863 GNDA.n1592 GNDA.n629 76.3222
R3864 GNDA.n1588 GNDA.n628 76.3222
R3865 GNDA.n1584 GNDA.n627 76.3222
R3866 GNDA.n1580 GNDA.n626 76.3222
R3867 GNDA.n947 GNDA.n719 76.3222
R3868 GNDA.n950 GNDA.n949 76.3222
R3869 GNDA.n945 GNDA.n944 76.3222
R3870 GNDA.n936 GNDA.n935 76.3222
R3871 GNDA.n933 GNDA.n932 76.3222
R3872 GNDA.n654 GNDA.n653 76.3222
R3873 GNDA.n651 GNDA.n650 76.3222
R3874 GNDA.n646 GNDA.n645 76.3222
R3875 GNDA.n643 GNDA.n642 76.3222
R3876 GNDA.n638 GNDA.n637 76.3222
R3877 GNDA.n1934 GNDA.n1933 76.3222
R3878 GNDA.n1923 GNDA.n1922 76.3222
R3879 GNDA.n1921 GNDA.n1920 76.3222
R3880 GNDA.n1910 GNDA.n582 76.3222
R3881 GNDA.n1909 GNDA.n1908 76.3222
R3882 GNDA.n929 GNDA.n728 76.3222
R3883 GNDA.n940 GNDA.n939 76.3222
R3884 GNDA.n941 GNDA.n724 76.3222
R3885 GNDA.n954 GNDA.n953 76.3222
R3886 GNDA.n957 GNDA.n956 76.3222
R3887 GNDA.n1575 GNDA.n636 76.3222
R3888 GNDA.n1573 GNDA.n1572 76.3222
R3889 GNDA.n1568 GNDA.n1567 76.3222
R3890 GNDA.n1565 GNDA.n1564 76.3222
R3891 GNDA.n1560 GNDA.n1559 76.3222
R3892 GNDA.n1904 GNDA.n584 76.3222
R3893 GNDA.n1915 GNDA.n1914 76.3222
R3894 GNDA.n1916 GNDA.n580 76.3222
R3895 GNDA.n1928 GNDA.n1927 76.3222
R3896 GNDA.n1931 GNDA.n1930 76.3222
R3897 GNDA.n1820 GNDA.n1819 76.3222
R3898 GNDA.n1273 GNDA.n1272 76.3222
R3899 GNDA.n1268 GNDA.n1219 76.3222
R3900 GNDA.n1264 GNDA.n1218 76.3222
R3901 GNDA.n1260 GNDA.n1217 76.3222
R3902 GNDA.n1256 GNDA.n1216 76.3222
R3903 GNDA.n1252 GNDA.n1215 76.3222
R3904 GNDA.n690 GNDA.n666 76.3222
R3905 GNDA.n683 GNDA.n665 76.3222
R3906 GNDA.n679 GNDA.n664 76.3222
R3907 GNDA.n675 GNDA.n663 76.3222
R3908 GNDA.n671 GNDA.n662 76.3222
R3909 GNDA.n667 GNDA.n661 76.3222
R3910 GNDA.n2334 GNDA.n148 76.3222
R3911 GNDA.n1229 GNDA.n165 76.3222
R3912 GNDA.n1227 GNDA.n164 76.3222
R3913 GNDA.n1225 GNDA.n163 76.3222
R3914 GNDA.n1223 GNDA.n162 76.3222
R3915 GNDA.n1247 GNDA.n204 76.3222
R3916 GNDA.n1243 GNDA.n203 76.3222
R3917 GNDA.n1239 GNDA.n202 76.3222
R3918 GNDA.n1235 GNDA.n201 76.3222
R3919 GNDA.n1231 GNDA.n200 76.3222
R3920 GNDA.n2027 GNDA.n205 76.3222
R3921 GNDA.n1203 GNDA.n1202 76.3222
R3922 GNDA.n1091 GNDA.n1084 76.3222
R3923 GNDA.n1192 GNDA.n1191 76.3222
R3924 GNDA.n1100 GNDA.n1093 76.3222
R3925 GNDA.n1181 GNDA.n1180 76.3222
R3926 GNDA.n1106 GNDA.n1102 76.3222
R3927 GNDA.n2154 GNDA.n2153 76.3222
R3928 GNDA.n2101 GNDA.n156 76.3222
R3929 GNDA.n1058 GNDA.n157 76.3222
R3930 GNDA.n1064 GNDA.n158 76.3222
R3931 GNDA.n1070 GNDA.n159 76.3222
R3932 GNDA.n1076 GNDA.n160 76.3222
R3933 GNDA.n1206 GNDA.n155 76.3222
R3934 GNDA.n1205 GNDA.n160 76.3222
R3935 GNDA.n1075 GNDA.n159 76.3222
R3936 GNDA.n1069 GNDA.n158 76.3222
R3937 GNDA.n1063 GNDA.n157 76.3222
R3938 GNDA.n1057 GNDA.n156 76.3222
R3939 GNDA.n1059 GNDA.n198 76.3222
R3940 GNDA.n1065 GNDA.n197 76.3222
R3941 GNDA.n1071 GNDA.n196 76.3222
R3942 GNDA.n1077 GNDA.n195 76.3222
R3943 GNDA.n1080 GNDA.n194 76.3222
R3944 GNDA.n1082 GNDA.n155 76.3222
R3945 GNDA.n1107 GNDA.n1106 76.3222
R3946 GNDA.n1180 GNDA.n1179 76.3222
R3947 GNDA.n1101 GNDA.n1100 76.3222
R3948 GNDA.n1191 GNDA.n1190 76.3222
R3949 GNDA.n1092 GNDA.n1091 76.3222
R3950 GNDA.n1202 GNDA.n1201 76.3222
R3951 GNDA.n961 GNDA.n960 76.3222
R3952 GNDA.n1213 GNDA.n697 76.3222
R3953 GNDA.n978 GNDA.n696 76.3222
R3954 GNDA.n983 GNDA.n695 76.3222
R3955 GNDA.n991 GNDA.n694 76.3222
R3956 GNDA.n996 GNDA.n693 76.3222
R3957 GNDA.n963 GNDA.n692 76.3222
R3958 GNDA.n1056 GNDA.n206 76.3222
R3959 GNDA.n882 GNDA.n881 76.3222
R3960 GNDA.n778 GNDA.n774 76.3222
R3961 GNDA.n857 GNDA.n856 76.3222
R3962 GNDA.n772 GNDA.n765 76.3222
R3963 GNDA.n868 GNDA.n867 76.3222
R3964 GNDA.n763 GNDA.n755 76.3222
R3965 GNDA.n879 GNDA.n878 76.3222
R3966 GNDA.n781 GNDA.n780 76.3222
R3967 GNDA.n276 GNDA.n154 76.3222
R3968 GNDA.n275 GNDA.n153 76.3222
R3969 GNDA.n269 GNDA.n152 76.3222
R3970 GNDA.n263 GNDA.n151 76.3222
R3971 GNDA.n258 GNDA.n150 76.3222
R3972 GNDA.n2303 GNDA.n186 76.3222
R3973 GNDA.n265 GNDA.n192 76.3222
R3974 GNDA.n271 GNDA.n191 76.3222
R3975 GNDA.n277 GNDA.n190 76.3222
R3976 GNDA.n280 GNDA.n189 76.3222
R3977 GNDA.n2307 GNDA.n181 76.3222
R3978 GNDA.n2314 GNDA.n2313 76.3222
R3979 GNDA.n2315 GNDA.n179 76.3222
R3980 GNDA.n2322 GNDA.n2321 76.3222
R3981 GNDA.n2323 GNDA.n177 76.3222
R3982 GNDA.n2330 GNDA.n2329 76.3222
R3983 GNDA.n282 GNDA.n149 76.3222
R3984 GNDA.n658 GNDA.n657 76.3222
R3985 GNDA.n1297 GNDA.n1294 76.3222
R3986 GNDA.n1372 GNDA.n1371 76.3222
R3987 GNDA.n1292 GNDA.n1285 76.3222
R3988 GNDA.n1383 GNDA.n1382 76.3222
R3989 GNDA.n1283 GNDA.n1276 76.3222
R3990 GNDA.n1394 GNDA.n1393 76.3222
R3991 GNDA.n2301 GNDA.n2300 76.3222
R3992 GNDA.n1453 GNDA.n1452 76.3222
R3993 GNDA.n1552 GNDA.n1551 76.3222
R3994 GNDA.n1469 GNDA.n1468 76.3222
R3995 GNDA.n1481 GNDA.n1480 76.3222
R3996 GNDA.n1466 GNDA.n1459 76.3222
R3997 GNDA.n1492 GNDA.n1491 76.3222
R3998 GNDA.n1457 GNDA.n1456 76.3222
R3999 GNDA.n1557 GNDA.n1398 76.3222
R4000 GNDA.n306 GNDA.n302 76.3222
R4001 GNDA.n2271 GNDA.n2270 76.3222
R4002 GNDA.n300 GNDA.n293 76.3222
R4003 GNDA.n2282 GNDA.n2281 76.3222
R4004 GNDA.n291 GNDA.n284 76.3222
R4005 GNDA.n2293 GNDA.n2292 76.3222
R4006 GNDA.n254 GNDA.n253 76.3222
R4007 GNDA.n249 GNDA.n210 76.3222
R4008 GNDA.n247 GNDA.n246 76.3222
R4009 GNDA.n242 GNDA.n241 76.3222
R4010 GNDA.n239 GNDA.n238 76.3222
R4011 GNDA.n234 GNDA.n233 76.3222
R4012 GNDA.n2153 GNDA.n524 76.3222
R4013 GNDA.n2195 GNDA.n307 76.3222
R4014 GNDA.n110 GNDA.n92 76.3222
R4015 GNDA.n1512 GNDA.n1412 76.062
R4016 GNDA.n1513 GNDA.n1512 76.062
R4017 GNDA.n1333 GNDA.n1332 76.062
R4018 GNDA.n1332 GNDA.n1331 76.062
R4019 GNDA.n2232 GNDA.n2231 76.062
R4020 GNDA.n2231 GNDA.n2230 76.062
R4021 GNDA.n818 GNDA.n817 76.062
R4022 GNDA.n817 GNDA.n816 76.062
R4023 GNDA.n1018 GNDA.n1017 76.062
R4024 GNDA.n1017 GNDA.n1016 76.062
R4025 GNDA.n1142 GNDA.n1141 76.062
R4026 GNDA.n1141 GNDA.n1140 76.062
R4027 GNDA.n1781 GNDA.n1760 76.062
R4028 GNDA.n1782 GNDA.n1781 76.062
R4029 GNDA.n1990 GNDA.n1971 76.062
R4030 GNDA.n1991 GNDA.n1990 76.062
R4031 GNDA.n2377 GNDA.n2376 76.062
R4032 GNDA.n2376 GNDA.n2375 76.062
R4033 GNDA.t305 GNDA.t299 75.8626
R4034 GNDA.t126 GNDA.t27 75.8626
R4035 GNDA.t315 GNDA.t302 75.8626
R4036 GNDA.n1711 GNDA.t187 75.8626
R4037 GNDA.n1727 GNDA.t22 75.8626
R4038 GNDA.n1727 GNDA.t185 75.8626
R4039 GNDA.n1652 GNDA.t172 75.8626
R4040 GNDA.n1652 GNDA.t320 75.8626
R4041 GNDA.n1702 GNDA.t171 75.8626
R4042 GNDA.n1496 GNDA.n1495 74.5978
R4043 GNDA.n1497 GNDA.n1496 74.5978
R4044 GNDA.n1389 GNDA.n1278 74.5978
R4045 GNDA.n1316 GNDA.n1278 74.5978
R4046 GNDA.n2288 GNDA.n286 74.5978
R4047 GNDA.n2215 GNDA.n286 74.5978
R4048 GNDA.n874 GNDA.n758 74.5978
R4049 GNDA.n801 GNDA.n758 74.5978
R4050 GNDA.n1000 GNDA.n999 74.5978
R4051 GNDA.n1001 GNDA.n1000 74.5978
R4052 GNDA.n1198 GNDA.n1086 74.5978
R4053 GNDA.n1125 GNDA.n1086 74.5978
R4054 GNDA.n1765 GNDA.n617 74.5978
R4055 GNDA.n1766 GNDA.n1765 74.5978
R4056 GNDA.n2060 GNDA.n1939 74.5978
R4057 GNDA.n1975 GNDA.n1939 74.5978
R4058 GNDA.n2359 GNDA.n2358 74.5978
R4059 GNDA.n2360 GNDA.n2359 74.5978
R4060 GNDA.n2441 GNDA.n94 73.3065
R4061 GNDA.n2471 GNDA.t337 72.3996
R4062 GNDA.n2457 GNDA.t114 72.3996
R4063 GNDA.n495 GNDA.t143 72.3996
R4064 GNDA.n403 GNDA.t6 72.3996
R4065 GNDA.t73 GNDA.n439 71.648
R4066 GNDA.n2465 GNDA.n62 70.0642
R4067 GNDA.n397 GNDA.n396 70.0642
R4068 GNDA.t58 GNDA.t184 69.5407
R4069 GNDA.t184 GNDA.t119 69.5407
R4070 GNDA.t121 GNDA.n1736 69.5407
R4071 GNDA.n1736 GNDA.t52 69.5407
R4072 GNDA.t174 GNDA.t165 69.5407
R4073 GNDA.t175 GNDA.t174 69.5407
R4074 GNDA.n1502 GNDA.t228 65.8183
R4075 GNDA.n1504 GNDA.t228 65.8183
R4076 GNDA.n1510 GNDA.t228 65.8183
R4077 GNDA.n1518 GNDA.t228 65.8183
R4078 GNDA.n1520 GNDA.t228 65.8183
R4079 GNDA.n1526 GNDA.t228 65.8183
R4080 GNDA.n1528 GNDA.t228 65.8183
R4081 GNDA.n1546 GNDA.t228 65.8183
R4082 GNDA.n1543 GNDA.t228 65.8183
R4083 GNDA.n1537 GNDA.t228 65.8183
R4084 GNDA.n1534 GNDA.t228 65.8183
R4085 GNDA.n1318 GNDA.t230 65.8183
R4086 GNDA.n1324 GNDA.t230 65.8183
R4087 GNDA.n1326 GNDA.t230 65.8183
R4088 GNDA.n1334 GNDA.t230 65.8183
R4089 GNDA.n1340 GNDA.t230 65.8183
R4090 GNDA.n1342 GNDA.t230 65.8183
R4091 GNDA.n1348 GNDA.t230 65.8183
R4092 GNDA.n1365 GNDA.t230 65.8183
R4093 GNDA.n1359 GNDA.t230 65.8183
R4094 GNDA.n1357 GNDA.t230 65.8183
R4095 GNDA.n1351 GNDA.t230 65.8183
R4096 GNDA.n2217 GNDA.t313 65.8183
R4097 GNDA.n2223 GNDA.t313 65.8183
R4098 GNDA.n2225 GNDA.t313 65.8183
R4099 GNDA.n2233 GNDA.t313 65.8183
R4100 GNDA.n2239 GNDA.t313 65.8183
R4101 GNDA.n2241 GNDA.t313 65.8183
R4102 GNDA.n2247 GNDA.t313 65.8183
R4103 GNDA.n2264 GNDA.t313 65.8183
R4104 GNDA.n2258 GNDA.t313 65.8183
R4105 GNDA.n2256 GNDA.t313 65.8183
R4106 GNDA.n2250 GNDA.t313 65.8183
R4107 GNDA.n803 GNDA.t279 65.8183
R4108 GNDA.n809 GNDA.t279 65.8183
R4109 GNDA.n811 GNDA.t279 65.8183
R4110 GNDA.n819 GNDA.t279 65.8183
R4111 GNDA.n825 GNDA.t279 65.8183
R4112 GNDA.n827 GNDA.t279 65.8183
R4113 GNDA.n833 GNDA.t279 65.8183
R4114 GNDA.n850 GNDA.t279 65.8183
R4115 GNDA.n844 GNDA.t279 65.8183
R4116 GNDA.n842 GNDA.t279 65.8183
R4117 GNDA.n836 GNDA.t279 65.8183
R4118 GNDA.n1003 GNDA.t283 65.8183
R4119 GNDA.n1009 GNDA.t283 65.8183
R4120 GNDA.n1011 GNDA.t283 65.8183
R4121 GNDA.n1019 GNDA.t283 65.8183
R4122 GNDA.n1025 GNDA.t283 65.8183
R4123 GNDA.n1027 GNDA.t283 65.8183
R4124 GNDA.n1033 GNDA.t283 65.8183
R4125 GNDA.n1050 GNDA.t283 65.8183
R4126 GNDA.n1044 GNDA.t283 65.8183
R4127 GNDA.n1042 GNDA.t283 65.8183
R4128 GNDA.n1036 GNDA.t283 65.8183
R4129 GNDA.n1127 GNDA.t261 65.8183
R4130 GNDA.n1133 GNDA.t261 65.8183
R4131 GNDA.n1135 GNDA.t261 65.8183
R4132 GNDA.n1143 GNDA.t261 65.8183
R4133 GNDA.n1149 GNDA.t261 65.8183
R4134 GNDA.n1151 GNDA.t261 65.8183
R4135 GNDA.n1157 GNDA.t261 65.8183
R4136 GNDA.n1174 GNDA.t261 65.8183
R4137 GNDA.n1168 GNDA.t261 65.8183
R4138 GNDA.n1166 GNDA.t261 65.8183
R4139 GNDA.n1160 GNDA.t261 65.8183
R4140 GNDA.n1771 GNDA.t260 65.8183
R4141 GNDA.n1773 GNDA.t260 65.8183
R4142 GNDA.n1779 GNDA.t260 65.8183
R4143 GNDA.n1787 GNDA.t260 65.8183
R4144 GNDA.n1789 GNDA.t260 65.8183
R4145 GNDA.n1795 GNDA.t260 65.8183
R4146 GNDA.n1797 GNDA.t260 65.8183
R4147 GNDA.n1815 GNDA.t260 65.8183
R4148 GNDA.n1812 GNDA.t260 65.8183
R4149 GNDA.n1806 GNDA.t260 65.8183
R4150 GNDA.n1803 GNDA.t260 65.8183
R4151 GNDA.n1980 GNDA.t262 65.8183
R4152 GNDA.n1982 GNDA.t262 65.8183
R4153 GNDA.n1988 GNDA.t262 65.8183
R4154 GNDA.n1996 GNDA.t262 65.8183
R4155 GNDA.n1998 GNDA.t262 65.8183
R4156 GNDA.n2004 GNDA.t262 65.8183
R4157 GNDA.n2006 GNDA.t262 65.8183
R4158 GNDA.n2024 GNDA.t262 65.8183
R4159 GNDA.n2021 GNDA.t262 65.8183
R4160 GNDA.n2015 GNDA.t262 65.8183
R4161 GNDA.n2012 GNDA.t262 65.8183
R4162 GNDA.n2362 GNDA.t247 65.8183
R4163 GNDA.n2368 GNDA.t247 65.8183
R4164 GNDA.n2370 GNDA.t247 65.8183
R4165 GNDA.n2378 GNDA.t247 65.8183
R4166 GNDA.n2384 GNDA.t247 65.8183
R4167 GNDA.n2386 GNDA.t247 65.8183
R4168 GNDA.n2392 GNDA.t247 65.8183
R4169 GNDA.n2409 GNDA.t247 65.8183
R4170 GNDA.n2403 GNDA.t247 65.8183
R4171 GNDA.n2401 GNDA.t247 65.8183
R4172 GNDA.n2395 GNDA.t247 65.8183
R4173 GNDA.n2412 GNDA.t247 65.8183
R4174 GNDA.n2421 GNDA.t247 65.8183
R4175 GNDA.n2347 GNDA.t247 65.8183
R4176 GNDA.n2345 GNDA.t247 65.8183
R4177 GNDA.n1961 GNDA.t262 65.8183
R4178 GNDA.n2043 GNDA.t262 65.8183
R4179 GNDA.n1947 GNDA.t262 65.8183
R4180 GNDA.n2058 GNDA.t262 65.8183
R4181 GNDA.n1750 GNDA.t260 65.8183
R4182 GNDA.n1834 GNDA.t260 65.8183
R4183 GNDA.n1610 GNDA.t260 65.8183
R4184 GNDA.n1846 GNDA.t260 65.8183
R4185 GNDA.n1104 GNDA.t261 65.8183
R4186 GNDA.n1185 GNDA.t261 65.8183
R4187 GNDA.n1095 GNDA.t261 65.8183
R4188 GNDA.n1196 GNDA.t261 65.8183
R4189 GNDA.t283 GNDA.n702 65.8183
R4190 GNDA.n973 GNDA.t283 65.8183
R4191 GNDA.n987 GNDA.t283 65.8183
R4192 GNDA.n969 GNDA.t283 65.8183
R4193 GNDA.n776 GNDA.t279 65.8183
R4194 GNDA.n861 GNDA.t279 65.8183
R4195 GNDA.n767 GNDA.t279 65.8183
R4196 GNDA.n872 GNDA.t279 65.8183
R4197 GNDA.n304 GNDA.t313 65.8183
R4198 GNDA.n2275 GNDA.t313 65.8183
R4199 GNDA.n295 GNDA.t313 65.8183
R4200 GNDA.n2286 GNDA.t313 65.8183
R4201 GNDA.n1296 GNDA.t230 65.8183
R4202 GNDA.n1376 GNDA.t230 65.8183
R4203 GNDA.n1287 GNDA.t230 65.8183
R4204 GNDA.n1387 GNDA.t230 65.8183
R4205 GNDA.n1474 GNDA.t228 65.8183
R4206 GNDA.n1471 GNDA.t228 65.8183
R4207 GNDA.n1485 GNDA.t228 65.8183
R4208 GNDA.n1461 GNDA.t228 65.8183
R4209 GNDA.n102 GNDA.n82 65.6476
R4210 GNDA.t229 GNDA.n621 65.4161
R4211 GNDA.n2077 GNDA.t231 65.4161
R4212 GNDA.n2112 GNDA.t248 65.4161
R4213 GNDA.n471 GNDA.n470 64.0005
R4214 GNDA.n470 GNDA.n346 64.0005
R4215 GNDA.t116 GNDA.t149 63.2189
R4216 GNDA.t64 GNDA.t86 63.2189
R4217 GNDA.t132 GNDA.t344 63.2189
R4218 GNDA.t146 GNDA.t92 63.2189
R4219 GNDA.t185 GNDA.n1726 63.2189
R4220 GNDA.t172 GNDA.n1651 63.2189
R4221 GNDA.t229 GNDA.n588 60.9488
R4222 GNDA.t231 GNDA.n187 60.9488
R4223 GNDA.n474 GNDA.t153 60.7372
R4224 GNDA.n440 GNDA.t333 60.7372
R4225 GNDA.t125 GNDA.n409 60.7372
R4226 GNDA.t239 GNDA.t217 59.0043
R4227 GNDA.t290 GNDA.t9 59.0043
R4228 GNDA.t308 GNDA.t186 56.897
R4229 GNDA.t61 GNDA.t169 56.897
R4230 GNDA.n1725 GNDA.t255 56.897
R4231 GNDA.n1650 GNDA.t277 56.897
R4232 GNDA.t319 GNDA.t35 56.897
R4233 GNDA.t285 GNDA.t182 56.897
R4234 GNDA.n522 GNDA.n172 55.2535
R4235 GNDA.n2194 GNDA.n169 55.2535
R4236 GNDA.n2442 GNDA.n93 55.2535
R4237 GNDA.n2359 GNDA.t247 55.2026
R4238 GNDA.t262 GNDA.n1939 55.2026
R4239 GNDA.n1765 GNDA.t260 55.2026
R4240 GNDA.t261 GNDA.n1086 55.2026
R4241 GNDA.n1000 GNDA.t283 55.2026
R4242 GNDA.t279 GNDA.n758 55.2026
R4243 GNDA.t313 GNDA.n286 55.2026
R4244 GNDA.t230 GNDA.n1278 55.2026
R4245 GNDA.n1496 GNDA.t228 55.2026
R4246 GNDA.n484 GNDA.t179 54.7898
R4247 GNDA.n2479 GNDA.t177 54.7898
R4248 GNDA.n1512 GNDA.t228 54.4705
R4249 GNDA.n1332 GNDA.t230 54.4705
R4250 GNDA.n2231 GNDA.t313 54.4705
R4251 GNDA.n817 GNDA.t279 54.4705
R4252 GNDA.n1017 GNDA.t283 54.4705
R4253 GNDA.n1141 GNDA.t261 54.4705
R4254 GNDA.n1781 GNDA.t260 54.4705
R4255 GNDA.n1990 GNDA.t262 54.4705
R4256 GNDA.n2376 GNDA.t247 54.4705
R4257 GNDA.n436 GNDA.n435 54.4005
R4258 GNDA.n1487 GNDA.n1461 53.3664
R4259 GNDA.n1485 GNDA.n1484 53.3664
R4260 GNDA.n1476 GNDA.n1471 53.3664
R4261 GNDA.n1474 GNDA.n1403 53.3664
R4262 GNDA.n1534 GNDA.n1533 53.3664
R4263 GNDA.n1538 GNDA.n1537 53.3664
R4264 GNDA.n1543 GNDA.n1542 53.3664
R4265 GNDA.n1546 GNDA.n1545 53.3664
R4266 GNDA.n1518 GNDA.n1517 53.3664
R4267 GNDA.n1521 GNDA.n1520 53.3664
R4268 GNDA.n1526 GNDA.n1525 53.3664
R4269 GNDA.n1529 GNDA.n1528 53.3664
R4270 GNDA.n1511 GNDA.n1510 53.3664
R4271 GNDA.n1504 GNDA.n1414 53.3664
R4272 GNDA.n1503 GNDA.n1502 53.3664
R4273 GNDA.n1502 GNDA.n1501 53.3664
R4274 GNDA.n1505 GNDA.n1504 53.3664
R4275 GNDA.n1510 GNDA.n1509 53.3664
R4276 GNDA.n1519 GNDA.n1518 53.3664
R4277 GNDA.n1520 GNDA.n1410 53.3664
R4278 GNDA.n1527 GNDA.n1526 53.3664
R4279 GNDA.n1528 GNDA.n1408 53.3664
R4280 GNDA.n1547 GNDA.n1546 53.3664
R4281 GNDA.n1544 GNDA.n1543 53.3664
R4282 GNDA.n1537 GNDA.n1405 53.3664
R4283 GNDA.n1535 GNDA.n1534 53.3664
R4284 GNDA.n1387 GNDA.n1386 53.3664
R4285 GNDA.n1378 GNDA.n1287 53.3664
R4286 GNDA.n1376 GNDA.n1375 53.3664
R4287 GNDA.n1367 GNDA.n1296 53.3664
R4288 GNDA.n1351 GNDA.n1350 53.3664
R4289 GNDA.n1357 GNDA.n1356 53.3664
R4290 GNDA.n1360 GNDA.n1359 53.3664
R4291 GNDA.n1365 GNDA.n1364 53.3664
R4292 GNDA.n1335 GNDA.n1334 53.3664
R4293 GNDA.n1340 GNDA.n1339 53.3664
R4294 GNDA.n1343 GNDA.n1342 53.3664
R4295 GNDA.n1348 GNDA.n1347 53.3664
R4296 GNDA.n1326 GNDA.n1311 53.3664
R4297 GNDA.n1325 GNDA.n1324 53.3664
R4298 GNDA.n1318 GNDA.n1313 53.3664
R4299 GNDA.n1319 GNDA.n1318 53.3664
R4300 GNDA.n1324 GNDA.n1323 53.3664
R4301 GNDA.n1327 GNDA.n1326 53.3664
R4302 GNDA.n1334 GNDA.n1309 53.3664
R4303 GNDA.n1341 GNDA.n1340 53.3664
R4304 GNDA.n1342 GNDA.n1307 53.3664
R4305 GNDA.n1349 GNDA.n1348 53.3664
R4306 GNDA.n1366 GNDA.n1365 53.3664
R4307 GNDA.n1359 GNDA.n1302 53.3664
R4308 GNDA.n1358 GNDA.n1357 53.3664
R4309 GNDA.n1352 GNDA.n1351 53.3664
R4310 GNDA.n2286 GNDA.n2285 53.3664
R4311 GNDA.n2277 GNDA.n295 53.3664
R4312 GNDA.n2275 GNDA.n2274 53.3664
R4313 GNDA.n2266 GNDA.n304 53.3664
R4314 GNDA.n2250 GNDA.n2249 53.3664
R4315 GNDA.n2256 GNDA.n2255 53.3664
R4316 GNDA.n2259 GNDA.n2258 53.3664
R4317 GNDA.n2264 GNDA.n2263 53.3664
R4318 GNDA.n2234 GNDA.n2233 53.3664
R4319 GNDA.n2239 GNDA.n2238 53.3664
R4320 GNDA.n2242 GNDA.n2241 53.3664
R4321 GNDA.n2247 GNDA.n2246 53.3664
R4322 GNDA.n2225 GNDA.n2210 53.3664
R4323 GNDA.n2224 GNDA.n2223 53.3664
R4324 GNDA.n2217 GNDA.n2212 53.3664
R4325 GNDA.n2218 GNDA.n2217 53.3664
R4326 GNDA.n2223 GNDA.n2222 53.3664
R4327 GNDA.n2226 GNDA.n2225 53.3664
R4328 GNDA.n2233 GNDA.n2208 53.3664
R4329 GNDA.n2240 GNDA.n2239 53.3664
R4330 GNDA.n2241 GNDA.n2206 53.3664
R4331 GNDA.n2248 GNDA.n2247 53.3664
R4332 GNDA.n2265 GNDA.n2264 53.3664
R4333 GNDA.n2258 GNDA.n2201 53.3664
R4334 GNDA.n2257 GNDA.n2256 53.3664
R4335 GNDA.n2251 GNDA.n2250 53.3664
R4336 GNDA.n872 GNDA.n871 53.3664
R4337 GNDA.n863 GNDA.n767 53.3664
R4338 GNDA.n861 GNDA.n860 53.3664
R4339 GNDA.n852 GNDA.n776 53.3664
R4340 GNDA.n836 GNDA.n835 53.3664
R4341 GNDA.n842 GNDA.n841 53.3664
R4342 GNDA.n845 GNDA.n844 53.3664
R4343 GNDA.n850 GNDA.n849 53.3664
R4344 GNDA.n820 GNDA.n819 53.3664
R4345 GNDA.n825 GNDA.n824 53.3664
R4346 GNDA.n828 GNDA.n827 53.3664
R4347 GNDA.n833 GNDA.n832 53.3664
R4348 GNDA.n811 GNDA.n796 53.3664
R4349 GNDA.n810 GNDA.n809 53.3664
R4350 GNDA.n803 GNDA.n798 53.3664
R4351 GNDA.n804 GNDA.n803 53.3664
R4352 GNDA.n809 GNDA.n808 53.3664
R4353 GNDA.n812 GNDA.n811 53.3664
R4354 GNDA.n819 GNDA.n794 53.3664
R4355 GNDA.n826 GNDA.n825 53.3664
R4356 GNDA.n827 GNDA.n792 53.3664
R4357 GNDA.n834 GNDA.n833 53.3664
R4358 GNDA.n851 GNDA.n850 53.3664
R4359 GNDA.n844 GNDA.n787 53.3664
R4360 GNDA.n843 GNDA.n842 53.3664
R4361 GNDA.n837 GNDA.n836 53.3664
R4362 GNDA.n970 GNDA.n969 53.3664
R4363 GNDA.n987 GNDA.n986 53.3664
R4364 GNDA.n974 GNDA.n973 53.3664
R4365 GNDA.n1052 GNDA.n702 53.3664
R4366 GNDA.n1036 GNDA.n1035 53.3664
R4367 GNDA.n1042 GNDA.n1041 53.3664
R4368 GNDA.n1045 GNDA.n1044 53.3664
R4369 GNDA.n1050 GNDA.n1049 53.3664
R4370 GNDA.n1020 GNDA.n1019 53.3664
R4371 GNDA.n1025 GNDA.n1024 53.3664
R4372 GNDA.n1028 GNDA.n1027 53.3664
R4373 GNDA.n1033 GNDA.n1032 53.3664
R4374 GNDA.n1011 GNDA.n712 53.3664
R4375 GNDA.n1010 GNDA.n1009 53.3664
R4376 GNDA.n1003 GNDA.n714 53.3664
R4377 GNDA.n1004 GNDA.n1003 53.3664
R4378 GNDA.n1009 GNDA.n1008 53.3664
R4379 GNDA.n1012 GNDA.n1011 53.3664
R4380 GNDA.n1019 GNDA.n710 53.3664
R4381 GNDA.n1026 GNDA.n1025 53.3664
R4382 GNDA.n1027 GNDA.n708 53.3664
R4383 GNDA.n1034 GNDA.n1033 53.3664
R4384 GNDA.n1051 GNDA.n1050 53.3664
R4385 GNDA.n1044 GNDA.n703 53.3664
R4386 GNDA.n1043 GNDA.n1042 53.3664
R4387 GNDA.n1037 GNDA.n1036 53.3664
R4388 GNDA.n1196 GNDA.n1195 53.3664
R4389 GNDA.n1187 GNDA.n1095 53.3664
R4390 GNDA.n1185 GNDA.n1184 53.3664
R4391 GNDA.n1176 GNDA.n1104 53.3664
R4392 GNDA.n1160 GNDA.n1159 53.3664
R4393 GNDA.n1166 GNDA.n1165 53.3664
R4394 GNDA.n1169 GNDA.n1168 53.3664
R4395 GNDA.n1174 GNDA.n1173 53.3664
R4396 GNDA.n1144 GNDA.n1143 53.3664
R4397 GNDA.n1149 GNDA.n1148 53.3664
R4398 GNDA.n1152 GNDA.n1151 53.3664
R4399 GNDA.n1157 GNDA.n1156 53.3664
R4400 GNDA.n1135 GNDA.n1120 53.3664
R4401 GNDA.n1134 GNDA.n1133 53.3664
R4402 GNDA.n1127 GNDA.n1122 53.3664
R4403 GNDA.n1128 GNDA.n1127 53.3664
R4404 GNDA.n1133 GNDA.n1132 53.3664
R4405 GNDA.n1136 GNDA.n1135 53.3664
R4406 GNDA.n1143 GNDA.n1118 53.3664
R4407 GNDA.n1150 GNDA.n1149 53.3664
R4408 GNDA.n1151 GNDA.n1116 53.3664
R4409 GNDA.n1158 GNDA.n1157 53.3664
R4410 GNDA.n1175 GNDA.n1174 53.3664
R4411 GNDA.n1168 GNDA.n1111 53.3664
R4412 GNDA.n1167 GNDA.n1166 53.3664
R4413 GNDA.n1161 GNDA.n1160 53.3664
R4414 GNDA.n1846 GNDA.n1845 53.3664
R4415 GNDA.n1611 GNDA.n1610 53.3664
R4416 GNDA.n1834 GNDA.n1833 53.3664
R4417 GNDA.n1751 GNDA.n1750 53.3664
R4418 GNDA.n1803 GNDA.n1802 53.3664
R4419 GNDA.n1807 GNDA.n1806 53.3664
R4420 GNDA.n1812 GNDA.n1811 53.3664
R4421 GNDA.n1815 GNDA.n1814 53.3664
R4422 GNDA.n1787 GNDA.n1786 53.3664
R4423 GNDA.n1790 GNDA.n1789 53.3664
R4424 GNDA.n1795 GNDA.n1794 53.3664
R4425 GNDA.n1798 GNDA.n1797 53.3664
R4426 GNDA.n1780 GNDA.n1779 53.3664
R4427 GNDA.n1773 GNDA.n1762 53.3664
R4428 GNDA.n1772 GNDA.n1771 53.3664
R4429 GNDA.n1771 GNDA.n1770 53.3664
R4430 GNDA.n1774 GNDA.n1773 53.3664
R4431 GNDA.n1779 GNDA.n1778 53.3664
R4432 GNDA.n1788 GNDA.n1787 53.3664
R4433 GNDA.n1789 GNDA.n1758 53.3664
R4434 GNDA.n1796 GNDA.n1795 53.3664
R4435 GNDA.n1797 GNDA.n1756 53.3664
R4436 GNDA.n1816 GNDA.n1815 53.3664
R4437 GNDA.n1813 GNDA.n1812 53.3664
R4438 GNDA.n1806 GNDA.n1753 53.3664
R4439 GNDA.n1804 GNDA.n1803 53.3664
R4440 GNDA.n2058 GNDA.n2057 53.3664
R4441 GNDA.n2045 GNDA.n1947 53.3664
R4442 GNDA.n2043 GNDA.n2042 53.3664
R4443 GNDA.n1962 GNDA.n1961 53.3664
R4444 GNDA.n2012 GNDA.n2011 53.3664
R4445 GNDA.n2016 GNDA.n2015 53.3664
R4446 GNDA.n2021 GNDA.n2020 53.3664
R4447 GNDA.n2024 GNDA.n2023 53.3664
R4448 GNDA.n1996 GNDA.n1995 53.3664
R4449 GNDA.n1999 GNDA.n1998 53.3664
R4450 GNDA.n2004 GNDA.n2003 53.3664
R4451 GNDA.n2007 GNDA.n2006 53.3664
R4452 GNDA.n1989 GNDA.n1988 53.3664
R4453 GNDA.n1982 GNDA.n1973 53.3664
R4454 GNDA.n1981 GNDA.n1980 53.3664
R4455 GNDA.n1980 GNDA.n1979 53.3664
R4456 GNDA.n1983 GNDA.n1982 53.3664
R4457 GNDA.n1988 GNDA.n1987 53.3664
R4458 GNDA.n1997 GNDA.n1996 53.3664
R4459 GNDA.n1998 GNDA.n1969 53.3664
R4460 GNDA.n2005 GNDA.n2004 53.3664
R4461 GNDA.n2006 GNDA.n1967 53.3664
R4462 GNDA.n2025 GNDA.n2024 53.3664
R4463 GNDA.n2022 GNDA.n2021 53.3664
R4464 GNDA.n2015 GNDA.n1964 53.3664
R4465 GNDA.n2013 GNDA.n2012 53.3664
R4466 GNDA.n2346 GNDA.n2345 53.3664
R4467 GNDA.n2347 GNDA.n125 53.3664
R4468 GNDA.n2421 GNDA.n2420 53.3664
R4469 GNDA.n2412 GNDA.n2411 53.3664
R4470 GNDA.n2395 GNDA.n2394 53.3664
R4471 GNDA.n2401 GNDA.n2400 53.3664
R4472 GNDA.n2404 GNDA.n2403 53.3664
R4473 GNDA.n2409 GNDA.n2408 53.3664
R4474 GNDA.n2379 GNDA.n2378 53.3664
R4475 GNDA.n2384 GNDA.n2383 53.3664
R4476 GNDA.n2387 GNDA.n2386 53.3664
R4477 GNDA.n2392 GNDA.n2391 53.3664
R4478 GNDA.n2370 GNDA.n135 53.3664
R4479 GNDA.n2369 GNDA.n2368 53.3664
R4480 GNDA.n2362 GNDA.n137 53.3664
R4481 GNDA.n2363 GNDA.n2362 53.3664
R4482 GNDA.n2368 GNDA.n2367 53.3664
R4483 GNDA.n2371 GNDA.n2370 53.3664
R4484 GNDA.n2378 GNDA.n133 53.3664
R4485 GNDA.n2385 GNDA.n2384 53.3664
R4486 GNDA.n2386 GNDA.n131 53.3664
R4487 GNDA.n2393 GNDA.n2392 53.3664
R4488 GNDA.n2410 GNDA.n2409 53.3664
R4489 GNDA.n2403 GNDA.n126 53.3664
R4490 GNDA.n2402 GNDA.n2401 53.3664
R4491 GNDA.n2396 GNDA.n2395 53.3664
R4492 GNDA.n2413 GNDA.n2412 53.3664
R4493 GNDA.n2422 GNDA.n2421 53.3664
R4494 GNDA.n2348 GNDA.n2347 53.3664
R4495 GNDA.n2345 GNDA.n140 53.3664
R4496 GNDA.n1961 GNDA.n1949 53.3664
R4497 GNDA.n2044 GNDA.n2043 53.3664
R4498 GNDA.n1947 GNDA.n1941 53.3664
R4499 GNDA.n2059 GNDA.n2058 53.3664
R4500 GNDA.n1750 GNDA.n1612 53.3664
R4501 GNDA.n1835 GNDA.n1834 53.3664
R4502 GNDA.n1610 GNDA.n618 53.3664
R4503 GNDA.n1847 GNDA.n1846 53.3664
R4504 GNDA.n1104 GNDA.n1097 53.3664
R4505 GNDA.n1186 GNDA.n1185 53.3664
R4506 GNDA.n1095 GNDA.n1088 53.3664
R4507 GNDA.n1197 GNDA.n1196 53.3664
R4508 GNDA.n975 GNDA.n702 53.3664
R4509 GNDA.n973 GNDA.n971 53.3664
R4510 GNDA.n988 GNDA.n987 53.3664
R4511 GNDA.n969 GNDA.n717 53.3664
R4512 GNDA.n776 GNDA.n769 53.3664
R4513 GNDA.n862 GNDA.n861 53.3664
R4514 GNDA.n767 GNDA.n760 53.3664
R4515 GNDA.n873 GNDA.n872 53.3664
R4516 GNDA.n304 GNDA.n297 53.3664
R4517 GNDA.n2276 GNDA.n2275 53.3664
R4518 GNDA.n295 GNDA.n288 53.3664
R4519 GNDA.n2287 GNDA.n2286 53.3664
R4520 GNDA.n1296 GNDA.n1289 53.3664
R4521 GNDA.n1377 GNDA.n1376 53.3664
R4522 GNDA.n1287 GNDA.n1280 53.3664
R4523 GNDA.n1388 GNDA.n1387 53.3664
R4524 GNDA.n1475 GNDA.n1474 53.3664
R4525 GNDA.n1471 GNDA.n1463 53.3664
R4526 GNDA.n1486 GNDA.n1485 53.3664
R4527 GNDA.n1461 GNDA.n1418 53.3664
R4528 GNDA.n2131 GNDA.n2128 52.5182
R4529 GNDA.n2332 GNDA.n173 52.5182
R4530 GNDA.n230 GNDA.n216 52.5182
R4531 GNDA.n472 GNDA.n471 51.2005
R4532 GNDA.n346 GNDA.n345 51.2005
R4533 GNDA.n403 GNDA.n370 50.5752
R4534 GNDA.n2472 GNDA.n2471 50.5752
R4535 GNDA.n2137 GNDA.n531 49.2359
R4536 GNDA.n2138 GNDA.n2137 49.2359
R4537 GNDA.n2140 GNDA.n2138 49.2359
R4538 GNDA.n2140 GNDA.n2139 49.2359
R4539 GNDA.n2147 GNDA.n2146 49.2359
R4540 GNDA.n2148 GNDA.n2147 49.2359
R4541 GNDA.n2148 GNDA.n519 49.2359
R4542 GNDA.n2155 GNDA.n522 49.2359
R4543 GNDA.n504 GNDA.n173 49.2359
R4544 GNDA.n510 GNDA.n504 49.2359
R4545 GNDA.n2166 GNDA.n2164 49.2359
R4546 GNDA.n2166 GNDA.n2165 49.2359
R4547 GNDA.n2190 GNDA.n2189 49.2359
R4548 GNDA.n2194 GNDA.n2193 49.2359
R4549 GNDA.n230 GNDA.n229 49.2359
R4550 GNDA.n229 GNDA.n228 49.2359
R4551 GNDA.n228 GNDA.n219 49.2359
R4552 GNDA.n222 GNDA.n219 49.2359
R4553 GNDA.n222 GNDA.n117 49.2359
R4554 GNDA.n2427 GNDA.n104 49.2359
R4555 GNDA.n2434 GNDA.n108 49.2359
R4556 GNDA.n111 GNDA.n108 49.2359
R4557 GNDA.n111 GNDA.n93 49.2359
R4558 GNDA.n78 GNDA.t12 49.0451
R4559 GNDA.t338 GNDA.n387 49.0451
R4560 GNDA.n354 GNDA.t210 48.0005
R4561 GNDA.n354 GNDA.t200 48.0005
R4562 GNDA.n351 GNDA.t212 48.0005
R4563 GNDA.n351 GNDA.t202 48.0005
R4564 GNDA.n350 GNDA.t208 48.0005
R4565 GNDA.n350 GNDA.t198 48.0005
R4566 GNDA.n348 GNDA.t214 48.0005
R4567 GNDA.n348 GNDA.t204 48.0005
R4568 GNDA.n347 GNDA.t216 48.0005
R4569 GNDA.n347 GNDA.t206 48.0005
R4570 GNDA.t248 GNDA.n2332 47.5947
R4571 GNDA.n2175 GNDA.n2174 47.5947
R4572 GNDA.t248 GNDA.n172 47.0476
R4573 GNDA.t248 GNDA.n169 47.0476
R4574 GNDA.t16 GNDA.t112 46.3607
R4575 GNDA.t112 GNDA.t50 46.3607
R4576 GNDA.n460 GNDA.t87 46.3607
R4577 GNDA.t83 GNDA.t45 46.3607
R4578 GNDA.t101 GNDA.t83 46.3607
R4579 GNDA.n391 GNDA.n385 44.8005
R4580 GNDA.n2462 GNDA.n2461 44.8005
R4581 GNDA.t99 GNDA.t39 44.2534
R4582 GNDA.t0 GNDA.t117 44.2534
R4583 GNDA.n120 GNDA.n118 43.0993
R4584 GNDA.t236 GNDA.t341 42.1461
R4585 GNDA.t85 GNDA.t157 42.1461
R4586 GNDA.t11 GNDA.t81 42.1461
R4587 GNDA.t326 GNDA.t181 42.1461
R4588 GNDA.t323 GNDA.t342 42.1461
R4589 GNDA.t98 GNDA.t137 42.1461
R4590 GNDA.t233 GNDA.t66 42.1461
R4591 GNDA.t41 GNDA.t296 42.1461
R4592 GNDA.t219 GNDA.t51 42.1461
R4593 GNDA.t151 GNDA.t1 42.1461
R4594 GNDA.t76 GNDA.t221 42.1461
R4595 GNDA.t324 GNDA.t180 42.1461
R4596 GNDA.t74 GNDA.t19 42.1461
R4597 GNDA.t346 GNDA.t147 42.1461
R4598 GNDA.t17 GNDA.t328 42.1461
R4599 GNDA.t264 GNDA.t331 42.1461
R4600 GNDA.n2163 GNDA.n510 42.1241
R4601 GNDA.t78 GNDA.n2464 39.7033
R4602 GNDA.n389 GNDA.t91 39.7033
R4603 GNDA.n484 GNDA.t50 37.9315
R4604 GNDA.n410 GNDA.t94 37.9315
R4605 GNDA.t159 GNDA.t97 37.9315
R4606 GNDA.n2479 GNDA.t45 37.9315
R4607 GNDA.n2190 GNDA.n308 36.6535
R4608 GNDA.n24 GNDA.n23 35.438
R4609 GNDA.n2497 GNDA.n12 35.438
R4610 GNDA.n2128 GNDA.n496 33.9182
R4611 GNDA.t130 GNDA.t236 33.717
R4612 GNDA.t68 GNDA.t62 33.717
R4613 GNDA.t157 GNDA.t26 33.717
R4614 GNDA.t81 GNDA.t115 33.717
R4615 GNDA.t140 GNDA.t326 33.717
R4616 GNDA.t342 GNDA.t339 33.717
R4617 GNDA.t66 GNDA.t239 33.717
R4618 GNDA.t290 GNDA.t41 33.717
R4619 GNDA.t5 GNDA.t151 33.717
R4620 GNDA.t332 GNDA.t76 33.717
R4621 GNDA.t340 GNDA.t324 33.717
R4622 GNDA.t141 GNDA.t74 33.717
R4623 GNDA.t139 GNDA.t346 33.717
R4624 GNDA.t111 GNDA.t17 33.717
R4625 GNDA.t79 GNDA.t264 33.717
R4626 GNDA.t187 GNDA.t56 31.6097
R4627 GNDA.t109 GNDA.t161 31.6097
R4628 GNDA.t7 GNDA.t167 31.6097
R4629 GNDA.t37 GNDA.t171 31.6097
R4630 GNDA.n2131 GNDA.n2130 31.1829
R4631 GNDA.n2188 GNDA.n312 31.1829
R4632 GNDA.n216 GNDA.n168 31.1829
R4633 GNDA.t229 GNDA.n622 31.0997
R4634 GNDA.n537 GNDA.t248 31.0997
R4635 GNDA.n64 GNDA.t337 30.3614
R4636 GNDA.n76 GNDA.t336 30.3614
R4637 GNDA.t70 GNDA.n388 30.3614
R4638 GNDA.n382 GNDA.t6 30.3614
R4639 GNDA.t149 GNDA.t105 29.5024
R4640 GNDA.t179 GNDA.t64 29.5024
R4641 GNDA.t344 GNDA.t177 29.5024
R4642 GNDA.t92 GNDA.t103 29.5024
R4643 GNDA.n491 GNDA.n490 28.413
R4644 GNDA.n72 GNDA.n49 28.413
R4645 GNDA.n2177 GNDA.n99 28.1318
R4646 GNDA.n380 GNDA.n379 28.038
R4647 GNDA.n60 GNDA.n39 28.038
R4648 GNDA.n1732 GNDA.n1628 27.8193
R4649 GNDA.n1730 GNDA.n1729 27.8193
R4650 GNDA.n1515 GNDA.n1514 27.5561
R4651 GNDA.n1330 GNDA.n1310 27.5561
R4652 GNDA.n2229 GNDA.n2209 27.5561
R4653 GNDA.n815 GNDA.n795 27.5561
R4654 GNDA.n1015 GNDA.n711 27.5561
R4655 GNDA.n1139 GNDA.n1119 27.5561
R4656 GNDA.n1784 GNDA.n1783 27.5561
R4657 GNDA.n1993 GNDA.n1992 27.5561
R4658 GNDA.n2374 GNDA.n134 27.5561
R4659 GNDA.n588 GNDA.n569 26.9584
R4660 GNDA.n2302 GNDA.n187 26.9584
R4661 GNDA.n2139 GNDA.t248 25.7123
R4662 GNDA.n2165 GNDA.t248 25.7123
R4663 GNDA.t248 GNDA.n117 25.7123
R4664 GNDA.t12 GNDA.n76 25.6905
R4665 GNDA.n388 GNDA.t338 25.6905
R4666 GNDA.n487 GNDA.n486 25.6005
R4667 GNDA.n2477 GNDA.n2476 25.6005
R4668 GNDA.n1713 GNDA.n1711 25.2879
R4669 GNDA.n1702 GNDA.n1647 25.2879
R4670 GNDA.n1677 GNDA.t166 24.0005
R4671 GNDA.n1677 GNDA.t176 24.0005
R4672 GNDA.n1675 GNDA.t118 24.0005
R4673 GNDA.n1675 GNDA.t36 24.0005
R4674 GNDA.n1673 GNDA.t168 24.0005
R4675 GNDA.n1673 GNDA.t38 24.0005
R4676 GNDA.n1671 GNDA.t124 24.0005
R4677 GNDA.n1671 GNDA.t55 24.0005
R4678 GNDA.n1669 GNDA.t53 24.0005
R4679 GNDA.n1669 GNDA.t108 24.0005
R4680 GNDA.n1667 GNDA.t164 24.0005
R4681 GNDA.n1667 GNDA.t122 24.0005
R4682 GNDA.n1665 GNDA.t44 24.0005
R4683 GNDA.n1665 GNDA.t34 24.0005
R4684 GNDA.n1663 GNDA.t57 24.0005
R4685 GNDA.n1663 GNDA.t110 24.0005
R4686 GNDA.n1661 GNDA.t170 24.0005
R4687 GNDA.n1661 GNDA.t40 24.0005
R4688 GNDA.n1660 GNDA.t59 24.0005
R4689 GNDA.n1660 GNDA.t120 24.0005
R4690 GNDA.n1532 GNDA.n1531 23.6449
R4691 GNDA.n1306 GNDA.n1305 23.6449
R4692 GNDA.n2205 GNDA.n2204 23.6449
R4693 GNDA.n791 GNDA.n790 23.6449
R4694 GNDA.n707 GNDA.n706 23.6449
R4695 GNDA.n1115 GNDA.n1114 23.6449
R4696 GNDA.n1801 GNDA.n1800 23.6449
R4697 GNDA.n2010 GNDA.n2009 23.6449
R4698 GNDA.n130 GNDA.n129 23.6449
R4699 GNDA.n2146 GNDA.t248 23.5241
R4700 GNDA.n2174 GNDA.t248 23.5241
R4701 GNDA.n2427 GNDA.t248 23.5241
R4702 GNDA.n401 GNDA.n380 22.4005
R4703 GNDA.n436 GNDA.n434 22.4005
R4704 GNDA.n2488 GNDA.n2487 22.4005
R4705 GNDA.n2469 GNDA.n60 22.4005
R4706 GNDA.t335 GNDA.t23 21.8829
R4707 GNDA.n560 GNDA.n499 21.4917
R4708 GNDA.n2085 GNDA.t231 21.4482
R4709 GNDA.n1658 GNDA.n1655 21.3338
R4710 GNDA.n1657 GNDA.n1656 21.3338
R4711 GNDA.n1733 GNDA.n1627 21.3338
R4712 GNDA.n1626 GNDA.n1625 21.3338
R4713 GNDA.n1630 GNDA.n1629 21.3338
R4714 GNDA.n1715 GNDA.n1714 21.3338
R4715 GNDA.n457 GNDA.n453 21.3338
R4716 GNDA.n452 GNDA.n451 21.3338
R4717 GNDA.n346 GNDA.n343 21.3338
R4718 GNDA.n345 GNDA.n344 21.3338
R4719 GNDA.n339 GNDA.n338 21.3338
R4720 GNDA.n473 GNDA.n340 21.3338
R4721 GNDA.n472 GNDA.n341 21.3338
R4722 GNDA.n471 GNDA.n342 21.3338
R4723 GNDA.n464 GNDA.n463 21.3338
R4724 GNDA.n359 GNDA.n358 21.3338
R4725 GNDA.n363 GNDA.n362 21.3338
R4726 GNDA.n364 GNDA.n361 21.3338
R4727 GNDA.n328 GNDA.n327 21.3338
R4728 GNDA.n324 GNDA.n323 21.3338
R4729 GNDA.n332 GNDA.n331 21.3338
R4730 GNDA.n330 GNDA.n329 21.3338
R4731 GNDA.n52 GNDA.n51 21.3338
R4732 GNDA.n47 GNDA.n46 21.3338
R4733 GNDA.n45 GNDA.n44 21.3338
R4734 GNDA.n43 GNDA.n42 21.3338
R4735 GNDA.n1683 GNDA.n1680 21.1792
R4736 GNDA.t137 GNDA.n447 21.0733
R4737 GNDA.n2492 GNDA.t25 21.0733
R4738 GNDA.n2461 GNDA.n2460 20.288
R4739 GNDA.n385 GNDA.n320 20.1943
R4740 GNDA.n2499 GNDA.n0 19.9817
R4741 GNDA.n488 GNDA.n487 19.7255
R4742 GNDA.n2476 GNDA.n2475 19.7255
R4743 GNDA.n22 GNDA.t178 19.7005
R4744 GNDA.n22 GNDA.t191 19.7005
R4745 GNDA.n20 GNDA.t131 19.7005
R4746 GNDA.n20 GNDA.t46 19.7005
R4747 GNDA.n18 GNDA.t133 19.7005
R4748 GNDA.n18 GNDA.t20 19.7005
R4749 GNDA.n16 GNDA.t47 19.7005
R4750 GNDA.n16 GNDA.t104 19.7005
R4751 GNDA.n14 GNDA.t145 19.7005
R4752 GNDA.n14 GNDA.t102 19.7005
R4753 GNDA.n13 GNDA.t189 19.7005
R4754 GNDA.n13 GNDA.t13 19.7005
R4755 GNDA.n11 GNDA.t190 19.7005
R4756 GNDA.n11 GNDA.t127 19.7005
R4757 GNDA.n9 GNDA.t329 19.7005
R4758 GNDA.n9 GNDA.t148 19.7005
R4759 GNDA.n7 GNDA.t334 19.7005
R4760 GNDA.n7 GNDA.t100 19.7005
R4761 GNDA.n5 GNDA.t49 19.7005
R4762 GNDA.n5 GNDA.t129 19.7005
R4763 GNDA.n3 GNDA.t48 19.7005
R4764 GNDA.n3 GNDA.t156 19.7005
R4765 GNDA.n2 GNDA.t21 19.7005
R4766 GNDA.n2 GNDA.t195 19.7005
R4767 GNDA.n557 GNDA.n556 19.4279
R4768 GNDA.n1706 GNDA.n1704 19.2005
R4769 GNDA.n2160 GNDA.n2159 19.2005
R4770 GNDA.n2438 GNDA.n2437 19.2005
R4771 GNDA.n520 GNDA.n499 19.2005
R4772 GNDA.n2178 GNDA.n316 19.2005
R4773 GNDA.n1639 GNDA.n1618 19.2005
R4774 GNDA.t183 GNDA.t109 18.966
R4775 GNDA.t167 GNDA.t173 18.966
R4776 GNDA.n65 GNDA.n64 18.6842
R4777 GNDA.n394 GNDA.n382 18.6842
R4778 GNDA.n2130 GNDA.n531 18.0535
R4779 GNDA.n2189 GNDA.n2188 18.0535
R4780 GNDA.n1708 GNDA.n1639 17.613
R4781 GNDA.n2083 GNDA.n561 17.4917
R4782 GNDA.n2081 GNDA.n2080 16.9605
R4783 GNDA.n1881 GNDA.n596 16.9379
R4784 GNDA.n1601 GNDA.n633 16.9379
R4785 GNDA.n904 GNDA.n903 16.9379
R4786 GNDA.n448 GNDA.t115 16.9236
R4787 GNDA.n444 GNDA.t203 16.9236
R4788 GNDA.n461 GNDA.t211 16.9236
R4789 GNDA.t340 GNDA.n29 16.9236
R4790 GNDA.t111 GNDA.n30 16.9236
R4791 GNDA.n2499 GNDA.n2498 16.883
R4792 GNDA.t333 GNDA.t73 16.8587
R4793 GNDA.t341 GNDA.t125 16.8587
R4794 GNDA.t130 GNDA.t94 16.8587
R4795 GNDA.t62 GNDA.t85 16.8587
R4796 GNDA.t26 GNDA.t11 16.8587
R4797 GNDA.t181 GNDA.t115 16.8587
R4798 GNDA.t140 GNDA.t323 16.8587
R4799 GNDA.t339 GNDA.t98 16.8587
R4800 GNDA.t330 GNDA.t233 16.8587
R4801 GNDA.t296 GNDA.t25 16.8587
R4802 GNDA.t51 GNDA.t5 16.8587
R4803 GNDA.t1 GNDA.t332 16.8587
R4804 GNDA.t221 GNDA.t340 16.8587
R4805 GNDA.t180 GNDA.t141 16.8587
R4806 GNDA.t19 GNDA.t139 16.8587
R4807 GNDA.t147 GNDA.t111 16.8587
R4808 GNDA.t328 GNDA.t79 16.8587
R4809 GNDA.t331 GNDA.t126 16.8587
R4810 GNDA.t248 GNDA.n168 16.4123
R4811 GNDA.n1514 GNDA.n1413 16.0005
R4812 GNDA.n1508 GNDA.n1413 16.0005
R4813 GNDA.n1508 GNDA.n1507 16.0005
R4814 GNDA.n1507 GNDA.n1506 16.0005
R4815 GNDA.n1506 GNDA.n1415 16.0005
R4816 GNDA.n1500 GNDA.n1415 16.0005
R4817 GNDA.n1500 GNDA.n1499 16.0005
R4818 GNDA.n1499 GNDA.n1498 16.0005
R4819 GNDA.n1516 GNDA.n1515 16.0005
R4820 GNDA.n1516 GNDA.n1411 16.0005
R4821 GNDA.n1522 GNDA.n1411 16.0005
R4822 GNDA.n1523 GNDA.n1522 16.0005
R4823 GNDA.n1524 GNDA.n1523 16.0005
R4824 GNDA.n1524 GNDA.n1409 16.0005
R4825 GNDA.n1530 GNDA.n1409 16.0005
R4826 GNDA.n1531 GNDA.n1530 16.0005
R4827 GNDA.n1532 GNDA.n1407 16.0005
R4828 GNDA.n1407 GNDA.n1406 16.0005
R4829 GNDA.n1539 GNDA.n1406 16.0005
R4830 GNDA.n1540 GNDA.n1539 16.0005
R4831 GNDA.n1541 GNDA.n1404 16.0005
R4832 GNDA.n1404 GNDA.n1402 16.0005
R4833 GNDA.n1548 GNDA.n1402 16.0005
R4834 GNDA.n1330 GNDA.n1329 16.0005
R4835 GNDA.n1329 GNDA.n1328 16.0005
R4836 GNDA.n1328 GNDA.n1312 16.0005
R4837 GNDA.n1322 GNDA.n1312 16.0005
R4838 GNDA.n1322 GNDA.n1321 16.0005
R4839 GNDA.n1321 GNDA.n1320 16.0005
R4840 GNDA.n1320 GNDA.n1314 16.0005
R4841 GNDA.n1315 GNDA.n1314 16.0005
R4842 GNDA.n1336 GNDA.n1310 16.0005
R4843 GNDA.n1337 GNDA.n1336 16.0005
R4844 GNDA.n1338 GNDA.n1337 16.0005
R4845 GNDA.n1338 GNDA.n1308 16.0005
R4846 GNDA.n1344 GNDA.n1308 16.0005
R4847 GNDA.n1345 GNDA.n1344 16.0005
R4848 GNDA.n1346 GNDA.n1345 16.0005
R4849 GNDA.n1346 GNDA.n1306 16.0005
R4850 GNDA.n1353 GNDA.n1305 16.0005
R4851 GNDA.n1354 GNDA.n1353 16.0005
R4852 GNDA.n1355 GNDA.n1354 16.0005
R4853 GNDA.n1355 GNDA.n1303 16.0005
R4854 GNDA.n1362 GNDA.n1361 16.0005
R4855 GNDA.n1363 GNDA.n1362 16.0005
R4856 GNDA.n1363 GNDA.n1301 16.0005
R4857 GNDA.n2229 GNDA.n2228 16.0005
R4858 GNDA.n2228 GNDA.n2227 16.0005
R4859 GNDA.n2227 GNDA.n2211 16.0005
R4860 GNDA.n2221 GNDA.n2211 16.0005
R4861 GNDA.n2221 GNDA.n2220 16.0005
R4862 GNDA.n2220 GNDA.n2219 16.0005
R4863 GNDA.n2219 GNDA.n2213 16.0005
R4864 GNDA.n2214 GNDA.n2213 16.0005
R4865 GNDA.n2235 GNDA.n2209 16.0005
R4866 GNDA.n2236 GNDA.n2235 16.0005
R4867 GNDA.n2237 GNDA.n2236 16.0005
R4868 GNDA.n2237 GNDA.n2207 16.0005
R4869 GNDA.n2243 GNDA.n2207 16.0005
R4870 GNDA.n2244 GNDA.n2243 16.0005
R4871 GNDA.n2245 GNDA.n2244 16.0005
R4872 GNDA.n2245 GNDA.n2205 16.0005
R4873 GNDA.n2252 GNDA.n2204 16.0005
R4874 GNDA.n2253 GNDA.n2252 16.0005
R4875 GNDA.n2254 GNDA.n2253 16.0005
R4876 GNDA.n2254 GNDA.n2202 16.0005
R4877 GNDA.n2261 GNDA.n2260 16.0005
R4878 GNDA.n2262 GNDA.n2261 16.0005
R4879 GNDA.n2262 GNDA.n2200 16.0005
R4880 GNDA.n815 GNDA.n814 16.0005
R4881 GNDA.n814 GNDA.n813 16.0005
R4882 GNDA.n813 GNDA.n797 16.0005
R4883 GNDA.n807 GNDA.n797 16.0005
R4884 GNDA.n807 GNDA.n806 16.0005
R4885 GNDA.n806 GNDA.n805 16.0005
R4886 GNDA.n805 GNDA.n799 16.0005
R4887 GNDA.n800 GNDA.n799 16.0005
R4888 GNDA.n821 GNDA.n795 16.0005
R4889 GNDA.n822 GNDA.n821 16.0005
R4890 GNDA.n823 GNDA.n822 16.0005
R4891 GNDA.n823 GNDA.n793 16.0005
R4892 GNDA.n829 GNDA.n793 16.0005
R4893 GNDA.n830 GNDA.n829 16.0005
R4894 GNDA.n831 GNDA.n830 16.0005
R4895 GNDA.n831 GNDA.n791 16.0005
R4896 GNDA.n838 GNDA.n790 16.0005
R4897 GNDA.n839 GNDA.n838 16.0005
R4898 GNDA.n840 GNDA.n839 16.0005
R4899 GNDA.n840 GNDA.n788 16.0005
R4900 GNDA.n847 GNDA.n846 16.0005
R4901 GNDA.n848 GNDA.n847 16.0005
R4902 GNDA.n848 GNDA.n786 16.0005
R4903 GNDA.n1015 GNDA.n1014 16.0005
R4904 GNDA.n1014 GNDA.n1013 16.0005
R4905 GNDA.n1013 GNDA.n713 16.0005
R4906 GNDA.n1007 GNDA.n713 16.0005
R4907 GNDA.n1007 GNDA.n1006 16.0005
R4908 GNDA.n1006 GNDA.n1005 16.0005
R4909 GNDA.n1005 GNDA.n715 16.0005
R4910 GNDA.n716 GNDA.n715 16.0005
R4911 GNDA.n1021 GNDA.n711 16.0005
R4912 GNDA.n1022 GNDA.n1021 16.0005
R4913 GNDA.n1023 GNDA.n1022 16.0005
R4914 GNDA.n1023 GNDA.n709 16.0005
R4915 GNDA.n1029 GNDA.n709 16.0005
R4916 GNDA.n1030 GNDA.n1029 16.0005
R4917 GNDA.n1031 GNDA.n1030 16.0005
R4918 GNDA.n1031 GNDA.n707 16.0005
R4919 GNDA.n1038 GNDA.n706 16.0005
R4920 GNDA.n1039 GNDA.n1038 16.0005
R4921 GNDA.n1040 GNDA.n1039 16.0005
R4922 GNDA.n1040 GNDA.n704 16.0005
R4923 GNDA.n1047 GNDA.n1046 16.0005
R4924 GNDA.n1048 GNDA.n1047 16.0005
R4925 GNDA.n1048 GNDA.n699 16.0005
R4926 GNDA.n1139 GNDA.n1138 16.0005
R4927 GNDA.n1138 GNDA.n1137 16.0005
R4928 GNDA.n1137 GNDA.n1121 16.0005
R4929 GNDA.n1131 GNDA.n1121 16.0005
R4930 GNDA.n1131 GNDA.n1130 16.0005
R4931 GNDA.n1130 GNDA.n1129 16.0005
R4932 GNDA.n1129 GNDA.n1123 16.0005
R4933 GNDA.n1124 GNDA.n1123 16.0005
R4934 GNDA.n1145 GNDA.n1119 16.0005
R4935 GNDA.n1146 GNDA.n1145 16.0005
R4936 GNDA.n1147 GNDA.n1146 16.0005
R4937 GNDA.n1147 GNDA.n1117 16.0005
R4938 GNDA.n1153 GNDA.n1117 16.0005
R4939 GNDA.n1154 GNDA.n1153 16.0005
R4940 GNDA.n1155 GNDA.n1154 16.0005
R4941 GNDA.n1155 GNDA.n1115 16.0005
R4942 GNDA.n1162 GNDA.n1114 16.0005
R4943 GNDA.n1163 GNDA.n1162 16.0005
R4944 GNDA.n1164 GNDA.n1163 16.0005
R4945 GNDA.n1164 GNDA.n1112 16.0005
R4946 GNDA.n1171 GNDA.n1170 16.0005
R4947 GNDA.n1172 GNDA.n1171 16.0005
R4948 GNDA.n1172 GNDA.n1110 16.0005
R4949 GNDA.n1783 GNDA.n1761 16.0005
R4950 GNDA.n1777 GNDA.n1761 16.0005
R4951 GNDA.n1777 GNDA.n1776 16.0005
R4952 GNDA.n1776 GNDA.n1775 16.0005
R4953 GNDA.n1775 GNDA.n1763 16.0005
R4954 GNDA.n1769 GNDA.n1763 16.0005
R4955 GNDA.n1769 GNDA.n1768 16.0005
R4956 GNDA.n1768 GNDA.n1767 16.0005
R4957 GNDA.n1785 GNDA.n1784 16.0005
R4958 GNDA.n1785 GNDA.n1759 16.0005
R4959 GNDA.n1791 GNDA.n1759 16.0005
R4960 GNDA.n1792 GNDA.n1791 16.0005
R4961 GNDA.n1793 GNDA.n1792 16.0005
R4962 GNDA.n1793 GNDA.n1757 16.0005
R4963 GNDA.n1799 GNDA.n1757 16.0005
R4964 GNDA.n1800 GNDA.n1799 16.0005
R4965 GNDA.n1801 GNDA.n1755 16.0005
R4966 GNDA.n1755 GNDA.n1754 16.0005
R4967 GNDA.n1808 GNDA.n1754 16.0005
R4968 GNDA.n1809 GNDA.n1808 16.0005
R4969 GNDA.n1810 GNDA.n1752 16.0005
R4970 GNDA.n1752 GNDA.n1749 16.0005
R4971 GNDA.n1817 GNDA.n1749 16.0005
R4972 GNDA.n1992 GNDA.n1972 16.0005
R4973 GNDA.n1986 GNDA.n1972 16.0005
R4974 GNDA.n1986 GNDA.n1985 16.0005
R4975 GNDA.n1985 GNDA.n1984 16.0005
R4976 GNDA.n1984 GNDA.n1974 16.0005
R4977 GNDA.n1978 GNDA.n1974 16.0005
R4978 GNDA.n1978 GNDA.n1977 16.0005
R4979 GNDA.n1977 GNDA.n1937 16.0005
R4980 GNDA.n1994 GNDA.n1993 16.0005
R4981 GNDA.n1994 GNDA.n1970 16.0005
R4982 GNDA.n2000 GNDA.n1970 16.0005
R4983 GNDA.n2001 GNDA.n2000 16.0005
R4984 GNDA.n2002 GNDA.n2001 16.0005
R4985 GNDA.n2002 GNDA.n1968 16.0005
R4986 GNDA.n2008 GNDA.n1968 16.0005
R4987 GNDA.n2009 GNDA.n2008 16.0005
R4988 GNDA.n2010 GNDA.n1966 16.0005
R4989 GNDA.n1966 GNDA.n1965 16.0005
R4990 GNDA.n2017 GNDA.n1965 16.0005
R4991 GNDA.n2018 GNDA.n2017 16.0005
R4992 GNDA.n2019 GNDA.n1963 16.0005
R4993 GNDA.n1963 GNDA.n1960 16.0005
R4994 GNDA.n2026 GNDA.n1960 16.0005
R4995 GNDA.n2374 GNDA.n2373 16.0005
R4996 GNDA.n2373 GNDA.n2372 16.0005
R4997 GNDA.n2372 GNDA.n136 16.0005
R4998 GNDA.n2366 GNDA.n136 16.0005
R4999 GNDA.n2366 GNDA.n2365 16.0005
R5000 GNDA.n2365 GNDA.n2364 16.0005
R5001 GNDA.n2364 GNDA.n138 16.0005
R5002 GNDA.n139 GNDA.n138 16.0005
R5003 GNDA.n2380 GNDA.n134 16.0005
R5004 GNDA.n2381 GNDA.n2380 16.0005
R5005 GNDA.n2382 GNDA.n2381 16.0005
R5006 GNDA.n2382 GNDA.n132 16.0005
R5007 GNDA.n2388 GNDA.n132 16.0005
R5008 GNDA.n2389 GNDA.n2388 16.0005
R5009 GNDA.n2390 GNDA.n2389 16.0005
R5010 GNDA.n2390 GNDA.n130 16.0005
R5011 GNDA.n2397 GNDA.n129 16.0005
R5012 GNDA.n2398 GNDA.n2397 16.0005
R5013 GNDA.n2399 GNDA.n2398 16.0005
R5014 GNDA.n2399 GNDA.n127 16.0005
R5015 GNDA.n2406 GNDA.n2405 16.0005
R5016 GNDA.n2407 GNDA.n2406 16.0005
R5017 GNDA.n2407 GNDA.n90 16.0005
R5018 GNDA.n2083 GNDA.n2082 16.0005
R5019 GNDA.n2082 GNDA.n2081 16.0005
R5020 GNDA.t336 GNDA.t2 15.8816
R5021 GNDA.t63 GNDA.t70 15.8816
R5022 GNDA.n1710 GNDA.n1636 15.363
R5023 GNDA.n1723 GNDA.n1710 15.363
R5024 GNDA.t3 GNDA.n2155 14.7711
R5025 GNDA.t23 GNDA.n2434 14.7711
R5026 GNDA.n2496 GNDA.n2495 14.6443
R5027 GNDA.n468 GNDA.n467 14.2068
R5028 GNDA.n468 GNDA.n357 14.2068
R5029 GNDA.n378 GNDA.n377 14.0505
R5030 GNDA.n2482 GNDA.n2481 14.0505
R5031 GNDA.n1541 GNDA 14.0449
R5032 GNDA.n1361 GNDA 14.0449
R5033 GNDA.n2260 GNDA 14.0449
R5034 GNDA.n846 GNDA 14.0449
R5035 GNDA.n1046 GNDA 14.0449
R5036 GNDA.n1170 GNDA 14.0449
R5037 GNDA.n1810 GNDA 14.0449
R5038 GNDA.n2019 GNDA 14.0449
R5039 GNDA.n2405 GNDA 14.0449
R5040 GNDA.n2487 GNDA.n2486 13.8005
R5041 GNDA.n434 GNDA.n433 13.8005
R5042 GNDA.n1707 GNDA.n1706 13.8005
R5043 GNDA.n1680 GNDA.n561 13.7706
R5044 GNDA.t305 GNDA.n440 13.4979
R5045 GNDA.n409 GNDA.t155 13.4979
R5046 GNDA.t302 GNDA.n474 13.4979
R5047 GNDA.n2298 GNDA.n257 12.9309
R5048 GNDA.n1397 GNDA.n656 12.9309
R5049 GNDA.n721 GNDA.n634 12.9309
R5050 GNDA.n1208 GNDA.n182 12.9309
R5051 GNDA.n321 GNDA.n320 12.8005
R5052 GNDA.n2460 GNDA.n69 12.8005
R5053 GNDA.n369 GNDA.t245 12.6442
R5054 GNDA.t226 GNDA.t30 12.6442
R5055 GNDA.t136 GNDA.t28 12.6442
R5056 GNDA.n447 GNDA.t330 12.6442
R5057 GNDA.n2492 GNDA.t219 12.6442
R5058 GNDA.t27 GNDA.n2491 12.6442
R5059 GNDA.t321 GNDA.t14 12.6442
R5060 GNDA.t258 GNDA.t134 12.6442
R5061 GNDA.n55 GNDA.t242 12.6442
R5062 GNDA.n2193 GNDA.n308 12.5829
R5063 GNDA.n218 GNDA.n215 12.4126
R5064 GNDA.n2133 GNDA.n533 12.4126
R5065 GNDA.n506 GNDA.n174 12.4126
R5066 GNDA.n1271 GNDA.n1221 11.6369
R5067 GNDA.n1271 GNDA.n1270 11.6369
R5068 GNDA.n1270 GNDA.n1269 11.6369
R5069 GNDA.n1269 GNDA.n1266 11.6369
R5070 GNDA.n1266 GNDA.n1265 11.6369
R5071 GNDA.n1265 GNDA.n1262 11.6369
R5072 GNDA.n1262 GNDA.n1261 11.6369
R5073 GNDA.n1261 GNDA.n1258 11.6369
R5074 GNDA.n1258 GNDA.n1257 11.6369
R5075 GNDA.n1257 GNDA.n1254 11.6369
R5076 GNDA.n1254 GNDA.n1253 11.6369
R5077 GNDA.n256 GNDA.n209 11.6369
R5078 GNDA.n251 GNDA.n209 11.6369
R5079 GNDA.n251 GNDA.n250 11.6369
R5080 GNDA.n250 GNDA.n211 11.6369
R5081 GNDA.n245 GNDA.n211 11.6369
R5082 GNDA.n245 GNDA.n244 11.6369
R5083 GNDA.n244 GNDA.n243 11.6369
R5084 GNDA.n243 GNDA.n213 11.6369
R5085 GNDA.n237 GNDA.n213 11.6369
R5086 GNDA.n237 GNDA.n236 11.6369
R5087 GNDA.n236 GNDA.n235 11.6369
R5088 GNDA.n221 GNDA.n218 11.6369
R5089 GNDA.n226 GNDA.n221 11.6369
R5090 GNDA.n226 GNDA.n225 11.6369
R5091 GNDA.n225 GNDA.n224 11.6369
R5092 GNDA.n224 GNDA.n114 11.6369
R5093 GNDA.n2429 GNDA.n114 11.6369
R5094 GNDA.n2432 GNDA.n2430 11.6369
R5095 GNDA.n2432 GNDA.n2431 11.6369
R5096 GNDA.n1882 GNDA.n1881 11.6369
R5097 GNDA.n1883 GNDA.n1882 11.6369
R5098 GNDA.n1883 GNDA.n594 11.6369
R5099 GNDA.n1889 GNDA.n594 11.6369
R5100 GNDA.n1890 GNDA.n1889 11.6369
R5101 GNDA.n1891 GNDA.n1890 11.6369
R5102 GNDA.n1891 GNDA.n592 11.6369
R5103 GNDA.n1897 GNDA.n592 11.6369
R5104 GNDA.n1898 GNDA.n1897 11.6369
R5105 GNDA.n1899 GNDA.n1898 11.6369
R5106 GNDA.n1899 GNDA.n589 11.6369
R5107 GNDA.n601 GNDA.n596 11.6369
R5108 GNDA.n1873 GNDA.n601 11.6369
R5109 GNDA.n1873 GNDA.n1872 11.6369
R5110 GNDA.n1872 GNDA.n1871 11.6369
R5111 GNDA.n1871 GNDA.n602 11.6369
R5112 GNDA.n1865 GNDA.n602 11.6369
R5113 GNDA.n1865 GNDA.n1864 11.6369
R5114 GNDA.n1864 GNDA.n1863 11.6369
R5115 GNDA.n1863 GNDA.n606 11.6369
R5116 GNDA.n688 GNDA.n687 11.6369
R5117 GNDA.n687 GNDA.n686 11.6369
R5118 GNDA.n686 GNDA.n684 11.6369
R5119 GNDA.n684 GNDA.n681 11.6369
R5120 GNDA.n681 GNDA.n680 11.6369
R5121 GNDA.n680 GNDA.n677 11.6369
R5122 GNDA.n677 GNDA.n676 11.6369
R5123 GNDA.n676 GNDA.n673 11.6369
R5124 GNDA.n673 GNDA.n672 11.6369
R5125 GNDA.n672 GNDA.n669 11.6369
R5126 GNDA.n669 GNDA.n668 11.6369
R5127 GNDA.n1601 GNDA.n1600 11.6369
R5128 GNDA.n1600 GNDA.n1599 11.6369
R5129 GNDA.n1599 GNDA.n1597 11.6369
R5130 GNDA.n1597 GNDA.n1594 11.6369
R5131 GNDA.n1594 GNDA.n1593 11.6369
R5132 GNDA.n1593 GNDA.n1590 11.6369
R5133 GNDA.n1590 GNDA.n1589 11.6369
R5134 GNDA.n1589 GNDA.n1586 11.6369
R5135 GNDA.n1586 GNDA.n1585 11.6369
R5136 GNDA.n1585 GNDA.n1582 11.6369
R5137 GNDA.n1582 GNDA.n1581 11.6369
R5138 GNDA.n1430 GNDA.n633 11.6369
R5139 GNDA.n1436 GNDA.n1430 11.6369
R5140 GNDA.n1437 GNDA.n1436 11.6369
R5141 GNDA.n1438 GNDA.n1437 11.6369
R5142 GNDA.n1438 GNDA.n1426 11.6369
R5143 GNDA.n1444 GNDA.n1426 11.6369
R5144 GNDA.n1445 GNDA.n1444 11.6369
R5145 GNDA.n1446 GNDA.n1445 11.6369
R5146 GNDA.n1446 GNDA.n1422 11.6369
R5147 GNDA.n903 GNDA.n742 11.6369
R5148 GNDA.n897 GNDA.n742 11.6369
R5149 GNDA.n897 GNDA.n896 11.6369
R5150 GNDA.n896 GNDA.n895 11.6369
R5151 GNDA.n895 GNDA.n746 11.6369
R5152 GNDA.n889 GNDA.n746 11.6369
R5153 GNDA.n889 GNDA.n888 11.6369
R5154 GNDA.n888 GNDA.n887 11.6369
R5155 GNDA.n887 GNDA.n750 11.6369
R5156 GNDA.n905 GNDA.n904 11.6369
R5157 GNDA.n905 GNDA.n738 11.6369
R5158 GNDA.n912 GNDA.n738 11.6369
R5159 GNDA.n913 GNDA.n912 11.6369
R5160 GNDA.n914 GNDA.n913 11.6369
R5161 GNDA.n914 GNDA.n736 11.6369
R5162 GNDA.n919 GNDA.n736 11.6369
R5163 GNDA.n920 GNDA.n919 11.6369
R5164 GNDA.n922 GNDA.n920 11.6369
R5165 GNDA.n922 GNDA.n921 11.6369
R5166 GNDA.n921 GNDA.n733 11.6369
R5167 GNDA.n2071 GNDA.n566 11.6369
R5168 GNDA.n2072 GNDA.n2071 11.6369
R5169 GNDA.n2073 GNDA.n2072 11.6369
R5170 GNDA.n2073 GNDA.n562 11.6369
R5171 GNDA.n2079 GNDA.n562 11.6369
R5172 GNDA.n2089 GNDA.n552 11.6369
R5173 GNDA.n2090 GNDA.n2089 11.6369
R5174 GNDA.n2092 GNDA.n2090 11.6369
R5175 GNDA.n2092 GNDA.n2091 11.6369
R5176 GNDA.n2091 GNDA.n549 11.6369
R5177 GNDA.n2106 GNDA.n543 11.6369
R5178 GNDA.n2107 GNDA.n2106 11.6369
R5179 GNDA.n2108 GNDA.n2107 11.6369
R5180 GNDA.n2108 GNDA.n539 11.6369
R5181 GNDA.n2114 GNDA.n539 11.6369
R5182 GNDA.n2115 GNDA.n2114 11.6369
R5183 GNDA.n2116 GNDA.n2115 11.6369
R5184 GNDA.n2116 GNDA.n535 11.6369
R5185 GNDA.n2123 GNDA.n535 11.6369
R5186 GNDA.n2124 GNDA.n2123 11.6369
R5187 GNDA.n2125 GNDA.n2124 11.6369
R5188 GNDA.n2134 GNDA.n2133 11.6369
R5189 GNDA.n2135 GNDA.n2134 11.6369
R5190 GNDA.n2135 GNDA.n529 11.6369
R5191 GNDA.n2142 GNDA.n529 11.6369
R5192 GNDA.n2143 GNDA.n2142 11.6369
R5193 GNDA.n2144 GNDA.n2143 11.6369
R5194 GNDA.n2150 GNDA.n526 11.6369
R5195 GNDA.n2151 GNDA.n2150 11.6369
R5196 GNDA.n2310 GNDA.n2309 11.6369
R5197 GNDA.n2311 GNDA.n2310 11.6369
R5198 GNDA.n2311 GNDA.n180 11.6369
R5199 GNDA.n2317 GNDA.n180 11.6369
R5200 GNDA.n2318 GNDA.n2317 11.6369
R5201 GNDA.n2319 GNDA.n2318 11.6369
R5202 GNDA.n2319 GNDA.n178 11.6369
R5203 GNDA.n2325 GNDA.n178 11.6369
R5204 GNDA.n2326 GNDA.n2325 11.6369
R5205 GNDA.n2327 GNDA.n2326 11.6369
R5206 GNDA.n2327 GNDA.n176 11.6369
R5207 GNDA.n507 GNDA.n506 11.6369
R5208 GNDA.n508 GNDA.n507 11.6369
R5209 GNDA.n508 GNDA.n502 11.6369
R5210 GNDA.n2168 GNDA.n502 11.6369
R5211 GNDA.n2169 GNDA.n2168 11.6369
R5212 GNDA.n2172 GNDA.n2169 11.6369
R5213 GNDA.n2171 GNDA.n2170 11.6369
R5214 GNDA.n2170 GNDA.n311 11.6369
R5215 GNDA.n2430 GNDA 11.5076
R5216 GNDA GNDA.n526 11.5076
R5217 GNDA GNDA.n2171 11.5076
R5218 GNDA.n2431 GNDA.n91 11.4026
R5219 GNDA.n2152 GNDA.n2151 11.4026
R5220 GNDA.n311 GNDA.n310 11.4026
R5221 GNDA.n1856 GNDA.n606 11.249
R5222 GNDA.n1454 GNDA.n1422 11.249
R5223 GNDA.n753 GNDA.n750 11.249
R5224 GNDA.n470 GNDA.n469 11.0505
R5225 GNDA.n2080 GNDA.n2079 10.4732
R5226 GNDA.n433 GNDA.n1 9.938
R5227 GNDA.n1709 GNDA.n1637 9.78488
R5228 GNDA GNDA.n0 9.67325
R5229 GNDA.n2086 GNDA.n2085 9.65197
R5230 GNDA.n2486 GNDA.n2485 9.6255
R5231 GNDA.n1705 GNDA.t192 9.6005
R5232 GNDA.n1705 GNDA.t194 9.6005
R5233 GNDA.n431 GNDA.t69 9.6005
R5234 GNDA.n431 GNDA.t158 9.6005
R5235 GNDA.n429 GNDA.t82 9.6005
R5236 GNDA.n429 GNDA.t327 9.6005
R5237 GNDA.n427 GNDA.t343 9.6005
R5238 GNDA.n427 GNDA.t138 9.6005
R5239 GNDA.n425 GNDA.t67 9.6005
R5240 GNDA.n425 GNDA.t218 9.6005
R5241 GNDA.n423 GNDA.t72 9.6005
R5242 GNDA.n423 GNDA.t88 9.6005
R5243 GNDA.n421 GNDA.t160 9.6005
R5244 GNDA.n421 GNDA.t32 9.6005
R5245 GNDA.n419 GNDA.t10 9.6005
R5246 GNDA.n419 GNDA.t42 9.6005
R5247 GNDA.n417 GNDA.t220 9.6005
R5248 GNDA.n417 GNDA.t152 9.6005
R5249 GNDA.n415 GNDA.t77 9.6005
R5250 GNDA.n415 GNDA.t325 9.6005
R5251 GNDA.n413 GNDA.t75 9.6005
R5252 GNDA.n413 GNDA.t347 9.6005
R5253 GNDA.n35 GNDA.t18 9.6005
R5254 GNDA.n35 GNDA.t265 9.6005
R5255 GNDA.n1638 GNDA.t188 9.6005
R5256 GNDA.n1638 GNDA.t196 9.6005
R5257 GNDA.n1707 GNDA.n1640 9.37925
R5258 GNDA.n2157 GNDA.n519 9.30051
R5259 GNDA.n2435 GNDA.n104 9.30051
R5260 GNDA.n455 GNDA.n356 9.3005
R5261 GNDA.n2156 GNDA.t3 8.75345
R5262 GNDA.n235 GNDA.n215 8.66313
R5263 GNDA.n2125 GNDA.n533 8.66313
R5264 GNDA.n176 GNDA.n174 8.66313
R5265 GNDA.n1253 GNDA.n257 8.53383
R5266 GNDA.n656 GNDA.n589 8.53383
R5267 GNDA.n668 GNDA.n182 8.53383
R5268 GNDA.n1581 GNDA.n634 8.53383
R5269 GNDA.n733 GNDA.n732 8.53383
R5270 GNDA.n549 GNDA.n548 8.53383
R5271 GNDA.n1679 GNDA.n1678 8.44175
R5272 GNDA.t97 GNDA.n460 8.42962
R5273 GNDA.n1498 GNDA.n1417 8.35606
R5274 GNDA.n1315 GNDA.n659 8.35606
R5275 GNDA.n2214 GNDA.n283 8.35606
R5276 GNDA.n800 GNDA.n756 8.35606
R5277 GNDA.n965 GNDA.n716 8.35606
R5278 GNDA.n1124 GNDA.n1083 8.35606
R5279 GNDA.n1767 GNDA.n610 8.35606
R5280 GNDA.n2063 GNDA.n1937 8.35606
R5281 GNDA.n2337 GNDA.n139 8.35606
R5282 GNDA.n1710 GNDA.n1709 7.71925
R5283 GNDA.t60 GNDA.n2156 7.65933
R5284 GNDA.n2164 GNDA.n2163 7.11227
R5285 GNDA.n65 GNDA.t142 7.00687
R5286 GNDA.t114 GNDA.n78 7.00687
R5287 GNDA.n387 GNDA.t143 7.00687
R5288 GNDA.t154 GNDA.n394 7.00687
R5289 GNDA.n2497 GNDA.n2496 6.7505
R5290 GNDA.n2496 GNDA.n24 6.688
R5291 GNDA.n376 GNDA.n1 6.563
R5292 GNDA.n2485 GNDA.n2484 6.563
R5293 GNDA.n2179 GNDA.n2178 6.4005
R5294 GNDA.n490 GNDA.n489 6.4005
R5295 GNDA.n2474 GNDA.n49 6.4005
R5296 GNDA.t39 GNDA.n1713 6.32234
R5297 GNDA.t162 GNDA.t293 6.32234
R5298 GNDA.n1737 GNDA.t121 6.32234
R5299 GNDA.n1649 GNDA.t52 6.32234
R5300 GNDA.t281 GNDA.t318 6.32234
R5301 GNDA.t117 GNDA.n1647 6.32234
R5302 GNDA.n2485 GNDA.n24 5.03175
R5303 GNDA.n557 GNDA.n0 5.02613
R5304 GNDA.n2157 GNDA.t96 4.92404
R5305 GNDA GNDA.n2499 4.8321
R5306 GNDA.n1823 GNDA.n1822 4.6085
R5307 GNDA.n2032 GNDA.n2031 4.6085
R5308 GNDA.n2445 GNDA.n2444 4.6085
R5309 GNDA.n784 GNDA.n777 4.6085
R5310 GNDA.n1211 GNDA.n1210 4.6085
R5311 GNDA.n1108 GNDA.n525 4.6085
R5312 GNDA.n1555 GNDA.n1399 4.6085
R5313 GNDA.n1299 GNDA.n208 4.6085
R5314 GNDA.n2198 GNDA.n305 4.6085
R5315 GNDA.n1249 GNDA.n1222 4.55161
R5316 GNDA.n1906 GNDA.n587 4.55161
R5317 GNDA.n1577 GNDA.n635 4.55161
R5318 GNDA.n931 GNDA.n730 4.55161
R5319 GNDA.n2100 GNDA.n544 4.55161
R5320 GNDA.n2305 GNDA.n183 4.55161
R5321 GNDA.n1818 GNDA.n575 4.5061
R5322 GNDA.n2028 GNDA.n147 4.5061
R5323 GNDA.n779 GNDA.n721 4.5061
R5324 GNDA.n1209 GNDA.n1208 4.5061
R5325 GNDA.n1556 GNDA.n1397 4.5061
R5326 GNDA.n2299 GNDA.n2298 4.5061
R5327 GNDA.n355 GNDA.n353 4.5005
R5328 GNDA.n469 GNDA.n468 4.5005
R5329 GNDA.n2498 GNDA.n2497 4.5005
R5330 GNDA.n1709 GNDA.n1708 4.5005
R5331 GNDA.n1221 GNDA.n656 4.39646
R5332 GNDA.n257 GNDA.n256 4.39646
R5333 GNDA.n688 GNDA.n634 4.39646
R5334 GNDA.n732 GNDA.n566 4.39646
R5335 GNDA.n548 GNDA.n543 4.39646
R5336 GNDA.n2309 GNDA.n182 4.39646
R5337 GNDA.n1936 GNDA.n575 4.3525
R5338 GNDA.n2336 GNDA.n147 4.3525
R5339 GNDA.n721 GNDA.n718 4.3525
R5340 GNDA.n1208 GNDA.n1207 4.3525
R5341 GNDA.n1397 GNDA.n1396 4.3525
R5342 GNDA.n2298 GNDA.n2297 4.3525
R5343 GNDA.n2064 GNDA.n1936 4.3013
R5344 GNDA.n2338 GNDA.n2336 4.3013
R5345 GNDA.n964 GNDA.n718 4.3013
R5346 GNDA.n1207 GNDA.n1204 4.3013
R5347 GNDA.n1396 GNDA.n1395 4.3013
R5348 GNDA.n2297 GNDA.n2294 4.3013
R5349 GNDA.n1249 GNDA.n1248 4.26717
R5350 GNDA.n1248 GNDA.n1245 4.26717
R5351 GNDA.n1245 GNDA.n1244 4.26717
R5352 GNDA.n1244 GNDA.n1241 4.26717
R5353 GNDA.n1241 GNDA.n1240 4.26717
R5354 GNDA.n1240 GNDA.n1237 4.26717
R5355 GNDA.n1236 GNDA.n1233 4.26717
R5356 GNDA.n1233 GNDA.n1232 4.26717
R5357 GNDA.n1906 GNDA.n585 4.26717
R5358 GNDA.n1912 GNDA.n585 4.26717
R5359 GNDA.n1912 GNDA.n583 4.26717
R5360 GNDA.n1918 GNDA.n583 4.26717
R5361 GNDA.n1918 GNDA.n581 4.26717
R5362 GNDA.n1925 GNDA.n581 4.26717
R5363 GNDA.n579 GNDA.n577 4.26717
R5364 GNDA.n1932 GNDA.n577 4.26717
R5365 GNDA.n1577 GNDA.n1576 4.26717
R5366 GNDA.n1576 GNDA.n640 4.26717
R5367 GNDA.n1571 GNDA.n640 4.26717
R5368 GNDA.n1571 GNDA.n1570 4.26717
R5369 GNDA.n1570 GNDA.n1569 4.26717
R5370 GNDA.n1569 GNDA.n648 4.26717
R5371 GNDA.n1563 GNDA.n1562 4.26717
R5372 GNDA.n1562 GNDA.n1561 4.26717
R5373 GNDA.n931 GNDA.n729 4.26717
R5374 GNDA.n937 GNDA.n729 4.26717
R5375 GNDA.n937 GNDA.n727 4.26717
R5376 GNDA.n943 GNDA.n727 4.26717
R5377 GNDA.n943 GNDA.n725 4.26717
R5378 GNDA.n951 GNDA.n725 4.26717
R5379 GNDA.n723 GNDA.n720 4.26717
R5380 GNDA.n958 GNDA.n720 4.26717
R5381 GNDA.n2100 GNDA.n545 4.26717
R5382 GNDA.n1061 GNDA.n545 4.26717
R5383 GNDA.n1062 GNDA.n1061 4.26717
R5384 GNDA.n1067 GNDA.n1062 4.26717
R5385 GNDA.n1068 GNDA.n1067 4.26717
R5386 GNDA.n1073 GNDA.n1068 4.26717
R5387 GNDA.n1079 GNDA.n1074 4.26717
R5388 GNDA.n1081 GNDA.n1079 4.26717
R5389 GNDA.n2305 GNDA.n184 4.26717
R5390 GNDA.n261 GNDA.n184 4.26717
R5391 GNDA.n262 GNDA.n261 4.26717
R5392 GNDA.n267 GNDA.n262 4.26717
R5393 GNDA.n268 GNDA.n267 4.26717
R5394 GNDA.n273 GNDA.n268 4.26717
R5395 GNDA.n279 GNDA.n274 4.26717
R5396 GNDA.n281 GNDA.n279 4.26717
R5397 GNDA.n754 GNDA.n753 4.2501
R5398 GNDA.n1455 GNDA.n1454 4.2501
R5399 GNDA GNDA.n1236 4.21976
R5400 GNDA GNDA.n579 4.21976
R5401 GNDA.n1563 GNDA 4.21976
R5402 GNDA GNDA.n723 4.21976
R5403 GNDA.n1074 GNDA 4.21976
R5404 GNDA.n274 GNDA 4.21976
R5405 GNDA.t311 GNDA.t252 4.21506
R5406 GNDA.n439 GNDA.t155 4.21506
R5407 GNDA.n410 GNDA.t68 4.21506
R5408 GNDA.n2491 GNDA.t153 4.21506
R5409 GNDA.t223 GNDA.t268 4.21506
R5410 GNDA.n1856 GNDA.n1855 4.1477
R5411 GNDA.n1232 GNDA.n147 4.12494
R5412 GNDA.n1932 GNDA.n575 4.12494
R5413 GNDA.n1561 GNDA.n1397 4.12494
R5414 GNDA.n958 GNDA.n721 4.12494
R5415 GNDA.n1208 GNDA.n1081 4.12494
R5416 GNDA.n2298 GNDA.n281 4.12494
R5417 GNDA.t96 GNDA.t60 3.82992
R5418 GNDA.n1708 GNDA.n1707 3.813
R5419 GNDA.n1640 GNDA 3.68412
R5420 GNDA.n615 GNDA.n614 3.5845
R5421 GNDA.n1849 GNDA.n1848 3.5845
R5422 GNDA.n1844 GNDA.n616 3.5845
R5423 GNDA.n1843 GNDA.n619 3.5845
R5424 GNDA.n1608 GNDA.n1607 3.5845
R5425 GNDA.n1837 GNDA.n1836 3.5845
R5426 GNDA.n1832 GNDA.n1609 3.5845
R5427 GNDA.n1831 GNDA.n1613 3.5845
R5428 GNDA.n1748 GNDA.n1747 3.5845
R5429 GNDA.n2062 GNDA.n2061 3.5845
R5430 GNDA.n1940 GNDA.n1938 3.5845
R5431 GNDA.n2056 GNDA.n1942 3.5845
R5432 GNDA.n2055 GNDA.n1943 3.5845
R5433 GNDA.n2047 GNDA.n2046 3.5845
R5434 GNDA.n1948 GNDA.n1946 3.5845
R5435 GNDA.n2041 GNDA.n1950 3.5845
R5436 GNDA.n2040 GNDA.n1951 3.5845
R5437 GNDA.n1959 GNDA.n1958 3.5845
R5438 GNDA.n2357 GNDA.n141 3.5845
R5439 GNDA.n2356 GNDA.n142 3.5845
R5440 GNDA.n2343 GNDA.n2342 3.5845
R5441 GNDA.n2350 GNDA.n2349 3.5845
R5442 GNDA.n2344 GNDA.n123 3.5845
R5443 GNDA.n2424 GNDA.n2423 3.5845
R5444 GNDA.n2419 GNDA.n124 3.5845
R5445 GNDA.n2418 GNDA.n2415 3.5845
R5446 GNDA.n2414 GNDA.n89 3.5845
R5447 GNDA.n876 GNDA.n875 3.5845
R5448 GNDA.n759 GNDA.n757 3.5845
R5449 GNDA.n870 GNDA.n761 3.5845
R5450 GNDA.n869 GNDA.n762 3.5845
R5451 GNDA.n865 GNDA.n864 3.5845
R5452 GNDA.n768 GNDA.n766 3.5845
R5453 GNDA.n859 GNDA.n770 3.5845
R5454 GNDA.n858 GNDA.n771 3.5845
R5455 GNDA.n854 GNDA.n853 3.5845
R5456 GNDA.n998 GNDA.n966 3.5845
R5457 GNDA.n997 GNDA.n994 3.5845
R5458 GNDA.n993 GNDA.n967 3.5845
R5459 GNDA.n990 GNDA.n989 3.5845
R5460 GNDA.n985 GNDA.n968 3.5845
R5461 GNDA.n984 GNDA.n981 3.5845
R5462 GNDA.n980 GNDA.n972 3.5845
R5463 GNDA.n977 GNDA.n976 3.5845
R5464 GNDA.n1053 GNDA.n701 3.5845
R5465 GNDA.n1200 GNDA.n1199 3.5845
R5466 GNDA.n1087 GNDA.n1085 3.5845
R5467 GNDA.n1194 GNDA.n1089 3.5845
R5468 GNDA.n1193 GNDA.n1090 3.5845
R5469 GNDA.n1189 GNDA.n1188 3.5845
R5470 GNDA.n1096 GNDA.n1094 3.5845
R5471 GNDA.n1183 GNDA.n1098 3.5845
R5472 GNDA.n1182 GNDA.n1099 3.5845
R5473 GNDA.n1178 GNDA.n1177 3.5845
R5474 GNDA.n1494 GNDA.n1419 3.5845
R5475 GNDA.n1493 GNDA.n1420 3.5845
R5476 GNDA.n1489 GNDA.n1488 3.5845
R5477 GNDA.n1462 GNDA.n1460 3.5845
R5478 GNDA.n1483 GNDA.n1464 3.5845
R5479 GNDA.n1482 GNDA.n1465 3.5845
R5480 GNDA.n1478 GNDA.n1477 3.5845
R5481 GNDA.n1473 GNDA.n1470 3.5845
R5482 GNDA.n1472 GNDA.n1401 3.5845
R5483 GNDA.n1391 GNDA.n1390 3.5845
R5484 GNDA.n1279 GNDA.n1277 3.5845
R5485 GNDA.n1385 GNDA.n1281 3.5845
R5486 GNDA.n1384 GNDA.n1282 3.5845
R5487 GNDA.n1380 GNDA.n1379 3.5845
R5488 GNDA.n1288 GNDA.n1286 3.5845
R5489 GNDA.n1374 GNDA.n1290 3.5845
R5490 GNDA.n1373 GNDA.n1291 3.5845
R5491 GNDA.n1369 GNDA.n1368 3.5845
R5492 GNDA.n2290 GNDA.n2289 3.5845
R5493 GNDA.n287 GNDA.n285 3.5845
R5494 GNDA.n2284 GNDA.n289 3.5845
R5495 GNDA.n2283 GNDA.n290 3.5845
R5496 GNDA.n2279 GNDA.n2278 3.5845
R5497 GNDA.n296 GNDA.n294 3.5845
R5498 GNDA.n2273 GNDA.n298 3.5845
R5499 GNDA.n2272 GNDA.n299 3.5845
R5500 GNDA.n2268 GNDA.n2267 3.5845
R5501 GNDA.n37 GNDA.t84 3.42907
R5502 GNDA.n37 GNDA.t93 3.42907
R5503 GNDA.n2483 GNDA.t322 3.42907
R5504 GNDA.n2483 GNDA.t345 3.42907
R5505 GNDA.n375 GNDA.t65 3.42907
R5506 GNDA.n375 GNDA.t29 3.42907
R5507 GNDA.n374 GNDA.t150 3.42907
R5508 GNDA.n374 GNDA.t113 3.42907
R5509 GNDA.n1855 GNDA.n610 3.3797
R5510 GNDA.n2064 GNDA.n2063 3.3797
R5511 GNDA.n2338 GNDA.n2337 3.3797
R5512 GNDA.n756 GNDA.n754 3.3797
R5513 GNDA.n965 GNDA.n964 3.3797
R5514 GNDA.n1204 GNDA.n1083 3.3797
R5515 GNDA.n1455 GNDA.n1417 3.3797
R5516 GNDA.n1395 GNDA.n659 3.3797
R5517 GNDA.n2294 GNDA.n283 3.3797
R5518 GNDA.n2435 GNDA.t335 3.28286
R5519 GNDA.n105 GNDA.n99 3.2005
R5520 GNDA.n316 GNDA.n315 3.2005
R5521 GNDA.n1825 GNDA.n1824 2.8677
R5522 GNDA.n2034 GNDA.n2033 2.8677
R5523 GNDA.n2447 GNDA.n2446 2.8677
R5524 GNDA.n785 GNDA.n775 2.8677
R5525 GNDA.n1055 GNDA.n1054 2.8677
R5526 GNDA.n1109 GNDA.n1103 2.8677
R5527 GNDA.n1550 GNDA.n1549 2.8677
R5528 GNDA.n1300 GNDA.n1295 2.8677
R5529 GNDA.n2199 GNDA.n303 2.8677
R5530 GNDA.n440 GNDA.t95 2.75116
R5531 GNDA.n409 GNDA.t317 2.75116
R5532 GNDA.n474 GNDA.t144 2.75116
R5533 GNDA.n1666 GNDA.n1664 2.34425
R5534 GNDA.n1674 GNDA.n1672 2.34425
R5535 GNDA.t142 GNDA.n62 2.33596
R5536 GNDA.n2465 GNDA.t78 2.33596
R5537 GNDA.n397 GNDA.t91 2.33596
R5538 GNDA.n396 GNDA.t154 2.33596
R5539 GNDA.n1549 GNDA.n1548 2.31161
R5540 GNDA.n1301 GNDA.n1300 2.31161
R5541 GNDA.n2200 GNDA.n2199 2.31161
R5542 GNDA.n786 GNDA.n785 2.31161
R5543 GNDA.n1055 GNDA.n699 2.31161
R5544 GNDA.n1110 GNDA.n1109 2.31161
R5545 GNDA.n1824 GNDA.n1817 2.31161
R5546 GNDA.n2033 GNDA.n2026 2.31161
R5547 GNDA.n2446 GNDA.n90 2.31161
R5548 GNDA GNDA.n1540 1.95606
R5549 GNDA.n1303 GNDA 1.95606
R5550 GNDA.n2202 GNDA 1.95606
R5551 GNDA.n788 GNDA 1.95606
R5552 GNDA.n704 GNDA 1.95606
R5553 GNDA.n1112 GNDA 1.95606
R5554 GNDA GNDA.n1809 1.95606
R5555 GNDA GNDA.n2018 1.95606
R5556 GNDA.n127 GNDA 1.95606
R5557 GNDA.n1824 GNDA.n1823 1.7413
R5558 GNDA.n2033 GNDA.n2032 1.7413
R5559 GNDA.n2446 GNDA.n2445 1.7413
R5560 GNDA.n785 GNDA.n784 1.7413
R5561 GNDA.n1211 GNDA.n1055 1.7413
R5562 GNDA.n1109 GNDA.n1108 1.7413
R5563 GNDA.n1549 GNDA.n1399 1.7413
R5564 GNDA.n1300 GNDA.n1299 1.7413
R5565 GNDA.n2199 GNDA.n2198 1.7413
R5566 GNDA.n561 GNDA.n560 1.73362
R5567 GNDA.n2175 GNDA.n312 1.64168
R5568 GNDA.n2495 GNDA.n25 1.6005
R5569 GNDA.n614 GNDA.n610 1.2293
R5570 GNDA.n2063 GNDA.n2062 1.2293
R5571 GNDA.n2337 GNDA.n141 1.2293
R5572 GNDA.n876 GNDA.n756 1.2293
R5573 GNDA.n966 GNDA.n965 1.2293
R5574 GNDA.n1200 GNDA.n1083 1.2293
R5575 GNDA.n1419 GNDA.n1417 1.2293
R5576 GNDA.n1391 GNDA.n659 1.2293
R5577 GNDA.n2290 GNDA.n283 1.2293
R5578 GNDA.n469 GNDA.n356 1.188
R5579 GNDA.n1822 GNDA.n1818 1.1781
R5580 GNDA.n2031 GNDA.n2028 1.1781
R5581 GNDA.n2444 GNDA.n91 1.1781
R5582 GNDA.n779 GNDA.n777 1.1781
R5583 GNDA.n1210 GNDA.n1209 1.1781
R5584 GNDA.n2152 GNDA.n525 1.1781
R5585 GNDA.n1556 GNDA.n1555 1.1781
R5586 GNDA.n2299 GNDA.n208 1.1781
R5587 GNDA.n310 GNDA.n305 1.1781
R5588 GNDA.n2080 GNDA.n552 1.16414
R5589 GNDA.n1849 GNDA.n615 1.0245
R5590 GNDA.n1848 GNDA.n616 1.0245
R5591 GNDA.n1844 GNDA.n1843 1.0245
R5592 GNDA.n1607 GNDA.n619 1.0245
R5593 GNDA.n1837 GNDA.n1608 1.0245
R5594 GNDA.n1836 GNDA.n1609 1.0245
R5595 GNDA.n1832 GNDA.n1831 1.0245
R5596 GNDA.n1747 GNDA.n1613 1.0245
R5597 GNDA.n1825 GNDA.n1748 1.0245
R5598 GNDA.n2061 GNDA.n1938 1.0245
R5599 GNDA.n1942 GNDA.n1940 1.0245
R5600 GNDA.n2056 GNDA.n2055 1.0245
R5601 GNDA.n2047 GNDA.n1943 1.0245
R5602 GNDA.n2046 GNDA.n1946 1.0245
R5603 GNDA.n1950 GNDA.n1948 1.0245
R5604 GNDA.n2041 GNDA.n2040 1.0245
R5605 GNDA.n1958 GNDA.n1951 1.0245
R5606 GNDA.n2034 GNDA.n1959 1.0245
R5607 GNDA.n2357 GNDA.n2356 1.0245
R5608 GNDA.n2342 GNDA.n142 1.0245
R5609 GNDA.n2350 GNDA.n2343 1.0245
R5610 GNDA.n2349 GNDA.n2344 1.0245
R5611 GNDA.n2424 GNDA.n123 1.0245
R5612 GNDA.n2423 GNDA.n124 1.0245
R5613 GNDA.n2419 GNDA.n2418 1.0245
R5614 GNDA.n2415 GNDA.n2414 1.0245
R5615 GNDA.n2447 GNDA.n89 1.0245
R5616 GNDA.n875 GNDA.n757 1.0245
R5617 GNDA.n761 GNDA.n759 1.0245
R5618 GNDA.n870 GNDA.n869 1.0245
R5619 GNDA.n865 GNDA.n762 1.0245
R5620 GNDA.n864 GNDA.n766 1.0245
R5621 GNDA.n770 GNDA.n768 1.0245
R5622 GNDA.n859 GNDA.n858 1.0245
R5623 GNDA.n854 GNDA.n771 1.0245
R5624 GNDA.n853 GNDA.n775 1.0245
R5625 GNDA.n998 GNDA.n997 1.0245
R5626 GNDA.n994 GNDA.n993 1.0245
R5627 GNDA.n990 GNDA.n967 1.0245
R5628 GNDA.n989 GNDA.n968 1.0245
R5629 GNDA.n985 GNDA.n984 1.0245
R5630 GNDA.n981 GNDA.n980 1.0245
R5631 GNDA.n977 GNDA.n972 1.0245
R5632 GNDA.n976 GNDA.n701 1.0245
R5633 GNDA.n1054 GNDA.n1053 1.0245
R5634 GNDA.n1199 GNDA.n1085 1.0245
R5635 GNDA.n1089 GNDA.n1087 1.0245
R5636 GNDA.n1194 GNDA.n1193 1.0245
R5637 GNDA.n1189 GNDA.n1090 1.0245
R5638 GNDA.n1188 GNDA.n1094 1.0245
R5639 GNDA.n1098 GNDA.n1096 1.0245
R5640 GNDA.n1183 GNDA.n1182 1.0245
R5641 GNDA.n1178 GNDA.n1099 1.0245
R5642 GNDA.n1177 GNDA.n1103 1.0245
R5643 GNDA.n1494 GNDA.n1493 1.0245
R5644 GNDA.n1489 GNDA.n1420 1.0245
R5645 GNDA.n1488 GNDA.n1460 1.0245
R5646 GNDA.n1464 GNDA.n1462 1.0245
R5647 GNDA.n1483 GNDA.n1482 1.0245
R5648 GNDA.n1478 GNDA.n1465 1.0245
R5649 GNDA.n1477 GNDA.n1470 1.0245
R5650 GNDA.n1473 GNDA.n1472 1.0245
R5651 GNDA.n1550 GNDA.n1401 1.0245
R5652 GNDA.n1390 GNDA.n1277 1.0245
R5653 GNDA.n1281 GNDA.n1279 1.0245
R5654 GNDA.n1385 GNDA.n1384 1.0245
R5655 GNDA.n1380 GNDA.n1282 1.0245
R5656 GNDA.n1379 GNDA.n1286 1.0245
R5657 GNDA.n1290 GNDA.n1288 1.0245
R5658 GNDA.n1374 GNDA.n1373 1.0245
R5659 GNDA.n1369 GNDA.n1291 1.0245
R5660 GNDA.n1368 GNDA.n1295 1.0245
R5661 GNDA.n2289 GNDA.n285 1.0245
R5662 GNDA.n289 GNDA.n287 1.0245
R5663 GNDA.n2284 GNDA.n2283 1.0245
R5664 GNDA.n2279 GNDA.n290 1.0245
R5665 GNDA.n2278 GNDA.n294 1.0245
R5666 GNDA.n298 GNDA.n296 1.0245
R5667 GNDA.n2273 GNDA.n2272 1.0245
R5668 GNDA.n2268 GNDA.n299 1.0245
R5669 GNDA.n2267 GNDA.n303 1.0245
R5670 GNDA.n433 GNDA.n432 0.59425
R5671 GNDA.n1664 GNDA.n1662 0.563
R5672 GNDA.n1668 GNDA.n1666 0.563
R5673 GNDA.n1670 GNDA.n1668 0.563
R5674 GNDA.n1672 GNDA.n1670 0.563
R5675 GNDA.n1676 GNDA.n1674 0.563
R5676 GNDA.n1678 GNDA.n1676 0.563
R5677 GNDA.n353 GNDA.n352 0.563
R5678 GNDA.n353 GNDA.n349 0.563
R5679 GNDA.n17 GNDA.n15 0.563
R5680 GNDA.n19 GNDA.n17 0.563
R5681 GNDA.n21 GNDA.n19 0.563
R5682 GNDA.n23 GNDA.n21 0.563
R5683 GNDA.n414 GNDA.n36 0.563
R5684 GNDA.n416 GNDA.n414 0.563
R5685 GNDA.n418 GNDA.n416 0.563
R5686 GNDA.n420 GNDA.n418 0.563
R5687 GNDA.n422 GNDA.n420 0.563
R5688 GNDA.n424 GNDA.n422 0.563
R5689 GNDA.n426 GNDA.n424 0.563
R5690 GNDA.n428 GNDA.n426 0.563
R5691 GNDA.n430 GNDA.n428 0.563
R5692 GNDA.n432 GNDA.n430 0.563
R5693 GNDA.n6 GNDA.n4 0.563
R5694 GNDA.n8 GNDA.n6 0.563
R5695 GNDA.n10 GNDA.n8 0.563
R5696 GNDA.n12 GNDA.n10 0.563
R5697 GNDA.n2498 GNDA.n1 0.53175
R5698 GNDA.n377 GNDA.n376 0.5005
R5699 GNDA.n2484 GNDA.n2482 0.5005
R5700 GNDA.n2464 GNDA.t2 0.467591
R5701 GNDA.n389 GNDA.t63 0.467591
R5702 GNDA.n558 GNDA.n557 0.41175
R5703 GNDA.n559 GNDA.n558 0.311875
R5704 GNDA.n2486 GNDA.n36 0.28175
R5705 GNDA.n1659 GNDA.n1640 0.276625
R5706 GNDA.n356 GNDA.n355 0.2505
R5707 GNDA.n1679 GNDA.n1659 0.22375
R5708 GNDA GNDA.n2429 0.129793
R5709 GNDA.n2144 GNDA 0.129793
R5710 GNDA.n2172 GNDA 0.129793
R5711 GNDA.n1680 GNDA.n1679 0.100375
R5712 GNDA.n560 GNDA.n559 0.076875
R5713 GNDA.n1222 GNDA.n257 0.0479074
R5714 GNDA.n1237 GNDA 0.0479074
R5715 GNDA.n656 GNDA.n587 0.0479074
R5716 GNDA.n1925 GNDA 0.0479074
R5717 GNDA.n635 GNDA.n634 0.0479074
R5718 GNDA GNDA.n648 0.0479074
R5719 GNDA.n732 GNDA.n730 0.0479074
R5720 GNDA.n951 GNDA 0.0479074
R5721 GNDA.n548 GNDA.n544 0.0479074
R5722 GNDA GNDA.n1073 0.0479074
R5723 GNDA.n183 GNDA.n182 0.0479074
R5724 GNDA GNDA.n273 0.0479074
R5725 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.t15 354.854
R5726 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.t30 346.8
R5727 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n4 339.522
R5728 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n11 339.522
R5729 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n9 335.022
R5730 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.t2 275.909
R5731 bgr_0.1st_Vout_1.n7 bgr_0.1st_Vout_1.n6 227.909
R5732 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n8 222.034
R5733 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t31 184.097
R5734 bgr_0.1st_Vout_1.n5 bgr_0.1st_Vout_1.t14 184.097
R5735 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t27 184.097
R5736 bgr_0.1st_Vout_1.n10 bgr_0.1st_Vout_1.t19 184.097
R5737 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n5 166.05
R5738 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n10 166.05
R5739 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t5 48.0005
R5740 bgr_0.1st_Vout_1.n8 bgr_0.1st_Vout_1.t7 48.0005
R5741 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t10 48.0005
R5742 bgr_0.1st_Vout_1.n6 bgr_0.1st_Vout_1.t3 48.0005
R5743 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t8 39.4005
R5744 bgr_0.1st_Vout_1.n9 bgr_0.1st_Vout_1.t1 39.4005
R5745 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t9 39.4005
R5746 bgr_0.1st_Vout_1.n11 bgr_0.1st_Vout_1.t6 39.4005
R5747 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t4 39.4005
R5748 bgr_0.1st_Vout_1.n4 bgr_0.1st_Vout_1.t0 39.4005
R5749 bgr_0.1st_Vout_1.n0 bgr_0.1st_Vout_1.n2 33.1711
R5750 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n0 5.6255
R5751 bgr_0.1st_Vout_1 bgr_0.1st_Vout_1.n3 5.28175
R5752 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t20 4.8295
R5753 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t29 4.8295
R5754 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t25 4.8295
R5755 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t35 4.8295
R5756 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t33 4.8295
R5757 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t17 4.8295
R5758 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t28 4.8295
R5759 bgr_0.1st_Vout_1.n3 bgr_0.1st_Vout_1.n7 4.5005
R5760 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t11 4.5005
R5761 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t32 4.5005
R5762 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t34 4.5005
R5763 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t21 4.5005
R5764 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t12 4.5005
R5765 bgr_0.1st_Vout_1.n1 bgr_0.1st_Vout_1.t16 4.5005
R5766 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t26 4.5005
R5767 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t22 4.5005
R5768 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t24 4.5005
R5769 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t23 4.5005
R5770 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t13 4.5005
R5771 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t18 4.5005
R5772 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.t36 4.5005
R5773 bgr_0.1st_Vout_1.n2 bgr_0.1st_Vout_1.n1 3.8075
R5774 bgr_0.cap_res1.t0 bgr_0.cap_res1.t18 178.633
R5775 bgr_0.cap_res1.t15 bgr_0.cap_res1.t1 0.1603
R5776 bgr_0.cap_res1.t11 bgr_0.cap_res1.t7 0.1603
R5777 bgr_0.cap_res1.t10 bgr_0.cap_res1.t16 0.1603
R5778 bgr_0.cap_res1.t8 bgr_0.cap_res1.t4 0.1603
R5779 bgr_0.cap_res1.t17 bgr_0.cap_res1.t2 0.1603
R5780 bgr_0.cap_res1.t13 bgr_0.cap_res1.t9 0.1603
R5781 bgr_0.cap_res1.t3 bgr_0.cap_res1.t6 0.1603
R5782 bgr_0.cap_res1.t20 bgr_0.cap_res1.t14 0.1603
R5783 bgr_0.cap_res1.n1 bgr_0.cap_res1.t5 0.159278
R5784 bgr_0.cap_res1.n2 bgr_0.cap_res1.t19 0.159278
R5785 bgr_0.cap_res1.n3 bgr_0.cap_res1.t12 0.159278
R5786 bgr_0.cap_res1.n3 bgr_0.cap_res1.t15 0.1368
R5787 bgr_0.cap_res1.n3 bgr_0.cap_res1.t11 0.1368
R5788 bgr_0.cap_res1.n2 bgr_0.cap_res1.t10 0.1368
R5789 bgr_0.cap_res1.n2 bgr_0.cap_res1.t8 0.1368
R5790 bgr_0.cap_res1.n1 bgr_0.cap_res1.t17 0.1368
R5791 bgr_0.cap_res1.n1 bgr_0.cap_res1.t13 0.1368
R5792 bgr_0.cap_res1.n0 bgr_0.cap_res1.t3 0.1368
R5793 bgr_0.cap_res1.n0 bgr_0.cap_res1.t20 0.1368
R5794 bgr_0.cap_res1.t5 bgr_0.cap_res1.n0 0.00152174
R5795 bgr_0.cap_res1.t19 bgr_0.cap_res1.n1 0.00152174
R5796 bgr_0.cap_res1.t12 bgr_0.cap_res1.n2 0.00152174
R5797 bgr_0.cap_res1.t18 bgr_0.cap_res1.n3 0.00152174
R5798 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.n7 114.719
R5799 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n6 114.719
R5800 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n10 114.156
R5801 two_stage_opamp_dummy_magic_0.VD2.n9 two_stage_opamp_dummy_magic_0.VD2.n8 114.156
R5802 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n0 112.456
R5803 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.n18 112.454
R5804 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n17 111.206
R5805 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n3 111.206
R5806 two_stage_opamp_dummy_magic_0.VD2.n2 two_stage_opamp_dummy_magic_0.VD2.n1 111.206
R5807 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n5 109.656
R5808 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n14 106.706
R5809 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t13 16.0005
R5810 two_stage_opamp_dummy_magic_0.VD2.n17 two_stage_opamp_dummy_magic_0.VD2.t19 16.0005
R5811 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t11 16.0005
R5812 two_stage_opamp_dummy_magic_0.VD2.n10 two_stage_opamp_dummy_magic_0.VD2.t10 16.0005
R5813 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.t8 16.0005
R5814 two_stage_opamp_dummy_magic_0.VD2.n8 two_stage_opamp_dummy_magic_0.VD2.t5 16.0005
R5815 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t9 16.0005
R5816 two_stage_opamp_dummy_magic_0.VD2.n7 two_stage_opamp_dummy_magic_0.VD2.t14 16.0005
R5817 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t3 16.0005
R5818 two_stage_opamp_dummy_magic_0.VD2.n6 two_stage_opamp_dummy_magic_0.VD2.t1 16.0005
R5819 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t20 16.0005
R5820 two_stage_opamp_dummy_magic_0.VD2.n5 two_stage_opamp_dummy_magic_0.VD2.t21 16.0005
R5821 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t0 16.0005
R5822 two_stage_opamp_dummy_magic_0.VD2.n14 two_stage_opamp_dummy_magic_0.VD2.t15 16.0005
R5823 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t7 16.0005
R5824 two_stage_opamp_dummy_magic_0.VD2.n3 two_stage_opamp_dummy_magic_0.VD2.t16 16.0005
R5825 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t6 16.0005
R5826 two_stage_opamp_dummy_magic_0.VD2.n1 two_stage_opamp_dummy_magic_0.VD2.t2 16.0005
R5827 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t4 16.0005
R5828 two_stage_opamp_dummy_magic_0.VD2.n0 two_stage_opamp_dummy_magic_0.VD2.t18 16.0005
R5829 two_stage_opamp_dummy_magic_0.VD2.n19 two_stage_opamp_dummy_magic_0.VD2.t12 16.0005
R5830 two_stage_opamp_dummy_magic_0.VD2.t17 two_stage_opamp_dummy_magic_0.VD2.n19 16.0005
R5831 two_stage_opamp_dummy_magic_0.VD2.n13 two_stage_opamp_dummy_magic_0.VD2.n12 4.5005
R5832 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n15 4.5005
R5833 two_stage_opamp_dummy_magic_0.VD2.n16 two_stage_opamp_dummy_magic_0.VD2.n4 3.6255
R5834 two_stage_opamp_dummy_magic_0.VD2.n4 two_stage_opamp_dummy_magic_0.VD2.n2 1.2505
R5835 two_stage_opamp_dummy_magic_0.VD2.n18 two_stage_opamp_dummy_magic_0.VD2.n16 1.2505
R5836 two_stage_opamp_dummy_magic_0.VD2.n15 two_stage_opamp_dummy_magic_0.VD2.n13 0.78175
R5837 two_stage_opamp_dummy_magic_0.VD2.n11 two_stage_opamp_dummy_magic_0.VD2.n9 0.563
R5838 two_stage_opamp_dummy_magic_0.VD2.n12 two_stage_opamp_dummy_magic_0.VD2.n11 0.563
R5839 two_stage_opamp_dummy_magic_0.VOUT+.n13 two_stage_opamp_dummy_magic_0.VOUT+.n5 145.989
R5840 two_stage_opamp_dummy_magic_0.VOUT+.n8 two_stage_opamp_dummy_magic_0.VOUT+.n6 145.989
R5841 two_stage_opamp_dummy_magic_0.VOUT+.n12 two_stage_opamp_dummy_magic_0.VOUT+.n11 145.427
R5842 two_stage_opamp_dummy_magic_0.VOUT+.n10 two_stage_opamp_dummy_magic_0.VOUT+.n9 145.427
R5843 two_stage_opamp_dummy_magic_0.VOUT+.n8 two_stage_opamp_dummy_magic_0.VOUT+.n7 145.427
R5844 two_stage_opamp_dummy_magic_0.VOUT+.n15 two_stage_opamp_dummy_magic_0.VOUT+.n14 140.927
R5845 two_stage_opamp_dummy_magic_0.VOUT+.t17 two_stage_opamp_dummy_magic_0.VOUT+.n96 113.192
R5846 two_stage_opamp_dummy_magic_0.VOUT+.n2 two_stage_opamp_dummy_magic_0.VOUT+.n0 95.7303
R5847 two_stage_opamp_dummy_magic_0.VOUT+.n4 two_stage_opamp_dummy_magic_0.VOUT+.n3 94.6053
R5848 two_stage_opamp_dummy_magic_0.VOUT+.n2 two_stage_opamp_dummy_magic_0.VOUT+.n1 94.6053
R5849 two_stage_opamp_dummy_magic_0.VOUT+.n95 two_stage_opamp_dummy_magic_0.VOUT+.n15 20.688
R5850 two_stage_opamp_dummy_magic_0.VOUT+.n95 two_stage_opamp_dummy_magic_0.VOUT+.n94 11.7059
R5851 two_stage_opamp_dummy_magic_0.VOUT+.n96 two_stage_opamp_dummy_magic_0.VOUT+.n95 11.063
R5852 two_stage_opamp_dummy_magic_0.VOUT+.n14 two_stage_opamp_dummy_magic_0.VOUT+.t11 6.56717
R5853 two_stage_opamp_dummy_magic_0.VOUT+.n14 two_stage_opamp_dummy_magic_0.VOUT+.t6 6.56717
R5854 two_stage_opamp_dummy_magic_0.VOUT+.n11 two_stage_opamp_dummy_magic_0.VOUT+.t1 6.56717
R5855 two_stage_opamp_dummy_magic_0.VOUT+.n11 two_stage_opamp_dummy_magic_0.VOUT+.t2 6.56717
R5856 two_stage_opamp_dummy_magic_0.VOUT+.n9 two_stage_opamp_dummy_magic_0.VOUT+.t10 6.56717
R5857 two_stage_opamp_dummy_magic_0.VOUT+.n9 two_stage_opamp_dummy_magic_0.VOUT+.t9 6.56717
R5858 two_stage_opamp_dummy_magic_0.VOUT+.n7 two_stage_opamp_dummy_magic_0.VOUT+.t5 6.56717
R5859 two_stage_opamp_dummy_magic_0.VOUT+.n7 two_stage_opamp_dummy_magic_0.VOUT+.t0 6.56717
R5860 two_stage_opamp_dummy_magic_0.VOUT+.n6 two_stage_opamp_dummy_magic_0.VOUT+.t8 6.56717
R5861 two_stage_opamp_dummy_magic_0.VOUT+.n6 two_stage_opamp_dummy_magic_0.VOUT+.t13 6.56717
R5862 two_stage_opamp_dummy_magic_0.VOUT+.n5 two_stage_opamp_dummy_magic_0.VOUT+.t12 6.56717
R5863 two_stage_opamp_dummy_magic_0.VOUT+.n5 two_stage_opamp_dummy_magic_0.VOUT+.t7 6.56717
R5864 two_stage_opamp_dummy_magic_0.VOUT+.n42 two_stage_opamp_dummy_magic_0.VOUT+.t85 4.8295
R5865 two_stage_opamp_dummy_magic_0.VOUT+.n44 two_stage_opamp_dummy_magic_0.VOUT+.t131 4.8295
R5866 two_stage_opamp_dummy_magic_0.VOUT+.n46 two_stage_opamp_dummy_magic_0.VOUT+.t31 4.8295
R5867 two_stage_opamp_dummy_magic_0.VOUT+.n48 two_stage_opamp_dummy_magic_0.VOUT+.t62 4.8295
R5868 two_stage_opamp_dummy_magic_0.VOUT+.n50 two_stage_opamp_dummy_magic_0.VOUT+.t114 4.8295
R5869 two_stage_opamp_dummy_magic_0.VOUT+.n62 two_stage_opamp_dummy_magic_0.VOUT+.t40 4.8295
R5870 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.t34 4.8295
R5871 two_stage_opamp_dummy_magic_0.VOUT+.n65 two_stage_opamp_dummy_magic_0.VOUT+.t136 4.8295
R5872 two_stage_opamp_dummy_magic_0.VOUT+.n67 two_stage_opamp_dummy_magic_0.VOUT+.t70 4.8295
R5873 two_stage_opamp_dummy_magic_0.VOUT+.n68 two_stage_opamp_dummy_magic_0.VOUT+.t36 4.8295
R5874 two_stage_opamp_dummy_magic_0.VOUT+.n70 two_stage_opamp_dummy_magic_0.VOUT+.t95 4.8295
R5875 two_stage_opamp_dummy_magic_0.VOUT+.n71 two_stage_opamp_dummy_magic_0.VOUT+.t66 4.8295
R5876 two_stage_opamp_dummy_magic_0.VOUT+.n73 two_stage_opamp_dummy_magic_0.VOUT+.t55 4.8295
R5877 two_stage_opamp_dummy_magic_0.VOUT+.n74 two_stage_opamp_dummy_magic_0.VOUT+.t29 4.8295
R5878 two_stage_opamp_dummy_magic_0.VOUT+.n76 two_stage_opamp_dummy_magic_0.VOUT+.t91 4.8295
R5879 two_stage_opamp_dummy_magic_0.VOUT+.n77 two_stage_opamp_dummy_magic_0.VOUT+.t58 4.8295
R5880 two_stage_opamp_dummy_magic_0.VOUT+.n79 two_stage_opamp_dummy_magic_0.VOUT+.t49 4.8295
R5881 two_stage_opamp_dummy_magic_0.VOUT+.n80 two_stage_opamp_dummy_magic_0.VOUT+.t20 4.8295
R5882 two_stage_opamp_dummy_magic_0.VOUT+.n82 two_stage_opamp_dummy_magic_0.VOUT+.t148 4.8295
R5883 two_stage_opamp_dummy_magic_0.VOUT+.n83 two_stage_opamp_dummy_magic_0.VOUT+.t122 4.8295
R5884 two_stage_opamp_dummy_magic_0.VOUT+.n85 two_stage_opamp_dummy_magic_0.VOUT+.t44 4.8295
R5885 two_stage_opamp_dummy_magic_0.VOUT+.n86 two_stage_opamp_dummy_magic_0.VOUT+.t152 4.8295
R5886 two_stage_opamp_dummy_magic_0.VOUT+.n88 two_stage_opamp_dummy_magic_0.VOUT+.t142 4.8295
R5887 two_stage_opamp_dummy_magic_0.VOUT+.n89 two_stage_opamp_dummy_magic_0.VOUT+.t116 4.8295
R5888 two_stage_opamp_dummy_magic_0.VOUT+.n16 two_stage_opamp_dummy_magic_0.VOUT+.t108 4.8295
R5889 two_stage_opamp_dummy_magic_0.VOUT+.n28 two_stage_opamp_dummy_magic_0.VOUT+.t28 4.8295
R5890 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.t24 4.8295
R5891 two_stage_opamp_dummy_magic_0.VOUT+.n31 two_stage_opamp_dummy_magic_0.VOUT+.t129 4.8295
R5892 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.t61 4.8295
R5893 two_stage_opamp_dummy_magic_0.VOUT+.n34 two_stage_opamp_dummy_magic_0.VOUT+.t32 4.8295
R5894 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.t100 4.8295
R5895 two_stage_opamp_dummy_magic_0.VOUT+.n37 two_stage_opamp_dummy_magic_0.VOUT+.t71 4.8295
R5896 two_stage_opamp_dummy_magic_0.VOUT+.n39 two_stage_opamp_dummy_magic_0.VOUT+.t69 4.8295
R5897 two_stage_opamp_dummy_magic_0.VOUT+.n40 two_stage_opamp_dummy_magic_0.VOUT+.t35 4.8295
R5898 two_stage_opamp_dummy_magic_0.VOUT+.n91 two_stage_opamp_dummy_magic_0.VOUT+.t77 4.8295
R5899 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.t26 4.8154
R5900 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.t59 4.8154
R5901 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.t37 4.8154
R5902 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.t81 4.8154
R5903 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.t132 4.806
R5904 two_stage_opamp_dummy_magic_0.VOUT+.n60 two_stage_opamp_dummy_magic_0.VOUT+.t115 4.806
R5905 two_stage_opamp_dummy_magic_0.VOUT+.n59 two_stage_opamp_dummy_magic_0.VOUT+.t146 4.806
R5906 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.t46 4.806
R5907 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.t87 4.806
R5908 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.t65 4.806
R5909 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.t102 4.806
R5910 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.t134 4.806
R5911 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.t120 4.806
R5912 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.t155 4.806
R5913 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.t48 4.806
R5914 two_stage_opamp_dummy_magic_0.VOUT+.n26 two_stage_opamp_dummy_magic_0.VOUT+.t92 4.806
R5915 two_stage_opamp_dummy_magic_0.VOUT+.n25 two_stage_opamp_dummy_magic_0.VOUT+.t42 4.806
R5916 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.t130 4.806
R5917 two_stage_opamp_dummy_magic_0.VOUT+.n23 two_stage_opamp_dummy_magic_0.VOUT+.t84 4.806
R5918 two_stage_opamp_dummy_magic_0.VOUT+.n22 two_stage_opamp_dummy_magic_0.VOUT+.t125 4.806
R5919 two_stage_opamp_dummy_magic_0.VOUT+.n21 two_stage_opamp_dummy_magic_0.VOUT+.t74 4.806
R5920 two_stage_opamp_dummy_magic_0.VOUT+.n20 two_stage_opamp_dummy_magic_0.VOUT+.t23 4.806
R5921 two_stage_opamp_dummy_magic_0.VOUT+.n19 two_stage_opamp_dummy_magic_0.VOUT+.t64 4.806
R5922 two_stage_opamp_dummy_magic_0.VOUT+.n18 two_stage_opamp_dummy_magic_0.VOUT+.t150 4.806
R5923 two_stage_opamp_dummy_magic_0.VOUT+.n43 two_stage_opamp_dummy_magic_0.VOUT+.t96 4.5005
R5924 two_stage_opamp_dummy_magic_0.VOUT+.n42 two_stage_opamp_dummy_magic_0.VOUT+.t57 4.5005
R5925 two_stage_opamp_dummy_magic_0.VOUT+.n44 two_stage_opamp_dummy_magic_0.VOUT+.t104 4.5005
R5926 two_stage_opamp_dummy_magic_0.VOUT+.n45 two_stage_opamp_dummy_magic_0.VOUT+.t73 4.5005
R5927 two_stage_opamp_dummy_magic_0.VOUT+.n46 two_stage_opamp_dummy_magic_0.VOUT+.t138 4.5005
R5928 two_stage_opamp_dummy_magic_0.VOUT+.n47 two_stage_opamp_dummy_magic_0.VOUT+.t107 4.5005
R5929 two_stage_opamp_dummy_magic_0.VOUT+.n48 two_stage_opamp_dummy_magic_0.VOUT+.t41 4.5005
R5930 two_stage_opamp_dummy_magic_0.VOUT+.n49 two_stage_opamp_dummy_magic_0.VOUT+.t143 4.5005
R5931 two_stage_opamp_dummy_magic_0.VOUT+.n50 two_stage_opamp_dummy_magic_0.VOUT+.t21 4.5005
R5932 two_stage_opamp_dummy_magic_0.VOUT+.n51 two_stage_opamp_dummy_magic_0.VOUT+.t126 4.5005
R5933 two_stage_opamp_dummy_magic_0.VOUT+.n52 two_stage_opamp_dummy_magic_0.VOUT+.t119 4.5005
R5934 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.t82 4.5005
R5935 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.t97 4.5005
R5936 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.t63 4.5005
R5937 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.t27 4.5005
R5938 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.t45 4.5005
R5939 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.t144 4.5005
R5940 two_stage_opamp_dummy_magic_0.VOUT+.n59 two_stage_opamp_dummy_magic_0.VOUT+.t112 4.5005
R5941 two_stage_opamp_dummy_magic_0.VOUT+.n60 two_stage_opamp_dummy_magic_0.VOUT+.t76 4.5005
R5942 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.t93 4.5005
R5943 two_stage_opamp_dummy_magic_0.VOUT+.n63 two_stage_opamp_dummy_magic_0.VOUT+.t56 4.5005
R5944 two_stage_opamp_dummy_magic_0.VOUT+.n62 two_stage_opamp_dummy_magic_0.VOUT+.t19 4.5005
R5945 two_stage_opamp_dummy_magic_0.VOUT+.n64 two_stage_opamp_dummy_magic_0.VOUT+.t52 4.5005
R5946 two_stage_opamp_dummy_magic_0.VOUT+.n66 two_stage_opamp_dummy_magic_0.VOUT+.t156 4.5005
R5947 two_stage_opamp_dummy_magic_0.VOUT+.n65 two_stage_opamp_dummy_magic_0.VOUT+.t121 4.5005
R5948 two_stage_opamp_dummy_magic_0.VOUT+.n67 two_stage_opamp_dummy_magic_0.VOUT+.t89 4.5005
R5949 two_stage_opamp_dummy_magic_0.VOUT+.n69 two_stage_opamp_dummy_magic_0.VOUT+.t50 4.5005
R5950 two_stage_opamp_dummy_magic_0.VOUT+.n68 two_stage_opamp_dummy_magic_0.VOUT+.t151 4.5005
R5951 two_stage_opamp_dummy_magic_0.VOUT+.n70 two_stage_opamp_dummy_magic_0.VOUT+.t43 4.5005
R5952 two_stage_opamp_dummy_magic_0.VOUT+.n72 two_stage_opamp_dummy_magic_0.VOUT+.t145 4.5005
R5953 two_stage_opamp_dummy_magic_0.VOUT+.n71 two_stage_opamp_dummy_magic_0.VOUT+.t118 4.5005
R5954 two_stage_opamp_dummy_magic_0.VOUT+.n73 two_stage_opamp_dummy_magic_0.VOUT+.t141 4.5005
R5955 two_stage_opamp_dummy_magic_0.VOUT+.n75 two_stage_opamp_dummy_magic_0.VOUT+.t111 4.5005
R5956 two_stage_opamp_dummy_magic_0.VOUT+.n74 two_stage_opamp_dummy_magic_0.VOUT+.t80 4.5005
R5957 two_stage_opamp_dummy_magic_0.VOUT+.n76 two_stage_opamp_dummy_magic_0.VOUT+.t39 4.5005
R5958 two_stage_opamp_dummy_magic_0.VOUT+.n78 two_stage_opamp_dummy_magic_0.VOUT+.t139 4.5005
R5959 two_stage_opamp_dummy_magic_0.VOUT+.n77 two_stage_opamp_dummy_magic_0.VOUT+.t109 4.5005
R5960 two_stage_opamp_dummy_magic_0.VOUT+.n79 two_stage_opamp_dummy_magic_0.VOUT+.t135 4.5005
R5961 two_stage_opamp_dummy_magic_0.VOUT+.n81 two_stage_opamp_dummy_magic_0.VOUT+.t103 4.5005
R5962 two_stage_opamp_dummy_magic_0.VOUT+.n80 two_stage_opamp_dummy_magic_0.VOUT+.t72 4.5005
R5963 two_stage_opamp_dummy_magic_0.VOUT+.n82 two_stage_opamp_dummy_magic_0.VOUT+.t99 4.5005
R5964 two_stage_opamp_dummy_magic_0.VOUT+.n84 two_stage_opamp_dummy_magic_0.VOUT+.t68 4.5005
R5965 two_stage_opamp_dummy_magic_0.VOUT+.n83 two_stage_opamp_dummy_magic_0.VOUT+.t33 4.5005
R5966 two_stage_opamp_dummy_magic_0.VOUT+.n85 two_stage_opamp_dummy_magic_0.VOUT+.t133 4.5005
R5967 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.t98 4.5005
R5968 two_stage_opamp_dummy_magic_0.VOUT+.n86 two_stage_opamp_dummy_magic_0.VOUT+.t67 4.5005
R5969 two_stage_opamp_dummy_magic_0.VOUT+.n88 two_stage_opamp_dummy_magic_0.VOUT+.t94 4.5005
R5970 two_stage_opamp_dummy_magic_0.VOUT+.n90 two_stage_opamp_dummy_magic_0.VOUT+.t60 4.5005
R5971 two_stage_opamp_dummy_magic_0.VOUT+.n89 two_stage_opamp_dummy_magic_0.VOUT+.t30 4.5005
R5972 two_stage_opamp_dummy_magic_0.VOUT+.n17 two_stage_opamp_dummy_magic_0.VOUT+.t101 4.5005
R5973 two_stage_opamp_dummy_magic_0.VOUT+.n16 two_stage_opamp_dummy_magic_0.VOUT+.t149 4.5005
R5974 two_stage_opamp_dummy_magic_0.VOUT+.n18 two_stage_opamp_dummy_magic_0.VOUT+.t88 4.5005
R5975 two_stage_opamp_dummy_magic_0.VOUT+.n19 two_stage_opamp_dummy_magic_0.VOUT+.t51 4.5005
R5976 two_stage_opamp_dummy_magic_0.VOUT+.n20 two_stage_opamp_dummy_magic_0.VOUT+.t137 4.5005
R5977 two_stage_opamp_dummy_magic_0.VOUT+.n21 two_stage_opamp_dummy_magic_0.VOUT+.t106 4.5005
R5978 two_stage_opamp_dummy_magic_0.VOUT+.n22 two_stage_opamp_dummy_magic_0.VOUT+.t75 4.5005
R5979 two_stage_opamp_dummy_magic_0.VOUT+.n23 two_stage_opamp_dummy_magic_0.VOUT+.t25 4.5005
R5980 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.t128 4.5005
R5981 two_stage_opamp_dummy_magic_0.VOUT+.n25 two_stage_opamp_dummy_magic_0.VOUT+.t90 4.5005
R5982 two_stage_opamp_dummy_magic_0.VOUT+.n26 two_stage_opamp_dummy_magic_0.VOUT+.t54 4.5005
R5983 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.t140 4.5005
R5984 two_stage_opamp_dummy_magic_0.VOUT+.n29 two_stage_opamp_dummy_magic_0.VOUT+.t110 4.5005
R5985 two_stage_opamp_dummy_magic_0.VOUT+.n28 two_stage_opamp_dummy_magic_0.VOUT+.t79 4.5005
R5986 two_stage_opamp_dummy_magic_0.VOUT+.n30 two_stage_opamp_dummy_magic_0.VOUT+.t113 4.5005
R5987 two_stage_opamp_dummy_magic_0.VOUT+.n32 two_stage_opamp_dummy_magic_0.VOUT+.t78 4.5005
R5988 two_stage_opamp_dummy_magic_0.VOUT+.n31 two_stage_opamp_dummy_magic_0.VOUT+.t38 4.5005
R5989 two_stage_opamp_dummy_magic_0.VOUT+.n33 two_stage_opamp_dummy_magic_0.VOUT+.t147 4.5005
R5990 two_stage_opamp_dummy_magic_0.VOUT+.n35 two_stage_opamp_dummy_magic_0.VOUT+.t117 4.5005
R5991 two_stage_opamp_dummy_magic_0.VOUT+.n34 two_stage_opamp_dummy_magic_0.VOUT+.t83 4.5005
R5992 two_stage_opamp_dummy_magic_0.VOUT+.n36 two_stage_opamp_dummy_magic_0.VOUT+.t47 4.5005
R5993 two_stage_opamp_dummy_magic_0.VOUT+.n38 two_stage_opamp_dummy_magic_0.VOUT+.t153 4.5005
R5994 two_stage_opamp_dummy_magic_0.VOUT+.n37 two_stage_opamp_dummy_magic_0.VOUT+.t123 4.5005
R5995 two_stage_opamp_dummy_magic_0.VOUT+.n39 two_stage_opamp_dummy_magic_0.VOUT+.t154 4.5005
R5996 two_stage_opamp_dummy_magic_0.VOUT+.n41 two_stage_opamp_dummy_magic_0.VOUT+.t124 4.5005
R5997 two_stage_opamp_dummy_magic_0.VOUT+.n40 two_stage_opamp_dummy_magic_0.VOUT+.t86 4.5005
R5998 two_stage_opamp_dummy_magic_0.VOUT+.n94 two_stage_opamp_dummy_magic_0.VOUT+.t105 4.5005
R5999 two_stage_opamp_dummy_magic_0.VOUT+.n93 two_stage_opamp_dummy_magic_0.VOUT+.t53 4.5005
R6000 two_stage_opamp_dummy_magic_0.VOUT+.n92 two_stage_opamp_dummy_magic_0.VOUT+.t22 4.5005
R6001 two_stage_opamp_dummy_magic_0.VOUT+.n91 two_stage_opamp_dummy_magic_0.VOUT+.t127 4.5005
R6002 two_stage_opamp_dummy_magic_0.VOUT+.n15 two_stage_opamp_dummy_magic_0.VOUT+.n13 4.5005
R6003 two_stage_opamp_dummy_magic_0.VOUT+.n3 two_stage_opamp_dummy_magic_0.VOUT+.t4 3.42907
R6004 two_stage_opamp_dummy_magic_0.VOUT+.n3 two_stage_opamp_dummy_magic_0.VOUT+.t14 3.42907
R6005 two_stage_opamp_dummy_magic_0.VOUT+.n1 two_stage_opamp_dummy_magic_0.VOUT+.t18 3.42907
R6006 two_stage_opamp_dummy_magic_0.VOUT+.n1 two_stage_opamp_dummy_magic_0.VOUT+.t3 3.42907
R6007 two_stage_opamp_dummy_magic_0.VOUT+.n0 two_stage_opamp_dummy_magic_0.VOUT+.t15 3.42907
R6008 two_stage_opamp_dummy_magic_0.VOUT+.n0 two_stage_opamp_dummy_magic_0.VOUT+.t16 3.42907
R6009 two_stage_opamp_dummy_magic_0.VOUT+.n96 two_stage_opamp_dummy_magic_0.VOUT+.n4 2.03175
R6010 two_stage_opamp_dummy_magic_0.VOUT+.n4 two_stage_opamp_dummy_magic_0.VOUT+.n2 1.1255
R6011 two_stage_opamp_dummy_magic_0.VOUT+.n10 two_stage_opamp_dummy_magic_0.VOUT+.n8 0.563
R6012 two_stage_opamp_dummy_magic_0.VOUT+.n12 two_stage_opamp_dummy_magic_0.VOUT+.n10 0.563
R6013 two_stage_opamp_dummy_magic_0.VOUT+.n13 two_stage_opamp_dummy_magic_0.VOUT+.n12 0.563
R6014 two_stage_opamp_dummy_magic_0.VOUT+.n43 two_stage_opamp_dummy_magic_0.VOUT+.n42 0.3295
R6015 two_stage_opamp_dummy_magic_0.VOUT+.n45 two_stage_opamp_dummy_magic_0.VOUT+.n44 0.3295
R6016 two_stage_opamp_dummy_magic_0.VOUT+.n47 two_stage_opamp_dummy_magic_0.VOUT+.n46 0.3295
R6017 two_stage_opamp_dummy_magic_0.VOUT+.n49 two_stage_opamp_dummy_magic_0.VOUT+.n48 0.3295
R6018 two_stage_opamp_dummy_magic_0.VOUT+.n51 two_stage_opamp_dummy_magic_0.VOUT+.n50 0.3295
R6019 two_stage_opamp_dummy_magic_0.VOUT+.n53 two_stage_opamp_dummy_magic_0.VOUT+.n52 0.3295
R6020 two_stage_opamp_dummy_magic_0.VOUT+.n54 two_stage_opamp_dummy_magic_0.VOUT+.n53 0.3295
R6021 two_stage_opamp_dummy_magic_0.VOUT+.n55 two_stage_opamp_dummy_magic_0.VOUT+.n54 0.3295
R6022 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.n55 0.3295
R6023 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.n56 0.3295
R6024 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.n57 0.3295
R6025 two_stage_opamp_dummy_magic_0.VOUT+.n59 two_stage_opamp_dummy_magic_0.VOUT+.n58 0.3295
R6026 two_stage_opamp_dummy_magic_0.VOUT+.n60 two_stage_opamp_dummy_magic_0.VOUT+.n59 0.3295
R6027 two_stage_opamp_dummy_magic_0.VOUT+.n61 two_stage_opamp_dummy_magic_0.VOUT+.n60 0.3295
R6028 two_stage_opamp_dummy_magic_0.VOUT+.n63 two_stage_opamp_dummy_magic_0.VOUT+.n61 0.3295
R6029 two_stage_opamp_dummy_magic_0.VOUT+.n63 two_stage_opamp_dummy_magic_0.VOUT+.n62 0.3295
R6030 two_stage_opamp_dummy_magic_0.VOUT+.n66 two_stage_opamp_dummy_magic_0.VOUT+.n64 0.3295
R6031 two_stage_opamp_dummy_magic_0.VOUT+.n66 two_stage_opamp_dummy_magic_0.VOUT+.n65 0.3295
R6032 two_stage_opamp_dummy_magic_0.VOUT+.n69 two_stage_opamp_dummy_magic_0.VOUT+.n67 0.3295
R6033 two_stage_opamp_dummy_magic_0.VOUT+.n69 two_stage_opamp_dummy_magic_0.VOUT+.n68 0.3295
R6034 two_stage_opamp_dummy_magic_0.VOUT+.n72 two_stage_opamp_dummy_magic_0.VOUT+.n70 0.3295
R6035 two_stage_opamp_dummy_magic_0.VOUT+.n72 two_stage_opamp_dummy_magic_0.VOUT+.n71 0.3295
R6036 two_stage_opamp_dummy_magic_0.VOUT+.n75 two_stage_opamp_dummy_magic_0.VOUT+.n73 0.3295
R6037 two_stage_opamp_dummy_magic_0.VOUT+.n75 two_stage_opamp_dummy_magic_0.VOUT+.n74 0.3295
R6038 two_stage_opamp_dummy_magic_0.VOUT+.n78 two_stage_opamp_dummy_magic_0.VOUT+.n76 0.3295
R6039 two_stage_opamp_dummy_magic_0.VOUT+.n78 two_stage_opamp_dummy_magic_0.VOUT+.n77 0.3295
R6040 two_stage_opamp_dummy_magic_0.VOUT+.n81 two_stage_opamp_dummy_magic_0.VOUT+.n79 0.3295
R6041 two_stage_opamp_dummy_magic_0.VOUT+.n81 two_stage_opamp_dummy_magic_0.VOUT+.n80 0.3295
R6042 two_stage_opamp_dummy_magic_0.VOUT+.n84 two_stage_opamp_dummy_magic_0.VOUT+.n82 0.3295
R6043 two_stage_opamp_dummy_magic_0.VOUT+.n84 two_stage_opamp_dummy_magic_0.VOUT+.n83 0.3295
R6044 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.n85 0.3295
R6045 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.n86 0.3295
R6046 two_stage_opamp_dummy_magic_0.VOUT+.n90 two_stage_opamp_dummy_magic_0.VOUT+.n88 0.3295
R6047 two_stage_opamp_dummy_magic_0.VOUT+.n90 two_stage_opamp_dummy_magic_0.VOUT+.n89 0.3295
R6048 two_stage_opamp_dummy_magic_0.VOUT+.n17 two_stage_opamp_dummy_magic_0.VOUT+.n16 0.3295
R6049 two_stage_opamp_dummy_magic_0.VOUT+.n19 two_stage_opamp_dummy_magic_0.VOUT+.n18 0.3295
R6050 two_stage_opamp_dummy_magic_0.VOUT+.n20 two_stage_opamp_dummy_magic_0.VOUT+.n19 0.3295
R6051 two_stage_opamp_dummy_magic_0.VOUT+.n21 two_stage_opamp_dummy_magic_0.VOUT+.n20 0.3295
R6052 two_stage_opamp_dummy_magic_0.VOUT+.n22 two_stage_opamp_dummy_magic_0.VOUT+.n21 0.3295
R6053 two_stage_opamp_dummy_magic_0.VOUT+.n23 two_stage_opamp_dummy_magic_0.VOUT+.n22 0.3295
R6054 two_stage_opamp_dummy_magic_0.VOUT+.n24 two_stage_opamp_dummy_magic_0.VOUT+.n23 0.3295
R6055 two_stage_opamp_dummy_magic_0.VOUT+.n25 two_stage_opamp_dummy_magic_0.VOUT+.n24 0.3295
R6056 two_stage_opamp_dummy_magic_0.VOUT+.n26 two_stage_opamp_dummy_magic_0.VOUT+.n25 0.3295
R6057 two_stage_opamp_dummy_magic_0.VOUT+.n27 two_stage_opamp_dummy_magic_0.VOUT+.n26 0.3295
R6058 two_stage_opamp_dummy_magic_0.VOUT+.n29 two_stage_opamp_dummy_magic_0.VOUT+.n27 0.3295
R6059 two_stage_opamp_dummy_magic_0.VOUT+.n29 two_stage_opamp_dummy_magic_0.VOUT+.n28 0.3295
R6060 two_stage_opamp_dummy_magic_0.VOUT+.n32 two_stage_opamp_dummy_magic_0.VOUT+.n30 0.3295
R6061 two_stage_opamp_dummy_magic_0.VOUT+.n32 two_stage_opamp_dummy_magic_0.VOUT+.n31 0.3295
R6062 two_stage_opamp_dummy_magic_0.VOUT+.n35 two_stage_opamp_dummy_magic_0.VOUT+.n33 0.3295
R6063 two_stage_opamp_dummy_magic_0.VOUT+.n35 two_stage_opamp_dummy_magic_0.VOUT+.n34 0.3295
R6064 two_stage_opamp_dummy_magic_0.VOUT+.n38 two_stage_opamp_dummy_magic_0.VOUT+.n36 0.3295
R6065 two_stage_opamp_dummy_magic_0.VOUT+.n38 two_stage_opamp_dummy_magic_0.VOUT+.n37 0.3295
R6066 two_stage_opamp_dummy_magic_0.VOUT+.n41 two_stage_opamp_dummy_magic_0.VOUT+.n39 0.3295
R6067 two_stage_opamp_dummy_magic_0.VOUT+.n41 two_stage_opamp_dummy_magic_0.VOUT+.n40 0.3295
R6068 two_stage_opamp_dummy_magic_0.VOUT+.n94 two_stage_opamp_dummy_magic_0.VOUT+.n93 0.3295
R6069 two_stage_opamp_dummy_magic_0.VOUT+.n93 two_stage_opamp_dummy_magic_0.VOUT+.n92 0.3295
R6070 two_stage_opamp_dummy_magic_0.VOUT+.n92 two_stage_opamp_dummy_magic_0.VOUT+.n91 0.3295
R6071 two_stage_opamp_dummy_magic_0.VOUT+.n59 two_stage_opamp_dummy_magic_0.VOUT+.n45 0.306
R6072 two_stage_opamp_dummy_magic_0.VOUT+.n58 two_stage_opamp_dummy_magic_0.VOUT+.n47 0.306
R6073 two_stage_opamp_dummy_magic_0.VOUT+.n57 two_stage_opamp_dummy_magic_0.VOUT+.n49 0.306
R6074 two_stage_opamp_dummy_magic_0.VOUT+.n56 two_stage_opamp_dummy_magic_0.VOUT+.n51 0.306
R6075 two_stage_opamp_dummy_magic_0.VOUT+.n63 two_stage_opamp_dummy_magic_0.VOUT+.n43 0.2825
R6076 two_stage_opamp_dummy_magic_0.VOUT+.n66 two_stage_opamp_dummy_magic_0.VOUT+.n63 0.2825
R6077 two_stage_opamp_dummy_magic_0.VOUT+.n69 two_stage_opamp_dummy_magic_0.VOUT+.n66 0.2825
R6078 two_stage_opamp_dummy_magic_0.VOUT+.n72 two_stage_opamp_dummy_magic_0.VOUT+.n69 0.2825
R6079 two_stage_opamp_dummy_magic_0.VOUT+.n75 two_stage_opamp_dummy_magic_0.VOUT+.n72 0.2825
R6080 two_stage_opamp_dummy_magic_0.VOUT+.n78 two_stage_opamp_dummy_magic_0.VOUT+.n75 0.2825
R6081 two_stage_opamp_dummy_magic_0.VOUT+.n81 two_stage_opamp_dummy_magic_0.VOUT+.n78 0.2825
R6082 two_stage_opamp_dummy_magic_0.VOUT+.n84 two_stage_opamp_dummy_magic_0.VOUT+.n81 0.2825
R6083 two_stage_opamp_dummy_magic_0.VOUT+.n87 two_stage_opamp_dummy_magic_0.VOUT+.n84 0.2825
R6084 two_stage_opamp_dummy_magic_0.VOUT+.n90 two_stage_opamp_dummy_magic_0.VOUT+.n87 0.2825
R6085 two_stage_opamp_dummy_magic_0.VOUT+.n29 two_stage_opamp_dummy_magic_0.VOUT+.n17 0.2825
R6086 two_stage_opamp_dummy_magic_0.VOUT+.n32 two_stage_opamp_dummy_magic_0.VOUT+.n29 0.2825
R6087 two_stage_opamp_dummy_magic_0.VOUT+.n35 two_stage_opamp_dummy_magic_0.VOUT+.n32 0.2825
R6088 two_stage_opamp_dummy_magic_0.VOUT+.n38 two_stage_opamp_dummy_magic_0.VOUT+.n35 0.2825
R6089 two_stage_opamp_dummy_magic_0.VOUT+.n41 two_stage_opamp_dummy_magic_0.VOUT+.n38 0.2825
R6090 two_stage_opamp_dummy_magic_0.VOUT+.n92 two_stage_opamp_dummy_magic_0.VOUT+.n41 0.2825
R6091 two_stage_opamp_dummy_magic_0.VOUT+.n92 two_stage_opamp_dummy_magic_0.VOUT+.n90 0.2825
R6092 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.cap_res_Y.t0 49.083
R6093 two_stage_opamp_dummy_magic_0.cap_res_Y two_stage_opamp_dummy_magic_0.cap_res_Y.t126 0.922875
R6094 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 0.1603
R6095 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 0.1603
R6096 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 0.1603
R6097 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 0.1603
R6098 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 0.1603
R6099 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 0.1603
R6100 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 0.1603
R6101 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 0.1603
R6102 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 0.1603
R6103 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 0.1603
R6104 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 0.1603
R6105 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 0.1603
R6106 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 0.1603
R6107 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 0.1603
R6108 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 0.1603
R6109 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 0.1603
R6110 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 0.1603
R6111 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 0.1603
R6112 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 0.1603
R6113 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 0.1603
R6114 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 0.1603
R6115 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 0.1603
R6116 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 0.1603
R6117 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 0.1603
R6118 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 0.1603
R6119 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 0.1603
R6120 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 0.1603
R6121 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 0.1603
R6122 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 0.1603
R6123 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 0.1603
R6124 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 0.1603
R6125 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 0.1603
R6126 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 0.1603
R6127 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 0.1603
R6128 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 0.1603
R6129 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 0.1603
R6130 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 0.1603
R6131 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 0.1603
R6132 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 0.1603
R6133 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 0.1603
R6134 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 0.1603
R6135 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 0.1603
R6136 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 0.1603
R6137 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 0.1603
R6138 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 0.1603
R6139 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 0.1603
R6140 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 0.1603
R6141 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 0.1603
R6142 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 0.1603
R6143 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 0.1603
R6144 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 0.1603
R6145 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 0.1603
R6146 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 0.1603
R6147 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 0.1603
R6148 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 0.1603
R6149 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 0.1603
R6150 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 0.1603
R6151 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 0.1603
R6152 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 0.159278
R6153 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 0.159278
R6154 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 0.159278
R6155 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 0.159278
R6156 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 0.159278
R6157 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 0.159278
R6158 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 0.159278
R6159 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 0.159278
R6160 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 0.159278
R6161 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 0.159278
R6162 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 0.159278
R6163 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 0.159278
R6164 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 0.159278
R6165 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 0.159278
R6166 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 0.159278
R6167 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 0.159278
R6168 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 0.159278
R6169 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 0.159278
R6170 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 0.159278
R6171 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 0.159278
R6172 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 0.159278
R6173 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 0.159278
R6174 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 0.159278
R6175 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 0.159278
R6176 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 0.159278
R6177 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 0.159278
R6178 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 0.159278
R6179 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 0.137822
R6180 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 0.1368
R6181 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 0.1368
R6182 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 0.1368
R6183 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 0.1368
R6184 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 0.1368
R6185 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 0.1368
R6186 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 0.1368
R6187 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 0.1368
R6188 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 0.1368
R6189 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 0.1368
R6190 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 0.1368
R6191 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 0.1368
R6192 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 0.1368
R6193 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 0.1368
R6194 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 0.1368
R6195 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 0.1368
R6196 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 0.1368
R6197 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 0.1368
R6198 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 0.1368
R6199 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 0.1368
R6200 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 0.1368
R6201 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 0.1368
R6202 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 0.1368
R6203 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 0.1368
R6204 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 0.1368
R6205 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 0.1368
R6206 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 0.1368
R6207 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 0.1368
R6208 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 0.1368
R6209 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 0.1368
R6210 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 0.1368
R6211 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 0.114322
R6212 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 0.1133
R6213 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 0.1133
R6214 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 0.1133
R6215 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 0.1133
R6216 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 0.1133
R6217 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 0.1133
R6218 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 0.1133
R6219 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 0.1133
R6220 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 0.1133
R6221 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 0.1133
R6222 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 0.1133
R6223 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 0.1133
R6224 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 0.1133
R6225 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 0.1133
R6226 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 0.1133
R6227 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 0.1133
R6228 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 0.1133
R6229 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 0.1133
R6230 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 0.1133
R6231 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 0.00152174
R6232 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 0.00152174
R6233 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 0.00152174
R6234 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 0.00152174
R6235 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 0.00152174
R6236 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 0.00152174
R6237 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 0.00152174
R6238 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 0.00152174
R6239 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 0.00152174
R6240 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 0.00152174
R6241 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 0.00152174
R6242 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 0.00152174
R6243 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 0.00152174
R6244 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 0.00152174
R6245 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 0.00152174
R6246 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 0.00152174
R6247 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 0.00152174
R6248 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 0.00152174
R6249 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 0.00152174
R6250 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 0.00152174
R6251 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 0.00152174
R6252 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 0.00152174
R6253 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 0.00152174
R6254 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 0.00152174
R6255 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 0.00152174
R6256 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 0.00152174
R6257 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 0.00152174
R6258 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 0.00152174
R6259 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 0.00152174
R6260 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 0.00152174
R6261 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 0.00152174
R6262 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 0.00152174
R6263 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 0.00152174
R6264 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 0.00152174
R6265 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 0.00152174
R6266 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 0.00152174
R6267 bgr_0.Vbe2.n145 bgr_0.Vbe2.n144 413.99
R6268 bgr_0.Vbe2.n136 bgr_0.Vbe2.t8 162.458
R6269 bgr_0.Vbe2.n146 bgr_0.Vbe2.n145 84.0884
R6270 bgr_0.Vbe2.n60 bgr_0.Vbe2.n59 83.5719
R6271 bgr_0.Vbe2.n55 bgr_0.Vbe2.n48 83.5719
R6272 bgr_0.Vbe2.n54 bgr_0.Vbe2.n53 83.5719
R6273 bgr_0.Vbe2.n127 bgr_0.Vbe2.n6 83.5719
R6274 bgr_0.Vbe2.n122 bgr_0.Vbe2.n7 83.5719
R6275 bgr_0.Vbe2.n45 bgr_0.Vbe2.n44 83.5719
R6276 bgr_0.Vbe2.n43 bgr_0.Vbe2.n42 83.5719
R6277 bgr_0.Vbe2.n41 bgr_0.Vbe2.n40 83.5719
R6278 bgr_0.Vbe2.n78 bgr_0.Vbe2.n77 83.5719
R6279 bgr_0.Vbe2.n76 bgr_0.Vbe2.n75 83.5719
R6280 bgr_0.Vbe2.n27 bgr_0.Vbe2.n26 83.5719
R6281 bgr_0.Vbe2.n86 bgr_0.Vbe2.n85 83.5719
R6282 bgr_0.Vbe2.n22 bgr_0.Vbe2.n20 83.5719
R6283 bgr_0.Vbe2.n91 bgr_0.Vbe2.n19 83.5719
R6284 bgr_0.Vbe2.n99 bgr_0.Vbe2.n98 83.5719
R6285 bgr_0.Vbe2.n17 bgr_0.Vbe2.n16 83.5719
R6286 bgr_0.Vbe2.n114 bgr_0.Vbe2.n113 83.5719
R6287 bgr_0.Vbe2.n112 bgr_0.Vbe2.n111 83.5719
R6288 bgr_0.Vbe2.n110 bgr_0.Vbe2.n109 83.5719
R6289 bgr_0.Vbe2.n143 bgr_0.Vbe2.n1 83.5719
R6290 bgr_0.Vbe2.n142 bgr_0.Vbe2.n0 83.5719
R6291 bgr_0.Vbe2.n141 bgr_0.Vbe2.n140 83.5719
R6292 bgr_0.Vbe2.n132 bgr_0.Vbe2.n4 83.5719
R6293 bgr_0.Vbe2.n72 bgr_0.Vbe2.n26 73.8495
R6294 bgr_0.Vbe2.n59 bgr_0.Vbe2.n58 73.3165
R6295 bgr_0.Vbe2.n129 bgr_0.Vbe2.n6 73.3165
R6296 bgr_0.Vbe2.n44 bgr_0.Vbe2.n36 73.3165
R6297 bgr_0.Vbe2.n85 bgr_0.Vbe2.n84 73.3165
R6298 bgr_0.Vbe2.n98 bgr_0.Vbe2.n97 73.3165
R6299 bgr_0.Vbe2.n115 bgr_0.Vbe2.n114 73.3165
R6300 bgr_0.Vbe2.n54 bgr_0.Vbe2.n49 73.19
R6301 bgr_0.Vbe2.n41 bgr_0.Vbe2.n39 73.19
R6302 bgr_0.Vbe2.n77 bgr_0.Vbe2.n23 73.19
R6303 bgr_0.Vbe2.n93 bgr_0.Vbe2.n19 73.19
R6304 bgr_0.Vbe2.n110 bgr_0.Vbe2.n13 73.19
R6305 bgr_0.Vbe2.n133 bgr_0.Vbe2.n132 73.19
R6306 bgr_0.Vbe2.n123 bgr_0.Vbe2.t4 65.0299
R6307 bgr_0.Vbe2.t6 bgr_0.Vbe2.n14 65.0299
R6308 bgr_0.Vbe2.n59 bgr_0.Vbe2.n55 26.074
R6309 bgr_0.Vbe2.n122 bgr_0.Vbe2.n6 26.074
R6310 bgr_0.Vbe2.n44 bgr_0.Vbe2.n43 26.074
R6311 bgr_0.Vbe2.n76 bgr_0.Vbe2.n26 26.074
R6312 bgr_0.Vbe2.n85 bgr_0.Vbe2.n22 26.074
R6313 bgr_0.Vbe2.n98 bgr_0.Vbe2.n17 26.074
R6314 bgr_0.Vbe2.n114 bgr_0.Vbe2.n112 26.074
R6315 bgr_0.Vbe2.n142 bgr_0.Vbe2.n141 26.074
R6316 bgr_0.Vbe2.n143 bgr_0.Vbe2.n142 26.074
R6317 bgr_0.Vbe2.n145 bgr_0.Vbe2.n143 26.074
R6318 bgr_0.Vbe2.t0 bgr_0.Vbe2.n54 25.7843
R6319 bgr_0.Vbe2.t2 bgr_0.Vbe2.n41 25.7843
R6320 bgr_0.Vbe2.n77 bgr_0.Vbe2.t3 25.7843
R6321 bgr_0.Vbe2.t1 bgr_0.Vbe2.n19 25.7843
R6322 bgr_0.Vbe2.t5 bgr_0.Vbe2.n110 25.7843
R6323 bgr_0.Vbe2.n132 bgr_0.Vbe2.t7 25.7843
R6324 bgr_0.Vbe2.n116 bgr_0.Vbe2.n104 9.3005
R6325 bgr_0.Vbe2.n104 bgr_0.Vbe2.n11 9.3005
R6326 bgr_0.Vbe2.n104 bgr_0.Vbe2.n12 9.3005
R6327 bgr_0.Vbe2.n120 bgr_0.Vbe2.n104 9.3005
R6328 bgr_0.Vbe2.n106 bgr_0.Vbe2.n11 9.3005
R6329 bgr_0.Vbe2.n106 bgr_0.Vbe2.n12 9.3005
R6330 bgr_0.Vbe2.n106 bgr_0.Vbe2.n9 9.3005
R6331 bgr_0.Vbe2.n120 bgr_0.Vbe2.n106 9.3005
R6332 bgr_0.Vbe2.n121 bgr_0.Vbe2.n11 9.3005
R6333 bgr_0.Vbe2.n121 bgr_0.Vbe2.n10 9.3005
R6334 bgr_0.Vbe2.n121 bgr_0.Vbe2.n12 9.3005
R6335 bgr_0.Vbe2.n121 bgr_0.Vbe2.n9 9.3005
R6336 bgr_0.Vbe2.n121 bgr_0.Vbe2.n120 9.3005
R6337 bgr_0.Vbe2.n120 bgr_0.Vbe2.n108 9.3005
R6338 bgr_0.Vbe2.n108 bgr_0.Vbe2.n9 9.3005
R6339 bgr_0.Vbe2.n108 bgr_0.Vbe2.n12 9.3005
R6340 bgr_0.Vbe2.n108 bgr_0.Vbe2.n10 9.3005
R6341 bgr_0.Vbe2.n120 bgr_0.Vbe2.n103 9.3005
R6342 bgr_0.Vbe2.n103 bgr_0.Vbe2.n9 9.3005
R6343 bgr_0.Vbe2.n103 bgr_0.Vbe2.n12 9.3005
R6344 bgr_0.Vbe2.n103 bgr_0.Vbe2.n10 9.3005
R6345 bgr_0.Vbe2.n116 bgr_0.Vbe2.n103 9.3005
R6346 bgr_0.Vbe2.n119 bgr_0.Vbe2.n11 9.3005
R6347 bgr_0.Vbe2.n119 bgr_0.Vbe2.n10 9.3005
R6348 bgr_0.Vbe2.n119 bgr_0.Vbe2.n12 9.3005
R6349 bgr_0.Vbe2.n120 bgr_0.Vbe2.n119 9.3005
R6350 bgr_0.Vbe2.n69 bgr_0.Vbe2.n68 9.3005
R6351 bgr_0.Vbe2.n68 bgr_0.Vbe2.n67 9.3005
R6352 bgr_0.Vbe2.n68 bgr_0.Vbe2.n29 9.3005
R6353 bgr_0.Vbe2.n68 bgr_0.Vbe2.n30 9.3005
R6354 bgr_0.Vbe2.n67 bgr_0.Vbe2.n65 9.3005
R6355 bgr_0.Vbe2.n65 bgr_0.Vbe2.n29 9.3005
R6356 bgr_0.Vbe2.n65 bgr_0.Vbe2.n31 9.3005
R6357 bgr_0.Vbe2.n65 bgr_0.Vbe2.n30 9.3005
R6358 bgr_0.Vbe2.n67 bgr_0.Vbe2.n64 9.3005
R6359 bgr_0.Vbe2.n64 bgr_0.Vbe2.n32 9.3005
R6360 bgr_0.Vbe2.n64 bgr_0.Vbe2.n29 9.3005
R6361 bgr_0.Vbe2.n64 bgr_0.Vbe2.n31 9.3005
R6362 bgr_0.Vbe2.n64 bgr_0.Vbe2.n30 9.3005
R6363 bgr_0.Vbe2.n33 bgr_0.Vbe2.n30 9.3005
R6364 bgr_0.Vbe2.n33 bgr_0.Vbe2.n31 9.3005
R6365 bgr_0.Vbe2.n33 bgr_0.Vbe2.n29 9.3005
R6366 bgr_0.Vbe2.n33 bgr_0.Vbe2.n32 9.3005
R6367 bgr_0.Vbe2.n70 bgr_0.Vbe2.n30 9.3005
R6368 bgr_0.Vbe2.n70 bgr_0.Vbe2.n31 9.3005
R6369 bgr_0.Vbe2.n70 bgr_0.Vbe2.n29 9.3005
R6370 bgr_0.Vbe2.n70 bgr_0.Vbe2.n32 9.3005
R6371 bgr_0.Vbe2.n70 bgr_0.Vbe2.n69 9.3005
R6372 bgr_0.Vbe2.n67 bgr_0.Vbe2.n66 9.3005
R6373 bgr_0.Vbe2.n66 bgr_0.Vbe2.n32 9.3005
R6374 bgr_0.Vbe2.n66 bgr_0.Vbe2.n29 9.3005
R6375 bgr_0.Vbe2.n66 bgr_0.Vbe2.n30 9.3005
R6376 bgr_0.Vbe2.n118 bgr_0.Vbe2.n9 4.64654
R6377 bgr_0.Vbe2.n105 bgr_0.Vbe2.n10 4.64654
R6378 bgr_0.Vbe2.n116 bgr_0.Vbe2.n8 4.64654
R6379 bgr_0.Vbe2.n107 bgr_0.Vbe2.n11 4.64654
R6380 bgr_0.Vbe2.n117 bgr_0.Vbe2.n116 4.64654
R6381 bgr_0.Vbe2.n37 bgr_0.Vbe2.n31 4.64654
R6382 bgr_0.Vbe2.n38 bgr_0.Vbe2.n32 4.64654
R6383 bgr_0.Vbe2.n69 bgr_0.Vbe2.n35 4.64654
R6384 bgr_0.Vbe2.n67 bgr_0.Vbe2.n28 4.64654
R6385 bgr_0.Vbe2.n69 bgr_0.Vbe2.n34 4.64654
R6386 bgr_0.Vbe2.n49 bgr_0.Vbe2.n3 2.36206
R6387 bgr_0.Vbe2.n81 bgr_0.Vbe2.n23 2.36206
R6388 bgr_0.Vbe2.n94 bgr_0.Vbe2.n93 2.36206
R6389 bgr_0.Vbe2.n133 bgr_0.Vbe2.n131 2.36206
R6390 bgr_0.Vbe2.n58 bgr_0.Vbe2.n56 2.19742
R6391 bgr_0.Vbe2.n130 bgr_0.Vbe2.n129 2.19742
R6392 bgr_0.Vbe2.n84 bgr_0.Vbe2.n82 2.19742
R6393 bgr_0.Vbe2.n97 bgr_0.Vbe2.n95 2.19742
R6394 bgr_0.Vbe2.n123 bgr_0.Vbe2.n7 1.56363
R6395 bgr_0.Vbe2.n16 bgr_0.Vbe2.n14 1.56363
R6396 bgr_0.Vbe2.n96 bgr_0.Vbe2.n15 1.5505
R6397 bgr_0.Vbe2.n101 bgr_0.Vbe2.n100 1.5505
R6398 bgr_0.Vbe2.n83 bgr_0.Vbe2.n21 1.5505
R6399 bgr_0.Vbe2.n88 bgr_0.Vbe2.n87 1.5505
R6400 bgr_0.Vbe2.n90 bgr_0.Vbe2.n89 1.5505
R6401 bgr_0.Vbe2.n92 bgr_0.Vbe2.n18 1.5505
R6402 bgr_0.Vbe2.n74 bgr_0.Vbe2.n73 1.5505
R6403 bgr_0.Vbe2.n80 bgr_0.Vbe2.n79 1.5505
R6404 bgr_0.Vbe2.n25 bgr_0.Vbe2.n24 1.5505
R6405 bgr_0.Vbe2.n128 bgr_0.Vbe2.n5 1.5505
R6406 bgr_0.Vbe2.n126 bgr_0.Vbe2.n125 1.5505
R6407 bgr_0.Vbe2.n57 bgr_0.Vbe2.n47 1.5505
R6408 bgr_0.Vbe2.n62 bgr_0.Vbe2.n61 1.5505
R6409 bgr_0.Vbe2.n52 bgr_0.Vbe2.n46 1.5505
R6410 bgr_0.Vbe2.n51 bgr_0.Vbe2.n50 1.5505
R6411 bgr_0.Vbe2.n147 bgr_0.Vbe2.n146 1.5505
R6412 bgr_0.Vbe2.n149 bgr_0.Vbe2.n148 1.5505
R6413 bgr_0.Vbe2.n139 bgr_0.Vbe2.n2 1.5505
R6414 bgr_0.Vbe2.n138 bgr_0.Vbe2.n137 1.5505
R6415 bgr_0.Vbe2.n135 bgr_0.Vbe2.n134 1.5505
R6416 bgr_0.Vbe2.n53 bgr_0.Vbe2.n51 1.25468
R6417 bgr_0.Vbe2.n40 bgr_0.Vbe2.n31 1.25468
R6418 bgr_0.Vbe2.n79 bgr_0.Vbe2.n78 1.25468
R6419 bgr_0.Vbe2.n92 bgr_0.Vbe2.n91 1.25468
R6420 bgr_0.Vbe2.n109 bgr_0.Vbe2.n9 1.25468
R6421 bgr_0.Vbe2.n134 bgr_0.Vbe2.n4 1.25468
R6422 bgr_0.Vbe2.n58 bgr_0.Vbe2.n57 1.19225
R6423 bgr_0.Vbe2.n129 bgr_0.Vbe2.n128 1.19225
R6424 bgr_0.Vbe2.n67 bgr_0.Vbe2.n36 1.19225
R6425 bgr_0.Vbe2.n84 bgr_0.Vbe2.n83 1.19225
R6426 bgr_0.Vbe2.n97 bgr_0.Vbe2.n96 1.19225
R6427 bgr_0.Vbe2.n115 bgr_0.Vbe2.n11 1.19225
R6428 bgr_0.Vbe2.n146 bgr_0.Vbe2.n1 1.14402
R6429 bgr_0.Vbe2.n52 bgr_0.Vbe2.n48 1.07024
R6430 bgr_0.Vbe2.n42 bgr_0.Vbe2.n29 1.07024
R6431 bgr_0.Vbe2.n75 bgr_0.Vbe2.n25 1.07024
R6432 bgr_0.Vbe2.n90 bgr_0.Vbe2.n20 1.07024
R6433 bgr_0.Vbe2.n111 bgr_0.Vbe2.n12 1.07024
R6434 bgr_0.Vbe2.n140 bgr_0.Vbe2.n138 1.07024
R6435 bgr_0.Vbe2.n51 bgr_0.Vbe2.n49 1.0237
R6436 bgr_0.Vbe2.n39 bgr_0.Vbe2.n31 1.0237
R6437 bgr_0.Vbe2.n79 bgr_0.Vbe2.n23 1.0237
R6438 bgr_0.Vbe2.n93 bgr_0.Vbe2.n92 1.0237
R6439 bgr_0.Vbe2.n13 bgr_0.Vbe2.n9 1.0237
R6440 bgr_0.Vbe2.n134 bgr_0.Vbe2.n133 1.0237
R6441 bgr_0.Vbe2.n61 bgr_0.Vbe2.n60 0.885803
R6442 bgr_0.Vbe2.n127 bgr_0.Vbe2.n126 0.885803
R6443 bgr_0.Vbe2.n45 bgr_0.Vbe2.n32 0.885803
R6444 bgr_0.Vbe2.n74 bgr_0.Vbe2.n27 0.885803
R6445 bgr_0.Vbe2.n87 bgr_0.Vbe2.n86 0.885803
R6446 bgr_0.Vbe2.n100 bgr_0.Vbe2.n99 0.885803
R6447 bgr_0.Vbe2.n113 bgr_0.Vbe2.n10 0.885803
R6448 bgr_0.Vbe2.n139 bgr_0.Vbe2.n0 0.885803
R6449 bgr_0.Vbe2.n39 bgr_0.Vbe2.n30 0.812055
R6450 bgr_0.Vbe2.n120 bgr_0.Vbe2.n13 0.812055
R6451 bgr_0.Vbe2.n61 bgr_0.Vbe2.n48 0.77514
R6452 bgr_0.Vbe2.n126 bgr_0.Vbe2.n7 0.77514
R6453 bgr_0.Vbe2.n42 bgr_0.Vbe2.n32 0.77514
R6454 bgr_0.Vbe2.n75 bgr_0.Vbe2.n74 0.77514
R6455 bgr_0.Vbe2.n87 bgr_0.Vbe2.n20 0.77514
R6456 bgr_0.Vbe2.n100 bgr_0.Vbe2.n16 0.77514
R6457 bgr_0.Vbe2.n111 bgr_0.Vbe2.n10 0.77514
R6458 bgr_0.Vbe2.n140 bgr_0.Vbe2.n139 0.77514
R6459 bgr_0.Vbe2.n60 bgr_0.Vbe2 0.756696
R6460 bgr_0.Vbe2 bgr_0.Vbe2.n127 0.756696
R6461 bgr_0.Vbe2 bgr_0.Vbe2.n45 0.756696
R6462 bgr_0.Vbe2 bgr_0.Vbe2.n27 0.756696
R6463 bgr_0.Vbe2.n86 bgr_0.Vbe2 0.756696
R6464 bgr_0.Vbe2.n99 bgr_0.Vbe2 0.756696
R6465 bgr_0.Vbe2.n113 bgr_0.Vbe2 0.756696
R6466 bgr_0.Vbe2 bgr_0.Vbe2.n0 0.756696
R6467 bgr_0.Vbe2.n73 bgr_0.Vbe2.n72 0.711459
R6468 bgr_0.Vbe2.n149 bgr_0.Vbe2.n1 0.701365
R6469 bgr_0.Vbe2.n69 bgr_0.Vbe2.n36 0.647417
R6470 bgr_0.Vbe2.n116 bgr_0.Vbe2.n115 0.647417
R6471 bgr_0.Vbe2.n53 bgr_0.Vbe2.n52 0.590702
R6472 bgr_0.Vbe2.n40 bgr_0.Vbe2.n29 0.590702
R6473 bgr_0.Vbe2.n78 bgr_0.Vbe2.n25 0.590702
R6474 bgr_0.Vbe2.n91 bgr_0.Vbe2.n90 0.590702
R6475 bgr_0.Vbe2.n109 bgr_0.Vbe2.n12 0.590702
R6476 bgr_0.Vbe2.n138 bgr_0.Vbe2.n4 0.590702
R6477 bgr_0.Vbe2.n72 bgr_0.Vbe2 0.576566
R6478 bgr_0.Vbe2.n102 bgr_0.Vbe2.n14 0.530034
R6479 bgr_0.Vbe2.n124 bgr_0.Vbe2.n123 0.530034
R6480 bgr_0.Vbe2.n55 bgr_0.Vbe2.t0 0.290206
R6481 bgr_0.Vbe2.t4 bgr_0.Vbe2.n122 0.290206
R6482 bgr_0.Vbe2.n43 bgr_0.Vbe2.t2 0.290206
R6483 bgr_0.Vbe2.t3 bgr_0.Vbe2.n76 0.290206
R6484 bgr_0.Vbe2.n22 bgr_0.Vbe2.t1 0.290206
R6485 bgr_0.Vbe2.n17 bgr_0.Vbe2.t6 0.290206
R6486 bgr_0.Vbe2.n112 bgr_0.Vbe2.t5 0.290206
R6487 bgr_0.Vbe2.n141 bgr_0.Vbe2.t7 0.290206
R6488 bgr_0.Vbe2.n57 bgr_0.Vbe2 0.203382
R6489 bgr_0.Vbe2.n128 bgr_0.Vbe2 0.203382
R6490 bgr_0.Vbe2.n67 bgr_0.Vbe2 0.203382
R6491 bgr_0.Vbe2.n83 bgr_0.Vbe2 0.203382
R6492 bgr_0.Vbe2.n96 bgr_0.Vbe2 0.203382
R6493 bgr_0.Vbe2 bgr_0.Vbe2.n11 0.203382
R6494 bgr_0.Vbe2 bgr_0.Vbe2.n149 0.203382
R6495 bgr_0.Vbe2.n95 bgr_0.Vbe2.n94 0.154071
R6496 bgr_0.Vbe2.n82 bgr_0.Vbe2.n81 0.154071
R6497 bgr_0.Vbe2.n131 bgr_0.Vbe2.n130 0.154071
R6498 bgr_0.Vbe2.n147 bgr_0.Vbe2.n3 0.154071
R6499 bgr_0.Vbe2.n124 bgr_0.Vbe2.n121 0.137464
R6500 bgr_0.Vbe2.n64 bgr_0.Vbe2.n63 0.137464
R6501 bgr_0.Vbe2.n103 bgr_0.Vbe2.n102 0.134964
R6502 bgr_0.Vbe2.n71 bgr_0.Vbe2.n70 0.134964
R6503 bgr_0.Vbe2.n56 bgr_0.Vbe2 0.0196071
R6504 bgr_0.Vbe2.n101 bgr_0.Vbe2.n15 0.0183571
R6505 bgr_0.Vbe2.n95 bgr_0.Vbe2.n15 0.0183571
R6506 bgr_0.Vbe2.n94 bgr_0.Vbe2.n18 0.0183571
R6507 bgr_0.Vbe2.n89 bgr_0.Vbe2.n18 0.0183571
R6508 bgr_0.Vbe2.n89 bgr_0.Vbe2.n88 0.0183571
R6509 bgr_0.Vbe2.n88 bgr_0.Vbe2.n21 0.0183571
R6510 bgr_0.Vbe2.n82 bgr_0.Vbe2.n21 0.0183571
R6511 bgr_0.Vbe2.n81 bgr_0.Vbe2.n80 0.0183571
R6512 bgr_0.Vbe2.n80 bgr_0.Vbe2.n24 0.0183571
R6513 bgr_0.Vbe2.n125 bgr_0.Vbe2.n5 0.0183571
R6514 bgr_0.Vbe2.n130 bgr_0.Vbe2.n5 0.0183571
R6515 bgr_0.Vbe2.n135 bgr_0.Vbe2.n131 0.0183571
R6516 bgr_0.Vbe2.n137 bgr_0.Vbe2.n135 0.0183571
R6517 bgr_0.Vbe2.n148 bgr_0.Vbe2.n2 0.0183571
R6518 bgr_0.Vbe2.n148 bgr_0.Vbe2.n147 0.0183571
R6519 bgr_0.Vbe2.n50 bgr_0.Vbe2.n3 0.0183571
R6520 bgr_0.Vbe2.n50 bgr_0.Vbe2.n46 0.0183571
R6521 bgr_0.Vbe2.n62 bgr_0.Vbe2.n47 0.0183571
R6522 bgr_0.Vbe2.n56 bgr_0.Vbe2.n47 0.0183571
R6523 bgr_0.Vbe2.n71 bgr_0.Vbe2.n24 0.0106786
R6524 bgr_0.Vbe2.n63 bgr_0.Vbe2.n46 0.0106786
R6525 bgr_0.Vbe2.n136 bgr_0.Vbe2.n2 0.00996429
R6526 bgr_0.Vbe2.n108 bgr_0.Vbe2.n107 0.00992001
R6527 bgr_0.Vbe2.n119 bgr_0.Vbe2.n117 0.00992001
R6528 bgr_0.Vbe2.n118 bgr_0.Vbe2.n104 0.00992001
R6529 bgr_0.Vbe2.n106 bgr_0.Vbe2.n105 0.00992001
R6530 bgr_0.Vbe2.n121 bgr_0.Vbe2.n8 0.00992001
R6531 bgr_0.Vbe2.n105 bgr_0.Vbe2.n104 0.00992001
R6532 bgr_0.Vbe2.n106 bgr_0.Vbe2.n8 0.00992001
R6533 bgr_0.Vbe2.n117 bgr_0.Vbe2.n108 0.00992001
R6534 bgr_0.Vbe2.n107 bgr_0.Vbe2.n103 0.00992001
R6535 bgr_0.Vbe2.n119 bgr_0.Vbe2.n118 0.00992001
R6536 bgr_0.Vbe2.n33 bgr_0.Vbe2.n28 0.00992001
R6537 bgr_0.Vbe2.n66 bgr_0.Vbe2.n34 0.00992001
R6538 bgr_0.Vbe2.n68 bgr_0.Vbe2.n37 0.00992001
R6539 bgr_0.Vbe2.n65 bgr_0.Vbe2.n38 0.00992001
R6540 bgr_0.Vbe2.n64 bgr_0.Vbe2.n35 0.00992001
R6541 bgr_0.Vbe2.n68 bgr_0.Vbe2.n38 0.00992001
R6542 bgr_0.Vbe2.n65 bgr_0.Vbe2.n35 0.00992001
R6543 bgr_0.Vbe2.n34 bgr_0.Vbe2.n33 0.00992001
R6544 bgr_0.Vbe2.n70 bgr_0.Vbe2.n28 0.00992001
R6545 bgr_0.Vbe2.n66 bgr_0.Vbe2.n37 0.00992001
R6546 bgr_0.Vbe2.n137 bgr_0.Vbe2.n136 0.00889286
R6547 bgr_0.Vbe2.n102 bgr_0.Vbe2.n101 0.00817857
R6548 bgr_0.Vbe2.n73 bgr_0.Vbe2.n71 0.00817857
R6549 bgr_0.Vbe2.n125 bgr_0.Vbe2.n124 0.00817857
R6550 bgr_0.Vbe2.n63 bgr_0.Vbe2.n62 0.00817857
R6551 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.t31 1172.87
R6552 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t40 1172.87
R6553 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.t50 996.134
R6554 two_stage_opamp_dummy_magic_0.Y.n49 two_stage_opamp_dummy_magic_0.Y.t39 996.134
R6555 two_stage_opamp_dummy_magic_0.Y.n43 two_stage_opamp_dummy_magic_0.Y.t53 996.134
R6556 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.t43 996.134
R6557 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.t26 996.134
R6558 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.t32 996.134
R6559 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.t48 996.134
R6560 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.t35 996.134
R6561 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t34 690.867
R6562 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t45 690.867
R6563 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t29 530.201
R6564 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t38 530.201
R6565 two_stage_opamp_dummy_magic_0.Y.n32 two_stage_opamp_dummy_magic_0.Y.t44 514.134
R6566 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.t54 514.134
R6567 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.t41 514.134
R6568 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.t51 514.134
R6569 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.t36 514.134
R6570 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.t28 514.134
R6571 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.t46 514.134
R6572 two_stage_opamp_dummy_magic_0.Y.n31 two_stage_opamp_dummy_magic_0.Y.t27 514.134
R6573 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.t42 353.467
R6574 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.t25 353.467
R6575 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.t30 353.467
R6576 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.t47 353.467
R6577 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.t33 353.467
R6578 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.t49 353.467
R6579 two_stage_opamp_dummy_magic_0.Y.n23 two_stage_opamp_dummy_magic_0.Y.t37 353.467
R6580 two_stage_opamp_dummy_magic_0.Y.n22 two_stage_opamp_dummy_magic_0.Y.t52 353.467
R6581 two_stage_opamp_dummy_magic_0.Y.n50 two_stage_opamp_dummy_magic_0.Y.n49 176.733
R6582 two_stage_opamp_dummy_magic_0.Y.n44 two_stage_opamp_dummy_magic_0.Y.n43 176.733
R6583 two_stage_opamp_dummy_magic_0.Y.n45 two_stage_opamp_dummy_magic_0.Y.n44 176.733
R6584 two_stage_opamp_dummy_magic_0.Y.n46 two_stage_opamp_dummy_magic_0.Y.n45 176.733
R6585 two_stage_opamp_dummy_magic_0.Y.n47 two_stage_opamp_dummy_magic_0.Y.n46 176.733
R6586 two_stage_opamp_dummy_magic_0.Y.n48 two_stage_opamp_dummy_magic_0.Y.n47 176.733
R6587 two_stage_opamp_dummy_magic_0.Y.n29 two_stage_opamp_dummy_magic_0.Y.n28 176.733
R6588 two_stage_opamp_dummy_magic_0.Y.n28 two_stage_opamp_dummy_magic_0.Y.n27 176.733
R6589 two_stage_opamp_dummy_magic_0.Y.n27 two_stage_opamp_dummy_magic_0.Y.n26 176.733
R6590 two_stage_opamp_dummy_magic_0.Y.n26 two_stage_opamp_dummy_magic_0.Y.n25 176.733
R6591 two_stage_opamp_dummy_magic_0.Y.n25 two_stage_opamp_dummy_magic_0.Y.n24 176.733
R6592 two_stage_opamp_dummy_magic_0.Y.n24 two_stage_opamp_dummy_magic_0.Y.n23 176.733
R6593 two_stage_opamp_dummy_magic_0.Y.n38 two_stage_opamp_dummy_magic_0.Y.n37 176.733
R6594 two_stage_opamp_dummy_magic_0.Y.n37 two_stage_opamp_dummy_magic_0.Y.n36 176.733
R6595 two_stage_opamp_dummy_magic_0.Y.n36 two_stage_opamp_dummy_magic_0.Y.n35 176.733
R6596 two_stage_opamp_dummy_magic_0.Y.n35 two_stage_opamp_dummy_magic_0.Y.n34 176.733
R6597 two_stage_opamp_dummy_magic_0.Y.n34 two_stage_opamp_dummy_magic_0.Y.n33 176.733
R6598 two_stage_opamp_dummy_magic_0.Y.n33 two_stage_opamp_dummy_magic_0.Y.n32 176.733
R6599 two_stage_opamp_dummy_magic_0.Y.n52 two_stage_opamp_dummy_magic_0.Y.n51 166.436
R6600 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n30 161.843
R6601 two_stage_opamp_dummy_magic_0.Y.n40 two_stage_opamp_dummy_magic_0.Y.n39 161.718
R6602 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.n11 160.427
R6603 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n18 159.802
R6604 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.n16 159.802
R6605 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.n14 159.802
R6606 two_stage_opamp_dummy_magic_0.Y.n13 two_stage_opamp_dummy_magic_0.Y.n12 159.802
R6607 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n20 155.302
R6608 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.n8 114.689
R6609 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.n1 114.689
R6610 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.n6 114.126
R6611 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.n4 114.126
R6612 two_stage_opamp_dummy_magic_0.Y.n3 two_stage_opamp_dummy_magic_0.Y.n2 114.126
R6613 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n0 109.626
R6614 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n50 51.9494
R6615 two_stage_opamp_dummy_magic_0.Y.n51 two_stage_opamp_dummy_magic_0.Y.n48 51.9494
R6616 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n29 51.9494
R6617 two_stage_opamp_dummy_magic_0.Y.n30 two_stage_opamp_dummy_magic_0.Y.n22 51.9494
R6618 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n38 51.9494
R6619 two_stage_opamp_dummy_magic_0.Y.n39 two_stage_opamp_dummy_magic_0.Y.n31 51.9494
R6620 two_stage_opamp_dummy_magic_0.Y.t0 two_stage_opamp_dummy_magic_0.Y.n52 49.3036
R6621 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n21 17.4067
R6622 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.t18 16.0005
R6623 two_stage_opamp_dummy_magic_0.Y.n8 two_stage_opamp_dummy_magic_0.Y.t20 16.0005
R6624 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.t14 16.0005
R6625 two_stage_opamp_dummy_magic_0.Y.n6 two_stage_opamp_dummy_magic_0.Y.t9 16.0005
R6626 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.t24 16.0005
R6627 two_stage_opamp_dummy_magic_0.Y.n4 two_stage_opamp_dummy_magic_0.Y.t15 16.0005
R6628 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.t1 16.0005
R6629 two_stage_opamp_dummy_magic_0.Y.n2 two_stage_opamp_dummy_magic_0.Y.t22 16.0005
R6630 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t19 16.0005
R6631 two_stage_opamp_dummy_magic_0.Y.n1 two_stage_opamp_dummy_magic_0.Y.t5 16.0005
R6632 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t6 16.0005
R6633 two_stage_opamp_dummy_magic_0.Y.n0 two_stage_opamp_dummy_magic_0.Y.t11 16.0005
R6634 two_stage_opamp_dummy_magic_0.Y.n41 two_stage_opamp_dummy_magic_0.Y.n40 13.9693
R6635 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.t10 11.2576
R6636 two_stage_opamp_dummy_magic_0.Y.n20 two_stage_opamp_dummy_magic_0.Y.t12 11.2576
R6637 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.t3 11.2576
R6638 two_stage_opamp_dummy_magic_0.Y.n18 two_stage_opamp_dummy_magic_0.Y.t8 11.2576
R6639 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.t23 11.2576
R6640 two_stage_opamp_dummy_magic_0.Y.n16 two_stage_opamp_dummy_magic_0.Y.t13 11.2576
R6641 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.t16 11.2576
R6642 two_stage_opamp_dummy_magic_0.Y.n14 two_stage_opamp_dummy_magic_0.Y.t21 11.2576
R6643 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t4 11.2576
R6644 two_stage_opamp_dummy_magic_0.Y.n12 two_stage_opamp_dummy_magic_0.Y.t2 11.2576
R6645 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t7 11.2576
R6646 two_stage_opamp_dummy_magic_0.Y.n11 two_stage_opamp_dummy_magic_0.Y.t17 11.2576
R6647 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.n10 9.28175
R6648 two_stage_opamp_dummy_magic_0.Y.n21 two_stage_opamp_dummy_magic_0.Y.n19 5.1255
R6649 two_stage_opamp_dummy_magic_0.Y.n10 two_stage_opamp_dummy_magic_0.Y.n9 4.5005
R6650 two_stage_opamp_dummy_magic_0.Y.n42 two_stage_opamp_dummy_magic_0.Y.n41 4.5005
R6651 two_stage_opamp_dummy_magic_0.Y.n52 two_stage_opamp_dummy_magic_0.Y.n42 3.40675
R6652 two_stage_opamp_dummy_magic_0.Y.n15 two_stage_opamp_dummy_magic_0.Y.n13 0.6255
R6653 two_stage_opamp_dummy_magic_0.Y.n17 two_stage_opamp_dummy_magic_0.Y.n15 0.6255
R6654 two_stage_opamp_dummy_magic_0.Y.n19 two_stage_opamp_dummy_magic_0.Y.n17 0.6255
R6655 two_stage_opamp_dummy_magic_0.Y.n5 two_stage_opamp_dummy_magic_0.Y.n3 0.563
R6656 two_stage_opamp_dummy_magic_0.Y.n7 two_stage_opamp_dummy_magic_0.Y.n5 0.563
R6657 two_stage_opamp_dummy_magic_0.Y.n9 two_stage_opamp_dummy_magic_0.Y.n7 0.563
R6658 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 345.264
R6659 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 344.7
R6660 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 344.7
R6661 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 206.052
R6662 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 205.488
R6663 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 205.488
R6664 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 205.488
R6665 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 205.488
R6666 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 122.504
R6667 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 57.1567
R6668 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 39.4005
R6669 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 39.4005
R6670 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 39.4005
R6671 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 39.4005
R6672 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 39.4005
R6673 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 39.4005
R6674 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 19.7005
R6675 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 19.7005
R6676 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 19.7005
R6677 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 19.7005
R6678 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 19.7005
R6679 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 19.7005
R6680 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 19.7005
R6681 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 19.7005
R6682 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 19.7005
R6683 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 19.7005
R6684 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 6.15675
R6685 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 6.09425
R6686 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 0.563
R6687 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 0.563
R6688 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 0.563
R6689 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 0.563
R6690 bgr_0.V_CMFB_S3 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 0.21925
R6691 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.t0 384.967
R6692 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t5 369.534
R6693 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t20 369.534
R6694 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t23 369.534
R6695 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t15 369.534
R6696 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t17 369.534
R6697 bgr_0.NFET_GATE_10uA.t0 bgr_0.NFET_GATE_10uA.n18 369.534
R6698 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n20 365.491
R6699 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.t12 192.8
R6700 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.t11 192.8
R6701 bgr_0.NFET_GATE_10uA.n10 bgr_0.NFET_GATE_10uA.t19 192.8
R6702 bgr_0.NFET_GATE_10uA.n9 bgr_0.NFET_GATE_10uA.t6 192.8
R6703 bgr_0.NFET_GATE_10uA.n7 bgr_0.NFET_GATE_10uA.t14 192.8
R6704 bgr_0.NFET_GATE_10uA.n4 bgr_0.NFET_GATE_10uA.t13 192.8
R6705 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.t21 192.8
R6706 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.t7 192.8
R6707 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.t16 192.8
R6708 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.t22 192.8
R6709 bgr_0.NFET_GATE_10uA.n1 bgr_0.NFET_GATE_10uA.t9 192.8
R6710 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.t10 192.8
R6711 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.t18 192.8
R6712 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.t8 192.8
R6713 bgr_0.NFET_GATE_10uA.n12 bgr_0.NFET_GATE_10uA.n11 176.733
R6714 bgr_0.NFET_GATE_10uA.n11 bgr_0.NFET_GATE_10uA.n10 176.733
R6715 bgr_0.NFET_GATE_10uA.n5 bgr_0.NFET_GATE_10uA.n4 176.733
R6716 bgr_0.NFET_GATE_10uA.n6 bgr_0.NFET_GATE_10uA.n5 176.733
R6717 bgr_0.NFET_GATE_10uA.n3 bgr_0.NFET_GATE_10uA.n2 176.733
R6718 bgr_0.NFET_GATE_10uA.n2 bgr_0.NFET_GATE_10uA.n1 176.733
R6719 bgr_0.NFET_GATE_10uA.n18 bgr_0.NFET_GATE_10uA.n17 176.733
R6720 bgr_0.NFET_GATE_10uA.n17 bgr_0.NFET_GATE_10uA.n16 176.733
R6721 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n13 169.852
R6722 bgr_0.NFET_GATE_10uA.n14 bgr_0.NFET_GATE_10uA.n8 169.852
R6723 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n14 166.133
R6724 bgr_0.NFET_GATE_10uA.n19 bgr_0.NFET_GATE_10uA.n0 126.877
R6725 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n12 56.2338
R6726 bgr_0.NFET_GATE_10uA.n13 bgr_0.NFET_GATE_10uA.n9 56.2338
R6727 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n7 56.2338
R6728 bgr_0.NFET_GATE_10uA.n8 bgr_0.NFET_GATE_10uA.n6 56.2338
R6729 bgr_0.NFET_GATE_10uA.n15 bgr_0.NFET_GATE_10uA.n3 56.2338
R6730 bgr_0.NFET_GATE_10uA.n16 bgr_0.NFET_GATE_10uA.n15 56.2338
R6731 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t2 39.4005
R6732 bgr_0.NFET_GATE_10uA.n20 bgr_0.NFET_GATE_10uA.t4 39.4005
R6733 bgr_0.NFET_GATE_10uA bgr_0.NFET_GATE_10uA.n19 28.6755
R6734 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t3 24.0005
R6735 bgr_0.NFET_GATE_10uA.n0 bgr_0.NFET_GATE_10uA.t1 24.0005
R6736 bgr_0.V_mir2.n20 bgr_0.V_mir2.n19 325.473
R6737 bgr_0.V_mir2.n13 bgr_0.V_mir2.n12 325.473
R6738 bgr_0.V_mir2.n4 bgr_0.V_mir2.n3 325.473
R6739 bgr_0.V_mir2.n16 bgr_0.V_mir2.t17 310.488
R6740 bgr_0.V_mir2.n9 bgr_0.V_mir2.t22 310.488
R6741 bgr_0.V_mir2.n0 bgr_0.V_mir2.t20 310.488
R6742 bgr_0.V_mir2.n7 bgr_0.V_mir2.t13 278.312
R6743 bgr_0.V_mir2.n7 bgr_0.V_mir2.n6 228.939
R6744 bgr_0.V_mir2.n8 bgr_0.V_mir2.n5 224.439
R6745 bgr_0.V_mir2.n18 bgr_0.V_mir2.t2 184.097
R6746 bgr_0.V_mir2.n11 bgr_0.V_mir2.t6 184.097
R6747 bgr_0.V_mir2.n2 bgr_0.V_mir2.t4 184.097
R6748 bgr_0.V_mir2.n17 bgr_0.V_mir2.n16 167.094
R6749 bgr_0.V_mir2.n10 bgr_0.V_mir2.n9 167.094
R6750 bgr_0.V_mir2.n1 bgr_0.V_mir2.n0 167.094
R6751 bgr_0.V_mir2.n13 bgr_0.V_mir2.n11 152
R6752 bgr_0.V_mir2.n4 bgr_0.V_mir2.n2 152
R6753 bgr_0.V_mir2.n19 bgr_0.V_mir2.n18 152
R6754 bgr_0.V_mir2.n16 bgr_0.V_mir2.t21 120.501
R6755 bgr_0.V_mir2.n17 bgr_0.V_mir2.t10 120.501
R6756 bgr_0.V_mir2.n9 bgr_0.V_mir2.t19 120.501
R6757 bgr_0.V_mir2.n10 bgr_0.V_mir2.t8 120.501
R6758 bgr_0.V_mir2.n0 bgr_0.V_mir2.t18 120.501
R6759 bgr_0.V_mir2.n1 bgr_0.V_mir2.t0 120.501
R6760 bgr_0.V_mir2.n6 bgr_0.V_mir2.t14 48.0005
R6761 bgr_0.V_mir2.n6 bgr_0.V_mir2.t12 48.0005
R6762 bgr_0.V_mir2.n5 bgr_0.V_mir2.t15 48.0005
R6763 bgr_0.V_mir2.n5 bgr_0.V_mir2.t16 48.0005
R6764 bgr_0.V_mir2.n18 bgr_0.V_mir2.n17 40.7027
R6765 bgr_0.V_mir2.n11 bgr_0.V_mir2.n10 40.7027
R6766 bgr_0.V_mir2.n2 bgr_0.V_mir2.n1 40.7027
R6767 bgr_0.V_mir2.n12 bgr_0.V_mir2.t9 39.4005
R6768 bgr_0.V_mir2.n12 bgr_0.V_mir2.t7 39.4005
R6769 bgr_0.V_mir2.n3 bgr_0.V_mir2.t1 39.4005
R6770 bgr_0.V_mir2.n3 bgr_0.V_mir2.t5 39.4005
R6771 bgr_0.V_mir2.t11 bgr_0.V_mir2.n20 39.4005
R6772 bgr_0.V_mir2.n20 bgr_0.V_mir2.t3 39.4005
R6773 bgr_0.V_mir2.n15 bgr_0.V_mir2.n4 15.8005
R6774 bgr_0.V_mir2.n19 bgr_0.V_mir2.n15 15.8005
R6775 bgr_0.V_mir2.n14 bgr_0.V_mir2.n13 9.3005
R6776 bgr_0.V_mir2.n8 bgr_0.V_mir2.n7 5.8755
R6777 bgr_0.V_mir2.n15 bgr_0.V_mir2.n14 4.5005
R6778 bgr_0.V_mir2.n14 bgr_0.V_mir2.n8 0.78175
R6779 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 688.859
R6780 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 514.134
R6781 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 323.491
R6782 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 322.692
R6783 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 270.591
R6784 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 270.591
R6785 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 270.591
R6786 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 270.591
R6787 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 233.374
R6788 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 233.374
R6789 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 233.374
R6790 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 233.374
R6791 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 208.838
R6792 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 197.964
R6793 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 174.726
R6794 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 174.726
R6795 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 174.726
R6796 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 174.726
R6797 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 169.216
R6798 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 169.216
R6799 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 169.216
R6800 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 129.24
R6801 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 129.24
R6802 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 129.24
R6803 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 129.24
R6804 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 128.534
R6805 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 128.534
R6806 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 16.8443
R6807 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 13.1338
R6808 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 13.1338
R6809 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 13.1338
R6810 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 13.1338
R6811 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 13.1338
R6812 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 13.1338
R6813 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 4.3755
R6814 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 4.3755
R6815 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 3.688
R6816 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 3.1255
R6817 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 2.0005
R6818 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 1.2755
R6819 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 1.2755
R6820 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 0.8005
R6821 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 632.186
R6822 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 630.264
R6823 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 630.264
R6824 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 630.264
R6825 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 628.003
R6826 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 628.003
R6827 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 626.753
R6828 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 626.753
R6829 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 625.756
R6830 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 622.231
R6831 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t11 78.8005
R6832 two_stage_opamp_dummy_magic_0.V_err_mir_p.n11 two_stage_opamp_dummy_magic_0.V_err_mir_p.t7 78.8005
R6833 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t9 78.8005
R6834 two_stage_opamp_dummy_magic_0.V_err_mir_p.n10 two_stage_opamp_dummy_magic_0.V_err_mir_p.t19 78.8005
R6835 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t18 78.8005
R6836 two_stage_opamp_dummy_magic_0.V_err_mir_p.n9 two_stage_opamp_dummy_magic_0.V_err_mir_p.t8 78.8005
R6837 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t5 78.8005
R6838 two_stage_opamp_dummy_magic_0.V_err_mir_p.n8 two_stage_opamp_dummy_magic_0.V_err_mir_p.t4 78.8005
R6839 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t1 78.8005
R6840 two_stage_opamp_dummy_magic_0.V_err_mir_p.n7 two_stage_opamp_dummy_magic_0.V_err_mir_p.t15 78.8005
R6841 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t12 78.8005
R6842 two_stage_opamp_dummy_magic_0.V_err_mir_p.n6 two_stage_opamp_dummy_magic_0.V_err_mir_p.t3 78.8005
R6843 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t13 78.8005
R6844 two_stage_opamp_dummy_magic_0.V_err_mir_p.n5 two_stage_opamp_dummy_magic_0.V_err_mir_p.t2 78.8005
R6845 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t16 78.8005
R6846 two_stage_opamp_dummy_magic_0.V_err_mir_p.n4 two_stage_opamp_dummy_magic_0.V_err_mir_p.t14 78.8005
R6847 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t10 78.8005
R6848 two_stage_opamp_dummy_magic_0.V_err_mir_p.n3 two_stage_opamp_dummy_magic_0.V_err_mir_p.t17 78.8005
R6849 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 two_stage_opamp_dummy_magic_0.V_err_mir_p.t6 78.8005
R6850 two_stage_opamp_dummy_magic_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_0.V_err_mir_p.n12 78.8005
R6851 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n0 8.22272
R6852 two_stage_opamp_dummy_magic_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_0.V_err_mir_p.n2 6.188
R6853 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n27 630.264
R6854 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n2 627.316
R6855 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n4 626.784
R6856 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n3 626.784
R6857 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n26 626.784
R6858 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate.n24 585
R6859 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t17 289.2
R6860 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t29 289.2
R6861 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.n21 176.733
R6862 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.n5 176.733
R6863 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.n6 176.733
R6864 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.n7 176.733
R6865 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.n8 176.733
R6866 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.n9 176.733
R6867 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.n10 176.733
R6868 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.n11 176.733
R6869 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.n12 176.733
R6870 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.n13 176.733
R6871 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.n14 176.733
R6872 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.n15 176.733
R6873 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.n16 176.733
R6874 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.n17 176.733
R6875 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.n18 176.733
R6876 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.n19 176.733
R6877 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n23 162.494
R6878 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n28 135.81
R6879 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.V_err_gate.n1 131.392
R6880 two_stage_opamp_dummy_magic_0.V_err_gate.n22 two_stage_opamp_dummy_magic_0.V_err_gate.t14 112.468
R6881 two_stage_opamp_dummy_magic_0.V_err_gate.n21 two_stage_opamp_dummy_magic_0.V_err_gate.t27 112.468
R6882 two_stage_opamp_dummy_magic_0.V_err_gate.n5 two_stage_opamp_dummy_magic_0.V_err_gate.t20 112.468
R6883 two_stage_opamp_dummy_magic_0.V_err_gate.n6 two_stage_opamp_dummy_magic_0.V_err_gate.t26 112.468
R6884 two_stage_opamp_dummy_magic_0.V_err_gate.n7 two_stage_opamp_dummy_magic_0.V_err_gate.t19 112.468
R6885 two_stage_opamp_dummy_magic_0.V_err_gate.n8 two_stage_opamp_dummy_magic_0.V_err_gate.t31 112.468
R6886 two_stage_opamp_dummy_magic_0.V_err_gate.n9 two_stage_opamp_dummy_magic_0.V_err_gate.t22 112.468
R6887 two_stage_opamp_dummy_magic_0.V_err_gate.n10 two_stage_opamp_dummy_magic_0.V_err_gate.t33 112.468
R6888 two_stage_opamp_dummy_magic_0.V_err_gate.n11 two_stage_opamp_dummy_magic_0.V_err_gate.t24 112.468
R6889 two_stage_opamp_dummy_magic_0.V_err_gate.n12 two_stage_opamp_dummy_magic_0.V_err_gate.t15 112.468
R6890 two_stage_opamp_dummy_magic_0.V_err_gate.n13 two_stage_opamp_dummy_magic_0.V_err_gate.t28 112.468
R6891 two_stage_opamp_dummy_magic_0.V_err_gate.n14 two_stage_opamp_dummy_magic_0.V_err_gate.t18 112.468
R6892 two_stage_opamp_dummy_magic_0.V_err_gate.n15 two_stage_opamp_dummy_magic_0.V_err_gate.t25 112.468
R6893 two_stage_opamp_dummy_magic_0.V_err_gate.n16 two_stage_opamp_dummy_magic_0.V_err_gate.t16 112.468
R6894 two_stage_opamp_dummy_magic_0.V_err_gate.n17 two_stage_opamp_dummy_magic_0.V_err_gate.t30 112.468
R6895 two_stage_opamp_dummy_magic_0.V_err_gate.n18 two_stage_opamp_dummy_magic_0.V_err_gate.t21 112.468
R6896 two_stage_opamp_dummy_magic_0.V_err_gate.n19 two_stage_opamp_dummy_magic_0.V_err_gate.t32 112.468
R6897 two_stage_opamp_dummy_magic_0.V_err_gate.n20 two_stage_opamp_dummy_magic_0.V_err_gate.t23 112.468
R6898 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t13 78.8005
R6899 two_stage_opamp_dummy_magic_0.V_err_gate.n4 two_stage_opamp_dummy_magic_0.V_err_gate.t10 78.8005
R6900 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t5 78.8005
R6901 two_stage_opamp_dummy_magic_0.V_err_gate.n3 two_stage_opamp_dummy_magic_0.V_err_gate.t2 78.8005
R6902 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t1 78.8005
R6903 two_stage_opamp_dummy_magic_0.V_err_gate.n2 two_stage_opamp_dummy_magic_0.V_err_gate.t11 78.8005
R6904 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t0 78.8005
R6905 two_stage_opamp_dummy_magic_0.V_err_gate.n26 two_stage_opamp_dummy_magic_0.V_err_gate.t9 78.8005
R6906 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t12 78.8005
R6907 two_stage_opamp_dummy_magic_0.V_err_gate.n27 two_stage_opamp_dummy_magic_0.V_err_gate.t3 78.8005
R6908 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t4 78.8005
R6909 two_stage_opamp_dummy_magic_0.V_err_gate.n24 two_stage_opamp_dummy_magic_0.V_err_gate.t6 78.8005
R6910 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n22 49.8072
R6911 two_stage_opamp_dummy_magic_0.V_err_gate.n23 two_stage_opamp_dummy_magic_0.V_err_gate.n20 49.8072
R6912 two_stage_opamp_dummy_magic_0.V_err_gate.n0 two_stage_opamp_dummy_magic_0.V_err_gate.n25 41.7838
R6913 two_stage_opamp_dummy_magic_0.V_err_gate.n25 two_stage_opamp_dummy_magic_0.V_err_gate 39.8442
R6914 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t8 24.0005
R6915 two_stage_opamp_dummy_magic_0.V_err_gate.n28 two_stage_opamp_dummy_magic_0.V_err_gate.t7 24.0005
R6916 two_stage_opamp_dummy_magic_0.V_err_gate.n1 two_stage_opamp_dummy_magic_0.V_err_gate.n0 2.313
R6917 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.t19 673.034
R6918 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.n0 620.841
R6919 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t28 611.739
R6920 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t16 611.739
R6921 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t22 611.739
R6922 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t31 611.739
R6923 two_stage_opamp_dummy_magic_0.Vb2.n15 two_stage_opamp_dummy_magic_0.Vb2.t11 421.75
R6924 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.t13 421.75
R6925 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.t15 421.75
R6926 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.t18 421.75
R6927 two_stage_opamp_dummy_magic_0.Vb2.n11 two_stage_opamp_dummy_magic_0.Vb2.t14 421.75
R6928 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.t12 421.75
R6929 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.t29 421.75
R6930 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.t24 421.75
R6931 two_stage_opamp_dummy_magic_0.Vb2.n6 two_stage_opamp_dummy_magic_0.Vb2.t27 421.75
R6932 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.t25 421.75
R6933 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.t30 421.75
R6934 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.t17 421.75
R6935 two_stage_opamp_dummy_magic_0.Vb2.n2 two_stage_opamp_dummy_magic_0.Vb2.t26 421.75
R6936 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.t21 421.75
R6937 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.t23 421.75
R6938 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.t20 421.75
R6939 two_stage_opamp_dummy_magic_0.Vb2.n1 two_stage_opamp_dummy_magic_0.Vb2.t0 288.166
R6940 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n10 169.311
R6941 two_stage_opamp_dummy_magic_0.Vb2.n20 two_stage_opamp_dummy_magic_0.Vb2.n19 168.936
R6942 two_stage_opamp_dummy_magic_0.Vb2.n16 two_stage_opamp_dummy_magic_0.Vb2.n15 167.094
R6943 two_stage_opamp_dummy_magic_0.Vb2.n17 two_stage_opamp_dummy_magic_0.Vb2.n16 167.094
R6944 two_stage_opamp_dummy_magic_0.Vb2.n18 two_stage_opamp_dummy_magic_0.Vb2.n17 167.094
R6945 two_stage_opamp_dummy_magic_0.Vb2.n12 two_stage_opamp_dummy_magic_0.Vb2.n11 167.094
R6946 two_stage_opamp_dummy_magic_0.Vb2.n13 two_stage_opamp_dummy_magic_0.Vb2.n12 167.094
R6947 two_stage_opamp_dummy_magic_0.Vb2.n14 two_stage_opamp_dummy_magic_0.Vb2.n13 167.094
R6948 two_stage_opamp_dummy_magic_0.Vb2.n7 two_stage_opamp_dummy_magic_0.Vb2.n6 167.094
R6949 two_stage_opamp_dummy_magic_0.Vb2.n8 two_stage_opamp_dummy_magic_0.Vb2.n7 167.094
R6950 two_stage_opamp_dummy_magic_0.Vb2.n9 two_stage_opamp_dummy_magic_0.Vb2.n8 167.094
R6951 two_stage_opamp_dummy_magic_0.Vb2.n3 two_stage_opamp_dummy_magic_0.Vb2.n2 167.094
R6952 two_stage_opamp_dummy_magic_0.Vb2.n4 two_stage_opamp_dummy_magic_0.Vb2.n3 167.094
R6953 two_stage_opamp_dummy_magic_0.Vb2.n5 two_stage_opamp_dummy_magic_0.Vb2.n4 167.094
R6954 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n24 139.639
R6955 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.n25 139.638
R6956 two_stage_opamp_dummy_magic_0.Vb2.n27 two_stage_opamp_dummy_magic_0.Vb2.n26 139.077
R6957 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n23 134.577
R6958 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n22 104.781
R6959 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t8 62.5402
R6960 two_stage_opamp_dummy_magic_0.Vb2.n0 two_stage_opamp_dummy_magic_0.Vb2.t1 62.5402
R6961 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.n18 47.1294
R6962 two_stage_opamp_dummy_magic_0.Vb2.n19 two_stage_opamp_dummy_magic_0.Vb2.n14 47.1294
R6963 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n9 47.1294
R6964 two_stage_opamp_dummy_magic_0.Vb2.n10 two_stage_opamp_dummy_magic_0.Vb2.n5 47.1294
R6965 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.t2 24.0005
R6966 two_stage_opamp_dummy_magic_0.Vb2.n25 two_stage_opamp_dummy_magic_0.Vb2.t9 24.0005
R6967 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t6 24.0005
R6968 two_stage_opamp_dummy_magic_0.Vb2.n23 two_stage_opamp_dummy_magic_0.Vb2.t3 24.0005
R6969 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.t10 24.0005
R6970 two_stage_opamp_dummy_magic_0.Vb2.n24 two_stage_opamp_dummy_magic_0.Vb2.t4 24.0005
R6971 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t7 24.0005
R6972 two_stage_opamp_dummy_magic_0.Vb2.n26 two_stage_opamp_dummy_magic_0.Vb2.t5 24.0005
R6973 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n1 18.0505
R6974 two_stage_opamp_dummy_magic_0.Vb2.n21 two_stage_opamp_dummy_magic_0.Vb2.n20 13.0943
R6975 two_stage_opamp_dummy_magic_0.Vb2.n29 two_stage_opamp_dummy_magic_0.Vb2.n28 4.5005
R6976 two_stage_opamp_dummy_magic_0.Vb2.n22 two_stage_opamp_dummy_magic_0.Vb2.n21 4.34425
R6977 bgr_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb2.n29 1.46925
R6978 two_stage_opamp_dummy_magic_0.Vb2.n28 two_stage_opamp_dummy_magic_0.Vb2.n27 0.563
R6979 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n4 4020
R6980 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.n4 4020
R6981 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n10 4020
R6982 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.n10 4020
R6983 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t35 660.109
R6984 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.t32 660.109
R6985 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n14 422.401
R6986 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n3 422.401
R6987 two_stage_opamp_dummy_magic_0.VD4.t36 two_stage_opamp_dummy_magic_0.VD4.n11 239.915
R6988 two_stage_opamp_dummy_magic_0.VD4.n13 two_stage_opamp_dummy_magic_0.VD4.t33 239.915
R6989 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n8 230.4
R6990 two_stage_opamp_dummy_magic_0.VD4.n9 two_stage_opamp_dummy_magic_0.VD4.n6 230.4
R6991 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.n6 198.4
R6992 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n3 198.4
R6993 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.n0 160.428
R6994 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n23 160.427
R6995 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n21 159.804
R6996 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.n19 159.803
R6997 two_stage_opamp_dummy_magic_0.VD4.n2 two_stage_opamp_dummy_magic_0.VD4.n1 159.803
R6998 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n32 159.802
R6999 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n30 159.802
R7000 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.n28 159.802
R7001 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n26 159.802
R7002 two_stage_opamp_dummy_magic_0.VD4.n25 two_stage_opamp_dummy_magic_0.VD4.n24 159.802
R7003 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n16 155.303
R7004 two_stage_opamp_dummy_magic_0.VD4.n7 two_stage_opamp_dummy_magic_0.VD4.t37 155.125
R7005 two_stage_opamp_dummy_magic_0.VD4.n5 two_stage_opamp_dummy_magic_0.VD4.t34 155.125
R7006 two_stage_opamp_dummy_magic_0.VD4.t9 two_stage_opamp_dummy_magic_0.VD4.t36 98.2764
R7007 two_stage_opamp_dummy_magic_0.VD4.t13 two_stage_opamp_dummy_magic_0.VD4.t9 98.2764
R7008 two_stage_opamp_dummy_magic_0.VD4.t17 two_stage_opamp_dummy_magic_0.VD4.t13 98.2764
R7009 two_stage_opamp_dummy_magic_0.VD4.t1 two_stage_opamp_dummy_magic_0.VD4.t17 98.2764
R7010 two_stage_opamp_dummy_magic_0.VD4.t5 two_stage_opamp_dummy_magic_0.VD4.t1 98.2764
R7011 two_stage_opamp_dummy_magic_0.VD4.t11 two_stage_opamp_dummy_magic_0.VD4.t7 98.2764
R7012 two_stage_opamp_dummy_magic_0.VD4.t15 two_stage_opamp_dummy_magic_0.VD4.t11 98.2764
R7013 two_stage_opamp_dummy_magic_0.VD4.t19 two_stage_opamp_dummy_magic_0.VD4.t15 98.2764
R7014 two_stage_opamp_dummy_magic_0.VD4.t3 two_stage_opamp_dummy_magic_0.VD4.t19 98.2764
R7015 two_stage_opamp_dummy_magic_0.VD4.t33 two_stage_opamp_dummy_magic_0.VD4.t3 98.2764
R7016 two_stage_opamp_dummy_magic_0.VD4.n14 two_stage_opamp_dummy_magic_0.VD4.n13 92.5005
R7017 two_stage_opamp_dummy_magic_0.VD4.n10 two_stage_opamp_dummy_magic_0.VD4.n9 92.5005
R7018 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n10 92.5005
R7019 two_stage_opamp_dummy_magic_0.VD4.n11 two_stage_opamp_dummy_magic_0.VD4.n3 92.5005
R7020 two_stage_opamp_dummy_magic_0.VD4.n15 two_stage_opamp_dummy_magic_0.VD4.n4 92.5005
R7021 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.n4 92.5005
R7022 two_stage_opamp_dummy_magic_0.VD4.n12 two_stage_opamp_dummy_magic_0.VD4.t5 49.1384
R7023 two_stage_opamp_dummy_magic_0.VD4.t7 two_stage_opamp_dummy_magic_0.VD4.n12 49.1384
R7024 two_stage_opamp_dummy_magic_0.VD4.n8 two_stage_opamp_dummy_magic_0.VD4.n7 21.3338
R7025 two_stage_opamp_dummy_magic_0.VD4.n6 two_stage_opamp_dummy_magic_0.VD4.n5 21.3338
R7026 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.t29 11.2576
R7027 two_stage_opamp_dummy_magic_0.VD4.n32 two_stage_opamp_dummy_magic_0.VD4.t27 11.2576
R7028 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.t0 11.2576
R7029 two_stage_opamp_dummy_magic_0.VD4.n30 two_stage_opamp_dummy_magic_0.VD4.t26 11.2576
R7030 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t21 11.2576
R7031 two_stage_opamp_dummy_magic_0.VD4.n28 two_stage_opamp_dummy_magic_0.VD4.t28 11.2576
R7032 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t31 11.2576
R7033 two_stage_opamp_dummy_magic_0.VD4.n26 two_stage_opamp_dummy_magic_0.VD4.t24 11.2576
R7034 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.t23 11.2576
R7035 two_stage_opamp_dummy_magic_0.VD4.n24 two_stage_opamp_dummy_magic_0.VD4.t22 11.2576
R7036 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t25 11.2576
R7037 two_stage_opamp_dummy_magic_0.VD4.n23 two_stage_opamp_dummy_magic_0.VD4.t30 11.2576
R7038 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.t12 11.2576
R7039 two_stage_opamp_dummy_magic_0.VD4.n19 two_stage_opamp_dummy_magic_0.VD4.t16 11.2576
R7040 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t6 11.2576
R7041 two_stage_opamp_dummy_magic_0.VD4.n16 two_stage_opamp_dummy_magic_0.VD4.t8 11.2576
R7042 two_stage_opamp_dummy_magic_0.VD4.n1 two_stage_opamp_dummy_magic_0.VD4.t18 11.2576
R7043 two_stage_opamp_dummy_magic_0.VD4.n1 two_stage_opamp_dummy_magic_0.VD4.t2 11.2576
R7044 two_stage_opamp_dummy_magic_0.VD4.n0 two_stage_opamp_dummy_magic_0.VD4.t10 11.2576
R7045 two_stage_opamp_dummy_magic_0.VD4.n0 two_stage_opamp_dummy_magic_0.VD4.t14 11.2576
R7046 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.t20 11.2576
R7047 two_stage_opamp_dummy_magic_0.VD4.n21 two_stage_opamp_dummy_magic_0.VD4.t4 11.2576
R7048 two_stage_opamp_dummy_magic_0.VD4.n17 two_stage_opamp_dummy_magic_0.VD4.n15 9.5505
R7049 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.VD4.n33 8.3755
R7050 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.VD4.n22 6.063
R7051 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.n17 4.5005
R7052 two_stage_opamp_dummy_magic_0.VD4.n27 two_stage_opamp_dummy_magic_0.VD4.n25 0.6255
R7053 two_stage_opamp_dummy_magic_0.VD4.n29 two_stage_opamp_dummy_magic_0.VD4.n27 0.6255
R7054 two_stage_opamp_dummy_magic_0.VD4.n31 two_stage_opamp_dummy_magic_0.VD4.n29 0.6255
R7055 two_stage_opamp_dummy_magic_0.VD4.n33 two_stage_opamp_dummy_magic_0.VD4.n31 0.6255
R7056 two_stage_opamp_dummy_magic_0.VD4.n18 two_stage_opamp_dummy_magic_0.VD4.n2 0.6255
R7057 two_stage_opamp_dummy_magic_0.VD4.n20 two_stage_opamp_dummy_magic_0.VD4.n18 0.6255
R7058 two_stage_opamp_dummy_magic_0.VD4.n22 two_stage_opamp_dummy_magic_0.VD4.n20 0.6255
R7059 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t29 1172.87
R7060 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t34 1172.87
R7061 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.t51 996.134
R7062 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.t39 996.134
R7063 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.t26 996.134
R7064 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.t44 996.134
R7065 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.t25 996.134
R7066 two_stage_opamp_dummy_magic_0.X.n13 two_stage_opamp_dummy_magic_0.X.t43 996.134
R7067 two_stage_opamp_dummy_magic_0.X.n11 two_stage_opamp_dummy_magic_0.X.t49 996.134
R7068 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.t36 996.134
R7069 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t32 690.867
R7070 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.t37 690.867
R7071 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.t28 530.201
R7072 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t33 530.201
R7073 two_stage_opamp_dummy_magic_0.X.n48 two_stage_opamp_dummy_magic_0.X.t46 514.134
R7074 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.t30 514.134
R7075 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.t47 514.134
R7076 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.t31 514.134
R7077 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.t45 514.134
R7078 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.t27 514.134
R7079 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.t40 514.134
R7080 two_stage_opamp_dummy_magic_0.X.n41 two_stage_opamp_dummy_magic_0.X.t52 514.134
R7081 two_stage_opamp_dummy_magic_0.X.n39 two_stage_opamp_dummy_magic_0.X.t41 353.467
R7082 two_stage_opamp_dummy_magic_0.X.n32 two_stage_opamp_dummy_magic_0.X.t48 353.467
R7083 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.t35 353.467
R7084 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.t50 353.467
R7085 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.t38 353.467
R7086 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.t54 353.467
R7087 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.t42 353.467
R7088 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.t53 353.467
R7089 two_stage_opamp_dummy_magic_0.X.n18 two_stage_opamp_dummy_magic_0.X.n17 176.733
R7090 two_stage_opamp_dummy_magic_0.X.n17 two_stage_opamp_dummy_magic_0.X.n16 176.733
R7091 two_stage_opamp_dummy_magic_0.X.n16 two_stage_opamp_dummy_magic_0.X.n15 176.733
R7092 two_stage_opamp_dummy_magic_0.X.n15 two_stage_opamp_dummy_magic_0.X.n14 176.733
R7093 two_stage_opamp_dummy_magic_0.X.n14 two_stage_opamp_dummy_magic_0.X.n13 176.733
R7094 two_stage_opamp_dummy_magic_0.X.n12 two_stage_opamp_dummy_magic_0.X.n11 176.733
R7095 two_stage_opamp_dummy_magic_0.X.n33 two_stage_opamp_dummy_magic_0.X.n32 176.733
R7096 two_stage_opamp_dummy_magic_0.X.n34 two_stage_opamp_dummy_magic_0.X.n33 176.733
R7097 two_stage_opamp_dummy_magic_0.X.n35 two_stage_opamp_dummy_magic_0.X.n34 176.733
R7098 two_stage_opamp_dummy_magic_0.X.n36 two_stage_opamp_dummy_magic_0.X.n35 176.733
R7099 two_stage_opamp_dummy_magic_0.X.n37 two_stage_opamp_dummy_magic_0.X.n36 176.733
R7100 two_stage_opamp_dummy_magic_0.X.n38 two_stage_opamp_dummy_magic_0.X.n37 176.733
R7101 two_stage_opamp_dummy_magic_0.X.n42 two_stage_opamp_dummy_magic_0.X.n41 176.733
R7102 two_stage_opamp_dummy_magic_0.X.n43 two_stage_opamp_dummy_magic_0.X.n42 176.733
R7103 two_stage_opamp_dummy_magic_0.X.n44 two_stage_opamp_dummy_magic_0.X.n43 176.733
R7104 two_stage_opamp_dummy_magic_0.X.n45 two_stage_opamp_dummy_magic_0.X.n44 176.733
R7105 two_stage_opamp_dummy_magic_0.X.n46 two_stage_opamp_dummy_magic_0.X.n45 176.733
R7106 two_stage_opamp_dummy_magic_0.X.n47 two_stage_opamp_dummy_magic_0.X.n46 176.733
R7107 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.n19 166.436
R7108 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n40 161.843
R7109 two_stage_opamp_dummy_magic_0.X.n50 two_stage_opamp_dummy_magic_0.X.n49 161.718
R7110 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.n21 160.427
R7111 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n28 159.802
R7112 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n26 159.802
R7113 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n24 159.802
R7114 two_stage_opamp_dummy_magic_0.X.n23 two_stage_opamp_dummy_magic_0.X.n22 159.802
R7115 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n30 155.302
R7116 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n2 114.689
R7117 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.n1 114.689
R7118 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n7 114.126
R7119 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n5 114.126
R7120 two_stage_opamp_dummy_magic_0.X.n4 two_stage_opamp_dummy_magic_0.X.n3 114.126
R7121 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n0 109.626
R7122 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n18 51.9494
R7123 two_stage_opamp_dummy_magic_0.X.n19 two_stage_opamp_dummy_magic_0.X.n12 51.9494
R7124 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n39 51.9494
R7125 two_stage_opamp_dummy_magic_0.X.n40 two_stage_opamp_dummy_magic_0.X.n38 51.9494
R7126 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.n48 51.9494
R7127 two_stage_opamp_dummy_magic_0.X.n49 two_stage_opamp_dummy_magic_0.X.n47 51.9494
R7128 two_stage_opamp_dummy_magic_0.X.n20 two_stage_opamp_dummy_magic_0.X.t12 49.3037
R7129 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n31 17.4067
R7130 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t15 16.0005
R7131 two_stage_opamp_dummy_magic_0.X.n7 two_stage_opamp_dummy_magic_0.X.t11 16.0005
R7132 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t10 16.0005
R7133 two_stage_opamp_dummy_magic_0.X.n5 two_stage_opamp_dummy_magic_0.X.t13 16.0005
R7134 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t16 16.0005
R7135 two_stage_opamp_dummy_magic_0.X.n3 two_stage_opamp_dummy_magic_0.X.t23 16.0005
R7136 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.t21 16.0005
R7137 two_stage_opamp_dummy_magic_0.X.n2 two_stage_opamp_dummy_magic_0.X.t19 16.0005
R7138 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t20 16.0005
R7139 two_stage_opamp_dummy_magic_0.X.n1 two_stage_opamp_dummy_magic_0.X.t22 16.0005
R7140 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t17 16.0005
R7141 two_stage_opamp_dummy_magic_0.X.n0 two_stage_opamp_dummy_magic_0.X.t14 16.0005
R7142 two_stage_opamp_dummy_magic_0.X.n51 two_stage_opamp_dummy_magic_0.X.n50 13.9693
R7143 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.t18 11.2576
R7144 two_stage_opamp_dummy_magic_0.X.n30 two_stage_opamp_dummy_magic_0.X.t1 11.2576
R7145 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.t0 11.2576
R7146 two_stage_opamp_dummy_magic_0.X.n28 two_stage_opamp_dummy_magic_0.X.t7 11.2576
R7147 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t5 11.2576
R7148 two_stage_opamp_dummy_magic_0.X.n26 two_stage_opamp_dummy_magic_0.X.t4 11.2576
R7149 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t3 11.2576
R7150 two_stage_opamp_dummy_magic_0.X.n24 two_stage_opamp_dummy_magic_0.X.t2 11.2576
R7151 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.t8 11.2576
R7152 two_stage_opamp_dummy_magic_0.X.n22 two_stage_opamp_dummy_magic_0.X.t9 11.2576
R7153 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.t6 11.2576
R7154 two_stage_opamp_dummy_magic_0.X.n21 two_stage_opamp_dummy_magic_0.X.t24 11.2576
R7155 two_stage_opamp_dummy_magic_0.X.n53 two_stage_opamp_dummy_magic_0.X.n52 7.5005
R7156 two_stage_opamp_dummy_magic_0.X.n31 two_stage_opamp_dummy_magic_0.X.n29 5.1255
R7157 two_stage_opamp_dummy_magic_0.X.n10 two_stage_opamp_dummy_magic_0.X.n9 4.5005
R7158 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n51 4.5005
R7159 two_stage_opamp_dummy_magic_0.X.n52 two_stage_opamp_dummy_magic_0.X.n20 3.40675
R7160 two_stage_opamp_dummy_magic_0.X.n53 two_stage_opamp_dummy_magic_0.X.n10 1.71925
R7161 two_stage_opamp_dummy_magic_0.X.n25 two_stage_opamp_dummy_magic_0.X.n23 0.6255
R7162 two_stage_opamp_dummy_magic_0.X.n27 two_stage_opamp_dummy_magic_0.X.n25 0.6255
R7163 two_stage_opamp_dummy_magic_0.X.n29 two_stage_opamp_dummy_magic_0.X.n27 0.6255
R7164 two_stage_opamp_dummy_magic_0.X.n6 two_stage_opamp_dummy_magic_0.X.n4 0.563
R7165 two_stage_opamp_dummy_magic_0.X.n8 two_stage_opamp_dummy_magic_0.X.n6 0.563
R7166 two_stage_opamp_dummy_magic_0.X.n9 two_stage_opamp_dummy_magic_0.X.n8 0.563
R7167 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.X.n53 0.063
R7168 two_stage_opamp_dummy_magic_0.VOUT-.n2 two_stage_opamp_dummy_magic_0.VOUT-.n0 145.989
R7169 two_stage_opamp_dummy_magic_0.VOUT-.n8 two_stage_opamp_dummy_magic_0.VOUT-.n7 145.989
R7170 two_stage_opamp_dummy_magic_0.VOUT-.n6 two_stage_opamp_dummy_magic_0.VOUT-.n5 145.427
R7171 two_stage_opamp_dummy_magic_0.VOUT-.n4 two_stage_opamp_dummy_magic_0.VOUT-.n3 145.427
R7172 two_stage_opamp_dummy_magic_0.VOUT-.n2 two_stage_opamp_dummy_magic_0.VOUT-.n1 145.427
R7173 two_stage_opamp_dummy_magic_0.VOUT-.n10 two_stage_opamp_dummy_magic_0.VOUT-.n9 140.927
R7174 two_stage_opamp_dummy_magic_0.VOUT-.t0 two_stage_opamp_dummy_magic_0.VOUT-.n96 113.192
R7175 two_stage_opamp_dummy_magic_0.VOUT-.n93 two_stage_opamp_dummy_magic_0.VOUT-.n91 95.7303
R7176 two_stage_opamp_dummy_magic_0.VOUT-.n95 two_stage_opamp_dummy_magic_0.VOUT-.n94 94.6053
R7177 two_stage_opamp_dummy_magic_0.VOUT-.n93 two_stage_opamp_dummy_magic_0.VOUT-.n92 94.6053
R7178 two_stage_opamp_dummy_magic_0.VOUT-.n90 two_stage_opamp_dummy_magic_0.VOUT-.n10 20.688
R7179 two_stage_opamp_dummy_magic_0.VOUT-.n90 two_stage_opamp_dummy_magic_0.VOUT-.n89 11.7059
R7180 two_stage_opamp_dummy_magic_0.VOUT-.n96 two_stage_opamp_dummy_magic_0.VOUT-.n90 11.063
R7181 two_stage_opamp_dummy_magic_0.VOUT-.n9 two_stage_opamp_dummy_magic_0.VOUT-.t13 6.56717
R7182 two_stage_opamp_dummy_magic_0.VOUT-.n9 two_stage_opamp_dummy_magic_0.VOUT-.t7 6.56717
R7183 two_stage_opamp_dummy_magic_0.VOUT-.n7 two_stage_opamp_dummy_magic_0.VOUT-.t11 6.56717
R7184 two_stage_opamp_dummy_magic_0.VOUT-.n7 two_stage_opamp_dummy_magic_0.VOUT-.t16 6.56717
R7185 two_stage_opamp_dummy_magic_0.VOUT-.n5 two_stage_opamp_dummy_magic_0.VOUT-.t12 6.56717
R7186 two_stage_opamp_dummy_magic_0.VOUT-.n5 two_stage_opamp_dummy_magic_0.VOUT-.t6 6.56717
R7187 two_stage_opamp_dummy_magic_0.VOUT-.n3 two_stage_opamp_dummy_magic_0.VOUT-.t4 6.56717
R7188 two_stage_opamp_dummy_magic_0.VOUT-.n3 two_stage_opamp_dummy_magic_0.VOUT-.t8 6.56717
R7189 two_stage_opamp_dummy_magic_0.VOUT-.n1 two_stage_opamp_dummy_magic_0.VOUT-.t5 6.56717
R7190 two_stage_opamp_dummy_magic_0.VOUT-.n1 two_stage_opamp_dummy_magic_0.VOUT-.t9 6.56717
R7191 two_stage_opamp_dummy_magic_0.VOUT-.n0 two_stage_opamp_dummy_magic_0.VOUT-.t15 6.56717
R7192 two_stage_opamp_dummy_magic_0.VOUT-.n0 two_stage_opamp_dummy_magic_0.VOUT-.t10 6.56717
R7193 two_stage_opamp_dummy_magic_0.VOUT-.n37 two_stage_opamp_dummy_magic_0.VOUT-.t108 4.8295
R7194 two_stage_opamp_dummy_magic_0.VOUT-.n46 two_stage_opamp_dummy_magic_0.VOUT-.t65 4.8295
R7195 two_stage_opamp_dummy_magic_0.VOUT-.n44 two_stage_opamp_dummy_magic_0.VOUT-.t118 4.8295
R7196 two_stage_opamp_dummy_magic_0.VOUT-.n42 two_stage_opamp_dummy_magic_0.VOUT-.t151 4.8295
R7197 two_stage_opamp_dummy_magic_0.VOUT-.n40 two_stage_opamp_dummy_magic_0.VOUT-.t44 4.8295
R7198 two_stage_opamp_dummy_magic_0.VOUT-.n39 two_stage_opamp_dummy_magic_0.VOUT-.t67 4.8295
R7199 two_stage_opamp_dummy_magic_0.VOUT-.n59 two_stage_opamp_dummy_magic_0.VOUT-.t27 4.8295
R7200 two_stage_opamp_dummy_magic_0.VOUT-.n60 two_stage_opamp_dummy_magic_0.VOUT-.t76 4.8295
R7201 two_stage_opamp_dummy_magic_0.VOUT-.n62 two_stage_opamp_dummy_magic_0.VOUT-.t62 4.8295
R7202 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.t112 4.8295
R7203 two_stage_opamp_dummy_magic_0.VOUT-.n65 two_stage_opamp_dummy_magic_0.VOUT-.t114 4.8295
R7204 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.t99 4.8295
R7205 two_stage_opamp_dummy_magic_0.VOUT-.n68 two_stage_opamp_dummy_magic_0.VOUT-.t74 4.8295
R7206 two_stage_opamp_dummy_magic_0.VOUT-.n69 two_stage_opamp_dummy_magic_0.VOUT-.t55 4.8295
R7207 two_stage_opamp_dummy_magic_0.VOUT-.n71 two_stage_opamp_dummy_magic_0.VOUT-.t109 4.8295
R7208 two_stage_opamp_dummy_magic_0.VOUT-.n72 two_stage_opamp_dummy_magic_0.VOUT-.t91 4.8295
R7209 two_stage_opamp_dummy_magic_0.VOUT-.n74 two_stage_opamp_dummy_magic_0.VOUT-.t68 4.8295
R7210 two_stage_opamp_dummy_magic_0.VOUT-.n75 two_stage_opamp_dummy_magic_0.VOUT-.t52 4.8295
R7211 two_stage_opamp_dummy_magic_0.VOUT-.n77 two_stage_opamp_dummy_magic_0.VOUT-.t29 4.8295
R7212 two_stage_opamp_dummy_magic_0.VOUT-.n78 two_stage_opamp_dummy_magic_0.VOUT-.t153 4.8295
R7213 two_stage_opamp_dummy_magic_0.VOUT-.n80 two_stage_opamp_dummy_magic_0.VOUT-.t63 4.8295
R7214 two_stage_opamp_dummy_magic_0.VOUT-.n81 two_stage_opamp_dummy_magic_0.VOUT-.t46 4.8295
R7215 two_stage_opamp_dummy_magic_0.VOUT-.n83 two_stage_opamp_dummy_magic_0.VOUT-.t22 4.8295
R7216 two_stage_opamp_dummy_magic_0.VOUT-.n84 two_stage_opamp_dummy_magic_0.VOUT-.t146 4.8295
R7217 two_stage_opamp_dummy_magic_0.VOUT-.n11 two_stage_opamp_dummy_magic_0.VOUT-.t117 4.8295
R7218 two_stage_opamp_dummy_magic_0.VOUT-.n13 two_stage_opamp_dummy_magic_0.VOUT-.t72 4.8295
R7219 two_stage_opamp_dummy_magic_0.VOUT-.n25 two_stage_opamp_dummy_magic_0.VOUT-.t37 4.8295
R7220 two_stage_opamp_dummy_magic_0.VOUT-.n26 two_stage_opamp_dummy_magic_0.VOUT-.t20 4.8295
R7221 two_stage_opamp_dummy_magic_0.VOUT-.n28 two_stage_opamp_dummy_magic_0.VOUT-.t79 4.8295
R7222 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.t60 4.8295
R7223 two_stage_opamp_dummy_magic_0.VOUT-.n31 two_stage_opamp_dummy_magic_0.VOUT-.t121 4.8295
R7224 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.t104 4.8295
R7225 two_stage_opamp_dummy_magic_0.VOUT-.n34 two_stage_opamp_dummy_magic_0.VOUT-.t84 4.8295
R7226 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.t66 4.8295
R7227 two_stage_opamp_dummy_magic_0.VOUT-.n86 two_stage_opamp_dummy_magic_0.VOUT-.t123 4.8295
R7228 two_stage_opamp_dummy_magic_0.VOUT-.n48 two_stage_opamp_dummy_magic_0.VOUT-.t95 4.8154
R7229 two_stage_opamp_dummy_magic_0.VOUT-.n49 two_stage_opamp_dummy_magic_0.VOUT-.t70 4.8154
R7230 two_stage_opamp_dummy_magic_0.VOUT-.n50 two_stage_opamp_dummy_magic_0.VOUT-.t110 4.8154
R7231 two_stage_opamp_dummy_magic_0.VOUT-.n51 two_stage_opamp_dummy_magic_0.VOUT-.t145 4.8154
R7232 two_stage_opamp_dummy_magic_0.VOUT-.n48 two_stage_opamp_dummy_magic_0.VOUT-.t32 4.806
R7233 two_stage_opamp_dummy_magic_0.VOUT-.n49 two_stage_opamp_dummy_magic_0.VOUT-.t150 4.806
R7234 two_stage_opamp_dummy_magic_0.VOUT-.n50 two_stage_opamp_dummy_magic_0.VOUT-.t50 4.806
R7235 two_stage_opamp_dummy_magic_0.VOUT-.n51 two_stage_opamp_dummy_magic_0.VOUT-.t87 4.806
R7236 two_stage_opamp_dummy_magic_0.VOUT-.n52 two_stage_opamp_dummy_magic_0.VOUT-.t125 4.806
R7237 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.t105 4.806
R7238 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.t140 4.806
R7239 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.t36 4.806
R7240 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.t156 4.806
R7241 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.t53 4.806
R7242 two_stage_opamp_dummy_magic_0.VOUT-.n14 two_stage_opamp_dummy_magic_0.VOUT-.t73 4.806
R7243 two_stage_opamp_dummy_magic_0.VOUT-.n15 two_stage_opamp_dummy_magic_0.VOUT-.t116 4.806
R7244 two_stage_opamp_dummy_magic_0.VOUT-.n16 two_stage_opamp_dummy_magic_0.VOUT-.t64 4.806
R7245 two_stage_opamp_dummy_magic_0.VOUT-.n17 two_stage_opamp_dummy_magic_0.VOUT-.t154 4.806
R7246 two_stage_opamp_dummy_magic_0.VOUT-.n18 two_stage_opamp_dummy_magic_0.VOUT-.t106 4.806
R7247 two_stage_opamp_dummy_magic_0.VOUT-.n19 two_stage_opamp_dummy_magic_0.VOUT-.t143 4.806
R7248 two_stage_opamp_dummy_magic_0.VOUT-.n20 two_stage_opamp_dummy_magic_0.VOUT-.t96 4.806
R7249 two_stage_opamp_dummy_magic_0.VOUT-.n21 two_stage_opamp_dummy_magic_0.VOUT-.t42 4.806
R7250 two_stage_opamp_dummy_magic_0.VOUT-.n22 two_stage_opamp_dummy_magic_0.VOUT-.t86 4.806
R7251 two_stage_opamp_dummy_magic_0.VOUT-.n23 two_stage_opamp_dummy_magic_0.VOUT-.t34 4.806
R7252 two_stage_opamp_dummy_magic_0.VOUT-.n37 two_stage_opamp_dummy_magic_0.VOUT-.t69 4.5005
R7253 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.t90 4.5005
R7254 two_stage_opamp_dummy_magic_0.VOUT-.n46 two_stage_opamp_dummy_magic_0.VOUT-.t80 4.5005
R7255 two_stage_opamp_dummy_magic_0.VOUT-.n47 two_stage_opamp_dummy_magic_0.VOUT-.t43 4.5005
R7256 two_stage_opamp_dummy_magic_0.VOUT-.n44 two_stage_opamp_dummy_magic_0.VOUT-.t56 4.5005
R7257 two_stage_opamp_dummy_magic_0.VOUT-.n45 two_stage_opamp_dummy_magic_0.VOUT-.t21 4.5005
R7258 two_stage_opamp_dummy_magic_0.VOUT-.n42 two_stage_opamp_dummy_magic_0.VOUT-.t98 4.5005
R7259 two_stage_opamp_dummy_magic_0.VOUT-.n43 two_stage_opamp_dummy_magic_0.VOUT-.t59 4.5005
R7260 two_stage_opamp_dummy_magic_0.VOUT-.n40 two_stage_opamp_dummy_magic_0.VOUT-.t136 4.5005
R7261 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.t101 4.5005
R7262 two_stage_opamp_dummy_magic_0.VOUT-.n39 two_stage_opamp_dummy_magic_0.VOUT-.t30 4.5005
R7263 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.t51 4.5005
R7264 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.t155 4.5005
R7265 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.t119 4.5005
R7266 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.t139 4.5005
R7267 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.t102 4.5005
R7268 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.t61 4.5005
R7269 two_stage_opamp_dummy_magic_0.VOUT-.n52 two_stage_opamp_dummy_magic_0.VOUT-.t85 4.5005
R7270 two_stage_opamp_dummy_magic_0.VOUT-.n51 two_stage_opamp_dummy_magic_0.VOUT-.t45 4.5005
R7271 two_stage_opamp_dummy_magic_0.VOUT-.n50 two_stage_opamp_dummy_magic_0.VOUT-.t147 4.5005
R7272 two_stage_opamp_dummy_magic_0.VOUT-.n49 two_stage_opamp_dummy_magic_0.VOUT-.t111 4.5005
R7273 two_stage_opamp_dummy_magic_0.VOUT-.n48 two_stage_opamp_dummy_magic_0.VOUT-.t134 4.5005
R7274 two_stage_opamp_dummy_magic_0.VOUT-.n59 two_stage_opamp_dummy_magic_0.VOUT-.t130 4.5005
R7275 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.t152 4.5005
R7276 two_stage_opamp_dummy_magic_0.VOUT-.n60 two_stage_opamp_dummy_magic_0.VOUT-.t115 4.5005
R7277 two_stage_opamp_dummy_magic_0.VOUT-.n62 two_stage_opamp_dummy_magic_0.VOUT-.t23 4.5005
R7278 two_stage_opamp_dummy_magic_0.VOUT-.n64 two_stage_opamp_dummy_magic_0.VOUT-.t47 4.5005
R7279 two_stage_opamp_dummy_magic_0.VOUT-.n63 two_stage_opamp_dummy_magic_0.VOUT-.t148 4.5005
R7280 two_stage_opamp_dummy_magic_0.VOUT-.n65 two_stage_opamp_dummy_magic_0.VOUT-.t78 4.5005
R7281 two_stage_opamp_dummy_magic_0.VOUT-.n67 two_stage_opamp_dummy_magic_0.VOUT-.t26 4.5005
R7282 two_stage_opamp_dummy_magic_0.VOUT-.n66 two_stage_opamp_dummy_magic_0.VOUT-.t132 4.5005
R7283 two_stage_opamp_dummy_magic_0.VOUT-.n68 two_stage_opamp_dummy_magic_0.VOUT-.t39 4.5005
R7284 two_stage_opamp_dummy_magic_0.VOUT-.n70 two_stage_opamp_dummy_magic_0.VOUT-.t128 4.5005
R7285 two_stage_opamp_dummy_magic_0.VOUT-.n69 two_stage_opamp_dummy_magic_0.VOUT-.t92 4.5005
R7286 two_stage_opamp_dummy_magic_0.VOUT-.n71 two_stage_opamp_dummy_magic_0.VOUT-.t71 4.5005
R7287 two_stage_opamp_dummy_magic_0.VOUT-.n73 two_stage_opamp_dummy_magic_0.VOUT-.t19 4.5005
R7288 two_stage_opamp_dummy_magic_0.VOUT-.n72 two_stage_opamp_dummy_magic_0.VOUT-.t126 4.5005
R7289 two_stage_opamp_dummy_magic_0.VOUT-.n74 two_stage_opamp_dummy_magic_0.VOUT-.t33 4.5005
R7290 two_stage_opamp_dummy_magic_0.VOUT-.n76 two_stage_opamp_dummy_magic_0.VOUT-.t122 4.5005
R7291 two_stage_opamp_dummy_magic_0.VOUT-.n75 two_stage_opamp_dummy_magic_0.VOUT-.t88 4.5005
R7292 two_stage_opamp_dummy_magic_0.VOUT-.n77 two_stage_opamp_dummy_magic_0.VOUT-.t135 4.5005
R7293 two_stage_opamp_dummy_magic_0.VOUT-.n79 two_stage_opamp_dummy_magic_0.VOUT-.t82 4.5005
R7294 two_stage_opamp_dummy_magic_0.VOUT-.n78 two_stage_opamp_dummy_magic_0.VOUT-.t48 4.5005
R7295 two_stage_opamp_dummy_magic_0.VOUT-.n80 two_stage_opamp_dummy_magic_0.VOUT-.t28 4.5005
R7296 two_stage_opamp_dummy_magic_0.VOUT-.n82 two_stage_opamp_dummy_magic_0.VOUT-.t120 4.5005
R7297 two_stage_opamp_dummy_magic_0.VOUT-.n81 two_stage_opamp_dummy_magic_0.VOUT-.t81 4.5005
R7298 two_stage_opamp_dummy_magic_0.VOUT-.n83 two_stage_opamp_dummy_magic_0.VOUT-.t129 4.5005
R7299 two_stage_opamp_dummy_magic_0.VOUT-.n85 two_stage_opamp_dummy_magic_0.VOUT-.t77 4.5005
R7300 two_stage_opamp_dummy_magic_0.VOUT-.n84 two_stage_opamp_dummy_magic_0.VOUT-.t40 4.5005
R7301 two_stage_opamp_dummy_magic_0.VOUT-.n11 two_stage_opamp_dummy_magic_0.VOUT-.t25 4.5005
R7302 two_stage_opamp_dummy_magic_0.VOUT-.n12 two_stage_opamp_dummy_magic_0.VOUT-.t124 4.5005
R7303 two_stage_opamp_dummy_magic_0.VOUT-.n13 two_stage_opamp_dummy_magic_0.VOUT-.t38 4.5005
R7304 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.t127 4.5005
R7305 two_stage_opamp_dummy_magic_0.VOUT-.n23 two_stage_opamp_dummy_magic_0.VOUT-.t94 4.5005
R7306 two_stage_opamp_dummy_magic_0.VOUT-.n22 two_stage_opamp_dummy_magic_0.VOUT-.t54 4.5005
R7307 two_stage_opamp_dummy_magic_0.VOUT-.n21 two_stage_opamp_dummy_magic_0.VOUT-.t144 4.5005
R7308 two_stage_opamp_dummy_magic_0.VOUT-.n20 two_stage_opamp_dummy_magic_0.VOUT-.t113 4.5005
R7309 two_stage_opamp_dummy_magic_0.VOUT-.n19 two_stage_opamp_dummy_magic_0.VOUT-.t75 4.5005
R7310 two_stage_opamp_dummy_magic_0.VOUT-.n18 two_stage_opamp_dummy_magic_0.VOUT-.t24 4.5005
R7311 two_stage_opamp_dummy_magic_0.VOUT-.n17 two_stage_opamp_dummy_magic_0.VOUT-.t131 4.5005
R7312 two_stage_opamp_dummy_magic_0.VOUT-.n16 two_stage_opamp_dummy_magic_0.VOUT-.t97 4.5005
R7313 two_stage_opamp_dummy_magic_0.VOUT-.n15 two_stage_opamp_dummy_magic_0.VOUT-.t58 4.5005
R7314 two_stage_opamp_dummy_magic_0.VOUT-.n14 two_stage_opamp_dummy_magic_0.VOUT-.t149 4.5005
R7315 two_stage_opamp_dummy_magic_0.VOUT-.n25 two_stage_opamp_dummy_magic_0.VOUT-.t142 4.5005
R7316 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.t93 4.5005
R7317 two_stage_opamp_dummy_magic_0.VOUT-.n26 two_stage_opamp_dummy_magic_0.VOUT-.t57 4.5005
R7318 two_stage_opamp_dummy_magic_0.VOUT-.n28 two_stage_opamp_dummy_magic_0.VOUT-.t41 4.5005
R7319 two_stage_opamp_dummy_magic_0.VOUT-.n30 two_stage_opamp_dummy_magic_0.VOUT-.t133 4.5005
R7320 two_stage_opamp_dummy_magic_0.VOUT-.n29 two_stage_opamp_dummy_magic_0.VOUT-.t100 4.5005
R7321 two_stage_opamp_dummy_magic_0.VOUT-.n31 two_stage_opamp_dummy_magic_0.VOUT-.t83 4.5005
R7322 two_stage_opamp_dummy_magic_0.VOUT-.n33 two_stage_opamp_dummy_magic_0.VOUT-.t31 4.5005
R7323 two_stage_opamp_dummy_magic_0.VOUT-.n32 two_stage_opamp_dummy_magic_0.VOUT-.t137 4.5005
R7324 two_stage_opamp_dummy_magic_0.VOUT-.n34 two_stage_opamp_dummy_magic_0.VOUT-.t49 4.5005
R7325 two_stage_opamp_dummy_magic_0.VOUT-.n36 two_stage_opamp_dummy_magic_0.VOUT-.t138 4.5005
R7326 two_stage_opamp_dummy_magic_0.VOUT-.n35 two_stage_opamp_dummy_magic_0.VOUT-.t103 4.5005
R7327 two_stage_opamp_dummy_magic_0.VOUT-.n86 two_stage_opamp_dummy_magic_0.VOUT-.t89 4.5005
R7328 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.t35 4.5005
R7329 two_stage_opamp_dummy_magic_0.VOUT-.n88 two_stage_opamp_dummy_magic_0.VOUT-.t141 4.5005
R7330 two_stage_opamp_dummy_magic_0.VOUT-.n89 two_stage_opamp_dummy_magic_0.VOUT-.t107 4.5005
R7331 two_stage_opamp_dummy_magic_0.VOUT-.n10 two_stage_opamp_dummy_magic_0.VOUT-.n8 4.5005
R7332 two_stage_opamp_dummy_magic_0.VOUT-.n94 two_stage_opamp_dummy_magic_0.VOUT-.t17 3.42907
R7333 two_stage_opamp_dummy_magic_0.VOUT-.n94 two_stage_opamp_dummy_magic_0.VOUT-.t14 3.42907
R7334 two_stage_opamp_dummy_magic_0.VOUT-.n92 two_stage_opamp_dummy_magic_0.VOUT-.t3 3.42907
R7335 two_stage_opamp_dummy_magic_0.VOUT-.n92 two_stage_opamp_dummy_magic_0.VOUT-.t2 3.42907
R7336 two_stage_opamp_dummy_magic_0.VOUT-.n91 two_stage_opamp_dummy_magic_0.VOUT-.t1 3.42907
R7337 two_stage_opamp_dummy_magic_0.VOUT-.n91 two_stage_opamp_dummy_magic_0.VOUT-.t18 3.42907
R7338 two_stage_opamp_dummy_magic_0.VOUT-.n96 two_stage_opamp_dummy_magic_0.VOUT-.n95 2.03175
R7339 two_stage_opamp_dummy_magic_0.VOUT-.n95 two_stage_opamp_dummy_magic_0.VOUT-.n93 1.1255
R7340 two_stage_opamp_dummy_magic_0.VOUT-.n4 two_stage_opamp_dummy_magic_0.VOUT-.n2 0.563
R7341 two_stage_opamp_dummy_magic_0.VOUT-.n6 two_stage_opamp_dummy_magic_0.VOUT-.n4 0.563
R7342 two_stage_opamp_dummy_magic_0.VOUT-.n8 two_stage_opamp_dummy_magic_0.VOUT-.n6 0.563
R7343 two_stage_opamp_dummy_magic_0.VOUT-.n38 two_stage_opamp_dummy_magic_0.VOUT-.n37 0.3295
R7344 two_stage_opamp_dummy_magic_0.VOUT-.n47 two_stage_opamp_dummy_magic_0.VOUT-.n46 0.3295
R7345 two_stage_opamp_dummy_magic_0.VOUT-.n45 two_stage_opamp_dummy_magic_0.VOUT-.n44 0.3295
R7346 two_stage_opamp_dummy_magic_0.VOUT-.n43 two_stage_opamp_dummy_magic_0.VOUT-.n42 0.3295
R7347 two_stage_opamp_dummy_magic_0.VOUT-.n41 two_stage_opamp_dummy_magic_0.VOUT-.n40 0.3295
R7348 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.n39 0.3295
R7349 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.n57 0.3295
R7350 two_stage_opamp_dummy_magic_0.VOUT-.n57 two_stage_opamp_dummy_magic_0.VOUT-.n56 0.3295
R7351 two_stage_opamp_dummy_magic_0.VOUT-.n56 two_stage_opamp_dummy_magic_0.VOUT-.n55 0.3295
R7352 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.n54 0.3295
R7353 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.n53 0.3295
R7354 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.n52 0.3295
R7355 two_stage_opamp_dummy_magic_0.VOUT-.n52 two_stage_opamp_dummy_magic_0.VOUT-.n51 0.3295
R7356 two_stage_opamp_dummy_magic_0.VOUT-.n51 two_stage_opamp_dummy_magic_0.VOUT-.n50 0.3295
R7357 two_stage_opamp_dummy_magic_0.VOUT-.n50 two_stage_opamp_dummy_magic_0.VOUT-.n49 0.3295
R7358 two_stage_opamp_dummy_magic_0.VOUT-.n49 two_stage_opamp_dummy_magic_0.VOUT-.n48 0.3295
R7359 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.n59 0.3295
R7360 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.n60 0.3295
R7361 two_stage_opamp_dummy_magic_0.VOUT-.n64 two_stage_opamp_dummy_magic_0.VOUT-.n62 0.3295
R7362 two_stage_opamp_dummy_magic_0.VOUT-.n64 two_stage_opamp_dummy_magic_0.VOUT-.n63 0.3295
R7363 two_stage_opamp_dummy_magic_0.VOUT-.n67 two_stage_opamp_dummy_magic_0.VOUT-.n65 0.3295
R7364 two_stage_opamp_dummy_magic_0.VOUT-.n67 two_stage_opamp_dummy_magic_0.VOUT-.n66 0.3295
R7365 two_stage_opamp_dummy_magic_0.VOUT-.n70 two_stage_opamp_dummy_magic_0.VOUT-.n68 0.3295
R7366 two_stage_opamp_dummy_magic_0.VOUT-.n70 two_stage_opamp_dummy_magic_0.VOUT-.n69 0.3295
R7367 two_stage_opamp_dummy_magic_0.VOUT-.n73 two_stage_opamp_dummy_magic_0.VOUT-.n71 0.3295
R7368 two_stage_opamp_dummy_magic_0.VOUT-.n73 two_stage_opamp_dummy_magic_0.VOUT-.n72 0.3295
R7369 two_stage_opamp_dummy_magic_0.VOUT-.n76 two_stage_opamp_dummy_magic_0.VOUT-.n74 0.3295
R7370 two_stage_opamp_dummy_magic_0.VOUT-.n76 two_stage_opamp_dummy_magic_0.VOUT-.n75 0.3295
R7371 two_stage_opamp_dummy_magic_0.VOUT-.n79 two_stage_opamp_dummy_magic_0.VOUT-.n77 0.3295
R7372 two_stage_opamp_dummy_magic_0.VOUT-.n79 two_stage_opamp_dummy_magic_0.VOUT-.n78 0.3295
R7373 two_stage_opamp_dummy_magic_0.VOUT-.n82 two_stage_opamp_dummy_magic_0.VOUT-.n80 0.3295
R7374 two_stage_opamp_dummy_magic_0.VOUT-.n82 two_stage_opamp_dummy_magic_0.VOUT-.n81 0.3295
R7375 two_stage_opamp_dummy_magic_0.VOUT-.n85 two_stage_opamp_dummy_magic_0.VOUT-.n83 0.3295
R7376 two_stage_opamp_dummy_magic_0.VOUT-.n85 two_stage_opamp_dummy_magic_0.VOUT-.n84 0.3295
R7377 two_stage_opamp_dummy_magic_0.VOUT-.n12 two_stage_opamp_dummy_magic_0.VOUT-.n11 0.3295
R7378 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.n13 0.3295
R7379 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.n23 0.3295
R7380 two_stage_opamp_dummy_magic_0.VOUT-.n23 two_stage_opamp_dummy_magic_0.VOUT-.n22 0.3295
R7381 two_stage_opamp_dummy_magic_0.VOUT-.n22 two_stage_opamp_dummy_magic_0.VOUT-.n21 0.3295
R7382 two_stage_opamp_dummy_magic_0.VOUT-.n21 two_stage_opamp_dummy_magic_0.VOUT-.n20 0.3295
R7383 two_stage_opamp_dummy_magic_0.VOUT-.n20 two_stage_opamp_dummy_magic_0.VOUT-.n19 0.3295
R7384 two_stage_opamp_dummy_magic_0.VOUT-.n19 two_stage_opamp_dummy_magic_0.VOUT-.n18 0.3295
R7385 two_stage_opamp_dummy_magic_0.VOUT-.n18 two_stage_opamp_dummy_magic_0.VOUT-.n17 0.3295
R7386 two_stage_opamp_dummy_magic_0.VOUT-.n17 two_stage_opamp_dummy_magic_0.VOUT-.n16 0.3295
R7387 two_stage_opamp_dummy_magic_0.VOUT-.n16 two_stage_opamp_dummy_magic_0.VOUT-.n15 0.3295
R7388 two_stage_opamp_dummy_magic_0.VOUT-.n15 two_stage_opamp_dummy_magic_0.VOUT-.n14 0.3295
R7389 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.n25 0.3295
R7390 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.n26 0.3295
R7391 two_stage_opamp_dummy_magic_0.VOUT-.n30 two_stage_opamp_dummy_magic_0.VOUT-.n28 0.3295
R7392 two_stage_opamp_dummy_magic_0.VOUT-.n30 two_stage_opamp_dummy_magic_0.VOUT-.n29 0.3295
R7393 two_stage_opamp_dummy_magic_0.VOUT-.n33 two_stage_opamp_dummy_magic_0.VOUT-.n31 0.3295
R7394 two_stage_opamp_dummy_magic_0.VOUT-.n33 two_stage_opamp_dummy_magic_0.VOUT-.n32 0.3295
R7395 two_stage_opamp_dummy_magic_0.VOUT-.n36 two_stage_opamp_dummy_magic_0.VOUT-.n34 0.3295
R7396 two_stage_opamp_dummy_magic_0.VOUT-.n36 two_stage_opamp_dummy_magic_0.VOUT-.n35 0.3295
R7397 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.n86 0.3295
R7398 two_stage_opamp_dummy_magic_0.VOUT-.n88 two_stage_opamp_dummy_magic_0.VOUT-.n87 0.3295
R7399 two_stage_opamp_dummy_magic_0.VOUT-.n89 two_stage_opamp_dummy_magic_0.VOUT-.n88 0.3295
R7400 two_stage_opamp_dummy_magic_0.VOUT-.n52 two_stage_opamp_dummy_magic_0.VOUT-.n47 0.306
R7401 two_stage_opamp_dummy_magic_0.VOUT-.n53 two_stage_opamp_dummy_magic_0.VOUT-.n45 0.306
R7402 two_stage_opamp_dummy_magic_0.VOUT-.n54 two_stage_opamp_dummy_magic_0.VOUT-.n43 0.306
R7403 two_stage_opamp_dummy_magic_0.VOUT-.n55 two_stage_opamp_dummy_magic_0.VOUT-.n41 0.306
R7404 two_stage_opamp_dummy_magic_0.VOUT-.n58 two_stage_opamp_dummy_magic_0.VOUT-.n38 0.2825
R7405 two_stage_opamp_dummy_magic_0.VOUT-.n61 two_stage_opamp_dummy_magic_0.VOUT-.n58 0.2825
R7406 two_stage_opamp_dummy_magic_0.VOUT-.n64 two_stage_opamp_dummy_magic_0.VOUT-.n61 0.2825
R7407 two_stage_opamp_dummy_magic_0.VOUT-.n67 two_stage_opamp_dummy_magic_0.VOUT-.n64 0.2825
R7408 two_stage_opamp_dummy_magic_0.VOUT-.n70 two_stage_opamp_dummy_magic_0.VOUT-.n67 0.2825
R7409 two_stage_opamp_dummy_magic_0.VOUT-.n73 two_stage_opamp_dummy_magic_0.VOUT-.n70 0.2825
R7410 two_stage_opamp_dummy_magic_0.VOUT-.n76 two_stage_opamp_dummy_magic_0.VOUT-.n73 0.2825
R7411 two_stage_opamp_dummy_magic_0.VOUT-.n79 two_stage_opamp_dummy_magic_0.VOUT-.n76 0.2825
R7412 two_stage_opamp_dummy_magic_0.VOUT-.n82 two_stage_opamp_dummy_magic_0.VOUT-.n79 0.2825
R7413 two_stage_opamp_dummy_magic_0.VOUT-.n85 two_stage_opamp_dummy_magic_0.VOUT-.n82 0.2825
R7414 two_stage_opamp_dummy_magic_0.VOUT-.n24 two_stage_opamp_dummy_magic_0.VOUT-.n12 0.2825
R7415 two_stage_opamp_dummy_magic_0.VOUT-.n27 two_stage_opamp_dummy_magic_0.VOUT-.n24 0.2825
R7416 two_stage_opamp_dummy_magic_0.VOUT-.n30 two_stage_opamp_dummy_magic_0.VOUT-.n27 0.2825
R7417 two_stage_opamp_dummy_magic_0.VOUT-.n33 two_stage_opamp_dummy_magic_0.VOUT-.n30 0.2825
R7418 two_stage_opamp_dummy_magic_0.VOUT-.n36 two_stage_opamp_dummy_magic_0.VOUT-.n33 0.2825
R7419 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.n36 0.2825
R7420 two_stage_opamp_dummy_magic_0.VOUT-.n87 two_stage_opamp_dummy_magic_0.VOUT-.n85 0.2825
R7421 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t16 449.868
R7422 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t21 449.868
R7423 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t13 449.868
R7424 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t17 449.868
R7425 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n0 339.961
R7426 two_stage_opamp_dummy_magic_0.Vb1.n2 two_stage_opamp_dummy_magic_0.Vb1.n1 339.272
R7427 two_stage_opamp_dummy_magic_0.Vb1.n16 two_stage_opamp_dummy_magic_0.Vb1.t6 273.134
R7428 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.t14 273.134
R7429 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.t25 273.134
R7430 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.t20 273.134
R7431 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.t9 273.134
R7432 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.t18 273.134
R7433 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.t23 273.134
R7434 two_stage_opamp_dummy_magic_0.Vb1.n12 two_stage_opamp_dummy_magic_0.Vb1.t11 273.134
R7435 two_stage_opamp_dummy_magic_0.Vb1.n7 two_stage_opamp_dummy_magic_0.Vb1.t24 273.134
R7436 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.t12 273.134
R7437 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.t22 273.134
R7438 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.t10 273.134
R7439 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.t7 273.134
R7440 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.t15 273.134
R7441 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.t19 273.134
R7442 two_stage_opamp_dummy_magic_0.Vb1.n3 two_stage_opamp_dummy_magic_0.Vb1.t8 273.134
R7443 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.t4 184.665
R7444 two_stage_opamp_dummy_magic_0.Vb1.n19 two_stage_opamp_dummy_magic_0.Vb1.n18 176.733
R7445 two_stage_opamp_dummy_magic_0.Vb1.n18 two_stage_opamp_dummy_magic_0.Vb1.n17 176.733
R7446 two_stage_opamp_dummy_magic_0.Vb1.n17 two_stage_opamp_dummy_magic_0.Vb1.n16 176.733
R7447 two_stage_opamp_dummy_magic_0.Vb1.n13 two_stage_opamp_dummy_magic_0.Vb1.n12 176.733
R7448 two_stage_opamp_dummy_magic_0.Vb1.n14 two_stage_opamp_dummy_magic_0.Vb1.n13 176.733
R7449 two_stage_opamp_dummy_magic_0.Vb1.n15 two_stage_opamp_dummy_magic_0.Vb1.n14 176.733
R7450 two_stage_opamp_dummy_magic_0.Vb1.n10 two_stage_opamp_dummy_magic_0.Vb1.n9 176.733
R7451 two_stage_opamp_dummy_magic_0.Vb1.n9 two_stage_opamp_dummy_magic_0.Vb1.n8 176.733
R7452 two_stage_opamp_dummy_magic_0.Vb1.n8 two_stage_opamp_dummy_magic_0.Vb1.n7 176.733
R7453 two_stage_opamp_dummy_magic_0.Vb1.n4 two_stage_opamp_dummy_magic_0.Vb1.n3 176.733
R7454 two_stage_opamp_dummy_magic_0.Vb1.n5 two_stage_opamp_dummy_magic_0.Vb1.n4 176.733
R7455 two_stage_opamp_dummy_magic_0.Vb1.n6 two_stage_opamp_dummy_magic_0.Vb1.n5 176.733
R7456 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n11 171.644
R7457 two_stage_opamp_dummy_magic_0.Vb1.n21 two_stage_opamp_dummy_magic_0.Vb1.n20 165.8
R7458 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n23 99.2817
R7459 two_stage_opamp_dummy_magic_0.Vb1.n22 two_stage_opamp_dummy_magic_0.Vb1.t3 62.0342
R7460 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n19 56.2338
R7461 two_stage_opamp_dummy_magic_0.Vb1.n20 two_stage_opamp_dummy_magic_0.Vb1.n15 56.2338
R7462 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n10 56.2338
R7463 two_stage_opamp_dummy_magic_0.Vb1.n11 two_stage_opamp_dummy_magic_0.Vb1.n6 56.2338
R7464 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t5 39.4005
R7465 two_stage_opamp_dummy_magic_0.Vb1.n1 two_stage_opamp_dummy_magic_0.Vb1.t1 39.4005
R7466 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t2 39.4005
R7467 two_stage_opamp_dummy_magic_0.Vb1.n0 two_stage_opamp_dummy_magic_0.Vb1.t0 39.4005
R7468 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n21 17.1724
R7469 two_stage_opamp_dummy_magic_0.Vb1.n23 two_stage_opamp_dummy_magic_0.Vb1.n22 14.2806
R7470 bgr_0.VB1_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb1.n2 4.46925
R7471 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t25 369.534
R7472 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t24 369.534
R7473 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t15 369.534
R7474 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t11 369.534
R7475 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t17 369.534
R7476 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t16 369.534
R7477 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n6 341.397
R7478 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n9 339.272
R7479 bgr_0.PFET_GATE_10uA.n8 bgr_0.PFET_GATE_10uA.n7 339.272
R7480 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n12 334.772
R7481 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t21 238.322
R7482 bgr_0.PFET_GATE_10uA.n15 bgr_0.PFET_GATE_10uA.t13 238.322
R7483 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.t3 194.895
R7484 bgr_0.PFET_GATE_10uA.n4 bgr_0.PFET_GATE_10uA.t18 192.8
R7485 bgr_0.PFET_GATE_10uA.n3 bgr_0.PFET_GATE_10uA.t10 192.8
R7486 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.t14 192.8
R7487 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.t22 192.8
R7488 bgr_0.PFET_GATE_10uA.n23 bgr_0.PFET_GATE_10uA.t28 192.8
R7489 bgr_0.PFET_GATE_10uA.n18 bgr_0.PFET_GATE_10uA.t19 192.8
R7490 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.t26 192.8
R7491 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.t12 192.8
R7492 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.t20 192.8
R7493 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.t27 192.8
R7494 bgr_0.PFET_GATE_10uA.n1 bgr_0.PFET_GATE_10uA.t29 192.8
R7495 bgr_0.PFET_GATE_10uA.n0 bgr_0.PFET_GATE_10uA.t23 192.8
R7496 bgr_0.PFET_GATE_10uA.n25 bgr_0.PFET_GATE_10uA.n24 176.733
R7497 bgr_0.PFET_GATE_10uA.n24 bgr_0.PFET_GATE_10uA.n23 176.733
R7498 bgr_0.PFET_GATE_10uA.n19 bgr_0.PFET_GATE_10uA.n18 176.733
R7499 bgr_0.PFET_GATE_10uA.n20 bgr_0.PFET_GATE_10uA.n19 176.733
R7500 bgr_0.PFET_GATE_10uA.n21 bgr_0.PFET_GATE_10uA.n20 176.733
R7501 bgr_0.PFET_GATE_10uA.n22 bgr_0.PFET_GATE_10uA.n21 176.733
R7502 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n2 171.321
R7503 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n15 169.394
R7504 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n5 168.166
R7505 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n26 166.071
R7506 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.t7 100.635
R7507 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n4 56.2338
R7508 bgr_0.PFET_GATE_10uA.n5 bgr_0.PFET_GATE_10uA.n3 56.2338
R7509 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n25 56.2338
R7510 bgr_0.PFET_GATE_10uA.n26 bgr_0.PFET_GATE_10uA.n22 56.2338
R7511 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n1 56.2338
R7512 bgr_0.PFET_GATE_10uA.n2 bgr_0.PFET_GATE_10uA.n0 56.2338
R7513 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t5 39.4005
R7514 bgr_0.PFET_GATE_10uA.n12 bgr_0.PFET_GATE_10uA.t9 39.4005
R7515 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t4 39.4005
R7516 bgr_0.PFET_GATE_10uA.n9 bgr_0.PFET_GATE_10uA.t0 39.4005
R7517 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t8 39.4005
R7518 bgr_0.PFET_GATE_10uA.n7 bgr_0.PFET_GATE_10uA.t1 39.4005
R7519 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t2 39.4005
R7520 bgr_0.PFET_GATE_10uA.n6 bgr_0.PFET_GATE_10uA.t6 39.4005
R7521 bgr_0.PFET_GATE_10uA.n17 bgr_0.PFET_GATE_10uA.n16 26.9067
R7522 bgr_0.PFET_GATE_10uA.n14 bgr_0.PFET_GATE_10uA.n13 5.15675
R7523 bgr_0.PFET_GATE_10uA.n13 bgr_0.PFET_GATE_10uA.n11 4.5005
R7524 bgr_0.PFET_GATE_10uA.n16 bgr_0.PFET_GATE_10uA.n14 4.188
R7525 bgr_0.PFET_GATE_10uA bgr_0.PFET_GATE_10uA.n17 3.03175
R7526 bgr_0.PFET_GATE_10uA.n10 bgr_0.PFET_GATE_10uA.n8 2.1255
R7527 bgr_0.PFET_GATE_10uA.n11 bgr_0.PFET_GATE_10uA.n10 2.1255
R7528 a_14520_5068.t0 a_14520_5068.t1 294.339
R7529 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 145.046
R7530 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 134.797
R7531 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 120.629
R7532 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 115.219
R7533 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 97.4009
R7534 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 96.8384
R7535 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 96.8384
R7536 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 96.8384
R7537 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 96.8384
R7538 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 24.0005
R7539 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 24.0005
R7540 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 24.0005
R7541 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 24.0005
R7542 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 8.0005
R7543 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 8.0005
R7544 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 8.0005
R7545 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 8.0005
R7546 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 8.0005
R7547 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 8.0005
R7548 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 8.0005
R7549 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 8.0005
R7550 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 8.0005
R7551 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 8.0005
R7552 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 5.84425
R7553 bgr_0.V_CMFB_S2 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 1.1255
R7554 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 0.563
R7555 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 0.563
R7556 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 0.563
R7557 bgr_0.V_mir1.n20 bgr_0.V_mir1.n19 325.473
R7558 bgr_0.V_mir1.n13 bgr_0.V_mir1.n12 325.473
R7559 bgr_0.V_mir1.n4 bgr_0.V_mir1.n3 325.473
R7560 bgr_0.V_mir1.n16 bgr_0.V_mir1.t22 310.488
R7561 bgr_0.V_mir1.n9 bgr_0.V_mir1.t21 310.488
R7562 bgr_0.V_mir1.n0 bgr_0.V_mir1.t20 310.488
R7563 bgr_0.V_mir1.n7 bgr_0.V_mir1.t14 278.312
R7564 bgr_0.V_mir1.n7 bgr_0.V_mir1.n6 228.939
R7565 bgr_0.V_mir1.n8 bgr_0.V_mir1.n5 224.439
R7566 bgr_0.V_mir1.n18 bgr_0.V_mir1.t10 184.097
R7567 bgr_0.V_mir1.n11 bgr_0.V_mir1.t0 184.097
R7568 bgr_0.V_mir1.n2 bgr_0.V_mir1.t8 184.097
R7569 bgr_0.V_mir1.n17 bgr_0.V_mir1.n16 167.094
R7570 bgr_0.V_mir1.n10 bgr_0.V_mir1.n9 167.094
R7571 bgr_0.V_mir1.n1 bgr_0.V_mir1.n0 167.094
R7572 bgr_0.V_mir1.n13 bgr_0.V_mir1.n11 152
R7573 bgr_0.V_mir1.n4 bgr_0.V_mir1.n2 152
R7574 bgr_0.V_mir1.n19 bgr_0.V_mir1.n18 152
R7575 bgr_0.V_mir1.n16 bgr_0.V_mir1.t19 120.501
R7576 bgr_0.V_mir1.n17 bgr_0.V_mir1.t2 120.501
R7577 bgr_0.V_mir1.n9 bgr_0.V_mir1.t18 120.501
R7578 bgr_0.V_mir1.n10 bgr_0.V_mir1.t4 120.501
R7579 bgr_0.V_mir1.n0 bgr_0.V_mir1.t17 120.501
R7580 bgr_0.V_mir1.n1 bgr_0.V_mir1.t6 120.501
R7581 bgr_0.V_mir1.n6 bgr_0.V_mir1.t16 48.0005
R7582 bgr_0.V_mir1.n6 bgr_0.V_mir1.t12 48.0005
R7583 bgr_0.V_mir1.n5 bgr_0.V_mir1.t15 48.0005
R7584 bgr_0.V_mir1.n5 bgr_0.V_mir1.t13 48.0005
R7585 bgr_0.V_mir1.n18 bgr_0.V_mir1.n17 40.7027
R7586 bgr_0.V_mir1.n11 bgr_0.V_mir1.n10 40.7027
R7587 bgr_0.V_mir1.n2 bgr_0.V_mir1.n1 40.7027
R7588 bgr_0.V_mir1.n12 bgr_0.V_mir1.t1 39.4005
R7589 bgr_0.V_mir1.n12 bgr_0.V_mir1.t5 39.4005
R7590 bgr_0.V_mir1.n3 bgr_0.V_mir1.t9 39.4005
R7591 bgr_0.V_mir1.n3 bgr_0.V_mir1.t7 39.4005
R7592 bgr_0.V_mir1.t11 bgr_0.V_mir1.n20 39.4005
R7593 bgr_0.V_mir1.n20 bgr_0.V_mir1.t3 39.4005
R7594 bgr_0.V_mir1.n15 bgr_0.V_mir1.n4 15.8005
R7595 bgr_0.V_mir1.n19 bgr_0.V_mir1.n15 15.8005
R7596 bgr_0.V_mir1.n14 bgr_0.V_mir1.n13 9.3005
R7597 bgr_0.V_mir1.n8 bgr_0.V_mir1.n7 5.8755
R7598 bgr_0.V_mir1.n15 bgr_0.V_mir1.n14 4.5005
R7599 bgr_0.V_mir1.n14 bgr_0.V_mir1.n8 0.78175
R7600 two_stage_opamp_dummy_magic_0.cap_res_X.t0 two_stage_opamp_dummy_magic_0.cap_res_X.t6 50.0055
R7601 two_stage_opamp_dummy_magic_0.cap_res_X.t23 two_stage_opamp_dummy_magic_0.cap_res_X.t62 0.1603
R7602 two_stage_opamp_dummy_magic_0.cap_res_X.t46 two_stage_opamp_dummy_magic_0.cap_res_X.t87 0.1603
R7603 two_stage_opamp_dummy_magic_0.cap_res_X.t10 two_stage_opamp_dummy_magic_0.cap_res_X.t47 0.1603
R7604 two_stage_opamp_dummy_magic_0.cap_res_X.t112 two_stage_opamp_dummy_magic_0.cap_res_X.t12 0.1603
R7605 two_stage_opamp_dummy_magic_0.cap_res_X.t77 two_stage_opamp_dummy_magic_0.cap_res_X.t92 0.1603
R7606 two_stage_opamp_dummy_magic_0.cap_res_X.t114 two_stage_opamp_dummy_magic_0.cap_res_X.t77 0.1603
R7607 two_stage_opamp_dummy_magic_0.cap_res_X.t72 two_stage_opamp_dummy_magic_0.cap_res_X.t114 0.1603
R7608 two_stage_opamp_dummy_magic_0.cap_res_X.t101 two_stage_opamp_dummy_magic_0.cap_res_X.t39 0.1603
R7609 two_stage_opamp_dummy_magic_0.cap_res_X.t136 two_stage_opamp_dummy_magic_0.cap_res_X.t101 0.1603
R7610 two_stage_opamp_dummy_magic_0.cap_res_X.t96 two_stage_opamp_dummy_magic_0.cap_res_X.t136 0.1603
R7611 two_stage_opamp_dummy_magic_0.cap_res_X.t127 two_stage_opamp_dummy_magic_0.cap_res_X.t90 0.1603
R7612 two_stage_opamp_dummy_magic_0.cap_res_X.t88 two_stage_opamp_dummy_magic_0.cap_res_X.t49 0.1603
R7613 two_stage_opamp_dummy_magic_0.cap_res_X.t42 two_stage_opamp_dummy_magic_0.cap_res_X.t81 0.1603
R7614 two_stage_opamp_dummy_magic_0.cap_res_X.t27 two_stage_opamp_dummy_magic_0.cap_res_X.t130 0.1603
R7615 two_stage_opamp_dummy_magic_0.cap_res_X.t9 two_stage_opamp_dummy_magic_0.cap_res_X.t45 0.1603
R7616 two_stage_opamp_dummy_magic_0.cap_res_X.t134 two_stage_opamp_dummy_magic_0.cap_res_X.t95 0.1603
R7617 two_stage_opamp_dummy_magic_0.cap_res_X.t25 two_stage_opamp_dummy_magic_0.cap_res_X.t58 0.1603
R7618 two_stage_opamp_dummy_magic_0.cap_res_X.t79 two_stage_opamp_dummy_magic_0.cap_res_X.t43 0.1603
R7619 two_stage_opamp_dummy_magic_0.cap_res_X.t65 two_stage_opamp_dummy_magic_0.cap_res_X.t102 0.1603
R7620 two_stage_opamp_dummy_magic_0.cap_res_X.t118 two_stage_opamp_dummy_magic_0.cap_res_X.t83 0.1603
R7621 two_stage_opamp_dummy_magic_0.cap_res_X.t31 two_stage_opamp_dummy_magic_0.cap_res_X.t66 0.1603
R7622 two_stage_opamp_dummy_magic_0.cap_res_X.t86 two_stage_opamp_dummy_magic_0.cap_res_X.t48 0.1603
R7623 two_stage_opamp_dummy_magic_0.cap_res_X.t69 two_stage_opamp_dummy_magic_0.cap_res_X.t105 0.1603
R7624 two_stage_opamp_dummy_magic_0.cap_res_X.t124 two_stage_opamp_dummy_magic_0.cap_res_X.t89 0.1603
R7625 two_stage_opamp_dummy_magic_0.cap_res_X.t109 two_stage_opamp_dummy_magic_0.cap_res_X.t4 0.1603
R7626 two_stage_opamp_dummy_magic_0.cap_res_X.t22 two_stage_opamp_dummy_magic_0.cap_res_X.t128 0.1603
R7627 two_stage_opamp_dummy_magic_0.cap_res_X.t76 two_stage_opamp_dummy_magic_0.cap_res_X.t111 0.1603
R7628 two_stage_opamp_dummy_magic_0.cap_res_X.t129 two_stage_opamp_dummy_magic_0.cap_res_X.t94 0.1603
R7629 two_stage_opamp_dummy_magic_0.cap_res_X.t117 two_stage_opamp_dummy_magic_0.cap_res_X.t11 0.1603
R7630 two_stage_opamp_dummy_magic_0.cap_res_X.t28 two_stage_opamp_dummy_magic_0.cap_res_X.t135 0.1603
R7631 two_stage_opamp_dummy_magic_0.cap_res_X.t16 two_stage_opamp_dummy_magic_0.cap_res_X.t50 0.1603
R7632 two_stage_opamp_dummy_magic_0.cap_res_X.t68 two_stage_opamp_dummy_magic_0.cap_res_X.t34 0.1603
R7633 two_stage_opamp_dummy_magic_0.cap_res_X.t54 two_stage_opamp_dummy_magic_0.cap_res_X.t91 0.1603
R7634 two_stage_opamp_dummy_magic_0.cap_res_X.t108 two_stage_opamp_dummy_magic_0.cap_res_X.t73 0.1603
R7635 two_stage_opamp_dummy_magic_0.cap_res_X.t20 two_stage_opamp_dummy_magic_0.cap_res_X.t53 0.1603
R7636 two_stage_opamp_dummy_magic_0.cap_res_X.t74 two_stage_opamp_dummy_magic_0.cap_res_X.t36 0.1603
R7637 two_stage_opamp_dummy_magic_0.cap_res_X.t57 two_stage_opamp_dummy_magic_0.cap_res_X.t97 0.1603
R7638 two_stage_opamp_dummy_magic_0.cap_res_X.t116 two_stage_opamp_dummy_magic_0.cap_res_X.t78 0.1603
R7639 two_stage_opamp_dummy_magic_0.cap_res_X.t100 two_stage_opamp_dummy_magic_0.cap_res_X.t137 0.1603
R7640 two_stage_opamp_dummy_magic_0.cap_res_X.t15 two_stage_opamp_dummy_magic_0.cap_res_X.t120 0.1603
R7641 two_stage_opamp_dummy_magic_0.cap_res_X.t8 two_stage_opamp_dummy_magic_0.cap_res_X.t84 0.1603
R7642 two_stage_opamp_dummy_magic_0.cap_res_X.t99 two_stage_opamp_dummy_magic_0.cap_res_X.t41 0.1603
R7643 two_stage_opamp_dummy_magic_0.cap_res_X.t60 two_stage_opamp_dummy_magic_0.cap_res_X.t93 0.1603
R7644 two_stage_opamp_dummy_magic_0.cap_res_X.t26 two_stage_opamp_dummy_magic_0.cap_res_X.t3 0.1603
R7645 two_stage_opamp_dummy_magic_0.cap_res_X.t133 two_stage_opamp_dummy_magic_0.cap_res_X.t51 0.1603
R7646 two_stage_opamp_dummy_magic_0.cap_res_X.t82 two_stage_opamp_dummy_magic_0.cap_res_X.t14 0.1603
R7647 two_stage_opamp_dummy_magic_0.cap_res_X.t44 two_stage_opamp_dummy_magic_0.cap_res_X.t61 0.1603
R7648 two_stage_opamp_dummy_magic_0.cap_res_X.t13 two_stage_opamp_dummy_magic_0.cap_res_X.t115 0.1603
R7649 two_stage_opamp_dummy_magic_0.cap_res_X.t103 two_stage_opamp_dummy_magic_0.cap_res_X.t71 0.1603
R7650 two_stage_opamp_dummy_magic_0.cap_res_X.t63 two_stage_opamp_dummy_magic_0.cap_res_X.t123 0.1603
R7651 two_stage_opamp_dummy_magic_0.cap_res_X.t119 two_stage_opamp_dummy_magic_0.cap_res_X.t85 0.1603
R7652 two_stage_opamp_dummy_magic_0.cap_res_X.t132 two_stage_opamp_dummy_magic_0.cap_res_X.t40 0.1603
R7653 two_stage_opamp_dummy_magic_0.cap_res_X.t21 two_stage_opamp_dummy_magic_0.cap_res_X.t113 0.1603
R7654 two_stage_opamp_dummy_magic_0.cap_res_X.t56 two_stage_opamp_dummy_magic_0.cap_res_X.t21 0.1603
R7655 two_stage_opamp_dummy_magic_0.cap_res_X.t18 two_stage_opamp_dummy_magic_0.cap_res_X.t56 0.1603
R7656 two_stage_opamp_dummy_magic_0.cap_res_X.t98 two_stage_opamp_dummy_magic_0.cap_res_X.t55 0.1603
R7657 two_stage_opamp_dummy_magic_0.cap_res_X.t59 two_stage_opamp_dummy_magic_0.cap_res_X.t98 0.1603
R7658 two_stage_opamp_dummy_magic_0.cap_res_X.t6 two_stage_opamp_dummy_magic_0.cap_res_X.t59 0.1603
R7659 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t125 0.159278
R7660 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t7 0.159278
R7661 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t107 0.159278
R7662 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t70 0.159278
R7663 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t32 0.159278
R7664 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t52 0.159278
R7665 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t67 0.159278
R7666 two_stage_opamp_dummy_magic_0.cap_res_X.t30 two_stage_opamp_dummy_magic_0.cap_res_X.n9 0.159278
R7667 two_stage_opamp_dummy_magic_0.cap_res_X.t64 two_stage_opamp_dummy_magic_0.cap_res_X.n10 0.159278
R7668 two_stage_opamp_dummy_magic_0.cap_res_X.t24 two_stage_opamp_dummy_magic_0.cap_res_X.n11 0.159278
R7669 two_stage_opamp_dummy_magic_0.cap_res_X.t126 two_stage_opamp_dummy_magic_0.cap_res_X.n12 0.159278
R7670 two_stage_opamp_dummy_magic_0.cap_res_X.t19 two_stage_opamp_dummy_magic_0.cap_res_X.n13 0.159278
R7671 two_stage_opamp_dummy_magic_0.cap_res_X.t122 two_stage_opamp_dummy_magic_0.cap_res_X.n14 0.159278
R7672 two_stage_opamp_dummy_magic_0.cap_res_X.t80 two_stage_opamp_dummy_magic_0.cap_res_X.n15 0.159278
R7673 two_stage_opamp_dummy_magic_0.cap_res_X.t37 two_stage_opamp_dummy_magic_0.cap_res_X.n16 0.159278
R7674 two_stage_opamp_dummy_magic_0.cap_res_X.t75 two_stage_opamp_dummy_magic_0.cap_res_X.n17 0.159278
R7675 two_stage_opamp_dummy_magic_0.cap_res_X.t35 two_stage_opamp_dummy_magic_0.cap_res_X.n18 0.159278
R7676 two_stage_opamp_dummy_magic_0.cap_res_X.t138 two_stage_opamp_dummy_magic_0.cap_res_X.n19 0.159278
R7677 two_stage_opamp_dummy_magic_0.cap_res_X.t29 two_stage_opamp_dummy_magic_0.cap_res_X.n20 0.159278
R7678 two_stage_opamp_dummy_magic_0.cap_res_X.t131 two_stage_opamp_dummy_magic_0.cap_res_X.n21 0.159278
R7679 two_stage_opamp_dummy_magic_0.cap_res_X.t110 two_stage_opamp_dummy_magic_0.cap_res_X.n22 0.159278
R7680 two_stage_opamp_dummy_magic_0.cap_res_X.t5 two_stage_opamp_dummy_magic_0.cap_res_X.n23 0.159278
R7681 two_stage_opamp_dummy_magic_0.cap_res_X.t106 two_stage_opamp_dummy_magic_0.cap_res_X.n24 0.159278
R7682 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t104 0.159278
R7683 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t1 0.159278
R7684 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t121 0.159278
R7685 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.t17 0.159278
R7686 two_stage_opamp_dummy_magic_0.cap_res_X.t67 two_stage_opamp_dummy_magic_0.cap_res_X.t88 0.137822
R7687 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t127 0.1368
R7688 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t42 0.1368
R7689 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t27 0.1368
R7690 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t9 0.1368
R7691 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t134 0.1368
R7692 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t25 0.1368
R7693 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t79 0.1368
R7694 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t65 0.1368
R7695 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t118 0.1368
R7696 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t31 0.1368
R7697 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t86 0.1368
R7698 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t69 0.1368
R7699 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t124 0.1368
R7700 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t109 0.1368
R7701 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t22 0.1368
R7702 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t76 0.1368
R7703 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t129 0.1368
R7704 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t117 0.1368
R7705 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t28 0.1368
R7706 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t16 0.1368
R7707 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t68 0.1368
R7708 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t54 0.1368
R7709 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t108 0.1368
R7710 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t20 0.1368
R7711 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t74 0.1368
R7712 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t57 0.1368
R7713 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t116 0.1368
R7714 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t100 0.1368
R7715 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t15 0.1368
R7716 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t119 0.1368
R7717 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t132 0.1368
R7718 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t8 0.114322
R7719 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.n29 0.1133
R7720 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.n30 0.1133
R7721 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.n31 0.1133
R7722 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.n32 0.1133
R7723 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.n33 0.1133
R7724 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.n0 0.1133
R7725 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.n1 0.1133
R7726 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.n2 0.1133
R7727 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.n3 0.1133
R7728 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.n4 0.1133
R7729 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.n5 0.1133
R7730 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.n6 0.1133
R7731 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.n7 0.1133
R7732 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.n8 0.1133
R7733 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.n25 0.1133
R7734 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.n26 0.1133
R7735 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.n27 0.1133
R7736 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n28 0.1133
R7737 two_stage_opamp_dummy_magic_0.cap_res_X.n35 two_stage_opamp_dummy_magic_0.cap_res_X.n34 0.1133
R7738 two_stage_opamp_dummy_magic_0.cap_res_X.n29 two_stage_opamp_dummy_magic_0.cap_res_X.t23 0.00152174
R7739 two_stage_opamp_dummy_magic_0.cap_res_X.n30 two_stage_opamp_dummy_magic_0.cap_res_X.t46 0.00152174
R7740 two_stage_opamp_dummy_magic_0.cap_res_X.n31 two_stage_opamp_dummy_magic_0.cap_res_X.t10 0.00152174
R7741 two_stage_opamp_dummy_magic_0.cap_res_X.n32 two_stage_opamp_dummy_magic_0.cap_res_X.t112 0.00152174
R7742 two_stage_opamp_dummy_magic_0.cap_res_X.n33 two_stage_opamp_dummy_magic_0.cap_res_X.t72 0.00152174
R7743 two_stage_opamp_dummy_magic_0.cap_res_X.n34 two_stage_opamp_dummy_magic_0.cap_res_X.t96 0.00152174
R7744 two_stage_opamp_dummy_magic_0.cap_res_X.n0 two_stage_opamp_dummy_magic_0.cap_res_X.t99 0.00152174
R7745 two_stage_opamp_dummy_magic_0.cap_res_X.n1 two_stage_opamp_dummy_magic_0.cap_res_X.t60 0.00152174
R7746 two_stage_opamp_dummy_magic_0.cap_res_X.n2 two_stage_opamp_dummy_magic_0.cap_res_X.t26 0.00152174
R7747 two_stage_opamp_dummy_magic_0.cap_res_X.n3 two_stage_opamp_dummy_magic_0.cap_res_X.t133 0.00152174
R7748 two_stage_opamp_dummy_magic_0.cap_res_X.n4 two_stage_opamp_dummy_magic_0.cap_res_X.t82 0.00152174
R7749 two_stage_opamp_dummy_magic_0.cap_res_X.n5 two_stage_opamp_dummy_magic_0.cap_res_X.t44 0.00152174
R7750 two_stage_opamp_dummy_magic_0.cap_res_X.n6 two_stage_opamp_dummy_magic_0.cap_res_X.t13 0.00152174
R7751 two_stage_opamp_dummy_magic_0.cap_res_X.n7 two_stage_opamp_dummy_magic_0.cap_res_X.t103 0.00152174
R7752 two_stage_opamp_dummy_magic_0.cap_res_X.n8 two_stage_opamp_dummy_magic_0.cap_res_X.t63 0.00152174
R7753 two_stage_opamp_dummy_magic_0.cap_res_X.n9 two_stage_opamp_dummy_magic_0.cap_res_X.t33 0.00152174
R7754 two_stage_opamp_dummy_magic_0.cap_res_X.n10 two_stage_opamp_dummy_magic_0.cap_res_X.t30 0.00152174
R7755 two_stage_opamp_dummy_magic_0.cap_res_X.n11 two_stage_opamp_dummy_magic_0.cap_res_X.t64 0.00152174
R7756 two_stage_opamp_dummy_magic_0.cap_res_X.n12 two_stage_opamp_dummy_magic_0.cap_res_X.t24 0.00152174
R7757 two_stage_opamp_dummy_magic_0.cap_res_X.n13 two_stage_opamp_dummy_magic_0.cap_res_X.t126 0.00152174
R7758 two_stage_opamp_dummy_magic_0.cap_res_X.n14 two_stage_opamp_dummy_magic_0.cap_res_X.t19 0.00152174
R7759 two_stage_opamp_dummy_magic_0.cap_res_X.n15 two_stage_opamp_dummy_magic_0.cap_res_X.t122 0.00152174
R7760 two_stage_opamp_dummy_magic_0.cap_res_X.n16 two_stage_opamp_dummy_magic_0.cap_res_X.t80 0.00152174
R7761 two_stage_opamp_dummy_magic_0.cap_res_X.n17 two_stage_opamp_dummy_magic_0.cap_res_X.t37 0.00152174
R7762 two_stage_opamp_dummy_magic_0.cap_res_X.n18 two_stage_opamp_dummy_magic_0.cap_res_X.t75 0.00152174
R7763 two_stage_opamp_dummy_magic_0.cap_res_X.n19 two_stage_opamp_dummy_magic_0.cap_res_X.t35 0.00152174
R7764 two_stage_opamp_dummy_magic_0.cap_res_X.n20 two_stage_opamp_dummy_magic_0.cap_res_X.t138 0.00152174
R7765 two_stage_opamp_dummy_magic_0.cap_res_X.n21 two_stage_opamp_dummy_magic_0.cap_res_X.t29 0.00152174
R7766 two_stage_opamp_dummy_magic_0.cap_res_X.n22 two_stage_opamp_dummy_magic_0.cap_res_X.t131 0.00152174
R7767 two_stage_opamp_dummy_magic_0.cap_res_X.n23 two_stage_opamp_dummy_magic_0.cap_res_X.t110 0.00152174
R7768 two_stage_opamp_dummy_magic_0.cap_res_X.n24 two_stage_opamp_dummy_magic_0.cap_res_X.t5 0.00152174
R7769 two_stage_opamp_dummy_magic_0.cap_res_X.n25 two_stage_opamp_dummy_magic_0.cap_res_X.t106 0.00152174
R7770 two_stage_opamp_dummy_magic_0.cap_res_X.n26 two_stage_opamp_dummy_magic_0.cap_res_X.t2 0.00152174
R7771 two_stage_opamp_dummy_magic_0.cap_res_X.n27 two_stage_opamp_dummy_magic_0.cap_res_X.t38 0.00152174
R7772 two_stage_opamp_dummy_magic_0.cap_res_X.n28 two_stage_opamp_dummy_magic_0.cap_res_X.t18 0.00152174
R7773 two_stage_opamp_dummy_magic_0.cap_res_X.t55 two_stage_opamp_dummy_magic_0.cap_res_X.n35 0.00152174
R7774 bgr_0.START_UP_NFET1 bgr_0.START_UP_NFET1.t0 141.653
R7775 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 610.534
R7776 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 610.534
R7777 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 433.8
R7778 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 433.8
R7779 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 433.8
R7780 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 433.8
R7781 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 433.8
R7782 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 433.8
R7783 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 433.8
R7784 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 433.8
R7785 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 433.8
R7786 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 433.8
R7787 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 433.8
R7788 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 433.8
R7789 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 433.8
R7790 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 433.8
R7791 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 433.8
R7792 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 433.8
R7793 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 433.8
R7794 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 433.8
R7795 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 339.836
R7796 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 339.834
R7797 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 339.272
R7798 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 334.772
R7799 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 221.293
R7800 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 176.733
R7801 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 176.733
R7802 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 176.733
R7803 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 176.733
R7804 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 176.733
R7805 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 176.733
R7806 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 176.733
R7807 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 176.733
R7808 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 176.733
R7809 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 176.733
R7810 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 176.733
R7811 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 176.733
R7812 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 176.733
R7813 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 176.733
R7814 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 176.733
R7815 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 176.733
R7816 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 118.45
R7817 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.V_tail_gate.n29 86.7036
R7818 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 64.5795
R7819 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 56.2338
R7820 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 56.2338
R7821 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 53.2453
R7822 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 39.4005
R7823 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 39.4005
R7824 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 39.4005
R7825 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 39.4005
R7826 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 39.4005
R7827 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 39.4005
R7828 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 39.4005
R7829 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 39.4005
R7830 bgr_0.TAIL_CUR_MIR_BIAS two_stage_opamp_dummy_magic_0.V_tail_gate.n6 18.3599
R7831 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 16.0005
R7832 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 16.0005
R7833 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 16.0005
R7834 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 16.0005
R7835 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 4.5005
R7836 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 0.563
R7837 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.n0 219.928
R7838 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t0 16.0005
R7839 two_stage_opamp_dummy_magic_0.V_p_mir.n0 two_stage_opamp_dummy_magic_0.V_p_mir.t1 16.0005
R7840 two_stage_opamp_dummy_magic_0.V_p_mir.t2 two_stage_opamp_dummy_magic_0.V_p_mir.n1 9.6005
R7841 two_stage_opamp_dummy_magic_0.V_p_mir.n1 two_stage_opamp_dummy_magic_0.V_p_mir.t3 9.6005
R7842 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 525.38
R7843 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 525.38
R7844 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 366.856
R7845 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 366.856
R7846 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 281.168
R7847 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 281.168
R7848 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 281.168
R7849 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 281.168
R7850 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 244.214
R7851 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 244.214
R7852 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 166.03
R7853 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 166.03
R7854 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 117.849
R7855 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 117.849
R7856 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 85.6894
R7857 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 85.6894
R7858 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 36.813
R7859 bgr_0.V_p_2.n0 bgr_0.V_p_2.n2 229.562
R7860 bgr_0.V_p_2.n1 bgr_0.V_p_2.n5 228.939
R7861 bgr_0.V_p_2.n0 bgr_0.V_p_2.n4 228.939
R7862 bgr_0.V_p_2.n0 bgr_0.V_p_2.n3 228.939
R7863 bgr_0.V_p_2.n6 bgr_0.V_p_2.n1 228.938
R7864 bgr_0.V_p_2.n1 bgr_0.V_p_2.t6 98.2279
R7865 bgr_0.V_p_2.n5 bgr_0.V_p_2.t8 48.0005
R7866 bgr_0.V_p_2.n5 bgr_0.V_p_2.t4 48.0005
R7867 bgr_0.V_p_2.n4 bgr_0.V_p_2.t1 48.0005
R7868 bgr_0.V_p_2.n4 bgr_0.V_p_2.t0 48.0005
R7869 bgr_0.V_p_2.n3 bgr_0.V_p_2.t7 48.0005
R7870 bgr_0.V_p_2.n3 bgr_0.V_p_2.t3 48.0005
R7871 bgr_0.V_p_2.n2 bgr_0.V_p_2.t2 48.0005
R7872 bgr_0.V_p_2.n2 bgr_0.V_p_2.t10 48.0005
R7873 bgr_0.V_p_2.t5 bgr_0.V_p_2.n6 48.0005
R7874 bgr_0.V_p_2.n6 bgr_0.V_p_2.t9 48.0005
R7875 bgr_0.V_p_2.n1 bgr_0.V_p_2.n0 1.8755
R7876 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n3 630.827
R7877 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n8 630.264
R7878 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n6 630.264
R7879 two_stage_opamp_dummy_magic_0.V_err_p.n5 two_stage_opamp_dummy_magic_0.V_err_p.n4 630.264
R7880 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n13 627.784
R7881 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n0 627.784
R7882 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n2 627.168
R7883 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n16 626.534
R7884 two_stage_opamp_dummy_magic_0.V_err_p.n15 two_stage_opamp_dummy_magic_0.V_err_p.n14 626.534
R7885 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.n18 626.534
R7886 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n1 622.034
R7887 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t13 78.8005
R7888 two_stage_opamp_dummy_magic_0.V_err_p.n16 two_stage_opamp_dummy_magic_0.V_err_p.t18 78.8005
R7889 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t10 78.8005
R7890 two_stage_opamp_dummy_magic_0.V_err_p.n14 two_stage_opamp_dummy_magic_0.V_err_p.t15 78.8005
R7891 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t17 78.8005
R7892 two_stage_opamp_dummy_magic_0.V_err_p.n13 two_stage_opamp_dummy_magic_0.V_err_p.t20 78.8005
R7893 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t16 78.8005
R7894 two_stage_opamp_dummy_magic_0.V_err_p.n1 two_stage_opamp_dummy_magic_0.V_err_p.t11 78.8005
R7895 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t1 78.8005
R7896 two_stage_opamp_dummy_magic_0.V_err_p.n8 two_stage_opamp_dummy_magic_0.V_err_p.t5 78.8005
R7897 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t6 78.8005
R7898 two_stage_opamp_dummy_magic_0.V_err_p.n6 two_stage_opamp_dummy_magic_0.V_err_p.t4 78.8005
R7899 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t3 78.8005
R7900 two_stage_opamp_dummy_magic_0.V_err_p.n4 two_stage_opamp_dummy_magic_0.V_err_p.t8 78.8005
R7901 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t9 78.8005
R7902 two_stage_opamp_dummy_magic_0.V_err_p.n3 two_stage_opamp_dummy_magic_0.V_err_p.t2 78.8005
R7903 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t7 78.8005
R7904 two_stage_opamp_dummy_magic_0.V_err_p.n2 two_stage_opamp_dummy_magic_0.V_err_p.t0 78.8005
R7905 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t21 78.8005
R7906 two_stage_opamp_dummy_magic_0.V_err_p.n0 two_stage_opamp_dummy_magic_0.V_err_p.t12 78.8005
R7907 two_stage_opamp_dummy_magic_0.V_err_p.n19 two_stage_opamp_dummy_magic_0.V_err_p.t14 78.8005
R7908 two_stage_opamp_dummy_magic_0.V_err_p.t19 two_stage_opamp_dummy_magic_0.V_err_p.n19 78.8005
R7909 two_stage_opamp_dummy_magic_0.V_err_p.n10 two_stage_opamp_dummy_magic_0.V_err_p.n9 5.0005
R7910 two_stage_opamp_dummy_magic_0.V_err_p.n12 two_stage_opamp_dummy_magic_0.V_err_p.n11 4.5005
R7911 two_stage_opamp_dummy_magic_0.V_err_p.n11 two_stage_opamp_dummy_magic_0.V_err_p.n10 1.60845
R7912 two_stage_opamp_dummy_magic_0.V_err_p.n17 two_stage_opamp_dummy_magic_0.V_err_p.n15 1.2505
R7913 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n17 1.2505
R7914 two_stage_opamp_dummy_magic_0.V_err_p.n18 two_stage_opamp_dummy_magic_0.V_err_p.n12 1.2505
R7915 two_stage_opamp_dummy_magic_0.V_err_p.n7 two_stage_opamp_dummy_magic_0.V_err_p.n5 0.563
R7916 two_stage_opamp_dummy_magic_0.V_err_p.n9 two_stage_opamp_dummy_magic_0.V_err_p.n7 0.563
R7917 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.t6 327.623
R7918 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.t4 326.365
R7919 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t10 168.701
R7920 two_stage_opamp_dummy_magic_0.V_tot.n5 two_stage_opamp_dummy_magic_0.V_tot.t9 168.701
R7921 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n1 167.05
R7922 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n7 165.8
R7923 two_stage_opamp_dummy_magic_0.V_tot.n6 two_stage_opamp_dummy_magic_0.V_tot.n5 165.8
R7924 two_stage_opamp_dummy_magic_0.V_tot.n3 two_stage_opamp_dummy_magic_0.V_tot.n2 165.8
R7925 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t13 157.989
R7926 two_stage_opamp_dummy_magic_0.V_tot.n7 two_stage_opamp_dummy_magic_0.V_tot.t7 157.989
R7927 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t8 157.989
R7928 two_stage_opamp_dummy_magic_0.V_tot.n2 two_stage_opamp_dummy_magic_0.V_tot.t12 157.989
R7929 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t5 157.989
R7930 two_stage_opamp_dummy_magic_0.V_tot.n1 two_stage_opamp_dummy_magic_0.V_tot.t11 157.989
R7931 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t3 117.591
R7932 two_stage_opamp_dummy_magic_0.V_tot.t0 two_stage_opamp_dummy_magic_0.V_tot.n11 117.591
R7933 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.t1 108.424
R7934 two_stage_opamp_dummy_magic_0.V_tot.n0 two_stage_opamp_dummy_magic_0.V_tot.t2 108.424
R7935 two_stage_opamp_dummy_magic_0.V_tot.n11 two_stage_opamp_dummy_magic_0.V_tot.n10 37.2371
R7936 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n0 37.1746
R7937 two_stage_opamp_dummy_magic_0.V_tot.n10 two_stage_opamp_dummy_magic_0.V_tot.n9 10.6255
R7938 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n8 1.8755
R7939 two_stage_opamp_dummy_magic_0.V_tot.n9 two_stage_opamp_dummy_magic_0.V_tot.n4 1.31612
R7940 two_stage_opamp_dummy_magic_0.V_tot.n8 two_stage_opamp_dummy_magic_0.V_tot.n6 1.26612
R7941 two_stage_opamp_dummy_magic_0.V_tot.n4 two_stage_opamp_dummy_magic_0.V_tot.n3 1.15363
R7942 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n9 114.719
R7943 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n4 114.719
R7944 two_stage_opamp_dummy_magic_0.VD1.n6 two_stage_opamp_dummy_magic_0.VD1.n5 114.156
R7945 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.n7 114.156
R7946 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n0 113.081
R7947 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n15 111.769
R7948 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n17 111.769
R7949 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n19 111.769
R7950 two_stage_opamp_dummy_magic_0.VD1.n2 two_stage_opamp_dummy_magic_0.VD1.n1 111.769
R7951 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n3 109.656
R7952 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n12 107.269
R7953 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t12 16.0005
R7954 two_stage_opamp_dummy_magic_0.VD1.n3 two_stage_opamp_dummy_magic_0.VD1.t17 16.0005
R7955 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t7 16.0005
R7956 two_stage_opamp_dummy_magic_0.VD1.n15 two_stage_opamp_dummy_magic_0.VD1.t2 16.0005
R7957 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t5 16.0005
R7958 two_stage_opamp_dummy_magic_0.VD1.n17 two_stage_opamp_dummy_magic_0.VD1.t0 16.0005
R7959 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t10 16.0005
R7960 two_stage_opamp_dummy_magic_0.VD1.n19 two_stage_opamp_dummy_magic_0.VD1.t1 16.0005
R7961 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t21 16.0005
R7962 two_stage_opamp_dummy_magic_0.VD1.n1 two_stage_opamp_dummy_magic_0.VD1.t3 16.0005
R7963 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t8 16.0005
R7964 two_stage_opamp_dummy_magic_0.VD1.n0 two_stage_opamp_dummy_magic_0.VD1.t4 16.0005
R7965 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t6 16.0005
R7966 two_stage_opamp_dummy_magic_0.VD1.n12 two_stage_opamp_dummy_magic_0.VD1.t9 16.0005
R7967 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.t11 16.0005
R7968 two_stage_opamp_dummy_magic_0.VD1.n9 two_stage_opamp_dummy_magic_0.VD1.t16 16.0005
R7969 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t13 16.0005
R7970 two_stage_opamp_dummy_magic_0.VD1.n5 two_stage_opamp_dummy_magic_0.VD1.t15 16.0005
R7971 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t14 16.0005
R7972 two_stage_opamp_dummy_magic_0.VD1.n4 two_stage_opamp_dummy_magic_0.VD1.t19 16.0005
R7973 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t20 16.0005
R7974 two_stage_opamp_dummy_magic_0.VD1.n7 two_stage_opamp_dummy_magic_0.VD1.t18 16.0005
R7975 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n13 4.5005
R7976 two_stage_opamp_dummy_magic_0.VD1.n11 two_stage_opamp_dummy_magic_0.VD1.n10 4.5005
R7977 two_stage_opamp_dummy_magic_0.VD1.n16 two_stage_opamp_dummy_magic_0.VD1.n14 3.563
R7978 two_stage_opamp_dummy_magic_0.VD1.n18 two_stage_opamp_dummy_magic_0.VD1.n16 1.313
R7979 two_stage_opamp_dummy_magic_0.VD1.n14 two_stage_opamp_dummy_magic_0.VD1.n2 1.2505
R7980 two_stage_opamp_dummy_magic_0.VD1 two_stage_opamp_dummy_magic_0.VD1.n18 1.2505
R7981 two_stage_opamp_dummy_magic_0.VD1.n10 two_stage_opamp_dummy_magic_0.VD1.n8 0.563
R7982 two_stage_opamp_dummy_magic_0.VD1.n8 two_stage_opamp_dummy_magic_0.VD1.n6 0.563
R7983 two_stage_opamp_dummy_magic_0.VD1.n13 two_stage_opamp_dummy_magic_0.VD1.n11 0.21925
R7984 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 344.837
R7985 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 344.274
R7986 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 292.5
R7987 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 206.052
R7988 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 205.488
R7989 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 205.488
R7990 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 205.488
R7991 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 205.488
R7992 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 122.474
R7993 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 80.6567
R7994 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 71.2813
R7995 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 52.3363
R7996 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 39.4005
R7997 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 39.4005
R7998 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 39.4005
R7999 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 39.4005
R8000 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 39.4005
R8001 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 39.4005
R8002 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 19.7005
R8003 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 19.7005
R8004 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 19.7005
R8005 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 19.7005
R8006 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 19.7005
R8007 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 19.7005
R8008 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 19.7005
R8009 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 19.7005
R8010 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 19.7005
R8011 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 19.7005
R8012 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 6.1255
R8013 bgr_0.V_CMFB_S1 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 1.15675
R8014 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 0.563
R8015 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 0.563
R8016 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 0.563
R8017 bgr_0.Vin+.n3 bgr_0.Vin+.n2 526.183
R8018 bgr_0.Vin+.n1 bgr_0.Vin+.n0 514.134
R8019 bgr_0.Vin+.n0 bgr_0.Vin+.t6 303.259
R8020 bgr_0.Vin+.n7 bgr_0.Vin+.n3 215.732
R8021 bgr_0.Vin+.n0 bgr_0.Vin+.t8 174.726
R8022 bgr_0.Vin+.n1 bgr_0.Vin+.t10 174.726
R8023 bgr_0.Vin+.n2 bgr_0.Vin+.t7 174.726
R8024 bgr_0.Vin+.n6 bgr_0.Vin+.n4 170.56
R8025 bgr_0.Vin+.n6 bgr_0.Vin+.n5 168.435
R8026 bgr_0.Vin+.n8 bgr_0.Vin+.t5 158.796
R8027 bgr_0.Vin+.t0 bgr_0.Vin+.n8 147.981
R8028 bgr_0.Vin+.n2 bgr_0.Vin+.n1 128.534
R8029 bgr_0.Vin+.n3 bgr_0.Vin+.t9 96.4005
R8030 bgr_0.Vin+.n7 bgr_0.Vin+.n6 13.5005
R8031 bgr_0.Vin+.n5 bgr_0.Vin+.t1 13.1338
R8032 bgr_0.Vin+.n5 bgr_0.Vin+.t4 13.1338
R8033 bgr_0.Vin+.n4 bgr_0.Vin+.t3 13.1338
R8034 bgr_0.Vin+.n4 bgr_0.Vin+.t2 13.1338
R8035 bgr_0.Vin+.n8 bgr_0.Vin+.n7 1.438
R8036 bgr_0.V_p_1.n6 bgr_0.V_p_1.n1 229.562
R8037 bgr_0.V_p_1.n1 bgr_0.V_p_1.n5 228.939
R8038 bgr_0.V_p_1.n1 bgr_0.V_p_1.n4 228.939
R8039 bgr_0.V_p_1.n0 bgr_0.V_p_1.n3 228.939
R8040 bgr_0.V_p_1.n0 bgr_0.V_p_1.n2 228.939
R8041 bgr_0.V_p_1.n0 bgr_0.V_p_1.t10 98.2279
R8042 bgr_0.V_p_1.n5 bgr_0.V_p_1.t5 48.0005
R8043 bgr_0.V_p_1.n5 bgr_0.V_p_1.t2 48.0005
R8044 bgr_0.V_p_1.n4 bgr_0.V_p_1.t0 48.0005
R8045 bgr_0.V_p_1.n4 bgr_0.V_p_1.t9 48.0005
R8046 bgr_0.V_p_1.n3 bgr_0.V_p_1.t6 48.0005
R8047 bgr_0.V_p_1.n3 bgr_0.V_p_1.t3 48.0005
R8048 bgr_0.V_p_1.n2 bgr_0.V_p_1.t1 48.0005
R8049 bgr_0.V_p_1.n2 bgr_0.V_p_1.t8 48.0005
R8050 bgr_0.V_p_1.t4 bgr_0.V_p_1.n6 48.0005
R8051 bgr_0.V_p_1.n6 bgr_0.V_p_1.t7 48.0005
R8052 bgr_0.V_p_1.n1 bgr_0.V_p_1.n0 1.8755
R8053 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.t13 355.293
R8054 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.t14 346.8
R8055 bgr_0.1st_Vout_2.n21 bgr_0.1st_Vout_2.n20 339.522
R8056 bgr_0.1st_Vout_2.n7 bgr_0.1st_Vout_2.n6 339.522
R8057 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.n14 335.022
R8058 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.t9 275.909
R8059 bgr_0.1st_Vout_2.n11 bgr_0.1st_Vout_2.n10 227.909
R8060 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n12 222.034
R8061 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t26 184.097
R8062 bgr_0.1st_Vout_2.n17 bgr_0.1st_Vout_2.t36 184.097
R8063 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t19 184.097
R8064 bgr_0.1st_Vout_2.n8 bgr_0.1st_Vout_2.t32 184.097
R8065 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n17 166.05
R8066 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.n8 166.05
R8067 bgr_0.1st_Vout_2.n19 bgr_0.1st_Vout_2.n4 57.7228
R8068 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t0 48.0005
R8069 bgr_0.1st_Vout_2.n12 bgr_0.1st_Vout_2.t8 48.0005
R8070 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t10 48.0005
R8071 bgr_0.1st_Vout_2.n10 bgr_0.1st_Vout_2.t7 48.0005
R8072 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.t1 39.4005
R8073 bgr_0.1st_Vout_2.n14 bgr_0.1st_Vout_2.t4 39.4005
R8074 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t3 39.4005
R8075 bgr_0.1st_Vout_2.n6 bgr_0.1st_Vout_2.t5 39.4005
R8076 bgr_0.1st_Vout_2.t6 bgr_0.1st_Vout_2.n21 39.4005
R8077 bgr_0.1st_Vout_2.n21 bgr_0.1st_Vout_2.t2 39.4005
R8078 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t17 4.8295
R8079 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t16 4.8295
R8080 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t27 4.8295
R8081 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t23 4.8295
R8082 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t35 4.8295
R8083 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t34 4.8295
R8084 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t28 4.8295
R8085 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t21 4.5005
R8086 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t15 4.5005
R8087 bgr_0.1st_Vout_2.n1 bgr_0.1st_Vout_2.t12 4.5005
R8088 bgr_0.1st_Vout_2.n5 bgr_0.1st_Vout_2.t30 4.5005
R8089 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t22 4.5005
R8090 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.t18 4.5005
R8091 bgr_0.1st_Vout_2.n3 bgr_0.1st_Vout_2.t11 4.5005
R8092 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t31 4.5005
R8093 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t29 4.5005
R8094 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t33 4.5005
R8095 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.t24 4.5005
R8096 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t20 4.5005
R8097 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.t25 4.5005
R8098 bgr_0.1st_Vout_2.n13 bgr_0.1st_Vout_2.n11 4.5005
R8099 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.n15 4.5005
R8100 bgr_0.1st_Vout_2.n9 bgr_0.1st_Vout_2.n7 1.3755
R8101 bgr_0.1st_Vout_2.n18 bgr_0.1st_Vout_2.n16 1.3755
R8102 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n19 1.188
R8103 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n5 0.9405
R8104 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n0 0.8935
R8105 bgr_0.1st_Vout_2.n15 bgr_0.1st_Vout_2.n13 0.78175
R8106 bgr_0.1st_Vout_2.n4 bgr_0.1st_Vout_2.n2 0.6585
R8107 bgr_0.1st_Vout_2.n2 bgr_0.1st_Vout_2.n3 0.6585
R8108 bgr_0.1st_Vout_2.n0 bgr_0.1st_Vout_2.n1 0.6585
R8109 bgr_0.1st_Vout_2.n16 bgr_0.1st_Vout_2.n9 0.6255
R8110 bgr_0.1st_Vout_2.n20 bgr_0.1st_Vout_2.n18 0.6255
R8111 bgr_0.cap_res2 bgr_0.cap_res2.t20 188.315
R8112 bgr_0.cap_res2 bgr_0.cap_res2.t9 0.259
R8113 bgr_0.cap_res2.t13 bgr_0.cap_res2.t8 0.1603
R8114 bgr_0.cap_res2.t2 bgr_0.cap_res2.t6 0.1603
R8115 bgr_0.cap_res2.t5 bgr_0.cap_res2.t1 0.1603
R8116 bgr_0.cap_res2.t19 bgr_0.cap_res2.t0 0.1603
R8117 bgr_0.cap_res2.t14 bgr_0.cap_res2.t10 0.1603
R8118 bgr_0.cap_res2.t4 bgr_0.cap_res2.t7 0.1603
R8119 bgr_0.cap_res2.t18 bgr_0.cap_res2.t16 0.1603
R8120 bgr_0.cap_res2.t12 bgr_0.cap_res2.t15 0.1603
R8121 bgr_0.cap_res2.n1 bgr_0.cap_res2.t17 0.159278
R8122 bgr_0.cap_res2.n2 bgr_0.cap_res2.t11 0.159278
R8123 bgr_0.cap_res2.n3 bgr_0.cap_res2.t3 0.159278
R8124 bgr_0.cap_res2.n3 bgr_0.cap_res2.t13 0.1368
R8125 bgr_0.cap_res2.n3 bgr_0.cap_res2.t2 0.1368
R8126 bgr_0.cap_res2.n2 bgr_0.cap_res2.t5 0.1368
R8127 bgr_0.cap_res2.n2 bgr_0.cap_res2.t19 0.1368
R8128 bgr_0.cap_res2.n1 bgr_0.cap_res2.t14 0.1368
R8129 bgr_0.cap_res2.n1 bgr_0.cap_res2.t4 0.1368
R8130 bgr_0.cap_res2.n0 bgr_0.cap_res2.t18 0.1368
R8131 bgr_0.cap_res2.n0 bgr_0.cap_res2.t12 0.1368
R8132 bgr_0.cap_res2.t17 bgr_0.cap_res2.n0 0.00152174
R8133 bgr_0.cap_res2.t11 bgr_0.cap_res2.n1 0.00152174
R8134 bgr_0.cap_res2.t3 bgr_0.cap_res2.n2 0.00152174
R8135 bgr_0.cap_res2.t9 bgr_0.cap_res2.n3 0.00152174
R8136 two_stage_opamp_dummy_magic_0.V_source.n9 two_stage_opamp_dummy_magic_0.V_source.t39 206.47
R8137 two_stage_opamp_dummy_magic_0.V_source.n28 two_stage_opamp_dummy_magic_0.V_source.n26 118.168
R8138 two_stage_opamp_dummy_magic_0.V_source.n21 two_stage_opamp_dummy_magic_0.V_source.n19 117.831
R8139 two_stage_opamp_dummy_magic_0.V_source.n34 two_stage_opamp_dummy_magic_0.V_source.n33 117.269
R8140 two_stage_opamp_dummy_magic_0.V_source.n32 two_stage_opamp_dummy_magic_0.V_source.n31 117.269
R8141 two_stage_opamp_dummy_magic_0.V_source.n30 two_stage_opamp_dummy_magic_0.V_source.n29 117.269
R8142 two_stage_opamp_dummy_magic_0.V_source.n28 two_stage_opamp_dummy_magic_0.V_source.n27 117.269
R8143 two_stage_opamp_dummy_magic_0.V_source.n25 two_stage_opamp_dummy_magic_0.V_source.n24 117.269
R8144 two_stage_opamp_dummy_magic_0.V_source.n23 two_stage_opamp_dummy_magic_0.V_source.n22 117.269
R8145 two_stage_opamp_dummy_magic_0.V_source.n21 two_stage_opamp_dummy_magic_0.V_source.n20 117.269
R8146 two_stage_opamp_dummy_magic_0.V_source.n36 two_stage_opamp_dummy_magic_0.V_source.n18 113.136
R8147 two_stage_opamp_dummy_magic_0.V_source.n2 two_stage_opamp_dummy_magic_0.V_source.n0 99.7407
R8148 two_stage_opamp_dummy_magic_0.V_source.n5 two_stage_opamp_dummy_magic_0.V_source.n3 99.647
R8149 two_stage_opamp_dummy_magic_0.V_source.n16 two_stage_opamp_dummy_magic_0.V_source.n15 99.0845
R8150 two_stage_opamp_dummy_magic_0.V_source.n14 two_stage_opamp_dummy_magic_0.V_source.n13 99.0845
R8151 two_stage_opamp_dummy_magic_0.V_source.n12 two_stage_opamp_dummy_magic_0.V_source.n11 99.0845
R8152 two_stage_opamp_dummy_magic_0.V_source.n7 two_stage_opamp_dummy_magic_0.V_source.n6 99.0845
R8153 two_stage_opamp_dummy_magic_0.V_source.n5 two_stage_opamp_dummy_magic_0.V_source.n4 99.0845
R8154 two_stage_opamp_dummy_magic_0.V_source.n2 two_stage_opamp_dummy_magic_0.V_source.n1 99.0845
R8155 two_stage_opamp_dummy_magic_0.V_source.n38 two_stage_opamp_dummy_magic_0.V_source.n37 94.5857
R8156 two_stage_opamp_dummy_magic_0.V_source.n9 two_stage_opamp_dummy_magic_0.V_source.n8 94.5845
R8157 two_stage_opamp_dummy_magic_0.V_source.n33 two_stage_opamp_dummy_magic_0.V_source.t4 16.0005
R8158 two_stage_opamp_dummy_magic_0.V_source.n33 two_stage_opamp_dummy_magic_0.V_source.t0 16.0005
R8159 two_stage_opamp_dummy_magic_0.V_source.n31 two_stage_opamp_dummy_magic_0.V_source.t15 16.0005
R8160 two_stage_opamp_dummy_magic_0.V_source.n31 two_stage_opamp_dummy_magic_0.V_source.t13 16.0005
R8161 two_stage_opamp_dummy_magic_0.V_source.n29 two_stage_opamp_dummy_magic_0.V_source.t2 16.0005
R8162 two_stage_opamp_dummy_magic_0.V_source.n29 two_stage_opamp_dummy_magic_0.V_source.t12 16.0005
R8163 two_stage_opamp_dummy_magic_0.V_source.n27 two_stage_opamp_dummy_magic_0.V_source.t19 16.0005
R8164 two_stage_opamp_dummy_magic_0.V_source.n27 two_stage_opamp_dummy_magic_0.V_source.t20 16.0005
R8165 two_stage_opamp_dummy_magic_0.V_source.n26 two_stage_opamp_dummy_magic_0.V_source.t3 16.0005
R8166 two_stage_opamp_dummy_magic_0.V_source.n26 two_stage_opamp_dummy_magic_0.V_source.t11 16.0005
R8167 two_stage_opamp_dummy_magic_0.V_source.n24 two_stage_opamp_dummy_magic_0.V_source.t1 16.0005
R8168 two_stage_opamp_dummy_magic_0.V_source.n24 two_stage_opamp_dummy_magic_0.V_source.t14 16.0005
R8169 two_stage_opamp_dummy_magic_0.V_source.n22 two_stage_opamp_dummy_magic_0.V_source.t8 16.0005
R8170 two_stage_opamp_dummy_magic_0.V_source.n22 two_stage_opamp_dummy_magic_0.V_source.t7 16.0005
R8171 two_stage_opamp_dummy_magic_0.V_source.n20 two_stage_opamp_dummy_magic_0.V_source.t17 16.0005
R8172 two_stage_opamp_dummy_magic_0.V_source.n20 two_stage_opamp_dummy_magic_0.V_source.t40 16.0005
R8173 two_stage_opamp_dummy_magic_0.V_source.n19 two_stage_opamp_dummy_magic_0.V_source.t9 16.0005
R8174 two_stage_opamp_dummy_magic_0.V_source.n19 two_stage_opamp_dummy_magic_0.V_source.t6 16.0005
R8175 two_stage_opamp_dummy_magic_0.V_source.n18 two_stage_opamp_dummy_magic_0.V_source.t18 16.0005
R8176 two_stage_opamp_dummy_magic_0.V_source.n18 two_stage_opamp_dummy_magic_0.V_source.t10 16.0005
R8177 two_stage_opamp_dummy_magic_0.V_source.n15 two_stage_opamp_dummy_magic_0.V_source.t35 9.6005
R8178 two_stage_opamp_dummy_magic_0.V_source.n15 two_stage_opamp_dummy_magic_0.V_source.t25 9.6005
R8179 two_stage_opamp_dummy_magic_0.V_source.n13 two_stage_opamp_dummy_magic_0.V_source.t33 9.6005
R8180 two_stage_opamp_dummy_magic_0.V_source.n13 two_stage_opamp_dummy_magic_0.V_source.t23 9.6005
R8181 two_stage_opamp_dummy_magic_0.V_source.n11 two_stage_opamp_dummy_magic_0.V_source.t29 9.6005
R8182 two_stage_opamp_dummy_magic_0.V_source.n11 two_stage_opamp_dummy_magic_0.V_source.t21 9.6005
R8183 two_stage_opamp_dummy_magic_0.V_source.n8 two_stage_opamp_dummy_magic_0.V_source.t32 9.6005
R8184 two_stage_opamp_dummy_magic_0.V_source.n8 two_stage_opamp_dummy_magic_0.V_source.t22 9.6005
R8185 two_stage_opamp_dummy_magic_0.V_source.n6 two_stage_opamp_dummy_magic_0.V_source.t28 9.6005
R8186 two_stage_opamp_dummy_magic_0.V_source.n6 two_stage_opamp_dummy_magic_0.V_source.t36 9.6005
R8187 two_stage_opamp_dummy_magic_0.V_source.n4 two_stage_opamp_dummy_magic_0.V_source.t26 9.6005
R8188 two_stage_opamp_dummy_magic_0.V_source.n4 two_stage_opamp_dummy_magic_0.V_source.t34 9.6005
R8189 two_stage_opamp_dummy_magic_0.V_source.n3 two_stage_opamp_dummy_magic_0.V_source.t24 9.6005
R8190 two_stage_opamp_dummy_magic_0.V_source.n3 two_stage_opamp_dummy_magic_0.V_source.t30 9.6005
R8191 two_stage_opamp_dummy_magic_0.V_source.n1 two_stage_opamp_dummy_magic_0.V_source.t37 9.6005
R8192 two_stage_opamp_dummy_magic_0.V_source.n1 two_stage_opamp_dummy_magic_0.V_source.t31 9.6005
R8193 two_stage_opamp_dummy_magic_0.V_source.n0 two_stage_opamp_dummy_magic_0.V_source.t16 9.6005
R8194 two_stage_opamp_dummy_magic_0.V_source.n0 two_stage_opamp_dummy_magic_0.V_source.t5 9.6005
R8195 two_stage_opamp_dummy_magic_0.V_source.t38 two_stage_opamp_dummy_magic_0.V_source.n38 9.6005
R8196 two_stage_opamp_dummy_magic_0.V_source.n38 two_stage_opamp_dummy_magic_0.V_source.t27 9.6005
R8197 two_stage_opamp_dummy_magic_0.V_source.n10 two_stage_opamp_dummy_magic_0.V_source.n9 4.5005
R8198 two_stage_opamp_dummy_magic_0.V_source.n36 two_stage_opamp_dummy_magic_0.V_source.n35 4.5005
R8199 two_stage_opamp_dummy_magic_0.V_source.n37 two_stage_opamp_dummy_magic_0.V_source.n17 4.5005
R8200 two_stage_opamp_dummy_magic_0.V_source.n35 two_stage_opamp_dummy_magic_0.V_source.n34 3.65675
R8201 two_stage_opamp_dummy_magic_0.V_source.n37 two_stage_opamp_dummy_magic_0.V_source.n36 1.28175
R8202 two_stage_opamp_dummy_magic_0.V_source.n7 two_stage_opamp_dummy_magic_0.V_source.n5 0.563
R8203 two_stage_opamp_dummy_magic_0.V_source.n10 two_stage_opamp_dummy_magic_0.V_source.n7 0.563
R8204 two_stage_opamp_dummy_magic_0.V_source.n12 two_stage_opamp_dummy_magic_0.V_source.n10 0.563
R8205 two_stage_opamp_dummy_magic_0.V_source.n14 two_stage_opamp_dummy_magic_0.V_source.n12 0.563
R8206 two_stage_opamp_dummy_magic_0.V_source.n16 two_stage_opamp_dummy_magic_0.V_source.n14 0.563
R8207 two_stage_opamp_dummy_magic_0.V_source.n17 two_stage_opamp_dummy_magic_0.V_source.n16 0.563
R8208 two_stage_opamp_dummy_magic_0.V_source.n17 two_stage_opamp_dummy_magic_0.V_source.n2 0.563
R8209 two_stage_opamp_dummy_magic_0.V_source.n30 two_stage_opamp_dummy_magic_0.V_source.n28 0.563
R8210 two_stage_opamp_dummy_magic_0.V_source.n32 two_stage_opamp_dummy_magic_0.V_source.n30 0.563
R8211 two_stage_opamp_dummy_magic_0.V_source.n34 two_stage_opamp_dummy_magic_0.V_source.n32 0.563
R8212 two_stage_opamp_dummy_magic_0.V_source.n23 two_stage_opamp_dummy_magic_0.V_source.n21 0.563
R8213 two_stage_opamp_dummy_magic_0.V_source.n25 two_stage_opamp_dummy_magic_0.V_source.n23 0.563
R8214 two_stage_opamp_dummy_magic_0.V_source.n35 two_stage_opamp_dummy_magic_0.V_source.n25 0.53175
R8215 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 144.827
R8216 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 134.577
R8217 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 120.66
R8218 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 97.4009
R8219 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 96.8384
R8220 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 96.8384
R8221 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 96.8384
R8222 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 96.8384
R8223 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 88.938
R8224 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 24.0005
R8225 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 24.0005
R8226 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 24.0005
R8227 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 24.0005
R8228 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 8.0005
R8229 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 8.0005
R8230 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 8.0005
R8231 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 8.0005
R8232 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 8.0005
R8233 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 8.0005
R8234 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 8.0005
R8235 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 8.0005
R8236 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 8.0005
R8237 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 8.0005
R8238 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 5.813
R8239 bgr_0.V_CMFB_S4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 1.46925
R8240 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 0.563
R8241 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 0.563
R8242 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 0.563
R8243 VIN-.n4 VIN-.t8 485.021
R8244 VIN-.n1 VIN-.t6 484.159
R8245 VIN-.n5 VIN-.t7 483.358
R8246 VIN-.n8 VIN-.t10 431.536
R8247 VIN-.n2 VIN-.t9 431.536
R8248 VIN-.n6 VIN-.t1 431.257
R8249 VIN-.n0 VIN-.t0 431.257
R8250 VIN-.n6 VIN-.t2 289.908
R8251 VIN-.n0 VIN-.t5 289.908
R8252 VIN-.n8 VIN-.t4 279.183
R8253 VIN-.n2 VIN-.t3 279.183
R8254 VIN-.n7 VIN-.n6 233.374
R8255 VIN-.n1 VIN-.n0 233.374
R8256 VIN-.n9 VIN-.n8 188.989
R8257 VIN-.n3 VIN-.n2 188.989
R8258 VIN-.n4 VIN-.n3 2.463
R8259 VIN- VIN-.n9 1.78175
R8260 VIN-.n5 VIN-.n4 1.563
R8261 VIN-.n3 VIN-.n1 1.2755
R8262 VIN-.n9 VIN-.n7 1.2755
R8263 VIN-.n7 VIN-.n5 0.8005
R8264 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.t12 670.048
R8265 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n0 631.982
R8266 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n3 627.128
R8267 two_stage_opamp_dummy_magic_0.err_amp_out.n2 two_stage_opamp_dummy_magic_0.err_amp_out.n1 627.128
R8268 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n7 226.534
R8269 two_stage_opamp_dummy_magic_0.err_amp_out.n6 two_stage_opamp_dummy_magic_0.err_amp_out.n5 226.534
R8270 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n4 222.034
R8271 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t0 78.8005
R8272 two_stage_opamp_dummy_magic_0.err_amp_out.n3 two_stage_opamp_dummy_magic_0.err_amp_out.t2 78.8005
R8273 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t1 78.8005
R8274 two_stage_opamp_dummy_magic_0.err_amp_out.n1 two_stage_opamp_dummy_magic_0.err_amp_out.t3 78.8005
R8275 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t5 78.8005
R8276 two_stage_opamp_dummy_magic_0.err_amp_out.n0 two_stage_opamp_dummy_magic_0.err_amp_out.t4 78.8005
R8277 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t7 48.0005
R8278 two_stage_opamp_dummy_magic_0.err_amp_out.n7 two_stage_opamp_dummy_magic_0.err_amp_out.t9 48.0005
R8279 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.t6 48.0005
R8280 two_stage_opamp_dummy_magic_0.err_amp_out.n4 two_stage_opamp_dummy_magic_0.err_amp_out.t11 48.0005
R8281 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t8 48.0005
R8282 two_stage_opamp_dummy_magic_0.err_amp_out.n5 two_stage_opamp_dummy_magic_0.err_amp_out.t10 48.0005
R8283 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n9 8.938
R8284 two_stage_opamp_dummy_magic_0.err_amp_out.n9 two_stage_opamp_dummy_magic_0.err_amp_out.n8 5.7505
R8285 two_stage_opamp_dummy_magic_0.err_amp_out two_stage_opamp_dummy_magic_0.err_amp_out.n2 1.313
R8286 two_stage_opamp_dummy_magic_0.err_amp_out.n8 two_stage_opamp_dummy_magic_0.err_amp_out.n6 1.2505
R8287 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n1 4020
R8288 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n1 4020
R8289 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n7 4020
R8290 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.n7 4020
R8291 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.t28 660.109
R8292 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.t25 660.109
R8293 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.n11 422.401
R8294 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.n0 422.401
R8295 two_stage_opamp_dummy_magic_0.VD3.t29 two_stage_opamp_dummy_magic_0.VD3.n8 239.915
R8296 two_stage_opamp_dummy_magic_0.VD3.n10 two_stage_opamp_dummy_magic_0.VD3.t26 239.915
R8297 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n5 230.4
R8298 two_stage_opamp_dummy_magic_0.VD3.n6 two_stage_opamp_dummy_magic_0.VD3.n3 230.4
R8299 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n3 198.4
R8300 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.n0 198.4
R8301 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.n28 160.428
R8302 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n13 160.427
R8303 two_stage_opamp_dummy_magic_0.VD3.n30 two_stage_opamp_dummy_magic_0.VD3.n29 159.803
R8304 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.n26 159.803
R8305 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n24 159.803
R8306 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n22 159.802
R8307 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n20 159.802
R8308 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n18 159.802
R8309 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n16 159.802
R8310 two_stage_opamp_dummy_magic_0.VD3.n15 two_stage_opamp_dummy_magic_0.VD3.n14 159.802
R8311 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.n32 155.304
R8312 two_stage_opamp_dummy_magic_0.VD3.n4 two_stage_opamp_dummy_magic_0.VD3.t30 155.125
R8313 two_stage_opamp_dummy_magic_0.VD3.n2 two_stage_opamp_dummy_magic_0.VD3.t27 155.125
R8314 two_stage_opamp_dummy_magic_0.VD3.t0 two_stage_opamp_dummy_magic_0.VD3.t29 98.2764
R8315 two_stage_opamp_dummy_magic_0.VD3.t6 two_stage_opamp_dummy_magic_0.VD3.t0 98.2764
R8316 two_stage_opamp_dummy_magic_0.VD3.t14 two_stage_opamp_dummy_magic_0.VD3.t6 98.2764
R8317 two_stage_opamp_dummy_magic_0.VD3.t10 two_stage_opamp_dummy_magic_0.VD3.t14 98.2764
R8318 two_stage_opamp_dummy_magic_0.VD3.t16 two_stage_opamp_dummy_magic_0.VD3.t10 98.2764
R8319 two_stage_opamp_dummy_magic_0.VD3.t2 two_stage_opamp_dummy_magic_0.VD3.t18 98.2764
R8320 two_stage_opamp_dummy_magic_0.VD3.t8 two_stage_opamp_dummy_magic_0.VD3.t2 98.2764
R8321 two_stage_opamp_dummy_magic_0.VD3.t4 two_stage_opamp_dummy_magic_0.VD3.t8 98.2764
R8322 two_stage_opamp_dummy_magic_0.VD3.t12 two_stage_opamp_dummy_magic_0.VD3.t4 98.2764
R8323 two_stage_opamp_dummy_magic_0.VD3.t26 two_stage_opamp_dummy_magic_0.VD3.t12 98.2764
R8324 two_stage_opamp_dummy_magic_0.VD3.n11 two_stage_opamp_dummy_magic_0.VD3.n10 92.5005
R8325 two_stage_opamp_dummy_magic_0.VD3.n7 two_stage_opamp_dummy_magic_0.VD3.n6 92.5005
R8326 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.n7 92.5005
R8327 two_stage_opamp_dummy_magic_0.VD3.n8 two_stage_opamp_dummy_magic_0.VD3.n0 92.5005
R8328 two_stage_opamp_dummy_magic_0.VD3.n12 two_stage_opamp_dummy_magic_0.VD3.n1 92.5005
R8329 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.n1 92.5005
R8330 two_stage_opamp_dummy_magic_0.VD3.n9 two_stage_opamp_dummy_magic_0.VD3.t16 49.1384
R8331 two_stage_opamp_dummy_magic_0.VD3.t18 two_stage_opamp_dummy_magic_0.VD3.n9 49.1384
R8332 two_stage_opamp_dummy_magic_0.VD3.n5 two_stage_opamp_dummy_magic_0.VD3.n4 21.3338
R8333 two_stage_opamp_dummy_magic_0.VD3.n3 two_stage_opamp_dummy_magic_0.VD3.n2 21.3338
R8334 two_stage_opamp_dummy_magic_0.VD3.n25 two_stage_opamp_dummy_magic_0.VD3.n23 14.438
R8335 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.t3 11.2576
R8336 two_stage_opamp_dummy_magic_0.VD3.n29 two_stage_opamp_dummy_magic_0.VD3.t9 11.2576
R8337 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.t5 11.2576
R8338 two_stage_opamp_dummy_magic_0.VD3.n28 two_stage_opamp_dummy_magic_0.VD3.t13 11.2576
R8339 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.t15 11.2576
R8340 two_stage_opamp_dummy_magic_0.VD3.n26 two_stage_opamp_dummy_magic_0.VD3.t11 11.2576
R8341 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t1 11.2576
R8342 two_stage_opamp_dummy_magic_0.VD3.n24 two_stage_opamp_dummy_magic_0.VD3.t7 11.2576
R8343 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.t21 11.2576
R8344 two_stage_opamp_dummy_magic_0.VD3.n22 two_stage_opamp_dummy_magic_0.VD3.t36 11.2576
R8345 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t34 11.2576
R8346 two_stage_opamp_dummy_magic_0.VD3.n20 two_stage_opamp_dummy_magic_0.VD3.t32 11.2576
R8347 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t24 11.2576
R8348 two_stage_opamp_dummy_magic_0.VD3.n18 two_stage_opamp_dummy_magic_0.VD3.t31 11.2576
R8349 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.t22 11.2576
R8350 two_stage_opamp_dummy_magic_0.VD3.n16 two_stage_opamp_dummy_magic_0.VD3.t37 11.2576
R8351 two_stage_opamp_dummy_magic_0.VD3.n14 two_stage_opamp_dummy_magic_0.VD3.t23 11.2576
R8352 two_stage_opamp_dummy_magic_0.VD3.n14 two_stage_opamp_dummy_magic_0.VD3.t20 11.2576
R8353 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.t35 11.2576
R8354 two_stage_opamp_dummy_magic_0.VD3.n13 two_stage_opamp_dummy_magic_0.VD3.t33 11.2576
R8355 two_stage_opamp_dummy_magic_0.VD3.n33 two_stage_opamp_dummy_magic_0.VD3.t17 11.2576
R8356 two_stage_opamp_dummy_magic_0.VD3.t19 two_stage_opamp_dummy_magic_0.VD3.n33 11.2576
R8357 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.n12 9.5505
R8358 two_stage_opamp_dummy_magic_0.VD3.n32 two_stage_opamp_dummy_magic_0.VD3.n31 4.5005
R8359 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n30 0.6255
R8360 two_stage_opamp_dummy_magic_0.VD3.n17 two_stage_opamp_dummy_magic_0.VD3.n15 0.6255
R8361 two_stage_opamp_dummy_magic_0.VD3.n19 two_stage_opamp_dummy_magic_0.VD3.n17 0.6255
R8362 two_stage_opamp_dummy_magic_0.VD3.n21 two_stage_opamp_dummy_magic_0.VD3.n19 0.6255
R8363 two_stage_opamp_dummy_magic_0.VD3.n23 two_stage_opamp_dummy_magic_0.VD3.n21 0.6255
R8364 two_stage_opamp_dummy_magic_0.VD3.n27 two_stage_opamp_dummy_magic_0.VD3.n25 0.6255
R8365 two_stage_opamp_dummy_magic_0.VD3.n31 two_stage_opamp_dummy_magic_0.VD3.n27 0.6255
R8366 a_14240_2076.t0 a_14240_2076.t1 169.905
R8367 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.t20 619.201
R8368 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t12 611.739
R8369 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t25 611.739
R8370 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t11 611.739
R8371 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t21 611.739
R8372 two_stage_opamp_dummy_magic_0.Vb3.n18 two_stage_opamp_dummy_magic_0.Vb3.t18 421.75
R8373 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.t22 421.75
R8374 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.t24 421.75
R8375 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.t27 421.75
R8376 two_stage_opamp_dummy_magic_0.Vb3.n14 two_stage_opamp_dummy_magic_0.Vb3.t23 421.75
R8377 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.t19 421.75
R8378 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.t14 421.75
R8379 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.t9 421.75
R8380 two_stage_opamp_dummy_magic_0.Vb3.n9 two_stage_opamp_dummy_magic_0.Vb3.t17 421.75
R8381 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.t15 421.75
R8382 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.t26 421.75
R8383 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.t28 421.75
R8384 two_stage_opamp_dummy_magic_0.Vb3.n5 two_stage_opamp_dummy_magic_0.Vb3.t16 421.75
R8385 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.t10 421.75
R8386 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.t13 421.75
R8387 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.t8 421.75
R8388 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n22 176.155
R8389 two_stage_opamp_dummy_magic_0.Vb3.n23 two_stage_opamp_dummy_magic_0.Vb3.n13 175.79
R8390 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n25 172.667
R8391 two_stage_opamp_dummy_magic_0.Vb3.n19 two_stage_opamp_dummy_magic_0.Vb3.n18 167.094
R8392 two_stage_opamp_dummy_magic_0.Vb3.n20 two_stage_opamp_dummy_magic_0.Vb3.n19 167.094
R8393 two_stage_opamp_dummy_magic_0.Vb3.n21 two_stage_opamp_dummy_magic_0.Vb3.n20 167.094
R8394 two_stage_opamp_dummy_magic_0.Vb3.n15 two_stage_opamp_dummy_magic_0.Vb3.n14 167.094
R8395 two_stage_opamp_dummy_magic_0.Vb3.n16 two_stage_opamp_dummy_magic_0.Vb3.n15 167.094
R8396 two_stage_opamp_dummy_magic_0.Vb3.n17 two_stage_opamp_dummy_magic_0.Vb3.n16 167.094
R8397 two_stage_opamp_dummy_magic_0.Vb3.n10 two_stage_opamp_dummy_magic_0.Vb3.n9 167.094
R8398 two_stage_opamp_dummy_magic_0.Vb3.n11 two_stage_opamp_dummy_magic_0.Vb3.n10 167.094
R8399 two_stage_opamp_dummy_magic_0.Vb3.n12 two_stage_opamp_dummy_magic_0.Vb3.n11 167.094
R8400 two_stage_opamp_dummy_magic_0.Vb3.n6 two_stage_opamp_dummy_magic_0.Vb3.n5 167.094
R8401 two_stage_opamp_dummy_magic_0.Vb3.n7 two_stage_opamp_dummy_magic_0.Vb3.n6 167.094
R8402 two_stage_opamp_dummy_magic_0.Vb3.n8 two_stage_opamp_dummy_magic_0.Vb3.n7 167.094
R8403 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n1 139.639
R8404 two_stage_opamp_dummy_magic_0.Vb3.n3 two_stage_opamp_dummy_magic_0.Vb3.n2 139.638
R8405 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n0 134.577
R8406 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n26 106.891
R8407 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n21 47.1294
R8408 two_stage_opamp_dummy_magic_0.Vb3.n22 two_stage_opamp_dummy_magic_0.Vb3.n17 47.1294
R8409 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n12 47.1294
R8410 two_stage_opamp_dummy_magic_0.Vb3.n13 two_stage_opamp_dummy_magic_0.Vb3.n8 47.1294
R8411 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t1 24.0005
R8412 two_stage_opamp_dummy_magic_0.Vb3.n0 two_stage_opamp_dummy_magic_0.Vb3.t4 24.0005
R8413 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t2 24.0005
R8414 two_stage_opamp_dummy_magic_0.Vb3.n2 two_stage_opamp_dummy_magic_0.Vb3.t7 24.0005
R8415 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t5 24.0005
R8416 two_stage_opamp_dummy_magic_0.Vb3.n1 two_stage_opamp_dummy_magic_0.Vb3.t3 24.0005
R8417 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t6 10.9449
R8418 two_stage_opamp_dummy_magic_0.Vb3.n25 two_stage_opamp_dummy_magic_0.Vb3.t0 10.9449
R8419 two_stage_opamp_dummy_magic_0.Vb3.n24 two_stage_opamp_dummy_magic_0.Vb3.n23 9.5005
R8420 two_stage_opamp_dummy_magic_0.Vb3.n26 two_stage_opamp_dummy_magic_0.Vb3.n24 8.79738
R8421 two_stage_opamp_dummy_magic_0.Vb3.n4 two_stage_opamp_dummy_magic_0.Vb3.n3 4.5005
R8422 bgr_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_0.Vb3.n4 0.96925
R8423 a_11220_17410.t0 a_11220_17410.t1 258.591
R8424 a_14640_5068.t0 a_14640_5068.t1 169.905
R8425 VIN+.n9 VIN+.t5 485.127
R8426 VIN+.n4 VIN+.t3 485.127
R8427 VIN+.n3 VIN+.t4 485.127
R8428 VIN+.n7 VIN+.t9 318.656
R8429 VIN+.n7 VIN+.t2 318.656
R8430 VIN+.n5 VIN+.t7 318.656
R8431 VIN+.n5 VIN+.t1 318.656
R8432 VIN+.n1 VIN+.t8 318.656
R8433 VIN+.n1 VIN+.t6 318.656
R8434 VIN+.n0 VIN+.t10 318.656
R8435 VIN+.n0 VIN+.t0 318.656
R8436 VIN+.n2 VIN+.n0 167.05
R8437 VIN+.n8 VIN+.n7 165.8
R8438 VIN+.n6 VIN+.n5 165.8
R8439 VIN+.n2 VIN+.n1 165.8
R8440 VIN+.n6 VIN+.n4 2.34425
R8441 VIN+.n4 VIN+.n3 1.3005
R8442 VIN+.n8 VIN+.n6 1.2505
R8443 VIN+.n3 VIN+.n2 1.15675
R8444 VIN+.n9 VIN+.n8 1.15675
R8445 VIN+ VIN+.n9 0.963
R8446 a_13730_17020.t0 a_13730_17020.t1 258.591
R8447 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.n2 526.183
R8448 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.n0 514.134
R8449 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t3 303.259
R8450 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n4 287.264
R8451 bgr_0.V_CUR_REF_REG.n5 bgr_0.V_CUR_REF_REG.n3 283.961
R8452 bgr_0.V_CUR_REF_REG.t0 bgr_0.V_CUR_REF_REG.n5 245.284
R8453 bgr_0.V_CUR_REF_REG.n0 bgr_0.V_CUR_REF_REG.t7 174.726
R8454 bgr_0.V_CUR_REF_REG.n1 bgr_0.V_CUR_REF_REG.t5 174.726
R8455 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.t6 174.726
R8456 bgr_0.V_CUR_REF_REG.n2 bgr_0.V_CUR_REF_REG.n1 128.534
R8457 bgr_0.V_CUR_REF_REG.n3 bgr_0.V_CUR_REF_REG.t4 96.4005
R8458 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t1 39.4005
R8459 bgr_0.V_CUR_REF_REG.n4 bgr_0.V_CUR_REF_REG.t2 39.4005
R8460 a_12828_17530.t0 a_12828_17530.t1 376.99
R8461 bgr_0.START_UP.n4 bgr_0.START_UP.t6 238.322
R8462 bgr_0.START_UP.n4 bgr_0.START_UP.t7 238.322
R8463 bgr_0.START_UP.n3 bgr_0.START_UP.n1 175.56
R8464 bgr_0.START_UP.n3 bgr_0.START_UP.n2 168.936
R8465 bgr_0.START_UP.n5 bgr_0.START_UP.n4 166.925
R8466 bgr_0.START_UP.n0 bgr_0.START_UP.t5 130.001
R8467 bgr_0.START_UP.n0 bgr_0.START_UP.t4 81.7074
R8468 bgr_0.START_UP bgr_0.START_UP.n0 38.2614
R8469 bgr_0.START_UP bgr_0.START_UP.n5 14.7817
R8470 bgr_0.START_UP.n1 bgr_0.START_UP.t0 13.1338
R8471 bgr_0.START_UP.n1 bgr_0.START_UP.t1 13.1338
R8472 bgr_0.START_UP.n2 bgr_0.START_UP.t2 13.1338
R8473 bgr_0.START_UP.n2 bgr_0.START_UP.t3 13.1338
R8474 bgr_0.START_UP.n5 bgr_0.START_UP.n3 4.21925
R8475 a_11220_17290.t0 a_11220_17290.t1 376.99
R8476 a_12828_17650.t0 a_12828_17650.t1 258.591
R8477 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2655
R8478 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2595
R8479 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 2280
R8480 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 2250
R8481 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t5 672.159
R8482 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t2 672.159
R8483 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 276.8
R8484 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 240
R8485 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 206.4
R8486 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 204.8
R8487 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 180.904
R8488 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 170.3
R8489 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 160.517
R8490 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 160.517
R8491 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 110.425
R8492 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 110.05
R8493 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t3 95.7988
R8494 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n3 92.5005
R8495 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n4 92.5005
R8496 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 92.5005
R8497 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n5 92.5005
R8498 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 89.6005
R8499 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 89.6005
R8500 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 76.8005
R8501 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t4 75.9449
R8502 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n15 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t8 75.9449
R8503 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t0 47.8997
R8504 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n10 47.8997
R8505 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n2 38.4005
R8506 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n6 24.5338
R8507 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n14 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n13 24.5338
R8508 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n8 16.8187
R8509 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n12 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n11 16.8187
R8510 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t9 12.313
R8511 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n18 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t10 12.313
R8512 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t1 10.9449
R8513 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_0.Vb2_Vb3.t7 10.9449
R8514 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 6.21925
R8515 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n17 two_stage_opamp_dummy_magic_0.Vb2_Vb3.n16 4.5005
R8516 a_5230_5068.t0 a_5230_5068.t1 294.339
R8517 a_5750_2076.t0 a_5750_2076.t1 169.905
R8518 a_13790_17550.t0 a_13790_17550.t1 258.591
R8519 a_5350_5068.t0 a_5350_5068.t1 169.905
C0 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.VD4 0.10263f
C1 bgr_0.PFET_GATE_10uA bgr_0.cap_res2 0.018633f
C2 bgr_0.Vbe2 bgr_0.NFET_GATE_10uA 0.021455f
C3 bgr_0.NFET_GATE_10uA VDDA 1.04957f
C4 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.cap_res_Y 0.790473f
C5 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.err_amp_out 0.253351f
C6 two_stage_opamp_dummy_magic_0.VD4 VDDA 4.37879f
C7 bgr_0.V_TOP two_stage_opamp_dummy_magic_0.V_err_amp_ref 1.13839f
C8 bgr_0.START_UP bgr_0.PFET_GATE_10uA 0.166283f
C9 two_stage_opamp_dummy_magic_0.Vb2_Vb3 VDDA 0.874875f
C10 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.1st_Vout_1 0.477103f
C11 two_stage_opamp_dummy_magic_0.cap_res_Y VDDA 0.921549f
C12 two_stage_opamp_dummy_magic_0.X VDDA 5.37188f
C13 bgr_0.Vbe2 bgr_0.V_TOP 0.285619f
C14 bgr_0.V_TOP VDDA 16.1464f
C15 bgr_0.1st_Vout_1 VDDA 2.06087f
C16 bgr_0.START_UP_NFET1 bgr_0.START_UP 0.145663f
C17 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.cap_res_Y 0.036092f
C18 bgr_0.V_TOP bgr_0.NFET_GATE_10uA 0.080353f
C19 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.cap_res2 0.551434f
C20 bgr_0.1st_Vout_1 bgr_0.NFET_GATE_10uA 1.02268f
C21 bgr_0.START_UP two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.09763f
C22 bgr_0.cap_res2 VDDA 0.586627f
C23 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.VD1 1.05329f
C24 two_stage_opamp_dummy_magic_0.VD1 VIN- 0.881216f
C25 bgr_0.V_TOP bgr_0.1st_Vout_1 0.925484f
C26 m2_8540_19780# VDDA 0.010446f
C27 bgr_0.START_UP bgr_0.Vbe2 0.193132f
C28 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.V_err_gate 1.3735f
C29 bgr_0.START_UP VDDA 1.37391f
C30 two_stage_opamp_dummy_magic_0.V_err_amp_ref two_stage_opamp_dummy_magic_0.err_amp_out 0.528215f
C31 VIN- VIN+ 0.562828f
C32 two_stage_opamp_dummy_magic_0.VD1 VIN+ 0.058217f
C33 bgr_0.START_UP bgr_0.NFET_GATE_10uA 0.518732f
C34 two_stage_opamp_dummy_magic_0.cap_res_Y bgr_0.cap_res2 0.048779f
C35 two_stage_opamp_dummy_magic_0.V_err_gate VDDA 4.87848f
C36 bgr_0.PFET_GATE_10uA m2_7180_19780# 0.012f
C37 two_stage_opamp_dummy_magic_0.err_amp_out VDDA 1.20093f
C38 bgr_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_amp_ref 2.46518f
C39 bgr_0.NFET_GATE_10uA two_stage_opamp_dummy_magic_0.V_err_gate 0.136183f
C40 bgr_0.1st_Vout_1 bgr_0.cap_res2 0.822981f
C41 bgr_0.V_TOP m2_8540_19780# 0.012f
C42 two_stage_opamp_dummy_magic_0.VD4 two_stage_opamp_dummy_magic_0.V_err_gate 0.013177f
C43 bgr_0.Vbe2 bgr_0.PFET_GATE_10uA 0.242909f
C44 bgr_0.START_UP bgr_0.V_TOP 0.815644f
C45 two_stage_opamp_dummy_magic_0.Vb2_Vb3 two_stage_opamp_dummy_magic_0.V_err_gate 0.065464f
C46 bgr_0.1st_Vout_1 m2_8540_19780# 0.075543f
C47 bgr_0.PFET_GATE_10uA VDDA 10.4831f
C48 bgr_0.START_UP bgr_0.1st_Vout_1 0.030647f
C49 two_stage_opamp_dummy_magic_0.V_err_gate two_stage_opamp_dummy_magic_0.X 0.166227f
C50 bgr_0.PFET_GATE_10uA bgr_0.NFET_GATE_10uA 0.050552f
C51 two_stage_opamp_dummy_magic_0.X two_stage_opamp_dummy_magic_0.err_amp_out 0.426362f
C52 bgr_0.START_UP_NFET1 VDDA 0.15057f
C53 bgr_0.PFET_GATE_10uA bgr_0.V_TOP 2.47366f
C54 bgr_0.START_UP_NFET1 bgr_0.NFET_GATE_10uA 0.318695f
C55 bgr_0.PFET_GATE_10uA bgr_0.1st_Vout_1 0.035393f
C56 m2_7180_19780# VDDA 0.010446f
C57 bgr_0.Vbe2 two_stage_opamp_dummy_magic_0.V_err_amp_ref 0.014154f
C58 two_stage_opamp_dummy_magic_0.V_err_amp_ref VDDA 4.36f
C59 two_stage_opamp_dummy_magic_0.V_err_amp_ref bgr_0.NFET_GATE_10uA 0.559544f
C60 bgr_0.Vbe2 VDDA 0.016701f
C61 VOUT+ GNDA 0.038801f
C62 VOUT- GNDA 0.038805f
C63 VIN+ GNDA 2.062214f
C64 VIN- GNDA 2.130657f
C65 VDDA GNDA 0.151768p
C66 two_stage_opamp_dummy_magic_0.VD1 GNDA 2.43523f
C67 two_stage_opamp_dummy_magic_0.err_amp_out GNDA 2.703803f
C68 two_stage_opamp_dummy_magic_0.cap_res_Y GNDA 33.253426f
C69 two_stage_opamp_dummy_magic_0.X GNDA 5.567724f
C70 bgr_0.cap_res2 GNDA 7.933997f
C71 bgr_0.1st_Vout_1 GNDA 4.989391f
C72 two_stage_opamp_dummy_magic_0.V_err_amp_ref GNDA 15.176401f
C73 bgr_0.V_TOP GNDA 6.831957f
C74 bgr_0.PFET_GATE_10uA GNDA 5.0864f
C75 bgr_0.Vbe2 GNDA 17.0659f
C76 bgr_0.START_UP GNDA 7.190113f
C77 bgr_0.START_UP_NFET1 GNDA 5.28334f
C78 two_stage_opamp_dummy_magic_0.V_err_gate GNDA 14.579249f
C79 bgr_0.NFET_GATE_10uA GNDA 7.22507f
C80 two_stage_opamp_dummy_magic_0.VD4 GNDA 6.478767f
C81 two_stage_opamp_dummy_magic_0.Vb2_Vb3 GNDA 3.6041f
C82 bgr_0.START_UP.t4 GNDA 1.6623f
C83 bgr_0.START_UP.t5 GNDA 0.043697f
C84 bgr_0.START_UP.n0 GNDA 1.12862f
C85 bgr_0.START_UP.t0 GNDA 0.041701f
C86 bgr_0.START_UP.t1 GNDA 0.041701f
C87 bgr_0.START_UP.n1 GNDA 0.151283f
C88 bgr_0.START_UP.t2 GNDA 0.041701f
C89 bgr_0.START_UP.t3 GNDA 0.041701f
C90 bgr_0.START_UP.n2 GNDA 0.139173f
C91 bgr_0.START_UP.n3 GNDA 0.720787f
C92 bgr_0.START_UP.t7 GNDA 0.01567f
C93 bgr_0.START_UP.t6 GNDA 0.01567f
C94 bgr_0.START_UP.n4 GNDA 0.044238f
C95 bgr_0.START_UP.n5 GNDA 0.445182f
C96 bgr_0.V_CUR_REF_REG.t3 GNDA 0.014208f
C97 bgr_0.V_CUR_REF_REG.n0 GNDA 0.030473f
C98 bgr_0.V_CUR_REF_REG.n1 GNDA 0.023714f
C99 bgr_0.V_CUR_REF_REG.n2 GNDA 0.024034f
C100 bgr_0.V_CUR_REF_REG.n3 GNDA 0.231183f
C101 bgr_0.V_CUR_REF_REG.n4 GNDA 0.01997f
C102 bgr_0.V_CUR_REF_REG.n5 GNDA 1.47498f
C103 bgr_0.V_CUR_REF_REG.t0 GNDA 0.42777f
C104 VIN+.t0 GNDA 0.042021f
C105 VIN+.t10 GNDA 0.042021f
C106 VIN+.n0 GNDA 0.086842f
C107 VIN+.t6 GNDA 0.042021f
C108 VIN+.t8 GNDA 0.042021f
C109 VIN+.n1 GNDA 0.085639f
C110 VIN+.n2 GNDA 0.361638f
C111 VIN+.t4 GNDA 0.059118f
C112 VIN+.n3 GNDA 0.216459f
C113 VIN+.t3 GNDA 0.059118f
C114 VIN+.n4 GNDA 0.263959f
C115 VIN+.t1 GNDA 0.042021f
C116 VIN+.t7 GNDA 0.042021f
C117 VIN+.n5 GNDA 0.085639f
C118 VIN+.n6 GNDA 0.249653f
C119 VIN+.t2 GNDA 0.042021f
C120 VIN+.t9 GNDA 0.042021f
C121 VIN+.n7 GNDA 0.085639f
C122 VIN+.n8 GNDA 0.202005f
C123 VIN+.t5 GNDA 0.059118f
C124 VIN+.n9 GNDA 0.202625f
C125 bgr_0.VB3_CUR_BIAS GNDA 4.82031f
C126 two_stage_opamp_dummy_magic_0.Vb3.t1 GNDA 0.032596f
C127 two_stage_opamp_dummy_magic_0.Vb3.t4 GNDA 0.032596f
C128 two_stage_opamp_dummy_magic_0.Vb3.n0 GNDA 0.098454f
C129 two_stage_opamp_dummy_magic_0.Vb3.t5 GNDA 0.032596f
C130 two_stage_opamp_dummy_magic_0.Vb3.t3 GNDA 0.032596f
C131 two_stage_opamp_dummy_magic_0.Vb3.n1 GNDA 0.104995f
C132 two_stage_opamp_dummy_magic_0.Vb3.t2 GNDA 0.032596f
C133 two_stage_opamp_dummy_magic_0.Vb3.t7 GNDA 0.032596f
C134 two_stage_opamp_dummy_magic_0.Vb3.n2 GNDA 0.104995f
C135 two_stage_opamp_dummy_magic_0.Vb3.n3 GNDA 0.578833f
C136 two_stage_opamp_dummy_magic_0.Vb3.n4 GNDA 0.216097f
C137 two_stage_opamp_dummy_magic_0.Vb3.t20 GNDA 0.185645f
C138 two_stage_opamp_dummy_magic_0.Vb3.t8 GNDA 0.16135f
C139 two_stage_opamp_dummy_magic_0.Vb3.t13 GNDA 0.16135f
C140 two_stage_opamp_dummy_magic_0.Vb3.t10 GNDA 0.16135f
C141 two_stage_opamp_dummy_magic_0.Vb3.t16 GNDA 0.16135f
C142 two_stage_opamp_dummy_magic_0.Vb3.t21 GNDA 0.186197f
C143 two_stage_opamp_dummy_magic_0.Vb3.n5 GNDA 0.151172f
C144 two_stage_opamp_dummy_magic_0.Vb3.n6 GNDA 0.092898f
C145 two_stage_opamp_dummy_magic_0.Vb3.n7 GNDA 0.092898f
C146 two_stage_opamp_dummy_magic_0.Vb3.n8 GNDA 0.086987f
C147 two_stage_opamp_dummy_magic_0.Vb3.t28 GNDA 0.16135f
C148 two_stage_opamp_dummy_magic_0.Vb3.t26 GNDA 0.16135f
C149 two_stage_opamp_dummy_magic_0.Vb3.t15 GNDA 0.16135f
C150 two_stage_opamp_dummy_magic_0.Vb3.t17 GNDA 0.16135f
C151 two_stage_opamp_dummy_magic_0.Vb3.t11 GNDA 0.186197f
C152 two_stage_opamp_dummy_magic_0.Vb3.n9 GNDA 0.151172f
C153 two_stage_opamp_dummy_magic_0.Vb3.n10 GNDA 0.092898f
C154 two_stage_opamp_dummy_magic_0.Vb3.n11 GNDA 0.092898f
C155 two_stage_opamp_dummy_magic_0.Vb3.n12 GNDA 0.086987f
C156 two_stage_opamp_dummy_magic_0.Vb3.n13 GNDA 0.090228f
C157 two_stage_opamp_dummy_magic_0.Vb3.t9 GNDA 0.16135f
C158 two_stage_opamp_dummy_magic_0.Vb3.t14 GNDA 0.16135f
C159 two_stage_opamp_dummy_magic_0.Vb3.t19 GNDA 0.16135f
C160 two_stage_opamp_dummy_magic_0.Vb3.t23 GNDA 0.16135f
C161 two_stage_opamp_dummy_magic_0.Vb3.t25 GNDA 0.186197f
C162 two_stage_opamp_dummy_magic_0.Vb3.n14 GNDA 0.151172f
C163 two_stage_opamp_dummy_magic_0.Vb3.n15 GNDA 0.092898f
C164 two_stage_opamp_dummy_magic_0.Vb3.n16 GNDA 0.092898f
C165 two_stage_opamp_dummy_magic_0.Vb3.n17 GNDA 0.086987f
C166 two_stage_opamp_dummy_magic_0.Vb3.t27 GNDA 0.16135f
C167 two_stage_opamp_dummy_magic_0.Vb3.t24 GNDA 0.16135f
C168 two_stage_opamp_dummy_magic_0.Vb3.t22 GNDA 0.16135f
C169 two_stage_opamp_dummy_magic_0.Vb3.t18 GNDA 0.16135f
C170 two_stage_opamp_dummy_magic_0.Vb3.t12 GNDA 0.186197f
C171 two_stage_opamp_dummy_magic_0.Vb3.n18 GNDA 0.151172f
C172 two_stage_opamp_dummy_magic_0.Vb3.n19 GNDA 0.092898f
C173 two_stage_opamp_dummy_magic_0.Vb3.n20 GNDA 0.092898f
C174 two_stage_opamp_dummy_magic_0.Vb3.n21 GNDA 0.086987f
C175 two_stage_opamp_dummy_magic_0.Vb3.n22 GNDA 0.093614f
C176 two_stage_opamp_dummy_magic_0.Vb3.n23 GNDA 2.5592f
C177 two_stage_opamp_dummy_magic_0.Vb3.n24 GNDA 0.713797f
C178 two_stage_opamp_dummy_magic_0.Vb3.t6 GNDA 0.117345f
C179 two_stage_opamp_dummy_magic_0.Vb3.t0 GNDA 0.117345f
C180 two_stage_opamp_dummy_magic_0.Vb3.n25 GNDA 0.419988f
C181 two_stage_opamp_dummy_magic_0.Vb3.n26 GNDA 5.16137f
C182 two_stage_opamp_dummy_magic_0.VD3.t17 GNDA 0.026025f
C183 two_stage_opamp_dummy_magic_0.VD3.n0 GNDA 0.073371f
C184 two_stage_opamp_dummy_magic_0.VD3.n1 GNDA 0.100747f
C185 two_stage_opamp_dummy_magic_0.VD3.t27 GNDA 0.128386f
C186 two_stage_opamp_dummy_magic_0.VD3.t25 GNDA 0.045318f
C187 two_stage_opamp_dummy_magic_0.VD3.n2 GNDA 0.083755f
C188 two_stage_opamp_dummy_magic_0.VD3.n3 GNDA 0.053992f
C189 two_stage_opamp_dummy_magic_0.VD3.t30 GNDA 0.128386f
C190 two_stage_opamp_dummy_magic_0.VD3.t28 GNDA 0.045318f
C191 two_stage_opamp_dummy_magic_0.VD3.n4 GNDA 0.083755f
C192 two_stage_opamp_dummy_magic_0.VD3.n5 GNDA 0.053992f
C193 two_stage_opamp_dummy_magic_0.VD3.n6 GNDA 0.053537f
C194 two_stage_opamp_dummy_magic_0.VD3.n7 GNDA 0.100747f
C195 two_stage_opamp_dummy_magic_0.VD3.n8 GNDA 0.300245f
C196 two_stage_opamp_dummy_magic_0.VD3.t29 GNDA 0.448159f
C197 two_stage_opamp_dummy_magic_0.VD3.t0 GNDA 0.25876f
C198 two_stage_opamp_dummy_magic_0.VD3.t6 GNDA 0.25876f
C199 two_stage_opamp_dummy_magic_0.VD3.t14 GNDA 0.25876f
C200 two_stage_opamp_dummy_magic_0.VD3.t10 GNDA 0.25876f
C201 two_stage_opamp_dummy_magic_0.VD3.t16 GNDA 0.19407f
C202 two_stage_opamp_dummy_magic_0.VD3.n9 GNDA 0.12938f
C203 two_stage_opamp_dummy_magic_0.VD3.t18 GNDA 0.19407f
C204 two_stage_opamp_dummy_magic_0.VD3.t2 GNDA 0.25876f
C205 two_stage_opamp_dummy_magic_0.VD3.t8 GNDA 0.25876f
C206 two_stage_opamp_dummy_magic_0.VD3.t4 GNDA 0.25876f
C207 two_stage_opamp_dummy_magic_0.VD3.t12 GNDA 0.25876f
C208 two_stage_opamp_dummy_magic_0.VD3.t26 GNDA 0.448159f
C209 two_stage_opamp_dummy_magic_0.VD3.n10 GNDA 0.300245f
C210 two_stage_opamp_dummy_magic_0.VD3.n11 GNDA 0.073371f
C211 two_stage_opamp_dummy_magic_0.VD3.n12 GNDA 0.108171f
C212 two_stage_opamp_dummy_magic_0.VD3.t35 GNDA 0.026025f
C213 two_stage_opamp_dummy_magic_0.VD3.t33 GNDA 0.026025f
C214 two_stage_opamp_dummy_magic_0.VD3.n13 GNDA 0.090509f
C215 two_stage_opamp_dummy_magic_0.VD3.t23 GNDA 0.026025f
C216 two_stage_opamp_dummy_magic_0.VD3.t20 GNDA 0.026025f
C217 two_stage_opamp_dummy_magic_0.VD3.n14 GNDA 0.090188f
C218 two_stage_opamp_dummy_magic_0.VD3.n15 GNDA 0.170266f
C219 two_stage_opamp_dummy_magic_0.VD3.t22 GNDA 0.026025f
C220 two_stage_opamp_dummy_magic_0.VD3.t37 GNDA 0.026025f
C221 two_stage_opamp_dummy_magic_0.VD3.n16 GNDA 0.090188f
C222 two_stage_opamp_dummy_magic_0.VD3.n17 GNDA 0.088268f
C223 two_stage_opamp_dummy_magic_0.VD3.t24 GNDA 0.026025f
C224 two_stage_opamp_dummy_magic_0.VD3.t31 GNDA 0.026025f
C225 two_stage_opamp_dummy_magic_0.VD3.n18 GNDA 0.090188f
C226 two_stage_opamp_dummy_magic_0.VD3.n19 GNDA 0.088268f
C227 two_stage_opamp_dummy_magic_0.VD3.t34 GNDA 0.026025f
C228 two_stage_opamp_dummy_magic_0.VD3.t32 GNDA 0.026025f
C229 two_stage_opamp_dummy_magic_0.VD3.n20 GNDA 0.090188f
C230 two_stage_opamp_dummy_magic_0.VD3.n21 GNDA 0.088268f
C231 two_stage_opamp_dummy_magic_0.VD3.t21 GNDA 0.026025f
C232 two_stage_opamp_dummy_magic_0.VD3.t36 GNDA 0.026025f
C233 two_stage_opamp_dummy_magic_0.VD3.n22 GNDA 0.090188f
C234 two_stage_opamp_dummy_magic_0.VD3.n23 GNDA 0.167835f
C235 two_stage_opamp_dummy_magic_0.VD3.t1 GNDA 0.026025f
C236 two_stage_opamp_dummy_magic_0.VD3.t7 GNDA 0.026025f
C237 two_stage_opamp_dummy_magic_0.VD3.n24 GNDA 0.090188f
C238 two_stage_opamp_dummy_magic_0.VD3.n25 GNDA 0.164848f
C239 two_stage_opamp_dummy_magic_0.VD3.t15 GNDA 0.026025f
C240 two_stage_opamp_dummy_magic_0.VD3.t11 GNDA 0.026025f
C241 two_stage_opamp_dummy_magic_0.VD3.n26 GNDA 0.090188f
C242 two_stage_opamp_dummy_magic_0.VD3.n27 GNDA 0.088268f
C243 two_stage_opamp_dummy_magic_0.VD3.t5 GNDA 0.026025f
C244 two_stage_opamp_dummy_magic_0.VD3.t13 GNDA 0.026025f
C245 two_stage_opamp_dummy_magic_0.VD3.n28 GNDA 0.090509f
C246 two_stage_opamp_dummy_magic_0.VD3.t3 GNDA 0.026025f
C247 two_stage_opamp_dummy_magic_0.VD3.t9 GNDA 0.026025f
C248 two_stage_opamp_dummy_magic_0.VD3.n29 GNDA 0.090188f
C249 two_stage_opamp_dummy_magic_0.VD3.n30 GNDA 0.170266f
C250 two_stage_opamp_dummy_magic_0.VD3.n31 GNDA 0.023794f
C251 two_stage_opamp_dummy_magic_0.VD3.n32 GNDA 0.069277f
C252 two_stage_opamp_dummy_magic_0.VD3.n33 GNDA 0.08832f
C253 two_stage_opamp_dummy_magic_0.VD3.t19 GNDA 0.026025f
C254 two_stage_opamp_dummy_magic_0.err_amp_out.n0 GNDA 0.018848f
C255 two_stage_opamp_dummy_magic_0.err_amp_out.n1 GNDA 0.018642f
C256 two_stage_opamp_dummy_magic_0.err_amp_out.n2 GNDA 0.371454f
C257 two_stage_opamp_dummy_magic_0.err_amp_out.n3 GNDA 0.018642f
C258 two_stage_opamp_dummy_magic_0.err_amp_out.n4 GNDA 0.020813f
C259 two_stage_opamp_dummy_magic_0.err_amp_out.t12 GNDA 0.074665f
C260 two_stage_opamp_dummy_magic_0.err_amp_out.n5 GNDA 0.022234f
C261 two_stage_opamp_dummy_magic_0.err_amp_out.n6 GNDA 1.11353f
C262 two_stage_opamp_dummy_magic_0.err_amp_out.n7 GNDA 0.022234f
C263 two_stage_opamp_dummy_magic_0.err_amp_out.n8 GNDA 0.195309f
C264 two_stage_opamp_dummy_magic_0.err_amp_out.n9 GNDA 0.190271f
C265 VIN-.t6 GNDA 0.050911f
C266 VIN-.t5 GNDA 0.03359f
C267 VIN-.t0 GNDA 0.04147f
C268 VIN-.n0 GNDA 0.05959f
C269 VIN-.n1 GNDA 0.281971f
C270 VIN-.t3 GNDA 0.033038f
C271 VIN-.t9 GNDA 0.041485f
C272 VIN-.n2 GNDA 0.065237f
C273 VIN-.n3 GNDA 0.201948f
C274 VIN-.t8 GNDA 0.050345f
C275 VIN-.n4 GNDA 0.237498f
C276 VIN-.t7 GNDA 0.050694f
C277 VIN-.n5 GNDA 0.181582f
C278 VIN-.t2 GNDA 0.03359f
C279 VIN-.t1 GNDA 0.04147f
C280 VIN-.n6 GNDA 0.05959f
C281 VIN-.n7 GNDA 0.150425f
C282 VIN-.t4 GNDA 0.033038f
C283 VIN-.t10 GNDA 0.041485f
C284 VIN-.n8 GNDA 0.065237f
C285 VIN-.n9 GNDA 0.178598f
C286 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t0 GNDA 0.472922f
C287 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t7 GNDA 0.113952f
C288 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t13 GNDA 0.113952f
C289 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n0 GNDA 0.471236f
C290 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t6 GNDA 0.113952f
C291 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t12 GNDA 0.113952f
C292 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n1 GNDA 0.469428f
C293 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n2 GNDA 0.650863f
C294 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t10 GNDA 0.113952f
C295 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t5 GNDA 0.113952f
C296 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n3 GNDA 0.469428f
C297 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n4 GNDA 0.33963f
C298 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t9 GNDA 0.113952f
C299 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t4 GNDA 0.113952f
C300 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n5 GNDA 0.469428f
C301 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n6 GNDA 0.33963f
C302 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t8 GNDA 0.113952f
C303 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t11 GNDA 0.113952f
C304 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n7 GNDA 0.469428f
C305 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n8 GNDA 0.488135f
C306 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n9 GNDA 5.6232f
C307 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t14 GNDA 0.037984f
C308 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t1 GNDA 0.037984f
C309 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n10 GNDA 0.138061f
C310 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t3 GNDA 0.037984f
C311 two_stage_opamp_dummy_magic_0.V_CMFB_S4.t2 GNDA 0.037984f
C312 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n11 GNDA 0.114728f
C313 two_stage_opamp_dummy_magic_0.V_CMFB_S4.n12 GNDA 0.717216f
C314 bgr_0.V_CMFB_S4 GNDA 4.37522f
C315 two_stage_opamp_dummy_magic_0.V_source.t27 GNDA 0.024498f
C316 two_stage_opamp_dummy_magic_0.V_source.t16 GNDA 0.024498f
C317 two_stage_opamp_dummy_magic_0.V_source.t5 GNDA 0.024498f
C318 two_stage_opamp_dummy_magic_0.V_source.n0 GNDA 0.097805f
C319 two_stage_opamp_dummy_magic_0.V_source.t37 GNDA 0.024498f
C320 two_stage_opamp_dummy_magic_0.V_source.t31 GNDA 0.024498f
C321 two_stage_opamp_dummy_magic_0.V_source.n1 GNDA 0.097268f
C322 two_stage_opamp_dummy_magic_0.V_source.n2 GNDA 0.169458f
C323 two_stage_opamp_dummy_magic_0.V_source.t24 GNDA 0.024498f
C324 two_stage_opamp_dummy_magic_0.V_source.t30 GNDA 0.024498f
C325 two_stage_opamp_dummy_magic_0.V_source.n3 GNDA 0.09772f
C326 two_stage_opamp_dummy_magic_0.V_source.t26 GNDA 0.024498f
C327 two_stage_opamp_dummy_magic_0.V_source.t34 GNDA 0.024498f
C328 two_stage_opamp_dummy_magic_0.V_source.n4 GNDA 0.097268f
C329 two_stage_opamp_dummy_magic_0.V_source.n5 GNDA 0.166602f
C330 two_stage_opamp_dummy_magic_0.V_source.t28 GNDA 0.024498f
C331 two_stage_opamp_dummy_magic_0.V_source.t36 GNDA 0.024498f
C332 two_stage_opamp_dummy_magic_0.V_source.n6 GNDA 0.097268f
C333 two_stage_opamp_dummy_magic_0.V_source.n7 GNDA 0.086957f
C334 two_stage_opamp_dummy_magic_0.V_source.t39 GNDA 0.102648f
C335 two_stage_opamp_dummy_magic_0.V_source.t32 GNDA 0.024498f
C336 two_stage_opamp_dummy_magic_0.V_source.t22 GNDA 0.024498f
C337 two_stage_opamp_dummy_magic_0.V_source.n8 GNDA 0.09453f
C338 two_stage_opamp_dummy_magic_0.V_source.n9 GNDA 0.675932f
C339 two_stage_opamp_dummy_magic_0.V_source.n10 GNDA 0.029398f
C340 two_stage_opamp_dummy_magic_0.V_source.t29 GNDA 0.024498f
C341 two_stage_opamp_dummy_magic_0.V_source.t21 GNDA 0.024498f
C342 two_stage_opamp_dummy_magic_0.V_source.n11 GNDA 0.097268f
C343 two_stage_opamp_dummy_magic_0.V_source.n12 GNDA 0.086957f
C344 two_stage_opamp_dummy_magic_0.V_source.t33 GNDA 0.024498f
C345 two_stage_opamp_dummy_magic_0.V_source.t23 GNDA 0.024498f
C346 two_stage_opamp_dummy_magic_0.V_source.n13 GNDA 0.097268f
C347 two_stage_opamp_dummy_magic_0.V_source.n14 GNDA 0.086957f
C348 two_stage_opamp_dummy_magic_0.V_source.t35 GNDA 0.024498f
C349 two_stage_opamp_dummy_magic_0.V_source.t25 GNDA 0.024498f
C350 two_stage_opamp_dummy_magic_0.V_source.n15 GNDA 0.097268f
C351 two_stage_opamp_dummy_magic_0.V_source.n16 GNDA 0.086957f
C352 two_stage_opamp_dummy_magic_0.V_source.n17 GNDA 0.029398f
C353 two_stage_opamp_dummy_magic_0.V_source.t18 GNDA 0.014699f
C354 two_stage_opamp_dummy_magic_0.V_source.t10 GNDA 0.014699f
C355 two_stage_opamp_dummy_magic_0.V_source.n18 GNDA 0.049939f
C356 two_stage_opamp_dummy_magic_0.V_source.t9 GNDA 0.014699f
C357 two_stage_opamp_dummy_magic_0.V_source.t6 GNDA 0.014699f
C358 two_stage_opamp_dummy_magic_0.V_source.n19 GNDA 0.052807f
C359 two_stage_opamp_dummy_magic_0.V_source.t17 GNDA 0.014699f
C360 two_stage_opamp_dummy_magic_0.V_source.t40 GNDA 0.014699f
C361 two_stage_opamp_dummy_magic_0.V_source.n20 GNDA 0.0524f
C362 two_stage_opamp_dummy_magic_0.V_source.n21 GNDA 0.177206f
C363 two_stage_opamp_dummy_magic_0.V_source.t8 GNDA 0.014699f
C364 two_stage_opamp_dummy_magic_0.V_source.t7 GNDA 0.014699f
C365 two_stage_opamp_dummy_magic_0.V_source.n22 GNDA 0.0524f
C366 two_stage_opamp_dummy_magic_0.V_source.n23 GNDA 0.092237f
C367 two_stage_opamp_dummy_magic_0.V_source.t1 GNDA 0.014699f
C368 two_stage_opamp_dummy_magic_0.V_source.t14 GNDA 0.014699f
C369 two_stage_opamp_dummy_magic_0.V_source.n24 GNDA 0.0524f
C370 two_stage_opamp_dummy_magic_0.V_source.n25 GNDA 0.091747f
C371 two_stage_opamp_dummy_magic_0.V_source.t3 GNDA 0.014699f
C372 two_stage_opamp_dummy_magic_0.V_source.t11 GNDA 0.014699f
C373 two_stage_opamp_dummy_magic_0.V_source.n26 GNDA 0.052785f
C374 two_stage_opamp_dummy_magic_0.V_source.t19 GNDA 0.014699f
C375 two_stage_opamp_dummy_magic_0.V_source.t20 GNDA 0.014699f
C376 two_stage_opamp_dummy_magic_0.V_source.n27 GNDA 0.0524f
C377 two_stage_opamp_dummy_magic_0.V_source.n28 GNDA 0.175465f
C378 two_stage_opamp_dummy_magic_0.V_source.t2 GNDA 0.014699f
C379 two_stage_opamp_dummy_magic_0.V_source.t12 GNDA 0.014699f
C380 two_stage_opamp_dummy_magic_0.V_source.n29 GNDA 0.0524f
C381 two_stage_opamp_dummy_magic_0.V_source.n30 GNDA 0.092237f
C382 two_stage_opamp_dummy_magic_0.V_source.t15 GNDA 0.014699f
C383 two_stage_opamp_dummy_magic_0.V_source.t13 GNDA 0.014699f
C384 two_stage_opamp_dummy_magic_0.V_source.n31 GNDA 0.0524f
C385 two_stage_opamp_dummy_magic_0.V_source.n32 GNDA 0.092237f
C386 two_stage_opamp_dummy_magic_0.V_source.t4 GNDA 0.014699f
C387 two_stage_opamp_dummy_magic_0.V_source.t0 GNDA 0.014699f
C388 two_stage_opamp_dummy_magic_0.V_source.n33 GNDA 0.0524f
C389 two_stage_opamp_dummy_magic_0.V_source.n34 GNDA 0.140743f
C390 two_stage_opamp_dummy_magic_0.V_source.n35 GNDA 0.077414f
C391 two_stage_opamp_dummy_magic_0.V_source.n36 GNDA 0.082836f
C392 two_stage_opamp_dummy_magic_0.V_source.n37 GNDA 0.082155f
C393 two_stage_opamp_dummy_magic_0.V_source.n38 GNDA 0.09453f
C394 two_stage_opamp_dummy_magic_0.V_source.t38 GNDA 0.024498f
C395 bgr_0.cap_res2.t6 GNDA 0.406156f
C396 bgr_0.cap_res2.t2 GNDA 0.407628f
C397 bgr_0.cap_res2.t8 GNDA 0.406156f
C398 bgr_0.cap_res2.t13 GNDA 0.407628f
C399 bgr_0.cap_res2.t0 GNDA 0.406156f
C400 bgr_0.cap_res2.t19 GNDA 0.407628f
C401 bgr_0.cap_res2.t1 GNDA 0.406156f
C402 bgr_0.cap_res2.t5 GNDA 0.407628f
C403 bgr_0.cap_res2.t7 GNDA 0.406156f
C404 bgr_0.cap_res2.t4 GNDA 0.407628f
C405 bgr_0.cap_res2.t10 GNDA 0.406156f
C406 bgr_0.cap_res2.t14 GNDA 0.407628f
C407 bgr_0.cap_res2.t15 GNDA 0.406156f
C408 bgr_0.cap_res2.t12 GNDA 0.407628f
C409 bgr_0.cap_res2.t16 GNDA 0.406156f
C410 bgr_0.cap_res2.t18 GNDA 0.407628f
C411 bgr_0.cap_res2.n0 GNDA 0.272247f
C412 bgr_0.cap_res2.t17 GNDA 0.216805f
C413 bgr_0.cap_res2.n1 GNDA 0.295394f
C414 bgr_0.cap_res2.t11 GNDA 0.216805f
C415 bgr_0.cap_res2.n2 GNDA 0.295394f
C416 bgr_0.cap_res2.t3 GNDA 0.216805f
C417 bgr_0.cap_res2.n3 GNDA 0.295394f
C418 bgr_0.cap_res2.t9 GNDA 0.214043f
C419 bgr_0.cap_res2.t20 GNDA 0.133038f
C420 bgr_0.1st_Vout_2.n0 GNDA 0.995956f
C421 bgr_0.1st_Vout_2.n1 GNDA 0.240335f
C422 bgr_0.1st_Vout_2.n2 GNDA 0.995956f
C423 bgr_0.1st_Vout_2.n3 GNDA 0.240335f
C424 bgr_0.1st_Vout_2.n4 GNDA 0.805677f
C425 bgr_0.1st_Vout_2.n5 GNDA 0.240335f
C426 bgr_0.1st_Vout_2.t13 GNDA 0.021508f
C427 bgr_0.1st_Vout_2.n6 GNDA 0.02259f
C428 bgr_0.1st_Vout_2.n7 GNDA 0.171874f
C429 bgr_0.1st_Vout_2.t32 GNDA 0.013652f
C430 bgr_0.1st_Vout_2.t19 GNDA 0.013652f
C431 bgr_0.1st_Vout_2.n8 GNDA 0.03037f
C432 bgr_0.1st_Vout_2.n9 GNDA 0.083918f
C433 bgr_0.1st_Vout_2.n10 GNDA 0.012945f
C434 bgr_0.1st_Vout_2.t9 GNDA 0.018875f
C435 bgr_0.1st_Vout_2.n11 GNDA 0.195802f
C436 bgr_0.1st_Vout_2.n12 GNDA 0.011712f
C437 bgr_0.1st_Vout_2.n13 GNDA 0.049674f
C438 bgr_0.1st_Vout_2.n14 GNDA 0.021654f
C439 bgr_0.1st_Vout_2.n15 GNDA 0.080059f
C440 bgr_0.1st_Vout_2.n16 GNDA 0.03943f
C441 bgr_0.1st_Vout_2.t36 GNDA 0.013652f
C442 bgr_0.1st_Vout_2.t26 GNDA 0.013652f
C443 bgr_0.1st_Vout_2.n17 GNDA 0.03037f
C444 bgr_0.1st_Vout_2.n18 GNDA 0.083918f
C445 bgr_0.1st_Vout_2.t17 GNDA 0.364565f
C446 bgr_0.1st_Vout_2.t21 GNDA 0.358459f
C447 bgr_0.1st_Vout_2.t15 GNDA 0.358459f
C448 bgr_0.1st_Vout_2.t16 GNDA 0.364565f
C449 bgr_0.1st_Vout_2.t12 GNDA 0.358459f
C450 bgr_0.1st_Vout_2.t27 GNDA 0.364565f
C451 bgr_0.1st_Vout_2.t30 GNDA 0.358459f
C452 bgr_0.1st_Vout_2.t22 GNDA 0.358459f
C453 bgr_0.1st_Vout_2.t23 GNDA 0.364565f
C454 bgr_0.1st_Vout_2.t18 GNDA 0.358459f
C455 bgr_0.1st_Vout_2.t35 GNDA 0.364565f
C456 bgr_0.1st_Vout_2.t11 GNDA 0.358459f
C457 bgr_0.1st_Vout_2.t31 GNDA 0.358459f
C458 bgr_0.1st_Vout_2.t34 GNDA 0.364565f
C459 bgr_0.1st_Vout_2.t29 GNDA 0.358459f
C460 bgr_0.1st_Vout_2.t28 GNDA 0.364565f
C461 bgr_0.1st_Vout_2.t33 GNDA 0.358459f
C462 bgr_0.1st_Vout_2.t24 GNDA 0.358459f
C463 bgr_0.1st_Vout_2.t20 GNDA 0.358459f
C464 bgr_0.1st_Vout_2.t25 GNDA 0.358459f
C465 bgr_0.1st_Vout_2.t14 GNDA 0.023417f
C466 bgr_0.1st_Vout_2.n19 GNDA 0.516024f
C467 bgr_0.1st_Vout_2.n20 GNDA 0.106455f
C468 bgr_0.1st_Vout_2.n21 GNDA 0.02259f
C469 bgr_0.Vin+.t6 GNDA 0.020459f
C470 bgr_0.Vin+.t8 GNDA 0.013299f
C471 bgr_0.Vin+.n0 GNDA 0.04388f
C472 bgr_0.Vin+.t10 GNDA 0.013299f
C473 bgr_0.Vin+.n1 GNDA 0.034146f
C474 bgr_0.Vin+.t7 GNDA 0.013299f
C475 bgr_0.Vin+.n2 GNDA 0.034607f
C476 bgr_0.Vin+.n3 GNDA 0.074523f
C477 bgr_0.Vin+.t3 GNDA 0.043132f
C478 bgr_0.Vin+.t2 GNDA 0.043132f
C479 bgr_0.Vin+.n4 GNDA 0.144858f
C480 bgr_0.Vin+.t1 GNDA 0.043132f
C481 bgr_0.Vin+.t4 GNDA 0.043132f
C482 bgr_0.Vin+.n5 GNDA 0.142495f
C483 bgr_0.Vin+.n6 GNDA 0.656763f
C484 bgr_0.Vin+.n7 GNDA 0.71769f
C485 bgr_0.Vin+.t5 GNDA 0.137433f
C486 bgr_0.Vin+.n8 GNDA 0.446219f
C487 bgr_0.Vin+.t0 GNDA 0.125873f
C488 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t15 GNDA 0.028956f
C489 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t4 GNDA 0.028956f
C490 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n0 GNDA 0.072583f
C491 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t2 GNDA 0.028956f
C492 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t1 GNDA 0.028956f
C493 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n1 GNDA 0.0722f
C494 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n2 GNDA 0.641714f
C495 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t3 GNDA 0.028956f
C496 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t16 GNDA 0.028956f
C497 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n3 GNDA 0.057912f
C498 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n4 GNDA 0.323662f
C499 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t0 GNDA 0.370568f
C500 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t10 GNDA 0.057912f
C501 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t14 GNDA 0.057912f
C502 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n5 GNDA 0.169912f
C503 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t9 GNDA 0.057912f
C504 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t6 GNDA 0.057912f
C505 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n6 GNDA 0.169141f
C506 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n7 GNDA 0.584649f
C507 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t11 GNDA 0.057912f
C508 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t5 GNDA 0.057912f
C509 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n8 GNDA 0.169141f
C510 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n9 GNDA 0.302845f
C511 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t12 GNDA 0.057912f
C512 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t7 GNDA 0.057912f
C513 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n10 GNDA 0.169141f
C514 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n11 GNDA 0.302845f
C515 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t13 GNDA 0.057912f
C516 two_stage_opamp_dummy_magic_0.V_CMFB_S1.t8 GNDA 0.057912f
C517 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n12 GNDA 0.169141f
C518 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n13 GNDA 0.437166f
C519 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n14 GNDA 4.23853f
C520 two_stage_opamp_dummy_magic_0.V_CMFB_S1.n15 GNDA 4.54194f
C521 bgr_0.V_CMFB_S1 GNDA 0.054039f
C522 two_stage_opamp_dummy_magic_0.V_tot.t1 GNDA 0.164536f
C523 two_stage_opamp_dummy_magic_0.V_tot.t3 GNDA 0.17527f
C524 two_stage_opamp_dummy_magic_0.V_tot.t2 GNDA 0.164536f
C525 two_stage_opamp_dummy_magic_0.V_tot.n0 GNDA 0.845382f
C526 two_stage_opamp_dummy_magic_0.V_tot.n1 GNDA 0.038722f
C527 two_stage_opamp_dummy_magic_0.V_tot.n2 GNDA 0.038019f
C528 two_stage_opamp_dummy_magic_0.V_tot.n3 GNDA 0.211094f
C529 two_stage_opamp_dummy_magic_0.V_tot.t4 GNDA 0.019739f
C530 two_stage_opamp_dummy_magic_0.V_tot.n4 GNDA 0.115272f
C531 two_stage_opamp_dummy_magic_0.V_tot.t6 GNDA 0.019871f
C532 two_stage_opamp_dummy_magic_0.V_tot.n5 GNDA 0.032356f
C533 two_stage_opamp_dummy_magic_0.V_tot.n6 GNDA 0.189211f
C534 two_stage_opamp_dummy_magic_0.V_tot.n7 GNDA 0.038019f
C535 two_stage_opamp_dummy_magic_0.V_tot.n8 GNDA 0.135136f
C536 two_stage_opamp_dummy_magic_0.V_tot.n9 GNDA 0.15059f
C537 two_stage_opamp_dummy_magic_0.V_tot.n10 GNDA 1.37135f
C538 two_stage_opamp_dummy_magic_0.V_tot.n11 GNDA 0.846166f
C539 two_stage_opamp_dummy_magic_0.V_tot.t0 GNDA 0.17529f
C540 two_stage_opamp_dummy_magic_0.V_err_p.n0 GNDA 0.021118f
C541 two_stage_opamp_dummy_magic_0.V_err_p.n1 GNDA 0.020212f
C542 two_stage_opamp_dummy_magic_0.V_err_p.n2 GNDA 0.020262f
C543 two_stage_opamp_dummy_magic_0.V_err_p.n3 GNDA 0.021093f
C544 two_stage_opamp_dummy_magic_0.V_err_p.n4 GNDA 0.020966f
C545 two_stage_opamp_dummy_magic_0.V_err_p.n5 GNDA 0.297859f
C546 two_stage_opamp_dummy_magic_0.V_err_p.n6 GNDA 0.020966f
C547 two_stage_opamp_dummy_magic_0.V_err_p.n7 GNDA 0.155369f
C548 two_stage_opamp_dummy_magic_0.V_err_p.n8 GNDA 0.020966f
C549 two_stage_opamp_dummy_magic_0.V_err_p.n9 GNDA 0.189616f
C550 two_stage_opamp_dummy_magic_0.V_err_p.n10 GNDA 0.160506f
C551 two_stage_opamp_dummy_magic_0.V_err_p.n11 GNDA 0.14076f
C552 two_stage_opamp_dummy_magic_0.V_err_p.n12 GNDA 0.241198f
C553 two_stage_opamp_dummy_magic_0.V_err_p.n13 GNDA 0.021118f
C554 two_stage_opamp_dummy_magic_0.V_err_p.n14 GNDA 0.020826f
C555 two_stage_opamp_dummy_magic_0.V_err_p.n15 GNDA 0.326026f
C556 two_stage_opamp_dummy_magic_0.V_err_p.n16 GNDA 0.020826f
C557 two_stage_opamp_dummy_magic_0.V_err_p.n17 GNDA 0.179554f
C558 two_stage_opamp_dummy_magic_0.V_err_p.n18 GNDA 0.179554f
C559 two_stage_opamp_dummy_magic_0.V_err_p.n19 GNDA 0.020826f
C560 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t1 GNDA 0.169032f
C561 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t4 GNDA 0.422255f
C562 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t9 GNDA 0.422255f
C563 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t5 GNDA 0.50115f
C564 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n0 GNDA 0.264704f
C565 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n1 GNDA 0.167525f
C566 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t7 GNDA 0.460418f
C567 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n2 GNDA 0.15482f
C568 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n3 GNDA 0.888114f
C569 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t2 GNDA 0.460418f
C570 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t6 GNDA 0.422255f
C571 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t8 GNDA 0.422255f
C572 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t3 GNDA 0.50115f
C573 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n4 GNDA 0.264704f
C574 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n5 GNDA 0.167525f
C575 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n6 GNDA 0.15482f
C576 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.n7 GNDA 0.88757f
C577 two_stage_opamp_dummy_magic_0.V_b_2nd_stage.t0 GNDA 0.169032f
C578 two_stage_opamp_dummy_magic_0.V_tail_gate.t1 GNDA 0.028044f
C579 two_stage_opamp_dummy_magic_0.V_tail_gate.t6 GNDA 0.028044f
C580 two_stage_opamp_dummy_magic_0.V_tail_gate.n0 GNDA 0.067636f
C581 two_stage_opamp_dummy_magic_0.V_tail_gate.t5 GNDA 0.028044f
C582 two_stage_opamp_dummy_magic_0.V_tail_gate.t2 GNDA 0.028044f
C583 two_stage_opamp_dummy_magic_0.V_tail_gate.n1 GNDA 0.070203f
C584 two_stage_opamp_dummy_magic_0.V_tail_gate.t7 GNDA 0.028044f
C585 two_stage_opamp_dummy_magic_0.V_tail_gate.t4 GNDA 0.028044f
C586 two_stage_opamp_dummy_magic_0.V_tail_gate.n2 GNDA 0.069827f
C587 two_stage_opamp_dummy_magic_0.V_tail_gate.n3 GNDA 0.474137f
C588 two_stage_opamp_dummy_magic_0.V_tail_gate.t3 GNDA 0.028044f
C589 two_stage_opamp_dummy_magic_0.V_tail_gate.t0 GNDA 0.028044f
C590 two_stage_opamp_dummy_magic_0.V_tail_gate.n4 GNDA 0.070203f
C591 two_stage_opamp_dummy_magic_0.V_tail_gate.n5 GNDA 0.311197f
C592 two_stage_opamp_dummy_magic_0.V_tail_gate.n6 GNDA 0.721672f
C593 two_stage_opamp_dummy_magic_0.V_tail_gate.t9 GNDA 0.042066f
C594 two_stage_opamp_dummy_magic_0.V_tail_gate.t8 GNDA 0.042066f
C595 two_stage_opamp_dummy_magic_0.V_tail_gate.n7 GNDA 0.152234f
C596 two_stage_opamp_dummy_magic_0.V_tail_gate.t31 GNDA 0.074668f
C597 two_stage_opamp_dummy_magic_0.V_tail_gate.t22 GNDA 0.074668f
C598 two_stage_opamp_dummy_magic_0.V_tail_gate.t28 GNDA 0.074668f
C599 two_stage_opamp_dummy_magic_0.V_tail_gate.t18 GNDA 0.074668f
C600 two_stage_opamp_dummy_magic_0.V_tail_gate.t26 GNDA 0.074668f
C601 two_stage_opamp_dummy_magic_0.V_tail_gate.t16 GNDA 0.074668f
C602 two_stage_opamp_dummy_magic_0.V_tail_gate.t24 GNDA 0.074668f
C603 two_stage_opamp_dummy_magic_0.V_tail_gate.t13 GNDA 0.074668f
C604 two_stage_opamp_dummy_magic_0.V_tail_gate.t20 GNDA 0.074668f
C605 two_stage_opamp_dummy_magic_0.V_tail_gate.t14 GNDA 0.087149f
C606 two_stage_opamp_dummy_magic_0.V_tail_gate.n8 GNDA 0.082168f
C607 two_stage_opamp_dummy_magic_0.V_tail_gate.n9 GNDA 0.051531f
C608 two_stage_opamp_dummy_magic_0.V_tail_gate.n10 GNDA 0.051531f
C609 two_stage_opamp_dummy_magic_0.V_tail_gate.n11 GNDA 0.051531f
C610 two_stage_opamp_dummy_magic_0.V_tail_gate.n12 GNDA 0.051531f
C611 two_stage_opamp_dummy_magic_0.V_tail_gate.n13 GNDA 0.051531f
C612 two_stage_opamp_dummy_magic_0.V_tail_gate.n14 GNDA 0.051531f
C613 two_stage_opamp_dummy_magic_0.V_tail_gate.n15 GNDA 0.051531f
C614 two_stage_opamp_dummy_magic_0.V_tail_gate.n16 GNDA 0.046048f
C615 two_stage_opamp_dummy_magic_0.V_tail_gate.t19 GNDA 0.074668f
C616 two_stage_opamp_dummy_magic_0.V_tail_gate.t29 GNDA 0.074668f
C617 two_stage_opamp_dummy_magic_0.V_tail_gate.t23 GNDA 0.074668f
C618 two_stage_opamp_dummy_magic_0.V_tail_gate.t15 GNDA 0.074668f
C619 two_stage_opamp_dummy_magic_0.V_tail_gate.t25 GNDA 0.074668f
C620 two_stage_opamp_dummy_magic_0.V_tail_gate.t17 GNDA 0.074668f
C621 two_stage_opamp_dummy_magic_0.V_tail_gate.t27 GNDA 0.074668f
C622 two_stage_opamp_dummy_magic_0.V_tail_gate.t21 GNDA 0.074668f
C623 two_stage_opamp_dummy_magic_0.V_tail_gate.t30 GNDA 0.074668f
C624 two_stage_opamp_dummy_magic_0.V_tail_gate.t12 GNDA 0.087149f
C625 two_stage_opamp_dummy_magic_0.V_tail_gate.n17 GNDA 0.082168f
C626 two_stage_opamp_dummy_magic_0.V_tail_gate.n18 GNDA 0.051531f
C627 two_stage_opamp_dummy_magic_0.V_tail_gate.n19 GNDA 0.051531f
C628 two_stage_opamp_dummy_magic_0.V_tail_gate.n20 GNDA 0.051531f
C629 two_stage_opamp_dummy_magic_0.V_tail_gate.n21 GNDA 0.051531f
C630 two_stage_opamp_dummy_magic_0.V_tail_gate.n22 GNDA 0.051531f
C631 two_stage_opamp_dummy_magic_0.V_tail_gate.n23 GNDA 0.051531f
C632 two_stage_opamp_dummy_magic_0.V_tail_gate.n24 GNDA 0.051531f
C633 two_stage_opamp_dummy_magic_0.V_tail_gate.n25 GNDA 0.046048f
C634 two_stage_opamp_dummy_magic_0.V_tail_gate.n26 GNDA 0.115078f
C635 two_stage_opamp_dummy_magic_0.V_tail_gate.t11 GNDA 0.042066f
C636 two_stage_opamp_dummy_magic_0.V_tail_gate.t10 GNDA 0.042066f
C637 two_stage_opamp_dummy_magic_0.V_tail_gate.n27 GNDA 0.084132f
C638 two_stage_opamp_dummy_magic_0.V_tail_gate.n28 GNDA 0.326114f
C639 two_stage_opamp_dummy_magic_0.V_tail_gate.n29 GNDA 3.33293f
C640 bgr_0.TAIL_CUR_MIR_BIAS GNDA 3.71584f
C641 two_stage_opamp_dummy_magic_0.cap_res_X.t90 GNDA 0.344645f
C642 two_stage_opamp_dummy_magic_0.cap_res_X.t127 GNDA 0.345894f
C643 two_stage_opamp_dummy_magic_0.cap_res_X.t49 GNDA 0.344645f
C644 two_stage_opamp_dummy_magic_0.cap_res_X.t88 GNDA 0.347347f
C645 two_stage_opamp_dummy_magic_0.cap_res_X.t67 GNDA 0.37779f
C646 two_stage_opamp_dummy_magic_0.cap_res_X.t130 GNDA 0.344645f
C647 two_stage_opamp_dummy_magic_0.cap_res_X.t27 GNDA 0.345894f
C648 two_stage_opamp_dummy_magic_0.cap_res_X.t81 GNDA 0.344645f
C649 two_stage_opamp_dummy_magic_0.cap_res_X.t42 GNDA 0.345894f
C650 two_stage_opamp_dummy_magic_0.cap_res_X.t95 GNDA 0.344645f
C651 two_stage_opamp_dummy_magic_0.cap_res_X.t134 GNDA 0.345894f
C652 two_stage_opamp_dummy_magic_0.cap_res_X.t45 GNDA 0.344645f
C653 two_stage_opamp_dummy_magic_0.cap_res_X.t9 GNDA 0.345894f
C654 two_stage_opamp_dummy_magic_0.cap_res_X.t43 GNDA 0.344645f
C655 two_stage_opamp_dummy_magic_0.cap_res_X.t79 GNDA 0.345894f
C656 two_stage_opamp_dummy_magic_0.cap_res_X.t58 GNDA 0.344645f
C657 two_stage_opamp_dummy_magic_0.cap_res_X.t25 GNDA 0.345894f
C658 two_stage_opamp_dummy_magic_0.cap_res_X.t83 GNDA 0.344645f
C659 two_stage_opamp_dummy_magic_0.cap_res_X.t118 GNDA 0.345894f
C660 two_stage_opamp_dummy_magic_0.cap_res_X.t102 GNDA 0.344645f
C661 two_stage_opamp_dummy_magic_0.cap_res_X.t65 GNDA 0.345894f
C662 two_stage_opamp_dummy_magic_0.cap_res_X.t48 GNDA 0.344645f
C663 two_stage_opamp_dummy_magic_0.cap_res_X.t86 GNDA 0.345894f
C664 two_stage_opamp_dummy_magic_0.cap_res_X.t66 GNDA 0.344645f
C665 two_stage_opamp_dummy_magic_0.cap_res_X.t31 GNDA 0.345894f
C666 two_stage_opamp_dummy_magic_0.cap_res_X.t89 GNDA 0.344645f
C667 two_stage_opamp_dummy_magic_0.cap_res_X.t124 GNDA 0.345894f
C668 two_stage_opamp_dummy_magic_0.cap_res_X.t105 GNDA 0.344645f
C669 two_stage_opamp_dummy_magic_0.cap_res_X.t69 GNDA 0.345894f
C670 two_stage_opamp_dummy_magic_0.cap_res_X.t128 GNDA 0.344645f
C671 two_stage_opamp_dummy_magic_0.cap_res_X.t22 GNDA 0.345894f
C672 two_stage_opamp_dummy_magic_0.cap_res_X.t4 GNDA 0.344645f
C673 two_stage_opamp_dummy_magic_0.cap_res_X.t109 GNDA 0.345894f
C674 two_stage_opamp_dummy_magic_0.cap_res_X.t94 GNDA 0.344645f
C675 two_stage_opamp_dummy_magic_0.cap_res_X.t129 GNDA 0.345894f
C676 two_stage_opamp_dummy_magic_0.cap_res_X.t111 GNDA 0.344645f
C677 two_stage_opamp_dummy_magic_0.cap_res_X.t76 GNDA 0.345894f
C678 two_stage_opamp_dummy_magic_0.cap_res_X.t135 GNDA 0.344645f
C679 two_stage_opamp_dummy_magic_0.cap_res_X.t28 GNDA 0.345894f
C680 two_stage_opamp_dummy_magic_0.cap_res_X.t11 GNDA 0.344645f
C681 two_stage_opamp_dummy_magic_0.cap_res_X.t117 GNDA 0.345894f
C682 two_stage_opamp_dummy_magic_0.cap_res_X.t34 GNDA 0.344645f
C683 two_stage_opamp_dummy_magic_0.cap_res_X.t68 GNDA 0.345894f
C684 two_stage_opamp_dummy_magic_0.cap_res_X.t50 GNDA 0.344645f
C685 two_stage_opamp_dummy_magic_0.cap_res_X.t16 GNDA 0.345894f
C686 two_stage_opamp_dummy_magic_0.cap_res_X.t73 GNDA 0.344645f
C687 two_stage_opamp_dummy_magic_0.cap_res_X.t108 GNDA 0.345894f
C688 two_stage_opamp_dummy_magic_0.cap_res_X.t91 GNDA 0.344645f
C689 two_stage_opamp_dummy_magic_0.cap_res_X.t54 GNDA 0.345894f
C690 two_stage_opamp_dummy_magic_0.cap_res_X.t36 GNDA 0.344645f
C691 two_stage_opamp_dummy_magic_0.cap_res_X.t74 GNDA 0.345894f
C692 two_stage_opamp_dummy_magic_0.cap_res_X.t53 GNDA 0.344645f
C693 two_stage_opamp_dummy_magic_0.cap_res_X.t20 GNDA 0.345894f
C694 two_stage_opamp_dummy_magic_0.cap_res_X.t78 GNDA 0.344645f
C695 two_stage_opamp_dummy_magic_0.cap_res_X.t116 GNDA 0.345894f
C696 two_stage_opamp_dummy_magic_0.cap_res_X.t97 GNDA 0.344645f
C697 two_stage_opamp_dummy_magic_0.cap_res_X.t57 GNDA 0.345894f
C698 two_stage_opamp_dummy_magic_0.cap_res_X.t120 GNDA 0.344645f
C699 two_stage_opamp_dummy_magic_0.cap_res_X.t15 GNDA 0.345894f
C700 two_stage_opamp_dummy_magic_0.cap_res_X.t137 GNDA 0.344645f
C701 two_stage_opamp_dummy_magic_0.cap_res_X.t100 GNDA 0.345894f
C702 two_stage_opamp_dummy_magic_0.cap_res_X.t85 GNDA 0.344645f
C703 two_stage_opamp_dummy_magic_0.cap_res_X.t119 GNDA 0.345894f
C704 two_stage_opamp_dummy_magic_0.cap_res_X.t84 GNDA 0.344645f
C705 two_stage_opamp_dummy_magic_0.cap_res_X.t8 GNDA 0.361543f
C706 two_stage_opamp_dummy_magic_0.cap_res_X.t41 GNDA 0.344645f
C707 two_stage_opamp_dummy_magic_0.cap_res_X.t99 GNDA 0.185116f
C708 two_stage_opamp_dummy_magic_0.cap_res_X.n0 GNDA 0.19812f
C709 two_stage_opamp_dummy_magic_0.cap_res_X.t93 GNDA 0.344645f
C710 two_stage_opamp_dummy_magic_0.cap_res_X.t60 GNDA 0.185116f
C711 two_stage_opamp_dummy_magic_0.cap_res_X.n1 GNDA 0.196522f
C712 two_stage_opamp_dummy_magic_0.cap_res_X.t3 GNDA 0.344645f
C713 two_stage_opamp_dummy_magic_0.cap_res_X.t26 GNDA 0.185116f
C714 two_stage_opamp_dummy_magic_0.cap_res_X.n2 GNDA 0.196522f
C715 two_stage_opamp_dummy_magic_0.cap_res_X.t51 GNDA 0.344645f
C716 two_stage_opamp_dummy_magic_0.cap_res_X.t133 GNDA 0.185116f
C717 two_stage_opamp_dummy_magic_0.cap_res_X.n3 GNDA 0.196522f
C718 two_stage_opamp_dummy_magic_0.cap_res_X.t14 GNDA 0.344645f
C719 two_stage_opamp_dummy_magic_0.cap_res_X.t82 GNDA 0.185116f
C720 two_stage_opamp_dummy_magic_0.cap_res_X.n4 GNDA 0.196522f
C721 two_stage_opamp_dummy_magic_0.cap_res_X.t61 GNDA 0.344645f
C722 two_stage_opamp_dummy_magic_0.cap_res_X.t44 GNDA 0.185116f
C723 two_stage_opamp_dummy_magic_0.cap_res_X.n5 GNDA 0.196522f
C724 two_stage_opamp_dummy_magic_0.cap_res_X.t115 GNDA 0.344645f
C725 two_stage_opamp_dummy_magic_0.cap_res_X.t13 GNDA 0.185116f
C726 two_stage_opamp_dummy_magic_0.cap_res_X.n6 GNDA 0.196522f
C727 two_stage_opamp_dummy_magic_0.cap_res_X.t71 GNDA 0.344645f
C728 two_stage_opamp_dummy_magic_0.cap_res_X.t103 GNDA 0.185116f
C729 two_stage_opamp_dummy_magic_0.cap_res_X.n7 GNDA 0.196522f
C730 two_stage_opamp_dummy_magic_0.cap_res_X.t123 GNDA 0.344645f
C731 two_stage_opamp_dummy_magic_0.cap_res_X.t63 GNDA 0.185116f
C732 two_stage_opamp_dummy_magic_0.cap_res_X.n8 GNDA 0.196522f
C733 two_stage_opamp_dummy_magic_0.cap_res_X.t40 GNDA 0.344645f
C734 two_stage_opamp_dummy_magic_0.cap_res_X.t132 GNDA 0.345894f
C735 two_stage_opamp_dummy_magic_0.cap_res_X.t33 GNDA 0.166619f
C736 two_stage_opamp_dummy_magic_0.cap_res_X.n9 GNDA 0.214914f
C737 two_stage_opamp_dummy_magic_0.cap_res_X.t30 GNDA 0.18397f
C738 two_stage_opamp_dummy_magic_0.cap_res_X.n10 GNDA 0.23341f
C739 two_stage_opamp_dummy_magic_0.cap_res_X.t64 GNDA 0.18397f
C740 two_stage_opamp_dummy_magic_0.cap_res_X.n11 GNDA 0.250658f
C741 two_stage_opamp_dummy_magic_0.cap_res_X.t24 GNDA 0.18397f
C742 two_stage_opamp_dummy_magic_0.cap_res_X.n12 GNDA 0.250658f
C743 two_stage_opamp_dummy_magic_0.cap_res_X.t126 GNDA 0.18397f
C744 two_stage_opamp_dummy_magic_0.cap_res_X.n13 GNDA 0.250658f
C745 two_stage_opamp_dummy_magic_0.cap_res_X.t19 GNDA 0.18397f
C746 two_stage_opamp_dummy_magic_0.cap_res_X.n14 GNDA 0.250658f
C747 two_stage_opamp_dummy_magic_0.cap_res_X.t122 GNDA 0.18397f
C748 two_stage_opamp_dummy_magic_0.cap_res_X.n15 GNDA 0.250658f
C749 two_stage_opamp_dummy_magic_0.cap_res_X.t80 GNDA 0.18397f
C750 two_stage_opamp_dummy_magic_0.cap_res_X.n16 GNDA 0.250658f
C751 two_stage_opamp_dummy_magic_0.cap_res_X.t37 GNDA 0.18397f
C752 two_stage_opamp_dummy_magic_0.cap_res_X.n17 GNDA 0.250658f
C753 two_stage_opamp_dummy_magic_0.cap_res_X.t75 GNDA 0.18397f
C754 two_stage_opamp_dummy_magic_0.cap_res_X.n18 GNDA 0.250658f
C755 two_stage_opamp_dummy_magic_0.cap_res_X.t35 GNDA 0.18397f
C756 two_stage_opamp_dummy_magic_0.cap_res_X.n19 GNDA 0.250658f
C757 two_stage_opamp_dummy_magic_0.cap_res_X.t138 GNDA 0.18397f
C758 two_stage_opamp_dummy_magic_0.cap_res_X.n20 GNDA 0.250658f
C759 two_stage_opamp_dummy_magic_0.cap_res_X.t29 GNDA 0.18397f
C760 two_stage_opamp_dummy_magic_0.cap_res_X.n21 GNDA 0.250658f
C761 two_stage_opamp_dummy_magic_0.cap_res_X.t131 GNDA 0.18397f
C762 two_stage_opamp_dummy_magic_0.cap_res_X.n22 GNDA 0.250658f
C763 two_stage_opamp_dummy_magic_0.cap_res_X.t110 GNDA 0.18397f
C764 two_stage_opamp_dummy_magic_0.cap_res_X.n23 GNDA 0.250658f
C765 two_stage_opamp_dummy_magic_0.cap_res_X.t5 GNDA 0.18397f
C766 two_stage_opamp_dummy_magic_0.cap_res_X.n24 GNDA 0.250658f
C767 two_stage_opamp_dummy_magic_0.cap_res_X.t106 GNDA 0.18397f
C768 two_stage_opamp_dummy_magic_0.cap_res_X.n25 GNDA 0.23341f
C769 two_stage_opamp_dummy_magic_0.cap_res_X.t104 GNDA 0.343499f
C770 two_stage_opamp_dummy_magic_0.cap_res_X.t2 GNDA 0.166619f
C771 two_stage_opamp_dummy_magic_0.cap_res_X.n26 GNDA 0.216163f
C772 two_stage_opamp_dummy_magic_0.cap_res_X.t1 GNDA 0.343499f
C773 two_stage_opamp_dummy_magic_0.cap_res_X.t38 GNDA 0.166619f
C774 two_stage_opamp_dummy_magic_0.cap_res_X.n27 GNDA 0.216163f
C775 two_stage_opamp_dummy_magic_0.cap_res_X.t121 GNDA 0.343499f
C776 two_stage_opamp_dummy_magic_0.cap_res_X.t113 GNDA 0.344645f
C777 two_stage_opamp_dummy_magic_0.cap_res_X.t21 GNDA 0.363141f
C778 two_stage_opamp_dummy_magic_0.cap_res_X.t56 GNDA 0.363141f
C779 two_stage_opamp_dummy_magic_0.cap_res_X.t18 GNDA 0.185116f
C780 two_stage_opamp_dummy_magic_0.cap_res_X.n28 GNDA 0.216163f
C781 two_stage_opamp_dummy_magic_0.cap_res_X.t125 GNDA 0.343499f
C782 two_stage_opamp_dummy_magic_0.cap_res_X.t62 GNDA 0.344645f
C783 two_stage_opamp_dummy_magic_0.cap_res_X.t23 GNDA 0.185116f
C784 two_stage_opamp_dummy_magic_0.cap_res_X.n29 GNDA 0.197667f
C785 two_stage_opamp_dummy_magic_0.cap_res_X.t7 GNDA 0.343499f
C786 two_stage_opamp_dummy_magic_0.cap_res_X.t87 GNDA 0.344645f
C787 two_stage_opamp_dummy_magic_0.cap_res_X.t46 GNDA 0.185116f
C788 two_stage_opamp_dummy_magic_0.cap_res_X.n30 GNDA 0.216163f
C789 two_stage_opamp_dummy_magic_0.cap_res_X.t107 GNDA 0.343499f
C790 two_stage_opamp_dummy_magic_0.cap_res_X.t47 GNDA 0.344645f
C791 two_stage_opamp_dummy_magic_0.cap_res_X.t10 GNDA 0.185116f
C792 two_stage_opamp_dummy_magic_0.cap_res_X.n31 GNDA 0.216163f
C793 two_stage_opamp_dummy_magic_0.cap_res_X.t70 GNDA 0.343499f
C794 two_stage_opamp_dummy_magic_0.cap_res_X.t12 GNDA 0.344645f
C795 two_stage_opamp_dummy_magic_0.cap_res_X.t112 GNDA 0.185116f
C796 two_stage_opamp_dummy_magic_0.cap_res_X.n32 GNDA 0.216163f
C797 two_stage_opamp_dummy_magic_0.cap_res_X.t32 GNDA 0.343499f
C798 two_stage_opamp_dummy_magic_0.cap_res_X.t92 GNDA 0.344645f
C799 two_stage_opamp_dummy_magic_0.cap_res_X.t77 GNDA 0.363141f
C800 two_stage_opamp_dummy_magic_0.cap_res_X.t114 GNDA 0.363141f
C801 two_stage_opamp_dummy_magic_0.cap_res_X.t72 GNDA 0.185116f
C802 two_stage_opamp_dummy_magic_0.cap_res_X.n33 GNDA 0.216163f
C803 two_stage_opamp_dummy_magic_0.cap_res_X.t52 GNDA 0.343499f
C804 two_stage_opamp_dummy_magic_0.cap_res_X.t39 GNDA 0.344645f
C805 two_stage_opamp_dummy_magic_0.cap_res_X.t101 GNDA 0.363141f
C806 two_stage_opamp_dummy_magic_0.cap_res_X.t136 GNDA 0.363141f
C807 two_stage_opamp_dummy_magic_0.cap_res_X.t96 GNDA 0.185116f
C808 two_stage_opamp_dummy_magic_0.cap_res_X.n34 GNDA 0.216163f
C809 two_stage_opamp_dummy_magic_0.cap_res_X.t17 GNDA 0.343499f
C810 two_stage_opamp_dummy_magic_0.cap_res_X.n35 GNDA 0.216163f
C811 two_stage_opamp_dummy_magic_0.cap_res_X.t55 GNDA 0.185116f
C812 two_stage_opamp_dummy_magic_0.cap_res_X.t98 GNDA 0.363141f
C813 two_stage_opamp_dummy_magic_0.cap_res_X.t59 GNDA 0.363141f
C814 two_stage_opamp_dummy_magic_0.cap_res_X.t6 GNDA 0.764814f
C815 two_stage_opamp_dummy_magic_0.cap_res_X.t0 GNDA 0.3034f
C816 bgr_0.V_mir1.t8 GNDA 0.053881f
C817 bgr_0.V_mir1.t6 GNDA 0.042444f
C818 bgr_0.V_mir1.t17 GNDA 0.042444f
C819 bgr_0.V_mir1.t20 GNDA 0.06851f
C820 bgr_0.V_mir1.n0 GNDA 0.076506f
C821 bgr_0.V_mir1.n1 GNDA 0.052264f
C822 bgr_0.V_mir1.n2 GNDA 0.081315f
C823 bgr_0.V_mir1.t9 GNDA 0.03537f
C824 bgr_0.V_mir1.t7 GNDA 0.03537f
C825 bgr_0.V_mir1.n3 GNDA 0.08097f
C826 bgr_0.V_mir1.n4 GNDA 0.203577f
C827 bgr_0.V_mir1.t15 GNDA 0.017685f
C828 bgr_0.V_mir1.t13 GNDA 0.017685f
C829 bgr_0.V_mir1.n5 GNDA 0.046242f
C830 bgr_0.V_mir1.t14 GNDA 0.075466f
C831 bgr_0.V_mir1.t16 GNDA 0.017685f
C832 bgr_0.V_mir1.t12 GNDA 0.017685f
C833 bgr_0.V_mir1.n6 GNDA 0.050199f
C834 bgr_0.V_mir1.n7 GNDA 0.827814f
C835 bgr_0.V_mir1.n8 GNDA 0.268286f
C836 bgr_0.V_mir1.t0 GNDA 0.053881f
C837 bgr_0.V_mir1.t4 GNDA 0.042444f
C838 bgr_0.V_mir1.t18 GNDA 0.042444f
C839 bgr_0.V_mir1.t21 GNDA 0.06851f
C840 bgr_0.V_mir1.n9 GNDA 0.076506f
C841 bgr_0.V_mir1.n10 GNDA 0.052264f
C842 bgr_0.V_mir1.n11 GNDA 0.081315f
C843 bgr_0.V_mir1.t1 GNDA 0.03537f
C844 bgr_0.V_mir1.t5 GNDA 0.03537f
C845 bgr_0.V_mir1.n12 GNDA 0.08097f
C846 bgr_0.V_mir1.n13 GNDA 0.156007f
C847 bgr_0.V_mir1.n14 GNDA 0.09373f
C848 bgr_0.V_mir1.n15 GNDA 0.699157f
C849 bgr_0.V_mir1.t10 GNDA 0.053881f
C850 bgr_0.V_mir1.t2 GNDA 0.042444f
C851 bgr_0.V_mir1.t19 GNDA 0.042444f
C852 bgr_0.V_mir1.t22 GNDA 0.06851f
C853 bgr_0.V_mir1.n16 GNDA 0.076506f
C854 bgr_0.V_mir1.n17 GNDA 0.052264f
C855 bgr_0.V_mir1.n18 GNDA 0.081315f
C856 bgr_0.V_mir1.n19 GNDA 0.201563f
C857 bgr_0.V_mir1.t3 GNDA 0.03537f
C858 bgr_0.V_mir1.n20 GNDA 0.08097f
C859 bgr_0.V_mir1.t11 GNDA 0.03537f
C860 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t0 GNDA 0.472675f
C861 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t6 GNDA 0.113969f
C862 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t10 GNDA 0.113969f
C863 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n0 GNDA 0.471306f
C864 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t5 GNDA 0.113969f
C865 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t12 GNDA 0.113969f
C866 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n1 GNDA 0.469498f
C867 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n2 GNDA 0.650959f
C868 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t7 GNDA 0.113969f
C869 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t11 GNDA 0.113969f
C870 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n3 GNDA 0.469498f
C871 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n4 GNDA 0.33968f
C872 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t8 GNDA 0.113969f
C873 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t13 GNDA 0.113969f
C874 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n5 GNDA 0.469498f
C875 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n6 GNDA 0.33968f
C876 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t9 GNDA 0.113969f
C877 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t4 GNDA 0.113969f
C878 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n7 GNDA 0.469498f
C879 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n8 GNDA 0.491019f
C880 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n9 GNDA 7.25939f
C881 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t2 GNDA 0.03799f
C882 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t1 GNDA 0.03799f
C883 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n10 GNDA 0.115079f
C884 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t3 GNDA 0.03799f
C885 two_stage_opamp_dummy_magic_0.V_CMFB_S2.t14 GNDA 0.03799f
C886 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n11 GNDA 0.143458f
C887 two_stage_opamp_dummy_magic_0.V_CMFB_S2.n12 GNDA 0.834929f
C888 bgr_0.V_CMFB_S2 GNDA 5.91219f
C889 bgr_0.PFET_GATE_10uA.t23 GNDA 0.039433f
C890 bgr_0.PFET_GATE_10uA.t16 GNDA 0.058292f
C891 bgr_0.PFET_GATE_10uA.n0 GNDA 0.064232f
C892 bgr_0.PFET_GATE_10uA.t29 GNDA 0.039433f
C893 bgr_0.PFET_GATE_10uA.t17 GNDA 0.058292f
C894 bgr_0.PFET_GATE_10uA.n1 GNDA 0.064232f
C895 bgr_0.PFET_GATE_10uA.n2 GNDA 0.077289f
C896 bgr_0.PFET_GATE_10uA.t10 GNDA 0.039433f
C897 bgr_0.PFET_GATE_10uA.t24 GNDA 0.058292f
C898 bgr_0.PFET_GATE_10uA.n3 GNDA 0.064232f
C899 bgr_0.PFET_GATE_10uA.t18 GNDA 0.039433f
C900 bgr_0.PFET_GATE_10uA.t25 GNDA 0.058292f
C901 bgr_0.PFET_GATE_10uA.n4 GNDA 0.064232f
C902 bgr_0.PFET_GATE_10uA.n5 GNDA 0.064438f
C903 bgr_0.PFET_GATE_10uA.t3 GNDA 0.786496f
C904 bgr_0.PFET_GATE_10uA.t7 GNDA 0.590788f
C905 bgr_0.PFET_GATE_10uA.t2 GNDA 0.040444f
C906 bgr_0.PFET_GATE_10uA.t6 GNDA 0.040444f
C907 bgr_0.PFET_GATE_10uA.n6 GNDA 0.103372f
C908 bgr_0.PFET_GATE_10uA.t8 GNDA 0.040444f
C909 bgr_0.PFET_GATE_10uA.t1 GNDA 0.040444f
C910 bgr_0.PFET_GATE_10uA.n7 GNDA 0.100701f
C911 bgr_0.PFET_GATE_10uA.n8 GNDA 0.984984f
C912 bgr_0.PFET_GATE_10uA.t4 GNDA 0.040444f
C913 bgr_0.PFET_GATE_10uA.t0 GNDA 0.040444f
C914 bgr_0.PFET_GATE_10uA.n9 GNDA 0.100701f
C915 bgr_0.PFET_GATE_10uA.n10 GNDA 0.558538f
C916 bgr_0.PFET_GATE_10uA.n11 GNDA 1.14022f
C917 bgr_0.PFET_GATE_10uA.t5 GNDA 0.040444f
C918 bgr_0.PFET_GATE_10uA.t9 GNDA 0.040444f
C919 bgr_0.PFET_GATE_10uA.n12 GNDA 0.097542f
C920 bgr_0.PFET_GATE_10uA.n13 GNDA 0.358998f
C921 bgr_0.PFET_GATE_10uA.n14 GNDA 3.87496f
C922 bgr_0.PFET_GATE_10uA.t13 GNDA 0.045593f
C923 bgr_0.PFET_GATE_10uA.t21 GNDA 0.045593f
C924 bgr_0.PFET_GATE_10uA.n15 GNDA 0.138029f
C925 bgr_0.PFET_GATE_10uA.n16 GNDA 1.80019f
C926 bgr_0.PFET_GATE_10uA.n17 GNDA 1.42645f
C927 bgr_0.PFET_GATE_10uA.t27 GNDA 0.039433f
C928 bgr_0.PFET_GATE_10uA.t20 GNDA 0.039433f
C929 bgr_0.PFET_GATE_10uA.t12 GNDA 0.039433f
C930 bgr_0.PFET_GATE_10uA.t26 GNDA 0.039433f
C931 bgr_0.PFET_GATE_10uA.t19 GNDA 0.039433f
C932 bgr_0.PFET_GATE_10uA.t11 GNDA 0.058292f
C933 bgr_0.PFET_GATE_10uA.n18 GNDA 0.07214f
C934 bgr_0.PFET_GATE_10uA.n19 GNDA 0.051566f
C935 bgr_0.PFET_GATE_10uA.n20 GNDA 0.051566f
C936 bgr_0.PFET_GATE_10uA.n21 GNDA 0.051566f
C937 bgr_0.PFET_GATE_10uA.n22 GNDA 0.043658f
C938 bgr_0.PFET_GATE_10uA.t14 GNDA 0.039433f
C939 bgr_0.PFET_GATE_10uA.t22 GNDA 0.039433f
C940 bgr_0.PFET_GATE_10uA.t28 GNDA 0.039433f
C941 bgr_0.PFET_GATE_10uA.t15 GNDA 0.058292f
C942 bgr_0.PFET_GATE_10uA.n23 GNDA 0.07214f
C943 bgr_0.PFET_GATE_10uA.n24 GNDA 0.051566f
C944 bgr_0.PFET_GATE_10uA.n25 GNDA 0.043658f
C945 bgr_0.PFET_GATE_10uA.n26 GNDA 0.059927f
C946 two_stage_opamp_dummy_magic_0.VOUT-.t15 GNDA 0.043622f
C947 two_stage_opamp_dummy_magic_0.VOUT-.t10 GNDA 0.043622f
C948 two_stage_opamp_dummy_magic_0.VOUT-.n0 GNDA 0.175328f
C949 two_stage_opamp_dummy_magic_0.VOUT-.t5 GNDA 0.043622f
C950 two_stage_opamp_dummy_magic_0.VOUT-.t9 GNDA 0.043622f
C951 two_stage_opamp_dummy_magic_0.VOUT-.n1 GNDA 0.175005f
C952 two_stage_opamp_dummy_magic_0.VOUT-.n2 GNDA 0.1724f
C953 two_stage_opamp_dummy_magic_0.VOUT-.t4 GNDA 0.043622f
C954 two_stage_opamp_dummy_magic_0.VOUT-.t8 GNDA 0.043622f
C955 two_stage_opamp_dummy_magic_0.VOUT-.n3 GNDA 0.175005f
C956 two_stage_opamp_dummy_magic_0.VOUT-.n4 GNDA 0.088906f
C957 two_stage_opamp_dummy_magic_0.VOUT-.t12 GNDA 0.043622f
C958 two_stage_opamp_dummy_magic_0.VOUT-.t6 GNDA 0.043622f
C959 two_stage_opamp_dummy_magic_0.VOUT-.n5 GNDA 0.175005f
C960 two_stage_opamp_dummy_magic_0.VOUT-.n6 GNDA 0.088906f
C961 two_stage_opamp_dummy_magic_0.VOUT-.t11 GNDA 0.043622f
C962 two_stage_opamp_dummy_magic_0.VOUT-.t16 GNDA 0.043622f
C963 two_stage_opamp_dummy_magic_0.VOUT-.n7 GNDA 0.175327f
C964 two_stage_opamp_dummy_magic_0.VOUT-.n8 GNDA 0.105305f
C965 two_stage_opamp_dummy_magic_0.VOUT-.t13 GNDA 0.043622f
C966 two_stage_opamp_dummy_magic_0.VOUT-.t7 GNDA 0.043622f
C967 two_stage_opamp_dummy_magic_0.VOUT-.n9 GNDA 0.172862f
C968 two_stage_opamp_dummy_magic_0.VOUT-.n10 GNDA 0.212252f
C969 two_stage_opamp_dummy_magic_0.VOUT-.t117 GNDA 0.295764f
C970 two_stage_opamp_dummy_magic_0.VOUT-.t25 GNDA 0.290811f
C971 two_stage_opamp_dummy_magic_0.VOUT-.n11 GNDA 0.194979f
C972 two_stage_opamp_dummy_magic_0.VOUT-.t124 GNDA 0.290811f
C973 two_stage_opamp_dummy_magic_0.VOUT-.n12 GNDA 0.12723f
C974 two_stage_opamp_dummy_magic_0.VOUT-.t72 GNDA 0.295764f
C975 two_stage_opamp_dummy_magic_0.VOUT-.t38 GNDA 0.290811f
C976 two_stage_opamp_dummy_magic_0.VOUT-.n13 GNDA 0.194979f
C977 two_stage_opamp_dummy_magic_0.VOUT-.t127 GNDA 0.290811f
C978 two_stage_opamp_dummy_magic_0.VOUT-.t34 GNDA 0.295144f
C979 two_stage_opamp_dummy_magic_0.VOUT-.t86 GNDA 0.295144f
C980 two_stage_opamp_dummy_magic_0.VOUT-.t42 GNDA 0.295144f
C981 two_stage_opamp_dummy_magic_0.VOUT-.t96 GNDA 0.295144f
C982 two_stage_opamp_dummy_magic_0.VOUT-.t143 GNDA 0.295144f
C983 two_stage_opamp_dummy_magic_0.VOUT-.t106 GNDA 0.295144f
C984 two_stage_opamp_dummy_magic_0.VOUT-.t154 GNDA 0.295144f
C985 two_stage_opamp_dummy_magic_0.VOUT-.t64 GNDA 0.295144f
C986 two_stage_opamp_dummy_magic_0.VOUT-.t116 GNDA 0.295144f
C987 two_stage_opamp_dummy_magic_0.VOUT-.t73 GNDA 0.295144f
C988 two_stage_opamp_dummy_magic_0.VOUT-.t149 GNDA 0.290811f
C989 two_stage_opamp_dummy_magic_0.VOUT-.n14 GNDA 0.195599f
C990 two_stage_opamp_dummy_magic_0.VOUT-.t58 GNDA 0.290811f
C991 two_stage_opamp_dummy_magic_0.VOUT-.n15 GNDA 0.250126f
C992 two_stage_opamp_dummy_magic_0.VOUT-.t97 GNDA 0.290811f
C993 two_stage_opamp_dummy_magic_0.VOUT-.n16 GNDA 0.250126f
C994 two_stage_opamp_dummy_magic_0.VOUT-.t131 GNDA 0.290811f
C995 two_stage_opamp_dummy_magic_0.VOUT-.n17 GNDA 0.250126f
C996 two_stage_opamp_dummy_magic_0.VOUT-.t24 GNDA 0.290811f
C997 two_stage_opamp_dummy_magic_0.VOUT-.n18 GNDA 0.250126f
C998 two_stage_opamp_dummy_magic_0.VOUT-.t75 GNDA 0.290811f
C999 two_stage_opamp_dummy_magic_0.VOUT-.n19 GNDA 0.250126f
C1000 two_stage_opamp_dummy_magic_0.VOUT-.t113 GNDA 0.290811f
C1001 two_stage_opamp_dummy_magic_0.VOUT-.n20 GNDA 0.250126f
C1002 two_stage_opamp_dummy_magic_0.VOUT-.t144 GNDA 0.290811f
C1003 two_stage_opamp_dummy_magic_0.VOUT-.n21 GNDA 0.250126f
C1004 two_stage_opamp_dummy_magic_0.VOUT-.t54 GNDA 0.290811f
C1005 two_stage_opamp_dummy_magic_0.VOUT-.n22 GNDA 0.250126f
C1006 two_stage_opamp_dummy_magic_0.VOUT-.t94 GNDA 0.290811f
C1007 two_stage_opamp_dummy_magic_0.VOUT-.n23 GNDA 0.250126f
C1008 two_stage_opamp_dummy_magic_0.VOUT-.n24 GNDA 0.236284f
C1009 two_stage_opamp_dummy_magic_0.VOUT-.t37 GNDA 0.295764f
C1010 two_stage_opamp_dummy_magic_0.VOUT-.t142 GNDA 0.290811f
C1011 two_stage_opamp_dummy_magic_0.VOUT-.n25 GNDA 0.194979f
C1012 two_stage_opamp_dummy_magic_0.VOUT-.t93 GNDA 0.290811f
C1013 two_stage_opamp_dummy_magic_0.VOUT-.t20 GNDA 0.295764f
C1014 two_stage_opamp_dummy_magic_0.VOUT-.t57 GNDA 0.290811f
C1015 two_stage_opamp_dummy_magic_0.VOUT-.n26 GNDA 0.194979f
C1016 two_stage_opamp_dummy_magic_0.VOUT-.n27 GNDA 0.236284f
C1017 two_stage_opamp_dummy_magic_0.VOUT-.t79 GNDA 0.295764f
C1018 two_stage_opamp_dummy_magic_0.VOUT-.t41 GNDA 0.290811f
C1019 two_stage_opamp_dummy_magic_0.VOUT-.n28 GNDA 0.194979f
C1020 two_stage_opamp_dummy_magic_0.VOUT-.t133 GNDA 0.290811f
C1021 two_stage_opamp_dummy_magic_0.VOUT-.t60 GNDA 0.295764f
C1022 two_stage_opamp_dummy_magic_0.VOUT-.t100 GNDA 0.290811f
C1023 two_stage_opamp_dummy_magic_0.VOUT-.n29 GNDA 0.194979f
C1024 two_stage_opamp_dummy_magic_0.VOUT-.n30 GNDA 0.236284f
C1025 two_stage_opamp_dummy_magic_0.VOUT-.t121 GNDA 0.295764f
C1026 two_stage_opamp_dummy_magic_0.VOUT-.t83 GNDA 0.290811f
C1027 two_stage_opamp_dummy_magic_0.VOUT-.n31 GNDA 0.194979f
C1028 two_stage_opamp_dummy_magic_0.VOUT-.t31 GNDA 0.290811f
C1029 two_stage_opamp_dummy_magic_0.VOUT-.t104 GNDA 0.295764f
C1030 two_stage_opamp_dummy_magic_0.VOUT-.t137 GNDA 0.290811f
C1031 two_stage_opamp_dummy_magic_0.VOUT-.n32 GNDA 0.194979f
C1032 two_stage_opamp_dummy_magic_0.VOUT-.n33 GNDA 0.236284f
C1033 two_stage_opamp_dummy_magic_0.VOUT-.t84 GNDA 0.295764f
C1034 two_stage_opamp_dummy_magic_0.VOUT-.t49 GNDA 0.290811f
C1035 two_stage_opamp_dummy_magic_0.VOUT-.n34 GNDA 0.194979f
C1036 two_stage_opamp_dummy_magic_0.VOUT-.t138 GNDA 0.290811f
C1037 two_stage_opamp_dummy_magic_0.VOUT-.t66 GNDA 0.295764f
C1038 two_stage_opamp_dummy_magic_0.VOUT-.t103 GNDA 0.290811f
C1039 two_stage_opamp_dummy_magic_0.VOUT-.n35 GNDA 0.194979f
C1040 two_stage_opamp_dummy_magic_0.VOUT-.n36 GNDA 0.236284f
C1041 two_stage_opamp_dummy_magic_0.VOUT-.t108 GNDA 0.295764f
C1042 two_stage_opamp_dummy_magic_0.VOUT-.t69 GNDA 0.290811f
C1043 two_stage_opamp_dummy_magic_0.VOUT-.n37 GNDA 0.194979f
C1044 two_stage_opamp_dummy_magic_0.VOUT-.t90 GNDA 0.290811f
C1045 two_stage_opamp_dummy_magic_0.VOUT-.n38 GNDA 0.12723f
C1046 two_stage_opamp_dummy_magic_0.VOUT-.t67 GNDA 0.295764f
C1047 two_stage_opamp_dummy_magic_0.VOUT-.t30 GNDA 0.290811f
C1048 two_stage_opamp_dummy_magic_0.VOUT-.n39 GNDA 0.194979f
C1049 two_stage_opamp_dummy_magic_0.VOUT-.t51 GNDA 0.290811f
C1050 two_stage_opamp_dummy_magic_0.VOUT-.t53 GNDA 0.295144f
C1051 two_stage_opamp_dummy_magic_0.VOUT-.t156 GNDA 0.295144f
C1052 two_stage_opamp_dummy_magic_0.VOUT-.t44 GNDA 0.295764f
C1053 two_stage_opamp_dummy_magic_0.VOUT-.t136 GNDA 0.290811f
C1054 two_stage_opamp_dummy_magic_0.VOUT-.n40 GNDA 0.194979f
C1055 two_stage_opamp_dummy_magic_0.VOUT-.t101 GNDA 0.290811f
C1056 two_stage_opamp_dummy_magic_0.VOUT-.n41 GNDA 0.122686f
C1057 two_stage_opamp_dummy_magic_0.VOUT-.t36 GNDA 0.295144f
C1058 two_stage_opamp_dummy_magic_0.VOUT-.t151 GNDA 0.295764f
C1059 two_stage_opamp_dummy_magic_0.VOUT-.t98 GNDA 0.290811f
C1060 two_stage_opamp_dummy_magic_0.VOUT-.n42 GNDA 0.194979f
C1061 two_stage_opamp_dummy_magic_0.VOUT-.t59 GNDA 0.290811f
C1062 two_stage_opamp_dummy_magic_0.VOUT-.n43 GNDA 0.122686f
C1063 two_stage_opamp_dummy_magic_0.VOUT-.t140 GNDA 0.295144f
C1064 two_stage_opamp_dummy_magic_0.VOUT-.t118 GNDA 0.295764f
C1065 two_stage_opamp_dummy_magic_0.VOUT-.t56 GNDA 0.290811f
C1066 two_stage_opamp_dummy_magic_0.VOUT-.n44 GNDA 0.194979f
C1067 two_stage_opamp_dummy_magic_0.VOUT-.t21 GNDA 0.290811f
C1068 two_stage_opamp_dummy_magic_0.VOUT-.n45 GNDA 0.122686f
C1069 two_stage_opamp_dummy_magic_0.VOUT-.t105 GNDA 0.295144f
C1070 two_stage_opamp_dummy_magic_0.VOUT-.t65 GNDA 0.295764f
C1071 two_stage_opamp_dummy_magic_0.VOUT-.t80 GNDA 0.290811f
C1072 two_stage_opamp_dummy_magic_0.VOUT-.n46 GNDA 0.194979f
C1073 two_stage_opamp_dummy_magic_0.VOUT-.t43 GNDA 0.290811f
C1074 two_stage_opamp_dummy_magic_0.VOUT-.n47 GNDA 0.122686f
C1075 two_stage_opamp_dummy_magic_0.VOUT-.t125 GNDA 0.295144f
C1076 two_stage_opamp_dummy_magic_0.VOUT-.t145 GNDA 0.295387f
C1077 two_stage_opamp_dummy_magic_0.VOUT-.t87 GNDA 0.295144f
C1078 two_stage_opamp_dummy_magic_0.VOUT-.t110 GNDA 0.295387f
C1079 two_stage_opamp_dummy_magic_0.VOUT-.t50 GNDA 0.295144f
C1080 two_stage_opamp_dummy_magic_0.VOUT-.t70 GNDA 0.295387f
C1081 two_stage_opamp_dummy_magic_0.VOUT-.t150 GNDA 0.295144f
C1082 two_stage_opamp_dummy_magic_0.VOUT-.t95 GNDA 0.295387f
C1083 two_stage_opamp_dummy_magic_0.VOUT-.t32 GNDA 0.295144f
C1084 two_stage_opamp_dummy_magic_0.VOUT-.t134 GNDA 0.290811f
C1085 two_stage_opamp_dummy_magic_0.VOUT-.n48 GNDA 0.321888f
C1086 two_stage_opamp_dummy_magic_0.VOUT-.t111 GNDA 0.290811f
C1087 two_stage_opamp_dummy_magic_0.VOUT-.n49 GNDA 0.376415f
C1088 two_stage_opamp_dummy_magic_0.VOUT-.t147 GNDA 0.290811f
C1089 two_stage_opamp_dummy_magic_0.VOUT-.n50 GNDA 0.376415f
C1090 two_stage_opamp_dummy_magic_0.VOUT-.t45 GNDA 0.290811f
C1091 two_stage_opamp_dummy_magic_0.VOUT-.n51 GNDA 0.376415f
C1092 two_stage_opamp_dummy_magic_0.VOUT-.t85 GNDA 0.290811f
C1093 two_stage_opamp_dummy_magic_0.VOUT-.n52 GNDA 0.309197f
C1094 two_stage_opamp_dummy_magic_0.VOUT-.t61 GNDA 0.290811f
C1095 two_stage_opamp_dummy_magic_0.VOUT-.n53 GNDA 0.309197f
C1096 two_stage_opamp_dummy_magic_0.VOUT-.t102 GNDA 0.290811f
C1097 two_stage_opamp_dummy_magic_0.VOUT-.n54 GNDA 0.309197f
C1098 two_stage_opamp_dummy_magic_0.VOUT-.t139 GNDA 0.290811f
C1099 two_stage_opamp_dummy_magic_0.VOUT-.n55 GNDA 0.309197f
C1100 two_stage_opamp_dummy_magic_0.VOUT-.t119 GNDA 0.290811f
C1101 two_stage_opamp_dummy_magic_0.VOUT-.n56 GNDA 0.250126f
C1102 two_stage_opamp_dummy_magic_0.VOUT-.t155 GNDA 0.290811f
C1103 two_stage_opamp_dummy_magic_0.VOUT-.n57 GNDA 0.250126f
C1104 two_stage_opamp_dummy_magic_0.VOUT-.n58 GNDA 0.236284f
C1105 two_stage_opamp_dummy_magic_0.VOUT-.t27 GNDA 0.295764f
C1106 two_stage_opamp_dummy_magic_0.VOUT-.t130 GNDA 0.290811f
C1107 two_stage_opamp_dummy_magic_0.VOUT-.n59 GNDA 0.194979f
C1108 two_stage_opamp_dummy_magic_0.VOUT-.t152 GNDA 0.290811f
C1109 two_stage_opamp_dummy_magic_0.VOUT-.t76 GNDA 0.295764f
C1110 two_stage_opamp_dummy_magic_0.VOUT-.t115 GNDA 0.290811f
C1111 two_stage_opamp_dummy_magic_0.VOUT-.n60 GNDA 0.194979f
C1112 two_stage_opamp_dummy_magic_0.VOUT-.n61 GNDA 0.236284f
C1113 two_stage_opamp_dummy_magic_0.VOUT-.t62 GNDA 0.295764f
C1114 two_stage_opamp_dummy_magic_0.VOUT-.t23 GNDA 0.290811f
C1115 two_stage_opamp_dummy_magic_0.VOUT-.n62 GNDA 0.194979f
C1116 two_stage_opamp_dummy_magic_0.VOUT-.t47 GNDA 0.290811f
C1117 two_stage_opamp_dummy_magic_0.VOUT-.t112 GNDA 0.295764f
C1118 two_stage_opamp_dummy_magic_0.VOUT-.t148 GNDA 0.290811f
C1119 two_stage_opamp_dummy_magic_0.VOUT-.n63 GNDA 0.194979f
C1120 two_stage_opamp_dummy_magic_0.VOUT-.n64 GNDA 0.236284f
C1121 two_stage_opamp_dummy_magic_0.VOUT-.t114 GNDA 0.295764f
C1122 two_stage_opamp_dummy_magic_0.VOUT-.t78 GNDA 0.290811f
C1123 two_stage_opamp_dummy_magic_0.VOUT-.n65 GNDA 0.194979f
C1124 two_stage_opamp_dummy_magic_0.VOUT-.t26 GNDA 0.290811f
C1125 two_stage_opamp_dummy_magic_0.VOUT-.t99 GNDA 0.295764f
C1126 two_stage_opamp_dummy_magic_0.VOUT-.t132 GNDA 0.290811f
C1127 two_stage_opamp_dummy_magic_0.VOUT-.n66 GNDA 0.194979f
C1128 two_stage_opamp_dummy_magic_0.VOUT-.n67 GNDA 0.236284f
C1129 two_stage_opamp_dummy_magic_0.VOUT-.t74 GNDA 0.295764f
C1130 two_stage_opamp_dummy_magic_0.VOUT-.t39 GNDA 0.290811f
C1131 two_stage_opamp_dummy_magic_0.VOUT-.n68 GNDA 0.194979f
C1132 two_stage_opamp_dummy_magic_0.VOUT-.t128 GNDA 0.290811f
C1133 two_stage_opamp_dummy_magic_0.VOUT-.t55 GNDA 0.295764f
C1134 two_stage_opamp_dummy_magic_0.VOUT-.t92 GNDA 0.290811f
C1135 two_stage_opamp_dummy_magic_0.VOUT-.n69 GNDA 0.194979f
C1136 two_stage_opamp_dummy_magic_0.VOUT-.n70 GNDA 0.236284f
C1137 two_stage_opamp_dummy_magic_0.VOUT-.t109 GNDA 0.295764f
C1138 two_stage_opamp_dummy_magic_0.VOUT-.t71 GNDA 0.290811f
C1139 two_stage_opamp_dummy_magic_0.VOUT-.n71 GNDA 0.194979f
C1140 two_stage_opamp_dummy_magic_0.VOUT-.t19 GNDA 0.290811f
C1141 two_stage_opamp_dummy_magic_0.VOUT-.t91 GNDA 0.295764f
C1142 two_stage_opamp_dummy_magic_0.VOUT-.t126 GNDA 0.290811f
C1143 two_stage_opamp_dummy_magic_0.VOUT-.n72 GNDA 0.194979f
C1144 two_stage_opamp_dummy_magic_0.VOUT-.n73 GNDA 0.236284f
C1145 two_stage_opamp_dummy_magic_0.VOUT-.t68 GNDA 0.295764f
C1146 two_stage_opamp_dummy_magic_0.VOUT-.t33 GNDA 0.290811f
C1147 two_stage_opamp_dummy_magic_0.VOUT-.n74 GNDA 0.194979f
C1148 two_stage_opamp_dummy_magic_0.VOUT-.t122 GNDA 0.290811f
C1149 two_stage_opamp_dummy_magic_0.VOUT-.t52 GNDA 0.295764f
C1150 two_stage_opamp_dummy_magic_0.VOUT-.t88 GNDA 0.290811f
C1151 two_stage_opamp_dummy_magic_0.VOUT-.n75 GNDA 0.194979f
C1152 two_stage_opamp_dummy_magic_0.VOUT-.n76 GNDA 0.236284f
C1153 two_stage_opamp_dummy_magic_0.VOUT-.t29 GNDA 0.295764f
C1154 two_stage_opamp_dummy_magic_0.VOUT-.t135 GNDA 0.290811f
C1155 two_stage_opamp_dummy_magic_0.VOUT-.n77 GNDA 0.194979f
C1156 two_stage_opamp_dummy_magic_0.VOUT-.t82 GNDA 0.290811f
C1157 two_stage_opamp_dummy_magic_0.VOUT-.t153 GNDA 0.295764f
C1158 two_stage_opamp_dummy_magic_0.VOUT-.t48 GNDA 0.290811f
C1159 two_stage_opamp_dummy_magic_0.VOUT-.n78 GNDA 0.194979f
C1160 two_stage_opamp_dummy_magic_0.VOUT-.n79 GNDA 0.236284f
C1161 two_stage_opamp_dummy_magic_0.VOUT-.t63 GNDA 0.295764f
C1162 two_stage_opamp_dummy_magic_0.VOUT-.t28 GNDA 0.290811f
C1163 two_stage_opamp_dummy_magic_0.VOUT-.n80 GNDA 0.194979f
C1164 two_stage_opamp_dummy_magic_0.VOUT-.t120 GNDA 0.290811f
C1165 two_stage_opamp_dummy_magic_0.VOUT-.t46 GNDA 0.295764f
C1166 two_stage_opamp_dummy_magic_0.VOUT-.t81 GNDA 0.290811f
C1167 two_stage_opamp_dummy_magic_0.VOUT-.n81 GNDA 0.194979f
C1168 two_stage_opamp_dummy_magic_0.VOUT-.n82 GNDA 0.236284f
C1169 two_stage_opamp_dummy_magic_0.VOUT-.t22 GNDA 0.295764f
C1170 two_stage_opamp_dummy_magic_0.VOUT-.t129 GNDA 0.290811f
C1171 two_stage_opamp_dummy_magic_0.VOUT-.n83 GNDA 0.194979f
C1172 two_stage_opamp_dummy_magic_0.VOUT-.t77 GNDA 0.290811f
C1173 two_stage_opamp_dummy_magic_0.VOUT-.t146 GNDA 0.295764f
C1174 two_stage_opamp_dummy_magic_0.VOUT-.t40 GNDA 0.290811f
C1175 two_stage_opamp_dummy_magic_0.VOUT-.n84 GNDA 0.194979f
C1176 two_stage_opamp_dummy_magic_0.VOUT-.n85 GNDA 0.236284f
C1177 two_stage_opamp_dummy_magic_0.VOUT-.t123 GNDA 0.295764f
C1178 two_stage_opamp_dummy_magic_0.VOUT-.t89 GNDA 0.290811f
C1179 two_stage_opamp_dummy_magic_0.VOUT-.n86 GNDA 0.194979f
C1180 two_stage_opamp_dummy_magic_0.VOUT-.t35 GNDA 0.290811f
C1181 two_stage_opamp_dummy_magic_0.VOUT-.n87 GNDA 0.236284f
C1182 two_stage_opamp_dummy_magic_0.VOUT-.t141 GNDA 0.290811f
C1183 two_stage_opamp_dummy_magic_0.VOUT-.n88 GNDA 0.12723f
C1184 two_stage_opamp_dummy_magic_0.VOUT-.t107 GNDA 0.290811f
C1185 two_stage_opamp_dummy_magic_0.VOUT-.n89 GNDA 0.23826f
C1186 two_stage_opamp_dummy_magic_0.VOUT-.n90 GNDA 0.300935f
C1187 two_stage_opamp_dummy_magic_0.VOUT-.t1 GNDA 0.050892f
C1188 two_stage_opamp_dummy_magic_0.VOUT-.t18 GNDA 0.050892f
C1189 two_stage_opamp_dummy_magic_0.VOUT-.n91 GNDA 0.235428f
C1190 two_stage_opamp_dummy_magic_0.VOUT-.t3 GNDA 0.050892f
C1191 two_stage_opamp_dummy_magic_0.VOUT-.t2 GNDA 0.050892f
C1192 two_stage_opamp_dummy_magic_0.VOUT-.n92 GNDA 0.23464f
C1193 two_stage_opamp_dummy_magic_0.VOUT-.n93 GNDA 0.144996f
C1194 two_stage_opamp_dummy_magic_0.VOUT-.t17 GNDA 0.050892f
C1195 two_stage_opamp_dummy_magic_0.VOUT-.t14 GNDA 0.050892f
C1196 two_stage_opamp_dummy_magic_0.VOUT-.n94 GNDA 0.23464f
C1197 two_stage_opamp_dummy_magic_0.VOUT-.n95 GNDA 0.08925f
C1198 two_stage_opamp_dummy_magic_0.VOUT-.n96 GNDA 0.170241f
C1199 two_stage_opamp_dummy_magic_0.VOUT-.t0 GNDA 0.084142f
C1200 two_stage_opamp_dummy_magic_0.X.t17 GNDA 0.024316f
C1201 two_stage_opamp_dummy_magic_0.X.t14 GNDA 0.024316f
C1202 two_stage_opamp_dummy_magic_0.X.n0 GNDA 0.082095f
C1203 two_stage_opamp_dummy_magic_0.X.t20 GNDA 0.024316f
C1204 two_stage_opamp_dummy_magic_0.X.t22 GNDA 0.024316f
C1205 two_stage_opamp_dummy_magic_0.X.n1 GNDA 0.087741f
C1206 two_stage_opamp_dummy_magic_0.X.t21 GNDA 0.024316f
C1207 two_stage_opamp_dummy_magic_0.X.t19 GNDA 0.024316f
C1208 two_stage_opamp_dummy_magic_0.X.n2 GNDA 0.087741f
C1209 two_stage_opamp_dummy_magic_0.X.t16 GNDA 0.024316f
C1210 two_stage_opamp_dummy_magic_0.X.t23 GNDA 0.024316f
C1211 two_stage_opamp_dummy_magic_0.X.n3 GNDA 0.086975f
C1212 two_stage_opamp_dummy_magic_0.X.n4 GNDA 0.32294f
C1213 two_stage_opamp_dummy_magic_0.X.t10 GNDA 0.024316f
C1214 two_stage_opamp_dummy_magic_0.X.t13 GNDA 0.024316f
C1215 two_stage_opamp_dummy_magic_0.X.n5 GNDA 0.086975f
C1216 two_stage_opamp_dummy_magic_0.X.n6 GNDA 0.167527f
C1217 two_stage_opamp_dummy_magic_0.X.t15 GNDA 0.024316f
C1218 two_stage_opamp_dummy_magic_0.X.t11 GNDA 0.024316f
C1219 two_stage_opamp_dummy_magic_0.X.n7 GNDA 0.086975f
C1220 two_stage_opamp_dummy_magic_0.X.n8 GNDA 0.167527f
C1221 two_stage_opamp_dummy_magic_0.X.n9 GNDA 0.204045f
C1222 two_stage_opamp_dummy_magic_0.X.n10 GNDA 0.164936f
C1223 two_stage_opamp_dummy_magic_0.X.t12 GNDA 0.79195f
C1224 two_stage_opamp_dummy_magic_0.X.t36 GNDA 0.106988f
C1225 two_stage_opamp_dummy_magic_0.X.t49 GNDA 0.106988f
C1226 two_stage_opamp_dummy_magic_0.X.t34 GNDA 0.11395f
C1227 two_stage_opamp_dummy_magic_0.X.n11 GNDA 0.0903f
C1228 two_stage_opamp_dummy_magic_0.X.n12 GNDA 0.048273f
C1229 two_stage_opamp_dummy_magic_0.X.t51 GNDA 0.106988f
C1230 two_stage_opamp_dummy_magic_0.X.t39 GNDA 0.106988f
C1231 two_stage_opamp_dummy_magic_0.X.t26 GNDA 0.106988f
C1232 two_stage_opamp_dummy_magic_0.X.t44 GNDA 0.106988f
C1233 two_stage_opamp_dummy_magic_0.X.t25 GNDA 0.106988f
C1234 two_stage_opamp_dummy_magic_0.X.t43 GNDA 0.106988f
C1235 two_stage_opamp_dummy_magic_0.X.t29 GNDA 0.11395f
C1236 two_stage_opamp_dummy_magic_0.X.n13 GNDA 0.0903f
C1237 two_stage_opamp_dummy_magic_0.X.n14 GNDA 0.051063f
C1238 two_stage_opamp_dummy_magic_0.X.n15 GNDA 0.051063f
C1239 two_stage_opamp_dummy_magic_0.X.n16 GNDA 0.051063f
C1240 two_stage_opamp_dummy_magic_0.X.n17 GNDA 0.051063f
C1241 two_stage_opamp_dummy_magic_0.X.n18 GNDA 0.048273f
C1242 two_stage_opamp_dummy_magic_0.X.n19 GNDA 0.026157f
C1243 two_stage_opamp_dummy_magic_0.X.n20 GNDA 0.942239f
C1244 two_stage_opamp_dummy_magic_0.X.t6 GNDA 0.056736f
C1245 two_stage_opamp_dummy_magic_0.X.t24 GNDA 0.056736f
C1246 two_stage_opamp_dummy_magic_0.X.n21 GNDA 0.197316f
C1247 two_stage_opamp_dummy_magic_0.X.t8 GNDA 0.056736f
C1248 two_stage_opamp_dummy_magic_0.X.t9 GNDA 0.056736f
C1249 two_stage_opamp_dummy_magic_0.X.n22 GNDA 0.196617f
C1250 two_stage_opamp_dummy_magic_0.X.n23 GNDA 0.371194f
C1251 two_stage_opamp_dummy_magic_0.X.t3 GNDA 0.056736f
C1252 two_stage_opamp_dummy_magic_0.X.t2 GNDA 0.056736f
C1253 two_stage_opamp_dummy_magic_0.X.n24 GNDA 0.196617f
C1254 two_stage_opamp_dummy_magic_0.X.n25 GNDA 0.19243f
C1255 two_stage_opamp_dummy_magic_0.X.t5 GNDA 0.056736f
C1256 two_stage_opamp_dummy_magic_0.X.t4 GNDA 0.056736f
C1257 two_stage_opamp_dummy_magic_0.X.n26 GNDA 0.196617f
C1258 two_stage_opamp_dummy_magic_0.X.n27 GNDA 0.19243f
C1259 two_stage_opamp_dummy_magic_0.X.t0 GNDA 0.056736f
C1260 two_stage_opamp_dummy_magic_0.X.t7 GNDA 0.056736f
C1261 two_stage_opamp_dummy_magic_0.X.n28 GNDA 0.196617f
C1262 two_stage_opamp_dummy_magic_0.X.n29 GNDA 0.226591f
C1263 two_stage_opamp_dummy_magic_0.X.t18 GNDA 0.056736f
C1264 two_stage_opamp_dummy_magic_0.X.t1 GNDA 0.056736f
C1265 two_stage_opamp_dummy_magic_0.X.n30 GNDA 0.192544f
C1266 two_stage_opamp_dummy_magic_0.X.n31 GNDA 0.383218f
C1267 two_stage_opamp_dummy_magic_0.X.t53 GNDA 0.034042f
C1268 two_stage_opamp_dummy_magic_0.X.t42 GNDA 0.034042f
C1269 two_stage_opamp_dummy_magic_0.X.t54 GNDA 0.034042f
C1270 two_stage_opamp_dummy_magic_0.X.t38 GNDA 0.034042f
C1271 two_stage_opamp_dummy_magic_0.X.t50 GNDA 0.034042f
C1272 two_stage_opamp_dummy_magic_0.X.t35 GNDA 0.034042f
C1273 two_stage_opamp_dummy_magic_0.X.t48 GNDA 0.034042f
C1274 two_stage_opamp_dummy_magic_0.X.t33 GNDA 0.041336f
C1275 two_stage_opamp_dummy_magic_0.X.n32 GNDA 0.041336f
C1276 two_stage_opamp_dummy_magic_0.X.n33 GNDA 0.026747f
C1277 two_stage_opamp_dummy_magic_0.X.n34 GNDA 0.026747f
C1278 two_stage_opamp_dummy_magic_0.X.n35 GNDA 0.026747f
C1279 two_stage_opamp_dummy_magic_0.X.n36 GNDA 0.026747f
C1280 two_stage_opamp_dummy_magic_0.X.n37 GNDA 0.026747f
C1281 two_stage_opamp_dummy_magic_0.X.n38 GNDA 0.023958f
C1282 two_stage_opamp_dummy_magic_0.X.t41 GNDA 0.034042f
C1283 two_stage_opamp_dummy_magic_0.X.t28 GNDA 0.041336f
C1284 two_stage_opamp_dummy_magic_0.X.n39 GNDA 0.038547f
C1285 two_stage_opamp_dummy_magic_0.X.n40 GNDA 0.023563f
C1286 two_stage_opamp_dummy_magic_0.X.t30 GNDA 0.052278f
C1287 two_stage_opamp_dummy_magic_0.X.t47 GNDA 0.052278f
C1288 two_stage_opamp_dummy_magic_0.X.t31 GNDA 0.052278f
C1289 two_stage_opamp_dummy_magic_0.X.t45 GNDA 0.052278f
C1290 two_stage_opamp_dummy_magic_0.X.t27 GNDA 0.052278f
C1291 two_stage_opamp_dummy_magic_0.X.t40 GNDA 0.052278f
C1292 two_stage_opamp_dummy_magic_0.X.t52 GNDA 0.052278f
C1293 two_stage_opamp_dummy_magic_0.X.t37 GNDA 0.059432f
C1294 two_stage_opamp_dummy_magic_0.X.n41 GNDA 0.053635f
C1295 two_stage_opamp_dummy_magic_0.X.n42 GNDA 0.032826f
C1296 two_stage_opamp_dummy_magic_0.X.n43 GNDA 0.032826f
C1297 two_stage_opamp_dummy_magic_0.X.n44 GNDA 0.032826f
C1298 two_stage_opamp_dummy_magic_0.X.n45 GNDA 0.032826f
C1299 two_stage_opamp_dummy_magic_0.X.n46 GNDA 0.032826f
C1300 two_stage_opamp_dummy_magic_0.X.n47 GNDA 0.030036f
C1301 two_stage_opamp_dummy_magic_0.X.t46 GNDA 0.052278f
C1302 two_stage_opamp_dummy_magic_0.X.t32 GNDA 0.059432f
C1303 two_stage_opamp_dummy_magic_0.X.n48 GNDA 0.050846f
C1304 two_stage_opamp_dummy_magic_0.X.n49 GNDA 0.023513f
C1305 two_stage_opamp_dummy_magic_0.X.n50 GNDA 0.25433f
C1306 two_stage_opamp_dummy_magic_0.X.n51 GNDA 0.527634f
C1307 two_stage_opamp_dummy_magic_0.X.n52 GNDA 0.245911f
C1308 two_stage_opamp_dummy_magic_0.X.n53 GNDA 0.104409f
C1309 two_stage_opamp_dummy_magic_0.VD4.t10 GNDA 0.026025f
C1310 two_stage_opamp_dummy_magic_0.VD4.t14 GNDA 0.026025f
C1311 two_stage_opamp_dummy_magic_0.VD4.n0 GNDA 0.090508f
C1312 two_stage_opamp_dummy_magic_0.VD4.t18 GNDA 0.026025f
C1313 two_stage_opamp_dummy_magic_0.VD4.t2 GNDA 0.026025f
C1314 two_stage_opamp_dummy_magic_0.VD4.n1 GNDA 0.090188f
C1315 two_stage_opamp_dummy_magic_0.VD4.n2 GNDA 0.170266f
C1316 two_stage_opamp_dummy_magic_0.VD4.n3 GNDA 0.073371f
C1317 two_stage_opamp_dummy_magic_0.VD4.n4 GNDA 0.100747f
C1318 two_stage_opamp_dummy_magic_0.VD4.t34 GNDA 0.128386f
C1319 two_stage_opamp_dummy_magic_0.VD4.t32 GNDA 0.045318f
C1320 two_stage_opamp_dummy_magic_0.VD4.n5 GNDA 0.083755f
C1321 two_stage_opamp_dummy_magic_0.VD4.n6 GNDA 0.053992f
C1322 two_stage_opamp_dummy_magic_0.VD4.t37 GNDA 0.128386f
C1323 two_stage_opamp_dummy_magic_0.VD4.t35 GNDA 0.045318f
C1324 two_stage_opamp_dummy_magic_0.VD4.n7 GNDA 0.083755f
C1325 two_stage_opamp_dummy_magic_0.VD4.n8 GNDA 0.053992f
C1326 two_stage_opamp_dummy_magic_0.VD4.n9 GNDA 0.053537f
C1327 two_stage_opamp_dummy_magic_0.VD4.n10 GNDA 0.100747f
C1328 two_stage_opamp_dummy_magic_0.VD4.n11 GNDA 0.300245f
C1329 two_stage_opamp_dummy_magic_0.VD4.t36 GNDA 0.448159f
C1330 two_stage_opamp_dummy_magic_0.VD4.t9 GNDA 0.25876f
C1331 two_stage_opamp_dummy_magic_0.VD4.t13 GNDA 0.25876f
C1332 two_stage_opamp_dummy_magic_0.VD4.t17 GNDA 0.25876f
C1333 two_stage_opamp_dummy_magic_0.VD4.t1 GNDA 0.25876f
C1334 two_stage_opamp_dummy_magic_0.VD4.t5 GNDA 0.19407f
C1335 two_stage_opamp_dummy_magic_0.VD4.n12 GNDA 0.12938f
C1336 two_stage_opamp_dummy_magic_0.VD4.t7 GNDA 0.19407f
C1337 two_stage_opamp_dummy_magic_0.VD4.t11 GNDA 0.25876f
C1338 two_stage_opamp_dummy_magic_0.VD4.t15 GNDA 0.25876f
C1339 two_stage_opamp_dummy_magic_0.VD4.t19 GNDA 0.25876f
C1340 two_stage_opamp_dummy_magic_0.VD4.t3 GNDA 0.25876f
C1341 two_stage_opamp_dummy_magic_0.VD4.t33 GNDA 0.448159f
C1342 two_stage_opamp_dummy_magic_0.VD4.n13 GNDA 0.300245f
C1343 two_stage_opamp_dummy_magic_0.VD4.n14 GNDA 0.073371f
C1344 two_stage_opamp_dummy_magic_0.VD4.n15 GNDA 0.108171f
C1345 two_stage_opamp_dummy_magic_0.VD4.t6 GNDA 0.026025f
C1346 two_stage_opamp_dummy_magic_0.VD4.t8 GNDA 0.026025f
C1347 two_stage_opamp_dummy_magic_0.VD4.n16 GNDA 0.08832f
C1348 two_stage_opamp_dummy_magic_0.VD4.n17 GNDA 0.069277f
C1349 two_stage_opamp_dummy_magic_0.VD4.n18 GNDA 0.023794f
C1350 two_stage_opamp_dummy_magic_0.VD4.t12 GNDA 0.026025f
C1351 two_stage_opamp_dummy_magic_0.VD4.t16 GNDA 0.026025f
C1352 two_stage_opamp_dummy_magic_0.VD4.n19 GNDA 0.090188f
C1353 two_stage_opamp_dummy_magic_0.VD4.n20 GNDA 0.088268f
C1354 two_stage_opamp_dummy_magic_0.VD4.t20 GNDA 0.026025f
C1355 two_stage_opamp_dummy_magic_0.VD4.t4 GNDA 0.026025f
C1356 two_stage_opamp_dummy_magic_0.VD4.n21 GNDA 0.090188f
C1357 two_stage_opamp_dummy_magic_0.VD4.n22 GNDA 0.117811f
C1358 two_stage_opamp_dummy_magic_0.VD4.t25 GNDA 0.026025f
C1359 two_stage_opamp_dummy_magic_0.VD4.t30 GNDA 0.026025f
C1360 two_stage_opamp_dummy_magic_0.VD4.n23 GNDA 0.090509f
C1361 two_stage_opamp_dummy_magic_0.VD4.t23 GNDA 0.026025f
C1362 two_stage_opamp_dummy_magic_0.VD4.t22 GNDA 0.026025f
C1363 two_stage_opamp_dummy_magic_0.VD4.n24 GNDA 0.090188f
C1364 two_stage_opamp_dummy_magic_0.VD4.n25 GNDA 0.170266f
C1365 two_stage_opamp_dummy_magic_0.VD4.t31 GNDA 0.026025f
C1366 two_stage_opamp_dummy_magic_0.VD4.t24 GNDA 0.026025f
C1367 two_stage_opamp_dummy_magic_0.VD4.n26 GNDA 0.090188f
C1368 two_stage_opamp_dummy_magic_0.VD4.n27 GNDA 0.088268f
C1369 two_stage_opamp_dummy_magic_0.VD4.t21 GNDA 0.026025f
C1370 two_stage_opamp_dummy_magic_0.VD4.t28 GNDA 0.026025f
C1371 two_stage_opamp_dummy_magic_0.VD4.n28 GNDA 0.090188f
C1372 two_stage_opamp_dummy_magic_0.VD4.n29 GNDA 0.088268f
C1373 two_stage_opamp_dummy_magic_0.VD4.t0 GNDA 0.026025f
C1374 two_stage_opamp_dummy_magic_0.VD4.t26 GNDA 0.026025f
C1375 two_stage_opamp_dummy_magic_0.VD4.n30 GNDA 0.090188f
C1376 two_stage_opamp_dummy_magic_0.VD4.n31 GNDA 0.088268f
C1377 two_stage_opamp_dummy_magic_0.VD4.t29 GNDA 0.026025f
C1378 two_stage_opamp_dummy_magic_0.VD4.t27 GNDA 0.026025f
C1379 two_stage_opamp_dummy_magic_0.VD4.n32 GNDA 0.090188f
C1380 two_stage_opamp_dummy_magic_0.VD4.n33 GNDA 0.133786f
C1381 two_stage_opamp_dummy_magic_0.Vb2.t8 GNDA 0.013856f
C1382 two_stage_opamp_dummy_magic_0.Vb2.t1 GNDA 0.013856f
C1383 two_stage_opamp_dummy_magic_0.Vb2.n0 GNDA 0.030075f
C1384 two_stage_opamp_dummy_magic_0.Vb2.t0 GNDA 0.043031f
C1385 two_stage_opamp_dummy_magic_0.Vb2.n1 GNDA 0.185079f
C1386 two_stage_opamp_dummy_magic_0.Vb2.t20 GNDA 0.108864f
C1387 two_stage_opamp_dummy_magic_0.Vb2.t23 GNDA 0.108864f
C1388 two_stage_opamp_dummy_magic_0.Vb2.t21 GNDA 0.108864f
C1389 two_stage_opamp_dummy_magic_0.Vb2.t26 GNDA 0.108864f
C1390 two_stage_opamp_dummy_magic_0.Vb2.t31 GNDA 0.125629f
C1391 two_stage_opamp_dummy_magic_0.Vb2.n2 GNDA 0.101997f
C1392 two_stage_opamp_dummy_magic_0.Vb2.n3 GNDA 0.062679f
C1393 two_stage_opamp_dummy_magic_0.Vb2.n4 GNDA 0.062679f
C1394 two_stage_opamp_dummy_magic_0.Vb2.n5 GNDA 0.058691f
C1395 two_stage_opamp_dummy_magic_0.Vb2.t17 GNDA 0.108864f
C1396 two_stage_opamp_dummy_magic_0.Vb2.t30 GNDA 0.108864f
C1397 two_stage_opamp_dummy_magic_0.Vb2.t25 GNDA 0.108864f
C1398 two_stage_opamp_dummy_magic_0.Vb2.t27 GNDA 0.108864f
C1399 two_stage_opamp_dummy_magic_0.Vb2.t22 GNDA 0.125629f
C1400 two_stage_opamp_dummy_magic_0.Vb2.n6 GNDA 0.101997f
C1401 two_stage_opamp_dummy_magic_0.Vb2.n7 GNDA 0.062679f
C1402 two_stage_opamp_dummy_magic_0.Vb2.n8 GNDA 0.062679f
C1403 two_stage_opamp_dummy_magic_0.Vb2.n9 GNDA 0.058691f
C1404 two_stage_opamp_dummy_magic_0.Vb2.n10 GNDA 0.039642f
C1405 two_stage_opamp_dummy_magic_0.Vb2.t24 GNDA 0.108864f
C1406 two_stage_opamp_dummy_magic_0.Vb2.t29 GNDA 0.108864f
C1407 two_stage_opamp_dummy_magic_0.Vb2.t12 GNDA 0.108864f
C1408 two_stage_opamp_dummy_magic_0.Vb2.t14 GNDA 0.108864f
C1409 two_stage_opamp_dummy_magic_0.Vb2.t16 GNDA 0.125629f
C1410 two_stage_opamp_dummy_magic_0.Vb2.n11 GNDA 0.101997f
C1411 two_stage_opamp_dummy_magic_0.Vb2.n12 GNDA 0.062679f
C1412 two_stage_opamp_dummy_magic_0.Vb2.n13 GNDA 0.062679f
C1413 two_stage_opamp_dummy_magic_0.Vb2.n14 GNDA 0.058691f
C1414 two_stage_opamp_dummy_magic_0.Vb2.t18 GNDA 0.108864f
C1415 two_stage_opamp_dummy_magic_0.Vb2.t15 GNDA 0.108864f
C1416 two_stage_opamp_dummy_magic_0.Vb2.t13 GNDA 0.108864f
C1417 two_stage_opamp_dummy_magic_0.Vb2.t11 GNDA 0.108864f
C1418 two_stage_opamp_dummy_magic_0.Vb2.t28 GNDA 0.125629f
C1419 two_stage_opamp_dummy_magic_0.Vb2.n15 GNDA 0.101997f
C1420 two_stage_opamp_dummy_magic_0.Vb2.n16 GNDA 0.062679f
C1421 two_stage_opamp_dummy_magic_0.Vb2.n17 GNDA 0.062679f
C1422 two_stage_opamp_dummy_magic_0.Vb2.n18 GNDA 0.058691f
C1423 two_stage_opamp_dummy_magic_0.Vb2.n19 GNDA 0.038886f
C1424 two_stage_opamp_dummy_magic_0.Vb2.n20 GNDA 0.883776f
C1425 two_stage_opamp_dummy_magic_0.Vb2.n21 GNDA 0.665732f
C1426 two_stage_opamp_dummy_magic_0.Vb2.t19 GNDA 0.131353f
C1427 two_stage_opamp_dummy_magic_0.Vb2.n22 GNDA 3.33247f
C1428 two_stage_opamp_dummy_magic_0.Vb2.t6 GNDA 0.021993f
C1429 two_stage_opamp_dummy_magic_0.Vb2.t3 GNDA 0.021993f
C1430 two_stage_opamp_dummy_magic_0.Vb2.n23 GNDA 0.066427f
C1431 two_stage_opamp_dummy_magic_0.Vb2.t10 GNDA 0.021993f
C1432 two_stage_opamp_dummy_magic_0.Vb2.t4 GNDA 0.021993f
C1433 two_stage_opamp_dummy_magic_0.Vb2.n24 GNDA 0.070841f
C1434 two_stage_opamp_dummy_magic_0.Vb2.t2 GNDA 0.021993f
C1435 two_stage_opamp_dummy_magic_0.Vb2.t9 GNDA 0.021993f
C1436 two_stage_opamp_dummy_magic_0.Vb2.n25 GNDA 0.070841f
C1437 two_stage_opamp_dummy_magic_0.Vb2.t7 GNDA 0.021993f
C1438 two_stage_opamp_dummy_magic_0.Vb2.t5 GNDA 0.021993f
C1439 two_stage_opamp_dummy_magic_0.Vb2.n26 GNDA 0.070184f
C1440 two_stage_opamp_dummy_magic_0.Vb2.n27 GNDA 0.340616f
C1441 two_stage_opamp_dummy_magic_0.Vb2.n28 GNDA 0.228261f
C1442 two_stage_opamp_dummy_magic_0.Vb2.n29 GNDA 0.163116f
C1443 bgr_0.VB2_CUR_BIAS GNDA 3.14749f
C1444 two_stage_opamp_dummy_magic_0.V_err_gate.n0 GNDA 1.72656f
C1445 two_stage_opamp_dummy_magic_0.V_err_gate.n1 GNDA 8.67705f
C1446 two_stage_opamp_dummy_magic_0.V_err_gate.t1 GNDA 0.02427f
C1447 two_stage_opamp_dummy_magic_0.V_err_gate.t11 GNDA 0.02427f
C1448 two_stage_opamp_dummy_magic_0.V_err_gate.n2 GNDA 0.05665f
C1449 two_stage_opamp_dummy_magic_0.V_err_gate.t5 GNDA 0.02427f
C1450 two_stage_opamp_dummy_magic_0.V_err_gate.t2 GNDA 0.02427f
C1451 two_stage_opamp_dummy_magic_0.V_err_gate.n3 GNDA 0.056284f
C1452 two_stage_opamp_dummy_magic_0.V_err_gate.t13 GNDA 0.02427f
C1453 two_stage_opamp_dummy_magic_0.V_err_gate.t10 GNDA 0.02427f
C1454 two_stage_opamp_dummy_magic_0.V_err_gate.n4 GNDA 0.056284f
C1455 two_stage_opamp_dummy_magic_0.V_err_gate.t23 GNDA 0.020022f
C1456 two_stage_opamp_dummy_magic_0.V_err_gate.t32 GNDA 0.020022f
C1457 two_stage_opamp_dummy_magic_0.V_err_gate.t21 GNDA 0.020022f
C1458 two_stage_opamp_dummy_magic_0.V_err_gate.t30 GNDA 0.020022f
C1459 two_stage_opamp_dummy_magic_0.V_err_gate.t16 GNDA 0.020022f
C1460 two_stage_opamp_dummy_magic_0.V_err_gate.t25 GNDA 0.020022f
C1461 two_stage_opamp_dummy_magic_0.V_err_gate.t18 GNDA 0.020022f
C1462 two_stage_opamp_dummy_magic_0.V_err_gate.t28 GNDA 0.020022f
C1463 two_stage_opamp_dummy_magic_0.V_err_gate.t15 GNDA 0.020022f
C1464 two_stage_opamp_dummy_magic_0.V_err_gate.t24 GNDA 0.020022f
C1465 two_stage_opamp_dummy_magic_0.V_err_gate.t33 GNDA 0.020022f
C1466 two_stage_opamp_dummy_magic_0.V_err_gate.t22 GNDA 0.020022f
C1467 two_stage_opamp_dummy_magic_0.V_err_gate.t31 GNDA 0.020022f
C1468 two_stage_opamp_dummy_magic_0.V_err_gate.t19 GNDA 0.020022f
C1469 two_stage_opamp_dummy_magic_0.V_err_gate.t26 GNDA 0.020022f
C1470 two_stage_opamp_dummy_magic_0.V_err_gate.t20 GNDA 0.020022f
C1471 two_stage_opamp_dummy_magic_0.V_err_gate.t29 GNDA 0.043382f
C1472 two_stage_opamp_dummy_magic_0.V_err_gate.n5 GNDA 0.067652f
C1473 two_stage_opamp_dummy_magic_0.V_err_gate.n6 GNDA 0.052787f
C1474 two_stage_opamp_dummy_magic_0.V_err_gate.n7 GNDA 0.052787f
C1475 two_stage_opamp_dummy_magic_0.V_err_gate.n8 GNDA 0.052787f
C1476 two_stage_opamp_dummy_magic_0.V_err_gate.n9 GNDA 0.052787f
C1477 two_stage_opamp_dummy_magic_0.V_err_gate.n10 GNDA 0.052787f
C1478 two_stage_opamp_dummy_magic_0.V_err_gate.n11 GNDA 0.052787f
C1479 two_stage_opamp_dummy_magic_0.V_err_gate.n12 GNDA 0.052787f
C1480 two_stage_opamp_dummy_magic_0.V_err_gate.n13 GNDA 0.052787f
C1481 two_stage_opamp_dummy_magic_0.V_err_gate.n14 GNDA 0.052787f
C1482 two_stage_opamp_dummy_magic_0.V_err_gate.n15 GNDA 0.052787f
C1483 two_stage_opamp_dummy_magic_0.V_err_gate.n16 GNDA 0.052787f
C1484 two_stage_opamp_dummy_magic_0.V_err_gate.n17 GNDA 0.052787f
C1485 two_stage_opamp_dummy_magic_0.V_err_gate.n18 GNDA 0.052787f
C1486 two_stage_opamp_dummy_magic_0.V_err_gate.n19 GNDA 0.052787f
C1487 two_stage_opamp_dummy_magic_0.V_err_gate.n20 GNDA 0.045171f
C1488 two_stage_opamp_dummy_magic_0.V_err_gate.t14 GNDA 0.020022f
C1489 two_stage_opamp_dummy_magic_0.V_err_gate.t27 GNDA 0.020022f
C1490 two_stage_opamp_dummy_magic_0.V_err_gate.t17 GNDA 0.043382f
C1491 two_stage_opamp_dummy_magic_0.V_err_gate.n21 GNDA 0.067652f
C1492 two_stage_opamp_dummy_magic_0.V_err_gate.n22 GNDA 0.045171f
C1493 two_stage_opamp_dummy_magic_0.V_err_gate.n23 GNDA 0.073284f
C1494 two_stage_opamp_dummy_magic_0.V_err_gate.t4 GNDA 0.02427f
C1495 two_stage_opamp_dummy_magic_0.V_err_gate.t6 GNDA 0.02427f
C1496 two_stage_opamp_dummy_magic_0.V_err_gate.n24 GNDA 0.04854f
C1497 two_stage_opamp_dummy_magic_0.V_err_gate.n25 GNDA 0.144588f
C1498 two_stage_opamp_dummy_magic_0.V_err_gate.t0 GNDA 0.02427f
C1499 two_stage_opamp_dummy_magic_0.V_err_gate.t9 GNDA 0.02427f
C1500 two_stage_opamp_dummy_magic_0.V_err_gate.n26 GNDA 0.056284f
C1501 two_stage_opamp_dummy_magic_0.V_err_gate.t12 GNDA 0.02427f
C1502 two_stage_opamp_dummy_magic_0.V_err_gate.t3 GNDA 0.02427f
C1503 two_stage_opamp_dummy_magic_0.V_err_gate.n27 GNDA 0.055865f
C1504 two_stage_opamp_dummy_magic_0.V_err_gate.t8 GNDA 0.04854f
C1505 two_stage_opamp_dummy_magic_0.V_err_gate.t7 GNDA 0.04854f
C1506 two_stage_opamp_dummy_magic_0.V_err_gate.n28 GNDA 0.149716f
C1507 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t17 GNDA 0.074255f
C1508 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t14 GNDA 0.027767f
C1509 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n0 GNDA 0.087091f
C1510 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t18 GNDA 0.027767f
C1511 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n1 GNDA 0.071293f
C1512 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t13 GNDA 0.027767f
C1513 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n2 GNDA 0.071293f
C1514 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t8 GNDA 0.027767f
C1515 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n3 GNDA 0.109376f
C1516 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t0 GNDA 0.709082f
C1517 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t5 GNDA 0.090054f
C1518 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t2 GNDA 0.090054f
C1519 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n4 GNDA 0.301772f
C1520 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n5 GNDA 3.40029f
C1521 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t4 GNDA 0.090054f
C1522 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t1 GNDA 0.090054f
C1523 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n6 GNDA 0.301772f
C1524 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n7 GNDA 0.814897f
C1525 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t3 GNDA 0.090054f
C1526 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t6 GNDA 0.090054f
C1527 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n8 GNDA 0.301772f
C1528 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n9 GNDA 1.16504f
C1529 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n10 GNDA 1.01344f
C1530 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t9 GNDA 0.043395f
C1531 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t20 GNDA 0.013631f
C1532 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t11 GNDA 0.025436f
C1533 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n11 GNDA 0.060728f
C1534 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n12 GNDA 0.379723f
C1535 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t21 GNDA 0.013631f
C1536 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t15 GNDA 0.025436f
C1537 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n13 GNDA 0.060728f
C1538 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n14 GNDA 0.350774f
C1539 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t16 GNDA 0.042979f
C1540 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n15 GNDA 0.341551f
C1541 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t12 GNDA 0.013631f
C1542 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t7 GNDA 0.025436f
C1543 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n16 GNDA 0.060728f
C1544 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n17 GNDA 0.212091f
C1545 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t10 GNDA 0.013631f
C1546 two_stage_opamp_dummy_magic_0.V_err_amp_ref.t19 GNDA 0.025436f
C1547 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n18 GNDA 0.060728f
C1548 two_stage_opamp_dummy_magic_0.V_err_amp_ref.n19 GNDA 0.269546f
C1549 bgr_0.V_mir2.t0 GNDA 0.042444f
C1550 bgr_0.V_mir2.t18 GNDA 0.042444f
C1551 bgr_0.V_mir2.t20 GNDA 0.06851f
C1552 bgr_0.V_mir2.n0 GNDA 0.076506f
C1553 bgr_0.V_mir2.n1 GNDA 0.052264f
C1554 bgr_0.V_mir2.t4 GNDA 0.053881f
C1555 bgr_0.V_mir2.n2 GNDA 0.081315f
C1556 bgr_0.V_mir2.t1 GNDA 0.03537f
C1557 bgr_0.V_mir2.t5 GNDA 0.03537f
C1558 bgr_0.V_mir2.n3 GNDA 0.08097f
C1559 bgr_0.V_mir2.n4 GNDA 0.201563f
C1560 bgr_0.V_mir2.t15 GNDA 0.017685f
C1561 bgr_0.V_mir2.t16 GNDA 0.017685f
C1562 bgr_0.V_mir2.n5 GNDA 0.046242f
C1563 bgr_0.V_mir2.t13 GNDA 0.075466f
C1564 bgr_0.V_mir2.t14 GNDA 0.017685f
C1565 bgr_0.V_mir2.t12 GNDA 0.017685f
C1566 bgr_0.V_mir2.n6 GNDA 0.050199f
C1567 bgr_0.V_mir2.n7 GNDA 0.827814f
C1568 bgr_0.V_mir2.n8 GNDA 0.268286f
C1569 bgr_0.V_mir2.t8 GNDA 0.042444f
C1570 bgr_0.V_mir2.t19 GNDA 0.042444f
C1571 bgr_0.V_mir2.t22 GNDA 0.06851f
C1572 bgr_0.V_mir2.n9 GNDA 0.076506f
C1573 bgr_0.V_mir2.n10 GNDA 0.052264f
C1574 bgr_0.V_mir2.t6 GNDA 0.053881f
C1575 bgr_0.V_mir2.n11 GNDA 0.081315f
C1576 bgr_0.V_mir2.t9 GNDA 0.03537f
C1577 bgr_0.V_mir2.t7 GNDA 0.03537f
C1578 bgr_0.V_mir2.n12 GNDA 0.08097f
C1579 bgr_0.V_mir2.n13 GNDA 0.156007f
C1580 bgr_0.V_mir2.n14 GNDA 0.09373f
C1581 bgr_0.V_mir2.n15 GNDA 0.699157f
C1582 bgr_0.V_mir2.t10 GNDA 0.042444f
C1583 bgr_0.V_mir2.t21 GNDA 0.042444f
C1584 bgr_0.V_mir2.t17 GNDA 0.06851f
C1585 bgr_0.V_mir2.n16 GNDA 0.076506f
C1586 bgr_0.V_mir2.n17 GNDA 0.052264f
C1587 bgr_0.V_mir2.t2 GNDA 0.053881f
C1588 bgr_0.V_mir2.n18 GNDA 0.081315f
C1589 bgr_0.V_mir2.n19 GNDA 0.203577f
C1590 bgr_0.V_mir2.t3 GNDA 0.03537f
C1591 bgr_0.V_mir2.n20 GNDA 0.08097f
C1592 bgr_0.V_mir2.t11 GNDA 0.03537f
C1593 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t15 GNDA 0.035433f
C1594 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t0 GNDA 0.035433f
C1595 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n0 GNDA 0.088857f
C1596 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t1 GNDA 0.035433f
C1597 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t3 GNDA 0.035433f
C1598 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n1 GNDA 0.088389f
C1599 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n2 GNDA 0.598744f
C1600 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t2 GNDA 0.035433f
C1601 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t14 GNDA 0.035433f
C1602 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n3 GNDA 0.088389f
C1603 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n4 GNDA 0.629136f
C1604 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t16 GNDA 0.453797f
C1605 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t8 GNDA 0.070867f
C1606 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t4 GNDA 0.070867f
C1607 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n5 GNDA 0.20792f
C1608 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t7 GNDA 0.070867f
C1609 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t13 GNDA 0.070867f
C1610 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n6 GNDA 0.206976f
C1611 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n7 GNDA 0.715428f
C1612 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t11 GNDA 0.070867f
C1613 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t6 GNDA 0.070867f
C1614 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n8 GNDA 0.206976f
C1615 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n9 GNDA 0.370588f
C1616 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t10 GNDA 0.070867f
C1617 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t5 GNDA 0.070867f
C1618 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n10 GNDA 0.206976f
C1619 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n11 GNDA 0.370588f
C1620 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t9 GNDA 0.070867f
C1621 two_stage_opamp_dummy_magic_0.V_CMFB_S3.t12 GNDA 0.070867f
C1622 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n12 GNDA 0.206976f
C1623 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n13 GNDA 0.532409f
C1624 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n14 GNDA 3.84512f
C1625 two_stage_opamp_dummy_magic_0.V_CMFB_S3.n15 GNDA 2.74603f
C1626 bgr_0.V_CMFB_S3 GNDA 0.015439f
C1627 two_stage_opamp_dummy_magic_0.Y.t6 GNDA 0.023873f
C1628 two_stage_opamp_dummy_magic_0.Y.t11 GNDA 0.023873f
C1629 two_stage_opamp_dummy_magic_0.Y.n0 GNDA 0.080602f
C1630 two_stage_opamp_dummy_magic_0.Y.t19 GNDA 0.023873f
C1631 two_stage_opamp_dummy_magic_0.Y.t5 GNDA 0.023873f
C1632 two_stage_opamp_dummy_magic_0.Y.n1 GNDA 0.086146f
C1633 two_stage_opamp_dummy_magic_0.Y.t1 GNDA 0.023873f
C1634 two_stage_opamp_dummy_magic_0.Y.t22 GNDA 0.023873f
C1635 two_stage_opamp_dummy_magic_0.Y.n2 GNDA 0.085394f
C1636 two_stage_opamp_dummy_magic_0.Y.n3 GNDA 0.317069f
C1637 two_stage_opamp_dummy_magic_0.Y.t24 GNDA 0.023873f
C1638 two_stage_opamp_dummy_magic_0.Y.t15 GNDA 0.023873f
C1639 two_stage_opamp_dummy_magic_0.Y.n4 GNDA 0.085394f
C1640 two_stage_opamp_dummy_magic_0.Y.n5 GNDA 0.164481f
C1641 two_stage_opamp_dummy_magic_0.Y.t14 GNDA 0.023873f
C1642 two_stage_opamp_dummy_magic_0.Y.t9 GNDA 0.023873f
C1643 two_stage_opamp_dummy_magic_0.Y.n6 GNDA 0.085394f
C1644 two_stage_opamp_dummy_magic_0.Y.n7 GNDA 0.164481f
C1645 two_stage_opamp_dummy_magic_0.Y.t18 GNDA 0.023873f
C1646 two_stage_opamp_dummy_magic_0.Y.t20 GNDA 0.023873f
C1647 two_stage_opamp_dummy_magic_0.Y.n8 GNDA 0.086146f
C1648 two_stage_opamp_dummy_magic_0.Y.n9 GNDA 0.200335f
C1649 two_stage_opamp_dummy_magic_0.Y.n10 GNDA 0.250257f
C1650 two_stage_opamp_dummy_magic_0.Y.t7 GNDA 0.055705f
C1651 two_stage_opamp_dummy_magic_0.Y.t17 GNDA 0.055705f
C1652 two_stage_opamp_dummy_magic_0.Y.n11 GNDA 0.193729f
C1653 two_stage_opamp_dummy_magic_0.Y.t4 GNDA 0.055705f
C1654 two_stage_opamp_dummy_magic_0.Y.t2 GNDA 0.055705f
C1655 two_stage_opamp_dummy_magic_0.Y.n12 GNDA 0.193042f
C1656 two_stage_opamp_dummy_magic_0.Y.n13 GNDA 0.364444f
C1657 two_stage_opamp_dummy_magic_0.Y.t16 GNDA 0.055705f
C1658 two_stage_opamp_dummy_magic_0.Y.t21 GNDA 0.055705f
C1659 two_stage_opamp_dummy_magic_0.Y.n14 GNDA 0.193042f
C1660 two_stage_opamp_dummy_magic_0.Y.n15 GNDA 0.188932f
C1661 two_stage_opamp_dummy_magic_0.Y.t23 GNDA 0.055705f
C1662 two_stage_opamp_dummy_magic_0.Y.t13 GNDA 0.055705f
C1663 two_stage_opamp_dummy_magic_0.Y.n16 GNDA 0.193042f
C1664 two_stage_opamp_dummy_magic_0.Y.n17 GNDA 0.188932f
C1665 two_stage_opamp_dummy_magic_0.Y.t3 GNDA 0.055705f
C1666 two_stage_opamp_dummy_magic_0.Y.t8 GNDA 0.055705f
C1667 two_stage_opamp_dummy_magic_0.Y.n18 GNDA 0.193042f
C1668 two_stage_opamp_dummy_magic_0.Y.n19 GNDA 0.222471f
C1669 two_stage_opamp_dummy_magic_0.Y.t10 GNDA 0.055705f
C1670 two_stage_opamp_dummy_magic_0.Y.t12 GNDA 0.055705f
C1671 two_stage_opamp_dummy_magic_0.Y.n20 GNDA 0.189043f
C1672 two_stage_opamp_dummy_magic_0.Y.n21 GNDA 0.376251f
C1673 two_stage_opamp_dummy_magic_0.Y.t52 GNDA 0.033423f
C1674 two_stage_opamp_dummy_magic_0.Y.t38 GNDA 0.040585f
C1675 two_stage_opamp_dummy_magic_0.Y.n22 GNDA 0.037846f
C1676 two_stage_opamp_dummy_magic_0.Y.t42 GNDA 0.033423f
C1677 two_stage_opamp_dummy_magic_0.Y.t25 GNDA 0.033423f
C1678 two_stage_opamp_dummy_magic_0.Y.t30 GNDA 0.033423f
C1679 two_stage_opamp_dummy_magic_0.Y.t47 GNDA 0.033423f
C1680 two_stage_opamp_dummy_magic_0.Y.t33 GNDA 0.033423f
C1681 two_stage_opamp_dummy_magic_0.Y.t49 GNDA 0.033423f
C1682 two_stage_opamp_dummy_magic_0.Y.t37 GNDA 0.033423f
C1683 two_stage_opamp_dummy_magic_0.Y.t29 GNDA 0.040585f
C1684 two_stage_opamp_dummy_magic_0.Y.n23 GNDA 0.040585f
C1685 two_stage_opamp_dummy_magic_0.Y.n24 GNDA 0.026261f
C1686 two_stage_opamp_dummy_magic_0.Y.n25 GNDA 0.026261f
C1687 two_stage_opamp_dummy_magic_0.Y.n26 GNDA 0.026261f
C1688 two_stage_opamp_dummy_magic_0.Y.n27 GNDA 0.026261f
C1689 two_stage_opamp_dummy_magic_0.Y.n28 GNDA 0.026261f
C1690 two_stage_opamp_dummy_magic_0.Y.n29 GNDA 0.023522f
C1691 two_stage_opamp_dummy_magic_0.Y.n30 GNDA 0.023134f
C1692 two_stage_opamp_dummy_magic_0.Y.t27 GNDA 0.051328f
C1693 two_stage_opamp_dummy_magic_0.Y.t45 GNDA 0.058351f
C1694 two_stage_opamp_dummy_magic_0.Y.n31 GNDA 0.049922f
C1695 two_stage_opamp_dummy_magic_0.Y.t46 GNDA 0.051328f
C1696 two_stage_opamp_dummy_magic_0.Y.t28 GNDA 0.051328f
C1697 two_stage_opamp_dummy_magic_0.Y.t36 GNDA 0.051328f
C1698 two_stage_opamp_dummy_magic_0.Y.t51 GNDA 0.051328f
C1699 two_stage_opamp_dummy_magic_0.Y.t41 GNDA 0.051328f
C1700 two_stage_opamp_dummy_magic_0.Y.t54 GNDA 0.051328f
C1701 two_stage_opamp_dummy_magic_0.Y.t44 GNDA 0.051328f
C1702 two_stage_opamp_dummy_magic_0.Y.t34 GNDA 0.058351f
C1703 two_stage_opamp_dummy_magic_0.Y.n32 GNDA 0.05266f
C1704 two_stage_opamp_dummy_magic_0.Y.n33 GNDA 0.032229f
C1705 two_stage_opamp_dummy_magic_0.Y.n34 GNDA 0.032229f
C1706 two_stage_opamp_dummy_magic_0.Y.n35 GNDA 0.032229f
C1707 two_stage_opamp_dummy_magic_0.Y.n36 GNDA 0.032229f
C1708 two_stage_opamp_dummy_magic_0.Y.n37 GNDA 0.032229f
C1709 two_stage_opamp_dummy_magic_0.Y.n38 GNDA 0.02949f
C1710 two_stage_opamp_dummy_magic_0.Y.n39 GNDA 0.023086f
C1711 two_stage_opamp_dummy_magic_0.Y.n40 GNDA 0.249706f
C1712 two_stage_opamp_dummy_magic_0.Y.n41 GNDA 0.51804f
C1713 two_stage_opamp_dummy_magic_0.Y.n42 GNDA 0.261996f
C1714 two_stage_opamp_dummy_magic_0.Y.t35 GNDA 0.105043f
C1715 two_stage_opamp_dummy_magic_0.Y.t48 GNDA 0.105043f
C1716 two_stage_opamp_dummy_magic_0.Y.t32 GNDA 0.105043f
C1717 two_stage_opamp_dummy_magic_0.Y.t26 GNDA 0.105043f
C1718 two_stage_opamp_dummy_magic_0.Y.t43 GNDA 0.105043f
C1719 two_stage_opamp_dummy_magic_0.Y.t53 GNDA 0.105043f
C1720 two_stage_opamp_dummy_magic_0.Y.t40 GNDA 0.111878f
C1721 two_stage_opamp_dummy_magic_0.Y.n43 GNDA 0.088659f
C1722 two_stage_opamp_dummy_magic_0.Y.n44 GNDA 0.050134f
C1723 two_stage_opamp_dummy_magic_0.Y.n45 GNDA 0.050134f
C1724 two_stage_opamp_dummy_magic_0.Y.n46 GNDA 0.050134f
C1725 two_stage_opamp_dummy_magic_0.Y.n47 GNDA 0.050134f
C1726 two_stage_opamp_dummy_magic_0.Y.n48 GNDA 0.047395f
C1727 two_stage_opamp_dummy_magic_0.Y.t50 GNDA 0.105043f
C1728 two_stage_opamp_dummy_magic_0.Y.t39 GNDA 0.105043f
C1729 two_stage_opamp_dummy_magic_0.Y.t31 GNDA 0.111878f
C1730 two_stage_opamp_dummy_magic_0.Y.n49 GNDA 0.088659f
C1731 two_stage_opamp_dummy_magic_0.Y.n50 GNDA 0.047395f
C1732 two_stage_opamp_dummy_magic_0.Y.n51 GNDA 0.025681f
C1733 two_stage_opamp_dummy_magic_0.Y.n52 GNDA 0.925108f
C1734 two_stage_opamp_dummy_magic_0.Y.t0 GNDA 0.777549f
C1735 two_stage_opamp_dummy_magic_0.cap_res_Y.t2 GNDA 0.343499f
C1736 two_stage_opamp_dummy_magic_0.cap_res_Y.t76 GNDA 0.344645f
C1737 two_stage_opamp_dummy_magic_0.cap_res_Y.t38 GNDA 0.185116f
C1738 two_stage_opamp_dummy_magic_0.cap_res_Y.n0 GNDA 0.197667f
C1739 two_stage_opamp_dummy_magic_0.cap_res_Y.t37 GNDA 0.343499f
C1740 two_stage_opamp_dummy_magic_0.cap_res_Y.t120 GNDA 0.344645f
C1741 two_stage_opamp_dummy_magic_0.cap_res_Y.t75 GNDA 0.185116f
C1742 two_stage_opamp_dummy_magic_0.cap_res_Y.n1 GNDA 0.216163f
C1743 two_stage_opamp_dummy_magic_0.cap_res_Y.t23 GNDA 0.343499f
C1744 two_stage_opamp_dummy_magic_0.cap_res_Y.t98 GNDA 0.344645f
C1745 two_stage_opamp_dummy_magic_0.cap_res_Y.t60 GNDA 0.185116f
C1746 two_stage_opamp_dummy_magic_0.cap_res_Y.n2 GNDA 0.216163f
C1747 two_stage_opamp_dummy_magic_0.cap_res_Y.t55 GNDA 0.343499f
C1748 two_stage_opamp_dummy_magic_0.cap_res_Y.t131 GNDA 0.344645f
C1749 two_stage_opamp_dummy_magic_0.cap_res_Y.t94 GNDA 0.185116f
C1750 two_stage_opamp_dummy_magic_0.cap_res_Y.n3 GNDA 0.216163f
C1751 two_stage_opamp_dummy_magic_0.cap_res_Y.t92 GNDA 0.343499f
C1752 two_stage_opamp_dummy_magic_0.cap_res_Y.t43 GNDA 0.344645f
C1753 two_stage_opamp_dummy_magic_0.cap_res_Y.t136 GNDA 0.363141f
C1754 two_stage_opamp_dummy_magic_0.cap_res_Y.t31 GNDA 0.363141f
C1755 two_stage_opamp_dummy_magic_0.cap_res_Y.t130 GNDA 0.185116f
C1756 two_stage_opamp_dummy_magic_0.cap_res_Y.n4 GNDA 0.216163f
C1757 two_stage_opamp_dummy_magic_0.cap_res_Y.t70 GNDA 0.343499f
C1758 two_stage_opamp_dummy_magic_0.cap_res_Y.t95 GNDA 0.344645f
C1759 two_stage_opamp_dummy_magic_0.cap_res_Y.t116 GNDA 0.363141f
C1760 two_stage_opamp_dummy_magic_0.cap_res_Y.t14 GNDA 0.363141f
C1761 two_stage_opamp_dummy_magic_0.cap_res_Y.t112 GNDA 0.185116f
C1762 two_stage_opamp_dummy_magic_0.cap_res_Y.n5 GNDA 0.216163f
C1763 two_stage_opamp_dummy_magic_0.cap_res_Y.t117 GNDA 0.344645f
C1764 two_stage_opamp_dummy_magic_0.cap_res_Y.t138 GNDA 0.345894f
C1765 two_stage_opamp_dummy_magic_0.cap_res_Y.t72 GNDA 0.344645f
C1766 two_stage_opamp_dummy_magic_0.cap_res_Y.t100 GNDA 0.347347f
C1767 two_stage_opamp_dummy_magic_0.cap_res_Y.t61 GNDA 0.377789f
C1768 two_stage_opamp_dummy_magic_0.cap_res_Y.t123 GNDA 0.344645f
C1769 two_stage_opamp_dummy_magic_0.cap_res_Y.t105 GNDA 0.345894f
C1770 two_stage_opamp_dummy_magic_0.cap_res_Y.t21 GNDA 0.344645f
C1771 two_stage_opamp_dummy_magic_0.cap_res_Y.t36 GNDA 0.345894f
C1772 two_stage_opamp_dummy_magic_0.cap_res_Y.t87 GNDA 0.344645f
C1773 two_stage_opamp_dummy_magic_0.cap_res_Y.t68 GNDA 0.345894f
C1774 two_stage_opamp_dummy_magic_0.cap_res_Y.t121 GNDA 0.344645f
C1775 two_stage_opamp_dummy_magic_0.cap_res_Y.t6 GNDA 0.345894f
C1776 two_stage_opamp_dummy_magic_0.cap_res_Y.t62 GNDA 0.344645f
C1777 two_stage_opamp_dummy_magic_0.cap_res_Y.t114 GNDA 0.345894f
C1778 two_stage_opamp_dummy_magic_0.cap_res_Y.t91 GNDA 0.344645f
C1779 two_stage_opamp_dummy_magic_0.cap_res_Y.t39 GNDA 0.345894f
C1780 two_stage_opamp_dummy_magic_0.cap_res_Y.t102 GNDA 0.344645f
C1781 two_stage_opamp_dummy_magic_0.cap_res_Y.t16 GNDA 0.345894f
C1782 two_stage_opamp_dummy_magic_0.cap_res_Y.t128 GNDA 0.344645f
C1783 two_stage_opamp_dummy_magic_0.cap_res_Y.t77 GNDA 0.345894f
C1784 two_stage_opamp_dummy_magic_0.cap_res_Y.t66 GNDA 0.344645f
C1785 two_stage_opamp_dummy_magic_0.cap_res_Y.t118 GNDA 0.345894f
C1786 two_stage_opamp_dummy_magic_0.cap_res_Y.t99 GNDA 0.344645f
C1787 two_stage_opamp_dummy_magic_0.cap_res_Y.t48 GNDA 0.345894f
C1788 two_stage_opamp_dummy_magic_0.cap_res_Y.t108 GNDA 0.344645f
C1789 two_stage_opamp_dummy_magic_0.cap_res_Y.t22 GNDA 0.345894f
C1790 two_stage_opamp_dummy_magic_0.cap_res_Y.t137 GNDA 0.344645f
C1791 two_stage_opamp_dummy_magic_0.cap_res_Y.t85 GNDA 0.345894f
C1792 two_stage_opamp_dummy_magic_0.cap_res_Y.t9 GNDA 0.344645f
C1793 two_stage_opamp_dummy_magic_0.cap_res_Y.t58 GNDA 0.345894f
C1794 two_stage_opamp_dummy_magic_0.cap_res_Y.t35 GNDA 0.344645f
C1795 two_stage_opamp_dummy_magic_0.cap_res_Y.t124 GNDA 0.345894f
C1796 two_stage_opamp_dummy_magic_0.cap_res_Y.t113 GNDA 0.344645f
C1797 two_stage_opamp_dummy_magic_0.cap_res_Y.t24 GNDA 0.345894f
C1798 two_stage_opamp_dummy_magic_0.cap_res_Y.t5 GNDA 0.344645f
C1799 two_stage_opamp_dummy_magic_0.cap_res_Y.t90 GNDA 0.345894f
C1800 two_stage_opamp_dummy_magic_0.cap_res_Y.t15 GNDA 0.344645f
C1801 two_stage_opamp_dummy_magic_0.cap_res_Y.t63 GNDA 0.345894f
C1802 two_stage_opamp_dummy_magic_0.cap_res_Y.t41 GNDA 0.344645f
C1803 two_stage_opamp_dummy_magic_0.cap_res_Y.t127 GNDA 0.345894f
C1804 two_stage_opamp_dummy_magic_0.cap_res_Y.t52 GNDA 0.344645f
C1805 two_stage_opamp_dummy_magic_0.cap_res_Y.t104 GNDA 0.345894f
C1806 two_stage_opamp_dummy_magic_0.cap_res_Y.t80 GNDA 0.344645f
C1807 two_stage_opamp_dummy_magic_0.cap_res_Y.t30 GNDA 0.345894f
C1808 two_stage_opamp_dummy_magic_0.cap_res_Y.t88 GNDA 0.344645f
C1809 two_stage_opamp_dummy_magic_0.cap_res_Y.t3 GNDA 0.345894f
C1810 two_stage_opamp_dummy_magic_0.cap_res_Y.t122 GNDA 0.344645f
C1811 two_stage_opamp_dummy_magic_0.cap_res_Y.t71 GNDA 0.345894f
C1812 two_stage_opamp_dummy_magic_0.cap_res_Y.t57 GNDA 0.344645f
C1813 two_stage_opamp_dummy_magic_0.cap_res_Y.t110 GNDA 0.345894f
C1814 two_stage_opamp_dummy_magic_0.cap_res_Y.t86 GNDA 0.344645f
C1815 two_stage_opamp_dummy_magic_0.cap_res_Y.t34 GNDA 0.345894f
C1816 two_stage_opamp_dummy_magic_0.cap_res_Y.t96 GNDA 0.344645f
C1817 two_stage_opamp_dummy_magic_0.cap_res_Y.t10 GNDA 0.345894f
C1818 two_stage_opamp_dummy_magic_0.cap_res_Y.t125 GNDA 0.344645f
C1819 two_stage_opamp_dummy_magic_0.cap_res_Y.t74 GNDA 0.345894f
C1820 two_stage_opamp_dummy_magic_0.cap_res_Y.t133 GNDA 0.344645f
C1821 two_stage_opamp_dummy_magic_0.cap_res_Y.t44 GNDA 0.345894f
C1822 two_stage_opamp_dummy_magic_0.cap_res_Y.t28 GNDA 0.344645f
C1823 two_stage_opamp_dummy_magic_0.cap_res_Y.t119 GNDA 0.345894f
C1824 two_stage_opamp_dummy_magic_0.cap_res_Y.t7 GNDA 0.344645f
C1825 two_stage_opamp_dummy_magic_0.cap_res_Y.t69 GNDA 0.361543f
C1826 two_stage_opamp_dummy_magic_0.cap_res_Y.t93 GNDA 0.344645f
C1827 two_stage_opamp_dummy_magic_0.cap_res_Y.t106 GNDA 0.185116f
C1828 two_stage_opamp_dummy_magic_0.cap_res_Y.n6 GNDA 0.19812f
C1829 two_stage_opamp_dummy_magic_0.cap_res_Y.t134 GNDA 0.344645f
C1830 two_stage_opamp_dummy_magic_0.cap_res_Y.t20 GNDA 0.185116f
C1831 two_stage_opamp_dummy_magic_0.cap_res_Y.n7 GNDA 0.196521f
C1832 two_stage_opamp_dummy_magic_0.cap_res_Y.t83 GNDA 0.344645f
C1833 two_stage_opamp_dummy_magic_0.cap_res_Y.t51 GNDA 0.185116f
C1834 two_stage_opamp_dummy_magic_0.cap_res_Y.n8 GNDA 0.196521f
C1835 two_stage_opamp_dummy_magic_0.cap_res_Y.t32 GNDA 0.344645f
C1836 two_stage_opamp_dummy_magic_0.cap_res_Y.t82 GNDA 0.185116f
C1837 two_stage_opamp_dummy_magic_0.cap_res_Y.n9 GNDA 0.196521f
C1838 two_stage_opamp_dummy_magic_0.cap_res_Y.t73 GNDA 0.344645f
C1839 two_stage_opamp_dummy_magic_0.cap_res_Y.t132 GNDA 0.185116f
C1840 two_stage_opamp_dummy_magic_0.cap_res_Y.n10 GNDA 0.196521f
C1841 two_stage_opamp_dummy_magic_0.cap_res_Y.t27 GNDA 0.344645f
C1842 two_stage_opamp_dummy_magic_0.cap_res_Y.t29 GNDA 0.185116f
C1843 two_stage_opamp_dummy_magic_0.cap_res_Y.n11 GNDA 0.196521f
C1844 two_stage_opamp_dummy_magic_0.cap_res_Y.t115 GNDA 0.344645f
C1845 two_stage_opamp_dummy_magic_0.cap_res_Y.t67 GNDA 0.185116f
C1846 two_stage_opamp_dummy_magic_0.cap_res_Y.n12 GNDA 0.196521f
C1847 two_stage_opamp_dummy_magic_0.cap_res_Y.t65 GNDA 0.344645f
C1848 two_stage_opamp_dummy_magic_0.cap_res_Y.t103 GNDA 0.185116f
C1849 two_stage_opamp_dummy_magic_0.cap_res_Y.n13 GNDA 0.196521f
C1850 two_stage_opamp_dummy_magic_0.cap_res_Y.t109 GNDA 0.344645f
C1851 two_stage_opamp_dummy_magic_0.cap_res_Y.t17 GNDA 0.185116f
C1852 two_stage_opamp_dummy_magic_0.cap_res_Y.n14 GNDA 0.196521f
C1853 two_stage_opamp_dummy_magic_0.cap_res_Y.t129 GNDA 0.344645f
C1854 two_stage_opamp_dummy_magic_0.cap_res_Y.t78 GNDA 0.345894f
C1855 two_stage_opamp_dummy_magic_0.cap_res_Y.t49 GNDA 0.344645f
C1856 two_stage_opamp_dummy_magic_0.cap_res_Y.t8 GNDA 0.345894f
C1857 two_stage_opamp_dummy_magic_0.cap_res_Y.t56 GNDA 0.166619f
C1858 two_stage_opamp_dummy_magic_0.cap_res_Y.n15 GNDA 0.214914f
C1859 two_stage_opamp_dummy_magic_0.cap_res_Y.t47 GNDA 0.18397f
C1860 two_stage_opamp_dummy_magic_0.cap_res_Y.n16 GNDA 0.23341f
C1861 two_stage_opamp_dummy_magic_0.cap_res_Y.t79 GNDA 0.18397f
C1862 two_stage_opamp_dummy_magic_0.cap_res_Y.n17 GNDA 0.250658f
C1863 two_stage_opamp_dummy_magic_0.cap_res_Y.t40 GNDA 0.18397f
C1864 two_stage_opamp_dummy_magic_0.cap_res_Y.n18 GNDA 0.250658f
C1865 two_stage_opamp_dummy_magic_0.cap_res_Y.t4 GNDA 0.18397f
C1866 two_stage_opamp_dummy_magic_0.cap_res_Y.n19 GNDA 0.250658f
C1867 two_stage_opamp_dummy_magic_0.cap_res_Y.t33 GNDA 0.18397f
C1868 two_stage_opamp_dummy_magic_0.cap_res_Y.n20 GNDA 0.250658f
C1869 two_stage_opamp_dummy_magic_0.cap_res_Y.t135 GNDA 0.18397f
C1870 two_stage_opamp_dummy_magic_0.cap_res_Y.n21 GNDA 0.250658f
C1871 two_stage_opamp_dummy_magic_0.cap_res_Y.t97 GNDA 0.18397f
C1872 two_stage_opamp_dummy_magic_0.cap_res_Y.n22 GNDA 0.250658f
C1873 two_stage_opamp_dummy_magic_0.cap_res_Y.t59 GNDA 0.18397f
C1874 two_stage_opamp_dummy_magic_0.cap_res_Y.n23 GNDA 0.250658f
C1875 two_stage_opamp_dummy_magic_0.cap_res_Y.t89 GNDA 0.18397f
C1876 two_stage_opamp_dummy_magic_0.cap_res_Y.n24 GNDA 0.250658f
C1877 two_stage_opamp_dummy_magic_0.cap_res_Y.t54 GNDA 0.18397f
C1878 two_stage_opamp_dummy_magic_0.cap_res_Y.n25 GNDA 0.250658f
C1879 two_stage_opamp_dummy_magic_0.cap_res_Y.t18 GNDA 0.18397f
C1880 two_stage_opamp_dummy_magic_0.cap_res_Y.n26 GNDA 0.250658f
C1881 two_stage_opamp_dummy_magic_0.cap_res_Y.t46 GNDA 0.18397f
C1882 two_stage_opamp_dummy_magic_0.cap_res_Y.n27 GNDA 0.250658f
C1883 two_stage_opamp_dummy_magic_0.cap_res_Y.t12 GNDA 0.18397f
C1884 two_stage_opamp_dummy_magic_0.cap_res_Y.n28 GNDA 0.250658f
C1885 two_stage_opamp_dummy_magic_0.cap_res_Y.t107 GNDA 0.18397f
C1886 two_stage_opamp_dummy_magic_0.cap_res_Y.n29 GNDA 0.250658f
C1887 two_stage_opamp_dummy_magic_0.cap_res_Y.t1 GNDA 0.18397f
C1888 two_stage_opamp_dummy_magic_0.cap_res_Y.n30 GNDA 0.250658f
C1889 two_stage_opamp_dummy_magic_0.cap_res_Y.t101 GNDA 0.18397f
C1890 two_stage_opamp_dummy_magic_0.cap_res_Y.n31 GNDA 0.23341f
C1891 two_stage_opamp_dummy_magic_0.cap_res_Y.t25 GNDA 0.343499f
C1892 two_stage_opamp_dummy_magic_0.cap_res_Y.t64 GNDA 0.166619f
C1893 two_stage_opamp_dummy_magic_0.cap_res_Y.n32 GNDA 0.216163f
C1894 two_stage_opamp_dummy_magic_0.cap_res_Y.t42 GNDA 0.343499f
C1895 two_stage_opamp_dummy_magic_0.cap_res_Y.t81 GNDA 0.166619f
C1896 two_stage_opamp_dummy_magic_0.cap_res_Y.n33 GNDA 0.216163f
C1897 two_stage_opamp_dummy_magic_0.cap_res_Y.t11 GNDA 0.343499f
C1898 two_stage_opamp_dummy_magic_0.cap_res_Y.t26 GNDA 0.344645f
C1899 two_stage_opamp_dummy_magic_0.cap_res_Y.t53 GNDA 0.363141f
C1900 two_stage_opamp_dummy_magic_0.cap_res_Y.t84 GNDA 0.363141f
C1901 two_stage_opamp_dummy_magic_0.cap_res_Y.t45 GNDA 0.185116f
C1902 two_stage_opamp_dummy_magic_0.cap_res_Y.n34 GNDA 0.216163f
C1903 two_stage_opamp_dummy_magic_0.cap_res_Y.t111 GNDA 0.343499f
C1904 two_stage_opamp_dummy_magic_0.cap_res_Y.n35 GNDA 0.216163f
C1905 two_stage_opamp_dummy_magic_0.cap_res_Y.t13 GNDA 0.185116f
C1906 two_stage_opamp_dummy_magic_0.cap_res_Y.t50 GNDA 0.363141f
C1907 two_stage_opamp_dummy_magic_0.cap_res_Y.t19 GNDA 0.363141f
C1908 two_stage_opamp_dummy_magic_0.cap_res_Y.t126 GNDA 0.434494f
C1909 two_stage_opamp_dummy_magic_0.cap_res_Y.t0 GNDA 0.297192f
C1910 two_stage_opamp_dummy_magic_0.VOUT+.t15 GNDA 0.050892f
C1911 two_stage_opamp_dummy_magic_0.VOUT+.t16 GNDA 0.050892f
C1912 two_stage_opamp_dummy_magic_0.VOUT+.n0 GNDA 0.235428f
C1913 two_stage_opamp_dummy_magic_0.VOUT+.t18 GNDA 0.050892f
C1914 two_stage_opamp_dummy_magic_0.VOUT+.t3 GNDA 0.050892f
C1915 two_stage_opamp_dummy_magic_0.VOUT+.n1 GNDA 0.23464f
C1916 two_stage_opamp_dummy_magic_0.VOUT+.n2 GNDA 0.144996f
C1917 two_stage_opamp_dummy_magic_0.VOUT+.t4 GNDA 0.050892f
C1918 two_stage_opamp_dummy_magic_0.VOUT+.t14 GNDA 0.050892f
C1919 two_stage_opamp_dummy_magic_0.VOUT+.n3 GNDA 0.23464f
C1920 two_stage_opamp_dummy_magic_0.VOUT+.n4 GNDA 0.08925f
C1921 two_stage_opamp_dummy_magic_0.VOUT+.t12 GNDA 0.043622f
C1922 two_stage_opamp_dummy_magic_0.VOUT+.t7 GNDA 0.043622f
C1923 two_stage_opamp_dummy_magic_0.VOUT+.n5 GNDA 0.175328f
C1924 two_stage_opamp_dummy_magic_0.VOUT+.t8 GNDA 0.043622f
C1925 two_stage_opamp_dummy_magic_0.VOUT+.t13 GNDA 0.043622f
C1926 two_stage_opamp_dummy_magic_0.VOUT+.n6 GNDA 0.175327f
C1927 two_stage_opamp_dummy_magic_0.VOUT+.t5 GNDA 0.043622f
C1928 two_stage_opamp_dummy_magic_0.VOUT+.t0 GNDA 0.043622f
C1929 two_stage_opamp_dummy_magic_0.VOUT+.n7 GNDA 0.175005f
C1930 two_stage_opamp_dummy_magic_0.VOUT+.n8 GNDA 0.1724f
C1931 two_stage_opamp_dummy_magic_0.VOUT+.t10 GNDA 0.043622f
C1932 two_stage_opamp_dummy_magic_0.VOUT+.t9 GNDA 0.043622f
C1933 two_stage_opamp_dummy_magic_0.VOUT+.n9 GNDA 0.175005f
C1934 two_stage_opamp_dummy_magic_0.VOUT+.n10 GNDA 0.088906f
C1935 two_stage_opamp_dummy_magic_0.VOUT+.t1 GNDA 0.043622f
C1936 two_stage_opamp_dummy_magic_0.VOUT+.t2 GNDA 0.043622f
C1937 two_stage_opamp_dummy_magic_0.VOUT+.n11 GNDA 0.175005f
C1938 two_stage_opamp_dummy_magic_0.VOUT+.n12 GNDA 0.088906f
C1939 two_stage_opamp_dummy_magic_0.VOUT+.n13 GNDA 0.105305f
C1940 two_stage_opamp_dummy_magic_0.VOUT+.t11 GNDA 0.043622f
C1941 two_stage_opamp_dummy_magic_0.VOUT+.t6 GNDA 0.043622f
C1942 two_stage_opamp_dummy_magic_0.VOUT+.n14 GNDA 0.172862f
C1943 two_stage_opamp_dummy_magic_0.VOUT+.n15 GNDA 0.212252f
C1944 two_stage_opamp_dummy_magic_0.VOUT+.t101 GNDA 0.290811f
C1945 two_stage_opamp_dummy_magic_0.VOUT+.t108 GNDA 0.295764f
C1946 two_stage_opamp_dummy_magic_0.VOUT+.t149 GNDA 0.290811f
C1947 two_stage_opamp_dummy_magic_0.VOUT+.n16 GNDA 0.194979f
C1948 two_stage_opamp_dummy_magic_0.VOUT+.n17 GNDA 0.12723f
C1949 two_stage_opamp_dummy_magic_0.VOUT+.t48 GNDA 0.295144f
C1950 two_stage_opamp_dummy_magic_0.VOUT+.t92 GNDA 0.295144f
C1951 two_stage_opamp_dummy_magic_0.VOUT+.t42 GNDA 0.295144f
C1952 two_stage_opamp_dummy_magic_0.VOUT+.t130 GNDA 0.295144f
C1953 two_stage_opamp_dummy_magic_0.VOUT+.t84 GNDA 0.295144f
C1954 two_stage_opamp_dummy_magic_0.VOUT+.t125 GNDA 0.295144f
C1955 two_stage_opamp_dummy_magic_0.VOUT+.t74 GNDA 0.295144f
C1956 two_stage_opamp_dummy_magic_0.VOUT+.t23 GNDA 0.295144f
C1957 two_stage_opamp_dummy_magic_0.VOUT+.t64 GNDA 0.295144f
C1958 two_stage_opamp_dummy_magic_0.VOUT+.t150 GNDA 0.295144f
C1959 two_stage_opamp_dummy_magic_0.VOUT+.t88 GNDA 0.290811f
C1960 two_stage_opamp_dummy_magic_0.VOUT+.n18 GNDA 0.195599f
C1961 two_stage_opamp_dummy_magic_0.VOUT+.t51 GNDA 0.290811f
C1962 two_stage_opamp_dummy_magic_0.VOUT+.n19 GNDA 0.250126f
C1963 two_stage_opamp_dummy_magic_0.VOUT+.t137 GNDA 0.290811f
C1964 two_stage_opamp_dummy_magic_0.VOUT+.n20 GNDA 0.250126f
C1965 two_stage_opamp_dummy_magic_0.VOUT+.t106 GNDA 0.290811f
C1966 two_stage_opamp_dummy_magic_0.VOUT+.n21 GNDA 0.250126f
C1967 two_stage_opamp_dummy_magic_0.VOUT+.t75 GNDA 0.290811f
C1968 two_stage_opamp_dummy_magic_0.VOUT+.n22 GNDA 0.250126f
C1969 two_stage_opamp_dummy_magic_0.VOUT+.t25 GNDA 0.290811f
C1970 two_stage_opamp_dummy_magic_0.VOUT+.n23 GNDA 0.250126f
C1971 two_stage_opamp_dummy_magic_0.VOUT+.t128 GNDA 0.290811f
C1972 two_stage_opamp_dummy_magic_0.VOUT+.n24 GNDA 0.250126f
C1973 two_stage_opamp_dummy_magic_0.VOUT+.t90 GNDA 0.290811f
C1974 two_stage_opamp_dummy_magic_0.VOUT+.n25 GNDA 0.250126f
C1975 two_stage_opamp_dummy_magic_0.VOUT+.t54 GNDA 0.290811f
C1976 two_stage_opamp_dummy_magic_0.VOUT+.n26 GNDA 0.250126f
C1977 two_stage_opamp_dummy_magic_0.VOUT+.t140 GNDA 0.290811f
C1978 two_stage_opamp_dummy_magic_0.VOUT+.n27 GNDA 0.250126f
C1979 two_stage_opamp_dummy_magic_0.VOUT+.t110 GNDA 0.290811f
C1980 two_stage_opamp_dummy_magic_0.VOUT+.t28 GNDA 0.295764f
C1981 two_stage_opamp_dummy_magic_0.VOUT+.t79 GNDA 0.290811f
C1982 two_stage_opamp_dummy_magic_0.VOUT+.n28 GNDA 0.194979f
C1983 two_stage_opamp_dummy_magic_0.VOUT+.n29 GNDA 0.236284f
C1984 two_stage_opamp_dummy_magic_0.VOUT+.t24 GNDA 0.295764f
C1985 two_stage_opamp_dummy_magic_0.VOUT+.t113 GNDA 0.290811f
C1986 two_stage_opamp_dummy_magic_0.VOUT+.n30 GNDA 0.194979f
C1987 two_stage_opamp_dummy_magic_0.VOUT+.t78 GNDA 0.290811f
C1988 two_stage_opamp_dummy_magic_0.VOUT+.t129 GNDA 0.295764f
C1989 two_stage_opamp_dummy_magic_0.VOUT+.t38 GNDA 0.290811f
C1990 two_stage_opamp_dummy_magic_0.VOUT+.n31 GNDA 0.194979f
C1991 two_stage_opamp_dummy_magic_0.VOUT+.n32 GNDA 0.236284f
C1992 two_stage_opamp_dummy_magic_0.VOUT+.t61 GNDA 0.295764f
C1993 two_stage_opamp_dummy_magic_0.VOUT+.t147 GNDA 0.290811f
C1994 two_stage_opamp_dummy_magic_0.VOUT+.n33 GNDA 0.194979f
C1995 two_stage_opamp_dummy_magic_0.VOUT+.t117 GNDA 0.290811f
C1996 two_stage_opamp_dummy_magic_0.VOUT+.t32 GNDA 0.295764f
C1997 two_stage_opamp_dummy_magic_0.VOUT+.t83 GNDA 0.290811f
C1998 two_stage_opamp_dummy_magic_0.VOUT+.n34 GNDA 0.194979f
C1999 two_stage_opamp_dummy_magic_0.VOUT+.n35 GNDA 0.236284f
C2000 two_stage_opamp_dummy_magic_0.VOUT+.t100 GNDA 0.295764f
C2001 two_stage_opamp_dummy_magic_0.VOUT+.t47 GNDA 0.290811f
C2002 two_stage_opamp_dummy_magic_0.VOUT+.n36 GNDA 0.194979f
C2003 two_stage_opamp_dummy_magic_0.VOUT+.t153 GNDA 0.290811f
C2004 two_stage_opamp_dummy_magic_0.VOUT+.t71 GNDA 0.295764f
C2005 two_stage_opamp_dummy_magic_0.VOUT+.t123 GNDA 0.290811f
C2006 two_stage_opamp_dummy_magic_0.VOUT+.n37 GNDA 0.194979f
C2007 two_stage_opamp_dummy_magic_0.VOUT+.n38 GNDA 0.236284f
C2008 two_stage_opamp_dummy_magic_0.VOUT+.t69 GNDA 0.295764f
C2009 two_stage_opamp_dummy_magic_0.VOUT+.t154 GNDA 0.290811f
C2010 two_stage_opamp_dummy_magic_0.VOUT+.n39 GNDA 0.194979f
C2011 two_stage_opamp_dummy_magic_0.VOUT+.t124 GNDA 0.290811f
C2012 two_stage_opamp_dummy_magic_0.VOUT+.t35 GNDA 0.295764f
C2013 two_stage_opamp_dummy_magic_0.VOUT+.t86 GNDA 0.290811f
C2014 two_stage_opamp_dummy_magic_0.VOUT+.n40 GNDA 0.194979f
C2015 two_stage_opamp_dummy_magic_0.VOUT+.n41 GNDA 0.236284f
C2016 two_stage_opamp_dummy_magic_0.VOUT+.t96 GNDA 0.290811f
C2017 two_stage_opamp_dummy_magic_0.VOUT+.t85 GNDA 0.295764f
C2018 two_stage_opamp_dummy_magic_0.VOUT+.t57 GNDA 0.290811f
C2019 two_stage_opamp_dummy_magic_0.VOUT+.n42 GNDA 0.194979f
C2020 two_stage_opamp_dummy_magic_0.VOUT+.n43 GNDA 0.12723f
C2021 two_stage_opamp_dummy_magic_0.VOUT+.t132 GNDA 0.295144f
C2022 two_stage_opamp_dummy_magic_0.VOUT+.t115 GNDA 0.295144f
C2023 two_stage_opamp_dummy_magic_0.VOUT+.t131 GNDA 0.295764f
C2024 two_stage_opamp_dummy_magic_0.VOUT+.t104 GNDA 0.290811f
C2025 two_stage_opamp_dummy_magic_0.VOUT+.n44 GNDA 0.194979f
C2026 two_stage_opamp_dummy_magic_0.VOUT+.t73 GNDA 0.290811f
C2027 two_stage_opamp_dummy_magic_0.VOUT+.n45 GNDA 0.122686f
C2028 two_stage_opamp_dummy_magic_0.VOUT+.t146 GNDA 0.295144f
C2029 two_stage_opamp_dummy_magic_0.VOUT+.t31 GNDA 0.295764f
C2030 two_stage_opamp_dummy_magic_0.VOUT+.t138 GNDA 0.290811f
C2031 two_stage_opamp_dummy_magic_0.VOUT+.n46 GNDA 0.194979f
C2032 two_stage_opamp_dummy_magic_0.VOUT+.t107 GNDA 0.290811f
C2033 two_stage_opamp_dummy_magic_0.VOUT+.n47 GNDA 0.122686f
C2034 two_stage_opamp_dummy_magic_0.VOUT+.t46 GNDA 0.295144f
C2035 two_stage_opamp_dummy_magic_0.VOUT+.t62 GNDA 0.295764f
C2036 two_stage_opamp_dummy_magic_0.VOUT+.t41 GNDA 0.290811f
C2037 two_stage_opamp_dummy_magic_0.VOUT+.n48 GNDA 0.194979f
C2038 two_stage_opamp_dummy_magic_0.VOUT+.t143 GNDA 0.290811f
C2039 two_stage_opamp_dummy_magic_0.VOUT+.n49 GNDA 0.122686f
C2040 two_stage_opamp_dummy_magic_0.VOUT+.t87 GNDA 0.295144f
C2041 two_stage_opamp_dummy_magic_0.VOUT+.t114 GNDA 0.295764f
C2042 two_stage_opamp_dummy_magic_0.VOUT+.t21 GNDA 0.290811f
C2043 two_stage_opamp_dummy_magic_0.VOUT+.n50 GNDA 0.194979f
C2044 two_stage_opamp_dummy_magic_0.VOUT+.t126 GNDA 0.290811f
C2045 two_stage_opamp_dummy_magic_0.VOUT+.n51 GNDA 0.122686f
C2046 two_stage_opamp_dummy_magic_0.VOUT+.t65 GNDA 0.295144f
C2047 two_stage_opamp_dummy_magic_0.VOUT+.t26 GNDA 0.295387f
C2048 two_stage_opamp_dummy_magic_0.VOUT+.t102 GNDA 0.295144f
C2049 two_stage_opamp_dummy_magic_0.VOUT+.t59 GNDA 0.295387f
C2050 two_stage_opamp_dummy_magic_0.VOUT+.t134 GNDA 0.295144f
C2051 two_stage_opamp_dummy_magic_0.VOUT+.t37 GNDA 0.295387f
C2052 two_stage_opamp_dummy_magic_0.VOUT+.t120 GNDA 0.295144f
C2053 two_stage_opamp_dummy_magic_0.VOUT+.t81 GNDA 0.295387f
C2054 two_stage_opamp_dummy_magic_0.VOUT+.t155 GNDA 0.295144f
C2055 two_stage_opamp_dummy_magic_0.VOUT+.t119 GNDA 0.290811f
C2056 two_stage_opamp_dummy_magic_0.VOUT+.n52 GNDA 0.321888f
C2057 two_stage_opamp_dummy_magic_0.VOUT+.t82 GNDA 0.290811f
C2058 two_stage_opamp_dummy_magic_0.VOUT+.n53 GNDA 0.376415f
C2059 two_stage_opamp_dummy_magic_0.VOUT+.t97 GNDA 0.290811f
C2060 two_stage_opamp_dummy_magic_0.VOUT+.n54 GNDA 0.376415f
C2061 two_stage_opamp_dummy_magic_0.VOUT+.t63 GNDA 0.290811f
C2062 two_stage_opamp_dummy_magic_0.VOUT+.n55 GNDA 0.376415f
C2063 two_stage_opamp_dummy_magic_0.VOUT+.t27 GNDA 0.290811f
C2064 two_stage_opamp_dummy_magic_0.VOUT+.n56 GNDA 0.309197f
C2065 two_stage_opamp_dummy_magic_0.VOUT+.t45 GNDA 0.290811f
C2066 two_stage_opamp_dummy_magic_0.VOUT+.n57 GNDA 0.309197f
C2067 two_stage_opamp_dummy_magic_0.VOUT+.t144 GNDA 0.290811f
C2068 two_stage_opamp_dummy_magic_0.VOUT+.n58 GNDA 0.309197f
C2069 two_stage_opamp_dummy_magic_0.VOUT+.t112 GNDA 0.290811f
C2070 two_stage_opamp_dummy_magic_0.VOUT+.n59 GNDA 0.309197f
C2071 two_stage_opamp_dummy_magic_0.VOUT+.t76 GNDA 0.290811f
C2072 two_stage_opamp_dummy_magic_0.VOUT+.n60 GNDA 0.250126f
C2073 two_stage_opamp_dummy_magic_0.VOUT+.t93 GNDA 0.290811f
C2074 two_stage_opamp_dummy_magic_0.VOUT+.n61 GNDA 0.250126f
C2075 two_stage_opamp_dummy_magic_0.VOUT+.t56 GNDA 0.290811f
C2076 two_stage_opamp_dummy_magic_0.VOUT+.t40 GNDA 0.295764f
C2077 two_stage_opamp_dummy_magic_0.VOUT+.t19 GNDA 0.290811f
C2078 two_stage_opamp_dummy_magic_0.VOUT+.n62 GNDA 0.194979f
C2079 two_stage_opamp_dummy_magic_0.VOUT+.n63 GNDA 0.236284f
C2080 two_stage_opamp_dummy_magic_0.VOUT+.t34 GNDA 0.295764f
C2081 two_stage_opamp_dummy_magic_0.VOUT+.t52 GNDA 0.290811f
C2082 two_stage_opamp_dummy_magic_0.VOUT+.n64 GNDA 0.194979f
C2083 two_stage_opamp_dummy_magic_0.VOUT+.t156 GNDA 0.290811f
C2084 two_stage_opamp_dummy_magic_0.VOUT+.t136 GNDA 0.295764f
C2085 two_stage_opamp_dummy_magic_0.VOUT+.t121 GNDA 0.290811f
C2086 two_stage_opamp_dummy_magic_0.VOUT+.n65 GNDA 0.194979f
C2087 two_stage_opamp_dummy_magic_0.VOUT+.n66 GNDA 0.236284f
C2088 two_stage_opamp_dummy_magic_0.VOUT+.t70 GNDA 0.295764f
C2089 two_stage_opamp_dummy_magic_0.VOUT+.t89 GNDA 0.290811f
C2090 two_stage_opamp_dummy_magic_0.VOUT+.n67 GNDA 0.194979f
C2091 two_stage_opamp_dummy_magic_0.VOUT+.t50 GNDA 0.290811f
C2092 two_stage_opamp_dummy_magic_0.VOUT+.t36 GNDA 0.295764f
C2093 two_stage_opamp_dummy_magic_0.VOUT+.t151 GNDA 0.290811f
C2094 two_stage_opamp_dummy_magic_0.VOUT+.n68 GNDA 0.194979f
C2095 two_stage_opamp_dummy_magic_0.VOUT+.n69 GNDA 0.236284f
C2096 two_stage_opamp_dummy_magic_0.VOUT+.t95 GNDA 0.295764f
C2097 two_stage_opamp_dummy_magic_0.VOUT+.t43 GNDA 0.290811f
C2098 two_stage_opamp_dummy_magic_0.VOUT+.n70 GNDA 0.194979f
C2099 two_stage_opamp_dummy_magic_0.VOUT+.t145 GNDA 0.290811f
C2100 two_stage_opamp_dummy_magic_0.VOUT+.t66 GNDA 0.295764f
C2101 two_stage_opamp_dummy_magic_0.VOUT+.t118 GNDA 0.290811f
C2102 two_stage_opamp_dummy_magic_0.VOUT+.n71 GNDA 0.194979f
C2103 two_stage_opamp_dummy_magic_0.VOUT+.n72 GNDA 0.236284f
C2104 two_stage_opamp_dummy_magic_0.VOUT+.t55 GNDA 0.295764f
C2105 two_stage_opamp_dummy_magic_0.VOUT+.t141 GNDA 0.290811f
C2106 two_stage_opamp_dummy_magic_0.VOUT+.n73 GNDA 0.194979f
C2107 two_stage_opamp_dummy_magic_0.VOUT+.t111 GNDA 0.290811f
C2108 two_stage_opamp_dummy_magic_0.VOUT+.t29 GNDA 0.295764f
C2109 two_stage_opamp_dummy_magic_0.VOUT+.t80 GNDA 0.290811f
C2110 two_stage_opamp_dummy_magic_0.VOUT+.n74 GNDA 0.194979f
C2111 two_stage_opamp_dummy_magic_0.VOUT+.n75 GNDA 0.236284f
C2112 two_stage_opamp_dummy_magic_0.VOUT+.t91 GNDA 0.295764f
C2113 two_stage_opamp_dummy_magic_0.VOUT+.t39 GNDA 0.290811f
C2114 two_stage_opamp_dummy_magic_0.VOUT+.n76 GNDA 0.194979f
C2115 two_stage_opamp_dummy_magic_0.VOUT+.t139 GNDA 0.290811f
C2116 two_stage_opamp_dummy_magic_0.VOUT+.t58 GNDA 0.295764f
C2117 two_stage_opamp_dummy_magic_0.VOUT+.t109 GNDA 0.290811f
C2118 two_stage_opamp_dummy_magic_0.VOUT+.n77 GNDA 0.194979f
C2119 two_stage_opamp_dummy_magic_0.VOUT+.n78 GNDA 0.236284f
C2120 two_stage_opamp_dummy_magic_0.VOUT+.t49 GNDA 0.295764f
C2121 two_stage_opamp_dummy_magic_0.VOUT+.t135 GNDA 0.290811f
C2122 two_stage_opamp_dummy_magic_0.VOUT+.n79 GNDA 0.194979f
C2123 two_stage_opamp_dummy_magic_0.VOUT+.t103 GNDA 0.290811f
C2124 two_stage_opamp_dummy_magic_0.VOUT+.t20 GNDA 0.295764f
C2125 two_stage_opamp_dummy_magic_0.VOUT+.t72 GNDA 0.290811f
C2126 two_stage_opamp_dummy_magic_0.VOUT+.n80 GNDA 0.194979f
C2127 two_stage_opamp_dummy_magic_0.VOUT+.n81 GNDA 0.236284f
C2128 two_stage_opamp_dummy_magic_0.VOUT+.t148 GNDA 0.295764f
C2129 two_stage_opamp_dummy_magic_0.VOUT+.t99 GNDA 0.290811f
C2130 two_stage_opamp_dummy_magic_0.VOUT+.n82 GNDA 0.194979f
C2131 two_stage_opamp_dummy_magic_0.VOUT+.t68 GNDA 0.290811f
C2132 two_stage_opamp_dummy_magic_0.VOUT+.t122 GNDA 0.295764f
C2133 two_stage_opamp_dummy_magic_0.VOUT+.t33 GNDA 0.290811f
C2134 two_stage_opamp_dummy_magic_0.VOUT+.n83 GNDA 0.194979f
C2135 two_stage_opamp_dummy_magic_0.VOUT+.n84 GNDA 0.236284f
C2136 two_stage_opamp_dummy_magic_0.VOUT+.t44 GNDA 0.295764f
C2137 two_stage_opamp_dummy_magic_0.VOUT+.t133 GNDA 0.290811f
C2138 two_stage_opamp_dummy_magic_0.VOUT+.n85 GNDA 0.194979f
C2139 two_stage_opamp_dummy_magic_0.VOUT+.t98 GNDA 0.290811f
C2140 two_stage_opamp_dummy_magic_0.VOUT+.t152 GNDA 0.295764f
C2141 two_stage_opamp_dummy_magic_0.VOUT+.t67 GNDA 0.290811f
C2142 two_stage_opamp_dummy_magic_0.VOUT+.n86 GNDA 0.194979f
C2143 two_stage_opamp_dummy_magic_0.VOUT+.n87 GNDA 0.236284f
C2144 two_stage_opamp_dummy_magic_0.VOUT+.t142 GNDA 0.295764f
C2145 two_stage_opamp_dummy_magic_0.VOUT+.t94 GNDA 0.290811f
C2146 two_stage_opamp_dummy_magic_0.VOUT+.n88 GNDA 0.194979f
C2147 two_stage_opamp_dummy_magic_0.VOUT+.t60 GNDA 0.290811f
C2148 two_stage_opamp_dummy_magic_0.VOUT+.t116 GNDA 0.295764f
C2149 two_stage_opamp_dummy_magic_0.VOUT+.t30 GNDA 0.290811f
C2150 two_stage_opamp_dummy_magic_0.VOUT+.n89 GNDA 0.194979f
C2151 two_stage_opamp_dummy_magic_0.VOUT+.n90 GNDA 0.236284f
C2152 two_stage_opamp_dummy_magic_0.VOUT+.t77 GNDA 0.295764f
C2153 two_stage_opamp_dummy_magic_0.VOUT+.t127 GNDA 0.290811f
C2154 two_stage_opamp_dummy_magic_0.VOUT+.n91 GNDA 0.194979f
C2155 two_stage_opamp_dummy_magic_0.VOUT+.t22 GNDA 0.290811f
C2156 two_stage_opamp_dummy_magic_0.VOUT+.n92 GNDA 0.236284f
C2157 two_stage_opamp_dummy_magic_0.VOUT+.t53 GNDA 0.290811f
C2158 two_stage_opamp_dummy_magic_0.VOUT+.n93 GNDA 0.12723f
C2159 two_stage_opamp_dummy_magic_0.VOUT+.t105 GNDA 0.290811f
C2160 two_stage_opamp_dummy_magic_0.VOUT+.n94 GNDA 0.23826f
C2161 two_stage_opamp_dummy_magic_0.VOUT+.n95 GNDA 0.300935f
C2162 two_stage_opamp_dummy_magic_0.VOUT+.n96 GNDA 0.170241f
C2163 two_stage_opamp_dummy_magic_0.VOUT+.t17 GNDA 0.084142f
C2164 two_stage_opamp_dummy_magic_0.VD2.t12 GNDA 0.013877f
C2165 two_stage_opamp_dummy_magic_0.VD2.t4 GNDA 0.013877f
C2166 two_stage_opamp_dummy_magic_0.VD2.t18 GNDA 0.013877f
C2167 two_stage_opamp_dummy_magic_0.VD2.n0 GNDA 0.048872f
C2168 two_stage_opamp_dummy_magic_0.VD2.t6 GNDA 0.013877f
C2169 two_stage_opamp_dummy_magic_0.VD2.t2 GNDA 0.013877f
C2170 two_stage_opamp_dummy_magic_0.VD2.n1 GNDA 0.047884f
C2171 two_stage_opamp_dummy_magic_0.VD2.n2 GNDA 0.193373f
C2172 two_stage_opamp_dummy_magic_0.VD2.t7 GNDA 0.013877f
C2173 two_stage_opamp_dummy_magic_0.VD2.t16 GNDA 0.013877f
C2174 two_stage_opamp_dummy_magic_0.VD2.n3 GNDA 0.047884f
C2175 two_stage_opamp_dummy_magic_0.VD2.n4 GNDA 0.140662f
C2176 two_stage_opamp_dummy_magic_0.VD2.t20 GNDA 0.013877f
C2177 two_stage_opamp_dummy_magic_0.VD2.t21 GNDA 0.013877f
C2178 two_stage_opamp_dummy_magic_0.VD2.n5 GNDA 0.04687f
C2179 two_stage_opamp_dummy_magic_0.VD2.t3 GNDA 0.013877f
C2180 two_stage_opamp_dummy_magic_0.VD2.t1 GNDA 0.013877f
C2181 two_stage_opamp_dummy_magic_0.VD2.n6 GNDA 0.050131f
C2182 two_stage_opamp_dummy_magic_0.VD2.t9 GNDA 0.013877f
C2183 two_stage_opamp_dummy_magic_0.VD2.t14 GNDA 0.013877f
C2184 two_stage_opamp_dummy_magic_0.VD2.n7 GNDA 0.050131f
C2185 two_stage_opamp_dummy_magic_0.VD2.t8 GNDA 0.013877f
C2186 two_stage_opamp_dummy_magic_0.VD2.t5 GNDA 0.013877f
C2187 two_stage_opamp_dummy_magic_0.VD2.n8 GNDA 0.04969f
C2188 two_stage_opamp_dummy_magic_0.VD2.n9 GNDA 0.186051f
C2189 two_stage_opamp_dummy_magic_0.VD2.t11 GNDA 0.013877f
C2190 two_stage_opamp_dummy_magic_0.VD2.t10 GNDA 0.013877f
C2191 two_stage_opamp_dummy_magic_0.VD2.n10 GNDA 0.04969f
C2192 two_stage_opamp_dummy_magic_0.VD2.n11 GNDA 0.096484f
C2193 two_stage_opamp_dummy_magic_0.VD2.n12 GNDA 0.117322f
C2194 two_stage_opamp_dummy_magic_0.VD2.n13 GNDA 0.081264f
C2195 two_stage_opamp_dummy_magic_0.VD2.t0 GNDA 0.013877f
C2196 two_stage_opamp_dummy_magic_0.VD2.t15 GNDA 0.013877f
C2197 two_stage_opamp_dummy_magic_0.VD2.n14 GNDA 0.045463f
C2198 two_stage_opamp_dummy_magic_0.VD2.n15 GNDA 0.069533f
C2199 two_stage_opamp_dummy_magic_0.VD2.n16 GNDA 0.083264f
C2200 two_stage_opamp_dummy_magic_0.VD2.t13 GNDA 0.013877f
C2201 two_stage_opamp_dummy_magic_0.VD2.t19 GNDA 0.013877f
C2202 two_stage_opamp_dummy_magic_0.VD2.n17 GNDA 0.047884f
C2203 two_stage_opamp_dummy_magic_0.VD2.n18 GNDA 0.193373f
C2204 two_stage_opamp_dummy_magic_0.VD2.n19 GNDA 0.048872f
C2205 two_stage_opamp_dummy_magic_0.VD2.t17 GNDA 0.013877f
C2206 bgr_0.cap_res1.t7 GNDA 0.417173f
C2207 bgr_0.cap_res1.t11 GNDA 0.418684f
C2208 bgr_0.cap_res1.t1 GNDA 0.417173f
C2209 bgr_0.cap_res1.t15 GNDA 0.418684f
C2210 bgr_0.cap_res1.t4 GNDA 0.417173f
C2211 bgr_0.cap_res1.t8 GNDA 0.418684f
C2212 bgr_0.cap_res1.t16 GNDA 0.417173f
C2213 bgr_0.cap_res1.t10 GNDA 0.418684f
C2214 bgr_0.cap_res1.t9 GNDA 0.417173f
C2215 bgr_0.cap_res1.t13 GNDA 0.418684f
C2216 bgr_0.cap_res1.t2 GNDA 0.417173f
C2217 bgr_0.cap_res1.t17 GNDA 0.418684f
C2218 bgr_0.cap_res1.t14 GNDA 0.417173f
C2219 bgr_0.cap_res1.t20 GNDA 0.418684f
C2220 bgr_0.cap_res1.t6 GNDA 0.417173f
C2221 bgr_0.cap_res1.t3 GNDA 0.418684f
C2222 bgr_0.cap_res1.n0 GNDA 0.279631f
C2223 bgr_0.cap_res1.t5 GNDA 0.222685f
C2224 bgr_0.cap_res1.n1 GNDA 0.303406f
C2225 bgr_0.cap_res1.t19 GNDA 0.222685f
C2226 bgr_0.cap_res1.n2 GNDA 0.303406f
C2227 bgr_0.cap_res1.t12 GNDA 0.222685f
C2228 bgr_0.cap_res1.n3 GNDA 0.303406f
C2229 bgr_0.cap_res1.t18 GNDA 0.649059f
C2230 bgr_0.cap_res1.t0 GNDA 0.10618f
C2231 bgr_0.1st_Vout_1.n0 GNDA 0.573726f
C2232 bgr_0.1st_Vout_1.n1 GNDA 1.42916f
C2233 bgr_0.1st_Vout_1.n2 GNDA 1.78489f
C2234 bgr_0.1st_Vout_1.n3 GNDA 0.125562f
C2235 bgr_0.1st_Vout_1.t20 GNDA 0.352846f
C2236 bgr_0.1st_Vout_1.t11 GNDA 0.346937f
C2237 bgr_0.1st_Vout_1.t32 GNDA 0.346937f
C2238 bgr_0.1st_Vout_1.t29 GNDA 0.352846f
C2239 bgr_0.1st_Vout_1.t34 GNDA 0.346937f
C2240 bgr_0.1st_Vout_1.t25 GNDA 0.352846f
C2241 bgr_0.1st_Vout_1.t21 GNDA 0.346937f
C2242 bgr_0.1st_Vout_1.t12 GNDA 0.346937f
C2243 bgr_0.1st_Vout_1.t35 GNDA 0.352846f
C2244 bgr_0.1st_Vout_1.t16 GNDA 0.346937f
C2245 bgr_0.1st_Vout_1.t33 GNDA 0.352846f
C2246 bgr_0.1st_Vout_1.t26 GNDA 0.346937f
C2247 bgr_0.1st_Vout_1.t22 GNDA 0.346937f
C2248 bgr_0.1st_Vout_1.t17 GNDA 0.352846f
C2249 bgr_0.1st_Vout_1.t24 GNDA 0.346937f
C2250 bgr_0.1st_Vout_1.t28 GNDA 0.352846f
C2251 bgr_0.1st_Vout_1.t23 GNDA 0.346937f
C2252 bgr_0.1st_Vout_1.t13 GNDA 0.346937f
C2253 bgr_0.1st_Vout_1.t18 GNDA 0.346937f
C2254 bgr_0.1st_Vout_1.t36 GNDA 0.346937f
C2255 bgr_0.1st_Vout_1.t30 GNDA 0.022665f
C2256 bgr_0.1st_Vout_1.n4 GNDA 0.021864f
C2257 bgr_0.1st_Vout_1.t14 GNDA 0.013213f
C2258 bgr_0.1st_Vout_1.t31 GNDA 0.013213f
C2259 bgr_0.1st_Vout_1.n5 GNDA 0.029393f
C2260 bgr_0.1st_Vout_1.t2 GNDA 0.018268f
C2261 bgr_0.1st_Vout_1.n6 GNDA 0.012529f
C2262 bgr_0.1st_Vout_1.n7 GNDA 0.189508f
C2263 bgr_0.1st_Vout_1.n8 GNDA 0.011336f
C2264 bgr_0.1st_Vout_1.n9 GNDA 0.020958f
C2265 bgr_0.1st_Vout_1.t19 GNDA 0.013213f
C2266 bgr_0.1st_Vout_1.t27 GNDA 0.013213f
C2267 bgr_0.1st_Vout_1.n10 GNDA 0.029393f
C2268 bgr_0.1st_Vout_1.n11 GNDA 0.021864f
C2269 bgr_0.1st_Vout_1.t15 GNDA 0.020738f
C2270 VDDA.t137 GNDA 0.020556f
C2271 VDDA.t34 GNDA 0.020556f
C2272 VDDA.n0 GNDA 0.085011f
C2273 VDDA.t212 GNDA 0.020556f
C2274 VDDA.t190 GNDA 0.020556f
C2275 VDDA.n1 GNDA 0.084685f
C2276 VDDA.n2 GNDA 0.117411f
C2277 VDDA.t118 GNDA 0.020556f
C2278 VDDA.t124 GNDA 0.020556f
C2279 VDDA.n3 GNDA 0.084685f
C2280 VDDA.n4 GNDA 0.061267f
C2281 VDDA.t254 GNDA 0.020556f
C2282 VDDA.t53 GNDA 0.020556f
C2283 VDDA.n5 GNDA 0.084685f
C2284 VDDA.n6 GNDA 0.061267f
C2285 VDDA.t15 GNDA 0.020556f
C2286 VDDA.t188 GNDA 0.020556f
C2287 VDDA.n7 GNDA 0.084685f
C2288 VDDA.n8 GNDA 0.061267f
C2289 VDDA.t232 GNDA 0.020556f
C2290 VDDA.t191 GNDA 0.020556f
C2291 VDDA.n9 GNDA 0.084685f
C2292 VDDA.n10 GNDA 0.145592f
C2293 VDDA.n11 GNDA 0.06638f
C2294 VDDA.n12 GNDA 0.177216f
C2295 VDDA.t321 GNDA 0.012911f
C2296 VDDA.n13 GNDA 0.027472f
C2297 VDDA.t430 GNDA 0.012911f
C2298 VDDA.n14 GNDA 0.027472f
C2299 VDDA.n15 GNDA 0.039889f
C2300 VDDA.n16 GNDA 0.067046f
C2301 VDDA.n17 GNDA 0.178679f
C2302 VDDA.t391 GNDA 0.012911f
C2303 VDDA.n18 GNDA 0.027472f
C2304 VDDA.t364 GNDA 0.012911f
C2305 VDDA.n19 GNDA 0.027472f
C2306 VDDA.n20 GNDA 0.037173f
C2307 VDDA.n21 GNDA 0.046144f
C2308 VDDA.n22 GNDA 0.178679f
C2309 VDDA.t363 GNDA 0.17382f
C2310 VDDA.t263 GNDA 0.107408f
C2311 VDDA.t48 GNDA 0.107408f
C2312 VDDA.t59 GNDA 0.107408f
C2313 VDDA.t86 GNDA 0.107408f
C2314 VDDA.t253 GNDA 0.080556f
C2315 VDDA.t390 GNDA 0.17382f
C2316 VDDA.t43 GNDA 0.107408f
C2317 VDDA.t250 GNDA 0.107408f
C2318 VDDA.t87 GNDA 0.107408f
C2319 VDDA.t45 GNDA 0.107408f
C2320 VDDA.t68 GNDA 0.080556f
C2321 VDDA.n23 GNDA 0.067711f
C2322 VDDA.n24 GNDA 0.053704f
C2323 VDDA.n25 GNDA 0.067711f
C2324 VDDA.n26 GNDA 0.045224f
C2325 VDDA.n27 GNDA 0.036591f
C2326 VDDA.n28 GNDA 0.085078f
C2327 VDDA.n29 GNDA 0.085078f
C2328 VDDA.n30 GNDA 0.177216f
C2329 VDDA.t429 GNDA 0.170315f
C2330 VDDA.t249 GNDA 0.105523f
C2331 VDDA.t27 GNDA 0.105523f
C2332 VDDA.t150 GNDA 0.105523f
C2333 VDDA.t251 GNDA 0.105523f
C2334 VDDA.t262 GNDA 0.079143f
C2335 VDDA.t320 GNDA 0.170315f
C2336 VDDA.t103 GNDA 0.105523f
C2337 VDDA.t248 GNDA 0.105523f
C2338 VDDA.t252 GNDA 0.105523f
C2339 VDDA.t257 GNDA 0.105523f
C2340 VDDA.t443 GNDA 0.079143f
C2341 VDDA.n31 GNDA 0.067711f
C2342 VDDA.n32 GNDA 0.052762f
C2343 VDDA.n33 GNDA 0.067711f
C2344 VDDA.n34 GNDA 0.045009f
C2345 VDDA.n35 GNDA 0.036591f
C2346 VDDA.n36 GNDA 0.070836f
C2347 VDDA.n37 GNDA 0.210513f
C2348 VDDA.t123 GNDA 0.041113f
C2349 VDDA.t211 GNDA 0.041113f
C2350 VDDA.n38 GNDA 0.16494f
C2351 VDDA.n39 GNDA 0.083794f
C2352 VDDA.t327 GNDA 0.040956f
C2353 VDDA.n40 GNDA 0.083113f
C2354 VDDA.n41 GNDA 0.055457f
C2355 VDDA.n42 GNDA 0.078279f
C2356 VDDA.t367 GNDA 0.045486f
C2357 VDDA.t365 GNDA 0.019919f
C2358 VDDA.n43 GNDA 0.072153f
C2359 VDDA.n44 GNDA 0.042476f
C2360 VDDA.t333 GNDA 0.045486f
C2361 VDDA.t331 GNDA 0.019919f
C2362 VDDA.n45 GNDA 0.072153f
C2363 VDDA.n46 GNDA 0.042476f
C2364 VDDA.n47 GNDA 0.045224f
C2365 VDDA.n48 GNDA 0.078279f
C2366 VDDA.n49 GNDA 0.226295f
C2367 VDDA.t332 GNDA 0.28026f
C2368 VDDA.t10 GNDA 0.162054f
C2369 VDDA.t209 GNDA 0.162054f
C2370 VDDA.t119 GNDA 0.162054f
C2371 VDDA.t55 GNDA 0.162054f
C2372 VDDA.t125 GNDA 0.12154f
C2373 VDDA.n50 GNDA 0.081027f
C2374 VDDA.t189 GNDA 0.12154f
C2375 VDDA.t21 GNDA 0.162054f
C2376 VDDA.t187 GNDA 0.162054f
C2377 VDDA.t54 GNDA 0.162054f
C2378 VDDA.t255 GNDA 0.162054f
C2379 VDDA.t366 GNDA 0.28026f
C2380 VDDA.n51 GNDA 0.226295f
C2381 VDDA.n52 GNDA 0.055457f
C2382 VDDA.n53 GNDA 0.104943f
C2383 VDDA.t355 GNDA 0.040956f
C2384 VDDA.t121 GNDA 0.041113f
C2385 VDDA.t14 GNDA 0.041113f
C2386 VDDA.n54 GNDA 0.16494f
C2387 VDDA.n55 GNDA 0.083794f
C2388 VDDA.t20 GNDA 0.041113f
C2389 VDDA.t186 GNDA 0.041113f
C2390 VDDA.n56 GNDA 0.16494f
C2391 VDDA.n57 GNDA 0.083794f
C2392 VDDA.t139 GNDA 0.041113f
C2393 VDDA.t117 GNDA 0.041113f
C2394 VDDA.n58 GNDA 0.16494f
C2395 VDDA.n59 GNDA 0.083794f
C2396 VDDA.t12 GNDA 0.041113f
C2397 VDDA.t127 GNDA 0.041113f
C2398 VDDA.n60 GNDA 0.16494f
C2399 VDDA.n61 GNDA 0.17608f
C2400 VDDA.n62 GNDA 0.132944f
C2401 VDDA.t353 GNDA 0.049694f
C2402 VDDA.n63 GNDA 0.095079f
C2403 VDDA.n64 GNDA 0.055548f
C2404 VDDA.n65 GNDA 0.365831f
C2405 VDDA.n66 GNDA 0.365831f
C2406 VDDA.t326 GNDA 0.565063f
C2407 VDDA.t122 GNDA 0.312802f
C2408 VDDA.t210 GNDA 0.312802f
C2409 VDDA.t120 GNDA 0.312802f
C2410 VDDA.t13 GNDA 0.312802f
C2411 VDDA.t19 GNDA 0.234601f
C2412 VDDA.n67 GNDA 0.083113f
C2413 VDDA.n68 GNDA 0.106529f
C2414 VDDA.n69 GNDA 0.106529f
C2415 VDDA.t354 GNDA 0.565063f
C2416 VDDA.t126 GNDA 0.312802f
C2417 VDDA.t11 GNDA 0.312802f
C2418 VDDA.t116 GNDA 0.312802f
C2419 VDDA.t138 GNDA 0.312802f
C2420 VDDA.t185 GNDA 0.234601f
C2421 VDDA.n70 GNDA 0.156401f
C2422 VDDA.n71 GNDA 0.105835f
C2423 VDDA.n72 GNDA 0.071819f
C2424 VDDA.n73 GNDA 0.055548f
C2425 VDDA.t325 GNDA 0.049694f
C2426 VDDA.n74 GNDA 0.095079f
C2427 VDDA.n75 GNDA 0.132601f
C2428 VDDA.n76 GNDA 0.117983f
C2429 VDDA.n77 GNDA 0.100384f
C2430 VDDA.t237 GNDA 0.023983f
C2431 VDDA.t136 GNDA 0.023983f
C2432 VDDA.n78 GNDA 0.083406f
C2433 VDDA.t33 GNDA 0.023983f
C2434 VDDA.t111 GNDA 0.023983f
C2435 VDDA.n79 GNDA 0.083111f
C2436 VDDA.n80 GNDA 0.156905f
C2437 VDDA.t208 GNDA 0.023983f
C2438 VDDA.t70 GNDA 0.023983f
C2439 VDDA.n81 GNDA 0.083406f
C2440 VDDA.t206 GNDA 0.023983f
C2441 VDDA.t259 GNDA 0.023983f
C2442 VDDA.n82 GNDA 0.083111f
C2443 VDDA.n83 GNDA 0.156905f
C2444 VDDA.n84 GNDA 0.021927f
C2445 VDDA.n85 GNDA 0.068276f
C2446 VDDA.n86 GNDA 0.092842f
C2447 VDDA.t421 GNDA 0.118311f
C2448 VDDA.t419 GNDA 0.041762f
C2449 VDDA.n87 GNDA 0.077183f
C2450 VDDA.n88 GNDA 0.049756f
C2451 VDDA.t376 GNDA 0.118311f
C2452 VDDA.t374 GNDA 0.041762f
C2453 VDDA.n89 GNDA 0.077183f
C2454 VDDA.n90 GNDA 0.049756f
C2455 VDDA.n91 GNDA 0.049336f
C2456 VDDA.n92 GNDA 0.092842f
C2457 VDDA.n93 GNDA 0.276684f
C2458 VDDA.t375 GNDA 0.412992f
C2459 VDDA.t236 GNDA 0.238456f
C2460 VDDA.t135 GNDA 0.238456f
C2461 VDDA.t32 GNDA 0.238456f
C2462 VDDA.t110 GNDA 0.238456f
C2463 VDDA.t449 GNDA 0.178842f
C2464 VDDA.n94 GNDA 0.119228f
C2465 VDDA.t172 GNDA 0.178842f
C2466 VDDA.t205 GNDA 0.238456f
C2467 VDDA.t258 GNDA 0.238456f
C2468 VDDA.t207 GNDA 0.238456f
C2469 VDDA.t69 GNDA 0.238456f
C2470 VDDA.t420 GNDA 0.412992f
C2471 VDDA.n95 GNDA 0.276684f
C2472 VDDA.n96 GNDA 0.068276f
C2473 VDDA.n97 GNDA 0.095583f
C2474 VDDA.t450 GNDA 0.023983f
C2475 VDDA.t173 GNDA 0.023983f
C2476 VDDA.n98 GNDA 0.078193f
C2477 VDDA.n99 GNDA 0.053368f
C2478 VDDA.n100 GNDA 0.044833f
C2479 VDDA.t35 GNDA 0.020556f
C2480 VDDA.t183 GNDA 0.020556f
C2481 VDDA.n101 GNDA 0.085011f
C2482 VDDA.t44 GNDA 0.020556f
C2483 VDDA.t169 GNDA 0.020556f
C2484 VDDA.n102 GNDA 0.084685f
C2485 VDDA.n103 GNDA 0.117411f
C2486 VDDA.t130 GNDA 0.020556f
C2487 VDDA.t18 GNDA 0.020556f
C2488 VDDA.n104 GNDA 0.084685f
C2489 VDDA.n105 GNDA 0.061267f
C2490 VDDA.t58 GNDA 0.020556f
C2491 VDDA.t256 GNDA 0.020556f
C2492 VDDA.n106 GNDA 0.084685f
C2493 VDDA.n107 GNDA 0.061267f
C2494 VDDA.t102 GNDA 0.020556f
C2495 VDDA.t192 GNDA 0.020556f
C2496 VDDA.n108 GNDA 0.084685f
C2497 VDDA.n109 GNDA 0.061267f
C2498 VDDA.t83 GNDA 0.020556f
C2499 VDDA.t112 GNDA 0.020556f
C2500 VDDA.n110 GNDA 0.084685f
C2501 VDDA.n111 GNDA 0.176944f
C2502 VDDA.t85 GNDA 0.041113f
C2503 VDDA.t115 GNDA 0.041113f
C2504 VDDA.n112 GNDA 0.16494f
C2505 VDDA.n113 GNDA 0.083794f
C2506 VDDA.t382 GNDA 0.040956f
C2507 VDDA.n114 GNDA 0.055457f
C2508 VDDA.n115 GNDA 0.078279f
C2509 VDDA.t388 GNDA 0.045486f
C2510 VDDA.t386 GNDA 0.019919f
C2511 VDDA.n116 GNDA 0.072153f
C2512 VDDA.n117 GNDA 0.042476f
C2513 VDDA.t361 GNDA 0.045486f
C2514 VDDA.t359 GNDA 0.019919f
C2515 VDDA.n118 GNDA 0.072153f
C2516 VDDA.n119 GNDA 0.042476f
C2517 VDDA.n120 GNDA 0.045224f
C2518 VDDA.n121 GNDA 0.078279f
C2519 VDDA.n122 GNDA 0.226295f
C2520 VDDA.t360 GNDA 0.28026f
C2521 VDDA.t182 GNDA 0.162054f
C2522 VDDA.t444 GNDA 0.162054f
C2523 VDDA.t221 GNDA 0.162054f
C2524 VDDA.t456 GNDA 0.162054f
C2525 VDDA.t113 GNDA 0.12154f
C2526 VDDA.n123 GNDA 0.081027f
C2527 VDDA.t57 GNDA 0.12154f
C2528 VDDA.t184 GNDA 0.162054f
C2529 VDDA.t56 GNDA 0.162054f
C2530 VDDA.t233 GNDA 0.162054f
C2531 VDDA.t26 GNDA 0.162054f
C2532 VDDA.t387 GNDA 0.28026f
C2533 VDDA.n124 GNDA 0.226295f
C2534 VDDA.n125 GNDA 0.055457f
C2535 VDDA.n126 GNDA 0.104943f
C2536 VDDA.n127 GNDA 0.071819f
C2537 VDDA.n128 GNDA 0.106529f
C2538 VDDA.n129 GNDA 0.106529f
C2539 VDDA.n130 GNDA 0.105835f
C2540 VDDA.t349 GNDA 0.040956f
C2541 VDDA.t17 GNDA 0.041113f
C2542 VDDA.t47 GNDA 0.041113f
C2543 VDDA.n131 GNDA 0.16494f
C2544 VDDA.n132 GNDA 0.083794f
C2545 VDDA.t129 GNDA 0.041113f
C2546 VDDA.t42 GNDA 0.041113f
C2547 VDDA.n133 GNDA 0.16494f
C2548 VDDA.n134 GNDA 0.083794f
C2549 VDDA.t223 GNDA 0.041113f
C2550 VDDA.t194 GNDA 0.041113f
C2551 VDDA.n135 GNDA 0.16494f
C2552 VDDA.n136 GNDA 0.083794f
C2553 VDDA.t171 GNDA 0.041113f
C2554 VDDA.t74 GNDA 0.041113f
C2555 VDDA.n137 GNDA 0.16494f
C2556 VDDA.n138 GNDA 0.17608f
C2557 VDDA.n139 GNDA 0.132944f
C2558 VDDA.t347 GNDA 0.049694f
C2559 VDDA.n140 GNDA 0.095079f
C2560 VDDA.n141 GNDA 0.055548f
C2561 VDDA.n142 GNDA 0.083113f
C2562 VDDA.n143 GNDA 0.365831f
C2563 VDDA.t348 GNDA 0.565063f
C2564 VDDA.t170 GNDA 0.312802f
C2565 VDDA.t73 GNDA 0.312802f
C2566 VDDA.t222 GNDA 0.312802f
C2567 VDDA.t193 GNDA 0.312802f
C2568 VDDA.t128 GNDA 0.234601f
C2569 VDDA.n144 GNDA 0.156401f
C2570 VDDA.t41 GNDA 0.234601f
C2571 VDDA.t16 GNDA 0.312802f
C2572 VDDA.t46 GNDA 0.312802f
C2573 VDDA.t84 GNDA 0.312802f
C2574 VDDA.t114 GNDA 0.312802f
C2575 VDDA.t381 GNDA 0.565063f
C2576 VDDA.n145 GNDA 0.365831f
C2577 VDDA.n146 GNDA 0.083113f
C2578 VDDA.n147 GNDA 0.055548f
C2579 VDDA.t380 GNDA 0.049694f
C2580 VDDA.n148 GNDA 0.095079f
C2581 VDDA.n149 GNDA 0.132601f
C2582 VDDA.n150 GNDA 0.101538f
C2583 VDDA.n152 GNDA 0.052465f
C2584 VDDA.n153 GNDA 0.065088f
C2585 VDDA.n155 GNDA 0.052465f
C2586 VDDA.n157 GNDA 0.052465f
C2587 VDDA.n159 GNDA 0.052465f
C2588 VDDA.n161 GNDA 0.052465f
C2589 VDDA.n163 GNDA 0.052465f
C2590 VDDA.n165 GNDA 0.052465f
C2591 VDDA.n167 GNDA 0.052465f
C2592 VDDA.n169 GNDA 0.052465f
C2593 VDDA.n171 GNDA 0.085855f
C2594 VDDA.t406 GNDA 0.012484f
C2595 VDDA.n172 GNDA 0.018537f
C2596 VDDA.n173 GNDA 0.016401f
C2597 VDDA.n174 GNDA 0.056016f
C2598 VDDA.n175 GNDA 0.215104f
C2599 VDDA.n176 GNDA 0.215104f
C2600 VDDA.t411 GNDA 0.170315f
C2601 VDDA.t153 GNDA 0.105523f
C2602 VDDA.t165 GNDA 0.105523f
C2603 VDDA.t161 GNDA 0.105523f
C2604 VDDA.t94 GNDA 0.105523f
C2605 VDDA.t148 GNDA 0.105523f
C2606 VDDA.t155 GNDA 0.105523f
C2607 VDDA.t90 GNDA 0.105523f
C2608 VDDA.t96 GNDA 0.105523f
C2609 VDDA.t66 GNDA 0.105523f
C2610 VDDA.t151 GNDA 0.079143f
C2611 VDDA.t405 GNDA 0.170315f
C2612 VDDA.t24 GNDA 0.105523f
C2613 VDDA.t163 GNDA 0.105523f
C2614 VDDA.t64 GNDA 0.105523f
C2615 VDDA.t157 GNDA 0.105523f
C2616 VDDA.t88 GNDA 0.105523f
C2617 VDDA.t167 GNDA 0.105523f
C2618 VDDA.t146 GNDA 0.105523f
C2619 VDDA.t22 GNDA 0.105523f
C2620 VDDA.t98 GNDA 0.105523f
C2621 VDDA.t92 GNDA 0.079143f
C2622 VDDA.n177 GNDA 0.065088f
C2623 VDDA.n178 GNDA 0.105196f
C2624 VDDA.n179 GNDA 0.105196f
C2625 VDDA.n180 GNDA 0.052762f
C2626 VDDA.n181 GNDA 0.105196f
C2627 VDDA.n182 GNDA 0.082911f
C2628 VDDA.n183 GNDA 0.056016f
C2629 VDDA.n184 GNDA 0.016401f
C2630 VDDA.t412 GNDA 0.012484f
C2631 VDDA.n185 GNDA 0.018084f
C2632 VDDA.n186 GNDA 0.064677f
C2633 VDDA.n187 GNDA 0.050706f
C2634 VDDA.n188 GNDA 0.261552f
C2635 VDDA.n189 GNDA 0.248765f
C2636 VDDA.t235 GNDA 0.023983f
C2637 VDDA.t1 GNDA 0.023983f
C2638 VDDA.n190 GNDA 0.083406f
C2639 VDDA.t231 GNDA 0.023983f
C2640 VDDA.t9 GNDA 0.023983f
C2641 VDDA.n191 GNDA 0.083111f
C2642 VDDA.n192 GNDA 0.156905f
C2643 VDDA.t40 GNDA 0.023983f
C2644 VDDA.t229 GNDA 0.023983f
C2645 VDDA.n193 GNDA 0.083406f
C2646 VDDA.t204 GNDA 0.023983f
C2647 VDDA.t78 GNDA 0.023983f
C2648 VDDA.n194 GNDA 0.083111f
C2649 VDDA.n195 GNDA 0.156905f
C2650 VDDA.n196 GNDA 0.021927f
C2651 VDDA.n197 GNDA 0.068276f
C2652 VDDA.n198 GNDA 0.092842f
C2653 VDDA.t397 GNDA 0.118311f
C2654 VDDA.t395 GNDA 0.041762f
C2655 VDDA.n199 GNDA 0.077183f
C2656 VDDA.n200 GNDA 0.049756f
C2657 VDDA.t370 GNDA 0.118311f
C2658 VDDA.t368 GNDA 0.041762f
C2659 VDDA.n201 GNDA 0.077183f
C2660 VDDA.n202 GNDA 0.049756f
C2661 VDDA.n203 GNDA 0.049336f
C2662 VDDA.n204 GNDA 0.092842f
C2663 VDDA.n205 GNDA 0.276684f
C2664 VDDA.t369 GNDA 0.412992f
C2665 VDDA.t234 GNDA 0.238456f
C2666 VDDA.t0 GNDA 0.238456f
C2667 VDDA.t230 GNDA 0.238456f
C2668 VDDA.t8 GNDA 0.238456f
C2669 VDDA.t260 GNDA 0.178842f
C2670 VDDA.n206 GNDA 0.119228f
C2671 VDDA.t445 GNDA 0.178842f
C2672 VDDA.t203 GNDA 0.238456f
C2673 VDDA.t77 GNDA 0.238456f
C2674 VDDA.t39 GNDA 0.238456f
C2675 VDDA.t228 GNDA 0.238456f
C2676 VDDA.t396 GNDA 0.412992f
C2677 VDDA.n207 GNDA 0.276684f
C2678 VDDA.n208 GNDA 0.068276f
C2679 VDDA.n209 GNDA 0.095583f
C2680 VDDA.t261 GNDA 0.023983f
C2681 VDDA.t446 GNDA 0.023983f
C2682 VDDA.n210 GNDA 0.078193f
C2683 VDDA.n211 GNDA 0.053368f
C2684 VDDA.n212 GNDA 0.044833f
C2685 VDDA.n213 GNDA 0.214864f
C2686 VDDA.n214 GNDA 0.084282f
C2687 VDDA.n216 GNDA 0.06687f
C2688 VDDA.n217 GNDA 0.012334f
C2689 VDDA.n218 GNDA 0.036433f
C2690 VDDA.n219 GNDA 0.036433f
C2691 VDDA.n220 GNDA 0.037149f
C2692 VDDA.n221 GNDA 0.093344f
C2693 VDDA.n222 GNDA 0.012334f
C2694 VDDA.n223 GNDA 0.053387f
C2695 VDDA.n224 GNDA 0.053387f
C2696 VDDA.n225 GNDA 0.056181f
C2697 VDDA.t241 GNDA 0.021927f
C2698 VDDA.n226 GNDA 0.07609f
C2699 VDDA.t379 GNDA 0.100155f
C2700 VDDA.n227 GNDA 0.049665f
C2701 VDDA.n228 GNDA 0.047678f
C2702 VDDA.t377 GNDA 0.038056f
C2703 VDDA.n229 GNDA 0.040291f
C2704 VDDA.n230 GNDA 0.031546f
C2705 VDDA.n231 GNDA 0.046872f
C2706 VDDA.n232 GNDA 0.309725f
C2707 VDDA.t378 GNDA 0.289526f
C2708 VDDA.n233 GNDA 0.095074f
C2709 VDDA.n234 GNDA 0.023768f
C2710 VDDA.t240 GNDA 0.133103f
C2711 VDDA.t399 GNDA 0.315801f
C2712 VDDA.n235 GNDA 0.310397f
C2713 VDDA.n236 GNDA 0.048626f
C2714 VDDA.n237 GNDA 0.031182f
C2715 VDDA.t398 GNDA 0.03874f
C2716 VDDA.n238 GNDA 0.040291f
C2717 VDDA.t400 GNDA 0.078228f
C2718 VDDA.n239 GNDA 0.053687f
C2719 VDDA.n240 GNDA 0.112868f
C2720 VDDA.n241 GNDA 0.073564f
C2721 VDDA.t330 GNDA 0.016017f
C2722 VDDA.n242 GNDA 0.017377f
C2723 VDDA.t328 GNDA 0.013437f
C2724 VDDA.n243 GNDA 0.017423f
C2725 VDDA.n244 GNDA 0.021905f
C2726 VDDA.n245 GNDA 0.030739f
C2727 VDDA.n246 GNDA 0.163961f
C2728 VDDA.t329 GNDA 0.181599f
C2729 VDDA.t62 GNDA 0.123339f
C2730 VDDA.t344 GNDA 0.181599f
C2731 VDDA.n247 GNDA 0.163961f
C2732 VDDA.n248 GNDA 0.030739f
C2733 VDDA.n249 GNDA 0.021905f
C2734 VDDA.t343 GNDA 0.013437f
C2735 VDDA.n250 GNDA 0.017423f
C2736 VDDA.t346 GNDA 0.016017f
C2737 VDDA.n251 GNDA 0.019437f
C2738 VDDA.n252 GNDA 0.075897f
C2739 VDDA.n253 GNDA 0.222153f
C2740 VDDA.n254 GNDA 4.5344f
C2741 VDDA.t470 GNDA 0.757536f
C2742 VDDA.t471 GNDA 0.807388f
C2743 VDDA.t469 GNDA 0.807388f
C2744 VDDA.t472 GNDA 0.774211f
C2745 VDDA.n255 GNDA 0.541196f
C2746 VDDA.n256 GNDA 0.262749f
C2747 VDDA.n257 GNDA 0.336861f
C2748 VDDA.n258 GNDA 2.4067f
C2749 VDDA.n259 GNDA 0.021927f
C2750 VDDA.n260 GNDA 0.016596f
C2751 VDDA.n261 GNDA 0.016596f
C2752 VDDA.n262 GNDA 0.0485f
C2753 VDDA.n263 GNDA 0.021927f
C2754 VDDA.t358 GNDA 0.025741f
C2755 VDDA.t356 GNDA 0.016962f
C2756 VDDA.n264 GNDA 0.04038f
C2757 VDDA.n265 GNDA 0.057456f
C2758 VDDA.n266 GNDA 0.108016f
C2759 VDDA.n267 GNDA 0.108016f
C2760 VDDA.t324 GNDA 0.025741f
C2761 VDDA.t322 GNDA 0.016962f
C2762 VDDA.n268 GNDA 0.04038f
C2763 VDDA.n269 GNDA 0.082226f
C2764 VDDA.n270 GNDA 0.057456f
C2765 VDDA.n271 GNDA 0.021927f
C2766 VDDA.n272 GNDA 0.016596f
C2767 VDDA.n273 GNDA 0.017352f
C2768 VDDA.n274 GNDA 0.017235f
C2769 VDDA.n275 GNDA 0.133977f
C2770 VDDA.n276 GNDA 0.017235f
C2771 VDDA.n277 GNDA 0.069788f
C2772 VDDA.n278 GNDA 0.017235f
C2773 VDDA.n279 GNDA 0.069788f
C2774 VDDA.n280 GNDA 0.016596f
C2775 VDDA.n281 GNDA 0.067401f
C2776 VDDA.n282 GNDA 0.108016f
C2777 VDDA.t373 GNDA 0.025741f
C2778 VDDA.t371 GNDA 0.016962f
C2779 VDDA.n283 GNDA 0.04038f
C2780 VDDA.n284 GNDA 0.057456f
C2781 VDDA.t427 GNDA 0.025741f
C2782 VDDA.t425 GNDA 0.016962f
C2783 VDDA.n285 GNDA 0.04038f
C2784 VDDA.n286 GNDA 0.057456f
C2785 VDDA.n287 GNDA 0.082226f
C2786 VDDA.n288 GNDA 0.108016f
C2787 VDDA.n289 GNDA 0.234857f
C2788 VDDA.t426 GNDA 0.214209f
C2789 VDDA.t431 GNDA 0.135673f
C2790 VDDA.t79 GNDA 0.135673f
C2791 VDDA.t106 GNDA 0.135673f
C2792 VDDA.t28 GNDA 0.135673f
C2793 VDDA.t2 GNDA 0.135673f
C2794 VDDA.t441 GNDA 0.135673f
C2795 VDDA.t433 GNDA 0.135673f
C2796 VDDA.t219 GNDA 0.135673f
C2797 VDDA.t81 GNDA 0.101755f
C2798 VDDA.n290 GNDA 0.067837f
C2799 VDDA.t178 GNDA 0.101755f
C2800 VDDA.t4 GNDA 0.135673f
C2801 VDDA.t437 GNDA 0.135673f
C2802 VDDA.t435 GNDA 0.135673f
C2803 VDDA.t217 GNDA 0.135673f
C2804 VDDA.t108 GNDA 0.135673f
C2805 VDDA.t180 GNDA 0.135673f
C2806 VDDA.t100 GNDA 0.135673f
C2807 VDDA.t439 GNDA 0.135673f
C2808 VDDA.t372 GNDA 0.214209f
C2809 VDDA.n291 GNDA 0.234857f
C2810 VDDA.n292 GNDA 0.067401f
C2811 VDDA.n293 GNDA 0.11482f
C2812 VDDA.n294 GNDA 0.0485f
C2813 VDDA.n295 GNDA 0.021927f
C2814 VDDA.n296 GNDA 0.017235f
C2815 VDDA.n297 GNDA 0.069788f
C2816 VDDA.n298 GNDA 0.017235f
C2817 VDDA.n299 GNDA 0.069788f
C2818 VDDA.n300 GNDA 0.017235f
C2819 VDDA.n301 GNDA 0.069788f
C2820 VDDA.n302 GNDA 0.017235f
C2821 VDDA.n303 GNDA 0.099937f
C2822 VDDA.n304 GNDA 0.021927f
C2823 VDDA.n305 GNDA 0.016596f
C2824 VDDA.n306 GNDA 0.016596f
C2825 VDDA.n307 GNDA 0.0485f
C2826 VDDA.n308 GNDA 0.021927f
C2827 VDDA.n309 GNDA 0.016596f
C2828 VDDA.n310 GNDA 0.021927f
C2829 VDDA.n311 GNDA 0.016596f
C2830 VDDA.n312 GNDA 0.0485f
C2831 VDDA.n313 GNDA 0.021927f
C2832 VDDA.n314 GNDA 0.021927f
C2833 VDDA.n315 GNDA 0.0485f
C2834 VDDA.n316 GNDA 0.021927f
C2835 VDDA.n317 GNDA 0.021927f
C2836 VDDA.n318 GNDA 0.016596f
C2837 VDDA.n319 GNDA 0.0485f
C2838 VDDA.n320 GNDA 0.021927f
C2839 VDDA.n321 GNDA 0.021927f
C2840 VDDA.n322 GNDA 0.0485f
C2841 VDDA.n323 GNDA 0.021927f
C2842 VDDA.n324 GNDA 0.016596f
C2843 VDDA.n325 GNDA 0.0485f
C2844 VDDA.n326 GNDA 0.021927f
C2845 VDDA.n327 GNDA 0.052076f
C2846 VDDA.n328 GNDA 0.0485f
C2847 VDDA.n329 GNDA 0.0358f
C2848 VDDA.n330 GNDA 0.034194f
C2849 VDDA.n331 GNDA 0.234857f
C2850 VDDA.t323 GNDA 0.214209f
C2851 VDDA.t465 GNDA 0.135673f
C2852 VDDA.t226 GNDA 0.135673f
C2853 VDDA.t133 GNDA 0.135673f
C2854 VDDA.t242 GNDA 0.135673f
C2855 VDDA.t246 GNDA 0.135673f
C2856 VDDA.t238 GNDA 0.135673f
C2857 VDDA.t6 GNDA 0.135673f
C2858 VDDA.t51 GNDA 0.135673f
C2859 VDDA.t224 GNDA 0.101755f
C2860 VDDA.n332 GNDA 0.067837f
C2861 VDDA.t461 GNDA 0.101755f
C2862 VDDA.t104 GNDA 0.135673f
C2863 VDDA.t459 GNDA 0.135673f
C2864 VDDA.t37 GNDA 0.135673f
C2865 VDDA.t131 GNDA 0.135673f
C2866 VDDA.t49 GNDA 0.135673f
C2867 VDDA.t201 GNDA 0.135673f
C2868 VDDA.t244 GNDA 0.135673f
C2869 VDDA.t60 GNDA 0.135673f
C2870 VDDA.t357 GNDA 0.214209f
C2871 VDDA.n333 GNDA 0.234857f
C2872 VDDA.n334 GNDA 0.034194f
C2873 VDDA.n335 GNDA 0.0358f
C2874 VDDA.n336 GNDA 0.0485f
C2875 VDDA.n337 GNDA 0.066382f
C2876 VDDA.n338 GNDA 0.201538f
C2877 VDDA.t291 GNDA 0.020556f
C2878 VDDA.t289 GNDA 0.020556f
C2879 VDDA.n339 GNDA 0.067912f
C2880 VDDA.n340 GNDA 0.087632f
C2881 VDDA.t409 GNDA 0.062997f
C2882 VDDA.n341 GNDA 0.111005f
C2883 VDDA.n342 GNDA 0.151321f
C2884 VDDA.n343 GNDA 0.151321f
C2885 VDDA.n344 GNDA 0.150626f
C2886 VDDA.t352 GNDA 0.062997f
C2887 VDDA.t350 GNDA 0.098022f
C2888 VDDA.t394 GNDA 0.025741f
C2889 VDDA.t392 GNDA 0.01299f
C2890 VDDA.n345 GNDA 0.040583f
C2891 VDDA.n346 GNDA 0.023401f
C2892 VDDA.n347 GNDA 0.041589f
C2893 VDDA.t415 GNDA 0.025741f
C2894 VDDA.t413 GNDA 0.01299f
C2895 VDDA.n348 GNDA 0.040583f
C2896 VDDA.n349 GNDA 0.041589f
C2897 VDDA.n350 GNDA 0.041589f
C2898 VDDA.n351 GNDA 0.034125f
C2899 VDDA.n352 GNDA 0.163981f
C2900 VDDA.t393 GNDA 0.205903f
C2901 VDDA.t36 GNDA 0.093275f
C2902 VDDA.n353 GNDA 0.062183f
C2903 VDDA.t455 GNDA 0.093275f
C2904 VDDA.t414 GNDA 0.208939f
C2905 VDDA.n354 GNDA 0.17225f
C2906 VDDA.n355 GNDA 0.034125f
C2907 VDDA.n356 GNDA 0.023401f
C2908 VDDA.n357 GNDA 0.032876f
C2909 VDDA.t310 GNDA 0.020556f
C2910 VDDA.t271 GNDA 0.020556f
C2911 VDDA.n358 GNDA 0.067912f
C2912 VDDA.n359 GNDA 0.087632f
C2913 VDDA.t282 GNDA 0.020556f
C2914 VDDA.t301 GNDA 0.020556f
C2915 VDDA.n360 GNDA 0.067912f
C2916 VDDA.n361 GNDA 0.087632f
C2917 VDDA.t266 GNDA 0.020556f
C2918 VDDA.t285 GNDA 0.020556f
C2919 VDDA.n362 GNDA 0.067912f
C2920 VDDA.n363 GNDA 0.087632f
C2921 VDDA.t299 GNDA 0.020556f
C2922 VDDA.t307 GNDA 0.020556f
C2923 VDDA.n364 GNDA 0.067912f
C2924 VDDA.n365 GNDA 0.087632f
C2925 VDDA.t280 GNDA 0.020556f
C2926 VDDA.t276 GNDA 0.020556f
C2927 VDDA.n366 GNDA 0.067912f
C2928 VDDA.n367 GNDA 0.087632f
C2929 VDDA.t305 GNDA 0.020556f
C2930 VDDA.t315 GNDA 0.020556f
C2931 VDDA.n368 GNDA 0.067912f
C2932 VDDA.n369 GNDA 0.087632f
C2933 VDDA.t273 GNDA 0.020556f
C2934 VDDA.t294 GNDA 0.020556f
C2935 VDDA.n370 GNDA 0.067912f
C2936 VDDA.n371 GNDA 0.087632f
C2937 VDDA.n372 GNDA 0.096756f
C2938 VDDA.n373 GNDA 0.116986f
C2939 VDDA.n374 GNDA 0.078854f
C2940 VDDA.n375 GNDA 0.096275f
C2941 VDDA.n376 GNDA 0.354727f
C2942 VDDA.t351 GNDA 0.457715f
C2943 VDDA.t272 GNDA 0.329932f
C2944 VDDA.t293 GNDA 0.329932f
C2945 VDDA.t304 GNDA 0.329932f
C2946 VDDA.t314 GNDA 0.329932f
C2947 VDDA.t279 GNDA 0.329932f
C2948 VDDA.t275 GNDA 0.329932f
C2949 VDDA.t298 GNDA 0.329932f
C2950 VDDA.t306 GNDA 0.247449f
C2951 VDDA.n377 GNDA 0.164966f
C2952 VDDA.t265 GNDA 0.247449f
C2953 VDDA.t284 GNDA 0.329932f
C2954 VDDA.t281 GNDA 0.329932f
C2955 VDDA.t300 GNDA 0.329932f
C2956 VDDA.t309 GNDA 0.329932f
C2957 VDDA.t270 GNDA 0.329932f
C2958 VDDA.t290 GNDA 0.329932f
C2959 VDDA.t288 GNDA 0.329932f
C2960 VDDA.t408 GNDA 0.457715f
C2961 VDDA.n378 GNDA 0.354727f
C2962 VDDA.n379 GNDA 0.096275f
C2963 VDDA.n380 GNDA 0.078854f
C2964 VDDA.t407 GNDA 0.098022f
C2965 VDDA.n381 GNDA 0.116986f
C2966 VDDA.n382 GNDA 0.053701f
C2967 VDDA.n383 GNDA 0.016549f
C2968 VDDA.t339 GNDA 0.025932f
C2969 VDDA.t337 GNDA 0.012654f
C2970 VDDA.n384 GNDA 0.038844f
C2971 VDDA.n385 GNDA 0.023293f
C2972 VDDA.n386 GNDA 0.041589f
C2973 VDDA.t336 GNDA 0.025932f
C2974 VDDA.t334 GNDA 0.012654f
C2975 VDDA.n387 GNDA 0.038844f
C2976 VDDA.n388 GNDA 0.041589f
C2977 VDDA.n389 GNDA 0.041589f
C2978 VDDA.n390 GNDA 0.034125f
C2979 VDDA.n391 GNDA 0.163981f
C2980 VDDA.t338 GNDA 0.205903f
C2981 VDDA.t71 GNDA 0.093275f
C2982 VDDA.n392 GNDA 0.062183f
C2983 VDDA.t463 GNDA 0.093275f
C2984 VDDA.t335 GNDA 0.205903f
C2985 VDDA.n393 GNDA 0.163981f
C2986 VDDA.n394 GNDA 0.034125f
C2987 VDDA.n395 GNDA 0.023293f
C2988 VDDA.n396 GNDA 0.024472f
C2989 VDDA.n397 GNDA 0.045806f
C2990 VDDA.n398 GNDA 0.096508f
C2991 VDDA.n399 GNDA 0.167583f
C2992 VDDA.n400 GNDA 0.017093f
C2993 VDDA.n401 GNDA 0.060337f
C2994 VDDA.t342 GNDA 0.027042f
C2995 VDDA.n402 GNDA 0.022612f
C2996 VDDA.n403 GNDA 0.048944f
C2997 VDDA.n404 GNDA 0.048944f
C2998 VDDA.n405 GNDA 0.048944f
C2999 VDDA.t403 GNDA 0.027042f
C3000 VDDA.t401 GNDA 0.013494f
C3001 VDDA.n406 GNDA 0.017061f
C3002 VDDA.n407 GNDA 0.060368f
C3003 VDDA.t418 GNDA 0.025806f
C3004 VDDA.n408 GNDA 0.045224f
C3005 VDDA.n409 GNDA 0.078716f
C3006 VDDA.n410 GNDA 0.078716f
C3007 VDDA.n411 GNDA 0.078716f
C3008 VDDA.t424 GNDA 0.025806f
C3009 VDDA.t422 GNDA 0.013494f
C3010 VDDA.n412 GNDA 0.0171f
C3011 VDDA.n413 GNDA 0.060329f
C3012 VDDA.t385 GNDA 0.027053f
C3013 VDDA.n414 GNDA 0.022612f
C3014 VDDA.n415 GNDA 0.048944f
C3015 VDDA.n416 GNDA 0.048944f
C3016 VDDA.n417 GNDA 0.048944f
C3017 VDDA.t318 GNDA 0.027053f
C3018 VDDA.t316 GNDA 0.013494f
C3019 VDDA.n418 GNDA 0.0171f
C3020 VDDA.n419 GNDA 0.082571f
C3021 VDDA.n420 GNDA 0.046331f
C3022 VDDA.n421 GNDA 0.027649f
C3023 VDDA.n422 GNDA 0.037985f
C3024 VDDA.n423 GNDA 0.173047f
C3025 VDDA.t317 GNDA 0.209524f
C3026 VDDA.t199 GNDA 0.126251f
C3027 VDDA.t195 GNDA 0.094688f
C3028 VDDA.n424 GNDA 0.063126f
C3029 VDDA.t142 GNDA 0.094688f
C3030 VDDA.t213 GNDA 0.126251f
C3031 VDDA.t384 GNDA 0.209524f
C3032 VDDA.n425 GNDA 0.173047f
C3033 VDDA.n426 GNDA 0.037985f
C3034 VDDA.n427 GNDA 0.027649f
C3035 VDDA.t383 GNDA 0.013922f
C3036 VDDA.n428 GNDA 0.045853f
C3037 VDDA.n429 GNDA 0.041649f
C3038 VDDA.n430 GNDA 0.017061f
C3039 VDDA.n431 GNDA 0.060368f
C3040 VDDA.n432 GNDA 0.017061f
C3041 VDDA.n433 GNDA 0.060368f
C3042 VDDA.n434 GNDA 0.017061f
C3043 VDDA.n435 GNDA 0.060368f
C3044 VDDA.n436 GNDA 0.017061f
C3045 VDDA.n437 GNDA 0.060368f
C3046 VDDA.n438 GNDA 0.041649f
C3047 VDDA.n439 GNDA 0.046672f
C3048 VDDA.n440 GNDA 0.042724f
C3049 VDDA.n441 GNDA 0.053248f
C3050 VDDA.n442 GNDA 0.203575f
C3051 VDDA.t423 GNDA 0.209524f
C3052 VDDA.t447 GNDA 0.126251f
C3053 VDDA.t467 GNDA 0.126251f
C3054 VDDA.t451 GNDA 0.126251f
C3055 VDDA.t30 GNDA 0.126251f
C3056 VDDA.t453 GNDA 0.126251f
C3057 VDDA.t457 GNDA 0.094688f
C3058 VDDA.n443 GNDA 0.063126f
C3059 VDDA.t176 GNDA 0.094688f
C3060 VDDA.t174 GNDA 0.126251f
C3061 VDDA.t140 GNDA 0.126251f
C3062 VDDA.t215 GNDA 0.126251f
C3063 VDDA.t417 GNDA 0.331696f
C3064 VDDA.n444 GNDA 0.333905f
C3065 VDDA.n445 GNDA 0.061131f
C3066 VDDA.n446 GNDA 0.042379f
C3067 VDDA.t416 GNDA 0.013494f
C3068 VDDA.n447 GNDA 0.046672f
C3069 VDDA.n448 GNDA 0.049187f
C3070 VDDA.n449 GNDA 0.017093f
C3071 VDDA.n450 GNDA 0.060337f
C3072 VDDA.n451 GNDA 0.049187f
C3073 VDDA.n452 GNDA 0.045436f
C3074 VDDA.n453 GNDA 0.027649f
C3075 VDDA.n454 GNDA 0.03746f
C3076 VDDA.n455 GNDA 0.171176f
C3077 VDDA.t402 GNDA 0.205903f
C3078 VDDA.t75 GNDA 0.124367f
C3079 VDDA.t144 GNDA 0.084796f
C3080 VDDA.n456 GNDA 0.031092f
C3081 VDDA.n457 GNDA 0.039571f
C3082 VDDA.t197 GNDA 0.093275f
C3083 VDDA.t159 GNDA 0.124367f
C3084 VDDA.t341 GNDA 0.205903f
C3085 VDDA.n458 GNDA 0.172225f
C3086 VDDA.n459 GNDA 0.038509f
C3087 VDDA.n460 GNDA 0.027649f
C3088 VDDA.t340 GNDA 0.013494f
C3089 VDDA.n461 GNDA 0.045436f
C3090 VDDA.n462 GNDA 0.090624f
C3091 VDDA.n463 GNDA 0.136034f
C3092 VDDA.t303 GNDA 0.383036f
C3093 VDDA.t311 GNDA 0.384424f
C3094 VDDA.t283 GNDA 0.383036f
C3095 VDDA.t267 GNDA 0.384424f
C3096 VDDA.t292 GNDA 0.383036f
C3097 VDDA.t296 GNDA 0.384424f
C3098 VDDA.t268 GNDA 0.383036f
C3099 VDDA.t308 GNDA 0.384424f
C3100 VDDA.t297 GNDA 0.383036f
C3101 VDDA.t313 GNDA 0.384424f
C3102 VDDA.t286 GNDA 0.383036f
C3103 VDDA.t269 GNDA 0.384424f
C3104 VDDA.t264 GNDA 0.383036f
C3105 VDDA.t278 GNDA 0.384424f
C3106 VDDA.t302 GNDA 0.383036f
C3107 VDDA.t287 GNDA 0.384424f
C3108 VDDA.n464 GNDA 0.25675f
C3109 VDDA.t295 GNDA 0.204463f
C3110 VDDA.n465 GNDA 0.278579f
C3111 VDDA.t277 GNDA 0.204463f
C3112 VDDA.n466 GNDA 0.278579f
C3113 VDDA.t312 GNDA 0.204463f
C3114 VDDA.n467 GNDA 0.278579f
C3115 VDDA.t274 GNDA 0.3051f
C3116 VDDA.n468 GNDA 0.265857f
C3117 VDDA.n469 GNDA 0.826218f
C3118 bgr_0.Vin-.n0 GNDA 0.073641f
C3119 bgr_0.Vin-.n1 GNDA 0.338979f
C3120 bgr_0.Vin-.n2 GNDA 0.510703f
C3121 bgr_0.Vin-.t2 GNDA 0.276239f
C3122 bgr_0.Vin-.n3 GNDA 0.331333f
C3123 bgr_0.Vin-.n4 GNDA 0.073776f
C3124 bgr_0.Vin-.n5 GNDA 0.12627f
C3125 bgr_0.Vin-.n6 GNDA 0.074468f
C3126 bgr_0.Vin-.n7 GNDA 0.998981f
C3127 bgr_0.Vin-.t3 GNDA 0.028614f
C3128 bgr_0.Vin-.t6 GNDA 0.028614f
C3129 bgr_0.Vin-.n8 GNDA 0.099613f
C3130 bgr_0.Vin-.t4 GNDA 0.028614f
C3131 bgr_0.Vin-.t5 GNDA 0.028614f
C3132 bgr_0.Vin-.n9 GNDA 0.095121f
C3133 bgr_0.Vin-.n10 GNDA 0.408067f
C3134 bgr_0.Vin-.t1 GNDA 0.098662f
C3135 bgr_0.Vin-.n11 GNDA 0.025702f
C3136 bgr_0.Vin-.n12 GNDA 0.469862f
C3137 bgr_0.Vin-.n13 GNDA 0.222852f
C3138 bgr_0.Vin-.t10 GNDA 0.023594f
C3139 bgr_0.Vin-.n14 GNDA 0.027673f
C3140 bgr_0.Vin-.n15 GNDA 0.022653f
C3141 bgr_0.Vin-.n16 GNDA 0.022653f
C3142 bgr_0.Vin-.n17 GNDA 0.040466f
C3143 bgr_0.Vin-.n18 GNDA 0.524007f
C3144 bgr_0.Vin-.n19 GNDA 0.461299f
C3145 bgr_0.Vin-.n20 GNDA 0.166915f
C3146 bgr_0.Vin-.n21 GNDA 0.074625f
C3147 bgr_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17.Emitter GNDA 0.043026f
C3148 bgr_0.V_TOP.t31 GNDA 0.115045f
C3149 bgr_0.V_TOP.t44 GNDA 0.115045f
C3150 bgr_0.V_TOP.t18 GNDA 0.115045f
C3151 bgr_0.V_TOP.t26 GNDA 0.115045f
C3152 bgr_0.V_TOP.t37 GNDA 0.115045f
C3153 bgr_0.V_TOP.t35 GNDA 0.115045f
C3154 bgr_0.V_TOP.t48 GNDA 0.115045f
C3155 bgr_0.V_TOP.t20 GNDA 0.115045f
C3156 bgr_0.V_TOP.t27 GNDA 0.115045f
C3157 bgr_0.V_TOP.t41 GNDA 0.115045f
C3158 bgr_0.V_TOP.t38 GNDA 0.115045f
C3159 bgr_0.V_TOP.t14 GNDA 0.115045f
C3160 bgr_0.V_TOP.t23 GNDA 0.115045f
C3161 bgr_0.V_TOP.t29 GNDA 0.115045f
C3162 bgr_0.V_TOP.t43 GNDA 0.150392f
C3163 bgr_0.V_TOP.n0 GNDA 0.084081f
C3164 bgr_0.V_TOP.n1 GNDA 0.061357f
C3165 bgr_0.V_TOP.n2 GNDA 0.061357f
C3166 bgr_0.V_TOP.n3 GNDA 0.061357f
C3167 bgr_0.V_TOP.n4 GNDA 0.061357f
C3168 bgr_0.V_TOP.n5 GNDA 0.057217f
C3169 bgr_0.V_TOP.t12 GNDA 0.147947f
C3170 bgr_0.V_TOP.t3 GNDA 0.155772f
C3171 bgr_0.V_TOP.t2 GNDA 0.010957f
C3172 bgr_0.V_TOP.t6 GNDA 0.010957f
C3173 bgr_0.V_TOP.n6 GNDA 0.027281f
C3174 bgr_0.V_TOP.n7 GNDA 0.726844f
C3175 bgr_0.V_TOP.t11 GNDA 0.010957f
C3176 bgr_0.V_TOP.t7 GNDA 0.010957f
C3177 bgr_0.V_TOP.n8 GNDA 0.026425f
C3178 bgr_0.V_TOP.t1 GNDA 0.010957f
C3179 bgr_0.V_TOP.t0 GNDA 0.010957f
C3180 bgr_0.V_TOP.n9 GNDA 0.027465f
C3181 bgr_0.V_TOP.t13 GNDA 0.010957f
C3182 bgr_0.V_TOP.t4 GNDA 0.010957f
C3183 bgr_0.V_TOP.n10 GNDA 0.027281f
C3184 bgr_0.V_TOP.n11 GNDA 0.252824f
C3185 bgr_0.V_TOP.n12 GNDA 0.153577f
C3186 bgr_0.V_TOP.n13 GNDA 0.087653f
C3187 bgr_0.V_TOP.t9 GNDA 0.010957f
C3188 bgr_0.V_TOP.t8 GNDA 0.010957f
C3189 bgr_0.V_TOP.n14 GNDA 0.027281f
C3190 bgr_0.V_TOP.n15 GNDA 0.151313f
C3191 bgr_0.V_TOP.t10 GNDA 0.010957f
C3192 bgr_0.V_TOP.t5 GNDA 0.010957f
C3193 bgr_0.V_TOP.n16 GNDA 0.027281f
C3194 bgr_0.V_TOP.n17 GNDA 0.149874f
C3195 bgr_0.V_TOP.n18 GNDA 0.329448f
C3196 bgr_0.V_TOP.n19 GNDA 0.023183f
C3197 bgr_0.V_TOP.n20 GNDA 0.057217f
C3198 bgr_0.V_TOP.n21 GNDA 0.061357f
C3199 bgr_0.V_TOP.n22 GNDA 0.061357f
C3200 bgr_0.V_TOP.n23 GNDA 0.061357f
C3201 bgr_0.V_TOP.n24 GNDA 0.061357f
C3202 bgr_0.V_TOP.n25 GNDA 0.061357f
C3203 bgr_0.V_TOP.n26 GNDA 0.061357f
C3204 bgr_0.V_TOP.n27 GNDA 0.057217f
C3205 bgr_0.V_TOP.t32 GNDA 0.132572f
C3206 bgr_0.V_TOP.t49 GNDA 0.445732f
C3207 bgr_0.V_TOP.t39 GNDA 0.438267f
C3208 bgr_0.V_TOP.n28 GNDA 0.293844f
C3209 bgr_0.V_TOP.t28 GNDA 0.438267f
C3210 bgr_0.V_TOP.t25 GNDA 0.445732f
C3211 bgr_0.V_TOP.t33 GNDA 0.438267f
C3212 bgr_0.V_TOP.n29 GNDA 0.293844f
C3213 bgr_0.V_TOP.n30 GNDA 0.273917f
C3214 bgr_0.V_TOP.t21 GNDA 0.445732f
C3215 bgr_0.V_TOP.t15 GNDA 0.438267f
C3216 bgr_0.V_TOP.n31 GNDA 0.293844f
C3217 bgr_0.V_TOP.t40 GNDA 0.438267f
C3218 bgr_0.V_TOP.t34 GNDA 0.445732f
C3219 bgr_0.V_TOP.t45 GNDA 0.438267f
C3220 bgr_0.V_TOP.n32 GNDA 0.293844f
C3221 bgr_0.V_TOP.n33 GNDA 0.356092f
C3222 bgr_0.V_TOP.t30 GNDA 0.445732f
C3223 bgr_0.V_TOP.t22 GNDA 0.438267f
C3224 bgr_0.V_TOP.n34 GNDA 0.293844f
C3225 bgr_0.V_TOP.t16 GNDA 0.438267f
C3226 bgr_0.V_TOP.t46 GNDA 0.445732f
C3227 bgr_0.V_TOP.t19 GNDA 0.438267f
C3228 bgr_0.V_TOP.n35 GNDA 0.293844f
C3229 bgr_0.V_TOP.n36 GNDA 0.356092f
C3230 bgr_0.V_TOP.t24 GNDA 0.445732f
C3231 bgr_0.V_TOP.t17 GNDA 0.438267f
C3232 bgr_0.V_TOP.n37 GNDA 0.293844f
C3233 bgr_0.V_TOP.t42 GNDA 0.438267f
C3234 bgr_0.V_TOP.n38 GNDA 0.273917f
C3235 bgr_0.V_TOP.t47 GNDA 0.438267f
C3236 bgr_0.V_TOP.n39 GNDA 0.191742f
C3237 bgr_0.V_TOP.t36 GNDA 0.438267f
C3238 bgr_0.V_TOP.n40 GNDA 0.893239f
.ends

