* PEX produced on Sat Feb  1 12:17:34 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from div5.ext - technology: sky130A

.subckt div5
X0 M.t3 Q2_b.t2 GNDA.t23 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X1 E.t1 VIN VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X2 D.t3 VIN GNDA.t37 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X3 I.t0 VOUT.t2 GNDA.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X4 Q2_b.t1 VIN VDDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X5 F.t1 E.t2 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X6 GNDA.t35 VIN J.t3 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X7 A.t2 Q2_b.t3 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X8 B.t1 VIN C.t1 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X9 I.t2 Q2_b.t4 H.t0 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X10 A.t0 Q2_b.t5 GNDA.t20 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X11 GNDA.t32 VIN D.t2 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X12 VDDA.t4 A.t3 B.t0 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X13 K.t1 Q2_b.t6 L.t1 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X14 GNDA.t30 VIN J.t2 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X15 GNDA.t17 Q2_b.t7 M.t2 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X16 VDDA.t1 VOUT.t3 K.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X17 GNDA.t15 Q2_b.t8 M.t1 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X18 G.t0 VOUT.t4 F.t0 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X19 GNDA.t28 VIN D.t1 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X20 GNDA.t9 E.t3 I.t1 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X21 J.t1 VIN GNDA.t26 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X22 E.t0 D.t4 GNDA.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X23 VDDA.t6 G.t3 J.t0 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X24 D.t0 B.t2 VDDA.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X25 VDDA.t18 Q2_b.t9 G.t1 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X26 VDDA.t16 Q2_b.t10 A.t1 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X27 C.t0 A.t4 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X28 H.t1 VIN G.t2 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X29 Q2_b.t0 J.t4 GNDA.t13 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X30 VOUT.t1 M.t4 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X31 M.t0 K.t2 VDDA.t12 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X32 VOUT.t0 Q2_b.t11 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X33 L.t0 VOUT.t5 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
R0 Q2_b.n6 Q2_b.t5 2779.53
R1 Q2_b.n7 Q2_b.n6 1206
R2 Q2_b.n4 Q2_b.t1 777.4
R3 Q2_b.t4 Q2_b.t9 514.134
R4 Q2_b.n3 Q2_b.n2 364.178
R5 Q2_b.n0 Q2_b.t11 353.467
R6 Q2_b.t5 Q2_b.n5 353.467
R7 Q2_b.n5 Q2_b.t3 289.2
R8 Q2_b.n4 Q2_b.n3 257.079
R9 Q2_b.t0 Q2_b.n7 233
R10 Q2_b.n6 Q2_b.t4 208.868
R11 Q2_b.n0 Q2_b.t7 192.8
R12 Q2_b.n2 Q2_b.n1 176.733
R13 Q2_b.n2 Q2_b.t8 112.468
R14 Q2_b.n1 Q2_b.t2 112.468
R15 Q2_b.n3 Q2_b.t6 112.468
R16 Q2_b.n5 Q2_b.t10 112.468
R17 Q2_b.n1 Q2_b.n0 96.4005
R18 Q2_b.n7 Q2_b.n4 21.3338
R19 GNDA.t10 GNDA.t24 3500
R20 GNDA.t12 GNDA.t0 3400
R21 GNDA.t2 GNDA.t34 3300
R22 GNDA.n10 GNDA.t19 3150
R23 GNDA.t18 GNDA.t14 2500
R24 GNDA.t33 GNDA.t27 2500
R25 GNDA.n10 GNDA.t4 1350
R26 GNDA.n2 GNDA.n10 1173.79
R27 GNDA.t16 GNDA.t6 1100
R28 GNDA.t22 GNDA.t16 1100
R29 GNDA.t14 GNDA.t22 1100
R30 GNDA.t0 GNDA.t18 1100
R31 GNDA.t29 GNDA.t12 1100
R32 GNDA.t25 GNDA.t29 1100
R33 GNDA.t34 GNDA.t25 1100
R34 GNDA.t8 GNDA.t2 1100
R35 GNDA.t21 GNDA.t8 1100
R36 GNDA.t24 GNDA.t21 1100
R37 GNDA.t31 GNDA.t10 1100
R38 GNDA.t36 GNDA.t31 1100
R39 GNDA.t27 GNDA.t36 1100
R40 GNDA.t4 GNDA.t33 1100
R41 GNDA GNDA.t20 242.3
R42 GNDA.n0 GNDA.t1 242.3
R43 GNDA.n2 GNDA.t5 236.792
R44 GNDA.n0 GNDA.n3 194.576
R45 GNDA.n1 GNDA.n9 194.3
R46 GNDA.n1 GNDA.n8 194.3
R47 GNDA.n1 GNDA.n7 194.3
R48 GNDA.n1 GNDA.n6 194.3
R49 GNDA.n1 GNDA.n5 194.3
R50 GNDA.n0 GNDA.n4 194.3
R51 GNDA.n9 GNDA.t37 48.0005
R52 GNDA.n9 GNDA.t28 48.0005
R53 GNDA.n8 GNDA.t11 48.0005
R54 GNDA.n8 GNDA.t32 48.0005
R55 GNDA.n7 GNDA.t3 48.0005
R56 GNDA.n7 GNDA.t9 48.0005
R57 GNDA.n6 GNDA.t26 48.0005
R58 GNDA.n6 GNDA.t35 48.0005
R59 GNDA.n5 GNDA.t13 48.0005
R60 GNDA.n5 GNDA.t30 48.0005
R61 GNDA.n4 GNDA.t23 48.0005
R62 GNDA.n4 GNDA.t15 48.0005
R63 GNDA.n3 GNDA.t7 48.0005
R64 GNDA.n3 GNDA.t17 48.0005
R65 GNDA.n2 GNDA 2.75546
R66 GNDA GNDA.n1 2.2755
R67 GNDA.n1 GNDA.n0 1.838
R68 M.n0 M.t0 761.4
R69 M.n1 M.t4 349.433
R70 M.n0 M.t1 254.333
R71 M.n2 M.n1 206.333
R72 M.n1 M.n0 70.4005
R73 M.n2 M.t2 48.0005
R74 M.t3 M.n2 48.0005
R75 VDDA.t23 VDDA.t17 2804.76
R76 VDDA.t21 VDDA.t0 2533.33
R77 VDDA.t3 VDDA.t19 1538.1
R78 VDDA.t2 VDDA.t5 1492.86
R79 VDDA.t11 VDDA.n7 1289.29
R80 VDDA.n8 VDDA.t7 1289.29
R81 VDDA.n6 VDDA.t14 667.62
R82 VDDA.n1 VDDA.t24 667.592
R83 VDDA.n7 VDDA.t13 610.715
R84 VDDA.n8 VDDA.t23 610.715
R85 VDDA VDDA.n10 594.301
R86 VDDA.n0 VDDA.n9 594.301
R87 VDDA.n0 VDDA.n2 594.301
R88 VDDA.n0 VDDA.n3 594.301
R89 VDDA.n5 VDDA.n4 594.301
R90 VDDA.t0 VDDA.t11 497.62
R91 VDDA.t5 VDDA.t21 497.62
R92 VDDA.t9 VDDA.t2 497.62
R93 VDDA.t17 VDDA.t9 497.62
R94 VDDA.t7 VDDA.t3 497.62
R95 VDDA.t19 VDDA.t15 497.62
R96 VDDA.n7 VDDA.n6 373.781
R97 VDDA.n10 VDDA.t20 78.8005
R98 VDDA.n10 VDDA.t16 78.8005
R99 VDDA.n9 VDDA.t8 78.8005
R100 VDDA.n9 VDDA.t4 78.8005
R101 VDDA.n2 VDDA.t10 78.8005
R102 VDDA.n2 VDDA.t18 78.8005
R103 VDDA.n3 VDDA.t22 78.8005
R104 VDDA.n3 VDDA.t6 78.8005
R105 VDDA.n4 VDDA.t12 78.8005
R106 VDDA.n4 VDDA.t1 78.8005
R107 VDDA.n1 VDDA.n0 2.75546
R108 VDDA.n1 VDDA.n8 373.793
R109 VDDA.n6 VDDA.n5 3.20124
R110 VDDA VDDA.n0 2.0005
R111 VDDA.n5 VDDA.n0 1.5255
R112 E.n0 E.t2 1207.57
R113 E.n0 E.t1 723
R114 E.t2 E.t3 514.134
R115 E.t0 E.n0 314.921
R116 D.n0 D.t0 761.4
R117 D.n1 D.t4 350.349
R118 D.n0 D.t1 254.333
R119 D.n2 D.n1 206.333
R120 D.n1 D.n0 70.4005
R121 D.n2 D.t2 48.0005
R122 D.t3 D.n2 48.0005
R123 VOUT.n2 VOUT.n1 2120.39
R124 VOUT.n1 VOUT.t4 1992.27
R125 VOUT.n2 VOUT.t0 796.388
R126 VOUT.t4 VOUT.t2 514.134
R127 VOUT.n0 VOUT.t5 289.2
R128 VOUT.t1 VOUT.n2 233
R129 VOUT.n1 VOUT.n0 208.868
R130 VOUT.n0 VOUT.t3 176.733
R131 I.t0 I.n0 531.067
R132 I.n0 I.t1 48.0005
R133 I.n0 I.t2 48.0005
R134 F.t0 F.t1 157.601
R135 J.n2 J.t0 723.534
R136 J.n1 J.t4 553.534
R137 J.t3 J.n2 254.333
R138 J.n1 J.n0 206.333
R139 J.n2 J.n1 70.4005
R140 J.n0 J.t2 48.0005
R141 J.n0 J.t1 48.0005
R142 A.n2 A.t1 755.534
R143 A.t2 A.n2 685.134
R144 A.n1 A.n0 389.733
R145 A.n1 A.t0 340.2
R146 A.n0 A.t4 321.334
R147 A.n0 A.t3 144.601
R148 A.n2 A.n1 19.2005
R149 C.t0 C.t1 96.0005
R150 B.n0 B.t0 663.801
R151 B.n0 B.t2 380.368
R152 B B.t1 282.921
R153 B B.n0 114.133
R154 H.t0 H.t1 96.0005
R155 L.t0 L.t1 96.0005
R156 K.n0 K.t0 663.801
R157 K.t1 K.n0 397.053
R158 K.n0 K.t2 380.368
R159 G.n0 G.t0 685.134
R160 G.n1 G.t1 685.134
R161 G.n0 G.t3 534.268
R162 G.t2 G.n1 340.521
R163 G.n1 G.n0 105.6
C0 VDDA VIN 0.290147f
C1 VIN B 0.143413f
C2 VDDA B 0.305296f
C3 VIN GNDA 1.85246f
C4 B GNDA 0.256727f
C5 VDDA GNDA 3.92947f
.ends

