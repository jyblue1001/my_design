magic
tech sky130A
timestamp 1755896225
<< metal1 >>
rect 2070 19310 2190 19325
rect 2070 19280 2115 19310
rect 2145 19280 2190 19310
rect 2070 19245 2190 19280
rect 2070 19215 2115 19245
rect 2145 19215 2190 19245
rect 2070 19175 2190 19215
rect 2070 19145 2115 19175
rect 2145 19145 2190 19175
rect 2070 19105 2190 19145
rect 2070 19075 2115 19105
rect 2145 19075 2190 19105
rect 2070 19035 2190 19075
rect 2070 19005 2115 19035
rect 2145 19005 2190 19035
rect 2070 18970 2190 19005
rect 2070 18940 2115 18970
rect 2145 18940 2190 18970
rect 2070 18910 2190 18940
rect 2070 18880 2115 18910
rect 2145 18880 2190 18910
rect 2070 18845 2190 18880
rect 2070 18815 2115 18845
rect 2145 18815 2190 18845
rect 2070 18775 2190 18815
rect 2070 18745 2115 18775
rect 2145 18745 2190 18775
rect 2070 18705 2190 18745
rect 2070 18675 2115 18705
rect 2145 18675 2190 18705
rect 2070 18635 2190 18675
rect 2070 18605 2115 18635
rect 2145 18605 2190 18635
rect 2070 18570 2190 18605
rect 2070 18540 2115 18570
rect 2145 18540 2190 18570
rect 2070 18510 2190 18540
rect 2070 18480 2115 18510
rect 2145 18480 2190 18510
rect 2070 18445 2190 18480
rect 2070 18415 2115 18445
rect 2145 18415 2190 18445
rect 2070 18375 2190 18415
rect 2070 18345 2115 18375
rect 2145 18345 2190 18375
rect 2070 18305 2190 18345
rect 2070 18275 2115 18305
rect 2145 18275 2190 18305
rect 2070 18235 2190 18275
rect 2070 18205 2115 18235
rect 2145 18205 2190 18235
rect 2070 18170 2190 18205
rect 2070 18140 2115 18170
rect 2145 18140 2190 18170
rect 2070 18110 2190 18140
rect 2070 18080 2115 18110
rect 2145 18080 2190 18110
rect 2070 18045 2190 18080
rect 2070 18015 2115 18045
rect 2145 18015 2190 18045
rect 2070 17975 2190 18015
rect 2070 17945 2115 17975
rect 2145 17945 2190 17975
rect 2070 17905 2190 17945
rect 2070 17875 2115 17905
rect 2145 17875 2190 17905
rect 2070 17835 2190 17875
rect 2070 17805 2115 17835
rect 2145 17805 2190 17835
rect 2070 17770 2190 17805
rect 2070 17740 2115 17770
rect 2145 17740 2190 17770
rect 2070 15690 2190 17740
rect 6690 19310 6750 19325
rect 6690 19280 6705 19310
rect 6735 19280 6750 19310
rect 6690 19245 6750 19280
rect 6690 19215 6705 19245
rect 6735 19215 6750 19245
rect 6690 19175 6750 19215
rect 6690 19145 6705 19175
rect 6735 19145 6750 19175
rect 6690 19105 6750 19145
rect 6690 19075 6705 19105
rect 6735 19075 6750 19105
rect 6690 19035 6750 19075
rect 6690 19005 6705 19035
rect 6735 19005 6750 19035
rect 6690 18970 6750 19005
rect 6690 18940 6705 18970
rect 6735 18940 6750 18970
rect 6690 18910 6750 18940
rect 6690 18880 6705 18910
rect 6735 18880 6750 18910
rect 6690 18845 6750 18880
rect 6690 18815 6705 18845
rect 6735 18815 6750 18845
rect 6690 18775 6750 18815
rect 6690 18745 6705 18775
rect 6735 18745 6750 18775
rect 6690 18705 6750 18745
rect 6690 18675 6705 18705
rect 6735 18675 6750 18705
rect 6690 18635 6750 18675
rect 6690 18605 6705 18635
rect 6735 18605 6750 18635
rect 6690 18570 6750 18605
rect 6690 18540 6705 18570
rect 6735 18540 6750 18570
rect 6690 18510 6750 18540
rect 6690 18480 6705 18510
rect 6735 18480 6750 18510
rect 6690 18445 6750 18480
rect 6690 18415 6705 18445
rect 6735 18415 6750 18445
rect 6690 18375 6750 18415
rect 6690 18345 6705 18375
rect 6735 18345 6750 18375
rect 6690 18305 6750 18345
rect 6690 18275 6705 18305
rect 6735 18275 6750 18305
rect 6690 18235 6750 18275
rect 6690 18205 6705 18235
rect 6735 18205 6750 18235
rect 6690 18170 6750 18205
rect 6690 18140 6705 18170
rect 6735 18140 6750 18170
rect 6690 18110 6750 18140
rect 6690 18080 6705 18110
rect 6735 18080 6750 18110
rect 6690 18045 6750 18080
rect 6690 18015 6705 18045
rect 6735 18015 6750 18045
rect 6690 17975 6750 18015
rect 6690 17945 6705 17975
rect 6735 17945 6750 17975
rect 6690 17905 6750 17945
rect 6690 17875 6705 17905
rect 6735 17875 6750 17905
rect 6690 17835 6750 17875
rect 6690 17805 6705 17835
rect 6735 17805 6750 17835
rect 6690 17770 6750 17805
rect 6690 17740 6705 17770
rect 6735 17740 6750 17770
rect 6690 17725 6750 17740
rect 2070 15660 2075 15690
rect 2105 15660 2115 15690
rect 2145 15660 2155 15690
rect 2185 15660 2190 15690
rect 2070 15650 2190 15660
rect 2070 15620 2075 15650
rect 2105 15620 2115 15650
rect 2145 15620 2155 15650
rect 2185 15620 2190 15650
rect 2070 15610 2190 15620
rect 2070 15580 2075 15610
rect 2105 15580 2115 15610
rect 2145 15580 2155 15610
rect 2185 15580 2190 15610
rect 2070 12710 2190 15580
rect 2070 12680 2075 12710
rect 2105 12680 2115 12710
rect 2145 12680 2155 12710
rect 2185 12680 2190 12710
rect 2070 12670 2190 12680
rect 2070 12640 2075 12670
rect 2105 12640 2115 12670
rect 2145 12640 2155 12670
rect 2185 12640 2190 12670
rect 2070 12550 2190 12640
rect 2070 12520 2075 12550
rect 2105 12520 2115 12550
rect 2145 12520 2155 12550
rect 2185 12520 2190 12550
rect 2070 12510 2190 12520
rect 2070 12480 2075 12510
rect 2105 12480 2115 12510
rect 2145 12480 2155 12510
rect 2185 12480 2190 12510
rect 2070 12470 2190 12480
rect 2070 12440 2075 12470
rect 2105 12440 2115 12470
rect 2145 12440 2155 12470
rect 2185 12440 2190 12470
rect 2070 12435 2190 12440
rect 2205 15925 2325 15930
rect 2205 15895 2210 15925
rect 2240 15895 2250 15925
rect 2280 15895 2290 15925
rect 2320 15895 2325 15925
rect -120 9635 0 9650
rect -120 9605 -75 9635
rect -45 9605 0 9635
rect -120 9570 0 9605
rect -120 9540 -75 9570
rect -45 9540 0 9570
rect -120 9500 0 9540
rect -120 9470 -75 9500
rect -45 9470 0 9500
rect -120 9430 0 9470
rect -120 9400 -75 9430
rect -45 9400 0 9430
rect -120 9360 0 9400
rect -120 9330 -75 9360
rect -45 9330 0 9360
rect -120 9295 0 9330
rect -120 9265 -75 9295
rect -45 9265 0 9295
rect -120 9235 0 9265
rect -120 9205 -75 9235
rect -45 9205 0 9235
rect -120 9170 0 9205
rect -120 9140 -75 9170
rect -45 9140 0 9170
rect -120 9100 0 9140
rect -120 9070 -75 9100
rect -45 9070 0 9100
rect -120 9030 0 9070
rect -120 9000 -75 9030
rect -45 9000 0 9030
rect -120 8960 0 9000
rect -120 8930 -75 8960
rect -45 8930 0 8960
rect -120 8895 0 8930
rect -120 8865 -75 8895
rect -45 8865 0 8895
rect -120 8835 0 8865
rect -120 8805 -75 8835
rect -45 8805 0 8835
rect -120 8770 0 8805
rect -120 8740 -75 8770
rect -45 8740 0 8770
rect -120 8700 0 8740
rect -120 8670 -75 8700
rect -45 8670 0 8700
rect -120 8630 0 8670
rect -120 8600 -75 8630
rect -45 8600 0 8630
rect -120 8560 0 8600
rect -120 8530 -75 8560
rect -45 8530 0 8560
rect -120 8495 0 8530
rect -120 8465 -75 8495
rect -45 8465 0 8495
rect -120 8435 0 8465
rect -120 8405 -75 8435
rect -45 8405 0 8435
rect -120 8370 0 8405
rect -120 8340 -75 8370
rect -45 8340 0 8370
rect -120 8300 0 8340
rect -120 8270 -75 8300
rect -45 8270 0 8300
rect -120 8230 0 8270
rect -120 8200 -75 8230
rect -45 8200 0 8230
rect -120 8160 0 8200
rect -120 8130 -75 8160
rect -45 8130 0 8160
rect -120 8095 0 8130
rect -120 8065 -75 8095
rect -45 8065 0 8095
rect -120 8035 0 8065
rect -120 8005 -75 8035
rect -45 8005 0 8035
rect -120 7970 0 8005
rect -120 7940 -75 7970
rect -45 7940 0 7970
rect -120 7900 0 7940
rect -120 7870 -75 7900
rect -45 7870 0 7900
rect -120 7830 0 7870
rect -120 7800 -75 7830
rect -45 7800 0 7830
rect -120 7760 0 7800
rect -120 7730 -75 7760
rect -45 7730 0 7760
rect -120 7695 0 7730
rect -120 7665 -75 7695
rect -45 7665 0 7695
rect -120 7635 0 7665
rect -120 7605 -75 7635
rect -45 7605 0 7635
rect -120 7570 0 7605
rect -120 7540 -75 7570
rect -45 7540 0 7570
rect -120 7500 0 7540
rect -120 7470 -75 7500
rect -45 7470 0 7500
rect -120 7430 0 7470
rect -120 7400 -75 7430
rect -45 7400 0 7430
rect -120 7360 0 7400
rect -120 7330 -75 7360
rect -45 7330 0 7360
rect -120 7295 0 7330
rect -120 7265 -75 7295
rect -45 7265 0 7295
rect -120 7235 0 7265
rect -120 7205 -75 7235
rect -45 7205 0 7235
rect -120 7170 0 7205
rect -120 7140 -75 7170
rect -45 7140 0 7170
rect -120 7100 0 7140
rect -120 7070 -75 7100
rect -45 7070 0 7100
rect -120 7030 0 7070
rect -120 7000 -75 7030
rect -45 7000 0 7030
rect -120 6960 0 7000
rect -120 6930 -75 6960
rect -45 6930 0 6960
rect -120 6895 0 6930
rect -120 6865 -75 6895
rect -45 6865 0 6895
rect -120 6835 0 6865
rect -120 6805 -75 6835
rect -45 6805 0 6835
rect -120 6770 0 6805
rect -120 6740 -75 6770
rect -45 6740 0 6770
rect -120 6700 0 6740
rect -120 6670 -75 6700
rect -45 6670 0 6700
rect -120 6630 0 6670
rect -120 6600 -75 6630
rect -45 6600 0 6630
rect -120 6560 0 6600
rect -120 6530 -75 6560
rect -45 6530 0 6560
rect -120 6495 0 6530
rect -120 6465 -75 6495
rect -45 6465 0 6495
rect -120 6210 0 6465
rect 230 9635 350 9650
rect 230 9605 275 9635
rect 305 9605 350 9635
rect 230 9570 350 9605
rect 230 9540 275 9570
rect 305 9540 350 9570
rect 230 9500 350 9540
rect 230 9470 275 9500
rect 305 9470 350 9500
rect 230 9430 350 9470
rect 230 9400 275 9430
rect 305 9400 350 9430
rect 230 9360 350 9400
rect 230 9330 275 9360
rect 305 9330 350 9360
rect 230 9295 350 9330
rect 230 9265 275 9295
rect 305 9265 350 9295
rect 230 9235 350 9265
rect 230 9205 275 9235
rect 305 9205 350 9235
rect 230 9170 350 9205
rect 230 9140 275 9170
rect 305 9140 350 9170
rect 230 9100 350 9140
rect 230 9070 275 9100
rect 305 9070 350 9100
rect 230 9030 350 9070
rect 230 9000 275 9030
rect 305 9000 350 9030
rect 230 8960 350 9000
rect 230 8930 275 8960
rect 305 8930 350 8960
rect 230 8895 350 8930
rect 230 8865 275 8895
rect 305 8865 350 8895
rect 230 8835 350 8865
rect 230 8805 275 8835
rect 305 8805 350 8835
rect 230 8770 350 8805
rect 230 8740 275 8770
rect 305 8740 350 8770
rect 230 8700 350 8740
rect 230 8670 275 8700
rect 305 8670 350 8700
rect 230 8630 350 8670
rect 230 8600 275 8630
rect 305 8600 350 8630
rect 230 8560 350 8600
rect 230 8530 275 8560
rect 305 8530 350 8560
rect 230 8495 350 8530
rect 230 8465 275 8495
rect 305 8465 350 8495
rect 230 8435 350 8465
rect 230 8405 275 8435
rect 305 8405 350 8435
rect 230 8370 350 8405
rect 230 8340 275 8370
rect 305 8340 350 8370
rect 230 8300 350 8340
rect 230 8270 275 8300
rect 305 8270 350 8300
rect 230 8230 350 8270
rect 230 8200 275 8230
rect 305 8200 350 8230
rect 230 8160 350 8200
rect 230 8130 275 8160
rect 305 8130 350 8160
rect 230 8095 350 8130
rect 230 8065 275 8095
rect 305 8065 350 8095
rect 230 8035 350 8065
rect 230 8005 275 8035
rect 305 8005 350 8035
rect 230 7970 350 8005
rect 230 7940 275 7970
rect 305 7940 350 7970
rect 230 7900 350 7940
rect 230 7870 275 7900
rect 305 7870 350 7900
rect 230 7830 350 7870
rect 230 7800 275 7830
rect 305 7800 350 7830
rect 230 7760 350 7800
rect 230 7730 275 7760
rect 305 7730 350 7760
rect 230 7695 350 7730
rect 230 7665 275 7695
rect 305 7665 350 7695
rect 230 7635 350 7665
rect 230 7605 275 7635
rect 305 7605 350 7635
rect 230 7570 350 7605
rect 230 7540 275 7570
rect 305 7540 350 7570
rect 230 7500 350 7540
rect 230 7470 275 7500
rect 305 7470 350 7500
rect 230 7430 350 7470
rect 230 7400 275 7430
rect 305 7400 350 7430
rect 230 7360 350 7400
rect 230 7330 275 7360
rect 305 7330 350 7360
rect 230 7295 350 7330
rect 230 7265 275 7295
rect 305 7265 350 7295
rect 230 7235 350 7265
rect 230 7205 275 7235
rect 305 7205 350 7235
rect 230 7170 350 7205
rect 230 7140 275 7170
rect 305 7140 350 7170
rect 230 7100 350 7140
rect 230 7070 275 7100
rect 305 7070 350 7100
rect 230 7030 350 7070
rect 230 7000 275 7030
rect 305 7000 350 7030
rect 230 6960 350 7000
rect 230 6930 275 6960
rect 305 6930 350 6960
rect 230 6895 350 6930
rect 230 6865 275 6895
rect 305 6865 350 6895
rect 230 6835 350 6865
rect 230 6805 275 6835
rect 305 6805 350 6835
rect 230 6770 350 6805
rect 230 6740 275 6770
rect 305 6740 350 6770
rect 230 6700 350 6740
rect 230 6670 275 6700
rect 305 6670 350 6700
rect 230 6630 350 6670
rect 230 6600 275 6630
rect 305 6600 350 6630
rect 230 6560 350 6600
rect 230 6530 275 6560
rect 305 6530 350 6560
rect 230 6495 350 6530
rect 230 6465 275 6495
rect 305 6465 350 6495
rect 230 6210 350 6465
rect 580 9635 700 9650
rect 580 9605 625 9635
rect 655 9605 700 9635
rect 580 9570 700 9605
rect 580 9540 625 9570
rect 655 9540 700 9570
rect 580 9500 700 9540
rect 580 9470 625 9500
rect 655 9470 700 9500
rect 580 9430 700 9470
rect 580 9400 625 9430
rect 655 9400 700 9430
rect 580 9360 700 9400
rect 580 9330 625 9360
rect 655 9330 700 9360
rect 580 9295 700 9330
rect 580 9265 625 9295
rect 655 9265 700 9295
rect 580 9235 700 9265
rect 580 9205 625 9235
rect 655 9205 700 9235
rect 580 9170 700 9205
rect 580 9140 625 9170
rect 655 9140 700 9170
rect 580 9100 700 9140
rect 580 9070 625 9100
rect 655 9070 700 9100
rect 580 9030 700 9070
rect 580 9000 625 9030
rect 655 9000 700 9030
rect 580 8960 700 9000
rect 580 8930 625 8960
rect 655 8930 700 8960
rect 580 8895 700 8930
rect 580 8865 625 8895
rect 655 8865 700 8895
rect 580 8835 700 8865
rect 580 8805 625 8835
rect 655 8805 700 8835
rect 580 8770 700 8805
rect 580 8740 625 8770
rect 655 8740 700 8770
rect 580 8700 700 8740
rect 580 8670 625 8700
rect 655 8670 700 8700
rect 580 8630 700 8670
rect 580 8600 625 8630
rect 655 8600 700 8630
rect 580 8560 700 8600
rect 580 8530 625 8560
rect 655 8530 700 8560
rect 580 8495 700 8530
rect 580 8465 625 8495
rect 655 8465 700 8495
rect 580 8435 700 8465
rect 580 8405 625 8435
rect 655 8405 700 8435
rect 580 8370 700 8405
rect 580 8340 625 8370
rect 655 8340 700 8370
rect 580 8300 700 8340
rect 580 8270 625 8300
rect 655 8270 700 8300
rect 580 8230 700 8270
rect 580 8200 625 8230
rect 655 8200 700 8230
rect 580 8160 700 8200
rect 580 8130 625 8160
rect 655 8130 700 8160
rect 580 8095 700 8130
rect 580 8065 625 8095
rect 655 8065 700 8095
rect 580 8035 700 8065
rect 580 8005 625 8035
rect 655 8005 700 8035
rect 580 7970 700 8005
rect 580 7940 625 7970
rect 655 7940 700 7970
rect 580 7900 700 7940
rect 580 7870 625 7900
rect 655 7870 700 7900
rect 580 7830 700 7870
rect 580 7800 625 7830
rect 655 7800 700 7830
rect 580 7760 700 7800
rect 580 7730 625 7760
rect 655 7730 700 7760
rect 580 7695 700 7730
rect 580 7665 625 7695
rect 655 7665 700 7695
rect 580 7635 700 7665
rect 580 7605 625 7635
rect 655 7605 700 7635
rect 580 7570 700 7605
rect 580 7540 625 7570
rect 655 7540 700 7570
rect 580 7500 700 7540
rect 580 7470 625 7500
rect 655 7470 700 7500
rect 580 7430 700 7470
rect 580 7400 625 7430
rect 655 7400 700 7430
rect 580 7360 700 7400
rect 580 7330 625 7360
rect 655 7330 700 7360
rect 580 7295 700 7330
rect 580 7265 625 7295
rect 655 7265 700 7295
rect 580 7235 700 7265
rect 580 7205 625 7235
rect 655 7205 700 7235
rect 580 7170 700 7205
rect 580 7140 625 7170
rect 655 7140 700 7170
rect 580 7100 700 7140
rect 580 7070 625 7100
rect 655 7070 700 7100
rect 580 7030 700 7070
rect 580 7000 625 7030
rect 655 7000 700 7030
rect 580 6960 700 7000
rect 580 6930 625 6960
rect 655 6930 700 6960
rect 580 6895 700 6930
rect 580 6865 625 6895
rect 655 6865 700 6895
rect 580 6835 700 6865
rect 580 6805 625 6835
rect 655 6805 700 6835
rect 580 6770 700 6805
rect 580 6740 625 6770
rect 655 6740 700 6770
rect 580 6700 700 6740
rect 580 6670 625 6700
rect 655 6670 700 6700
rect 580 6630 700 6670
rect 580 6600 625 6630
rect 655 6600 700 6630
rect 580 6560 700 6600
rect 580 6530 625 6560
rect 655 6530 700 6560
rect 580 6495 700 6530
rect 580 6465 625 6495
rect 655 6465 700 6495
rect 580 6210 700 6465
rect 930 9635 1050 9650
rect 930 9605 975 9635
rect 1005 9605 1050 9635
rect 930 9570 1050 9605
rect 930 9540 975 9570
rect 1005 9540 1050 9570
rect 930 9500 1050 9540
rect 930 9470 975 9500
rect 1005 9470 1050 9500
rect 930 9430 1050 9470
rect 930 9400 975 9430
rect 1005 9400 1050 9430
rect 930 9360 1050 9400
rect 930 9330 975 9360
rect 1005 9330 1050 9360
rect 930 9295 1050 9330
rect 930 9265 975 9295
rect 1005 9265 1050 9295
rect 930 9235 1050 9265
rect 930 9205 975 9235
rect 1005 9205 1050 9235
rect 930 9170 1050 9205
rect 930 9140 975 9170
rect 1005 9140 1050 9170
rect 930 9100 1050 9140
rect 930 9070 975 9100
rect 1005 9070 1050 9100
rect 930 9030 1050 9070
rect 930 9000 975 9030
rect 1005 9000 1050 9030
rect 930 8960 1050 9000
rect 930 8930 975 8960
rect 1005 8930 1050 8960
rect 930 8895 1050 8930
rect 930 8865 975 8895
rect 1005 8865 1050 8895
rect 930 8835 1050 8865
rect 930 8805 975 8835
rect 1005 8805 1050 8835
rect 930 8770 1050 8805
rect 930 8740 975 8770
rect 1005 8740 1050 8770
rect 930 8700 1050 8740
rect 930 8670 975 8700
rect 1005 8670 1050 8700
rect 930 8630 1050 8670
rect 930 8600 975 8630
rect 1005 8600 1050 8630
rect 930 8560 1050 8600
rect 930 8530 975 8560
rect 1005 8530 1050 8560
rect 930 8495 1050 8530
rect 930 8465 975 8495
rect 1005 8465 1050 8495
rect 930 8435 1050 8465
rect 930 8405 975 8435
rect 1005 8405 1050 8435
rect 930 8370 1050 8405
rect 930 8340 975 8370
rect 1005 8340 1050 8370
rect 930 8300 1050 8340
rect 930 8270 975 8300
rect 1005 8270 1050 8300
rect 930 8230 1050 8270
rect 930 8200 975 8230
rect 1005 8200 1050 8230
rect 930 8160 1050 8200
rect 930 8130 975 8160
rect 1005 8130 1050 8160
rect 930 8095 1050 8130
rect 930 8065 975 8095
rect 1005 8065 1050 8095
rect 930 8035 1050 8065
rect 930 8005 975 8035
rect 1005 8005 1050 8035
rect 930 7970 1050 8005
rect 930 7940 975 7970
rect 1005 7940 1050 7970
rect 930 7900 1050 7940
rect 930 7870 975 7900
rect 1005 7870 1050 7900
rect 930 7830 1050 7870
rect 930 7800 975 7830
rect 1005 7800 1050 7830
rect 930 7760 1050 7800
rect 930 7730 975 7760
rect 1005 7730 1050 7760
rect 930 7695 1050 7730
rect 930 7665 975 7695
rect 1005 7665 1050 7695
rect 930 7635 1050 7665
rect 930 7605 975 7635
rect 1005 7605 1050 7635
rect 930 7570 1050 7605
rect 930 7540 975 7570
rect 1005 7540 1050 7570
rect 930 7500 1050 7540
rect 930 7470 975 7500
rect 1005 7470 1050 7500
rect 930 7430 1050 7470
rect 930 7400 975 7430
rect 1005 7400 1050 7430
rect 930 7360 1050 7400
rect 930 7330 975 7360
rect 1005 7330 1050 7360
rect 930 7295 1050 7330
rect 930 7265 975 7295
rect 1005 7265 1050 7295
rect 930 7235 1050 7265
rect 930 7205 975 7235
rect 1005 7205 1050 7235
rect 930 7170 1050 7205
rect 930 7140 975 7170
rect 1005 7140 1050 7170
rect 930 7100 1050 7140
rect 930 7070 975 7100
rect 1005 7070 1050 7100
rect 930 7030 1050 7070
rect 930 7000 975 7030
rect 1005 7000 1050 7030
rect 930 6960 1050 7000
rect 930 6930 975 6960
rect 1005 6930 1050 6960
rect 930 6895 1050 6930
rect 930 6865 975 6895
rect 1005 6865 1050 6895
rect 930 6835 1050 6865
rect 930 6805 975 6835
rect 1005 6805 1050 6835
rect 930 6770 1050 6805
rect 930 6740 975 6770
rect 1005 6740 1050 6770
rect 930 6700 1050 6740
rect 930 6670 975 6700
rect 1005 6670 1050 6700
rect 930 6630 1050 6670
rect 930 6600 975 6630
rect 1005 6600 1050 6630
rect 930 6560 1050 6600
rect 930 6530 975 6560
rect 1005 6530 1050 6560
rect 930 6495 1050 6530
rect 930 6465 975 6495
rect 1005 6465 1050 6495
rect 930 6210 1050 6465
rect 1630 9635 1750 9650
rect 1630 9605 1675 9635
rect 1705 9605 1750 9635
rect 1630 9570 1750 9605
rect 1630 9540 1675 9570
rect 1705 9540 1750 9570
rect 1630 9500 1750 9540
rect 1630 9470 1675 9500
rect 1705 9470 1750 9500
rect 1630 9430 1750 9470
rect 1630 9400 1675 9430
rect 1705 9400 1750 9430
rect 1630 9360 1750 9400
rect 1630 9330 1675 9360
rect 1705 9330 1750 9360
rect 1630 9295 1750 9330
rect 1630 9265 1675 9295
rect 1705 9265 1750 9295
rect 1630 9235 1750 9265
rect 1630 9205 1675 9235
rect 1705 9205 1750 9235
rect 1630 9170 1750 9205
rect 1630 9140 1675 9170
rect 1705 9140 1750 9170
rect 1630 9100 1750 9140
rect 1630 9070 1675 9100
rect 1705 9070 1750 9100
rect 1630 9030 1750 9070
rect 1630 9000 1675 9030
rect 1705 9000 1750 9030
rect 1630 8960 1750 9000
rect 1630 8930 1675 8960
rect 1705 8930 1750 8960
rect 1630 8895 1750 8930
rect 1630 8865 1675 8895
rect 1705 8865 1750 8895
rect 1630 8835 1750 8865
rect 1630 8805 1675 8835
rect 1705 8805 1750 8835
rect 1630 8770 1750 8805
rect 1630 8740 1675 8770
rect 1705 8740 1750 8770
rect 1630 8700 1750 8740
rect 1630 8670 1675 8700
rect 1705 8670 1750 8700
rect 1630 8630 1750 8670
rect 1630 8600 1675 8630
rect 1705 8600 1750 8630
rect 1630 8560 1750 8600
rect 1630 8530 1675 8560
rect 1705 8530 1750 8560
rect 1630 8495 1750 8530
rect 1630 8465 1675 8495
rect 1705 8465 1750 8495
rect 1630 8435 1750 8465
rect 1630 8405 1675 8435
rect 1705 8405 1750 8435
rect 1630 8370 1750 8405
rect 1630 8340 1675 8370
rect 1705 8340 1750 8370
rect 1630 8300 1750 8340
rect 1630 8270 1675 8300
rect 1705 8270 1750 8300
rect 1630 8230 1750 8270
rect 1630 8200 1675 8230
rect 1705 8200 1750 8230
rect 1630 8160 1750 8200
rect 1630 8130 1675 8160
rect 1705 8130 1750 8160
rect 1630 8095 1750 8130
rect 1630 8065 1675 8095
rect 1705 8065 1750 8095
rect 1630 8035 1750 8065
rect 1630 8005 1675 8035
rect 1705 8005 1750 8035
rect 1630 7970 1750 8005
rect 1630 7940 1675 7970
rect 1705 7940 1750 7970
rect 1630 7900 1750 7940
rect 1630 7870 1675 7900
rect 1705 7870 1750 7900
rect 1630 7830 1750 7870
rect 1630 7800 1675 7830
rect 1705 7800 1750 7830
rect 1630 7760 1750 7800
rect 1630 7730 1675 7760
rect 1705 7730 1750 7760
rect 1630 7695 1750 7730
rect 1630 7665 1675 7695
rect 1705 7665 1750 7695
rect 1630 7635 1750 7665
rect 1630 7605 1675 7635
rect 1705 7605 1750 7635
rect 1630 7570 1750 7605
rect 1630 7540 1675 7570
rect 1705 7540 1750 7570
rect 1630 7500 1750 7540
rect 1630 7470 1675 7500
rect 1705 7470 1750 7500
rect 1630 7430 1750 7470
rect 1630 7400 1675 7430
rect 1705 7400 1750 7430
rect 1630 7360 1750 7400
rect 1630 7330 1675 7360
rect 1705 7330 1750 7360
rect 1630 7295 1750 7330
rect 1630 7265 1675 7295
rect 1705 7265 1750 7295
rect 1630 7235 1750 7265
rect 1630 7205 1675 7235
rect 1705 7205 1750 7235
rect 1630 7170 1750 7205
rect 1630 7140 1675 7170
rect 1705 7140 1750 7170
rect 1630 7100 1750 7140
rect 1630 7070 1675 7100
rect 1705 7070 1750 7100
rect 1630 7030 1750 7070
rect 1630 7000 1675 7030
rect 1705 7000 1750 7030
rect 1630 6960 1750 7000
rect 1630 6930 1675 6960
rect 1705 6930 1750 6960
rect 1630 6895 1750 6930
rect 1630 6865 1675 6895
rect 1705 6865 1750 6895
rect 1630 6835 1750 6865
rect 1630 6805 1675 6835
rect 1705 6805 1750 6835
rect 1630 6770 1750 6805
rect 1630 6740 1675 6770
rect 1705 6740 1750 6770
rect 1630 6700 1750 6740
rect 1630 6670 1675 6700
rect 1705 6670 1750 6700
rect 1630 6630 1750 6670
rect 1630 6600 1675 6630
rect 1705 6600 1750 6630
rect 1630 6560 1750 6600
rect 1630 6530 1675 6560
rect 1705 6530 1750 6560
rect 1630 6495 1750 6530
rect 1630 6465 1675 6495
rect 1705 6465 1750 6495
rect 1630 6210 1750 6465
rect 2205 9635 2325 15895
rect 6660 15595 6780 17725
rect 6660 15565 6665 15595
rect 6695 15565 6705 15595
rect 6735 15565 6745 15595
rect 6775 15565 6780 15595
rect 6660 15555 6780 15565
rect 6660 15525 6665 15555
rect 6695 15525 6705 15555
rect 6735 15525 6745 15555
rect 6775 15525 6780 15555
rect 6660 15515 6780 15525
rect 6660 15485 6665 15515
rect 6695 15485 6705 15515
rect 6735 15485 6745 15515
rect 6775 15485 6780 15515
rect 6660 12925 6780 15485
rect 6660 12895 6665 12925
rect 6695 12895 6705 12925
rect 6735 12895 6745 12925
rect 6775 12895 6780 12925
rect 6660 12885 6780 12895
rect 6660 12855 6665 12885
rect 6695 12855 6705 12885
rect 6735 12855 6745 12885
rect 6775 12855 6780 12885
rect 6660 12845 6780 12855
rect 6660 12815 6665 12845
rect 6695 12815 6705 12845
rect 6735 12815 6745 12845
rect 6775 12815 6780 12845
rect 6660 12810 6780 12815
rect 6660 12150 6780 12155
rect 6660 12120 6665 12150
rect 6695 12120 6705 12150
rect 6735 12120 6745 12150
rect 6775 12120 6780 12150
rect 6660 12110 6780 12120
rect 6660 12080 6665 12110
rect 6695 12080 6705 12110
rect 6735 12080 6745 12110
rect 6775 12080 6780 12110
rect 6660 12070 6780 12080
rect 6660 12040 6665 12070
rect 6695 12040 6705 12070
rect 6735 12040 6745 12070
rect 6775 12040 6780 12070
rect 6660 11165 6780 12040
rect 6660 11135 6665 11165
rect 6695 11135 6705 11165
rect 6735 11135 6745 11165
rect 6775 11135 6780 11165
rect 6660 11125 6780 11135
rect 6660 11095 6665 11125
rect 6695 11095 6705 11125
rect 6735 11095 6745 11125
rect 6775 11095 6780 11125
rect 6660 11085 6780 11095
rect 6660 11055 6665 11085
rect 6695 11055 6705 11085
rect 6735 11055 6745 11085
rect 6775 11055 6780 11085
rect 6660 10440 6780 11055
rect 6660 10410 6665 10440
rect 6695 10410 6705 10440
rect 6735 10410 6745 10440
rect 6775 10410 6780 10440
rect 6660 10400 6780 10410
rect 6660 10370 6665 10400
rect 6695 10370 6705 10400
rect 6735 10370 6745 10400
rect 6775 10370 6780 10400
rect 6660 10360 6780 10370
rect 6660 10330 6665 10360
rect 6695 10330 6705 10360
rect 6735 10330 6745 10360
rect 6775 10330 6780 10360
rect 2205 9605 2250 9635
rect 2280 9605 2325 9635
rect 2205 9570 2325 9605
rect 2205 9540 2250 9570
rect 2280 9540 2325 9570
rect 2205 9500 2325 9540
rect 2205 9470 2250 9500
rect 2280 9470 2325 9500
rect 2205 9430 2325 9470
rect 2205 9400 2250 9430
rect 2280 9400 2325 9430
rect 2205 9360 2325 9400
rect 2205 9330 2250 9360
rect 2280 9330 2325 9360
rect 2205 9295 2325 9330
rect 2205 9265 2250 9295
rect 2280 9265 2325 9295
rect 2205 9235 2325 9265
rect 2205 9205 2250 9235
rect 2280 9205 2325 9235
rect 2205 9170 2325 9205
rect 2205 9140 2250 9170
rect 2280 9140 2325 9170
rect 2205 9100 2325 9140
rect 2205 9070 2250 9100
rect 2280 9070 2325 9100
rect 2205 9030 2325 9070
rect 2205 9000 2250 9030
rect 2280 9000 2325 9030
rect 2205 8960 2325 9000
rect 2205 8930 2250 8960
rect 2280 8930 2325 8960
rect 2205 8895 2325 8930
rect 2205 8865 2250 8895
rect 2280 8865 2325 8895
rect 2205 8835 2325 8865
rect 2205 8805 2250 8835
rect 2280 8805 2325 8835
rect 2205 8770 2325 8805
rect 2205 8740 2250 8770
rect 2280 8740 2325 8770
rect 2205 8700 2325 8740
rect 2205 8670 2250 8700
rect 2280 8670 2325 8700
rect 2205 8630 2325 8670
rect 2205 8600 2250 8630
rect 2280 8600 2325 8630
rect 2205 8560 2325 8600
rect 2205 8530 2250 8560
rect 2280 8530 2325 8560
rect 2205 8495 2325 8530
rect 2205 8465 2250 8495
rect 2280 8465 2325 8495
rect 2205 8435 2325 8465
rect 2205 8405 2250 8435
rect 2280 8405 2325 8435
rect 2205 8370 2325 8405
rect 2205 8340 2250 8370
rect 2280 8340 2325 8370
rect 2205 8300 2325 8340
rect 2205 8270 2250 8300
rect 2280 8270 2325 8300
rect 2205 8230 2325 8270
rect 2205 8200 2250 8230
rect 2280 8200 2325 8230
rect 2205 8160 2325 8200
rect 2205 8130 2250 8160
rect 2280 8130 2325 8160
rect 2205 8095 2325 8130
rect 2205 8065 2250 8095
rect 2280 8065 2325 8095
rect 2205 8035 2325 8065
rect 2205 8005 2250 8035
rect 2280 8005 2325 8035
rect 2205 7970 2325 8005
rect 2205 7940 2250 7970
rect 2280 7940 2325 7970
rect 2205 7900 2325 7940
rect 2205 7870 2250 7900
rect 2280 7870 2325 7900
rect 2205 7830 2325 7870
rect 2205 7800 2250 7830
rect 2280 7800 2325 7830
rect 2205 7760 2325 7800
rect 2205 7730 2250 7760
rect 2280 7730 2325 7760
rect 2205 7695 2325 7730
rect 2205 7665 2250 7695
rect 2280 7665 2325 7695
rect 2205 7635 2325 7665
rect 2205 7605 2250 7635
rect 2280 7605 2325 7635
rect 2205 7570 2325 7605
rect 2205 7540 2250 7570
rect 2280 7540 2325 7570
rect 2205 7500 2325 7540
rect 2205 7470 2250 7500
rect 2280 7470 2325 7500
rect 2205 7430 2325 7470
rect 2205 7400 2250 7430
rect 2280 7400 2325 7430
rect 2205 7360 2325 7400
rect 2205 7330 2250 7360
rect 2280 7330 2325 7360
rect 2205 7295 2325 7330
rect 2205 7265 2250 7295
rect 2280 7265 2325 7295
rect 2205 7235 2325 7265
rect 2205 7205 2250 7235
rect 2280 7205 2325 7235
rect 2205 7170 2325 7205
rect 2205 7140 2250 7170
rect 2280 7140 2325 7170
rect 2205 7100 2325 7140
rect 2205 7070 2250 7100
rect 2280 7070 2325 7100
rect 2205 7030 2325 7070
rect 2205 7000 2250 7030
rect 2280 7000 2325 7030
rect 2205 6960 2325 7000
rect 2205 6930 2250 6960
rect 2280 6930 2325 6960
rect 2205 6895 2325 6930
rect 2205 6865 2250 6895
rect 2280 6865 2325 6895
rect 2205 6835 2325 6865
rect 2205 6805 2250 6835
rect 2280 6805 2325 6835
rect 2205 6770 2325 6805
rect 2205 6740 2250 6770
rect 2280 6740 2325 6770
rect 2205 6700 2325 6740
rect 2205 6670 2250 6700
rect 2280 6670 2325 6700
rect 2205 6630 2325 6670
rect 2205 6600 2250 6630
rect 2280 6600 2325 6630
rect 2205 6560 2325 6600
rect 2205 6530 2250 6560
rect 2280 6530 2325 6560
rect 2205 6495 2325 6530
rect 2205 6465 2250 6495
rect 2280 6465 2325 6495
rect 2205 6450 2325 6465
rect 2485 6435 2505 9735
rect 2045 6430 2085 6435
rect 2045 6400 2050 6430
rect 2080 6400 2085 6430
rect 2045 6395 2085 6400
rect 2475 6430 2515 6435
rect 2475 6400 2480 6430
rect 2510 6400 2515 6430
rect 2475 6395 2515 6400
rect 2000 6375 2040 6380
rect 2000 6345 2005 6375
rect 2035 6345 2040 6375
rect 2000 6340 2040 6345
rect 1280 6205 1400 6210
rect 1280 6175 1285 6205
rect 1315 6175 1325 6205
rect 1355 6175 1365 6205
rect 1395 6175 1400 6205
rect 1280 6165 1400 6175
rect 1280 6135 1285 6165
rect 1315 6135 1325 6165
rect 1355 6135 1365 6165
rect 1395 6135 1400 6165
rect 1280 6125 1400 6135
rect 1280 6095 1285 6125
rect 1315 6095 1325 6125
rect 1355 6095 1365 6125
rect 1395 6095 1400 6125
rect 1280 1160 1400 6095
rect 2010 2265 2030 6340
rect 2055 2320 2075 6395
rect 2725 6335 2745 9735
rect 2855 6435 2875 9735
rect 3175 9650 3215 10325
rect 3235 9650 3275 10325
rect 3165 9635 3280 9650
rect 3165 9605 3180 9635
rect 3210 9605 3240 9635
rect 3270 9605 3280 9635
rect 3165 9570 3280 9605
rect 3165 9540 3180 9570
rect 3210 9540 3240 9570
rect 3270 9540 3280 9570
rect 3165 9500 3280 9540
rect 3165 9470 3180 9500
rect 3210 9470 3240 9500
rect 3270 9470 3280 9500
rect 3165 9430 3280 9470
rect 3165 9400 3180 9430
rect 3210 9400 3240 9430
rect 3270 9400 3280 9430
rect 3165 9360 3280 9400
rect 3165 9330 3180 9360
rect 3210 9330 3240 9360
rect 3270 9330 3280 9360
rect 3165 9295 3280 9330
rect 3165 9265 3180 9295
rect 3210 9265 3240 9295
rect 3270 9265 3280 9295
rect 3165 9235 3280 9265
rect 3165 9205 3180 9235
rect 3210 9205 3240 9235
rect 3270 9205 3280 9235
rect 3165 9170 3280 9205
rect 3165 9140 3180 9170
rect 3210 9140 3240 9170
rect 3270 9140 3280 9170
rect 3165 9100 3280 9140
rect 3165 9070 3180 9100
rect 3210 9070 3240 9100
rect 3270 9070 3280 9100
rect 3165 9030 3280 9070
rect 3165 9000 3180 9030
rect 3210 9000 3240 9030
rect 3270 9000 3280 9030
rect 3165 8960 3280 9000
rect 3165 8930 3180 8960
rect 3210 8930 3240 8960
rect 3270 8930 3280 8960
rect 3165 8895 3280 8930
rect 3165 8865 3180 8895
rect 3210 8865 3240 8895
rect 3270 8865 3280 8895
rect 3165 8835 3280 8865
rect 3165 8805 3180 8835
rect 3210 8805 3240 8835
rect 3270 8805 3280 8835
rect 3165 8770 3280 8805
rect 3165 8740 3180 8770
rect 3210 8740 3240 8770
rect 3270 8740 3280 8770
rect 3165 8700 3280 8740
rect 3165 8670 3180 8700
rect 3210 8670 3240 8700
rect 3270 8670 3280 8700
rect 3165 8630 3280 8670
rect 3165 8600 3180 8630
rect 3210 8600 3240 8630
rect 3270 8600 3280 8630
rect 3165 8560 3280 8600
rect 3165 8530 3180 8560
rect 3210 8530 3240 8560
rect 3270 8530 3280 8560
rect 3165 8495 3280 8530
rect 3165 8465 3180 8495
rect 3210 8465 3240 8495
rect 3270 8465 3280 8495
rect 3165 8435 3280 8465
rect 3165 8405 3180 8435
rect 3210 8405 3240 8435
rect 3270 8405 3280 8435
rect 3165 8370 3280 8405
rect 3165 8340 3180 8370
rect 3210 8340 3240 8370
rect 3270 8340 3280 8370
rect 3165 8300 3280 8340
rect 3165 8270 3180 8300
rect 3210 8270 3240 8300
rect 3270 8270 3280 8300
rect 3165 8230 3280 8270
rect 3165 8200 3180 8230
rect 3210 8200 3240 8230
rect 3270 8200 3280 8230
rect 3165 8160 3280 8200
rect 3165 8130 3180 8160
rect 3210 8130 3240 8160
rect 3270 8130 3280 8160
rect 3165 8095 3280 8130
rect 3165 8065 3180 8095
rect 3210 8065 3240 8095
rect 3270 8065 3280 8095
rect 3165 8035 3280 8065
rect 3165 8005 3180 8035
rect 3210 8005 3240 8035
rect 3270 8005 3280 8035
rect 3165 7970 3280 8005
rect 3165 7940 3180 7970
rect 3210 7940 3240 7970
rect 3270 7940 3280 7970
rect 3165 7900 3280 7940
rect 3165 7870 3180 7900
rect 3210 7870 3240 7900
rect 3270 7870 3280 7900
rect 3165 7830 3280 7870
rect 3165 7800 3180 7830
rect 3210 7800 3240 7830
rect 3270 7800 3280 7830
rect 3165 7760 3280 7800
rect 3165 7730 3180 7760
rect 3210 7730 3240 7760
rect 3270 7730 3280 7760
rect 3165 7695 3280 7730
rect 3165 7665 3180 7695
rect 3210 7665 3240 7695
rect 3270 7665 3280 7695
rect 3165 7635 3280 7665
rect 3165 7605 3180 7635
rect 3210 7605 3240 7635
rect 3270 7605 3280 7635
rect 3165 7570 3280 7605
rect 3165 7540 3180 7570
rect 3210 7540 3240 7570
rect 3270 7540 3280 7570
rect 3165 7500 3280 7540
rect 3165 7470 3180 7500
rect 3210 7470 3240 7500
rect 3270 7470 3280 7500
rect 3165 7430 3280 7470
rect 3165 7400 3180 7430
rect 3210 7400 3240 7430
rect 3270 7400 3280 7430
rect 3165 7360 3280 7400
rect 3165 7330 3180 7360
rect 3210 7330 3240 7360
rect 3270 7330 3280 7360
rect 3165 7295 3280 7330
rect 3165 7265 3180 7295
rect 3210 7265 3240 7295
rect 3270 7265 3280 7295
rect 3165 7235 3280 7265
rect 3165 7205 3180 7235
rect 3210 7205 3240 7235
rect 3270 7205 3280 7235
rect 3165 7170 3280 7205
rect 3165 7140 3180 7170
rect 3210 7140 3240 7170
rect 3270 7140 3280 7170
rect 3165 7100 3280 7140
rect 3165 7070 3180 7100
rect 3210 7070 3240 7100
rect 3270 7070 3280 7100
rect 3165 7030 3280 7070
rect 3165 7000 3180 7030
rect 3210 7000 3240 7030
rect 3270 7000 3280 7030
rect 3165 6960 3280 7000
rect 3165 6930 3180 6960
rect 3210 6930 3240 6960
rect 3270 6930 3280 6960
rect 3165 6895 3280 6930
rect 3165 6865 3180 6895
rect 3210 6865 3240 6895
rect 3270 6865 3280 6895
rect 3165 6835 3280 6865
rect 3165 6805 3180 6835
rect 3210 6805 3240 6835
rect 3270 6805 3280 6835
rect 3165 6770 3280 6805
rect 3165 6740 3180 6770
rect 3210 6740 3240 6770
rect 3270 6740 3280 6770
rect 3165 6700 3280 6740
rect 3165 6670 3180 6700
rect 3210 6670 3240 6700
rect 3270 6670 3280 6700
rect 3165 6630 3280 6670
rect 3165 6600 3180 6630
rect 3210 6600 3240 6630
rect 3270 6600 3280 6630
rect 3165 6560 3280 6600
rect 3165 6530 3180 6560
rect 3210 6530 3240 6560
rect 3270 6530 3280 6560
rect 3165 6495 3280 6530
rect 3165 6465 3180 6495
rect 3210 6465 3240 6495
rect 3270 6465 3280 6495
rect 3165 6450 3280 6465
rect 2845 6430 2885 6435
rect 2845 6400 2850 6430
rect 2880 6400 2885 6430
rect 2845 6395 2885 6400
rect 2715 6330 2755 6335
rect 2715 6300 2720 6330
rect 2750 6300 2755 6330
rect 2715 6295 2755 6300
rect 3075 6330 3115 6335
rect 3075 6300 3080 6330
rect 3110 6300 3115 6330
rect 3295 6320 3325 9740
rect 3345 9650 3385 10325
rect 6660 10080 6780 10330
rect 6660 10050 6665 10080
rect 6695 10050 6705 10080
rect 6735 10050 6745 10080
rect 6775 10050 6780 10080
rect 6660 10040 6780 10050
rect 6660 10010 6665 10040
rect 6695 10010 6705 10040
rect 6735 10010 6745 10040
rect 6775 10010 6780 10040
rect 6660 10000 6780 10010
rect 6660 9970 6665 10000
rect 6695 9970 6705 10000
rect 6735 9970 6745 10000
rect 6775 9970 6780 10000
rect 3740 9910 3780 9920
rect 3340 9635 3395 9650
rect 3340 9605 3350 9635
rect 3380 9605 3395 9635
rect 3340 9570 3395 9605
rect 3340 9540 3350 9570
rect 3380 9540 3395 9570
rect 3340 9500 3395 9540
rect 3340 9470 3350 9500
rect 3380 9470 3395 9500
rect 3340 9430 3395 9470
rect 3340 9400 3350 9430
rect 3380 9400 3395 9430
rect 3340 9360 3395 9400
rect 3340 9330 3350 9360
rect 3380 9330 3395 9360
rect 3340 9295 3395 9330
rect 3340 9265 3350 9295
rect 3380 9265 3395 9295
rect 3340 9235 3395 9265
rect 3340 9205 3350 9235
rect 3380 9205 3395 9235
rect 3340 9170 3395 9205
rect 3340 9140 3350 9170
rect 3380 9140 3395 9170
rect 3340 9100 3395 9140
rect 3340 9070 3350 9100
rect 3380 9070 3395 9100
rect 3340 9030 3395 9070
rect 3340 9000 3350 9030
rect 3380 9000 3395 9030
rect 3340 8960 3395 9000
rect 3340 8930 3350 8960
rect 3380 8930 3395 8960
rect 3340 8895 3395 8930
rect 3340 8865 3350 8895
rect 3380 8865 3395 8895
rect 3340 8835 3395 8865
rect 3340 8805 3350 8835
rect 3380 8805 3395 8835
rect 3340 8770 3395 8805
rect 3340 8740 3350 8770
rect 3380 8740 3395 8770
rect 3340 8700 3395 8740
rect 3340 8670 3350 8700
rect 3380 8670 3395 8700
rect 3340 8630 3395 8670
rect 3340 8600 3350 8630
rect 3380 8600 3395 8630
rect 3340 8560 3395 8600
rect 3340 8530 3350 8560
rect 3380 8530 3395 8560
rect 3340 8495 3395 8530
rect 3340 8465 3350 8495
rect 3380 8465 3395 8495
rect 3340 8435 3395 8465
rect 3340 8405 3350 8435
rect 3380 8405 3395 8435
rect 3340 8370 3395 8405
rect 3340 8340 3350 8370
rect 3380 8340 3395 8370
rect 3340 8300 3395 8340
rect 3340 8270 3350 8300
rect 3380 8270 3395 8300
rect 3340 8230 3395 8270
rect 3340 8200 3350 8230
rect 3380 8200 3395 8230
rect 3340 8160 3395 8200
rect 3340 8130 3350 8160
rect 3380 8130 3395 8160
rect 3340 8095 3395 8130
rect 3340 8065 3350 8095
rect 3380 8065 3395 8095
rect 3340 8035 3395 8065
rect 3340 8005 3350 8035
rect 3380 8005 3395 8035
rect 3340 7970 3395 8005
rect 3340 7940 3350 7970
rect 3380 7940 3395 7970
rect 3340 7900 3395 7940
rect 3340 7870 3350 7900
rect 3380 7870 3395 7900
rect 3340 7830 3395 7870
rect 3340 7800 3350 7830
rect 3380 7800 3395 7830
rect 3340 7760 3395 7800
rect 3340 7730 3350 7760
rect 3380 7730 3395 7760
rect 3340 7695 3395 7730
rect 3340 7665 3350 7695
rect 3380 7665 3395 7695
rect 3340 7635 3395 7665
rect 3340 7605 3350 7635
rect 3380 7605 3395 7635
rect 3340 7570 3395 7605
rect 3340 7540 3350 7570
rect 3380 7540 3395 7570
rect 3340 7500 3395 7540
rect 3340 7470 3350 7500
rect 3380 7470 3395 7500
rect 3340 7430 3395 7470
rect 3340 7400 3350 7430
rect 3380 7400 3395 7430
rect 3340 7360 3395 7400
rect 3340 7330 3350 7360
rect 3380 7330 3395 7360
rect 3340 7295 3395 7330
rect 3340 7265 3350 7295
rect 3380 7265 3395 7295
rect 3340 7235 3395 7265
rect 3340 7205 3350 7235
rect 3380 7205 3395 7235
rect 3340 7170 3395 7205
rect 3340 7140 3350 7170
rect 3380 7140 3395 7170
rect 3340 7100 3395 7140
rect 3340 7070 3350 7100
rect 3380 7070 3395 7100
rect 3340 7030 3395 7070
rect 3340 7000 3350 7030
rect 3380 7000 3395 7030
rect 3640 7010 3660 9740
rect 3340 6960 3395 7000
rect 3340 6930 3350 6960
rect 3380 6930 3395 6960
rect 3340 6895 3395 6930
rect 3340 6865 3350 6895
rect 3380 6865 3395 6895
rect 3340 6835 3395 6865
rect 3340 6805 3350 6835
rect 3380 6805 3395 6835
rect 3340 6770 3395 6805
rect 3340 6740 3350 6770
rect 3380 6740 3395 6770
rect 3340 6700 3395 6740
rect 3340 6670 3350 6700
rect 3380 6670 3395 6700
rect 3340 6630 3395 6670
rect 3340 6600 3350 6630
rect 3380 6600 3395 6630
rect 3340 6560 3395 6600
rect 3340 6530 3350 6560
rect 3380 6530 3395 6560
rect 3340 6495 3395 6530
rect 3340 6465 3350 6495
rect 3380 6465 3395 6495
rect 3340 6450 3395 6465
rect 3380 6430 3420 6435
rect 3380 6400 3385 6430
rect 3415 6400 3420 6430
rect 3380 6395 3420 6400
rect 3075 6295 3115 6300
rect 3290 6315 3330 6320
rect 3085 5095 3105 6295
rect 3290 6285 3295 6315
rect 3325 6285 3330 6315
rect 3290 6280 3330 6285
rect 3075 5090 3115 5095
rect 3075 5060 3080 5090
rect 3110 5060 3115 5090
rect 3075 5055 3115 5060
rect 3390 3810 3410 6395
rect 3630 6375 3670 7010
rect 3630 6345 3635 6375
rect 3665 6345 3670 6375
rect 3630 6340 3670 6345
rect 3435 6260 3475 6265
rect 3435 6230 3440 6260
rect 3470 6230 3475 6260
rect 3380 3805 3420 3810
rect 3380 3775 3385 3805
rect 3415 3775 3420 3805
rect 3380 3770 3420 3775
rect 3435 3125 3475 6230
rect 4310 6205 4340 9740
rect 4310 6165 4340 6175
rect 4310 6125 4340 6135
rect 4310 6090 4340 6095
rect 4420 6205 4450 9740
rect 4470 6315 4510 6320
rect 4470 6285 4475 6315
rect 4505 6285 4510 6315
rect 4470 6260 4510 6285
rect 4470 6230 4475 6260
rect 4505 6230 4510 6260
rect 4470 6225 4510 6230
rect 4420 6165 4450 6175
rect 4420 6125 4450 6135
rect 4420 6090 4450 6095
rect 4530 6205 4560 9740
rect 4530 6165 4560 6175
rect 4530 6125 4560 6135
rect 4530 6090 4560 6095
rect 4640 6205 4670 9740
rect 5320 6380 5340 9740
rect 6155 6435 6175 9740
rect 5470 6430 5510 6435
rect 5470 6400 5475 6430
rect 5505 6400 5510 6430
rect 5470 6395 5510 6400
rect 6145 6430 6185 6435
rect 6145 6400 6150 6430
rect 6180 6400 6185 6430
rect 6145 6395 6185 6400
rect 5310 6375 5350 6380
rect 5310 6345 5315 6375
rect 5345 6345 5350 6375
rect 5310 6340 5350 6345
rect 4640 6165 4670 6175
rect 4640 6125 4670 6135
rect 4640 6090 4670 6095
rect 5480 3870 5500 6395
rect 5520 6260 5560 6265
rect 5520 6230 5525 6260
rect 5555 6230 5560 6260
rect 5475 3865 5505 3870
rect 5475 3830 5505 3835
rect 3435 3095 3440 3125
rect 3470 3095 3475 3125
rect 3435 3090 3475 3095
rect 4470 3125 4510 3130
rect 4470 3095 4475 3125
rect 4505 3095 4510 3125
rect 4470 3015 4510 3095
rect 5520 3125 5560 6230
rect 6230 5440 6250 9740
rect 6475 6435 6500 9740
rect 6660 9570 6780 9970
rect 6660 9540 6705 9570
rect 6735 9540 6780 9570
rect 6660 9500 6780 9540
rect 6660 9470 6705 9500
rect 6735 9470 6780 9500
rect 6660 9430 6780 9470
rect 6660 9400 6705 9430
rect 6735 9400 6780 9430
rect 6660 9360 6780 9400
rect 6660 9330 6705 9360
rect 6735 9330 6780 9360
rect 6660 9295 6780 9330
rect 6660 9265 6705 9295
rect 6735 9265 6780 9295
rect 6660 9235 6780 9265
rect 6660 9205 6705 9235
rect 6735 9205 6780 9235
rect 6660 9170 6780 9205
rect 6660 9140 6705 9170
rect 6735 9140 6780 9170
rect 6660 9100 6780 9140
rect 6660 9070 6705 9100
rect 6735 9070 6780 9100
rect 6660 9030 6780 9070
rect 6660 9000 6705 9030
rect 6735 9000 6780 9030
rect 6660 8960 6780 9000
rect 6660 8930 6705 8960
rect 6735 8930 6780 8960
rect 6660 8895 6780 8930
rect 6660 8865 6705 8895
rect 6735 8865 6780 8895
rect 6660 8835 6780 8865
rect 6660 8805 6705 8835
rect 6735 8805 6780 8835
rect 6660 8770 6780 8805
rect 6660 8740 6705 8770
rect 6735 8740 6780 8770
rect 6660 8700 6780 8740
rect 6660 8670 6705 8700
rect 6735 8670 6780 8700
rect 6660 8630 6780 8670
rect 6660 8600 6705 8630
rect 6735 8600 6780 8630
rect 6660 8560 6780 8600
rect 6660 8530 6705 8560
rect 6735 8530 6780 8560
rect 6660 8495 6780 8530
rect 6660 8465 6705 8495
rect 6735 8465 6780 8495
rect 6660 8435 6780 8465
rect 6660 8405 6705 8435
rect 6735 8405 6780 8435
rect 6660 8370 6780 8405
rect 6660 8340 6705 8370
rect 6735 8340 6780 8370
rect 6660 8300 6780 8340
rect 6660 8270 6705 8300
rect 6735 8270 6780 8300
rect 6660 8230 6780 8270
rect 6660 8200 6705 8230
rect 6735 8200 6780 8230
rect 6660 8160 6780 8200
rect 6660 8130 6705 8160
rect 6735 8130 6780 8160
rect 6660 8095 6780 8130
rect 6660 8065 6705 8095
rect 6735 8065 6780 8095
rect 6660 8035 6780 8065
rect 6660 8005 6705 8035
rect 6735 8005 6780 8035
rect 6660 7970 6780 8005
rect 6660 7940 6705 7970
rect 6735 7940 6780 7970
rect 6660 7900 6780 7940
rect 6660 7870 6705 7900
rect 6735 7870 6780 7900
rect 6660 7830 6780 7870
rect 6660 7800 6705 7830
rect 6735 7800 6780 7830
rect 6660 7760 6780 7800
rect 6660 7730 6705 7760
rect 6735 7730 6780 7760
rect 6660 7695 6780 7730
rect 6660 7665 6705 7695
rect 6735 7665 6780 7695
rect 6660 7635 6780 7665
rect 6660 7605 6705 7635
rect 6735 7605 6780 7635
rect 6660 7570 6780 7605
rect 6660 7540 6705 7570
rect 6735 7540 6780 7570
rect 6660 7500 6780 7540
rect 6660 7470 6705 7500
rect 6735 7470 6780 7500
rect 6660 7430 6780 7470
rect 6660 7400 6705 7430
rect 6735 7400 6780 7430
rect 6660 7360 6780 7400
rect 6660 7330 6705 7360
rect 6735 7330 6780 7360
rect 6660 7295 6780 7330
rect 6660 7265 6705 7295
rect 6735 7265 6780 7295
rect 6660 7235 6780 7265
rect 6660 7205 6705 7235
rect 6735 7205 6780 7235
rect 6660 7170 6780 7205
rect 6660 7140 6705 7170
rect 6735 7140 6780 7170
rect 6660 7100 6780 7140
rect 6660 7070 6705 7100
rect 6735 7070 6780 7100
rect 6660 7030 6780 7070
rect 6660 7000 6705 7030
rect 6735 7000 6780 7030
rect 6660 6960 6780 7000
rect 6660 6930 6705 6960
rect 6735 6930 6780 6960
rect 6660 6895 6780 6930
rect 6660 6865 6705 6895
rect 6735 6865 6780 6895
rect 6660 6835 6780 6865
rect 6660 6805 6705 6835
rect 6735 6805 6780 6835
rect 6660 6770 6780 6805
rect 6660 6740 6705 6770
rect 6735 6740 6780 6770
rect 6660 6700 6780 6740
rect 6660 6670 6705 6700
rect 6735 6670 6780 6700
rect 6660 6630 6780 6670
rect 6660 6600 6705 6630
rect 6735 6600 6780 6630
rect 6660 6560 6780 6600
rect 6660 6530 6705 6560
rect 6735 6530 6780 6560
rect 6660 6495 6780 6530
rect 6660 6465 6705 6495
rect 6735 6465 6780 6495
rect 6660 6450 6780 6465
rect 7230 9635 7350 9650
rect 7230 9605 7275 9635
rect 7305 9605 7350 9635
rect 7230 9570 7350 9605
rect 7230 9540 7275 9570
rect 7305 9540 7350 9570
rect 7230 9500 7350 9540
rect 7230 9470 7275 9500
rect 7305 9470 7350 9500
rect 7230 9430 7350 9470
rect 7230 9400 7275 9430
rect 7305 9400 7350 9430
rect 7230 9360 7350 9400
rect 7230 9330 7275 9360
rect 7305 9330 7350 9360
rect 7230 9295 7350 9330
rect 7230 9265 7275 9295
rect 7305 9265 7350 9295
rect 7230 9235 7350 9265
rect 7230 9205 7275 9235
rect 7305 9205 7350 9235
rect 7230 9170 7350 9205
rect 7230 9140 7275 9170
rect 7305 9140 7350 9170
rect 7230 9100 7350 9140
rect 7230 9070 7275 9100
rect 7305 9070 7350 9100
rect 7230 9030 7350 9070
rect 7230 9000 7275 9030
rect 7305 9000 7350 9030
rect 7230 8960 7350 9000
rect 7230 8930 7275 8960
rect 7305 8930 7350 8960
rect 7230 8895 7350 8930
rect 7230 8865 7275 8895
rect 7305 8865 7350 8895
rect 7230 8835 7350 8865
rect 7230 8805 7275 8835
rect 7305 8805 7350 8835
rect 7230 8770 7350 8805
rect 7230 8740 7275 8770
rect 7305 8740 7350 8770
rect 7230 8700 7350 8740
rect 7230 8670 7275 8700
rect 7305 8670 7350 8700
rect 7230 8630 7350 8670
rect 7230 8600 7275 8630
rect 7305 8600 7350 8630
rect 7230 8560 7350 8600
rect 7230 8530 7275 8560
rect 7305 8530 7350 8560
rect 7230 8495 7350 8530
rect 7230 8465 7275 8495
rect 7305 8465 7350 8495
rect 7230 8435 7350 8465
rect 7230 8405 7275 8435
rect 7305 8405 7350 8435
rect 7230 8370 7350 8405
rect 7230 8340 7275 8370
rect 7305 8340 7350 8370
rect 7230 8300 7350 8340
rect 7230 8270 7275 8300
rect 7305 8270 7350 8300
rect 7230 8230 7350 8270
rect 7230 8200 7275 8230
rect 7305 8200 7350 8230
rect 7230 8160 7350 8200
rect 7230 8130 7275 8160
rect 7305 8130 7350 8160
rect 7230 8095 7350 8130
rect 7230 8065 7275 8095
rect 7305 8065 7350 8095
rect 7230 8035 7350 8065
rect 7230 8005 7275 8035
rect 7305 8005 7350 8035
rect 7230 7970 7350 8005
rect 7230 7940 7275 7970
rect 7305 7940 7350 7970
rect 7230 7900 7350 7940
rect 7230 7870 7275 7900
rect 7305 7870 7350 7900
rect 7230 7830 7350 7870
rect 7230 7800 7275 7830
rect 7305 7800 7350 7830
rect 7230 7760 7350 7800
rect 7230 7730 7275 7760
rect 7305 7730 7350 7760
rect 7230 7695 7350 7730
rect 7230 7665 7275 7695
rect 7305 7665 7350 7695
rect 7230 7635 7350 7665
rect 7230 7605 7275 7635
rect 7305 7605 7350 7635
rect 7230 7570 7350 7605
rect 7230 7540 7275 7570
rect 7305 7540 7350 7570
rect 7230 7500 7350 7540
rect 7230 7470 7275 7500
rect 7305 7470 7350 7500
rect 7230 7430 7350 7470
rect 7230 7400 7275 7430
rect 7305 7400 7350 7430
rect 7230 7360 7350 7400
rect 7230 7330 7275 7360
rect 7305 7330 7350 7360
rect 7230 7295 7350 7330
rect 7230 7265 7275 7295
rect 7305 7265 7350 7295
rect 7230 7235 7350 7265
rect 7230 7205 7275 7235
rect 7305 7205 7350 7235
rect 7230 7170 7350 7205
rect 7230 7140 7275 7170
rect 7305 7140 7350 7170
rect 7230 7100 7350 7140
rect 7230 7070 7275 7100
rect 7305 7070 7350 7100
rect 7230 7030 7350 7070
rect 7230 7000 7275 7030
rect 7305 7000 7350 7030
rect 7230 6960 7350 7000
rect 7230 6930 7275 6960
rect 7305 6930 7350 6960
rect 7230 6895 7350 6930
rect 7230 6865 7275 6895
rect 7305 6865 7350 6895
rect 7230 6835 7350 6865
rect 7230 6805 7275 6835
rect 7305 6805 7350 6835
rect 7230 6770 7350 6805
rect 7230 6740 7275 6770
rect 7305 6740 7350 6770
rect 7230 6700 7350 6740
rect 7230 6670 7275 6700
rect 7305 6670 7350 6700
rect 7230 6630 7350 6670
rect 7230 6600 7275 6630
rect 7305 6600 7350 6630
rect 7230 6560 7350 6600
rect 7230 6530 7275 6560
rect 7305 6530 7350 6560
rect 7230 6495 7350 6530
rect 7230 6465 7275 6495
rect 7305 6465 7350 6495
rect 6465 6430 6505 6435
rect 6465 6400 6470 6430
rect 6500 6400 6505 6430
rect 6465 6395 6505 6400
rect 6895 6430 6935 6435
rect 6895 6400 6900 6430
rect 6930 6400 6935 6430
rect 6895 6395 6935 6400
rect 5575 5435 5605 5440
rect 5575 5400 5605 5405
rect 6220 5435 6260 5440
rect 6220 5405 6225 5435
rect 6255 5405 6260 5435
rect 6220 5400 6260 5405
rect 5580 4445 5600 5400
rect 5575 4440 5605 4445
rect 5575 4405 5605 4410
rect 5520 3095 5525 3125
rect 5555 3095 5560 3125
rect 5520 3090 5560 3095
rect 4470 2985 4475 3015
rect 4505 2985 4510 3015
rect 4470 2980 4510 2985
rect 6905 2320 6925 6395
rect 6940 6375 6980 6380
rect 6940 6345 6945 6375
rect 6975 6345 6980 6375
rect 6940 6340 6980 6345
rect 2045 2315 2085 2320
rect 2045 2285 2050 2315
rect 2080 2285 2085 2315
rect 2045 2280 2085 2285
rect 2120 2315 2160 2320
rect 2120 2285 2125 2315
rect 2155 2285 2160 2315
rect 2120 2280 2160 2285
rect 6820 2315 6860 2320
rect 6820 2285 6825 2315
rect 6855 2285 6860 2315
rect 6820 2280 6860 2285
rect 6895 2315 6935 2320
rect 6895 2285 6900 2315
rect 6930 2285 6935 2315
rect 6895 2280 6935 2285
rect 2000 2260 2040 2265
rect 2000 2230 2005 2260
rect 2035 2230 2040 2260
rect 2000 2225 2040 2230
rect 2075 2260 2115 2265
rect 2075 2230 2080 2260
rect 2110 2230 2115 2260
rect 2075 2225 2115 2230
rect 2085 2075 2105 2225
rect 2130 1890 2150 2280
rect 6830 1890 6850 2280
rect 6950 2265 6970 6340
rect 7230 6210 7350 6465
rect 7930 9635 8050 9650
rect 7930 9605 7975 9635
rect 8005 9605 8050 9635
rect 7930 9570 8050 9605
rect 7930 9540 7975 9570
rect 8005 9540 8050 9570
rect 7930 9500 8050 9540
rect 7930 9470 7975 9500
rect 8005 9470 8050 9500
rect 7930 9430 8050 9470
rect 7930 9400 7975 9430
rect 8005 9400 8050 9430
rect 7930 9360 8050 9400
rect 7930 9330 7975 9360
rect 8005 9330 8050 9360
rect 7930 9295 8050 9330
rect 7930 9265 7975 9295
rect 8005 9265 8050 9295
rect 7930 9235 8050 9265
rect 7930 9205 7975 9235
rect 8005 9205 8050 9235
rect 7930 9170 8050 9205
rect 7930 9140 7975 9170
rect 8005 9140 8050 9170
rect 7930 9100 8050 9140
rect 7930 9070 7975 9100
rect 8005 9070 8050 9100
rect 7930 9030 8050 9070
rect 7930 9000 7975 9030
rect 8005 9000 8050 9030
rect 7930 8960 8050 9000
rect 7930 8930 7975 8960
rect 8005 8930 8050 8960
rect 7930 8895 8050 8930
rect 7930 8865 7975 8895
rect 8005 8865 8050 8895
rect 7930 8835 8050 8865
rect 7930 8805 7975 8835
rect 8005 8805 8050 8835
rect 7930 8770 8050 8805
rect 7930 8740 7975 8770
rect 8005 8740 8050 8770
rect 7930 8700 8050 8740
rect 7930 8670 7975 8700
rect 8005 8670 8050 8700
rect 7930 8630 8050 8670
rect 7930 8600 7975 8630
rect 8005 8600 8050 8630
rect 7930 8560 8050 8600
rect 7930 8530 7975 8560
rect 8005 8530 8050 8560
rect 7930 8495 8050 8530
rect 7930 8465 7975 8495
rect 8005 8465 8050 8495
rect 7930 8435 8050 8465
rect 7930 8405 7975 8435
rect 8005 8405 8050 8435
rect 7930 8370 8050 8405
rect 7930 8340 7975 8370
rect 8005 8340 8050 8370
rect 7930 8300 8050 8340
rect 7930 8270 7975 8300
rect 8005 8270 8050 8300
rect 7930 8230 8050 8270
rect 7930 8200 7975 8230
rect 8005 8200 8050 8230
rect 7930 8160 8050 8200
rect 7930 8130 7975 8160
rect 8005 8130 8050 8160
rect 7930 8095 8050 8130
rect 7930 8065 7975 8095
rect 8005 8065 8050 8095
rect 7930 8035 8050 8065
rect 7930 8005 7975 8035
rect 8005 8005 8050 8035
rect 7930 7970 8050 8005
rect 7930 7940 7975 7970
rect 8005 7940 8050 7970
rect 7930 7900 8050 7940
rect 7930 7870 7975 7900
rect 8005 7870 8050 7900
rect 7930 7830 8050 7870
rect 7930 7800 7975 7830
rect 8005 7800 8050 7830
rect 7930 7760 8050 7800
rect 7930 7730 7975 7760
rect 8005 7730 8050 7760
rect 7930 7695 8050 7730
rect 7930 7665 7975 7695
rect 8005 7665 8050 7695
rect 7930 7635 8050 7665
rect 7930 7605 7975 7635
rect 8005 7605 8050 7635
rect 7930 7570 8050 7605
rect 7930 7540 7975 7570
rect 8005 7540 8050 7570
rect 7930 7500 8050 7540
rect 7930 7470 7975 7500
rect 8005 7470 8050 7500
rect 7930 7430 8050 7470
rect 7930 7400 7975 7430
rect 8005 7400 8050 7430
rect 7930 7360 8050 7400
rect 7930 7330 7975 7360
rect 8005 7330 8050 7360
rect 7930 7295 8050 7330
rect 7930 7265 7975 7295
rect 8005 7265 8050 7295
rect 7930 7235 8050 7265
rect 7930 7205 7975 7235
rect 8005 7205 8050 7235
rect 7930 7170 8050 7205
rect 7930 7140 7975 7170
rect 8005 7140 8050 7170
rect 7930 7100 8050 7140
rect 7930 7070 7975 7100
rect 8005 7070 8050 7100
rect 7930 7030 8050 7070
rect 7930 7000 7975 7030
rect 8005 7000 8050 7030
rect 7930 6960 8050 7000
rect 7930 6930 7975 6960
rect 8005 6930 8050 6960
rect 7930 6895 8050 6930
rect 7930 6865 7975 6895
rect 8005 6865 8050 6895
rect 7930 6835 8050 6865
rect 7930 6805 7975 6835
rect 8005 6805 8050 6835
rect 7930 6770 8050 6805
rect 7930 6740 7975 6770
rect 8005 6740 8050 6770
rect 7930 6700 8050 6740
rect 7930 6670 7975 6700
rect 8005 6670 8050 6700
rect 7930 6630 8050 6670
rect 7930 6600 7975 6630
rect 8005 6600 8050 6630
rect 7930 6560 8050 6600
rect 7930 6530 7975 6560
rect 8005 6530 8050 6560
rect 7930 6495 8050 6530
rect 7930 6465 7975 6495
rect 8005 6465 8050 6495
rect 7580 6205 7700 6210
rect 7580 6175 7585 6205
rect 7615 6175 7625 6205
rect 7655 6175 7665 6205
rect 7695 6175 7700 6205
rect 7930 6195 8050 6465
rect 8280 9635 8400 9650
rect 8280 9605 8325 9635
rect 8355 9605 8400 9635
rect 8280 9570 8400 9605
rect 8280 9540 8325 9570
rect 8355 9540 8400 9570
rect 8280 9500 8400 9540
rect 8280 9470 8325 9500
rect 8355 9470 8400 9500
rect 8280 9430 8400 9470
rect 8280 9400 8325 9430
rect 8355 9400 8400 9430
rect 8280 9360 8400 9400
rect 8280 9330 8325 9360
rect 8355 9330 8400 9360
rect 8280 9295 8400 9330
rect 8280 9265 8325 9295
rect 8355 9265 8400 9295
rect 8280 9235 8400 9265
rect 8280 9205 8325 9235
rect 8355 9205 8400 9235
rect 8280 9170 8400 9205
rect 8280 9140 8325 9170
rect 8355 9140 8400 9170
rect 8280 9100 8400 9140
rect 8280 9070 8325 9100
rect 8355 9070 8400 9100
rect 8280 9030 8400 9070
rect 8280 9000 8325 9030
rect 8355 9000 8400 9030
rect 8280 8960 8400 9000
rect 8280 8930 8325 8960
rect 8355 8930 8400 8960
rect 8280 8895 8400 8930
rect 8280 8865 8325 8895
rect 8355 8865 8400 8895
rect 8280 8835 8400 8865
rect 8280 8805 8325 8835
rect 8355 8805 8400 8835
rect 8280 8770 8400 8805
rect 8280 8740 8325 8770
rect 8355 8740 8400 8770
rect 8280 8700 8400 8740
rect 8280 8670 8325 8700
rect 8355 8670 8400 8700
rect 8280 8630 8400 8670
rect 8280 8600 8325 8630
rect 8355 8600 8400 8630
rect 8280 8560 8400 8600
rect 8280 8530 8325 8560
rect 8355 8530 8400 8560
rect 8280 8495 8400 8530
rect 8280 8465 8325 8495
rect 8355 8465 8400 8495
rect 8280 8435 8400 8465
rect 8280 8405 8325 8435
rect 8355 8405 8400 8435
rect 8280 8370 8400 8405
rect 8280 8340 8325 8370
rect 8355 8340 8400 8370
rect 8280 8300 8400 8340
rect 8280 8270 8325 8300
rect 8355 8270 8400 8300
rect 8280 8230 8400 8270
rect 8280 8200 8325 8230
rect 8355 8200 8400 8230
rect 8280 8160 8400 8200
rect 8280 8130 8325 8160
rect 8355 8130 8400 8160
rect 8280 8095 8400 8130
rect 8280 8065 8325 8095
rect 8355 8065 8400 8095
rect 8280 8035 8400 8065
rect 8280 8005 8325 8035
rect 8355 8005 8400 8035
rect 8280 7970 8400 8005
rect 8280 7940 8325 7970
rect 8355 7940 8400 7970
rect 8280 7900 8400 7940
rect 8280 7870 8325 7900
rect 8355 7870 8400 7900
rect 8280 7830 8400 7870
rect 8280 7800 8325 7830
rect 8355 7800 8400 7830
rect 8280 7760 8400 7800
rect 8280 7730 8325 7760
rect 8355 7730 8400 7760
rect 8280 7695 8400 7730
rect 8280 7665 8325 7695
rect 8355 7665 8400 7695
rect 8280 7635 8400 7665
rect 8280 7605 8325 7635
rect 8355 7605 8400 7635
rect 8280 7570 8400 7605
rect 8280 7540 8325 7570
rect 8355 7540 8400 7570
rect 8280 7500 8400 7540
rect 8280 7470 8325 7500
rect 8355 7470 8400 7500
rect 8280 7430 8400 7470
rect 8280 7400 8325 7430
rect 8355 7400 8400 7430
rect 8280 7360 8400 7400
rect 8280 7330 8325 7360
rect 8355 7330 8400 7360
rect 8280 7295 8400 7330
rect 8280 7265 8325 7295
rect 8355 7265 8400 7295
rect 8280 7235 8400 7265
rect 8280 7205 8325 7235
rect 8355 7205 8400 7235
rect 8280 7170 8400 7205
rect 8280 7140 8325 7170
rect 8355 7140 8400 7170
rect 8280 7100 8400 7140
rect 8280 7070 8325 7100
rect 8355 7070 8400 7100
rect 8280 7030 8400 7070
rect 8280 7000 8325 7030
rect 8355 7000 8400 7030
rect 8280 6960 8400 7000
rect 8280 6930 8325 6960
rect 8355 6930 8400 6960
rect 8280 6895 8400 6930
rect 8280 6865 8325 6895
rect 8355 6865 8400 6895
rect 8280 6835 8400 6865
rect 8280 6805 8325 6835
rect 8355 6805 8400 6835
rect 8280 6770 8400 6805
rect 8280 6740 8325 6770
rect 8355 6740 8400 6770
rect 8280 6700 8400 6740
rect 8280 6670 8325 6700
rect 8355 6670 8400 6700
rect 8280 6630 8400 6670
rect 8280 6600 8325 6630
rect 8355 6600 8400 6630
rect 8280 6560 8400 6600
rect 8280 6530 8325 6560
rect 8355 6530 8400 6560
rect 8280 6495 8400 6530
rect 8280 6465 8325 6495
rect 8355 6465 8400 6495
rect 8280 6210 8400 6465
rect 8630 9635 8750 9650
rect 8630 9605 8675 9635
rect 8705 9605 8750 9635
rect 8630 9570 8750 9605
rect 8630 9540 8675 9570
rect 8705 9540 8750 9570
rect 8630 9500 8750 9540
rect 8630 9470 8675 9500
rect 8705 9470 8750 9500
rect 8630 9430 8750 9470
rect 8630 9400 8675 9430
rect 8705 9400 8750 9430
rect 8630 9360 8750 9400
rect 8630 9330 8675 9360
rect 8705 9330 8750 9360
rect 8630 9295 8750 9330
rect 8630 9265 8675 9295
rect 8705 9265 8750 9295
rect 8630 9235 8750 9265
rect 8630 9205 8675 9235
rect 8705 9205 8750 9235
rect 8630 9170 8750 9205
rect 8630 9140 8675 9170
rect 8705 9140 8750 9170
rect 8630 9100 8750 9140
rect 8630 9070 8675 9100
rect 8705 9070 8750 9100
rect 8630 9030 8750 9070
rect 8630 9000 8675 9030
rect 8705 9000 8750 9030
rect 8630 8960 8750 9000
rect 8630 8930 8675 8960
rect 8705 8930 8750 8960
rect 8630 8895 8750 8930
rect 8630 8865 8675 8895
rect 8705 8865 8750 8895
rect 8630 8835 8750 8865
rect 8630 8805 8675 8835
rect 8705 8805 8750 8835
rect 8630 8770 8750 8805
rect 8630 8740 8675 8770
rect 8705 8740 8750 8770
rect 8630 8700 8750 8740
rect 8630 8670 8675 8700
rect 8705 8670 8750 8700
rect 8630 8630 8750 8670
rect 8630 8600 8675 8630
rect 8705 8600 8750 8630
rect 8630 8560 8750 8600
rect 8630 8530 8675 8560
rect 8705 8530 8750 8560
rect 8630 8495 8750 8530
rect 8630 8465 8675 8495
rect 8705 8465 8750 8495
rect 8630 8435 8750 8465
rect 8630 8405 8675 8435
rect 8705 8405 8750 8435
rect 8630 8370 8750 8405
rect 8630 8340 8675 8370
rect 8705 8340 8750 8370
rect 8630 8300 8750 8340
rect 8630 8270 8675 8300
rect 8705 8270 8750 8300
rect 8630 8230 8750 8270
rect 8630 8200 8675 8230
rect 8705 8200 8750 8230
rect 8630 8160 8750 8200
rect 8630 8130 8675 8160
rect 8705 8130 8750 8160
rect 8630 8095 8750 8130
rect 8630 8065 8675 8095
rect 8705 8065 8750 8095
rect 8630 8035 8750 8065
rect 8630 8005 8675 8035
rect 8705 8005 8750 8035
rect 8630 7970 8750 8005
rect 8630 7940 8675 7970
rect 8705 7940 8750 7970
rect 8630 7900 8750 7940
rect 8630 7870 8675 7900
rect 8705 7870 8750 7900
rect 8630 7830 8750 7870
rect 8630 7800 8675 7830
rect 8705 7800 8750 7830
rect 8630 7760 8750 7800
rect 8630 7730 8675 7760
rect 8705 7730 8750 7760
rect 8630 7695 8750 7730
rect 8630 7665 8675 7695
rect 8705 7665 8750 7695
rect 8630 7635 8750 7665
rect 8630 7605 8675 7635
rect 8705 7605 8750 7635
rect 8630 7570 8750 7605
rect 8630 7540 8675 7570
rect 8705 7540 8750 7570
rect 8630 7500 8750 7540
rect 8630 7470 8675 7500
rect 8705 7470 8750 7500
rect 8630 7430 8750 7470
rect 8630 7400 8675 7430
rect 8705 7400 8750 7430
rect 8630 7360 8750 7400
rect 8630 7330 8675 7360
rect 8705 7330 8750 7360
rect 8630 7295 8750 7330
rect 8630 7265 8675 7295
rect 8705 7265 8750 7295
rect 8630 7235 8750 7265
rect 8630 7205 8675 7235
rect 8705 7205 8750 7235
rect 8630 7170 8750 7205
rect 8630 7140 8675 7170
rect 8705 7140 8750 7170
rect 8630 7100 8750 7140
rect 8630 7070 8675 7100
rect 8705 7070 8750 7100
rect 8630 7030 8750 7070
rect 8630 7000 8675 7030
rect 8705 7000 8750 7030
rect 8630 6960 8750 7000
rect 8630 6930 8675 6960
rect 8705 6930 8750 6960
rect 8630 6895 8750 6930
rect 8630 6865 8675 6895
rect 8705 6865 8750 6895
rect 8630 6835 8750 6865
rect 8630 6805 8675 6835
rect 8705 6805 8750 6835
rect 8630 6770 8750 6805
rect 8630 6740 8675 6770
rect 8705 6740 8750 6770
rect 8630 6700 8750 6740
rect 8630 6670 8675 6700
rect 8705 6670 8750 6700
rect 8630 6630 8750 6670
rect 8630 6600 8675 6630
rect 8705 6600 8750 6630
rect 8630 6560 8750 6600
rect 8630 6530 8675 6560
rect 8705 6530 8750 6560
rect 8630 6495 8750 6530
rect 8630 6465 8675 6495
rect 8705 6465 8750 6495
rect 8630 6210 8750 6465
rect 8980 9635 9100 9650
rect 8980 9605 9025 9635
rect 9055 9605 9100 9635
rect 8980 9570 9100 9605
rect 8980 9540 9025 9570
rect 9055 9540 9100 9570
rect 8980 9500 9100 9540
rect 8980 9470 9025 9500
rect 9055 9470 9100 9500
rect 8980 9430 9100 9470
rect 8980 9400 9025 9430
rect 9055 9400 9100 9430
rect 8980 9360 9100 9400
rect 8980 9330 9025 9360
rect 9055 9330 9100 9360
rect 8980 9295 9100 9330
rect 8980 9265 9025 9295
rect 9055 9265 9100 9295
rect 8980 9235 9100 9265
rect 8980 9205 9025 9235
rect 9055 9205 9100 9235
rect 8980 9170 9100 9205
rect 8980 9140 9025 9170
rect 9055 9140 9100 9170
rect 8980 9100 9100 9140
rect 8980 9070 9025 9100
rect 9055 9070 9100 9100
rect 8980 9030 9100 9070
rect 8980 9000 9025 9030
rect 9055 9000 9100 9030
rect 8980 8960 9100 9000
rect 8980 8930 9025 8960
rect 9055 8930 9100 8960
rect 8980 8895 9100 8930
rect 8980 8865 9025 8895
rect 9055 8865 9100 8895
rect 8980 8835 9100 8865
rect 8980 8805 9025 8835
rect 9055 8805 9100 8835
rect 8980 8770 9100 8805
rect 8980 8740 9025 8770
rect 9055 8740 9100 8770
rect 8980 8700 9100 8740
rect 8980 8670 9025 8700
rect 9055 8670 9100 8700
rect 8980 8630 9100 8670
rect 8980 8600 9025 8630
rect 9055 8600 9100 8630
rect 8980 8560 9100 8600
rect 8980 8530 9025 8560
rect 9055 8530 9100 8560
rect 8980 8495 9100 8530
rect 8980 8465 9025 8495
rect 9055 8465 9100 8495
rect 8980 8435 9100 8465
rect 8980 8405 9025 8435
rect 9055 8405 9100 8435
rect 8980 8370 9100 8405
rect 8980 8340 9025 8370
rect 9055 8340 9100 8370
rect 8980 8300 9100 8340
rect 8980 8270 9025 8300
rect 9055 8270 9100 8300
rect 8980 8230 9100 8270
rect 8980 8200 9025 8230
rect 9055 8200 9100 8230
rect 8980 8160 9100 8200
rect 8980 8130 9025 8160
rect 9055 8130 9100 8160
rect 8980 8095 9100 8130
rect 8980 8065 9025 8095
rect 9055 8065 9100 8095
rect 8980 8035 9100 8065
rect 8980 8005 9025 8035
rect 9055 8005 9100 8035
rect 8980 7970 9100 8005
rect 8980 7940 9025 7970
rect 9055 7940 9100 7970
rect 8980 7900 9100 7940
rect 8980 7870 9025 7900
rect 9055 7870 9100 7900
rect 8980 7830 9100 7870
rect 8980 7800 9025 7830
rect 9055 7800 9100 7830
rect 8980 7760 9100 7800
rect 8980 7730 9025 7760
rect 9055 7730 9100 7760
rect 8980 7695 9100 7730
rect 8980 7665 9025 7695
rect 9055 7665 9100 7695
rect 8980 7635 9100 7665
rect 8980 7605 9025 7635
rect 9055 7605 9100 7635
rect 8980 7570 9100 7605
rect 8980 7540 9025 7570
rect 9055 7540 9100 7570
rect 8980 7500 9100 7540
rect 8980 7470 9025 7500
rect 9055 7470 9100 7500
rect 8980 7430 9100 7470
rect 8980 7400 9025 7430
rect 9055 7400 9100 7430
rect 8980 7360 9100 7400
rect 8980 7330 9025 7360
rect 9055 7330 9100 7360
rect 8980 7295 9100 7330
rect 8980 7265 9025 7295
rect 9055 7265 9100 7295
rect 8980 7235 9100 7265
rect 8980 7205 9025 7235
rect 9055 7205 9100 7235
rect 8980 7170 9100 7205
rect 8980 7140 9025 7170
rect 9055 7140 9100 7170
rect 8980 7100 9100 7140
rect 8980 7070 9025 7100
rect 9055 7070 9100 7100
rect 8980 7030 9100 7070
rect 8980 7000 9025 7030
rect 9055 7000 9100 7030
rect 8980 6960 9100 7000
rect 8980 6930 9025 6960
rect 9055 6930 9100 6960
rect 8980 6895 9100 6930
rect 8980 6865 9025 6895
rect 9055 6865 9100 6895
rect 8980 6835 9100 6865
rect 8980 6805 9025 6835
rect 9055 6805 9100 6835
rect 8980 6770 9100 6805
rect 8980 6740 9025 6770
rect 9055 6740 9100 6770
rect 8980 6700 9100 6740
rect 8980 6670 9025 6700
rect 9055 6670 9100 6700
rect 8980 6630 9100 6670
rect 8980 6600 9025 6630
rect 9055 6600 9100 6630
rect 8980 6560 9100 6600
rect 8980 6530 9025 6560
rect 9055 6530 9100 6560
rect 8980 6495 9100 6530
rect 8980 6465 9025 6495
rect 9055 6465 9100 6495
rect 8980 6210 9100 6465
rect 7580 6165 7700 6175
rect 7580 6135 7585 6165
rect 7615 6135 7625 6165
rect 7655 6135 7665 6165
rect 7695 6135 7700 6165
rect 7580 6125 7700 6135
rect 7580 6095 7585 6125
rect 7615 6095 7625 6125
rect 7655 6095 7665 6125
rect 7695 6095 7700 6125
rect 6865 2260 6905 2265
rect 6865 2230 6870 2260
rect 6900 2230 6905 2260
rect 6865 2225 6905 2230
rect 6940 2260 6980 2265
rect 6940 2230 6945 2260
rect 6975 2230 6980 2260
rect 6940 2225 6980 2230
rect 6875 2075 6895 2225
rect 1280 1130 1285 1160
rect 1315 1130 1325 1160
rect 1355 1130 1365 1160
rect 1395 1130 1400 1160
rect 1280 1120 1400 1130
rect 1280 1090 1285 1120
rect 1315 1090 1325 1120
rect 1355 1090 1365 1120
rect 1395 1090 1400 1120
rect 1280 1080 1400 1090
rect 1280 1050 1285 1080
rect 1315 1050 1325 1080
rect 1355 1050 1365 1080
rect 1395 1050 1400 1080
rect 1280 1045 1400 1050
rect 4415 1160 4455 1165
rect 4415 1130 4420 1160
rect 4450 1130 4455 1160
rect 4415 1120 4455 1130
rect 4415 1090 4420 1120
rect 4450 1090 4455 1120
rect 4415 1080 4455 1090
rect 4415 1050 4420 1080
rect 4450 1050 4455 1080
rect 4415 1045 4455 1050
rect 4525 1160 4565 1165
rect 4525 1130 4530 1160
rect 4560 1130 4565 1160
rect 4525 1120 4565 1130
rect 4525 1090 4530 1120
rect 4560 1090 4565 1120
rect 4525 1080 4565 1090
rect 4525 1050 4530 1080
rect 4560 1050 4565 1080
rect 4525 1045 4565 1050
rect 7580 1160 7700 6095
rect 7580 1130 7585 1160
rect 7615 1130 7625 1160
rect 7655 1130 7665 1160
rect 7695 1130 7700 1160
rect 7580 1120 7700 1130
rect 7580 1090 7585 1120
rect 7615 1090 7625 1120
rect 7655 1090 7665 1120
rect 7695 1090 7700 1120
rect 7580 1080 7700 1090
rect 7580 1050 7585 1080
rect 7615 1050 7625 1080
rect 7655 1050 7665 1080
rect 7695 1050 7700 1080
rect 7580 1045 7700 1050
rect -120 -1305 0 -1240
rect -120 -1335 -75 -1305
rect -45 -1335 0 -1305
rect -120 -1370 0 -1335
rect -120 -1400 -75 -1370
rect -45 -1400 0 -1370
rect -120 -1440 0 -1400
rect -120 -1470 -75 -1440
rect -45 -1470 0 -1440
rect -120 -1510 0 -1470
rect -120 -1540 -75 -1510
rect -45 -1540 0 -1510
rect -120 -1580 0 -1540
rect -120 -1610 -75 -1580
rect -45 -1610 0 -1580
rect -120 -1645 0 -1610
rect -120 -1675 -75 -1645
rect -45 -1675 0 -1645
rect -120 -1705 0 -1675
rect -120 -1735 -75 -1705
rect -45 -1735 0 -1705
rect -120 -1770 0 -1735
rect -120 -1800 -75 -1770
rect -45 -1800 0 -1770
rect -120 -1840 0 -1800
rect -120 -1870 -75 -1840
rect -45 -1870 0 -1840
rect -120 -1910 0 -1870
rect -120 -1940 -75 -1910
rect -45 -1940 0 -1910
rect -120 -1980 0 -1940
rect -120 -2010 -75 -1980
rect -45 -2010 0 -1980
rect -120 -2045 0 -2010
rect -120 -2075 -75 -2045
rect -45 -2075 0 -2045
rect -120 -2105 0 -2075
rect -120 -2135 -75 -2105
rect -45 -2135 0 -2105
rect -120 -2170 0 -2135
rect -120 -2200 -75 -2170
rect -45 -2200 0 -2170
rect -120 -2240 0 -2200
rect -120 -2270 -75 -2240
rect -45 -2270 0 -2240
rect -120 -2310 0 -2270
rect -120 -2340 -75 -2310
rect -45 -2340 0 -2310
rect -120 -2380 0 -2340
rect -120 -2410 -75 -2380
rect -45 -2410 0 -2380
rect -120 -2445 0 -2410
rect -120 -2475 -75 -2445
rect -45 -2475 0 -2445
rect -120 -2505 0 -2475
rect -120 -2535 -75 -2505
rect -45 -2535 0 -2505
rect -120 -2570 0 -2535
rect -120 -2600 -75 -2570
rect -45 -2600 0 -2570
rect -120 -2640 0 -2600
rect -120 -2670 -75 -2640
rect -45 -2670 0 -2640
rect -120 -2710 0 -2670
rect -120 -2740 -75 -2710
rect -45 -2740 0 -2710
rect -120 -2780 0 -2740
rect -120 -2810 -75 -2780
rect -45 -2810 0 -2780
rect -120 -2845 0 -2810
rect -120 -2875 -75 -2845
rect -45 -2875 0 -2845
rect -120 -2890 0 -2875
rect 230 -1305 350 -1240
rect 230 -1335 275 -1305
rect 305 -1335 350 -1305
rect 230 -1370 350 -1335
rect 230 -1400 275 -1370
rect 305 -1400 350 -1370
rect 230 -1440 350 -1400
rect 230 -1470 275 -1440
rect 305 -1470 350 -1440
rect 230 -1510 350 -1470
rect 230 -1540 275 -1510
rect 305 -1540 350 -1510
rect 230 -1580 350 -1540
rect 230 -1610 275 -1580
rect 305 -1610 350 -1580
rect 230 -1645 350 -1610
rect 230 -1675 275 -1645
rect 305 -1675 350 -1645
rect 230 -1705 350 -1675
rect 230 -1735 275 -1705
rect 305 -1735 350 -1705
rect 230 -1770 350 -1735
rect 230 -1800 275 -1770
rect 305 -1800 350 -1770
rect 230 -1840 350 -1800
rect 230 -1870 275 -1840
rect 305 -1870 350 -1840
rect 230 -1910 350 -1870
rect 230 -1940 275 -1910
rect 305 -1940 350 -1910
rect 230 -1980 350 -1940
rect 230 -2010 275 -1980
rect 305 -2010 350 -1980
rect 230 -2045 350 -2010
rect 230 -2075 275 -2045
rect 305 -2075 350 -2045
rect 230 -2105 350 -2075
rect 230 -2135 275 -2105
rect 305 -2135 350 -2105
rect 230 -2170 350 -2135
rect 230 -2200 275 -2170
rect 305 -2200 350 -2170
rect 230 -2240 350 -2200
rect 230 -2270 275 -2240
rect 305 -2270 350 -2240
rect 230 -2310 350 -2270
rect 230 -2340 275 -2310
rect 305 -2340 350 -2310
rect 230 -2380 350 -2340
rect 230 -2410 275 -2380
rect 305 -2410 350 -2380
rect 230 -2445 350 -2410
rect 230 -2475 275 -2445
rect 305 -2475 350 -2445
rect 230 -2505 350 -2475
rect 230 -2535 275 -2505
rect 305 -2535 350 -2505
rect 230 -2570 350 -2535
rect 230 -2600 275 -2570
rect 305 -2600 350 -2570
rect 230 -2640 350 -2600
rect 230 -2670 275 -2640
rect 305 -2670 350 -2640
rect 230 -2710 350 -2670
rect 230 -2740 275 -2710
rect 305 -2740 350 -2710
rect 230 -2780 350 -2740
rect 230 -2810 275 -2780
rect 305 -2810 350 -2780
rect 230 -2845 350 -2810
rect 230 -2875 275 -2845
rect 305 -2875 350 -2845
rect 230 -2890 350 -2875
rect 580 -1305 700 -1240
rect 580 -1335 625 -1305
rect 655 -1335 700 -1305
rect 580 -1370 700 -1335
rect 580 -1400 625 -1370
rect 655 -1400 700 -1370
rect 580 -1440 700 -1400
rect 580 -1470 625 -1440
rect 655 -1470 700 -1440
rect 580 -1510 700 -1470
rect 580 -1540 625 -1510
rect 655 -1540 700 -1510
rect 580 -1580 700 -1540
rect 580 -1610 625 -1580
rect 655 -1610 700 -1580
rect 580 -1645 700 -1610
rect 580 -1675 625 -1645
rect 655 -1675 700 -1645
rect 580 -1705 700 -1675
rect 580 -1735 625 -1705
rect 655 -1735 700 -1705
rect 580 -1770 700 -1735
rect 580 -1800 625 -1770
rect 655 -1800 700 -1770
rect 580 -1840 700 -1800
rect 580 -1870 625 -1840
rect 655 -1870 700 -1840
rect 580 -1910 700 -1870
rect 580 -1940 625 -1910
rect 655 -1940 700 -1910
rect 580 -1980 700 -1940
rect 580 -2010 625 -1980
rect 655 -2010 700 -1980
rect 580 -2045 700 -2010
rect 580 -2075 625 -2045
rect 655 -2075 700 -2045
rect 580 -2105 700 -2075
rect 580 -2135 625 -2105
rect 655 -2135 700 -2105
rect 580 -2170 700 -2135
rect 580 -2200 625 -2170
rect 655 -2200 700 -2170
rect 580 -2240 700 -2200
rect 580 -2270 625 -2240
rect 655 -2270 700 -2240
rect 580 -2310 700 -2270
rect 580 -2340 625 -2310
rect 655 -2340 700 -2310
rect 580 -2380 700 -2340
rect 580 -2410 625 -2380
rect 655 -2410 700 -2380
rect 580 -2445 700 -2410
rect 580 -2475 625 -2445
rect 655 -2475 700 -2445
rect 580 -2505 700 -2475
rect 580 -2535 625 -2505
rect 655 -2535 700 -2505
rect 580 -2570 700 -2535
rect 580 -2600 625 -2570
rect 655 -2600 700 -2570
rect 580 -2640 700 -2600
rect 580 -2670 625 -2640
rect 655 -2670 700 -2640
rect 580 -2710 700 -2670
rect 580 -2740 625 -2710
rect 655 -2740 700 -2710
rect 580 -2780 700 -2740
rect 580 -2810 625 -2780
rect 655 -2810 700 -2780
rect 580 -2845 700 -2810
rect 580 -2875 625 -2845
rect 655 -2875 700 -2845
rect 580 -2890 700 -2875
rect 930 -1305 1050 -1240
rect 930 -1335 975 -1305
rect 1005 -1335 1050 -1305
rect 930 -1370 1050 -1335
rect 930 -1400 975 -1370
rect 1005 -1400 1050 -1370
rect 930 -1440 1050 -1400
rect 930 -1470 975 -1440
rect 1005 -1470 1050 -1440
rect 930 -1510 1050 -1470
rect 930 -1540 975 -1510
rect 1005 -1540 1050 -1510
rect 930 -1580 1050 -1540
rect 930 -1610 975 -1580
rect 1005 -1610 1050 -1580
rect 930 -1645 1050 -1610
rect 930 -1675 975 -1645
rect 1005 -1675 1050 -1645
rect 930 -1705 1050 -1675
rect 930 -1735 975 -1705
rect 1005 -1735 1050 -1705
rect 930 -1770 1050 -1735
rect 930 -1800 975 -1770
rect 1005 -1800 1050 -1770
rect 930 -1840 1050 -1800
rect 930 -1870 975 -1840
rect 1005 -1870 1050 -1840
rect 930 -1910 1050 -1870
rect 930 -1940 975 -1910
rect 1005 -1940 1050 -1910
rect 930 -1980 1050 -1940
rect 930 -2010 975 -1980
rect 1005 -2010 1050 -1980
rect 930 -2045 1050 -2010
rect 930 -2075 975 -2045
rect 1005 -2075 1050 -2045
rect 930 -2105 1050 -2075
rect 930 -2135 975 -2105
rect 1005 -2135 1050 -2105
rect 930 -2170 1050 -2135
rect 930 -2200 975 -2170
rect 1005 -2200 1050 -2170
rect 930 -2240 1050 -2200
rect 930 -2270 975 -2240
rect 1005 -2270 1050 -2240
rect 930 -2310 1050 -2270
rect 930 -2340 975 -2310
rect 1005 -2340 1050 -2310
rect 930 -2380 1050 -2340
rect 930 -2410 975 -2380
rect 1005 -2410 1050 -2380
rect 930 -2445 1050 -2410
rect 930 -2475 975 -2445
rect 1005 -2475 1050 -2445
rect 930 -2505 1050 -2475
rect 930 -2535 975 -2505
rect 1005 -2535 1050 -2505
rect 930 -2570 1050 -2535
rect 930 -2600 975 -2570
rect 1005 -2600 1050 -2570
rect 930 -2640 1050 -2600
rect 930 -2670 975 -2640
rect 1005 -2670 1050 -2640
rect 930 -2710 1050 -2670
rect 930 -2740 975 -2710
rect 1005 -2740 1050 -2710
rect 930 -2780 1050 -2740
rect 930 -2810 975 -2780
rect 1005 -2810 1050 -2780
rect 930 -2845 1050 -2810
rect 930 -2875 975 -2845
rect 1005 -2875 1050 -2845
rect 930 -2890 1050 -2875
rect 1280 -1305 1400 -1240
rect 1280 -1335 1325 -1305
rect 1355 -1335 1400 -1305
rect 1280 -1370 1400 -1335
rect 1280 -1400 1325 -1370
rect 1355 -1400 1400 -1370
rect 1280 -1440 1400 -1400
rect 1280 -1470 1325 -1440
rect 1355 -1470 1400 -1440
rect 1280 -1510 1400 -1470
rect 1280 -1540 1325 -1510
rect 1355 -1540 1400 -1510
rect 1280 -1580 1400 -1540
rect 1280 -1610 1325 -1580
rect 1355 -1610 1400 -1580
rect 1280 -1645 1400 -1610
rect 1280 -1675 1325 -1645
rect 1355 -1675 1400 -1645
rect 1280 -1705 1400 -1675
rect 1280 -1735 1325 -1705
rect 1355 -1735 1400 -1705
rect 1280 -1770 1400 -1735
rect 1280 -1800 1325 -1770
rect 1355 -1800 1400 -1770
rect 1280 -1840 1400 -1800
rect 1280 -1870 1325 -1840
rect 1355 -1870 1400 -1840
rect 1280 -1910 1400 -1870
rect 1280 -1940 1325 -1910
rect 1355 -1940 1400 -1910
rect 1280 -1980 1400 -1940
rect 1280 -2010 1325 -1980
rect 1355 -2010 1400 -1980
rect 1280 -2045 1400 -2010
rect 1280 -2075 1325 -2045
rect 1355 -2075 1400 -2045
rect 1280 -2105 1400 -2075
rect 1280 -2135 1325 -2105
rect 1355 -2135 1400 -2105
rect 1280 -2170 1400 -2135
rect 1280 -2200 1325 -2170
rect 1355 -2200 1400 -2170
rect 1280 -2240 1400 -2200
rect 1280 -2270 1325 -2240
rect 1355 -2270 1400 -2240
rect 1280 -2310 1400 -2270
rect 1280 -2340 1325 -2310
rect 1355 -2340 1400 -2310
rect 1280 -2380 1400 -2340
rect 1280 -2410 1325 -2380
rect 1355 -2410 1400 -2380
rect 1280 -2445 1400 -2410
rect 1280 -2475 1325 -2445
rect 1355 -2475 1400 -2445
rect 1280 -2505 1400 -2475
rect 1280 -2535 1325 -2505
rect 1355 -2535 1400 -2505
rect 1280 -2570 1400 -2535
rect 1280 -2600 1325 -2570
rect 1355 -2600 1400 -2570
rect 1280 -2640 1400 -2600
rect 1280 -2670 1325 -2640
rect 1355 -2670 1400 -2640
rect 1280 -2710 1400 -2670
rect 1280 -2740 1325 -2710
rect 1355 -2740 1400 -2710
rect 1280 -2780 1400 -2740
rect 1280 -2810 1325 -2780
rect 1355 -2810 1400 -2780
rect 1280 -2845 1400 -2810
rect 1280 -2875 1325 -2845
rect 1355 -2875 1400 -2845
rect 1280 -2890 1400 -2875
rect 1630 -1305 1750 -1240
rect 1630 -1335 1675 -1305
rect 1705 -1335 1750 -1305
rect 1630 -1370 1750 -1335
rect 1630 -1400 1675 -1370
rect 1705 -1400 1750 -1370
rect 1630 -1440 1750 -1400
rect 1630 -1470 1675 -1440
rect 1705 -1470 1750 -1440
rect 1630 -1510 1750 -1470
rect 1630 -1540 1675 -1510
rect 1705 -1540 1750 -1510
rect 1630 -1580 1750 -1540
rect 1630 -1610 1675 -1580
rect 1705 -1610 1750 -1580
rect 1630 -1645 1750 -1610
rect 1630 -1675 1675 -1645
rect 1705 -1675 1750 -1645
rect 1630 -1705 1750 -1675
rect 1630 -1735 1675 -1705
rect 1705 -1735 1750 -1705
rect 1630 -1770 1750 -1735
rect 1630 -1800 1675 -1770
rect 1705 -1800 1750 -1770
rect 1630 -1840 1750 -1800
rect 1630 -1870 1675 -1840
rect 1705 -1870 1750 -1840
rect 1630 -1910 1750 -1870
rect 1630 -1940 1675 -1910
rect 1705 -1940 1750 -1910
rect 1630 -1980 1750 -1940
rect 1630 -2010 1675 -1980
rect 1705 -2010 1750 -1980
rect 1630 -2045 1750 -2010
rect 1630 -2075 1675 -2045
rect 1705 -2075 1750 -2045
rect 1630 -2105 1750 -2075
rect 1630 -2135 1675 -2105
rect 1705 -2135 1750 -2105
rect 1630 -2170 1750 -2135
rect 1630 -2200 1675 -2170
rect 1705 -2200 1750 -2170
rect 1630 -2240 1750 -2200
rect 1630 -2270 1675 -2240
rect 1705 -2270 1750 -2240
rect 1630 -2310 1750 -2270
rect 1630 -2340 1675 -2310
rect 1705 -2340 1750 -2310
rect 1630 -2380 1750 -2340
rect 1630 -2410 1675 -2380
rect 1705 -2410 1750 -2380
rect 1630 -2445 1750 -2410
rect 1630 -2475 1675 -2445
rect 1705 -2475 1750 -2445
rect 1630 -2505 1750 -2475
rect 1630 -2535 1675 -2505
rect 1705 -2535 1750 -2505
rect 1630 -2570 1750 -2535
rect 1630 -2600 1675 -2570
rect 1705 -2600 1750 -2570
rect 1630 -2640 1750 -2600
rect 1630 -2670 1675 -2640
rect 1705 -2670 1750 -2640
rect 1630 -2710 1750 -2670
rect 1630 -2740 1675 -2710
rect 1705 -2740 1750 -2710
rect 1630 -2780 1750 -2740
rect 1630 -2810 1675 -2780
rect 1705 -2810 1750 -2780
rect 1630 -2845 1750 -2810
rect 1630 -2875 1675 -2845
rect 1705 -2875 1750 -2845
rect 1630 -2890 1750 -2875
rect 1980 -1305 2100 -1240
rect 1980 -1335 2025 -1305
rect 2055 -1335 2100 -1305
rect 1980 -1370 2100 -1335
rect 1980 -1400 2025 -1370
rect 2055 -1400 2100 -1370
rect 1980 -1440 2100 -1400
rect 1980 -1470 2025 -1440
rect 2055 -1470 2100 -1440
rect 1980 -1510 2100 -1470
rect 1980 -1540 2025 -1510
rect 2055 -1540 2100 -1510
rect 1980 -1580 2100 -1540
rect 1980 -1610 2025 -1580
rect 2055 -1610 2100 -1580
rect 1980 -1645 2100 -1610
rect 1980 -1675 2025 -1645
rect 2055 -1675 2100 -1645
rect 1980 -1705 2100 -1675
rect 1980 -1735 2025 -1705
rect 2055 -1735 2100 -1705
rect 1980 -1770 2100 -1735
rect 1980 -1800 2025 -1770
rect 2055 -1800 2100 -1770
rect 1980 -1840 2100 -1800
rect 1980 -1870 2025 -1840
rect 2055 -1870 2100 -1840
rect 1980 -1910 2100 -1870
rect 1980 -1940 2025 -1910
rect 2055 -1940 2100 -1910
rect 1980 -1980 2100 -1940
rect 1980 -2010 2025 -1980
rect 2055 -2010 2100 -1980
rect 1980 -2045 2100 -2010
rect 1980 -2075 2025 -2045
rect 2055 -2075 2100 -2045
rect 1980 -2105 2100 -2075
rect 1980 -2135 2025 -2105
rect 2055 -2135 2100 -2105
rect 1980 -2170 2100 -2135
rect 1980 -2200 2025 -2170
rect 2055 -2200 2100 -2170
rect 1980 -2240 2100 -2200
rect 1980 -2270 2025 -2240
rect 2055 -2270 2100 -2240
rect 1980 -2310 2100 -2270
rect 1980 -2340 2025 -2310
rect 2055 -2340 2100 -2310
rect 1980 -2380 2100 -2340
rect 1980 -2410 2025 -2380
rect 2055 -2410 2100 -2380
rect 1980 -2445 2100 -2410
rect 1980 -2475 2025 -2445
rect 2055 -2475 2100 -2445
rect 1980 -2505 2100 -2475
rect 1980 -2535 2025 -2505
rect 2055 -2535 2100 -2505
rect 1980 -2570 2100 -2535
rect 1980 -2600 2025 -2570
rect 2055 -2600 2100 -2570
rect 1980 -2640 2100 -2600
rect 1980 -2670 2025 -2640
rect 2055 -2670 2100 -2640
rect 1980 -2710 2100 -2670
rect 1980 -2740 2025 -2710
rect 2055 -2740 2100 -2710
rect 1980 -2780 2100 -2740
rect 1980 -2810 2025 -2780
rect 2055 -2810 2100 -2780
rect 1980 -2845 2100 -2810
rect 1980 -2875 2025 -2845
rect 2055 -2875 2100 -2845
rect 1980 -2890 2100 -2875
rect 2330 -1305 2450 -1240
rect 2330 -1335 2375 -1305
rect 2405 -1335 2450 -1305
rect 2330 -1370 2450 -1335
rect 2330 -1400 2375 -1370
rect 2405 -1400 2450 -1370
rect 2330 -1440 2450 -1400
rect 2330 -1470 2375 -1440
rect 2405 -1470 2450 -1440
rect 2330 -1510 2450 -1470
rect 2330 -1540 2375 -1510
rect 2405 -1540 2450 -1510
rect 2330 -1580 2450 -1540
rect 2330 -1610 2375 -1580
rect 2405 -1610 2450 -1580
rect 2330 -1645 2450 -1610
rect 2330 -1675 2375 -1645
rect 2405 -1675 2450 -1645
rect 2330 -1705 2450 -1675
rect 2330 -1735 2375 -1705
rect 2405 -1735 2450 -1705
rect 2330 -1770 2450 -1735
rect 2330 -1800 2375 -1770
rect 2405 -1800 2450 -1770
rect 2330 -1840 2450 -1800
rect 2330 -1870 2375 -1840
rect 2405 -1870 2450 -1840
rect 2330 -1910 2450 -1870
rect 2330 -1940 2375 -1910
rect 2405 -1940 2450 -1910
rect 2330 -1980 2450 -1940
rect 2330 -2010 2375 -1980
rect 2405 -2010 2450 -1980
rect 2330 -2045 2450 -2010
rect 2330 -2075 2375 -2045
rect 2405 -2075 2450 -2045
rect 2330 -2105 2450 -2075
rect 2330 -2135 2375 -2105
rect 2405 -2135 2450 -2105
rect 2330 -2170 2450 -2135
rect 2330 -2200 2375 -2170
rect 2405 -2200 2450 -2170
rect 2330 -2240 2450 -2200
rect 2330 -2270 2375 -2240
rect 2405 -2270 2450 -2240
rect 2330 -2310 2450 -2270
rect 2330 -2340 2375 -2310
rect 2405 -2340 2450 -2310
rect 2330 -2380 2450 -2340
rect 2330 -2410 2375 -2380
rect 2405 -2410 2450 -2380
rect 2330 -2445 2450 -2410
rect 2330 -2475 2375 -2445
rect 2405 -2475 2450 -2445
rect 2330 -2505 2450 -2475
rect 2330 -2535 2375 -2505
rect 2405 -2535 2450 -2505
rect 2330 -2570 2450 -2535
rect 2330 -2600 2375 -2570
rect 2405 -2600 2450 -2570
rect 2330 -2640 2450 -2600
rect 2330 -2670 2375 -2640
rect 2405 -2670 2450 -2640
rect 2330 -2710 2450 -2670
rect 2330 -2740 2375 -2710
rect 2405 -2740 2450 -2710
rect 2330 -2780 2450 -2740
rect 2330 -2810 2375 -2780
rect 2405 -2810 2450 -2780
rect 2330 -2845 2450 -2810
rect 2330 -2875 2375 -2845
rect 2405 -2875 2450 -2845
rect 2330 -2890 2450 -2875
rect 2680 -1305 2800 -1240
rect 2680 -1335 2725 -1305
rect 2755 -1335 2800 -1305
rect 2680 -1370 2800 -1335
rect 2680 -1400 2725 -1370
rect 2755 -1400 2800 -1370
rect 2680 -1440 2800 -1400
rect 2680 -1470 2725 -1440
rect 2755 -1470 2800 -1440
rect 2680 -1510 2800 -1470
rect 2680 -1540 2725 -1510
rect 2755 -1540 2800 -1510
rect 2680 -1580 2800 -1540
rect 2680 -1610 2725 -1580
rect 2755 -1610 2800 -1580
rect 2680 -1645 2800 -1610
rect 2680 -1675 2725 -1645
rect 2755 -1675 2800 -1645
rect 2680 -1705 2800 -1675
rect 2680 -1735 2725 -1705
rect 2755 -1735 2800 -1705
rect 2680 -1770 2800 -1735
rect 2680 -1800 2725 -1770
rect 2755 -1800 2800 -1770
rect 2680 -1840 2800 -1800
rect 2680 -1870 2725 -1840
rect 2755 -1870 2800 -1840
rect 2680 -1910 2800 -1870
rect 2680 -1940 2725 -1910
rect 2755 -1940 2800 -1910
rect 2680 -1980 2800 -1940
rect 2680 -2010 2725 -1980
rect 2755 -2010 2800 -1980
rect 2680 -2045 2800 -2010
rect 2680 -2075 2725 -2045
rect 2755 -2075 2800 -2045
rect 2680 -2105 2800 -2075
rect 2680 -2135 2725 -2105
rect 2755 -2135 2800 -2105
rect 2680 -2170 2800 -2135
rect 2680 -2200 2725 -2170
rect 2755 -2200 2800 -2170
rect 2680 -2240 2800 -2200
rect 2680 -2270 2725 -2240
rect 2755 -2270 2800 -2240
rect 2680 -2310 2800 -2270
rect 2680 -2340 2725 -2310
rect 2755 -2340 2800 -2310
rect 2680 -2380 2800 -2340
rect 2680 -2410 2725 -2380
rect 2755 -2410 2800 -2380
rect 2680 -2445 2800 -2410
rect 2680 -2475 2725 -2445
rect 2755 -2475 2800 -2445
rect 2680 -2505 2800 -2475
rect 2680 -2535 2725 -2505
rect 2755 -2535 2800 -2505
rect 2680 -2570 2800 -2535
rect 2680 -2600 2725 -2570
rect 2755 -2600 2800 -2570
rect 2680 -2640 2800 -2600
rect 2680 -2670 2725 -2640
rect 2755 -2670 2800 -2640
rect 2680 -2710 2800 -2670
rect 2680 -2740 2725 -2710
rect 2755 -2740 2800 -2710
rect 2680 -2780 2800 -2740
rect 2680 -2810 2725 -2780
rect 2755 -2810 2800 -2780
rect 2680 -2845 2800 -2810
rect 2680 -2875 2725 -2845
rect 2755 -2875 2800 -2845
rect 2680 -2890 2800 -2875
rect 3030 -1305 3150 -1240
rect 3030 -1335 3075 -1305
rect 3105 -1335 3150 -1305
rect 3030 -1370 3150 -1335
rect 3030 -1400 3075 -1370
rect 3105 -1400 3150 -1370
rect 3030 -1440 3150 -1400
rect 3030 -1470 3075 -1440
rect 3105 -1470 3150 -1440
rect 3030 -1510 3150 -1470
rect 3030 -1540 3075 -1510
rect 3105 -1540 3150 -1510
rect 3030 -1580 3150 -1540
rect 3030 -1610 3075 -1580
rect 3105 -1610 3150 -1580
rect 3030 -1645 3150 -1610
rect 3030 -1675 3075 -1645
rect 3105 -1675 3150 -1645
rect 3030 -1705 3150 -1675
rect 3030 -1735 3075 -1705
rect 3105 -1735 3150 -1705
rect 3030 -1770 3150 -1735
rect 3030 -1800 3075 -1770
rect 3105 -1800 3150 -1770
rect 3030 -1840 3150 -1800
rect 3030 -1870 3075 -1840
rect 3105 -1870 3150 -1840
rect 3030 -1910 3150 -1870
rect 3030 -1940 3075 -1910
rect 3105 -1940 3150 -1910
rect 3030 -1980 3150 -1940
rect 3030 -2010 3075 -1980
rect 3105 -2010 3150 -1980
rect 3030 -2045 3150 -2010
rect 3030 -2075 3075 -2045
rect 3105 -2075 3150 -2045
rect 3030 -2105 3150 -2075
rect 3030 -2135 3075 -2105
rect 3105 -2135 3150 -2105
rect 3030 -2170 3150 -2135
rect 3030 -2200 3075 -2170
rect 3105 -2200 3150 -2170
rect 3030 -2240 3150 -2200
rect 3030 -2270 3075 -2240
rect 3105 -2270 3150 -2240
rect 3030 -2310 3150 -2270
rect 3030 -2340 3075 -2310
rect 3105 -2340 3150 -2310
rect 3030 -2380 3150 -2340
rect 3030 -2410 3075 -2380
rect 3105 -2410 3150 -2380
rect 3030 -2445 3150 -2410
rect 3030 -2475 3075 -2445
rect 3105 -2475 3150 -2445
rect 3030 -2505 3150 -2475
rect 3030 -2535 3075 -2505
rect 3105 -2535 3150 -2505
rect 3030 -2570 3150 -2535
rect 3030 -2600 3075 -2570
rect 3105 -2600 3150 -2570
rect 3030 -2640 3150 -2600
rect 3030 -2670 3075 -2640
rect 3105 -2670 3150 -2640
rect 3030 -2710 3150 -2670
rect 3030 -2740 3075 -2710
rect 3105 -2740 3150 -2710
rect 3030 -2780 3150 -2740
rect 3030 -2810 3075 -2780
rect 3105 -2810 3150 -2780
rect 3030 -2845 3150 -2810
rect 3030 -2875 3075 -2845
rect 3105 -2875 3150 -2845
rect 3030 -2890 3150 -2875
rect 3380 -1305 3500 -1240
rect 3380 -1335 3425 -1305
rect 3455 -1335 3500 -1305
rect 3380 -1370 3500 -1335
rect 3380 -1400 3425 -1370
rect 3455 -1400 3500 -1370
rect 3380 -1440 3500 -1400
rect 3380 -1470 3425 -1440
rect 3455 -1470 3500 -1440
rect 3380 -1510 3500 -1470
rect 3380 -1540 3425 -1510
rect 3455 -1540 3500 -1510
rect 3380 -1580 3500 -1540
rect 3380 -1610 3425 -1580
rect 3455 -1610 3500 -1580
rect 3380 -1645 3500 -1610
rect 3380 -1675 3425 -1645
rect 3455 -1675 3500 -1645
rect 3380 -1705 3500 -1675
rect 3380 -1735 3425 -1705
rect 3455 -1735 3500 -1705
rect 3380 -1770 3500 -1735
rect 3380 -1800 3425 -1770
rect 3455 -1800 3500 -1770
rect 3380 -1840 3500 -1800
rect 3380 -1870 3425 -1840
rect 3455 -1870 3500 -1840
rect 3380 -1910 3500 -1870
rect 3380 -1940 3425 -1910
rect 3455 -1940 3500 -1910
rect 3380 -1980 3500 -1940
rect 3380 -2010 3425 -1980
rect 3455 -2010 3500 -1980
rect 3380 -2045 3500 -2010
rect 3380 -2075 3425 -2045
rect 3455 -2075 3500 -2045
rect 3380 -2105 3500 -2075
rect 3380 -2135 3425 -2105
rect 3455 -2135 3500 -2105
rect 3380 -2170 3500 -2135
rect 3380 -2200 3425 -2170
rect 3455 -2200 3500 -2170
rect 3380 -2240 3500 -2200
rect 3380 -2270 3425 -2240
rect 3455 -2270 3500 -2240
rect 3380 -2310 3500 -2270
rect 3380 -2340 3425 -2310
rect 3455 -2340 3500 -2310
rect 3380 -2380 3500 -2340
rect 3380 -2410 3425 -2380
rect 3455 -2410 3500 -2380
rect 3380 -2445 3500 -2410
rect 3380 -2475 3425 -2445
rect 3455 -2475 3500 -2445
rect 3380 -2505 3500 -2475
rect 3380 -2535 3425 -2505
rect 3455 -2535 3500 -2505
rect 3380 -2570 3500 -2535
rect 3380 -2600 3425 -2570
rect 3455 -2600 3500 -2570
rect 3380 -2640 3500 -2600
rect 3380 -2670 3425 -2640
rect 3455 -2670 3500 -2640
rect 3380 -2710 3500 -2670
rect 3380 -2740 3425 -2710
rect 3455 -2740 3500 -2710
rect 3380 -2780 3500 -2740
rect 3380 -2810 3425 -2780
rect 3455 -2810 3500 -2780
rect 3380 -2845 3500 -2810
rect 3380 -2875 3425 -2845
rect 3455 -2875 3500 -2845
rect 3380 -2890 3500 -2875
rect 3730 -1305 3850 -1240
rect 3730 -1335 3775 -1305
rect 3805 -1335 3850 -1305
rect 3730 -1370 3850 -1335
rect 3730 -1400 3775 -1370
rect 3805 -1400 3850 -1370
rect 3730 -1440 3850 -1400
rect 3730 -1470 3775 -1440
rect 3805 -1470 3850 -1440
rect 3730 -1510 3850 -1470
rect 3730 -1540 3775 -1510
rect 3805 -1540 3850 -1510
rect 3730 -1580 3850 -1540
rect 3730 -1610 3775 -1580
rect 3805 -1610 3850 -1580
rect 3730 -1645 3850 -1610
rect 3730 -1675 3775 -1645
rect 3805 -1675 3850 -1645
rect 3730 -1705 3850 -1675
rect 3730 -1735 3775 -1705
rect 3805 -1735 3850 -1705
rect 3730 -1770 3850 -1735
rect 3730 -1800 3775 -1770
rect 3805 -1800 3850 -1770
rect 3730 -1840 3850 -1800
rect 3730 -1870 3775 -1840
rect 3805 -1870 3850 -1840
rect 3730 -1910 3850 -1870
rect 3730 -1940 3775 -1910
rect 3805 -1940 3850 -1910
rect 3730 -1980 3850 -1940
rect 3730 -2010 3775 -1980
rect 3805 -2010 3850 -1980
rect 3730 -2045 3850 -2010
rect 3730 -2075 3775 -2045
rect 3805 -2075 3850 -2045
rect 3730 -2105 3850 -2075
rect 3730 -2135 3775 -2105
rect 3805 -2135 3850 -2105
rect 3730 -2170 3850 -2135
rect 3730 -2200 3775 -2170
rect 3805 -2200 3850 -2170
rect 3730 -2240 3850 -2200
rect 3730 -2270 3775 -2240
rect 3805 -2270 3850 -2240
rect 3730 -2310 3850 -2270
rect 3730 -2340 3775 -2310
rect 3805 -2340 3850 -2310
rect 3730 -2380 3850 -2340
rect 3730 -2410 3775 -2380
rect 3805 -2410 3850 -2380
rect 3730 -2445 3850 -2410
rect 3730 -2475 3775 -2445
rect 3805 -2475 3850 -2445
rect 3730 -2505 3850 -2475
rect 3730 -2535 3775 -2505
rect 3805 -2535 3850 -2505
rect 3730 -2570 3850 -2535
rect 3730 -2600 3775 -2570
rect 3805 -2600 3850 -2570
rect 3730 -2640 3850 -2600
rect 3730 -2670 3775 -2640
rect 3805 -2670 3850 -2640
rect 3730 -2710 3850 -2670
rect 3730 -2740 3775 -2710
rect 3805 -2740 3850 -2710
rect 3730 -2780 3850 -2740
rect 3730 -2810 3775 -2780
rect 3805 -2810 3850 -2780
rect 3730 -2845 3850 -2810
rect 3730 -2875 3775 -2845
rect 3805 -2875 3850 -2845
rect 3730 -2890 3850 -2875
rect 4080 -1305 4200 -1240
rect 4080 -1335 4125 -1305
rect 4155 -1335 4200 -1305
rect 4080 -1370 4200 -1335
rect 4080 -1400 4125 -1370
rect 4155 -1400 4200 -1370
rect 4080 -1440 4200 -1400
rect 4080 -1470 4125 -1440
rect 4155 -1470 4200 -1440
rect 4080 -1510 4200 -1470
rect 4080 -1540 4125 -1510
rect 4155 -1540 4200 -1510
rect 4080 -1580 4200 -1540
rect 4080 -1610 4125 -1580
rect 4155 -1610 4200 -1580
rect 4080 -1645 4200 -1610
rect 4080 -1675 4125 -1645
rect 4155 -1675 4200 -1645
rect 4080 -1705 4200 -1675
rect 4080 -1735 4125 -1705
rect 4155 -1735 4200 -1705
rect 4080 -1770 4200 -1735
rect 4080 -1800 4125 -1770
rect 4155 -1800 4200 -1770
rect 4080 -1840 4200 -1800
rect 4080 -1870 4125 -1840
rect 4155 -1870 4200 -1840
rect 4080 -1910 4200 -1870
rect 4080 -1940 4125 -1910
rect 4155 -1940 4200 -1910
rect 4080 -1980 4200 -1940
rect 4080 -2010 4125 -1980
rect 4155 -2010 4200 -1980
rect 4080 -2045 4200 -2010
rect 4080 -2075 4125 -2045
rect 4155 -2075 4200 -2045
rect 4080 -2105 4200 -2075
rect 4080 -2135 4125 -2105
rect 4155 -2135 4200 -2105
rect 4080 -2170 4200 -2135
rect 4080 -2200 4125 -2170
rect 4155 -2200 4200 -2170
rect 4080 -2240 4200 -2200
rect 4080 -2270 4125 -2240
rect 4155 -2270 4200 -2240
rect 4080 -2310 4200 -2270
rect 4080 -2340 4125 -2310
rect 4155 -2340 4200 -2310
rect 4080 -2380 4200 -2340
rect 4080 -2410 4125 -2380
rect 4155 -2410 4200 -2380
rect 4080 -2445 4200 -2410
rect 4080 -2475 4125 -2445
rect 4155 -2475 4200 -2445
rect 4080 -2505 4200 -2475
rect 4080 -2535 4125 -2505
rect 4155 -2535 4200 -2505
rect 4080 -2570 4200 -2535
rect 4080 -2600 4125 -2570
rect 4155 -2600 4200 -2570
rect 4080 -2640 4200 -2600
rect 4080 -2670 4125 -2640
rect 4155 -2670 4200 -2640
rect 4080 -2710 4200 -2670
rect 4080 -2740 4125 -2710
rect 4155 -2740 4200 -2710
rect 4080 -2780 4200 -2740
rect 4080 -2810 4125 -2780
rect 4155 -2810 4200 -2780
rect 4080 -2845 4200 -2810
rect 4080 -2875 4125 -2845
rect 4155 -2875 4200 -2845
rect 4080 -2890 4200 -2875
rect 4430 -1305 4550 -1240
rect 4430 -1335 4475 -1305
rect 4505 -1335 4550 -1305
rect 4430 -1370 4550 -1335
rect 4430 -1400 4475 -1370
rect 4505 -1400 4550 -1370
rect 4430 -1440 4550 -1400
rect 4430 -1470 4475 -1440
rect 4505 -1470 4550 -1440
rect 4430 -1510 4550 -1470
rect 4430 -1540 4475 -1510
rect 4505 -1540 4550 -1510
rect 4430 -1580 4550 -1540
rect 4430 -1610 4475 -1580
rect 4505 -1610 4550 -1580
rect 4430 -1645 4550 -1610
rect 4430 -1675 4475 -1645
rect 4505 -1675 4550 -1645
rect 4430 -1705 4550 -1675
rect 4430 -1735 4475 -1705
rect 4505 -1735 4550 -1705
rect 4430 -1770 4550 -1735
rect 4430 -1800 4475 -1770
rect 4505 -1800 4550 -1770
rect 4430 -1840 4550 -1800
rect 4430 -1870 4475 -1840
rect 4505 -1870 4550 -1840
rect 4430 -1910 4550 -1870
rect 4430 -1940 4475 -1910
rect 4505 -1940 4550 -1910
rect 4430 -1980 4550 -1940
rect 4430 -2010 4475 -1980
rect 4505 -2010 4550 -1980
rect 4430 -2045 4550 -2010
rect 4430 -2075 4475 -2045
rect 4505 -2075 4550 -2045
rect 4430 -2105 4550 -2075
rect 4430 -2135 4475 -2105
rect 4505 -2135 4550 -2105
rect 4430 -2170 4550 -2135
rect 4430 -2200 4475 -2170
rect 4505 -2200 4550 -2170
rect 4430 -2240 4550 -2200
rect 4430 -2270 4475 -2240
rect 4505 -2270 4550 -2240
rect 4430 -2310 4550 -2270
rect 4430 -2340 4475 -2310
rect 4505 -2340 4550 -2310
rect 4430 -2380 4550 -2340
rect 4430 -2410 4475 -2380
rect 4505 -2410 4550 -2380
rect 4430 -2445 4550 -2410
rect 4430 -2475 4475 -2445
rect 4505 -2475 4550 -2445
rect 4430 -2505 4550 -2475
rect 4430 -2535 4475 -2505
rect 4505 -2535 4550 -2505
rect 4430 -2570 4550 -2535
rect 4430 -2600 4475 -2570
rect 4505 -2600 4550 -2570
rect 4430 -2640 4550 -2600
rect 4430 -2670 4475 -2640
rect 4505 -2670 4550 -2640
rect 4430 -2710 4550 -2670
rect 4430 -2740 4475 -2710
rect 4505 -2740 4550 -2710
rect 4430 -2780 4550 -2740
rect 4430 -2810 4475 -2780
rect 4505 -2810 4550 -2780
rect 4430 -2845 4550 -2810
rect 4430 -2875 4475 -2845
rect 4505 -2875 4550 -2845
rect 4430 -2890 4550 -2875
rect 4780 -1305 4900 -1240
rect 4780 -1335 4825 -1305
rect 4855 -1335 4900 -1305
rect 4780 -1370 4900 -1335
rect 4780 -1400 4825 -1370
rect 4855 -1400 4900 -1370
rect 4780 -1440 4900 -1400
rect 4780 -1470 4825 -1440
rect 4855 -1470 4900 -1440
rect 4780 -1510 4900 -1470
rect 4780 -1540 4825 -1510
rect 4855 -1540 4900 -1510
rect 4780 -1580 4900 -1540
rect 4780 -1610 4825 -1580
rect 4855 -1610 4900 -1580
rect 4780 -1645 4900 -1610
rect 4780 -1675 4825 -1645
rect 4855 -1675 4900 -1645
rect 4780 -1705 4900 -1675
rect 4780 -1735 4825 -1705
rect 4855 -1735 4900 -1705
rect 4780 -1770 4900 -1735
rect 4780 -1800 4825 -1770
rect 4855 -1800 4900 -1770
rect 4780 -1840 4900 -1800
rect 4780 -1870 4825 -1840
rect 4855 -1870 4900 -1840
rect 4780 -1910 4900 -1870
rect 4780 -1940 4825 -1910
rect 4855 -1940 4900 -1910
rect 4780 -1980 4900 -1940
rect 4780 -2010 4825 -1980
rect 4855 -2010 4900 -1980
rect 4780 -2045 4900 -2010
rect 4780 -2075 4825 -2045
rect 4855 -2075 4900 -2045
rect 4780 -2105 4900 -2075
rect 4780 -2135 4825 -2105
rect 4855 -2135 4900 -2105
rect 4780 -2170 4900 -2135
rect 4780 -2200 4825 -2170
rect 4855 -2200 4900 -2170
rect 4780 -2240 4900 -2200
rect 4780 -2270 4825 -2240
rect 4855 -2270 4900 -2240
rect 4780 -2310 4900 -2270
rect 4780 -2340 4825 -2310
rect 4855 -2340 4900 -2310
rect 4780 -2380 4900 -2340
rect 4780 -2410 4825 -2380
rect 4855 -2410 4900 -2380
rect 4780 -2445 4900 -2410
rect 4780 -2475 4825 -2445
rect 4855 -2475 4900 -2445
rect 4780 -2505 4900 -2475
rect 4780 -2535 4825 -2505
rect 4855 -2535 4900 -2505
rect 4780 -2570 4900 -2535
rect 4780 -2600 4825 -2570
rect 4855 -2600 4900 -2570
rect 4780 -2640 4900 -2600
rect 4780 -2670 4825 -2640
rect 4855 -2670 4900 -2640
rect 4780 -2710 4900 -2670
rect 4780 -2740 4825 -2710
rect 4855 -2740 4900 -2710
rect 4780 -2780 4900 -2740
rect 4780 -2810 4825 -2780
rect 4855 -2810 4900 -2780
rect 4780 -2845 4900 -2810
rect 4780 -2875 4825 -2845
rect 4855 -2875 4900 -2845
rect 4780 -2890 4900 -2875
rect 5130 -1305 5250 -1240
rect 5130 -1335 5175 -1305
rect 5205 -1335 5250 -1305
rect 5130 -1370 5250 -1335
rect 5130 -1400 5175 -1370
rect 5205 -1400 5250 -1370
rect 5130 -1440 5250 -1400
rect 5130 -1470 5175 -1440
rect 5205 -1470 5250 -1440
rect 5130 -1510 5250 -1470
rect 5130 -1540 5175 -1510
rect 5205 -1540 5250 -1510
rect 5130 -1580 5250 -1540
rect 5130 -1610 5175 -1580
rect 5205 -1610 5250 -1580
rect 5130 -1645 5250 -1610
rect 5130 -1675 5175 -1645
rect 5205 -1675 5250 -1645
rect 5130 -1705 5250 -1675
rect 5130 -1735 5175 -1705
rect 5205 -1735 5250 -1705
rect 5130 -1770 5250 -1735
rect 5130 -1800 5175 -1770
rect 5205 -1800 5250 -1770
rect 5130 -1840 5250 -1800
rect 5130 -1870 5175 -1840
rect 5205 -1870 5250 -1840
rect 5130 -1910 5250 -1870
rect 5130 -1940 5175 -1910
rect 5205 -1940 5250 -1910
rect 5130 -1980 5250 -1940
rect 5130 -2010 5175 -1980
rect 5205 -2010 5250 -1980
rect 5130 -2045 5250 -2010
rect 5130 -2075 5175 -2045
rect 5205 -2075 5250 -2045
rect 5130 -2105 5250 -2075
rect 5130 -2135 5175 -2105
rect 5205 -2135 5250 -2105
rect 5130 -2170 5250 -2135
rect 5130 -2200 5175 -2170
rect 5205 -2200 5250 -2170
rect 5130 -2240 5250 -2200
rect 5130 -2270 5175 -2240
rect 5205 -2270 5250 -2240
rect 5130 -2310 5250 -2270
rect 5130 -2340 5175 -2310
rect 5205 -2340 5250 -2310
rect 5130 -2380 5250 -2340
rect 5130 -2410 5175 -2380
rect 5205 -2410 5250 -2380
rect 5130 -2445 5250 -2410
rect 5130 -2475 5175 -2445
rect 5205 -2475 5250 -2445
rect 5130 -2505 5250 -2475
rect 5130 -2535 5175 -2505
rect 5205 -2535 5250 -2505
rect 5130 -2570 5250 -2535
rect 5130 -2600 5175 -2570
rect 5205 -2600 5250 -2570
rect 5130 -2640 5250 -2600
rect 5130 -2670 5175 -2640
rect 5205 -2670 5250 -2640
rect 5130 -2710 5250 -2670
rect 5130 -2740 5175 -2710
rect 5205 -2740 5250 -2710
rect 5130 -2780 5250 -2740
rect 5130 -2810 5175 -2780
rect 5205 -2810 5250 -2780
rect 5130 -2845 5250 -2810
rect 5130 -2875 5175 -2845
rect 5205 -2875 5250 -2845
rect 5130 -2890 5250 -2875
rect 5480 -1305 5600 -1240
rect 5480 -1335 5525 -1305
rect 5555 -1335 5600 -1305
rect 5480 -1370 5600 -1335
rect 5480 -1400 5525 -1370
rect 5555 -1400 5600 -1370
rect 5480 -1440 5600 -1400
rect 5480 -1470 5525 -1440
rect 5555 -1470 5600 -1440
rect 5480 -1510 5600 -1470
rect 5480 -1540 5525 -1510
rect 5555 -1540 5600 -1510
rect 5480 -1580 5600 -1540
rect 5480 -1610 5525 -1580
rect 5555 -1610 5600 -1580
rect 5480 -1645 5600 -1610
rect 5480 -1675 5525 -1645
rect 5555 -1675 5600 -1645
rect 5480 -1705 5600 -1675
rect 5480 -1735 5525 -1705
rect 5555 -1735 5600 -1705
rect 5480 -1770 5600 -1735
rect 5480 -1800 5525 -1770
rect 5555 -1800 5600 -1770
rect 5480 -1840 5600 -1800
rect 5480 -1870 5525 -1840
rect 5555 -1870 5600 -1840
rect 5480 -1910 5600 -1870
rect 5480 -1940 5525 -1910
rect 5555 -1940 5600 -1910
rect 5480 -1980 5600 -1940
rect 5480 -2010 5525 -1980
rect 5555 -2010 5600 -1980
rect 5480 -2045 5600 -2010
rect 5480 -2075 5525 -2045
rect 5555 -2075 5600 -2045
rect 5480 -2105 5600 -2075
rect 5480 -2135 5525 -2105
rect 5555 -2135 5600 -2105
rect 5480 -2170 5600 -2135
rect 5480 -2200 5525 -2170
rect 5555 -2200 5600 -2170
rect 5480 -2240 5600 -2200
rect 5480 -2270 5525 -2240
rect 5555 -2270 5600 -2240
rect 5480 -2310 5600 -2270
rect 5480 -2340 5525 -2310
rect 5555 -2340 5600 -2310
rect 5480 -2380 5600 -2340
rect 5480 -2410 5525 -2380
rect 5555 -2410 5600 -2380
rect 5480 -2445 5600 -2410
rect 5480 -2475 5525 -2445
rect 5555 -2475 5600 -2445
rect 5480 -2505 5600 -2475
rect 5480 -2535 5525 -2505
rect 5555 -2535 5600 -2505
rect 5480 -2570 5600 -2535
rect 5480 -2600 5525 -2570
rect 5555 -2600 5600 -2570
rect 5480 -2640 5600 -2600
rect 5480 -2670 5525 -2640
rect 5555 -2670 5600 -2640
rect 5480 -2710 5600 -2670
rect 5480 -2740 5525 -2710
rect 5555 -2740 5600 -2710
rect 5480 -2780 5600 -2740
rect 5480 -2810 5525 -2780
rect 5555 -2810 5600 -2780
rect 5480 -2845 5600 -2810
rect 5480 -2875 5525 -2845
rect 5555 -2875 5600 -2845
rect 5480 -2890 5600 -2875
rect 5830 -1305 5950 -1240
rect 5830 -1335 5875 -1305
rect 5905 -1335 5950 -1305
rect 5830 -1370 5950 -1335
rect 5830 -1400 5875 -1370
rect 5905 -1400 5950 -1370
rect 5830 -1440 5950 -1400
rect 5830 -1470 5875 -1440
rect 5905 -1470 5950 -1440
rect 5830 -1510 5950 -1470
rect 5830 -1540 5875 -1510
rect 5905 -1540 5950 -1510
rect 5830 -1580 5950 -1540
rect 5830 -1610 5875 -1580
rect 5905 -1610 5950 -1580
rect 5830 -1645 5950 -1610
rect 5830 -1675 5875 -1645
rect 5905 -1675 5950 -1645
rect 5830 -1705 5950 -1675
rect 5830 -1735 5875 -1705
rect 5905 -1735 5950 -1705
rect 5830 -1770 5950 -1735
rect 5830 -1800 5875 -1770
rect 5905 -1800 5950 -1770
rect 5830 -1840 5950 -1800
rect 5830 -1870 5875 -1840
rect 5905 -1870 5950 -1840
rect 5830 -1910 5950 -1870
rect 5830 -1940 5875 -1910
rect 5905 -1940 5950 -1910
rect 5830 -1980 5950 -1940
rect 5830 -2010 5875 -1980
rect 5905 -2010 5950 -1980
rect 5830 -2045 5950 -2010
rect 5830 -2075 5875 -2045
rect 5905 -2075 5950 -2045
rect 5830 -2105 5950 -2075
rect 5830 -2135 5875 -2105
rect 5905 -2135 5950 -2105
rect 5830 -2170 5950 -2135
rect 5830 -2200 5875 -2170
rect 5905 -2200 5950 -2170
rect 5830 -2240 5950 -2200
rect 5830 -2270 5875 -2240
rect 5905 -2270 5950 -2240
rect 5830 -2310 5950 -2270
rect 5830 -2340 5875 -2310
rect 5905 -2340 5950 -2310
rect 5830 -2380 5950 -2340
rect 5830 -2410 5875 -2380
rect 5905 -2410 5950 -2380
rect 5830 -2445 5950 -2410
rect 5830 -2475 5875 -2445
rect 5905 -2475 5950 -2445
rect 5830 -2505 5950 -2475
rect 5830 -2535 5875 -2505
rect 5905 -2535 5950 -2505
rect 5830 -2570 5950 -2535
rect 5830 -2600 5875 -2570
rect 5905 -2600 5950 -2570
rect 5830 -2640 5950 -2600
rect 5830 -2670 5875 -2640
rect 5905 -2670 5950 -2640
rect 5830 -2710 5950 -2670
rect 5830 -2740 5875 -2710
rect 5905 -2740 5950 -2710
rect 5830 -2780 5950 -2740
rect 5830 -2810 5875 -2780
rect 5905 -2810 5950 -2780
rect 5830 -2845 5950 -2810
rect 5830 -2875 5875 -2845
rect 5905 -2875 5950 -2845
rect 5830 -2890 5950 -2875
rect 6180 -1305 6300 -1240
rect 6180 -1335 6225 -1305
rect 6255 -1335 6300 -1305
rect 6180 -1370 6300 -1335
rect 6180 -1400 6225 -1370
rect 6255 -1400 6300 -1370
rect 6180 -1440 6300 -1400
rect 6180 -1470 6225 -1440
rect 6255 -1470 6300 -1440
rect 6180 -1510 6300 -1470
rect 6180 -1540 6225 -1510
rect 6255 -1540 6300 -1510
rect 6180 -1580 6300 -1540
rect 6180 -1610 6225 -1580
rect 6255 -1610 6300 -1580
rect 6180 -1645 6300 -1610
rect 6180 -1675 6225 -1645
rect 6255 -1675 6300 -1645
rect 6180 -1705 6300 -1675
rect 6180 -1735 6225 -1705
rect 6255 -1735 6300 -1705
rect 6180 -1770 6300 -1735
rect 6180 -1800 6225 -1770
rect 6255 -1800 6300 -1770
rect 6180 -1840 6300 -1800
rect 6180 -1870 6225 -1840
rect 6255 -1870 6300 -1840
rect 6180 -1910 6300 -1870
rect 6180 -1940 6225 -1910
rect 6255 -1940 6300 -1910
rect 6180 -1980 6300 -1940
rect 6180 -2010 6225 -1980
rect 6255 -2010 6300 -1980
rect 6180 -2045 6300 -2010
rect 6180 -2075 6225 -2045
rect 6255 -2075 6300 -2045
rect 6180 -2105 6300 -2075
rect 6180 -2135 6225 -2105
rect 6255 -2135 6300 -2105
rect 6180 -2170 6300 -2135
rect 6180 -2200 6225 -2170
rect 6255 -2200 6300 -2170
rect 6180 -2240 6300 -2200
rect 6180 -2270 6225 -2240
rect 6255 -2270 6300 -2240
rect 6180 -2310 6300 -2270
rect 6180 -2340 6225 -2310
rect 6255 -2340 6300 -2310
rect 6180 -2380 6300 -2340
rect 6180 -2410 6225 -2380
rect 6255 -2410 6300 -2380
rect 6180 -2445 6300 -2410
rect 6180 -2475 6225 -2445
rect 6255 -2475 6300 -2445
rect 6180 -2505 6300 -2475
rect 6180 -2535 6225 -2505
rect 6255 -2535 6300 -2505
rect 6180 -2570 6300 -2535
rect 6180 -2600 6225 -2570
rect 6255 -2600 6300 -2570
rect 6180 -2640 6300 -2600
rect 6180 -2670 6225 -2640
rect 6255 -2670 6300 -2640
rect 6180 -2710 6300 -2670
rect 6180 -2740 6225 -2710
rect 6255 -2740 6300 -2710
rect 6180 -2780 6300 -2740
rect 6180 -2810 6225 -2780
rect 6255 -2810 6300 -2780
rect 6180 -2845 6300 -2810
rect 6180 -2875 6225 -2845
rect 6255 -2875 6300 -2845
rect 6180 -2890 6300 -2875
rect 6530 -1305 6650 -1240
rect 6530 -1335 6575 -1305
rect 6605 -1335 6650 -1305
rect 6530 -1370 6650 -1335
rect 6530 -1400 6575 -1370
rect 6605 -1400 6650 -1370
rect 6530 -1440 6650 -1400
rect 6530 -1470 6575 -1440
rect 6605 -1470 6650 -1440
rect 6530 -1510 6650 -1470
rect 6530 -1540 6575 -1510
rect 6605 -1540 6650 -1510
rect 6530 -1580 6650 -1540
rect 6530 -1610 6575 -1580
rect 6605 -1610 6650 -1580
rect 6530 -1645 6650 -1610
rect 6530 -1675 6575 -1645
rect 6605 -1675 6650 -1645
rect 6530 -1705 6650 -1675
rect 6530 -1735 6575 -1705
rect 6605 -1735 6650 -1705
rect 6530 -1770 6650 -1735
rect 6530 -1800 6575 -1770
rect 6605 -1800 6650 -1770
rect 6530 -1840 6650 -1800
rect 6530 -1870 6575 -1840
rect 6605 -1870 6650 -1840
rect 6530 -1910 6650 -1870
rect 6530 -1940 6575 -1910
rect 6605 -1940 6650 -1910
rect 6530 -1980 6650 -1940
rect 6530 -2010 6575 -1980
rect 6605 -2010 6650 -1980
rect 6530 -2045 6650 -2010
rect 6530 -2075 6575 -2045
rect 6605 -2075 6650 -2045
rect 6530 -2105 6650 -2075
rect 6530 -2135 6575 -2105
rect 6605 -2135 6650 -2105
rect 6530 -2170 6650 -2135
rect 6530 -2200 6575 -2170
rect 6605 -2200 6650 -2170
rect 6530 -2240 6650 -2200
rect 6530 -2270 6575 -2240
rect 6605 -2270 6650 -2240
rect 6530 -2310 6650 -2270
rect 6530 -2340 6575 -2310
rect 6605 -2340 6650 -2310
rect 6530 -2380 6650 -2340
rect 6530 -2410 6575 -2380
rect 6605 -2410 6650 -2380
rect 6530 -2445 6650 -2410
rect 6530 -2475 6575 -2445
rect 6605 -2475 6650 -2445
rect 6530 -2505 6650 -2475
rect 6530 -2535 6575 -2505
rect 6605 -2535 6650 -2505
rect 6530 -2570 6650 -2535
rect 6530 -2600 6575 -2570
rect 6605 -2600 6650 -2570
rect 6530 -2640 6650 -2600
rect 6530 -2670 6575 -2640
rect 6605 -2670 6650 -2640
rect 6530 -2710 6650 -2670
rect 6530 -2740 6575 -2710
rect 6605 -2740 6650 -2710
rect 6530 -2780 6650 -2740
rect 6530 -2810 6575 -2780
rect 6605 -2810 6650 -2780
rect 6530 -2845 6650 -2810
rect 6530 -2875 6575 -2845
rect 6605 -2875 6650 -2845
rect 6530 -2890 6650 -2875
rect 6880 -1305 7000 -1240
rect 6880 -1335 6925 -1305
rect 6955 -1335 7000 -1305
rect 6880 -1370 7000 -1335
rect 6880 -1400 6925 -1370
rect 6955 -1400 7000 -1370
rect 6880 -1440 7000 -1400
rect 6880 -1470 6925 -1440
rect 6955 -1470 7000 -1440
rect 6880 -1510 7000 -1470
rect 6880 -1540 6925 -1510
rect 6955 -1540 7000 -1510
rect 6880 -1580 7000 -1540
rect 6880 -1610 6925 -1580
rect 6955 -1610 7000 -1580
rect 6880 -1645 7000 -1610
rect 6880 -1675 6925 -1645
rect 6955 -1675 7000 -1645
rect 6880 -1705 7000 -1675
rect 6880 -1735 6925 -1705
rect 6955 -1735 7000 -1705
rect 6880 -1770 7000 -1735
rect 6880 -1800 6925 -1770
rect 6955 -1800 7000 -1770
rect 6880 -1840 7000 -1800
rect 6880 -1870 6925 -1840
rect 6955 -1870 7000 -1840
rect 6880 -1910 7000 -1870
rect 6880 -1940 6925 -1910
rect 6955 -1940 7000 -1910
rect 6880 -1980 7000 -1940
rect 6880 -2010 6925 -1980
rect 6955 -2010 7000 -1980
rect 6880 -2045 7000 -2010
rect 6880 -2075 6925 -2045
rect 6955 -2075 7000 -2045
rect 6880 -2105 7000 -2075
rect 6880 -2135 6925 -2105
rect 6955 -2135 7000 -2105
rect 6880 -2170 7000 -2135
rect 6880 -2200 6925 -2170
rect 6955 -2200 7000 -2170
rect 6880 -2240 7000 -2200
rect 6880 -2270 6925 -2240
rect 6955 -2270 7000 -2240
rect 6880 -2310 7000 -2270
rect 6880 -2340 6925 -2310
rect 6955 -2340 7000 -2310
rect 6880 -2380 7000 -2340
rect 6880 -2410 6925 -2380
rect 6955 -2410 7000 -2380
rect 6880 -2445 7000 -2410
rect 6880 -2475 6925 -2445
rect 6955 -2475 7000 -2445
rect 6880 -2505 7000 -2475
rect 6880 -2535 6925 -2505
rect 6955 -2535 7000 -2505
rect 6880 -2570 7000 -2535
rect 6880 -2600 6925 -2570
rect 6955 -2600 7000 -2570
rect 6880 -2640 7000 -2600
rect 6880 -2670 6925 -2640
rect 6955 -2670 7000 -2640
rect 6880 -2710 7000 -2670
rect 6880 -2740 6925 -2710
rect 6955 -2740 7000 -2710
rect 6880 -2780 7000 -2740
rect 6880 -2810 6925 -2780
rect 6955 -2810 7000 -2780
rect 6880 -2845 7000 -2810
rect 6880 -2875 6925 -2845
rect 6955 -2875 7000 -2845
rect 6880 -2890 7000 -2875
rect 7230 -1305 7350 -1240
rect 7230 -1335 7275 -1305
rect 7305 -1335 7350 -1305
rect 7230 -1370 7350 -1335
rect 7230 -1400 7275 -1370
rect 7305 -1400 7350 -1370
rect 7230 -1440 7350 -1400
rect 7230 -1470 7275 -1440
rect 7305 -1470 7350 -1440
rect 7230 -1510 7350 -1470
rect 7230 -1540 7275 -1510
rect 7305 -1540 7350 -1510
rect 7230 -1580 7350 -1540
rect 7230 -1610 7275 -1580
rect 7305 -1610 7350 -1580
rect 7230 -1645 7350 -1610
rect 7230 -1675 7275 -1645
rect 7305 -1675 7350 -1645
rect 7230 -1705 7350 -1675
rect 7230 -1735 7275 -1705
rect 7305 -1735 7350 -1705
rect 7230 -1770 7350 -1735
rect 7230 -1800 7275 -1770
rect 7305 -1800 7350 -1770
rect 7230 -1840 7350 -1800
rect 7230 -1870 7275 -1840
rect 7305 -1870 7350 -1840
rect 7230 -1910 7350 -1870
rect 7230 -1940 7275 -1910
rect 7305 -1940 7350 -1910
rect 7230 -1980 7350 -1940
rect 7230 -2010 7275 -1980
rect 7305 -2010 7350 -1980
rect 7230 -2045 7350 -2010
rect 7230 -2075 7275 -2045
rect 7305 -2075 7350 -2045
rect 7230 -2105 7350 -2075
rect 7230 -2135 7275 -2105
rect 7305 -2135 7350 -2105
rect 7230 -2170 7350 -2135
rect 7230 -2200 7275 -2170
rect 7305 -2200 7350 -2170
rect 7230 -2240 7350 -2200
rect 7230 -2270 7275 -2240
rect 7305 -2270 7350 -2240
rect 7230 -2310 7350 -2270
rect 7230 -2340 7275 -2310
rect 7305 -2340 7350 -2310
rect 7230 -2380 7350 -2340
rect 7230 -2410 7275 -2380
rect 7305 -2410 7350 -2380
rect 7230 -2445 7350 -2410
rect 7230 -2475 7275 -2445
rect 7305 -2475 7350 -2445
rect 7230 -2505 7350 -2475
rect 7230 -2535 7275 -2505
rect 7305 -2535 7350 -2505
rect 7230 -2570 7350 -2535
rect 7230 -2600 7275 -2570
rect 7305 -2600 7350 -2570
rect 7230 -2640 7350 -2600
rect 7230 -2670 7275 -2640
rect 7305 -2670 7350 -2640
rect 7230 -2710 7350 -2670
rect 7230 -2740 7275 -2710
rect 7305 -2740 7350 -2710
rect 7230 -2780 7350 -2740
rect 7230 -2810 7275 -2780
rect 7305 -2810 7350 -2780
rect 7230 -2845 7350 -2810
rect 7230 -2875 7275 -2845
rect 7305 -2875 7350 -2845
rect 7230 -2890 7350 -2875
rect 7580 -1305 7700 -1240
rect 7580 -1335 7625 -1305
rect 7655 -1335 7700 -1305
rect 7580 -1370 7700 -1335
rect 7580 -1400 7625 -1370
rect 7655 -1400 7700 -1370
rect 7580 -1440 7700 -1400
rect 7580 -1470 7625 -1440
rect 7655 -1470 7700 -1440
rect 7580 -1510 7700 -1470
rect 7580 -1540 7625 -1510
rect 7655 -1540 7700 -1510
rect 7580 -1580 7700 -1540
rect 7580 -1610 7625 -1580
rect 7655 -1610 7700 -1580
rect 7580 -1645 7700 -1610
rect 7580 -1675 7625 -1645
rect 7655 -1675 7700 -1645
rect 7580 -1705 7700 -1675
rect 7580 -1735 7625 -1705
rect 7655 -1735 7700 -1705
rect 7580 -1770 7700 -1735
rect 7580 -1800 7625 -1770
rect 7655 -1800 7700 -1770
rect 7580 -1840 7700 -1800
rect 7580 -1870 7625 -1840
rect 7655 -1870 7700 -1840
rect 7580 -1910 7700 -1870
rect 7580 -1940 7625 -1910
rect 7655 -1940 7700 -1910
rect 7580 -1980 7700 -1940
rect 7580 -2010 7625 -1980
rect 7655 -2010 7700 -1980
rect 7580 -2045 7700 -2010
rect 7580 -2075 7625 -2045
rect 7655 -2075 7700 -2045
rect 7580 -2105 7700 -2075
rect 7580 -2135 7625 -2105
rect 7655 -2135 7700 -2105
rect 7580 -2170 7700 -2135
rect 7580 -2200 7625 -2170
rect 7655 -2200 7700 -2170
rect 7580 -2240 7700 -2200
rect 7580 -2270 7625 -2240
rect 7655 -2270 7700 -2240
rect 7580 -2310 7700 -2270
rect 7580 -2340 7625 -2310
rect 7655 -2340 7700 -2310
rect 7580 -2380 7700 -2340
rect 7580 -2410 7625 -2380
rect 7655 -2410 7700 -2380
rect 7580 -2445 7700 -2410
rect 7580 -2475 7625 -2445
rect 7655 -2475 7700 -2445
rect 7580 -2505 7700 -2475
rect 7580 -2535 7625 -2505
rect 7655 -2535 7700 -2505
rect 7580 -2570 7700 -2535
rect 7580 -2600 7625 -2570
rect 7655 -2600 7700 -2570
rect 7580 -2640 7700 -2600
rect 7580 -2670 7625 -2640
rect 7655 -2670 7700 -2640
rect 7580 -2710 7700 -2670
rect 7580 -2740 7625 -2710
rect 7655 -2740 7700 -2710
rect 7580 -2780 7700 -2740
rect 7580 -2810 7625 -2780
rect 7655 -2810 7700 -2780
rect 7580 -2845 7700 -2810
rect 7580 -2875 7625 -2845
rect 7655 -2875 7700 -2845
rect 7580 -2890 7700 -2875
rect 7930 -1305 8050 -1240
rect 7930 -1335 7975 -1305
rect 8005 -1335 8050 -1305
rect 7930 -1370 8050 -1335
rect 7930 -1400 7975 -1370
rect 8005 -1400 8050 -1370
rect 7930 -1440 8050 -1400
rect 7930 -1470 7975 -1440
rect 8005 -1470 8050 -1440
rect 7930 -1510 8050 -1470
rect 7930 -1540 7975 -1510
rect 8005 -1540 8050 -1510
rect 7930 -1580 8050 -1540
rect 7930 -1610 7975 -1580
rect 8005 -1610 8050 -1580
rect 7930 -1645 8050 -1610
rect 7930 -1675 7975 -1645
rect 8005 -1675 8050 -1645
rect 7930 -1705 8050 -1675
rect 7930 -1735 7975 -1705
rect 8005 -1735 8050 -1705
rect 7930 -1770 8050 -1735
rect 7930 -1800 7975 -1770
rect 8005 -1800 8050 -1770
rect 7930 -1840 8050 -1800
rect 7930 -1870 7975 -1840
rect 8005 -1870 8050 -1840
rect 7930 -1910 8050 -1870
rect 7930 -1940 7975 -1910
rect 8005 -1940 8050 -1910
rect 7930 -1980 8050 -1940
rect 7930 -2010 7975 -1980
rect 8005 -2010 8050 -1980
rect 7930 -2045 8050 -2010
rect 7930 -2075 7975 -2045
rect 8005 -2075 8050 -2045
rect 7930 -2105 8050 -2075
rect 7930 -2135 7975 -2105
rect 8005 -2135 8050 -2105
rect 7930 -2170 8050 -2135
rect 7930 -2200 7975 -2170
rect 8005 -2200 8050 -2170
rect 7930 -2240 8050 -2200
rect 7930 -2270 7975 -2240
rect 8005 -2270 8050 -2240
rect 7930 -2310 8050 -2270
rect 7930 -2340 7975 -2310
rect 8005 -2340 8050 -2310
rect 7930 -2380 8050 -2340
rect 7930 -2410 7975 -2380
rect 8005 -2410 8050 -2380
rect 7930 -2445 8050 -2410
rect 7930 -2475 7975 -2445
rect 8005 -2475 8050 -2445
rect 7930 -2505 8050 -2475
rect 7930 -2535 7975 -2505
rect 8005 -2535 8050 -2505
rect 7930 -2570 8050 -2535
rect 7930 -2600 7975 -2570
rect 8005 -2600 8050 -2570
rect 7930 -2640 8050 -2600
rect 7930 -2670 7975 -2640
rect 8005 -2670 8050 -2640
rect 7930 -2710 8050 -2670
rect 7930 -2740 7975 -2710
rect 8005 -2740 8050 -2710
rect 7930 -2780 8050 -2740
rect 7930 -2810 7975 -2780
rect 8005 -2810 8050 -2780
rect 7930 -2845 8050 -2810
rect 7930 -2875 7975 -2845
rect 8005 -2875 8050 -2845
rect 7930 -2890 8050 -2875
rect 8280 -1305 8400 -1240
rect 8280 -1335 8325 -1305
rect 8355 -1335 8400 -1305
rect 8280 -1370 8400 -1335
rect 8280 -1400 8325 -1370
rect 8355 -1400 8400 -1370
rect 8280 -1440 8400 -1400
rect 8280 -1470 8325 -1440
rect 8355 -1470 8400 -1440
rect 8280 -1510 8400 -1470
rect 8280 -1540 8325 -1510
rect 8355 -1540 8400 -1510
rect 8280 -1580 8400 -1540
rect 8280 -1610 8325 -1580
rect 8355 -1610 8400 -1580
rect 8280 -1645 8400 -1610
rect 8280 -1675 8325 -1645
rect 8355 -1675 8400 -1645
rect 8280 -1705 8400 -1675
rect 8280 -1735 8325 -1705
rect 8355 -1735 8400 -1705
rect 8280 -1770 8400 -1735
rect 8280 -1800 8325 -1770
rect 8355 -1800 8400 -1770
rect 8280 -1840 8400 -1800
rect 8280 -1870 8325 -1840
rect 8355 -1870 8400 -1840
rect 8280 -1910 8400 -1870
rect 8280 -1940 8325 -1910
rect 8355 -1940 8400 -1910
rect 8280 -1980 8400 -1940
rect 8280 -2010 8325 -1980
rect 8355 -2010 8400 -1980
rect 8280 -2045 8400 -2010
rect 8280 -2075 8325 -2045
rect 8355 -2075 8400 -2045
rect 8280 -2105 8400 -2075
rect 8280 -2135 8325 -2105
rect 8355 -2135 8400 -2105
rect 8280 -2170 8400 -2135
rect 8280 -2200 8325 -2170
rect 8355 -2200 8400 -2170
rect 8280 -2240 8400 -2200
rect 8280 -2270 8325 -2240
rect 8355 -2270 8400 -2240
rect 8280 -2310 8400 -2270
rect 8280 -2340 8325 -2310
rect 8355 -2340 8400 -2310
rect 8280 -2380 8400 -2340
rect 8280 -2410 8325 -2380
rect 8355 -2410 8400 -2380
rect 8280 -2445 8400 -2410
rect 8280 -2475 8325 -2445
rect 8355 -2475 8400 -2445
rect 8280 -2505 8400 -2475
rect 8280 -2535 8325 -2505
rect 8355 -2535 8400 -2505
rect 8280 -2570 8400 -2535
rect 8280 -2600 8325 -2570
rect 8355 -2600 8400 -2570
rect 8280 -2640 8400 -2600
rect 8280 -2670 8325 -2640
rect 8355 -2670 8400 -2640
rect 8280 -2710 8400 -2670
rect 8280 -2740 8325 -2710
rect 8355 -2740 8400 -2710
rect 8280 -2780 8400 -2740
rect 8280 -2810 8325 -2780
rect 8355 -2810 8400 -2780
rect 8280 -2845 8400 -2810
rect 8280 -2875 8325 -2845
rect 8355 -2875 8400 -2845
rect 8280 -2890 8400 -2875
rect 8630 -1305 8750 -1240
rect 8630 -1335 8675 -1305
rect 8705 -1335 8750 -1305
rect 8630 -1370 8750 -1335
rect 8630 -1400 8675 -1370
rect 8705 -1400 8750 -1370
rect 8630 -1440 8750 -1400
rect 8630 -1470 8675 -1440
rect 8705 -1470 8750 -1440
rect 8630 -1510 8750 -1470
rect 8630 -1540 8675 -1510
rect 8705 -1540 8750 -1510
rect 8630 -1580 8750 -1540
rect 8630 -1610 8675 -1580
rect 8705 -1610 8750 -1580
rect 8630 -1645 8750 -1610
rect 8630 -1675 8675 -1645
rect 8705 -1675 8750 -1645
rect 8630 -1705 8750 -1675
rect 8630 -1735 8675 -1705
rect 8705 -1735 8750 -1705
rect 8630 -1770 8750 -1735
rect 8630 -1800 8675 -1770
rect 8705 -1800 8750 -1770
rect 8630 -1840 8750 -1800
rect 8630 -1870 8675 -1840
rect 8705 -1870 8750 -1840
rect 8630 -1910 8750 -1870
rect 8630 -1940 8675 -1910
rect 8705 -1940 8750 -1910
rect 8630 -1980 8750 -1940
rect 8630 -2010 8675 -1980
rect 8705 -2010 8750 -1980
rect 8630 -2045 8750 -2010
rect 8630 -2075 8675 -2045
rect 8705 -2075 8750 -2045
rect 8630 -2105 8750 -2075
rect 8630 -2135 8675 -2105
rect 8705 -2135 8750 -2105
rect 8630 -2170 8750 -2135
rect 8630 -2200 8675 -2170
rect 8705 -2200 8750 -2170
rect 8630 -2240 8750 -2200
rect 8630 -2270 8675 -2240
rect 8705 -2270 8750 -2240
rect 8630 -2310 8750 -2270
rect 8630 -2340 8675 -2310
rect 8705 -2340 8750 -2310
rect 8630 -2380 8750 -2340
rect 8630 -2410 8675 -2380
rect 8705 -2410 8750 -2380
rect 8630 -2445 8750 -2410
rect 8630 -2475 8675 -2445
rect 8705 -2475 8750 -2445
rect 8630 -2505 8750 -2475
rect 8630 -2535 8675 -2505
rect 8705 -2535 8750 -2505
rect 8630 -2570 8750 -2535
rect 8630 -2600 8675 -2570
rect 8705 -2600 8750 -2570
rect 8630 -2640 8750 -2600
rect 8630 -2670 8675 -2640
rect 8705 -2670 8750 -2640
rect 8630 -2710 8750 -2670
rect 8630 -2740 8675 -2710
rect 8705 -2740 8750 -2710
rect 8630 -2780 8750 -2740
rect 8630 -2810 8675 -2780
rect 8705 -2810 8750 -2780
rect 8630 -2845 8750 -2810
rect 8630 -2875 8675 -2845
rect 8705 -2875 8750 -2845
rect 8630 -2890 8750 -2875
rect 8980 -1305 9100 -1290
rect 8980 -1335 9025 -1305
rect 9055 -1335 9100 -1305
rect 8980 -1370 9100 -1335
rect 8980 -1400 9025 -1370
rect 9055 -1400 9100 -1370
rect 8980 -1440 9100 -1400
rect 8980 -1470 9025 -1440
rect 9055 -1470 9100 -1440
rect 8980 -1510 9100 -1470
rect 8980 -1540 9025 -1510
rect 9055 -1540 9100 -1510
rect 8980 -1580 9100 -1540
rect 8980 -1610 9025 -1580
rect 9055 -1610 9100 -1580
rect 8980 -1645 9100 -1610
rect 8980 -1675 9025 -1645
rect 9055 -1675 9100 -1645
rect 8980 -1705 9100 -1675
rect 8980 -1735 9025 -1705
rect 9055 -1735 9100 -1705
rect 8980 -1770 9100 -1735
rect 8980 -1800 9025 -1770
rect 9055 -1800 9100 -1770
rect 8980 -1840 9100 -1800
rect 8980 -1870 9025 -1840
rect 9055 -1870 9100 -1840
rect 8980 -1910 9100 -1870
rect 8980 -1940 9025 -1910
rect 9055 -1940 9100 -1910
rect 8980 -1980 9100 -1940
rect 8980 -2010 9025 -1980
rect 9055 -2010 9100 -1980
rect 8980 -2045 9100 -2010
rect 8980 -2075 9025 -2045
rect 9055 -2075 9100 -2045
rect 8980 -2105 9100 -2075
rect 8980 -2135 9025 -2105
rect 9055 -2135 9100 -2105
rect 8980 -2170 9100 -2135
rect 8980 -2200 9025 -2170
rect 9055 -2200 9100 -2170
rect 8980 -2240 9100 -2200
rect 8980 -2270 9025 -2240
rect 9055 -2270 9100 -2240
rect 8980 -2310 9100 -2270
rect 8980 -2340 9025 -2310
rect 9055 -2340 9100 -2310
rect 8980 -2380 9100 -2340
rect 8980 -2410 9025 -2380
rect 9055 -2410 9100 -2380
rect 8980 -2445 9100 -2410
rect 8980 -2475 9025 -2445
rect 9055 -2475 9100 -2445
rect 8980 -2505 9100 -2475
rect 8980 -2535 9025 -2505
rect 9055 -2535 9100 -2505
rect 8980 -2570 9100 -2535
rect 8980 -2600 9025 -2570
rect 9055 -2600 9100 -2570
rect 8980 -2640 9100 -2600
rect 8980 -2670 9025 -2640
rect 9055 -2670 9100 -2640
rect 8980 -2710 9100 -2670
rect 8980 -2740 9025 -2710
rect 9055 -2740 9100 -2710
rect 8980 -2780 9100 -2740
rect 8980 -2810 9025 -2780
rect 9055 -2810 9100 -2780
rect 8980 -2845 9100 -2810
rect 8980 -2875 9025 -2845
rect 9055 -2875 9100 -2845
rect 8980 -2890 9100 -2875
<< via1 >>
rect 2115 19280 2145 19310
rect 2115 19215 2145 19245
rect 2115 19145 2145 19175
rect 2115 19075 2145 19105
rect 2115 19005 2145 19035
rect 2115 18940 2145 18970
rect 2115 18880 2145 18910
rect 2115 18815 2145 18845
rect 2115 18745 2145 18775
rect 2115 18675 2145 18705
rect 2115 18605 2145 18635
rect 2115 18540 2145 18570
rect 2115 18480 2145 18510
rect 2115 18415 2145 18445
rect 2115 18345 2145 18375
rect 2115 18275 2145 18305
rect 2115 18205 2145 18235
rect 2115 18140 2145 18170
rect 2115 18080 2145 18110
rect 2115 18015 2145 18045
rect 2115 17945 2145 17975
rect 2115 17875 2145 17905
rect 2115 17805 2145 17835
rect 2115 17740 2145 17770
rect 6705 19280 6735 19310
rect 6705 19215 6735 19245
rect 6705 19145 6735 19175
rect 6705 19075 6735 19105
rect 6705 19005 6735 19035
rect 6705 18940 6735 18970
rect 6705 18880 6735 18910
rect 6705 18815 6735 18845
rect 6705 18745 6735 18775
rect 6705 18675 6735 18705
rect 6705 18605 6735 18635
rect 6705 18540 6735 18570
rect 6705 18480 6735 18510
rect 6705 18415 6735 18445
rect 6705 18345 6735 18375
rect 6705 18275 6735 18305
rect 6705 18205 6735 18235
rect 6705 18140 6735 18170
rect 6705 18080 6735 18110
rect 6705 18015 6735 18045
rect 6705 17945 6735 17975
rect 6705 17875 6735 17905
rect 6705 17805 6735 17835
rect 6705 17740 6735 17770
rect 2075 15660 2105 15690
rect 2115 15660 2145 15690
rect 2155 15660 2185 15690
rect 2075 15620 2105 15650
rect 2115 15620 2145 15650
rect 2155 15620 2185 15650
rect 2075 15580 2105 15610
rect 2115 15580 2145 15610
rect 2155 15580 2185 15610
rect 2075 12680 2105 12710
rect 2115 12680 2145 12710
rect 2155 12680 2185 12710
rect 2075 12640 2105 12670
rect 2115 12640 2145 12670
rect 2155 12640 2185 12670
rect 2075 12520 2105 12550
rect 2115 12520 2145 12550
rect 2155 12520 2185 12550
rect 2075 12480 2105 12510
rect 2115 12480 2145 12510
rect 2155 12480 2185 12510
rect 2075 12440 2105 12470
rect 2115 12440 2145 12470
rect 2155 12440 2185 12470
rect 2210 15895 2240 15925
rect 2250 15895 2280 15925
rect 2290 15895 2320 15925
rect -75 9605 -45 9635
rect -75 9540 -45 9570
rect -75 9470 -45 9500
rect -75 9400 -45 9430
rect -75 9330 -45 9360
rect -75 9265 -45 9295
rect -75 9205 -45 9235
rect -75 9140 -45 9170
rect -75 9070 -45 9100
rect -75 9000 -45 9030
rect -75 8930 -45 8960
rect -75 8865 -45 8895
rect -75 8805 -45 8835
rect -75 8740 -45 8770
rect -75 8670 -45 8700
rect -75 8600 -45 8630
rect -75 8530 -45 8560
rect -75 8465 -45 8495
rect -75 8405 -45 8435
rect -75 8340 -45 8370
rect -75 8270 -45 8300
rect -75 8200 -45 8230
rect -75 8130 -45 8160
rect -75 8065 -45 8095
rect -75 8005 -45 8035
rect -75 7940 -45 7970
rect -75 7870 -45 7900
rect -75 7800 -45 7830
rect -75 7730 -45 7760
rect -75 7665 -45 7695
rect -75 7605 -45 7635
rect -75 7540 -45 7570
rect -75 7470 -45 7500
rect -75 7400 -45 7430
rect -75 7330 -45 7360
rect -75 7265 -45 7295
rect -75 7205 -45 7235
rect -75 7140 -45 7170
rect -75 7070 -45 7100
rect -75 7000 -45 7030
rect -75 6930 -45 6960
rect -75 6865 -45 6895
rect -75 6805 -45 6835
rect -75 6740 -45 6770
rect -75 6670 -45 6700
rect -75 6600 -45 6630
rect -75 6530 -45 6560
rect -75 6465 -45 6495
rect 275 9605 305 9635
rect 275 9540 305 9570
rect 275 9470 305 9500
rect 275 9400 305 9430
rect 275 9330 305 9360
rect 275 9265 305 9295
rect 275 9205 305 9235
rect 275 9140 305 9170
rect 275 9070 305 9100
rect 275 9000 305 9030
rect 275 8930 305 8960
rect 275 8865 305 8895
rect 275 8805 305 8835
rect 275 8740 305 8770
rect 275 8670 305 8700
rect 275 8600 305 8630
rect 275 8530 305 8560
rect 275 8465 305 8495
rect 275 8405 305 8435
rect 275 8340 305 8370
rect 275 8270 305 8300
rect 275 8200 305 8230
rect 275 8130 305 8160
rect 275 8065 305 8095
rect 275 8005 305 8035
rect 275 7940 305 7970
rect 275 7870 305 7900
rect 275 7800 305 7830
rect 275 7730 305 7760
rect 275 7665 305 7695
rect 275 7605 305 7635
rect 275 7540 305 7570
rect 275 7470 305 7500
rect 275 7400 305 7430
rect 275 7330 305 7360
rect 275 7265 305 7295
rect 275 7205 305 7235
rect 275 7140 305 7170
rect 275 7070 305 7100
rect 275 7000 305 7030
rect 275 6930 305 6960
rect 275 6865 305 6895
rect 275 6805 305 6835
rect 275 6740 305 6770
rect 275 6670 305 6700
rect 275 6600 305 6630
rect 275 6530 305 6560
rect 275 6465 305 6495
rect 625 9605 655 9635
rect 625 9540 655 9570
rect 625 9470 655 9500
rect 625 9400 655 9430
rect 625 9330 655 9360
rect 625 9265 655 9295
rect 625 9205 655 9235
rect 625 9140 655 9170
rect 625 9070 655 9100
rect 625 9000 655 9030
rect 625 8930 655 8960
rect 625 8865 655 8895
rect 625 8805 655 8835
rect 625 8740 655 8770
rect 625 8670 655 8700
rect 625 8600 655 8630
rect 625 8530 655 8560
rect 625 8465 655 8495
rect 625 8405 655 8435
rect 625 8340 655 8370
rect 625 8270 655 8300
rect 625 8200 655 8230
rect 625 8130 655 8160
rect 625 8065 655 8095
rect 625 8005 655 8035
rect 625 7940 655 7970
rect 625 7870 655 7900
rect 625 7800 655 7830
rect 625 7730 655 7760
rect 625 7665 655 7695
rect 625 7605 655 7635
rect 625 7540 655 7570
rect 625 7470 655 7500
rect 625 7400 655 7430
rect 625 7330 655 7360
rect 625 7265 655 7295
rect 625 7205 655 7235
rect 625 7140 655 7170
rect 625 7070 655 7100
rect 625 7000 655 7030
rect 625 6930 655 6960
rect 625 6865 655 6895
rect 625 6805 655 6835
rect 625 6740 655 6770
rect 625 6670 655 6700
rect 625 6600 655 6630
rect 625 6530 655 6560
rect 625 6465 655 6495
rect 975 9605 1005 9635
rect 975 9540 1005 9570
rect 975 9470 1005 9500
rect 975 9400 1005 9430
rect 975 9330 1005 9360
rect 975 9265 1005 9295
rect 975 9205 1005 9235
rect 975 9140 1005 9170
rect 975 9070 1005 9100
rect 975 9000 1005 9030
rect 975 8930 1005 8960
rect 975 8865 1005 8895
rect 975 8805 1005 8835
rect 975 8740 1005 8770
rect 975 8670 1005 8700
rect 975 8600 1005 8630
rect 975 8530 1005 8560
rect 975 8465 1005 8495
rect 975 8405 1005 8435
rect 975 8340 1005 8370
rect 975 8270 1005 8300
rect 975 8200 1005 8230
rect 975 8130 1005 8160
rect 975 8065 1005 8095
rect 975 8005 1005 8035
rect 975 7940 1005 7970
rect 975 7870 1005 7900
rect 975 7800 1005 7830
rect 975 7730 1005 7760
rect 975 7665 1005 7695
rect 975 7605 1005 7635
rect 975 7540 1005 7570
rect 975 7470 1005 7500
rect 975 7400 1005 7430
rect 975 7330 1005 7360
rect 975 7265 1005 7295
rect 975 7205 1005 7235
rect 975 7140 1005 7170
rect 975 7070 1005 7100
rect 975 7000 1005 7030
rect 975 6930 1005 6960
rect 975 6865 1005 6895
rect 975 6805 1005 6835
rect 975 6740 1005 6770
rect 975 6670 1005 6700
rect 975 6600 1005 6630
rect 975 6530 1005 6560
rect 975 6465 1005 6495
rect 1675 9605 1705 9635
rect 1675 9540 1705 9570
rect 1675 9470 1705 9500
rect 1675 9400 1705 9430
rect 1675 9330 1705 9360
rect 1675 9265 1705 9295
rect 1675 9205 1705 9235
rect 1675 9140 1705 9170
rect 1675 9070 1705 9100
rect 1675 9000 1705 9030
rect 1675 8930 1705 8960
rect 1675 8865 1705 8895
rect 1675 8805 1705 8835
rect 1675 8740 1705 8770
rect 1675 8670 1705 8700
rect 1675 8600 1705 8630
rect 1675 8530 1705 8560
rect 1675 8465 1705 8495
rect 1675 8405 1705 8435
rect 1675 8340 1705 8370
rect 1675 8270 1705 8300
rect 1675 8200 1705 8230
rect 1675 8130 1705 8160
rect 1675 8065 1705 8095
rect 1675 8005 1705 8035
rect 1675 7940 1705 7970
rect 1675 7870 1705 7900
rect 1675 7800 1705 7830
rect 1675 7730 1705 7760
rect 1675 7665 1705 7695
rect 1675 7605 1705 7635
rect 1675 7540 1705 7570
rect 1675 7470 1705 7500
rect 1675 7400 1705 7430
rect 1675 7330 1705 7360
rect 1675 7265 1705 7295
rect 1675 7205 1705 7235
rect 1675 7140 1705 7170
rect 1675 7070 1705 7100
rect 1675 7000 1705 7030
rect 1675 6930 1705 6960
rect 1675 6865 1705 6895
rect 1675 6805 1705 6835
rect 1675 6740 1705 6770
rect 1675 6670 1705 6700
rect 1675 6600 1705 6630
rect 1675 6530 1705 6560
rect 1675 6465 1705 6495
rect 6665 15565 6695 15595
rect 6705 15565 6735 15595
rect 6745 15565 6775 15595
rect 6665 15525 6695 15555
rect 6705 15525 6735 15555
rect 6745 15525 6775 15555
rect 6665 15485 6695 15515
rect 6705 15485 6735 15515
rect 6745 15485 6775 15515
rect 6665 12895 6695 12925
rect 6705 12895 6735 12925
rect 6745 12895 6775 12925
rect 6665 12855 6695 12885
rect 6705 12855 6735 12885
rect 6745 12855 6775 12885
rect 6665 12815 6695 12845
rect 6705 12815 6735 12845
rect 6745 12815 6775 12845
rect 6665 12120 6695 12150
rect 6705 12120 6735 12150
rect 6745 12120 6775 12150
rect 6665 12080 6695 12110
rect 6705 12080 6735 12110
rect 6745 12080 6775 12110
rect 6665 12040 6695 12070
rect 6705 12040 6735 12070
rect 6745 12040 6775 12070
rect 6665 11135 6695 11165
rect 6705 11135 6735 11165
rect 6745 11135 6775 11165
rect 6665 11095 6695 11125
rect 6705 11095 6735 11125
rect 6745 11095 6775 11125
rect 6665 11055 6695 11085
rect 6705 11055 6735 11085
rect 6745 11055 6775 11085
rect 6665 10410 6695 10440
rect 6705 10410 6735 10440
rect 6745 10410 6775 10440
rect 6665 10370 6695 10400
rect 6705 10370 6735 10400
rect 6745 10370 6775 10400
rect 6665 10330 6695 10360
rect 6705 10330 6735 10360
rect 6745 10330 6775 10360
rect 2250 9605 2280 9635
rect 2250 9540 2280 9570
rect 2250 9470 2280 9500
rect 2250 9400 2280 9430
rect 2250 9330 2280 9360
rect 2250 9265 2280 9295
rect 2250 9205 2280 9235
rect 2250 9140 2280 9170
rect 2250 9070 2280 9100
rect 2250 9000 2280 9030
rect 2250 8930 2280 8960
rect 2250 8865 2280 8895
rect 2250 8805 2280 8835
rect 2250 8740 2280 8770
rect 2250 8670 2280 8700
rect 2250 8600 2280 8630
rect 2250 8530 2280 8560
rect 2250 8465 2280 8495
rect 2250 8405 2280 8435
rect 2250 8340 2280 8370
rect 2250 8270 2280 8300
rect 2250 8200 2280 8230
rect 2250 8130 2280 8160
rect 2250 8065 2280 8095
rect 2250 8005 2280 8035
rect 2250 7940 2280 7970
rect 2250 7870 2280 7900
rect 2250 7800 2280 7830
rect 2250 7730 2280 7760
rect 2250 7665 2280 7695
rect 2250 7605 2280 7635
rect 2250 7540 2280 7570
rect 2250 7470 2280 7500
rect 2250 7400 2280 7430
rect 2250 7330 2280 7360
rect 2250 7265 2280 7295
rect 2250 7205 2280 7235
rect 2250 7140 2280 7170
rect 2250 7070 2280 7100
rect 2250 7000 2280 7030
rect 2250 6930 2280 6960
rect 2250 6865 2280 6895
rect 2250 6805 2280 6835
rect 2250 6740 2280 6770
rect 2250 6670 2280 6700
rect 2250 6600 2280 6630
rect 2250 6530 2280 6560
rect 2250 6465 2280 6495
rect 2050 6400 2080 6430
rect 2480 6400 2510 6430
rect 2005 6345 2035 6375
rect 1285 6175 1315 6205
rect 1325 6175 1355 6205
rect 1365 6175 1395 6205
rect 1285 6135 1315 6165
rect 1325 6135 1355 6165
rect 1365 6135 1395 6165
rect 1285 6095 1315 6125
rect 1325 6095 1355 6125
rect 1365 6095 1395 6125
rect 3180 9605 3210 9635
rect 3240 9605 3270 9635
rect 3180 9540 3210 9570
rect 3240 9540 3270 9570
rect 3180 9470 3210 9500
rect 3240 9470 3270 9500
rect 3180 9400 3210 9430
rect 3240 9400 3270 9430
rect 3180 9330 3210 9360
rect 3240 9330 3270 9360
rect 3180 9265 3210 9295
rect 3240 9265 3270 9295
rect 3180 9205 3210 9235
rect 3240 9205 3270 9235
rect 3180 9140 3210 9170
rect 3240 9140 3270 9170
rect 3180 9070 3210 9100
rect 3240 9070 3270 9100
rect 3180 9000 3210 9030
rect 3240 9000 3270 9030
rect 3180 8930 3210 8960
rect 3240 8930 3270 8960
rect 3180 8865 3210 8895
rect 3240 8865 3270 8895
rect 3180 8805 3210 8835
rect 3240 8805 3270 8835
rect 3180 8740 3210 8770
rect 3240 8740 3270 8770
rect 3180 8670 3210 8700
rect 3240 8670 3270 8700
rect 3180 8600 3210 8630
rect 3240 8600 3270 8630
rect 3180 8530 3210 8560
rect 3240 8530 3270 8560
rect 3180 8465 3210 8495
rect 3240 8465 3270 8495
rect 3180 8405 3210 8435
rect 3240 8405 3270 8435
rect 3180 8340 3210 8370
rect 3240 8340 3270 8370
rect 3180 8270 3210 8300
rect 3240 8270 3270 8300
rect 3180 8200 3210 8230
rect 3240 8200 3270 8230
rect 3180 8130 3210 8160
rect 3240 8130 3270 8160
rect 3180 8065 3210 8095
rect 3240 8065 3270 8095
rect 3180 8005 3210 8035
rect 3240 8005 3270 8035
rect 3180 7940 3210 7970
rect 3240 7940 3270 7970
rect 3180 7870 3210 7900
rect 3240 7870 3270 7900
rect 3180 7800 3210 7830
rect 3240 7800 3270 7830
rect 3180 7730 3210 7760
rect 3240 7730 3270 7760
rect 3180 7665 3210 7695
rect 3240 7665 3270 7695
rect 3180 7605 3210 7635
rect 3240 7605 3270 7635
rect 3180 7540 3210 7570
rect 3240 7540 3270 7570
rect 3180 7470 3210 7500
rect 3240 7470 3270 7500
rect 3180 7400 3210 7430
rect 3240 7400 3270 7430
rect 3180 7330 3210 7360
rect 3240 7330 3270 7360
rect 3180 7265 3210 7295
rect 3240 7265 3270 7295
rect 3180 7205 3210 7235
rect 3240 7205 3270 7235
rect 3180 7140 3210 7170
rect 3240 7140 3270 7170
rect 3180 7070 3210 7100
rect 3240 7070 3270 7100
rect 3180 7000 3210 7030
rect 3240 7000 3270 7030
rect 3180 6930 3210 6960
rect 3240 6930 3270 6960
rect 3180 6865 3210 6895
rect 3240 6865 3270 6895
rect 3180 6805 3210 6835
rect 3240 6805 3270 6835
rect 3180 6740 3210 6770
rect 3240 6740 3270 6770
rect 3180 6670 3210 6700
rect 3240 6670 3270 6700
rect 3180 6600 3210 6630
rect 3240 6600 3270 6630
rect 3180 6530 3210 6560
rect 3240 6530 3270 6560
rect 3180 6465 3210 6495
rect 3240 6465 3270 6495
rect 2850 6400 2880 6430
rect 2720 6300 2750 6330
rect 3080 6300 3110 6330
rect 6665 10050 6695 10080
rect 6705 10050 6735 10080
rect 6745 10050 6775 10080
rect 6665 10010 6695 10040
rect 6705 10010 6735 10040
rect 6745 10010 6775 10040
rect 6665 9970 6695 10000
rect 6705 9970 6735 10000
rect 6745 9970 6775 10000
rect 3350 9605 3380 9635
rect 3350 9540 3380 9570
rect 3350 9470 3380 9500
rect 3350 9400 3380 9430
rect 3350 9330 3380 9360
rect 3350 9265 3380 9295
rect 3350 9205 3380 9235
rect 3350 9140 3380 9170
rect 3350 9070 3380 9100
rect 3350 9000 3380 9030
rect 3350 8930 3380 8960
rect 3350 8865 3380 8895
rect 3350 8805 3380 8835
rect 3350 8740 3380 8770
rect 3350 8670 3380 8700
rect 3350 8600 3380 8630
rect 3350 8530 3380 8560
rect 3350 8465 3380 8495
rect 3350 8405 3380 8435
rect 3350 8340 3380 8370
rect 3350 8270 3380 8300
rect 3350 8200 3380 8230
rect 3350 8130 3380 8160
rect 3350 8065 3380 8095
rect 3350 8005 3380 8035
rect 3350 7940 3380 7970
rect 3350 7870 3380 7900
rect 3350 7800 3380 7830
rect 3350 7730 3380 7760
rect 3350 7665 3380 7695
rect 3350 7605 3380 7635
rect 3350 7540 3380 7570
rect 3350 7470 3380 7500
rect 3350 7400 3380 7430
rect 3350 7330 3380 7360
rect 3350 7265 3380 7295
rect 3350 7205 3380 7235
rect 3350 7140 3380 7170
rect 3350 7070 3380 7100
rect 3350 7000 3380 7030
rect 3350 6930 3380 6960
rect 3350 6865 3380 6895
rect 3350 6805 3380 6835
rect 3350 6740 3380 6770
rect 3350 6670 3380 6700
rect 3350 6600 3380 6630
rect 3350 6530 3380 6560
rect 3350 6465 3380 6495
rect 3385 6400 3415 6430
rect 3295 6285 3325 6315
rect 3080 5060 3110 5090
rect 3635 6345 3665 6375
rect 3440 6230 3470 6260
rect 3385 3775 3415 3805
rect 4310 6175 4340 6205
rect 4310 6135 4340 6165
rect 4310 6095 4340 6125
rect 4475 6285 4505 6315
rect 4475 6230 4505 6260
rect 4420 6175 4450 6205
rect 4420 6135 4450 6165
rect 4420 6095 4450 6125
rect 4530 6175 4560 6205
rect 4530 6135 4560 6165
rect 4530 6095 4560 6125
rect 5475 6400 5505 6430
rect 6150 6400 6180 6430
rect 5315 6345 5345 6375
rect 4640 6175 4670 6205
rect 4640 6135 4670 6165
rect 4640 6095 4670 6125
rect 5525 6230 5555 6260
rect 5475 3835 5505 3865
rect 3440 3095 3470 3125
rect 4475 3095 4505 3125
rect 6705 9540 6735 9570
rect 6705 9470 6735 9500
rect 6705 9400 6735 9430
rect 6705 9330 6735 9360
rect 6705 9265 6735 9295
rect 6705 9205 6735 9235
rect 6705 9140 6735 9170
rect 6705 9070 6735 9100
rect 6705 9000 6735 9030
rect 6705 8930 6735 8960
rect 6705 8865 6735 8895
rect 6705 8805 6735 8835
rect 6705 8740 6735 8770
rect 6705 8670 6735 8700
rect 6705 8600 6735 8630
rect 6705 8530 6735 8560
rect 6705 8465 6735 8495
rect 6705 8405 6735 8435
rect 6705 8340 6735 8370
rect 6705 8270 6735 8300
rect 6705 8200 6735 8230
rect 6705 8130 6735 8160
rect 6705 8065 6735 8095
rect 6705 8005 6735 8035
rect 6705 7940 6735 7970
rect 6705 7870 6735 7900
rect 6705 7800 6735 7830
rect 6705 7730 6735 7760
rect 6705 7665 6735 7695
rect 6705 7605 6735 7635
rect 6705 7540 6735 7570
rect 6705 7470 6735 7500
rect 6705 7400 6735 7430
rect 6705 7330 6735 7360
rect 6705 7265 6735 7295
rect 6705 7205 6735 7235
rect 6705 7140 6735 7170
rect 6705 7070 6735 7100
rect 6705 7000 6735 7030
rect 6705 6930 6735 6960
rect 6705 6865 6735 6895
rect 6705 6805 6735 6835
rect 6705 6740 6735 6770
rect 6705 6670 6735 6700
rect 6705 6600 6735 6630
rect 6705 6530 6735 6560
rect 6705 6465 6735 6495
rect 7275 9605 7305 9635
rect 7275 9540 7305 9570
rect 7275 9470 7305 9500
rect 7275 9400 7305 9430
rect 7275 9330 7305 9360
rect 7275 9265 7305 9295
rect 7275 9205 7305 9235
rect 7275 9140 7305 9170
rect 7275 9070 7305 9100
rect 7275 9000 7305 9030
rect 7275 8930 7305 8960
rect 7275 8865 7305 8895
rect 7275 8805 7305 8835
rect 7275 8740 7305 8770
rect 7275 8670 7305 8700
rect 7275 8600 7305 8630
rect 7275 8530 7305 8560
rect 7275 8465 7305 8495
rect 7275 8405 7305 8435
rect 7275 8340 7305 8370
rect 7275 8270 7305 8300
rect 7275 8200 7305 8230
rect 7275 8130 7305 8160
rect 7275 8065 7305 8095
rect 7275 8005 7305 8035
rect 7275 7940 7305 7970
rect 7275 7870 7305 7900
rect 7275 7800 7305 7830
rect 7275 7730 7305 7760
rect 7275 7665 7305 7695
rect 7275 7605 7305 7635
rect 7275 7540 7305 7570
rect 7275 7470 7305 7500
rect 7275 7400 7305 7430
rect 7275 7330 7305 7360
rect 7275 7265 7305 7295
rect 7275 7205 7305 7235
rect 7275 7140 7305 7170
rect 7275 7070 7305 7100
rect 7275 7000 7305 7030
rect 7275 6930 7305 6960
rect 7275 6865 7305 6895
rect 7275 6805 7305 6835
rect 7275 6740 7305 6770
rect 7275 6670 7305 6700
rect 7275 6600 7305 6630
rect 7275 6530 7305 6560
rect 7275 6465 7305 6495
rect 6470 6400 6500 6430
rect 6900 6400 6930 6430
rect 5575 5405 5605 5435
rect 6225 5405 6255 5435
rect 5575 4410 5605 4440
rect 5525 3095 5555 3125
rect 4475 2985 4505 3015
rect 6945 6345 6975 6375
rect 2050 2285 2080 2315
rect 2125 2285 2155 2315
rect 6825 2285 6855 2315
rect 6900 2285 6930 2315
rect 2005 2230 2035 2260
rect 2080 2230 2110 2260
rect 7975 9605 8005 9635
rect 7975 9540 8005 9570
rect 7975 9470 8005 9500
rect 7975 9400 8005 9430
rect 7975 9330 8005 9360
rect 7975 9265 8005 9295
rect 7975 9205 8005 9235
rect 7975 9140 8005 9170
rect 7975 9070 8005 9100
rect 7975 9000 8005 9030
rect 7975 8930 8005 8960
rect 7975 8865 8005 8895
rect 7975 8805 8005 8835
rect 7975 8740 8005 8770
rect 7975 8670 8005 8700
rect 7975 8600 8005 8630
rect 7975 8530 8005 8560
rect 7975 8465 8005 8495
rect 7975 8405 8005 8435
rect 7975 8340 8005 8370
rect 7975 8270 8005 8300
rect 7975 8200 8005 8230
rect 7975 8130 8005 8160
rect 7975 8065 8005 8095
rect 7975 8005 8005 8035
rect 7975 7940 8005 7970
rect 7975 7870 8005 7900
rect 7975 7800 8005 7830
rect 7975 7730 8005 7760
rect 7975 7665 8005 7695
rect 7975 7605 8005 7635
rect 7975 7540 8005 7570
rect 7975 7470 8005 7500
rect 7975 7400 8005 7430
rect 7975 7330 8005 7360
rect 7975 7265 8005 7295
rect 7975 7205 8005 7235
rect 7975 7140 8005 7170
rect 7975 7070 8005 7100
rect 7975 7000 8005 7030
rect 7975 6930 8005 6960
rect 7975 6865 8005 6895
rect 7975 6805 8005 6835
rect 7975 6740 8005 6770
rect 7975 6670 8005 6700
rect 7975 6600 8005 6630
rect 7975 6530 8005 6560
rect 7975 6465 8005 6495
rect 7585 6175 7615 6205
rect 7625 6175 7655 6205
rect 7665 6175 7695 6205
rect 8325 9605 8355 9635
rect 8325 9540 8355 9570
rect 8325 9470 8355 9500
rect 8325 9400 8355 9430
rect 8325 9330 8355 9360
rect 8325 9265 8355 9295
rect 8325 9205 8355 9235
rect 8325 9140 8355 9170
rect 8325 9070 8355 9100
rect 8325 9000 8355 9030
rect 8325 8930 8355 8960
rect 8325 8865 8355 8895
rect 8325 8805 8355 8835
rect 8325 8740 8355 8770
rect 8325 8670 8355 8700
rect 8325 8600 8355 8630
rect 8325 8530 8355 8560
rect 8325 8465 8355 8495
rect 8325 8405 8355 8435
rect 8325 8340 8355 8370
rect 8325 8270 8355 8300
rect 8325 8200 8355 8230
rect 8325 8130 8355 8160
rect 8325 8065 8355 8095
rect 8325 8005 8355 8035
rect 8325 7940 8355 7970
rect 8325 7870 8355 7900
rect 8325 7800 8355 7830
rect 8325 7730 8355 7760
rect 8325 7665 8355 7695
rect 8325 7605 8355 7635
rect 8325 7540 8355 7570
rect 8325 7470 8355 7500
rect 8325 7400 8355 7430
rect 8325 7330 8355 7360
rect 8325 7265 8355 7295
rect 8325 7205 8355 7235
rect 8325 7140 8355 7170
rect 8325 7070 8355 7100
rect 8325 7000 8355 7030
rect 8325 6930 8355 6960
rect 8325 6865 8355 6895
rect 8325 6805 8355 6835
rect 8325 6740 8355 6770
rect 8325 6670 8355 6700
rect 8325 6600 8355 6630
rect 8325 6530 8355 6560
rect 8325 6465 8355 6495
rect 8675 9605 8705 9635
rect 8675 9540 8705 9570
rect 8675 9470 8705 9500
rect 8675 9400 8705 9430
rect 8675 9330 8705 9360
rect 8675 9265 8705 9295
rect 8675 9205 8705 9235
rect 8675 9140 8705 9170
rect 8675 9070 8705 9100
rect 8675 9000 8705 9030
rect 8675 8930 8705 8960
rect 8675 8865 8705 8895
rect 8675 8805 8705 8835
rect 8675 8740 8705 8770
rect 8675 8670 8705 8700
rect 8675 8600 8705 8630
rect 8675 8530 8705 8560
rect 8675 8465 8705 8495
rect 8675 8405 8705 8435
rect 8675 8340 8705 8370
rect 8675 8270 8705 8300
rect 8675 8200 8705 8230
rect 8675 8130 8705 8160
rect 8675 8065 8705 8095
rect 8675 8005 8705 8035
rect 8675 7940 8705 7970
rect 8675 7870 8705 7900
rect 8675 7800 8705 7830
rect 8675 7730 8705 7760
rect 8675 7665 8705 7695
rect 8675 7605 8705 7635
rect 8675 7540 8705 7570
rect 8675 7470 8705 7500
rect 8675 7400 8705 7430
rect 8675 7330 8705 7360
rect 8675 7265 8705 7295
rect 8675 7205 8705 7235
rect 8675 7140 8705 7170
rect 8675 7070 8705 7100
rect 8675 7000 8705 7030
rect 8675 6930 8705 6960
rect 8675 6865 8705 6895
rect 8675 6805 8705 6835
rect 8675 6740 8705 6770
rect 8675 6670 8705 6700
rect 8675 6600 8705 6630
rect 8675 6530 8705 6560
rect 8675 6465 8705 6495
rect 9025 9605 9055 9635
rect 9025 9540 9055 9570
rect 9025 9470 9055 9500
rect 9025 9400 9055 9430
rect 9025 9330 9055 9360
rect 9025 9265 9055 9295
rect 9025 9205 9055 9235
rect 9025 9140 9055 9170
rect 9025 9070 9055 9100
rect 9025 9000 9055 9030
rect 9025 8930 9055 8960
rect 9025 8865 9055 8895
rect 9025 8805 9055 8835
rect 9025 8740 9055 8770
rect 9025 8670 9055 8700
rect 9025 8600 9055 8630
rect 9025 8530 9055 8560
rect 9025 8465 9055 8495
rect 9025 8405 9055 8435
rect 9025 8340 9055 8370
rect 9025 8270 9055 8300
rect 9025 8200 9055 8230
rect 9025 8130 9055 8160
rect 9025 8065 9055 8095
rect 9025 8005 9055 8035
rect 9025 7940 9055 7970
rect 9025 7870 9055 7900
rect 9025 7800 9055 7830
rect 9025 7730 9055 7760
rect 9025 7665 9055 7695
rect 9025 7605 9055 7635
rect 9025 7540 9055 7570
rect 9025 7470 9055 7500
rect 9025 7400 9055 7430
rect 9025 7330 9055 7360
rect 9025 7265 9055 7295
rect 9025 7205 9055 7235
rect 9025 7140 9055 7170
rect 9025 7070 9055 7100
rect 9025 7000 9055 7030
rect 9025 6930 9055 6960
rect 9025 6865 9055 6895
rect 9025 6805 9055 6835
rect 9025 6740 9055 6770
rect 9025 6670 9055 6700
rect 9025 6600 9055 6630
rect 9025 6530 9055 6560
rect 9025 6465 9055 6495
rect 7585 6135 7615 6165
rect 7625 6135 7655 6165
rect 7665 6135 7695 6165
rect 7585 6095 7615 6125
rect 7625 6095 7655 6125
rect 7665 6095 7695 6125
rect 6870 2230 6900 2260
rect 6945 2230 6975 2260
rect 1285 1130 1315 1160
rect 1325 1130 1355 1160
rect 1365 1130 1395 1160
rect 1285 1090 1315 1120
rect 1325 1090 1355 1120
rect 1365 1090 1395 1120
rect 1285 1050 1315 1080
rect 1325 1050 1355 1080
rect 1365 1050 1395 1080
rect 4420 1130 4450 1160
rect 4420 1090 4450 1120
rect 4420 1050 4450 1080
rect 4530 1130 4560 1160
rect 4530 1090 4560 1120
rect 4530 1050 4560 1080
rect 7585 1130 7615 1160
rect 7625 1130 7655 1160
rect 7665 1130 7695 1160
rect 7585 1090 7615 1120
rect 7625 1090 7655 1120
rect 7665 1090 7695 1120
rect 7585 1050 7615 1080
rect 7625 1050 7655 1080
rect 7665 1050 7695 1080
rect -75 -1335 -45 -1305
rect -75 -1400 -45 -1370
rect -75 -1470 -45 -1440
rect -75 -1540 -45 -1510
rect -75 -1610 -45 -1580
rect -75 -1675 -45 -1645
rect -75 -1735 -45 -1705
rect -75 -1800 -45 -1770
rect -75 -1870 -45 -1840
rect -75 -1940 -45 -1910
rect -75 -2010 -45 -1980
rect -75 -2075 -45 -2045
rect -75 -2135 -45 -2105
rect -75 -2200 -45 -2170
rect -75 -2270 -45 -2240
rect -75 -2340 -45 -2310
rect -75 -2410 -45 -2380
rect -75 -2475 -45 -2445
rect -75 -2535 -45 -2505
rect -75 -2600 -45 -2570
rect -75 -2670 -45 -2640
rect -75 -2740 -45 -2710
rect -75 -2810 -45 -2780
rect -75 -2875 -45 -2845
rect 275 -1335 305 -1305
rect 275 -1400 305 -1370
rect 275 -1470 305 -1440
rect 275 -1540 305 -1510
rect 275 -1610 305 -1580
rect 275 -1675 305 -1645
rect 275 -1735 305 -1705
rect 275 -1800 305 -1770
rect 275 -1870 305 -1840
rect 275 -1940 305 -1910
rect 275 -2010 305 -1980
rect 275 -2075 305 -2045
rect 275 -2135 305 -2105
rect 275 -2200 305 -2170
rect 275 -2270 305 -2240
rect 275 -2340 305 -2310
rect 275 -2410 305 -2380
rect 275 -2475 305 -2445
rect 275 -2535 305 -2505
rect 275 -2600 305 -2570
rect 275 -2670 305 -2640
rect 275 -2740 305 -2710
rect 275 -2810 305 -2780
rect 275 -2875 305 -2845
rect 625 -1335 655 -1305
rect 625 -1400 655 -1370
rect 625 -1470 655 -1440
rect 625 -1540 655 -1510
rect 625 -1610 655 -1580
rect 625 -1675 655 -1645
rect 625 -1735 655 -1705
rect 625 -1800 655 -1770
rect 625 -1870 655 -1840
rect 625 -1940 655 -1910
rect 625 -2010 655 -1980
rect 625 -2075 655 -2045
rect 625 -2135 655 -2105
rect 625 -2200 655 -2170
rect 625 -2270 655 -2240
rect 625 -2340 655 -2310
rect 625 -2410 655 -2380
rect 625 -2475 655 -2445
rect 625 -2535 655 -2505
rect 625 -2600 655 -2570
rect 625 -2670 655 -2640
rect 625 -2740 655 -2710
rect 625 -2810 655 -2780
rect 625 -2875 655 -2845
rect 975 -1335 1005 -1305
rect 975 -1400 1005 -1370
rect 975 -1470 1005 -1440
rect 975 -1540 1005 -1510
rect 975 -1610 1005 -1580
rect 975 -1675 1005 -1645
rect 975 -1735 1005 -1705
rect 975 -1800 1005 -1770
rect 975 -1870 1005 -1840
rect 975 -1940 1005 -1910
rect 975 -2010 1005 -1980
rect 975 -2075 1005 -2045
rect 975 -2135 1005 -2105
rect 975 -2200 1005 -2170
rect 975 -2270 1005 -2240
rect 975 -2340 1005 -2310
rect 975 -2410 1005 -2380
rect 975 -2475 1005 -2445
rect 975 -2535 1005 -2505
rect 975 -2600 1005 -2570
rect 975 -2670 1005 -2640
rect 975 -2740 1005 -2710
rect 975 -2810 1005 -2780
rect 975 -2875 1005 -2845
rect 1325 -1335 1355 -1305
rect 1325 -1400 1355 -1370
rect 1325 -1470 1355 -1440
rect 1325 -1540 1355 -1510
rect 1325 -1610 1355 -1580
rect 1325 -1675 1355 -1645
rect 1325 -1735 1355 -1705
rect 1325 -1800 1355 -1770
rect 1325 -1870 1355 -1840
rect 1325 -1940 1355 -1910
rect 1325 -2010 1355 -1980
rect 1325 -2075 1355 -2045
rect 1325 -2135 1355 -2105
rect 1325 -2200 1355 -2170
rect 1325 -2270 1355 -2240
rect 1325 -2340 1355 -2310
rect 1325 -2410 1355 -2380
rect 1325 -2475 1355 -2445
rect 1325 -2535 1355 -2505
rect 1325 -2600 1355 -2570
rect 1325 -2670 1355 -2640
rect 1325 -2740 1355 -2710
rect 1325 -2810 1355 -2780
rect 1325 -2875 1355 -2845
rect 1675 -1335 1705 -1305
rect 1675 -1400 1705 -1370
rect 1675 -1470 1705 -1440
rect 1675 -1540 1705 -1510
rect 1675 -1610 1705 -1580
rect 1675 -1675 1705 -1645
rect 1675 -1735 1705 -1705
rect 1675 -1800 1705 -1770
rect 1675 -1870 1705 -1840
rect 1675 -1940 1705 -1910
rect 1675 -2010 1705 -1980
rect 1675 -2075 1705 -2045
rect 1675 -2135 1705 -2105
rect 1675 -2200 1705 -2170
rect 1675 -2270 1705 -2240
rect 1675 -2340 1705 -2310
rect 1675 -2410 1705 -2380
rect 1675 -2475 1705 -2445
rect 1675 -2535 1705 -2505
rect 1675 -2600 1705 -2570
rect 1675 -2670 1705 -2640
rect 1675 -2740 1705 -2710
rect 1675 -2810 1705 -2780
rect 1675 -2875 1705 -2845
rect 2025 -1335 2055 -1305
rect 2025 -1400 2055 -1370
rect 2025 -1470 2055 -1440
rect 2025 -1540 2055 -1510
rect 2025 -1610 2055 -1580
rect 2025 -1675 2055 -1645
rect 2025 -1735 2055 -1705
rect 2025 -1800 2055 -1770
rect 2025 -1870 2055 -1840
rect 2025 -1940 2055 -1910
rect 2025 -2010 2055 -1980
rect 2025 -2075 2055 -2045
rect 2025 -2135 2055 -2105
rect 2025 -2200 2055 -2170
rect 2025 -2270 2055 -2240
rect 2025 -2340 2055 -2310
rect 2025 -2410 2055 -2380
rect 2025 -2475 2055 -2445
rect 2025 -2535 2055 -2505
rect 2025 -2600 2055 -2570
rect 2025 -2670 2055 -2640
rect 2025 -2740 2055 -2710
rect 2025 -2810 2055 -2780
rect 2025 -2875 2055 -2845
rect 2375 -1335 2405 -1305
rect 2375 -1400 2405 -1370
rect 2375 -1470 2405 -1440
rect 2375 -1540 2405 -1510
rect 2375 -1610 2405 -1580
rect 2375 -1675 2405 -1645
rect 2375 -1735 2405 -1705
rect 2375 -1800 2405 -1770
rect 2375 -1870 2405 -1840
rect 2375 -1940 2405 -1910
rect 2375 -2010 2405 -1980
rect 2375 -2075 2405 -2045
rect 2375 -2135 2405 -2105
rect 2375 -2200 2405 -2170
rect 2375 -2270 2405 -2240
rect 2375 -2340 2405 -2310
rect 2375 -2410 2405 -2380
rect 2375 -2475 2405 -2445
rect 2375 -2535 2405 -2505
rect 2375 -2600 2405 -2570
rect 2375 -2670 2405 -2640
rect 2375 -2740 2405 -2710
rect 2375 -2810 2405 -2780
rect 2375 -2875 2405 -2845
rect 2725 -1335 2755 -1305
rect 2725 -1400 2755 -1370
rect 2725 -1470 2755 -1440
rect 2725 -1540 2755 -1510
rect 2725 -1610 2755 -1580
rect 2725 -1675 2755 -1645
rect 2725 -1735 2755 -1705
rect 2725 -1800 2755 -1770
rect 2725 -1870 2755 -1840
rect 2725 -1940 2755 -1910
rect 2725 -2010 2755 -1980
rect 2725 -2075 2755 -2045
rect 2725 -2135 2755 -2105
rect 2725 -2200 2755 -2170
rect 2725 -2270 2755 -2240
rect 2725 -2340 2755 -2310
rect 2725 -2410 2755 -2380
rect 2725 -2475 2755 -2445
rect 2725 -2535 2755 -2505
rect 2725 -2600 2755 -2570
rect 2725 -2670 2755 -2640
rect 2725 -2740 2755 -2710
rect 2725 -2810 2755 -2780
rect 2725 -2875 2755 -2845
rect 3075 -1335 3105 -1305
rect 3075 -1400 3105 -1370
rect 3075 -1470 3105 -1440
rect 3075 -1540 3105 -1510
rect 3075 -1610 3105 -1580
rect 3075 -1675 3105 -1645
rect 3075 -1735 3105 -1705
rect 3075 -1800 3105 -1770
rect 3075 -1870 3105 -1840
rect 3075 -1940 3105 -1910
rect 3075 -2010 3105 -1980
rect 3075 -2075 3105 -2045
rect 3075 -2135 3105 -2105
rect 3075 -2200 3105 -2170
rect 3075 -2270 3105 -2240
rect 3075 -2340 3105 -2310
rect 3075 -2410 3105 -2380
rect 3075 -2475 3105 -2445
rect 3075 -2535 3105 -2505
rect 3075 -2600 3105 -2570
rect 3075 -2670 3105 -2640
rect 3075 -2740 3105 -2710
rect 3075 -2810 3105 -2780
rect 3075 -2875 3105 -2845
rect 3425 -1335 3455 -1305
rect 3425 -1400 3455 -1370
rect 3425 -1470 3455 -1440
rect 3425 -1540 3455 -1510
rect 3425 -1610 3455 -1580
rect 3425 -1675 3455 -1645
rect 3425 -1735 3455 -1705
rect 3425 -1800 3455 -1770
rect 3425 -1870 3455 -1840
rect 3425 -1940 3455 -1910
rect 3425 -2010 3455 -1980
rect 3425 -2075 3455 -2045
rect 3425 -2135 3455 -2105
rect 3425 -2200 3455 -2170
rect 3425 -2270 3455 -2240
rect 3425 -2340 3455 -2310
rect 3425 -2410 3455 -2380
rect 3425 -2475 3455 -2445
rect 3425 -2535 3455 -2505
rect 3425 -2600 3455 -2570
rect 3425 -2670 3455 -2640
rect 3425 -2740 3455 -2710
rect 3425 -2810 3455 -2780
rect 3425 -2875 3455 -2845
rect 3775 -1335 3805 -1305
rect 3775 -1400 3805 -1370
rect 3775 -1470 3805 -1440
rect 3775 -1540 3805 -1510
rect 3775 -1610 3805 -1580
rect 3775 -1675 3805 -1645
rect 3775 -1735 3805 -1705
rect 3775 -1800 3805 -1770
rect 3775 -1870 3805 -1840
rect 3775 -1940 3805 -1910
rect 3775 -2010 3805 -1980
rect 3775 -2075 3805 -2045
rect 3775 -2135 3805 -2105
rect 3775 -2200 3805 -2170
rect 3775 -2270 3805 -2240
rect 3775 -2340 3805 -2310
rect 3775 -2410 3805 -2380
rect 3775 -2475 3805 -2445
rect 3775 -2535 3805 -2505
rect 3775 -2600 3805 -2570
rect 3775 -2670 3805 -2640
rect 3775 -2740 3805 -2710
rect 3775 -2810 3805 -2780
rect 3775 -2875 3805 -2845
rect 4125 -1335 4155 -1305
rect 4125 -1400 4155 -1370
rect 4125 -1470 4155 -1440
rect 4125 -1540 4155 -1510
rect 4125 -1610 4155 -1580
rect 4125 -1675 4155 -1645
rect 4125 -1735 4155 -1705
rect 4125 -1800 4155 -1770
rect 4125 -1870 4155 -1840
rect 4125 -1940 4155 -1910
rect 4125 -2010 4155 -1980
rect 4125 -2075 4155 -2045
rect 4125 -2135 4155 -2105
rect 4125 -2200 4155 -2170
rect 4125 -2270 4155 -2240
rect 4125 -2340 4155 -2310
rect 4125 -2410 4155 -2380
rect 4125 -2475 4155 -2445
rect 4125 -2535 4155 -2505
rect 4125 -2600 4155 -2570
rect 4125 -2670 4155 -2640
rect 4125 -2740 4155 -2710
rect 4125 -2810 4155 -2780
rect 4125 -2875 4155 -2845
rect 4475 -1335 4505 -1305
rect 4475 -1400 4505 -1370
rect 4475 -1470 4505 -1440
rect 4475 -1540 4505 -1510
rect 4475 -1610 4505 -1580
rect 4475 -1675 4505 -1645
rect 4475 -1735 4505 -1705
rect 4475 -1800 4505 -1770
rect 4475 -1870 4505 -1840
rect 4475 -1940 4505 -1910
rect 4475 -2010 4505 -1980
rect 4475 -2075 4505 -2045
rect 4475 -2135 4505 -2105
rect 4475 -2200 4505 -2170
rect 4475 -2270 4505 -2240
rect 4475 -2340 4505 -2310
rect 4475 -2410 4505 -2380
rect 4475 -2475 4505 -2445
rect 4475 -2535 4505 -2505
rect 4475 -2600 4505 -2570
rect 4475 -2670 4505 -2640
rect 4475 -2740 4505 -2710
rect 4475 -2810 4505 -2780
rect 4475 -2875 4505 -2845
rect 4825 -1335 4855 -1305
rect 4825 -1400 4855 -1370
rect 4825 -1470 4855 -1440
rect 4825 -1540 4855 -1510
rect 4825 -1610 4855 -1580
rect 4825 -1675 4855 -1645
rect 4825 -1735 4855 -1705
rect 4825 -1800 4855 -1770
rect 4825 -1870 4855 -1840
rect 4825 -1940 4855 -1910
rect 4825 -2010 4855 -1980
rect 4825 -2075 4855 -2045
rect 4825 -2135 4855 -2105
rect 4825 -2200 4855 -2170
rect 4825 -2270 4855 -2240
rect 4825 -2340 4855 -2310
rect 4825 -2410 4855 -2380
rect 4825 -2475 4855 -2445
rect 4825 -2535 4855 -2505
rect 4825 -2600 4855 -2570
rect 4825 -2670 4855 -2640
rect 4825 -2740 4855 -2710
rect 4825 -2810 4855 -2780
rect 4825 -2875 4855 -2845
rect 5175 -1335 5205 -1305
rect 5175 -1400 5205 -1370
rect 5175 -1470 5205 -1440
rect 5175 -1540 5205 -1510
rect 5175 -1610 5205 -1580
rect 5175 -1675 5205 -1645
rect 5175 -1735 5205 -1705
rect 5175 -1800 5205 -1770
rect 5175 -1870 5205 -1840
rect 5175 -1940 5205 -1910
rect 5175 -2010 5205 -1980
rect 5175 -2075 5205 -2045
rect 5175 -2135 5205 -2105
rect 5175 -2200 5205 -2170
rect 5175 -2270 5205 -2240
rect 5175 -2340 5205 -2310
rect 5175 -2410 5205 -2380
rect 5175 -2475 5205 -2445
rect 5175 -2535 5205 -2505
rect 5175 -2600 5205 -2570
rect 5175 -2670 5205 -2640
rect 5175 -2740 5205 -2710
rect 5175 -2810 5205 -2780
rect 5175 -2875 5205 -2845
rect 5525 -1335 5555 -1305
rect 5525 -1400 5555 -1370
rect 5525 -1470 5555 -1440
rect 5525 -1540 5555 -1510
rect 5525 -1610 5555 -1580
rect 5525 -1675 5555 -1645
rect 5525 -1735 5555 -1705
rect 5525 -1800 5555 -1770
rect 5525 -1870 5555 -1840
rect 5525 -1940 5555 -1910
rect 5525 -2010 5555 -1980
rect 5525 -2075 5555 -2045
rect 5525 -2135 5555 -2105
rect 5525 -2200 5555 -2170
rect 5525 -2270 5555 -2240
rect 5525 -2340 5555 -2310
rect 5525 -2410 5555 -2380
rect 5525 -2475 5555 -2445
rect 5525 -2535 5555 -2505
rect 5525 -2600 5555 -2570
rect 5525 -2670 5555 -2640
rect 5525 -2740 5555 -2710
rect 5525 -2810 5555 -2780
rect 5525 -2875 5555 -2845
rect 5875 -1335 5905 -1305
rect 5875 -1400 5905 -1370
rect 5875 -1470 5905 -1440
rect 5875 -1540 5905 -1510
rect 5875 -1610 5905 -1580
rect 5875 -1675 5905 -1645
rect 5875 -1735 5905 -1705
rect 5875 -1800 5905 -1770
rect 5875 -1870 5905 -1840
rect 5875 -1940 5905 -1910
rect 5875 -2010 5905 -1980
rect 5875 -2075 5905 -2045
rect 5875 -2135 5905 -2105
rect 5875 -2200 5905 -2170
rect 5875 -2270 5905 -2240
rect 5875 -2340 5905 -2310
rect 5875 -2410 5905 -2380
rect 5875 -2475 5905 -2445
rect 5875 -2535 5905 -2505
rect 5875 -2600 5905 -2570
rect 5875 -2670 5905 -2640
rect 5875 -2740 5905 -2710
rect 5875 -2810 5905 -2780
rect 5875 -2875 5905 -2845
rect 6225 -1335 6255 -1305
rect 6225 -1400 6255 -1370
rect 6225 -1470 6255 -1440
rect 6225 -1540 6255 -1510
rect 6225 -1610 6255 -1580
rect 6225 -1675 6255 -1645
rect 6225 -1735 6255 -1705
rect 6225 -1800 6255 -1770
rect 6225 -1870 6255 -1840
rect 6225 -1940 6255 -1910
rect 6225 -2010 6255 -1980
rect 6225 -2075 6255 -2045
rect 6225 -2135 6255 -2105
rect 6225 -2200 6255 -2170
rect 6225 -2270 6255 -2240
rect 6225 -2340 6255 -2310
rect 6225 -2410 6255 -2380
rect 6225 -2475 6255 -2445
rect 6225 -2535 6255 -2505
rect 6225 -2600 6255 -2570
rect 6225 -2670 6255 -2640
rect 6225 -2740 6255 -2710
rect 6225 -2810 6255 -2780
rect 6225 -2875 6255 -2845
rect 6575 -1335 6605 -1305
rect 6575 -1400 6605 -1370
rect 6575 -1470 6605 -1440
rect 6575 -1540 6605 -1510
rect 6575 -1610 6605 -1580
rect 6575 -1675 6605 -1645
rect 6575 -1735 6605 -1705
rect 6575 -1800 6605 -1770
rect 6575 -1870 6605 -1840
rect 6575 -1940 6605 -1910
rect 6575 -2010 6605 -1980
rect 6575 -2075 6605 -2045
rect 6575 -2135 6605 -2105
rect 6575 -2200 6605 -2170
rect 6575 -2270 6605 -2240
rect 6575 -2340 6605 -2310
rect 6575 -2410 6605 -2380
rect 6575 -2475 6605 -2445
rect 6575 -2535 6605 -2505
rect 6575 -2600 6605 -2570
rect 6575 -2670 6605 -2640
rect 6575 -2740 6605 -2710
rect 6575 -2810 6605 -2780
rect 6575 -2875 6605 -2845
rect 6925 -1335 6955 -1305
rect 6925 -1400 6955 -1370
rect 6925 -1470 6955 -1440
rect 6925 -1540 6955 -1510
rect 6925 -1610 6955 -1580
rect 6925 -1675 6955 -1645
rect 6925 -1735 6955 -1705
rect 6925 -1800 6955 -1770
rect 6925 -1870 6955 -1840
rect 6925 -1940 6955 -1910
rect 6925 -2010 6955 -1980
rect 6925 -2075 6955 -2045
rect 6925 -2135 6955 -2105
rect 6925 -2200 6955 -2170
rect 6925 -2270 6955 -2240
rect 6925 -2340 6955 -2310
rect 6925 -2410 6955 -2380
rect 6925 -2475 6955 -2445
rect 6925 -2535 6955 -2505
rect 6925 -2600 6955 -2570
rect 6925 -2670 6955 -2640
rect 6925 -2740 6955 -2710
rect 6925 -2810 6955 -2780
rect 6925 -2875 6955 -2845
rect 7275 -1335 7305 -1305
rect 7275 -1400 7305 -1370
rect 7275 -1470 7305 -1440
rect 7275 -1540 7305 -1510
rect 7275 -1610 7305 -1580
rect 7275 -1675 7305 -1645
rect 7275 -1735 7305 -1705
rect 7275 -1800 7305 -1770
rect 7275 -1870 7305 -1840
rect 7275 -1940 7305 -1910
rect 7275 -2010 7305 -1980
rect 7275 -2075 7305 -2045
rect 7275 -2135 7305 -2105
rect 7275 -2200 7305 -2170
rect 7275 -2270 7305 -2240
rect 7275 -2340 7305 -2310
rect 7275 -2410 7305 -2380
rect 7275 -2475 7305 -2445
rect 7275 -2535 7305 -2505
rect 7275 -2600 7305 -2570
rect 7275 -2670 7305 -2640
rect 7275 -2740 7305 -2710
rect 7275 -2810 7305 -2780
rect 7275 -2875 7305 -2845
rect 7625 -1335 7655 -1305
rect 7625 -1400 7655 -1370
rect 7625 -1470 7655 -1440
rect 7625 -1540 7655 -1510
rect 7625 -1610 7655 -1580
rect 7625 -1675 7655 -1645
rect 7625 -1735 7655 -1705
rect 7625 -1800 7655 -1770
rect 7625 -1870 7655 -1840
rect 7625 -1940 7655 -1910
rect 7625 -2010 7655 -1980
rect 7625 -2075 7655 -2045
rect 7625 -2135 7655 -2105
rect 7625 -2200 7655 -2170
rect 7625 -2270 7655 -2240
rect 7625 -2340 7655 -2310
rect 7625 -2410 7655 -2380
rect 7625 -2475 7655 -2445
rect 7625 -2535 7655 -2505
rect 7625 -2600 7655 -2570
rect 7625 -2670 7655 -2640
rect 7625 -2740 7655 -2710
rect 7625 -2810 7655 -2780
rect 7625 -2875 7655 -2845
rect 7975 -1335 8005 -1305
rect 7975 -1400 8005 -1370
rect 7975 -1470 8005 -1440
rect 7975 -1540 8005 -1510
rect 7975 -1610 8005 -1580
rect 7975 -1675 8005 -1645
rect 7975 -1735 8005 -1705
rect 7975 -1800 8005 -1770
rect 7975 -1870 8005 -1840
rect 7975 -1940 8005 -1910
rect 7975 -2010 8005 -1980
rect 7975 -2075 8005 -2045
rect 7975 -2135 8005 -2105
rect 7975 -2200 8005 -2170
rect 7975 -2270 8005 -2240
rect 7975 -2340 8005 -2310
rect 7975 -2410 8005 -2380
rect 7975 -2475 8005 -2445
rect 7975 -2535 8005 -2505
rect 7975 -2600 8005 -2570
rect 7975 -2670 8005 -2640
rect 7975 -2740 8005 -2710
rect 7975 -2810 8005 -2780
rect 7975 -2875 8005 -2845
rect 8325 -1335 8355 -1305
rect 8325 -1400 8355 -1370
rect 8325 -1470 8355 -1440
rect 8325 -1540 8355 -1510
rect 8325 -1610 8355 -1580
rect 8325 -1675 8355 -1645
rect 8325 -1735 8355 -1705
rect 8325 -1800 8355 -1770
rect 8325 -1870 8355 -1840
rect 8325 -1940 8355 -1910
rect 8325 -2010 8355 -1980
rect 8325 -2075 8355 -2045
rect 8325 -2135 8355 -2105
rect 8325 -2200 8355 -2170
rect 8325 -2270 8355 -2240
rect 8325 -2340 8355 -2310
rect 8325 -2410 8355 -2380
rect 8325 -2475 8355 -2445
rect 8325 -2535 8355 -2505
rect 8325 -2600 8355 -2570
rect 8325 -2670 8355 -2640
rect 8325 -2740 8355 -2710
rect 8325 -2810 8355 -2780
rect 8325 -2875 8355 -2845
rect 8675 -1335 8705 -1305
rect 8675 -1400 8705 -1370
rect 8675 -1470 8705 -1440
rect 8675 -1540 8705 -1510
rect 8675 -1610 8705 -1580
rect 8675 -1675 8705 -1645
rect 8675 -1735 8705 -1705
rect 8675 -1800 8705 -1770
rect 8675 -1870 8705 -1840
rect 8675 -1940 8705 -1910
rect 8675 -2010 8705 -1980
rect 8675 -2075 8705 -2045
rect 8675 -2135 8705 -2105
rect 8675 -2200 8705 -2170
rect 8675 -2270 8705 -2240
rect 8675 -2340 8705 -2310
rect 8675 -2410 8705 -2380
rect 8675 -2475 8705 -2445
rect 8675 -2535 8705 -2505
rect 8675 -2600 8705 -2570
rect 8675 -2670 8705 -2640
rect 8675 -2740 8705 -2710
rect 8675 -2810 8705 -2780
rect 8675 -2875 8705 -2845
rect 9025 -1335 9055 -1305
rect 9025 -1400 9055 -1370
rect 9025 -1470 9055 -1440
rect 9025 -1540 9055 -1510
rect 9025 -1610 9055 -1580
rect 9025 -1675 9055 -1645
rect 9025 -1735 9055 -1705
rect 9025 -1800 9055 -1770
rect 9025 -1870 9055 -1840
rect 9025 -1940 9055 -1910
rect 9025 -2010 9055 -1980
rect 9025 -2075 9055 -2045
rect 9025 -2135 9055 -2105
rect 9025 -2200 9055 -2170
rect 9025 -2270 9055 -2240
rect 9025 -2340 9055 -2310
rect 9025 -2410 9055 -2380
rect 9025 -2475 9055 -2445
rect 9025 -2535 9055 -2505
rect 9025 -2600 9055 -2570
rect 9025 -2670 9055 -2640
rect 9025 -2740 9055 -2710
rect 9025 -2810 9055 -2780
rect 9025 -2875 9055 -2845
<< metal2 >>
rect 2100 19310 2160 19325
rect 2100 19280 2115 19310
rect 2145 19280 2160 19310
rect 2100 19245 2160 19280
rect 2100 19215 2115 19245
rect 2145 19215 2160 19245
rect 2100 19175 2160 19215
rect 2100 19145 2115 19175
rect 2145 19145 2160 19175
rect 2100 19105 2160 19145
rect 2100 19075 2115 19105
rect 2145 19075 2160 19105
rect 2100 19035 2160 19075
rect 2100 19005 2115 19035
rect 2145 19005 2160 19035
rect 2100 18970 2160 19005
rect 2100 18940 2115 18970
rect 2145 18940 2160 18970
rect 2100 18910 2160 18940
rect 2100 18880 2115 18910
rect 2145 18880 2160 18910
rect 2100 18845 2160 18880
rect 2100 18815 2115 18845
rect 2145 18815 2160 18845
rect 2100 18775 2160 18815
rect 2100 18745 2115 18775
rect 2145 18745 2160 18775
rect 2100 18705 2160 18745
rect 2100 18675 2115 18705
rect 2145 18675 2160 18705
rect 2100 18635 2160 18675
rect 2100 18605 2115 18635
rect 2145 18605 2160 18635
rect 2100 18570 2160 18605
rect 2100 18540 2115 18570
rect 2145 18540 2160 18570
rect 2100 18510 2160 18540
rect 2100 18480 2115 18510
rect 2145 18480 2160 18510
rect 2100 18445 2160 18480
rect 2100 18415 2115 18445
rect 2145 18415 2160 18445
rect 2100 18375 2160 18415
rect 2100 18345 2115 18375
rect 2145 18345 2160 18375
rect 2100 18305 2160 18345
rect 2100 18275 2115 18305
rect 2145 18275 2160 18305
rect 2100 18235 2160 18275
rect 2100 18205 2115 18235
rect 2145 18205 2160 18235
rect 2100 18170 2160 18205
rect 2100 18140 2115 18170
rect 2145 18140 2160 18170
rect 2100 18110 2160 18140
rect 2100 18080 2115 18110
rect 2145 18080 2160 18110
rect 2100 18045 2160 18080
rect 2100 18015 2115 18045
rect 2145 18015 2160 18045
rect 2100 17975 2160 18015
rect 2100 17945 2115 17975
rect 2145 17945 2160 17975
rect 2100 17905 2160 17945
rect 2100 17875 2115 17905
rect 2145 17875 2160 17905
rect 2100 17835 2160 17875
rect 2100 17805 2115 17835
rect 2145 17805 2160 17835
rect 2100 17770 2160 17805
rect 2100 17740 2115 17770
rect 2145 17740 2160 17770
rect 2100 17725 2160 17740
rect 6690 19310 6750 19325
rect 6690 19280 6705 19310
rect 6735 19280 6750 19310
rect 6690 19245 6750 19280
rect 6690 19215 6705 19245
rect 6735 19215 6750 19245
rect 6690 19175 6750 19215
rect 6690 19145 6705 19175
rect 6735 19145 6750 19175
rect 6690 19105 6750 19145
rect 6690 19075 6705 19105
rect 6735 19075 6750 19105
rect 6690 19035 6750 19075
rect 6690 19005 6705 19035
rect 6735 19005 6750 19035
rect 6690 18970 6750 19005
rect 6690 18940 6705 18970
rect 6735 18940 6750 18970
rect 6690 18910 6750 18940
rect 6690 18880 6705 18910
rect 6735 18880 6750 18910
rect 6690 18845 6750 18880
rect 6690 18815 6705 18845
rect 6735 18815 6750 18845
rect 6690 18775 6750 18815
rect 6690 18745 6705 18775
rect 6735 18745 6750 18775
rect 6690 18705 6750 18745
rect 6690 18675 6705 18705
rect 6735 18675 6750 18705
rect 6690 18635 6750 18675
rect 6690 18605 6705 18635
rect 6735 18605 6750 18635
rect 6690 18570 6750 18605
rect 6690 18540 6705 18570
rect 6735 18540 6750 18570
rect 6690 18510 6750 18540
rect 6690 18480 6705 18510
rect 6735 18480 6750 18510
rect 6690 18445 6750 18480
rect 6690 18415 6705 18445
rect 6735 18415 6750 18445
rect 6690 18375 6750 18415
rect 6690 18345 6705 18375
rect 6735 18345 6750 18375
rect 6690 18305 6750 18345
rect 6690 18275 6705 18305
rect 6735 18275 6750 18305
rect 6690 18235 6750 18275
rect 6690 18205 6705 18235
rect 6735 18205 6750 18235
rect 6690 18170 6750 18205
rect 6690 18140 6705 18170
rect 6735 18140 6750 18170
rect 6690 18110 6750 18140
rect 6690 18080 6705 18110
rect 6735 18080 6750 18110
rect 6690 18045 6750 18080
rect 6690 18015 6705 18045
rect 6735 18015 6750 18045
rect 6690 17975 6750 18015
rect 6690 17945 6705 17975
rect 6735 17945 6750 17975
rect 6690 17905 6750 17945
rect 6690 17875 6705 17905
rect 6735 17875 6750 17905
rect 6690 17835 6750 17875
rect 6690 17805 6705 17835
rect 6735 17805 6750 17835
rect 6690 17770 6750 17805
rect 6690 17740 6705 17770
rect 6735 17740 6750 17770
rect 6690 17725 6750 17740
rect 2205 15925 2325 15930
rect 2205 15895 2210 15925
rect 2240 15895 2250 15925
rect 2280 15895 2290 15925
rect 2320 15920 2325 15925
rect 2320 15900 2385 15920
rect 2320 15895 2325 15900
rect 2205 15890 2325 15895
rect 2070 15690 2970 15695
rect 2070 15660 2075 15690
rect 2105 15660 2115 15690
rect 2145 15660 2155 15690
rect 2185 15660 2970 15690
rect 2070 15650 2970 15660
rect 2070 15620 2075 15650
rect 2105 15620 2115 15650
rect 2145 15620 2155 15650
rect 2185 15620 2970 15650
rect 2070 15610 2970 15620
rect 2070 15580 2075 15610
rect 2105 15580 2115 15610
rect 2145 15580 2155 15610
rect 2185 15580 2970 15610
rect 2070 15575 2970 15580
rect 6650 15595 6780 15600
rect 6650 15565 6665 15595
rect 6695 15565 6705 15595
rect 6735 15565 6745 15595
rect 6775 15565 6780 15595
rect 6650 15555 6780 15565
rect 6650 15525 6665 15555
rect 6695 15525 6705 15555
rect 6735 15525 6745 15555
rect 6775 15525 6780 15555
rect 6650 15515 6780 15525
rect 6650 15485 6665 15515
rect 6695 15485 6705 15515
rect 6735 15485 6745 15515
rect 6775 15485 6780 15515
rect 6650 15480 6780 15485
rect 5690 12925 6780 12930
rect 5690 12895 6665 12925
rect 6695 12895 6705 12925
rect 6735 12895 6745 12925
rect 6775 12895 6780 12925
rect 5690 12885 6780 12895
rect 5690 12855 6665 12885
rect 6695 12855 6705 12885
rect 6735 12855 6745 12885
rect 6775 12855 6780 12885
rect 5690 12845 6780 12855
rect 5690 12815 6665 12845
rect 6695 12815 6705 12845
rect 6735 12815 6745 12845
rect 6775 12815 6780 12845
rect 5690 12810 6780 12815
rect 2070 12710 3355 12715
rect 2070 12680 2075 12710
rect 2105 12680 2115 12710
rect 2145 12680 2155 12710
rect 2185 12680 3355 12710
rect 2070 12670 3355 12680
rect 2070 12640 2075 12670
rect 2105 12640 2115 12670
rect 2145 12640 2155 12670
rect 2185 12640 3355 12670
rect 2070 12635 3355 12640
rect 2070 12550 3800 12555
rect 2070 12520 2075 12550
rect 2105 12520 2115 12550
rect 2145 12520 2155 12550
rect 2185 12520 3800 12550
rect 2070 12510 3800 12520
rect 2070 12480 2075 12510
rect 2105 12480 2115 12510
rect 2145 12480 2155 12510
rect 2185 12480 3800 12510
rect 2070 12470 3800 12480
rect 2070 12440 2075 12470
rect 2105 12440 2115 12470
rect 2145 12440 2155 12470
rect 2185 12440 3800 12470
rect 2070 12435 3800 12440
rect 5670 12150 6780 12155
rect 5670 12120 6665 12150
rect 6695 12120 6705 12150
rect 6735 12120 6745 12150
rect 6775 12120 6780 12150
rect 5670 12110 6780 12120
rect 5670 12080 6665 12110
rect 6695 12080 6705 12110
rect 6735 12080 6745 12110
rect 6775 12080 6780 12110
rect 5670 12070 6780 12080
rect 5670 12040 6665 12070
rect 6695 12040 6705 12070
rect 6735 12040 6745 12070
rect 6775 12040 6780 12070
rect 5670 12035 6780 12040
rect 5870 11165 6780 11170
rect 5870 11135 6665 11165
rect 6695 11135 6705 11165
rect 6735 11135 6745 11165
rect 6775 11135 6780 11165
rect 5870 11125 6780 11135
rect 5870 11095 6665 11125
rect 6695 11095 6705 11125
rect 6735 11095 6745 11125
rect 6775 11095 6780 11125
rect 5870 11085 6780 11095
rect 5870 11055 6665 11085
rect 6695 11055 6705 11085
rect 6735 11055 6745 11085
rect 6775 11055 6780 11085
rect 5870 11050 6780 11055
rect 5855 10440 6780 10445
rect 5855 10410 6665 10440
rect 6695 10410 6705 10440
rect 6735 10410 6745 10440
rect 6775 10410 6780 10440
rect 5855 10400 6780 10410
rect 5855 10370 6665 10400
rect 6695 10370 6705 10400
rect 6735 10370 6745 10400
rect 6775 10370 6780 10400
rect 5855 10360 6780 10370
rect 5855 10330 6665 10360
rect 6695 10330 6705 10360
rect 6735 10330 6745 10360
rect 6775 10330 6780 10360
rect 5855 10325 6780 10330
rect 5925 10080 6780 10085
rect 5925 10050 6665 10080
rect 6695 10050 6705 10080
rect 6735 10050 6745 10080
rect 6775 10050 6780 10080
rect 5925 10040 6780 10050
rect 5925 10010 6665 10040
rect 6695 10010 6705 10040
rect 6735 10010 6745 10040
rect 6775 10010 6780 10040
rect 5925 10000 6780 10010
rect 5925 9970 6665 10000
rect 6695 9970 6705 10000
rect 6735 9970 6745 10000
rect 6775 9970 6780 10000
rect 5925 9965 6780 9970
rect 3740 9915 3780 9920
rect 3700 9910 3790 9915
rect -90 9635 -30 9650
rect -90 9605 -75 9635
rect -45 9605 -30 9635
rect -90 9570 -30 9605
rect -90 9540 -75 9570
rect -45 9540 -30 9570
rect -90 9500 -30 9540
rect -90 9470 -75 9500
rect -45 9470 -30 9500
rect -90 9430 -30 9470
rect -90 9400 -75 9430
rect -45 9400 -30 9430
rect -90 9360 -30 9400
rect -90 9330 -75 9360
rect -45 9330 -30 9360
rect -90 9295 -30 9330
rect -90 9265 -75 9295
rect -45 9265 -30 9295
rect -90 9235 -30 9265
rect -90 9205 -75 9235
rect -45 9205 -30 9235
rect -90 9170 -30 9205
rect -90 9140 -75 9170
rect -45 9140 -30 9170
rect -90 9100 -30 9140
rect -90 9070 -75 9100
rect -45 9070 -30 9100
rect -90 9030 -30 9070
rect -90 9000 -75 9030
rect -45 9000 -30 9030
rect -90 8960 -30 9000
rect -90 8930 -75 8960
rect -45 8930 -30 8960
rect -90 8895 -30 8930
rect -90 8865 -75 8895
rect -45 8865 -30 8895
rect -90 8835 -30 8865
rect -90 8805 -75 8835
rect -45 8805 -30 8835
rect -90 8770 -30 8805
rect -90 8740 -75 8770
rect -45 8740 -30 8770
rect -90 8700 -30 8740
rect -90 8670 -75 8700
rect -45 8670 -30 8700
rect -90 8630 -30 8670
rect -90 8600 -75 8630
rect -45 8600 -30 8630
rect -90 8560 -30 8600
rect -90 8530 -75 8560
rect -45 8530 -30 8560
rect -90 8495 -30 8530
rect -90 8465 -75 8495
rect -45 8465 -30 8495
rect -90 8435 -30 8465
rect -90 8405 -75 8435
rect -45 8405 -30 8435
rect -90 8370 -30 8405
rect -90 8340 -75 8370
rect -45 8340 -30 8370
rect -90 8300 -30 8340
rect -90 8270 -75 8300
rect -45 8270 -30 8300
rect -90 8230 -30 8270
rect -90 8200 -75 8230
rect -45 8200 -30 8230
rect -90 8160 -30 8200
rect -90 8130 -75 8160
rect -45 8130 -30 8160
rect -90 8095 -30 8130
rect -90 8065 -75 8095
rect -45 8065 -30 8095
rect -90 8035 -30 8065
rect -90 8005 -75 8035
rect -45 8005 -30 8035
rect -90 7970 -30 8005
rect -90 7940 -75 7970
rect -45 7940 -30 7970
rect -90 7900 -30 7940
rect -90 7870 -75 7900
rect -45 7870 -30 7900
rect -90 7830 -30 7870
rect -90 7800 -75 7830
rect -45 7800 -30 7830
rect -90 7760 -30 7800
rect -90 7730 -75 7760
rect -45 7730 -30 7760
rect -90 7695 -30 7730
rect -90 7665 -75 7695
rect -45 7665 -30 7695
rect -90 7635 -30 7665
rect -90 7605 -75 7635
rect -45 7605 -30 7635
rect -90 7570 -30 7605
rect -90 7540 -75 7570
rect -45 7540 -30 7570
rect -90 7500 -30 7540
rect -90 7470 -75 7500
rect -45 7470 -30 7500
rect -90 7430 -30 7470
rect -90 7400 -75 7430
rect -45 7400 -30 7430
rect -90 7360 -30 7400
rect -90 7330 -75 7360
rect -45 7330 -30 7360
rect -90 7295 -30 7330
rect -90 7265 -75 7295
rect -45 7265 -30 7295
rect -90 7235 -30 7265
rect -90 7205 -75 7235
rect -45 7205 -30 7235
rect -90 7170 -30 7205
rect -90 7140 -75 7170
rect -45 7140 -30 7170
rect -90 7100 -30 7140
rect -90 7070 -75 7100
rect -45 7070 -30 7100
rect -90 7030 -30 7070
rect -90 7000 -75 7030
rect -45 7000 -30 7030
rect -90 6960 -30 7000
rect -90 6930 -75 6960
rect -45 6930 -30 6960
rect -90 6895 -30 6930
rect -90 6865 -75 6895
rect -45 6865 -30 6895
rect -90 6835 -30 6865
rect -90 6805 -75 6835
rect -45 6805 -30 6835
rect -90 6770 -30 6805
rect -90 6740 -75 6770
rect -45 6740 -30 6770
rect -90 6700 -30 6740
rect -90 6670 -75 6700
rect -45 6670 -30 6700
rect -90 6630 -30 6670
rect -90 6600 -75 6630
rect -45 6600 -30 6630
rect -90 6560 -30 6600
rect -90 6530 -75 6560
rect -45 6530 -30 6560
rect -90 6495 -30 6530
rect -90 6465 -75 6495
rect -45 6465 -30 6495
rect -90 6450 -30 6465
rect 260 9635 320 9650
rect 260 9605 275 9635
rect 305 9605 320 9635
rect 260 9570 320 9605
rect 260 9540 275 9570
rect 305 9540 320 9570
rect 260 9500 320 9540
rect 260 9470 275 9500
rect 305 9470 320 9500
rect 260 9430 320 9470
rect 260 9400 275 9430
rect 305 9400 320 9430
rect 260 9360 320 9400
rect 260 9330 275 9360
rect 305 9330 320 9360
rect 260 9295 320 9330
rect 260 9265 275 9295
rect 305 9265 320 9295
rect 260 9235 320 9265
rect 260 9205 275 9235
rect 305 9205 320 9235
rect 260 9170 320 9205
rect 260 9140 275 9170
rect 305 9140 320 9170
rect 260 9100 320 9140
rect 260 9070 275 9100
rect 305 9070 320 9100
rect 260 9030 320 9070
rect 260 9000 275 9030
rect 305 9000 320 9030
rect 260 8960 320 9000
rect 260 8930 275 8960
rect 305 8930 320 8960
rect 260 8895 320 8930
rect 260 8865 275 8895
rect 305 8865 320 8895
rect 260 8835 320 8865
rect 260 8805 275 8835
rect 305 8805 320 8835
rect 260 8770 320 8805
rect 260 8740 275 8770
rect 305 8740 320 8770
rect 260 8700 320 8740
rect 260 8670 275 8700
rect 305 8670 320 8700
rect 260 8630 320 8670
rect 260 8600 275 8630
rect 305 8600 320 8630
rect 260 8560 320 8600
rect 260 8530 275 8560
rect 305 8530 320 8560
rect 260 8495 320 8530
rect 260 8465 275 8495
rect 305 8465 320 8495
rect 260 8435 320 8465
rect 260 8405 275 8435
rect 305 8405 320 8435
rect 260 8370 320 8405
rect 260 8340 275 8370
rect 305 8340 320 8370
rect 260 8300 320 8340
rect 260 8270 275 8300
rect 305 8270 320 8300
rect 260 8230 320 8270
rect 260 8200 275 8230
rect 305 8200 320 8230
rect 260 8160 320 8200
rect 260 8130 275 8160
rect 305 8130 320 8160
rect 260 8095 320 8130
rect 260 8065 275 8095
rect 305 8065 320 8095
rect 260 8035 320 8065
rect 260 8005 275 8035
rect 305 8005 320 8035
rect 260 7970 320 8005
rect 260 7940 275 7970
rect 305 7940 320 7970
rect 260 7900 320 7940
rect 260 7870 275 7900
rect 305 7870 320 7900
rect 260 7830 320 7870
rect 260 7800 275 7830
rect 305 7800 320 7830
rect 260 7760 320 7800
rect 260 7730 275 7760
rect 305 7730 320 7760
rect 260 7695 320 7730
rect 260 7665 275 7695
rect 305 7665 320 7695
rect 260 7635 320 7665
rect 260 7605 275 7635
rect 305 7605 320 7635
rect 260 7570 320 7605
rect 260 7540 275 7570
rect 305 7540 320 7570
rect 260 7500 320 7540
rect 260 7470 275 7500
rect 305 7470 320 7500
rect 260 7430 320 7470
rect 260 7400 275 7430
rect 305 7400 320 7430
rect 260 7360 320 7400
rect 260 7330 275 7360
rect 305 7330 320 7360
rect 260 7295 320 7330
rect 260 7265 275 7295
rect 305 7265 320 7295
rect 260 7235 320 7265
rect 260 7205 275 7235
rect 305 7205 320 7235
rect 260 7170 320 7205
rect 260 7140 275 7170
rect 305 7140 320 7170
rect 260 7100 320 7140
rect 260 7070 275 7100
rect 305 7070 320 7100
rect 260 7030 320 7070
rect 260 7000 275 7030
rect 305 7000 320 7030
rect 260 6960 320 7000
rect 260 6930 275 6960
rect 305 6930 320 6960
rect 260 6895 320 6930
rect 260 6865 275 6895
rect 305 6865 320 6895
rect 260 6835 320 6865
rect 260 6805 275 6835
rect 305 6805 320 6835
rect 260 6770 320 6805
rect 260 6740 275 6770
rect 305 6740 320 6770
rect 260 6700 320 6740
rect 260 6670 275 6700
rect 305 6670 320 6700
rect 260 6630 320 6670
rect 260 6600 275 6630
rect 305 6600 320 6630
rect 260 6560 320 6600
rect 260 6530 275 6560
rect 305 6530 320 6560
rect 260 6495 320 6530
rect 260 6465 275 6495
rect 305 6465 320 6495
rect 260 6450 320 6465
rect 610 9635 670 9650
rect 610 9605 625 9635
rect 655 9605 670 9635
rect 610 9570 670 9605
rect 610 9540 625 9570
rect 655 9540 670 9570
rect 610 9500 670 9540
rect 610 9470 625 9500
rect 655 9470 670 9500
rect 610 9430 670 9470
rect 610 9400 625 9430
rect 655 9400 670 9430
rect 610 9360 670 9400
rect 610 9330 625 9360
rect 655 9330 670 9360
rect 610 9295 670 9330
rect 610 9265 625 9295
rect 655 9265 670 9295
rect 610 9235 670 9265
rect 610 9205 625 9235
rect 655 9205 670 9235
rect 610 9170 670 9205
rect 610 9140 625 9170
rect 655 9140 670 9170
rect 610 9100 670 9140
rect 610 9070 625 9100
rect 655 9070 670 9100
rect 610 9030 670 9070
rect 610 9000 625 9030
rect 655 9000 670 9030
rect 610 8960 670 9000
rect 610 8930 625 8960
rect 655 8930 670 8960
rect 610 8895 670 8930
rect 610 8865 625 8895
rect 655 8865 670 8895
rect 610 8835 670 8865
rect 610 8805 625 8835
rect 655 8805 670 8835
rect 610 8770 670 8805
rect 610 8740 625 8770
rect 655 8740 670 8770
rect 610 8700 670 8740
rect 610 8670 625 8700
rect 655 8670 670 8700
rect 610 8630 670 8670
rect 610 8600 625 8630
rect 655 8600 670 8630
rect 610 8560 670 8600
rect 610 8530 625 8560
rect 655 8530 670 8560
rect 610 8495 670 8530
rect 610 8465 625 8495
rect 655 8465 670 8495
rect 610 8435 670 8465
rect 610 8405 625 8435
rect 655 8405 670 8435
rect 610 8370 670 8405
rect 610 8340 625 8370
rect 655 8340 670 8370
rect 610 8300 670 8340
rect 610 8270 625 8300
rect 655 8270 670 8300
rect 610 8230 670 8270
rect 610 8200 625 8230
rect 655 8200 670 8230
rect 610 8160 670 8200
rect 610 8130 625 8160
rect 655 8130 670 8160
rect 610 8095 670 8130
rect 610 8065 625 8095
rect 655 8065 670 8095
rect 610 8035 670 8065
rect 610 8005 625 8035
rect 655 8005 670 8035
rect 610 7970 670 8005
rect 610 7940 625 7970
rect 655 7940 670 7970
rect 610 7900 670 7940
rect 610 7870 625 7900
rect 655 7870 670 7900
rect 610 7830 670 7870
rect 610 7800 625 7830
rect 655 7800 670 7830
rect 610 7760 670 7800
rect 610 7730 625 7760
rect 655 7730 670 7760
rect 610 7695 670 7730
rect 610 7665 625 7695
rect 655 7665 670 7695
rect 610 7635 670 7665
rect 610 7605 625 7635
rect 655 7605 670 7635
rect 610 7570 670 7605
rect 610 7540 625 7570
rect 655 7540 670 7570
rect 610 7500 670 7540
rect 610 7470 625 7500
rect 655 7470 670 7500
rect 610 7430 670 7470
rect 610 7400 625 7430
rect 655 7400 670 7430
rect 610 7360 670 7400
rect 610 7330 625 7360
rect 655 7330 670 7360
rect 610 7295 670 7330
rect 610 7265 625 7295
rect 655 7265 670 7295
rect 610 7235 670 7265
rect 610 7205 625 7235
rect 655 7205 670 7235
rect 610 7170 670 7205
rect 610 7140 625 7170
rect 655 7140 670 7170
rect 610 7100 670 7140
rect 610 7070 625 7100
rect 655 7070 670 7100
rect 610 7030 670 7070
rect 610 7000 625 7030
rect 655 7000 670 7030
rect 610 6960 670 7000
rect 610 6930 625 6960
rect 655 6930 670 6960
rect 610 6895 670 6930
rect 610 6865 625 6895
rect 655 6865 670 6895
rect 610 6835 670 6865
rect 610 6805 625 6835
rect 655 6805 670 6835
rect 610 6770 670 6805
rect 610 6740 625 6770
rect 655 6740 670 6770
rect 610 6700 670 6740
rect 610 6670 625 6700
rect 655 6670 670 6700
rect 610 6630 670 6670
rect 610 6600 625 6630
rect 655 6600 670 6630
rect 610 6560 670 6600
rect 610 6530 625 6560
rect 655 6530 670 6560
rect 610 6495 670 6530
rect 610 6465 625 6495
rect 655 6465 670 6495
rect 610 6450 670 6465
rect 960 9635 1020 9650
rect 960 9605 975 9635
rect 1005 9605 1020 9635
rect 960 9570 1020 9605
rect 960 9540 975 9570
rect 1005 9540 1020 9570
rect 960 9500 1020 9540
rect 960 9470 975 9500
rect 1005 9470 1020 9500
rect 960 9430 1020 9470
rect 960 9400 975 9430
rect 1005 9400 1020 9430
rect 960 9360 1020 9400
rect 960 9330 975 9360
rect 1005 9330 1020 9360
rect 960 9295 1020 9330
rect 960 9265 975 9295
rect 1005 9265 1020 9295
rect 960 9235 1020 9265
rect 960 9205 975 9235
rect 1005 9205 1020 9235
rect 960 9170 1020 9205
rect 960 9140 975 9170
rect 1005 9140 1020 9170
rect 960 9100 1020 9140
rect 960 9070 975 9100
rect 1005 9070 1020 9100
rect 960 9030 1020 9070
rect 960 9000 975 9030
rect 1005 9000 1020 9030
rect 960 8960 1020 9000
rect 960 8930 975 8960
rect 1005 8930 1020 8960
rect 960 8895 1020 8930
rect 960 8865 975 8895
rect 1005 8865 1020 8895
rect 960 8835 1020 8865
rect 960 8805 975 8835
rect 1005 8805 1020 8835
rect 960 8770 1020 8805
rect 960 8740 975 8770
rect 1005 8740 1020 8770
rect 960 8700 1020 8740
rect 960 8670 975 8700
rect 1005 8670 1020 8700
rect 960 8630 1020 8670
rect 960 8600 975 8630
rect 1005 8600 1020 8630
rect 960 8560 1020 8600
rect 960 8530 975 8560
rect 1005 8530 1020 8560
rect 960 8495 1020 8530
rect 960 8465 975 8495
rect 1005 8465 1020 8495
rect 960 8435 1020 8465
rect 960 8405 975 8435
rect 1005 8405 1020 8435
rect 960 8370 1020 8405
rect 960 8340 975 8370
rect 1005 8340 1020 8370
rect 960 8300 1020 8340
rect 960 8270 975 8300
rect 1005 8270 1020 8300
rect 960 8230 1020 8270
rect 960 8200 975 8230
rect 1005 8200 1020 8230
rect 960 8160 1020 8200
rect 960 8130 975 8160
rect 1005 8130 1020 8160
rect 960 8095 1020 8130
rect 960 8065 975 8095
rect 1005 8065 1020 8095
rect 960 8035 1020 8065
rect 960 8005 975 8035
rect 1005 8005 1020 8035
rect 960 7970 1020 8005
rect 960 7940 975 7970
rect 1005 7940 1020 7970
rect 960 7900 1020 7940
rect 960 7870 975 7900
rect 1005 7870 1020 7900
rect 960 7830 1020 7870
rect 960 7800 975 7830
rect 1005 7800 1020 7830
rect 960 7760 1020 7800
rect 960 7730 975 7760
rect 1005 7730 1020 7760
rect 960 7695 1020 7730
rect 960 7665 975 7695
rect 1005 7665 1020 7695
rect 960 7635 1020 7665
rect 960 7605 975 7635
rect 1005 7605 1020 7635
rect 960 7570 1020 7605
rect 960 7540 975 7570
rect 1005 7540 1020 7570
rect 960 7500 1020 7540
rect 960 7470 975 7500
rect 1005 7470 1020 7500
rect 960 7430 1020 7470
rect 960 7400 975 7430
rect 1005 7400 1020 7430
rect 960 7360 1020 7400
rect 960 7330 975 7360
rect 1005 7330 1020 7360
rect 960 7295 1020 7330
rect 960 7265 975 7295
rect 1005 7265 1020 7295
rect 960 7235 1020 7265
rect 960 7205 975 7235
rect 1005 7205 1020 7235
rect 960 7170 1020 7205
rect 960 7140 975 7170
rect 1005 7140 1020 7170
rect 960 7100 1020 7140
rect 960 7070 975 7100
rect 1005 7070 1020 7100
rect 960 7030 1020 7070
rect 960 7000 975 7030
rect 1005 7000 1020 7030
rect 960 6960 1020 7000
rect 960 6930 975 6960
rect 1005 6930 1020 6960
rect 960 6895 1020 6930
rect 960 6865 975 6895
rect 1005 6865 1020 6895
rect 960 6835 1020 6865
rect 960 6805 975 6835
rect 1005 6805 1020 6835
rect 960 6770 1020 6805
rect 960 6740 975 6770
rect 1005 6740 1020 6770
rect 960 6700 1020 6740
rect 960 6670 975 6700
rect 1005 6670 1020 6700
rect 960 6630 1020 6670
rect 960 6600 975 6630
rect 1005 6600 1020 6630
rect 960 6560 1020 6600
rect 960 6530 975 6560
rect 1005 6530 1020 6560
rect 960 6495 1020 6530
rect 960 6465 975 6495
rect 1005 6465 1020 6495
rect 960 6450 1020 6465
rect 1660 9635 1720 9650
rect 1660 9605 1675 9635
rect 1705 9605 1720 9635
rect 1660 9570 1720 9605
rect 1660 9540 1675 9570
rect 1705 9540 1720 9570
rect 1660 9500 1720 9540
rect 1660 9470 1675 9500
rect 1705 9470 1720 9500
rect 1660 9430 1720 9470
rect 1660 9400 1675 9430
rect 1705 9400 1720 9430
rect 1660 9360 1720 9400
rect 1660 9330 1675 9360
rect 1705 9330 1720 9360
rect 1660 9295 1720 9330
rect 1660 9265 1675 9295
rect 1705 9265 1720 9295
rect 1660 9235 1720 9265
rect 1660 9205 1675 9235
rect 1705 9205 1720 9235
rect 1660 9170 1720 9205
rect 1660 9140 1675 9170
rect 1705 9140 1720 9170
rect 1660 9100 1720 9140
rect 1660 9070 1675 9100
rect 1705 9070 1720 9100
rect 1660 9030 1720 9070
rect 1660 9000 1675 9030
rect 1705 9000 1720 9030
rect 1660 8960 1720 9000
rect 1660 8930 1675 8960
rect 1705 8930 1720 8960
rect 1660 8895 1720 8930
rect 1660 8865 1675 8895
rect 1705 8865 1720 8895
rect 1660 8835 1720 8865
rect 1660 8805 1675 8835
rect 1705 8805 1720 8835
rect 1660 8770 1720 8805
rect 1660 8740 1675 8770
rect 1705 8740 1720 8770
rect 1660 8700 1720 8740
rect 1660 8670 1675 8700
rect 1705 8670 1720 8700
rect 1660 8630 1720 8670
rect 1660 8600 1675 8630
rect 1705 8600 1720 8630
rect 1660 8560 1720 8600
rect 1660 8530 1675 8560
rect 1705 8530 1720 8560
rect 1660 8495 1720 8530
rect 1660 8465 1675 8495
rect 1705 8465 1720 8495
rect 1660 8435 1720 8465
rect 1660 8405 1675 8435
rect 1705 8405 1720 8435
rect 1660 8370 1720 8405
rect 1660 8340 1675 8370
rect 1705 8340 1720 8370
rect 1660 8300 1720 8340
rect 1660 8270 1675 8300
rect 1705 8270 1720 8300
rect 1660 8230 1720 8270
rect 1660 8200 1675 8230
rect 1705 8200 1720 8230
rect 1660 8160 1720 8200
rect 1660 8130 1675 8160
rect 1705 8130 1720 8160
rect 1660 8095 1720 8130
rect 1660 8065 1675 8095
rect 1705 8065 1720 8095
rect 1660 8035 1720 8065
rect 1660 8005 1675 8035
rect 1705 8005 1720 8035
rect 1660 7970 1720 8005
rect 1660 7940 1675 7970
rect 1705 7940 1720 7970
rect 1660 7900 1720 7940
rect 1660 7870 1675 7900
rect 1705 7870 1720 7900
rect 1660 7830 1720 7870
rect 1660 7800 1675 7830
rect 1705 7800 1720 7830
rect 1660 7760 1720 7800
rect 1660 7730 1675 7760
rect 1705 7730 1720 7760
rect 1660 7695 1720 7730
rect 1660 7665 1675 7695
rect 1705 7665 1720 7695
rect 1660 7635 1720 7665
rect 1660 7605 1675 7635
rect 1705 7605 1720 7635
rect 1660 7570 1720 7605
rect 1660 7540 1675 7570
rect 1705 7540 1720 7570
rect 1660 7500 1720 7540
rect 1660 7470 1675 7500
rect 1705 7470 1720 7500
rect 1660 7430 1720 7470
rect 1660 7400 1675 7430
rect 1705 7400 1720 7430
rect 1660 7360 1720 7400
rect 1660 7330 1675 7360
rect 1705 7330 1720 7360
rect 1660 7295 1720 7330
rect 1660 7265 1675 7295
rect 1705 7265 1720 7295
rect 1660 7235 1720 7265
rect 1660 7205 1675 7235
rect 1705 7205 1720 7235
rect 1660 7170 1720 7205
rect 1660 7140 1675 7170
rect 1705 7140 1720 7170
rect 1660 7100 1720 7140
rect 1660 7070 1675 7100
rect 1705 7070 1720 7100
rect 1660 7030 1720 7070
rect 1660 7000 1675 7030
rect 1705 7000 1720 7030
rect 1660 6960 1720 7000
rect 1660 6930 1675 6960
rect 1705 6930 1720 6960
rect 1660 6895 1720 6930
rect 1660 6865 1675 6895
rect 1705 6865 1720 6895
rect 1660 6835 1720 6865
rect 1660 6805 1675 6835
rect 1705 6805 1720 6835
rect 1660 6770 1720 6805
rect 1660 6740 1675 6770
rect 1705 6740 1720 6770
rect 1660 6700 1720 6740
rect 1660 6670 1675 6700
rect 1705 6670 1720 6700
rect 1660 6630 1720 6670
rect 1660 6600 1675 6630
rect 1705 6600 1720 6630
rect 1660 6560 1720 6600
rect 1660 6530 1675 6560
rect 1705 6530 1720 6560
rect 1660 6495 1720 6530
rect 1660 6465 1675 6495
rect 1705 6465 1720 6495
rect 1660 6450 1720 6465
rect 2235 9635 2295 9650
rect 2235 9605 2250 9635
rect 2280 9605 2295 9635
rect 2235 9570 2295 9605
rect 2235 9540 2250 9570
rect 2280 9540 2295 9570
rect 2235 9500 2295 9540
rect 2235 9470 2250 9500
rect 2280 9470 2295 9500
rect 2235 9430 2295 9470
rect 2235 9400 2250 9430
rect 2280 9400 2295 9430
rect 2235 9360 2295 9400
rect 2235 9330 2250 9360
rect 2280 9330 2295 9360
rect 2235 9295 2295 9330
rect 2235 9265 2250 9295
rect 2280 9265 2295 9295
rect 2235 9235 2295 9265
rect 2235 9205 2250 9235
rect 2280 9205 2295 9235
rect 2235 9170 2295 9205
rect 2235 9140 2250 9170
rect 2280 9140 2295 9170
rect 2235 9100 2295 9140
rect 2235 9070 2250 9100
rect 2280 9070 2295 9100
rect 2235 9030 2295 9070
rect 2235 9000 2250 9030
rect 2280 9000 2295 9030
rect 2235 8960 2295 9000
rect 2235 8930 2250 8960
rect 2280 8930 2295 8960
rect 2235 8895 2295 8930
rect 2235 8865 2250 8895
rect 2280 8865 2295 8895
rect 2235 8835 2295 8865
rect 2235 8805 2250 8835
rect 2280 8805 2295 8835
rect 2235 8770 2295 8805
rect 2235 8740 2250 8770
rect 2280 8740 2295 8770
rect 2235 8700 2295 8740
rect 2235 8670 2250 8700
rect 2280 8670 2295 8700
rect 2235 8630 2295 8670
rect 2235 8600 2250 8630
rect 2280 8600 2295 8630
rect 2235 8560 2295 8600
rect 2235 8530 2250 8560
rect 2280 8530 2295 8560
rect 2235 8495 2295 8530
rect 2235 8465 2250 8495
rect 2280 8465 2295 8495
rect 2235 8435 2295 8465
rect 2235 8405 2250 8435
rect 2280 8405 2295 8435
rect 2235 8370 2295 8405
rect 2235 8340 2250 8370
rect 2280 8340 2295 8370
rect 2235 8300 2295 8340
rect 2235 8270 2250 8300
rect 2280 8270 2295 8300
rect 2235 8230 2295 8270
rect 2235 8200 2250 8230
rect 2280 8200 2295 8230
rect 2235 8160 2295 8200
rect 2235 8130 2250 8160
rect 2280 8130 2295 8160
rect 2235 8095 2295 8130
rect 2235 8065 2250 8095
rect 2280 8065 2295 8095
rect 2235 8035 2295 8065
rect 2235 8005 2250 8035
rect 2280 8005 2295 8035
rect 2235 7970 2295 8005
rect 2235 7940 2250 7970
rect 2280 7940 2295 7970
rect 2235 7900 2295 7940
rect 2235 7870 2250 7900
rect 2280 7870 2295 7900
rect 2235 7830 2295 7870
rect 2235 7800 2250 7830
rect 2280 7800 2295 7830
rect 2235 7760 2295 7800
rect 2235 7730 2250 7760
rect 2280 7730 2295 7760
rect 2235 7695 2295 7730
rect 2235 7665 2250 7695
rect 2280 7665 2295 7695
rect 2235 7635 2295 7665
rect 2235 7605 2250 7635
rect 2280 7605 2295 7635
rect 2235 7570 2295 7605
rect 2235 7540 2250 7570
rect 2280 7540 2295 7570
rect 2235 7500 2295 7540
rect 2235 7470 2250 7500
rect 2280 7470 2295 7500
rect 2235 7430 2295 7470
rect 2235 7400 2250 7430
rect 2280 7400 2295 7430
rect 2235 7360 2295 7400
rect 2235 7330 2250 7360
rect 2280 7330 2295 7360
rect 2235 7295 2295 7330
rect 2235 7265 2250 7295
rect 2280 7265 2295 7295
rect 2235 7235 2295 7265
rect 2235 7205 2250 7235
rect 2280 7205 2295 7235
rect 2235 7170 2295 7205
rect 2235 7140 2250 7170
rect 2280 7140 2295 7170
rect 2235 7100 2295 7140
rect 2235 7070 2250 7100
rect 2280 7070 2295 7100
rect 2235 7030 2295 7070
rect 2235 7000 2250 7030
rect 2280 7000 2295 7030
rect 2235 6960 2295 7000
rect 2235 6930 2250 6960
rect 2280 6930 2295 6960
rect 2235 6895 2295 6930
rect 2235 6865 2250 6895
rect 2280 6865 2295 6895
rect 2235 6835 2295 6865
rect 2235 6805 2250 6835
rect 2280 6805 2295 6835
rect 2235 6770 2295 6805
rect 2235 6740 2250 6770
rect 2280 6740 2295 6770
rect 2235 6700 2295 6740
rect 2235 6670 2250 6700
rect 2280 6670 2295 6700
rect 2235 6630 2295 6670
rect 2235 6600 2250 6630
rect 2280 6600 2295 6630
rect 2235 6560 2295 6600
rect 2235 6530 2250 6560
rect 2280 6530 2295 6560
rect 2235 6495 2295 6530
rect 2235 6465 2250 6495
rect 2280 6465 2295 6495
rect 2235 6450 2295 6465
rect 3165 9635 3280 9650
rect 3165 9605 3180 9635
rect 3210 9605 3240 9635
rect 3270 9605 3280 9635
rect 3165 9570 3280 9605
rect 3165 9540 3180 9570
rect 3210 9540 3240 9570
rect 3270 9540 3280 9570
rect 3165 9500 3280 9540
rect 3165 9470 3180 9500
rect 3210 9470 3240 9500
rect 3270 9470 3280 9500
rect 3165 9430 3280 9470
rect 3165 9400 3180 9430
rect 3210 9400 3240 9430
rect 3270 9400 3280 9430
rect 3165 9360 3280 9400
rect 3165 9330 3180 9360
rect 3210 9330 3240 9360
rect 3270 9330 3280 9360
rect 3165 9295 3280 9330
rect 3165 9265 3180 9295
rect 3210 9265 3240 9295
rect 3270 9265 3280 9295
rect 3165 9235 3280 9265
rect 3165 9205 3180 9235
rect 3210 9205 3240 9235
rect 3270 9205 3280 9235
rect 3165 9170 3280 9205
rect 3165 9140 3180 9170
rect 3210 9140 3240 9170
rect 3270 9140 3280 9170
rect 3165 9100 3280 9140
rect 3165 9070 3180 9100
rect 3210 9070 3240 9100
rect 3270 9070 3280 9100
rect 3165 9030 3280 9070
rect 3165 9000 3180 9030
rect 3210 9000 3240 9030
rect 3270 9000 3280 9030
rect 3165 8960 3280 9000
rect 3165 8930 3180 8960
rect 3210 8930 3240 8960
rect 3270 8930 3280 8960
rect 3165 8895 3280 8930
rect 3165 8865 3180 8895
rect 3210 8865 3240 8895
rect 3270 8865 3280 8895
rect 3165 8835 3280 8865
rect 3165 8805 3180 8835
rect 3210 8805 3240 8835
rect 3270 8805 3280 8835
rect 3165 8770 3280 8805
rect 3165 8740 3180 8770
rect 3210 8740 3240 8770
rect 3270 8740 3280 8770
rect 3165 8700 3280 8740
rect 3165 8670 3180 8700
rect 3210 8670 3240 8700
rect 3270 8670 3280 8700
rect 3165 8630 3280 8670
rect 3165 8600 3180 8630
rect 3210 8600 3240 8630
rect 3270 8600 3280 8630
rect 3165 8560 3280 8600
rect 3165 8530 3180 8560
rect 3210 8530 3240 8560
rect 3270 8530 3280 8560
rect 3165 8495 3280 8530
rect 3165 8465 3180 8495
rect 3210 8465 3240 8495
rect 3270 8465 3280 8495
rect 3165 8435 3280 8465
rect 3165 8405 3180 8435
rect 3210 8405 3240 8435
rect 3270 8405 3280 8435
rect 3165 8370 3280 8405
rect 3165 8340 3180 8370
rect 3210 8340 3240 8370
rect 3270 8340 3280 8370
rect 3165 8300 3280 8340
rect 3165 8270 3180 8300
rect 3210 8270 3240 8300
rect 3270 8270 3280 8300
rect 3165 8230 3280 8270
rect 3165 8200 3180 8230
rect 3210 8200 3240 8230
rect 3270 8200 3280 8230
rect 3165 8160 3280 8200
rect 3165 8130 3180 8160
rect 3210 8130 3240 8160
rect 3270 8130 3280 8160
rect 3165 8095 3280 8130
rect 3165 8065 3180 8095
rect 3210 8065 3240 8095
rect 3270 8065 3280 8095
rect 3165 8035 3280 8065
rect 3165 8005 3180 8035
rect 3210 8005 3240 8035
rect 3270 8005 3280 8035
rect 3165 7970 3280 8005
rect 3165 7940 3180 7970
rect 3210 7940 3240 7970
rect 3270 7940 3280 7970
rect 3165 7900 3280 7940
rect 3165 7870 3180 7900
rect 3210 7870 3240 7900
rect 3270 7870 3280 7900
rect 3165 7830 3280 7870
rect 3165 7800 3180 7830
rect 3210 7800 3240 7830
rect 3270 7800 3280 7830
rect 3165 7760 3280 7800
rect 3165 7730 3180 7760
rect 3210 7730 3240 7760
rect 3270 7730 3280 7760
rect 3165 7695 3280 7730
rect 3165 7665 3180 7695
rect 3210 7665 3240 7695
rect 3270 7665 3280 7695
rect 3165 7635 3280 7665
rect 3165 7605 3180 7635
rect 3210 7605 3240 7635
rect 3270 7605 3280 7635
rect 3165 7570 3280 7605
rect 3165 7540 3180 7570
rect 3210 7540 3240 7570
rect 3270 7540 3280 7570
rect 3165 7500 3280 7540
rect 3165 7470 3180 7500
rect 3210 7470 3240 7500
rect 3270 7470 3280 7500
rect 3165 7430 3280 7470
rect 3165 7400 3180 7430
rect 3210 7400 3240 7430
rect 3270 7400 3280 7430
rect 3165 7360 3280 7400
rect 3165 7330 3180 7360
rect 3210 7330 3240 7360
rect 3270 7330 3280 7360
rect 3165 7295 3280 7330
rect 3165 7265 3180 7295
rect 3210 7265 3240 7295
rect 3270 7265 3280 7295
rect 3165 7235 3280 7265
rect 3165 7205 3180 7235
rect 3210 7205 3240 7235
rect 3270 7205 3280 7235
rect 3165 7170 3280 7205
rect 3165 7140 3180 7170
rect 3210 7140 3240 7170
rect 3270 7140 3280 7170
rect 3165 7100 3280 7140
rect 3165 7070 3180 7100
rect 3210 7070 3240 7100
rect 3270 7070 3280 7100
rect 3165 7030 3280 7070
rect 3165 7000 3180 7030
rect 3210 7000 3240 7030
rect 3270 7000 3280 7030
rect 3165 6960 3280 7000
rect 3165 6930 3180 6960
rect 3210 6930 3240 6960
rect 3270 6930 3280 6960
rect 3165 6895 3280 6930
rect 3165 6865 3180 6895
rect 3210 6865 3240 6895
rect 3270 6865 3280 6895
rect 3165 6835 3280 6865
rect 3165 6805 3180 6835
rect 3210 6805 3240 6835
rect 3270 6805 3280 6835
rect 3165 6770 3280 6805
rect 3165 6740 3180 6770
rect 3210 6740 3240 6770
rect 3270 6740 3280 6770
rect 3165 6700 3280 6740
rect 3165 6670 3180 6700
rect 3210 6670 3240 6700
rect 3270 6670 3280 6700
rect 3165 6630 3280 6670
rect 3165 6600 3180 6630
rect 3210 6600 3240 6630
rect 3270 6600 3280 6630
rect 3165 6560 3280 6600
rect 3165 6530 3180 6560
rect 3210 6530 3240 6560
rect 3270 6530 3280 6560
rect 3165 6495 3280 6530
rect 3165 6465 3180 6495
rect 3210 6465 3240 6495
rect 3270 6465 3280 6495
rect 3165 6450 3280 6465
rect 3340 9635 3395 9650
rect 3340 9605 3350 9635
rect 3380 9605 3395 9635
rect 3340 9570 3395 9605
rect 3340 9540 3350 9570
rect 3380 9540 3395 9570
rect 3340 9500 3395 9540
rect 3340 9470 3350 9500
rect 3380 9470 3395 9500
rect 3340 9430 3395 9470
rect 3340 9400 3350 9430
rect 3380 9400 3395 9430
rect 3340 9360 3395 9400
rect 3340 9330 3350 9360
rect 3380 9330 3395 9360
rect 3340 9295 3395 9330
rect 3340 9265 3350 9295
rect 3380 9265 3395 9295
rect 3340 9235 3395 9265
rect 3340 9205 3350 9235
rect 3380 9205 3395 9235
rect 3340 9170 3395 9205
rect 3340 9140 3350 9170
rect 3380 9140 3395 9170
rect 3340 9100 3395 9140
rect 3340 9070 3350 9100
rect 3380 9070 3395 9100
rect 3340 9030 3395 9070
rect 3340 9000 3350 9030
rect 3380 9000 3395 9030
rect 3340 8960 3395 9000
rect 3340 8930 3350 8960
rect 3380 8930 3395 8960
rect 3340 8895 3395 8930
rect 3340 8865 3350 8895
rect 3380 8865 3395 8895
rect 3340 8835 3395 8865
rect 3340 8805 3350 8835
rect 3380 8805 3395 8835
rect 3340 8770 3395 8805
rect 3340 8740 3350 8770
rect 3380 8740 3395 8770
rect 3340 8700 3395 8740
rect 3340 8670 3350 8700
rect 3380 8670 3395 8700
rect 3340 8630 3395 8670
rect 3340 8600 3350 8630
rect 3380 8600 3395 8630
rect 3340 8560 3395 8600
rect 3340 8530 3350 8560
rect 3380 8530 3395 8560
rect 3340 8495 3395 8530
rect 3340 8465 3350 8495
rect 3380 8465 3395 8495
rect 3340 8435 3395 8465
rect 3340 8405 3350 8435
rect 3380 8405 3395 8435
rect 3340 8370 3395 8405
rect 3340 8340 3350 8370
rect 3380 8340 3395 8370
rect 3340 8300 3395 8340
rect 3340 8270 3350 8300
rect 3380 8270 3395 8300
rect 3340 8230 3395 8270
rect 3340 8200 3350 8230
rect 3380 8200 3395 8230
rect 3340 8160 3395 8200
rect 3340 8130 3350 8160
rect 3380 8130 3395 8160
rect 3340 8095 3395 8130
rect 3340 8065 3350 8095
rect 3380 8065 3395 8095
rect 3340 8035 3395 8065
rect 3340 8005 3350 8035
rect 3380 8005 3395 8035
rect 3340 7970 3395 8005
rect 3340 7940 3350 7970
rect 3380 7940 3395 7970
rect 3340 7900 3395 7940
rect 3340 7870 3350 7900
rect 3380 7870 3395 7900
rect 3340 7830 3395 7870
rect 3340 7800 3350 7830
rect 3380 7800 3395 7830
rect 3340 7760 3395 7800
rect 3340 7730 3350 7760
rect 3380 7730 3395 7760
rect 3340 7695 3395 7730
rect 3340 7665 3350 7695
rect 3380 7665 3395 7695
rect 3340 7635 3395 7665
rect 3340 7605 3350 7635
rect 3380 7605 3395 7635
rect 3340 7570 3395 7605
rect 3340 7540 3350 7570
rect 3380 7540 3395 7570
rect 3340 7500 3395 7540
rect 3340 7470 3350 7500
rect 3380 7470 3395 7500
rect 3340 7430 3395 7470
rect 3340 7400 3350 7430
rect 3380 7400 3395 7430
rect 3340 7360 3395 7400
rect 3340 7330 3350 7360
rect 3380 7330 3395 7360
rect 3340 7295 3395 7330
rect 3340 7265 3350 7295
rect 3380 7265 3395 7295
rect 3340 7235 3395 7265
rect 3340 7205 3350 7235
rect 3380 7205 3395 7235
rect 3340 7170 3395 7205
rect 3340 7140 3350 7170
rect 3380 7140 3395 7170
rect 3340 7100 3395 7140
rect 3340 7070 3350 7100
rect 3380 7070 3395 7100
rect 3340 7030 3395 7070
rect 3340 7000 3350 7030
rect 3380 7000 3395 7030
rect 3340 6960 3395 7000
rect 3340 6930 3350 6960
rect 3380 6930 3395 6960
rect 3340 6895 3395 6930
rect 3340 6865 3350 6895
rect 3380 6865 3395 6895
rect 3340 6835 3395 6865
rect 3340 6805 3350 6835
rect 3380 6805 3395 6835
rect 3340 6770 3395 6805
rect 3340 6740 3350 6770
rect 3380 6740 3395 6770
rect 3340 6700 3395 6740
rect 3340 6670 3350 6700
rect 3380 6670 3395 6700
rect 3340 6630 3395 6670
rect 3340 6600 3350 6630
rect 3380 6600 3395 6630
rect 3340 6560 3395 6600
rect 3340 6530 3350 6560
rect 3380 6530 3395 6560
rect 3340 6495 3395 6530
rect 3340 6465 3350 6495
rect 3380 6465 3395 6495
rect 3340 6450 3395 6465
rect 6690 9635 6750 9650
rect 6690 9605 6705 9635
rect 6735 9605 6750 9635
rect 6690 9570 6750 9605
rect 6690 9540 6705 9570
rect 6735 9540 6750 9570
rect 6690 9500 6750 9540
rect 6690 9470 6705 9500
rect 6735 9470 6750 9500
rect 6690 9430 6750 9470
rect 6690 9400 6705 9430
rect 6735 9400 6750 9430
rect 6690 9360 6750 9400
rect 6690 9330 6705 9360
rect 6735 9330 6750 9360
rect 6690 9295 6750 9330
rect 6690 9265 6705 9295
rect 6735 9265 6750 9295
rect 6690 9235 6750 9265
rect 6690 9205 6705 9235
rect 6735 9205 6750 9235
rect 6690 9170 6750 9205
rect 6690 9140 6705 9170
rect 6735 9140 6750 9170
rect 6690 9100 6750 9140
rect 6690 9070 6705 9100
rect 6735 9070 6750 9100
rect 6690 9030 6750 9070
rect 6690 9000 6705 9030
rect 6735 9000 6750 9030
rect 6690 8960 6750 9000
rect 6690 8930 6705 8960
rect 6735 8930 6750 8960
rect 6690 8895 6750 8930
rect 6690 8865 6705 8895
rect 6735 8865 6750 8895
rect 6690 8835 6750 8865
rect 6690 8805 6705 8835
rect 6735 8805 6750 8835
rect 6690 8770 6750 8805
rect 6690 8740 6705 8770
rect 6735 8740 6750 8770
rect 6690 8700 6750 8740
rect 6690 8670 6705 8700
rect 6735 8670 6750 8700
rect 6690 8630 6750 8670
rect 6690 8600 6705 8630
rect 6735 8600 6750 8630
rect 6690 8560 6750 8600
rect 6690 8530 6705 8560
rect 6735 8530 6750 8560
rect 6690 8495 6750 8530
rect 6690 8465 6705 8495
rect 6735 8465 6750 8495
rect 6690 8435 6750 8465
rect 6690 8405 6705 8435
rect 6735 8405 6750 8435
rect 6690 8370 6750 8405
rect 6690 8340 6705 8370
rect 6735 8340 6750 8370
rect 6690 8300 6750 8340
rect 6690 8270 6705 8300
rect 6735 8270 6750 8300
rect 6690 8230 6750 8270
rect 6690 8200 6705 8230
rect 6735 8200 6750 8230
rect 6690 8160 6750 8200
rect 6690 8130 6705 8160
rect 6735 8130 6750 8160
rect 6690 8095 6750 8130
rect 6690 8065 6705 8095
rect 6735 8065 6750 8095
rect 6690 8035 6750 8065
rect 6690 8005 6705 8035
rect 6735 8005 6750 8035
rect 6690 7970 6750 8005
rect 6690 7940 6705 7970
rect 6735 7940 6750 7970
rect 6690 7900 6750 7940
rect 6690 7870 6705 7900
rect 6735 7870 6750 7900
rect 6690 7830 6750 7870
rect 6690 7800 6705 7830
rect 6735 7800 6750 7830
rect 6690 7760 6750 7800
rect 6690 7730 6705 7760
rect 6735 7730 6750 7760
rect 6690 7695 6750 7730
rect 6690 7665 6705 7695
rect 6735 7665 6750 7695
rect 6690 7635 6750 7665
rect 6690 7605 6705 7635
rect 6735 7605 6750 7635
rect 6690 7570 6750 7605
rect 6690 7540 6705 7570
rect 6735 7540 6750 7570
rect 6690 7500 6750 7540
rect 6690 7470 6705 7500
rect 6735 7470 6750 7500
rect 6690 7430 6750 7470
rect 6690 7400 6705 7430
rect 6735 7400 6750 7430
rect 6690 7360 6750 7400
rect 6690 7330 6705 7360
rect 6735 7330 6750 7360
rect 6690 7295 6750 7330
rect 6690 7265 6705 7295
rect 6735 7265 6750 7295
rect 6690 7235 6750 7265
rect 6690 7205 6705 7235
rect 6735 7205 6750 7235
rect 6690 7170 6750 7205
rect 6690 7140 6705 7170
rect 6735 7140 6750 7170
rect 6690 7100 6750 7140
rect 6690 7070 6705 7100
rect 6735 7070 6750 7100
rect 6690 7030 6750 7070
rect 6690 7000 6705 7030
rect 6735 7000 6750 7030
rect 6690 6960 6750 7000
rect 6690 6930 6705 6960
rect 6735 6930 6750 6960
rect 6690 6895 6750 6930
rect 6690 6865 6705 6895
rect 6735 6865 6750 6895
rect 6690 6835 6750 6865
rect 6690 6805 6705 6835
rect 6735 6805 6750 6835
rect 6690 6770 6750 6805
rect 6690 6740 6705 6770
rect 6735 6740 6750 6770
rect 6690 6700 6750 6740
rect 6690 6670 6705 6700
rect 6735 6670 6750 6700
rect 6690 6630 6750 6670
rect 6690 6600 6705 6630
rect 6735 6600 6750 6630
rect 6690 6560 6750 6600
rect 6690 6530 6705 6560
rect 6735 6530 6750 6560
rect 6690 6495 6750 6530
rect 6690 6465 6705 6495
rect 6735 6465 6750 6495
rect 6690 6450 6750 6465
rect 7260 9635 7320 9650
rect 7260 9605 7275 9635
rect 7305 9605 7320 9635
rect 7260 9570 7320 9605
rect 7260 9540 7275 9570
rect 7305 9540 7320 9570
rect 7260 9500 7320 9540
rect 7260 9470 7275 9500
rect 7305 9470 7320 9500
rect 7260 9430 7320 9470
rect 7260 9400 7275 9430
rect 7305 9400 7320 9430
rect 7260 9360 7320 9400
rect 7260 9330 7275 9360
rect 7305 9330 7320 9360
rect 7260 9295 7320 9330
rect 7260 9265 7275 9295
rect 7305 9265 7320 9295
rect 7260 9235 7320 9265
rect 7260 9205 7275 9235
rect 7305 9205 7320 9235
rect 7260 9170 7320 9205
rect 7260 9140 7275 9170
rect 7305 9140 7320 9170
rect 7260 9100 7320 9140
rect 7260 9070 7275 9100
rect 7305 9070 7320 9100
rect 7260 9030 7320 9070
rect 7260 9000 7275 9030
rect 7305 9000 7320 9030
rect 7260 8960 7320 9000
rect 7260 8930 7275 8960
rect 7305 8930 7320 8960
rect 7260 8895 7320 8930
rect 7260 8865 7275 8895
rect 7305 8865 7320 8895
rect 7260 8835 7320 8865
rect 7260 8805 7275 8835
rect 7305 8805 7320 8835
rect 7260 8770 7320 8805
rect 7260 8740 7275 8770
rect 7305 8740 7320 8770
rect 7260 8700 7320 8740
rect 7260 8670 7275 8700
rect 7305 8670 7320 8700
rect 7260 8630 7320 8670
rect 7260 8600 7275 8630
rect 7305 8600 7320 8630
rect 7260 8560 7320 8600
rect 7260 8530 7275 8560
rect 7305 8530 7320 8560
rect 7260 8495 7320 8530
rect 7260 8465 7275 8495
rect 7305 8465 7320 8495
rect 7260 8435 7320 8465
rect 7260 8405 7275 8435
rect 7305 8405 7320 8435
rect 7260 8370 7320 8405
rect 7260 8340 7275 8370
rect 7305 8340 7320 8370
rect 7260 8300 7320 8340
rect 7260 8270 7275 8300
rect 7305 8270 7320 8300
rect 7260 8230 7320 8270
rect 7260 8200 7275 8230
rect 7305 8200 7320 8230
rect 7260 8160 7320 8200
rect 7260 8130 7275 8160
rect 7305 8130 7320 8160
rect 7260 8095 7320 8130
rect 7260 8065 7275 8095
rect 7305 8065 7320 8095
rect 7260 8035 7320 8065
rect 7260 8005 7275 8035
rect 7305 8005 7320 8035
rect 7260 7970 7320 8005
rect 7260 7940 7275 7970
rect 7305 7940 7320 7970
rect 7260 7900 7320 7940
rect 7260 7870 7275 7900
rect 7305 7870 7320 7900
rect 7260 7830 7320 7870
rect 7260 7800 7275 7830
rect 7305 7800 7320 7830
rect 7260 7760 7320 7800
rect 7260 7730 7275 7760
rect 7305 7730 7320 7760
rect 7260 7695 7320 7730
rect 7260 7665 7275 7695
rect 7305 7665 7320 7695
rect 7260 7635 7320 7665
rect 7260 7605 7275 7635
rect 7305 7605 7320 7635
rect 7260 7570 7320 7605
rect 7260 7540 7275 7570
rect 7305 7540 7320 7570
rect 7260 7500 7320 7540
rect 7260 7470 7275 7500
rect 7305 7470 7320 7500
rect 7260 7430 7320 7470
rect 7260 7400 7275 7430
rect 7305 7400 7320 7430
rect 7260 7360 7320 7400
rect 7260 7330 7275 7360
rect 7305 7330 7320 7360
rect 7260 7295 7320 7330
rect 7260 7265 7275 7295
rect 7305 7265 7320 7295
rect 7260 7235 7320 7265
rect 7260 7205 7275 7235
rect 7305 7205 7320 7235
rect 7260 7170 7320 7205
rect 7260 7140 7275 7170
rect 7305 7140 7320 7170
rect 7260 7100 7320 7140
rect 7260 7070 7275 7100
rect 7305 7070 7320 7100
rect 7260 7030 7320 7070
rect 7260 7000 7275 7030
rect 7305 7000 7320 7030
rect 7260 6960 7320 7000
rect 7260 6930 7275 6960
rect 7305 6930 7320 6960
rect 7260 6895 7320 6930
rect 7260 6865 7275 6895
rect 7305 6865 7320 6895
rect 7260 6835 7320 6865
rect 7260 6805 7275 6835
rect 7305 6805 7320 6835
rect 7260 6770 7320 6805
rect 7260 6740 7275 6770
rect 7305 6740 7320 6770
rect 7260 6700 7320 6740
rect 7260 6670 7275 6700
rect 7305 6670 7320 6700
rect 7260 6630 7320 6670
rect 7260 6600 7275 6630
rect 7305 6600 7320 6630
rect 7260 6560 7320 6600
rect 7260 6530 7275 6560
rect 7305 6530 7320 6560
rect 7260 6495 7320 6530
rect 7260 6465 7275 6495
rect 7305 6465 7320 6495
rect 7260 6450 7320 6465
rect 7960 9635 8020 9650
rect 7960 9605 7975 9635
rect 8005 9605 8020 9635
rect 7960 9570 8020 9605
rect 7960 9540 7975 9570
rect 8005 9540 8020 9570
rect 7960 9500 8020 9540
rect 7960 9470 7975 9500
rect 8005 9470 8020 9500
rect 7960 9430 8020 9470
rect 7960 9400 7975 9430
rect 8005 9400 8020 9430
rect 7960 9360 8020 9400
rect 7960 9330 7975 9360
rect 8005 9330 8020 9360
rect 7960 9295 8020 9330
rect 7960 9265 7975 9295
rect 8005 9265 8020 9295
rect 7960 9235 8020 9265
rect 7960 9205 7975 9235
rect 8005 9205 8020 9235
rect 7960 9170 8020 9205
rect 7960 9140 7975 9170
rect 8005 9140 8020 9170
rect 7960 9100 8020 9140
rect 7960 9070 7975 9100
rect 8005 9070 8020 9100
rect 7960 9030 8020 9070
rect 7960 9000 7975 9030
rect 8005 9000 8020 9030
rect 7960 8960 8020 9000
rect 7960 8930 7975 8960
rect 8005 8930 8020 8960
rect 7960 8895 8020 8930
rect 7960 8865 7975 8895
rect 8005 8865 8020 8895
rect 7960 8835 8020 8865
rect 7960 8805 7975 8835
rect 8005 8805 8020 8835
rect 7960 8770 8020 8805
rect 7960 8740 7975 8770
rect 8005 8740 8020 8770
rect 7960 8700 8020 8740
rect 7960 8670 7975 8700
rect 8005 8670 8020 8700
rect 7960 8630 8020 8670
rect 7960 8600 7975 8630
rect 8005 8600 8020 8630
rect 7960 8560 8020 8600
rect 7960 8530 7975 8560
rect 8005 8530 8020 8560
rect 7960 8495 8020 8530
rect 7960 8465 7975 8495
rect 8005 8465 8020 8495
rect 7960 8435 8020 8465
rect 7960 8405 7975 8435
rect 8005 8405 8020 8435
rect 7960 8370 8020 8405
rect 7960 8340 7975 8370
rect 8005 8340 8020 8370
rect 7960 8300 8020 8340
rect 7960 8270 7975 8300
rect 8005 8270 8020 8300
rect 7960 8230 8020 8270
rect 7960 8200 7975 8230
rect 8005 8200 8020 8230
rect 7960 8160 8020 8200
rect 7960 8130 7975 8160
rect 8005 8130 8020 8160
rect 7960 8095 8020 8130
rect 7960 8065 7975 8095
rect 8005 8065 8020 8095
rect 7960 8035 8020 8065
rect 7960 8005 7975 8035
rect 8005 8005 8020 8035
rect 7960 7970 8020 8005
rect 7960 7940 7975 7970
rect 8005 7940 8020 7970
rect 7960 7900 8020 7940
rect 7960 7870 7975 7900
rect 8005 7870 8020 7900
rect 7960 7830 8020 7870
rect 7960 7800 7975 7830
rect 8005 7800 8020 7830
rect 7960 7760 8020 7800
rect 7960 7730 7975 7760
rect 8005 7730 8020 7760
rect 7960 7695 8020 7730
rect 7960 7665 7975 7695
rect 8005 7665 8020 7695
rect 7960 7635 8020 7665
rect 7960 7605 7975 7635
rect 8005 7605 8020 7635
rect 7960 7570 8020 7605
rect 7960 7540 7975 7570
rect 8005 7540 8020 7570
rect 7960 7500 8020 7540
rect 7960 7470 7975 7500
rect 8005 7470 8020 7500
rect 7960 7430 8020 7470
rect 7960 7400 7975 7430
rect 8005 7400 8020 7430
rect 7960 7360 8020 7400
rect 7960 7330 7975 7360
rect 8005 7330 8020 7360
rect 7960 7295 8020 7330
rect 7960 7265 7975 7295
rect 8005 7265 8020 7295
rect 7960 7235 8020 7265
rect 7960 7205 7975 7235
rect 8005 7205 8020 7235
rect 7960 7170 8020 7205
rect 7960 7140 7975 7170
rect 8005 7140 8020 7170
rect 7960 7100 8020 7140
rect 7960 7070 7975 7100
rect 8005 7070 8020 7100
rect 7960 7030 8020 7070
rect 7960 7000 7975 7030
rect 8005 7000 8020 7030
rect 7960 6960 8020 7000
rect 7960 6930 7975 6960
rect 8005 6930 8020 6960
rect 7960 6895 8020 6930
rect 7960 6865 7975 6895
rect 8005 6865 8020 6895
rect 7960 6835 8020 6865
rect 7960 6805 7975 6835
rect 8005 6805 8020 6835
rect 7960 6770 8020 6805
rect 7960 6740 7975 6770
rect 8005 6740 8020 6770
rect 7960 6700 8020 6740
rect 7960 6670 7975 6700
rect 8005 6670 8020 6700
rect 7960 6630 8020 6670
rect 7960 6600 7975 6630
rect 8005 6600 8020 6630
rect 7960 6560 8020 6600
rect 7960 6530 7975 6560
rect 8005 6530 8020 6560
rect 7960 6495 8020 6530
rect 7960 6465 7975 6495
rect 8005 6465 8020 6495
rect 7960 6450 8020 6465
rect 8310 9635 8370 9650
rect 8310 9605 8325 9635
rect 8355 9605 8370 9635
rect 8310 9570 8370 9605
rect 8310 9540 8325 9570
rect 8355 9540 8370 9570
rect 8310 9500 8370 9540
rect 8310 9470 8325 9500
rect 8355 9470 8370 9500
rect 8310 9430 8370 9470
rect 8310 9400 8325 9430
rect 8355 9400 8370 9430
rect 8310 9360 8370 9400
rect 8310 9330 8325 9360
rect 8355 9330 8370 9360
rect 8310 9295 8370 9330
rect 8310 9265 8325 9295
rect 8355 9265 8370 9295
rect 8310 9235 8370 9265
rect 8310 9205 8325 9235
rect 8355 9205 8370 9235
rect 8310 9170 8370 9205
rect 8310 9140 8325 9170
rect 8355 9140 8370 9170
rect 8310 9100 8370 9140
rect 8310 9070 8325 9100
rect 8355 9070 8370 9100
rect 8310 9030 8370 9070
rect 8310 9000 8325 9030
rect 8355 9000 8370 9030
rect 8310 8960 8370 9000
rect 8310 8930 8325 8960
rect 8355 8930 8370 8960
rect 8310 8895 8370 8930
rect 8310 8865 8325 8895
rect 8355 8865 8370 8895
rect 8310 8835 8370 8865
rect 8310 8805 8325 8835
rect 8355 8805 8370 8835
rect 8310 8770 8370 8805
rect 8310 8740 8325 8770
rect 8355 8740 8370 8770
rect 8310 8700 8370 8740
rect 8310 8670 8325 8700
rect 8355 8670 8370 8700
rect 8310 8630 8370 8670
rect 8310 8600 8325 8630
rect 8355 8600 8370 8630
rect 8310 8560 8370 8600
rect 8310 8530 8325 8560
rect 8355 8530 8370 8560
rect 8310 8495 8370 8530
rect 8310 8465 8325 8495
rect 8355 8465 8370 8495
rect 8310 8435 8370 8465
rect 8310 8405 8325 8435
rect 8355 8405 8370 8435
rect 8310 8370 8370 8405
rect 8310 8340 8325 8370
rect 8355 8340 8370 8370
rect 8310 8300 8370 8340
rect 8310 8270 8325 8300
rect 8355 8270 8370 8300
rect 8310 8230 8370 8270
rect 8310 8200 8325 8230
rect 8355 8200 8370 8230
rect 8310 8160 8370 8200
rect 8310 8130 8325 8160
rect 8355 8130 8370 8160
rect 8310 8095 8370 8130
rect 8310 8065 8325 8095
rect 8355 8065 8370 8095
rect 8310 8035 8370 8065
rect 8310 8005 8325 8035
rect 8355 8005 8370 8035
rect 8310 7970 8370 8005
rect 8310 7940 8325 7970
rect 8355 7940 8370 7970
rect 8310 7900 8370 7940
rect 8310 7870 8325 7900
rect 8355 7870 8370 7900
rect 8310 7830 8370 7870
rect 8310 7800 8325 7830
rect 8355 7800 8370 7830
rect 8310 7760 8370 7800
rect 8310 7730 8325 7760
rect 8355 7730 8370 7760
rect 8310 7695 8370 7730
rect 8310 7665 8325 7695
rect 8355 7665 8370 7695
rect 8310 7635 8370 7665
rect 8310 7605 8325 7635
rect 8355 7605 8370 7635
rect 8310 7570 8370 7605
rect 8310 7540 8325 7570
rect 8355 7540 8370 7570
rect 8310 7500 8370 7540
rect 8310 7470 8325 7500
rect 8355 7470 8370 7500
rect 8310 7430 8370 7470
rect 8310 7400 8325 7430
rect 8355 7400 8370 7430
rect 8310 7360 8370 7400
rect 8310 7330 8325 7360
rect 8355 7330 8370 7360
rect 8310 7295 8370 7330
rect 8310 7265 8325 7295
rect 8355 7265 8370 7295
rect 8310 7235 8370 7265
rect 8310 7205 8325 7235
rect 8355 7205 8370 7235
rect 8310 7170 8370 7205
rect 8310 7140 8325 7170
rect 8355 7140 8370 7170
rect 8310 7100 8370 7140
rect 8310 7070 8325 7100
rect 8355 7070 8370 7100
rect 8310 7030 8370 7070
rect 8310 7000 8325 7030
rect 8355 7000 8370 7030
rect 8310 6960 8370 7000
rect 8310 6930 8325 6960
rect 8355 6930 8370 6960
rect 8310 6895 8370 6930
rect 8310 6865 8325 6895
rect 8355 6865 8370 6895
rect 8310 6835 8370 6865
rect 8310 6805 8325 6835
rect 8355 6805 8370 6835
rect 8310 6770 8370 6805
rect 8310 6740 8325 6770
rect 8355 6740 8370 6770
rect 8310 6700 8370 6740
rect 8310 6670 8325 6700
rect 8355 6670 8370 6700
rect 8310 6630 8370 6670
rect 8310 6600 8325 6630
rect 8355 6600 8370 6630
rect 8310 6560 8370 6600
rect 8310 6530 8325 6560
rect 8355 6530 8370 6560
rect 8310 6495 8370 6530
rect 8310 6465 8325 6495
rect 8355 6465 8370 6495
rect 8310 6450 8370 6465
rect 8660 9635 8720 9650
rect 8660 9605 8675 9635
rect 8705 9605 8720 9635
rect 8660 9570 8720 9605
rect 8660 9540 8675 9570
rect 8705 9540 8720 9570
rect 8660 9500 8720 9540
rect 8660 9470 8675 9500
rect 8705 9470 8720 9500
rect 8660 9430 8720 9470
rect 8660 9400 8675 9430
rect 8705 9400 8720 9430
rect 8660 9360 8720 9400
rect 8660 9330 8675 9360
rect 8705 9330 8720 9360
rect 8660 9295 8720 9330
rect 8660 9265 8675 9295
rect 8705 9265 8720 9295
rect 8660 9235 8720 9265
rect 8660 9205 8675 9235
rect 8705 9205 8720 9235
rect 8660 9170 8720 9205
rect 8660 9140 8675 9170
rect 8705 9140 8720 9170
rect 8660 9100 8720 9140
rect 8660 9070 8675 9100
rect 8705 9070 8720 9100
rect 8660 9030 8720 9070
rect 8660 9000 8675 9030
rect 8705 9000 8720 9030
rect 8660 8960 8720 9000
rect 8660 8930 8675 8960
rect 8705 8930 8720 8960
rect 8660 8895 8720 8930
rect 8660 8865 8675 8895
rect 8705 8865 8720 8895
rect 8660 8835 8720 8865
rect 8660 8805 8675 8835
rect 8705 8805 8720 8835
rect 8660 8770 8720 8805
rect 8660 8740 8675 8770
rect 8705 8740 8720 8770
rect 8660 8700 8720 8740
rect 8660 8670 8675 8700
rect 8705 8670 8720 8700
rect 8660 8630 8720 8670
rect 8660 8600 8675 8630
rect 8705 8600 8720 8630
rect 8660 8560 8720 8600
rect 8660 8530 8675 8560
rect 8705 8530 8720 8560
rect 8660 8495 8720 8530
rect 8660 8465 8675 8495
rect 8705 8465 8720 8495
rect 8660 8435 8720 8465
rect 8660 8405 8675 8435
rect 8705 8405 8720 8435
rect 8660 8370 8720 8405
rect 8660 8340 8675 8370
rect 8705 8340 8720 8370
rect 8660 8300 8720 8340
rect 8660 8270 8675 8300
rect 8705 8270 8720 8300
rect 8660 8230 8720 8270
rect 8660 8200 8675 8230
rect 8705 8200 8720 8230
rect 8660 8160 8720 8200
rect 8660 8130 8675 8160
rect 8705 8130 8720 8160
rect 8660 8095 8720 8130
rect 8660 8065 8675 8095
rect 8705 8065 8720 8095
rect 8660 8035 8720 8065
rect 8660 8005 8675 8035
rect 8705 8005 8720 8035
rect 8660 7970 8720 8005
rect 8660 7940 8675 7970
rect 8705 7940 8720 7970
rect 8660 7900 8720 7940
rect 8660 7870 8675 7900
rect 8705 7870 8720 7900
rect 8660 7830 8720 7870
rect 8660 7800 8675 7830
rect 8705 7800 8720 7830
rect 8660 7760 8720 7800
rect 8660 7730 8675 7760
rect 8705 7730 8720 7760
rect 8660 7695 8720 7730
rect 8660 7665 8675 7695
rect 8705 7665 8720 7695
rect 8660 7635 8720 7665
rect 8660 7605 8675 7635
rect 8705 7605 8720 7635
rect 8660 7570 8720 7605
rect 8660 7540 8675 7570
rect 8705 7540 8720 7570
rect 8660 7500 8720 7540
rect 8660 7470 8675 7500
rect 8705 7470 8720 7500
rect 8660 7430 8720 7470
rect 8660 7400 8675 7430
rect 8705 7400 8720 7430
rect 8660 7360 8720 7400
rect 8660 7330 8675 7360
rect 8705 7330 8720 7360
rect 8660 7295 8720 7330
rect 8660 7265 8675 7295
rect 8705 7265 8720 7295
rect 8660 7235 8720 7265
rect 8660 7205 8675 7235
rect 8705 7205 8720 7235
rect 8660 7170 8720 7205
rect 8660 7140 8675 7170
rect 8705 7140 8720 7170
rect 8660 7100 8720 7140
rect 8660 7070 8675 7100
rect 8705 7070 8720 7100
rect 8660 7030 8720 7070
rect 8660 7000 8675 7030
rect 8705 7000 8720 7030
rect 8660 6960 8720 7000
rect 8660 6930 8675 6960
rect 8705 6930 8720 6960
rect 8660 6895 8720 6930
rect 8660 6865 8675 6895
rect 8705 6865 8720 6895
rect 8660 6835 8720 6865
rect 8660 6805 8675 6835
rect 8705 6805 8720 6835
rect 8660 6770 8720 6805
rect 8660 6740 8675 6770
rect 8705 6740 8720 6770
rect 8660 6700 8720 6740
rect 8660 6670 8675 6700
rect 8705 6670 8720 6700
rect 8660 6630 8720 6670
rect 8660 6600 8675 6630
rect 8705 6600 8720 6630
rect 8660 6560 8720 6600
rect 8660 6530 8675 6560
rect 8705 6530 8720 6560
rect 8660 6495 8720 6530
rect 8660 6465 8675 6495
rect 8705 6465 8720 6495
rect 8660 6450 8720 6465
rect 9010 9635 9070 9650
rect 9010 9605 9025 9635
rect 9055 9605 9070 9635
rect 9010 9570 9070 9605
rect 9010 9540 9025 9570
rect 9055 9540 9070 9570
rect 9010 9500 9070 9540
rect 9010 9470 9025 9500
rect 9055 9470 9070 9500
rect 9010 9430 9070 9470
rect 9010 9400 9025 9430
rect 9055 9400 9070 9430
rect 9010 9360 9070 9400
rect 9010 9330 9025 9360
rect 9055 9330 9070 9360
rect 9010 9295 9070 9330
rect 9010 9265 9025 9295
rect 9055 9265 9070 9295
rect 9010 9235 9070 9265
rect 9010 9205 9025 9235
rect 9055 9205 9070 9235
rect 9010 9170 9070 9205
rect 9010 9140 9025 9170
rect 9055 9140 9070 9170
rect 9010 9100 9070 9140
rect 9010 9070 9025 9100
rect 9055 9070 9070 9100
rect 9010 9030 9070 9070
rect 9010 9000 9025 9030
rect 9055 9000 9070 9030
rect 9010 8960 9070 9000
rect 9010 8930 9025 8960
rect 9055 8930 9070 8960
rect 9010 8895 9070 8930
rect 9010 8865 9025 8895
rect 9055 8865 9070 8895
rect 9010 8835 9070 8865
rect 9010 8805 9025 8835
rect 9055 8805 9070 8835
rect 9010 8770 9070 8805
rect 9010 8740 9025 8770
rect 9055 8740 9070 8770
rect 9010 8700 9070 8740
rect 9010 8670 9025 8700
rect 9055 8670 9070 8700
rect 9010 8630 9070 8670
rect 9010 8600 9025 8630
rect 9055 8600 9070 8630
rect 9010 8560 9070 8600
rect 9010 8530 9025 8560
rect 9055 8530 9070 8560
rect 9010 8495 9070 8530
rect 9010 8465 9025 8495
rect 9055 8465 9070 8495
rect 9010 8435 9070 8465
rect 9010 8405 9025 8435
rect 9055 8405 9070 8435
rect 9010 8370 9070 8405
rect 9010 8340 9025 8370
rect 9055 8340 9070 8370
rect 9010 8300 9070 8340
rect 9010 8270 9025 8300
rect 9055 8270 9070 8300
rect 9010 8230 9070 8270
rect 9010 8200 9025 8230
rect 9055 8200 9070 8230
rect 9010 8160 9070 8200
rect 9010 8130 9025 8160
rect 9055 8130 9070 8160
rect 9010 8095 9070 8130
rect 9010 8065 9025 8095
rect 9055 8065 9070 8095
rect 9010 8035 9070 8065
rect 9010 8005 9025 8035
rect 9055 8005 9070 8035
rect 9010 7970 9070 8005
rect 9010 7940 9025 7970
rect 9055 7940 9070 7970
rect 9010 7900 9070 7940
rect 9010 7870 9025 7900
rect 9055 7870 9070 7900
rect 9010 7830 9070 7870
rect 9010 7800 9025 7830
rect 9055 7800 9070 7830
rect 9010 7760 9070 7800
rect 9010 7730 9025 7760
rect 9055 7730 9070 7760
rect 9010 7695 9070 7730
rect 9010 7665 9025 7695
rect 9055 7665 9070 7695
rect 9010 7635 9070 7665
rect 9010 7605 9025 7635
rect 9055 7605 9070 7635
rect 9010 7570 9070 7605
rect 9010 7540 9025 7570
rect 9055 7540 9070 7570
rect 9010 7500 9070 7540
rect 9010 7470 9025 7500
rect 9055 7470 9070 7500
rect 9010 7430 9070 7470
rect 9010 7400 9025 7430
rect 9055 7400 9070 7430
rect 9010 7360 9070 7400
rect 9010 7330 9025 7360
rect 9055 7330 9070 7360
rect 9010 7295 9070 7330
rect 9010 7265 9025 7295
rect 9055 7265 9070 7295
rect 9010 7235 9070 7265
rect 9010 7205 9025 7235
rect 9055 7205 9070 7235
rect 9010 7170 9070 7205
rect 9010 7140 9025 7170
rect 9055 7140 9070 7170
rect 9010 7100 9070 7140
rect 9010 7070 9025 7100
rect 9055 7070 9070 7100
rect 9010 7030 9070 7070
rect 9010 7000 9025 7030
rect 9055 7000 9070 7030
rect 9010 6960 9070 7000
rect 9010 6930 9025 6960
rect 9055 6930 9070 6960
rect 9010 6895 9070 6930
rect 9010 6865 9025 6895
rect 9055 6865 9070 6895
rect 9010 6835 9070 6865
rect 9010 6805 9025 6835
rect 9055 6805 9070 6835
rect 9010 6770 9070 6805
rect 9010 6740 9025 6770
rect 9055 6740 9070 6770
rect 9010 6700 9070 6740
rect 9010 6670 9025 6700
rect 9055 6670 9070 6700
rect 9010 6630 9070 6670
rect 9010 6600 9025 6630
rect 9055 6600 9070 6630
rect 9010 6560 9070 6600
rect 9010 6530 9025 6560
rect 9055 6530 9070 6560
rect 9010 6495 9070 6530
rect 9010 6465 9025 6495
rect 9055 6465 9070 6495
rect 9010 6450 9070 6465
rect 2045 6430 2515 6435
rect 2045 6400 2050 6430
rect 2080 6400 2480 6430
rect 2510 6400 2515 6430
rect 2045 6395 2515 6400
rect 2845 6430 2885 6435
rect 2845 6400 2850 6430
rect 2880 6425 2885 6430
rect 3380 6430 3420 6435
rect 3380 6425 3385 6430
rect 2880 6405 3385 6425
rect 2880 6400 2885 6405
rect 2845 6395 2885 6400
rect 3380 6400 3385 6405
rect 3415 6400 3420 6430
rect 3380 6395 3420 6400
rect 5470 6430 5510 6435
rect 5470 6400 5475 6430
rect 5505 6425 5510 6430
rect 6145 6430 6185 6435
rect 6145 6425 6150 6430
rect 5505 6405 6150 6425
rect 5505 6400 5510 6405
rect 5470 6395 5510 6400
rect 6145 6400 6150 6405
rect 6180 6400 6185 6430
rect 6145 6395 6185 6400
rect 6465 6430 6935 6435
rect 6465 6400 6470 6430
rect 6500 6400 6900 6430
rect 6930 6400 6935 6430
rect 6465 6395 6935 6400
rect 2000 6375 2040 6380
rect 2000 6345 2005 6375
rect 2035 6370 2040 6375
rect 3630 6375 3670 6380
rect 3630 6370 3635 6375
rect 2035 6350 3635 6370
rect 2035 6345 2040 6350
rect 2000 6340 2040 6345
rect 3630 6345 3635 6350
rect 3665 6345 3670 6375
rect 3630 6340 3670 6345
rect 5310 6375 5350 6380
rect 5310 6345 5315 6375
rect 5345 6370 5350 6375
rect 6940 6375 6980 6380
rect 6940 6370 6945 6375
rect 5345 6350 6945 6370
rect 5345 6345 5350 6350
rect 5310 6340 5350 6345
rect 6940 6345 6945 6350
rect 6975 6345 6980 6375
rect 6940 6340 6980 6345
rect 2715 6330 2755 6335
rect 2715 6300 2720 6330
rect 2750 6325 2755 6330
rect 3075 6330 3115 6335
rect 3075 6325 3080 6330
rect 2750 6305 3080 6325
rect 2750 6300 2755 6305
rect 2715 6295 2755 6300
rect 3075 6300 3080 6305
rect 3110 6300 3115 6330
rect 3075 6295 3115 6300
rect 3290 6315 4510 6320
rect 3290 6285 3295 6315
rect 3325 6285 4475 6315
rect 4505 6285 4510 6315
rect 3290 6280 4510 6285
rect 3435 6260 5560 6265
rect 3435 6230 3440 6260
rect 3470 6230 4475 6260
rect 4505 6230 5525 6260
rect 5555 6230 5560 6260
rect 3435 6225 5560 6230
rect 1280 6205 7700 6210
rect 1280 6175 1285 6205
rect 1315 6175 1325 6205
rect 1355 6175 1365 6205
rect 1395 6175 4310 6205
rect 4340 6175 4420 6205
rect 4450 6175 4530 6205
rect 4560 6175 4640 6205
rect 4670 6175 7585 6205
rect 7615 6175 7625 6205
rect 7655 6175 7665 6205
rect 7695 6175 7700 6205
rect 1280 6165 7700 6175
rect 1280 6135 1285 6165
rect 1315 6135 1325 6165
rect 1355 6135 1365 6165
rect 1395 6135 4310 6165
rect 4340 6135 4420 6165
rect 4450 6135 4530 6165
rect 4560 6135 4640 6165
rect 4670 6135 7585 6165
rect 7615 6135 7625 6165
rect 7655 6135 7665 6165
rect 7695 6135 7700 6165
rect 1280 6125 7700 6135
rect 1280 6095 1285 6125
rect 1315 6095 1325 6125
rect 1355 6095 1365 6125
rect 1395 6095 4310 6125
rect 4340 6095 4420 6125
rect 4450 6095 4530 6125
rect 4560 6095 4640 6125
rect 4670 6095 7585 6125
rect 7615 6095 7625 6125
rect 7655 6095 7665 6125
rect 7695 6095 7700 6125
rect 1280 6090 7700 6095
rect 5575 5435 5605 5440
rect 6220 5435 6260 5440
rect 6220 5430 6225 5435
rect 5605 5410 6225 5430
rect 5575 5400 5605 5405
rect 6220 5405 6225 5410
rect 6255 5405 6260 5435
rect 6220 5400 6260 5405
rect 3075 5090 3115 5095
rect 3075 5060 3080 5090
rect 3110 5060 3115 5090
rect 3075 5055 3115 5060
rect 5575 4440 5605 4445
rect 5575 4405 5605 4410
rect 5475 3865 5505 3870
rect 4720 3840 5475 3860
rect 5475 3830 5505 3835
rect 3380 3805 3420 3810
rect 3380 3775 3385 3805
rect 3415 3800 3420 3805
rect 3415 3780 3955 3800
rect 3415 3775 3420 3780
rect 3380 3770 3420 3775
rect 3435 3125 5560 3130
rect 3435 3095 3440 3125
rect 3470 3095 4475 3125
rect 4505 3095 5525 3125
rect 5555 3095 5560 3125
rect 3435 3090 5560 3095
rect 4470 3015 4510 3020
rect 4470 2985 4475 3015
rect 4505 2985 4510 3015
rect 4470 2980 4510 2985
rect 2045 2315 2085 2320
rect 2045 2285 2050 2315
rect 2080 2310 2085 2315
rect 2120 2315 2160 2320
rect 2120 2310 2125 2315
rect 2080 2290 2125 2310
rect 2080 2285 2085 2290
rect 2045 2280 2085 2285
rect 2120 2285 2125 2290
rect 2155 2285 2160 2315
rect 2120 2280 2160 2285
rect 6820 2315 6860 2320
rect 6820 2285 6825 2315
rect 6855 2310 6860 2315
rect 6895 2315 6935 2320
rect 6895 2310 6900 2315
rect 6855 2290 6900 2310
rect 6855 2285 6860 2290
rect 6820 2280 6860 2285
rect 6895 2285 6900 2290
rect 6930 2285 6935 2315
rect 6895 2280 6935 2285
rect 2000 2260 2040 2265
rect 2000 2230 2005 2260
rect 2035 2255 2040 2260
rect 2075 2260 2115 2265
rect 2075 2255 2080 2260
rect 2035 2235 2080 2255
rect 2035 2230 2040 2235
rect 2000 2225 2040 2230
rect 2075 2230 2080 2235
rect 2110 2230 2115 2260
rect 2075 2225 2115 2230
rect 6865 2260 6905 2265
rect 6865 2230 6870 2260
rect 6900 2255 6905 2260
rect 6940 2260 6980 2265
rect 6940 2255 6945 2260
rect 6900 2235 6945 2255
rect 6900 2230 6905 2235
rect 6865 2225 6905 2230
rect 6940 2230 6945 2235
rect 6975 2230 6980 2260
rect 6940 2225 6980 2230
rect 3605 2080 3625 2100
rect 5355 2080 5375 2100
rect 1280 1160 7700 1165
rect 1280 1130 1285 1160
rect 1315 1130 1325 1160
rect 1355 1130 1365 1160
rect 1395 1130 4420 1160
rect 4450 1130 4530 1160
rect 4560 1130 7585 1160
rect 7615 1130 7625 1160
rect 7655 1130 7665 1160
rect 7695 1130 7700 1160
rect 1280 1120 7700 1130
rect 1280 1090 1285 1120
rect 1315 1090 1325 1120
rect 1355 1090 1365 1120
rect 1395 1090 4420 1120
rect 4450 1090 4530 1120
rect 4560 1090 7585 1120
rect 7615 1090 7625 1120
rect 7655 1090 7665 1120
rect 7695 1090 7700 1120
rect 1280 1080 7700 1090
rect 1280 1050 1285 1080
rect 1315 1050 1325 1080
rect 1355 1050 1365 1080
rect 1395 1050 4420 1080
rect 4450 1050 4530 1080
rect 4560 1050 7585 1080
rect 7615 1050 7625 1080
rect 7655 1050 7665 1080
rect 7695 1050 7700 1080
rect 1280 1045 7700 1050
rect 2175 855 2195 875
rect 6785 855 6805 875
rect -90 -1305 -30 -1290
rect -90 -1335 -75 -1305
rect -45 -1335 -30 -1305
rect -90 -1370 -30 -1335
rect -90 -1400 -75 -1370
rect -45 -1400 -30 -1370
rect -90 -1440 -30 -1400
rect -90 -1470 -75 -1440
rect -45 -1470 -30 -1440
rect -90 -1510 -30 -1470
rect -90 -1540 -75 -1510
rect -45 -1540 -30 -1510
rect -90 -1580 -30 -1540
rect -90 -1610 -75 -1580
rect -45 -1610 -30 -1580
rect -90 -1645 -30 -1610
rect -90 -1675 -75 -1645
rect -45 -1675 -30 -1645
rect -90 -1705 -30 -1675
rect -90 -1735 -75 -1705
rect -45 -1735 -30 -1705
rect -90 -1770 -30 -1735
rect -90 -1800 -75 -1770
rect -45 -1800 -30 -1770
rect -90 -1840 -30 -1800
rect -90 -1870 -75 -1840
rect -45 -1870 -30 -1840
rect -90 -1910 -30 -1870
rect -90 -1940 -75 -1910
rect -45 -1940 -30 -1910
rect -90 -1980 -30 -1940
rect -90 -2010 -75 -1980
rect -45 -2010 -30 -1980
rect -90 -2045 -30 -2010
rect -90 -2075 -75 -2045
rect -45 -2075 -30 -2045
rect -90 -2105 -30 -2075
rect -90 -2135 -75 -2105
rect -45 -2135 -30 -2105
rect -90 -2170 -30 -2135
rect -90 -2200 -75 -2170
rect -45 -2200 -30 -2170
rect -90 -2240 -30 -2200
rect -90 -2270 -75 -2240
rect -45 -2270 -30 -2240
rect -90 -2310 -30 -2270
rect -90 -2340 -75 -2310
rect -45 -2340 -30 -2310
rect -90 -2380 -30 -2340
rect -90 -2410 -75 -2380
rect -45 -2410 -30 -2380
rect -90 -2445 -30 -2410
rect -90 -2475 -75 -2445
rect -45 -2475 -30 -2445
rect -90 -2505 -30 -2475
rect -90 -2535 -75 -2505
rect -45 -2535 -30 -2505
rect -90 -2570 -30 -2535
rect -90 -2600 -75 -2570
rect -45 -2600 -30 -2570
rect -90 -2640 -30 -2600
rect -90 -2670 -75 -2640
rect -45 -2670 -30 -2640
rect -90 -2710 -30 -2670
rect -90 -2740 -75 -2710
rect -45 -2740 -30 -2710
rect -90 -2780 -30 -2740
rect -90 -2810 -75 -2780
rect -45 -2810 -30 -2780
rect -90 -2845 -30 -2810
rect -90 -2875 -75 -2845
rect -45 -2875 -30 -2845
rect -90 -2890 -30 -2875
rect 260 -1305 320 -1290
rect 260 -1335 275 -1305
rect 305 -1335 320 -1305
rect 260 -1370 320 -1335
rect 260 -1400 275 -1370
rect 305 -1400 320 -1370
rect 260 -1440 320 -1400
rect 260 -1470 275 -1440
rect 305 -1470 320 -1440
rect 260 -1510 320 -1470
rect 260 -1540 275 -1510
rect 305 -1540 320 -1510
rect 260 -1580 320 -1540
rect 260 -1610 275 -1580
rect 305 -1610 320 -1580
rect 260 -1645 320 -1610
rect 260 -1675 275 -1645
rect 305 -1675 320 -1645
rect 260 -1705 320 -1675
rect 260 -1735 275 -1705
rect 305 -1735 320 -1705
rect 260 -1770 320 -1735
rect 260 -1800 275 -1770
rect 305 -1800 320 -1770
rect 260 -1840 320 -1800
rect 260 -1870 275 -1840
rect 305 -1870 320 -1840
rect 260 -1910 320 -1870
rect 260 -1940 275 -1910
rect 305 -1940 320 -1910
rect 260 -1980 320 -1940
rect 260 -2010 275 -1980
rect 305 -2010 320 -1980
rect 260 -2045 320 -2010
rect 260 -2075 275 -2045
rect 305 -2075 320 -2045
rect 260 -2105 320 -2075
rect 260 -2135 275 -2105
rect 305 -2135 320 -2105
rect 260 -2170 320 -2135
rect 260 -2200 275 -2170
rect 305 -2200 320 -2170
rect 260 -2240 320 -2200
rect 260 -2270 275 -2240
rect 305 -2270 320 -2240
rect 260 -2310 320 -2270
rect 260 -2340 275 -2310
rect 305 -2340 320 -2310
rect 260 -2380 320 -2340
rect 260 -2410 275 -2380
rect 305 -2410 320 -2380
rect 260 -2445 320 -2410
rect 260 -2475 275 -2445
rect 305 -2475 320 -2445
rect 260 -2505 320 -2475
rect 260 -2535 275 -2505
rect 305 -2535 320 -2505
rect 260 -2570 320 -2535
rect 260 -2600 275 -2570
rect 305 -2600 320 -2570
rect 260 -2640 320 -2600
rect 260 -2670 275 -2640
rect 305 -2670 320 -2640
rect 260 -2710 320 -2670
rect 260 -2740 275 -2710
rect 305 -2740 320 -2710
rect 260 -2780 320 -2740
rect 260 -2810 275 -2780
rect 305 -2810 320 -2780
rect 260 -2845 320 -2810
rect 260 -2875 275 -2845
rect 305 -2875 320 -2845
rect 260 -2890 320 -2875
rect 610 -1305 670 -1290
rect 610 -1335 625 -1305
rect 655 -1335 670 -1305
rect 610 -1370 670 -1335
rect 610 -1400 625 -1370
rect 655 -1400 670 -1370
rect 610 -1440 670 -1400
rect 610 -1470 625 -1440
rect 655 -1470 670 -1440
rect 610 -1510 670 -1470
rect 610 -1540 625 -1510
rect 655 -1540 670 -1510
rect 610 -1580 670 -1540
rect 610 -1610 625 -1580
rect 655 -1610 670 -1580
rect 610 -1645 670 -1610
rect 610 -1675 625 -1645
rect 655 -1675 670 -1645
rect 610 -1705 670 -1675
rect 610 -1735 625 -1705
rect 655 -1735 670 -1705
rect 610 -1770 670 -1735
rect 610 -1800 625 -1770
rect 655 -1800 670 -1770
rect 610 -1840 670 -1800
rect 610 -1870 625 -1840
rect 655 -1870 670 -1840
rect 610 -1910 670 -1870
rect 610 -1940 625 -1910
rect 655 -1940 670 -1910
rect 610 -1980 670 -1940
rect 610 -2010 625 -1980
rect 655 -2010 670 -1980
rect 610 -2045 670 -2010
rect 610 -2075 625 -2045
rect 655 -2075 670 -2045
rect 610 -2105 670 -2075
rect 610 -2135 625 -2105
rect 655 -2135 670 -2105
rect 610 -2170 670 -2135
rect 610 -2200 625 -2170
rect 655 -2200 670 -2170
rect 610 -2240 670 -2200
rect 610 -2270 625 -2240
rect 655 -2270 670 -2240
rect 610 -2310 670 -2270
rect 610 -2340 625 -2310
rect 655 -2340 670 -2310
rect 610 -2380 670 -2340
rect 610 -2410 625 -2380
rect 655 -2410 670 -2380
rect 610 -2445 670 -2410
rect 610 -2475 625 -2445
rect 655 -2475 670 -2445
rect 610 -2505 670 -2475
rect 610 -2535 625 -2505
rect 655 -2535 670 -2505
rect 610 -2570 670 -2535
rect 610 -2600 625 -2570
rect 655 -2600 670 -2570
rect 610 -2640 670 -2600
rect 610 -2670 625 -2640
rect 655 -2670 670 -2640
rect 610 -2710 670 -2670
rect 610 -2740 625 -2710
rect 655 -2740 670 -2710
rect 610 -2780 670 -2740
rect 610 -2810 625 -2780
rect 655 -2810 670 -2780
rect 610 -2845 670 -2810
rect 610 -2875 625 -2845
rect 655 -2875 670 -2845
rect 610 -2890 670 -2875
rect 960 -1305 1020 -1290
rect 960 -1335 975 -1305
rect 1005 -1335 1020 -1305
rect 960 -1370 1020 -1335
rect 960 -1400 975 -1370
rect 1005 -1400 1020 -1370
rect 960 -1440 1020 -1400
rect 960 -1470 975 -1440
rect 1005 -1470 1020 -1440
rect 960 -1510 1020 -1470
rect 960 -1540 975 -1510
rect 1005 -1540 1020 -1510
rect 960 -1580 1020 -1540
rect 960 -1610 975 -1580
rect 1005 -1610 1020 -1580
rect 960 -1645 1020 -1610
rect 960 -1675 975 -1645
rect 1005 -1675 1020 -1645
rect 960 -1705 1020 -1675
rect 960 -1735 975 -1705
rect 1005 -1735 1020 -1705
rect 960 -1770 1020 -1735
rect 960 -1800 975 -1770
rect 1005 -1800 1020 -1770
rect 960 -1840 1020 -1800
rect 960 -1870 975 -1840
rect 1005 -1870 1020 -1840
rect 960 -1910 1020 -1870
rect 960 -1940 975 -1910
rect 1005 -1940 1020 -1910
rect 960 -1980 1020 -1940
rect 960 -2010 975 -1980
rect 1005 -2010 1020 -1980
rect 960 -2045 1020 -2010
rect 960 -2075 975 -2045
rect 1005 -2075 1020 -2045
rect 960 -2105 1020 -2075
rect 960 -2135 975 -2105
rect 1005 -2135 1020 -2105
rect 960 -2170 1020 -2135
rect 960 -2200 975 -2170
rect 1005 -2200 1020 -2170
rect 960 -2240 1020 -2200
rect 960 -2270 975 -2240
rect 1005 -2270 1020 -2240
rect 960 -2310 1020 -2270
rect 960 -2340 975 -2310
rect 1005 -2340 1020 -2310
rect 960 -2380 1020 -2340
rect 960 -2410 975 -2380
rect 1005 -2410 1020 -2380
rect 960 -2445 1020 -2410
rect 960 -2475 975 -2445
rect 1005 -2475 1020 -2445
rect 960 -2505 1020 -2475
rect 960 -2535 975 -2505
rect 1005 -2535 1020 -2505
rect 960 -2570 1020 -2535
rect 960 -2600 975 -2570
rect 1005 -2600 1020 -2570
rect 960 -2640 1020 -2600
rect 960 -2670 975 -2640
rect 1005 -2670 1020 -2640
rect 960 -2710 1020 -2670
rect 960 -2740 975 -2710
rect 1005 -2740 1020 -2710
rect 960 -2780 1020 -2740
rect 960 -2810 975 -2780
rect 1005 -2810 1020 -2780
rect 960 -2845 1020 -2810
rect 960 -2875 975 -2845
rect 1005 -2875 1020 -2845
rect 960 -2890 1020 -2875
rect 1310 -1305 1370 -1290
rect 1310 -1335 1325 -1305
rect 1355 -1335 1370 -1305
rect 1310 -1370 1370 -1335
rect 1310 -1400 1325 -1370
rect 1355 -1400 1370 -1370
rect 1310 -1440 1370 -1400
rect 1310 -1470 1325 -1440
rect 1355 -1470 1370 -1440
rect 1310 -1510 1370 -1470
rect 1310 -1540 1325 -1510
rect 1355 -1540 1370 -1510
rect 1310 -1580 1370 -1540
rect 1310 -1610 1325 -1580
rect 1355 -1610 1370 -1580
rect 1310 -1645 1370 -1610
rect 1310 -1675 1325 -1645
rect 1355 -1675 1370 -1645
rect 1310 -1705 1370 -1675
rect 1310 -1735 1325 -1705
rect 1355 -1735 1370 -1705
rect 1310 -1770 1370 -1735
rect 1310 -1800 1325 -1770
rect 1355 -1800 1370 -1770
rect 1310 -1840 1370 -1800
rect 1310 -1870 1325 -1840
rect 1355 -1870 1370 -1840
rect 1310 -1910 1370 -1870
rect 1310 -1940 1325 -1910
rect 1355 -1940 1370 -1910
rect 1310 -1980 1370 -1940
rect 1310 -2010 1325 -1980
rect 1355 -2010 1370 -1980
rect 1310 -2045 1370 -2010
rect 1310 -2075 1325 -2045
rect 1355 -2075 1370 -2045
rect 1310 -2105 1370 -2075
rect 1310 -2135 1325 -2105
rect 1355 -2135 1370 -2105
rect 1310 -2170 1370 -2135
rect 1310 -2200 1325 -2170
rect 1355 -2200 1370 -2170
rect 1310 -2240 1370 -2200
rect 1310 -2270 1325 -2240
rect 1355 -2270 1370 -2240
rect 1310 -2310 1370 -2270
rect 1310 -2340 1325 -2310
rect 1355 -2340 1370 -2310
rect 1310 -2380 1370 -2340
rect 1310 -2410 1325 -2380
rect 1355 -2410 1370 -2380
rect 1310 -2445 1370 -2410
rect 1310 -2475 1325 -2445
rect 1355 -2475 1370 -2445
rect 1310 -2505 1370 -2475
rect 1310 -2535 1325 -2505
rect 1355 -2535 1370 -2505
rect 1310 -2570 1370 -2535
rect 1310 -2600 1325 -2570
rect 1355 -2600 1370 -2570
rect 1310 -2640 1370 -2600
rect 1310 -2670 1325 -2640
rect 1355 -2670 1370 -2640
rect 1310 -2710 1370 -2670
rect 1310 -2740 1325 -2710
rect 1355 -2740 1370 -2710
rect 1310 -2780 1370 -2740
rect 1310 -2810 1325 -2780
rect 1355 -2810 1370 -2780
rect 1310 -2845 1370 -2810
rect 1310 -2875 1325 -2845
rect 1355 -2875 1370 -2845
rect 1310 -2890 1370 -2875
rect 1660 -1305 1720 -1290
rect 1660 -1335 1675 -1305
rect 1705 -1335 1720 -1305
rect 1660 -1370 1720 -1335
rect 1660 -1400 1675 -1370
rect 1705 -1400 1720 -1370
rect 1660 -1440 1720 -1400
rect 1660 -1470 1675 -1440
rect 1705 -1470 1720 -1440
rect 1660 -1510 1720 -1470
rect 1660 -1540 1675 -1510
rect 1705 -1540 1720 -1510
rect 1660 -1580 1720 -1540
rect 1660 -1610 1675 -1580
rect 1705 -1610 1720 -1580
rect 1660 -1645 1720 -1610
rect 1660 -1675 1675 -1645
rect 1705 -1675 1720 -1645
rect 1660 -1705 1720 -1675
rect 1660 -1735 1675 -1705
rect 1705 -1735 1720 -1705
rect 1660 -1770 1720 -1735
rect 1660 -1800 1675 -1770
rect 1705 -1800 1720 -1770
rect 1660 -1840 1720 -1800
rect 1660 -1870 1675 -1840
rect 1705 -1870 1720 -1840
rect 1660 -1910 1720 -1870
rect 1660 -1940 1675 -1910
rect 1705 -1940 1720 -1910
rect 1660 -1980 1720 -1940
rect 1660 -2010 1675 -1980
rect 1705 -2010 1720 -1980
rect 1660 -2045 1720 -2010
rect 1660 -2075 1675 -2045
rect 1705 -2075 1720 -2045
rect 1660 -2105 1720 -2075
rect 1660 -2135 1675 -2105
rect 1705 -2135 1720 -2105
rect 1660 -2170 1720 -2135
rect 1660 -2200 1675 -2170
rect 1705 -2200 1720 -2170
rect 1660 -2240 1720 -2200
rect 1660 -2270 1675 -2240
rect 1705 -2270 1720 -2240
rect 1660 -2310 1720 -2270
rect 1660 -2340 1675 -2310
rect 1705 -2340 1720 -2310
rect 1660 -2380 1720 -2340
rect 1660 -2410 1675 -2380
rect 1705 -2410 1720 -2380
rect 1660 -2445 1720 -2410
rect 1660 -2475 1675 -2445
rect 1705 -2475 1720 -2445
rect 1660 -2505 1720 -2475
rect 1660 -2535 1675 -2505
rect 1705 -2535 1720 -2505
rect 1660 -2570 1720 -2535
rect 1660 -2600 1675 -2570
rect 1705 -2600 1720 -2570
rect 1660 -2640 1720 -2600
rect 1660 -2670 1675 -2640
rect 1705 -2670 1720 -2640
rect 1660 -2710 1720 -2670
rect 1660 -2740 1675 -2710
rect 1705 -2740 1720 -2710
rect 1660 -2780 1720 -2740
rect 1660 -2810 1675 -2780
rect 1705 -2810 1720 -2780
rect 1660 -2845 1720 -2810
rect 1660 -2875 1675 -2845
rect 1705 -2875 1720 -2845
rect 1660 -2890 1720 -2875
rect 2010 -1305 2070 -1290
rect 2010 -1335 2025 -1305
rect 2055 -1335 2070 -1305
rect 2010 -1370 2070 -1335
rect 2010 -1400 2025 -1370
rect 2055 -1400 2070 -1370
rect 2010 -1440 2070 -1400
rect 2010 -1470 2025 -1440
rect 2055 -1470 2070 -1440
rect 2010 -1510 2070 -1470
rect 2010 -1540 2025 -1510
rect 2055 -1540 2070 -1510
rect 2010 -1580 2070 -1540
rect 2010 -1610 2025 -1580
rect 2055 -1610 2070 -1580
rect 2010 -1645 2070 -1610
rect 2010 -1675 2025 -1645
rect 2055 -1675 2070 -1645
rect 2010 -1705 2070 -1675
rect 2010 -1735 2025 -1705
rect 2055 -1735 2070 -1705
rect 2010 -1770 2070 -1735
rect 2010 -1800 2025 -1770
rect 2055 -1800 2070 -1770
rect 2010 -1840 2070 -1800
rect 2010 -1870 2025 -1840
rect 2055 -1870 2070 -1840
rect 2010 -1910 2070 -1870
rect 2010 -1940 2025 -1910
rect 2055 -1940 2070 -1910
rect 2010 -1980 2070 -1940
rect 2010 -2010 2025 -1980
rect 2055 -2010 2070 -1980
rect 2010 -2045 2070 -2010
rect 2010 -2075 2025 -2045
rect 2055 -2075 2070 -2045
rect 2010 -2105 2070 -2075
rect 2010 -2135 2025 -2105
rect 2055 -2135 2070 -2105
rect 2010 -2170 2070 -2135
rect 2010 -2200 2025 -2170
rect 2055 -2200 2070 -2170
rect 2010 -2240 2070 -2200
rect 2010 -2270 2025 -2240
rect 2055 -2270 2070 -2240
rect 2010 -2310 2070 -2270
rect 2010 -2340 2025 -2310
rect 2055 -2340 2070 -2310
rect 2010 -2380 2070 -2340
rect 2010 -2410 2025 -2380
rect 2055 -2410 2070 -2380
rect 2010 -2445 2070 -2410
rect 2010 -2475 2025 -2445
rect 2055 -2475 2070 -2445
rect 2010 -2505 2070 -2475
rect 2010 -2535 2025 -2505
rect 2055 -2535 2070 -2505
rect 2010 -2570 2070 -2535
rect 2010 -2600 2025 -2570
rect 2055 -2600 2070 -2570
rect 2010 -2640 2070 -2600
rect 2010 -2670 2025 -2640
rect 2055 -2670 2070 -2640
rect 2010 -2710 2070 -2670
rect 2010 -2740 2025 -2710
rect 2055 -2740 2070 -2710
rect 2010 -2780 2070 -2740
rect 2010 -2810 2025 -2780
rect 2055 -2810 2070 -2780
rect 2010 -2845 2070 -2810
rect 2010 -2875 2025 -2845
rect 2055 -2875 2070 -2845
rect 2010 -2890 2070 -2875
rect 2360 -1305 2420 -1290
rect 2360 -1335 2375 -1305
rect 2405 -1335 2420 -1305
rect 2360 -1370 2420 -1335
rect 2360 -1400 2375 -1370
rect 2405 -1400 2420 -1370
rect 2360 -1440 2420 -1400
rect 2360 -1470 2375 -1440
rect 2405 -1470 2420 -1440
rect 2360 -1510 2420 -1470
rect 2360 -1540 2375 -1510
rect 2405 -1540 2420 -1510
rect 2360 -1580 2420 -1540
rect 2360 -1610 2375 -1580
rect 2405 -1610 2420 -1580
rect 2360 -1645 2420 -1610
rect 2360 -1675 2375 -1645
rect 2405 -1675 2420 -1645
rect 2360 -1705 2420 -1675
rect 2360 -1735 2375 -1705
rect 2405 -1735 2420 -1705
rect 2360 -1770 2420 -1735
rect 2360 -1800 2375 -1770
rect 2405 -1800 2420 -1770
rect 2360 -1840 2420 -1800
rect 2360 -1870 2375 -1840
rect 2405 -1870 2420 -1840
rect 2360 -1910 2420 -1870
rect 2360 -1940 2375 -1910
rect 2405 -1940 2420 -1910
rect 2360 -1980 2420 -1940
rect 2360 -2010 2375 -1980
rect 2405 -2010 2420 -1980
rect 2360 -2045 2420 -2010
rect 2360 -2075 2375 -2045
rect 2405 -2075 2420 -2045
rect 2360 -2105 2420 -2075
rect 2360 -2135 2375 -2105
rect 2405 -2135 2420 -2105
rect 2360 -2170 2420 -2135
rect 2360 -2200 2375 -2170
rect 2405 -2200 2420 -2170
rect 2360 -2240 2420 -2200
rect 2360 -2270 2375 -2240
rect 2405 -2270 2420 -2240
rect 2360 -2310 2420 -2270
rect 2360 -2340 2375 -2310
rect 2405 -2340 2420 -2310
rect 2360 -2380 2420 -2340
rect 2360 -2410 2375 -2380
rect 2405 -2410 2420 -2380
rect 2360 -2445 2420 -2410
rect 2360 -2475 2375 -2445
rect 2405 -2475 2420 -2445
rect 2360 -2505 2420 -2475
rect 2360 -2535 2375 -2505
rect 2405 -2535 2420 -2505
rect 2360 -2570 2420 -2535
rect 2360 -2600 2375 -2570
rect 2405 -2600 2420 -2570
rect 2360 -2640 2420 -2600
rect 2360 -2670 2375 -2640
rect 2405 -2670 2420 -2640
rect 2360 -2710 2420 -2670
rect 2360 -2740 2375 -2710
rect 2405 -2740 2420 -2710
rect 2360 -2780 2420 -2740
rect 2360 -2810 2375 -2780
rect 2405 -2810 2420 -2780
rect 2360 -2845 2420 -2810
rect 2360 -2875 2375 -2845
rect 2405 -2875 2420 -2845
rect 2360 -2890 2420 -2875
rect 2710 -1305 2770 -1290
rect 2710 -1335 2725 -1305
rect 2755 -1335 2770 -1305
rect 2710 -1370 2770 -1335
rect 2710 -1400 2725 -1370
rect 2755 -1400 2770 -1370
rect 2710 -1440 2770 -1400
rect 2710 -1470 2725 -1440
rect 2755 -1470 2770 -1440
rect 2710 -1510 2770 -1470
rect 2710 -1540 2725 -1510
rect 2755 -1540 2770 -1510
rect 2710 -1580 2770 -1540
rect 2710 -1610 2725 -1580
rect 2755 -1610 2770 -1580
rect 2710 -1645 2770 -1610
rect 2710 -1675 2725 -1645
rect 2755 -1675 2770 -1645
rect 2710 -1705 2770 -1675
rect 2710 -1735 2725 -1705
rect 2755 -1735 2770 -1705
rect 2710 -1770 2770 -1735
rect 2710 -1800 2725 -1770
rect 2755 -1800 2770 -1770
rect 2710 -1840 2770 -1800
rect 2710 -1870 2725 -1840
rect 2755 -1870 2770 -1840
rect 2710 -1910 2770 -1870
rect 2710 -1940 2725 -1910
rect 2755 -1940 2770 -1910
rect 2710 -1980 2770 -1940
rect 2710 -2010 2725 -1980
rect 2755 -2010 2770 -1980
rect 2710 -2045 2770 -2010
rect 2710 -2075 2725 -2045
rect 2755 -2075 2770 -2045
rect 2710 -2105 2770 -2075
rect 2710 -2135 2725 -2105
rect 2755 -2135 2770 -2105
rect 2710 -2170 2770 -2135
rect 2710 -2200 2725 -2170
rect 2755 -2200 2770 -2170
rect 2710 -2240 2770 -2200
rect 2710 -2270 2725 -2240
rect 2755 -2270 2770 -2240
rect 2710 -2310 2770 -2270
rect 2710 -2340 2725 -2310
rect 2755 -2340 2770 -2310
rect 2710 -2380 2770 -2340
rect 2710 -2410 2725 -2380
rect 2755 -2410 2770 -2380
rect 2710 -2445 2770 -2410
rect 2710 -2475 2725 -2445
rect 2755 -2475 2770 -2445
rect 2710 -2505 2770 -2475
rect 2710 -2535 2725 -2505
rect 2755 -2535 2770 -2505
rect 2710 -2570 2770 -2535
rect 2710 -2600 2725 -2570
rect 2755 -2600 2770 -2570
rect 2710 -2640 2770 -2600
rect 2710 -2670 2725 -2640
rect 2755 -2670 2770 -2640
rect 2710 -2710 2770 -2670
rect 2710 -2740 2725 -2710
rect 2755 -2740 2770 -2710
rect 2710 -2780 2770 -2740
rect 2710 -2810 2725 -2780
rect 2755 -2810 2770 -2780
rect 2710 -2845 2770 -2810
rect 2710 -2875 2725 -2845
rect 2755 -2875 2770 -2845
rect 2710 -2890 2770 -2875
rect 3060 -1305 3120 -1290
rect 3060 -1335 3075 -1305
rect 3105 -1335 3120 -1305
rect 3060 -1370 3120 -1335
rect 3060 -1400 3075 -1370
rect 3105 -1400 3120 -1370
rect 3060 -1440 3120 -1400
rect 3060 -1470 3075 -1440
rect 3105 -1470 3120 -1440
rect 3060 -1510 3120 -1470
rect 3060 -1540 3075 -1510
rect 3105 -1540 3120 -1510
rect 3060 -1580 3120 -1540
rect 3060 -1610 3075 -1580
rect 3105 -1610 3120 -1580
rect 3060 -1645 3120 -1610
rect 3060 -1675 3075 -1645
rect 3105 -1675 3120 -1645
rect 3060 -1705 3120 -1675
rect 3060 -1735 3075 -1705
rect 3105 -1735 3120 -1705
rect 3060 -1770 3120 -1735
rect 3060 -1800 3075 -1770
rect 3105 -1800 3120 -1770
rect 3060 -1840 3120 -1800
rect 3060 -1870 3075 -1840
rect 3105 -1870 3120 -1840
rect 3060 -1910 3120 -1870
rect 3060 -1940 3075 -1910
rect 3105 -1940 3120 -1910
rect 3060 -1980 3120 -1940
rect 3060 -2010 3075 -1980
rect 3105 -2010 3120 -1980
rect 3060 -2045 3120 -2010
rect 3060 -2075 3075 -2045
rect 3105 -2075 3120 -2045
rect 3060 -2105 3120 -2075
rect 3060 -2135 3075 -2105
rect 3105 -2135 3120 -2105
rect 3060 -2170 3120 -2135
rect 3060 -2200 3075 -2170
rect 3105 -2200 3120 -2170
rect 3060 -2240 3120 -2200
rect 3060 -2270 3075 -2240
rect 3105 -2270 3120 -2240
rect 3060 -2310 3120 -2270
rect 3060 -2340 3075 -2310
rect 3105 -2340 3120 -2310
rect 3060 -2380 3120 -2340
rect 3060 -2410 3075 -2380
rect 3105 -2410 3120 -2380
rect 3060 -2445 3120 -2410
rect 3060 -2475 3075 -2445
rect 3105 -2475 3120 -2445
rect 3060 -2505 3120 -2475
rect 3060 -2535 3075 -2505
rect 3105 -2535 3120 -2505
rect 3060 -2570 3120 -2535
rect 3060 -2600 3075 -2570
rect 3105 -2600 3120 -2570
rect 3060 -2640 3120 -2600
rect 3060 -2670 3075 -2640
rect 3105 -2670 3120 -2640
rect 3060 -2710 3120 -2670
rect 3060 -2740 3075 -2710
rect 3105 -2740 3120 -2710
rect 3060 -2780 3120 -2740
rect 3060 -2810 3075 -2780
rect 3105 -2810 3120 -2780
rect 3060 -2845 3120 -2810
rect 3060 -2875 3075 -2845
rect 3105 -2875 3120 -2845
rect 3060 -2890 3120 -2875
rect 3410 -1305 3470 -1290
rect 3410 -1335 3425 -1305
rect 3455 -1335 3470 -1305
rect 3410 -1370 3470 -1335
rect 3410 -1400 3425 -1370
rect 3455 -1400 3470 -1370
rect 3410 -1440 3470 -1400
rect 3410 -1470 3425 -1440
rect 3455 -1470 3470 -1440
rect 3410 -1510 3470 -1470
rect 3410 -1540 3425 -1510
rect 3455 -1540 3470 -1510
rect 3410 -1580 3470 -1540
rect 3410 -1610 3425 -1580
rect 3455 -1610 3470 -1580
rect 3410 -1645 3470 -1610
rect 3410 -1675 3425 -1645
rect 3455 -1675 3470 -1645
rect 3410 -1705 3470 -1675
rect 3410 -1735 3425 -1705
rect 3455 -1735 3470 -1705
rect 3410 -1770 3470 -1735
rect 3410 -1800 3425 -1770
rect 3455 -1800 3470 -1770
rect 3410 -1840 3470 -1800
rect 3410 -1870 3425 -1840
rect 3455 -1870 3470 -1840
rect 3410 -1910 3470 -1870
rect 3410 -1940 3425 -1910
rect 3455 -1940 3470 -1910
rect 3410 -1980 3470 -1940
rect 3410 -2010 3425 -1980
rect 3455 -2010 3470 -1980
rect 3410 -2045 3470 -2010
rect 3410 -2075 3425 -2045
rect 3455 -2075 3470 -2045
rect 3410 -2105 3470 -2075
rect 3410 -2135 3425 -2105
rect 3455 -2135 3470 -2105
rect 3410 -2170 3470 -2135
rect 3410 -2200 3425 -2170
rect 3455 -2200 3470 -2170
rect 3410 -2240 3470 -2200
rect 3410 -2270 3425 -2240
rect 3455 -2270 3470 -2240
rect 3410 -2310 3470 -2270
rect 3410 -2340 3425 -2310
rect 3455 -2340 3470 -2310
rect 3410 -2380 3470 -2340
rect 3410 -2410 3425 -2380
rect 3455 -2410 3470 -2380
rect 3410 -2445 3470 -2410
rect 3410 -2475 3425 -2445
rect 3455 -2475 3470 -2445
rect 3410 -2505 3470 -2475
rect 3410 -2535 3425 -2505
rect 3455 -2535 3470 -2505
rect 3410 -2570 3470 -2535
rect 3410 -2600 3425 -2570
rect 3455 -2600 3470 -2570
rect 3410 -2640 3470 -2600
rect 3410 -2670 3425 -2640
rect 3455 -2670 3470 -2640
rect 3410 -2710 3470 -2670
rect 3410 -2740 3425 -2710
rect 3455 -2740 3470 -2710
rect 3410 -2780 3470 -2740
rect 3410 -2810 3425 -2780
rect 3455 -2810 3470 -2780
rect 3410 -2845 3470 -2810
rect 3410 -2875 3425 -2845
rect 3455 -2875 3470 -2845
rect 3410 -2890 3470 -2875
rect 3760 -1305 3820 -1290
rect 3760 -1335 3775 -1305
rect 3805 -1335 3820 -1305
rect 3760 -1370 3820 -1335
rect 3760 -1400 3775 -1370
rect 3805 -1400 3820 -1370
rect 3760 -1440 3820 -1400
rect 3760 -1470 3775 -1440
rect 3805 -1470 3820 -1440
rect 3760 -1510 3820 -1470
rect 3760 -1540 3775 -1510
rect 3805 -1540 3820 -1510
rect 3760 -1580 3820 -1540
rect 3760 -1610 3775 -1580
rect 3805 -1610 3820 -1580
rect 3760 -1645 3820 -1610
rect 3760 -1675 3775 -1645
rect 3805 -1675 3820 -1645
rect 3760 -1705 3820 -1675
rect 3760 -1735 3775 -1705
rect 3805 -1735 3820 -1705
rect 3760 -1770 3820 -1735
rect 3760 -1800 3775 -1770
rect 3805 -1800 3820 -1770
rect 3760 -1840 3820 -1800
rect 3760 -1870 3775 -1840
rect 3805 -1870 3820 -1840
rect 3760 -1910 3820 -1870
rect 3760 -1940 3775 -1910
rect 3805 -1940 3820 -1910
rect 3760 -1980 3820 -1940
rect 3760 -2010 3775 -1980
rect 3805 -2010 3820 -1980
rect 3760 -2045 3820 -2010
rect 3760 -2075 3775 -2045
rect 3805 -2075 3820 -2045
rect 3760 -2105 3820 -2075
rect 3760 -2135 3775 -2105
rect 3805 -2135 3820 -2105
rect 3760 -2170 3820 -2135
rect 3760 -2200 3775 -2170
rect 3805 -2200 3820 -2170
rect 3760 -2240 3820 -2200
rect 3760 -2270 3775 -2240
rect 3805 -2270 3820 -2240
rect 3760 -2310 3820 -2270
rect 3760 -2340 3775 -2310
rect 3805 -2340 3820 -2310
rect 3760 -2380 3820 -2340
rect 3760 -2410 3775 -2380
rect 3805 -2410 3820 -2380
rect 3760 -2445 3820 -2410
rect 3760 -2475 3775 -2445
rect 3805 -2475 3820 -2445
rect 3760 -2505 3820 -2475
rect 3760 -2535 3775 -2505
rect 3805 -2535 3820 -2505
rect 3760 -2570 3820 -2535
rect 3760 -2600 3775 -2570
rect 3805 -2600 3820 -2570
rect 3760 -2640 3820 -2600
rect 3760 -2670 3775 -2640
rect 3805 -2670 3820 -2640
rect 3760 -2710 3820 -2670
rect 3760 -2740 3775 -2710
rect 3805 -2740 3820 -2710
rect 3760 -2780 3820 -2740
rect 3760 -2810 3775 -2780
rect 3805 -2810 3820 -2780
rect 3760 -2845 3820 -2810
rect 3760 -2875 3775 -2845
rect 3805 -2875 3820 -2845
rect 3760 -2890 3820 -2875
rect 4110 -1305 4170 -1290
rect 4110 -1335 4125 -1305
rect 4155 -1335 4170 -1305
rect 4110 -1370 4170 -1335
rect 4110 -1400 4125 -1370
rect 4155 -1400 4170 -1370
rect 4110 -1440 4170 -1400
rect 4110 -1470 4125 -1440
rect 4155 -1470 4170 -1440
rect 4110 -1510 4170 -1470
rect 4110 -1540 4125 -1510
rect 4155 -1540 4170 -1510
rect 4110 -1580 4170 -1540
rect 4110 -1610 4125 -1580
rect 4155 -1610 4170 -1580
rect 4110 -1645 4170 -1610
rect 4110 -1675 4125 -1645
rect 4155 -1675 4170 -1645
rect 4110 -1705 4170 -1675
rect 4110 -1735 4125 -1705
rect 4155 -1735 4170 -1705
rect 4110 -1770 4170 -1735
rect 4110 -1800 4125 -1770
rect 4155 -1800 4170 -1770
rect 4110 -1840 4170 -1800
rect 4110 -1870 4125 -1840
rect 4155 -1870 4170 -1840
rect 4110 -1910 4170 -1870
rect 4110 -1940 4125 -1910
rect 4155 -1940 4170 -1910
rect 4110 -1980 4170 -1940
rect 4110 -2010 4125 -1980
rect 4155 -2010 4170 -1980
rect 4110 -2045 4170 -2010
rect 4110 -2075 4125 -2045
rect 4155 -2075 4170 -2045
rect 4110 -2105 4170 -2075
rect 4110 -2135 4125 -2105
rect 4155 -2135 4170 -2105
rect 4110 -2170 4170 -2135
rect 4110 -2200 4125 -2170
rect 4155 -2200 4170 -2170
rect 4110 -2240 4170 -2200
rect 4110 -2270 4125 -2240
rect 4155 -2270 4170 -2240
rect 4110 -2310 4170 -2270
rect 4110 -2340 4125 -2310
rect 4155 -2340 4170 -2310
rect 4110 -2380 4170 -2340
rect 4110 -2410 4125 -2380
rect 4155 -2410 4170 -2380
rect 4110 -2445 4170 -2410
rect 4110 -2475 4125 -2445
rect 4155 -2475 4170 -2445
rect 4110 -2505 4170 -2475
rect 4110 -2535 4125 -2505
rect 4155 -2535 4170 -2505
rect 4110 -2570 4170 -2535
rect 4110 -2600 4125 -2570
rect 4155 -2600 4170 -2570
rect 4110 -2640 4170 -2600
rect 4110 -2670 4125 -2640
rect 4155 -2670 4170 -2640
rect 4110 -2710 4170 -2670
rect 4110 -2740 4125 -2710
rect 4155 -2740 4170 -2710
rect 4110 -2780 4170 -2740
rect 4110 -2810 4125 -2780
rect 4155 -2810 4170 -2780
rect 4110 -2845 4170 -2810
rect 4110 -2875 4125 -2845
rect 4155 -2875 4170 -2845
rect 4110 -2890 4170 -2875
rect 4460 -1305 4520 -1290
rect 4460 -1335 4475 -1305
rect 4505 -1335 4520 -1305
rect 4460 -1370 4520 -1335
rect 4460 -1400 4475 -1370
rect 4505 -1400 4520 -1370
rect 4460 -1440 4520 -1400
rect 4460 -1470 4475 -1440
rect 4505 -1470 4520 -1440
rect 4460 -1510 4520 -1470
rect 4460 -1540 4475 -1510
rect 4505 -1540 4520 -1510
rect 4460 -1580 4520 -1540
rect 4460 -1610 4475 -1580
rect 4505 -1610 4520 -1580
rect 4460 -1645 4520 -1610
rect 4460 -1675 4475 -1645
rect 4505 -1675 4520 -1645
rect 4460 -1705 4520 -1675
rect 4460 -1735 4475 -1705
rect 4505 -1735 4520 -1705
rect 4460 -1770 4520 -1735
rect 4460 -1800 4475 -1770
rect 4505 -1800 4520 -1770
rect 4460 -1840 4520 -1800
rect 4460 -1870 4475 -1840
rect 4505 -1870 4520 -1840
rect 4460 -1910 4520 -1870
rect 4460 -1940 4475 -1910
rect 4505 -1940 4520 -1910
rect 4460 -1980 4520 -1940
rect 4460 -2010 4475 -1980
rect 4505 -2010 4520 -1980
rect 4460 -2045 4520 -2010
rect 4460 -2075 4475 -2045
rect 4505 -2075 4520 -2045
rect 4460 -2105 4520 -2075
rect 4460 -2135 4475 -2105
rect 4505 -2135 4520 -2105
rect 4460 -2170 4520 -2135
rect 4460 -2200 4475 -2170
rect 4505 -2200 4520 -2170
rect 4460 -2240 4520 -2200
rect 4460 -2270 4475 -2240
rect 4505 -2270 4520 -2240
rect 4460 -2310 4520 -2270
rect 4460 -2340 4475 -2310
rect 4505 -2340 4520 -2310
rect 4460 -2380 4520 -2340
rect 4460 -2410 4475 -2380
rect 4505 -2410 4520 -2380
rect 4460 -2445 4520 -2410
rect 4460 -2475 4475 -2445
rect 4505 -2475 4520 -2445
rect 4460 -2505 4520 -2475
rect 4460 -2535 4475 -2505
rect 4505 -2535 4520 -2505
rect 4460 -2570 4520 -2535
rect 4460 -2600 4475 -2570
rect 4505 -2600 4520 -2570
rect 4460 -2640 4520 -2600
rect 4460 -2670 4475 -2640
rect 4505 -2670 4520 -2640
rect 4460 -2710 4520 -2670
rect 4460 -2740 4475 -2710
rect 4505 -2740 4520 -2710
rect 4460 -2780 4520 -2740
rect 4460 -2810 4475 -2780
rect 4505 -2810 4520 -2780
rect 4460 -2845 4520 -2810
rect 4460 -2875 4475 -2845
rect 4505 -2875 4520 -2845
rect 4460 -2890 4520 -2875
rect 4810 -1305 4870 -1290
rect 4810 -1335 4825 -1305
rect 4855 -1335 4870 -1305
rect 4810 -1370 4870 -1335
rect 4810 -1400 4825 -1370
rect 4855 -1400 4870 -1370
rect 4810 -1440 4870 -1400
rect 4810 -1470 4825 -1440
rect 4855 -1470 4870 -1440
rect 4810 -1510 4870 -1470
rect 4810 -1540 4825 -1510
rect 4855 -1540 4870 -1510
rect 4810 -1580 4870 -1540
rect 4810 -1610 4825 -1580
rect 4855 -1610 4870 -1580
rect 4810 -1645 4870 -1610
rect 4810 -1675 4825 -1645
rect 4855 -1675 4870 -1645
rect 4810 -1705 4870 -1675
rect 4810 -1735 4825 -1705
rect 4855 -1735 4870 -1705
rect 4810 -1770 4870 -1735
rect 4810 -1800 4825 -1770
rect 4855 -1800 4870 -1770
rect 4810 -1840 4870 -1800
rect 4810 -1870 4825 -1840
rect 4855 -1870 4870 -1840
rect 4810 -1910 4870 -1870
rect 4810 -1940 4825 -1910
rect 4855 -1940 4870 -1910
rect 4810 -1980 4870 -1940
rect 4810 -2010 4825 -1980
rect 4855 -2010 4870 -1980
rect 4810 -2045 4870 -2010
rect 4810 -2075 4825 -2045
rect 4855 -2075 4870 -2045
rect 4810 -2105 4870 -2075
rect 4810 -2135 4825 -2105
rect 4855 -2135 4870 -2105
rect 4810 -2170 4870 -2135
rect 4810 -2200 4825 -2170
rect 4855 -2200 4870 -2170
rect 4810 -2240 4870 -2200
rect 4810 -2270 4825 -2240
rect 4855 -2270 4870 -2240
rect 4810 -2310 4870 -2270
rect 4810 -2340 4825 -2310
rect 4855 -2340 4870 -2310
rect 4810 -2380 4870 -2340
rect 4810 -2410 4825 -2380
rect 4855 -2410 4870 -2380
rect 4810 -2445 4870 -2410
rect 4810 -2475 4825 -2445
rect 4855 -2475 4870 -2445
rect 4810 -2505 4870 -2475
rect 4810 -2535 4825 -2505
rect 4855 -2535 4870 -2505
rect 4810 -2570 4870 -2535
rect 4810 -2600 4825 -2570
rect 4855 -2600 4870 -2570
rect 4810 -2640 4870 -2600
rect 4810 -2670 4825 -2640
rect 4855 -2670 4870 -2640
rect 4810 -2710 4870 -2670
rect 4810 -2740 4825 -2710
rect 4855 -2740 4870 -2710
rect 4810 -2780 4870 -2740
rect 4810 -2810 4825 -2780
rect 4855 -2810 4870 -2780
rect 4810 -2845 4870 -2810
rect 4810 -2875 4825 -2845
rect 4855 -2875 4870 -2845
rect 4810 -2890 4870 -2875
rect 5160 -1305 5220 -1290
rect 5160 -1335 5175 -1305
rect 5205 -1335 5220 -1305
rect 5160 -1370 5220 -1335
rect 5160 -1400 5175 -1370
rect 5205 -1400 5220 -1370
rect 5160 -1440 5220 -1400
rect 5160 -1470 5175 -1440
rect 5205 -1470 5220 -1440
rect 5160 -1510 5220 -1470
rect 5160 -1540 5175 -1510
rect 5205 -1540 5220 -1510
rect 5160 -1580 5220 -1540
rect 5160 -1610 5175 -1580
rect 5205 -1610 5220 -1580
rect 5160 -1645 5220 -1610
rect 5160 -1675 5175 -1645
rect 5205 -1675 5220 -1645
rect 5160 -1705 5220 -1675
rect 5160 -1735 5175 -1705
rect 5205 -1735 5220 -1705
rect 5160 -1770 5220 -1735
rect 5160 -1800 5175 -1770
rect 5205 -1800 5220 -1770
rect 5160 -1840 5220 -1800
rect 5160 -1870 5175 -1840
rect 5205 -1870 5220 -1840
rect 5160 -1910 5220 -1870
rect 5160 -1940 5175 -1910
rect 5205 -1940 5220 -1910
rect 5160 -1980 5220 -1940
rect 5160 -2010 5175 -1980
rect 5205 -2010 5220 -1980
rect 5160 -2045 5220 -2010
rect 5160 -2075 5175 -2045
rect 5205 -2075 5220 -2045
rect 5160 -2105 5220 -2075
rect 5160 -2135 5175 -2105
rect 5205 -2135 5220 -2105
rect 5160 -2170 5220 -2135
rect 5160 -2200 5175 -2170
rect 5205 -2200 5220 -2170
rect 5160 -2240 5220 -2200
rect 5160 -2270 5175 -2240
rect 5205 -2270 5220 -2240
rect 5160 -2310 5220 -2270
rect 5160 -2340 5175 -2310
rect 5205 -2340 5220 -2310
rect 5160 -2380 5220 -2340
rect 5160 -2410 5175 -2380
rect 5205 -2410 5220 -2380
rect 5160 -2445 5220 -2410
rect 5160 -2475 5175 -2445
rect 5205 -2475 5220 -2445
rect 5160 -2505 5220 -2475
rect 5160 -2535 5175 -2505
rect 5205 -2535 5220 -2505
rect 5160 -2570 5220 -2535
rect 5160 -2600 5175 -2570
rect 5205 -2600 5220 -2570
rect 5160 -2640 5220 -2600
rect 5160 -2670 5175 -2640
rect 5205 -2670 5220 -2640
rect 5160 -2710 5220 -2670
rect 5160 -2740 5175 -2710
rect 5205 -2740 5220 -2710
rect 5160 -2780 5220 -2740
rect 5160 -2810 5175 -2780
rect 5205 -2810 5220 -2780
rect 5160 -2845 5220 -2810
rect 5160 -2875 5175 -2845
rect 5205 -2875 5220 -2845
rect 5160 -2890 5220 -2875
rect 5510 -1305 5570 -1290
rect 5510 -1335 5525 -1305
rect 5555 -1335 5570 -1305
rect 5510 -1370 5570 -1335
rect 5510 -1400 5525 -1370
rect 5555 -1400 5570 -1370
rect 5510 -1440 5570 -1400
rect 5510 -1470 5525 -1440
rect 5555 -1470 5570 -1440
rect 5510 -1510 5570 -1470
rect 5510 -1540 5525 -1510
rect 5555 -1540 5570 -1510
rect 5510 -1580 5570 -1540
rect 5510 -1610 5525 -1580
rect 5555 -1610 5570 -1580
rect 5510 -1645 5570 -1610
rect 5510 -1675 5525 -1645
rect 5555 -1675 5570 -1645
rect 5510 -1705 5570 -1675
rect 5510 -1735 5525 -1705
rect 5555 -1735 5570 -1705
rect 5510 -1770 5570 -1735
rect 5510 -1800 5525 -1770
rect 5555 -1800 5570 -1770
rect 5510 -1840 5570 -1800
rect 5510 -1870 5525 -1840
rect 5555 -1870 5570 -1840
rect 5510 -1910 5570 -1870
rect 5510 -1940 5525 -1910
rect 5555 -1940 5570 -1910
rect 5510 -1980 5570 -1940
rect 5510 -2010 5525 -1980
rect 5555 -2010 5570 -1980
rect 5510 -2045 5570 -2010
rect 5510 -2075 5525 -2045
rect 5555 -2075 5570 -2045
rect 5510 -2105 5570 -2075
rect 5510 -2135 5525 -2105
rect 5555 -2135 5570 -2105
rect 5510 -2170 5570 -2135
rect 5510 -2200 5525 -2170
rect 5555 -2200 5570 -2170
rect 5510 -2240 5570 -2200
rect 5510 -2270 5525 -2240
rect 5555 -2270 5570 -2240
rect 5510 -2310 5570 -2270
rect 5510 -2340 5525 -2310
rect 5555 -2340 5570 -2310
rect 5510 -2380 5570 -2340
rect 5510 -2410 5525 -2380
rect 5555 -2410 5570 -2380
rect 5510 -2445 5570 -2410
rect 5510 -2475 5525 -2445
rect 5555 -2475 5570 -2445
rect 5510 -2505 5570 -2475
rect 5510 -2535 5525 -2505
rect 5555 -2535 5570 -2505
rect 5510 -2570 5570 -2535
rect 5510 -2600 5525 -2570
rect 5555 -2600 5570 -2570
rect 5510 -2640 5570 -2600
rect 5510 -2670 5525 -2640
rect 5555 -2670 5570 -2640
rect 5510 -2710 5570 -2670
rect 5510 -2740 5525 -2710
rect 5555 -2740 5570 -2710
rect 5510 -2780 5570 -2740
rect 5510 -2810 5525 -2780
rect 5555 -2810 5570 -2780
rect 5510 -2845 5570 -2810
rect 5510 -2875 5525 -2845
rect 5555 -2875 5570 -2845
rect 5510 -2890 5570 -2875
rect 5860 -1305 5920 -1290
rect 5860 -1335 5875 -1305
rect 5905 -1335 5920 -1305
rect 5860 -1370 5920 -1335
rect 5860 -1400 5875 -1370
rect 5905 -1400 5920 -1370
rect 5860 -1440 5920 -1400
rect 5860 -1470 5875 -1440
rect 5905 -1470 5920 -1440
rect 5860 -1510 5920 -1470
rect 5860 -1540 5875 -1510
rect 5905 -1540 5920 -1510
rect 5860 -1580 5920 -1540
rect 5860 -1610 5875 -1580
rect 5905 -1610 5920 -1580
rect 5860 -1645 5920 -1610
rect 5860 -1675 5875 -1645
rect 5905 -1675 5920 -1645
rect 5860 -1705 5920 -1675
rect 5860 -1735 5875 -1705
rect 5905 -1735 5920 -1705
rect 5860 -1770 5920 -1735
rect 5860 -1800 5875 -1770
rect 5905 -1800 5920 -1770
rect 5860 -1840 5920 -1800
rect 5860 -1870 5875 -1840
rect 5905 -1870 5920 -1840
rect 5860 -1910 5920 -1870
rect 5860 -1940 5875 -1910
rect 5905 -1940 5920 -1910
rect 5860 -1980 5920 -1940
rect 5860 -2010 5875 -1980
rect 5905 -2010 5920 -1980
rect 5860 -2045 5920 -2010
rect 5860 -2075 5875 -2045
rect 5905 -2075 5920 -2045
rect 5860 -2105 5920 -2075
rect 5860 -2135 5875 -2105
rect 5905 -2135 5920 -2105
rect 5860 -2170 5920 -2135
rect 5860 -2200 5875 -2170
rect 5905 -2200 5920 -2170
rect 5860 -2240 5920 -2200
rect 5860 -2270 5875 -2240
rect 5905 -2270 5920 -2240
rect 5860 -2310 5920 -2270
rect 5860 -2340 5875 -2310
rect 5905 -2340 5920 -2310
rect 5860 -2380 5920 -2340
rect 5860 -2410 5875 -2380
rect 5905 -2410 5920 -2380
rect 5860 -2445 5920 -2410
rect 5860 -2475 5875 -2445
rect 5905 -2475 5920 -2445
rect 5860 -2505 5920 -2475
rect 5860 -2535 5875 -2505
rect 5905 -2535 5920 -2505
rect 5860 -2570 5920 -2535
rect 5860 -2600 5875 -2570
rect 5905 -2600 5920 -2570
rect 5860 -2640 5920 -2600
rect 5860 -2670 5875 -2640
rect 5905 -2670 5920 -2640
rect 5860 -2710 5920 -2670
rect 5860 -2740 5875 -2710
rect 5905 -2740 5920 -2710
rect 5860 -2780 5920 -2740
rect 5860 -2810 5875 -2780
rect 5905 -2810 5920 -2780
rect 5860 -2845 5920 -2810
rect 5860 -2875 5875 -2845
rect 5905 -2875 5920 -2845
rect 5860 -2890 5920 -2875
rect 6210 -1305 6270 -1290
rect 6210 -1335 6225 -1305
rect 6255 -1335 6270 -1305
rect 6210 -1370 6270 -1335
rect 6210 -1400 6225 -1370
rect 6255 -1400 6270 -1370
rect 6210 -1440 6270 -1400
rect 6210 -1470 6225 -1440
rect 6255 -1470 6270 -1440
rect 6210 -1510 6270 -1470
rect 6210 -1540 6225 -1510
rect 6255 -1540 6270 -1510
rect 6210 -1580 6270 -1540
rect 6210 -1610 6225 -1580
rect 6255 -1610 6270 -1580
rect 6210 -1645 6270 -1610
rect 6210 -1675 6225 -1645
rect 6255 -1675 6270 -1645
rect 6210 -1705 6270 -1675
rect 6210 -1735 6225 -1705
rect 6255 -1735 6270 -1705
rect 6210 -1770 6270 -1735
rect 6210 -1800 6225 -1770
rect 6255 -1800 6270 -1770
rect 6210 -1840 6270 -1800
rect 6210 -1870 6225 -1840
rect 6255 -1870 6270 -1840
rect 6210 -1910 6270 -1870
rect 6210 -1940 6225 -1910
rect 6255 -1940 6270 -1910
rect 6210 -1980 6270 -1940
rect 6210 -2010 6225 -1980
rect 6255 -2010 6270 -1980
rect 6210 -2045 6270 -2010
rect 6210 -2075 6225 -2045
rect 6255 -2075 6270 -2045
rect 6210 -2105 6270 -2075
rect 6210 -2135 6225 -2105
rect 6255 -2135 6270 -2105
rect 6210 -2170 6270 -2135
rect 6210 -2200 6225 -2170
rect 6255 -2200 6270 -2170
rect 6210 -2240 6270 -2200
rect 6210 -2270 6225 -2240
rect 6255 -2270 6270 -2240
rect 6210 -2310 6270 -2270
rect 6210 -2340 6225 -2310
rect 6255 -2340 6270 -2310
rect 6210 -2380 6270 -2340
rect 6210 -2410 6225 -2380
rect 6255 -2410 6270 -2380
rect 6210 -2445 6270 -2410
rect 6210 -2475 6225 -2445
rect 6255 -2475 6270 -2445
rect 6210 -2505 6270 -2475
rect 6210 -2535 6225 -2505
rect 6255 -2535 6270 -2505
rect 6210 -2570 6270 -2535
rect 6210 -2600 6225 -2570
rect 6255 -2600 6270 -2570
rect 6210 -2640 6270 -2600
rect 6210 -2670 6225 -2640
rect 6255 -2670 6270 -2640
rect 6210 -2710 6270 -2670
rect 6210 -2740 6225 -2710
rect 6255 -2740 6270 -2710
rect 6210 -2780 6270 -2740
rect 6210 -2810 6225 -2780
rect 6255 -2810 6270 -2780
rect 6210 -2845 6270 -2810
rect 6210 -2875 6225 -2845
rect 6255 -2875 6270 -2845
rect 6210 -2890 6270 -2875
rect 6560 -1305 6620 -1290
rect 6560 -1335 6575 -1305
rect 6605 -1335 6620 -1305
rect 6560 -1370 6620 -1335
rect 6560 -1400 6575 -1370
rect 6605 -1400 6620 -1370
rect 6560 -1440 6620 -1400
rect 6560 -1470 6575 -1440
rect 6605 -1470 6620 -1440
rect 6560 -1510 6620 -1470
rect 6560 -1540 6575 -1510
rect 6605 -1540 6620 -1510
rect 6560 -1580 6620 -1540
rect 6560 -1610 6575 -1580
rect 6605 -1610 6620 -1580
rect 6560 -1645 6620 -1610
rect 6560 -1675 6575 -1645
rect 6605 -1675 6620 -1645
rect 6560 -1705 6620 -1675
rect 6560 -1735 6575 -1705
rect 6605 -1735 6620 -1705
rect 6560 -1770 6620 -1735
rect 6560 -1800 6575 -1770
rect 6605 -1800 6620 -1770
rect 6560 -1840 6620 -1800
rect 6560 -1870 6575 -1840
rect 6605 -1870 6620 -1840
rect 6560 -1910 6620 -1870
rect 6560 -1940 6575 -1910
rect 6605 -1940 6620 -1910
rect 6560 -1980 6620 -1940
rect 6560 -2010 6575 -1980
rect 6605 -2010 6620 -1980
rect 6560 -2045 6620 -2010
rect 6560 -2075 6575 -2045
rect 6605 -2075 6620 -2045
rect 6560 -2105 6620 -2075
rect 6560 -2135 6575 -2105
rect 6605 -2135 6620 -2105
rect 6560 -2170 6620 -2135
rect 6560 -2200 6575 -2170
rect 6605 -2200 6620 -2170
rect 6560 -2240 6620 -2200
rect 6560 -2270 6575 -2240
rect 6605 -2270 6620 -2240
rect 6560 -2310 6620 -2270
rect 6560 -2340 6575 -2310
rect 6605 -2340 6620 -2310
rect 6560 -2380 6620 -2340
rect 6560 -2410 6575 -2380
rect 6605 -2410 6620 -2380
rect 6560 -2445 6620 -2410
rect 6560 -2475 6575 -2445
rect 6605 -2475 6620 -2445
rect 6560 -2505 6620 -2475
rect 6560 -2535 6575 -2505
rect 6605 -2535 6620 -2505
rect 6560 -2570 6620 -2535
rect 6560 -2600 6575 -2570
rect 6605 -2600 6620 -2570
rect 6560 -2640 6620 -2600
rect 6560 -2670 6575 -2640
rect 6605 -2670 6620 -2640
rect 6560 -2710 6620 -2670
rect 6560 -2740 6575 -2710
rect 6605 -2740 6620 -2710
rect 6560 -2780 6620 -2740
rect 6560 -2810 6575 -2780
rect 6605 -2810 6620 -2780
rect 6560 -2845 6620 -2810
rect 6560 -2875 6575 -2845
rect 6605 -2875 6620 -2845
rect 6560 -2890 6620 -2875
rect 6910 -1305 6970 -1290
rect 6910 -1335 6925 -1305
rect 6955 -1335 6970 -1305
rect 6910 -1370 6970 -1335
rect 6910 -1400 6925 -1370
rect 6955 -1400 6970 -1370
rect 6910 -1440 6970 -1400
rect 6910 -1470 6925 -1440
rect 6955 -1470 6970 -1440
rect 6910 -1510 6970 -1470
rect 6910 -1540 6925 -1510
rect 6955 -1540 6970 -1510
rect 6910 -1580 6970 -1540
rect 6910 -1610 6925 -1580
rect 6955 -1610 6970 -1580
rect 6910 -1645 6970 -1610
rect 6910 -1675 6925 -1645
rect 6955 -1675 6970 -1645
rect 6910 -1705 6970 -1675
rect 6910 -1735 6925 -1705
rect 6955 -1735 6970 -1705
rect 6910 -1770 6970 -1735
rect 6910 -1800 6925 -1770
rect 6955 -1800 6970 -1770
rect 6910 -1840 6970 -1800
rect 6910 -1870 6925 -1840
rect 6955 -1870 6970 -1840
rect 6910 -1910 6970 -1870
rect 6910 -1940 6925 -1910
rect 6955 -1940 6970 -1910
rect 6910 -1980 6970 -1940
rect 6910 -2010 6925 -1980
rect 6955 -2010 6970 -1980
rect 6910 -2045 6970 -2010
rect 6910 -2075 6925 -2045
rect 6955 -2075 6970 -2045
rect 6910 -2105 6970 -2075
rect 6910 -2135 6925 -2105
rect 6955 -2135 6970 -2105
rect 6910 -2170 6970 -2135
rect 6910 -2200 6925 -2170
rect 6955 -2200 6970 -2170
rect 6910 -2240 6970 -2200
rect 6910 -2270 6925 -2240
rect 6955 -2270 6970 -2240
rect 6910 -2310 6970 -2270
rect 6910 -2340 6925 -2310
rect 6955 -2340 6970 -2310
rect 6910 -2380 6970 -2340
rect 6910 -2410 6925 -2380
rect 6955 -2410 6970 -2380
rect 6910 -2445 6970 -2410
rect 6910 -2475 6925 -2445
rect 6955 -2475 6970 -2445
rect 6910 -2505 6970 -2475
rect 6910 -2535 6925 -2505
rect 6955 -2535 6970 -2505
rect 6910 -2570 6970 -2535
rect 6910 -2600 6925 -2570
rect 6955 -2600 6970 -2570
rect 6910 -2640 6970 -2600
rect 6910 -2670 6925 -2640
rect 6955 -2670 6970 -2640
rect 6910 -2710 6970 -2670
rect 6910 -2740 6925 -2710
rect 6955 -2740 6970 -2710
rect 6910 -2780 6970 -2740
rect 6910 -2810 6925 -2780
rect 6955 -2810 6970 -2780
rect 6910 -2845 6970 -2810
rect 6910 -2875 6925 -2845
rect 6955 -2875 6970 -2845
rect 6910 -2890 6970 -2875
rect 7260 -1305 7320 -1290
rect 7260 -1335 7275 -1305
rect 7305 -1335 7320 -1305
rect 7260 -1370 7320 -1335
rect 7260 -1400 7275 -1370
rect 7305 -1400 7320 -1370
rect 7260 -1440 7320 -1400
rect 7260 -1470 7275 -1440
rect 7305 -1470 7320 -1440
rect 7260 -1510 7320 -1470
rect 7260 -1540 7275 -1510
rect 7305 -1540 7320 -1510
rect 7260 -1580 7320 -1540
rect 7260 -1610 7275 -1580
rect 7305 -1610 7320 -1580
rect 7260 -1645 7320 -1610
rect 7260 -1675 7275 -1645
rect 7305 -1675 7320 -1645
rect 7260 -1705 7320 -1675
rect 7260 -1735 7275 -1705
rect 7305 -1735 7320 -1705
rect 7260 -1770 7320 -1735
rect 7260 -1800 7275 -1770
rect 7305 -1800 7320 -1770
rect 7260 -1840 7320 -1800
rect 7260 -1870 7275 -1840
rect 7305 -1870 7320 -1840
rect 7260 -1910 7320 -1870
rect 7260 -1940 7275 -1910
rect 7305 -1940 7320 -1910
rect 7260 -1980 7320 -1940
rect 7260 -2010 7275 -1980
rect 7305 -2010 7320 -1980
rect 7260 -2045 7320 -2010
rect 7260 -2075 7275 -2045
rect 7305 -2075 7320 -2045
rect 7260 -2105 7320 -2075
rect 7260 -2135 7275 -2105
rect 7305 -2135 7320 -2105
rect 7260 -2170 7320 -2135
rect 7260 -2200 7275 -2170
rect 7305 -2200 7320 -2170
rect 7260 -2240 7320 -2200
rect 7260 -2270 7275 -2240
rect 7305 -2270 7320 -2240
rect 7260 -2310 7320 -2270
rect 7260 -2340 7275 -2310
rect 7305 -2340 7320 -2310
rect 7260 -2380 7320 -2340
rect 7260 -2410 7275 -2380
rect 7305 -2410 7320 -2380
rect 7260 -2445 7320 -2410
rect 7260 -2475 7275 -2445
rect 7305 -2475 7320 -2445
rect 7260 -2505 7320 -2475
rect 7260 -2535 7275 -2505
rect 7305 -2535 7320 -2505
rect 7260 -2570 7320 -2535
rect 7260 -2600 7275 -2570
rect 7305 -2600 7320 -2570
rect 7260 -2640 7320 -2600
rect 7260 -2670 7275 -2640
rect 7305 -2670 7320 -2640
rect 7260 -2710 7320 -2670
rect 7260 -2740 7275 -2710
rect 7305 -2740 7320 -2710
rect 7260 -2780 7320 -2740
rect 7260 -2810 7275 -2780
rect 7305 -2810 7320 -2780
rect 7260 -2845 7320 -2810
rect 7260 -2875 7275 -2845
rect 7305 -2875 7320 -2845
rect 7260 -2890 7320 -2875
rect 7610 -1305 7670 -1290
rect 7610 -1335 7625 -1305
rect 7655 -1335 7670 -1305
rect 7610 -1370 7670 -1335
rect 7610 -1400 7625 -1370
rect 7655 -1400 7670 -1370
rect 7610 -1440 7670 -1400
rect 7610 -1470 7625 -1440
rect 7655 -1470 7670 -1440
rect 7610 -1510 7670 -1470
rect 7610 -1540 7625 -1510
rect 7655 -1540 7670 -1510
rect 7610 -1580 7670 -1540
rect 7610 -1610 7625 -1580
rect 7655 -1610 7670 -1580
rect 7610 -1645 7670 -1610
rect 7610 -1675 7625 -1645
rect 7655 -1675 7670 -1645
rect 7610 -1705 7670 -1675
rect 7610 -1735 7625 -1705
rect 7655 -1735 7670 -1705
rect 7610 -1770 7670 -1735
rect 7610 -1800 7625 -1770
rect 7655 -1800 7670 -1770
rect 7610 -1840 7670 -1800
rect 7610 -1870 7625 -1840
rect 7655 -1870 7670 -1840
rect 7610 -1910 7670 -1870
rect 7610 -1940 7625 -1910
rect 7655 -1940 7670 -1910
rect 7610 -1980 7670 -1940
rect 7610 -2010 7625 -1980
rect 7655 -2010 7670 -1980
rect 7610 -2045 7670 -2010
rect 7610 -2075 7625 -2045
rect 7655 -2075 7670 -2045
rect 7610 -2105 7670 -2075
rect 7610 -2135 7625 -2105
rect 7655 -2135 7670 -2105
rect 7610 -2170 7670 -2135
rect 7610 -2200 7625 -2170
rect 7655 -2200 7670 -2170
rect 7610 -2240 7670 -2200
rect 7610 -2270 7625 -2240
rect 7655 -2270 7670 -2240
rect 7610 -2310 7670 -2270
rect 7610 -2340 7625 -2310
rect 7655 -2340 7670 -2310
rect 7610 -2380 7670 -2340
rect 7610 -2410 7625 -2380
rect 7655 -2410 7670 -2380
rect 7610 -2445 7670 -2410
rect 7610 -2475 7625 -2445
rect 7655 -2475 7670 -2445
rect 7610 -2505 7670 -2475
rect 7610 -2535 7625 -2505
rect 7655 -2535 7670 -2505
rect 7610 -2570 7670 -2535
rect 7610 -2600 7625 -2570
rect 7655 -2600 7670 -2570
rect 7610 -2640 7670 -2600
rect 7610 -2670 7625 -2640
rect 7655 -2670 7670 -2640
rect 7610 -2710 7670 -2670
rect 7610 -2740 7625 -2710
rect 7655 -2740 7670 -2710
rect 7610 -2780 7670 -2740
rect 7610 -2810 7625 -2780
rect 7655 -2810 7670 -2780
rect 7610 -2845 7670 -2810
rect 7610 -2875 7625 -2845
rect 7655 -2875 7670 -2845
rect 7610 -2890 7670 -2875
rect 7960 -1305 8020 -1290
rect 7960 -1335 7975 -1305
rect 8005 -1335 8020 -1305
rect 7960 -1370 8020 -1335
rect 7960 -1400 7975 -1370
rect 8005 -1400 8020 -1370
rect 7960 -1440 8020 -1400
rect 7960 -1470 7975 -1440
rect 8005 -1470 8020 -1440
rect 7960 -1510 8020 -1470
rect 7960 -1540 7975 -1510
rect 8005 -1540 8020 -1510
rect 7960 -1580 8020 -1540
rect 7960 -1610 7975 -1580
rect 8005 -1610 8020 -1580
rect 7960 -1645 8020 -1610
rect 7960 -1675 7975 -1645
rect 8005 -1675 8020 -1645
rect 7960 -1705 8020 -1675
rect 7960 -1735 7975 -1705
rect 8005 -1735 8020 -1705
rect 7960 -1770 8020 -1735
rect 7960 -1800 7975 -1770
rect 8005 -1800 8020 -1770
rect 7960 -1840 8020 -1800
rect 7960 -1870 7975 -1840
rect 8005 -1870 8020 -1840
rect 7960 -1910 8020 -1870
rect 7960 -1940 7975 -1910
rect 8005 -1940 8020 -1910
rect 7960 -1980 8020 -1940
rect 7960 -2010 7975 -1980
rect 8005 -2010 8020 -1980
rect 7960 -2045 8020 -2010
rect 7960 -2075 7975 -2045
rect 8005 -2075 8020 -2045
rect 7960 -2105 8020 -2075
rect 7960 -2135 7975 -2105
rect 8005 -2135 8020 -2105
rect 7960 -2170 8020 -2135
rect 7960 -2200 7975 -2170
rect 8005 -2200 8020 -2170
rect 7960 -2240 8020 -2200
rect 7960 -2270 7975 -2240
rect 8005 -2270 8020 -2240
rect 7960 -2310 8020 -2270
rect 7960 -2340 7975 -2310
rect 8005 -2340 8020 -2310
rect 7960 -2380 8020 -2340
rect 7960 -2410 7975 -2380
rect 8005 -2410 8020 -2380
rect 7960 -2445 8020 -2410
rect 7960 -2475 7975 -2445
rect 8005 -2475 8020 -2445
rect 7960 -2505 8020 -2475
rect 7960 -2535 7975 -2505
rect 8005 -2535 8020 -2505
rect 7960 -2570 8020 -2535
rect 7960 -2600 7975 -2570
rect 8005 -2600 8020 -2570
rect 7960 -2640 8020 -2600
rect 7960 -2670 7975 -2640
rect 8005 -2670 8020 -2640
rect 7960 -2710 8020 -2670
rect 7960 -2740 7975 -2710
rect 8005 -2740 8020 -2710
rect 7960 -2780 8020 -2740
rect 7960 -2810 7975 -2780
rect 8005 -2810 8020 -2780
rect 7960 -2845 8020 -2810
rect 7960 -2875 7975 -2845
rect 8005 -2875 8020 -2845
rect 7960 -2890 8020 -2875
rect 8310 -1305 8370 -1290
rect 8310 -1335 8325 -1305
rect 8355 -1335 8370 -1305
rect 8310 -1370 8370 -1335
rect 8310 -1400 8325 -1370
rect 8355 -1400 8370 -1370
rect 8310 -1440 8370 -1400
rect 8310 -1470 8325 -1440
rect 8355 -1470 8370 -1440
rect 8310 -1510 8370 -1470
rect 8310 -1540 8325 -1510
rect 8355 -1540 8370 -1510
rect 8310 -1580 8370 -1540
rect 8310 -1610 8325 -1580
rect 8355 -1610 8370 -1580
rect 8310 -1645 8370 -1610
rect 8310 -1675 8325 -1645
rect 8355 -1675 8370 -1645
rect 8310 -1705 8370 -1675
rect 8310 -1735 8325 -1705
rect 8355 -1735 8370 -1705
rect 8310 -1770 8370 -1735
rect 8310 -1800 8325 -1770
rect 8355 -1800 8370 -1770
rect 8310 -1840 8370 -1800
rect 8310 -1870 8325 -1840
rect 8355 -1870 8370 -1840
rect 8310 -1910 8370 -1870
rect 8310 -1940 8325 -1910
rect 8355 -1940 8370 -1910
rect 8310 -1980 8370 -1940
rect 8310 -2010 8325 -1980
rect 8355 -2010 8370 -1980
rect 8310 -2045 8370 -2010
rect 8310 -2075 8325 -2045
rect 8355 -2075 8370 -2045
rect 8310 -2105 8370 -2075
rect 8310 -2135 8325 -2105
rect 8355 -2135 8370 -2105
rect 8310 -2170 8370 -2135
rect 8310 -2200 8325 -2170
rect 8355 -2200 8370 -2170
rect 8310 -2240 8370 -2200
rect 8310 -2270 8325 -2240
rect 8355 -2270 8370 -2240
rect 8310 -2310 8370 -2270
rect 8310 -2340 8325 -2310
rect 8355 -2340 8370 -2310
rect 8310 -2380 8370 -2340
rect 8310 -2410 8325 -2380
rect 8355 -2410 8370 -2380
rect 8310 -2445 8370 -2410
rect 8310 -2475 8325 -2445
rect 8355 -2475 8370 -2445
rect 8310 -2505 8370 -2475
rect 8310 -2535 8325 -2505
rect 8355 -2535 8370 -2505
rect 8310 -2570 8370 -2535
rect 8310 -2600 8325 -2570
rect 8355 -2600 8370 -2570
rect 8310 -2640 8370 -2600
rect 8310 -2670 8325 -2640
rect 8355 -2670 8370 -2640
rect 8310 -2710 8370 -2670
rect 8310 -2740 8325 -2710
rect 8355 -2740 8370 -2710
rect 8310 -2780 8370 -2740
rect 8310 -2810 8325 -2780
rect 8355 -2810 8370 -2780
rect 8310 -2845 8370 -2810
rect 8310 -2875 8325 -2845
rect 8355 -2875 8370 -2845
rect 8310 -2890 8370 -2875
rect 8660 -1305 8720 -1290
rect 8660 -1335 8675 -1305
rect 8705 -1335 8720 -1305
rect 8660 -1370 8720 -1335
rect 8660 -1400 8675 -1370
rect 8705 -1400 8720 -1370
rect 8660 -1440 8720 -1400
rect 8660 -1470 8675 -1440
rect 8705 -1470 8720 -1440
rect 8660 -1510 8720 -1470
rect 8660 -1540 8675 -1510
rect 8705 -1540 8720 -1510
rect 8660 -1580 8720 -1540
rect 8660 -1610 8675 -1580
rect 8705 -1610 8720 -1580
rect 8660 -1645 8720 -1610
rect 8660 -1675 8675 -1645
rect 8705 -1675 8720 -1645
rect 8660 -1705 8720 -1675
rect 8660 -1735 8675 -1705
rect 8705 -1735 8720 -1705
rect 8660 -1770 8720 -1735
rect 8660 -1800 8675 -1770
rect 8705 -1800 8720 -1770
rect 8660 -1840 8720 -1800
rect 8660 -1870 8675 -1840
rect 8705 -1870 8720 -1840
rect 8660 -1910 8720 -1870
rect 8660 -1940 8675 -1910
rect 8705 -1940 8720 -1910
rect 8660 -1980 8720 -1940
rect 8660 -2010 8675 -1980
rect 8705 -2010 8720 -1980
rect 8660 -2045 8720 -2010
rect 8660 -2075 8675 -2045
rect 8705 -2075 8720 -2045
rect 8660 -2105 8720 -2075
rect 8660 -2135 8675 -2105
rect 8705 -2135 8720 -2105
rect 8660 -2170 8720 -2135
rect 8660 -2200 8675 -2170
rect 8705 -2200 8720 -2170
rect 8660 -2240 8720 -2200
rect 8660 -2270 8675 -2240
rect 8705 -2270 8720 -2240
rect 8660 -2310 8720 -2270
rect 8660 -2340 8675 -2310
rect 8705 -2340 8720 -2310
rect 8660 -2380 8720 -2340
rect 8660 -2410 8675 -2380
rect 8705 -2410 8720 -2380
rect 8660 -2445 8720 -2410
rect 8660 -2475 8675 -2445
rect 8705 -2475 8720 -2445
rect 8660 -2505 8720 -2475
rect 8660 -2535 8675 -2505
rect 8705 -2535 8720 -2505
rect 8660 -2570 8720 -2535
rect 8660 -2600 8675 -2570
rect 8705 -2600 8720 -2570
rect 8660 -2640 8720 -2600
rect 8660 -2670 8675 -2640
rect 8705 -2670 8720 -2640
rect 8660 -2710 8720 -2670
rect 8660 -2740 8675 -2710
rect 8705 -2740 8720 -2710
rect 8660 -2780 8720 -2740
rect 8660 -2810 8675 -2780
rect 8705 -2810 8720 -2780
rect 8660 -2845 8720 -2810
rect 8660 -2875 8675 -2845
rect 8705 -2875 8720 -2845
rect 8660 -2890 8720 -2875
rect 9010 -1305 9070 -1290
rect 9010 -1335 9025 -1305
rect 9055 -1335 9070 -1305
rect 9010 -1370 9070 -1335
rect 9010 -1400 9025 -1370
rect 9055 -1400 9070 -1370
rect 9010 -1440 9070 -1400
rect 9010 -1470 9025 -1440
rect 9055 -1470 9070 -1440
rect 9010 -1510 9070 -1470
rect 9010 -1540 9025 -1510
rect 9055 -1540 9070 -1510
rect 9010 -1580 9070 -1540
rect 9010 -1610 9025 -1580
rect 9055 -1610 9070 -1580
rect 9010 -1645 9070 -1610
rect 9010 -1675 9025 -1645
rect 9055 -1675 9070 -1645
rect 9010 -1705 9070 -1675
rect 9010 -1735 9025 -1705
rect 9055 -1735 9070 -1705
rect 9010 -1770 9070 -1735
rect 9010 -1800 9025 -1770
rect 9055 -1800 9070 -1770
rect 9010 -1840 9070 -1800
rect 9010 -1870 9025 -1840
rect 9055 -1870 9070 -1840
rect 9010 -1910 9070 -1870
rect 9010 -1940 9025 -1910
rect 9055 -1940 9070 -1910
rect 9010 -1980 9070 -1940
rect 9010 -2010 9025 -1980
rect 9055 -2010 9070 -1980
rect 9010 -2045 9070 -2010
rect 9010 -2075 9025 -2045
rect 9055 -2075 9070 -2045
rect 9010 -2105 9070 -2075
rect 9010 -2135 9025 -2105
rect 9055 -2135 9070 -2105
rect 9010 -2170 9070 -2135
rect 9010 -2200 9025 -2170
rect 9055 -2200 9070 -2170
rect 9010 -2240 9070 -2200
rect 9010 -2270 9025 -2240
rect 9055 -2270 9070 -2240
rect 9010 -2310 9070 -2270
rect 9010 -2340 9025 -2310
rect 9055 -2340 9070 -2310
rect 9010 -2380 9070 -2340
rect 9010 -2410 9025 -2380
rect 9055 -2410 9070 -2380
rect 9010 -2445 9070 -2410
rect 9010 -2475 9025 -2445
rect 9055 -2475 9070 -2445
rect 9010 -2505 9070 -2475
rect 9010 -2535 9025 -2505
rect 9055 -2535 9070 -2505
rect 9010 -2570 9070 -2535
rect 9010 -2600 9025 -2570
rect 9055 -2600 9070 -2570
rect 9010 -2640 9070 -2600
rect 9010 -2670 9025 -2640
rect 9055 -2670 9070 -2640
rect 9010 -2710 9070 -2670
rect 9010 -2740 9025 -2710
rect 9055 -2740 9070 -2710
rect 9010 -2780 9070 -2740
rect 9010 -2810 9025 -2780
rect 9055 -2810 9070 -2780
rect 9010 -2845 9070 -2810
rect 9010 -2875 9025 -2845
rect 9055 -2875 9070 -2845
rect 9010 -2890 9070 -2875
<< via2 >>
rect 2115 19280 2145 19310
rect 2115 19215 2145 19245
rect 2115 19145 2145 19175
rect 2115 19075 2145 19105
rect 2115 19005 2145 19035
rect 2115 18940 2145 18970
rect 2115 18880 2145 18910
rect 2115 18815 2145 18845
rect 2115 18745 2145 18775
rect 2115 18675 2145 18705
rect 2115 18605 2145 18635
rect 2115 18540 2145 18570
rect 2115 18480 2145 18510
rect 2115 18415 2145 18445
rect 2115 18345 2145 18375
rect 2115 18275 2145 18305
rect 2115 18205 2145 18235
rect 2115 18140 2145 18170
rect 2115 18080 2145 18110
rect 2115 18015 2145 18045
rect 2115 17945 2145 17975
rect 2115 17875 2145 17905
rect 2115 17805 2145 17835
rect 2115 17740 2145 17770
rect 6705 19280 6735 19310
rect 6705 19215 6735 19245
rect 6705 19145 6735 19175
rect 6705 19075 6735 19105
rect 6705 19005 6735 19035
rect 6705 18940 6735 18970
rect 6705 18880 6735 18910
rect 6705 18815 6735 18845
rect 6705 18745 6735 18775
rect 6705 18675 6735 18705
rect 6705 18605 6735 18635
rect 6705 18540 6735 18570
rect 6705 18480 6735 18510
rect 6705 18415 6735 18445
rect 6705 18345 6735 18375
rect 6705 18275 6735 18305
rect 6705 18205 6735 18235
rect 6705 18140 6735 18170
rect 6705 18080 6735 18110
rect 6705 18015 6735 18045
rect 6705 17945 6735 17975
rect 6705 17875 6735 17905
rect 6705 17805 6735 17835
rect 6705 17740 6735 17770
rect -75 9605 -45 9635
rect -75 9540 -45 9570
rect -75 9470 -45 9500
rect -75 9400 -45 9430
rect -75 9330 -45 9360
rect -75 9265 -45 9295
rect -75 9205 -45 9235
rect -75 9140 -45 9170
rect -75 9070 -45 9100
rect -75 9000 -45 9030
rect -75 8930 -45 8960
rect -75 8865 -45 8895
rect -75 8805 -45 8835
rect -75 8740 -45 8770
rect -75 8670 -45 8700
rect -75 8600 -45 8630
rect -75 8530 -45 8560
rect -75 8465 -45 8495
rect -75 8405 -45 8435
rect -75 8340 -45 8370
rect -75 8270 -45 8300
rect -75 8200 -45 8230
rect -75 8130 -45 8160
rect -75 8065 -45 8095
rect -75 8005 -45 8035
rect -75 7940 -45 7970
rect -75 7870 -45 7900
rect -75 7800 -45 7830
rect -75 7730 -45 7760
rect -75 7665 -45 7695
rect -75 7605 -45 7635
rect -75 7540 -45 7570
rect -75 7470 -45 7500
rect -75 7400 -45 7430
rect -75 7330 -45 7360
rect -75 7265 -45 7295
rect -75 7205 -45 7235
rect -75 7140 -45 7170
rect -75 7070 -45 7100
rect -75 7000 -45 7030
rect -75 6930 -45 6960
rect -75 6865 -45 6895
rect -75 6805 -45 6835
rect -75 6740 -45 6770
rect -75 6670 -45 6700
rect -75 6600 -45 6630
rect -75 6530 -45 6560
rect -75 6465 -45 6495
rect 275 9605 305 9635
rect 275 9540 305 9570
rect 275 9470 305 9500
rect 275 9400 305 9430
rect 275 9330 305 9360
rect 275 9265 305 9295
rect 275 9205 305 9235
rect 275 9140 305 9170
rect 275 9070 305 9100
rect 275 9000 305 9030
rect 275 8930 305 8960
rect 275 8865 305 8895
rect 275 8805 305 8835
rect 275 8740 305 8770
rect 275 8670 305 8700
rect 275 8600 305 8630
rect 275 8530 305 8560
rect 275 8465 305 8495
rect 275 8405 305 8435
rect 275 8340 305 8370
rect 275 8270 305 8300
rect 275 8200 305 8230
rect 275 8130 305 8160
rect 275 8065 305 8095
rect 275 8005 305 8035
rect 275 7940 305 7970
rect 275 7870 305 7900
rect 275 7800 305 7830
rect 275 7730 305 7760
rect 275 7665 305 7695
rect 275 7605 305 7635
rect 275 7540 305 7570
rect 275 7470 305 7500
rect 275 7400 305 7430
rect 275 7330 305 7360
rect 275 7265 305 7295
rect 275 7205 305 7235
rect 275 7140 305 7170
rect 275 7070 305 7100
rect 275 7000 305 7030
rect 275 6930 305 6960
rect 275 6865 305 6895
rect 275 6805 305 6835
rect 275 6740 305 6770
rect 275 6670 305 6700
rect 275 6600 305 6630
rect 275 6530 305 6560
rect 275 6465 305 6495
rect 625 9605 655 9635
rect 625 9540 655 9570
rect 625 9470 655 9500
rect 625 9400 655 9430
rect 625 9330 655 9360
rect 625 9265 655 9295
rect 625 9205 655 9235
rect 625 9140 655 9170
rect 625 9070 655 9100
rect 625 9000 655 9030
rect 625 8930 655 8960
rect 625 8865 655 8895
rect 625 8805 655 8835
rect 625 8740 655 8770
rect 625 8670 655 8700
rect 625 8600 655 8630
rect 625 8530 655 8560
rect 625 8465 655 8495
rect 625 8405 655 8435
rect 625 8340 655 8370
rect 625 8270 655 8300
rect 625 8200 655 8230
rect 625 8130 655 8160
rect 625 8065 655 8095
rect 625 8005 655 8035
rect 625 7940 655 7970
rect 625 7870 655 7900
rect 625 7800 655 7830
rect 625 7730 655 7760
rect 625 7665 655 7695
rect 625 7605 655 7635
rect 625 7540 655 7570
rect 625 7470 655 7500
rect 625 7400 655 7430
rect 625 7330 655 7360
rect 625 7265 655 7295
rect 625 7205 655 7235
rect 625 7140 655 7170
rect 625 7070 655 7100
rect 625 7000 655 7030
rect 625 6930 655 6960
rect 625 6865 655 6895
rect 625 6805 655 6835
rect 625 6740 655 6770
rect 625 6670 655 6700
rect 625 6600 655 6630
rect 625 6530 655 6560
rect 625 6465 655 6495
rect 975 9605 1005 9635
rect 975 9540 1005 9570
rect 975 9470 1005 9500
rect 975 9400 1005 9430
rect 975 9330 1005 9360
rect 975 9265 1005 9295
rect 975 9205 1005 9235
rect 975 9140 1005 9170
rect 975 9070 1005 9100
rect 975 9000 1005 9030
rect 975 8930 1005 8960
rect 975 8865 1005 8895
rect 975 8805 1005 8835
rect 975 8740 1005 8770
rect 975 8670 1005 8700
rect 975 8600 1005 8630
rect 975 8530 1005 8560
rect 975 8465 1005 8495
rect 975 8405 1005 8435
rect 975 8340 1005 8370
rect 975 8270 1005 8300
rect 975 8200 1005 8230
rect 975 8130 1005 8160
rect 975 8065 1005 8095
rect 975 8005 1005 8035
rect 975 7940 1005 7970
rect 975 7870 1005 7900
rect 975 7800 1005 7830
rect 975 7730 1005 7760
rect 975 7665 1005 7695
rect 975 7605 1005 7635
rect 975 7540 1005 7570
rect 975 7470 1005 7500
rect 975 7400 1005 7430
rect 975 7330 1005 7360
rect 975 7265 1005 7295
rect 975 7205 1005 7235
rect 975 7140 1005 7170
rect 975 7070 1005 7100
rect 975 7000 1005 7030
rect 975 6930 1005 6960
rect 975 6865 1005 6895
rect 975 6805 1005 6835
rect 975 6740 1005 6770
rect 975 6670 1005 6700
rect 975 6600 1005 6630
rect 975 6530 1005 6560
rect 975 6465 1005 6495
rect 1675 9605 1705 9635
rect 1675 9540 1705 9570
rect 1675 9470 1705 9500
rect 1675 9400 1705 9430
rect 1675 9330 1705 9360
rect 1675 9265 1705 9295
rect 1675 9205 1705 9235
rect 1675 9140 1705 9170
rect 1675 9070 1705 9100
rect 1675 9000 1705 9030
rect 1675 8930 1705 8960
rect 1675 8865 1705 8895
rect 1675 8805 1705 8835
rect 1675 8740 1705 8770
rect 1675 8670 1705 8700
rect 1675 8600 1705 8630
rect 1675 8530 1705 8560
rect 1675 8465 1705 8495
rect 1675 8405 1705 8435
rect 1675 8340 1705 8370
rect 1675 8270 1705 8300
rect 1675 8200 1705 8230
rect 1675 8130 1705 8160
rect 1675 8065 1705 8095
rect 1675 8005 1705 8035
rect 1675 7940 1705 7970
rect 1675 7870 1705 7900
rect 1675 7800 1705 7830
rect 1675 7730 1705 7760
rect 1675 7665 1705 7695
rect 1675 7605 1705 7635
rect 1675 7540 1705 7570
rect 1675 7470 1705 7500
rect 1675 7400 1705 7430
rect 1675 7330 1705 7360
rect 1675 7265 1705 7295
rect 1675 7205 1705 7235
rect 1675 7140 1705 7170
rect 1675 7070 1705 7100
rect 1675 7000 1705 7030
rect 1675 6930 1705 6960
rect 1675 6865 1705 6895
rect 1675 6805 1705 6835
rect 1675 6740 1705 6770
rect 1675 6670 1705 6700
rect 1675 6600 1705 6630
rect 1675 6530 1705 6560
rect 1675 6465 1705 6495
rect 2250 9605 2280 9635
rect 2250 9540 2280 9570
rect 2250 9470 2280 9500
rect 2250 9400 2280 9430
rect 2250 9330 2280 9360
rect 2250 9265 2280 9295
rect 2250 9205 2280 9235
rect 2250 9140 2280 9170
rect 2250 9070 2280 9100
rect 2250 9000 2280 9030
rect 2250 8930 2280 8960
rect 2250 8865 2280 8895
rect 2250 8805 2280 8835
rect 2250 8740 2280 8770
rect 2250 8670 2280 8700
rect 2250 8600 2280 8630
rect 2250 8530 2280 8560
rect 2250 8465 2280 8495
rect 2250 8405 2280 8435
rect 2250 8340 2280 8370
rect 2250 8270 2280 8300
rect 2250 8200 2280 8230
rect 2250 8130 2280 8160
rect 2250 8065 2280 8095
rect 2250 8005 2280 8035
rect 2250 7940 2280 7970
rect 2250 7870 2280 7900
rect 2250 7800 2280 7830
rect 2250 7730 2280 7760
rect 2250 7665 2280 7695
rect 2250 7605 2280 7635
rect 2250 7540 2280 7570
rect 2250 7470 2280 7500
rect 2250 7400 2280 7430
rect 2250 7330 2280 7360
rect 2250 7265 2280 7295
rect 2250 7205 2280 7235
rect 2250 7140 2280 7170
rect 2250 7070 2280 7100
rect 2250 7000 2280 7030
rect 2250 6930 2280 6960
rect 2250 6865 2280 6895
rect 2250 6805 2280 6835
rect 2250 6740 2280 6770
rect 2250 6670 2280 6700
rect 2250 6600 2280 6630
rect 2250 6530 2280 6560
rect 2250 6465 2280 6495
rect 3180 9605 3210 9635
rect 3240 9605 3270 9635
rect 3180 9540 3210 9570
rect 3240 9540 3270 9570
rect 3180 9470 3210 9500
rect 3240 9470 3270 9500
rect 3180 9400 3210 9430
rect 3240 9400 3270 9430
rect 3180 9330 3210 9360
rect 3240 9330 3270 9360
rect 3180 9265 3210 9295
rect 3240 9265 3270 9295
rect 3180 9205 3210 9235
rect 3240 9205 3270 9235
rect 3180 9140 3210 9170
rect 3240 9140 3270 9170
rect 3180 9070 3210 9100
rect 3240 9070 3270 9100
rect 3180 9000 3210 9030
rect 3240 9000 3270 9030
rect 3180 8930 3210 8960
rect 3240 8930 3270 8960
rect 3180 8865 3210 8895
rect 3240 8865 3270 8895
rect 3180 8805 3210 8835
rect 3240 8805 3270 8835
rect 3180 8740 3210 8770
rect 3240 8740 3270 8770
rect 3180 8670 3210 8700
rect 3240 8670 3270 8700
rect 3180 8600 3210 8630
rect 3240 8600 3270 8630
rect 3180 8530 3210 8560
rect 3240 8530 3270 8560
rect 3180 8465 3210 8495
rect 3240 8465 3270 8495
rect 3180 8405 3210 8435
rect 3240 8405 3270 8435
rect 3180 8340 3210 8370
rect 3240 8340 3270 8370
rect 3180 8270 3210 8300
rect 3240 8270 3270 8300
rect 3180 8200 3210 8230
rect 3240 8200 3270 8230
rect 3180 8130 3210 8160
rect 3240 8130 3270 8160
rect 3180 8065 3210 8095
rect 3240 8065 3270 8095
rect 3180 8005 3210 8035
rect 3240 8005 3270 8035
rect 3180 7940 3210 7970
rect 3240 7940 3270 7970
rect 3180 7870 3210 7900
rect 3240 7870 3270 7900
rect 3180 7800 3210 7830
rect 3240 7800 3270 7830
rect 3180 7730 3210 7760
rect 3240 7730 3270 7760
rect 3180 7665 3210 7695
rect 3240 7665 3270 7695
rect 3180 7605 3210 7635
rect 3240 7605 3270 7635
rect 3180 7540 3210 7570
rect 3240 7540 3270 7570
rect 3180 7470 3210 7500
rect 3240 7470 3270 7500
rect 3180 7400 3210 7430
rect 3240 7400 3270 7430
rect 3180 7330 3210 7360
rect 3240 7330 3270 7360
rect 3180 7265 3210 7295
rect 3240 7265 3270 7295
rect 3180 7205 3210 7235
rect 3240 7205 3270 7235
rect 3180 7140 3210 7170
rect 3240 7140 3270 7170
rect 3180 7070 3210 7100
rect 3240 7070 3270 7100
rect 3180 7000 3210 7030
rect 3240 7000 3270 7030
rect 3180 6930 3210 6960
rect 3240 6930 3270 6960
rect 3180 6865 3210 6895
rect 3240 6865 3270 6895
rect 3180 6805 3210 6835
rect 3240 6805 3270 6835
rect 3180 6740 3210 6770
rect 3240 6740 3270 6770
rect 3180 6670 3210 6700
rect 3240 6670 3270 6700
rect 3180 6600 3210 6630
rect 3240 6600 3270 6630
rect 3180 6530 3210 6560
rect 3240 6530 3270 6560
rect 3180 6465 3210 6495
rect 3240 6465 3270 6495
rect 3350 9605 3380 9635
rect 3350 9540 3380 9570
rect 3350 9470 3380 9500
rect 3350 9400 3380 9430
rect 3350 9330 3380 9360
rect 3350 9265 3380 9295
rect 3350 9205 3380 9235
rect 3350 9140 3380 9170
rect 3350 9070 3380 9100
rect 3350 9000 3380 9030
rect 3350 8930 3380 8960
rect 3350 8865 3380 8895
rect 3350 8805 3380 8835
rect 3350 8740 3380 8770
rect 3350 8670 3380 8700
rect 3350 8600 3380 8630
rect 3350 8530 3380 8560
rect 3350 8465 3380 8495
rect 3350 8405 3380 8435
rect 3350 8340 3380 8370
rect 3350 8270 3380 8300
rect 3350 8200 3380 8230
rect 3350 8130 3380 8160
rect 3350 8065 3380 8095
rect 3350 8005 3380 8035
rect 3350 7940 3380 7970
rect 3350 7870 3380 7900
rect 3350 7800 3380 7830
rect 3350 7730 3380 7760
rect 3350 7665 3380 7695
rect 3350 7605 3380 7635
rect 3350 7540 3380 7570
rect 3350 7470 3380 7500
rect 3350 7400 3380 7430
rect 3350 7330 3380 7360
rect 3350 7265 3380 7295
rect 3350 7205 3380 7235
rect 3350 7140 3380 7170
rect 3350 7070 3380 7100
rect 3350 7000 3380 7030
rect 3350 6930 3380 6960
rect 3350 6865 3380 6895
rect 3350 6805 3380 6835
rect 3350 6740 3380 6770
rect 3350 6670 3380 6700
rect 3350 6600 3380 6630
rect 3350 6530 3380 6560
rect 3350 6465 3380 6495
rect 6705 9605 6735 9635
rect 6705 9540 6735 9570
rect 6705 9470 6735 9500
rect 6705 9400 6735 9430
rect 6705 9330 6735 9360
rect 6705 9265 6735 9295
rect 6705 9205 6735 9235
rect 6705 9140 6735 9170
rect 6705 9070 6735 9100
rect 6705 9000 6735 9030
rect 6705 8930 6735 8960
rect 6705 8865 6735 8895
rect 6705 8805 6735 8835
rect 6705 8740 6735 8770
rect 6705 8670 6735 8700
rect 6705 8600 6735 8630
rect 6705 8530 6735 8560
rect 6705 8465 6735 8495
rect 6705 8405 6735 8435
rect 6705 8340 6735 8370
rect 6705 8270 6735 8300
rect 6705 8200 6735 8230
rect 6705 8130 6735 8160
rect 6705 8065 6735 8095
rect 6705 8005 6735 8035
rect 6705 7940 6735 7970
rect 6705 7870 6735 7900
rect 6705 7800 6735 7830
rect 6705 7730 6735 7760
rect 6705 7665 6735 7695
rect 6705 7605 6735 7635
rect 6705 7540 6735 7570
rect 6705 7470 6735 7500
rect 6705 7400 6735 7430
rect 6705 7330 6735 7360
rect 6705 7265 6735 7295
rect 6705 7205 6735 7235
rect 6705 7140 6735 7170
rect 6705 7070 6735 7100
rect 6705 7000 6735 7030
rect 6705 6930 6735 6960
rect 6705 6865 6735 6895
rect 6705 6805 6735 6835
rect 6705 6740 6735 6770
rect 6705 6670 6735 6700
rect 6705 6600 6735 6630
rect 6705 6530 6735 6560
rect 6705 6465 6735 6495
rect 7275 9605 7305 9635
rect 7275 9540 7305 9570
rect 7275 9470 7305 9500
rect 7275 9400 7305 9430
rect 7275 9330 7305 9360
rect 7275 9265 7305 9295
rect 7275 9205 7305 9235
rect 7275 9140 7305 9170
rect 7275 9070 7305 9100
rect 7275 9000 7305 9030
rect 7275 8930 7305 8960
rect 7275 8865 7305 8895
rect 7275 8805 7305 8835
rect 7275 8740 7305 8770
rect 7275 8670 7305 8700
rect 7275 8600 7305 8630
rect 7275 8530 7305 8560
rect 7275 8465 7305 8495
rect 7275 8405 7305 8435
rect 7275 8340 7305 8370
rect 7275 8270 7305 8300
rect 7275 8200 7305 8230
rect 7275 8130 7305 8160
rect 7275 8065 7305 8095
rect 7275 8005 7305 8035
rect 7275 7940 7305 7970
rect 7275 7870 7305 7900
rect 7275 7800 7305 7830
rect 7275 7730 7305 7760
rect 7275 7665 7305 7695
rect 7275 7605 7305 7635
rect 7275 7540 7305 7570
rect 7275 7470 7305 7500
rect 7275 7400 7305 7430
rect 7275 7330 7305 7360
rect 7275 7265 7305 7295
rect 7275 7205 7305 7235
rect 7275 7140 7305 7170
rect 7275 7070 7305 7100
rect 7275 7000 7305 7030
rect 7275 6930 7305 6960
rect 7275 6865 7305 6895
rect 7275 6805 7305 6835
rect 7275 6740 7305 6770
rect 7275 6670 7305 6700
rect 7275 6600 7305 6630
rect 7275 6530 7305 6560
rect 7275 6465 7305 6495
rect 7975 9605 8005 9635
rect 7975 9540 8005 9570
rect 7975 9470 8005 9500
rect 7975 9400 8005 9430
rect 7975 9330 8005 9360
rect 7975 9265 8005 9295
rect 7975 9205 8005 9235
rect 7975 9140 8005 9170
rect 7975 9070 8005 9100
rect 7975 9000 8005 9030
rect 7975 8930 8005 8960
rect 7975 8865 8005 8895
rect 7975 8805 8005 8835
rect 7975 8740 8005 8770
rect 7975 8670 8005 8700
rect 7975 8600 8005 8630
rect 7975 8530 8005 8560
rect 7975 8465 8005 8495
rect 7975 8405 8005 8435
rect 7975 8340 8005 8370
rect 7975 8270 8005 8300
rect 7975 8200 8005 8230
rect 7975 8130 8005 8160
rect 7975 8065 8005 8095
rect 7975 8005 8005 8035
rect 7975 7940 8005 7970
rect 7975 7870 8005 7900
rect 7975 7800 8005 7830
rect 7975 7730 8005 7760
rect 7975 7665 8005 7695
rect 7975 7605 8005 7635
rect 7975 7540 8005 7570
rect 7975 7470 8005 7500
rect 7975 7400 8005 7430
rect 7975 7330 8005 7360
rect 7975 7265 8005 7295
rect 7975 7205 8005 7235
rect 7975 7140 8005 7170
rect 7975 7070 8005 7100
rect 7975 7000 8005 7030
rect 7975 6930 8005 6960
rect 7975 6865 8005 6895
rect 7975 6805 8005 6835
rect 7975 6740 8005 6770
rect 7975 6670 8005 6700
rect 7975 6600 8005 6630
rect 7975 6530 8005 6560
rect 7975 6465 8005 6495
rect 8325 9605 8355 9635
rect 8325 9540 8355 9570
rect 8325 9470 8355 9500
rect 8325 9400 8355 9430
rect 8325 9330 8355 9360
rect 8325 9265 8355 9295
rect 8325 9205 8355 9235
rect 8325 9140 8355 9170
rect 8325 9070 8355 9100
rect 8325 9000 8355 9030
rect 8325 8930 8355 8960
rect 8325 8865 8355 8895
rect 8325 8805 8355 8835
rect 8325 8740 8355 8770
rect 8325 8670 8355 8700
rect 8325 8600 8355 8630
rect 8325 8530 8355 8560
rect 8325 8465 8355 8495
rect 8325 8405 8355 8435
rect 8325 8340 8355 8370
rect 8325 8270 8355 8300
rect 8325 8200 8355 8230
rect 8325 8130 8355 8160
rect 8325 8065 8355 8095
rect 8325 8005 8355 8035
rect 8325 7940 8355 7970
rect 8325 7870 8355 7900
rect 8325 7800 8355 7830
rect 8325 7730 8355 7760
rect 8325 7665 8355 7695
rect 8325 7605 8355 7635
rect 8325 7540 8355 7570
rect 8325 7470 8355 7500
rect 8325 7400 8355 7430
rect 8325 7330 8355 7360
rect 8325 7265 8355 7295
rect 8325 7205 8355 7235
rect 8325 7140 8355 7170
rect 8325 7070 8355 7100
rect 8325 7000 8355 7030
rect 8325 6930 8355 6960
rect 8325 6865 8355 6895
rect 8325 6805 8355 6835
rect 8325 6740 8355 6770
rect 8325 6670 8355 6700
rect 8325 6600 8355 6630
rect 8325 6530 8355 6560
rect 8325 6465 8355 6495
rect 8675 9605 8705 9635
rect 8675 9540 8705 9570
rect 8675 9470 8705 9500
rect 8675 9400 8705 9430
rect 8675 9330 8705 9360
rect 8675 9265 8705 9295
rect 8675 9205 8705 9235
rect 8675 9140 8705 9170
rect 8675 9070 8705 9100
rect 8675 9000 8705 9030
rect 8675 8930 8705 8960
rect 8675 8865 8705 8895
rect 8675 8805 8705 8835
rect 8675 8740 8705 8770
rect 8675 8670 8705 8700
rect 8675 8600 8705 8630
rect 8675 8530 8705 8560
rect 8675 8465 8705 8495
rect 8675 8405 8705 8435
rect 8675 8340 8705 8370
rect 8675 8270 8705 8300
rect 8675 8200 8705 8230
rect 8675 8130 8705 8160
rect 8675 8065 8705 8095
rect 8675 8005 8705 8035
rect 8675 7940 8705 7970
rect 8675 7870 8705 7900
rect 8675 7800 8705 7830
rect 8675 7730 8705 7760
rect 8675 7665 8705 7695
rect 8675 7605 8705 7635
rect 8675 7540 8705 7570
rect 8675 7470 8705 7500
rect 8675 7400 8705 7430
rect 8675 7330 8705 7360
rect 8675 7265 8705 7295
rect 8675 7205 8705 7235
rect 8675 7140 8705 7170
rect 8675 7070 8705 7100
rect 8675 7000 8705 7030
rect 8675 6930 8705 6960
rect 8675 6865 8705 6895
rect 8675 6805 8705 6835
rect 8675 6740 8705 6770
rect 8675 6670 8705 6700
rect 8675 6600 8705 6630
rect 8675 6530 8705 6560
rect 8675 6465 8705 6495
rect 9025 9605 9055 9635
rect 9025 9540 9055 9570
rect 9025 9470 9055 9500
rect 9025 9400 9055 9430
rect 9025 9330 9055 9360
rect 9025 9265 9055 9295
rect 9025 9205 9055 9235
rect 9025 9140 9055 9170
rect 9025 9070 9055 9100
rect 9025 9000 9055 9030
rect 9025 8930 9055 8960
rect 9025 8865 9055 8895
rect 9025 8805 9055 8835
rect 9025 8740 9055 8770
rect 9025 8670 9055 8700
rect 9025 8600 9055 8630
rect 9025 8530 9055 8560
rect 9025 8465 9055 8495
rect 9025 8405 9055 8435
rect 9025 8340 9055 8370
rect 9025 8270 9055 8300
rect 9025 8200 9055 8230
rect 9025 8130 9055 8160
rect 9025 8065 9055 8095
rect 9025 8005 9055 8035
rect 9025 7940 9055 7970
rect 9025 7870 9055 7900
rect 9025 7800 9055 7830
rect 9025 7730 9055 7760
rect 9025 7665 9055 7695
rect 9025 7605 9055 7635
rect 9025 7540 9055 7570
rect 9025 7470 9055 7500
rect 9025 7400 9055 7430
rect 9025 7330 9055 7360
rect 9025 7265 9055 7295
rect 9025 7205 9055 7235
rect 9025 7140 9055 7170
rect 9025 7070 9055 7100
rect 9025 7000 9055 7030
rect 9025 6930 9055 6960
rect 9025 6865 9055 6895
rect 9025 6805 9055 6835
rect 9025 6740 9055 6770
rect 9025 6670 9055 6700
rect 9025 6600 9055 6630
rect 9025 6530 9055 6560
rect 9025 6465 9055 6495
rect -75 -1335 -45 -1305
rect -75 -1400 -45 -1370
rect -75 -1470 -45 -1440
rect -75 -1540 -45 -1510
rect -75 -1610 -45 -1580
rect -75 -1675 -45 -1645
rect -75 -1735 -45 -1705
rect -75 -1800 -45 -1770
rect -75 -1870 -45 -1840
rect -75 -1940 -45 -1910
rect -75 -2010 -45 -1980
rect -75 -2075 -45 -2045
rect -75 -2135 -45 -2105
rect -75 -2200 -45 -2170
rect -75 -2270 -45 -2240
rect -75 -2340 -45 -2310
rect -75 -2410 -45 -2380
rect -75 -2475 -45 -2445
rect -75 -2535 -45 -2505
rect -75 -2600 -45 -2570
rect -75 -2670 -45 -2640
rect -75 -2740 -45 -2710
rect -75 -2810 -45 -2780
rect -75 -2875 -45 -2845
rect 275 -1335 305 -1305
rect 275 -1400 305 -1370
rect 275 -1470 305 -1440
rect 275 -1540 305 -1510
rect 275 -1610 305 -1580
rect 275 -1675 305 -1645
rect 275 -1735 305 -1705
rect 275 -1800 305 -1770
rect 275 -1870 305 -1840
rect 275 -1940 305 -1910
rect 275 -2010 305 -1980
rect 275 -2075 305 -2045
rect 275 -2135 305 -2105
rect 275 -2200 305 -2170
rect 275 -2270 305 -2240
rect 275 -2340 305 -2310
rect 275 -2410 305 -2380
rect 275 -2475 305 -2445
rect 275 -2535 305 -2505
rect 275 -2600 305 -2570
rect 275 -2670 305 -2640
rect 275 -2740 305 -2710
rect 275 -2810 305 -2780
rect 275 -2875 305 -2845
rect 625 -1335 655 -1305
rect 625 -1400 655 -1370
rect 625 -1470 655 -1440
rect 625 -1540 655 -1510
rect 625 -1610 655 -1580
rect 625 -1675 655 -1645
rect 625 -1735 655 -1705
rect 625 -1800 655 -1770
rect 625 -1870 655 -1840
rect 625 -1940 655 -1910
rect 625 -2010 655 -1980
rect 625 -2075 655 -2045
rect 625 -2135 655 -2105
rect 625 -2200 655 -2170
rect 625 -2270 655 -2240
rect 625 -2340 655 -2310
rect 625 -2410 655 -2380
rect 625 -2475 655 -2445
rect 625 -2535 655 -2505
rect 625 -2600 655 -2570
rect 625 -2670 655 -2640
rect 625 -2740 655 -2710
rect 625 -2810 655 -2780
rect 625 -2875 655 -2845
rect 975 -1335 1005 -1305
rect 975 -1400 1005 -1370
rect 975 -1470 1005 -1440
rect 975 -1540 1005 -1510
rect 975 -1610 1005 -1580
rect 975 -1675 1005 -1645
rect 975 -1735 1005 -1705
rect 975 -1800 1005 -1770
rect 975 -1870 1005 -1840
rect 975 -1940 1005 -1910
rect 975 -2010 1005 -1980
rect 975 -2075 1005 -2045
rect 975 -2135 1005 -2105
rect 975 -2200 1005 -2170
rect 975 -2270 1005 -2240
rect 975 -2340 1005 -2310
rect 975 -2410 1005 -2380
rect 975 -2475 1005 -2445
rect 975 -2535 1005 -2505
rect 975 -2600 1005 -2570
rect 975 -2670 1005 -2640
rect 975 -2740 1005 -2710
rect 975 -2810 1005 -2780
rect 975 -2875 1005 -2845
rect 1325 -1335 1355 -1305
rect 1325 -1400 1355 -1370
rect 1325 -1470 1355 -1440
rect 1325 -1540 1355 -1510
rect 1325 -1610 1355 -1580
rect 1325 -1675 1355 -1645
rect 1325 -1735 1355 -1705
rect 1325 -1800 1355 -1770
rect 1325 -1870 1355 -1840
rect 1325 -1940 1355 -1910
rect 1325 -2010 1355 -1980
rect 1325 -2075 1355 -2045
rect 1325 -2135 1355 -2105
rect 1325 -2200 1355 -2170
rect 1325 -2270 1355 -2240
rect 1325 -2340 1355 -2310
rect 1325 -2410 1355 -2380
rect 1325 -2475 1355 -2445
rect 1325 -2535 1355 -2505
rect 1325 -2600 1355 -2570
rect 1325 -2670 1355 -2640
rect 1325 -2740 1355 -2710
rect 1325 -2810 1355 -2780
rect 1325 -2875 1355 -2845
rect 1675 -1335 1705 -1305
rect 1675 -1400 1705 -1370
rect 1675 -1470 1705 -1440
rect 1675 -1540 1705 -1510
rect 1675 -1610 1705 -1580
rect 1675 -1675 1705 -1645
rect 1675 -1735 1705 -1705
rect 1675 -1800 1705 -1770
rect 1675 -1870 1705 -1840
rect 1675 -1940 1705 -1910
rect 1675 -2010 1705 -1980
rect 1675 -2075 1705 -2045
rect 1675 -2135 1705 -2105
rect 1675 -2200 1705 -2170
rect 1675 -2270 1705 -2240
rect 1675 -2340 1705 -2310
rect 1675 -2410 1705 -2380
rect 1675 -2475 1705 -2445
rect 1675 -2535 1705 -2505
rect 1675 -2600 1705 -2570
rect 1675 -2670 1705 -2640
rect 1675 -2740 1705 -2710
rect 1675 -2810 1705 -2780
rect 1675 -2875 1705 -2845
rect 2025 -1335 2055 -1305
rect 2025 -1400 2055 -1370
rect 2025 -1470 2055 -1440
rect 2025 -1540 2055 -1510
rect 2025 -1610 2055 -1580
rect 2025 -1675 2055 -1645
rect 2025 -1735 2055 -1705
rect 2025 -1800 2055 -1770
rect 2025 -1870 2055 -1840
rect 2025 -1940 2055 -1910
rect 2025 -2010 2055 -1980
rect 2025 -2075 2055 -2045
rect 2025 -2135 2055 -2105
rect 2025 -2200 2055 -2170
rect 2025 -2270 2055 -2240
rect 2025 -2340 2055 -2310
rect 2025 -2410 2055 -2380
rect 2025 -2475 2055 -2445
rect 2025 -2535 2055 -2505
rect 2025 -2600 2055 -2570
rect 2025 -2670 2055 -2640
rect 2025 -2740 2055 -2710
rect 2025 -2810 2055 -2780
rect 2025 -2875 2055 -2845
rect 2375 -1335 2405 -1305
rect 2375 -1400 2405 -1370
rect 2375 -1470 2405 -1440
rect 2375 -1540 2405 -1510
rect 2375 -1610 2405 -1580
rect 2375 -1675 2405 -1645
rect 2375 -1735 2405 -1705
rect 2375 -1800 2405 -1770
rect 2375 -1870 2405 -1840
rect 2375 -1940 2405 -1910
rect 2375 -2010 2405 -1980
rect 2375 -2075 2405 -2045
rect 2375 -2135 2405 -2105
rect 2375 -2200 2405 -2170
rect 2375 -2270 2405 -2240
rect 2375 -2340 2405 -2310
rect 2375 -2410 2405 -2380
rect 2375 -2475 2405 -2445
rect 2375 -2535 2405 -2505
rect 2375 -2600 2405 -2570
rect 2375 -2670 2405 -2640
rect 2375 -2740 2405 -2710
rect 2375 -2810 2405 -2780
rect 2375 -2875 2405 -2845
rect 2725 -1335 2755 -1305
rect 2725 -1400 2755 -1370
rect 2725 -1470 2755 -1440
rect 2725 -1540 2755 -1510
rect 2725 -1610 2755 -1580
rect 2725 -1675 2755 -1645
rect 2725 -1735 2755 -1705
rect 2725 -1800 2755 -1770
rect 2725 -1870 2755 -1840
rect 2725 -1940 2755 -1910
rect 2725 -2010 2755 -1980
rect 2725 -2075 2755 -2045
rect 2725 -2135 2755 -2105
rect 2725 -2200 2755 -2170
rect 2725 -2270 2755 -2240
rect 2725 -2340 2755 -2310
rect 2725 -2410 2755 -2380
rect 2725 -2475 2755 -2445
rect 2725 -2535 2755 -2505
rect 2725 -2600 2755 -2570
rect 2725 -2670 2755 -2640
rect 2725 -2740 2755 -2710
rect 2725 -2810 2755 -2780
rect 2725 -2875 2755 -2845
rect 3075 -1335 3105 -1305
rect 3075 -1400 3105 -1370
rect 3075 -1470 3105 -1440
rect 3075 -1540 3105 -1510
rect 3075 -1610 3105 -1580
rect 3075 -1675 3105 -1645
rect 3075 -1735 3105 -1705
rect 3075 -1800 3105 -1770
rect 3075 -1870 3105 -1840
rect 3075 -1940 3105 -1910
rect 3075 -2010 3105 -1980
rect 3075 -2075 3105 -2045
rect 3075 -2135 3105 -2105
rect 3075 -2200 3105 -2170
rect 3075 -2270 3105 -2240
rect 3075 -2340 3105 -2310
rect 3075 -2410 3105 -2380
rect 3075 -2475 3105 -2445
rect 3075 -2535 3105 -2505
rect 3075 -2600 3105 -2570
rect 3075 -2670 3105 -2640
rect 3075 -2740 3105 -2710
rect 3075 -2810 3105 -2780
rect 3075 -2875 3105 -2845
rect 3425 -1335 3455 -1305
rect 3425 -1400 3455 -1370
rect 3425 -1470 3455 -1440
rect 3425 -1540 3455 -1510
rect 3425 -1610 3455 -1580
rect 3425 -1675 3455 -1645
rect 3425 -1735 3455 -1705
rect 3425 -1800 3455 -1770
rect 3425 -1870 3455 -1840
rect 3425 -1940 3455 -1910
rect 3425 -2010 3455 -1980
rect 3425 -2075 3455 -2045
rect 3425 -2135 3455 -2105
rect 3425 -2200 3455 -2170
rect 3425 -2270 3455 -2240
rect 3425 -2340 3455 -2310
rect 3425 -2410 3455 -2380
rect 3425 -2475 3455 -2445
rect 3425 -2535 3455 -2505
rect 3425 -2600 3455 -2570
rect 3425 -2670 3455 -2640
rect 3425 -2740 3455 -2710
rect 3425 -2810 3455 -2780
rect 3425 -2875 3455 -2845
rect 3775 -1335 3805 -1305
rect 3775 -1400 3805 -1370
rect 3775 -1470 3805 -1440
rect 3775 -1540 3805 -1510
rect 3775 -1610 3805 -1580
rect 3775 -1675 3805 -1645
rect 3775 -1735 3805 -1705
rect 3775 -1800 3805 -1770
rect 3775 -1870 3805 -1840
rect 3775 -1940 3805 -1910
rect 3775 -2010 3805 -1980
rect 3775 -2075 3805 -2045
rect 3775 -2135 3805 -2105
rect 3775 -2200 3805 -2170
rect 3775 -2270 3805 -2240
rect 3775 -2340 3805 -2310
rect 3775 -2410 3805 -2380
rect 3775 -2475 3805 -2445
rect 3775 -2535 3805 -2505
rect 3775 -2600 3805 -2570
rect 3775 -2670 3805 -2640
rect 3775 -2740 3805 -2710
rect 3775 -2810 3805 -2780
rect 3775 -2875 3805 -2845
rect 4125 -1335 4155 -1305
rect 4125 -1400 4155 -1370
rect 4125 -1470 4155 -1440
rect 4125 -1540 4155 -1510
rect 4125 -1610 4155 -1580
rect 4125 -1675 4155 -1645
rect 4125 -1735 4155 -1705
rect 4125 -1800 4155 -1770
rect 4125 -1870 4155 -1840
rect 4125 -1940 4155 -1910
rect 4125 -2010 4155 -1980
rect 4125 -2075 4155 -2045
rect 4125 -2135 4155 -2105
rect 4125 -2200 4155 -2170
rect 4125 -2270 4155 -2240
rect 4125 -2340 4155 -2310
rect 4125 -2410 4155 -2380
rect 4125 -2475 4155 -2445
rect 4125 -2535 4155 -2505
rect 4125 -2600 4155 -2570
rect 4125 -2670 4155 -2640
rect 4125 -2740 4155 -2710
rect 4125 -2810 4155 -2780
rect 4125 -2875 4155 -2845
rect 4475 -1335 4505 -1305
rect 4475 -1400 4505 -1370
rect 4475 -1470 4505 -1440
rect 4475 -1540 4505 -1510
rect 4475 -1610 4505 -1580
rect 4475 -1675 4505 -1645
rect 4475 -1735 4505 -1705
rect 4475 -1800 4505 -1770
rect 4475 -1870 4505 -1840
rect 4475 -1940 4505 -1910
rect 4475 -2010 4505 -1980
rect 4475 -2075 4505 -2045
rect 4475 -2135 4505 -2105
rect 4475 -2200 4505 -2170
rect 4475 -2270 4505 -2240
rect 4475 -2340 4505 -2310
rect 4475 -2410 4505 -2380
rect 4475 -2475 4505 -2445
rect 4475 -2535 4505 -2505
rect 4475 -2600 4505 -2570
rect 4475 -2670 4505 -2640
rect 4475 -2740 4505 -2710
rect 4475 -2810 4505 -2780
rect 4475 -2875 4505 -2845
rect 4825 -1335 4855 -1305
rect 4825 -1400 4855 -1370
rect 4825 -1470 4855 -1440
rect 4825 -1540 4855 -1510
rect 4825 -1610 4855 -1580
rect 4825 -1675 4855 -1645
rect 4825 -1735 4855 -1705
rect 4825 -1800 4855 -1770
rect 4825 -1870 4855 -1840
rect 4825 -1940 4855 -1910
rect 4825 -2010 4855 -1980
rect 4825 -2075 4855 -2045
rect 4825 -2135 4855 -2105
rect 4825 -2200 4855 -2170
rect 4825 -2270 4855 -2240
rect 4825 -2340 4855 -2310
rect 4825 -2410 4855 -2380
rect 4825 -2475 4855 -2445
rect 4825 -2535 4855 -2505
rect 4825 -2600 4855 -2570
rect 4825 -2670 4855 -2640
rect 4825 -2740 4855 -2710
rect 4825 -2810 4855 -2780
rect 4825 -2875 4855 -2845
rect 5175 -1335 5205 -1305
rect 5175 -1400 5205 -1370
rect 5175 -1470 5205 -1440
rect 5175 -1540 5205 -1510
rect 5175 -1610 5205 -1580
rect 5175 -1675 5205 -1645
rect 5175 -1735 5205 -1705
rect 5175 -1800 5205 -1770
rect 5175 -1870 5205 -1840
rect 5175 -1940 5205 -1910
rect 5175 -2010 5205 -1980
rect 5175 -2075 5205 -2045
rect 5175 -2135 5205 -2105
rect 5175 -2200 5205 -2170
rect 5175 -2270 5205 -2240
rect 5175 -2340 5205 -2310
rect 5175 -2410 5205 -2380
rect 5175 -2475 5205 -2445
rect 5175 -2535 5205 -2505
rect 5175 -2600 5205 -2570
rect 5175 -2670 5205 -2640
rect 5175 -2740 5205 -2710
rect 5175 -2810 5205 -2780
rect 5175 -2875 5205 -2845
rect 5525 -1335 5555 -1305
rect 5525 -1400 5555 -1370
rect 5525 -1470 5555 -1440
rect 5525 -1540 5555 -1510
rect 5525 -1610 5555 -1580
rect 5525 -1675 5555 -1645
rect 5525 -1735 5555 -1705
rect 5525 -1800 5555 -1770
rect 5525 -1870 5555 -1840
rect 5525 -1940 5555 -1910
rect 5525 -2010 5555 -1980
rect 5525 -2075 5555 -2045
rect 5525 -2135 5555 -2105
rect 5525 -2200 5555 -2170
rect 5525 -2270 5555 -2240
rect 5525 -2340 5555 -2310
rect 5525 -2410 5555 -2380
rect 5525 -2475 5555 -2445
rect 5525 -2535 5555 -2505
rect 5525 -2600 5555 -2570
rect 5525 -2670 5555 -2640
rect 5525 -2740 5555 -2710
rect 5525 -2810 5555 -2780
rect 5525 -2875 5555 -2845
rect 5875 -1335 5905 -1305
rect 5875 -1400 5905 -1370
rect 5875 -1470 5905 -1440
rect 5875 -1540 5905 -1510
rect 5875 -1610 5905 -1580
rect 5875 -1675 5905 -1645
rect 5875 -1735 5905 -1705
rect 5875 -1800 5905 -1770
rect 5875 -1870 5905 -1840
rect 5875 -1940 5905 -1910
rect 5875 -2010 5905 -1980
rect 5875 -2075 5905 -2045
rect 5875 -2135 5905 -2105
rect 5875 -2200 5905 -2170
rect 5875 -2270 5905 -2240
rect 5875 -2340 5905 -2310
rect 5875 -2410 5905 -2380
rect 5875 -2475 5905 -2445
rect 5875 -2535 5905 -2505
rect 5875 -2600 5905 -2570
rect 5875 -2670 5905 -2640
rect 5875 -2740 5905 -2710
rect 5875 -2810 5905 -2780
rect 5875 -2875 5905 -2845
rect 6225 -1335 6255 -1305
rect 6225 -1400 6255 -1370
rect 6225 -1470 6255 -1440
rect 6225 -1540 6255 -1510
rect 6225 -1610 6255 -1580
rect 6225 -1675 6255 -1645
rect 6225 -1735 6255 -1705
rect 6225 -1800 6255 -1770
rect 6225 -1870 6255 -1840
rect 6225 -1940 6255 -1910
rect 6225 -2010 6255 -1980
rect 6225 -2075 6255 -2045
rect 6225 -2135 6255 -2105
rect 6225 -2200 6255 -2170
rect 6225 -2270 6255 -2240
rect 6225 -2340 6255 -2310
rect 6225 -2410 6255 -2380
rect 6225 -2475 6255 -2445
rect 6225 -2535 6255 -2505
rect 6225 -2600 6255 -2570
rect 6225 -2670 6255 -2640
rect 6225 -2740 6255 -2710
rect 6225 -2810 6255 -2780
rect 6225 -2875 6255 -2845
rect 6575 -1335 6605 -1305
rect 6575 -1400 6605 -1370
rect 6575 -1470 6605 -1440
rect 6575 -1540 6605 -1510
rect 6575 -1610 6605 -1580
rect 6575 -1675 6605 -1645
rect 6575 -1735 6605 -1705
rect 6575 -1800 6605 -1770
rect 6575 -1870 6605 -1840
rect 6575 -1940 6605 -1910
rect 6575 -2010 6605 -1980
rect 6575 -2075 6605 -2045
rect 6575 -2135 6605 -2105
rect 6575 -2200 6605 -2170
rect 6575 -2270 6605 -2240
rect 6575 -2340 6605 -2310
rect 6575 -2410 6605 -2380
rect 6575 -2475 6605 -2445
rect 6575 -2535 6605 -2505
rect 6575 -2600 6605 -2570
rect 6575 -2670 6605 -2640
rect 6575 -2740 6605 -2710
rect 6575 -2810 6605 -2780
rect 6575 -2875 6605 -2845
rect 6925 -1335 6955 -1305
rect 6925 -1400 6955 -1370
rect 6925 -1470 6955 -1440
rect 6925 -1540 6955 -1510
rect 6925 -1610 6955 -1580
rect 6925 -1675 6955 -1645
rect 6925 -1735 6955 -1705
rect 6925 -1800 6955 -1770
rect 6925 -1870 6955 -1840
rect 6925 -1940 6955 -1910
rect 6925 -2010 6955 -1980
rect 6925 -2075 6955 -2045
rect 6925 -2135 6955 -2105
rect 6925 -2200 6955 -2170
rect 6925 -2270 6955 -2240
rect 6925 -2340 6955 -2310
rect 6925 -2410 6955 -2380
rect 6925 -2475 6955 -2445
rect 6925 -2535 6955 -2505
rect 6925 -2600 6955 -2570
rect 6925 -2670 6955 -2640
rect 6925 -2740 6955 -2710
rect 6925 -2810 6955 -2780
rect 6925 -2875 6955 -2845
rect 7275 -1335 7305 -1305
rect 7275 -1400 7305 -1370
rect 7275 -1470 7305 -1440
rect 7275 -1540 7305 -1510
rect 7275 -1610 7305 -1580
rect 7275 -1675 7305 -1645
rect 7275 -1735 7305 -1705
rect 7275 -1800 7305 -1770
rect 7275 -1870 7305 -1840
rect 7275 -1940 7305 -1910
rect 7275 -2010 7305 -1980
rect 7275 -2075 7305 -2045
rect 7275 -2135 7305 -2105
rect 7275 -2200 7305 -2170
rect 7275 -2270 7305 -2240
rect 7275 -2340 7305 -2310
rect 7275 -2410 7305 -2380
rect 7275 -2475 7305 -2445
rect 7275 -2535 7305 -2505
rect 7275 -2600 7305 -2570
rect 7275 -2670 7305 -2640
rect 7275 -2740 7305 -2710
rect 7275 -2810 7305 -2780
rect 7275 -2875 7305 -2845
rect 7625 -1335 7655 -1305
rect 7625 -1400 7655 -1370
rect 7625 -1470 7655 -1440
rect 7625 -1540 7655 -1510
rect 7625 -1610 7655 -1580
rect 7625 -1675 7655 -1645
rect 7625 -1735 7655 -1705
rect 7625 -1800 7655 -1770
rect 7625 -1870 7655 -1840
rect 7625 -1940 7655 -1910
rect 7625 -2010 7655 -1980
rect 7625 -2075 7655 -2045
rect 7625 -2135 7655 -2105
rect 7625 -2200 7655 -2170
rect 7625 -2270 7655 -2240
rect 7625 -2340 7655 -2310
rect 7625 -2410 7655 -2380
rect 7625 -2475 7655 -2445
rect 7625 -2535 7655 -2505
rect 7625 -2600 7655 -2570
rect 7625 -2670 7655 -2640
rect 7625 -2740 7655 -2710
rect 7625 -2810 7655 -2780
rect 7625 -2875 7655 -2845
rect 7975 -1335 8005 -1305
rect 7975 -1400 8005 -1370
rect 7975 -1470 8005 -1440
rect 7975 -1540 8005 -1510
rect 7975 -1610 8005 -1580
rect 7975 -1675 8005 -1645
rect 7975 -1735 8005 -1705
rect 7975 -1800 8005 -1770
rect 7975 -1870 8005 -1840
rect 7975 -1940 8005 -1910
rect 7975 -2010 8005 -1980
rect 7975 -2075 8005 -2045
rect 7975 -2135 8005 -2105
rect 7975 -2200 8005 -2170
rect 7975 -2270 8005 -2240
rect 7975 -2340 8005 -2310
rect 7975 -2410 8005 -2380
rect 7975 -2475 8005 -2445
rect 7975 -2535 8005 -2505
rect 7975 -2600 8005 -2570
rect 7975 -2670 8005 -2640
rect 7975 -2740 8005 -2710
rect 7975 -2810 8005 -2780
rect 7975 -2875 8005 -2845
rect 8325 -1335 8355 -1305
rect 8325 -1400 8355 -1370
rect 8325 -1470 8355 -1440
rect 8325 -1540 8355 -1510
rect 8325 -1610 8355 -1580
rect 8325 -1675 8355 -1645
rect 8325 -1735 8355 -1705
rect 8325 -1800 8355 -1770
rect 8325 -1870 8355 -1840
rect 8325 -1940 8355 -1910
rect 8325 -2010 8355 -1980
rect 8325 -2075 8355 -2045
rect 8325 -2135 8355 -2105
rect 8325 -2200 8355 -2170
rect 8325 -2270 8355 -2240
rect 8325 -2340 8355 -2310
rect 8325 -2410 8355 -2380
rect 8325 -2475 8355 -2445
rect 8325 -2535 8355 -2505
rect 8325 -2600 8355 -2570
rect 8325 -2670 8355 -2640
rect 8325 -2740 8355 -2710
rect 8325 -2810 8355 -2780
rect 8325 -2875 8355 -2845
rect 8675 -1335 8705 -1305
rect 8675 -1400 8705 -1370
rect 8675 -1470 8705 -1440
rect 8675 -1540 8705 -1510
rect 8675 -1610 8705 -1580
rect 8675 -1675 8705 -1645
rect 8675 -1735 8705 -1705
rect 8675 -1800 8705 -1770
rect 8675 -1870 8705 -1840
rect 8675 -1940 8705 -1910
rect 8675 -2010 8705 -1980
rect 8675 -2075 8705 -2045
rect 8675 -2135 8705 -2105
rect 8675 -2200 8705 -2170
rect 8675 -2270 8705 -2240
rect 8675 -2340 8705 -2310
rect 8675 -2410 8705 -2380
rect 8675 -2475 8705 -2445
rect 8675 -2535 8705 -2505
rect 8675 -2600 8705 -2570
rect 8675 -2670 8705 -2640
rect 8675 -2740 8705 -2710
rect 8675 -2810 8705 -2780
rect 8675 -2875 8705 -2845
rect 9025 -1335 9055 -1305
rect 9025 -1400 9055 -1370
rect 9025 -1470 9055 -1440
rect 9025 -1540 9055 -1510
rect 9025 -1610 9055 -1580
rect 9025 -1675 9055 -1645
rect 9025 -1735 9055 -1705
rect 9025 -1800 9055 -1770
rect 9025 -1870 9055 -1840
rect 9025 -1940 9055 -1910
rect 9025 -2010 9055 -1980
rect 9025 -2075 9055 -2045
rect 9025 -2135 9055 -2105
rect 9025 -2200 9055 -2170
rect 9025 -2270 9055 -2240
rect 9025 -2340 9055 -2310
rect 9025 -2410 9055 -2380
rect 9025 -2475 9055 -2445
rect 9025 -2535 9055 -2505
rect 9025 -2600 9055 -2570
rect 9025 -2670 9055 -2640
rect 9025 -2740 9055 -2710
rect 9025 -2810 9055 -2780
rect 9025 -2875 9055 -2845
<< metal3 >>
rect 2100 19315 2160 19325
rect 2100 19275 2110 19315
rect 2150 19275 2160 19315
rect 2100 19250 2160 19275
rect 2100 19210 2110 19250
rect 2150 19210 2160 19250
rect 2100 19180 2160 19210
rect 2100 19140 2110 19180
rect 2150 19140 2160 19180
rect 2100 19110 2160 19140
rect 2100 19070 2110 19110
rect 2150 19070 2160 19110
rect 2100 19040 2160 19070
rect 2100 19000 2110 19040
rect 2150 19000 2160 19040
rect 2100 18975 2160 19000
rect 2100 18935 2110 18975
rect 2150 18935 2160 18975
rect 2100 18915 2160 18935
rect 2100 18875 2110 18915
rect 2150 18875 2160 18915
rect 2100 18850 2160 18875
rect 2100 18810 2110 18850
rect 2150 18810 2160 18850
rect 2100 18780 2160 18810
rect 2100 18740 2110 18780
rect 2150 18740 2160 18780
rect 2100 18710 2160 18740
rect 2100 18670 2110 18710
rect 2150 18670 2160 18710
rect 2100 18640 2160 18670
rect 2100 18600 2110 18640
rect 2150 18600 2160 18640
rect 2100 18575 2160 18600
rect 2100 18535 2110 18575
rect 2150 18535 2160 18575
rect 2100 18515 2160 18535
rect 2100 18475 2110 18515
rect 2150 18475 2160 18515
rect 2100 18450 2160 18475
rect 2100 18410 2110 18450
rect 2150 18410 2160 18450
rect 2100 18380 2160 18410
rect 2100 18340 2110 18380
rect 2150 18340 2160 18380
rect 2100 18310 2160 18340
rect 2100 18270 2110 18310
rect 2150 18270 2160 18310
rect 2100 18240 2160 18270
rect 2100 18200 2110 18240
rect 2150 18200 2160 18240
rect 2100 18175 2160 18200
rect 2100 18135 2110 18175
rect 2150 18135 2160 18175
rect 2100 18115 2160 18135
rect 2100 18075 2110 18115
rect 2150 18075 2160 18115
rect 2100 18050 2160 18075
rect 2100 18010 2110 18050
rect 2150 18010 2160 18050
rect 2100 17980 2160 18010
rect 2100 17940 2110 17980
rect 2150 17940 2160 17980
rect 2100 17910 2160 17940
rect 2100 17870 2110 17910
rect 2150 17870 2160 17910
rect 2100 17840 2160 17870
rect 2100 17800 2110 17840
rect 2150 17800 2160 17840
rect 2100 17775 2160 17800
rect 2100 17735 2110 17775
rect 2150 17735 2160 17775
rect 2100 17725 2160 17735
rect 6690 19315 6750 19325
rect 6690 19275 6700 19315
rect 6740 19275 6750 19315
rect 6690 19250 6750 19275
rect 6690 19210 6700 19250
rect 6740 19210 6750 19250
rect 6690 19180 6750 19210
rect 6690 19140 6700 19180
rect 6740 19140 6750 19180
rect 6690 19110 6750 19140
rect 6690 19070 6700 19110
rect 6740 19070 6750 19110
rect 6690 19040 6750 19070
rect 6690 19000 6700 19040
rect 6740 19000 6750 19040
rect 6690 18975 6750 19000
rect 6690 18935 6700 18975
rect 6740 18935 6750 18975
rect 6690 18915 6750 18935
rect 6690 18875 6700 18915
rect 6740 18875 6750 18915
rect 6690 18850 6750 18875
rect 6690 18810 6700 18850
rect 6740 18810 6750 18850
rect 6690 18780 6750 18810
rect 6690 18740 6700 18780
rect 6740 18740 6750 18780
rect 6690 18710 6750 18740
rect 6690 18670 6700 18710
rect 6740 18670 6750 18710
rect 6690 18640 6750 18670
rect 6690 18600 6700 18640
rect 6740 18600 6750 18640
rect 6690 18575 6750 18600
rect 6690 18535 6700 18575
rect 6740 18535 6750 18575
rect 6690 18515 6750 18535
rect 6690 18475 6700 18515
rect 6740 18475 6750 18515
rect 6690 18450 6750 18475
rect 6690 18410 6700 18450
rect 6740 18410 6750 18450
rect 6690 18380 6750 18410
rect 6690 18340 6700 18380
rect 6740 18340 6750 18380
rect 6690 18310 6750 18340
rect 6690 18270 6700 18310
rect 6740 18270 6750 18310
rect 6690 18240 6750 18270
rect 6690 18200 6700 18240
rect 6740 18200 6750 18240
rect 6690 18175 6750 18200
rect 6690 18135 6700 18175
rect 6740 18135 6750 18175
rect 6690 18115 6750 18135
rect 6690 18075 6700 18115
rect 6740 18075 6750 18115
rect 6690 18050 6750 18075
rect 6690 18010 6700 18050
rect 6740 18010 6750 18050
rect 6690 17980 6750 18010
rect 6690 17940 6700 17980
rect 6740 17940 6750 17980
rect 6690 17910 6750 17940
rect 6690 17870 6700 17910
rect 6740 17870 6750 17910
rect 6690 17840 6750 17870
rect 6690 17800 6700 17840
rect 6740 17800 6750 17840
rect 6690 17775 6750 17800
rect 6690 17735 6700 17775
rect 6740 17735 6750 17775
rect 6690 17725 6750 17735
rect 31290 19305 32890 19325
rect 31290 19270 31305 19305
rect 31340 19270 31350 19305
rect 31385 19270 31395 19305
rect 31430 19270 31440 19305
rect 31475 19270 31485 19305
rect 31520 19270 31530 19305
rect 31565 19270 31575 19305
rect 31610 19270 31620 19305
rect 31655 19270 31665 19305
rect 31700 19270 31710 19305
rect 31745 19270 31755 19305
rect 31790 19270 31800 19305
rect 31835 19270 31845 19305
rect 31880 19270 31890 19305
rect 31925 19270 31935 19305
rect 31970 19270 31980 19305
rect 32015 19270 32025 19305
rect 32060 19270 32070 19305
rect 32105 19270 32115 19305
rect 32150 19270 32160 19305
rect 32195 19270 32205 19305
rect 32240 19270 32250 19305
rect 32285 19270 32295 19305
rect 32330 19270 32340 19305
rect 32375 19270 32385 19305
rect 32420 19270 32430 19305
rect 32465 19270 32475 19305
rect 32510 19270 32520 19305
rect 32555 19270 32565 19305
rect 32600 19270 32610 19305
rect 32645 19270 32655 19305
rect 32690 19270 32700 19305
rect 32735 19270 32745 19305
rect 32780 19270 32790 19305
rect 32825 19270 32835 19305
rect 32870 19270 32890 19305
rect 31290 19260 32890 19270
rect 31290 19225 31305 19260
rect 31340 19225 31350 19260
rect 31385 19225 31395 19260
rect 31430 19225 31440 19260
rect 31475 19225 31485 19260
rect 31520 19225 31530 19260
rect 31565 19225 31575 19260
rect 31610 19225 31620 19260
rect 31655 19225 31665 19260
rect 31700 19225 31710 19260
rect 31745 19225 31755 19260
rect 31790 19225 31800 19260
rect 31835 19225 31845 19260
rect 31880 19225 31890 19260
rect 31925 19225 31935 19260
rect 31970 19225 31980 19260
rect 32015 19225 32025 19260
rect 32060 19225 32070 19260
rect 32105 19225 32115 19260
rect 32150 19225 32160 19260
rect 32195 19225 32205 19260
rect 32240 19225 32250 19260
rect 32285 19225 32295 19260
rect 32330 19225 32340 19260
rect 32375 19225 32385 19260
rect 32420 19225 32430 19260
rect 32465 19225 32475 19260
rect 32510 19225 32520 19260
rect 32555 19225 32565 19260
rect 32600 19225 32610 19260
rect 32645 19225 32655 19260
rect 32690 19225 32700 19260
rect 32735 19225 32745 19260
rect 32780 19225 32790 19260
rect 32825 19225 32835 19260
rect 32870 19225 32890 19260
rect 31290 19215 32890 19225
rect 31290 19180 31305 19215
rect 31340 19180 31350 19215
rect 31385 19180 31395 19215
rect 31430 19180 31440 19215
rect 31475 19180 31485 19215
rect 31520 19180 31530 19215
rect 31565 19180 31575 19215
rect 31610 19180 31620 19215
rect 31655 19180 31665 19215
rect 31700 19180 31710 19215
rect 31745 19180 31755 19215
rect 31790 19180 31800 19215
rect 31835 19180 31845 19215
rect 31880 19180 31890 19215
rect 31925 19180 31935 19215
rect 31970 19180 31980 19215
rect 32015 19180 32025 19215
rect 32060 19180 32070 19215
rect 32105 19180 32115 19215
rect 32150 19180 32160 19215
rect 32195 19180 32205 19215
rect 32240 19180 32250 19215
rect 32285 19180 32295 19215
rect 32330 19180 32340 19215
rect 32375 19180 32385 19215
rect 32420 19180 32430 19215
rect 32465 19180 32475 19215
rect 32510 19180 32520 19215
rect 32555 19180 32565 19215
rect 32600 19180 32610 19215
rect 32645 19180 32655 19215
rect 32690 19180 32700 19215
rect 32735 19180 32745 19215
rect 32780 19180 32790 19215
rect 32825 19180 32835 19215
rect 32870 19180 32890 19215
rect 31290 19170 32890 19180
rect 31290 19135 31305 19170
rect 31340 19135 31350 19170
rect 31385 19135 31395 19170
rect 31430 19135 31440 19170
rect 31475 19135 31485 19170
rect 31520 19135 31530 19170
rect 31565 19135 31575 19170
rect 31610 19135 31620 19170
rect 31655 19135 31665 19170
rect 31700 19135 31710 19170
rect 31745 19135 31755 19170
rect 31790 19135 31800 19170
rect 31835 19135 31845 19170
rect 31880 19135 31890 19170
rect 31925 19135 31935 19170
rect 31970 19135 31980 19170
rect 32015 19135 32025 19170
rect 32060 19135 32070 19170
rect 32105 19135 32115 19170
rect 32150 19135 32160 19170
rect 32195 19135 32205 19170
rect 32240 19135 32250 19170
rect 32285 19135 32295 19170
rect 32330 19135 32340 19170
rect 32375 19135 32385 19170
rect 32420 19135 32430 19170
rect 32465 19135 32475 19170
rect 32510 19135 32520 19170
rect 32555 19135 32565 19170
rect 32600 19135 32610 19170
rect 32645 19135 32655 19170
rect 32690 19135 32700 19170
rect 32735 19135 32745 19170
rect 32780 19135 32790 19170
rect 32825 19135 32835 19170
rect 32870 19135 32890 19170
rect 31290 19125 32890 19135
rect 31290 19090 31305 19125
rect 31340 19090 31350 19125
rect 31385 19090 31395 19125
rect 31430 19090 31440 19125
rect 31475 19090 31485 19125
rect 31520 19090 31530 19125
rect 31565 19090 31575 19125
rect 31610 19090 31620 19125
rect 31655 19090 31665 19125
rect 31700 19090 31710 19125
rect 31745 19090 31755 19125
rect 31790 19090 31800 19125
rect 31835 19090 31845 19125
rect 31880 19090 31890 19125
rect 31925 19090 31935 19125
rect 31970 19090 31980 19125
rect 32015 19090 32025 19125
rect 32060 19090 32070 19125
rect 32105 19090 32115 19125
rect 32150 19090 32160 19125
rect 32195 19090 32205 19125
rect 32240 19090 32250 19125
rect 32285 19090 32295 19125
rect 32330 19090 32340 19125
rect 32375 19090 32385 19125
rect 32420 19090 32430 19125
rect 32465 19090 32475 19125
rect 32510 19090 32520 19125
rect 32555 19090 32565 19125
rect 32600 19090 32610 19125
rect 32645 19090 32655 19125
rect 32690 19090 32700 19125
rect 32735 19090 32745 19125
rect 32780 19090 32790 19125
rect 32825 19090 32835 19125
rect 32870 19090 32890 19125
rect 31290 19080 32890 19090
rect 31290 19045 31305 19080
rect 31340 19045 31350 19080
rect 31385 19045 31395 19080
rect 31430 19045 31440 19080
rect 31475 19045 31485 19080
rect 31520 19045 31530 19080
rect 31565 19045 31575 19080
rect 31610 19045 31620 19080
rect 31655 19045 31665 19080
rect 31700 19045 31710 19080
rect 31745 19045 31755 19080
rect 31790 19045 31800 19080
rect 31835 19045 31845 19080
rect 31880 19045 31890 19080
rect 31925 19045 31935 19080
rect 31970 19045 31980 19080
rect 32015 19045 32025 19080
rect 32060 19045 32070 19080
rect 32105 19045 32115 19080
rect 32150 19045 32160 19080
rect 32195 19045 32205 19080
rect 32240 19045 32250 19080
rect 32285 19045 32295 19080
rect 32330 19045 32340 19080
rect 32375 19045 32385 19080
rect 32420 19045 32430 19080
rect 32465 19045 32475 19080
rect 32510 19045 32520 19080
rect 32555 19045 32565 19080
rect 32600 19045 32610 19080
rect 32645 19045 32655 19080
rect 32690 19045 32700 19080
rect 32735 19045 32745 19080
rect 32780 19045 32790 19080
rect 32825 19045 32835 19080
rect 32870 19045 32890 19080
rect 31290 19035 32890 19045
rect 31290 19000 31305 19035
rect 31340 19000 31350 19035
rect 31385 19000 31395 19035
rect 31430 19000 31440 19035
rect 31475 19000 31485 19035
rect 31520 19000 31530 19035
rect 31565 19000 31575 19035
rect 31610 19000 31620 19035
rect 31655 19000 31665 19035
rect 31700 19000 31710 19035
rect 31745 19000 31755 19035
rect 31790 19000 31800 19035
rect 31835 19000 31845 19035
rect 31880 19000 31890 19035
rect 31925 19000 31935 19035
rect 31970 19000 31980 19035
rect 32015 19000 32025 19035
rect 32060 19000 32070 19035
rect 32105 19000 32115 19035
rect 32150 19000 32160 19035
rect 32195 19000 32205 19035
rect 32240 19000 32250 19035
rect 32285 19000 32295 19035
rect 32330 19000 32340 19035
rect 32375 19000 32385 19035
rect 32420 19000 32430 19035
rect 32465 19000 32475 19035
rect 32510 19000 32520 19035
rect 32555 19000 32565 19035
rect 32600 19000 32610 19035
rect 32645 19000 32655 19035
rect 32690 19000 32700 19035
rect 32735 19000 32745 19035
rect 32780 19000 32790 19035
rect 32825 19000 32835 19035
rect 32870 19000 32890 19035
rect 31290 18990 32890 19000
rect 31290 18955 31305 18990
rect 31340 18955 31350 18990
rect 31385 18955 31395 18990
rect 31430 18955 31440 18990
rect 31475 18955 31485 18990
rect 31520 18955 31530 18990
rect 31565 18955 31575 18990
rect 31610 18955 31620 18990
rect 31655 18955 31665 18990
rect 31700 18955 31710 18990
rect 31745 18955 31755 18990
rect 31790 18955 31800 18990
rect 31835 18955 31845 18990
rect 31880 18955 31890 18990
rect 31925 18955 31935 18990
rect 31970 18955 31980 18990
rect 32015 18955 32025 18990
rect 32060 18955 32070 18990
rect 32105 18955 32115 18990
rect 32150 18955 32160 18990
rect 32195 18955 32205 18990
rect 32240 18955 32250 18990
rect 32285 18955 32295 18990
rect 32330 18955 32340 18990
rect 32375 18955 32385 18990
rect 32420 18955 32430 18990
rect 32465 18955 32475 18990
rect 32510 18955 32520 18990
rect 32555 18955 32565 18990
rect 32600 18955 32610 18990
rect 32645 18955 32655 18990
rect 32690 18955 32700 18990
rect 32735 18955 32745 18990
rect 32780 18955 32790 18990
rect 32825 18955 32835 18990
rect 32870 18955 32890 18990
rect 31290 18945 32890 18955
rect 31290 18910 31305 18945
rect 31340 18910 31350 18945
rect 31385 18910 31395 18945
rect 31430 18910 31440 18945
rect 31475 18910 31485 18945
rect 31520 18910 31530 18945
rect 31565 18910 31575 18945
rect 31610 18910 31620 18945
rect 31655 18910 31665 18945
rect 31700 18910 31710 18945
rect 31745 18910 31755 18945
rect 31790 18910 31800 18945
rect 31835 18910 31845 18945
rect 31880 18910 31890 18945
rect 31925 18910 31935 18945
rect 31970 18910 31980 18945
rect 32015 18910 32025 18945
rect 32060 18910 32070 18945
rect 32105 18910 32115 18945
rect 32150 18910 32160 18945
rect 32195 18910 32205 18945
rect 32240 18910 32250 18945
rect 32285 18910 32295 18945
rect 32330 18910 32340 18945
rect 32375 18910 32385 18945
rect 32420 18910 32430 18945
rect 32465 18910 32475 18945
rect 32510 18910 32520 18945
rect 32555 18910 32565 18945
rect 32600 18910 32610 18945
rect 32645 18910 32655 18945
rect 32690 18910 32700 18945
rect 32735 18910 32745 18945
rect 32780 18910 32790 18945
rect 32825 18910 32835 18945
rect 32870 18910 32890 18945
rect 31290 18900 32890 18910
rect 31290 18865 31305 18900
rect 31340 18865 31350 18900
rect 31385 18865 31395 18900
rect 31430 18865 31440 18900
rect 31475 18865 31485 18900
rect 31520 18865 31530 18900
rect 31565 18865 31575 18900
rect 31610 18865 31620 18900
rect 31655 18865 31665 18900
rect 31700 18865 31710 18900
rect 31745 18865 31755 18900
rect 31790 18865 31800 18900
rect 31835 18865 31845 18900
rect 31880 18865 31890 18900
rect 31925 18865 31935 18900
rect 31970 18865 31980 18900
rect 32015 18865 32025 18900
rect 32060 18865 32070 18900
rect 32105 18865 32115 18900
rect 32150 18865 32160 18900
rect 32195 18865 32205 18900
rect 32240 18865 32250 18900
rect 32285 18865 32295 18900
rect 32330 18865 32340 18900
rect 32375 18865 32385 18900
rect 32420 18865 32430 18900
rect 32465 18865 32475 18900
rect 32510 18865 32520 18900
rect 32555 18865 32565 18900
rect 32600 18865 32610 18900
rect 32645 18865 32655 18900
rect 32690 18865 32700 18900
rect 32735 18865 32745 18900
rect 32780 18865 32790 18900
rect 32825 18865 32835 18900
rect 32870 18865 32890 18900
rect 31290 18855 32890 18865
rect 31290 18820 31305 18855
rect 31340 18820 31350 18855
rect 31385 18820 31395 18855
rect 31430 18820 31440 18855
rect 31475 18820 31485 18855
rect 31520 18820 31530 18855
rect 31565 18820 31575 18855
rect 31610 18820 31620 18855
rect 31655 18820 31665 18855
rect 31700 18820 31710 18855
rect 31745 18820 31755 18855
rect 31790 18820 31800 18855
rect 31835 18820 31845 18855
rect 31880 18820 31890 18855
rect 31925 18820 31935 18855
rect 31970 18820 31980 18855
rect 32015 18820 32025 18855
rect 32060 18820 32070 18855
rect 32105 18820 32115 18855
rect 32150 18820 32160 18855
rect 32195 18820 32205 18855
rect 32240 18820 32250 18855
rect 32285 18820 32295 18855
rect 32330 18820 32340 18855
rect 32375 18820 32385 18855
rect 32420 18820 32430 18855
rect 32465 18820 32475 18855
rect 32510 18820 32520 18855
rect 32555 18820 32565 18855
rect 32600 18820 32610 18855
rect 32645 18820 32655 18855
rect 32690 18820 32700 18855
rect 32735 18820 32745 18855
rect 32780 18820 32790 18855
rect 32825 18820 32835 18855
rect 32870 18820 32890 18855
rect 31290 18810 32890 18820
rect 31290 18775 31305 18810
rect 31340 18775 31350 18810
rect 31385 18775 31395 18810
rect 31430 18775 31440 18810
rect 31475 18775 31485 18810
rect 31520 18775 31530 18810
rect 31565 18775 31575 18810
rect 31610 18775 31620 18810
rect 31655 18775 31665 18810
rect 31700 18775 31710 18810
rect 31745 18775 31755 18810
rect 31790 18775 31800 18810
rect 31835 18775 31845 18810
rect 31880 18775 31890 18810
rect 31925 18775 31935 18810
rect 31970 18775 31980 18810
rect 32015 18775 32025 18810
rect 32060 18775 32070 18810
rect 32105 18775 32115 18810
rect 32150 18775 32160 18810
rect 32195 18775 32205 18810
rect 32240 18775 32250 18810
rect 32285 18775 32295 18810
rect 32330 18775 32340 18810
rect 32375 18775 32385 18810
rect 32420 18775 32430 18810
rect 32465 18775 32475 18810
rect 32510 18775 32520 18810
rect 32555 18775 32565 18810
rect 32600 18775 32610 18810
rect 32645 18775 32655 18810
rect 32690 18775 32700 18810
rect 32735 18775 32745 18810
rect 32780 18775 32790 18810
rect 32825 18775 32835 18810
rect 32870 18775 32890 18810
rect 31290 18765 32890 18775
rect 31290 18730 31305 18765
rect 31340 18730 31350 18765
rect 31385 18730 31395 18765
rect 31430 18730 31440 18765
rect 31475 18730 31485 18765
rect 31520 18730 31530 18765
rect 31565 18730 31575 18765
rect 31610 18730 31620 18765
rect 31655 18730 31665 18765
rect 31700 18730 31710 18765
rect 31745 18730 31755 18765
rect 31790 18730 31800 18765
rect 31835 18730 31845 18765
rect 31880 18730 31890 18765
rect 31925 18730 31935 18765
rect 31970 18730 31980 18765
rect 32015 18730 32025 18765
rect 32060 18730 32070 18765
rect 32105 18730 32115 18765
rect 32150 18730 32160 18765
rect 32195 18730 32205 18765
rect 32240 18730 32250 18765
rect 32285 18730 32295 18765
rect 32330 18730 32340 18765
rect 32375 18730 32385 18765
rect 32420 18730 32430 18765
rect 32465 18730 32475 18765
rect 32510 18730 32520 18765
rect 32555 18730 32565 18765
rect 32600 18730 32610 18765
rect 32645 18730 32655 18765
rect 32690 18730 32700 18765
rect 32735 18730 32745 18765
rect 32780 18730 32790 18765
rect 32825 18730 32835 18765
rect 32870 18730 32890 18765
rect 31290 18720 32890 18730
rect 31290 18685 31305 18720
rect 31340 18685 31350 18720
rect 31385 18685 31395 18720
rect 31430 18685 31440 18720
rect 31475 18685 31485 18720
rect 31520 18685 31530 18720
rect 31565 18685 31575 18720
rect 31610 18685 31620 18720
rect 31655 18685 31665 18720
rect 31700 18685 31710 18720
rect 31745 18685 31755 18720
rect 31790 18685 31800 18720
rect 31835 18685 31845 18720
rect 31880 18685 31890 18720
rect 31925 18685 31935 18720
rect 31970 18685 31980 18720
rect 32015 18685 32025 18720
rect 32060 18685 32070 18720
rect 32105 18685 32115 18720
rect 32150 18685 32160 18720
rect 32195 18685 32205 18720
rect 32240 18685 32250 18720
rect 32285 18685 32295 18720
rect 32330 18685 32340 18720
rect 32375 18685 32385 18720
rect 32420 18685 32430 18720
rect 32465 18685 32475 18720
rect 32510 18685 32520 18720
rect 32555 18685 32565 18720
rect 32600 18685 32610 18720
rect 32645 18685 32655 18720
rect 32690 18685 32700 18720
rect 32735 18685 32745 18720
rect 32780 18685 32790 18720
rect 32825 18685 32835 18720
rect 32870 18685 32890 18720
rect 31290 18675 32890 18685
rect 31290 18640 31305 18675
rect 31340 18640 31350 18675
rect 31385 18640 31395 18675
rect 31430 18640 31440 18675
rect 31475 18640 31485 18675
rect 31520 18640 31530 18675
rect 31565 18640 31575 18675
rect 31610 18640 31620 18675
rect 31655 18640 31665 18675
rect 31700 18640 31710 18675
rect 31745 18640 31755 18675
rect 31790 18640 31800 18675
rect 31835 18640 31845 18675
rect 31880 18640 31890 18675
rect 31925 18640 31935 18675
rect 31970 18640 31980 18675
rect 32015 18640 32025 18675
rect 32060 18640 32070 18675
rect 32105 18640 32115 18675
rect 32150 18640 32160 18675
rect 32195 18640 32205 18675
rect 32240 18640 32250 18675
rect 32285 18640 32295 18675
rect 32330 18640 32340 18675
rect 32375 18640 32385 18675
rect 32420 18640 32430 18675
rect 32465 18640 32475 18675
rect 32510 18640 32520 18675
rect 32555 18640 32565 18675
rect 32600 18640 32610 18675
rect 32645 18640 32655 18675
rect 32690 18640 32700 18675
rect 32735 18640 32745 18675
rect 32780 18640 32790 18675
rect 32825 18640 32835 18675
rect 32870 18640 32890 18675
rect 31290 18630 32890 18640
rect 31290 18595 31305 18630
rect 31340 18595 31350 18630
rect 31385 18595 31395 18630
rect 31430 18595 31440 18630
rect 31475 18595 31485 18630
rect 31520 18595 31530 18630
rect 31565 18595 31575 18630
rect 31610 18595 31620 18630
rect 31655 18595 31665 18630
rect 31700 18595 31710 18630
rect 31745 18595 31755 18630
rect 31790 18595 31800 18630
rect 31835 18595 31845 18630
rect 31880 18595 31890 18630
rect 31925 18595 31935 18630
rect 31970 18595 31980 18630
rect 32015 18595 32025 18630
rect 32060 18595 32070 18630
rect 32105 18595 32115 18630
rect 32150 18595 32160 18630
rect 32195 18595 32205 18630
rect 32240 18595 32250 18630
rect 32285 18595 32295 18630
rect 32330 18595 32340 18630
rect 32375 18595 32385 18630
rect 32420 18595 32430 18630
rect 32465 18595 32475 18630
rect 32510 18595 32520 18630
rect 32555 18595 32565 18630
rect 32600 18595 32610 18630
rect 32645 18595 32655 18630
rect 32690 18595 32700 18630
rect 32735 18595 32745 18630
rect 32780 18595 32790 18630
rect 32825 18595 32835 18630
rect 32870 18595 32890 18630
rect 31290 18585 32890 18595
rect 31290 18550 31305 18585
rect 31340 18550 31350 18585
rect 31385 18550 31395 18585
rect 31430 18550 31440 18585
rect 31475 18550 31485 18585
rect 31520 18550 31530 18585
rect 31565 18550 31575 18585
rect 31610 18550 31620 18585
rect 31655 18550 31665 18585
rect 31700 18550 31710 18585
rect 31745 18550 31755 18585
rect 31790 18550 31800 18585
rect 31835 18550 31845 18585
rect 31880 18550 31890 18585
rect 31925 18550 31935 18585
rect 31970 18550 31980 18585
rect 32015 18550 32025 18585
rect 32060 18550 32070 18585
rect 32105 18550 32115 18585
rect 32150 18550 32160 18585
rect 32195 18550 32205 18585
rect 32240 18550 32250 18585
rect 32285 18550 32295 18585
rect 32330 18550 32340 18585
rect 32375 18550 32385 18585
rect 32420 18550 32430 18585
rect 32465 18550 32475 18585
rect 32510 18550 32520 18585
rect 32555 18550 32565 18585
rect 32600 18550 32610 18585
rect 32645 18550 32655 18585
rect 32690 18550 32700 18585
rect 32735 18550 32745 18585
rect 32780 18550 32790 18585
rect 32825 18550 32835 18585
rect 32870 18550 32890 18585
rect 31290 18540 32890 18550
rect 31290 18505 31305 18540
rect 31340 18505 31350 18540
rect 31385 18505 31395 18540
rect 31430 18505 31440 18540
rect 31475 18505 31485 18540
rect 31520 18505 31530 18540
rect 31565 18505 31575 18540
rect 31610 18505 31620 18540
rect 31655 18505 31665 18540
rect 31700 18505 31710 18540
rect 31745 18505 31755 18540
rect 31790 18505 31800 18540
rect 31835 18505 31845 18540
rect 31880 18505 31890 18540
rect 31925 18505 31935 18540
rect 31970 18505 31980 18540
rect 32015 18505 32025 18540
rect 32060 18505 32070 18540
rect 32105 18505 32115 18540
rect 32150 18505 32160 18540
rect 32195 18505 32205 18540
rect 32240 18505 32250 18540
rect 32285 18505 32295 18540
rect 32330 18505 32340 18540
rect 32375 18505 32385 18540
rect 32420 18505 32430 18540
rect 32465 18505 32475 18540
rect 32510 18505 32520 18540
rect 32555 18505 32565 18540
rect 32600 18505 32610 18540
rect 32645 18505 32655 18540
rect 32690 18505 32700 18540
rect 32735 18505 32745 18540
rect 32780 18505 32790 18540
rect 32825 18505 32835 18540
rect 32870 18505 32890 18540
rect 31290 18495 32890 18505
rect 31290 18460 31305 18495
rect 31340 18460 31350 18495
rect 31385 18460 31395 18495
rect 31430 18460 31440 18495
rect 31475 18460 31485 18495
rect 31520 18460 31530 18495
rect 31565 18460 31575 18495
rect 31610 18460 31620 18495
rect 31655 18460 31665 18495
rect 31700 18460 31710 18495
rect 31745 18460 31755 18495
rect 31790 18460 31800 18495
rect 31835 18460 31845 18495
rect 31880 18460 31890 18495
rect 31925 18460 31935 18495
rect 31970 18460 31980 18495
rect 32015 18460 32025 18495
rect 32060 18460 32070 18495
rect 32105 18460 32115 18495
rect 32150 18460 32160 18495
rect 32195 18460 32205 18495
rect 32240 18460 32250 18495
rect 32285 18460 32295 18495
rect 32330 18460 32340 18495
rect 32375 18460 32385 18495
rect 32420 18460 32430 18495
rect 32465 18460 32475 18495
rect 32510 18460 32520 18495
rect 32555 18460 32565 18495
rect 32600 18460 32610 18495
rect 32645 18460 32655 18495
rect 32690 18460 32700 18495
rect 32735 18460 32745 18495
rect 32780 18460 32790 18495
rect 32825 18460 32835 18495
rect 32870 18460 32890 18495
rect 31290 18450 32890 18460
rect 31290 18415 31305 18450
rect 31340 18415 31350 18450
rect 31385 18415 31395 18450
rect 31430 18415 31440 18450
rect 31475 18415 31485 18450
rect 31520 18415 31530 18450
rect 31565 18415 31575 18450
rect 31610 18415 31620 18450
rect 31655 18415 31665 18450
rect 31700 18415 31710 18450
rect 31745 18415 31755 18450
rect 31790 18415 31800 18450
rect 31835 18415 31845 18450
rect 31880 18415 31890 18450
rect 31925 18415 31935 18450
rect 31970 18415 31980 18450
rect 32015 18415 32025 18450
rect 32060 18415 32070 18450
rect 32105 18415 32115 18450
rect 32150 18415 32160 18450
rect 32195 18415 32205 18450
rect 32240 18415 32250 18450
rect 32285 18415 32295 18450
rect 32330 18415 32340 18450
rect 32375 18415 32385 18450
rect 32420 18415 32430 18450
rect 32465 18415 32475 18450
rect 32510 18415 32520 18450
rect 32555 18415 32565 18450
rect 32600 18415 32610 18450
rect 32645 18415 32655 18450
rect 32690 18415 32700 18450
rect 32735 18415 32745 18450
rect 32780 18415 32790 18450
rect 32825 18415 32835 18450
rect 32870 18415 32890 18450
rect 31290 18405 32890 18415
rect 31290 18370 31305 18405
rect 31340 18370 31350 18405
rect 31385 18370 31395 18405
rect 31430 18370 31440 18405
rect 31475 18370 31485 18405
rect 31520 18370 31530 18405
rect 31565 18370 31575 18405
rect 31610 18370 31620 18405
rect 31655 18370 31665 18405
rect 31700 18370 31710 18405
rect 31745 18370 31755 18405
rect 31790 18370 31800 18405
rect 31835 18370 31845 18405
rect 31880 18370 31890 18405
rect 31925 18370 31935 18405
rect 31970 18370 31980 18405
rect 32015 18370 32025 18405
rect 32060 18370 32070 18405
rect 32105 18370 32115 18405
rect 32150 18370 32160 18405
rect 32195 18370 32205 18405
rect 32240 18370 32250 18405
rect 32285 18370 32295 18405
rect 32330 18370 32340 18405
rect 32375 18370 32385 18405
rect 32420 18370 32430 18405
rect 32465 18370 32475 18405
rect 32510 18370 32520 18405
rect 32555 18370 32565 18405
rect 32600 18370 32610 18405
rect 32645 18370 32655 18405
rect 32690 18370 32700 18405
rect 32735 18370 32745 18405
rect 32780 18370 32790 18405
rect 32825 18370 32835 18405
rect 32870 18370 32890 18405
rect 31290 18360 32890 18370
rect 31290 18325 31305 18360
rect 31340 18325 31350 18360
rect 31385 18325 31395 18360
rect 31430 18325 31440 18360
rect 31475 18325 31485 18360
rect 31520 18325 31530 18360
rect 31565 18325 31575 18360
rect 31610 18325 31620 18360
rect 31655 18325 31665 18360
rect 31700 18325 31710 18360
rect 31745 18325 31755 18360
rect 31790 18325 31800 18360
rect 31835 18325 31845 18360
rect 31880 18325 31890 18360
rect 31925 18325 31935 18360
rect 31970 18325 31980 18360
rect 32015 18325 32025 18360
rect 32060 18325 32070 18360
rect 32105 18325 32115 18360
rect 32150 18325 32160 18360
rect 32195 18325 32205 18360
rect 32240 18325 32250 18360
rect 32285 18325 32295 18360
rect 32330 18325 32340 18360
rect 32375 18325 32385 18360
rect 32420 18325 32430 18360
rect 32465 18325 32475 18360
rect 32510 18325 32520 18360
rect 32555 18325 32565 18360
rect 32600 18325 32610 18360
rect 32645 18325 32655 18360
rect 32690 18325 32700 18360
rect 32735 18325 32745 18360
rect 32780 18325 32790 18360
rect 32825 18325 32835 18360
rect 32870 18325 32890 18360
rect 31290 18315 32890 18325
rect 31290 18280 31305 18315
rect 31340 18280 31350 18315
rect 31385 18280 31395 18315
rect 31430 18280 31440 18315
rect 31475 18280 31485 18315
rect 31520 18280 31530 18315
rect 31565 18280 31575 18315
rect 31610 18280 31620 18315
rect 31655 18280 31665 18315
rect 31700 18280 31710 18315
rect 31745 18280 31755 18315
rect 31790 18280 31800 18315
rect 31835 18280 31845 18315
rect 31880 18280 31890 18315
rect 31925 18280 31935 18315
rect 31970 18280 31980 18315
rect 32015 18280 32025 18315
rect 32060 18280 32070 18315
rect 32105 18280 32115 18315
rect 32150 18280 32160 18315
rect 32195 18280 32205 18315
rect 32240 18280 32250 18315
rect 32285 18280 32295 18315
rect 32330 18280 32340 18315
rect 32375 18280 32385 18315
rect 32420 18280 32430 18315
rect 32465 18280 32475 18315
rect 32510 18280 32520 18315
rect 32555 18280 32565 18315
rect 32600 18280 32610 18315
rect 32645 18280 32655 18315
rect 32690 18280 32700 18315
rect 32735 18280 32745 18315
rect 32780 18280 32790 18315
rect 32825 18280 32835 18315
rect 32870 18280 32890 18315
rect 31290 18270 32890 18280
rect 31290 18235 31305 18270
rect 31340 18235 31350 18270
rect 31385 18235 31395 18270
rect 31430 18235 31440 18270
rect 31475 18235 31485 18270
rect 31520 18235 31530 18270
rect 31565 18235 31575 18270
rect 31610 18235 31620 18270
rect 31655 18235 31665 18270
rect 31700 18235 31710 18270
rect 31745 18235 31755 18270
rect 31790 18235 31800 18270
rect 31835 18235 31845 18270
rect 31880 18235 31890 18270
rect 31925 18235 31935 18270
rect 31970 18235 31980 18270
rect 32015 18235 32025 18270
rect 32060 18235 32070 18270
rect 32105 18235 32115 18270
rect 32150 18235 32160 18270
rect 32195 18235 32205 18270
rect 32240 18235 32250 18270
rect 32285 18235 32295 18270
rect 32330 18235 32340 18270
rect 32375 18235 32385 18270
rect 32420 18235 32430 18270
rect 32465 18235 32475 18270
rect 32510 18235 32520 18270
rect 32555 18235 32565 18270
rect 32600 18235 32610 18270
rect 32645 18235 32655 18270
rect 32690 18235 32700 18270
rect 32735 18235 32745 18270
rect 32780 18235 32790 18270
rect 32825 18235 32835 18270
rect 32870 18235 32890 18270
rect 31290 18225 32890 18235
rect 31290 18190 31305 18225
rect 31340 18190 31350 18225
rect 31385 18190 31395 18225
rect 31430 18190 31440 18225
rect 31475 18190 31485 18225
rect 31520 18190 31530 18225
rect 31565 18190 31575 18225
rect 31610 18190 31620 18225
rect 31655 18190 31665 18225
rect 31700 18190 31710 18225
rect 31745 18190 31755 18225
rect 31790 18190 31800 18225
rect 31835 18190 31845 18225
rect 31880 18190 31890 18225
rect 31925 18190 31935 18225
rect 31970 18190 31980 18225
rect 32015 18190 32025 18225
rect 32060 18190 32070 18225
rect 32105 18190 32115 18225
rect 32150 18190 32160 18225
rect 32195 18190 32205 18225
rect 32240 18190 32250 18225
rect 32285 18190 32295 18225
rect 32330 18190 32340 18225
rect 32375 18190 32385 18225
rect 32420 18190 32430 18225
rect 32465 18190 32475 18225
rect 32510 18190 32520 18225
rect 32555 18190 32565 18225
rect 32600 18190 32610 18225
rect 32645 18190 32655 18225
rect 32690 18190 32700 18225
rect 32735 18190 32745 18225
rect 32780 18190 32790 18225
rect 32825 18190 32835 18225
rect 32870 18190 32890 18225
rect 31290 18180 32890 18190
rect 31290 18145 31305 18180
rect 31340 18145 31350 18180
rect 31385 18145 31395 18180
rect 31430 18145 31440 18180
rect 31475 18145 31485 18180
rect 31520 18145 31530 18180
rect 31565 18145 31575 18180
rect 31610 18145 31620 18180
rect 31655 18145 31665 18180
rect 31700 18145 31710 18180
rect 31745 18145 31755 18180
rect 31790 18145 31800 18180
rect 31835 18145 31845 18180
rect 31880 18145 31890 18180
rect 31925 18145 31935 18180
rect 31970 18145 31980 18180
rect 32015 18145 32025 18180
rect 32060 18145 32070 18180
rect 32105 18145 32115 18180
rect 32150 18145 32160 18180
rect 32195 18145 32205 18180
rect 32240 18145 32250 18180
rect 32285 18145 32295 18180
rect 32330 18145 32340 18180
rect 32375 18145 32385 18180
rect 32420 18145 32430 18180
rect 32465 18145 32475 18180
rect 32510 18145 32520 18180
rect 32555 18145 32565 18180
rect 32600 18145 32610 18180
rect 32645 18145 32655 18180
rect 32690 18145 32700 18180
rect 32735 18145 32745 18180
rect 32780 18145 32790 18180
rect 32825 18145 32835 18180
rect 32870 18145 32890 18180
rect 31290 18135 32890 18145
rect 31290 18100 31305 18135
rect 31340 18100 31350 18135
rect 31385 18100 31395 18135
rect 31430 18100 31440 18135
rect 31475 18100 31485 18135
rect 31520 18100 31530 18135
rect 31565 18100 31575 18135
rect 31610 18100 31620 18135
rect 31655 18100 31665 18135
rect 31700 18100 31710 18135
rect 31745 18100 31755 18135
rect 31790 18100 31800 18135
rect 31835 18100 31845 18135
rect 31880 18100 31890 18135
rect 31925 18100 31935 18135
rect 31970 18100 31980 18135
rect 32015 18100 32025 18135
rect 32060 18100 32070 18135
rect 32105 18100 32115 18135
rect 32150 18100 32160 18135
rect 32195 18100 32205 18135
rect 32240 18100 32250 18135
rect 32285 18100 32295 18135
rect 32330 18100 32340 18135
rect 32375 18100 32385 18135
rect 32420 18100 32430 18135
rect 32465 18100 32475 18135
rect 32510 18100 32520 18135
rect 32555 18100 32565 18135
rect 32600 18100 32610 18135
rect 32645 18100 32655 18135
rect 32690 18100 32700 18135
rect 32735 18100 32745 18135
rect 32780 18100 32790 18135
rect 32825 18100 32835 18135
rect 32870 18100 32890 18135
rect 31290 18090 32890 18100
rect 31290 18055 31305 18090
rect 31340 18055 31350 18090
rect 31385 18055 31395 18090
rect 31430 18055 31440 18090
rect 31475 18055 31485 18090
rect 31520 18055 31530 18090
rect 31565 18055 31575 18090
rect 31610 18055 31620 18090
rect 31655 18055 31665 18090
rect 31700 18055 31710 18090
rect 31745 18055 31755 18090
rect 31790 18055 31800 18090
rect 31835 18055 31845 18090
rect 31880 18055 31890 18090
rect 31925 18055 31935 18090
rect 31970 18055 31980 18090
rect 32015 18055 32025 18090
rect 32060 18055 32070 18090
rect 32105 18055 32115 18090
rect 32150 18055 32160 18090
rect 32195 18055 32205 18090
rect 32240 18055 32250 18090
rect 32285 18055 32295 18090
rect 32330 18055 32340 18090
rect 32375 18055 32385 18090
rect 32420 18055 32430 18090
rect 32465 18055 32475 18090
rect 32510 18055 32520 18090
rect 32555 18055 32565 18090
rect 32600 18055 32610 18090
rect 32645 18055 32655 18090
rect 32690 18055 32700 18090
rect 32735 18055 32745 18090
rect 32780 18055 32790 18090
rect 32825 18055 32835 18090
rect 32870 18055 32890 18090
rect 31290 18045 32890 18055
rect 31290 18010 31305 18045
rect 31340 18010 31350 18045
rect 31385 18010 31395 18045
rect 31430 18010 31440 18045
rect 31475 18010 31485 18045
rect 31520 18010 31530 18045
rect 31565 18010 31575 18045
rect 31610 18010 31620 18045
rect 31655 18010 31665 18045
rect 31700 18010 31710 18045
rect 31745 18010 31755 18045
rect 31790 18010 31800 18045
rect 31835 18010 31845 18045
rect 31880 18010 31890 18045
rect 31925 18010 31935 18045
rect 31970 18010 31980 18045
rect 32015 18010 32025 18045
rect 32060 18010 32070 18045
rect 32105 18010 32115 18045
rect 32150 18010 32160 18045
rect 32195 18010 32205 18045
rect 32240 18010 32250 18045
rect 32285 18010 32295 18045
rect 32330 18010 32340 18045
rect 32375 18010 32385 18045
rect 32420 18010 32430 18045
rect 32465 18010 32475 18045
rect 32510 18010 32520 18045
rect 32555 18010 32565 18045
rect 32600 18010 32610 18045
rect 32645 18010 32655 18045
rect 32690 18010 32700 18045
rect 32735 18010 32745 18045
rect 32780 18010 32790 18045
rect 32825 18010 32835 18045
rect 32870 18010 32890 18045
rect 31290 18000 32890 18010
rect 31290 17965 31305 18000
rect 31340 17965 31350 18000
rect 31385 17965 31395 18000
rect 31430 17965 31440 18000
rect 31475 17965 31485 18000
rect 31520 17965 31530 18000
rect 31565 17965 31575 18000
rect 31610 17965 31620 18000
rect 31655 17965 31665 18000
rect 31700 17965 31710 18000
rect 31745 17965 31755 18000
rect 31790 17965 31800 18000
rect 31835 17965 31845 18000
rect 31880 17965 31890 18000
rect 31925 17965 31935 18000
rect 31970 17965 31980 18000
rect 32015 17965 32025 18000
rect 32060 17965 32070 18000
rect 32105 17965 32115 18000
rect 32150 17965 32160 18000
rect 32195 17965 32205 18000
rect 32240 17965 32250 18000
rect 32285 17965 32295 18000
rect 32330 17965 32340 18000
rect 32375 17965 32385 18000
rect 32420 17965 32430 18000
rect 32465 17965 32475 18000
rect 32510 17965 32520 18000
rect 32555 17965 32565 18000
rect 32600 17965 32610 18000
rect 32645 17965 32655 18000
rect 32690 17965 32700 18000
rect 32735 17965 32745 18000
rect 32780 17965 32790 18000
rect 32825 17965 32835 18000
rect 32870 17965 32890 18000
rect 31290 17955 32890 17965
rect 31290 17920 31305 17955
rect 31340 17920 31350 17955
rect 31385 17920 31395 17955
rect 31430 17920 31440 17955
rect 31475 17920 31485 17955
rect 31520 17920 31530 17955
rect 31565 17920 31575 17955
rect 31610 17920 31620 17955
rect 31655 17920 31665 17955
rect 31700 17920 31710 17955
rect 31745 17920 31755 17955
rect 31790 17920 31800 17955
rect 31835 17920 31845 17955
rect 31880 17920 31890 17955
rect 31925 17920 31935 17955
rect 31970 17920 31980 17955
rect 32015 17920 32025 17955
rect 32060 17920 32070 17955
rect 32105 17920 32115 17955
rect 32150 17920 32160 17955
rect 32195 17920 32205 17955
rect 32240 17920 32250 17955
rect 32285 17920 32295 17955
rect 32330 17920 32340 17955
rect 32375 17920 32385 17955
rect 32420 17920 32430 17955
rect 32465 17920 32475 17955
rect 32510 17920 32520 17955
rect 32555 17920 32565 17955
rect 32600 17920 32610 17955
rect 32645 17920 32655 17955
rect 32690 17920 32700 17955
rect 32735 17920 32745 17955
rect 32780 17920 32790 17955
rect 32825 17920 32835 17955
rect 32870 17920 32890 17955
rect 31290 17910 32890 17920
rect 31290 17875 31305 17910
rect 31340 17875 31350 17910
rect 31385 17875 31395 17910
rect 31430 17875 31440 17910
rect 31475 17875 31485 17910
rect 31520 17875 31530 17910
rect 31565 17875 31575 17910
rect 31610 17875 31620 17910
rect 31655 17875 31665 17910
rect 31700 17875 31710 17910
rect 31745 17875 31755 17910
rect 31790 17875 31800 17910
rect 31835 17875 31845 17910
rect 31880 17875 31890 17910
rect 31925 17875 31935 17910
rect 31970 17875 31980 17910
rect 32015 17875 32025 17910
rect 32060 17875 32070 17910
rect 32105 17875 32115 17910
rect 32150 17875 32160 17910
rect 32195 17875 32205 17910
rect 32240 17875 32250 17910
rect 32285 17875 32295 17910
rect 32330 17875 32340 17910
rect 32375 17875 32385 17910
rect 32420 17875 32430 17910
rect 32465 17875 32475 17910
rect 32510 17875 32520 17910
rect 32555 17875 32565 17910
rect 32600 17875 32610 17910
rect 32645 17875 32655 17910
rect 32690 17875 32700 17910
rect 32735 17875 32745 17910
rect 32780 17875 32790 17910
rect 32825 17875 32835 17910
rect 32870 17875 32890 17910
rect 31290 17865 32890 17875
rect 31290 17830 31305 17865
rect 31340 17830 31350 17865
rect 31385 17830 31395 17865
rect 31430 17830 31440 17865
rect 31475 17830 31485 17865
rect 31520 17830 31530 17865
rect 31565 17830 31575 17865
rect 31610 17830 31620 17865
rect 31655 17830 31665 17865
rect 31700 17830 31710 17865
rect 31745 17830 31755 17865
rect 31790 17830 31800 17865
rect 31835 17830 31845 17865
rect 31880 17830 31890 17865
rect 31925 17830 31935 17865
rect 31970 17830 31980 17865
rect 32015 17830 32025 17865
rect 32060 17830 32070 17865
rect 32105 17830 32115 17865
rect 32150 17830 32160 17865
rect 32195 17830 32205 17865
rect 32240 17830 32250 17865
rect 32285 17830 32295 17865
rect 32330 17830 32340 17865
rect 32375 17830 32385 17865
rect 32420 17830 32430 17865
rect 32465 17830 32475 17865
rect 32510 17830 32520 17865
rect 32555 17830 32565 17865
rect 32600 17830 32610 17865
rect 32645 17830 32655 17865
rect 32690 17830 32700 17865
rect 32735 17830 32745 17865
rect 32780 17830 32790 17865
rect 32825 17830 32835 17865
rect 32870 17830 32890 17865
rect 31290 17820 32890 17830
rect 31290 17785 31305 17820
rect 31340 17785 31350 17820
rect 31385 17785 31395 17820
rect 31430 17785 31440 17820
rect 31475 17785 31485 17820
rect 31520 17785 31530 17820
rect 31565 17785 31575 17820
rect 31610 17785 31620 17820
rect 31655 17785 31665 17820
rect 31700 17785 31710 17820
rect 31745 17785 31755 17820
rect 31790 17785 31800 17820
rect 31835 17785 31845 17820
rect 31880 17785 31890 17820
rect 31925 17785 31935 17820
rect 31970 17785 31980 17820
rect 32015 17785 32025 17820
rect 32060 17785 32070 17820
rect 32105 17785 32115 17820
rect 32150 17785 32160 17820
rect 32195 17785 32205 17820
rect 32240 17785 32250 17820
rect 32285 17785 32295 17820
rect 32330 17785 32340 17820
rect 32375 17785 32385 17820
rect 32420 17785 32430 17820
rect 32465 17785 32475 17820
rect 32510 17785 32520 17820
rect 32555 17785 32565 17820
rect 32600 17785 32610 17820
rect 32645 17785 32655 17820
rect 32690 17785 32700 17820
rect 32735 17785 32745 17820
rect 32780 17785 32790 17820
rect 32825 17785 32835 17820
rect 32870 17785 32890 17820
rect 31290 17775 32890 17785
rect 31290 17740 31305 17775
rect 31340 17740 31350 17775
rect 31385 17740 31395 17775
rect 31430 17740 31440 17775
rect 31475 17740 31485 17775
rect 31520 17740 31530 17775
rect 31565 17740 31575 17775
rect 31610 17740 31620 17775
rect 31655 17740 31665 17775
rect 31700 17740 31710 17775
rect 31745 17740 31755 17775
rect 31790 17740 31800 17775
rect 31835 17740 31845 17775
rect 31880 17740 31890 17775
rect 31925 17740 31935 17775
rect 31970 17740 31980 17775
rect 32015 17740 32025 17775
rect 32060 17740 32070 17775
rect 32105 17740 32115 17775
rect 32150 17740 32160 17775
rect 32195 17740 32205 17775
rect 32240 17740 32250 17775
rect 32285 17740 32295 17775
rect 32330 17740 32340 17775
rect 32375 17740 32385 17775
rect 32420 17740 32430 17775
rect 32465 17740 32475 17775
rect 32510 17740 32520 17775
rect 32555 17740 32565 17775
rect 32600 17740 32610 17775
rect 32645 17740 32655 17775
rect 32690 17740 32700 17775
rect 32735 17740 32745 17775
rect 32780 17740 32790 17775
rect 32825 17740 32835 17775
rect 32870 17740 32890 17775
rect -38770 9630 -37170 10155
rect -38770 9595 -38755 9630
rect -38720 9595 -38710 9630
rect -38675 9595 -38665 9630
rect -38630 9595 -38620 9630
rect -38585 9595 -38575 9630
rect -38540 9595 -38530 9630
rect -38495 9595 -38485 9630
rect -38450 9595 -38440 9630
rect -38405 9595 -38395 9630
rect -38360 9595 -38350 9630
rect -38315 9595 -38305 9630
rect -38270 9595 -38260 9630
rect -38225 9595 -38215 9630
rect -38180 9595 -38170 9630
rect -38135 9595 -38125 9630
rect -38090 9595 -38080 9630
rect -38045 9595 -38035 9630
rect -38000 9595 -37990 9630
rect -37955 9595 -37945 9630
rect -37910 9595 -37900 9630
rect -37865 9595 -37855 9630
rect -37820 9595 -37810 9630
rect -37775 9595 -37765 9630
rect -37730 9595 -37720 9630
rect -37685 9595 -37675 9630
rect -37640 9595 -37630 9630
rect -37595 9595 -37585 9630
rect -37550 9595 -37540 9630
rect -37505 9595 -37495 9630
rect -37460 9595 -37450 9630
rect -37415 9595 -37405 9630
rect -37370 9595 -37360 9630
rect -37325 9595 -37315 9630
rect -37280 9595 -37270 9630
rect -37235 9595 -37225 9630
rect -37190 9595 -37170 9630
rect -38770 9585 -37170 9595
rect -38770 9550 -38755 9585
rect -38720 9550 -38710 9585
rect -38675 9550 -38665 9585
rect -38630 9550 -38620 9585
rect -38585 9550 -38575 9585
rect -38540 9550 -38530 9585
rect -38495 9550 -38485 9585
rect -38450 9550 -38440 9585
rect -38405 9550 -38395 9585
rect -38360 9550 -38350 9585
rect -38315 9550 -38305 9585
rect -38270 9550 -38260 9585
rect -38225 9550 -38215 9585
rect -38180 9550 -38170 9585
rect -38135 9550 -38125 9585
rect -38090 9550 -38080 9585
rect -38045 9550 -38035 9585
rect -38000 9550 -37990 9585
rect -37955 9550 -37945 9585
rect -37910 9550 -37900 9585
rect -37865 9550 -37855 9585
rect -37820 9550 -37810 9585
rect -37775 9550 -37765 9585
rect -37730 9550 -37720 9585
rect -37685 9550 -37675 9585
rect -37640 9550 -37630 9585
rect -37595 9550 -37585 9585
rect -37550 9550 -37540 9585
rect -37505 9550 -37495 9585
rect -37460 9550 -37450 9585
rect -37415 9550 -37405 9585
rect -37370 9550 -37360 9585
rect -37325 9550 -37315 9585
rect -37280 9550 -37270 9585
rect -37235 9550 -37225 9585
rect -37190 9550 -37170 9585
rect -38770 9540 -37170 9550
rect -38770 9505 -38755 9540
rect -38720 9505 -38710 9540
rect -38675 9505 -38665 9540
rect -38630 9505 -38620 9540
rect -38585 9505 -38575 9540
rect -38540 9505 -38530 9540
rect -38495 9505 -38485 9540
rect -38450 9505 -38440 9540
rect -38405 9505 -38395 9540
rect -38360 9505 -38350 9540
rect -38315 9505 -38305 9540
rect -38270 9505 -38260 9540
rect -38225 9505 -38215 9540
rect -38180 9505 -38170 9540
rect -38135 9505 -38125 9540
rect -38090 9505 -38080 9540
rect -38045 9505 -38035 9540
rect -38000 9505 -37990 9540
rect -37955 9505 -37945 9540
rect -37910 9505 -37900 9540
rect -37865 9505 -37855 9540
rect -37820 9505 -37810 9540
rect -37775 9505 -37765 9540
rect -37730 9505 -37720 9540
rect -37685 9505 -37675 9540
rect -37640 9505 -37630 9540
rect -37595 9505 -37585 9540
rect -37550 9505 -37540 9540
rect -37505 9505 -37495 9540
rect -37460 9505 -37450 9540
rect -37415 9505 -37405 9540
rect -37370 9505 -37360 9540
rect -37325 9505 -37315 9540
rect -37280 9505 -37270 9540
rect -37235 9505 -37225 9540
rect -37190 9505 -37170 9540
rect -38770 9495 -37170 9505
rect -38770 9460 -38755 9495
rect -38720 9460 -38710 9495
rect -38675 9460 -38665 9495
rect -38630 9460 -38620 9495
rect -38585 9460 -38575 9495
rect -38540 9460 -38530 9495
rect -38495 9460 -38485 9495
rect -38450 9460 -38440 9495
rect -38405 9460 -38395 9495
rect -38360 9460 -38350 9495
rect -38315 9460 -38305 9495
rect -38270 9460 -38260 9495
rect -38225 9460 -38215 9495
rect -38180 9460 -38170 9495
rect -38135 9460 -38125 9495
rect -38090 9460 -38080 9495
rect -38045 9460 -38035 9495
rect -38000 9460 -37990 9495
rect -37955 9460 -37945 9495
rect -37910 9460 -37900 9495
rect -37865 9460 -37855 9495
rect -37820 9460 -37810 9495
rect -37775 9460 -37765 9495
rect -37730 9460 -37720 9495
rect -37685 9460 -37675 9495
rect -37640 9460 -37630 9495
rect -37595 9460 -37585 9495
rect -37550 9460 -37540 9495
rect -37505 9460 -37495 9495
rect -37460 9460 -37450 9495
rect -37415 9460 -37405 9495
rect -37370 9460 -37360 9495
rect -37325 9460 -37315 9495
rect -37280 9460 -37270 9495
rect -37235 9460 -37225 9495
rect -37190 9460 -37170 9495
rect -38770 9450 -37170 9460
rect -38770 9415 -38755 9450
rect -38720 9415 -38710 9450
rect -38675 9415 -38665 9450
rect -38630 9415 -38620 9450
rect -38585 9415 -38575 9450
rect -38540 9415 -38530 9450
rect -38495 9415 -38485 9450
rect -38450 9415 -38440 9450
rect -38405 9415 -38395 9450
rect -38360 9415 -38350 9450
rect -38315 9415 -38305 9450
rect -38270 9415 -38260 9450
rect -38225 9415 -38215 9450
rect -38180 9415 -38170 9450
rect -38135 9415 -38125 9450
rect -38090 9415 -38080 9450
rect -38045 9415 -38035 9450
rect -38000 9415 -37990 9450
rect -37955 9415 -37945 9450
rect -37910 9415 -37900 9450
rect -37865 9415 -37855 9450
rect -37820 9415 -37810 9450
rect -37775 9415 -37765 9450
rect -37730 9415 -37720 9450
rect -37685 9415 -37675 9450
rect -37640 9415 -37630 9450
rect -37595 9415 -37585 9450
rect -37550 9415 -37540 9450
rect -37505 9415 -37495 9450
rect -37460 9415 -37450 9450
rect -37415 9415 -37405 9450
rect -37370 9415 -37360 9450
rect -37325 9415 -37315 9450
rect -37280 9415 -37270 9450
rect -37235 9415 -37225 9450
rect -37190 9415 -37170 9450
rect -38770 9405 -37170 9415
rect -38770 9370 -38755 9405
rect -38720 9370 -38710 9405
rect -38675 9370 -38665 9405
rect -38630 9370 -38620 9405
rect -38585 9370 -38575 9405
rect -38540 9370 -38530 9405
rect -38495 9370 -38485 9405
rect -38450 9370 -38440 9405
rect -38405 9370 -38395 9405
rect -38360 9370 -38350 9405
rect -38315 9370 -38305 9405
rect -38270 9370 -38260 9405
rect -38225 9370 -38215 9405
rect -38180 9370 -38170 9405
rect -38135 9370 -38125 9405
rect -38090 9370 -38080 9405
rect -38045 9370 -38035 9405
rect -38000 9370 -37990 9405
rect -37955 9370 -37945 9405
rect -37910 9370 -37900 9405
rect -37865 9370 -37855 9405
rect -37820 9370 -37810 9405
rect -37775 9370 -37765 9405
rect -37730 9370 -37720 9405
rect -37685 9370 -37675 9405
rect -37640 9370 -37630 9405
rect -37595 9370 -37585 9405
rect -37550 9370 -37540 9405
rect -37505 9370 -37495 9405
rect -37460 9370 -37450 9405
rect -37415 9370 -37405 9405
rect -37370 9370 -37360 9405
rect -37325 9370 -37315 9405
rect -37280 9370 -37270 9405
rect -37235 9370 -37225 9405
rect -37190 9370 -37170 9405
rect -38770 9360 -37170 9370
rect -38770 9325 -38755 9360
rect -38720 9325 -38710 9360
rect -38675 9325 -38665 9360
rect -38630 9325 -38620 9360
rect -38585 9325 -38575 9360
rect -38540 9325 -38530 9360
rect -38495 9325 -38485 9360
rect -38450 9325 -38440 9360
rect -38405 9325 -38395 9360
rect -38360 9325 -38350 9360
rect -38315 9325 -38305 9360
rect -38270 9325 -38260 9360
rect -38225 9325 -38215 9360
rect -38180 9325 -38170 9360
rect -38135 9325 -38125 9360
rect -38090 9325 -38080 9360
rect -38045 9325 -38035 9360
rect -38000 9325 -37990 9360
rect -37955 9325 -37945 9360
rect -37910 9325 -37900 9360
rect -37865 9325 -37855 9360
rect -37820 9325 -37810 9360
rect -37775 9325 -37765 9360
rect -37730 9325 -37720 9360
rect -37685 9325 -37675 9360
rect -37640 9325 -37630 9360
rect -37595 9325 -37585 9360
rect -37550 9325 -37540 9360
rect -37505 9325 -37495 9360
rect -37460 9325 -37450 9360
rect -37415 9325 -37405 9360
rect -37370 9325 -37360 9360
rect -37325 9325 -37315 9360
rect -37280 9325 -37270 9360
rect -37235 9325 -37225 9360
rect -37190 9325 -37170 9360
rect -38770 9315 -37170 9325
rect -38770 9280 -38755 9315
rect -38720 9280 -38710 9315
rect -38675 9280 -38665 9315
rect -38630 9280 -38620 9315
rect -38585 9280 -38575 9315
rect -38540 9280 -38530 9315
rect -38495 9280 -38485 9315
rect -38450 9280 -38440 9315
rect -38405 9280 -38395 9315
rect -38360 9280 -38350 9315
rect -38315 9280 -38305 9315
rect -38270 9280 -38260 9315
rect -38225 9280 -38215 9315
rect -38180 9280 -38170 9315
rect -38135 9280 -38125 9315
rect -38090 9280 -38080 9315
rect -38045 9280 -38035 9315
rect -38000 9280 -37990 9315
rect -37955 9280 -37945 9315
rect -37910 9280 -37900 9315
rect -37865 9280 -37855 9315
rect -37820 9280 -37810 9315
rect -37775 9280 -37765 9315
rect -37730 9280 -37720 9315
rect -37685 9280 -37675 9315
rect -37640 9280 -37630 9315
rect -37595 9280 -37585 9315
rect -37550 9280 -37540 9315
rect -37505 9280 -37495 9315
rect -37460 9280 -37450 9315
rect -37415 9280 -37405 9315
rect -37370 9280 -37360 9315
rect -37325 9280 -37315 9315
rect -37280 9280 -37270 9315
rect -37235 9280 -37225 9315
rect -37190 9280 -37170 9315
rect -38770 9270 -37170 9280
rect -38770 9235 -38755 9270
rect -38720 9235 -38710 9270
rect -38675 9235 -38665 9270
rect -38630 9235 -38620 9270
rect -38585 9235 -38575 9270
rect -38540 9235 -38530 9270
rect -38495 9235 -38485 9270
rect -38450 9235 -38440 9270
rect -38405 9235 -38395 9270
rect -38360 9235 -38350 9270
rect -38315 9235 -38305 9270
rect -38270 9235 -38260 9270
rect -38225 9235 -38215 9270
rect -38180 9235 -38170 9270
rect -38135 9235 -38125 9270
rect -38090 9235 -38080 9270
rect -38045 9235 -38035 9270
rect -38000 9235 -37990 9270
rect -37955 9235 -37945 9270
rect -37910 9235 -37900 9270
rect -37865 9235 -37855 9270
rect -37820 9235 -37810 9270
rect -37775 9235 -37765 9270
rect -37730 9235 -37720 9270
rect -37685 9235 -37675 9270
rect -37640 9235 -37630 9270
rect -37595 9235 -37585 9270
rect -37550 9235 -37540 9270
rect -37505 9235 -37495 9270
rect -37460 9235 -37450 9270
rect -37415 9235 -37405 9270
rect -37370 9235 -37360 9270
rect -37325 9235 -37315 9270
rect -37280 9235 -37270 9270
rect -37235 9235 -37225 9270
rect -37190 9235 -37170 9270
rect -38770 9225 -37170 9235
rect -38770 9190 -38755 9225
rect -38720 9190 -38710 9225
rect -38675 9190 -38665 9225
rect -38630 9190 -38620 9225
rect -38585 9190 -38575 9225
rect -38540 9190 -38530 9225
rect -38495 9190 -38485 9225
rect -38450 9190 -38440 9225
rect -38405 9190 -38395 9225
rect -38360 9190 -38350 9225
rect -38315 9190 -38305 9225
rect -38270 9190 -38260 9225
rect -38225 9190 -38215 9225
rect -38180 9190 -38170 9225
rect -38135 9190 -38125 9225
rect -38090 9190 -38080 9225
rect -38045 9190 -38035 9225
rect -38000 9190 -37990 9225
rect -37955 9190 -37945 9225
rect -37910 9190 -37900 9225
rect -37865 9190 -37855 9225
rect -37820 9190 -37810 9225
rect -37775 9190 -37765 9225
rect -37730 9190 -37720 9225
rect -37685 9190 -37675 9225
rect -37640 9190 -37630 9225
rect -37595 9190 -37585 9225
rect -37550 9190 -37540 9225
rect -37505 9190 -37495 9225
rect -37460 9190 -37450 9225
rect -37415 9190 -37405 9225
rect -37370 9190 -37360 9225
rect -37325 9190 -37315 9225
rect -37280 9190 -37270 9225
rect -37235 9190 -37225 9225
rect -37190 9190 -37170 9225
rect -38770 9180 -37170 9190
rect -38770 9145 -38755 9180
rect -38720 9145 -38710 9180
rect -38675 9145 -38665 9180
rect -38630 9145 -38620 9180
rect -38585 9145 -38575 9180
rect -38540 9145 -38530 9180
rect -38495 9145 -38485 9180
rect -38450 9145 -38440 9180
rect -38405 9145 -38395 9180
rect -38360 9145 -38350 9180
rect -38315 9145 -38305 9180
rect -38270 9145 -38260 9180
rect -38225 9145 -38215 9180
rect -38180 9145 -38170 9180
rect -38135 9145 -38125 9180
rect -38090 9145 -38080 9180
rect -38045 9145 -38035 9180
rect -38000 9145 -37990 9180
rect -37955 9145 -37945 9180
rect -37910 9145 -37900 9180
rect -37865 9145 -37855 9180
rect -37820 9145 -37810 9180
rect -37775 9145 -37765 9180
rect -37730 9145 -37720 9180
rect -37685 9145 -37675 9180
rect -37640 9145 -37630 9180
rect -37595 9145 -37585 9180
rect -37550 9145 -37540 9180
rect -37505 9145 -37495 9180
rect -37460 9145 -37450 9180
rect -37415 9145 -37405 9180
rect -37370 9145 -37360 9180
rect -37325 9145 -37315 9180
rect -37280 9145 -37270 9180
rect -37235 9145 -37225 9180
rect -37190 9145 -37170 9180
rect -38770 9135 -37170 9145
rect -38770 9100 -38755 9135
rect -38720 9100 -38710 9135
rect -38675 9100 -38665 9135
rect -38630 9100 -38620 9135
rect -38585 9100 -38575 9135
rect -38540 9100 -38530 9135
rect -38495 9100 -38485 9135
rect -38450 9100 -38440 9135
rect -38405 9100 -38395 9135
rect -38360 9100 -38350 9135
rect -38315 9100 -38305 9135
rect -38270 9100 -38260 9135
rect -38225 9100 -38215 9135
rect -38180 9100 -38170 9135
rect -38135 9100 -38125 9135
rect -38090 9100 -38080 9135
rect -38045 9100 -38035 9135
rect -38000 9100 -37990 9135
rect -37955 9100 -37945 9135
rect -37910 9100 -37900 9135
rect -37865 9100 -37855 9135
rect -37820 9100 -37810 9135
rect -37775 9100 -37765 9135
rect -37730 9100 -37720 9135
rect -37685 9100 -37675 9135
rect -37640 9100 -37630 9135
rect -37595 9100 -37585 9135
rect -37550 9100 -37540 9135
rect -37505 9100 -37495 9135
rect -37460 9100 -37450 9135
rect -37415 9100 -37405 9135
rect -37370 9100 -37360 9135
rect -37325 9100 -37315 9135
rect -37280 9100 -37270 9135
rect -37235 9100 -37225 9135
rect -37190 9100 -37170 9135
rect -38770 9090 -37170 9100
rect -38770 9055 -38755 9090
rect -38720 9055 -38710 9090
rect -38675 9055 -38665 9090
rect -38630 9055 -38620 9090
rect -38585 9055 -38575 9090
rect -38540 9055 -38530 9090
rect -38495 9055 -38485 9090
rect -38450 9055 -38440 9090
rect -38405 9055 -38395 9090
rect -38360 9055 -38350 9090
rect -38315 9055 -38305 9090
rect -38270 9055 -38260 9090
rect -38225 9055 -38215 9090
rect -38180 9055 -38170 9090
rect -38135 9055 -38125 9090
rect -38090 9055 -38080 9090
rect -38045 9055 -38035 9090
rect -38000 9055 -37990 9090
rect -37955 9055 -37945 9090
rect -37910 9055 -37900 9090
rect -37865 9055 -37855 9090
rect -37820 9055 -37810 9090
rect -37775 9055 -37765 9090
rect -37730 9055 -37720 9090
rect -37685 9055 -37675 9090
rect -37640 9055 -37630 9090
rect -37595 9055 -37585 9090
rect -37550 9055 -37540 9090
rect -37505 9055 -37495 9090
rect -37460 9055 -37450 9090
rect -37415 9055 -37405 9090
rect -37370 9055 -37360 9090
rect -37325 9055 -37315 9090
rect -37280 9055 -37270 9090
rect -37235 9055 -37225 9090
rect -37190 9055 -37170 9090
rect -38770 9045 -37170 9055
rect -38770 9010 -38755 9045
rect -38720 9010 -38710 9045
rect -38675 9010 -38665 9045
rect -38630 9010 -38620 9045
rect -38585 9010 -38575 9045
rect -38540 9010 -38530 9045
rect -38495 9010 -38485 9045
rect -38450 9010 -38440 9045
rect -38405 9010 -38395 9045
rect -38360 9010 -38350 9045
rect -38315 9010 -38305 9045
rect -38270 9010 -38260 9045
rect -38225 9010 -38215 9045
rect -38180 9010 -38170 9045
rect -38135 9010 -38125 9045
rect -38090 9010 -38080 9045
rect -38045 9010 -38035 9045
rect -38000 9010 -37990 9045
rect -37955 9010 -37945 9045
rect -37910 9010 -37900 9045
rect -37865 9010 -37855 9045
rect -37820 9010 -37810 9045
rect -37775 9010 -37765 9045
rect -37730 9010 -37720 9045
rect -37685 9010 -37675 9045
rect -37640 9010 -37630 9045
rect -37595 9010 -37585 9045
rect -37550 9010 -37540 9045
rect -37505 9010 -37495 9045
rect -37460 9010 -37450 9045
rect -37415 9010 -37405 9045
rect -37370 9010 -37360 9045
rect -37325 9010 -37315 9045
rect -37280 9010 -37270 9045
rect -37235 9010 -37225 9045
rect -37190 9010 -37170 9045
rect -38770 9000 -37170 9010
rect -38770 8965 -38755 9000
rect -38720 8965 -38710 9000
rect -38675 8965 -38665 9000
rect -38630 8965 -38620 9000
rect -38585 8965 -38575 9000
rect -38540 8965 -38530 9000
rect -38495 8965 -38485 9000
rect -38450 8965 -38440 9000
rect -38405 8965 -38395 9000
rect -38360 8965 -38350 9000
rect -38315 8965 -38305 9000
rect -38270 8965 -38260 9000
rect -38225 8965 -38215 9000
rect -38180 8965 -38170 9000
rect -38135 8965 -38125 9000
rect -38090 8965 -38080 9000
rect -38045 8965 -38035 9000
rect -38000 8965 -37990 9000
rect -37955 8965 -37945 9000
rect -37910 8965 -37900 9000
rect -37865 8965 -37855 9000
rect -37820 8965 -37810 9000
rect -37775 8965 -37765 9000
rect -37730 8965 -37720 9000
rect -37685 8965 -37675 9000
rect -37640 8965 -37630 9000
rect -37595 8965 -37585 9000
rect -37550 8965 -37540 9000
rect -37505 8965 -37495 9000
rect -37460 8965 -37450 9000
rect -37415 8965 -37405 9000
rect -37370 8965 -37360 9000
rect -37325 8965 -37315 9000
rect -37280 8965 -37270 9000
rect -37235 8965 -37225 9000
rect -37190 8965 -37170 9000
rect -38770 8955 -37170 8965
rect -38770 8920 -38755 8955
rect -38720 8920 -38710 8955
rect -38675 8920 -38665 8955
rect -38630 8920 -38620 8955
rect -38585 8920 -38575 8955
rect -38540 8920 -38530 8955
rect -38495 8920 -38485 8955
rect -38450 8920 -38440 8955
rect -38405 8920 -38395 8955
rect -38360 8920 -38350 8955
rect -38315 8920 -38305 8955
rect -38270 8920 -38260 8955
rect -38225 8920 -38215 8955
rect -38180 8920 -38170 8955
rect -38135 8920 -38125 8955
rect -38090 8920 -38080 8955
rect -38045 8920 -38035 8955
rect -38000 8920 -37990 8955
rect -37955 8920 -37945 8955
rect -37910 8920 -37900 8955
rect -37865 8920 -37855 8955
rect -37820 8920 -37810 8955
rect -37775 8920 -37765 8955
rect -37730 8920 -37720 8955
rect -37685 8920 -37675 8955
rect -37640 8920 -37630 8955
rect -37595 8920 -37585 8955
rect -37550 8920 -37540 8955
rect -37505 8920 -37495 8955
rect -37460 8920 -37450 8955
rect -37415 8920 -37405 8955
rect -37370 8920 -37360 8955
rect -37325 8920 -37315 8955
rect -37280 8920 -37270 8955
rect -37235 8920 -37225 8955
rect -37190 8920 -37170 8955
rect -38770 8910 -37170 8920
rect -38770 8875 -38755 8910
rect -38720 8875 -38710 8910
rect -38675 8875 -38665 8910
rect -38630 8875 -38620 8910
rect -38585 8875 -38575 8910
rect -38540 8875 -38530 8910
rect -38495 8875 -38485 8910
rect -38450 8875 -38440 8910
rect -38405 8875 -38395 8910
rect -38360 8875 -38350 8910
rect -38315 8875 -38305 8910
rect -38270 8875 -38260 8910
rect -38225 8875 -38215 8910
rect -38180 8875 -38170 8910
rect -38135 8875 -38125 8910
rect -38090 8875 -38080 8910
rect -38045 8875 -38035 8910
rect -38000 8875 -37990 8910
rect -37955 8875 -37945 8910
rect -37910 8875 -37900 8910
rect -37865 8875 -37855 8910
rect -37820 8875 -37810 8910
rect -37775 8875 -37765 8910
rect -37730 8875 -37720 8910
rect -37685 8875 -37675 8910
rect -37640 8875 -37630 8910
rect -37595 8875 -37585 8910
rect -37550 8875 -37540 8910
rect -37505 8875 -37495 8910
rect -37460 8875 -37450 8910
rect -37415 8875 -37405 8910
rect -37370 8875 -37360 8910
rect -37325 8875 -37315 8910
rect -37280 8875 -37270 8910
rect -37235 8875 -37225 8910
rect -37190 8875 -37170 8910
rect -38770 8865 -37170 8875
rect -38770 8830 -38755 8865
rect -38720 8830 -38710 8865
rect -38675 8830 -38665 8865
rect -38630 8830 -38620 8865
rect -38585 8830 -38575 8865
rect -38540 8830 -38530 8865
rect -38495 8830 -38485 8865
rect -38450 8830 -38440 8865
rect -38405 8830 -38395 8865
rect -38360 8830 -38350 8865
rect -38315 8830 -38305 8865
rect -38270 8830 -38260 8865
rect -38225 8830 -38215 8865
rect -38180 8830 -38170 8865
rect -38135 8830 -38125 8865
rect -38090 8830 -38080 8865
rect -38045 8830 -38035 8865
rect -38000 8830 -37990 8865
rect -37955 8830 -37945 8865
rect -37910 8830 -37900 8865
rect -37865 8830 -37855 8865
rect -37820 8830 -37810 8865
rect -37775 8830 -37765 8865
rect -37730 8830 -37720 8865
rect -37685 8830 -37675 8865
rect -37640 8830 -37630 8865
rect -37595 8830 -37585 8865
rect -37550 8830 -37540 8865
rect -37505 8830 -37495 8865
rect -37460 8830 -37450 8865
rect -37415 8830 -37405 8865
rect -37370 8830 -37360 8865
rect -37325 8830 -37315 8865
rect -37280 8830 -37270 8865
rect -37235 8830 -37225 8865
rect -37190 8830 -37170 8865
rect -38770 8820 -37170 8830
rect -38770 8785 -38755 8820
rect -38720 8785 -38710 8820
rect -38675 8785 -38665 8820
rect -38630 8785 -38620 8820
rect -38585 8785 -38575 8820
rect -38540 8785 -38530 8820
rect -38495 8785 -38485 8820
rect -38450 8785 -38440 8820
rect -38405 8785 -38395 8820
rect -38360 8785 -38350 8820
rect -38315 8785 -38305 8820
rect -38270 8785 -38260 8820
rect -38225 8785 -38215 8820
rect -38180 8785 -38170 8820
rect -38135 8785 -38125 8820
rect -38090 8785 -38080 8820
rect -38045 8785 -38035 8820
rect -38000 8785 -37990 8820
rect -37955 8785 -37945 8820
rect -37910 8785 -37900 8820
rect -37865 8785 -37855 8820
rect -37820 8785 -37810 8820
rect -37775 8785 -37765 8820
rect -37730 8785 -37720 8820
rect -37685 8785 -37675 8820
rect -37640 8785 -37630 8820
rect -37595 8785 -37585 8820
rect -37550 8785 -37540 8820
rect -37505 8785 -37495 8820
rect -37460 8785 -37450 8820
rect -37415 8785 -37405 8820
rect -37370 8785 -37360 8820
rect -37325 8785 -37315 8820
rect -37280 8785 -37270 8820
rect -37235 8785 -37225 8820
rect -37190 8785 -37170 8820
rect -38770 8775 -37170 8785
rect -38770 8740 -38755 8775
rect -38720 8740 -38710 8775
rect -38675 8740 -38665 8775
rect -38630 8740 -38620 8775
rect -38585 8740 -38575 8775
rect -38540 8740 -38530 8775
rect -38495 8740 -38485 8775
rect -38450 8740 -38440 8775
rect -38405 8740 -38395 8775
rect -38360 8740 -38350 8775
rect -38315 8740 -38305 8775
rect -38270 8740 -38260 8775
rect -38225 8740 -38215 8775
rect -38180 8740 -38170 8775
rect -38135 8740 -38125 8775
rect -38090 8740 -38080 8775
rect -38045 8740 -38035 8775
rect -38000 8740 -37990 8775
rect -37955 8740 -37945 8775
rect -37910 8740 -37900 8775
rect -37865 8740 -37855 8775
rect -37820 8740 -37810 8775
rect -37775 8740 -37765 8775
rect -37730 8740 -37720 8775
rect -37685 8740 -37675 8775
rect -37640 8740 -37630 8775
rect -37595 8740 -37585 8775
rect -37550 8740 -37540 8775
rect -37505 8740 -37495 8775
rect -37460 8740 -37450 8775
rect -37415 8740 -37405 8775
rect -37370 8740 -37360 8775
rect -37325 8740 -37315 8775
rect -37280 8740 -37270 8775
rect -37235 8740 -37225 8775
rect -37190 8740 -37170 8775
rect -38770 8730 -37170 8740
rect -38770 8695 -38755 8730
rect -38720 8695 -38710 8730
rect -38675 8695 -38665 8730
rect -38630 8695 -38620 8730
rect -38585 8695 -38575 8730
rect -38540 8695 -38530 8730
rect -38495 8695 -38485 8730
rect -38450 8695 -38440 8730
rect -38405 8695 -38395 8730
rect -38360 8695 -38350 8730
rect -38315 8695 -38305 8730
rect -38270 8695 -38260 8730
rect -38225 8695 -38215 8730
rect -38180 8695 -38170 8730
rect -38135 8695 -38125 8730
rect -38090 8695 -38080 8730
rect -38045 8695 -38035 8730
rect -38000 8695 -37990 8730
rect -37955 8695 -37945 8730
rect -37910 8695 -37900 8730
rect -37865 8695 -37855 8730
rect -37820 8695 -37810 8730
rect -37775 8695 -37765 8730
rect -37730 8695 -37720 8730
rect -37685 8695 -37675 8730
rect -37640 8695 -37630 8730
rect -37595 8695 -37585 8730
rect -37550 8695 -37540 8730
rect -37505 8695 -37495 8730
rect -37460 8695 -37450 8730
rect -37415 8695 -37405 8730
rect -37370 8695 -37360 8730
rect -37325 8695 -37315 8730
rect -37280 8695 -37270 8730
rect -37235 8695 -37225 8730
rect -37190 8695 -37170 8730
rect -38770 8685 -37170 8695
rect -38770 8650 -38755 8685
rect -38720 8650 -38710 8685
rect -38675 8650 -38665 8685
rect -38630 8650 -38620 8685
rect -38585 8650 -38575 8685
rect -38540 8650 -38530 8685
rect -38495 8650 -38485 8685
rect -38450 8650 -38440 8685
rect -38405 8650 -38395 8685
rect -38360 8650 -38350 8685
rect -38315 8650 -38305 8685
rect -38270 8650 -38260 8685
rect -38225 8650 -38215 8685
rect -38180 8650 -38170 8685
rect -38135 8650 -38125 8685
rect -38090 8650 -38080 8685
rect -38045 8650 -38035 8685
rect -38000 8650 -37990 8685
rect -37955 8650 -37945 8685
rect -37910 8650 -37900 8685
rect -37865 8650 -37855 8685
rect -37820 8650 -37810 8685
rect -37775 8650 -37765 8685
rect -37730 8650 -37720 8685
rect -37685 8650 -37675 8685
rect -37640 8650 -37630 8685
rect -37595 8650 -37585 8685
rect -37550 8650 -37540 8685
rect -37505 8650 -37495 8685
rect -37460 8650 -37450 8685
rect -37415 8650 -37405 8685
rect -37370 8650 -37360 8685
rect -37325 8650 -37315 8685
rect -37280 8650 -37270 8685
rect -37235 8650 -37225 8685
rect -37190 8650 -37170 8685
rect -38770 8640 -37170 8650
rect -38770 8605 -38755 8640
rect -38720 8605 -38710 8640
rect -38675 8605 -38665 8640
rect -38630 8605 -38620 8640
rect -38585 8605 -38575 8640
rect -38540 8605 -38530 8640
rect -38495 8605 -38485 8640
rect -38450 8605 -38440 8640
rect -38405 8605 -38395 8640
rect -38360 8605 -38350 8640
rect -38315 8605 -38305 8640
rect -38270 8605 -38260 8640
rect -38225 8605 -38215 8640
rect -38180 8605 -38170 8640
rect -38135 8605 -38125 8640
rect -38090 8605 -38080 8640
rect -38045 8605 -38035 8640
rect -38000 8605 -37990 8640
rect -37955 8605 -37945 8640
rect -37910 8605 -37900 8640
rect -37865 8605 -37855 8640
rect -37820 8605 -37810 8640
rect -37775 8605 -37765 8640
rect -37730 8605 -37720 8640
rect -37685 8605 -37675 8640
rect -37640 8605 -37630 8640
rect -37595 8605 -37585 8640
rect -37550 8605 -37540 8640
rect -37505 8605 -37495 8640
rect -37460 8605 -37450 8640
rect -37415 8605 -37405 8640
rect -37370 8605 -37360 8640
rect -37325 8605 -37315 8640
rect -37280 8605 -37270 8640
rect -37235 8605 -37225 8640
rect -37190 8605 -37170 8640
rect -38770 8595 -37170 8605
rect -38770 8560 -38755 8595
rect -38720 8560 -38710 8595
rect -38675 8560 -38665 8595
rect -38630 8560 -38620 8595
rect -38585 8560 -38575 8595
rect -38540 8560 -38530 8595
rect -38495 8560 -38485 8595
rect -38450 8560 -38440 8595
rect -38405 8560 -38395 8595
rect -38360 8560 -38350 8595
rect -38315 8560 -38305 8595
rect -38270 8560 -38260 8595
rect -38225 8560 -38215 8595
rect -38180 8560 -38170 8595
rect -38135 8560 -38125 8595
rect -38090 8560 -38080 8595
rect -38045 8560 -38035 8595
rect -38000 8560 -37990 8595
rect -37955 8560 -37945 8595
rect -37910 8560 -37900 8595
rect -37865 8560 -37855 8595
rect -37820 8560 -37810 8595
rect -37775 8560 -37765 8595
rect -37730 8560 -37720 8595
rect -37685 8560 -37675 8595
rect -37640 8560 -37630 8595
rect -37595 8560 -37585 8595
rect -37550 8560 -37540 8595
rect -37505 8560 -37495 8595
rect -37460 8560 -37450 8595
rect -37415 8560 -37405 8595
rect -37370 8560 -37360 8595
rect -37325 8560 -37315 8595
rect -37280 8560 -37270 8595
rect -37235 8560 -37225 8595
rect -37190 8560 -37170 8595
rect -38770 8550 -37170 8560
rect -38770 8515 -38755 8550
rect -38720 8515 -38710 8550
rect -38675 8515 -38665 8550
rect -38630 8515 -38620 8550
rect -38585 8515 -38575 8550
rect -38540 8515 -38530 8550
rect -38495 8515 -38485 8550
rect -38450 8515 -38440 8550
rect -38405 8515 -38395 8550
rect -38360 8515 -38350 8550
rect -38315 8515 -38305 8550
rect -38270 8515 -38260 8550
rect -38225 8515 -38215 8550
rect -38180 8515 -38170 8550
rect -38135 8515 -38125 8550
rect -38090 8515 -38080 8550
rect -38045 8515 -38035 8550
rect -38000 8515 -37990 8550
rect -37955 8515 -37945 8550
rect -37910 8515 -37900 8550
rect -37865 8515 -37855 8550
rect -37820 8515 -37810 8550
rect -37775 8515 -37765 8550
rect -37730 8515 -37720 8550
rect -37685 8515 -37675 8550
rect -37640 8515 -37630 8550
rect -37595 8515 -37585 8550
rect -37550 8515 -37540 8550
rect -37505 8515 -37495 8550
rect -37460 8515 -37450 8550
rect -37415 8515 -37405 8550
rect -37370 8515 -37360 8550
rect -37325 8515 -37315 8550
rect -37280 8515 -37270 8550
rect -37235 8515 -37225 8550
rect -37190 8515 -37170 8550
rect -38770 8505 -37170 8515
rect -38770 8470 -38755 8505
rect -38720 8470 -38710 8505
rect -38675 8470 -38665 8505
rect -38630 8470 -38620 8505
rect -38585 8470 -38575 8505
rect -38540 8470 -38530 8505
rect -38495 8470 -38485 8505
rect -38450 8470 -38440 8505
rect -38405 8470 -38395 8505
rect -38360 8470 -38350 8505
rect -38315 8470 -38305 8505
rect -38270 8470 -38260 8505
rect -38225 8470 -38215 8505
rect -38180 8470 -38170 8505
rect -38135 8470 -38125 8505
rect -38090 8470 -38080 8505
rect -38045 8470 -38035 8505
rect -38000 8470 -37990 8505
rect -37955 8470 -37945 8505
rect -37910 8470 -37900 8505
rect -37865 8470 -37855 8505
rect -37820 8470 -37810 8505
rect -37775 8470 -37765 8505
rect -37730 8470 -37720 8505
rect -37685 8470 -37675 8505
rect -37640 8470 -37630 8505
rect -37595 8470 -37585 8505
rect -37550 8470 -37540 8505
rect -37505 8470 -37495 8505
rect -37460 8470 -37450 8505
rect -37415 8470 -37405 8505
rect -37370 8470 -37360 8505
rect -37325 8470 -37315 8505
rect -37280 8470 -37270 8505
rect -37235 8470 -37225 8505
rect -37190 8470 -37170 8505
rect -38770 8460 -37170 8470
rect -38770 8425 -38755 8460
rect -38720 8425 -38710 8460
rect -38675 8425 -38665 8460
rect -38630 8425 -38620 8460
rect -38585 8425 -38575 8460
rect -38540 8425 -38530 8460
rect -38495 8425 -38485 8460
rect -38450 8425 -38440 8460
rect -38405 8425 -38395 8460
rect -38360 8425 -38350 8460
rect -38315 8425 -38305 8460
rect -38270 8425 -38260 8460
rect -38225 8425 -38215 8460
rect -38180 8425 -38170 8460
rect -38135 8425 -38125 8460
rect -38090 8425 -38080 8460
rect -38045 8425 -38035 8460
rect -38000 8425 -37990 8460
rect -37955 8425 -37945 8460
rect -37910 8425 -37900 8460
rect -37865 8425 -37855 8460
rect -37820 8425 -37810 8460
rect -37775 8425 -37765 8460
rect -37730 8425 -37720 8460
rect -37685 8425 -37675 8460
rect -37640 8425 -37630 8460
rect -37595 8425 -37585 8460
rect -37550 8425 -37540 8460
rect -37505 8425 -37495 8460
rect -37460 8425 -37450 8460
rect -37415 8425 -37405 8460
rect -37370 8425 -37360 8460
rect -37325 8425 -37315 8460
rect -37280 8425 -37270 8460
rect -37235 8425 -37225 8460
rect -37190 8425 -37170 8460
rect -38770 8415 -37170 8425
rect -38770 8380 -38755 8415
rect -38720 8380 -38710 8415
rect -38675 8380 -38665 8415
rect -38630 8380 -38620 8415
rect -38585 8380 -38575 8415
rect -38540 8380 -38530 8415
rect -38495 8380 -38485 8415
rect -38450 8380 -38440 8415
rect -38405 8380 -38395 8415
rect -38360 8380 -38350 8415
rect -38315 8380 -38305 8415
rect -38270 8380 -38260 8415
rect -38225 8380 -38215 8415
rect -38180 8380 -38170 8415
rect -38135 8380 -38125 8415
rect -38090 8380 -38080 8415
rect -38045 8380 -38035 8415
rect -38000 8380 -37990 8415
rect -37955 8380 -37945 8415
rect -37910 8380 -37900 8415
rect -37865 8380 -37855 8415
rect -37820 8380 -37810 8415
rect -37775 8380 -37765 8415
rect -37730 8380 -37720 8415
rect -37685 8380 -37675 8415
rect -37640 8380 -37630 8415
rect -37595 8380 -37585 8415
rect -37550 8380 -37540 8415
rect -37505 8380 -37495 8415
rect -37460 8380 -37450 8415
rect -37415 8380 -37405 8415
rect -37370 8380 -37360 8415
rect -37325 8380 -37315 8415
rect -37280 8380 -37270 8415
rect -37235 8380 -37225 8415
rect -37190 8380 -37170 8415
rect -38770 8370 -37170 8380
rect -38770 8335 -38755 8370
rect -38720 8335 -38710 8370
rect -38675 8335 -38665 8370
rect -38630 8335 -38620 8370
rect -38585 8335 -38575 8370
rect -38540 8335 -38530 8370
rect -38495 8335 -38485 8370
rect -38450 8335 -38440 8370
rect -38405 8335 -38395 8370
rect -38360 8335 -38350 8370
rect -38315 8335 -38305 8370
rect -38270 8335 -38260 8370
rect -38225 8335 -38215 8370
rect -38180 8335 -38170 8370
rect -38135 8335 -38125 8370
rect -38090 8335 -38080 8370
rect -38045 8335 -38035 8370
rect -38000 8335 -37990 8370
rect -37955 8335 -37945 8370
rect -37910 8335 -37900 8370
rect -37865 8335 -37855 8370
rect -37820 8335 -37810 8370
rect -37775 8335 -37765 8370
rect -37730 8335 -37720 8370
rect -37685 8335 -37675 8370
rect -37640 8335 -37630 8370
rect -37595 8335 -37585 8370
rect -37550 8335 -37540 8370
rect -37505 8335 -37495 8370
rect -37460 8335 -37450 8370
rect -37415 8335 -37405 8370
rect -37370 8335 -37360 8370
rect -37325 8335 -37315 8370
rect -37280 8335 -37270 8370
rect -37235 8335 -37225 8370
rect -37190 8335 -37170 8370
rect -38770 8325 -37170 8335
rect -38770 8290 -38755 8325
rect -38720 8290 -38710 8325
rect -38675 8290 -38665 8325
rect -38630 8290 -38620 8325
rect -38585 8290 -38575 8325
rect -38540 8290 -38530 8325
rect -38495 8290 -38485 8325
rect -38450 8290 -38440 8325
rect -38405 8290 -38395 8325
rect -38360 8290 -38350 8325
rect -38315 8290 -38305 8325
rect -38270 8290 -38260 8325
rect -38225 8290 -38215 8325
rect -38180 8290 -38170 8325
rect -38135 8290 -38125 8325
rect -38090 8290 -38080 8325
rect -38045 8290 -38035 8325
rect -38000 8290 -37990 8325
rect -37955 8290 -37945 8325
rect -37910 8290 -37900 8325
rect -37865 8290 -37855 8325
rect -37820 8290 -37810 8325
rect -37775 8290 -37765 8325
rect -37730 8290 -37720 8325
rect -37685 8290 -37675 8325
rect -37640 8290 -37630 8325
rect -37595 8290 -37585 8325
rect -37550 8290 -37540 8325
rect -37505 8290 -37495 8325
rect -37460 8290 -37450 8325
rect -37415 8290 -37405 8325
rect -37370 8290 -37360 8325
rect -37325 8290 -37315 8325
rect -37280 8290 -37270 8325
rect -37235 8290 -37225 8325
rect -37190 8290 -37170 8325
rect -38770 8280 -37170 8290
rect -38770 8245 -38755 8280
rect -38720 8245 -38710 8280
rect -38675 8245 -38665 8280
rect -38630 8245 -38620 8280
rect -38585 8245 -38575 8280
rect -38540 8245 -38530 8280
rect -38495 8245 -38485 8280
rect -38450 8245 -38440 8280
rect -38405 8245 -38395 8280
rect -38360 8245 -38350 8280
rect -38315 8245 -38305 8280
rect -38270 8245 -38260 8280
rect -38225 8245 -38215 8280
rect -38180 8245 -38170 8280
rect -38135 8245 -38125 8280
rect -38090 8245 -38080 8280
rect -38045 8245 -38035 8280
rect -38000 8245 -37990 8280
rect -37955 8245 -37945 8280
rect -37910 8245 -37900 8280
rect -37865 8245 -37855 8280
rect -37820 8245 -37810 8280
rect -37775 8245 -37765 8280
rect -37730 8245 -37720 8280
rect -37685 8245 -37675 8280
rect -37640 8245 -37630 8280
rect -37595 8245 -37585 8280
rect -37550 8245 -37540 8280
rect -37505 8245 -37495 8280
rect -37460 8245 -37450 8280
rect -37415 8245 -37405 8280
rect -37370 8245 -37360 8280
rect -37325 8245 -37315 8280
rect -37280 8245 -37270 8280
rect -37235 8245 -37225 8280
rect -37190 8245 -37170 8280
rect -38770 8235 -37170 8245
rect -38770 8200 -38755 8235
rect -38720 8200 -38710 8235
rect -38675 8200 -38665 8235
rect -38630 8200 -38620 8235
rect -38585 8200 -38575 8235
rect -38540 8200 -38530 8235
rect -38495 8200 -38485 8235
rect -38450 8200 -38440 8235
rect -38405 8200 -38395 8235
rect -38360 8200 -38350 8235
rect -38315 8200 -38305 8235
rect -38270 8200 -38260 8235
rect -38225 8200 -38215 8235
rect -38180 8200 -38170 8235
rect -38135 8200 -38125 8235
rect -38090 8200 -38080 8235
rect -38045 8200 -38035 8235
rect -38000 8200 -37990 8235
rect -37955 8200 -37945 8235
rect -37910 8200 -37900 8235
rect -37865 8200 -37855 8235
rect -37820 8200 -37810 8235
rect -37775 8200 -37765 8235
rect -37730 8200 -37720 8235
rect -37685 8200 -37675 8235
rect -37640 8200 -37630 8235
rect -37595 8200 -37585 8235
rect -37550 8200 -37540 8235
rect -37505 8200 -37495 8235
rect -37460 8200 -37450 8235
rect -37415 8200 -37405 8235
rect -37370 8200 -37360 8235
rect -37325 8200 -37315 8235
rect -37280 8200 -37270 8235
rect -37235 8200 -37225 8235
rect -37190 8200 -37170 8235
rect -38770 8190 -37170 8200
rect -38770 8155 -38755 8190
rect -38720 8155 -38710 8190
rect -38675 8155 -38665 8190
rect -38630 8155 -38620 8190
rect -38585 8155 -38575 8190
rect -38540 8155 -38530 8190
rect -38495 8155 -38485 8190
rect -38450 8155 -38440 8190
rect -38405 8155 -38395 8190
rect -38360 8155 -38350 8190
rect -38315 8155 -38305 8190
rect -38270 8155 -38260 8190
rect -38225 8155 -38215 8190
rect -38180 8155 -38170 8190
rect -38135 8155 -38125 8190
rect -38090 8155 -38080 8190
rect -38045 8155 -38035 8190
rect -38000 8155 -37990 8190
rect -37955 8155 -37945 8190
rect -37910 8155 -37900 8190
rect -37865 8155 -37855 8190
rect -37820 8155 -37810 8190
rect -37775 8155 -37765 8190
rect -37730 8155 -37720 8190
rect -37685 8155 -37675 8190
rect -37640 8155 -37630 8190
rect -37595 8155 -37585 8190
rect -37550 8155 -37540 8190
rect -37505 8155 -37495 8190
rect -37460 8155 -37450 8190
rect -37415 8155 -37405 8190
rect -37370 8155 -37360 8190
rect -37325 8155 -37315 8190
rect -37280 8155 -37270 8190
rect -37235 8155 -37225 8190
rect -37190 8155 -37170 8190
rect -38770 8145 -37170 8155
rect -38770 8110 -38755 8145
rect -38720 8110 -38710 8145
rect -38675 8110 -38665 8145
rect -38630 8110 -38620 8145
rect -38585 8110 -38575 8145
rect -38540 8110 -38530 8145
rect -38495 8110 -38485 8145
rect -38450 8110 -38440 8145
rect -38405 8110 -38395 8145
rect -38360 8110 -38350 8145
rect -38315 8110 -38305 8145
rect -38270 8110 -38260 8145
rect -38225 8110 -38215 8145
rect -38180 8110 -38170 8145
rect -38135 8110 -38125 8145
rect -38090 8110 -38080 8145
rect -38045 8110 -38035 8145
rect -38000 8110 -37990 8145
rect -37955 8110 -37945 8145
rect -37910 8110 -37900 8145
rect -37865 8110 -37855 8145
rect -37820 8110 -37810 8145
rect -37775 8110 -37765 8145
rect -37730 8110 -37720 8145
rect -37685 8110 -37675 8145
rect -37640 8110 -37630 8145
rect -37595 8110 -37585 8145
rect -37550 8110 -37540 8145
rect -37505 8110 -37495 8145
rect -37460 8110 -37450 8145
rect -37415 8110 -37405 8145
rect -37370 8110 -37360 8145
rect -37325 8110 -37315 8145
rect -37280 8110 -37270 8145
rect -37235 8110 -37225 8145
rect -37190 8110 -37170 8145
rect -38770 8100 -37170 8110
rect -38770 8065 -38755 8100
rect -38720 8065 -38710 8100
rect -38675 8065 -38665 8100
rect -38630 8065 -38620 8100
rect -38585 8065 -38575 8100
rect -38540 8065 -38530 8100
rect -38495 8065 -38485 8100
rect -38450 8065 -38440 8100
rect -38405 8065 -38395 8100
rect -38360 8065 -38350 8100
rect -38315 8065 -38305 8100
rect -38270 8065 -38260 8100
rect -38225 8065 -38215 8100
rect -38180 8065 -38170 8100
rect -38135 8065 -38125 8100
rect -38090 8065 -38080 8100
rect -38045 8065 -38035 8100
rect -38000 8065 -37990 8100
rect -37955 8065 -37945 8100
rect -37910 8065 -37900 8100
rect -37865 8065 -37855 8100
rect -37820 8065 -37810 8100
rect -37775 8065 -37765 8100
rect -37730 8065 -37720 8100
rect -37685 8065 -37675 8100
rect -37640 8065 -37630 8100
rect -37595 8065 -37585 8100
rect -37550 8065 -37540 8100
rect -37505 8065 -37495 8100
rect -37460 8065 -37450 8100
rect -37415 8065 -37405 8100
rect -37370 8065 -37360 8100
rect -37325 8065 -37315 8100
rect -37280 8065 -37270 8100
rect -37235 8065 -37225 8100
rect -37190 8065 -37170 8100
rect -38770 8030 -37170 8065
rect -38770 7995 -38755 8030
rect -38720 7995 -38710 8030
rect -38675 7995 -38665 8030
rect -38630 7995 -38620 8030
rect -38585 7995 -38575 8030
rect -38540 7995 -38530 8030
rect -38495 7995 -38485 8030
rect -38450 7995 -38440 8030
rect -38405 7995 -38395 8030
rect -38360 7995 -38350 8030
rect -38315 7995 -38305 8030
rect -38270 7995 -38260 8030
rect -38225 7995 -38215 8030
rect -38180 7995 -38170 8030
rect -38135 7995 -38125 8030
rect -38090 7995 -38080 8030
rect -38045 7995 -38035 8030
rect -38000 7995 -37990 8030
rect -37955 7995 -37945 8030
rect -37910 7995 -37900 8030
rect -37865 7995 -37855 8030
rect -37820 7995 -37810 8030
rect -37775 7995 -37765 8030
rect -37730 7995 -37720 8030
rect -37685 7995 -37675 8030
rect -37640 7995 -37630 8030
rect -37595 7995 -37585 8030
rect -37550 7995 -37540 8030
rect -37505 7995 -37495 8030
rect -37460 7995 -37450 8030
rect -37415 7995 -37405 8030
rect -37370 7995 -37360 8030
rect -37325 7995 -37315 8030
rect -37280 7995 -37270 8030
rect -37235 7995 -37225 8030
rect -37190 7995 -37170 8030
rect -38770 7985 -37170 7995
rect -38770 7950 -38755 7985
rect -38720 7950 -38710 7985
rect -38675 7950 -38665 7985
rect -38630 7950 -38620 7985
rect -38585 7950 -38575 7985
rect -38540 7950 -38530 7985
rect -38495 7950 -38485 7985
rect -38450 7950 -38440 7985
rect -38405 7950 -38395 7985
rect -38360 7950 -38350 7985
rect -38315 7950 -38305 7985
rect -38270 7950 -38260 7985
rect -38225 7950 -38215 7985
rect -38180 7950 -38170 7985
rect -38135 7950 -38125 7985
rect -38090 7950 -38080 7985
rect -38045 7950 -38035 7985
rect -38000 7950 -37990 7985
rect -37955 7950 -37945 7985
rect -37910 7950 -37900 7985
rect -37865 7950 -37855 7985
rect -37820 7950 -37810 7985
rect -37775 7950 -37765 7985
rect -37730 7950 -37720 7985
rect -37685 7950 -37675 7985
rect -37640 7950 -37630 7985
rect -37595 7950 -37585 7985
rect -37550 7950 -37540 7985
rect -37505 7950 -37495 7985
rect -37460 7950 -37450 7985
rect -37415 7950 -37405 7985
rect -37370 7950 -37360 7985
rect -37325 7950 -37315 7985
rect -37280 7950 -37270 7985
rect -37235 7950 -37225 7985
rect -37190 7950 -37170 7985
rect -38770 7940 -37170 7950
rect -38770 7905 -38755 7940
rect -38720 7905 -38710 7940
rect -38675 7905 -38665 7940
rect -38630 7905 -38620 7940
rect -38585 7905 -38575 7940
rect -38540 7905 -38530 7940
rect -38495 7905 -38485 7940
rect -38450 7905 -38440 7940
rect -38405 7905 -38395 7940
rect -38360 7905 -38350 7940
rect -38315 7905 -38305 7940
rect -38270 7905 -38260 7940
rect -38225 7905 -38215 7940
rect -38180 7905 -38170 7940
rect -38135 7905 -38125 7940
rect -38090 7905 -38080 7940
rect -38045 7905 -38035 7940
rect -38000 7905 -37990 7940
rect -37955 7905 -37945 7940
rect -37910 7905 -37900 7940
rect -37865 7905 -37855 7940
rect -37820 7905 -37810 7940
rect -37775 7905 -37765 7940
rect -37730 7905 -37720 7940
rect -37685 7905 -37675 7940
rect -37640 7905 -37630 7940
rect -37595 7905 -37585 7940
rect -37550 7905 -37540 7940
rect -37505 7905 -37495 7940
rect -37460 7905 -37450 7940
rect -37415 7905 -37405 7940
rect -37370 7905 -37360 7940
rect -37325 7905 -37315 7940
rect -37280 7905 -37270 7940
rect -37235 7905 -37225 7940
rect -37190 7905 -37170 7940
rect -38770 7895 -37170 7905
rect -38770 7860 -38755 7895
rect -38720 7860 -38710 7895
rect -38675 7860 -38665 7895
rect -38630 7860 -38620 7895
rect -38585 7860 -38575 7895
rect -38540 7860 -38530 7895
rect -38495 7860 -38485 7895
rect -38450 7860 -38440 7895
rect -38405 7860 -38395 7895
rect -38360 7860 -38350 7895
rect -38315 7860 -38305 7895
rect -38270 7860 -38260 7895
rect -38225 7860 -38215 7895
rect -38180 7860 -38170 7895
rect -38135 7860 -38125 7895
rect -38090 7860 -38080 7895
rect -38045 7860 -38035 7895
rect -38000 7860 -37990 7895
rect -37955 7860 -37945 7895
rect -37910 7860 -37900 7895
rect -37865 7860 -37855 7895
rect -37820 7860 -37810 7895
rect -37775 7860 -37765 7895
rect -37730 7860 -37720 7895
rect -37685 7860 -37675 7895
rect -37640 7860 -37630 7895
rect -37595 7860 -37585 7895
rect -37550 7860 -37540 7895
rect -37505 7860 -37495 7895
rect -37460 7860 -37450 7895
rect -37415 7860 -37405 7895
rect -37370 7860 -37360 7895
rect -37325 7860 -37315 7895
rect -37280 7860 -37270 7895
rect -37235 7860 -37225 7895
rect -37190 7860 -37170 7895
rect -38770 7850 -37170 7860
rect -38770 7815 -38755 7850
rect -38720 7815 -38710 7850
rect -38675 7815 -38665 7850
rect -38630 7815 -38620 7850
rect -38585 7815 -38575 7850
rect -38540 7815 -38530 7850
rect -38495 7815 -38485 7850
rect -38450 7815 -38440 7850
rect -38405 7815 -38395 7850
rect -38360 7815 -38350 7850
rect -38315 7815 -38305 7850
rect -38270 7815 -38260 7850
rect -38225 7815 -38215 7850
rect -38180 7815 -38170 7850
rect -38135 7815 -38125 7850
rect -38090 7815 -38080 7850
rect -38045 7815 -38035 7850
rect -38000 7815 -37990 7850
rect -37955 7815 -37945 7850
rect -37910 7815 -37900 7850
rect -37865 7815 -37855 7850
rect -37820 7815 -37810 7850
rect -37775 7815 -37765 7850
rect -37730 7815 -37720 7850
rect -37685 7815 -37675 7850
rect -37640 7815 -37630 7850
rect -37595 7815 -37585 7850
rect -37550 7815 -37540 7850
rect -37505 7815 -37495 7850
rect -37460 7815 -37450 7850
rect -37415 7815 -37405 7850
rect -37370 7815 -37360 7850
rect -37325 7815 -37315 7850
rect -37280 7815 -37270 7850
rect -37235 7815 -37225 7850
rect -37190 7815 -37170 7850
rect -38770 7805 -37170 7815
rect -38770 7770 -38755 7805
rect -38720 7770 -38710 7805
rect -38675 7770 -38665 7805
rect -38630 7770 -38620 7805
rect -38585 7770 -38575 7805
rect -38540 7770 -38530 7805
rect -38495 7770 -38485 7805
rect -38450 7770 -38440 7805
rect -38405 7770 -38395 7805
rect -38360 7770 -38350 7805
rect -38315 7770 -38305 7805
rect -38270 7770 -38260 7805
rect -38225 7770 -38215 7805
rect -38180 7770 -38170 7805
rect -38135 7770 -38125 7805
rect -38090 7770 -38080 7805
rect -38045 7770 -38035 7805
rect -38000 7770 -37990 7805
rect -37955 7770 -37945 7805
rect -37910 7770 -37900 7805
rect -37865 7770 -37855 7805
rect -37820 7770 -37810 7805
rect -37775 7770 -37765 7805
rect -37730 7770 -37720 7805
rect -37685 7770 -37675 7805
rect -37640 7770 -37630 7805
rect -37595 7770 -37585 7805
rect -37550 7770 -37540 7805
rect -37505 7770 -37495 7805
rect -37460 7770 -37450 7805
rect -37415 7770 -37405 7805
rect -37370 7770 -37360 7805
rect -37325 7770 -37315 7805
rect -37280 7770 -37270 7805
rect -37235 7770 -37225 7805
rect -37190 7770 -37170 7805
rect -38770 7760 -37170 7770
rect -38770 7725 -38755 7760
rect -38720 7725 -38710 7760
rect -38675 7725 -38665 7760
rect -38630 7725 -38620 7760
rect -38585 7725 -38575 7760
rect -38540 7725 -38530 7760
rect -38495 7725 -38485 7760
rect -38450 7725 -38440 7760
rect -38405 7725 -38395 7760
rect -38360 7725 -38350 7760
rect -38315 7725 -38305 7760
rect -38270 7725 -38260 7760
rect -38225 7725 -38215 7760
rect -38180 7725 -38170 7760
rect -38135 7725 -38125 7760
rect -38090 7725 -38080 7760
rect -38045 7725 -38035 7760
rect -38000 7725 -37990 7760
rect -37955 7725 -37945 7760
rect -37910 7725 -37900 7760
rect -37865 7725 -37855 7760
rect -37820 7725 -37810 7760
rect -37775 7725 -37765 7760
rect -37730 7725 -37720 7760
rect -37685 7725 -37675 7760
rect -37640 7725 -37630 7760
rect -37595 7725 -37585 7760
rect -37550 7725 -37540 7760
rect -37505 7725 -37495 7760
rect -37460 7725 -37450 7760
rect -37415 7725 -37405 7760
rect -37370 7725 -37360 7760
rect -37325 7725 -37315 7760
rect -37280 7725 -37270 7760
rect -37235 7725 -37225 7760
rect -37190 7725 -37170 7760
rect -38770 7715 -37170 7725
rect -38770 7680 -38755 7715
rect -38720 7680 -38710 7715
rect -38675 7680 -38665 7715
rect -38630 7680 -38620 7715
rect -38585 7680 -38575 7715
rect -38540 7680 -38530 7715
rect -38495 7680 -38485 7715
rect -38450 7680 -38440 7715
rect -38405 7680 -38395 7715
rect -38360 7680 -38350 7715
rect -38315 7680 -38305 7715
rect -38270 7680 -38260 7715
rect -38225 7680 -38215 7715
rect -38180 7680 -38170 7715
rect -38135 7680 -38125 7715
rect -38090 7680 -38080 7715
rect -38045 7680 -38035 7715
rect -38000 7680 -37990 7715
rect -37955 7680 -37945 7715
rect -37910 7680 -37900 7715
rect -37865 7680 -37855 7715
rect -37820 7680 -37810 7715
rect -37775 7680 -37765 7715
rect -37730 7680 -37720 7715
rect -37685 7680 -37675 7715
rect -37640 7680 -37630 7715
rect -37595 7680 -37585 7715
rect -37550 7680 -37540 7715
rect -37505 7680 -37495 7715
rect -37460 7680 -37450 7715
rect -37415 7680 -37405 7715
rect -37370 7680 -37360 7715
rect -37325 7680 -37315 7715
rect -37280 7680 -37270 7715
rect -37235 7680 -37225 7715
rect -37190 7680 -37170 7715
rect -38770 7670 -37170 7680
rect -38770 7635 -38755 7670
rect -38720 7635 -38710 7670
rect -38675 7635 -38665 7670
rect -38630 7635 -38620 7670
rect -38585 7635 -38575 7670
rect -38540 7635 -38530 7670
rect -38495 7635 -38485 7670
rect -38450 7635 -38440 7670
rect -38405 7635 -38395 7670
rect -38360 7635 -38350 7670
rect -38315 7635 -38305 7670
rect -38270 7635 -38260 7670
rect -38225 7635 -38215 7670
rect -38180 7635 -38170 7670
rect -38135 7635 -38125 7670
rect -38090 7635 -38080 7670
rect -38045 7635 -38035 7670
rect -38000 7635 -37990 7670
rect -37955 7635 -37945 7670
rect -37910 7635 -37900 7670
rect -37865 7635 -37855 7670
rect -37820 7635 -37810 7670
rect -37775 7635 -37765 7670
rect -37730 7635 -37720 7670
rect -37685 7635 -37675 7670
rect -37640 7635 -37630 7670
rect -37595 7635 -37585 7670
rect -37550 7635 -37540 7670
rect -37505 7635 -37495 7670
rect -37460 7635 -37450 7670
rect -37415 7635 -37405 7670
rect -37370 7635 -37360 7670
rect -37325 7635 -37315 7670
rect -37280 7635 -37270 7670
rect -37235 7635 -37225 7670
rect -37190 7635 -37170 7670
rect -38770 7625 -37170 7635
rect -38770 7590 -38755 7625
rect -38720 7590 -38710 7625
rect -38675 7590 -38665 7625
rect -38630 7590 -38620 7625
rect -38585 7590 -38575 7625
rect -38540 7590 -38530 7625
rect -38495 7590 -38485 7625
rect -38450 7590 -38440 7625
rect -38405 7590 -38395 7625
rect -38360 7590 -38350 7625
rect -38315 7590 -38305 7625
rect -38270 7590 -38260 7625
rect -38225 7590 -38215 7625
rect -38180 7590 -38170 7625
rect -38135 7590 -38125 7625
rect -38090 7590 -38080 7625
rect -38045 7590 -38035 7625
rect -38000 7590 -37990 7625
rect -37955 7590 -37945 7625
rect -37910 7590 -37900 7625
rect -37865 7590 -37855 7625
rect -37820 7590 -37810 7625
rect -37775 7590 -37765 7625
rect -37730 7590 -37720 7625
rect -37685 7590 -37675 7625
rect -37640 7590 -37630 7625
rect -37595 7590 -37585 7625
rect -37550 7590 -37540 7625
rect -37505 7590 -37495 7625
rect -37460 7590 -37450 7625
rect -37415 7590 -37405 7625
rect -37370 7590 -37360 7625
rect -37325 7590 -37315 7625
rect -37280 7590 -37270 7625
rect -37235 7590 -37225 7625
rect -37190 7590 -37170 7625
rect -38770 7580 -37170 7590
rect -38770 7545 -38755 7580
rect -38720 7545 -38710 7580
rect -38675 7545 -38665 7580
rect -38630 7545 -38620 7580
rect -38585 7545 -38575 7580
rect -38540 7545 -38530 7580
rect -38495 7545 -38485 7580
rect -38450 7545 -38440 7580
rect -38405 7545 -38395 7580
rect -38360 7545 -38350 7580
rect -38315 7545 -38305 7580
rect -38270 7545 -38260 7580
rect -38225 7545 -38215 7580
rect -38180 7545 -38170 7580
rect -38135 7545 -38125 7580
rect -38090 7545 -38080 7580
rect -38045 7545 -38035 7580
rect -38000 7545 -37990 7580
rect -37955 7545 -37945 7580
rect -37910 7545 -37900 7580
rect -37865 7545 -37855 7580
rect -37820 7545 -37810 7580
rect -37775 7545 -37765 7580
rect -37730 7545 -37720 7580
rect -37685 7545 -37675 7580
rect -37640 7545 -37630 7580
rect -37595 7545 -37585 7580
rect -37550 7545 -37540 7580
rect -37505 7545 -37495 7580
rect -37460 7545 -37450 7580
rect -37415 7545 -37405 7580
rect -37370 7545 -37360 7580
rect -37325 7545 -37315 7580
rect -37280 7545 -37270 7580
rect -37235 7545 -37225 7580
rect -37190 7545 -37170 7580
rect -38770 7535 -37170 7545
rect -38770 7500 -38755 7535
rect -38720 7500 -38710 7535
rect -38675 7500 -38665 7535
rect -38630 7500 -38620 7535
rect -38585 7500 -38575 7535
rect -38540 7500 -38530 7535
rect -38495 7500 -38485 7535
rect -38450 7500 -38440 7535
rect -38405 7500 -38395 7535
rect -38360 7500 -38350 7535
rect -38315 7500 -38305 7535
rect -38270 7500 -38260 7535
rect -38225 7500 -38215 7535
rect -38180 7500 -38170 7535
rect -38135 7500 -38125 7535
rect -38090 7500 -38080 7535
rect -38045 7500 -38035 7535
rect -38000 7500 -37990 7535
rect -37955 7500 -37945 7535
rect -37910 7500 -37900 7535
rect -37865 7500 -37855 7535
rect -37820 7500 -37810 7535
rect -37775 7500 -37765 7535
rect -37730 7500 -37720 7535
rect -37685 7500 -37675 7535
rect -37640 7500 -37630 7535
rect -37595 7500 -37585 7535
rect -37550 7500 -37540 7535
rect -37505 7500 -37495 7535
rect -37460 7500 -37450 7535
rect -37415 7500 -37405 7535
rect -37370 7500 -37360 7535
rect -37325 7500 -37315 7535
rect -37280 7500 -37270 7535
rect -37235 7500 -37225 7535
rect -37190 7500 -37170 7535
rect -38770 7490 -37170 7500
rect -38770 7455 -38755 7490
rect -38720 7455 -38710 7490
rect -38675 7455 -38665 7490
rect -38630 7455 -38620 7490
rect -38585 7455 -38575 7490
rect -38540 7455 -38530 7490
rect -38495 7455 -38485 7490
rect -38450 7455 -38440 7490
rect -38405 7455 -38395 7490
rect -38360 7455 -38350 7490
rect -38315 7455 -38305 7490
rect -38270 7455 -38260 7490
rect -38225 7455 -38215 7490
rect -38180 7455 -38170 7490
rect -38135 7455 -38125 7490
rect -38090 7455 -38080 7490
rect -38045 7455 -38035 7490
rect -38000 7455 -37990 7490
rect -37955 7455 -37945 7490
rect -37910 7455 -37900 7490
rect -37865 7455 -37855 7490
rect -37820 7455 -37810 7490
rect -37775 7455 -37765 7490
rect -37730 7455 -37720 7490
rect -37685 7455 -37675 7490
rect -37640 7455 -37630 7490
rect -37595 7455 -37585 7490
rect -37550 7455 -37540 7490
rect -37505 7455 -37495 7490
rect -37460 7455 -37450 7490
rect -37415 7455 -37405 7490
rect -37370 7455 -37360 7490
rect -37325 7455 -37315 7490
rect -37280 7455 -37270 7490
rect -37235 7455 -37225 7490
rect -37190 7455 -37170 7490
rect -38770 7445 -37170 7455
rect -38770 7410 -38755 7445
rect -38720 7410 -38710 7445
rect -38675 7410 -38665 7445
rect -38630 7410 -38620 7445
rect -38585 7410 -38575 7445
rect -38540 7410 -38530 7445
rect -38495 7410 -38485 7445
rect -38450 7410 -38440 7445
rect -38405 7410 -38395 7445
rect -38360 7410 -38350 7445
rect -38315 7410 -38305 7445
rect -38270 7410 -38260 7445
rect -38225 7410 -38215 7445
rect -38180 7410 -38170 7445
rect -38135 7410 -38125 7445
rect -38090 7410 -38080 7445
rect -38045 7410 -38035 7445
rect -38000 7410 -37990 7445
rect -37955 7410 -37945 7445
rect -37910 7410 -37900 7445
rect -37865 7410 -37855 7445
rect -37820 7410 -37810 7445
rect -37775 7410 -37765 7445
rect -37730 7410 -37720 7445
rect -37685 7410 -37675 7445
rect -37640 7410 -37630 7445
rect -37595 7410 -37585 7445
rect -37550 7410 -37540 7445
rect -37505 7410 -37495 7445
rect -37460 7410 -37450 7445
rect -37415 7410 -37405 7445
rect -37370 7410 -37360 7445
rect -37325 7410 -37315 7445
rect -37280 7410 -37270 7445
rect -37235 7410 -37225 7445
rect -37190 7410 -37170 7445
rect -38770 7400 -37170 7410
rect -38770 7365 -38755 7400
rect -38720 7365 -38710 7400
rect -38675 7365 -38665 7400
rect -38630 7365 -38620 7400
rect -38585 7365 -38575 7400
rect -38540 7365 -38530 7400
rect -38495 7365 -38485 7400
rect -38450 7365 -38440 7400
rect -38405 7365 -38395 7400
rect -38360 7365 -38350 7400
rect -38315 7365 -38305 7400
rect -38270 7365 -38260 7400
rect -38225 7365 -38215 7400
rect -38180 7365 -38170 7400
rect -38135 7365 -38125 7400
rect -38090 7365 -38080 7400
rect -38045 7365 -38035 7400
rect -38000 7365 -37990 7400
rect -37955 7365 -37945 7400
rect -37910 7365 -37900 7400
rect -37865 7365 -37855 7400
rect -37820 7365 -37810 7400
rect -37775 7365 -37765 7400
rect -37730 7365 -37720 7400
rect -37685 7365 -37675 7400
rect -37640 7365 -37630 7400
rect -37595 7365 -37585 7400
rect -37550 7365 -37540 7400
rect -37505 7365 -37495 7400
rect -37460 7365 -37450 7400
rect -37415 7365 -37405 7400
rect -37370 7365 -37360 7400
rect -37325 7365 -37315 7400
rect -37280 7365 -37270 7400
rect -37235 7365 -37225 7400
rect -37190 7365 -37170 7400
rect -38770 7355 -37170 7365
rect -38770 7320 -38755 7355
rect -38720 7320 -38710 7355
rect -38675 7320 -38665 7355
rect -38630 7320 -38620 7355
rect -38585 7320 -38575 7355
rect -38540 7320 -38530 7355
rect -38495 7320 -38485 7355
rect -38450 7320 -38440 7355
rect -38405 7320 -38395 7355
rect -38360 7320 -38350 7355
rect -38315 7320 -38305 7355
rect -38270 7320 -38260 7355
rect -38225 7320 -38215 7355
rect -38180 7320 -38170 7355
rect -38135 7320 -38125 7355
rect -38090 7320 -38080 7355
rect -38045 7320 -38035 7355
rect -38000 7320 -37990 7355
rect -37955 7320 -37945 7355
rect -37910 7320 -37900 7355
rect -37865 7320 -37855 7355
rect -37820 7320 -37810 7355
rect -37775 7320 -37765 7355
rect -37730 7320 -37720 7355
rect -37685 7320 -37675 7355
rect -37640 7320 -37630 7355
rect -37595 7320 -37585 7355
rect -37550 7320 -37540 7355
rect -37505 7320 -37495 7355
rect -37460 7320 -37450 7355
rect -37415 7320 -37405 7355
rect -37370 7320 -37360 7355
rect -37325 7320 -37315 7355
rect -37280 7320 -37270 7355
rect -37235 7320 -37225 7355
rect -37190 7320 -37170 7355
rect -38770 7310 -37170 7320
rect -38770 7275 -38755 7310
rect -38720 7275 -38710 7310
rect -38675 7275 -38665 7310
rect -38630 7275 -38620 7310
rect -38585 7275 -38575 7310
rect -38540 7275 -38530 7310
rect -38495 7275 -38485 7310
rect -38450 7275 -38440 7310
rect -38405 7275 -38395 7310
rect -38360 7275 -38350 7310
rect -38315 7275 -38305 7310
rect -38270 7275 -38260 7310
rect -38225 7275 -38215 7310
rect -38180 7275 -38170 7310
rect -38135 7275 -38125 7310
rect -38090 7275 -38080 7310
rect -38045 7275 -38035 7310
rect -38000 7275 -37990 7310
rect -37955 7275 -37945 7310
rect -37910 7275 -37900 7310
rect -37865 7275 -37855 7310
rect -37820 7275 -37810 7310
rect -37775 7275 -37765 7310
rect -37730 7275 -37720 7310
rect -37685 7275 -37675 7310
rect -37640 7275 -37630 7310
rect -37595 7275 -37585 7310
rect -37550 7275 -37540 7310
rect -37505 7275 -37495 7310
rect -37460 7275 -37450 7310
rect -37415 7275 -37405 7310
rect -37370 7275 -37360 7310
rect -37325 7275 -37315 7310
rect -37280 7275 -37270 7310
rect -37235 7275 -37225 7310
rect -37190 7275 -37170 7310
rect -38770 7265 -37170 7275
rect -38770 7230 -38755 7265
rect -38720 7230 -38710 7265
rect -38675 7230 -38665 7265
rect -38630 7230 -38620 7265
rect -38585 7230 -38575 7265
rect -38540 7230 -38530 7265
rect -38495 7230 -38485 7265
rect -38450 7230 -38440 7265
rect -38405 7230 -38395 7265
rect -38360 7230 -38350 7265
rect -38315 7230 -38305 7265
rect -38270 7230 -38260 7265
rect -38225 7230 -38215 7265
rect -38180 7230 -38170 7265
rect -38135 7230 -38125 7265
rect -38090 7230 -38080 7265
rect -38045 7230 -38035 7265
rect -38000 7230 -37990 7265
rect -37955 7230 -37945 7265
rect -37910 7230 -37900 7265
rect -37865 7230 -37855 7265
rect -37820 7230 -37810 7265
rect -37775 7230 -37765 7265
rect -37730 7230 -37720 7265
rect -37685 7230 -37675 7265
rect -37640 7230 -37630 7265
rect -37595 7230 -37585 7265
rect -37550 7230 -37540 7265
rect -37505 7230 -37495 7265
rect -37460 7230 -37450 7265
rect -37415 7230 -37405 7265
rect -37370 7230 -37360 7265
rect -37325 7230 -37315 7265
rect -37280 7230 -37270 7265
rect -37235 7230 -37225 7265
rect -37190 7230 -37170 7265
rect -38770 7220 -37170 7230
rect -38770 7185 -38755 7220
rect -38720 7185 -38710 7220
rect -38675 7185 -38665 7220
rect -38630 7185 -38620 7220
rect -38585 7185 -38575 7220
rect -38540 7185 -38530 7220
rect -38495 7185 -38485 7220
rect -38450 7185 -38440 7220
rect -38405 7185 -38395 7220
rect -38360 7185 -38350 7220
rect -38315 7185 -38305 7220
rect -38270 7185 -38260 7220
rect -38225 7185 -38215 7220
rect -38180 7185 -38170 7220
rect -38135 7185 -38125 7220
rect -38090 7185 -38080 7220
rect -38045 7185 -38035 7220
rect -38000 7185 -37990 7220
rect -37955 7185 -37945 7220
rect -37910 7185 -37900 7220
rect -37865 7185 -37855 7220
rect -37820 7185 -37810 7220
rect -37775 7185 -37765 7220
rect -37730 7185 -37720 7220
rect -37685 7185 -37675 7220
rect -37640 7185 -37630 7220
rect -37595 7185 -37585 7220
rect -37550 7185 -37540 7220
rect -37505 7185 -37495 7220
rect -37460 7185 -37450 7220
rect -37415 7185 -37405 7220
rect -37370 7185 -37360 7220
rect -37325 7185 -37315 7220
rect -37280 7185 -37270 7220
rect -37235 7185 -37225 7220
rect -37190 7185 -37170 7220
rect -38770 7175 -37170 7185
rect -38770 7140 -38755 7175
rect -38720 7140 -38710 7175
rect -38675 7140 -38665 7175
rect -38630 7140 -38620 7175
rect -38585 7140 -38575 7175
rect -38540 7140 -38530 7175
rect -38495 7140 -38485 7175
rect -38450 7140 -38440 7175
rect -38405 7140 -38395 7175
rect -38360 7140 -38350 7175
rect -38315 7140 -38305 7175
rect -38270 7140 -38260 7175
rect -38225 7140 -38215 7175
rect -38180 7140 -38170 7175
rect -38135 7140 -38125 7175
rect -38090 7140 -38080 7175
rect -38045 7140 -38035 7175
rect -38000 7140 -37990 7175
rect -37955 7140 -37945 7175
rect -37910 7140 -37900 7175
rect -37865 7140 -37855 7175
rect -37820 7140 -37810 7175
rect -37775 7140 -37765 7175
rect -37730 7140 -37720 7175
rect -37685 7140 -37675 7175
rect -37640 7140 -37630 7175
rect -37595 7140 -37585 7175
rect -37550 7140 -37540 7175
rect -37505 7140 -37495 7175
rect -37460 7140 -37450 7175
rect -37415 7140 -37405 7175
rect -37370 7140 -37360 7175
rect -37325 7140 -37315 7175
rect -37280 7140 -37270 7175
rect -37235 7140 -37225 7175
rect -37190 7140 -37170 7175
rect -38770 7130 -37170 7140
rect -38770 7095 -38755 7130
rect -38720 7095 -38710 7130
rect -38675 7095 -38665 7130
rect -38630 7095 -38620 7130
rect -38585 7095 -38575 7130
rect -38540 7095 -38530 7130
rect -38495 7095 -38485 7130
rect -38450 7095 -38440 7130
rect -38405 7095 -38395 7130
rect -38360 7095 -38350 7130
rect -38315 7095 -38305 7130
rect -38270 7095 -38260 7130
rect -38225 7095 -38215 7130
rect -38180 7095 -38170 7130
rect -38135 7095 -38125 7130
rect -38090 7095 -38080 7130
rect -38045 7095 -38035 7130
rect -38000 7095 -37990 7130
rect -37955 7095 -37945 7130
rect -37910 7095 -37900 7130
rect -37865 7095 -37855 7130
rect -37820 7095 -37810 7130
rect -37775 7095 -37765 7130
rect -37730 7095 -37720 7130
rect -37685 7095 -37675 7130
rect -37640 7095 -37630 7130
rect -37595 7095 -37585 7130
rect -37550 7095 -37540 7130
rect -37505 7095 -37495 7130
rect -37460 7095 -37450 7130
rect -37415 7095 -37405 7130
rect -37370 7095 -37360 7130
rect -37325 7095 -37315 7130
rect -37280 7095 -37270 7130
rect -37235 7095 -37225 7130
rect -37190 7095 -37170 7130
rect -38770 7085 -37170 7095
rect -38770 7050 -38755 7085
rect -38720 7050 -38710 7085
rect -38675 7050 -38665 7085
rect -38630 7050 -38620 7085
rect -38585 7050 -38575 7085
rect -38540 7050 -38530 7085
rect -38495 7050 -38485 7085
rect -38450 7050 -38440 7085
rect -38405 7050 -38395 7085
rect -38360 7050 -38350 7085
rect -38315 7050 -38305 7085
rect -38270 7050 -38260 7085
rect -38225 7050 -38215 7085
rect -38180 7050 -38170 7085
rect -38135 7050 -38125 7085
rect -38090 7050 -38080 7085
rect -38045 7050 -38035 7085
rect -38000 7050 -37990 7085
rect -37955 7050 -37945 7085
rect -37910 7050 -37900 7085
rect -37865 7050 -37855 7085
rect -37820 7050 -37810 7085
rect -37775 7050 -37765 7085
rect -37730 7050 -37720 7085
rect -37685 7050 -37675 7085
rect -37640 7050 -37630 7085
rect -37595 7050 -37585 7085
rect -37550 7050 -37540 7085
rect -37505 7050 -37495 7085
rect -37460 7050 -37450 7085
rect -37415 7050 -37405 7085
rect -37370 7050 -37360 7085
rect -37325 7050 -37315 7085
rect -37280 7050 -37270 7085
rect -37235 7050 -37225 7085
rect -37190 7050 -37170 7085
rect -38770 7040 -37170 7050
rect -38770 7005 -38755 7040
rect -38720 7005 -38710 7040
rect -38675 7005 -38665 7040
rect -38630 7005 -38620 7040
rect -38585 7005 -38575 7040
rect -38540 7005 -38530 7040
rect -38495 7005 -38485 7040
rect -38450 7005 -38440 7040
rect -38405 7005 -38395 7040
rect -38360 7005 -38350 7040
rect -38315 7005 -38305 7040
rect -38270 7005 -38260 7040
rect -38225 7005 -38215 7040
rect -38180 7005 -38170 7040
rect -38135 7005 -38125 7040
rect -38090 7005 -38080 7040
rect -38045 7005 -38035 7040
rect -38000 7005 -37990 7040
rect -37955 7005 -37945 7040
rect -37910 7005 -37900 7040
rect -37865 7005 -37855 7040
rect -37820 7005 -37810 7040
rect -37775 7005 -37765 7040
rect -37730 7005 -37720 7040
rect -37685 7005 -37675 7040
rect -37640 7005 -37630 7040
rect -37595 7005 -37585 7040
rect -37550 7005 -37540 7040
rect -37505 7005 -37495 7040
rect -37460 7005 -37450 7040
rect -37415 7005 -37405 7040
rect -37370 7005 -37360 7040
rect -37325 7005 -37315 7040
rect -37280 7005 -37270 7040
rect -37235 7005 -37225 7040
rect -37190 7005 -37170 7040
rect -38770 6995 -37170 7005
rect -38770 6960 -38755 6995
rect -38720 6960 -38710 6995
rect -38675 6960 -38665 6995
rect -38630 6960 -38620 6995
rect -38585 6960 -38575 6995
rect -38540 6960 -38530 6995
rect -38495 6960 -38485 6995
rect -38450 6960 -38440 6995
rect -38405 6960 -38395 6995
rect -38360 6960 -38350 6995
rect -38315 6960 -38305 6995
rect -38270 6960 -38260 6995
rect -38225 6960 -38215 6995
rect -38180 6960 -38170 6995
rect -38135 6960 -38125 6995
rect -38090 6960 -38080 6995
rect -38045 6960 -38035 6995
rect -38000 6960 -37990 6995
rect -37955 6960 -37945 6995
rect -37910 6960 -37900 6995
rect -37865 6960 -37855 6995
rect -37820 6960 -37810 6995
rect -37775 6960 -37765 6995
rect -37730 6960 -37720 6995
rect -37685 6960 -37675 6995
rect -37640 6960 -37630 6995
rect -37595 6960 -37585 6995
rect -37550 6960 -37540 6995
rect -37505 6960 -37495 6995
rect -37460 6960 -37450 6995
rect -37415 6960 -37405 6995
rect -37370 6960 -37360 6995
rect -37325 6960 -37315 6995
rect -37280 6960 -37270 6995
rect -37235 6960 -37225 6995
rect -37190 6960 -37170 6995
rect -38770 6950 -37170 6960
rect -38770 6915 -38755 6950
rect -38720 6915 -38710 6950
rect -38675 6915 -38665 6950
rect -38630 6915 -38620 6950
rect -38585 6915 -38575 6950
rect -38540 6915 -38530 6950
rect -38495 6915 -38485 6950
rect -38450 6915 -38440 6950
rect -38405 6915 -38395 6950
rect -38360 6915 -38350 6950
rect -38315 6915 -38305 6950
rect -38270 6915 -38260 6950
rect -38225 6915 -38215 6950
rect -38180 6915 -38170 6950
rect -38135 6915 -38125 6950
rect -38090 6915 -38080 6950
rect -38045 6915 -38035 6950
rect -38000 6915 -37990 6950
rect -37955 6915 -37945 6950
rect -37910 6915 -37900 6950
rect -37865 6915 -37855 6950
rect -37820 6915 -37810 6950
rect -37775 6915 -37765 6950
rect -37730 6915 -37720 6950
rect -37685 6915 -37675 6950
rect -37640 6915 -37630 6950
rect -37595 6915 -37585 6950
rect -37550 6915 -37540 6950
rect -37505 6915 -37495 6950
rect -37460 6915 -37450 6950
rect -37415 6915 -37405 6950
rect -37370 6915 -37360 6950
rect -37325 6915 -37315 6950
rect -37280 6915 -37270 6950
rect -37235 6915 -37225 6950
rect -37190 6915 -37170 6950
rect -38770 6905 -37170 6915
rect -38770 6870 -38755 6905
rect -38720 6870 -38710 6905
rect -38675 6870 -38665 6905
rect -38630 6870 -38620 6905
rect -38585 6870 -38575 6905
rect -38540 6870 -38530 6905
rect -38495 6870 -38485 6905
rect -38450 6870 -38440 6905
rect -38405 6870 -38395 6905
rect -38360 6870 -38350 6905
rect -38315 6870 -38305 6905
rect -38270 6870 -38260 6905
rect -38225 6870 -38215 6905
rect -38180 6870 -38170 6905
rect -38135 6870 -38125 6905
rect -38090 6870 -38080 6905
rect -38045 6870 -38035 6905
rect -38000 6870 -37990 6905
rect -37955 6870 -37945 6905
rect -37910 6870 -37900 6905
rect -37865 6870 -37855 6905
rect -37820 6870 -37810 6905
rect -37775 6870 -37765 6905
rect -37730 6870 -37720 6905
rect -37685 6870 -37675 6905
rect -37640 6870 -37630 6905
rect -37595 6870 -37585 6905
rect -37550 6870 -37540 6905
rect -37505 6870 -37495 6905
rect -37460 6870 -37450 6905
rect -37415 6870 -37405 6905
rect -37370 6870 -37360 6905
rect -37325 6870 -37315 6905
rect -37280 6870 -37270 6905
rect -37235 6870 -37225 6905
rect -37190 6870 -37170 6905
rect -38770 6860 -37170 6870
rect -38770 6825 -38755 6860
rect -38720 6825 -38710 6860
rect -38675 6825 -38665 6860
rect -38630 6825 -38620 6860
rect -38585 6825 -38575 6860
rect -38540 6825 -38530 6860
rect -38495 6825 -38485 6860
rect -38450 6825 -38440 6860
rect -38405 6825 -38395 6860
rect -38360 6825 -38350 6860
rect -38315 6825 -38305 6860
rect -38270 6825 -38260 6860
rect -38225 6825 -38215 6860
rect -38180 6825 -38170 6860
rect -38135 6825 -38125 6860
rect -38090 6825 -38080 6860
rect -38045 6825 -38035 6860
rect -38000 6825 -37990 6860
rect -37955 6825 -37945 6860
rect -37910 6825 -37900 6860
rect -37865 6825 -37855 6860
rect -37820 6825 -37810 6860
rect -37775 6825 -37765 6860
rect -37730 6825 -37720 6860
rect -37685 6825 -37675 6860
rect -37640 6825 -37630 6860
rect -37595 6825 -37585 6860
rect -37550 6825 -37540 6860
rect -37505 6825 -37495 6860
rect -37460 6825 -37450 6860
rect -37415 6825 -37405 6860
rect -37370 6825 -37360 6860
rect -37325 6825 -37315 6860
rect -37280 6825 -37270 6860
rect -37235 6825 -37225 6860
rect -37190 6825 -37170 6860
rect -38770 6815 -37170 6825
rect -38770 6780 -38755 6815
rect -38720 6780 -38710 6815
rect -38675 6780 -38665 6815
rect -38630 6780 -38620 6815
rect -38585 6780 -38575 6815
rect -38540 6780 -38530 6815
rect -38495 6780 -38485 6815
rect -38450 6780 -38440 6815
rect -38405 6780 -38395 6815
rect -38360 6780 -38350 6815
rect -38315 6780 -38305 6815
rect -38270 6780 -38260 6815
rect -38225 6780 -38215 6815
rect -38180 6780 -38170 6815
rect -38135 6780 -38125 6815
rect -38090 6780 -38080 6815
rect -38045 6780 -38035 6815
rect -38000 6780 -37990 6815
rect -37955 6780 -37945 6815
rect -37910 6780 -37900 6815
rect -37865 6780 -37855 6815
rect -37820 6780 -37810 6815
rect -37775 6780 -37765 6815
rect -37730 6780 -37720 6815
rect -37685 6780 -37675 6815
rect -37640 6780 -37630 6815
rect -37595 6780 -37585 6815
rect -37550 6780 -37540 6815
rect -37505 6780 -37495 6815
rect -37460 6780 -37450 6815
rect -37415 6780 -37405 6815
rect -37370 6780 -37360 6815
rect -37325 6780 -37315 6815
rect -37280 6780 -37270 6815
rect -37235 6780 -37225 6815
rect -37190 6780 -37170 6815
rect -38770 6770 -37170 6780
rect -38770 6735 -38755 6770
rect -38720 6735 -38710 6770
rect -38675 6735 -38665 6770
rect -38630 6735 -38620 6770
rect -38585 6735 -38575 6770
rect -38540 6735 -38530 6770
rect -38495 6735 -38485 6770
rect -38450 6735 -38440 6770
rect -38405 6735 -38395 6770
rect -38360 6735 -38350 6770
rect -38315 6735 -38305 6770
rect -38270 6735 -38260 6770
rect -38225 6735 -38215 6770
rect -38180 6735 -38170 6770
rect -38135 6735 -38125 6770
rect -38090 6735 -38080 6770
rect -38045 6735 -38035 6770
rect -38000 6735 -37990 6770
rect -37955 6735 -37945 6770
rect -37910 6735 -37900 6770
rect -37865 6735 -37855 6770
rect -37820 6735 -37810 6770
rect -37775 6735 -37765 6770
rect -37730 6735 -37720 6770
rect -37685 6735 -37675 6770
rect -37640 6735 -37630 6770
rect -37595 6735 -37585 6770
rect -37550 6735 -37540 6770
rect -37505 6735 -37495 6770
rect -37460 6735 -37450 6770
rect -37415 6735 -37405 6770
rect -37370 6735 -37360 6770
rect -37325 6735 -37315 6770
rect -37280 6735 -37270 6770
rect -37235 6735 -37225 6770
rect -37190 6735 -37170 6770
rect -38770 6725 -37170 6735
rect -38770 6690 -38755 6725
rect -38720 6690 -38710 6725
rect -38675 6690 -38665 6725
rect -38630 6690 -38620 6725
rect -38585 6690 -38575 6725
rect -38540 6690 -38530 6725
rect -38495 6690 -38485 6725
rect -38450 6690 -38440 6725
rect -38405 6690 -38395 6725
rect -38360 6690 -38350 6725
rect -38315 6690 -38305 6725
rect -38270 6690 -38260 6725
rect -38225 6690 -38215 6725
rect -38180 6690 -38170 6725
rect -38135 6690 -38125 6725
rect -38090 6690 -38080 6725
rect -38045 6690 -38035 6725
rect -38000 6690 -37990 6725
rect -37955 6690 -37945 6725
rect -37910 6690 -37900 6725
rect -37865 6690 -37855 6725
rect -37820 6690 -37810 6725
rect -37775 6690 -37765 6725
rect -37730 6690 -37720 6725
rect -37685 6690 -37675 6725
rect -37640 6690 -37630 6725
rect -37595 6690 -37585 6725
rect -37550 6690 -37540 6725
rect -37505 6690 -37495 6725
rect -37460 6690 -37450 6725
rect -37415 6690 -37405 6725
rect -37370 6690 -37360 6725
rect -37325 6690 -37315 6725
rect -37280 6690 -37270 6725
rect -37235 6690 -37225 6725
rect -37190 6690 -37170 6725
rect -38770 6680 -37170 6690
rect -38770 6645 -38755 6680
rect -38720 6645 -38710 6680
rect -38675 6645 -38665 6680
rect -38630 6645 -38620 6680
rect -38585 6645 -38575 6680
rect -38540 6645 -38530 6680
rect -38495 6645 -38485 6680
rect -38450 6645 -38440 6680
rect -38405 6645 -38395 6680
rect -38360 6645 -38350 6680
rect -38315 6645 -38305 6680
rect -38270 6645 -38260 6680
rect -38225 6645 -38215 6680
rect -38180 6645 -38170 6680
rect -38135 6645 -38125 6680
rect -38090 6645 -38080 6680
rect -38045 6645 -38035 6680
rect -38000 6645 -37990 6680
rect -37955 6645 -37945 6680
rect -37910 6645 -37900 6680
rect -37865 6645 -37855 6680
rect -37820 6645 -37810 6680
rect -37775 6645 -37765 6680
rect -37730 6645 -37720 6680
rect -37685 6645 -37675 6680
rect -37640 6645 -37630 6680
rect -37595 6645 -37585 6680
rect -37550 6645 -37540 6680
rect -37505 6645 -37495 6680
rect -37460 6645 -37450 6680
rect -37415 6645 -37405 6680
rect -37370 6645 -37360 6680
rect -37325 6645 -37315 6680
rect -37280 6645 -37270 6680
rect -37235 6645 -37225 6680
rect -37190 6645 -37170 6680
rect -38770 6635 -37170 6645
rect -38770 6600 -38755 6635
rect -38720 6600 -38710 6635
rect -38675 6600 -38665 6635
rect -38630 6600 -38620 6635
rect -38585 6600 -38575 6635
rect -38540 6600 -38530 6635
rect -38495 6600 -38485 6635
rect -38450 6600 -38440 6635
rect -38405 6600 -38395 6635
rect -38360 6600 -38350 6635
rect -38315 6600 -38305 6635
rect -38270 6600 -38260 6635
rect -38225 6600 -38215 6635
rect -38180 6600 -38170 6635
rect -38135 6600 -38125 6635
rect -38090 6600 -38080 6635
rect -38045 6600 -38035 6635
rect -38000 6600 -37990 6635
rect -37955 6600 -37945 6635
rect -37910 6600 -37900 6635
rect -37865 6600 -37855 6635
rect -37820 6600 -37810 6635
rect -37775 6600 -37765 6635
rect -37730 6600 -37720 6635
rect -37685 6600 -37675 6635
rect -37640 6600 -37630 6635
rect -37595 6600 -37585 6635
rect -37550 6600 -37540 6635
rect -37505 6600 -37495 6635
rect -37460 6600 -37450 6635
rect -37415 6600 -37405 6635
rect -37370 6600 -37360 6635
rect -37325 6600 -37315 6635
rect -37280 6600 -37270 6635
rect -37235 6600 -37225 6635
rect -37190 6600 -37170 6635
rect -38770 6590 -37170 6600
rect -38770 6555 -38755 6590
rect -38720 6555 -38710 6590
rect -38675 6555 -38665 6590
rect -38630 6555 -38620 6590
rect -38585 6555 -38575 6590
rect -38540 6555 -38530 6590
rect -38495 6555 -38485 6590
rect -38450 6555 -38440 6590
rect -38405 6555 -38395 6590
rect -38360 6555 -38350 6590
rect -38315 6555 -38305 6590
rect -38270 6555 -38260 6590
rect -38225 6555 -38215 6590
rect -38180 6555 -38170 6590
rect -38135 6555 -38125 6590
rect -38090 6555 -38080 6590
rect -38045 6555 -38035 6590
rect -38000 6555 -37990 6590
rect -37955 6555 -37945 6590
rect -37910 6555 -37900 6590
rect -37865 6555 -37855 6590
rect -37820 6555 -37810 6590
rect -37775 6555 -37765 6590
rect -37730 6555 -37720 6590
rect -37685 6555 -37675 6590
rect -37640 6555 -37630 6590
rect -37595 6555 -37585 6590
rect -37550 6555 -37540 6590
rect -37505 6555 -37495 6590
rect -37460 6555 -37450 6590
rect -37415 6555 -37405 6590
rect -37370 6555 -37360 6590
rect -37325 6555 -37315 6590
rect -37280 6555 -37270 6590
rect -37235 6555 -37225 6590
rect -37190 6555 -37170 6590
rect -38770 6545 -37170 6555
rect -38770 6510 -38755 6545
rect -38720 6510 -38710 6545
rect -38675 6510 -38665 6545
rect -38630 6510 -38620 6545
rect -38585 6510 -38575 6545
rect -38540 6510 -38530 6545
rect -38495 6510 -38485 6545
rect -38450 6510 -38440 6545
rect -38405 6510 -38395 6545
rect -38360 6510 -38350 6545
rect -38315 6510 -38305 6545
rect -38270 6510 -38260 6545
rect -38225 6510 -38215 6545
rect -38180 6510 -38170 6545
rect -38135 6510 -38125 6545
rect -38090 6510 -38080 6545
rect -38045 6510 -38035 6545
rect -38000 6510 -37990 6545
rect -37955 6510 -37945 6545
rect -37910 6510 -37900 6545
rect -37865 6510 -37855 6545
rect -37820 6510 -37810 6545
rect -37775 6510 -37765 6545
rect -37730 6510 -37720 6545
rect -37685 6510 -37675 6545
rect -37640 6510 -37630 6545
rect -37595 6510 -37585 6545
rect -37550 6510 -37540 6545
rect -37505 6510 -37495 6545
rect -37460 6510 -37450 6545
rect -37415 6510 -37405 6545
rect -37370 6510 -37360 6545
rect -37325 6510 -37315 6545
rect -37280 6510 -37270 6545
rect -37235 6510 -37225 6545
rect -37190 6510 -37170 6545
rect -38770 6500 -37170 6510
rect -38770 6465 -38755 6500
rect -38720 6465 -38710 6500
rect -38675 6465 -38665 6500
rect -38630 6465 -38620 6500
rect -38585 6465 -38575 6500
rect -38540 6465 -38530 6500
rect -38495 6465 -38485 6500
rect -38450 6465 -38440 6500
rect -38405 6465 -38395 6500
rect -38360 6465 -38350 6500
rect -38315 6465 -38305 6500
rect -38270 6465 -38260 6500
rect -38225 6465 -38215 6500
rect -38180 6465 -38170 6500
rect -38135 6465 -38125 6500
rect -38090 6465 -38080 6500
rect -38045 6465 -38035 6500
rect -38000 6465 -37990 6500
rect -37955 6465 -37945 6500
rect -37910 6465 -37900 6500
rect -37865 6465 -37855 6500
rect -37820 6465 -37810 6500
rect -37775 6465 -37765 6500
rect -37730 6465 -37720 6500
rect -37685 6465 -37675 6500
rect -37640 6465 -37630 6500
rect -37595 6465 -37585 6500
rect -37550 6465 -37540 6500
rect -37505 6465 -37495 6500
rect -37460 6465 -37450 6500
rect -37415 6465 -37405 6500
rect -37370 6465 -37360 6500
rect -37325 6465 -37315 6500
rect -37280 6465 -37270 6500
rect -37235 6465 -37225 6500
rect -37190 6465 -37170 6500
rect -38770 6450 -37170 6465
rect -90 9640 -30 9650
rect -90 9600 -80 9640
rect -40 9600 -30 9640
rect -90 9575 -30 9600
rect -90 9535 -80 9575
rect -40 9535 -30 9575
rect -90 9505 -30 9535
rect -90 9465 -80 9505
rect -40 9465 -30 9505
rect -90 9435 -30 9465
rect -90 9395 -80 9435
rect -40 9395 -30 9435
rect -90 9365 -30 9395
rect -90 9325 -80 9365
rect -40 9325 -30 9365
rect -90 9300 -30 9325
rect -90 9260 -80 9300
rect -40 9260 -30 9300
rect -90 9240 -30 9260
rect -90 9200 -80 9240
rect -40 9200 -30 9240
rect -90 9175 -30 9200
rect -90 9135 -80 9175
rect -40 9135 -30 9175
rect -90 9105 -30 9135
rect -90 9065 -80 9105
rect -40 9065 -30 9105
rect -90 9035 -30 9065
rect -90 8995 -80 9035
rect -40 8995 -30 9035
rect -90 8965 -30 8995
rect -90 8925 -80 8965
rect -40 8925 -30 8965
rect -90 8900 -30 8925
rect -90 8860 -80 8900
rect -40 8860 -30 8900
rect -90 8840 -30 8860
rect -90 8800 -80 8840
rect -40 8800 -30 8840
rect -90 8775 -30 8800
rect -90 8735 -80 8775
rect -40 8735 -30 8775
rect -90 8705 -30 8735
rect -90 8665 -80 8705
rect -40 8665 -30 8705
rect -90 8635 -30 8665
rect -90 8595 -80 8635
rect -40 8595 -30 8635
rect -90 8565 -30 8595
rect -90 8525 -80 8565
rect -40 8525 -30 8565
rect -90 8500 -30 8525
rect -90 8460 -80 8500
rect -40 8460 -30 8500
rect -90 8440 -30 8460
rect -90 8400 -80 8440
rect -40 8400 -30 8440
rect -90 8375 -30 8400
rect -90 8335 -80 8375
rect -40 8335 -30 8375
rect -90 8305 -30 8335
rect -90 8265 -80 8305
rect -40 8265 -30 8305
rect -90 8235 -30 8265
rect -90 8195 -80 8235
rect -40 8195 -30 8235
rect -90 8165 -30 8195
rect -90 8125 -80 8165
rect -40 8125 -30 8165
rect -90 8100 -30 8125
rect -90 8060 -80 8100
rect -40 8060 -30 8100
rect -90 8040 -30 8060
rect -90 8000 -80 8040
rect -40 8000 -30 8040
rect -90 7975 -30 8000
rect -90 7935 -80 7975
rect -40 7935 -30 7975
rect -90 7905 -30 7935
rect -90 7865 -80 7905
rect -40 7865 -30 7905
rect -90 7835 -30 7865
rect -90 7795 -80 7835
rect -40 7795 -30 7835
rect -90 7765 -30 7795
rect -90 7725 -80 7765
rect -40 7725 -30 7765
rect -90 7700 -30 7725
rect -90 7660 -80 7700
rect -40 7660 -30 7700
rect -90 7640 -30 7660
rect -90 7600 -80 7640
rect -40 7600 -30 7640
rect -90 7575 -30 7600
rect -90 7535 -80 7575
rect -40 7535 -30 7575
rect -90 7505 -30 7535
rect -90 7465 -80 7505
rect -40 7465 -30 7505
rect -90 7435 -30 7465
rect -90 7395 -80 7435
rect -40 7395 -30 7435
rect -90 7365 -30 7395
rect -90 7325 -80 7365
rect -40 7325 -30 7365
rect -90 7300 -30 7325
rect -90 7260 -80 7300
rect -40 7260 -30 7300
rect -90 7240 -30 7260
rect -90 7200 -80 7240
rect -40 7200 -30 7240
rect -90 7175 -30 7200
rect -90 7135 -80 7175
rect -40 7135 -30 7175
rect -90 7105 -30 7135
rect -90 7065 -80 7105
rect -40 7065 -30 7105
rect -90 7035 -30 7065
rect -90 6995 -80 7035
rect -40 6995 -30 7035
rect -90 6965 -30 6995
rect -90 6925 -80 6965
rect -40 6925 -30 6965
rect -90 6900 -30 6925
rect -90 6860 -80 6900
rect -40 6860 -30 6900
rect -90 6840 -30 6860
rect -90 6800 -80 6840
rect -40 6800 -30 6840
rect -90 6775 -30 6800
rect -90 6735 -80 6775
rect -40 6735 -30 6775
rect -90 6705 -30 6735
rect -90 6665 -80 6705
rect -40 6665 -30 6705
rect -90 6635 -30 6665
rect -90 6595 -80 6635
rect -40 6595 -30 6635
rect -90 6565 -30 6595
rect -90 6525 -80 6565
rect -40 6525 -30 6565
rect -90 6500 -30 6525
rect -90 6460 -80 6500
rect -40 6460 -30 6500
rect -90 6450 -30 6460
rect 260 9640 320 9650
rect 260 9600 270 9640
rect 310 9600 320 9640
rect 260 9575 320 9600
rect 260 9535 270 9575
rect 310 9535 320 9575
rect 260 9505 320 9535
rect 260 9465 270 9505
rect 310 9465 320 9505
rect 260 9435 320 9465
rect 260 9395 270 9435
rect 310 9395 320 9435
rect 260 9365 320 9395
rect 260 9325 270 9365
rect 310 9325 320 9365
rect 260 9300 320 9325
rect 260 9260 270 9300
rect 310 9260 320 9300
rect 260 9240 320 9260
rect 260 9200 270 9240
rect 310 9200 320 9240
rect 260 9175 320 9200
rect 260 9135 270 9175
rect 310 9135 320 9175
rect 260 9105 320 9135
rect 260 9065 270 9105
rect 310 9065 320 9105
rect 260 9035 320 9065
rect 260 8995 270 9035
rect 310 8995 320 9035
rect 260 8965 320 8995
rect 260 8925 270 8965
rect 310 8925 320 8965
rect 260 8900 320 8925
rect 260 8860 270 8900
rect 310 8860 320 8900
rect 260 8840 320 8860
rect 260 8800 270 8840
rect 310 8800 320 8840
rect 260 8775 320 8800
rect 260 8735 270 8775
rect 310 8735 320 8775
rect 260 8705 320 8735
rect 260 8665 270 8705
rect 310 8665 320 8705
rect 260 8635 320 8665
rect 260 8595 270 8635
rect 310 8595 320 8635
rect 260 8565 320 8595
rect 260 8525 270 8565
rect 310 8525 320 8565
rect 260 8500 320 8525
rect 260 8460 270 8500
rect 310 8460 320 8500
rect 260 8440 320 8460
rect 260 8400 270 8440
rect 310 8400 320 8440
rect 260 8375 320 8400
rect 260 8335 270 8375
rect 310 8335 320 8375
rect 260 8305 320 8335
rect 260 8265 270 8305
rect 310 8265 320 8305
rect 260 8235 320 8265
rect 260 8195 270 8235
rect 310 8195 320 8235
rect 260 8165 320 8195
rect 260 8125 270 8165
rect 310 8125 320 8165
rect 260 8100 320 8125
rect 260 8060 270 8100
rect 310 8060 320 8100
rect 260 8040 320 8060
rect 260 8000 270 8040
rect 310 8000 320 8040
rect 260 7975 320 8000
rect 260 7935 270 7975
rect 310 7935 320 7975
rect 260 7905 320 7935
rect 260 7865 270 7905
rect 310 7865 320 7905
rect 260 7835 320 7865
rect 260 7795 270 7835
rect 310 7795 320 7835
rect 260 7765 320 7795
rect 260 7725 270 7765
rect 310 7725 320 7765
rect 260 7700 320 7725
rect 260 7660 270 7700
rect 310 7660 320 7700
rect 260 7640 320 7660
rect 260 7600 270 7640
rect 310 7600 320 7640
rect 260 7575 320 7600
rect 260 7535 270 7575
rect 310 7535 320 7575
rect 260 7505 320 7535
rect 260 7465 270 7505
rect 310 7465 320 7505
rect 260 7435 320 7465
rect 260 7395 270 7435
rect 310 7395 320 7435
rect 260 7365 320 7395
rect 260 7325 270 7365
rect 310 7325 320 7365
rect 260 7300 320 7325
rect 260 7260 270 7300
rect 310 7260 320 7300
rect 260 7240 320 7260
rect 260 7200 270 7240
rect 310 7200 320 7240
rect 260 7175 320 7200
rect 260 7135 270 7175
rect 310 7135 320 7175
rect 260 7105 320 7135
rect 260 7065 270 7105
rect 310 7065 320 7105
rect 260 7035 320 7065
rect 260 6995 270 7035
rect 310 6995 320 7035
rect 260 6965 320 6995
rect 260 6925 270 6965
rect 310 6925 320 6965
rect 260 6900 320 6925
rect 260 6860 270 6900
rect 310 6860 320 6900
rect 260 6840 320 6860
rect 260 6800 270 6840
rect 310 6800 320 6840
rect 260 6775 320 6800
rect 260 6735 270 6775
rect 310 6735 320 6775
rect 260 6705 320 6735
rect 260 6665 270 6705
rect 310 6665 320 6705
rect 260 6635 320 6665
rect 260 6595 270 6635
rect 310 6595 320 6635
rect 260 6565 320 6595
rect 260 6525 270 6565
rect 310 6525 320 6565
rect 260 6500 320 6525
rect 260 6460 270 6500
rect 310 6460 320 6500
rect 260 6450 320 6460
rect 610 9640 670 9650
rect 610 9600 620 9640
rect 660 9600 670 9640
rect 610 9575 670 9600
rect 610 9535 620 9575
rect 660 9535 670 9575
rect 610 9505 670 9535
rect 610 9465 620 9505
rect 660 9465 670 9505
rect 610 9435 670 9465
rect 610 9395 620 9435
rect 660 9395 670 9435
rect 610 9365 670 9395
rect 610 9325 620 9365
rect 660 9325 670 9365
rect 610 9300 670 9325
rect 610 9260 620 9300
rect 660 9260 670 9300
rect 610 9240 670 9260
rect 610 9200 620 9240
rect 660 9200 670 9240
rect 610 9175 670 9200
rect 610 9135 620 9175
rect 660 9135 670 9175
rect 610 9105 670 9135
rect 610 9065 620 9105
rect 660 9065 670 9105
rect 610 9035 670 9065
rect 610 8995 620 9035
rect 660 8995 670 9035
rect 610 8965 670 8995
rect 610 8925 620 8965
rect 660 8925 670 8965
rect 610 8900 670 8925
rect 610 8860 620 8900
rect 660 8860 670 8900
rect 610 8840 670 8860
rect 610 8800 620 8840
rect 660 8800 670 8840
rect 610 8775 670 8800
rect 610 8735 620 8775
rect 660 8735 670 8775
rect 610 8705 670 8735
rect 610 8665 620 8705
rect 660 8665 670 8705
rect 610 8635 670 8665
rect 610 8595 620 8635
rect 660 8595 670 8635
rect 610 8565 670 8595
rect 610 8525 620 8565
rect 660 8525 670 8565
rect 610 8500 670 8525
rect 610 8460 620 8500
rect 660 8460 670 8500
rect 610 8440 670 8460
rect 610 8400 620 8440
rect 660 8400 670 8440
rect 610 8375 670 8400
rect 610 8335 620 8375
rect 660 8335 670 8375
rect 610 8305 670 8335
rect 610 8265 620 8305
rect 660 8265 670 8305
rect 610 8235 670 8265
rect 610 8195 620 8235
rect 660 8195 670 8235
rect 610 8165 670 8195
rect 610 8125 620 8165
rect 660 8125 670 8165
rect 610 8100 670 8125
rect 610 8060 620 8100
rect 660 8060 670 8100
rect 610 8040 670 8060
rect 610 8000 620 8040
rect 660 8000 670 8040
rect 610 7975 670 8000
rect 610 7935 620 7975
rect 660 7935 670 7975
rect 610 7905 670 7935
rect 610 7865 620 7905
rect 660 7865 670 7905
rect 610 7835 670 7865
rect 610 7795 620 7835
rect 660 7795 670 7835
rect 610 7765 670 7795
rect 610 7725 620 7765
rect 660 7725 670 7765
rect 610 7700 670 7725
rect 610 7660 620 7700
rect 660 7660 670 7700
rect 610 7640 670 7660
rect 610 7600 620 7640
rect 660 7600 670 7640
rect 610 7575 670 7600
rect 610 7535 620 7575
rect 660 7535 670 7575
rect 610 7505 670 7535
rect 610 7465 620 7505
rect 660 7465 670 7505
rect 610 7435 670 7465
rect 610 7395 620 7435
rect 660 7395 670 7435
rect 610 7365 670 7395
rect 610 7325 620 7365
rect 660 7325 670 7365
rect 610 7300 670 7325
rect 610 7260 620 7300
rect 660 7260 670 7300
rect 610 7240 670 7260
rect 610 7200 620 7240
rect 660 7200 670 7240
rect 610 7175 670 7200
rect 610 7135 620 7175
rect 660 7135 670 7175
rect 610 7105 670 7135
rect 610 7065 620 7105
rect 660 7065 670 7105
rect 610 7035 670 7065
rect 610 6995 620 7035
rect 660 6995 670 7035
rect 610 6965 670 6995
rect 610 6925 620 6965
rect 660 6925 670 6965
rect 610 6900 670 6925
rect 610 6860 620 6900
rect 660 6860 670 6900
rect 610 6840 670 6860
rect 610 6800 620 6840
rect 660 6800 670 6840
rect 610 6775 670 6800
rect 610 6735 620 6775
rect 660 6735 670 6775
rect 610 6705 670 6735
rect 610 6665 620 6705
rect 660 6665 670 6705
rect 610 6635 670 6665
rect 610 6595 620 6635
rect 660 6595 670 6635
rect 610 6565 670 6595
rect 610 6525 620 6565
rect 660 6525 670 6565
rect 610 6500 670 6525
rect 610 6460 620 6500
rect 660 6460 670 6500
rect 610 6450 670 6460
rect 960 9640 1020 9650
rect 960 9600 970 9640
rect 1010 9600 1020 9640
rect 960 9575 1020 9600
rect 960 9535 970 9575
rect 1010 9535 1020 9575
rect 960 9505 1020 9535
rect 960 9465 970 9505
rect 1010 9465 1020 9505
rect 960 9435 1020 9465
rect 960 9395 970 9435
rect 1010 9395 1020 9435
rect 960 9365 1020 9395
rect 960 9325 970 9365
rect 1010 9325 1020 9365
rect 960 9300 1020 9325
rect 960 9260 970 9300
rect 1010 9260 1020 9300
rect 960 9240 1020 9260
rect 960 9200 970 9240
rect 1010 9200 1020 9240
rect 960 9175 1020 9200
rect 960 9135 970 9175
rect 1010 9135 1020 9175
rect 960 9105 1020 9135
rect 960 9065 970 9105
rect 1010 9065 1020 9105
rect 960 9035 1020 9065
rect 960 8995 970 9035
rect 1010 8995 1020 9035
rect 960 8965 1020 8995
rect 960 8925 970 8965
rect 1010 8925 1020 8965
rect 960 8900 1020 8925
rect 960 8860 970 8900
rect 1010 8860 1020 8900
rect 960 8840 1020 8860
rect 960 8800 970 8840
rect 1010 8800 1020 8840
rect 960 8775 1020 8800
rect 960 8735 970 8775
rect 1010 8735 1020 8775
rect 960 8705 1020 8735
rect 960 8665 970 8705
rect 1010 8665 1020 8705
rect 960 8635 1020 8665
rect 960 8595 970 8635
rect 1010 8595 1020 8635
rect 960 8565 1020 8595
rect 960 8525 970 8565
rect 1010 8525 1020 8565
rect 960 8500 1020 8525
rect 960 8460 970 8500
rect 1010 8460 1020 8500
rect 960 8440 1020 8460
rect 960 8400 970 8440
rect 1010 8400 1020 8440
rect 960 8375 1020 8400
rect 960 8335 970 8375
rect 1010 8335 1020 8375
rect 960 8305 1020 8335
rect 960 8265 970 8305
rect 1010 8265 1020 8305
rect 960 8235 1020 8265
rect 960 8195 970 8235
rect 1010 8195 1020 8235
rect 960 8165 1020 8195
rect 960 8125 970 8165
rect 1010 8125 1020 8165
rect 960 8100 1020 8125
rect 960 8060 970 8100
rect 1010 8060 1020 8100
rect 960 8040 1020 8060
rect 960 8000 970 8040
rect 1010 8000 1020 8040
rect 960 7975 1020 8000
rect 960 7935 970 7975
rect 1010 7935 1020 7975
rect 960 7905 1020 7935
rect 960 7865 970 7905
rect 1010 7865 1020 7905
rect 960 7835 1020 7865
rect 960 7795 970 7835
rect 1010 7795 1020 7835
rect 960 7765 1020 7795
rect 960 7725 970 7765
rect 1010 7725 1020 7765
rect 960 7700 1020 7725
rect 960 7660 970 7700
rect 1010 7660 1020 7700
rect 960 7640 1020 7660
rect 960 7600 970 7640
rect 1010 7600 1020 7640
rect 960 7575 1020 7600
rect 960 7535 970 7575
rect 1010 7535 1020 7575
rect 960 7505 1020 7535
rect 960 7465 970 7505
rect 1010 7465 1020 7505
rect 960 7435 1020 7465
rect 960 7395 970 7435
rect 1010 7395 1020 7435
rect 960 7365 1020 7395
rect 960 7325 970 7365
rect 1010 7325 1020 7365
rect 960 7300 1020 7325
rect 960 7260 970 7300
rect 1010 7260 1020 7300
rect 960 7240 1020 7260
rect 960 7200 970 7240
rect 1010 7200 1020 7240
rect 960 7175 1020 7200
rect 960 7135 970 7175
rect 1010 7135 1020 7175
rect 960 7105 1020 7135
rect 960 7065 970 7105
rect 1010 7065 1020 7105
rect 960 7035 1020 7065
rect 960 6995 970 7035
rect 1010 6995 1020 7035
rect 960 6965 1020 6995
rect 960 6925 970 6965
rect 1010 6925 1020 6965
rect 960 6900 1020 6925
rect 960 6860 970 6900
rect 1010 6860 1020 6900
rect 960 6840 1020 6860
rect 960 6800 970 6840
rect 1010 6800 1020 6840
rect 960 6775 1020 6800
rect 960 6735 970 6775
rect 1010 6735 1020 6775
rect 960 6705 1020 6735
rect 960 6665 970 6705
rect 1010 6665 1020 6705
rect 960 6635 1020 6665
rect 960 6595 970 6635
rect 1010 6595 1020 6635
rect 960 6565 1020 6595
rect 960 6525 970 6565
rect 1010 6525 1020 6565
rect 960 6500 1020 6525
rect 960 6460 970 6500
rect 1010 6460 1020 6500
rect 960 6450 1020 6460
rect 1660 9640 1720 9650
rect 1660 9600 1670 9640
rect 1710 9600 1720 9640
rect 1660 9575 1720 9600
rect 1660 9535 1670 9575
rect 1710 9535 1720 9575
rect 1660 9505 1720 9535
rect 1660 9465 1670 9505
rect 1710 9465 1720 9505
rect 1660 9435 1720 9465
rect 1660 9395 1670 9435
rect 1710 9395 1720 9435
rect 1660 9365 1720 9395
rect 1660 9325 1670 9365
rect 1710 9325 1720 9365
rect 1660 9300 1720 9325
rect 1660 9260 1670 9300
rect 1710 9260 1720 9300
rect 1660 9240 1720 9260
rect 1660 9200 1670 9240
rect 1710 9200 1720 9240
rect 1660 9175 1720 9200
rect 1660 9135 1670 9175
rect 1710 9135 1720 9175
rect 1660 9105 1720 9135
rect 1660 9065 1670 9105
rect 1710 9065 1720 9105
rect 1660 9035 1720 9065
rect 1660 8995 1670 9035
rect 1710 8995 1720 9035
rect 1660 8965 1720 8995
rect 1660 8925 1670 8965
rect 1710 8925 1720 8965
rect 1660 8900 1720 8925
rect 1660 8860 1670 8900
rect 1710 8860 1720 8900
rect 1660 8840 1720 8860
rect 1660 8800 1670 8840
rect 1710 8800 1720 8840
rect 1660 8775 1720 8800
rect 1660 8735 1670 8775
rect 1710 8735 1720 8775
rect 1660 8705 1720 8735
rect 1660 8665 1670 8705
rect 1710 8665 1720 8705
rect 1660 8635 1720 8665
rect 1660 8595 1670 8635
rect 1710 8595 1720 8635
rect 1660 8565 1720 8595
rect 1660 8525 1670 8565
rect 1710 8525 1720 8565
rect 1660 8500 1720 8525
rect 1660 8460 1670 8500
rect 1710 8460 1720 8500
rect 1660 8440 1720 8460
rect 1660 8400 1670 8440
rect 1710 8400 1720 8440
rect 1660 8375 1720 8400
rect 1660 8335 1670 8375
rect 1710 8335 1720 8375
rect 1660 8305 1720 8335
rect 1660 8265 1670 8305
rect 1710 8265 1720 8305
rect 1660 8235 1720 8265
rect 1660 8195 1670 8235
rect 1710 8195 1720 8235
rect 1660 8165 1720 8195
rect 1660 8125 1670 8165
rect 1710 8125 1720 8165
rect 1660 8100 1720 8125
rect 1660 8060 1670 8100
rect 1710 8060 1720 8100
rect 1660 8040 1720 8060
rect 1660 8000 1670 8040
rect 1710 8000 1720 8040
rect 1660 7975 1720 8000
rect 1660 7935 1670 7975
rect 1710 7935 1720 7975
rect 1660 7905 1720 7935
rect 1660 7865 1670 7905
rect 1710 7865 1720 7905
rect 1660 7835 1720 7865
rect 1660 7795 1670 7835
rect 1710 7795 1720 7835
rect 1660 7765 1720 7795
rect 1660 7725 1670 7765
rect 1710 7725 1720 7765
rect 1660 7700 1720 7725
rect 1660 7660 1670 7700
rect 1710 7660 1720 7700
rect 1660 7640 1720 7660
rect 1660 7600 1670 7640
rect 1710 7600 1720 7640
rect 1660 7575 1720 7600
rect 1660 7535 1670 7575
rect 1710 7535 1720 7575
rect 1660 7505 1720 7535
rect 1660 7465 1670 7505
rect 1710 7465 1720 7505
rect 1660 7435 1720 7465
rect 1660 7395 1670 7435
rect 1710 7395 1720 7435
rect 1660 7365 1720 7395
rect 1660 7325 1670 7365
rect 1710 7325 1720 7365
rect 1660 7300 1720 7325
rect 1660 7260 1670 7300
rect 1710 7260 1720 7300
rect 1660 7240 1720 7260
rect 1660 7200 1670 7240
rect 1710 7200 1720 7240
rect 1660 7175 1720 7200
rect 1660 7135 1670 7175
rect 1710 7135 1720 7175
rect 1660 7105 1720 7135
rect 1660 7065 1670 7105
rect 1710 7065 1720 7105
rect 1660 7035 1720 7065
rect 1660 6995 1670 7035
rect 1710 6995 1720 7035
rect 1660 6965 1720 6995
rect 1660 6925 1670 6965
rect 1710 6925 1720 6965
rect 1660 6900 1720 6925
rect 1660 6860 1670 6900
rect 1710 6860 1720 6900
rect 1660 6840 1720 6860
rect 1660 6800 1670 6840
rect 1710 6800 1720 6840
rect 1660 6775 1720 6800
rect 1660 6735 1670 6775
rect 1710 6735 1720 6775
rect 1660 6705 1720 6735
rect 1660 6665 1670 6705
rect 1710 6665 1720 6705
rect 1660 6635 1720 6665
rect 1660 6595 1670 6635
rect 1710 6595 1720 6635
rect 1660 6565 1720 6595
rect 1660 6525 1670 6565
rect 1710 6525 1720 6565
rect 1660 6500 1720 6525
rect 1660 6460 1670 6500
rect 1710 6460 1720 6500
rect 1660 6450 1720 6460
rect 2235 9640 2295 9650
rect 2235 9600 2245 9640
rect 2285 9600 2295 9640
rect 2235 9575 2295 9600
rect 2235 9535 2245 9575
rect 2285 9535 2295 9575
rect 2235 9505 2295 9535
rect 2235 9465 2245 9505
rect 2285 9465 2295 9505
rect 2235 9435 2295 9465
rect 2235 9395 2245 9435
rect 2285 9395 2295 9435
rect 2235 9365 2295 9395
rect 2235 9325 2245 9365
rect 2285 9325 2295 9365
rect 2235 9300 2295 9325
rect 2235 9260 2245 9300
rect 2285 9260 2295 9300
rect 2235 9240 2295 9260
rect 2235 9200 2245 9240
rect 2285 9200 2295 9240
rect 2235 9175 2295 9200
rect 2235 9135 2245 9175
rect 2285 9135 2295 9175
rect 2235 9105 2295 9135
rect 2235 9065 2245 9105
rect 2285 9065 2295 9105
rect 2235 9035 2295 9065
rect 2235 8995 2245 9035
rect 2285 8995 2295 9035
rect 2235 8965 2295 8995
rect 2235 8925 2245 8965
rect 2285 8925 2295 8965
rect 2235 8900 2295 8925
rect 2235 8860 2245 8900
rect 2285 8860 2295 8900
rect 2235 8840 2295 8860
rect 2235 8800 2245 8840
rect 2285 8800 2295 8840
rect 2235 8775 2295 8800
rect 2235 8735 2245 8775
rect 2285 8735 2295 8775
rect 2235 8705 2295 8735
rect 2235 8665 2245 8705
rect 2285 8665 2295 8705
rect 2235 8635 2295 8665
rect 2235 8595 2245 8635
rect 2285 8595 2295 8635
rect 2235 8565 2295 8595
rect 2235 8525 2245 8565
rect 2285 8525 2295 8565
rect 2235 8500 2295 8525
rect 2235 8460 2245 8500
rect 2285 8460 2295 8500
rect 2235 8440 2295 8460
rect 2235 8400 2245 8440
rect 2285 8400 2295 8440
rect 2235 8375 2295 8400
rect 2235 8335 2245 8375
rect 2285 8335 2295 8375
rect 2235 8305 2295 8335
rect 2235 8265 2245 8305
rect 2285 8265 2295 8305
rect 2235 8235 2295 8265
rect 2235 8195 2245 8235
rect 2285 8195 2295 8235
rect 2235 8165 2295 8195
rect 2235 8125 2245 8165
rect 2285 8125 2295 8165
rect 2235 8100 2295 8125
rect 2235 8060 2245 8100
rect 2285 8060 2295 8100
rect 2235 8040 2295 8060
rect 2235 8000 2245 8040
rect 2285 8000 2295 8040
rect 2235 7975 2295 8000
rect 2235 7935 2245 7975
rect 2285 7935 2295 7975
rect 2235 7905 2295 7935
rect 2235 7865 2245 7905
rect 2285 7865 2295 7905
rect 2235 7835 2295 7865
rect 2235 7795 2245 7835
rect 2285 7795 2295 7835
rect 2235 7765 2295 7795
rect 2235 7725 2245 7765
rect 2285 7725 2295 7765
rect 2235 7700 2295 7725
rect 2235 7660 2245 7700
rect 2285 7660 2295 7700
rect 2235 7640 2295 7660
rect 2235 7600 2245 7640
rect 2285 7600 2295 7640
rect 2235 7575 2295 7600
rect 2235 7535 2245 7575
rect 2285 7535 2295 7575
rect 2235 7505 2295 7535
rect 2235 7465 2245 7505
rect 2285 7465 2295 7505
rect 2235 7435 2295 7465
rect 2235 7395 2245 7435
rect 2285 7395 2295 7435
rect 2235 7365 2295 7395
rect 2235 7325 2245 7365
rect 2285 7325 2295 7365
rect 2235 7300 2295 7325
rect 2235 7260 2245 7300
rect 2285 7260 2295 7300
rect 2235 7240 2295 7260
rect 2235 7200 2245 7240
rect 2285 7200 2295 7240
rect 2235 7175 2295 7200
rect 2235 7135 2245 7175
rect 2285 7135 2295 7175
rect 2235 7105 2295 7135
rect 2235 7065 2245 7105
rect 2285 7065 2295 7105
rect 2235 7035 2295 7065
rect 2235 6995 2245 7035
rect 2285 6995 2295 7035
rect 2235 6965 2295 6995
rect 2235 6925 2245 6965
rect 2285 6925 2295 6965
rect 2235 6900 2295 6925
rect 2235 6860 2245 6900
rect 2285 6860 2295 6900
rect 2235 6840 2295 6860
rect 2235 6800 2245 6840
rect 2285 6800 2295 6840
rect 2235 6775 2295 6800
rect 2235 6735 2245 6775
rect 2285 6735 2295 6775
rect 2235 6705 2295 6735
rect 2235 6665 2245 6705
rect 2285 6665 2295 6705
rect 2235 6635 2295 6665
rect 2235 6595 2245 6635
rect 2285 6595 2295 6635
rect 2235 6565 2295 6595
rect 2235 6525 2245 6565
rect 2285 6525 2295 6565
rect 2235 6500 2295 6525
rect 2235 6460 2245 6500
rect 2285 6460 2295 6500
rect 2235 6450 2295 6460
rect 3165 9640 3280 9650
rect 3165 9600 3175 9640
rect 3215 9600 3235 9640
rect 3275 9600 3280 9640
rect 3165 9575 3280 9600
rect 3165 9535 3175 9575
rect 3215 9535 3235 9575
rect 3275 9535 3280 9575
rect 3165 9505 3280 9535
rect 3165 9465 3175 9505
rect 3215 9465 3235 9505
rect 3275 9465 3280 9505
rect 3165 9435 3280 9465
rect 3165 9395 3175 9435
rect 3215 9395 3235 9435
rect 3275 9395 3280 9435
rect 3165 9365 3280 9395
rect 3165 9325 3175 9365
rect 3215 9325 3235 9365
rect 3275 9325 3280 9365
rect 3165 9300 3280 9325
rect 3165 9260 3175 9300
rect 3215 9260 3235 9300
rect 3275 9260 3280 9300
rect 3165 9240 3280 9260
rect 3165 9200 3175 9240
rect 3215 9200 3235 9240
rect 3275 9200 3280 9240
rect 3165 9175 3280 9200
rect 3165 9135 3175 9175
rect 3215 9135 3235 9175
rect 3275 9135 3280 9175
rect 3165 9105 3280 9135
rect 3165 9065 3175 9105
rect 3215 9065 3235 9105
rect 3275 9065 3280 9105
rect 3165 9035 3280 9065
rect 3165 8995 3175 9035
rect 3215 8995 3235 9035
rect 3275 8995 3280 9035
rect 3165 8965 3280 8995
rect 3165 8925 3175 8965
rect 3215 8925 3235 8965
rect 3275 8925 3280 8965
rect 3165 8900 3280 8925
rect 3165 8860 3175 8900
rect 3215 8860 3235 8900
rect 3275 8860 3280 8900
rect 3165 8840 3280 8860
rect 3165 8800 3175 8840
rect 3215 8800 3235 8840
rect 3275 8800 3280 8840
rect 3165 8775 3280 8800
rect 3165 8735 3175 8775
rect 3215 8735 3235 8775
rect 3275 8735 3280 8775
rect 3165 8705 3280 8735
rect 3165 8665 3175 8705
rect 3215 8665 3235 8705
rect 3275 8665 3280 8705
rect 3165 8635 3280 8665
rect 3165 8595 3175 8635
rect 3215 8595 3235 8635
rect 3275 8595 3280 8635
rect 3165 8565 3280 8595
rect 3165 8525 3175 8565
rect 3215 8525 3235 8565
rect 3275 8525 3280 8565
rect 3165 8500 3280 8525
rect 3165 8460 3175 8500
rect 3215 8460 3235 8500
rect 3275 8460 3280 8500
rect 3165 8440 3280 8460
rect 3165 8400 3175 8440
rect 3215 8400 3235 8440
rect 3275 8400 3280 8440
rect 3165 8375 3280 8400
rect 3165 8335 3175 8375
rect 3215 8335 3235 8375
rect 3275 8335 3280 8375
rect 3165 8305 3280 8335
rect 3165 8265 3175 8305
rect 3215 8265 3235 8305
rect 3275 8265 3280 8305
rect 3165 8235 3280 8265
rect 3165 8195 3175 8235
rect 3215 8195 3235 8235
rect 3275 8195 3280 8235
rect 3165 8165 3280 8195
rect 3165 8125 3175 8165
rect 3215 8125 3235 8165
rect 3275 8125 3280 8165
rect 3165 8100 3280 8125
rect 3165 8060 3175 8100
rect 3215 8060 3235 8100
rect 3275 8060 3280 8100
rect 3165 8040 3280 8060
rect 3165 8000 3175 8040
rect 3215 8000 3235 8040
rect 3275 8000 3280 8040
rect 3165 7975 3280 8000
rect 3165 7935 3175 7975
rect 3215 7935 3235 7975
rect 3275 7935 3280 7975
rect 3165 7905 3280 7935
rect 3165 7865 3175 7905
rect 3215 7865 3235 7905
rect 3275 7865 3280 7905
rect 3165 7835 3280 7865
rect 3165 7795 3175 7835
rect 3215 7795 3235 7835
rect 3275 7795 3280 7835
rect 3165 7765 3280 7795
rect 3165 7725 3175 7765
rect 3215 7725 3235 7765
rect 3275 7725 3280 7765
rect 3165 7700 3280 7725
rect 3165 7660 3175 7700
rect 3215 7660 3235 7700
rect 3275 7660 3280 7700
rect 3165 7640 3280 7660
rect 3165 7600 3175 7640
rect 3215 7600 3235 7640
rect 3275 7600 3280 7640
rect 3165 7575 3280 7600
rect 3165 7535 3175 7575
rect 3215 7535 3235 7575
rect 3275 7535 3280 7575
rect 3165 7505 3280 7535
rect 3165 7465 3175 7505
rect 3215 7465 3235 7505
rect 3275 7465 3280 7505
rect 3165 7435 3280 7465
rect 3165 7395 3175 7435
rect 3215 7395 3235 7435
rect 3275 7395 3280 7435
rect 3165 7365 3280 7395
rect 3165 7325 3175 7365
rect 3215 7325 3235 7365
rect 3275 7325 3280 7365
rect 3165 7300 3280 7325
rect 3165 7260 3175 7300
rect 3215 7260 3235 7300
rect 3275 7260 3280 7300
rect 3165 7240 3280 7260
rect 3165 7200 3175 7240
rect 3215 7200 3235 7240
rect 3275 7200 3280 7240
rect 3165 7175 3280 7200
rect 3165 7135 3175 7175
rect 3215 7135 3235 7175
rect 3275 7135 3280 7175
rect 3165 7105 3280 7135
rect 3165 7065 3175 7105
rect 3215 7065 3235 7105
rect 3275 7065 3280 7105
rect 3165 7035 3280 7065
rect 3165 6995 3175 7035
rect 3215 6995 3235 7035
rect 3275 6995 3280 7035
rect 3165 6965 3280 6995
rect 3165 6925 3175 6965
rect 3215 6925 3235 6965
rect 3275 6925 3280 6965
rect 3165 6900 3280 6925
rect 3165 6860 3175 6900
rect 3215 6860 3235 6900
rect 3275 6860 3280 6900
rect 3165 6840 3280 6860
rect 3165 6800 3175 6840
rect 3215 6800 3235 6840
rect 3275 6800 3280 6840
rect 3165 6775 3280 6800
rect 3165 6735 3175 6775
rect 3215 6735 3235 6775
rect 3275 6735 3280 6775
rect 3165 6705 3280 6735
rect 3165 6665 3175 6705
rect 3215 6665 3235 6705
rect 3275 6665 3280 6705
rect 3165 6635 3280 6665
rect 3165 6595 3175 6635
rect 3215 6595 3235 6635
rect 3275 6595 3280 6635
rect 3165 6565 3280 6595
rect 3165 6525 3175 6565
rect 3215 6525 3235 6565
rect 3275 6525 3280 6565
rect 3165 6500 3280 6525
rect 3165 6460 3175 6500
rect 3215 6460 3235 6500
rect 3275 6460 3280 6500
rect 3165 6450 3280 6460
rect 3340 9640 3395 9650
rect 3340 9600 3345 9640
rect 3385 9600 3395 9640
rect 3340 9575 3395 9600
rect 3340 9535 3345 9575
rect 3385 9535 3395 9575
rect 3340 9505 3395 9535
rect 3340 9465 3345 9505
rect 3385 9465 3395 9505
rect 3340 9435 3395 9465
rect 3340 9395 3345 9435
rect 3385 9395 3395 9435
rect 3340 9365 3395 9395
rect 3340 9325 3345 9365
rect 3385 9325 3395 9365
rect 3340 9300 3395 9325
rect 3340 9260 3345 9300
rect 3385 9260 3395 9300
rect 3340 9240 3395 9260
rect 3340 9200 3345 9240
rect 3385 9200 3395 9240
rect 3340 9175 3395 9200
rect 3340 9135 3345 9175
rect 3385 9135 3395 9175
rect 3340 9105 3395 9135
rect 3340 9065 3345 9105
rect 3385 9065 3395 9105
rect 3340 9035 3395 9065
rect 3340 8995 3345 9035
rect 3385 8995 3395 9035
rect 3340 8965 3395 8995
rect 3340 8925 3345 8965
rect 3385 8925 3395 8965
rect 3340 8900 3395 8925
rect 3340 8860 3345 8900
rect 3385 8860 3395 8900
rect 3340 8840 3395 8860
rect 3340 8800 3345 8840
rect 3385 8800 3395 8840
rect 3340 8775 3395 8800
rect 3340 8735 3345 8775
rect 3385 8735 3395 8775
rect 3340 8705 3395 8735
rect 3340 8665 3345 8705
rect 3385 8665 3395 8705
rect 3340 8635 3395 8665
rect 3340 8595 3345 8635
rect 3385 8595 3395 8635
rect 3340 8565 3395 8595
rect 3340 8525 3345 8565
rect 3385 8525 3395 8565
rect 3340 8500 3395 8525
rect 3340 8460 3345 8500
rect 3385 8460 3395 8500
rect 3340 8440 3395 8460
rect 3340 8400 3345 8440
rect 3385 8400 3395 8440
rect 3340 8375 3395 8400
rect 3340 8335 3345 8375
rect 3385 8335 3395 8375
rect 3340 8305 3395 8335
rect 3340 8265 3345 8305
rect 3385 8265 3395 8305
rect 3340 8235 3395 8265
rect 3340 8195 3345 8235
rect 3385 8195 3395 8235
rect 3340 8165 3395 8195
rect 3340 8125 3345 8165
rect 3385 8125 3395 8165
rect 3340 8100 3395 8125
rect 3340 8060 3345 8100
rect 3385 8060 3395 8100
rect 3340 8040 3395 8060
rect 3340 8000 3345 8040
rect 3385 8000 3395 8040
rect 3340 7975 3395 8000
rect 3340 7935 3345 7975
rect 3385 7935 3395 7975
rect 3340 7905 3395 7935
rect 3340 7865 3345 7905
rect 3385 7865 3395 7905
rect 3340 7835 3395 7865
rect 3340 7795 3345 7835
rect 3385 7795 3395 7835
rect 3340 7765 3395 7795
rect 3340 7725 3345 7765
rect 3385 7725 3395 7765
rect 3340 7700 3395 7725
rect 3340 7660 3345 7700
rect 3385 7660 3395 7700
rect 3340 7640 3395 7660
rect 3340 7600 3345 7640
rect 3385 7600 3395 7640
rect 3340 7575 3395 7600
rect 3340 7535 3345 7575
rect 3385 7535 3395 7575
rect 3340 7505 3395 7535
rect 3340 7465 3345 7505
rect 3385 7465 3395 7505
rect 3340 7435 3395 7465
rect 3340 7395 3345 7435
rect 3385 7395 3395 7435
rect 3340 7365 3395 7395
rect 3340 7325 3345 7365
rect 3385 7325 3395 7365
rect 3340 7300 3395 7325
rect 3340 7260 3345 7300
rect 3385 7260 3395 7300
rect 3340 7240 3395 7260
rect 3340 7200 3345 7240
rect 3385 7200 3395 7240
rect 3340 7175 3395 7200
rect 3340 7135 3345 7175
rect 3385 7135 3395 7175
rect 3340 7105 3395 7135
rect 3340 7065 3345 7105
rect 3385 7065 3395 7105
rect 3340 7035 3395 7065
rect 3340 6995 3345 7035
rect 3385 6995 3395 7035
rect 3340 6965 3395 6995
rect 3340 6925 3345 6965
rect 3385 6925 3395 6965
rect 3340 6900 3395 6925
rect 3340 6860 3345 6900
rect 3385 6860 3395 6900
rect 3340 6840 3395 6860
rect 3340 6800 3345 6840
rect 3385 6800 3395 6840
rect 3340 6775 3395 6800
rect 3340 6735 3345 6775
rect 3385 6735 3395 6775
rect 3340 6705 3395 6735
rect 3340 6665 3345 6705
rect 3385 6665 3395 6705
rect 3340 6635 3395 6665
rect 3340 6595 3345 6635
rect 3385 6595 3395 6635
rect 3340 6565 3395 6595
rect 3340 6525 3345 6565
rect 3385 6525 3395 6565
rect 3340 6500 3395 6525
rect 3340 6460 3345 6500
rect 3385 6460 3395 6500
rect 3340 6450 3395 6460
rect 6690 9640 6750 9650
rect 6690 9600 6700 9640
rect 6740 9600 6750 9640
rect 6690 9575 6750 9600
rect 6690 9535 6700 9575
rect 6740 9535 6750 9575
rect 6690 9505 6750 9535
rect 6690 9465 6700 9505
rect 6740 9465 6750 9505
rect 6690 9435 6750 9465
rect 6690 9395 6700 9435
rect 6740 9395 6750 9435
rect 6690 9365 6750 9395
rect 6690 9325 6700 9365
rect 6740 9325 6750 9365
rect 6690 9300 6750 9325
rect 6690 9260 6700 9300
rect 6740 9260 6750 9300
rect 6690 9240 6750 9260
rect 6690 9200 6700 9240
rect 6740 9200 6750 9240
rect 6690 9175 6750 9200
rect 6690 9135 6700 9175
rect 6740 9135 6750 9175
rect 6690 9105 6750 9135
rect 6690 9065 6700 9105
rect 6740 9065 6750 9105
rect 6690 9035 6750 9065
rect 6690 8995 6700 9035
rect 6740 8995 6750 9035
rect 6690 8965 6750 8995
rect 6690 8925 6700 8965
rect 6740 8925 6750 8965
rect 6690 8900 6750 8925
rect 6690 8860 6700 8900
rect 6740 8860 6750 8900
rect 6690 8840 6750 8860
rect 6690 8800 6700 8840
rect 6740 8800 6750 8840
rect 6690 8775 6750 8800
rect 6690 8735 6700 8775
rect 6740 8735 6750 8775
rect 6690 8705 6750 8735
rect 6690 8665 6700 8705
rect 6740 8665 6750 8705
rect 6690 8635 6750 8665
rect 6690 8595 6700 8635
rect 6740 8595 6750 8635
rect 6690 8565 6750 8595
rect 6690 8525 6700 8565
rect 6740 8525 6750 8565
rect 6690 8500 6750 8525
rect 6690 8460 6700 8500
rect 6740 8460 6750 8500
rect 6690 8440 6750 8460
rect 6690 8400 6700 8440
rect 6740 8400 6750 8440
rect 6690 8375 6750 8400
rect 6690 8335 6700 8375
rect 6740 8335 6750 8375
rect 6690 8305 6750 8335
rect 6690 8265 6700 8305
rect 6740 8265 6750 8305
rect 6690 8235 6750 8265
rect 6690 8195 6700 8235
rect 6740 8195 6750 8235
rect 6690 8165 6750 8195
rect 6690 8125 6700 8165
rect 6740 8125 6750 8165
rect 6690 8100 6750 8125
rect 6690 8060 6700 8100
rect 6740 8060 6750 8100
rect 6690 8040 6750 8060
rect 6690 8000 6700 8040
rect 6740 8000 6750 8040
rect 6690 7975 6750 8000
rect 6690 7935 6700 7975
rect 6740 7935 6750 7975
rect 6690 7905 6750 7935
rect 6690 7865 6700 7905
rect 6740 7865 6750 7905
rect 6690 7835 6750 7865
rect 6690 7795 6700 7835
rect 6740 7795 6750 7835
rect 6690 7765 6750 7795
rect 6690 7725 6700 7765
rect 6740 7725 6750 7765
rect 6690 7700 6750 7725
rect 6690 7660 6700 7700
rect 6740 7660 6750 7700
rect 6690 7640 6750 7660
rect 6690 7600 6700 7640
rect 6740 7600 6750 7640
rect 6690 7575 6750 7600
rect 6690 7535 6700 7575
rect 6740 7535 6750 7575
rect 6690 7505 6750 7535
rect 6690 7465 6700 7505
rect 6740 7465 6750 7505
rect 6690 7435 6750 7465
rect 6690 7395 6700 7435
rect 6740 7395 6750 7435
rect 6690 7365 6750 7395
rect 6690 7325 6700 7365
rect 6740 7325 6750 7365
rect 6690 7300 6750 7325
rect 6690 7260 6700 7300
rect 6740 7260 6750 7300
rect 6690 7240 6750 7260
rect 6690 7200 6700 7240
rect 6740 7200 6750 7240
rect 6690 7175 6750 7200
rect 6690 7135 6700 7175
rect 6740 7135 6750 7175
rect 6690 7105 6750 7135
rect 6690 7065 6700 7105
rect 6740 7065 6750 7105
rect 6690 7035 6750 7065
rect 6690 6995 6700 7035
rect 6740 6995 6750 7035
rect 6690 6965 6750 6995
rect 6690 6925 6700 6965
rect 6740 6925 6750 6965
rect 6690 6900 6750 6925
rect 6690 6860 6700 6900
rect 6740 6860 6750 6900
rect 6690 6840 6750 6860
rect 6690 6800 6700 6840
rect 6740 6800 6750 6840
rect 6690 6775 6750 6800
rect 6690 6735 6700 6775
rect 6740 6735 6750 6775
rect 6690 6705 6750 6735
rect 6690 6665 6700 6705
rect 6740 6665 6750 6705
rect 6690 6635 6750 6665
rect 6690 6595 6700 6635
rect 6740 6595 6750 6635
rect 6690 6565 6750 6595
rect 6690 6525 6700 6565
rect 6740 6525 6750 6565
rect 6690 6500 6750 6525
rect 6690 6460 6700 6500
rect 6740 6460 6750 6500
rect 6690 6450 6750 6460
rect 7260 9640 7320 9650
rect 7260 9600 7270 9640
rect 7310 9600 7320 9640
rect 7260 9575 7320 9600
rect 7260 9535 7270 9575
rect 7310 9535 7320 9575
rect 7260 9505 7320 9535
rect 7260 9465 7270 9505
rect 7310 9465 7320 9505
rect 7260 9435 7320 9465
rect 7260 9395 7270 9435
rect 7310 9395 7320 9435
rect 7260 9365 7320 9395
rect 7260 9325 7270 9365
rect 7310 9325 7320 9365
rect 7260 9300 7320 9325
rect 7260 9260 7270 9300
rect 7310 9260 7320 9300
rect 7260 9240 7320 9260
rect 7260 9200 7270 9240
rect 7310 9200 7320 9240
rect 7260 9175 7320 9200
rect 7260 9135 7270 9175
rect 7310 9135 7320 9175
rect 7260 9105 7320 9135
rect 7260 9065 7270 9105
rect 7310 9065 7320 9105
rect 7260 9035 7320 9065
rect 7260 8995 7270 9035
rect 7310 8995 7320 9035
rect 7260 8965 7320 8995
rect 7260 8925 7270 8965
rect 7310 8925 7320 8965
rect 7260 8900 7320 8925
rect 7260 8860 7270 8900
rect 7310 8860 7320 8900
rect 7260 8840 7320 8860
rect 7260 8800 7270 8840
rect 7310 8800 7320 8840
rect 7260 8775 7320 8800
rect 7260 8735 7270 8775
rect 7310 8735 7320 8775
rect 7260 8705 7320 8735
rect 7260 8665 7270 8705
rect 7310 8665 7320 8705
rect 7260 8635 7320 8665
rect 7260 8595 7270 8635
rect 7310 8595 7320 8635
rect 7260 8565 7320 8595
rect 7260 8525 7270 8565
rect 7310 8525 7320 8565
rect 7260 8500 7320 8525
rect 7260 8460 7270 8500
rect 7310 8460 7320 8500
rect 7260 8440 7320 8460
rect 7260 8400 7270 8440
rect 7310 8400 7320 8440
rect 7260 8375 7320 8400
rect 7260 8335 7270 8375
rect 7310 8335 7320 8375
rect 7260 8305 7320 8335
rect 7260 8265 7270 8305
rect 7310 8265 7320 8305
rect 7260 8235 7320 8265
rect 7260 8195 7270 8235
rect 7310 8195 7320 8235
rect 7260 8165 7320 8195
rect 7260 8125 7270 8165
rect 7310 8125 7320 8165
rect 7260 8100 7320 8125
rect 7260 8060 7270 8100
rect 7310 8060 7320 8100
rect 7260 8040 7320 8060
rect 7260 8000 7270 8040
rect 7310 8000 7320 8040
rect 7260 7975 7320 8000
rect 7260 7935 7270 7975
rect 7310 7935 7320 7975
rect 7260 7905 7320 7935
rect 7260 7865 7270 7905
rect 7310 7865 7320 7905
rect 7260 7835 7320 7865
rect 7260 7795 7270 7835
rect 7310 7795 7320 7835
rect 7260 7765 7320 7795
rect 7260 7725 7270 7765
rect 7310 7725 7320 7765
rect 7260 7700 7320 7725
rect 7260 7660 7270 7700
rect 7310 7660 7320 7700
rect 7260 7640 7320 7660
rect 7260 7600 7270 7640
rect 7310 7600 7320 7640
rect 7260 7575 7320 7600
rect 7260 7535 7270 7575
rect 7310 7535 7320 7575
rect 7260 7505 7320 7535
rect 7260 7465 7270 7505
rect 7310 7465 7320 7505
rect 7260 7435 7320 7465
rect 7260 7395 7270 7435
rect 7310 7395 7320 7435
rect 7260 7365 7320 7395
rect 7260 7325 7270 7365
rect 7310 7325 7320 7365
rect 7260 7300 7320 7325
rect 7260 7260 7270 7300
rect 7310 7260 7320 7300
rect 7260 7240 7320 7260
rect 7260 7200 7270 7240
rect 7310 7200 7320 7240
rect 7260 7175 7320 7200
rect 7260 7135 7270 7175
rect 7310 7135 7320 7175
rect 7260 7105 7320 7135
rect 7260 7065 7270 7105
rect 7310 7065 7320 7105
rect 7260 7035 7320 7065
rect 7260 6995 7270 7035
rect 7310 6995 7320 7035
rect 7260 6965 7320 6995
rect 7260 6925 7270 6965
rect 7310 6925 7320 6965
rect 7260 6900 7320 6925
rect 7260 6860 7270 6900
rect 7310 6860 7320 6900
rect 7260 6840 7320 6860
rect 7260 6800 7270 6840
rect 7310 6800 7320 6840
rect 7260 6775 7320 6800
rect 7260 6735 7270 6775
rect 7310 6735 7320 6775
rect 7260 6705 7320 6735
rect 7260 6665 7270 6705
rect 7310 6665 7320 6705
rect 7260 6635 7320 6665
rect 7260 6595 7270 6635
rect 7310 6595 7320 6635
rect 7260 6565 7320 6595
rect 7260 6525 7270 6565
rect 7310 6525 7320 6565
rect 7260 6500 7320 6525
rect 7260 6460 7270 6500
rect 7310 6460 7320 6500
rect 7260 6450 7320 6460
rect 7960 9640 8020 9650
rect 7960 9600 7970 9640
rect 8010 9600 8020 9640
rect 7960 9575 8020 9600
rect 7960 9535 7970 9575
rect 8010 9535 8020 9575
rect 7960 9505 8020 9535
rect 7960 9465 7970 9505
rect 8010 9465 8020 9505
rect 7960 9435 8020 9465
rect 7960 9395 7970 9435
rect 8010 9395 8020 9435
rect 7960 9365 8020 9395
rect 7960 9325 7970 9365
rect 8010 9325 8020 9365
rect 7960 9300 8020 9325
rect 7960 9260 7970 9300
rect 8010 9260 8020 9300
rect 7960 9240 8020 9260
rect 7960 9200 7970 9240
rect 8010 9200 8020 9240
rect 7960 9175 8020 9200
rect 7960 9135 7970 9175
rect 8010 9135 8020 9175
rect 7960 9105 8020 9135
rect 7960 9065 7970 9105
rect 8010 9065 8020 9105
rect 7960 9035 8020 9065
rect 7960 8995 7970 9035
rect 8010 8995 8020 9035
rect 7960 8965 8020 8995
rect 7960 8925 7970 8965
rect 8010 8925 8020 8965
rect 7960 8900 8020 8925
rect 7960 8860 7970 8900
rect 8010 8860 8020 8900
rect 7960 8840 8020 8860
rect 7960 8800 7970 8840
rect 8010 8800 8020 8840
rect 7960 8775 8020 8800
rect 7960 8735 7970 8775
rect 8010 8735 8020 8775
rect 7960 8705 8020 8735
rect 7960 8665 7970 8705
rect 8010 8665 8020 8705
rect 7960 8635 8020 8665
rect 7960 8595 7970 8635
rect 8010 8595 8020 8635
rect 7960 8565 8020 8595
rect 7960 8525 7970 8565
rect 8010 8525 8020 8565
rect 7960 8500 8020 8525
rect 7960 8460 7970 8500
rect 8010 8460 8020 8500
rect 7960 8440 8020 8460
rect 7960 8400 7970 8440
rect 8010 8400 8020 8440
rect 7960 8375 8020 8400
rect 7960 8335 7970 8375
rect 8010 8335 8020 8375
rect 7960 8305 8020 8335
rect 7960 8265 7970 8305
rect 8010 8265 8020 8305
rect 7960 8235 8020 8265
rect 7960 8195 7970 8235
rect 8010 8195 8020 8235
rect 7960 8165 8020 8195
rect 7960 8125 7970 8165
rect 8010 8125 8020 8165
rect 7960 8100 8020 8125
rect 7960 8060 7970 8100
rect 8010 8060 8020 8100
rect 7960 8040 8020 8060
rect 7960 8000 7970 8040
rect 8010 8000 8020 8040
rect 7960 7975 8020 8000
rect 7960 7935 7970 7975
rect 8010 7935 8020 7975
rect 7960 7905 8020 7935
rect 7960 7865 7970 7905
rect 8010 7865 8020 7905
rect 7960 7835 8020 7865
rect 7960 7795 7970 7835
rect 8010 7795 8020 7835
rect 7960 7765 8020 7795
rect 7960 7725 7970 7765
rect 8010 7725 8020 7765
rect 7960 7700 8020 7725
rect 7960 7660 7970 7700
rect 8010 7660 8020 7700
rect 7960 7640 8020 7660
rect 7960 7600 7970 7640
rect 8010 7600 8020 7640
rect 7960 7575 8020 7600
rect 7960 7535 7970 7575
rect 8010 7535 8020 7575
rect 7960 7505 8020 7535
rect 7960 7465 7970 7505
rect 8010 7465 8020 7505
rect 7960 7435 8020 7465
rect 7960 7395 7970 7435
rect 8010 7395 8020 7435
rect 7960 7365 8020 7395
rect 7960 7325 7970 7365
rect 8010 7325 8020 7365
rect 7960 7300 8020 7325
rect 7960 7260 7970 7300
rect 8010 7260 8020 7300
rect 7960 7240 8020 7260
rect 7960 7200 7970 7240
rect 8010 7200 8020 7240
rect 7960 7175 8020 7200
rect 7960 7135 7970 7175
rect 8010 7135 8020 7175
rect 7960 7105 8020 7135
rect 7960 7065 7970 7105
rect 8010 7065 8020 7105
rect 7960 7035 8020 7065
rect 7960 6995 7970 7035
rect 8010 6995 8020 7035
rect 7960 6965 8020 6995
rect 7960 6925 7970 6965
rect 8010 6925 8020 6965
rect 7960 6900 8020 6925
rect 7960 6860 7970 6900
rect 8010 6860 8020 6900
rect 7960 6840 8020 6860
rect 7960 6800 7970 6840
rect 8010 6800 8020 6840
rect 7960 6775 8020 6800
rect 7960 6735 7970 6775
rect 8010 6735 8020 6775
rect 7960 6705 8020 6735
rect 7960 6665 7970 6705
rect 8010 6665 8020 6705
rect 7960 6635 8020 6665
rect 7960 6595 7970 6635
rect 8010 6595 8020 6635
rect 7960 6565 8020 6595
rect 7960 6525 7970 6565
rect 8010 6525 8020 6565
rect 7960 6500 8020 6525
rect 7960 6460 7970 6500
rect 8010 6460 8020 6500
rect 7960 6450 8020 6460
rect 8310 9640 8370 9650
rect 8310 9600 8320 9640
rect 8360 9600 8370 9640
rect 8310 9575 8370 9600
rect 8310 9535 8320 9575
rect 8360 9535 8370 9575
rect 8310 9505 8370 9535
rect 8310 9465 8320 9505
rect 8360 9465 8370 9505
rect 8310 9435 8370 9465
rect 8310 9395 8320 9435
rect 8360 9395 8370 9435
rect 8310 9365 8370 9395
rect 8310 9325 8320 9365
rect 8360 9325 8370 9365
rect 8310 9300 8370 9325
rect 8310 9260 8320 9300
rect 8360 9260 8370 9300
rect 8310 9240 8370 9260
rect 8310 9200 8320 9240
rect 8360 9200 8370 9240
rect 8310 9175 8370 9200
rect 8310 9135 8320 9175
rect 8360 9135 8370 9175
rect 8310 9105 8370 9135
rect 8310 9065 8320 9105
rect 8360 9065 8370 9105
rect 8310 9035 8370 9065
rect 8310 8995 8320 9035
rect 8360 8995 8370 9035
rect 8310 8965 8370 8995
rect 8310 8925 8320 8965
rect 8360 8925 8370 8965
rect 8310 8900 8370 8925
rect 8310 8860 8320 8900
rect 8360 8860 8370 8900
rect 8310 8840 8370 8860
rect 8310 8800 8320 8840
rect 8360 8800 8370 8840
rect 8310 8775 8370 8800
rect 8310 8735 8320 8775
rect 8360 8735 8370 8775
rect 8310 8705 8370 8735
rect 8310 8665 8320 8705
rect 8360 8665 8370 8705
rect 8310 8635 8370 8665
rect 8310 8595 8320 8635
rect 8360 8595 8370 8635
rect 8310 8565 8370 8595
rect 8310 8525 8320 8565
rect 8360 8525 8370 8565
rect 8310 8500 8370 8525
rect 8310 8460 8320 8500
rect 8360 8460 8370 8500
rect 8310 8440 8370 8460
rect 8310 8400 8320 8440
rect 8360 8400 8370 8440
rect 8310 8375 8370 8400
rect 8310 8335 8320 8375
rect 8360 8335 8370 8375
rect 8310 8305 8370 8335
rect 8310 8265 8320 8305
rect 8360 8265 8370 8305
rect 8310 8235 8370 8265
rect 8310 8195 8320 8235
rect 8360 8195 8370 8235
rect 8310 8165 8370 8195
rect 8310 8125 8320 8165
rect 8360 8125 8370 8165
rect 8310 8100 8370 8125
rect 8310 8060 8320 8100
rect 8360 8060 8370 8100
rect 8310 8040 8370 8060
rect 8310 8000 8320 8040
rect 8360 8000 8370 8040
rect 8310 7975 8370 8000
rect 8310 7935 8320 7975
rect 8360 7935 8370 7975
rect 8310 7905 8370 7935
rect 8310 7865 8320 7905
rect 8360 7865 8370 7905
rect 8310 7835 8370 7865
rect 8310 7795 8320 7835
rect 8360 7795 8370 7835
rect 8310 7765 8370 7795
rect 8310 7725 8320 7765
rect 8360 7725 8370 7765
rect 8310 7700 8370 7725
rect 8310 7660 8320 7700
rect 8360 7660 8370 7700
rect 8310 7640 8370 7660
rect 8310 7600 8320 7640
rect 8360 7600 8370 7640
rect 8310 7575 8370 7600
rect 8310 7535 8320 7575
rect 8360 7535 8370 7575
rect 8310 7505 8370 7535
rect 8310 7465 8320 7505
rect 8360 7465 8370 7505
rect 8310 7435 8370 7465
rect 8310 7395 8320 7435
rect 8360 7395 8370 7435
rect 8310 7365 8370 7395
rect 8310 7325 8320 7365
rect 8360 7325 8370 7365
rect 8310 7300 8370 7325
rect 8310 7260 8320 7300
rect 8360 7260 8370 7300
rect 8310 7240 8370 7260
rect 8310 7200 8320 7240
rect 8360 7200 8370 7240
rect 8310 7175 8370 7200
rect 8310 7135 8320 7175
rect 8360 7135 8370 7175
rect 8310 7105 8370 7135
rect 8310 7065 8320 7105
rect 8360 7065 8370 7105
rect 8310 7035 8370 7065
rect 8310 6995 8320 7035
rect 8360 6995 8370 7035
rect 8310 6965 8370 6995
rect 8310 6925 8320 6965
rect 8360 6925 8370 6965
rect 8310 6900 8370 6925
rect 8310 6860 8320 6900
rect 8360 6860 8370 6900
rect 8310 6840 8370 6860
rect 8310 6800 8320 6840
rect 8360 6800 8370 6840
rect 8310 6775 8370 6800
rect 8310 6735 8320 6775
rect 8360 6735 8370 6775
rect 8310 6705 8370 6735
rect 8310 6665 8320 6705
rect 8360 6665 8370 6705
rect 8310 6635 8370 6665
rect 8310 6595 8320 6635
rect 8360 6595 8370 6635
rect 8310 6565 8370 6595
rect 8310 6525 8320 6565
rect 8360 6525 8370 6565
rect 8310 6500 8370 6525
rect 8310 6460 8320 6500
rect 8360 6460 8370 6500
rect 8310 6450 8370 6460
rect 8660 9640 8720 9650
rect 8660 9600 8670 9640
rect 8710 9600 8720 9640
rect 8660 9575 8720 9600
rect 8660 9535 8670 9575
rect 8710 9535 8720 9575
rect 8660 9505 8720 9535
rect 8660 9465 8670 9505
rect 8710 9465 8720 9505
rect 8660 9435 8720 9465
rect 8660 9395 8670 9435
rect 8710 9395 8720 9435
rect 8660 9365 8720 9395
rect 8660 9325 8670 9365
rect 8710 9325 8720 9365
rect 8660 9300 8720 9325
rect 8660 9260 8670 9300
rect 8710 9260 8720 9300
rect 8660 9240 8720 9260
rect 8660 9200 8670 9240
rect 8710 9200 8720 9240
rect 8660 9175 8720 9200
rect 8660 9135 8670 9175
rect 8710 9135 8720 9175
rect 8660 9105 8720 9135
rect 8660 9065 8670 9105
rect 8710 9065 8720 9105
rect 8660 9035 8720 9065
rect 8660 8995 8670 9035
rect 8710 8995 8720 9035
rect 8660 8965 8720 8995
rect 8660 8925 8670 8965
rect 8710 8925 8720 8965
rect 8660 8900 8720 8925
rect 8660 8860 8670 8900
rect 8710 8860 8720 8900
rect 8660 8840 8720 8860
rect 8660 8800 8670 8840
rect 8710 8800 8720 8840
rect 8660 8775 8720 8800
rect 8660 8735 8670 8775
rect 8710 8735 8720 8775
rect 8660 8705 8720 8735
rect 8660 8665 8670 8705
rect 8710 8665 8720 8705
rect 8660 8635 8720 8665
rect 8660 8595 8670 8635
rect 8710 8595 8720 8635
rect 8660 8565 8720 8595
rect 8660 8525 8670 8565
rect 8710 8525 8720 8565
rect 8660 8500 8720 8525
rect 8660 8460 8670 8500
rect 8710 8460 8720 8500
rect 8660 8440 8720 8460
rect 8660 8400 8670 8440
rect 8710 8400 8720 8440
rect 8660 8375 8720 8400
rect 8660 8335 8670 8375
rect 8710 8335 8720 8375
rect 8660 8305 8720 8335
rect 8660 8265 8670 8305
rect 8710 8265 8720 8305
rect 8660 8235 8720 8265
rect 8660 8195 8670 8235
rect 8710 8195 8720 8235
rect 8660 8165 8720 8195
rect 8660 8125 8670 8165
rect 8710 8125 8720 8165
rect 8660 8100 8720 8125
rect 8660 8060 8670 8100
rect 8710 8060 8720 8100
rect 8660 8040 8720 8060
rect 8660 8000 8670 8040
rect 8710 8000 8720 8040
rect 8660 7975 8720 8000
rect 8660 7935 8670 7975
rect 8710 7935 8720 7975
rect 8660 7905 8720 7935
rect 8660 7865 8670 7905
rect 8710 7865 8720 7905
rect 8660 7835 8720 7865
rect 8660 7795 8670 7835
rect 8710 7795 8720 7835
rect 8660 7765 8720 7795
rect 8660 7725 8670 7765
rect 8710 7725 8720 7765
rect 8660 7700 8720 7725
rect 8660 7660 8670 7700
rect 8710 7660 8720 7700
rect 8660 7640 8720 7660
rect 8660 7600 8670 7640
rect 8710 7600 8720 7640
rect 8660 7575 8720 7600
rect 8660 7535 8670 7575
rect 8710 7535 8720 7575
rect 8660 7505 8720 7535
rect 8660 7465 8670 7505
rect 8710 7465 8720 7505
rect 8660 7435 8720 7465
rect 8660 7395 8670 7435
rect 8710 7395 8720 7435
rect 8660 7365 8720 7395
rect 8660 7325 8670 7365
rect 8710 7325 8720 7365
rect 8660 7300 8720 7325
rect 8660 7260 8670 7300
rect 8710 7260 8720 7300
rect 8660 7240 8720 7260
rect 8660 7200 8670 7240
rect 8710 7200 8720 7240
rect 8660 7175 8720 7200
rect 8660 7135 8670 7175
rect 8710 7135 8720 7175
rect 8660 7105 8720 7135
rect 8660 7065 8670 7105
rect 8710 7065 8720 7105
rect 8660 7035 8720 7065
rect 8660 6995 8670 7035
rect 8710 6995 8720 7035
rect 8660 6965 8720 6995
rect 8660 6925 8670 6965
rect 8710 6925 8720 6965
rect 8660 6900 8720 6925
rect 8660 6860 8670 6900
rect 8710 6860 8720 6900
rect 8660 6840 8720 6860
rect 8660 6800 8670 6840
rect 8710 6800 8720 6840
rect 8660 6775 8720 6800
rect 8660 6735 8670 6775
rect 8710 6735 8720 6775
rect 8660 6705 8720 6735
rect 8660 6665 8670 6705
rect 8710 6665 8720 6705
rect 8660 6635 8720 6665
rect 8660 6595 8670 6635
rect 8710 6595 8720 6635
rect 8660 6565 8720 6595
rect 8660 6525 8670 6565
rect 8710 6525 8720 6565
rect 8660 6500 8720 6525
rect 8660 6460 8670 6500
rect 8710 6460 8720 6500
rect 8660 6450 8720 6460
rect 9010 9640 9070 9650
rect 9010 9600 9020 9640
rect 9060 9600 9070 9640
rect 9010 9575 9070 9600
rect 9010 9535 9020 9575
rect 9060 9535 9070 9575
rect 9010 9505 9070 9535
rect 9010 9465 9020 9505
rect 9060 9465 9070 9505
rect 9010 9435 9070 9465
rect 9010 9395 9020 9435
rect 9060 9395 9070 9435
rect 9010 9365 9070 9395
rect 9010 9325 9020 9365
rect 9060 9325 9070 9365
rect 9010 9300 9070 9325
rect 9010 9260 9020 9300
rect 9060 9260 9070 9300
rect 9010 9240 9070 9260
rect 9010 9200 9020 9240
rect 9060 9200 9070 9240
rect 9010 9175 9070 9200
rect 9010 9135 9020 9175
rect 9060 9135 9070 9175
rect 9010 9105 9070 9135
rect 9010 9065 9020 9105
rect 9060 9065 9070 9105
rect 9010 9035 9070 9065
rect 9010 8995 9020 9035
rect 9060 8995 9070 9035
rect 9010 8965 9070 8995
rect 9010 8925 9020 8965
rect 9060 8925 9070 8965
rect 9010 8900 9070 8925
rect 9010 8860 9020 8900
rect 9060 8860 9070 8900
rect 9010 8840 9070 8860
rect 9010 8800 9020 8840
rect 9060 8800 9070 8840
rect 9010 8775 9070 8800
rect 9010 8735 9020 8775
rect 9060 8735 9070 8775
rect 9010 8705 9070 8735
rect 9010 8665 9020 8705
rect 9060 8665 9070 8705
rect 9010 8635 9070 8665
rect 9010 8595 9020 8635
rect 9060 8595 9070 8635
rect 9010 8565 9070 8595
rect 9010 8525 9020 8565
rect 9060 8525 9070 8565
rect 9010 8500 9070 8525
rect 9010 8460 9020 8500
rect 9060 8460 9070 8500
rect 9010 8440 9070 8460
rect 9010 8400 9020 8440
rect 9060 8400 9070 8440
rect 9010 8375 9070 8400
rect 9010 8335 9020 8375
rect 9060 8335 9070 8375
rect 9010 8305 9070 8335
rect 9010 8265 9020 8305
rect 9060 8265 9070 8305
rect 9010 8235 9070 8265
rect 9010 8195 9020 8235
rect 9060 8195 9070 8235
rect 9010 8165 9070 8195
rect 9010 8125 9020 8165
rect 9060 8125 9070 8165
rect 9010 8100 9070 8125
rect 9010 8060 9020 8100
rect 9060 8060 9070 8100
rect 9010 8040 9070 8060
rect 9010 8000 9020 8040
rect 9060 8000 9070 8040
rect 9010 7975 9070 8000
rect 9010 7935 9020 7975
rect 9060 7935 9070 7975
rect 9010 7905 9070 7935
rect 9010 7865 9020 7905
rect 9060 7865 9070 7905
rect 9010 7835 9070 7865
rect 9010 7795 9020 7835
rect 9060 7795 9070 7835
rect 9010 7765 9070 7795
rect 9010 7725 9020 7765
rect 9060 7725 9070 7765
rect 9010 7700 9070 7725
rect 9010 7660 9020 7700
rect 9060 7660 9070 7700
rect 9010 7640 9070 7660
rect 9010 7600 9020 7640
rect 9060 7600 9070 7640
rect 9010 7575 9070 7600
rect 9010 7535 9020 7575
rect 9060 7535 9070 7575
rect 9010 7505 9070 7535
rect 9010 7465 9020 7505
rect 9060 7465 9070 7505
rect 9010 7435 9070 7465
rect 9010 7395 9020 7435
rect 9060 7395 9070 7435
rect 9010 7365 9070 7395
rect 9010 7325 9020 7365
rect 9060 7325 9070 7365
rect 9010 7300 9070 7325
rect 9010 7260 9020 7300
rect 9060 7260 9070 7300
rect 9010 7240 9070 7260
rect 9010 7200 9020 7240
rect 9060 7200 9070 7240
rect 9010 7175 9070 7200
rect 9010 7135 9020 7175
rect 9060 7135 9070 7175
rect 9010 7105 9070 7135
rect 9010 7065 9020 7105
rect 9060 7065 9070 7105
rect 9010 7035 9070 7065
rect 9010 6995 9020 7035
rect 9060 6995 9070 7035
rect 9010 6965 9070 6995
rect 9010 6925 9020 6965
rect 9060 6925 9070 6965
rect 9010 6900 9070 6925
rect 9010 6860 9020 6900
rect 9060 6860 9070 6900
rect 9010 6840 9070 6860
rect 9010 6800 9020 6840
rect 9060 6800 9070 6840
rect 9010 6775 9070 6800
rect 9010 6735 9020 6775
rect 9060 6735 9070 6775
rect 9010 6705 9070 6735
rect 9010 6665 9020 6705
rect 9060 6665 9070 6705
rect 9010 6635 9070 6665
rect 9010 6595 9020 6635
rect 9060 6595 9070 6635
rect 9010 6565 9070 6595
rect 9010 6525 9020 6565
rect 9060 6525 9070 6565
rect 9010 6500 9070 6525
rect 9010 6460 9020 6500
rect 9060 6460 9070 6500
rect 9010 6450 9070 6460
rect 31290 8030 32890 17740
rect 31290 7995 31305 8030
rect 31340 7995 31350 8030
rect 31385 7995 31395 8030
rect 31430 7995 31440 8030
rect 31475 7995 31485 8030
rect 31520 7995 31530 8030
rect 31565 7995 31575 8030
rect 31610 7995 31620 8030
rect 31655 7995 31665 8030
rect 31700 7995 31710 8030
rect 31745 7995 31755 8030
rect 31790 7995 31800 8030
rect 31835 7995 31845 8030
rect 31880 7995 31890 8030
rect 31925 7995 31935 8030
rect 31970 7995 31980 8030
rect 32015 7995 32025 8030
rect 32060 7995 32070 8030
rect 32105 7995 32115 8030
rect 32150 7995 32160 8030
rect 32195 7995 32205 8030
rect 32240 7995 32250 8030
rect 32285 7995 32295 8030
rect 32330 7995 32340 8030
rect 32375 7995 32385 8030
rect 32420 7995 32430 8030
rect 32465 7995 32475 8030
rect 32510 7995 32520 8030
rect 32555 7995 32565 8030
rect 32600 7995 32610 8030
rect 32645 7995 32655 8030
rect 32690 7995 32700 8030
rect 32735 7995 32745 8030
rect 32780 7995 32790 8030
rect 32825 7995 32835 8030
rect 32870 7995 32890 8030
rect 31290 7985 32890 7995
rect 31290 7950 31305 7985
rect 31340 7950 31350 7985
rect 31385 7950 31395 7985
rect 31430 7950 31440 7985
rect 31475 7950 31485 7985
rect 31520 7950 31530 7985
rect 31565 7950 31575 7985
rect 31610 7950 31620 7985
rect 31655 7950 31665 7985
rect 31700 7950 31710 7985
rect 31745 7950 31755 7985
rect 31790 7950 31800 7985
rect 31835 7950 31845 7985
rect 31880 7950 31890 7985
rect 31925 7950 31935 7985
rect 31970 7950 31980 7985
rect 32015 7950 32025 7985
rect 32060 7950 32070 7985
rect 32105 7950 32115 7985
rect 32150 7950 32160 7985
rect 32195 7950 32205 7985
rect 32240 7950 32250 7985
rect 32285 7950 32295 7985
rect 32330 7950 32340 7985
rect 32375 7950 32385 7985
rect 32420 7950 32430 7985
rect 32465 7950 32475 7985
rect 32510 7950 32520 7985
rect 32555 7950 32565 7985
rect 32600 7950 32610 7985
rect 32645 7950 32655 7985
rect 32690 7950 32700 7985
rect 32735 7950 32745 7985
rect 32780 7950 32790 7985
rect 32825 7950 32835 7985
rect 32870 7950 32890 7985
rect 31290 7940 32890 7950
rect 31290 7905 31305 7940
rect 31340 7905 31350 7940
rect 31385 7905 31395 7940
rect 31430 7905 31440 7940
rect 31475 7905 31485 7940
rect 31520 7905 31530 7940
rect 31565 7905 31575 7940
rect 31610 7905 31620 7940
rect 31655 7905 31665 7940
rect 31700 7905 31710 7940
rect 31745 7905 31755 7940
rect 31790 7905 31800 7940
rect 31835 7905 31845 7940
rect 31880 7905 31890 7940
rect 31925 7905 31935 7940
rect 31970 7905 31980 7940
rect 32015 7905 32025 7940
rect 32060 7905 32070 7940
rect 32105 7905 32115 7940
rect 32150 7905 32160 7940
rect 32195 7905 32205 7940
rect 32240 7905 32250 7940
rect 32285 7905 32295 7940
rect 32330 7905 32340 7940
rect 32375 7905 32385 7940
rect 32420 7905 32430 7940
rect 32465 7905 32475 7940
rect 32510 7905 32520 7940
rect 32555 7905 32565 7940
rect 32600 7905 32610 7940
rect 32645 7905 32655 7940
rect 32690 7905 32700 7940
rect 32735 7905 32745 7940
rect 32780 7905 32790 7940
rect 32825 7905 32835 7940
rect 32870 7905 32890 7940
rect 31290 7895 32890 7905
rect 31290 7860 31305 7895
rect 31340 7860 31350 7895
rect 31385 7860 31395 7895
rect 31430 7860 31440 7895
rect 31475 7860 31485 7895
rect 31520 7860 31530 7895
rect 31565 7860 31575 7895
rect 31610 7860 31620 7895
rect 31655 7860 31665 7895
rect 31700 7860 31710 7895
rect 31745 7860 31755 7895
rect 31790 7860 31800 7895
rect 31835 7860 31845 7895
rect 31880 7860 31890 7895
rect 31925 7860 31935 7895
rect 31970 7860 31980 7895
rect 32015 7860 32025 7895
rect 32060 7860 32070 7895
rect 32105 7860 32115 7895
rect 32150 7860 32160 7895
rect 32195 7860 32205 7895
rect 32240 7860 32250 7895
rect 32285 7860 32295 7895
rect 32330 7860 32340 7895
rect 32375 7860 32385 7895
rect 32420 7860 32430 7895
rect 32465 7860 32475 7895
rect 32510 7860 32520 7895
rect 32555 7860 32565 7895
rect 32600 7860 32610 7895
rect 32645 7860 32655 7895
rect 32690 7860 32700 7895
rect 32735 7860 32745 7895
rect 32780 7860 32790 7895
rect 32825 7860 32835 7895
rect 32870 7860 32890 7895
rect 31290 7850 32890 7860
rect 31290 7815 31305 7850
rect 31340 7815 31350 7850
rect 31385 7815 31395 7850
rect 31430 7815 31440 7850
rect 31475 7815 31485 7850
rect 31520 7815 31530 7850
rect 31565 7815 31575 7850
rect 31610 7815 31620 7850
rect 31655 7815 31665 7850
rect 31700 7815 31710 7850
rect 31745 7815 31755 7850
rect 31790 7815 31800 7850
rect 31835 7815 31845 7850
rect 31880 7815 31890 7850
rect 31925 7815 31935 7850
rect 31970 7815 31980 7850
rect 32015 7815 32025 7850
rect 32060 7815 32070 7850
rect 32105 7815 32115 7850
rect 32150 7815 32160 7850
rect 32195 7815 32205 7850
rect 32240 7815 32250 7850
rect 32285 7815 32295 7850
rect 32330 7815 32340 7850
rect 32375 7815 32385 7850
rect 32420 7815 32430 7850
rect 32465 7815 32475 7850
rect 32510 7815 32520 7850
rect 32555 7815 32565 7850
rect 32600 7815 32610 7850
rect 32645 7815 32655 7850
rect 32690 7815 32700 7850
rect 32735 7815 32745 7850
rect 32780 7815 32790 7850
rect 32825 7815 32835 7850
rect 32870 7815 32890 7850
rect 31290 7805 32890 7815
rect 31290 7770 31305 7805
rect 31340 7770 31350 7805
rect 31385 7770 31395 7805
rect 31430 7770 31440 7805
rect 31475 7770 31485 7805
rect 31520 7770 31530 7805
rect 31565 7770 31575 7805
rect 31610 7770 31620 7805
rect 31655 7770 31665 7805
rect 31700 7770 31710 7805
rect 31745 7770 31755 7805
rect 31790 7770 31800 7805
rect 31835 7770 31845 7805
rect 31880 7770 31890 7805
rect 31925 7770 31935 7805
rect 31970 7770 31980 7805
rect 32015 7770 32025 7805
rect 32060 7770 32070 7805
rect 32105 7770 32115 7805
rect 32150 7770 32160 7805
rect 32195 7770 32205 7805
rect 32240 7770 32250 7805
rect 32285 7770 32295 7805
rect 32330 7770 32340 7805
rect 32375 7770 32385 7805
rect 32420 7770 32430 7805
rect 32465 7770 32475 7805
rect 32510 7770 32520 7805
rect 32555 7770 32565 7805
rect 32600 7770 32610 7805
rect 32645 7770 32655 7805
rect 32690 7770 32700 7805
rect 32735 7770 32745 7805
rect 32780 7770 32790 7805
rect 32825 7770 32835 7805
rect 32870 7770 32890 7805
rect 31290 7760 32890 7770
rect 31290 7725 31305 7760
rect 31340 7725 31350 7760
rect 31385 7725 31395 7760
rect 31430 7725 31440 7760
rect 31475 7725 31485 7760
rect 31520 7725 31530 7760
rect 31565 7725 31575 7760
rect 31610 7725 31620 7760
rect 31655 7725 31665 7760
rect 31700 7725 31710 7760
rect 31745 7725 31755 7760
rect 31790 7725 31800 7760
rect 31835 7725 31845 7760
rect 31880 7725 31890 7760
rect 31925 7725 31935 7760
rect 31970 7725 31980 7760
rect 32015 7725 32025 7760
rect 32060 7725 32070 7760
rect 32105 7725 32115 7760
rect 32150 7725 32160 7760
rect 32195 7725 32205 7760
rect 32240 7725 32250 7760
rect 32285 7725 32295 7760
rect 32330 7725 32340 7760
rect 32375 7725 32385 7760
rect 32420 7725 32430 7760
rect 32465 7725 32475 7760
rect 32510 7725 32520 7760
rect 32555 7725 32565 7760
rect 32600 7725 32610 7760
rect 32645 7725 32655 7760
rect 32690 7725 32700 7760
rect 32735 7725 32745 7760
rect 32780 7725 32790 7760
rect 32825 7725 32835 7760
rect 32870 7725 32890 7760
rect 31290 7715 32890 7725
rect 31290 7680 31305 7715
rect 31340 7680 31350 7715
rect 31385 7680 31395 7715
rect 31430 7680 31440 7715
rect 31475 7680 31485 7715
rect 31520 7680 31530 7715
rect 31565 7680 31575 7715
rect 31610 7680 31620 7715
rect 31655 7680 31665 7715
rect 31700 7680 31710 7715
rect 31745 7680 31755 7715
rect 31790 7680 31800 7715
rect 31835 7680 31845 7715
rect 31880 7680 31890 7715
rect 31925 7680 31935 7715
rect 31970 7680 31980 7715
rect 32015 7680 32025 7715
rect 32060 7680 32070 7715
rect 32105 7680 32115 7715
rect 32150 7680 32160 7715
rect 32195 7680 32205 7715
rect 32240 7680 32250 7715
rect 32285 7680 32295 7715
rect 32330 7680 32340 7715
rect 32375 7680 32385 7715
rect 32420 7680 32430 7715
rect 32465 7680 32475 7715
rect 32510 7680 32520 7715
rect 32555 7680 32565 7715
rect 32600 7680 32610 7715
rect 32645 7680 32655 7715
rect 32690 7680 32700 7715
rect 32735 7680 32745 7715
rect 32780 7680 32790 7715
rect 32825 7680 32835 7715
rect 32870 7680 32890 7715
rect 31290 7670 32890 7680
rect 31290 7635 31305 7670
rect 31340 7635 31350 7670
rect 31385 7635 31395 7670
rect 31430 7635 31440 7670
rect 31475 7635 31485 7670
rect 31520 7635 31530 7670
rect 31565 7635 31575 7670
rect 31610 7635 31620 7670
rect 31655 7635 31665 7670
rect 31700 7635 31710 7670
rect 31745 7635 31755 7670
rect 31790 7635 31800 7670
rect 31835 7635 31845 7670
rect 31880 7635 31890 7670
rect 31925 7635 31935 7670
rect 31970 7635 31980 7670
rect 32015 7635 32025 7670
rect 32060 7635 32070 7670
rect 32105 7635 32115 7670
rect 32150 7635 32160 7670
rect 32195 7635 32205 7670
rect 32240 7635 32250 7670
rect 32285 7635 32295 7670
rect 32330 7635 32340 7670
rect 32375 7635 32385 7670
rect 32420 7635 32430 7670
rect 32465 7635 32475 7670
rect 32510 7635 32520 7670
rect 32555 7635 32565 7670
rect 32600 7635 32610 7670
rect 32645 7635 32655 7670
rect 32690 7635 32700 7670
rect 32735 7635 32745 7670
rect 32780 7635 32790 7670
rect 32825 7635 32835 7670
rect 32870 7635 32890 7670
rect 31290 7625 32890 7635
rect 31290 7590 31305 7625
rect 31340 7590 31350 7625
rect 31385 7590 31395 7625
rect 31430 7590 31440 7625
rect 31475 7590 31485 7625
rect 31520 7590 31530 7625
rect 31565 7590 31575 7625
rect 31610 7590 31620 7625
rect 31655 7590 31665 7625
rect 31700 7590 31710 7625
rect 31745 7590 31755 7625
rect 31790 7590 31800 7625
rect 31835 7590 31845 7625
rect 31880 7590 31890 7625
rect 31925 7590 31935 7625
rect 31970 7590 31980 7625
rect 32015 7590 32025 7625
rect 32060 7590 32070 7625
rect 32105 7590 32115 7625
rect 32150 7590 32160 7625
rect 32195 7590 32205 7625
rect 32240 7590 32250 7625
rect 32285 7590 32295 7625
rect 32330 7590 32340 7625
rect 32375 7590 32385 7625
rect 32420 7590 32430 7625
rect 32465 7590 32475 7625
rect 32510 7590 32520 7625
rect 32555 7590 32565 7625
rect 32600 7590 32610 7625
rect 32645 7590 32655 7625
rect 32690 7590 32700 7625
rect 32735 7590 32745 7625
rect 32780 7590 32790 7625
rect 32825 7590 32835 7625
rect 32870 7590 32890 7625
rect 31290 7580 32890 7590
rect 31290 7545 31305 7580
rect 31340 7545 31350 7580
rect 31385 7545 31395 7580
rect 31430 7545 31440 7580
rect 31475 7545 31485 7580
rect 31520 7545 31530 7580
rect 31565 7545 31575 7580
rect 31610 7545 31620 7580
rect 31655 7545 31665 7580
rect 31700 7545 31710 7580
rect 31745 7545 31755 7580
rect 31790 7545 31800 7580
rect 31835 7545 31845 7580
rect 31880 7545 31890 7580
rect 31925 7545 31935 7580
rect 31970 7545 31980 7580
rect 32015 7545 32025 7580
rect 32060 7545 32070 7580
rect 32105 7545 32115 7580
rect 32150 7545 32160 7580
rect 32195 7545 32205 7580
rect 32240 7545 32250 7580
rect 32285 7545 32295 7580
rect 32330 7545 32340 7580
rect 32375 7545 32385 7580
rect 32420 7545 32430 7580
rect 32465 7545 32475 7580
rect 32510 7545 32520 7580
rect 32555 7545 32565 7580
rect 32600 7545 32610 7580
rect 32645 7545 32655 7580
rect 32690 7545 32700 7580
rect 32735 7545 32745 7580
rect 32780 7545 32790 7580
rect 32825 7545 32835 7580
rect 32870 7545 32890 7580
rect 31290 7535 32890 7545
rect 31290 7500 31305 7535
rect 31340 7500 31350 7535
rect 31385 7500 31395 7535
rect 31430 7500 31440 7535
rect 31475 7500 31485 7535
rect 31520 7500 31530 7535
rect 31565 7500 31575 7535
rect 31610 7500 31620 7535
rect 31655 7500 31665 7535
rect 31700 7500 31710 7535
rect 31745 7500 31755 7535
rect 31790 7500 31800 7535
rect 31835 7500 31845 7535
rect 31880 7500 31890 7535
rect 31925 7500 31935 7535
rect 31970 7500 31980 7535
rect 32015 7500 32025 7535
rect 32060 7500 32070 7535
rect 32105 7500 32115 7535
rect 32150 7500 32160 7535
rect 32195 7500 32205 7535
rect 32240 7500 32250 7535
rect 32285 7500 32295 7535
rect 32330 7500 32340 7535
rect 32375 7500 32385 7535
rect 32420 7500 32430 7535
rect 32465 7500 32475 7535
rect 32510 7500 32520 7535
rect 32555 7500 32565 7535
rect 32600 7500 32610 7535
rect 32645 7500 32655 7535
rect 32690 7500 32700 7535
rect 32735 7500 32745 7535
rect 32780 7500 32790 7535
rect 32825 7500 32835 7535
rect 32870 7500 32890 7535
rect 31290 7490 32890 7500
rect 31290 7455 31305 7490
rect 31340 7455 31350 7490
rect 31385 7455 31395 7490
rect 31430 7455 31440 7490
rect 31475 7455 31485 7490
rect 31520 7455 31530 7490
rect 31565 7455 31575 7490
rect 31610 7455 31620 7490
rect 31655 7455 31665 7490
rect 31700 7455 31710 7490
rect 31745 7455 31755 7490
rect 31790 7455 31800 7490
rect 31835 7455 31845 7490
rect 31880 7455 31890 7490
rect 31925 7455 31935 7490
rect 31970 7455 31980 7490
rect 32015 7455 32025 7490
rect 32060 7455 32070 7490
rect 32105 7455 32115 7490
rect 32150 7455 32160 7490
rect 32195 7455 32205 7490
rect 32240 7455 32250 7490
rect 32285 7455 32295 7490
rect 32330 7455 32340 7490
rect 32375 7455 32385 7490
rect 32420 7455 32430 7490
rect 32465 7455 32475 7490
rect 32510 7455 32520 7490
rect 32555 7455 32565 7490
rect 32600 7455 32610 7490
rect 32645 7455 32655 7490
rect 32690 7455 32700 7490
rect 32735 7455 32745 7490
rect 32780 7455 32790 7490
rect 32825 7455 32835 7490
rect 32870 7455 32890 7490
rect 31290 7445 32890 7455
rect 31290 7410 31305 7445
rect 31340 7410 31350 7445
rect 31385 7410 31395 7445
rect 31430 7410 31440 7445
rect 31475 7410 31485 7445
rect 31520 7410 31530 7445
rect 31565 7410 31575 7445
rect 31610 7410 31620 7445
rect 31655 7410 31665 7445
rect 31700 7410 31710 7445
rect 31745 7410 31755 7445
rect 31790 7410 31800 7445
rect 31835 7410 31845 7445
rect 31880 7410 31890 7445
rect 31925 7410 31935 7445
rect 31970 7410 31980 7445
rect 32015 7410 32025 7445
rect 32060 7410 32070 7445
rect 32105 7410 32115 7445
rect 32150 7410 32160 7445
rect 32195 7410 32205 7445
rect 32240 7410 32250 7445
rect 32285 7410 32295 7445
rect 32330 7410 32340 7445
rect 32375 7410 32385 7445
rect 32420 7410 32430 7445
rect 32465 7410 32475 7445
rect 32510 7410 32520 7445
rect 32555 7410 32565 7445
rect 32600 7410 32610 7445
rect 32645 7410 32655 7445
rect 32690 7410 32700 7445
rect 32735 7410 32745 7445
rect 32780 7410 32790 7445
rect 32825 7410 32835 7445
rect 32870 7410 32890 7445
rect 31290 7400 32890 7410
rect 31290 7365 31305 7400
rect 31340 7365 31350 7400
rect 31385 7365 31395 7400
rect 31430 7365 31440 7400
rect 31475 7365 31485 7400
rect 31520 7365 31530 7400
rect 31565 7365 31575 7400
rect 31610 7365 31620 7400
rect 31655 7365 31665 7400
rect 31700 7365 31710 7400
rect 31745 7365 31755 7400
rect 31790 7365 31800 7400
rect 31835 7365 31845 7400
rect 31880 7365 31890 7400
rect 31925 7365 31935 7400
rect 31970 7365 31980 7400
rect 32015 7365 32025 7400
rect 32060 7365 32070 7400
rect 32105 7365 32115 7400
rect 32150 7365 32160 7400
rect 32195 7365 32205 7400
rect 32240 7365 32250 7400
rect 32285 7365 32295 7400
rect 32330 7365 32340 7400
rect 32375 7365 32385 7400
rect 32420 7365 32430 7400
rect 32465 7365 32475 7400
rect 32510 7365 32520 7400
rect 32555 7365 32565 7400
rect 32600 7365 32610 7400
rect 32645 7365 32655 7400
rect 32690 7365 32700 7400
rect 32735 7365 32745 7400
rect 32780 7365 32790 7400
rect 32825 7365 32835 7400
rect 32870 7365 32890 7400
rect 31290 7355 32890 7365
rect 31290 7320 31305 7355
rect 31340 7320 31350 7355
rect 31385 7320 31395 7355
rect 31430 7320 31440 7355
rect 31475 7320 31485 7355
rect 31520 7320 31530 7355
rect 31565 7320 31575 7355
rect 31610 7320 31620 7355
rect 31655 7320 31665 7355
rect 31700 7320 31710 7355
rect 31745 7320 31755 7355
rect 31790 7320 31800 7355
rect 31835 7320 31845 7355
rect 31880 7320 31890 7355
rect 31925 7320 31935 7355
rect 31970 7320 31980 7355
rect 32015 7320 32025 7355
rect 32060 7320 32070 7355
rect 32105 7320 32115 7355
rect 32150 7320 32160 7355
rect 32195 7320 32205 7355
rect 32240 7320 32250 7355
rect 32285 7320 32295 7355
rect 32330 7320 32340 7355
rect 32375 7320 32385 7355
rect 32420 7320 32430 7355
rect 32465 7320 32475 7355
rect 32510 7320 32520 7355
rect 32555 7320 32565 7355
rect 32600 7320 32610 7355
rect 32645 7320 32655 7355
rect 32690 7320 32700 7355
rect 32735 7320 32745 7355
rect 32780 7320 32790 7355
rect 32825 7320 32835 7355
rect 32870 7320 32890 7355
rect 31290 7310 32890 7320
rect 31290 7275 31305 7310
rect 31340 7275 31350 7310
rect 31385 7275 31395 7310
rect 31430 7275 31440 7310
rect 31475 7275 31485 7310
rect 31520 7275 31530 7310
rect 31565 7275 31575 7310
rect 31610 7275 31620 7310
rect 31655 7275 31665 7310
rect 31700 7275 31710 7310
rect 31745 7275 31755 7310
rect 31790 7275 31800 7310
rect 31835 7275 31845 7310
rect 31880 7275 31890 7310
rect 31925 7275 31935 7310
rect 31970 7275 31980 7310
rect 32015 7275 32025 7310
rect 32060 7275 32070 7310
rect 32105 7275 32115 7310
rect 32150 7275 32160 7310
rect 32195 7275 32205 7310
rect 32240 7275 32250 7310
rect 32285 7275 32295 7310
rect 32330 7275 32340 7310
rect 32375 7275 32385 7310
rect 32420 7275 32430 7310
rect 32465 7275 32475 7310
rect 32510 7275 32520 7310
rect 32555 7275 32565 7310
rect 32600 7275 32610 7310
rect 32645 7275 32655 7310
rect 32690 7275 32700 7310
rect 32735 7275 32745 7310
rect 32780 7275 32790 7310
rect 32825 7275 32835 7310
rect 32870 7275 32890 7310
rect 31290 7265 32890 7275
rect 31290 7230 31305 7265
rect 31340 7230 31350 7265
rect 31385 7230 31395 7265
rect 31430 7230 31440 7265
rect 31475 7230 31485 7265
rect 31520 7230 31530 7265
rect 31565 7230 31575 7265
rect 31610 7230 31620 7265
rect 31655 7230 31665 7265
rect 31700 7230 31710 7265
rect 31745 7230 31755 7265
rect 31790 7230 31800 7265
rect 31835 7230 31845 7265
rect 31880 7230 31890 7265
rect 31925 7230 31935 7265
rect 31970 7230 31980 7265
rect 32015 7230 32025 7265
rect 32060 7230 32070 7265
rect 32105 7230 32115 7265
rect 32150 7230 32160 7265
rect 32195 7230 32205 7265
rect 32240 7230 32250 7265
rect 32285 7230 32295 7265
rect 32330 7230 32340 7265
rect 32375 7230 32385 7265
rect 32420 7230 32430 7265
rect 32465 7230 32475 7265
rect 32510 7230 32520 7265
rect 32555 7230 32565 7265
rect 32600 7230 32610 7265
rect 32645 7230 32655 7265
rect 32690 7230 32700 7265
rect 32735 7230 32745 7265
rect 32780 7230 32790 7265
rect 32825 7230 32835 7265
rect 32870 7230 32890 7265
rect 31290 7220 32890 7230
rect 31290 7185 31305 7220
rect 31340 7185 31350 7220
rect 31385 7185 31395 7220
rect 31430 7185 31440 7220
rect 31475 7185 31485 7220
rect 31520 7185 31530 7220
rect 31565 7185 31575 7220
rect 31610 7185 31620 7220
rect 31655 7185 31665 7220
rect 31700 7185 31710 7220
rect 31745 7185 31755 7220
rect 31790 7185 31800 7220
rect 31835 7185 31845 7220
rect 31880 7185 31890 7220
rect 31925 7185 31935 7220
rect 31970 7185 31980 7220
rect 32015 7185 32025 7220
rect 32060 7185 32070 7220
rect 32105 7185 32115 7220
rect 32150 7185 32160 7220
rect 32195 7185 32205 7220
rect 32240 7185 32250 7220
rect 32285 7185 32295 7220
rect 32330 7185 32340 7220
rect 32375 7185 32385 7220
rect 32420 7185 32430 7220
rect 32465 7185 32475 7220
rect 32510 7185 32520 7220
rect 32555 7185 32565 7220
rect 32600 7185 32610 7220
rect 32645 7185 32655 7220
rect 32690 7185 32700 7220
rect 32735 7185 32745 7220
rect 32780 7185 32790 7220
rect 32825 7185 32835 7220
rect 32870 7185 32890 7220
rect 31290 7175 32890 7185
rect 31290 7140 31305 7175
rect 31340 7140 31350 7175
rect 31385 7140 31395 7175
rect 31430 7140 31440 7175
rect 31475 7140 31485 7175
rect 31520 7140 31530 7175
rect 31565 7140 31575 7175
rect 31610 7140 31620 7175
rect 31655 7140 31665 7175
rect 31700 7140 31710 7175
rect 31745 7140 31755 7175
rect 31790 7140 31800 7175
rect 31835 7140 31845 7175
rect 31880 7140 31890 7175
rect 31925 7140 31935 7175
rect 31970 7140 31980 7175
rect 32015 7140 32025 7175
rect 32060 7140 32070 7175
rect 32105 7140 32115 7175
rect 32150 7140 32160 7175
rect 32195 7140 32205 7175
rect 32240 7140 32250 7175
rect 32285 7140 32295 7175
rect 32330 7140 32340 7175
rect 32375 7140 32385 7175
rect 32420 7140 32430 7175
rect 32465 7140 32475 7175
rect 32510 7140 32520 7175
rect 32555 7140 32565 7175
rect 32600 7140 32610 7175
rect 32645 7140 32655 7175
rect 32690 7140 32700 7175
rect 32735 7140 32745 7175
rect 32780 7140 32790 7175
rect 32825 7140 32835 7175
rect 32870 7140 32890 7175
rect 31290 7130 32890 7140
rect 31290 7095 31305 7130
rect 31340 7095 31350 7130
rect 31385 7095 31395 7130
rect 31430 7095 31440 7130
rect 31475 7095 31485 7130
rect 31520 7095 31530 7130
rect 31565 7095 31575 7130
rect 31610 7095 31620 7130
rect 31655 7095 31665 7130
rect 31700 7095 31710 7130
rect 31745 7095 31755 7130
rect 31790 7095 31800 7130
rect 31835 7095 31845 7130
rect 31880 7095 31890 7130
rect 31925 7095 31935 7130
rect 31970 7095 31980 7130
rect 32015 7095 32025 7130
rect 32060 7095 32070 7130
rect 32105 7095 32115 7130
rect 32150 7095 32160 7130
rect 32195 7095 32205 7130
rect 32240 7095 32250 7130
rect 32285 7095 32295 7130
rect 32330 7095 32340 7130
rect 32375 7095 32385 7130
rect 32420 7095 32430 7130
rect 32465 7095 32475 7130
rect 32510 7095 32520 7130
rect 32555 7095 32565 7130
rect 32600 7095 32610 7130
rect 32645 7095 32655 7130
rect 32690 7095 32700 7130
rect 32735 7095 32745 7130
rect 32780 7095 32790 7130
rect 32825 7095 32835 7130
rect 32870 7095 32890 7130
rect 31290 7085 32890 7095
rect 31290 7050 31305 7085
rect 31340 7050 31350 7085
rect 31385 7050 31395 7085
rect 31430 7050 31440 7085
rect 31475 7050 31485 7085
rect 31520 7050 31530 7085
rect 31565 7050 31575 7085
rect 31610 7050 31620 7085
rect 31655 7050 31665 7085
rect 31700 7050 31710 7085
rect 31745 7050 31755 7085
rect 31790 7050 31800 7085
rect 31835 7050 31845 7085
rect 31880 7050 31890 7085
rect 31925 7050 31935 7085
rect 31970 7050 31980 7085
rect 32015 7050 32025 7085
rect 32060 7050 32070 7085
rect 32105 7050 32115 7085
rect 32150 7050 32160 7085
rect 32195 7050 32205 7085
rect 32240 7050 32250 7085
rect 32285 7050 32295 7085
rect 32330 7050 32340 7085
rect 32375 7050 32385 7085
rect 32420 7050 32430 7085
rect 32465 7050 32475 7085
rect 32510 7050 32520 7085
rect 32555 7050 32565 7085
rect 32600 7050 32610 7085
rect 32645 7050 32655 7085
rect 32690 7050 32700 7085
rect 32735 7050 32745 7085
rect 32780 7050 32790 7085
rect 32825 7050 32835 7085
rect 32870 7050 32890 7085
rect 31290 7040 32890 7050
rect 31290 7005 31305 7040
rect 31340 7005 31350 7040
rect 31385 7005 31395 7040
rect 31430 7005 31440 7040
rect 31475 7005 31485 7040
rect 31520 7005 31530 7040
rect 31565 7005 31575 7040
rect 31610 7005 31620 7040
rect 31655 7005 31665 7040
rect 31700 7005 31710 7040
rect 31745 7005 31755 7040
rect 31790 7005 31800 7040
rect 31835 7005 31845 7040
rect 31880 7005 31890 7040
rect 31925 7005 31935 7040
rect 31970 7005 31980 7040
rect 32015 7005 32025 7040
rect 32060 7005 32070 7040
rect 32105 7005 32115 7040
rect 32150 7005 32160 7040
rect 32195 7005 32205 7040
rect 32240 7005 32250 7040
rect 32285 7005 32295 7040
rect 32330 7005 32340 7040
rect 32375 7005 32385 7040
rect 32420 7005 32430 7040
rect 32465 7005 32475 7040
rect 32510 7005 32520 7040
rect 32555 7005 32565 7040
rect 32600 7005 32610 7040
rect 32645 7005 32655 7040
rect 32690 7005 32700 7040
rect 32735 7005 32745 7040
rect 32780 7005 32790 7040
rect 32825 7005 32835 7040
rect 32870 7005 32890 7040
rect 31290 6995 32890 7005
rect 31290 6960 31305 6995
rect 31340 6960 31350 6995
rect 31385 6960 31395 6995
rect 31430 6960 31440 6995
rect 31475 6960 31485 6995
rect 31520 6960 31530 6995
rect 31565 6960 31575 6995
rect 31610 6960 31620 6995
rect 31655 6960 31665 6995
rect 31700 6960 31710 6995
rect 31745 6960 31755 6995
rect 31790 6960 31800 6995
rect 31835 6960 31845 6995
rect 31880 6960 31890 6995
rect 31925 6960 31935 6995
rect 31970 6960 31980 6995
rect 32015 6960 32025 6995
rect 32060 6960 32070 6995
rect 32105 6960 32115 6995
rect 32150 6960 32160 6995
rect 32195 6960 32205 6995
rect 32240 6960 32250 6995
rect 32285 6960 32295 6995
rect 32330 6960 32340 6995
rect 32375 6960 32385 6995
rect 32420 6960 32430 6995
rect 32465 6960 32475 6995
rect 32510 6960 32520 6995
rect 32555 6960 32565 6995
rect 32600 6960 32610 6995
rect 32645 6960 32655 6995
rect 32690 6960 32700 6995
rect 32735 6960 32745 6995
rect 32780 6960 32790 6995
rect 32825 6960 32835 6995
rect 32870 6960 32890 6995
rect 31290 6950 32890 6960
rect 31290 6915 31305 6950
rect 31340 6915 31350 6950
rect 31385 6915 31395 6950
rect 31430 6915 31440 6950
rect 31475 6915 31485 6950
rect 31520 6915 31530 6950
rect 31565 6915 31575 6950
rect 31610 6915 31620 6950
rect 31655 6915 31665 6950
rect 31700 6915 31710 6950
rect 31745 6915 31755 6950
rect 31790 6915 31800 6950
rect 31835 6915 31845 6950
rect 31880 6915 31890 6950
rect 31925 6915 31935 6950
rect 31970 6915 31980 6950
rect 32015 6915 32025 6950
rect 32060 6915 32070 6950
rect 32105 6915 32115 6950
rect 32150 6915 32160 6950
rect 32195 6915 32205 6950
rect 32240 6915 32250 6950
rect 32285 6915 32295 6950
rect 32330 6915 32340 6950
rect 32375 6915 32385 6950
rect 32420 6915 32430 6950
rect 32465 6915 32475 6950
rect 32510 6915 32520 6950
rect 32555 6915 32565 6950
rect 32600 6915 32610 6950
rect 32645 6915 32655 6950
rect 32690 6915 32700 6950
rect 32735 6915 32745 6950
rect 32780 6915 32790 6950
rect 32825 6915 32835 6950
rect 32870 6915 32890 6950
rect 31290 6905 32890 6915
rect 31290 6870 31305 6905
rect 31340 6870 31350 6905
rect 31385 6870 31395 6905
rect 31430 6870 31440 6905
rect 31475 6870 31485 6905
rect 31520 6870 31530 6905
rect 31565 6870 31575 6905
rect 31610 6870 31620 6905
rect 31655 6870 31665 6905
rect 31700 6870 31710 6905
rect 31745 6870 31755 6905
rect 31790 6870 31800 6905
rect 31835 6870 31845 6905
rect 31880 6870 31890 6905
rect 31925 6870 31935 6905
rect 31970 6870 31980 6905
rect 32015 6870 32025 6905
rect 32060 6870 32070 6905
rect 32105 6870 32115 6905
rect 32150 6870 32160 6905
rect 32195 6870 32205 6905
rect 32240 6870 32250 6905
rect 32285 6870 32295 6905
rect 32330 6870 32340 6905
rect 32375 6870 32385 6905
rect 32420 6870 32430 6905
rect 32465 6870 32475 6905
rect 32510 6870 32520 6905
rect 32555 6870 32565 6905
rect 32600 6870 32610 6905
rect 32645 6870 32655 6905
rect 32690 6870 32700 6905
rect 32735 6870 32745 6905
rect 32780 6870 32790 6905
rect 32825 6870 32835 6905
rect 32870 6870 32890 6905
rect 31290 6860 32890 6870
rect 31290 6825 31305 6860
rect 31340 6825 31350 6860
rect 31385 6825 31395 6860
rect 31430 6825 31440 6860
rect 31475 6825 31485 6860
rect 31520 6825 31530 6860
rect 31565 6825 31575 6860
rect 31610 6825 31620 6860
rect 31655 6825 31665 6860
rect 31700 6825 31710 6860
rect 31745 6825 31755 6860
rect 31790 6825 31800 6860
rect 31835 6825 31845 6860
rect 31880 6825 31890 6860
rect 31925 6825 31935 6860
rect 31970 6825 31980 6860
rect 32015 6825 32025 6860
rect 32060 6825 32070 6860
rect 32105 6825 32115 6860
rect 32150 6825 32160 6860
rect 32195 6825 32205 6860
rect 32240 6825 32250 6860
rect 32285 6825 32295 6860
rect 32330 6825 32340 6860
rect 32375 6825 32385 6860
rect 32420 6825 32430 6860
rect 32465 6825 32475 6860
rect 32510 6825 32520 6860
rect 32555 6825 32565 6860
rect 32600 6825 32610 6860
rect 32645 6825 32655 6860
rect 32690 6825 32700 6860
rect 32735 6825 32745 6860
rect 32780 6825 32790 6860
rect 32825 6825 32835 6860
rect 32870 6825 32890 6860
rect 31290 6815 32890 6825
rect 31290 6780 31305 6815
rect 31340 6780 31350 6815
rect 31385 6780 31395 6815
rect 31430 6780 31440 6815
rect 31475 6780 31485 6815
rect 31520 6780 31530 6815
rect 31565 6780 31575 6815
rect 31610 6780 31620 6815
rect 31655 6780 31665 6815
rect 31700 6780 31710 6815
rect 31745 6780 31755 6815
rect 31790 6780 31800 6815
rect 31835 6780 31845 6815
rect 31880 6780 31890 6815
rect 31925 6780 31935 6815
rect 31970 6780 31980 6815
rect 32015 6780 32025 6815
rect 32060 6780 32070 6815
rect 32105 6780 32115 6815
rect 32150 6780 32160 6815
rect 32195 6780 32205 6815
rect 32240 6780 32250 6815
rect 32285 6780 32295 6815
rect 32330 6780 32340 6815
rect 32375 6780 32385 6815
rect 32420 6780 32430 6815
rect 32465 6780 32475 6815
rect 32510 6780 32520 6815
rect 32555 6780 32565 6815
rect 32600 6780 32610 6815
rect 32645 6780 32655 6815
rect 32690 6780 32700 6815
rect 32735 6780 32745 6815
rect 32780 6780 32790 6815
rect 32825 6780 32835 6815
rect 32870 6780 32890 6815
rect 31290 6770 32890 6780
rect 31290 6735 31305 6770
rect 31340 6735 31350 6770
rect 31385 6735 31395 6770
rect 31430 6735 31440 6770
rect 31475 6735 31485 6770
rect 31520 6735 31530 6770
rect 31565 6735 31575 6770
rect 31610 6735 31620 6770
rect 31655 6735 31665 6770
rect 31700 6735 31710 6770
rect 31745 6735 31755 6770
rect 31790 6735 31800 6770
rect 31835 6735 31845 6770
rect 31880 6735 31890 6770
rect 31925 6735 31935 6770
rect 31970 6735 31980 6770
rect 32015 6735 32025 6770
rect 32060 6735 32070 6770
rect 32105 6735 32115 6770
rect 32150 6735 32160 6770
rect 32195 6735 32205 6770
rect 32240 6735 32250 6770
rect 32285 6735 32295 6770
rect 32330 6735 32340 6770
rect 32375 6735 32385 6770
rect 32420 6735 32430 6770
rect 32465 6735 32475 6770
rect 32510 6735 32520 6770
rect 32555 6735 32565 6770
rect 32600 6735 32610 6770
rect 32645 6735 32655 6770
rect 32690 6735 32700 6770
rect 32735 6735 32745 6770
rect 32780 6735 32790 6770
rect 32825 6735 32835 6770
rect 32870 6735 32890 6770
rect 31290 6725 32890 6735
rect 31290 6690 31305 6725
rect 31340 6690 31350 6725
rect 31385 6690 31395 6725
rect 31430 6690 31440 6725
rect 31475 6690 31485 6725
rect 31520 6690 31530 6725
rect 31565 6690 31575 6725
rect 31610 6690 31620 6725
rect 31655 6690 31665 6725
rect 31700 6690 31710 6725
rect 31745 6690 31755 6725
rect 31790 6690 31800 6725
rect 31835 6690 31845 6725
rect 31880 6690 31890 6725
rect 31925 6690 31935 6725
rect 31970 6690 31980 6725
rect 32015 6690 32025 6725
rect 32060 6690 32070 6725
rect 32105 6690 32115 6725
rect 32150 6690 32160 6725
rect 32195 6690 32205 6725
rect 32240 6690 32250 6725
rect 32285 6690 32295 6725
rect 32330 6690 32340 6725
rect 32375 6690 32385 6725
rect 32420 6690 32430 6725
rect 32465 6690 32475 6725
rect 32510 6690 32520 6725
rect 32555 6690 32565 6725
rect 32600 6690 32610 6725
rect 32645 6690 32655 6725
rect 32690 6690 32700 6725
rect 32735 6690 32745 6725
rect 32780 6690 32790 6725
rect 32825 6690 32835 6725
rect 32870 6690 32890 6725
rect 31290 6680 32890 6690
rect 31290 6645 31305 6680
rect 31340 6645 31350 6680
rect 31385 6645 31395 6680
rect 31430 6645 31440 6680
rect 31475 6645 31485 6680
rect 31520 6645 31530 6680
rect 31565 6645 31575 6680
rect 31610 6645 31620 6680
rect 31655 6645 31665 6680
rect 31700 6645 31710 6680
rect 31745 6645 31755 6680
rect 31790 6645 31800 6680
rect 31835 6645 31845 6680
rect 31880 6645 31890 6680
rect 31925 6645 31935 6680
rect 31970 6645 31980 6680
rect 32015 6645 32025 6680
rect 32060 6645 32070 6680
rect 32105 6645 32115 6680
rect 32150 6645 32160 6680
rect 32195 6645 32205 6680
rect 32240 6645 32250 6680
rect 32285 6645 32295 6680
rect 32330 6645 32340 6680
rect 32375 6645 32385 6680
rect 32420 6645 32430 6680
rect 32465 6645 32475 6680
rect 32510 6645 32520 6680
rect 32555 6645 32565 6680
rect 32600 6645 32610 6680
rect 32645 6645 32655 6680
rect 32690 6645 32700 6680
rect 32735 6645 32745 6680
rect 32780 6645 32790 6680
rect 32825 6645 32835 6680
rect 32870 6645 32890 6680
rect 31290 6635 32890 6645
rect 31290 6600 31305 6635
rect 31340 6600 31350 6635
rect 31385 6600 31395 6635
rect 31430 6600 31440 6635
rect 31475 6600 31485 6635
rect 31520 6600 31530 6635
rect 31565 6600 31575 6635
rect 31610 6600 31620 6635
rect 31655 6600 31665 6635
rect 31700 6600 31710 6635
rect 31745 6600 31755 6635
rect 31790 6600 31800 6635
rect 31835 6600 31845 6635
rect 31880 6600 31890 6635
rect 31925 6600 31935 6635
rect 31970 6600 31980 6635
rect 32015 6600 32025 6635
rect 32060 6600 32070 6635
rect 32105 6600 32115 6635
rect 32150 6600 32160 6635
rect 32195 6600 32205 6635
rect 32240 6600 32250 6635
rect 32285 6600 32295 6635
rect 32330 6600 32340 6635
rect 32375 6600 32385 6635
rect 32420 6600 32430 6635
rect 32465 6600 32475 6635
rect 32510 6600 32520 6635
rect 32555 6600 32565 6635
rect 32600 6600 32610 6635
rect 32645 6600 32655 6635
rect 32690 6600 32700 6635
rect 32735 6600 32745 6635
rect 32780 6600 32790 6635
rect 32825 6600 32835 6635
rect 32870 6600 32890 6635
rect 31290 6590 32890 6600
rect 31290 6555 31305 6590
rect 31340 6555 31350 6590
rect 31385 6555 31395 6590
rect 31430 6555 31440 6590
rect 31475 6555 31485 6590
rect 31520 6555 31530 6590
rect 31565 6555 31575 6590
rect 31610 6555 31620 6590
rect 31655 6555 31665 6590
rect 31700 6555 31710 6590
rect 31745 6555 31755 6590
rect 31790 6555 31800 6590
rect 31835 6555 31845 6590
rect 31880 6555 31890 6590
rect 31925 6555 31935 6590
rect 31970 6555 31980 6590
rect 32015 6555 32025 6590
rect 32060 6555 32070 6590
rect 32105 6555 32115 6590
rect 32150 6555 32160 6590
rect 32195 6555 32205 6590
rect 32240 6555 32250 6590
rect 32285 6555 32295 6590
rect 32330 6555 32340 6590
rect 32375 6555 32385 6590
rect 32420 6555 32430 6590
rect 32465 6555 32475 6590
rect 32510 6555 32520 6590
rect 32555 6555 32565 6590
rect 32600 6555 32610 6590
rect 32645 6555 32655 6590
rect 32690 6555 32700 6590
rect 32735 6555 32745 6590
rect 32780 6555 32790 6590
rect 32825 6555 32835 6590
rect 32870 6555 32890 6590
rect 31290 6545 32890 6555
rect 31290 6510 31305 6545
rect 31340 6510 31350 6545
rect 31385 6510 31395 6545
rect 31430 6510 31440 6545
rect 31475 6510 31485 6545
rect 31520 6510 31530 6545
rect 31565 6510 31575 6545
rect 31610 6510 31620 6545
rect 31655 6510 31665 6545
rect 31700 6510 31710 6545
rect 31745 6510 31755 6545
rect 31790 6510 31800 6545
rect 31835 6510 31845 6545
rect 31880 6510 31890 6545
rect 31925 6510 31935 6545
rect 31970 6510 31980 6545
rect 32015 6510 32025 6545
rect 32060 6510 32070 6545
rect 32105 6510 32115 6545
rect 32150 6510 32160 6545
rect 32195 6510 32205 6545
rect 32240 6510 32250 6545
rect 32285 6510 32295 6545
rect 32330 6510 32340 6545
rect 32375 6510 32385 6545
rect 32420 6510 32430 6545
rect 32465 6510 32475 6545
rect 32510 6510 32520 6545
rect 32555 6510 32565 6545
rect 32600 6510 32610 6545
rect 32645 6510 32655 6545
rect 32690 6510 32700 6545
rect 32735 6510 32745 6545
rect 32780 6510 32790 6545
rect 32825 6510 32835 6545
rect 32870 6510 32890 6545
rect 31290 6500 32890 6510
rect 31290 6465 31305 6500
rect 31340 6465 31350 6500
rect 31385 6465 31395 6500
rect 31430 6465 31440 6500
rect 31475 6465 31485 6500
rect 31520 6465 31530 6500
rect 31565 6465 31575 6500
rect 31610 6465 31620 6500
rect 31655 6465 31665 6500
rect 31700 6465 31710 6500
rect 31745 6465 31755 6500
rect 31790 6465 31800 6500
rect 31835 6465 31845 6500
rect 31880 6465 31890 6500
rect 31925 6465 31935 6500
rect 31970 6465 31980 6500
rect 32015 6465 32025 6500
rect 32060 6465 32070 6500
rect 32105 6465 32115 6500
rect 32150 6465 32160 6500
rect 32195 6465 32205 6500
rect 32240 6465 32250 6500
rect 32285 6465 32295 6500
rect 32330 6465 32340 6500
rect 32375 6465 32385 6500
rect 32420 6465 32430 6500
rect 32465 6465 32475 6500
rect 32510 6465 32520 6500
rect 32555 6465 32565 6500
rect 32600 6465 32610 6500
rect 32645 6465 32655 6500
rect 32690 6465 32700 6500
rect 32735 6465 32745 6500
rect 32780 6465 32790 6500
rect 32825 6465 32835 6500
rect 32870 6465 32890 6500
rect -90 -1300 -30 -1290
rect -90 -1340 -80 -1300
rect -40 -1340 -30 -1300
rect -90 -1365 -30 -1340
rect -90 -1405 -80 -1365
rect -40 -1405 -30 -1365
rect -90 -1435 -30 -1405
rect -90 -1475 -80 -1435
rect -40 -1475 -30 -1435
rect -90 -1505 -30 -1475
rect -90 -1545 -80 -1505
rect -40 -1545 -30 -1505
rect -90 -1575 -30 -1545
rect -90 -1615 -80 -1575
rect -40 -1615 -30 -1575
rect -90 -1640 -30 -1615
rect -90 -1680 -80 -1640
rect -40 -1680 -30 -1640
rect -90 -1700 -30 -1680
rect -90 -1740 -80 -1700
rect -40 -1740 -30 -1700
rect -90 -1765 -30 -1740
rect -90 -1805 -80 -1765
rect -40 -1805 -30 -1765
rect -90 -1835 -30 -1805
rect -90 -1875 -80 -1835
rect -40 -1875 -30 -1835
rect -90 -1905 -30 -1875
rect -90 -1945 -80 -1905
rect -40 -1945 -30 -1905
rect -90 -1975 -30 -1945
rect -90 -2015 -80 -1975
rect -40 -2015 -30 -1975
rect -90 -2040 -30 -2015
rect -90 -2080 -80 -2040
rect -40 -2080 -30 -2040
rect -90 -2100 -30 -2080
rect -90 -2140 -80 -2100
rect -40 -2140 -30 -2100
rect -90 -2165 -30 -2140
rect -90 -2205 -80 -2165
rect -40 -2205 -30 -2165
rect -90 -2235 -30 -2205
rect -90 -2275 -80 -2235
rect -40 -2275 -30 -2235
rect -90 -2305 -30 -2275
rect -90 -2345 -80 -2305
rect -40 -2345 -30 -2305
rect -90 -2375 -30 -2345
rect -90 -2415 -80 -2375
rect -40 -2415 -30 -2375
rect -90 -2440 -30 -2415
rect -90 -2480 -80 -2440
rect -40 -2480 -30 -2440
rect -90 -2500 -30 -2480
rect -90 -2540 -80 -2500
rect -40 -2540 -30 -2500
rect -90 -2565 -30 -2540
rect -90 -2605 -80 -2565
rect -40 -2605 -30 -2565
rect -90 -2635 -30 -2605
rect -90 -2675 -80 -2635
rect -40 -2675 -30 -2635
rect -90 -2705 -30 -2675
rect -90 -2745 -80 -2705
rect -40 -2745 -30 -2705
rect -90 -2775 -30 -2745
rect -90 -2815 -80 -2775
rect -40 -2815 -30 -2775
rect -90 -2840 -30 -2815
rect -90 -2880 -80 -2840
rect -40 -2880 -30 -2840
rect -90 -2890 -30 -2880
rect 260 -1300 320 -1290
rect 260 -1340 270 -1300
rect 310 -1340 320 -1300
rect 260 -1365 320 -1340
rect 260 -1405 270 -1365
rect 310 -1405 320 -1365
rect 260 -1435 320 -1405
rect 260 -1475 270 -1435
rect 310 -1475 320 -1435
rect 260 -1505 320 -1475
rect 260 -1545 270 -1505
rect 310 -1545 320 -1505
rect 260 -1575 320 -1545
rect 260 -1615 270 -1575
rect 310 -1615 320 -1575
rect 260 -1640 320 -1615
rect 260 -1680 270 -1640
rect 310 -1680 320 -1640
rect 260 -1700 320 -1680
rect 260 -1740 270 -1700
rect 310 -1740 320 -1700
rect 260 -1765 320 -1740
rect 260 -1805 270 -1765
rect 310 -1805 320 -1765
rect 260 -1835 320 -1805
rect 260 -1875 270 -1835
rect 310 -1875 320 -1835
rect 260 -1905 320 -1875
rect 260 -1945 270 -1905
rect 310 -1945 320 -1905
rect 260 -1975 320 -1945
rect 260 -2015 270 -1975
rect 310 -2015 320 -1975
rect 260 -2040 320 -2015
rect 260 -2080 270 -2040
rect 310 -2080 320 -2040
rect 260 -2100 320 -2080
rect 260 -2140 270 -2100
rect 310 -2140 320 -2100
rect 260 -2165 320 -2140
rect 260 -2205 270 -2165
rect 310 -2205 320 -2165
rect 260 -2235 320 -2205
rect 260 -2275 270 -2235
rect 310 -2275 320 -2235
rect 260 -2305 320 -2275
rect 260 -2345 270 -2305
rect 310 -2345 320 -2305
rect 260 -2375 320 -2345
rect 260 -2415 270 -2375
rect 310 -2415 320 -2375
rect 260 -2440 320 -2415
rect 260 -2480 270 -2440
rect 310 -2480 320 -2440
rect 260 -2500 320 -2480
rect 260 -2540 270 -2500
rect 310 -2540 320 -2500
rect 260 -2565 320 -2540
rect 260 -2605 270 -2565
rect 310 -2605 320 -2565
rect 260 -2635 320 -2605
rect 260 -2675 270 -2635
rect 310 -2675 320 -2635
rect 260 -2705 320 -2675
rect 260 -2745 270 -2705
rect 310 -2745 320 -2705
rect 260 -2775 320 -2745
rect 260 -2815 270 -2775
rect 310 -2815 320 -2775
rect 260 -2840 320 -2815
rect 260 -2880 270 -2840
rect 310 -2880 320 -2840
rect 260 -2890 320 -2880
rect 610 -1300 670 -1290
rect 610 -1340 620 -1300
rect 660 -1340 670 -1300
rect 610 -1365 670 -1340
rect 610 -1405 620 -1365
rect 660 -1405 670 -1365
rect 610 -1435 670 -1405
rect 610 -1475 620 -1435
rect 660 -1475 670 -1435
rect 610 -1505 670 -1475
rect 610 -1545 620 -1505
rect 660 -1545 670 -1505
rect 610 -1575 670 -1545
rect 610 -1615 620 -1575
rect 660 -1615 670 -1575
rect 610 -1640 670 -1615
rect 610 -1680 620 -1640
rect 660 -1680 670 -1640
rect 610 -1700 670 -1680
rect 610 -1740 620 -1700
rect 660 -1740 670 -1700
rect 610 -1765 670 -1740
rect 610 -1805 620 -1765
rect 660 -1805 670 -1765
rect 610 -1835 670 -1805
rect 610 -1875 620 -1835
rect 660 -1875 670 -1835
rect 610 -1905 670 -1875
rect 610 -1945 620 -1905
rect 660 -1945 670 -1905
rect 610 -1975 670 -1945
rect 610 -2015 620 -1975
rect 660 -2015 670 -1975
rect 610 -2040 670 -2015
rect 610 -2080 620 -2040
rect 660 -2080 670 -2040
rect 610 -2100 670 -2080
rect 610 -2140 620 -2100
rect 660 -2140 670 -2100
rect 610 -2165 670 -2140
rect 610 -2205 620 -2165
rect 660 -2205 670 -2165
rect 610 -2235 670 -2205
rect 610 -2275 620 -2235
rect 660 -2275 670 -2235
rect 610 -2305 670 -2275
rect 610 -2345 620 -2305
rect 660 -2345 670 -2305
rect 610 -2375 670 -2345
rect 610 -2415 620 -2375
rect 660 -2415 670 -2375
rect 610 -2440 670 -2415
rect 610 -2480 620 -2440
rect 660 -2480 670 -2440
rect 610 -2500 670 -2480
rect 610 -2540 620 -2500
rect 660 -2540 670 -2500
rect 610 -2565 670 -2540
rect 610 -2605 620 -2565
rect 660 -2605 670 -2565
rect 610 -2635 670 -2605
rect 610 -2675 620 -2635
rect 660 -2675 670 -2635
rect 610 -2705 670 -2675
rect 610 -2745 620 -2705
rect 660 -2745 670 -2705
rect 610 -2775 670 -2745
rect 610 -2815 620 -2775
rect 660 -2815 670 -2775
rect 610 -2840 670 -2815
rect 610 -2880 620 -2840
rect 660 -2880 670 -2840
rect 610 -2890 670 -2880
rect 960 -1300 1020 -1290
rect 960 -1340 970 -1300
rect 1010 -1340 1020 -1300
rect 960 -1365 1020 -1340
rect 960 -1405 970 -1365
rect 1010 -1405 1020 -1365
rect 960 -1435 1020 -1405
rect 960 -1475 970 -1435
rect 1010 -1475 1020 -1435
rect 960 -1505 1020 -1475
rect 960 -1545 970 -1505
rect 1010 -1545 1020 -1505
rect 960 -1575 1020 -1545
rect 960 -1615 970 -1575
rect 1010 -1615 1020 -1575
rect 960 -1640 1020 -1615
rect 960 -1680 970 -1640
rect 1010 -1680 1020 -1640
rect 960 -1700 1020 -1680
rect 960 -1740 970 -1700
rect 1010 -1740 1020 -1700
rect 960 -1765 1020 -1740
rect 960 -1805 970 -1765
rect 1010 -1805 1020 -1765
rect 960 -1835 1020 -1805
rect 960 -1875 970 -1835
rect 1010 -1875 1020 -1835
rect 960 -1905 1020 -1875
rect 960 -1945 970 -1905
rect 1010 -1945 1020 -1905
rect 960 -1975 1020 -1945
rect 960 -2015 970 -1975
rect 1010 -2015 1020 -1975
rect 960 -2040 1020 -2015
rect 960 -2080 970 -2040
rect 1010 -2080 1020 -2040
rect 960 -2100 1020 -2080
rect 960 -2140 970 -2100
rect 1010 -2140 1020 -2100
rect 960 -2165 1020 -2140
rect 960 -2205 970 -2165
rect 1010 -2205 1020 -2165
rect 960 -2235 1020 -2205
rect 960 -2275 970 -2235
rect 1010 -2275 1020 -2235
rect 960 -2305 1020 -2275
rect 960 -2345 970 -2305
rect 1010 -2345 1020 -2305
rect 960 -2375 1020 -2345
rect 960 -2415 970 -2375
rect 1010 -2415 1020 -2375
rect 960 -2440 1020 -2415
rect 960 -2480 970 -2440
rect 1010 -2480 1020 -2440
rect 960 -2500 1020 -2480
rect 960 -2540 970 -2500
rect 1010 -2540 1020 -2500
rect 960 -2565 1020 -2540
rect 960 -2605 970 -2565
rect 1010 -2605 1020 -2565
rect 960 -2635 1020 -2605
rect 960 -2675 970 -2635
rect 1010 -2675 1020 -2635
rect 960 -2705 1020 -2675
rect 960 -2745 970 -2705
rect 1010 -2745 1020 -2705
rect 960 -2775 1020 -2745
rect 960 -2815 970 -2775
rect 1010 -2815 1020 -2775
rect 960 -2840 1020 -2815
rect 960 -2880 970 -2840
rect 1010 -2880 1020 -2840
rect 960 -2890 1020 -2880
rect 1310 -1300 1370 -1290
rect 1310 -1340 1320 -1300
rect 1360 -1340 1370 -1300
rect 1310 -1365 1370 -1340
rect 1310 -1405 1320 -1365
rect 1360 -1405 1370 -1365
rect 1310 -1435 1370 -1405
rect 1310 -1475 1320 -1435
rect 1360 -1475 1370 -1435
rect 1310 -1505 1370 -1475
rect 1310 -1545 1320 -1505
rect 1360 -1545 1370 -1505
rect 1310 -1575 1370 -1545
rect 1310 -1615 1320 -1575
rect 1360 -1615 1370 -1575
rect 1310 -1640 1370 -1615
rect 1310 -1680 1320 -1640
rect 1360 -1680 1370 -1640
rect 1310 -1700 1370 -1680
rect 1310 -1740 1320 -1700
rect 1360 -1740 1370 -1700
rect 1310 -1765 1370 -1740
rect 1310 -1805 1320 -1765
rect 1360 -1805 1370 -1765
rect 1310 -1835 1370 -1805
rect 1310 -1875 1320 -1835
rect 1360 -1875 1370 -1835
rect 1310 -1905 1370 -1875
rect 1310 -1945 1320 -1905
rect 1360 -1945 1370 -1905
rect 1310 -1975 1370 -1945
rect 1310 -2015 1320 -1975
rect 1360 -2015 1370 -1975
rect 1310 -2040 1370 -2015
rect 1310 -2080 1320 -2040
rect 1360 -2080 1370 -2040
rect 1310 -2100 1370 -2080
rect 1310 -2140 1320 -2100
rect 1360 -2140 1370 -2100
rect 1310 -2165 1370 -2140
rect 1310 -2205 1320 -2165
rect 1360 -2205 1370 -2165
rect 1310 -2235 1370 -2205
rect 1310 -2275 1320 -2235
rect 1360 -2275 1370 -2235
rect 1310 -2305 1370 -2275
rect 1310 -2345 1320 -2305
rect 1360 -2345 1370 -2305
rect 1310 -2375 1370 -2345
rect 1310 -2415 1320 -2375
rect 1360 -2415 1370 -2375
rect 1310 -2440 1370 -2415
rect 1310 -2480 1320 -2440
rect 1360 -2480 1370 -2440
rect 1310 -2500 1370 -2480
rect 1310 -2540 1320 -2500
rect 1360 -2540 1370 -2500
rect 1310 -2565 1370 -2540
rect 1310 -2605 1320 -2565
rect 1360 -2605 1370 -2565
rect 1310 -2635 1370 -2605
rect 1310 -2675 1320 -2635
rect 1360 -2675 1370 -2635
rect 1310 -2705 1370 -2675
rect 1310 -2745 1320 -2705
rect 1360 -2745 1370 -2705
rect 1310 -2775 1370 -2745
rect 1310 -2815 1320 -2775
rect 1360 -2815 1370 -2775
rect 1310 -2840 1370 -2815
rect 1310 -2880 1320 -2840
rect 1360 -2880 1370 -2840
rect 1310 -2890 1370 -2880
rect 1660 -1300 1720 -1290
rect 1660 -1340 1670 -1300
rect 1710 -1340 1720 -1300
rect 1660 -1365 1720 -1340
rect 1660 -1405 1670 -1365
rect 1710 -1405 1720 -1365
rect 1660 -1435 1720 -1405
rect 1660 -1475 1670 -1435
rect 1710 -1475 1720 -1435
rect 1660 -1505 1720 -1475
rect 1660 -1545 1670 -1505
rect 1710 -1545 1720 -1505
rect 1660 -1575 1720 -1545
rect 1660 -1615 1670 -1575
rect 1710 -1615 1720 -1575
rect 1660 -1640 1720 -1615
rect 1660 -1680 1670 -1640
rect 1710 -1680 1720 -1640
rect 1660 -1700 1720 -1680
rect 1660 -1740 1670 -1700
rect 1710 -1740 1720 -1700
rect 1660 -1765 1720 -1740
rect 1660 -1805 1670 -1765
rect 1710 -1805 1720 -1765
rect 1660 -1835 1720 -1805
rect 1660 -1875 1670 -1835
rect 1710 -1875 1720 -1835
rect 1660 -1905 1720 -1875
rect 1660 -1945 1670 -1905
rect 1710 -1945 1720 -1905
rect 1660 -1975 1720 -1945
rect 1660 -2015 1670 -1975
rect 1710 -2015 1720 -1975
rect 1660 -2040 1720 -2015
rect 1660 -2080 1670 -2040
rect 1710 -2080 1720 -2040
rect 1660 -2100 1720 -2080
rect 1660 -2140 1670 -2100
rect 1710 -2140 1720 -2100
rect 1660 -2165 1720 -2140
rect 1660 -2205 1670 -2165
rect 1710 -2205 1720 -2165
rect 1660 -2235 1720 -2205
rect 1660 -2275 1670 -2235
rect 1710 -2275 1720 -2235
rect 1660 -2305 1720 -2275
rect 1660 -2345 1670 -2305
rect 1710 -2345 1720 -2305
rect 1660 -2375 1720 -2345
rect 1660 -2415 1670 -2375
rect 1710 -2415 1720 -2375
rect 1660 -2440 1720 -2415
rect 1660 -2480 1670 -2440
rect 1710 -2480 1720 -2440
rect 1660 -2500 1720 -2480
rect 1660 -2540 1670 -2500
rect 1710 -2540 1720 -2500
rect 1660 -2565 1720 -2540
rect 1660 -2605 1670 -2565
rect 1710 -2605 1720 -2565
rect 1660 -2635 1720 -2605
rect 1660 -2675 1670 -2635
rect 1710 -2675 1720 -2635
rect 1660 -2705 1720 -2675
rect 1660 -2745 1670 -2705
rect 1710 -2745 1720 -2705
rect 1660 -2775 1720 -2745
rect 1660 -2815 1670 -2775
rect 1710 -2815 1720 -2775
rect 1660 -2840 1720 -2815
rect 1660 -2880 1670 -2840
rect 1710 -2880 1720 -2840
rect 1660 -2890 1720 -2880
rect 2010 -1300 2070 -1290
rect 2010 -1340 2020 -1300
rect 2060 -1340 2070 -1300
rect 2010 -1365 2070 -1340
rect 2010 -1405 2020 -1365
rect 2060 -1405 2070 -1365
rect 2010 -1435 2070 -1405
rect 2010 -1475 2020 -1435
rect 2060 -1475 2070 -1435
rect 2010 -1505 2070 -1475
rect 2010 -1545 2020 -1505
rect 2060 -1545 2070 -1505
rect 2010 -1575 2070 -1545
rect 2010 -1615 2020 -1575
rect 2060 -1615 2070 -1575
rect 2010 -1640 2070 -1615
rect 2010 -1680 2020 -1640
rect 2060 -1680 2070 -1640
rect 2010 -1700 2070 -1680
rect 2010 -1740 2020 -1700
rect 2060 -1740 2070 -1700
rect 2010 -1765 2070 -1740
rect 2010 -1805 2020 -1765
rect 2060 -1805 2070 -1765
rect 2010 -1835 2070 -1805
rect 2010 -1875 2020 -1835
rect 2060 -1875 2070 -1835
rect 2010 -1905 2070 -1875
rect 2010 -1945 2020 -1905
rect 2060 -1945 2070 -1905
rect 2010 -1975 2070 -1945
rect 2010 -2015 2020 -1975
rect 2060 -2015 2070 -1975
rect 2010 -2040 2070 -2015
rect 2010 -2080 2020 -2040
rect 2060 -2080 2070 -2040
rect 2010 -2100 2070 -2080
rect 2010 -2140 2020 -2100
rect 2060 -2140 2070 -2100
rect 2010 -2165 2070 -2140
rect 2010 -2205 2020 -2165
rect 2060 -2205 2070 -2165
rect 2010 -2235 2070 -2205
rect 2010 -2275 2020 -2235
rect 2060 -2275 2070 -2235
rect 2010 -2305 2070 -2275
rect 2010 -2345 2020 -2305
rect 2060 -2345 2070 -2305
rect 2010 -2375 2070 -2345
rect 2010 -2415 2020 -2375
rect 2060 -2415 2070 -2375
rect 2010 -2440 2070 -2415
rect 2010 -2480 2020 -2440
rect 2060 -2480 2070 -2440
rect 2010 -2500 2070 -2480
rect 2010 -2540 2020 -2500
rect 2060 -2540 2070 -2500
rect 2010 -2565 2070 -2540
rect 2010 -2605 2020 -2565
rect 2060 -2605 2070 -2565
rect 2010 -2635 2070 -2605
rect 2010 -2675 2020 -2635
rect 2060 -2675 2070 -2635
rect 2010 -2705 2070 -2675
rect 2010 -2745 2020 -2705
rect 2060 -2745 2070 -2705
rect 2010 -2775 2070 -2745
rect 2010 -2815 2020 -2775
rect 2060 -2815 2070 -2775
rect 2010 -2840 2070 -2815
rect 2010 -2880 2020 -2840
rect 2060 -2880 2070 -2840
rect 2010 -2890 2070 -2880
rect 2360 -1300 2420 -1290
rect 2360 -1340 2370 -1300
rect 2410 -1340 2420 -1300
rect 2360 -1365 2420 -1340
rect 2360 -1405 2370 -1365
rect 2410 -1405 2420 -1365
rect 2360 -1435 2420 -1405
rect 2360 -1475 2370 -1435
rect 2410 -1475 2420 -1435
rect 2360 -1505 2420 -1475
rect 2360 -1545 2370 -1505
rect 2410 -1545 2420 -1505
rect 2360 -1575 2420 -1545
rect 2360 -1615 2370 -1575
rect 2410 -1615 2420 -1575
rect 2360 -1640 2420 -1615
rect 2360 -1680 2370 -1640
rect 2410 -1680 2420 -1640
rect 2360 -1700 2420 -1680
rect 2360 -1740 2370 -1700
rect 2410 -1740 2420 -1700
rect 2360 -1765 2420 -1740
rect 2360 -1805 2370 -1765
rect 2410 -1805 2420 -1765
rect 2360 -1835 2420 -1805
rect 2360 -1875 2370 -1835
rect 2410 -1875 2420 -1835
rect 2360 -1905 2420 -1875
rect 2360 -1945 2370 -1905
rect 2410 -1945 2420 -1905
rect 2360 -1975 2420 -1945
rect 2360 -2015 2370 -1975
rect 2410 -2015 2420 -1975
rect 2360 -2040 2420 -2015
rect 2360 -2080 2370 -2040
rect 2410 -2080 2420 -2040
rect 2360 -2100 2420 -2080
rect 2360 -2140 2370 -2100
rect 2410 -2140 2420 -2100
rect 2360 -2165 2420 -2140
rect 2360 -2205 2370 -2165
rect 2410 -2205 2420 -2165
rect 2360 -2235 2420 -2205
rect 2360 -2275 2370 -2235
rect 2410 -2275 2420 -2235
rect 2360 -2305 2420 -2275
rect 2360 -2345 2370 -2305
rect 2410 -2345 2420 -2305
rect 2360 -2375 2420 -2345
rect 2360 -2415 2370 -2375
rect 2410 -2415 2420 -2375
rect 2360 -2440 2420 -2415
rect 2360 -2480 2370 -2440
rect 2410 -2480 2420 -2440
rect 2360 -2500 2420 -2480
rect 2360 -2540 2370 -2500
rect 2410 -2540 2420 -2500
rect 2360 -2565 2420 -2540
rect 2360 -2605 2370 -2565
rect 2410 -2605 2420 -2565
rect 2360 -2635 2420 -2605
rect 2360 -2675 2370 -2635
rect 2410 -2675 2420 -2635
rect 2360 -2705 2420 -2675
rect 2360 -2745 2370 -2705
rect 2410 -2745 2420 -2705
rect 2360 -2775 2420 -2745
rect 2360 -2815 2370 -2775
rect 2410 -2815 2420 -2775
rect 2360 -2840 2420 -2815
rect 2360 -2880 2370 -2840
rect 2410 -2880 2420 -2840
rect 2360 -2890 2420 -2880
rect 2710 -1300 2770 -1290
rect 2710 -1340 2720 -1300
rect 2760 -1340 2770 -1300
rect 2710 -1365 2770 -1340
rect 2710 -1405 2720 -1365
rect 2760 -1405 2770 -1365
rect 2710 -1435 2770 -1405
rect 2710 -1475 2720 -1435
rect 2760 -1475 2770 -1435
rect 2710 -1505 2770 -1475
rect 2710 -1545 2720 -1505
rect 2760 -1545 2770 -1505
rect 2710 -1575 2770 -1545
rect 2710 -1615 2720 -1575
rect 2760 -1615 2770 -1575
rect 2710 -1640 2770 -1615
rect 2710 -1680 2720 -1640
rect 2760 -1680 2770 -1640
rect 2710 -1700 2770 -1680
rect 2710 -1740 2720 -1700
rect 2760 -1740 2770 -1700
rect 2710 -1765 2770 -1740
rect 2710 -1805 2720 -1765
rect 2760 -1805 2770 -1765
rect 2710 -1835 2770 -1805
rect 2710 -1875 2720 -1835
rect 2760 -1875 2770 -1835
rect 2710 -1905 2770 -1875
rect 2710 -1945 2720 -1905
rect 2760 -1945 2770 -1905
rect 2710 -1975 2770 -1945
rect 2710 -2015 2720 -1975
rect 2760 -2015 2770 -1975
rect 2710 -2040 2770 -2015
rect 2710 -2080 2720 -2040
rect 2760 -2080 2770 -2040
rect 2710 -2100 2770 -2080
rect 2710 -2140 2720 -2100
rect 2760 -2140 2770 -2100
rect 2710 -2165 2770 -2140
rect 2710 -2205 2720 -2165
rect 2760 -2205 2770 -2165
rect 2710 -2235 2770 -2205
rect 2710 -2275 2720 -2235
rect 2760 -2275 2770 -2235
rect 2710 -2305 2770 -2275
rect 2710 -2345 2720 -2305
rect 2760 -2345 2770 -2305
rect 2710 -2375 2770 -2345
rect 2710 -2415 2720 -2375
rect 2760 -2415 2770 -2375
rect 2710 -2440 2770 -2415
rect 2710 -2480 2720 -2440
rect 2760 -2480 2770 -2440
rect 2710 -2500 2770 -2480
rect 2710 -2540 2720 -2500
rect 2760 -2540 2770 -2500
rect 2710 -2565 2770 -2540
rect 2710 -2605 2720 -2565
rect 2760 -2605 2770 -2565
rect 2710 -2635 2770 -2605
rect 2710 -2675 2720 -2635
rect 2760 -2675 2770 -2635
rect 2710 -2705 2770 -2675
rect 2710 -2745 2720 -2705
rect 2760 -2745 2770 -2705
rect 2710 -2775 2770 -2745
rect 2710 -2815 2720 -2775
rect 2760 -2815 2770 -2775
rect 2710 -2840 2770 -2815
rect 2710 -2880 2720 -2840
rect 2760 -2880 2770 -2840
rect 2710 -2890 2770 -2880
rect 3060 -1300 3120 -1290
rect 3060 -1340 3070 -1300
rect 3110 -1340 3120 -1300
rect 3060 -1365 3120 -1340
rect 3060 -1405 3070 -1365
rect 3110 -1405 3120 -1365
rect 3060 -1435 3120 -1405
rect 3060 -1475 3070 -1435
rect 3110 -1475 3120 -1435
rect 3060 -1505 3120 -1475
rect 3060 -1545 3070 -1505
rect 3110 -1545 3120 -1505
rect 3060 -1575 3120 -1545
rect 3060 -1615 3070 -1575
rect 3110 -1615 3120 -1575
rect 3060 -1640 3120 -1615
rect 3060 -1680 3070 -1640
rect 3110 -1680 3120 -1640
rect 3060 -1700 3120 -1680
rect 3060 -1740 3070 -1700
rect 3110 -1740 3120 -1700
rect 3060 -1765 3120 -1740
rect 3060 -1805 3070 -1765
rect 3110 -1805 3120 -1765
rect 3060 -1835 3120 -1805
rect 3060 -1875 3070 -1835
rect 3110 -1875 3120 -1835
rect 3060 -1905 3120 -1875
rect 3060 -1945 3070 -1905
rect 3110 -1945 3120 -1905
rect 3060 -1975 3120 -1945
rect 3060 -2015 3070 -1975
rect 3110 -2015 3120 -1975
rect 3060 -2040 3120 -2015
rect 3060 -2080 3070 -2040
rect 3110 -2080 3120 -2040
rect 3060 -2100 3120 -2080
rect 3060 -2140 3070 -2100
rect 3110 -2140 3120 -2100
rect 3060 -2165 3120 -2140
rect 3060 -2205 3070 -2165
rect 3110 -2205 3120 -2165
rect 3060 -2235 3120 -2205
rect 3060 -2275 3070 -2235
rect 3110 -2275 3120 -2235
rect 3060 -2305 3120 -2275
rect 3060 -2345 3070 -2305
rect 3110 -2345 3120 -2305
rect 3060 -2375 3120 -2345
rect 3060 -2415 3070 -2375
rect 3110 -2415 3120 -2375
rect 3060 -2440 3120 -2415
rect 3060 -2480 3070 -2440
rect 3110 -2480 3120 -2440
rect 3060 -2500 3120 -2480
rect 3060 -2540 3070 -2500
rect 3110 -2540 3120 -2500
rect 3060 -2565 3120 -2540
rect 3060 -2605 3070 -2565
rect 3110 -2605 3120 -2565
rect 3060 -2635 3120 -2605
rect 3060 -2675 3070 -2635
rect 3110 -2675 3120 -2635
rect 3060 -2705 3120 -2675
rect 3060 -2745 3070 -2705
rect 3110 -2745 3120 -2705
rect 3060 -2775 3120 -2745
rect 3060 -2815 3070 -2775
rect 3110 -2815 3120 -2775
rect 3060 -2840 3120 -2815
rect 3060 -2880 3070 -2840
rect 3110 -2880 3120 -2840
rect 3060 -2890 3120 -2880
rect 3410 -1300 3470 -1290
rect 3410 -1340 3420 -1300
rect 3460 -1340 3470 -1300
rect 3410 -1365 3470 -1340
rect 3410 -1405 3420 -1365
rect 3460 -1405 3470 -1365
rect 3410 -1435 3470 -1405
rect 3410 -1475 3420 -1435
rect 3460 -1475 3470 -1435
rect 3410 -1505 3470 -1475
rect 3410 -1545 3420 -1505
rect 3460 -1545 3470 -1505
rect 3410 -1575 3470 -1545
rect 3410 -1615 3420 -1575
rect 3460 -1615 3470 -1575
rect 3410 -1640 3470 -1615
rect 3410 -1680 3420 -1640
rect 3460 -1680 3470 -1640
rect 3410 -1700 3470 -1680
rect 3410 -1740 3420 -1700
rect 3460 -1740 3470 -1700
rect 3410 -1765 3470 -1740
rect 3410 -1805 3420 -1765
rect 3460 -1805 3470 -1765
rect 3410 -1835 3470 -1805
rect 3410 -1875 3420 -1835
rect 3460 -1875 3470 -1835
rect 3410 -1905 3470 -1875
rect 3410 -1945 3420 -1905
rect 3460 -1945 3470 -1905
rect 3410 -1975 3470 -1945
rect 3410 -2015 3420 -1975
rect 3460 -2015 3470 -1975
rect 3410 -2040 3470 -2015
rect 3410 -2080 3420 -2040
rect 3460 -2080 3470 -2040
rect 3410 -2100 3470 -2080
rect 3410 -2140 3420 -2100
rect 3460 -2140 3470 -2100
rect 3410 -2165 3470 -2140
rect 3410 -2205 3420 -2165
rect 3460 -2205 3470 -2165
rect 3410 -2235 3470 -2205
rect 3410 -2275 3420 -2235
rect 3460 -2275 3470 -2235
rect 3410 -2305 3470 -2275
rect 3410 -2345 3420 -2305
rect 3460 -2345 3470 -2305
rect 3410 -2375 3470 -2345
rect 3410 -2415 3420 -2375
rect 3460 -2415 3470 -2375
rect 3410 -2440 3470 -2415
rect 3410 -2480 3420 -2440
rect 3460 -2480 3470 -2440
rect 3410 -2500 3470 -2480
rect 3410 -2540 3420 -2500
rect 3460 -2540 3470 -2500
rect 3410 -2565 3470 -2540
rect 3410 -2605 3420 -2565
rect 3460 -2605 3470 -2565
rect 3410 -2635 3470 -2605
rect 3410 -2675 3420 -2635
rect 3460 -2675 3470 -2635
rect 3410 -2705 3470 -2675
rect 3410 -2745 3420 -2705
rect 3460 -2745 3470 -2705
rect 3410 -2775 3470 -2745
rect 3410 -2815 3420 -2775
rect 3460 -2815 3470 -2775
rect 3410 -2840 3470 -2815
rect 3410 -2880 3420 -2840
rect 3460 -2880 3470 -2840
rect 3410 -2890 3470 -2880
rect 3760 -1300 3820 -1290
rect 3760 -1340 3770 -1300
rect 3810 -1340 3820 -1300
rect 3760 -1365 3820 -1340
rect 3760 -1405 3770 -1365
rect 3810 -1405 3820 -1365
rect 3760 -1435 3820 -1405
rect 3760 -1475 3770 -1435
rect 3810 -1475 3820 -1435
rect 3760 -1505 3820 -1475
rect 3760 -1545 3770 -1505
rect 3810 -1545 3820 -1505
rect 3760 -1575 3820 -1545
rect 3760 -1615 3770 -1575
rect 3810 -1615 3820 -1575
rect 3760 -1640 3820 -1615
rect 3760 -1680 3770 -1640
rect 3810 -1680 3820 -1640
rect 3760 -1700 3820 -1680
rect 3760 -1740 3770 -1700
rect 3810 -1740 3820 -1700
rect 3760 -1765 3820 -1740
rect 3760 -1805 3770 -1765
rect 3810 -1805 3820 -1765
rect 3760 -1835 3820 -1805
rect 3760 -1875 3770 -1835
rect 3810 -1875 3820 -1835
rect 3760 -1905 3820 -1875
rect 3760 -1945 3770 -1905
rect 3810 -1945 3820 -1905
rect 3760 -1975 3820 -1945
rect 3760 -2015 3770 -1975
rect 3810 -2015 3820 -1975
rect 3760 -2040 3820 -2015
rect 3760 -2080 3770 -2040
rect 3810 -2080 3820 -2040
rect 3760 -2100 3820 -2080
rect 3760 -2140 3770 -2100
rect 3810 -2140 3820 -2100
rect 3760 -2165 3820 -2140
rect 3760 -2205 3770 -2165
rect 3810 -2205 3820 -2165
rect 3760 -2235 3820 -2205
rect 3760 -2275 3770 -2235
rect 3810 -2275 3820 -2235
rect 3760 -2305 3820 -2275
rect 3760 -2345 3770 -2305
rect 3810 -2345 3820 -2305
rect 3760 -2375 3820 -2345
rect 3760 -2415 3770 -2375
rect 3810 -2415 3820 -2375
rect 3760 -2440 3820 -2415
rect 3760 -2480 3770 -2440
rect 3810 -2480 3820 -2440
rect 3760 -2500 3820 -2480
rect 3760 -2540 3770 -2500
rect 3810 -2540 3820 -2500
rect 3760 -2565 3820 -2540
rect 3760 -2605 3770 -2565
rect 3810 -2605 3820 -2565
rect 3760 -2635 3820 -2605
rect 3760 -2675 3770 -2635
rect 3810 -2675 3820 -2635
rect 3760 -2705 3820 -2675
rect 3760 -2745 3770 -2705
rect 3810 -2745 3820 -2705
rect 3760 -2775 3820 -2745
rect 3760 -2815 3770 -2775
rect 3810 -2815 3820 -2775
rect 3760 -2840 3820 -2815
rect 3760 -2880 3770 -2840
rect 3810 -2880 3820 -2840
rect 3760 -2890 3820 -2880
rect 4110 -1300 4170 -1290
rect 4110 -1340 4120 -1300
rect 4160 -1340 4170 -1300
rect 4110 -1365 4170 -1340
rect 4110 -1405 4120 -1365
rect 4160 -1405 4170 -1365
rect 4110 -1435 4170 -1405
rect 4110 -1475 4120 -1435
rect 4160 -1475 4170 -1435
rect 4110 -1505 4170 -1475
rect 4110 -1545 4120 -1505
rect 4160 -1545 4170 -1505
rect 4110 -1575 4170 -1545
rect 4110 -1615 4120 -1575
rect 4160 -1615 4170 -1575
rect 4110 -1640 4170 -1615
rect 4110 -1680 4120 -1640
rect 4160 -1680 4170 -1640
rect 4110 -1700 4170 -1680
rect 4110 -1740 4120 -1700
rect 4160 -1740 4170 -1700
rect 4110 -1765 4170 -1740
rect 4110 -1805 4120 -1765
rect 4160 -1805 4170 -1765
rect 4110 -1835 4170 -1805
rect 4110 -1875 4120 -1835
rect 4160 -1875 4170 -1835
rect 4110 -1905 4170 -1875
rect 4110 -1945 4120 -1905
rect 4160 -1945 4170 -1905
rect 4110 -1975 4170 -1945
rect 4110 -2015 4120 -1975
rect 4160 -2015 4170 -1975
rect 4110 -2040 4170 -2015
rect 4110 -2080 4120 -2040
rect 4160 -2080 4170 -2040
rect 4110 -2100 4170 -2080
rect 4110 -2140 4120 -2100
rect 4160 -2140 4170 -2100
rect 4110 -2165 4170 -2140
rect 4110 -2205 4120 -2165
rect 4160 -2205 4170 -2165
rect 4110 -2235 4170 -2205
rect 4110 -2275 4120 -2235
rect 4160 -2275 4170 -2235
rect 4110 -2305 4170 -2275
rect 4110 -2345 4120 -2305
rect 4160 -2345 4170 -2305
rect 4110 -2375 4170 -2345
rect 4110 -2415 4120 -2375
rect 4160 -2415 4170 -2375
rect 4110 -2440 4170 -2415
rect 4110 -2480 4120 -2440
rect 4160 -2480 4170 -2440
rect 4110 -2500 4170 -2480
rect 4110 -2540 4120 -2500
rect 4160 -2540 4170 -2500
rect 4110 -2565 4170 -2540
rect 4110 -2605 4120 -2565
rect 4160 -2605 4170 -2565
rect 4110 -2635 4170 -2605
rect 4110 -2675 4120 -2635
rect 4160 -2675 4170 -2635
rect 4110 -2705 4170 -2675
rect 4110 -2745 4120 -2705
rect 4160 -2745 4170 -2705
rect 4110 -2775 4170 -2745
rect 4110 -2815 4120 -2775
rect 4160 -2815 4170 -2775
rect 4110 -2840 4170 -2815
rect 4110 -2880 4120 -2840
rect 4160 -2880 4170 -2840
rect 4110 -2890 4170 -2880
rect 4460 -1300 4520 -1290
rect 4460 -1340 4470 -1300
rect 4510 -1340 4520 -1300
rect 4460 -1365 4520 -1340
rect 4460 -1405 4470 -1365
rect 4510 -1405 4520 -1365
rect 4460 -1435 4520 -1405
rect 4460 -1475 4470 -1435
rect 4510 -1475 4520 -1435
rect 4460 -1505 4520 -1475
rect 4460 -1545 4470 -1505
rect 4510 -1545 4520 -1505
rect 4460 -1575 4520 -1545
rect 4460 -1615 4470 -1575
rect 4510 -1615 4520 -1575
rect 4460 -1640 4520 -1615
rect 4460 -1680 4470 -1640
rect 4510 -1680 4520 -1640
rect 4460 -1700 4520 -1680
rect 4460 -1740 4470 -1700
rect 4510 -1740 4520 -1700
rect 4460 -1765 4520 -1740
rect 4460 -1805 4470 -1765
rect 4510 -1805 4520 -1765
rect 4460 -1835 4520 -1805
rect 4460 -1875 4470 -1835
rect 4510 -1875 4520 -1835
rect 4460 -1905 4520 -1875
rect 4460 -1945 4470 -1905
rect 4510 -1945 4520 -1905
rect 4460 -1975 4520 -1945
rect 4460 -2015 4470 -1975
rect 4510 -2015 4520 -1975
rect 4460 -2040 4520 -2015
rect 4460 -2080 4470 -2040
rect 4510 -2080 4520 -2040
rect 4460 -2100 4520 -2080
rect 4460 -2140 4470 -2100
rect 4510 -2140 4520 -2100
rect 4460 -2165 4520 -2140
rect 4460 -2205 4470 -2165
rect 4510 -2205 4520 -2165
rect 4460 -2235 4520 -2205
rect 4460 -2275 4470 -2235
rect 4510 -2275 4520 -2235
rect 4460 -2305 4520 -2275
rect 4460 -2345 4470 -2305
rect 4510 -2345 4520 -2305
rect 4460 -2375 4520 -2345
rect 4460 -2415 4470 -2375
rect 4510 -2415 4520 -2375
rect 4460 -2440 4520 -2415
rect 4460 -2480 4470 -2440
rect 4510 -2480 4520 -2440
rect 4460 -2500 4520 -2480
rect 4460 -2540 4470 -2500
rect 4510 -2540 4520 -2500
rect 4460 -2565 4520 -2540
rect 4460 -2605 4470 -2565
rect 4510 -2605 4520 -2565
rect 4460 -2635 4520 -2605
rect 4460 -2675 4470 -2635
rect 4510 -2675 4520 -2635
rect 4460 -2705 4520 -2675
rect 4460 -2745 4470 -2705
rect 4510 -2745 4520 -2705
rect 4460 -2775 4520 -2745
rect 4460 -2815 4470 -2775
rect 4510 -2815 4520 -2775
rect 4460 -2840 4520 -2815
rect 4460 -2880 4470 -2840
rect 4510 -2880 4520 -2840
rect 4460 -2890 4520 -2880
rect 4810 -1300 4870 -1290
rect 4810 -1340 4820 -1300
rect 4860 -1340 4870 -1300
rect 4810 -1365 4870 -1340
rect 4810 -1405 4820 -1365
rect 4860 -1405 4870 -1365
rect 4810 -1435 4870 -1405
rect 4810 -1475 4820 -1435
rect 4860 -1475 4870 -1435
rect 4810 -1505 4870 -1475
rect 4810 -1545 4820 -1505
rect 4860 -1545 4870 -1505
rect 4810 -1575 4870 -1545
rect 4810 -1615 4820 -1575
rect 4860 -1615 4870 -1575
rect 4810 -1640 4870 -1615
rect 4810 -1680 4820 -1640
rect 4860 -1680 4870 -1640
rect 4810 -1700 4870 -1680
rect 4810 -1740 4820 -1700
rect 4860 -1740 4870 -1700
rect 4810 -1765 4870 -1740
rect 4810 -1805 4820 -1765
rect 4860 -1805 4870 -1765
rect 4810 -1835 4870 -1805
rect 4810 -1875 4820 -1835
rect 4860 -1875 4870 -1835
rect 4810 -1905 4870 -1875
rect 4810 -1945 4820 -1905
rect 4860 -1945 4870 -1905
rect 4810 -1975 4870 -1945
rect 4810 -2015 4820 -1975
rect 4860 -2015 4870 -1975
rect 4810 -2040 4870 -2015
rect 4810 -2080 4820 -2040
rect 4860 -2080 4870 -2040
rect 4810 -2100 4870 -2080
rect 4810 -2140 4820 -2100
rect 4860 -2140 4870 -2100
rect 4810 -2165 4870 -2140
rect 4810 -2205 4820 -2165
rect 4860 -2205 4870 -2165
rect 4810 -2235 4870 -2205
rect 4810 -2275 4820 -2235
rect 4860 -2275 4870 -2235
rect 4810 -2305 4870 -2275
rect 4810 -2345 4820 -2305
rect 4860 -2345 4870 -2305
rect 4810 -2375 4870 -2345
rect 4810 -2415 4820 -2375
rect 4860 -2415 4870 -2375
rect 4810 -2440 4870 -2415
rect 4810 -2480 4820 -2440
rect 4860 -2480 4870 -2440
rect 4810 -2500 4870 -2480
rect 4810 -2540 4820 -2500
rect 4860 -2540 4870 -2500
rect 4810 -2565 4870 -2540
rect 4810 -2605 4820 -2565
rect 4860 -2605 4870 -2565
rect 4810 -2635 4870 -2605
rect 4810 -2675 4820 -2635
rect 4860 -2675 4870 -2635
rect 4810 -2705 4870 -2675
rect 4810 -2745 4820 -2705
rect 4860 -2745 4870 -2705
rect 4810 -2775 4870 -2745
rect 4810 -2815 4820 -2775
rect 4860 -2815 4870 -2775
rect 4810 -2840 4870 -2815
rect 4810 -2880 4820 -2840
rect 4860 -2880 4870 -2840
rect 4810 -2890 4870 -2880
rect 5160 -1300 5220 -1290
rect 5160 -1340 5170 -1300
rect 5210 -1340 5220 -1300
rect 5160 -1365 5220 -1340
rect 5160 -1405 5170 -1365
rect 5210 -1405 5220 -1365
rect 5160 -1435 5220 -1405
rect 5160 -1475 5170 -1435
rect 5210 -1475 5220 -1435
rect 5160 -1505 5220 -1475
rect 5160 -1545 5170 -1505
rect 5210 -1545 5220 -1505
rect 5160 -1575 5220 -1545
rect 5160 -1615 5170 -1575
rect 5210 -1615 5220 -1575
rect 5160 -1640 5220 -1615
rect 5160 -1680 5170 -1640
rect 5210 -1680 5220 -1640
rect 5160 -1700 5220 -1680
rect 5160 -1740 5170 -1700
rect 5210 -1740 5220 -1700
rect 5160 -1765 5220 -1740
rect 5160 -1805 5170 -1765
rect 5210 -1805 5220 -1765
rect 5160 -1835 5220 -1805
rect 5160 -1875 5170 -1835
rect 5210 -1875 5220 -1835
rect 5160 -1905 5220 -1875
rect 5160 -1945 5170 -1905
rect 5210 -1945 5220 -1905
rect 5160 -1975 5220 -1945
rect 5160 -2015 5170 -1975
rect 5210 -2015 5220 -1975
rect 5160 -2040 5220 -2015
rect 5160 -2080 5170 -2040
rect 5210 -2080 5220 -2040
rect 5160 -2100 5220 -2080
rect 5160 -2140 5170 -2100
rect 5210 -2140 5220 -2100
rect 5160 -2165 5220 -2140
rect 5160 -2205 5170 -2165
rect 5210 -2205 5220 -2165
rect 5160 -2235 5220 -2205
rect 5160 -2275 5170 -2235
rect 5210 -2275 5220 -2235
rect 5160 -2305 5220 -2275
rect 5160 -2345 5170 -2305
rect 5210 -2345 5220 -2305
rect 5160 -2375 5220 -2345
rect 5160 -2415 5170 -2375
rect 5210 -2415 5220 -2375
rect 5160 -2440 5220 -2415
rect 5160 -2480 5170 -2440
rect 5210 -2480 5220 -2440
rect 5160 -2500 5220 -2480
rect 5160 -2540 5170 -2500
rect 5210 -2540 5220 -2500
rect 5160 -2565 5220 -2540
rect 5160 -2605 5170 -2565
rect 5210 -2605 5220 -2565
rect 5160 -2635 5220 -2605
rect 5160 -2675 5170 -2635
rect 5210 -2675 5220 -2635
rect 5160 -2705 5220 -2675
rect 5160 -2745 5170 -2705
rect 5210 -2745 5220 -2705
rect 5160 -2775 5220 -2745
rect 5160 -2815 5170 -2775
rect 5210 -2815 5220 -2775
rect 5160 -2840 5220 -2815
rect 5160 -2880 5170 -2840
rect 5210 -2880 5220 -2840
rect 5160 -2890 5220 -2880
rect 5510 -1300 5570 -1290
rect 5510 -1340 5520 -1300
rect 5560 -1340 5570 -1300
rect 5510 -1365 5570 -1340
rect 5510 -1405 5520 -1365
rect 5560 -1405 5570 -1365
rect 5510 -1435 5570 -1405
rect 5510 -1475 5520 -1435
rect 5560 -1475 5570 -1435
rect 5510 -1505 5570 -1475
rect 5510 -1545 5520 -1505
rect 5560 -1545 5570 -1505
rect 5510 -1575 5570 -1545
rect 5510 -1615 5520 -1575
rect 5560 -1615 5570 -1575
rect 5510 -1640 5570 -1615
rect 5510 -1680 5520 -1640
rect 5560 -1680 5570 -1640
rect 5510 -1700 5570 -1680
rect 5510 -1740 5520 -1700
rect 5560 -1740 5570 -1700
rect 5510 -1765 5570 -1740
rect 5510 -1805 5520 -1765
rect 5560 -1805 5570 -1765
rect 5510 -1835 5570 -1805
rect 5510 -1875 5520 -1835
rect 5560 -1875 5570 -1835
rect 5510 -1905 5570 -1875
rect 5510 -1945 5520 -1905
rect 5560 -1945 5570 -1905
rect 5510 -1975 5570 -1945
rect 5510 -2015 5520 -1975
rect 5560 -2015 5570 -1975
rect 5510 -2040 5570 -2015
rect 5510 -2080 5520 -2040
rect 5560 -2080 5570 -2040
rect 5510 -2100 5570 -2080
rect 5510 -2140 5520 -2100
rect 5560 -2140 5570 -2100
rect 5510 -2165 5570 -2140
rect 5510 -2205 5520 -2165
rect 5560 -2205 5570 -2165
rect 5510 -2235 5570 -2205
rect 5510 -2275 5520 -2235
rect 5560 -2275 5570 -2235
rect 5510 -2305 5570 -2275
rect 5510 -2345 5520 -2305
rect 5560 -2345 5570 -2305
rect 5510 -2375 5570 -2345
rect 5510 -2415 5520 -2375
rect 5560 -2415 5570 -2375
rect 5510 -2440 5570 -2415
rect 5510 -2480 5520 -2440
rect 5560 -2480 5570 -2440
rect 5510 -2500 5570 -2480
rect 5510 -2540 5520 -2500
rect 5560 -2540 5570 -2500
rect 5510 -2565 5570 -2540
rect 5510 -2605 5520 -2565
rect 5560 -2605 5570 -2565
rect 5510 -2635 5570 -2605
rect 5510 -2675 5520 -2635
rect 5560 -2675 5570 -2635
rect 5510 -2705 5570 -2675
rect 5510 -2745 5520 -2705
rect 5560 -2745 5570 -2705
rect 5510 -2775 5570 -2745
rect 5510 -2815 5520 -2775
rect 5560 -2815 5570 -2775
rect 5510 -2840 5570 -2815
rect 5510 -2880 5520 -2840
rect 5560 -2880 5570 -2840
rect 5510 -2890 5570 -2880
rect 5860 -1300 5920 -1290
rect 5860 -1340 5870 -1300
rect 5910 -1340 5920 -1300
rect 5860 -1365 5920 -1340
rect 5860 -1405 5870 -1365
rect 5910 -1405 5920 -1365
rect 5860 -1435 5920 -1405
rect 5860 -1475 5870 -1435
rect 5910 -1475 5920 -1435
rect 5860 -1505 5920 -1475
rect 5860 -1545 5870 -1505
rect 5910 -1545 5920 -1505
rect 5860 -1575 5920 -1545
rect 5860 -1615 5870 -1575
rect 5910 -1615 5920 -1575
rect 5860 -1640 5920 -1615
rect 5860 -1680 5870 -1640
rect 5910 -1680 5920 -1640
rect 5860 -1700 5920 -1680
rect 5860 -1740 5870 -1700
rect 5910 -1740 5920 -1700
rect 5860 -1765 5920 -1740
rect 5860 -1805 5870 -1765
rect 5910 -1805 5920 -1765
rect 5860 -1835 5920 -1805
rect 5860 -1875 5870 -1835
rect 5910 -1875 5920 -1835
rect 5860 -1905 5920 -1875
rect 5860 -1945 5870 -1905
rect 5910 -1945 5920 -1905
rect 5860 -1975 5920 -1945
rect 5860 -2015 5870 -1975
rect 5910 -2015 5920 -1975
rect 5860 -2040 5920 -2015
rect 5860 -2080 5870 -2040
rect 5910 -2080 5920 -2040
rect 5860 -2100 5920 -2080
rect 5860 -2140 5870 -2100
rect 5910 -2140 5920 -2100
rect 5860 -2165 5920 -2140
rect 5860 -2205 5870 -2165
rect 5910 -2205 5920 -2165
rect 5860 -2235 5920 -2205
rect 5860 -2275 5870 -2235
rect 5910 -2275 5920 -2235
rect 5860 -2305 5920 -2275
rect 5860 -2345 5870 -2305
rect 5910 -2345 5920 -2305
rect 5860 -2375 5920 -2345
rect 5860 -2415 5870 -2375
rect 5910 -2415 5920 -2375
rect 5860 -2440 5920 -2415
rect 5860 -2480 5870 -2440
rect 5910 -2480 5920 -2440
rect 5860 -2500 5920 -2480
rect 5860 -2540 5870 -2500
rect 5910 -2540 5920 -2500
rect 5860 -2565 5920 -2540
rect 5860 -2605 5870 -2565
rect 5910 -2605 5920 -2565
rect 5860 -2635 5920 -2605
rect 5860 -2675 5870 -2635
rect 5910 -2675 5920 -2635
rect 5860 -2705 5920 -2675
rect 5860 -2745 5870 -2705
rect 5910 -2745 5920 -2705
rect 5860 -2775 5920 -2745
rect 5860 -2815 5870 -2775
rect 5910 -2815 5920 -2775
rect 5860 -2840 5920 -2815
rect 5860 -2880 5870 -2840
rect 5910 -2880 5920 -2840
rect 5860 -2890 5920 -2880
rect 6210 -1300 6270 -1290
rect 6210 -1340 6220 -1300
rect 6260 -1340 6270 -1300
rect 6210 -1365 6270 -1340
rect 6210 -1405 6220 -1365
rect 6260 -1405 6270 -1365
rect 6210 -1435 6270 -1405
rect 6210 -1475 6220 -1435
rect 6260 -1475 6270 -1435
rect 6210 -1505 6270 -1475
rect 6210 -1545 6220 -1505
rect 6260 -1545 6270 -1505
rect 6210 -1575 6270 -1545
rect 6210 -1615 6220 -1575
rect 6260 -1615 6270 -1575
rect 6210 -1640 6270 -1615
rect 6210 -1680 6220 -1640
rect 6260 -1680 6270 -1640
rect 6210 -1700 6270 -1680
rect 6210 -1740 6220 -1700
rect 6260 -1740 6270 -1700
rect 6210 -1765 6270 -1740
rect 6210 -1805 6220 -1765
rect 6260 -1805 6270 -1765
rect 6210 -1835 6270 -1805
rect 6210 -1875 6220 -1835
rect 6260 -1875 6270 -1835
rect 6210 -1905 6270 -1875
rect 6210 -1945 6220 -1905
rect 6260 -1945 6270 -1905
rect 6210 -1975 6270 -1945
rect 6210 -2015 6220 -1975
rect 6260 -2015 6270 -1975
rect 6210 -2040 6270 -2015
rect 6210 -2080 6220 -2040
rect 6260 -2080 6270 -2040
rect 6210 -2100 6270 -2080
rect 6210 -2140 6220 -2100
rect 6260 -2140 6270 -2100
rect 6210 -2165 6270 -2140
rect 6210 -2205 6220 -2165
rect 6260 -2205 6270 -2165
rect 6210 -2235 6270 -2205
rect 6210 -2275 6220 -2235
rect 6260 -2275 6270 -2235
rect 6210 -2305 6270 -2275
rect 6210 -2345 6220 -2305
rect 6260 -2345 6270 -2305
rect 6210 -2375 6270 -2345
rect 6210 -2415 6220 -2375
rect 6260 -2415 6270 -2375
rect 6210 -2440 6270 -2415
rect 6210 -2480 6220 -2440
rect 6260 -2480 6270 -2440
rect 6210 -2500 6270 -2480
rect 6210 -2540 6220 -2500
rect 6260 -2540 6270 -2500
rect 6210 -2565 6270 -2540
rect 6210 -2605 6220 -2565
rect 6260 -2605 6270 -2565
rect 6210 -2635 6270 -2605
rect 6210 -2675 6220 -2635
rect 6260 -2675 6270 -2635
rect 6210 -2705 6270 -2675
rect 6210 -2745 6220 -2705
rect 6260 -2745 6270 -2705
rect 6210 -2775 6270 -2745
rect 6210 -2815 6220 -2775
rect 6260 -2815 6270 -2775
rect 6210 -2840 6270 -2815
rect 6210 -2880 6220 -2840
rect 6260 -2880 6270 -2840
rect 6210 -2890 6270 -2880
rect 6560 -1300 6620 -1290
rect 6560 -1340 6570 -1300
rect 6610 -1340 6620 -1300
rect 6560 -1365 6620 -1340
rect 6560 -1405 6570 -1365
rect 6610 -1405 6620 -1365
rect 6560 -1435 6620 -1405
rect 6560 -1475 6570 -1435
rect 6610 -1475 6620 -1435
rect 6560 -1505 6620 -1475
rect 6560 -1545 6570 -1505
rect 6610 -1545 6620 -1505
rect 6560 -1575 6620 -1545
rect 6560 -1615 6570 -1575
rect 6610 -1615 6620 -1575
rect 6560 -1640 6620 -1615
rect 6560 -1680 6570 -1640
rect 6610 -1680 6620 -1640
rect 6560 -1700 6620 -1680
rect 6560 -1740 6570 -1700
rect 6610 -1740 6620 -1700
rect 6560 -1765 6620 -1740
rect 6560 -1805 6570 -1765
rect 6610 -1805 6620 -1765
rect 6560 -1835 6620 -1805
rect 6560 -1875 6570 -1835
rect 6610 -1875 6620 -1835
rect 6560 -1905 6620 -1875
rect 6560 -1945 6570 -1905
rect 6610 -1945 6620 -1905
rect 6560 -1975 6620 -1945
rect 6560 -2015 6570 -1975
rect 6610 -2015 6620 -1975
rect 6560 -2040 6620 -2015
rect 6560 -2080 6570 -2040
rect 6610 -2080 6620 -2040
rect 6560 -2100 6620 -2080
rect 6560 -2140 6570 -2100
rect 6610 -2140 6620 -2100
rect 6560 -2165 6620 -2140
rect 6560 -2205 6570 -2165
rect 6610 -2205 6620 -2165
rect 6560 -2235 6620 -2205
rect 6560 -2275 6570 -2235
rect 6610 -2275 6620 -2235
rect 6560 -2305 6620 -2275
rect 6560 -2345 6570 -2305
rect 6610 -2345 6620 -2305
rect 6560 -2375 6620 -2345
rect 6560 -2415 6570 -2375
rect 6610 -2415 6620 -2375
rect 6560 -2440 6620 -2415
rect 6560 -2480 6570 -2440
rect 6610 -2480 6620 -2440
rect 6560 -2500 6620 -2480
rect 6560 -2540 6570 -2500
rect 6610 -2540 6620 -2500
rect 6560 -2565 6620 -2540
rect 6560 -2605 6570 -2565
rect 6610 -2605 6620 -2565
rect 6560 -2635 6620 -2605
rect 6560 -2675 6570 -2635
rect 6610 -2675 6620 -2635
rect 6560 -2705 6620 -2675
rect 6560 -2745 6570 -2705
rect 6610 -2745 6620 -2705
rect 6560 -2775 6620 -2745
rect 6560 -2815 6570 -2775
rect 6610 -2815 6620 -2775
rect 6560 -2840 6620 -2815
rect 6560 -2880 6570 -2840
rect 6610 -2880 6620 -2840
rect 6560 -2890 6620 -2880
rect 6910 -1300 6970 -1290
rect 6910 -1340 6920 -1300
rect 6960 -1340 6970 -1300
rect 6910 -1365 6970 -1340
rect 6910 -1405 6920 -1365
rect 6960 -1405 6970 -1365
rect 6910 -1435 6970 -1405
rect 6910 -1475 6920 -1435
rect 6960 -1475 6970 -1435
rect 6910 -1505 6970 -1475
rect 6910 -1545 6920 -1505
rect 6960 -1545 6970 -1505
rect 6910 -1575 6970 -1545
rect 6910 -1615 6920 -1575
rect 6960 -1615 6970 -1575
rect 6910 -1640 6970 -1615
rect 6910 -1680 6920 -1640
rect 6960 -1680 6970 -1640
rect 6910 -1700 6970 -1680
rect 6910 -1740 6920 -1700
rect 6960 -1740 6970 -1700
rect 6910 -1765 6970 -1740
rect 6910 -1805 6920 -1765
rect 6960 -1805 6970 -1765
rect 6910 -1835 6970 -1805
rect 6910 -1875 6920 -1835
rect 6960 -1875 6970 -1835
rect 6910 -1905 6970 -1875
rect 6910 -1945 6920 -1905
rect 6960 -1945 6970 -1905
rect 6910 -1975 6970 -1945
rect 6910 -2015 6920 -1975
rect 6960 -2015 6970 -1975
rect 6910 -2040 6970 -2015
rect 6910 -2080 6920 -2040
rect 6960 -2080 6970 -2040
rect 6910 -2100 6970 -2080
rect 6910 -2140 6920 -2100
rect 6960 -2140 6970 -2100
rect 6910 -2165 6970 -2140
rect 6910 -2205 6920 -2165
rect 6960 -2205 6970 -2165
rect 6910 -2235 6970 -2205
rect 6910 -2275 6920 -2235
rect 6960 -2275 6970 -2235
rect 6910 -2305 6970 -2275
rect 6910 -2345 6920 -2305
rect 6960 -2345 6970 -2305
rect 6910 -2375 6970 -2345
rect 6910 -2415 6920 -2375
rect 6960 -2415 6970 -2375
rect 6910 -2440 6970 -2415
rect 6910 -2480 6920 -2440
rect 6960 -2480 6970 -2440
rect 6910 -2500 6970 -2480
rect 6910 -2540 6920 -2500
rect 6960 -2540 6970 -2500
rect 6910 -2565 6970 -2540
rect 6910 -2605 6920 -2565
rect 6960 -2605 6970 -2565
rect 6910 -2635 6970 -2605
rect 6910 -2675 6920 -2635
rect 6960 -2675 6970 -2635
rect 6910 -2705 6970 -2675
rect 6910 -2745 6920 -2705
rect 6960 -2745 6970 -2705
rect 6910 -2775 6970 -2745
rect 6910 -2815 6920 -2775
rect 6960 -2815 6970 -2775
rect 6910 -2840 6970 -2815
rect 6910 -2880 6920 -2840
rect 6960 -2880 6970 -2840
rect 6910 -2890 6970 -2880
rect 7260 -1300 7320 -1290
rect 7260 -1340 7270 -1300
rect 7310 -1340 7320 -1300
rect 7260 -1365 7320 -1340
rect 7260 -1405 7270 -1365
rect 7310 -1405 7320 -1365
rect 7260 -1435 7320 -1405
rect 7260 -1475 7270 -1435
rect 7310 -1475 7320 -1435
rect 7260 -1505 7320 -1475
rect 7260 -1545 7270 -1505
rect 7310 -1545 7320 -1505
rect 7260 -1575 7320 -1545
rect 7260 -1615 7270 -1575
rect 7310 -1615 7320 -1575
rect 7260 -1640 7320 -1615
rect 7260 -1680 7270 -1640
rect 7310 -1680 7320 -1640
rect 7260 -1700 7320 -1680
rect 7260 -1740 7270 -1700
rect 7310 -1740 7320 -1700
rect 7260 -1765 7320 -1740
rect 7260 -1805 7270 -1765
rect 7310 -1805 7320 -1765
rect 7260 -1835 7320 -1805
rect 7260 -1875 7270 -1835
rect 7310 -1875 7320 -1835
rect 7260 -1905 7320 -1875
rect 7260 -1945 7270 -1905
rect 7310 -1945 7320 -1905
rect 7260 -1975 7320 -1945
rect 7260 -2015 7270 -1975
rect 7310 -2015 7320 -1975
rect 7260 -2040 7320 -2015
rect 7260 -2080 7270 -2040
rect 7310 -2080 7320 -2040
rect 7260 -2100 7320 -2080
rect 7260 -2140 7270 -2100
rect 7310 -2140 7320 -2100
rect 7260 -2165 7320 -2140
rect 7260 -2205 7270 -2165
rect 7310 -2205 7320 -2165
rect 7260 -2235 7320 -2205
rect 7260 -2275 7270 -2235
rect 7310 -2275 7320 -2235
rect 7260 -2305 7320 -2275
rect 7260 -2345 7270 -2305
rect 7310 -2345 7320 -2305
rect 7260 -2375 7320 -2345
rect 7260 -2415 7270 -2375
rect 7310 -2415 7320 -2375
rect 7260 -2440 7320 -2415
rect 7260 -2480 7270 -2440
rect 7310 -2480 7320 -2440
rect 7260 -2500 7320 -2480
rect 7260 -2540 7270 -2500
rect 7310 -2540 7320 -2500
rect 7260 -2565 7320 -2540
rect 7260 -2605 7270 -2565
rect 7310 -2605 7320 -2565
rect 7260 -2635 7320 -2605
rect 7260 -2675 7270 -2635
rect 7310 -2675 7320 -2635
rect 7260 -2705 7320 -2675
rect 7260 -2745 7270 -2705
rect 7310 -2745 7320 -2705
rect 7260 -2775 7320 -2745
rect 7260 -2815 7270 -2775
rect 7310 -2815 7320 -2775
rect 7260 -2840 7320 -2815
rect 7260 -2880 7270 -2840
rect 7310 -2880 7320 -2840
rect 7260 -2890 7320 -2880
rect 7610 -1300 7670 -1290
rect 7610 -1340 7620 -1300
rect 7660 -1340 7670 -1300
rect 7610 -1365 7670 -1340
rect 7610 -1405 7620 -1365
rect 7660 -1405 7670 -1365
rect 7610 -1435 7670 -1405
rect 7610 -1475 7620 -1435
rect 7660 -1475 7670 -1435
rect 7610 -1505 7670 -1475
rect 7610 -1545 7620 -1505
rect 7660 -1545 7670 -1505
rect 7610 -1575 7670 -1545
rect 7610 -1615 7620 -1575
rect 7660 -1615 7670 -1575
rect 7610 -1640 7670 -1615
rect 7610 -1680 7620 -1640
rect 7660 -1680 7670 -1640
rect 7610 -1700 7670 -1680
rect 7610 -1740 7620 -1700
rect 7660 -1740 7670 -1700
rect 7610 -1765 7670 -1740
rect 7610 -1805 7620 -1765
rect 7660 -1805 7670 -1765
rect 7610 -1835 7670 -1805
rect 7610 -1875 7620 -1835
rect 7660 -1875 7670 -1835
rect 7610 -1905 7670 -1875
rect 7610 -1945 7620 -1905
rect 7660 -1945 7670 -1905
rect 7610 -1975 7670 -1945
rect 7610 -2015 7620 -1975
rect 7660 -2015 7670 -1975
rect 7610 -2040 7670 -2015
rect 7610 -2080 7620 -2040
rect 7660 -2080 7670 -2040
rect 7610 -2100 7670 -2080
rect 7610 -2140 7620 -2100
rect 7660 -2140 7670 -2100
rect 7610 -2165 7670 -2140
rect 7610 -2205 7620 -2165
rect 7660 -2205 7670 -2165
rect 7610 -2235 7670 -2205
rect 7610 -2275 7620 -2235
rect 7660 -2275 7670 -2235
rect 7610 -2305 7670 -2275
rect 7610 -2345 7620 -2305
rect 7660 -2345 7670 -2305
rect 7610 -2375 7670 -2345
rect 7610 -2415 7620 -2375
rect 7660 -2415 7670 -2375
rect 7610 -2440 7670 -2415
rect 7610 -2480 7620 -2440
rect 7660 -2480 7670 -2440
rect 7610 -2500 7670 -2480
rect 7610 -2540 7620 -2500
rect 7660 -2540 7670 -2500
rect 7610 -2565 7670 -2540
rect 7610 -2605 7620 -2565
rect 7660 -2605 7670 -2565
rect 7610 -2635 7670 -2605
rect 7610 -2675 7620 -2635
rect 7660 -2675 7670 -2635
rect 7610 -2705 7670 -2675
rect 7610 -2745 7620 -2705
rect 7660 -2745 7670 -2705
rect 7610 -2775 7670 -2745
rect 7610 -2815 7620 -2775
rect 7660 -2815 7670 -2775
rect 7610 -2840 7670 -2815
rect 7610 -2880 7620 -2840
rect 7660 -2880 7670 -2840
rect 7610 -2890 7670 -2880
rect 7960 -1300 8020 -1290
rect 7960 -1340 7970 -1300
rect 8010 -1340 8020 -1300
rect 7960 -1365 8020 -1340
rect 7960 -1405 7970 -1365
rect 8010 -1405 8020 -1365
rect 7960 -1435 8020 -1405
rect 7960 -1475 7970 -1435
rect 8010 -1475 8020 -1435
rect 7960 -1505 8020 -1475
rect 7960 -1545 7970 -1505
rect 8010 -1545 8020 -1505
rect 7960 -1575 8020 -1545
rect 7960 -1615 7970 -1575
rect 8010 -1615 8020 -1575
rect 7960 -1640 8020 -1615
rect 7960 -1680 7970 -1640
rect 8010 -1680 8020 -1640
rect 7960 -1700 8020 -1680
rect 7960 -1740 7970 -1700
rect 8010 -1740 8020 -1700
rect 7960 -1765 8020 -1740
rect 7960 -1805 7970 -1765
rect 8010 -1805 8020 -1765
rect 7960 -1835 8020 -1805
rect 7960 -1875 7970 -1835
rect 8010 -1875 8020 -1835
rect 7960 -1905 8020 -1875
rect 7960 -1945 7970 -1905
rect 8010 -1945 8020 -1905
rect 7960 -1975 8020 -1945
rect 7960 -2015 7970 -1975
rect 8010 -2015 8020 -1975
rect 7960 -2040 8020 -2015
rect 7960 -2080 7970 -2040
rect 8010 -2080 8020 -2040
rect 7960 -2100 8020 -2080
rect 7960 -2140 7970 -2100
rect 8010 -2140 8020 -2100
rect 7960 -2165 8020 -2140
rect 7960 -2205 7970 -2165
rect 8010 -2205 8020 -2165
rect 7960 -2235 8020 -2205
rect 7960 -2275 7970 -2235
rect 8010 -2275 8020 -2235
rect 7960 -2305 8020 -2275
rect 7960 -2345 7970 -2305
rect 8010 -2345 8020 -2305
rect 7960 -2375 8020 -2345
rect 7960 -2415 7970 -2375
rect 8010 -2415 8020 -2375
rect 7960 -2440 8020 -2415
rect 7960 -2480 7970 -2440
rect 8010 -2480 8020 -2440
rect 7960 -2500 8020 -2480
rect 7960 -2540 7970 -2500
rect 8010 -2540 8020 -2500
rect 7960 -2565 8020 -2540
rect 7960 -2605 7970 -2565
rect 8010 -2605 8020 -2565
rect 7960 -2635 8020 -2605
rect 7960 -2675 7970 -2635
rect 8010 -2675 8020 -2635
rect 7960 -2705 8020 -2675
rect 7960 -2745 7970 -2705
rect 8010 -2745 8020 -2705
rect 7960 -2775 8020 -2745
rect 7960 -2815 7970 -2775
rect 8010 -2815 8020 -2775
rect 7960 -2840 8020 -2815
rect 7960 -2880 7970 -2840
rect 8010 -2880 8020 -2840
rect 7960 -2890 8020 -2880
rect 8310 -1300 8370 -1290
rect 8310 -1340 8320 -1300
rect 8360 -1340 8370 -1300
rect 8310 -1365 8370 -1340
rect 8310 -1405 8320 -1365
rect 8360 -1405 8370 -1365
rect 8310 -1435 8370 -1405
rect 8310 -1475 8320 -1435
rect 8360 -1475 8370 -1435
rect 8310 -1505 8370 -1475
rect 8310 -1545 8320 -1505
rect 8360 -1545 8370 -1505
rect 8310 -1575 8370 -1545
rect 8310 -1615 8320 -1575
rect 8360 -1615 8370 -1575
rect 8310 -1640 8370 -1615
rect 8310 -1680 8320 -1640
rect 8360 -1680 8370 -1640
rect 8310 -1700 8370 -1680
rect 8310 -1740 8320 -1700
rect 8360 -1740 8370 -1700
rect 8310 -1765 8370 -1740
rect 8310 -1805 8320 -1765
rect 8360 -1805 8370 -1765
rect 8310 -1835 8370 -1805
rect 8310 -1875 8320 -1835
rect 8360 -1875 8370 -1835
rect 8310 -1905 8370 -1875
rect 8310 -1945 8320 -1905
rect 8360 -1945 8370 -1905
rect 8310 -1975 8370 -1945
rect 8310 -2015 8320 -1975
rect 8360 -2015 8370 -1975
rect 8310 -2040 8370 -2015
rect 8310 -2080 8320 -2040
rect 8360 -2080 8370 -2040
rect 8310 -2100 8370 -2080
rect 8310 -2140 8320 -2100
rect 8360 -2140 8370 -2100
rect 8310 -2165 8370 -2140
rect 8310 -2205 8320 -2165
rect 8360 -2205 8370 -2165
rect 8310 -2235 8370 -2205
rect 8310 -2275 8320 -2235
rect 8360 -2275 8370 -2235
rect 8310 -2305 8370 -2275
rect 8310 -2345 8320 -2305
rect 8360 -2345 8370 -2305
rect 8310 -2375 8370 -2345
rect 8310 -2415 8320 -2375
rect 8360 -2415 8370 -2375
rect 8310 -2440 8370 -2415
rect 8310 -2480 8320 -2440
rect 8360 -2480 8370 -2440
rect 8310 -2500 8370 -2480
rect 8310 -2540 8320 -2500
rect 8360 -2540 8370 -2500
rect 8310 -2565 8370 -2540
rect 8310 -2605 8320 -2565
rect 8360 -2605 8370 -2565
rect 8310 -2635 8370 -2605
rect 8310 -2675 8320 -2635
rect 8360 -2675 8370 -2635
rect 8310 -2705 8370 -2675
rect 8310 -2745 8320 -2705
rect 8360 -2745 8370 -2705
rect 8310 -2775 8370 -2745
rect 8310 -2815 8320 -2775
rect 8360 -2815 8370 -2775
rect 8310 -2840 8370 -2815
rect 8310 -2880 8320 -2840
rect 8360 -2880 8370 -2840
rect 8310 -2890 8370 -2880
rect 8660 -1305 8720 -1290
rect 8660 -1335 8675 -1305
rect 8705 -1335 8720 -1305
rect 8660 -1370 8720 -1335
rect 8660 -1400 8675 -1370
rect 8705 -1400 8720 -1370
rect 8660 -1440 8720 -1400
rect 8660 -1470 8675 -1440
rect 8705 -1470 8720 -1440
rect 8660 -1510 8720 -1470
rect 8660 -1540 8675 -1510
rect 8705 -1540 8720 -1510
rect 8660 -1580 8720 -1540
rect 8660 -1610 8675 -1580
rect 8705 -1610 8720 -1580
rect 8660 -1645 8720 -1610
rect 8660 -1675 8675 -1645
rect 8705 -1675 8720 -1645
rect 8660 -1705 8720 -1675
rect 8660 -1735 8675 -1705
rect 8705 -1735 8720 -1705
rect 8660 -1770 8720 -1735
rect 8660 -1800 8675 -1770
rect 8705 -1800 8720 -1770
rect 8660 -1840 8720 -1800
rect 8660 -1870 8675 -1840
rect 8705 -1870 8720 -1840
rect 8660 -1910 8720 -1870
rect 8660 -1940 8675 -1910
rect 8705 -1940 8720 -1910
rect 8660 -1980 8720 -1940
rect 8660 -2010 8675 -1980
rect 8705 -2010 8720 -1980
rect 8660 -2045 8720 -2010
rect 8660 -2075 8675 -2045
rect 8705 -2075 8720 -2045
rect 8660 -2105 8720 -2075
rect 8660 -2135 8675 -2105
rect 8705 -2135 8720 -2105
rect 8660 -2170 8720 -2135
rect 8660 -2200 8675 -2170
rect 8705 -2200 8720 -2170
rect 8660 -2240 8720 -2200
rect 8660 -2270 8675 -2240
rect 8705 -2270 8720 -2240
rect 8660 -2310 8720 -2270
rect 8660 -2340 8675 -2310
rect 8705 -2340 8720 -2310
rect 8660 -2380 8720 -2340
rect 8660 -2410 8675 -2380
rect 8705 -2410 8720 -2380
rect 8660 -2445 8720 -2410
rect 8660 -2475 8675 -2445
rect 8705 -2475 8720 -2445
rect 8660 -2505 8720 -2475
rect 8660 -2535 8675 -2505
rect 8705 -2535 8720 -2505
rect 8660 -2570 8720 -2535
rect 8660 -2600 8675 -2570
rect 8705 -2600 8720 -2570
rect 8660 -2640 8720 -2600
rect 8660 -2670 8675 -2640
rect 8705 -2670 8720 -2640
rect 8660 -2710 8720 -2670
rect 8660 -2740 8675 -2710
rect 8705 -2740 8720 -2710
rect 8660 -2780 8720 -2740
rect 8660 -2810 8675 -2780
rect 8705 -2810 8720 -2780
rect 8660 -2845 8720 -2810
rect 8660 -2875 8675 -2845
rect 8705 -2875 8720 -2845
rect 8660 -2890 8720 -2875
rect 9010 -1305 9070 -1290
rect 9010 -1335 9025 -1305
rect 9055 -1335 9070 -1305
rect 9010 -1370 9070 -1335
rect 9010 -1400 9025 -1370
rect 9055 -1400 9070 -1370
rect 9010 -1440 9070 -1400
rect 9010 -1470 9025 -1440
rect 9055 -1470 9070 -1440
rect 9010 -1510 9070 -1470
rect 9010 -1540 9025 -1510
rect 9055 -1540 9070 -1510
rect 9010 -1580 9070 -1540
rect 9010 -1610 9025 -1580
rect 9055 -1610 9070 -1580
rect 9010 -1645 9070 -1610
rect 9010 -1675 9025 -1645
rect 9055 -1675 9070 -1645
rect 9010 -1705 9070 -1675
rect 9010 -1735 9025 -1705
rect 9055 -1735 9070 -1705
rect 9010 -1770 9070 -1735
rect 9010 -1800 9025 -1770
rect 9055 -1800 9070 -1770
rect 9010 -1840 9070 -1800
rect 9010 -1870 9025 -1840
rect 9055 -1870 9070 -1840
rect 9010 -1910 9070 -1870
rect 9010 -1940 9025 -1910
rect 9055 -1940 9070 -1910
rect 9010 -1980 9070 -1940
rect 9010 -2010 9025 -1980
rect 9055 -2010 9070 -1980
rect 9010 -2045 9070 -2010
rect 9010 -2075 9025 -2045
rect 9055 -2075 9070 -2045
rect 9010 -2105 9070 -2075
rect 9010 -2135 9025 -2105
rect 9055 -2135 9070 -2105
rect 9010 -2170 9070 -2135
rect 9010 -2200 9025 -2170
rect 9055 -2200 9070 -2170
rect 9010 -2240 9070 -2200
rect 9010 -2270 9025 -2240
rect 9055 -2270 9070 -2240
rect 9010 -2310 9070 -2270
rect 9010 -2340 9025 -2310
rect 9055 -2340 9070 -2310
rect 9010 -2380 9070 -2340
rect 9010 -2410 9025 -2380
rect 9055 -2410 9070 -2380
rect 9010 -2445 9070 -2410
rect 9010 -2475 9025 -2445
rect 9055 -2475 9070 -2445
rect 9010 -2505 9070 -2475
rect 9010 -2535 9025 -2505
rect 9055 -2535 9070 -2505
rect 9010 -2570 9070 -2535
rect 9010 -2600 9025 -2570
rect 9055 -2600 9070 -2570
rect 9010 -2640 9070 -2600
rect 9010 -2670 9025 -2640
rect 9055 -2670 9070 -2640
rect 9010 -2710 9070 -2670
rect 9010 -2740 9025 -2710
rect 9055 -2740 9070 -2710
rect 9010 -2780 9070 -2740
rect 9010 -2810 9025 -2780
rect 9055 -2810 9070 -2780
rect 9010 -2845 9070 -2810
rect 9010 -2875 9025 -2845
rect 9055 -2875 9070 -2845
rect 9010 -2890 9070 -2875
rect 31290 -1310 32890 6465
rect 31290 -1345 31305 -1310
rect 31340 -1345 31350 -1310
rect 31385 -1345 31395 -1310
rect 31430 -1345 31440 -1310
rect 31475 -1345 31485 -1310
rect 31520 -1345 31530 -1310
rect 31565 -1345 31575 -1310
rect 31610 -1345 31620 -1310
rect 31655 -1345 31665 -1310
rect 31700 -1345 31710 -1310
rect 31745 -1345 31755 -1310
rect 31790 -1345 31800 -1310
rect 31835 -1345 31845 -1310
rect 31880 -1345 31890 -1310
rect 31925 -1345 31935 -1310
rect 31970 -1345 31980 -1310
rect 32015 -1345 32025 -1310
rect 32060 -1345 32070 -1310
rect 32105 -1345 32115 -1310
rect 32150 -1345 32160 -1310
rect 32195 -1345 32205 -1310
rect 32240 -1345 32250 -1310
rect 32285 -1345 32295 -1310
rect 32330 -1345 32340 -1310
rect 32375 -1345 32385 -1310
rect 32420 -1345 32430 -1310
rect 32465 -1345 32475 -1310
rect 32510 -1345 32520 -1310
rect 32555 -1345 32565 -1310
rect 32600 -1345 32610 -1310
rect 32645 -1345 32655 -1310
rect 32690 -1345 32700 -1310
rect 32735 -1345 32745 -1310
rect 32780 -1345 32790 -1310
rect 32825 -1345 32835 -1310
rect 32870 -1345 32890 -1310
rect 31290 -1355 32890 -1345
rect 31290 -1390 31305 -1355
rect 31340 -1390 31350 -1355
rect 31385 -1390 31395 -1355
rect 31430 -1390 31440 -1355
rect 31475 -1390 31485 -1355
rect 31520 -1390 31530 -1355
rect 31565 -1390 31575 -1355
rect 31610 -1390 31620 -1355
rect 31655 -1390 31665 -1355
rect 31700 -1390 31710 -1355
rect 31745 -1390 31755 -1355
rect 31790 -1390 31800 -1355
rect 31835 -1390 31845 -1355
rect 31880 -1390 31890 -1355
rect 31925 -1390 31935 -1355
rect 31970 -1390 31980 -1355
rect 32015 -1390 32025 -1355
rect 32060 -1390 32070 -1355
rect 32105 -1390 32115 -1355
rect 32150 -1390 32160 -1355
rect 32195 -1390 32205 -1355
rect 32240 -1390 32250 -1355
rect 32285 -1390 32295 -1355
rect 32330 -1390 32340 -1355
rect 32375 -1390 32385 -1355
rect 32420 -1390 32430 -1355
rect 32465 -1390 32475 -1355
rect 32510 -1390 32520 -1355
rect 32555 -1390 32565 -1355
rect 32600 -1390 32610 -1355
rect 32645 -1390 32655 -1355
rect 32690 -1390 32700 -1355
rect 32735 -1390 32745 -1355
rect 32780 -1390 32790 -1355
rect 32825 -1390 32835 -1355
rect 32870 -1390 32890 -1355
rect 31290 -1400 32890 -1390
rect 31290 -1435 31305 -1400
rect 31340 -1435 31350 -1400
rect 31385 -1435 31395 -1400
rect 31430 -1435 31440 -1400
rect 31475 -1435 31485 -1400
rect 31520 -1435 31530 -1400
rect 31565 -1435 31575 -1400
rect 31610 -1435 31620 -1400
rect 31655 -1435 31665 -1400
rect 31700 -1435 31710 -1400
rect 31745 -1435 31755 -1400
rect 31790 -1435 31800 -1400
rect 31835 -1435 31845 -1400
rect 31880 -1435 31890 -1400
rect 31925 -1435 31935 -1400
rect 31970 -1435 31980 -1400
rect 32015 -1435 32025 -1400
rect 32060 -1435 32070 -1400
rect 32105 -1435 32115 -1400
rect 32150 -1435 32160 -1400
rect 32195 -1435 32205 -1400
rect 32240 -1435 32250 -1400
rect 32285 -1435 32295 -1400
rect 32330 -1435 32340 -1400
rect 32375 -1435 32385 -1400
rect 32420 -1435 32430 -1400
rect 32465 -1435 32475 -1400
rect 32510 -1435 32520 -1400
rect 32555 -1435 32565 -1400
rect 32600 -1435 32610 -1400
rect 32645 -1435 32655 -1400
rect 32690 -1435 32700 -1400
rect 32735 -1435 32745 -1400
rect 32780 -1435 32790 -1400
rect 32825 -1435 32835 -1400
rect 32870 -1435 32890 -1400
rect 31290 -1445 32890 -1435
rect 31290 -1480 31305 -1445
rect 31340 -1480 31350 -1445
rect 31385 -1480 31395 -1445
rect 31430 -1480 31440 -1445
rect 31475 -1480 31485 -1445
rect 31520 -1480 31530 -1445
rect 31565 -1480 31575 -1445
rect 31610 -1480 31620 -1445
rect 31655 -1480 31665 -1445
rect 31700 -1480 31710 -1445
rect 31745 -1480 31755 -1445
rect 31790 -1480 31800 -1445
rect 31835 -1480 31845 -1445
rect 31880 -1480 31890 -1445
rect 31925 -1480 31935 -1445
rect 31970 -1480 31980 -1445
rect 32015 -1480 32025 -1445
rect 32060 -1480 32070 -1445
rect 32105 -1480 32115 -1445
rect 32150 -1480 32160 -1445
rect 32195 -1480 32205 -1445
rect 32240 -1480 32250 -1445
rect 32285 -1480 32295 -1445
rect 32330 -1480 32340 -1445
rect 32375 -1480 32385 -1445
rect 32420 -1480 32430 -1445
rect 32465 -1480 32475 -1445
rect 32510 -1480 32520 -1445
rect 32555 -1480 32565 -1445
rect 32600 -1480 32610 -1445
rect 32645 -1480 32655 -1445
rect 32690 -1480 32700 -1445
rect 32735 -1480 32745 -1445
rect 32780 -1480 32790 -1445
rect 32825 -1480 32835 -1445
rect 32870 -1480 32890 -1445
rect 31290 -1490 32890 -1480
rect 31290 -1525 31305 -1490
rect 31340 -1525 31350 -1490
rect 31385 -1525 31395 -1490
rect 31430 -1525 31440 -1490
rect 31475 -1525 31485 -1490
rect 31520 -1525 31530 -1490
rect 31565 -1525 31575 -1490
rect 31610 -1525 31620 -1490
rect 31655 -1525 31665 -1490
rect 31700 -1525 31710 -1490
rect 31745 -1525 31755 -1490
rect 31790 -1525 31800 -1490
rect 31835 -1525 31845 -1490
rect 31880 -1525 31890 -1490
rect 31925 -1525 31935 -1490
rect 31970 -1525 31980 -1490
rect 32015 -1525 32025 -1490
rect 32060 -1525 32070 -1490
rect 32105 -1525 32115 -1490
rect 32150 -1525 32160 -1490
rect 32195 -1525 32205 -1490
rect 32240 -1525 32250 -1490
rect 32285 -1525 32295 -1490
rect 32330 -1525 32340 -1490
rect 32375 -1525 32385 -1490
rect 32420 -1525 32430 -1490
rect 32465 -1525 32475 -1490
rect 32510 -1525 32520 -1490
rect 32555 -1525 32565 -1490
rect 32600 -1525 32610 -1490
rect 32645 -1525 32655 -1490
rect 32690 -1525 32700 -1490
rect 32735 -1525 32745 -1490
rect 32780 -1525 32790 -1490
rect 32825 -1525 32835 -1490
rect 32870 -1525 32890 -1490
rect 31290 -1535 32890 -1525
rect 31290 -1570 31305 -1535
rect 31340 -1570 31350 -1535
rect 31385 -1570 31395 -1535
rect 31430 -1570 31440 -1535
rect 31475 -1570 31485 -1535
rect 31520 -1570 31530 -1535
rect 31565 -1570 31575 -1535
rect 31610 -1570 31620 -1535
rect 31655 -1570 31665 -1535
rect 31700 -1570 31710 -1535
rect 31745 -1570 31755 -1535
rect 31790 -1570 31800 -1535
rect 31835 -1570 31845 -1535
rect 31880 -1570 31890 -1535
rect 31925 -1570 31935 -1535
rect 31970 -1570 31980 -1535
rect 32015 -1570 32025 -1535
rect 32060 -1570 32070 -1535
rect 32105 -1570 32115 -1535
rect 32150 -1570 32160 -1535
rect 32195 -1570 32205 -1535
rect 32240 -1570 32250 -1535
rect 32285 -1570 32295 -1535
rect 32330 -1570 32340 -1535
rect 32375 -1570 32385 -1535
rect 32420 -1570 32430 -1535
rect 32465 -1570 32475 -1535
rect 32510 -1570 32520 -1535
rect 32555 -1570 32565 -1535
rect 32600 -1570 32610 -1535
rect 32645 -1570 32655 -1535
rect 32690 -1570 32700 -1535
rect 32735 -1570 32745 -1535
rect 32780 -1570 32790 -1535
rect 32825 -1570 32835 -1535
rect 32870 -1570 32890 -1535
rect 31290 -1580 32890 -1570
rect 31290 -1615 31305 -1580
rect 31340 -1615 31350 -1580
rect 31385 -1615 31395 -1580
rect 31430 -1615 31440 -1580
rect 31475 -1615 31485 -1580
rect 31520 -1615 31530 -1580
rect 31565 -1615 31575 -1580
rect 31610 -1615 31620 -1580
rect 31655 -1615 31665 -1580
rect 31700 -1615 31710 -1580
rect 31745 -1615 31755 -1580
rect 31790 -1615 31800 -1580
rect 31835 -1615 31845 -1580
rect 31880 -1615 31890 -1580
rect 31925 -1615 31935 -1580
rect 31970 -1615 31980 -1580
rect 32015 -1615 32025 -1580
rect 32060 -1615 32070 -1580
rect 32105 -1615 32115 -1580
rect 32150 -1615 32160 -1580
rect 32195 -1615 32205 -1580
rect 32240 -1615 32250 -1580
rect 32285 -1615 32295 -1580
rect 32330 -1615 32340 -1580
rect 32375 -1615 32385 -1580
rect 32420 -1615 32430 -1580
rect 32465 -1615 32475 -1580
rect 32510 -1615 32520 -1580
rect 32555 -1615 32565 -1580
rect 32600 -1615 32610 -1580
rect 32645 -1615 32655 -1580
rect 32690 -1615 32700 -1580
rect 32735 -1615 32745 -1580
rect 32780 -1615 32790 -1580
rect 32825 -1615 32835 -1580
rect 32870 -1615 32890 -1580
rect 31290 -1625 32890 -1615
rect 31290 -1660 31305 -1625
rect 31340 -1660 31350 -1625
rect 31385 -1660 31395 -1625
rect 31430 -1660 31440 -1625
rect 31475 -1660 31485 -1625
rect 31520 -1660 31530 -1625
rect 31565 -1660 31575 -1625
rect 31610 -1660 31620 -1625
rect 31655 -1660 31665 -1625
rect 31700 -1660 31710 -1625
rect 31745 -1660 31755 -1625
rect 31790 -1660 31800 -1625
rect 31835 -1660 31845 -1625
rect 31880 -1660 31890 -1625
rect 31925 -1660 31935 -1625
rect 31970 -1660 31980 -1625
rect 32015 -1660 32025 -1625
rect 32060 -1660 32070 -1625
rect 32105 -1660 32115 -1625
rect 32150 -1660 32160 -1625
rect 32195 -1660 32205 -1625
rect 32240 -1660 32250 -1625
rect 32285 -1660 32295 -1625
rect 32330 -1660 32340 -1625
rect 32375 -1660 32385 -1625
rect 32420 -1660 32430 -1625
rect 32465 -1660 32475 -1625
rect 32510 -1660 32520 -1625
rect 32555 -1660 32565 -1625
rect 32600 -1660 32610 -1625
rect 32645 -1660 32655 -1625
rect 32690 -1660 32700 -1625
rect 32735 -1660 32745 -1625
rect 32780 -1660 32790 -1625
rect 32825 -1660 32835 -1625
rect 32870 -1660 32890 -1625
rect 31290 -1670 32890 -1660
rect 31290 -1705 31305 -1670
rect 31340 -1705 31350 -1670
rect 31385 -1705 31395 -1670
rect 31430 -1705 31440 -1670
rect 31475 -1705 31485 -1670
rect 31520 -1705 31530 -1670
rect 31565 -1705 31575 -1670
rect 31610 -1705 31620 -1670
rect 31655 -1705 31665 -1670
rect 31700 -1705 31710 -1670
rect 31745 -1705 31755 -1670
rect 31790 -1705 31800 -1670
rect 31835 -1705 31845 -1670
rect 31880 -1705 31890 -1670
rect 31925 -1705 31935 -1670
rect 31970 -1705 31980 -1670
rect 32015 -1705 32025 -1670
rect 32060 -1705 32070 -1670
rect 32105 -1705 32115 -1670
rect 32150 -1705 32160 -1670
rect 32195 -1705 32205 -1670
rect 32240 -1705 32250 -1670
rect 32285 -1705 32295 -1670
rect 32330 -1705 32340 -1670
rect 32375 -1705 32385 -1670
rect 32420 -1705 32430 -1670
rect 32465 -1705 32475 -1670
rect 32510 -1705 32520 -1670
rect 32555 -1705 32565 -1670
rect 32600 -1705 32610 -1670
rect 32645 -1705 32655 -1670
rect 32690 -1705 32700 -1670
rect 32735 -1705 32745 -1670
rect 32780 -1705 32790 -1670
rect 32825 -1705 32835 -1670
rect 32870 -1705 32890 -1670
rect 31290 -1715 32890 -1705
rect 31290 -1750 31305 -1715
rect 31340 -1750 31350 -1715
rect 31385 -1750 31395 -1715
rect 31430 -1750 31440 -1715
rect 31475 -1750 31485 -1715
rect 31520 -1750 31530 -1715
rect 31565 -1750 31575 -1715
rect 31610 -1750 31620 -1715
rect 31655 -1750 31665 -1715
rect 31700 -1750 31710 -1715
rect 31745 -1750 31755 -1715
rect 31790 -1750 31800 -1715
rect 31835 -1750 31845 -1715
rect 31880 -1750 31890 -1715
rect 31925 -1750 31935 -1715
rect 31970 -1750 31980 -1715
rect 32015 -1750 32025 -1715
rect 32060 -1750 32070 -1715
rect 32105 -1750 32115 -1715
rect 32150 -1750 32160 -1715
rect 32195 -1750 32205 -1715
rect 32240 -1750 32250 -1715
rect 32285 -1750 32295 -1715
rect 32330 -1750 32340 -1715
rect 32375 -1750 32385 -1715
rect 32420 -1750 32430 -1715
rect 32465 -1750 32475 -1715
rect 32510 -1750 32520 -1715
rect 32555 -1750 32565 -1715
rect 32600 -1750 32610 -1715
rect 32645 -1750 32655 -1715
rect 32690 -1750 32700 -1715
rect 32735 -1750 32745 -1715
rect 32780 -1750 32790 -1715
rect 32825 -1750 32835 -1715
rect 32870 -1750 32890 -1715
rect 31290 -1760 32890 -1750
rect 31290 -1795 31305 -1760
rect 31340 -1795 31350 -1760
rect 31385 -1795 31395 -1760
rect 31430 -1795 31440 -1760
rect 31475 -1795 31485 -1760
rect 31520 -1795 31530 -1760
rect 31565 -1795 31575 -1760
rect 31610 -1795 31620 -1760
rect 31655 -1795 31665 -1760
rect 31700 -1795 31710 -1760
rect 31745 -1795 31755 -1760
rect 31790 -1795 31800 -1760
rect 31835 -1795 31845 -1760
rect 31880 -1795 31890 -1760
rect 31925 -1795 31935 -1760
rect 31970 -1795 31980 -1760
rect 32015 -1795 32025 -1760
rect 32060 -1795 32070 -1760
rect 32105 -1795 32115 -1760
rect 32150 -1795 32160 -1760
rect 32195 -1795 32205 -1760
rect 32240 -1795 32250 -1760
rect 32285 -1795 32295 -1760
rect 32330 -1795 32340 -1760
rect 32375 -1795 32385 -1760
rect 32420 -1795 32430 -1760
rect 32465 -1795 32475 -1760
rect 32510 -1795 32520 -1760
rect 32555 -1795 32565 -1760
rect 32600 -1795 32610 -1760
rect 32645 -1795 32655 -1760
rect 32690 -1795 32700 -1760
rect 32735 -1795 32745 -1760
rect 32780 -1795 32790 -1760
rect 32825 -1795 32835 -1760
rect 32870 -1795 32890 -1760
rect 31290 -1805 32890 -1795
rect 31290 -1840 31305 -1805
rect 31340 -1840 31350 -1805
rect 31385 -1840 31395 -1805
rect 31430 -1840 31440 -1805
rect 31475 -1840 31485 -1805
rect 31520 -1840 31530 -1805
rect 31565 -1840 31575 -1805
rect 31610 -1840 31620 -1805
rect 31655 -1840 31665 -1805
rect 31700 -1840 31710 -1805
rect 31745 -1840 31755 -1805
rect 31790 -1840 31800 -1805
rect 31835 -1840 31845 -1805
rect 31880 -1840 31890 -1805
rect 31925 -1840 31935 -1805
rect 31970 -1840 31980 -1805
rect 32015 -1840 32025 -1805
rect 32060 -1840 32070 -1805
rect 32105 -1840 32115 -1805
rect 32150 -1840 32160 -1805
rect 32195 -1840 32205 -1805
rect 32240 -1840 32250 -1805
rect 32285 -1840 32295 -1805
rect 32330 -1840 32340 -1805
rect 32375 -1840 32385 -1805
rect 32420 -1840 32430 -1805
rect 32465 -1840 32475 -1805
rect 32510 -1840 32520 -1805
rect 32555 -1840 32565 -1805
rect 32600 -1840 32610 -1805
rect 32645 -1840 32655 -1805
rect 32690 -1840 32700 -1805
rect 32735 -1840 32745 -1805
rect 32780 -1840 32790 -1805
rect 32825 -1840 32835 -1805
rect 32870 -1840 32890 -1805
rect 31290 -1850 32890 -1840
rect 31290 -1885 31305 -1850
rect 31340 -1885 31350 -1850
rect 31385 -1885 31395 -1850
rect 31430 -1885 31440 -1850
rect 31475 -1885 31485 -1850
rect 31520 -1885 31530 -1850
rect 31565 -1885 31575 -1850
rect 31610 -1885 31620 -1850
rect 31655 -1885 31665 -1850
rect 31700 -1885 31710 -1850
rect 31745 -1885 31755 -1850
rect 31790 -1885 31800 -1850
rect 31835 -1885 31845 -1850
rect 31880 -1885 31890 -1850
rect 31925 -1885 31935 -1850
rect 31970 -1885 31980 -1850
rect 32015 -1885 32025 -1850
rect 32060 -1885 32070 -1850
rect 32105 -1885 32115 -1850
rect 32150 -1885 32160 -1850
rect 32195 -1885 32205 -1850
rect 32240 -1885 32250 -1850
rect 32285 -1885 32295 -1850
rect 32330 -1885 32340 -1850
rect 32375 -1885 32385 -1850
rect 32420 -1885 32430 -1850
rect 32465 -1885 32475 -1850
rect 32510 -1885 32520 -1850
rect 32555 -1885 32565 -1850
rect 32600 -1885 32610 -1850
rect 32645 -1885 32655 -1850
rect 32690 -1885 32700 -1850
rect 32735 -1885 32745 -1850
rect 32780 -1885 32790 -1850
rect 32825 -1885 32835 -1850
rect 32870 -1885 32890 -1850
rect 31290 -1895 32890 -1885
rect 31290 -1930 31305 -1895
rect 31340 -1930 31350 -1895
rect 31385 -1930 31395 -1895
rect 31430 -1930 31440 -1895
rect 31475 -1930 31485 -1895
rect 31520 -1930 31530 -1895
rect 31565 -1930 31575 -1895
rect 31610 -1930 31620 -1895
rect 31655 -1930 31665 -1895
rect 31700 -1930 31710 -1895
rect 31745 -1930 31755 -1895
rect 31790 -1930 31800 -1895
rect 31835 -1930 31845 -1895
rect 31880 -1930 31890 -1895
rect 31925 -1930 31935 -1895
rect 31970 -1930 31980 -1895
rect 32015 -1930 32025 -1895
rect 32060 -1930 32070 -1895
rect 32105 -1930 32115 -1895
rect 32150 -1930 32160 -1895
rect 32195 -1930 32205 -1895
rect 32240 -1930 32250 -1895
rect 32285 -1930 32295 -1895
rect 32330 -1930 32340 -1895
rect 32375 -1930 32385 -1895
rect 32420 -1930 32430 -1895
rect 32465 -1930 32475 -1895
rect 32510 -1930 32520 -1895
rect 32555 -1930 32565 -1895
rect 32600 -1930 32610 -1895
rect 32645 -1930 32655 -1895
rect 32690 -1930 32700 -1895
rect 32735 -1930 32745 -1895
rect 32780 -1930 32790 -1895
rect 32825 -1930 32835 -1895
rect 32870 -1930 32890 -1895
rect 31290 -1940 32890 -1930
rect 31290 -1975 31305 -1940
rect 31340 -1975 31350 -1940
rect 31385 -1975 31395 -1940
rect 31430 -1975 31440 -1940
rect 31475 -1975 31485 -1940
rect 31520 -1975 31530 -1940
rect 31565 -1975 31575 -1940
rect 31610 -1975 31620 -1940
rect 31655 -1975 31665 -1940
rect 31700 -1975 31710 -1940
rect 31745 -1975 31755 -1940
rect 31790 -1975 31800 -1940
rect 31835 -1975 31845 -1940
rect 31880 -1975 31890 -1940
rect 31925 -1975 31935 -1940
rect 31970 -1975 31980 -1940
rect 32015 -1975 32025 -1940
rect 32060 -1975 32070 -1940
rect 32105 -1975 32115 -1940
rect 32150 -1975 32160 -1940
rect 32195 -1975 32205 -1940
rect 32240 -1975 32250 -1940
rect 32285 -1975 32295 -1940
rect 32330 -1975 32340 -1940
rect 32375 -1975 32385 -1940
rect 32420 -1975 32430 -1940
rect 32465 -1975 32475 -1940
rect 32510 -1975 32520 -1940
rect 32555 -1975 32565 -1940
rect 32600 -1975 32610 -1940
rect 32645 -1975 32655 -1940
rect 32690 -1975 32700 -1940
rect 32735 -1975 32745 -1940
rect 32780 -1975 32790 -1940
rect 32825 -1975 32835 -1940
rect 32870 -1975 32890 -1940
rect 31290 -1985 32890 -1975
rect 31290 -2020 31305 -1985
rect 31340 -2020 31350 -1985
rect 31385 -2020 31395 -1985
rect 31430 -2020 31440 -1985
rect 31475 -2020 31485 -1985
rect 31520 -2020 31530 -1985
rect 31565 -2020 31575 -1985
rect 31610 -2020 31620 -1985
rect 31655 -2020 31665 -1985
rect 31700 -2020 31710 -1985
rect 31745 -2020 31755 -1985
rect 31790 -2020 31800 -1985
rect 31835 -2020 31845 -1985
rect 31880 -2020 31890 -1985
rect 31925 -2020 31935 -1985
rect 31970 -2020 31980 -1985
rect 32015 -2020 32025 -1985
rect 32060 -2020 32070 -1985
rect 32105 -2020 32115 -1985
rect 32150 -2020 32160 -1985
rect 32195 -2020 32205 -1985
rect 32240 -2020 32250 -1985
rect 32285 -2020 32295 -1985
rect 32330 -2020 32340 -1985
rect 32375 -2020 32385 -1985
rect 32420 -2020 32430 -1985
rect 32465 -2020 32475 -1985
rect 32510 -2020 32520 -1985
rect 32555 -2020 32565 -1985
rect 32600 -2020 32610 -1985
rect 32645 -2020 32655 -1985
rect 32690 -2020 32700 -1985
rect 32735 -2020 32745 -1985
rect 32780 -2020 32790 -1985
rect 32825 -2020 32835 -1985
rect 32870 -2020 32890 -1985
rect 31290 -2030 32890 -2020
rect 31290 -2065 31305 -2030
rect 31340 -2065 31350 -2030
rect 31385 -2065 31395 -2030
rect 31430 -2065 31440 -2030
rect 31475 -2065 31485 -2030
rect 31520 -2065 31530 -2030
rect 31565 -2065 31575 -2030
rect 31610 -2065 31620 -2030
rect 31655 -2065 31665 -2030
rect 31700 -2065 31710 -2030
rect 31745 -2065 31755 -2030
rect 31790 -2065 31800 -2030
rect 31835 -2065 31845 -2030
rect 31880 -2065 31890 -2030
rect 31925 -2065 31935 -2030
rect 31970 -2065 31980 -2030
rect 32015 -2065 32025 -2030
rect 32060 -2065 32070 -2030
rect 32105 -2065 32115 -2030
rect 32150 -2065 32160 -2030
rect 32195 -2065 32205 -2030
rect 32240 -2065 32250 -2030
rect 32285 -2065 32295 -2030
rect 32330 -2065 32340 -2030
rect 32375 -2065 32385 -2030
rect 32420 -2065 32430 -2030
rect 32465 -2065 32475 -2030
rect 32510 -2065 32520 -2030
rect 32555 -2065 32565 -2030
rect 32600 -2065 32610 -2030
rect 32645 -2065 32655 -2030
rect 32690 -2065 32700 -2030
rect 32735 -2065 32745 -2030
rect 32780 -2065 32790 -2030
rect 32825 -2065 32835 -2030
rect 32870 -2065 32890 -2030
rect 31290 -2075 32890 -2065
rect 31290 -2110 31305 -2075
rect 31340 -2110 31350 -2075
rect 31385 -2110 31395 -2075
rect 31430 -2110 31440 -2075
rect 31475 -2110 31485 -2075
rect 31520 -2110 31530 -2075
rect 31565 -2110 31575 -2075
rect 31610 -2110 31620 -2075
rect 31655 -2110 31665 -2075
rect 31700 -2110 31710 -2075
rect 31745 -2110 31755 -2075
rect 31790 -2110 31800 -2075
rect 31835 -2110 31845 -2075
rect 31880 -2110 31890 -2075
rect 31925 -2110 31935 -2075
rect 31970 -2110 31980 -2075
rect 32015 -2110 32025 -2075
rect 32060 -2110 32070 -2075
rect 32105 -2110 32115 -2075
rect 32150 -2110 32160 -2075
rect 32195 -2110 32205 -2075
rect 32240 -2110 32250 -2075
rect 32285 -2110 32295 -2075
rect 32330 -2110 32340 -2075
rect 32375 -2110 32385 -2075
rect 32420 -2110 32430 -2075
rect 32465 -2110 32475 -2075
rect 32510 -2110 32520 -2075
rect 32555 -2110 32565 -2075
rect 32600 -2110 32610 -2075
rect 32645 -2110 32655 -2075
rect 32690 -2110 32700 -2075
rect 32735 -2110 32745 -2075
rect 32780 -2110 32790 -2075
rect 32825 -2110 32835 -2075
rect 32870 -2110 32890 -2075
rect 31290 -2120 32890 -2110
rect 31290 -2155 31305 -2120
rect 31340 -2155 31350 -2120
rect 31385 -2155 31395 -2120
rect 31430 -2155 31440 -2120
rect 31475 -2155 31485 -2120
rect 31520 -2155 31530 -2120
rect 31565 -2155 31575 -2120
rect 31610 -2155 31620 -2120
rect 31655 -2155 31665 -2120
rect 31700 -2155 31710 -2120
rect 31745 -2155 31755 -2120
rect 31790 -2155 31800 -2120
rect 31835 -2155 31845 -2120
rect 31880 -2155 31890 -2120
rect 31925 -2155 31935 -2120
rect 31970 -2155 31980 -2120
rect 32015 -2155 32025 -2120
rect 32060 -2155 32070 -2120
rect 32105 -2155 32115 -2120
rect 32150 -2155 32160 -2120
rect 32195 -2155 32205 -2120
rect 32240 -2155 32250 -2120
rect 32285 -2155 32295 -2120
rect 32330 -2155 32340 -2120
rect 32375 -2155 32385 -2120
rect 32420 -2155 32430 -2120
rect 32465 -2155 32475 -2120
rect 32510 -2155 32520 -2120
rect 32555 -2155 32565 -2120
rect 32600 -2155 32610 -2120
rect 32645 -2155 32655 -2120
rect 32690 -2155 32700 -2120
rect 32735 -2155 32745 -2120
rect 32780 -2155 32790 -2120
rect 32825 -2155 32835 -2120
rect 32870 -2155 32890 -2120
rect 31290 -2165 32890 -2155
rect 31290 -2200 31305 -2165
rect 31340 -2200 31350 -2165
rect 31385 -2200 31395 -2165
rect 31430 -2200 31440 -2165
rect 31475 -2200 31485 -2165
rect 31520 -2200 31530 -2165
rect 31565 -2200 31575 -2165
rect 31610 -2200 31620 -2165
rect 31655 -2200 31665 -2165
rect 31700 -2200 31710 -2165
rect 31745 -2200 31755 -2165
rect 31790 -2200 31800 -2165
rect 31835 -2200 31845 -2165
rect 31880 -2200 31890 -2165
rect 31925 -2200 31935 -2165
rect 31970 -2200 31980 -2165
rect 32015 -2200 32025 -2165
rect 32060 -2200 32070 -2165
rect 32105 -2200 32115 -2165
rect 32150 -2200 32160 -2165
rect 32195 -2200 32205 -2165
rect 32240 -2200 32250 -2165
rect 32285 -2200 32295 -2165
rect 32330 -2200 32340 -2165
rect 32375 -2200 32385 -2165
rect 32420 -2200 32430 -2165
rect 32465 -2200 32475 -2165
rect 32510 -2200 32520 -2165
rect 32555 -2200 32565 -2165
rect 32600 -2200 32610 -2165
rect 32645 -2200 32655 -2165
rect 32690 -2200 32700 -2165
rect 32735 -2200 32745 -2165
rect 32780 -2200 32790 -2165
rect 32825 -2200 32835 -2165
rect 32870 -2200 32890 -2165
rect 31290 -2210 32890 -2200
rect 31290 -2245 31305 -2210
rect 31340 -2245 31350 -2210
rect 31385 -2245 31395 -2210
rect 31430 -2245 31440 -2210
rect 31475 -2245 31485 -2210
rect 31520 -2245 31530 -2210
rect 31565 -2245 31575 -2210
rect 31610 -2245 31620 -2210
rect 31655 -2245 31665 -2210
rect 31700 -2245 31710 -2210
rect 31745 -2245 31755 -2210
rect 31790 -2245 31800 -2210
rect 31835 -2245 31845 -2210
rect 31880 -2245 31890 -2210
rect 31925 -2245 31935 -2210
rect 31970 -2245 31980 -2210
rect 32015 -2245 32025 -2210
rect 32060 -2245 32070 -2210
rect 32105 -2245 32115 -2210
rect 32150 -2245 32160 -2210
rect 32195 -2245 32205 -2210
rect 32240 -2245 32250 -2210
rect 32285 -2245 32295 -2210
rect 32330 -2245 32340 -2210
rect 32375 -2245 32385 -2210
rect 32420 -2245 32430 -2210
rect 32465 -2245 32475 -2210
rect 32510 -2245 32520 -2210
rect 32555 -2245 32565 -2210
rect 32600 -2245 32610 -2210
rect 32645 -2245 32655 -2210
rect 32690 -2245 32700 -2210
rect 32735 -2245 32745 -2210
rect 32780 -2245 32790 -2210
rect 32825 -2245 32835 -2210
rect 32870 -2245 32890 -2210
rect 31290 -2255 32890 -2245
rect 31290 -2290 31305 -2255
rect 31340 -2290 31350 -2255
rect 31385 -2290 31395 -2255
rect 31430 -2290 31440 -2255
rect 31475 -2290 31485 -2255
rect 31520 -2290 31530 -2255
rect 31565 -2290 31575 -2255
rect 31610 -2290 31620 -2255
rect 31655 -2290 31665 -2255
rect 31700 -2290 31710 -2255
rect 31745 -2290 31755 -2255
rect 31790 -2290 31800 -2255
rect 31835 -2290 31845 -2255
rect 31880 -2290 31890 -2255
rect 31925 -2290 31935 -2255
rect 31970 -2290 31980 -2255
rect 32015 -2290 32025 -2255
rect 32060 -2290 32070 -2255
rect 32105 -2290 32115 -2255
rect 32150 -2290 32160 -2255
rect 32195 -2290 32205 -2255
rect 32240 -2290 32250 -2255
rect 32285 -2290 32295 -2255
rect 32330 -2290 32340 -2255
rect 32375 -2290 32385 -2255
rect 32420 -2290 32430 -2255
rect 32465 -2290 32475 -2255
rect 32510 -2290 32520 -2255
rect 32555 -2290 32565 -2255
rect 32600 -2290 32610 -2255
rect 32645 -2290 32655 -2255
rect 32690 -2290 32700 -2255
rect 32735 -2290 32745 -2255
rect 32780 -2290 32790 -2255
rect 32825 -2290 32835 -2255
rect 32870 -2290 32890 -2255
rect 31290 -2300 32890 -2290
rect 31290 -2335 31305 -2300
rect 31340 -2335 31350 -2300
rect 31385 -2335 31395 -2300
rect 31430 -2335 31440 -2300
rect 31475 -2335 31485 -2300
rect 31520 -2335 31530 -2300
rect 31565 -2335 31575 -2300
rect 31610 -2335 31620 -2300
rect 31655 -2335 31665 -2300
rect 31700 -2335 31710 -2300
rect 31745 -2335 31755 -2300
rect 31790 -2335 31800 -2300
rect 31835 -2335 31845 -2300
rect 31880 -2335 31890 -2300
rect 31925 -2335 31935 -2300
rect 31970 -2335 31980 -2300
rect 32015 -2335 32025 -2300
rect 32060 -2335 32070 -2300
rect 32105 -2335 32115 -2300
rect 32150 -2335 32160 -2300
rect 32195 -2335 32205 -2300
rect 32240 -2335 32250 -2300
rect 32285 -2335 32295 -2300
rect 32330 -2335 32340 -2300
rect 32375 -2335 32385 -2300
rect 32420 -2335 32430 -2300
rect 32465 -2335 32475 -2300
rect 32510 -2335 32520 -2300
rect 32555 -2335 32565 -2300
rect 32600 -2335 32610 -2300
rect 32645 -2335 32655 -2300
rect 32690 -2335 32700 -2300
rect 32735 -2335 32745 -2300
rect 32780 -2335 32790 -2300
rect 32825 -2335 32835 -2300
rect 32870 -2335 32890 -2300
rect 31290 -2345 32890 -2335
rect 31290 -2380 31305 -2345
rect 31340 -2380 31350 -2345
rect 31385 -2380 31395 -2345
rect 31430 -2380 31440 -2345
rect 31475 -2380 31485 -2345
rect 31520 -2380 31530 -2345
rect 31565 -2380 31575 -2345
rect 31610 -2380 31620 -2345
rect 31655 -2380 31665 -2345
rect 31700 -2380 31710 -2345
rect 31745 -2380 31755 -2345
rect 31790 -2380 31800 -2345
rect 31835 -2380 31845 -2345
rect 31880 -2380 31890 -2345
rect 31925 -2380 31935 -2345
rect 31970 -2380 31980 -2345
rect 32015 -2380 32025 -2345
rect 32060 -2380 32070 -2345
rect 32105 -2380 32115 -2345
rect 32150 -2380 32160 -2345
rect 32195 -2380 32205 -2345
rect 32240 -2380 32250 -2345
rect 32285 -2380 32295 -2345
rect 32330 -2380 32340 -2345
rect 32375 -2380 32385 -2345
rect 32420 -2380 32430 -2345
rect 32465 -2380 32475 -2345
rect 32510 -2380 32520 -2345
rect 32555 -2380 32565 -2345
rect 32600 -2380 32610 -2345
rect 32645 -2380 32655 -2345
rect 32690 -2380 32700 -2345
rect 32735 -2380 32745 -2345
rect 32780 -2380 32790 -2345
rect 32825 -2380 32835 -2345
rect 32870 -2380 32890 -2345
rect 31290 -2390 32890 -2380
rect 31290 -2425 31305 -2390
rect 31340 -2425 31350 -2390
rect 31385 -2425 31395 -2390
rect 31430 -2425 31440 -2390
rect 31475 -2425 31485 -2390
rect 31520 -2425 31530 -2390
rect 31565 -2425 31575 -2390
rect 31610 -2425 31620 -2390
rect 31655 -2425 31665 -2390
rect 31700 -2425 31710 -2390
rect 31745 -2425 31755 -2390
rect 31790 -2425 31800 -2390
rect 31835 -2425 31845 -2390
rect 31880 -2425 31890 -2390
rect 31925 -2425 31935 -2390
rect 31970 -2425 31980 -2390
rect 32015 -2425 32025 -2390
rect 32060 -2425 32070 -2390
rect 32105 -2425 32115 -2390
rect 32150 -2425 32160 -2390
rect 32195 -2425 32205 -2390
rect 32240 -2425 32250 -2390
rect 32285 -2425 32295 -2390
rect 32330 -2425 32340 -2390
rect 32375 -2425 32385 -2390
rect 32420 -2425 32430 -2390
rect 32465 -2425 32475 -2390
rect 32510 -2425 32520 -2390
rect 32555 -2425 32565 -2390
rect 32600 -2425 32610 -2390
rect 32645 -2425 32655 -2390
rect 32690 -2425 32700 -2390
rect 32735 -2425 32745 -2390
rect 32780 -2425 32790 -2390
rect 32825 -2425 32835 -2390
rect 32870 -2425 32890 -2390
rect 31290 -2435 32890 -2425
rect 31290 -2470 31305 -2435
rect 31340 -2470 31350 -2435
rect 31385 -2470 31395 -2435
rect 31430 -2470 31440 -2435
rect 31475 -2470 31485 -2435
rect 31520 -2470 31530 -2435
rect 31565 -2470 31575 -2435
rect 31610 -2470 31620 -2435
rect 31655 -2470 31665 -2435
rect 31700 -2470 31710 -2435
rect 31745 -2470 31755 -2435
rect 31790 -2470 31800 -2435
rect 31835 -2470 31845 -2435
rect 31880 -2470 31890 -2435
rect 31925 -2470 31935 -2435
rect 31970 -2470 31980 -2435
rect 32015 -2470 32025 -2435
rect 32060 -2470 32070 -2435
rect 32105 -2470 32115 -2435
rect 32150 -2470 32160 -2435
rect 32195 -2470 32205 -2435
rect 32240 -2470 32250 -2435
rect 32285 -2470 32295 -2435
rect 32330 -2470 32340 -2435
rect 32375 -2470 32385 -2435
rect 32420 -2470 32430 -2435
rect 32465 -2470 32475 -2435
rect 32510 -2470 32520 -2435
rect 32555 -2470 32565 -2435
rect 32600 -2470 32610 -2435
rect 32645 -2470 32655 -2435
rect 32690 -2470 32700 -2435
rect 32735 -2470 32745 -2435
rect 32780 -2470 32790 -2435
rect 32825 -2470 32835 -2435
rect 32870 -2470 32890 -2435
rect 31290 -2480 32890 -2470
rect 31290 -2515 31305 -2480
rect 31340 -2515 31350 -2480
rect 31385 -2515 31395 -2480
rect 31430 -2515 31440 -2480
rect 31475 -2515 31485 -2480
rect 31520 -2515 31530 -2480
rect 31565 -2515 31575 -2480
rect 31610 -2515 31620 -2480
rect 31655 -2515 31665 -2480
rect 31700 -2515 31710 -2480
rect 31745 -2515 31755 -2480
rect 31790 -2515 31800 -2480
rect 31835 -2515 31845 -2480
rect 31880 -2515 31890 -2480
rect 31925 -2515 31935 -2480
rect 31970 -2515 31980 -2480
rect 32015 -2515 32025 -2480
rect 32060 -2515 32070 -2480
rect 32105 -2515 32115 -2480
rect 32150 -2515 32160 -2480
rect 32195 -2515 32205 -2480
rect 32240 -2515 32250 -2480
rect 32285 -2515 32295 -2480
rect 32330 -2515 32340 -2480
rect 32375 -2515 32385 -2480
rect 32420 -2515 32430 -2480
rect 32465 -2515 32475 -2480
rect 32510 -2515 32520 -2480
rect 32555 -2515 32565 -2480
rect 32600 -2515 32610 -2480
rect 32645 -2515 32655 -2480
rect 32690 -2515 32700 -2480
rect 32735 -2515 32745 -2480
rect 32780 -2515 32790 -2480
rect 32825 -2515 32835 -2480
rect 32870 -2515 32890 -2480
rect 31290 -2525 32890 -2515
rect 31290 -2560 31305 -2525
rect 31340 -2560 31350 -2525
rect 31385 -2560 31395 -2525
rect 31430 -2560 31440 -2525
rect 31475 -2560 31485 -2525
rect 31520 -2560 31530 -2525
rect 31565 -2560 31575 -2525
rect 31610 -2560 31620 -2525
rect 31655 -2560 31665 -2525
rect 31700 -2560 31710 -2525
rect 31745 -2560 31755 -2525
rect 31790 -2560 31800 -2525
rect 31835 -2560 31845 -2525
rect 31880 -2560 31890 -2525
rect 31925 -2560 31935 -2525
rect 31970 -2560 31980 -2525
rect 32015 -2560 32025 -2525
rect 32060 -2560 32070 -2525
rect 32105 -2560 32115 -2525
rect 32150 -2560 32160 -2525
rect 32195 -2560 32205 -2525
rect 32240 -2560 32250 -2525
rect 32285 -2560 32295 -2525
rect 32330 -2560 32340 -2525
rect 32375 -2560 32385 -2525
rect 32420 -2560 32430 -2525
rect 32465 -2560 32475 -2525
rect 32510 -2560 32520 -2525
rect 32555 -2560 32565 -2525
rect 32600 -2560 32610 -2525
rect 32645 -2560 32655 -2525
rect 32690 -2560 32700 -2525
rect 32735 -2560 32745 -2525
rect 32780 -2560 32790 -2525
rect 32825 -2560 32835 -2525
rect 32870 -2560 32890 -2525
rect 31290 -2570 32890 -2560
rect 31290 -2605 31305 -2570
rect 31340 -2605 31350 -2570
rect 31385 -2605 31395 -2570
rect 31430 -2605 31440 -2570
rect 31475 -2605 31485 -2570
rect 31520 -2605 31530 -2570
rect 31565 -2605 31575 -2570
rect 31610 -2605 31620 -2570
rect 31655 -2605 31665 -2570
rect 31700 -2605 31710 -2570
rect 31745 -2605 31755 -2570
rect 31790 -2605 31800 -2570
rect 31835 -2605 31845 -2570
rect 31880 -2605 31890 -2570
rect 31925 -2605 31935 -2570
rect 31970 -2605 31980 -2570
rect 32015 -2605 32025 -2570
rect 32060 -2605 32070 -2570
rect 32105 -2605 32115 -2570
rect 32150 -2605 32160 -2570
rect 32195 -2605 32205 -2570
rect 32240 -2605 32250 -2570
rect 32285 -2605 32295 -2570
rect 32330 -2605 32340 -2570
rect 32375 -2605 32385 -2570
rect 32420 -2605 32430 -2570
rect 32465 -2605 32475 -2570
rect 32510 -2605 32520 -2570
rect 32555 -2605 32565 -2570
rect 32600 -2605 32610 -2570
rect 32645 -2605 32655 -2570
rect 32690 -2605 32700 -2570
rect 32735 -2605 32745 -2570
rect 32780 -2605 32790 -2570
rect 32825 -2605 32835 -2570
rect 32870 -2605 32890 -2570
rect 31290 -2615 32890 -2605
rect 31290 -2650 31305 -2615
rect 31340 -2650 31350 -2615
rect 31385 -2650 31395 -2615
rect 31430 -2650 31440 -2615
rect 31475 -2650 31485 -2615
rect 31520 -2650 31530 -2615
rect 31565 -2650 31575 -2615
rect 31610 -2650 31620 -2615
rect 31655 -2650 31665 -2615
rect 31700 -2650 31710 -2615
rect 31745 -2650 31755 -2615
rect 31790 -2650 31800 -2615
rect 31835 -2650 31845 -2615
rect 31880 -2650 31890 -2615
rect 31925 -2650 31935 -2615
rect 31970 -2650 31980 -2615
rect 32015 -2650 32025 -2615
rect 32060 -2650 32070 -2615
rect 32105 -2650 32115 -2615
rect 32150 -2650 32160 -2615
rect 32195 -2650 32205 -2615
rect 32240 -2650 32250 -2615
rect 32285 -2650 32295 -2615
rect 32330 -2650 32340 -2615
rect 32375 -2650 32385 -2615
rect 32420 -2650 32430 -2615
rect 32465 -2650 32475 -2615
rect 32510 -2650 32520 -2615
rect 32555 -2650 32565 -2615
rect 32600 -2650 32610 -2615
rect 32645 -2650 32655 -2615
rect 32690 -2650 32700 -2615
rect 32735 -2650 32745 -2615
rect 32780 -2650 32790 -2615
rect 32825 -2650 32835 -2615
rect 32870 -2650 32890 -2615
rect 31290 -2660 32890 -2650
rect 31290 -2695 31305 -2660
rect 31340 -2695 31350 -2660
rect 31385 -2695 31395 -2660
rect 31430 -2695 31440 -2660
rect 31475 -2695 31485 -2660
rect 31520 -2695 31530 -2660
rect 31565 -2695 31575 -2660
rect 31610 -2695 31620 -2660
rect 31655 -2695 31665 -2660
rect 31700 -2695 31710 -2660
rect 31745 -2695 31755 -2660
rect 31790 -2695 31800 -2660
rect 31835 -2695 31845 -2660
rect 31880 -2695 31890 -2660
rect 31925 -2695 31935 -2660
rect 31970 -2695 31980 -2660
rect 32015 -2695 32025 -2660
rect 32060 -2695 32070 -2660
rect 32105 -2695 32115 -2660
rect 32150 -2695 32160 -2660
rect 32195 -2695 32205 -2660
rect 32240 -2695 32250 -2660
rect 32285 -2695 32295 -2660
rect 32330 -2695 32340 -2660
rect 32375 -2695 32385 -2660
rect 32420 -2695 32430 -2660
rect 32465 -2695 32475 -2660
rect 32510 -2695 32520 -2660
rect 32555 -2695 32565 -2660
rect 32600 -2695 32610 -2660
rect 32645 -2695 32655 -2660
rect 32690 -2695 32700 -2660
rect 32735 -2695 32745 -2660
rect 32780 -2695 32790 -2660
rect 32825 -2695 32835 -2660
rect 32870 -2695 32890 -2660
rect 31290 -2705 32890 -2695
rect 31290 -2740 31305 -2705
rect 31340 -2740 31350 -2705
rect 31385 -2740 31395 -2705
rect 31430 -2740 31440 -2705
rect 31475 -2740 31485 -2705
rect 31520 -2740 31530 -2705
rect 31565 -2740 31575 -2705
rect 31610 -2740 31620 -2705
rect 31655 -2740 31665 -2705
rect 31700 -2740 31710 -2705
rect 31745 -2740 31755 -2705
rect 31790 -2740 31800 -2705
rect 31835 -2740 31845 -2705
rect 31880 -2740 31890 -2705
rect 31925 -2740 31935 -2705
rect 31970 -2740 31980 -2705
rect 32015 -2740 32025 -2705
rect 32060 -2740 32070 -2705
rect 32105 -2740 32115 -2705
rect 32150 -2740 32160 -2705
rect 32195 -2740 32205 -2705
rect 32240 -2740 32250 -2705
rect 32285 -2740 32295 -2705
rect 32330 -2740 32340 -2705
rect 32375 -2740 32385 -2705
rect 32420 -2740 32430 -2705
rect 32465 -2740 32475 -2705
rect 32510 -2740 32520 -2705
rect 32555 -2740 32565 -2705
rect 32600 -2740 32610 -2705
rect 32645 -2740 32655 -2705
rect 32690 -2740 32700 -2705
rect 32735 -2740 32745 -2705
rect 32780 -2740 32790 -2705
rect 32825 -2740 32835 -2705
rect 32870 -2740 32890 -2705
rect 31290 -2750 32890 -2740
rect 31290 -2785 31305 -2750
rect 31340 -2785 31350 -2750
rect 31385 -2785 31395 -2750
rect 31430 -2785 31440 -2750
rect 31475 -2785 31485 -2750
rect 31520 -2785 31530 -2750
rect 31565 -2785 31575 -2750
rect 31610 -2785 31620 -2750
rect 31655 -2785 31665 -2750
rect 31700 -2785 31710 -2750
rect 31745 -2785 31755 -2750
rect 31790 -2785 31800 -2750
rect 31835 -2785 31845 -2750
rect 31880 -2785 31890 -2750
rect 31925 -2785 31935 -2750
rect 31970 -2785 31980 -2750
rect 32015 -2785 32025 -2750
rect 32060 -2785 32070 -2750
rect 32105 -2785 32115 -2750
rect 32150 -2785 32160 -2750
rect 32195 -2785 32205 -2750
rect 32240 -2785 32250 -2750
rect 32285 -2785 32295 -2750
rect 32330 -2785 32340 -2750
rect 32375 -2785 32385 -2750
rect 32420 -2785 32430 -2750
rect 32465 -2785 32475 -2750
rect 32510 -2785 32520 -2750
rect 32555 -2785 32565 -2750
rect 32600 -2785 32610 -2750
rect 32645 -2785 32655 -2750
rect 32690 -2785 32700 -2750
rect 32735 -2785 32745 -2750
rect 32780 -2785 32790 -2750
rect 32825 -2785 32835 -2750
rect 32870 -2785 32890 -2750
rect 31290 -2795 32890 -2785
rect 31290 -2830 31305 -2795
rect 31340 -2830 31350 -2795
rect 31385 -2830 31395 -2795
rect 31430 -2830 31440 -2795
rect 31475 -2830 31485 -2795
rect 31520 -2830 31530 -2795
rect 31565 -2830 31575 -2795
rect 31610 -2830 31620 -2795
rect 31655 -2830 31665 -2795
rect 31700 -2830 31710 -2795
rect 31745 -2830 31755 -2795
rect 31790 -2830 31800 -2795
rect 31835 -2830 31845 -2795
rect 31880 -2830 31890 -2795
rect 31925 -2830 31935 -2795
rect 31970 -2830 31980 -2795
rect 32015 -2830 32025 -2795
rect 32060 -2830 32070 -2795
rect 32105 -2830 32115 -2795
rect 32150 -2830 32160 -2795
rect 32195 -2830 32205 -2795
rect 32240 -2830 32250 -2795
rect 32285 -2830 32295 -2795
rect 32330 -2830 32340 -2795
rect 32375 -2830 32385 -2795
rect 32420 -2830 32430 -2795
rect 32465 -2830 32475 -2795
rect 32510 -2830 32520 -2795
rect 32555 -2830 32565 -2795
rect 32600 -2830 32610 -2795
rect 32645 -2830 32655 -2795
rect 32690 -2830 32700 -2795
rect 32735 -2830 32745 -2795
rect 32780 -2830 32790 -2795
rect 32825 -2830 32835 -2795
rect 32870 -2830 32890 -2795
rect 31290 -2840 32890 -2830
rect 31290 -2875 31305 -2840
rect 31340 -2875 31350 -2840
rect 31385 -2875 31395 -2840
rect 31430 -2875 31440 -2840
rect 31475 -2875 31485 -2840
rect 31520 -2875 31530 -2840
rect 31565 -2875 31575 -2840
rect 31610 -2875 31620 -2840
rect 31655 -2875 31665 -2840
rect 31700 -2875 31710 -2840
rect 31745 -2875 31755 -2840
rect 31790 -2875 31800 -2840
rect 31835 -2875 31845 -2840
rect 31880 -2875 31890 -2840
rect 31925 -2875 31935 -2840
rect 31970 -2875 31980 -2840
rect 32015 -2875 32025 -2840
rect 32060 -2875 32070 -2840
rect 32105 -2875 32115 -2840
rect 32150 -2875 32160 -2840
rect 32195 -2875 32205 -2840
rect 32240 -2875 32250 -2840
rect 32285 -2875 32295 -2840
rect 32330 -2875 32340 -2840
rect 32375 -2875 32385 -2840
rect 32420 -2875 32430 -2840
rect 32465 -2875 32475 -2840
rect 32510 -2875 32520 -2840
rect 32555 -2875 32565 -2840
rect 32600 -2875 32610 -2840
rect 32645 -2875 32655 -2840
rect 32690 -2875 32700 -2840
rect 32735 -2875 32745 -2840
rect 32780 -2875 32790 -2840
rect 32825 -2875 32835 -2840
rect 32870 -2875 32890 -2840
rect 31290 -2890 32890 -2875
<< via3 >>
rect 2110 19310 2150 19315
rect 2110 19280 2115 19310
rect 2115 19280 2145 19310
rect 2145 19280 2150 19310
rect 2110 19275 2150 19280
rect 2110 19245 2150 19250
rect 2110 19215 2115 19245
rect 2115 19215 2145 19245
rect 2145 19215 2150 19245
rect 2110 19210 2150 19215
rect 2110 19175 2150 19180
rect 2110 19145 2115 19175
rect 2115 19145 2145 19175
rect 2145 19145 2150 19175
rect 2110 19140 2150 19145
rect 2110 19105 2150 19110
rect 2110 19075 2115 19105
rect 2115 19075 2145 19105
rect 2145 19075 2150 19105
rect 2110 19070 2150 19075
rect 2110 19035 2150 19040
rect 2110 19005 2115 19035
rect 2115 19005 2145 19035
rect 2145 19005 2150 19035
rect 2110 19000 2150 19005
rect 2110 18970 2150 18975
rect 2110 18940 2115 18970
rect 2115 18940 2145 18970
rect 2145 18940 2150 18970
rect 2110 18935 2150 18940
rect 2110 18910 2150 18915
rect 2110 18880 2115 18910
rect 2115 18880 2145 18910
rect 2145 18880 2150 18910
rect 2110 18875 2150 18880
rect 2110 18845 2150 18850
rect 2110 18815 2115 18845
rect 2115 18815 2145 18845
rect 2145 18815 2150 18845
rect 2110 18810 2150 18815
rect 2110 18775 2150 18780
rect 2110 18745 2115 18775
rect 2115 18745 2145 18775
rect 2145 18745 2150 18775
rect 2110 18740 2150 18745
rect 2110 18705 2150 18710
rect 2110 18675 2115 18705
rect 2115 18675 2145 18705
rect 2145 18675 2150 18705
rect 2110 18670 2150 18675
rect 2110 18635 2150 18640
rect 2110 18605 2115 18635
rect 2115 18605 2145 18635
rect 2145 18605 2150 18635
rect 2110 18600 2150 18605
rect 2110 18570 2150 18575
rect 2110 18540 2115 18570
rect 2115 18540 2145 18570
rect 2145 18540 2150 18570
rect 2110 18535 2150 18540
rect 2110 18510 2150 18515
rect 2110 18480 2115 18510
rect 2115 18480 2145 18510
rect 2145 18480 2150 18510
rect 2110 18475 2150 18480
rect 2110 18445 2150 18450
rect 2110 18415 2115 18445
rect 2115 18415 2145 18445
rect 2145 18415 2150 18445
rect 2110 18410 2150 18415
rect 2110 18375 2150 18380
rect 2110 18345 2115 18375
rect 2115 18345 2145 18375
rect 2145 18345 2150 18375
rect 2110 18340 2150 18345
rect 2110 18305 2150 18310
rect 2110 18275 2115 18305
rect 2115 18275 2145 18305
rect 2145 18275 2150 18305
rect 2110 18270 2150 18275
rect 2110 18235 2150 18240
rect 2110 18205 2115 18235
rect 2115 18205 2145 18235
rect 2145 18205 2150 18235
rect 2110 18200 2150 18205
rect 2110 18170 2150 18175
rect 2110 18140 2115 18170
rect 2115 18140 2145 18170
rect 2145 18140 2150 18170
rect 2110 18135 2150 18140
rect 2110 18110 2150 18115
rect 2110 18080 2115 18110
rect 2115 18080 2145 18110
rect 2145 18080 2150 18110
rect 2110 18075 2150 18080
rect 2110 18045 2150 18050
rect 2110 18015 2115 18045
rect 2115 18015 2145 18045
rect 2145 18015 2150 18045
rect 2110 18010 2150 18015
rect 2110 17975 2150 17980
rect 2110 17945 2115 17975
rect 2115 17945 2145 17975
rect 2145 17945 2150 17975
rect 2110 17940 2150 17945
rect 2110 17905 2150 17910
rect 2110 17875 2115 17905
rect 2115 17875 2145 17905
rect 2145 17875 2150 17905
rect 2110 17870 2150 17875
rect 2110 17835 2150 17840
rect 2110 17805 2115 17835
rect 2115 17805 2145 17835
rect 2145 17805 2150 17835
rect 2110 17800 2150 17805
rect 2110 17770 2150 17775
rect 2110 17740 2115 17770
rect 2115 17740 2145 17770
rect 2145 17740 2150 17770
rect 2110 17735 2150 17740
rect 6700 19310 6740 19315
rect 6700 19280 6705 19310
rect 6705 19280 6735 19310
rect 6735 19280 6740 19310
rect 6700 19275 6740 19280
rect 6700 19245 6740 19250
rect 6700 19215 6705 19245
rect 6705 19215 6735 19245
rect 6735 19215 6740 19245
rect 6700 19210 6740 19215
rect 6700 19175 6740 19180
rect 6700 19145 6705 19175
rect 6705 19145 6735 19175
rect 6735 19145 6740 19175
rect 6700 19140 6740 19145
rect 6700 19105 6740 19110
rect 6700 19075 6705 19105
rect 6705 19075 6735 19105
rect 6735 19075 6740 19105
rect 6700 19070 6740 19075
rect 6700 19035 6740 19040
rect 6700 19005 6705 19035
rect 6705 19005 6735 19035
rect 6735 19005 6740 19035
rect 6700 19000 6740 19005
rect 6700 18970 6740 18975
rect 6700 18940 6705 18970
rect 6705 18940 6735 18970
rect 6735 18940 6740 18970
rect 6700 18935 6740 18940
rect 6700 18910 6740 18915
rect 6700 18880 6705 18910
rect 6705 18880 6735 18910
rect 6735 18880 6740 18910
rect 6700 18875 6740 18880
rect 6700 18845 6740 18850
rect 6700 18815 6705 18845
rect 6705 18815 6735 18845
rect 6735 18815 6740 18845
rect 6700 18810 6740 18815
rect 6700 18775 6740 18780
rect 6700 18745 6705 18775
rect 6705 18745 6735 18775
rect 6735 18745 6740 18775
rect 6700 18740 6740 18745
rect 6700 18705 6740 18710
rect 6700 18675 6705 18705
rect 6705 18675 6735 18705
rect 6735 18675 6740 18705
rect 6700 18670 6740 18675
rect 6700 18635 6740 18640
rect 6700 18605 6705 18635
rect 6705 18605 6735 18635
rect 6735 18605 6740 18635
rect 6700 18600 6740 18605
rect 6700 18570 6740 18575
rect 6700 18540 6705 18570
rect 6705 18540 6735 18570
rect 6735 18540 6740 18570
rect 6700 18535 6740 18540
rect 6700 18510 6740 18515
rect 6700 18480 6705 18510
rect 6705 18480 6735 18510
rect 6735 18480 6740 18510
rect 6700 18475 6740 18480
rect 6700 18445 6740 18450
rect 6700 18415 6705 18445
rect 6705 18415 6735 18445
rect 6735 18415 6740 18445
rect 6700 18410 6740 18415
rect 6700 18375 6740 18380
rect 6700 18345 6705 18375
rect 6705 18345 6735 18375
rect 6735 18345 6740 18375
rect 6700 18340 6740 18345
rect 6700 18305 6740 18310
rect 6700 18275 6705 18305
rect 6705 18275 6735 18305
rect 6735 18275 6740 18305
rect 6700 18270 6740 18275
rect 6700 18235 6740 18240
rect 6700 18205 6705 18235
rect 6705 18205 6735 18235
rect 6735 18205 6740 18235
rect 6700 18200 6740 18205
rect 6700 18170 6740 18175
rect 6700 18140 6705 18170
rect 6705 18140 6735 18170
rect 6735 18140 6740 18170
rect 6700 18135 6740 18140
rect 6700 18110 6740 18115
rect 6700 18080 6705 18110
rect 6705 18080 6735 18110
rect 6735 18080 6740 18110
rect 6700 18075 6740 18080
rect 6700 18045 6740 18050
rect 6700 18015 6705 18045
rect 6705 18015 6735 18045
rect 6735 18015 6740 18045
rect 6700 18010 6740 18015
rect 6700 17975 6740 17980
rect 6700 17945 6705 17975
rect 6705 17945 6735 17975
rect 6735 17945 6740 17975
rect 6700 17940 6740 17945
rect 6700 17905 6740 17910
rect 6700 17875 6705 17905
rect 6705 17875 6735 17905
rect 6735 17875 6740 17905
rect 6700 17870 6740 17875
rect 6700 17835 6740 17840
rect 6700 17805 6705 17835
rect 6705 17805 6735 17835
rect 6735 17805 6740 17835
rect 6700 17800 6740 17805
rect 6700 17770 6740 17775
rect 6700 17740 6705 17770
rect 6705 17740 6735 17770
rect 6735 17740 6740 17770
rect 6700 17735 6740 17740
rect 31305 19270 31340 19305
rect 31350 19270 31385 19305
rect 31395 19270 31430 19305
rect 31440 19270 31475 19305
rect 31485 19270 31520 19305
rect 31530 19270 31565 19305
rect 31575 19270 31610 19305
rect 31620 19270 31655 19305
rect 31665 19270 31700 19305
rect 31710 19270 31745 19305
rect 31755 19270 31790 19305
rect 31800 19270 31835 19305
rect 31845 19270 31880 19305
rect 31890 19270 31925 19305
rect 31935 19270 31970 19305
rect 31980 19270 32015 19305
rect 32025 19270 32060 19305
rect 32070 19270 32105 19305
rect 32115 19270 32150 19305
rect 32160 19270 32195 19305
rect 32205 19270 32240 19305
rect 32250 19270 32285 19305
rect 32295 19270 32330 19305
rect 32340 19270 32375 19305
rect 32385 19270 32420 19305
rect 32430 19270 32465 19305
rect 32475 19270 32510 19305
rect 32520 19270 32555 19305
rect 32565 19270 32600 19305
rect 32610 19270 32645 19305
rect 32655 19270 32690 19305
rect 32700 19270 32735 19305
rect 32745 19270 32780 19305
rect 32790 19270 32825 19305
rect 32835 19270 32870 19305
rect 31305 19225 31340 19260
rect 31350 19225 31385 19260
rect 31395 19225 31430 19260
rect 31440 19225 31475 19260
rect 31485 19225 31520 19260
rect 31530 19225 31565 19260
rect 31575 19225 31610 19260
rect 31620 19225 31655 19260
rect 31665 19225 31700 19260
rect 31710 19225 31745 19260
rect 31755 19225 31790 19260
rect 31800 19225 31835 19260
rect 31845 19225 31880 19260
rect 31890 19225 31925 19260
rect 31935 19225 31970 19260
rect 31980 19225 32015 19260
rect 32025 19225 32060 19260
rect 32070 19225 32105 19260
rect 32115 19225 32150 19260
rect 32160 19225 32195 19260
rect 32205 19225 32240 19260
rect 32250 19225 32285 19260
rect 32295 19225 32330 19260
rect 32340 19225 32375 19260
rect 32385 19225 32420 19260
rect 32430 19225 32465 19260
rect 32475 19225 32510 19260
rect 32520 19225 32555 19260
rect 32565 19225 32600 19260
rect 32610 19225 32645 19260
rect 32655 19225 32690 19260
rect 32700 19225 32735 19260
rect 32745 19225 32780 19260
rect 32790 19225 32825 19260
rect 32835 19225 32870 19260
rect 31305 19180 31340 19215
rect 31350 19180 31385 19215
rect 31395 19180 31430 19215
rect 31440 19180 31475 19215
rect 31485 19180 31520 19215
rect 31530 19180 31565 19215
rect 31575 19180 31610 19215
rect 31620 19180 31655 19215
rect 31665 19180 31700 19215
rect 31710 19180 31745 19215
rect 31755 19180 31790 19215
rect 31800 19180 31835 19215
rect 31845 19180 31880 19215
rect 31890 19180 31925 19215
rect 31935 19180 31970 19215
rect 31980 19180 32015 19215
rect 32025 19180 32060 19215
rect 32070 19180 32105 19215
rect 32115 19180 32150 19215
rect 32160 19180 32195 19215
rect 32205 19180 32240 19215
rect 32250 19180 32285 19215
rect 32295 19180 32330 19215
rect 32340 19180 32375 19215
rect 32385 19180 32420 19215
rect 32430 19180 32465 19215
rect 32475 19180 32510 19215
rect 32520 19180 32555 19215
rect 32565 19180 32600 19215
rect 32610 19180 32645 19215
rect 32655 19180 32690 19215
rect 32700 19180 32735 19215
rect 32745 19180 32780 19215
rect 32790 19180 32825 19215
rect 32835 19180 32870 19215
rect 31305 19135 31340 19170
rect 31350 19135 31385 19170
rect 31395 19135 31430 19170
rect 31440 19135 31475 19170
rect 31485 19135 31520 19170
rect 31530 19135 31565 19170
rect 31575 19135 31610 19170
rect 31620 19135 31655 19170
rect 31665 19135 31700 19170
rect 31710 19135 31745 19170
rect 31755 19135 31790 19170
rect 31800 19135 31835 19170
rect 31845 19135 31880 19170
rect 31890 19135 31925 19170
rect 31935 19135 31970 19170
rect 31980 19135 32015 19170
rect 32025 19135 32060 19170
rect 32070 19135 32105 19170
rect 32115 19135 32150 19170
rect 32160 19135 32195 19170
rect 32205 19135 32240 19170
rect 32250 19135 32285 19170
rect 32295 19135 32330 19170
rect 32340 19135 32375 19170
rect 32385 19135 32420 19170
rect 32430 19135 32465 19170
rect 32475 19135 32510 19170
rect 32520 19135 32555 19170
rect 32565 19135 32600 19170
rect 32610 19135 32645 19170
rect 32655 19135 32690 19170
rect 32700 19135 32735 19170
rect 32745 19135 32780 19170
rect 32790 19135 32825 19170
rect 32835 19135 32870 19170
rect 31305 19090 31340 19125
rect 31350 19090 31385 19125
rect 31395 19090 31430 19125
rect 31440 19090 31475 19125
rect 31485 19090 31520 19125
rect 31530 19090 31565 19125
rect 31575 19090 31610 19125
rect 31620 19090 31655 19125
rect 31665 19090 31700 19125
rect 31710 19090 31745 19125
rect 31755 19090 31790 19125
rect 31800 19090 31835 19125
rect 31845 19090 31880 19125
rect 31890 19090 31925 19125
rect 31935 19090 31970 19125
rect 31980 19090 32015 19125
rect 32025 19090 32060 19125
rect 32070 19090 32105 19125
rect 32115 19090 32150 19125
rect 32160 19090 32195 19125
rect 32205 19090 32240 19125
rect 32250 19090 32285 19125
rect 32295 19090 32330 19125
rect 32340 19090 32375 19125
rect 32385 19090 32420 19125
rect 32430 19090 32465 19125
rect 32475 19090 32510 19125
rect 32520 19090 32555 19125
rect 32565 19090 32600 19125
rect 32610 19090 32645 19125
rect 32655 19090 32690 19125
rect 32700 19090 32735 19125
rect 32745 19090 32780 19125
rect 32790 19090 32825 19125
rect 32835 19090 32870 19125
rect 31305 19045 31340 19080
rect 31350 19045 31385 19080
rect 31395 19045 31430 19080
rect 31440 19045 31475 19080
rect 31485 19045 31520 19080
rect 31530 19045 31565 19080
rect 31575 19045 31610 19080
rect 31620 19045 31655 19080
rect 31665 19045 31700 19080
rect 31710 19045 31745 19080
rect 31755 19045 31790 19080
rect 31800 19045 31835 19080
rect 31845 19045 31880 19080
rect 31890 19045 31925 19080
rect 31935 19045 31970 19080
rect 31980 19045 32015 19080
rect 32025 19045 32060 19080
rect 32070 19045 32105 19080
rect 32115 19045 32150 19080
rect 32160 19045 32195 19080
rect 32205 19045 32240 19080
rect 32250 19045 32285 19080
rect 32295 19045 32330 19080
rect 32340 19045 32375 19080
rect 32385 19045 32420 19080
rect 32430 19045 32465 19080
rect 32475 19045 32510 19080
rect 32520 19045 32555 19080
rect 32565 19045 32600 19080
rect 32610 19045 32645 19080
rect 32655 19045 32690 19080
rect 32700 19045 32735 19080
rect 32745 19045 32780 19080
rect 32790 19045 32825 19080
rect 32835 19045 32870 19080
rect 31305 19000 31340 19035
rect 31350 19000 31385 19035
rect 31395 19000 31430 19035
rect 31440 19000 31475 19035
rect 31485 19000 31520 19035
rect 31530 19000 31565 19035
rect 31575 19000 31610 19035
rect 31620 19000 31655 19035
rect 31665 19000 31700 19035
rect 31710 19000 31745 19035
rect 31755 19000 31790 19035
rect 31800 19000 31835 19035
rect 31845 19000 31880 19035
rect 31890 19000 31925 19035
rect 31935 19000 31970 19035
rect 31980 19000 32015 19035
rect 32025 19000 32060 19035
rect 32070 19000 32105 19035
rect 32115 19000 32150 19035
rect 32160 19000 32195 19035
rect 32205 19000 32240 19035
rect 32250 19000 32285 19035
rect 32295 19000 32330 19035
rect 32340 19000 32375 19035
rect 32385 19000 32420 19035
rect 32430 19000 32465 19035
rect 32475 19000 32510 19035
rect 32520 19000 32555 19035
rect 32565 19000 32600 19035
rect 32610 19000 32645 19035
rect 32655 19000 32690 19035
rect 32700 19000 32735 19035
rect 32745 19000 32780 19035
rect 32790 19000 32825 19035
rect 32835 19000 32870 19035
rect 31305 18955 31340 18990
rect 31350 18955 31385 18990
rect 31395 18955 31430 18990
rect 31440 18955 31475 18990
rect 31485 18955 31520 18990
rect 31530 18955 31565 18990
rect 31575 18955 31610 18990
rect 31620 18955 31655 18990
rect 31665 18955 31700 18990
rect 31710 18955 31745 18990
rect 31755 18955 31790 18990
rect 31800 18955 31835 18990
rect 31845 18955 31880 18990
rect 31890 18955 31925 18990
rect 31935 18955 31970 18990
rect 31980 18955 32015 18990
rect 32025 18955 32060 18990
rect 32070 18955 32105 18990
rect 32115 18955 32150 18990
rect 32160 18955 32195 18990
rect 32205 18955 32240 18990
rect 32250 18955 32285 18990
rect 32295 18955 32330 18990
rect 32340 18955 32375 18990
rect 32385 18955 32420 18990
rect 32430 18955 32465 18990
rect 32475 18955 32510 18990
rect 32520 18955 32555 18990
rect 32565 18955 32600 18990
rect 32610 18955 32645 18990
rect 32655 18955 32690 18990
rect 32700 18955 32735 18990
rect 32745 18955 32780 18990
rect 32790 18955 32825 18990
rect 32835 18955 32870 18990
rect 31305 18910 31340 18945
rect 31350 18910 31385 18945
rect 31395 18910 31430 18945
rect 31440 18910 31475 18945
rect 31485 18910 31520 18945
rect 31530 18910 31565 18945
rect 31575 18910 31610 18945
rect 31620 18910 31655 18945
rect 31665 18910 31700 18945
rect 31710 18910 31745 18945
rect 31755 18910 31790 18945
rect 31800 18910 31835 18945
rect 31845 18910 31880 18945
rect 31890 18910 31925 18945
rect 31935 18910 31970 18945
rect 31980 18910 32015 18945
rect 32025 18910 32060 18945
rect 32070 18910 32105 18945
rect 32115 18910 32150 18945
rect 32160 18910 32195 18945
rect 32205 18910 32240 18945
rect 32250 18910 32285 18945
rect 32295 18910 32330 18945
rect 32340 18910 32375 18945
rect 32385 18910 32420 18945
rect 32430 18910 32465 18945
rect 32475 18910 32510 18945
rect 32520 18910 32555 18945
rect 32565 18910 32600 18945
rect 32610 18910 32645 18945
rect 32655 18910 32690 18945
rect 32700 18910 32735 18945
rect 32745 18910 32780 18945
rect 32790 18910 32825 18945
rect 32835 18910 32870 18945
rect 31305 18865 31340 18900
rect 31350 18865 31385 18900
rect 31395 18865 31430 18900
rect 31440 18865 31475 18900
rect 31485 18865 31520 18900
rect 31530 18865 31565 18900
rect 31575 18865 31610 18900
rect 31620 18865 31655 18900
rect 31665 18865 31700 18900
rect 31710 18865 31745 18900
rect 31755 18865 31790 18900
rect 31800 18865 31835 18900
rect 31845 18865 31880 18900
rect 31890 18865 31925 18900
rect 31935 18865 31970 18900
rect 31980 18865 32015 18900
rect 32025 18865 32060 18900
rect 32070 18865 32105 18900
rect 32115 18865 32150 18900
rect 32160 18865 32195 18900
rect 32205 18865 32240 18900
rect 32250 18865 32285 18900
rect 32295 18865 32330 18900
rect 32340 18865 32375 18900
rect 32385 18865 32420 18900
rect 32430 18865 32465 18900
rect 32475 18865 32510 18900
rect 32520 18865 32555 18900
rect 32565 18865 32600 18900
rect 32610 18865 32645 18900
rect 32655 18865 32690 18900
rect 32700 18865 32735 18900
rect 32745 18865 32780 18900
rect 32790 18865 32825 18900
rect 32835 18865 32870 18900
rect 31305 18820 31340 18855
rect 31350 18820 31385 18855
rect 31395 18820 31430 18855
rect 31440 18820 31475 18855
rect 31485 18820 31520 18855
rect 31530 18820 31565 18855
rect 31575 18820 31610 18855
rect 31620 18820 31655 18855
rect 31665 18820 31700 18855
rect 31710 18820 31745 18855
rect 31755 18820 31790 18855
rect 31800 18820 31835 18855
rect 31845 18820 31880 18855
rect 31890 18820 31925 18855
rect 31935 18820 31970 18855
rect 31980 18820 32015 18855
rect 32025 18820 32060 18855
rect 32070 18820 32105 18855
rect 32115 18820 32150 18855
rect 32160 18820 32195 18855
rect 32205 18820 32240 18855
rect 32250 18820 32285 18855
rect 32295 18820 32330 18855
rect 32340 18820 32375 18855
rect 32385 18820 32420 18855
rect 32430 18820 32465 18855
rect 32475 18820 32510 18855
rect 32520 18820 32555 18855
rect 32565 18820 32600 18855
rect 32610 18820 32645 18855
rect 32655 18820 32690 18855
rect 32700 18820 32735 18855
rect 32745 18820 32780 18855
rect 32790 18820 32825 18855
rect 32835 18820 32870 18855
rect 31305 18775 31340 18810
rect 31350 18775 31385 18810
rect 31395 18775 31430 18810
rect 31440 18775 31475 18810
rect 31485 18775 31520 18810
rect 31530 18775 31565 18810
rect 31575 18775 31610 18810
rect 31620 18775 31655 18810
rect 31665 18775 31700 18810
rect 31710 18775 31745 18810
rect 31755 18775 31790 18810
rect 31800 18775 31835 18810
rect 31845 18775 31880 18810
rect 31890 18775 31925 18810
rect 31935 18775 31970 18810
rect 31980 18775 32015 18810
rect 32025 18775 32060 18810
rect 32070 18775 32105 18810
rect 32115 18775 32150 18810
rect 32160 18775 32195 18810
rect 32205 18775 32240 18810
rect 32250 18775 32285 18810
rect 32295 18775 32330 18810
rect 32340 18775 32375 18810
rect 32385 18775 32420 18810
rect 32430 18775 32465 18810
rect 32475 18775 32510 18810
rect 32520 18775 32555 18810
rect 32565 18775 32600 18810
rect 32610 18775 32645 18810
rect 32655 18775 32690 18810
rect 32700 18775 32735 18810
rect 32745 18775 32780 18810
rect 32790 18775 32825 18810
rect 32835 18775 32870 18810
rect 31305 18730 31340 18765
rect 31350 18730 31385 18765
rect 31395 18730 31430 18765
rect 31440 18730 31475 18765
rect 31485 18730 31520 18765
rect 31530 18730 31565 18765
rect 31575 18730 31610 18765
rect 31620 18730 31655 18765
rect 31665 18730 31700 18765
rect 31710 18730 31745 18765
rect 31755 18730 31790 18765
rect 31800 18730 31835 18765
rect 31845 18730 31880 18765
rect 31890 18730 31925 18765
rect 31935 18730 31970 18765
rect 31980 18730 32015 18765
rect 32025 18730 32060 18765
rect 32070 18730 32105 18765
rect 32115 18730 32150 18765
rect 32160 18730 32195 18765
rect 32205 18730 32240 18765
rect 32250 18730 32285 18765
rect 32295 18730 32330 18765
rect 32340 18730 32375 18765
rect 32385 18730 32420 18765
rect 32430 18730 32465 18765
rect 32475 18730 32510 18765
rect 32520 18730 32555 18765
rect 32565 18730 32600 18765
rect 32610 18730 32645 18765
rect 32655 18730 32690 18765
rect 32700 18730 32735 18765
rect 32745 18730 32780 18765
rect 32790 18730 32825 18765
rect 32835 18730 32870 18765
rect 31305 18685 31340 18720
rect 31350 18685 31385 18720
rect 31395 18685 31430 18720
rect 31440 18685 31475 18720
rect 31485 18685 31520 18720
rect 31530 18685 31565 18720
rect 31575 18685 31610 18720
rect 31620 18685 31655 18720
rect 31665 18685 31700 18720
rect 31710 18685 31745 18720
rect 31755 18685 31790 18720
rect 31800 18685 31835 18720
rect 31845 18685 31880 18720
rect 31890 18685 31925 18720
rect 31935 18685 31970 18720
rect 31980 18685 32015 18720
rect 32025 18685 32060 18720
rect 32070 18685 32105 18720
rect 32115 18685 32150 18720
rect 32160 18685 32195 18720
rect 32205 18685 32240 18720
rect 32250 18685 32285 18720
rect 32295 18685 32330 18720
rect 32340 18685 32375 18720
rect 32385 18685 32420 18720
rect 32430 18685 32465 18720
rect 32475 18685 32510 18720
rect 32520 18685 32555 18720
rect 32565 18685 32600 18720
rect 32610 18685 32645 18720
rect 32655 18685 32690 18720
rect 32700 18685 32735 18720
rect 32745 18685 32780 18720
rect 32790 18685 32825 18720
rect 32835 18685 32870 18720
rect 31305 18640 31340 18675
rect 31350 18640 31385 18675
rect 31395 18640 31430 18675
rect 31440 18640 31475 18675
rect 31485 18640 31520 18675
rect 31530 18640 31565 18675
rect 31575 18640 31610 18675
rect 31620 18640 31655 18675
rect 31665 18640 31700 18675
rect 31710 18640 31745 18675
rect 31755 18640 31790 18675
rect 31800 18640 31835 18675
rect 31845 18640 31880 18675
rect 31890 18640 31925 18675
rect 31935 18640 31970 18675
rect 31980 18640 32015 18675
rect 32025 18640 32060 18675
rect 32070 18640 32105 18675
rect 32115 18640 32150 18675
rect 32160 18640 32195 18675
rect 32205 18640 32240 18675
rect 32250 18640 32285 18675
rect 32295 18640 32330 18675
rect 32340 18640 32375 18675
rect 32385 18640 32420 18675
rect 32430 18640 32465 18675
rect 32475 18640 32510 18675
rect 32520 18640 32555 18675
rect 32565 18640 32600 18675
rect 32610 18640 32645 18675
rect 32655 18640 32690 18675
rect 32700 18640 32735 18675
rect 32745 18640 32780 18675
rect 32790 18640 32825 18675
rect 32835 18640 32870 18675
rect 31305 18595 31340 18630
rect 31350 18595 31385 18630
rect 31395 18595 31430 18630
rect 31440 18595 31475 18630
rect 31485 18595 31520 18630
rect 31530 18595 31565 18630
rect 31575 18595 31610 18630
rect 31620 18595 31655 18630
rect 31665 18595 31700 18630
rect 31710 18595 31745 18630
rect 31755 18595 31790 18630
rect 31800 18595 31835 18630
rect 31845 18595 31880 18630
rect 31890 18595 31925 18630
rect 31935 18595 31970 18630
rect 31980 18595 32015 18630
rect 32025 18595 32060 18630
rect 32070 18595 32105 18630
rect 32115 18595 32150 18630
rect 32160 18595 32195 18630
rect 32205 18595 32240 18630
rect 32250 18595 32285 18630
rect 32295 18595 32330 18630
rect 32340 18595 32375 18630
rect 32385 18595 32420 18630
rect 32430 18595 32465 18630
rect 32475 18595 32510 18630
rect 32520 18595 32555 18630
rect 32565 18595 32600 18630
rect 32610 18595 32645 18630
rect 32655 18595 32690 18630
rect 32700 18595 32735 18630
rect 32745 18595 32780 18630
rect 32790 18595 32825 18630
rect 32835 18595 32870 18630
rect 31305 18550 31340 18585
rect 31350 18550 31385 18585
rect 31395 18550 31430 18585
rect 31440 18550 31475 18585
rect 31485 18550 31520 18585
rect 31530 18550 31565 18585
rect 31575 18550 31610 18585
rect 31620 18550 31655 18585
rect 31665 18550 31700 18585
rect 31710 18550 31745 18585
rect 31755 18550 31790 18585
rect 31800 18550 31835 18585
rect 31845 18550 31880 18585
rect 31890 18550 31925 18585
rect 31935 18550 31970 18585
rect 31980 18550 32015 18585
rect 32025 18550 32060 18585
rect 32070 18550 32105 18585
rect 32115 18550 32150 18585
rect 32160 18550 32195 18585
rect 32205 18550 32240 18585
rect 32250 18550 32285 18585
rect 32295 18550 32330 18585
rect 32340 18550 32375 18585
rect 32385 18550 32420 18585
rect 32430 18550 32465 18585
rect 32475 18550 32510 18585
rect 32520 18550 32555 18585
rect 32565 18550 32600 18585
rect 32610 18550 32645 18585
rect 32655 18550 32690 18585
rect 32700 18550 32735 18585
rect 32745 18550 32780 18585
rect 32790 18550 32825 18585
rect 32835 18550 32870 18585
rect 31305 18505 31340 18540
rect 31350 18505 31385 18540
rect 31395 18505 31430 18540
rect 31440 18505 31475 18540
rect 31485 18505 31520 18540
rect 31530 18505 31565 18540
rect 31575 18505 31610 18540
rect 31620 18505 31655 18540
rect 31665 18505 31700 18540
rect 31710 18505 31745 18540
rect 31755 18505 31790 18540
rect 31800 18505 31835 18540
rect 31845 18505 31880 18540
rect 31890 18505 31925 18540
rect 31935 18505 31970 18540
rect 31980 18505 32015 18540
rect 32025 18505 32060 18540
rect 32070 18505 32105 18540
rect 32115 18505 32150 18540
rect 32160 18505 32195 18540
rect 32205 18505 32240 18540
rect 32250 18505 32285 18540
rect 32295 18505 32330 18540
rect 32340 18505 32375 18540
rect 32385 18505 32420 18540
rect 32430 18505 32465 18540
rect 32475 18505 32510 18540
rect 32520 18505 32555 18540
rect 32565 18505 32600 18540
rect 32610 18505 32645 18540
rect 32655 18505 32690 18540
rect 32700 18505 32735 18540
rect 32745 18505 32780 18540
rect 32790 18505 32825 18540
rect 32835 18505 32870 18540
rect 31305 18460 31340 18495
rect 31350 18460 31385 18495
rect 31395 18460 31430 18495
rect 31440 18460 31475 18495
rect 31485 18460 31520 18495
rect 31530 18460 31565 18495
rect 31575 18460 31610 18495
rect 31620 18460 31655 18495
rect 31665 18460 31700 18495
rect 31710 18460 31745 18495
rect 31755 18460 31790 18495
rect 31800 18460 31835 18495
rect 31845 18460 31880 18495
rect 31890 18460 31925 18495
rect 31935 18460 31970 18495
rect 31980 18460 32015 18495
rect 32025 18460 32060 18495
rect 32070 18460 32105 18495
rect 32115 18460 32150 18495
rect 32160 18460 32195 18495
rect 32205 18460 32240 18495
rect 32250 18460 32285 18495
rect 32295 18460 32330 18495
rect 32340 18460 32375 18495
rect 32385 18460 32420 18495
rect 32430 18460 32465 18495
rect 32475 18460 32510 18495
rect 32520 18460 32555 18495
rect 32565 18460 32600 18495
rect 32610 18460 32645 18495
rect 32655 18460 32690 18495
rect 32700 18460 32735 18495
rect 32745 18460 32780 18495
rect 32790 18460 32825 18495
rect 32835 18460 32870 18495
rect 31305 18415 31340 18450
rect 31350 18415 31385 18450
rect 31395 18415 31430 18450
rect 31440 18415 31475 18450
rect 31485 18415 31520 18450
rect 31530 18415 31565 18450
rect 31575 18415 31610 18450
rect 31620 18415 31655 18450
rect 31665 18415 31700 18450
rect 31710 18415 31745 18450
rect 31755 18415 31790 18450
rect 31800 18415 31835 18450
rect 31845 18415 31880 18450
rect 31890 18415 31925 18450
rect 31935 18415 31970 18450
rect 31980 18415 32015 18450
rect 32025 18415 32060 18450
rect 32070 18415 32105 18450
rect 32115 18415 32150 18450
rect 32160 18415 32195 18450
rect 32205 18415 32240 18450
rect 32250 18415 32285 18450
rect 32295 18415 32330 18450
rect 32340 18415 32375 18450
rect 32385 18415 32420 18450
rect 32430 18415 32465 18450
rect 32475 18415 32510 18450
rect 32520 18415 32555 18450
rect 32565 18415 32600 18450
rect 32610 18415 32645 18450
rect 32655 18415 32690 18450
rect 32700 18415 32735 18450
rect 32745 18415 32780 18450
rect 32790 18415 32825 18450
rect 32835 18415 32870 18450
rect 31305 18370 31340 18405
rect 31350 18370 31385 18405
rect 31395 18370 31430 18405
rect 31440 18370 31475 18405
rect 31485 18370 31520 18405
rect 31530 18370 31565 18405
rect 31575 18370 31610 18405
rect 31620 18370 31655 18405
rect 31665 18370 31700 18405
rect 31710 18370 31745 18405
rect 31755 18370 31790 18405
rect 31800 18370 31835 18405
rect 31845 18370 31880 18405
rect 31890 18370 31925 18405
rect 31935 18370 31970 18405
rect 31980 18370 32015 18405
rect 32025 18370 32060 18405
rect 32070 18370 32105 18405
rect 32115 18370 32150 18405
rect 32160 18370 32195 18405
rect 32205 18370 32240 18405
rect 32250 18370 32285 18405
rect 32295 18370 32330 18405
rect 32340 18370 32375 18405
rect 32385 18370 32420 18405
rect 32430 18370 32465 18405
rect 32475 18370 32510 18405
rect 32520 18370 32555 18405
rect 32565 18370 32600 18405
rect 32610 18370 32645 18405
rect 32655 18370 32690 18405
rect 32700 18370 32735 18405
rect 32745 18370 32780 18405
rect 32790 18370 32825 18405
rect 32835 18370 32870 18405
rect 31305 18325 31340 18360
rect 31350 18325 31385 18360
rect 31395 18325 31430 18360
rect 31440 18325 31475 18360
rect 31485 18325 31520 18360
rect 31530 18325 31565 18360
rect 31575 18325 31610 18360
rect 31620 18325 31655 18360
rect 31665 18325 31700 18360
rect 31710 18325 31745 18360
rect 31755 18325 31790 18360
rect 31800 18325 31835 18360
rect 31845 18325 31880 18360
rect 31890 18325 31925 18360
rect 31935 18325 31970 18360
rect 31980 18325 32015 18360
rect 32025 18325 32060 18360
rect 32070 18325 32105 18360
rect 32115 18325 32150 18360
rect 32160 18325 32195 18360
rect 32205 18325 32240 18360
rect 32250 18325 32285 18360
rect 32295 18325 32330 18360
rect 32340 18325 32375 18360
rect 32385 18325 32420 18360
rect 32430 18325 32465 18360
rect 32475 18325 32510 18360
rect 32520 18325 32555 18360
rect 32565 18325 32600 18360
rect 32610 18325 32645 18360
rect 32655 18325 32690 18360
rect 32700 18325 32735 18360
rect 32745 18325 32780 18360
rect 32790 18325 32825 18360
rect 32835 18325 32870 18360
rect 31305 18280 31340 18315
rect 31350 18280 31385 18315
rect 31395 18280 31430 18315
rect 31440 18280 31475 18315
rect 31485 18280 31520 18315
rect 31530 18280 31565 18315
rect 31575 18280 31610 18315
rect 31620 18280 31655 18315
rect 31665 18280 31700 18315
rect 31710 18280 31745 18315
rect 31755 18280 31790 18315
rect 31800 18280 31835 18315
rect 31845 18280 31880 18315
rect 31890 18280 31925 18315
rect 31935 18280 31970 18315
rect 31980 18280 32015 18315
rect 32025 18280 32060 18315
rect 32070 18280 32105 18315
rect 32115 18280 32150 18315
rect 32160 18280 32195 18315
rect 32205 18280 32240 18315
rect 32250 18280 32285 18315
rect 32295 18280 32330 18315
rect 32340 18280 32375 18315
rect 32385 18280 32420 18315
rect 32430 18280 32465 18315
rect 32475 18280 32510 18315
rect 32520 18280 32555 18315
rect 32565 18280 32600 18315
rect 32610 18280 32645 18315
rect 32655 18280 32690 18315
rect 32700 18280 32735 18315
rect 32745 18280 32780 18315
rect 32790 18280 32825 18315
rect 32835 18280 32870 18315
rect 31305 18235 31340 18270
rect 31350 18235 31385 18270
rect 31395 18235 31430 18270
rect 31440 18235 31475 18270
rect 31485 18235 31520 18270
rect 31530 18235 31565 18270
rect 31575 18235 31610 18270
rect 31620 18235 31655 18270
rect 31665 18235 31700 18270
rect 31710 18235 31745 18270
rect 31755 18235 31790 18270
rect 31800 18235 31835 18270
rect 31845 18235 31880 18270
rect 31890 18235 31925 18270
rect 31935 18235 31970 18270
rect 31980 18235 32015 18270
rect 32025 18235 32060 18270
rect 32070 18235 32105 18270
rect 32115 18235 32150 18270
rect 32160 18235 32195 18270
rect 32205 18235 32240 18270
rect 32250 18235 32285 18270
rect 32295 18235 32330 18270
rect 32340 18235 32375 18270
rect 32385 18235 32420 18270
rect 32430 18235 32465 18270
rect 32475 18235 32510 18270
rect 32520 18235 32555 18270
rect 32565 18235 32600 18270
rect 32610 18235 32645 18270
rect 32655 18235 32690 18270
rect 32700 18235 32735 18270
rect 32745 18235 32780 18270
rect 32790 18235 32825 18270
rect 32835 18235 32870 18270
rect 31305 18190 31340 18225
rect 31350 18190 31385 18225
rect 31395 18190 31430 18225
rect 31440 18190 31475 18225
rect 31485 18190 31520 18225
rect 31530 18190 31565 18225
rect 31575 18190 31610 18225
rect 31620 18190 31655 18225
rect 31665 18190 31700 18225
rect 31710 18190 31745 18225
rect 31755 18190 31790 18225
rect 31800 18190 31835 18225
rect 31845 18190 31880 18225
rect 31890 18190 31925 18225
rect 31935 18190 31970 18225
rect 31980 18190 32015 18225
rect 32025 18190 32060 18225
rect 32070 18190 32105 18225
rect 32115 18190 32150 18225
rect 32160 18190 32195 18225
rect 32205 18190 32240 18225
rect 32250 18190 32285 18225
rect 32295 18190 32330 18225
rect 32340 18190 32375 18225
rect 32385 18190 32420 18225
rect 32430 18190 32465 18225
rect 32475 18190 32510 18225
rect 32520 18190 32555 18225
rect 32565 18190 32600 18225
rect 32610 18190 32645 18225
rect 32655 18190 32690 18225
rect 32700 18190 32735 18225
rect 32745 18190 32780 18225
rect 32790 18190 32825 18225
rect 32835 18190 32870 18225
rect 31305 18145 31340 18180
rect 31350 18145 31385 18180
rect 31395 18145 31430 18180
rect 31440 18145 31475 18180
rect 31485 18145 31520 18180
rect 31530 18145 31565 18180
rect 31575 18145 31610 18180
rect 31620 18145 31655 18180
rect 31665 18145 31700 18180
rect 31710 18145 31745 18180
rect 31755 18145 31790 18180
rect 31800 18145 31835 18180
rect 31845 18145 31880 18180
rect 31890 18145 31925 18180
rect 31935 18145 31970 18180
rect 31980 18145 32015 18180
rect 32025 18145 32060 18180
rect 32070 18145 32105 18180
rect 32115 18145 32150 18180
rect 32160 18145 32195 18180
rect 32205 18145 32240 18180
rect 32250 18145 32285 18180
rect 32295 18145 32330 18180
rect 32340 18145 32375 18180
rect 32385 18145 32420 18180
rect 32430 18145 32465 18180
rect 32475 18145 32510 18180
rect 32520 18145 32555 18180
rect 32565 18145 32600 18180
rect 32610 18145 32645 18180
rect 32655 18145 32690 18180
rect 32700 18145 32735 18180
rect 32745 18145 32780 18180
rect 32790 18145 32825 18180
rect 32835 18145 32870 18180
rect 31305 18100 31340 18135
rect 31350 18100 31385 18135
rect 31395 18100 31430 18135
rect 31440 18100 31475 18135
rect 31485 18100 31520 18135
rect 31530 18100 31565 18135
rect 31575 18100 31610 18135
rect 31620 18100 31655 18135
rect 31665 18100 31700 18135
rect 31710 18100 31745 18135
rect 31755 18100 31790 18135
rect 31800 18100 31835 18135
rect 31845 18100 31880 18135
rect 31890 18100 31925 18135
rect 31935 18100 31970 18135
rect 31980 18100 32015 18135
rect 32025 18100 32060 18135
rect 32070 18100 32105 18135
rect 32115 18100 32150 18135
rect 32160 18100 32195 18135
rect 32205 18100 32240 18135
rect 32250 18100 32285 18135
rect 32295 18100 32330 18135
rect 32340 18100 32375 18135
rect 32385 18100 32420 18135
rect 32430 18100 32465 18135
rect 32475 18100 32510 18135
rect 32520 18100 32555 18135
rect 32565 18100 32600 18135
rect 32610 18100 32645 18135
rect 32655 18100 32690 18135
rect 32700 18100 32735 18135
rect 32745 18100 32780 18135
rect 32790 18100 32825 18135
rect 32835 18100 32870 18135
rect 31305 18055 31340 18090
rect 31350 18055 31385 18090
rect 31395 18055 31430 18090
rect 31440 18055 31475 18090
rect 31485 18055 31520 18090
rect 31530 18055 31565 18090
rect 31575 18055 31610 18090
rect 31620 18055 31655 18090
rect 31665 18055 31700 18090
rect 31710 18055 31745 18090
rect 31755 18055 31790 18090
rect 31800 18055 31835 18090
rect 31845 18055 31880 18090
rect 31890 18055 31925 18090
rect 31935 18055 31970 18090
rect 31980 18055 32015 18090
rect 32025 18055 32060 18090
rect 32070 18055 32105 18090
rect 32115 18055 32150 18090
rect 32160 18055 32195 18090
rect 32205 18055 32240 18090
rect 32250 18055 32285 18090
rect 32295 18055 32330 18090
rect 32340 18055 32375 18090
rect 32385 18055 32420 18090
rect 32430 18055 32465 18090
rect 32475 18055 32510 18090
rect 32520 18055 32555 18090
rect 32565 18055 32600 18090
rect 32610 18055 32645 18090
rect 32655 18055 32690 18090
rect 32700 18055 32735 18090
rect 32745 18055 32780 18090
rect 32790 18055 32825 18090
rect 32835 18055 32870 18090
rect 31305 18010 31340 18045
rect 31350 18010 31385 18045
rect 31395 18010 31430 18045
rect 31440 18010 31475 18045
rect 31485 18010 31520 18045
rect 31530 18010 31565 18045
rect 31575 18010 31610 18045
rect 31620 18010 31655 18045
rect 31665 18010 31700 18045
rect 31710 18010 31745 18045
rect 31755 18010 31790 18045
rect 31800 18010 31835 18045
rect 31845 18010 31880 18045
rect 31890 18010 31925 18045
rect 31935 18010 31970 18045
rect 31980 18010 32015 18045
rect 32025 18010 32060 18045
rect 32070 18010 32105 18045
rect 32115 18010 32150 18045
rect 32160 18010 32195 18045
rect 32205 18010 32240 18045
rect 32250 18010 32285 18045
rect 32295 18010 32330 18045
rect 32340 18010 32375 18045
rect 32385 18010 32420 18045
rect 32430 18010 32465 18045
rect 32475 18010 32510 18045
rect 32520 18010 32555 18045
rect 32565 18010 32600 18045
rect 32610 18010 32645 18045
rect 32655 18010 32690 18045
rect 32700 18010 32735 18045
rect 32745 18010 32780 18045
rect 32790 18010 32825 18045
rect 32835 18010 32870 18045
rect 31305 17965 31340 18000
rect 31350 17965 31385 18000
rect 31395 17965 31430 18000
rect 31440 17965 31475 18000
rect 31485 17965 31520 18000
rect 31530 17965 31565 18000
rect 31575 17965 31610 18000
rect 31620 17965 31655 18000
rect 31665 17965 31700 18000
rect 31710 17965 31745 18000
rect 31755 17965 31790 18000
rect 31800 17965 31835 18000
rect 31845 17965 31880 18000
rect 31890 17965 31925 18000
rect 31935 17965 31970 18000
rect 31980 17965 32015 18000
rect 32025 17965 32060 18000
rect 32070 17965 32105 18000
rect 32115 17965 32150 18000
rect 32160 17965 32195 18000
rect 32205 17965 32240 18000
rect 32250 17965 32285 18000
rect 32295 17965 32330 18000
rect 32340 17965 32375 18000
rect 32385 17965 32420 18000
rect 32430 17965 32465 18000
rect 32475 17965 32510 18000
rect 32520 17965 32555 18000
rect 32565 17965 32600 18000
rect 32610 17965 32645 18000
rect 32655 17965 32690 18000
rect 32700 17965 32735 18000
rect 32745 17965 32780 18000
rect 32790 17965 32825 18000
rect 32835 17965 32870 18000
rect 31305 17920 31340 17955
rect 31350 17920 31385 17955
rect 31395 17920 31430 17955
rect 31440 17920 31475 17955
rect 31485 17920 31520 17955
rect 31530 17920 31565 17955
rect 31575 17920 31610 17955
rect 31620 17920 31655 17955
rect 31665 17920 31700 17955
rect 31710 17920 31745 17955
rect 31755 17920 31790 17955
rect 31800 17920 31835 17955
rect 31845 17920 31880 17955
rect 31890 17920 31925 17955
rect 31935 17920 31970 17955
rect 31980 17920 32015 17955
rect 32025 17920 32060 17955
rect 32070 17920 32105 17955
rect 32115 17920 32150 17955
rect 32160 17920 32195 17955
rect 32205 17920 32240 17955
rect 32250 17920 32285 17955
rect 32295 17920 32330 17955
rect 32340 17920 32375 17955
rect 32385 17920 32420 17955
rect 32430 17920 32465 17955
rect 32475 17920 32510 17955
rect 32520 17920 32555 17955
rect 32565 17920 32600 17955
rect 32610 17920 32645 17955
rect 32655 17920 32690 17955
rect 32700 17920 32735 17955
rect 32745 17920 32780 17955
rect 32790 17920 32825 17955
rect 32835 17920 32870 17955
rect 31305 17875 31340 17910
rect 31350 17875 31385 17910
rect 31395 17875 31430 17910
rect 31440 17875 31475 17910
rect 31485 17875 31520 17910
rect 31530 17875 31565 17910
rect 31575 17875 31610 17910
rect 31620 17875 31655 17910
rect 31665 17875 31700 17910
rect 31710 17875 31745 17910
rect 31755 17875 31790 17910
rect 31800 17875 31835 17910
rect 31845 17875 31880 17910
rect 31890 17875 31925 17910
rect 31935 17875 31970 17910
rect 31980 17875 32015 17910
rect 32025 17875 32060 17910
rect 32070 17875 32105 17910
rect 32115 17875 32150 17910
rect 32160 17875 32195 17910
rect 32205 17875 32240 17910
rect 32250 17875 32285 17910
rect 32295 17875 32330 17910
rect 32340 17875 32375 17910
rect 32385 17875 32420 17910
rect 32430 17875 32465 17910
rect 32475 17875 32510 17910
rect 32520 17875 32555 17910
rect 32565 17875 32600 17910
rect 32610 17875 32645 17910
rect 32655 17875 32690 17910
rect 32700 17875 32735 17910
rect 32745 17875 32780 17910
rect 32790 17875 32825 17910
rect 32835 17875 32870 17910
rect 31305 17830 31340 17865
rect 31350 17830 31385 17865
rect 31395 17830 31430 17865
rect 31440 17830 31475 17865
rect 31485 17830 31520 17865
rect 31530 17830 31565 17865
rect 31575 17830 31610 17865
rect 31620 17830 31655 17865
rect 31665 17830 31700 17865
rect 31710 17830 31745 17865
rect 31755 17830 31790 17865
rect 31800 17830 31835 17865
rect 31845 17830 31880 17865
rect 31890 17830 31925 17865
rect 31935 17830 31970 17865
rect 31980 17830 32015 17865
rect 32025 17830 32060 17865
rect 32070 17830 32105 17865
rect 32115 17830 32150 17865
rect 32160 17830 32195 17865
rect 32205 17830 32240 17865
rect 32250 17830 32285 17865
rect 32295 17830 32330 17865
rect 32340 17830 32375 17865
rect 32385 17830 32420 17865
rect 32430 17830 32465 17865
rect 32475 17830 32510 17865
rect 32520 17830 32555 17865
rect 32565 17830 32600 17865
rect 32610 17830 32645 17865
rect 32655 17830 32690 17865
rect 32700 17830 32735 17865
rect 32745 17830 32780 17865
rect 32790 17830 32825 17865
rect 32835 17830 32870 17865
rect 31305 17785 31340 17820
rect 31350 17785 31385 17820
rect 31395 17785 31430 17820
rect 31440 17785 31475 17820
rect 31485 17785 31520 17820
rect 31530 17785 31565 17820
rect 31575 17785 31610 17820
rect 31620 17785 31655 17820
rect 31665 17785 31700 17820
rect 31710 17785 31745 17820
rect 31755 17785 31790 17820
rect 31800 17785 31835 17820
rect 31845 17785 31880 17820
rect 31890 17785 31925 17820
rect 31935 17785 31970 17820
rect 31980 17785 32015 17820
rect 32025 17785 32060 17820
rect 32070 17785 32105 17820
rect 32115 17785 32150 17820
rect 32160 17785 32195 17820
rect 32205 17785 32240 17820
rect 32250 17785 32285 17820
rect 32295 17785 32330 17820
rect 32340 17785 32375 17820
rect 32385 17785 32420 17820
rect 32430 17785 32465 17820
rect 32475 17785 32510 17820
rect 32520 17785 32555 17820
rect 32565 17785 32600 17820
rect 32610 17785 32645 17820
rect 32655 17785 32690 17820
rect 32700 17785 32735 17820
rect 32745 17785 32780 17820
rect 32790 17785 32825 17820
rect 32835 17785 32870 17820
rect 31305 17740 31340 17775
rect 31350 17740 31385 17775
rect 31395 17740 31430 17775
rect 31440 17740 31475 17775
rect 31485 17740 31520 17775
rect 31530 17740 31565 17775
rect 31575 17740 31610 17775
rect 31620 17740 31655 17775
rect 31665 17740 31700 17775
rect 31710 17740 31745 17775
rect 31755 17740 31790 17775
rect 31800 17740 31835 17775
rect 31845 17740 31880 17775
rect 31890 17740 31925 17775
rect 31935 17740 31970 17775
rect 31980 17740 32015 17775
rect 32025 17740 32060 17775
rect 32070 17740 32105 17775
rect 32115 17740 32150 17775
rect 32160 17740 32195 17775
rect 32205 17740 32240 17775
rect 32250 17740 32285 17775
rect 32295 17740 32330 17775
rect 32340 17740 32375 17775
rect 32385 17740 32420 17775
rect 32430 17740 32465 17775
rect 32475 17740 32510 17775
rect 32520 17740 32555 17775
rect 32565 17740 32600 17775
rect 32610 17740 32645 17775
rect 32655 17740 32690 17775
rect 32700 17740 32735 17775
rect 32745 17740 32780 17775
rect 32790 17740 32825 17775
rect 32835 17740 32870 17775
rect -38755 9595 -38720 9630
rect -38710 9595 -38675 9630
rect -38665 9595 -38630 9630
rect -38620 9595 -38585 9630
rect -38575 9595 -38540 9630
rect -38530 9595 -38495 9630
rect -38485 9595 -38450 9630
rect -38440 9595 -38405 9630
rect -38395 9595 -38360 9630
rect -38350 9595 -38315 9630
rect -38305 9595 -38270 9630
rect -38260 9595 -38225 9630
rect -38215 9595 -38180 9630
rect -38170 9595 -38135 9630
rect -38125 9595 -38090 9630
rect -38080 9595 -38045 9630
rect -38035 9595 -38000 9630
rect -37990 9595 -37955 9630
rect -37945 9595 -37910 9630
rect -37900 9595 -37865 9630
rect -37855 9595 -37820 9630
rect -37810 9595 -37775 9630
rect -37765 9595 -37730 9630
rect -37720 9595 -37685 9630
rect -37675 9595 -37640 9630
rect -37630 9595 -37595 9630
rect -37585 9595 -37550 9630
rect -37540 9595 -37505 9630
rect -37495 9595 -37460 9630
rect -37450 9595 -37415 9630
rect -37405 9595 -37370 9630
rect -37360 9595 -37325 9630
rect -37315 9595 -37280 9630
rect -37270 9595 -37235 9630
rect -37225 9595 -37190 9630
rect -38755 9550 -38720 9585
rect -38710 9550 -38675 9585
rect -38665 9550 -38630 9585
rect -38620 9550 -38585 9585
rect -38575 9550 -38540 9585
rect -38530 9550 -38495 9585
rect -38485 9550 -38450 9585
rect -38440 9550 -38405 9585
rect -38395 9550 -38360 9585
rect -38350 9550 -38315 9585
rect -38305 9550 -38270 9585
rect -38260 9550 -38225 9585
rect -38215 9550 -38180 9585
rect -38170 9550 -38135 9585
rect -38125 9550 -38090 9585
rect -38080 9550 -38045 9585
rect -38035 9550 -38000 9585
rect -37990 9550 -37955 9585
rect -37945 9550 -37910 9585
rect -37900 9550 -37865 9585
rect -37855 9550 -37820 9585
rect -37810 9550 -37775 9585
rect -37765 9550 -37730 9585
rect -37720 9550 -37685 9585
rect -37675 9550 -37640 9585
rect -37630 9550 -37595 9585
rect -37585 9550 -37550 9585
rect -37540 9550 -37505 9585
rect -37495 9550 -37460 9585
rect -37450 9550 -37415 9585
rect -37405 9550 -37370 9585
rect -37360 9550 -37325 9585
rect -37315 9550 -37280 9585
rect -37270 9550 -37235 9585
rect -37225 9550 -37190 9585
rect -38755 9505 -38720 9540
rect -38710 9505 -38675 9540
rect -38665 9505 -38630 9540
rect -38620 9505 -38585 9540
rect -38575 9505 -38540 9540
rect -38530 9505 -38495 9540
rect -38485 9505 -38450 9540
rect -38440 9505 -38405 9540
rect -38395 9505 -38360 9540
rect -38350 9505 -38315 9540
rect -38305 9505 -38270 9540
rect -38260 9505 -38225 9540
rect -38215 9505 -38180 9540
rect -38170 9505 -38135 9540
rect -38125 9505 -38090 9540
rect -38080 9505 -38045 9540
rect -38035 9505 -38000 9540
rect -37990 9505 -37955 9540
rect -37945 9505 -37910 9540
rect -37900 9505 -37865 9540
rect -37855 9505 -37820 9540
rect -37810 9505 -37775 9540
rect -37765 9505 -37730 9540
rect -37720 9505 -37685 9540
rect -37675 9505 -37640 9540
rect -37630 9505 -37595 9540
rect -37585 9505 -37550 9540
rect -37540 9505 -37505 9540
rect -37495 9505 -37460 9540
rect -37450 9505 -37415 9540
rect -37405 9505 -37370 9540
rect -37360 9505 -37325 9540
rect -37315 9505 -37280 9540
rect -37270 9505 -37235 9540
rect -37225 9505 -37190 9540
rect -38755 9460 -38720 9495
rect -38710 9460 -38675 9495
rect -38665 9460 -38630 9495
rect -38620 9460 -38585 9495
rect -38575 9460 -38540 9495
rect -38530 9460 -38495 9495
rect -38485 9460 -38450 9495
rect -38440 9460 -38405 9495
rect -38395 9460 -38360 9495
rect -38350 9460 -38315 9495
rect -38305 9460 -38270 9495
rect -38260 9460 -38225 9495
rect -38215 9460 -38180 9495
rect -38170 9460 -38135 9495
rect -38125 9460 -38090 9495
rect -38080 9460 -38045 9495
rect -38035 9460 -38000 9495
rect -37990 9460 -37955 9495
rect -37945 9460 -37910 9495
rect -37900 9460 -37865 9495
rect -37855 9460 -37820 9495
rect -37810 9460 -37775 9495
rect -37765 9460 -37730 9495
rect -37720 9460 -37685 9495
rect -37675 9460 -37640 9495
rect -37630 9460 -37595 9495
rect -37585 9460 -37550 9495
rect -37540 9460 -37505 9495
rect -37495 9460 -37460 9495
rect -37450 9460 -37415 9495
rect -37405 9460 -37370 9495
rect -37360 9460 -37325 9495
rect -37315 9460 -37280 9495
rect -37270 9460 -37235 9495
rect -37225 9460 -37190 9495
rect -38755 9415 -38720 9450
rect -38710 9415 -38675 9450
rect -38665 9415 -38630 9450
rect -38620 9415 -38585 9450
rect -38575 9415 -38540 9450
rect -38530 9415 -38495 9450
rect -38485 9415 -38450 9450
rect -38440 9415 -38405 9450
rect -38395 9415 -38360 9450
rect -38350 9415 -38315 9450
rect -38305 9415 -38270 9450
rect -38260 9415 -38225 9450
rect -38215 9415 -38180 9450
rect -38170 9415 -38135 9450
rect -38125 9415 -38090 9450
rect -38080 9415 -38045 9450
rect -38035 9415 -38000 9450
rect -37990 9415 -37955 9450
rect -37945 9415 -37910 9450
rect -37900 9415 -37865 9450
rect -37855 9415 -37820 9450
rect -37810 9415 -37775 9450
rect -37765 9415 -37730 9450
rect -37720 9415 -37685 9450
rect -37675 9415 -37640 9450
rect -37630 9415 -37595 9450
rect -37585 9415 -37550 9450
rect -37540 9415 -37505 9450
rect -37495 9415 -37460 9450
rect -37450 9415 -37415 9450
rect -37405 9415 -37370 9450
rect -37360 9415 -37325 9450
rect -37315 9415 -37280 9450
rect -37270 9415 -37235 9450
rect -37225 9415 -37190 9450
rect -38755 9370 -38720 9405
rect -38710 9370 -38675 9405
rect -38665 9370 -38630 9405
rect -38620 9370 -38585 9405
rect -38575 9370 -38540 9405
rect -38530 9370 -38495 9405
rect -38485 9370 -38450 9405
rect -38440 9370 -38405 9405
rect -38395 9370 -38360 9405
rect -38350 9370 -38315 9405
rect -38305 9370 -38270 9405
rect -38260 9370 -38225 9405
rect -38215 9370 -38180 9405
rect -38170 9370 -38135 9405
rect -38125 9370 -38090 9405
rect -38080 9370 -38045 9405
rect -38035 9370 -38000 9405
rect -37990 9370 -37955 9405
rect -37945 9370 -37910 9405
rect -37900 9370 -37865 9405
rect -37855 9370 -37820 9405
rect -37810 9370 -37775 9405
rect -37765 9370 -37730 9405
rect -37720 9370 -37685 9405
rect -37675 9370 -37640 9405
rect -37630 9370 -37595 9405
rect -37585 9370 -37550 9405
rect -37540 9370 -37505 9405
rect -37495 9370 -37460 9405
rect -37450 9370 -37415 9405
rect -37405 9370 -37370 9405
rect -37360 9370 -37325 9405
rect -37315 9370 -37280 9405
rect -37270 9370 -37235 9405
rect -37225 9370 -37190 9405
rect -38755 9325 -38720 9360
rect -38710 9325 -38675 9360
rect -38665 9325 -38630 9360
rect -38620 9325 -38585 9360
rect -38575 9325 -38540 9360
rect -38530 9325 -38495 9360
rect -38485 9325 -38450 9360
rect -38440 9325 -38405 9360
rect -38395 9325 -38360 9360
rect -38350 9325 -38315 9360
rect -38305 9325 -38270 9360
rect -38260 9325 -38225 9360
rect -38215 9325 -38180 9360
rect -38170 9325 -38135 9360
rect -38125 9325 -38090 9360
rect -38080 9325 -38045 9360
rect -38035 9325 -38000 9360
rect -37990 9325 -37955 9360
rect -37945 9325 -37910 9360
rect -37900 9325 -37865 9360
rect -37855 9325 -37820 9360
rect -37810 9325 -37775 9360
rect -37765 9325 -37730 9360
rect -37720 9325 -37685 9360
rect -37675 9325 -37640 9360
rect -37630 9325 -37595 9360
rect -37585 9325 -37550 9360
rect -37540 9325 -37505 9360
rect -37495 9325 -37460 9360
rect -37450 9325 -37415 9360
rect -37405 9325 -37370 9360
rect -37360 9325 -37325 9360
rect -37315 9325 -37280 9360
rect -37270 9325 -37235 9360
rect -37225 9325 -37190 9360
rect -38755 9280 -38720 9315
rect -38710 9280 -38675 9315
rect -38665 9280 -38630 9315
rect -38620 9280 -38585 9315
rect -38575 9280 -38540 9315
rect -38530 9280 -38495 9315
rect -38485 9280 -38450 9315
rect -38440 9280 -38405 9315
rect -38395 9280 -38360 9315
rect -38350 9280 -38315 9315
rect -38305 9280 -38270 9315
rect -38260 9280 -38225 9315
rect -38215 9280 -38180 9315
rect -38170 9280 -38135 9315
rect -38125 9280 -38090 9315
rect -38080 9280 -38045 9315
rect -38035 9280 -38000 9315
rect -37990 9280 -37955 9315
rect -37945 9280 -37910 9315
rect -37900 9280 -37865 9315
rect -37855 9280 -37820 9315
rect -37810 9280 -37775 9315
rect -37765 9280 -37730 9315
rect -37720 9280 -37685 9315
rect -37675 9280 -37640 9315
rect -37630 9280 -37595 9315
rect -37585 9280 -37550 9315
rect -37540 9280 -37505 9315
rect -37495 9280 -37460 9315
rect -37450 9280 -37415 9315
rect -37405 9280 -37370 9315
rect -37360 9280 -37325 9315
rect -37315 9280 -37280 9315
rect -37270 9280 -37235 9315
rect -37225 9280 -37190 9315
rect -38755 9235 -38720 9270
rect -38710 9235 -38675 9270
rect -38665 9235 -38630 9270
rect -38620 9235 -38585 9270
rect -38575 9235 -38540 9270
rect -38530 9235 -38495 9270
rect -38485 9235 -38450 9270
rect -38440 9235 -38405 9270
rect -38395 9235 -38360 9270
rect -38350 9235 -38315 9270
rect -38305 9235 -38270 9270
rect -38260 9235 -38225 9270
rect -38215 9235 -38180 9270
rect -38170 9235 -38135 9270
rect -38125 9235 -38090 9270
rect -38080 9235 -38045 9270
rect -38035 9235 -38000 9270
rect -37990 9235 -37955 9270
rect -37945 9235 -37910 9270
rect -37900 9235 -37865 9270
rect -37855 9235 -37820 9270
rect -37810 9235 -37775 9270
rect -37765 9235 -37730 9270
rect -37720 9235 -37685 9270
rect -37675 9235 -37640 9270
rect -37630 9235 -37595 9270
rect -37585 9235 -37550 9270
rect -37540 9235 -37505 9270
rect -37495 9235 -37460 9270
rect -37450 9235 -37415 9270
rect -37405 9235 -37370 9270
rect -37360 9235 -37325 9270
rect -37315 9235 -37280 9270
rect -37270 9235 -37235 9270
rect -37225 9235 -37190 9270
rect -38755 9190 -38720 9225
rect -38710 9190 -38675 9225
rect -38665 9190 -38630 9225
rect -38620 9190 -38585 9225
rect -38575 9190 -38540 9225
rect -38530 9190 -38495 9225
rect -38485 9190 -38450 9225
rect -38440 9190 -38405 9225
rect -38395 9190 -38360 9225
rect -38350 9190 -38315 9225
rect -38305 9190 -38270 9225
rect -38260 9190 -38225 9225
rect -38215 9190 -38180 9225
rect -38170 9190 -38135 9225
rect -38125 9190 -38090 9225
rect -38080 9190 -38045 9225
rect -38035 9190 -38000 9225
rect -37990 9190 -37955 9225
rect -37945 9190 -37910 9225
rect -37900 9190 -37865 9225
rect -37855 9190 -37820 9225
rect -37810 9190 -37775 9225
rect -37765 9190 -37730 9225
rect -37720 9190 -37685 9225
rect -37675 9190 -37640 9225
rect -37630 9190 -37595 9225
rect -37585 9190 -37550 9225
rect -37540 9190 -37505 9225
rect -37495 9190 -37460 9225
rect -37450 9190 -37415 9225
rect -37405 9190 -37370 9225
rect -37360 9190 -37325 9225
rect -37315 9190 -37280 9225
rect -37270 9190 -37235 9225
rect -37225 9190 -37190 9225
rect -38755 9145 -38720 9180
rect -38710 9145 -38675 9180
rect -38665 9145 -38630 9180
rect -38620 9145 -38585 9180
rect -38575 9145 -38540 9180
rect -38530 9145 -38495 9180
rect -38485 9145 -38450 9180
rect -38440 9145 -38405 9180
rect -38395 9145 -38360 9180
rect -38350 9145 -38315 9180
rect -38305 9145 -38270 9180
rect -38260 9145 -38225 9180
rect -38215 9145 -38180 9180
rect -38170 9145 -38135 9180
rect -38125 9145 -38090 9180
rect -38080 9145 -38045 9180
rect -38035 9145 -38000 9180
rect -37990 9145 -37955 9180
rect -37945 9145 -37910 9180
rect -37900 9145 -37865 9180
rect -37855 9145 -37820 9180
rect -37810 9145 -37775 9180
rect -37765 9145 -37730 9180
rect -37720 9145 -37685 9180
rect -37675 9145 -37640 9180
rect -37630 9145 -37595 9180
rect -37585 9145 -37550 9180
rect -37540 9145 -37505 9180
rect -37495 9145 -37460 9180
rect -37450 9145 -37415 9180
rect -37405 9145 -37370 9180
rect -37360 9145 -37325 9180
rect -37315 9145 -37280 9180
rect -37270 9145 -37235 9180
rect -37225 9145 -37190 9180
rect -38755 9100 -38720 9135
rect -38710 9100 -38675 9135
rect -38665 9100 -38630 9135
rect -38620 9100 -38585 9135
rect -38575 9100 -38540 9135
rect -38530 9100 -38495 9135
rect -38485 9100 -38450 9135
rect -38440 9100 -38405 9135
rect -38395 9100 -38360 9135
rect -38350 9100 -38315 9135
rect -38305 9100 -38270 9135
rect -38260 9100 -38225 9135
rect -38215 9100 -38180 9135
rect -38170 9100 -38135 9135
rect -38125 9100 -38090 9135
rect -38080 9100 -38045 9135
rect -38035 9100 -38000 9135
rect -37990 9100 -37955 9135
rect -37945 9100 -37910 9135
rect -37900 9100 -37865 9135
rect -37855 9100 -37820 9135
rect -37810 9100 -37775 9135
rect -37765 9100 -37730 9135
rect -37720 9100 -37685 9135
rect -37675 9100 -37640 9135
rect -37630 9100 -37595 9135
rect -37585 9100 -37550 9135
rect -37540 9100 -37505 9135
rect -37495 9100 -37460 9135
rect -37450 9100 -37415 9135
rect -37405 9100 -37370 9135
rect -37360 9100 -37325 9135
rect -37315 9100 -37280 9135
rect -37270 9100 -37235 9135
rect -37225 9100 -37190 9135
rect -38755 9055 -38720 9090
rect -38710 9055 -38675 9090
rect -38665 9055 -38630 9090
rect -38620 9055 -38585 9090
rect -38575 9055 -38540 9090
rect -38530 9055 -38495 9090
rect -38485 9055 -38450 9090
rect -38440 9055 -38405 9090
rect -38395 9055 -38360 9090
rect -38350 9055 -38315 9090
rect -38305 9055 -38270 9090
rect -38260 9055 -38225 9090
rect -38215 9055 -38180 9090
rect -38170 9055 -38135 9090
rect -38125 9055 -38090 9090
rect -38080 9055 -38045 9090
rect -38035 9055 -38000 9090
rect -37990 9055 -37955 9090
rect -37945 9055 -37910 9090
rect -37900 9055 -37865 9090
rect -37855 9055 -37820 9090
rect -37810 9055 -37775 9090
rect -37765 9055 -37730 9090
rect -37720 9055 -37685 9090
rect -37675 9055 -37640 9090
rect -37630 9055 -37595 9090
rect -37585 9055 -37550 9090
rect -37540 9055 -37505 9090
rect -37495 9055 -37460 9090
rect -37450 9055 -37415 9090
rect -37405 9055 -37370 9090
rect -37360 9055 -37325 9090
rect -37315 9055 -37280 9090
rect -37270 9055 -37235 9090
rect -37225 9055 -37190 9090
rect -38755 9010 -38720 9045
rect -38710 9010 -38675 9045
rect -38665 9010 -38630 9045
rect -38620 9010 -38585 9045
rect -38575 9010 -38540 9045
rect -38530 9010 -38495 9045
rect -38485 9010 -38450 9045
rect -38440 9010 -38405 9045
rect -38395 9010 -38360 9045
rect -38350 9010 -38315 9045
rect -38305 9010 -38270 9045
rect -38260 9010 -38225 9045
rect -38215 9010 -38180 9045
rect -38170 9010 -38135 9045
rect -38125 9010 -38090 9045
rect -38080 9010 -38045 9045
rect -38035 9010 -38000 9045
rect -37990 9010 -37955 9045
rect -37945 9010 -37910 9045
rect -37900 9010 -37865 9045
rect -37855 9010 -37820 9045
rect -37810 9010 -37775 9045
rect -37765 9010 -37730 9045
rect -37720 9010 -37685 9045
rect -37675 9010 -37640 9045
rect -37630 9010 -37595 9045
rect -37585 9010 -37550 9045
rect -37540 9010 -37505 9045
rect -37495 9010 -37460 9045
rect -37450 9010 -37415 9045
rect -37405 9010 -37370 9045
rect -37360 9010 -37325 9045
rect -37315 9010 -37280 9045
rect -37270 9010 -37235 9045
rect -37225 9010 -37190 9045
rect -38755 8965 -38720 9000
rect -38710 8965 -38675 9000
rect -38665 8965 -38630 9000
rect -38620 8965 -38585 9000
rect -38575 8965 -38540 9000
rect -38530 8965 -38495 9000
rect -38485 8965 -38450 9000
rect -38440 8965 -38405 9000
rect -38395 8965 -38360 9000
rect -38350 8965 -38315 9000
rect -38305 8965 -38270 9000
rect -38260 8965 -38225 9000
rect -38215 8965 -38180 9000
rect -38170 8965 -38135 9000
rect -38125 8965 -38090 9000
rect -38080 8965 -38045 9000
rect -38035 8965 -38000 9000
rect -37990 8965 -37955 9000
rect -37945 8965 -37910 9000
rect -37900 8965 -37865 9000
rect -37855 8965 -37820 9000
rect -37810 8965 -37775 9000
rect -37765 8965 -37730 9000
rect -37720 8965 -37685 9000
rect -37675 8965 -37640 9000
rect -37630 8965 -37595 9000
rect -37585 8965 -37550 9000
rect -37540 8965 -37505 9000
rect -37495 8965 -37460 9000
rect -37450 8965 -37415 9000
rect -37405 8965 -37370 9000
rect -37360 8965 -37325 9000
rect -37315 8965 -37280 9000
rect -37270 8965 -37235 9000
rect -37225 8965 -37190 9000
rect -38755 8920 -38720 8955
rect -38710 8920 -38675 8955
rect -38665 8920 -38630 8955
rect -38620 8920 -38585 8955
rect -38575 8920 -38540 8955
rect -38530 8920 -38495 8955
rect -38485 8920 -38450 8955
rect -38440 8920 -38405 8955
rect -38395 8920 -38360 8955
rect -38350 8920 -38315 8955
rect -38305 8920 -38270 8955
rect -38260 8920 -38225 8955
rect -38215 8920 -38180 8955
rect -38170 8920 -38135 8955
rect -38125 8920 -38090 8955
rect -38080 8920 -38045 8955
rect -38035 8920 -38000 8955
rect -37990 8920 -37955 8955
rect -37945 8920 -37910 8955
rect -37900 8920 -37865 8955
rect -37855 8920 -37820 8955
rect -37810 8920 -37775 8955
rect -37765 8920 -37730 8955
rect -37720 8920 -37685 8955
rect -37675 8920 -37640 8955
rect -37630 8920 -37595 8955
rect -37585 8920 -37550 8955
rect -37540 8920 -37505 8955
rect -37495 8920 -37460 8955
rect -37450 8920 -37415 8955
rect -37405 8920 -37370 8955
rect -37360 8920 -37325 8955
rect -37315 8920 -37280 8955
rect -37270 8920 -37235 8955
rect -37225 8920 -37190 8955
rect -38755 8875 -38720 8910
rect -38710 8875 -38675 8910
rect -38665 8875 -38630 8910
rect -38620 8875 -38585 8910
rect -38575 8875 -38540 8910
rect -38530 8875 -38495 8910
rect -38485 8875 -38450 8910
rect -38440 8875 -38405 8910
rect -38395 8875 -38360 8910
rect -38350 8875 -38315 8910
rect -38305 8875 -38270 8910
rect -38260 8875 -38225 8910
rect -38215 8875 -38180 8910
rect -38170 8875 -38135 8910
rect -38125 8875 -38090 8910
rect -38080 8875 -38045 8910
rect -38035 8875 -38000 8910
rect -37990 8875 -37955 8910
rect -37945 8875 -37910 8910
rect -37900 8875 -37865 8910
rect -37855 8875 -37820 8910
rect -37810 8875 -37775 8910
rect -37765 8875 -37730 8910
rect -37720 8875 -37685 8910
rect -37675 8875 -37640 8910
rect -37630 8875 -37595 8910
rect -37585 8875 -37550 8910
rect -37540 8875 -37505 8910
rect -37495 8875 -37460 8910
rect -37450 8875 -37415 8910
rect -37405 8875 -37370 8910
rect -37360 8875 -37325 8910
rect -37315 8875 -37280 8910
rect -37270 8875 -37235 8910
rect -37225 8875 -37190 8910
rect -38755 8830 -38720 8865
rect -38710 8830 -38675 8865
rect -38665 8830 -38630 8865
rect -38620 8830 -38585 8865
rect -38575 8830 -38540 8865
rect -38530 8830 -38495 8865
rect -38485 8830 -38450 8865
rect -38440 8830 -38405 8865
rect -38395 8830 -38360 8865
rect -38350 8830 -38315 8865
rect -38305 8830 -38270 8865
rect -38260 8830 -38225 8865
rect -38215 8830 -38180 8865
rect -38170 8830 -38135 8865
rect -38125 8830 -38090 8865
rect -38080 8830 -38045 8865
rect -38035 8830 -38000 8865
rect -37990 8830 -37955 8865
rect -37945 8830 -37910 8865
rect -37900 8830 -37865 8865
rect -37855 8830 -37820 8865
rect -37810 8830 -37775 8865
rect -37765 8830 -37730 8865
rect -37720 8830 -37685 8865
rect -37675 8830 -37640 8865
rect -37630 8830 -37595 8865
rect -37585 8830 -37550 8865
rect -37540 8830 -37505 8865
rect -37495 8830 -37460 8865
rect -37450 8830 -37415 8865
rect -37405 8830 -37370 8865
rect -37360 8830 -37325 8865
rect -37315 8830 -37280 8865
rect -37270 8830 -37235 8865
rect -37225 8830 -37190 8865
rect -38755 8785 -38720 8820
rect -38710 8785 -38675 8820
rect -38665 8785 -38630 8820
rect -38620 8785 -38585 8820
rect -38575 8785 -38540 8820
rect -38530 8785 -38495 8820
rect -38485 8785 -38450 8820
rect -38440 8785 -38405 8820
rect -38395 8785 -38360 8820
rect -38350 8785 -38315 8820
rect -38305 8785 -38270 8820
rect -38260 8785 -38225 8820
rect -38215 8785 -38180 8820
rect -38170 8785 -38135 8820
rect -38125 8785 -38090 8820
rect -38080 8785 -38045 8820
rect -38035 8785 -38000 8820
rect -37990 8785 -37955 8820
rect -37945 8785 -37910 8820
rect -37900 8785 -37865 8820
rect -37855 8785 -37820 8820
rect -37810 8785 -37775 8820
rect -37765 8785 -37730 8820
rect -37720 8785 -37685 8820
rect -37675 8785 -37640 8820
rect -37630 8785 -37595 8820
rect -37585 8785 -37550 8820
rect -37540 8785 -37505 8820
rect -37495 8785 -37460 8820
rect -37450 8785 -37415 8820
rect -37405 8785 -37370 8820
rect -37360 8785 -37325 8820
rect -37315 8785 -37280 8820
rect -37270 8785 -37235 8820
rect -37225 8785 -37190 8820
rect -38755 8740 -38720 8775
rect -38710 8740 -38675 8775
rect -38665 8740 -38630 8775
rect -38620 8740 -38585 8775
rect -38575 8740 -38540 8775
rect -38530 8740 -38495 8775
rect -38485 8740 -38450 8775
rect -38440 8740 -38405 8775
rect -38395 8740 -38360 8775
rect -38350 8740 -38315 8775
rect -38305 8740 -38270 8775
rect -38260 8740 -38225 8775
rect -38215 8740 -38180 8775
rect -38170 8740 -38135 8775
rect -38125 8740 -38090 8775
rect -38080 8740 -38045 8775
rect -38035 8740 -38000 8775
rect -37990 8740 -37955 8775
rect -37945 8740 -37910 8775
rect -37900 8740 -37865 8775
rect -37855 8740 -37820 8775
rect -37810 8740 -37775 8775
rect -37765 8740 -37730 8775
rect -37720 8740 -37685 8775
rect -37675 8740 -37640 8775
rect -37630 8740 -37595 8775
rect -37585 8740 -37550 8775
rect -37540 8740 -37505 8775
rect -37495 8740 -37460 8775
rect -37450 8740 -37415 8775
rect -37405 8740 -37370 8775
rect -37360 8740 -37325 8775
rect -37315 8740 -37280 8775
rect -37270 8740 -37235 8775
rect -37225 8740 -37190 8775
rect -38755 8695 -38720 8730
rect -38710 8695 -38675 8730
rect -38665 8695 -38630 8730
rect -38620 8695 -38585 8730
rect -38575 8695 -38540 8730
rect -38530 8695 -38495 8730
rect -38485 8695 -38450 8730
rect -38440 8695 -38405 8730
rect -38395 8695 -38360 8730
rect -38350 8695 -38315 8730
rect -38305 8695 -38270 8730
rect -38260 8695 -38225 8730
rect -38215 8695 -38180 8730
rect -38170 8695 -38135 8730
rect -38125 8695 -38090 8730
rect -38080 8695 -38045 8730
rect -38035 8695 -38000 8730
rect -37990 8695 -37955 8730
rect -37945 8695 -37910 8730
rect -37900 8695 -37865 8730
rect -37855 8695 -37820 8730
rect -37810 8695 -37775 8730
rect -37765 8695 -37730 8730
rect -37720 8695 -37685 8730
rect -37675 8695 -37640 8730
rect -37630 8695 -37595 8730
rect -37585 8695 -37550 8730
rect -37540 8695 -37505 8730
rect -37495 8695 -37460 8730
rect -37450 8695 -37415 8730
rect -37405 8695 -37370 8730
rect -37360 8695 -37325 8730
rect -37315 8695 -37280 8730
rect -37270 8695 -37235 8730
rect -37225 8695 -37190 8730
rect -38755 8650 -38720 8685
rect -38710 8650 -38675 8685
rect -38665 8650 -38630 8685
rect -38620 8650 -38585 8685
rect -38575 8650 -38540 8685
rect -38530 8650 -38495 8685
rect -38485 8650 -38450 8685
rect -38440 8650 -38405 8685
rect -38395 8650 -38360 8685
rect -38350 8650 -38315 8685
rect -38305 8650 -38270 8685
rect -38260 8650 -38225 8685
rect -38215 8650 -38180 8685
rect -38170 8650 -38135 8685
rect -38125 8650 -38090 8685
rect -38080 8650 -38045 8685
rect -38035 8650 -38000 8685
rect -37990 8650 -37955 8685
rect -37945 8650 -37910 8685
rect -37900 8650 -37865 8685
rect -37855 8650 -37820 8685
rect -37810 8650 -37775 8685
rect -37765 8650 -37730 8685
rect -37720 8650 -37685 8685
rect -37675 8650 -37640 8685
rect -37630 8650 -37595 8685
rect -37585 8650 -37550 8685
rect -37540 8650 -37505 8685
rect -37495 8650 -37460 8685
rect -37450 8650 -37415 8685
rect -37405 8650 -37370 8685
rect -37360 8650 -37325 8685
rect -37315 8650 -37280 8685
rect -37270 8650 -37235 8685
rect -37225 8650 -37190 8685
rect -38755 8605 -38720 8640
rect -38710 8605 -38675 8640
rect -38665 8605 -38630 8640
rect -38620 8605 -38585 8640
rect -38575 8605 -38540 8640
rect -38530 8605 -38495 8640
rect -38485 8605 -38450 8640
rect -38440 8605 -38405 8640
rect -38395 8605 -38360 8640
rect -38350 8605 -38315 8640
rect -38305 8605 -38270 8640
rect -38260 8605 -38225 8640
rect -38215 8605 -38180 8640
rect -38170 8605 -38135 8640
rect -38125 8605 -38090 8640
rect -38080 8605 -38045 8640
rect -38035 8605 -38000 8640
rect -37990 8605 -37955 8640
rect -37945 8605 -37910 8640
rect -37900 8605 -37865 8640
rect -37855 8605 -37820 8640
rect -37810 8605 -37775 8640
rect -37765 8605 -37730 8640
rect -37720 8605 -37685 8640
rect -37675 8605 -37640 8640
rect -37630 8605 -37595 8640
rect -37585 8605 -37550 8640
rect -37540 8605 -37505 8640
rect -37495 8605 -37460 8640
rect -37450 8605 -37415 8640
rect -37405 8605 -37370 8640
rect -37360 8605 -37325 8640
rect -37315 8605 -37280 8640
rect -37270 8605 -37235 8640
rect -37225 8605 -37190 8640
rect -38755 8560 -38720 8595
rect -38710 8560 -38675 8595
rect -38665 8560 -38630 8595
rect -38620 8560 -38585 8595
rect -38575 8560 -38540 8595
rect -38530 8560 -38495 8595
rect -38485 8560 -38450 8595
rect -38440 8560 -38405 8595
rect -38395 8560 -38360 8595
rect -38350 8560 -38315 8595
rect -38305 8560 -38270 8595
rect -38260 8560 -38225 8595
rect -38215 8560 -38180 8595
rect -38170 8560 -38135 8595
rect -38125 8560 -38090 8595
rect -38080 8560 -38045 8595
rect -38035 8560 -38000 8595
rect -37990 8560 -37955 8595
rect -37945 8560 -37910 8595
rect -37900 8560 -37865 8595
rect -37855 8560 -37820 8595
rect -37810 8560 -37775 8595
rect -37765 8560 -37730 8595
rect -37720 8560 -37685 8595
rect -37675 8560 -37640 8595
rect -37630 8560 -37595 8595
rect -37585 8560 -37550 8595
rect -37540 8560 -37505 8595
rect -37495 8560 -37460 8595
rect -37450 8560 -37415 8595
rect -37405 8560 -37370 8595
rect -37360 8560 -37325 8595
rect -37315 8560 -37280 8595
rect -37270 8560 -37235 8595
rect -37225 8560 -37190 8595
rect -38755 8515 -38720 8550
rect -38710 8515 -38675 8550
rect -38665 8515 -38630 8550
rect -38620 8515 -38585 8550
rect -38575 8515 -38540 8550
rect -38530 8515 -38495 8550
rect -38485 8515 -38450 8550
rect -38440 8515 -38405 8550
rect -38395 8515 -38360 8550
rect -38350 8515 -38315 8550
rect -38305 8515 -38270 8550
rect -38260 8515 -38225 8550
rect -38215 8515 -38180 8550
rect -38170 8515 -38135 8550
rect -38125 8515 -38090 8550
rect -38080 8515 -38045 8550
rect -38035 8515 -38000 8550
rect -37990 8515 -37955 8550
rect -37945 8515 -37910 8550
rect -37900 8515 -37865 8550
rect -37855 8515 -37820 8550
rect -37810 8515 -37775 8550
rect -37765 8515 -37730 8550
rect -37720 8515 -37685 8550
rect -37675 8515 -37640 8550
rect -37630 8515 -37595 8550
rect -37585 8515 -37550 8550
rect -37540 8515 -37505 8550
rect -37495 8515 -37460 8550
rect -37450 8515 -37415 8550
rect -37405 8515 -37370 8550
rect -37360 8515 -37325 8550
rect -37315 8515 -37280 8550
rect -37270 8515 -37235 8550
rect -37225 8515 -37190 8550
rect -38755 8470 -38720 8505
rect -38710 8470 -38675 8505
rect -38665 8470 -38630 8505
rect -38620 8470 -38585 8505
rect -38575 8470 -38540 8505
rect -38530 8470 -38495 8505
rect -38485 8470 -38450 8505
rect -38440 8470 -38405 8505
rect -38395 8470 -38360 8505
rect -38350 8470 -38315 8505
rect -38305 8470 -38270 8505
rect -38260 8470 -38225 8505
rect -38215 8470 -38180 8505
rect -38170 8470 -38135 8505
rect -38125 8470 -38090 8505
rect -38080 8470 -38045 8505
rect -38035 8470 -38000 8505
rect -37990 8470 -37955 8505
rect -37945 8470 -37910 8505
rect -37900 8470 -37865 8505
rect -37855 8470 -37820 8505
rect -37810 8470 -37775 8505
rect -37765 8470 -37730 8505
rect -37720 8470 -37685 8505
rect -37675 8470 -37640 8505
rect -37630 8470 -37595 8505
rect -37585 8470 -37550 8505
rect -37540 8470 -37505 8505
rect -37495 8470 -37460 8505
rect -37450 8470 -37415 8505
rect -37405 8470 -37370 8505
rect -37360 8470 -37325 8505
rect -37315 8470 -37280 8505
rect -37270 8470 -37235 8505
rect -37225 8470 -37190 8505
rect -38755 8425 -38720 8460
rect -38710 8425 -38675 8460
rect -38665 8425 -38630 8460
rect -38620 8425 -38585 8460
rect -38575 8425 -38540 8460
rect -38530 8425 -38495 8460
rect -38485 8425 -38450 8460
rect -38440 8425 -38405 8460
rect -38395 8425 -38360 8460
rect -38350 8425 -38315 8460
rect -38305 8425 -38270 8460
rect -38260 8425 -38225 8460
rect -38215 8425 -38180 8460
rect -38170 8425 -38135 8460
rect -38125 8425 -38090 8460
rect -38080 8425 -38045 8460
rect -38035 8425 -38000 8460
rect -37990 8425 -37955 8460
rect -37945 8425 -37910 8460
rect -37900 8425 -37865 8460
rect -37855 8425 -37820 8460
rect -37810 8425 -37775 8460
rect -37765 8425 -37730 8460
rect -37720 8425 -37685 8460
rect -37675 8425 -37640 8460
rect -37630 8425 -37595 8460
rect -37585 8425 -37550 8460
rect -37540 8425 -37505 8460
rect -37495 8425 -37460 8460
rect -37450 8425 -37415 8460
rect -37405 8425 -37370 8460
rect -37360 8425 -37325 8460
rect -37315 8425 -37280 8460
rect -37270 8425 -37235 8460
rect -37225 8425 -37190 8460
rect -38755 8380 -38720 8415
rect -38710 8380 -38675 8415
rect -38665 8380 -38630 8415
rect -38620 8380 -38585 8415
rect -38575 8380 -38540 8415
rect -38530 8380 -38495 8415
rect -38485 8380 -38450 8415
rect -38440 8380 -38405 8415
rect -38395 8380 -38360 8415
rect -38350 8380 -38315 8415
rect -38305 8380 -38270 8415
rect -38260 8380 -38225 8415
rect -38215 8380 -38180 8415
rect -38170 8380 -38135 8415
rect -38125 8380 -38090 8415
rect -38080 8380 -38045 8415
rect -38035 8380 -38000 8415
rect -37990 8380 -37955 8415
rect -37945 8380 -37910 8415
rect -37900 8380 -37865 8415
rect -37855 8380 -37820 8415
rect -37810 8380 -37775 8415
rect -37765 8380 -37730 8415
rect -37720 8380 -37685 8415
rect -37675 8380 -37640 8415
rect -37630 8380 -37595 8415
rect -37585 8380 -37550 8415
rect -37540 8380 -37505 8415
rect -37495 8380 -37460 8415
rect -37450 8380 -37415 8415
rect -37405 8380 -37370 8415
rect -37360 8380 -37325 8415
rect -37315 8380 -37280 8415
rect -37270 8380 -37235 8415
rect -37225 8380 -37190 8415
rect -38755 8335 -38720 8370
rect -38710 8335 -38675 8370
rect -38665 8335 -38630 8370
rect -38620 8335 -38585 8370
rect -38575 8335 -38540 8370
rect -38530 8335 -38495 8370
rect -38485 8335 -38450 8370
rect -38440 8335 -38405 8370
rect -38395 8335 -38360 8370
rect -38350 8335 -38315 8370
rect -38305 8335 -38270 8370
rect -38260 8335 -38225 8370
rect -38215 8335 -38180 8370
rect -38170 8335 -38135 8370
rect -38125 8335 -38090 8370
rect -38080 8335 -38045 8370
rect -38035 8335 -38000 8370
rect -37990 8335 -37955 8370
rect -37945 8335 -37910 8370
rect -37900 8335 -37865 8370
rect -37855 8335 -37820 8370
rect -37810 8335 -37775 8370
rect -37765 8335 -37730 8370
rect -37720 8335 -37685 8370
rect -37675 8335 -37640 8370
rect -37630 8335 -37595 8370
rect -37585 8335 -37550 8370
rect -37540 8335 -37505 8370
rect -37495 8335 -37460 8370
rect -37450 8335 -37415 8370
rect -37405 8335 -37370 8370
rect -37360 8335 -37325 8370
rect -37315 8335 -37280 8370
rect -37270 8335 -37235 8370
rect -37225 8335 -37190 8370
rect -38755 8290 -38720 8325
rect -38710 8290 -38675 8325
rect -38665 8290 -38630 8325
rect -38620 8290 -38585 8325
rect -38575 8290 -38540 8325
rect -38530 8290 -38495 8325
rect -38485 8290 -38450 8325
rect -38440 8290 -38405 8325
rect -38395 8290 -38360 8325
rect -38350 8290 -38315 8325
rect -38305 8290 -38270 8325
rect -38260 8290 -38225 8325
rect -38215 8290 -38180 8325
rect -38170 8290 -38135 8325
rect -38125 8290 -38090 8325
rect -38080 8290 -38045 8325
rect -38035 8290 -38000 8325
rect -37990 8290 -37955 8325
rect -37945 8290 -37910 8325
rect -37900 8290 -37865 8325
rect -37855 8290 -37820 8325
rect -37810 8290 -37775 8325
rect -37765 8290 -37730 8325
rect -37720 8290 -37685 8325
rect -37675 8290 -37640 8325
rect -37630 8290 -37595 8325
rect -37585 8290 -37550 8325
rect -37540 8290 -37505 8325
rect -37495 8290 -37460 8325
rect -37450 8290 -37415 8325
rect -37405 8290 -37370 8325
rect -37360 8290 -37325 8325
rect -37315 8290 -37280 8325
rect -37270 8290 -37235 8325
rect -37225 8290 -37190 8325
rect -38755 8245 -38720 8280
rect -38710 8245 -38675 8280
rect -38665 8245 -38630 8280
rect -38620 8245 -38585 8280
rect -38575 8245 -38540 8280
rect -38530 8245 -38495 8280
rect -38485 8245 -38450 8280
rect -38440 8245 -38405 8280
rect -38395 8245 -38360 8280
rect -38350 8245 -38315 8280
rect -38305 8245 -38270 8280
rect -38260 8245 -38225 8280
rect -38215 8245 -38180 8280
rect -38170 8245 -38135 8280
rect -38125 8245 -38090 8280
rect -38080 8245 -38045 8280
rect -38035 8245 -38000 8280
rect -37990 8245 -37955 8280
rect -37945 8245 -37910 8280
rect -37900 8245 -37865 8280
rect -37855 8245 -37820 8280
rect -37810 8245 -37775 8280
rect -37765 8245 -37730 8280
rect -37720 8245 -37685 8280
rect -37675 8245 -37640 8280
rect -37630 8245 -37595 8280
rect -37585 8245 -37550 8280
rect -37540 8245 -37505 8280
rect -37495 8245 -37460 8280
rect -37450 8245 -37415 8280
rect -37405 8245 -37370 8280
rect -37360 8245 -37325 8280
rect -37315 8245 -37280 8280
rect -37270 8245 -37235 8280
rect -37225 8245 -37190 8280
rect -38755 8200 -38720 8235
rect -38710 8200 -38675 8235
rect -38665 8200 -38630 8235
rect -38620 8200 -38585 8235
rect -38575 8200 -38540 8235
rect -38530 8200 -38495 8235
rect -38485 8200 -38450 8235
rect -38440 8200 -38405 8235
rect -38395 8200 -38360 8235
rect -38350 8200 -38315 8235
rect -38305 8200 -38270 8235
rect -38260 8200 -38225 8235
rect -38215 8200 -38180 8235
rect -38170 8200 -38135 8235
rect -38125 8200 -38090 8235
rect -38080 8200 -38045 8235
rect -38035 8200 -38000 8235
rect -37990 8200 -37955 8235
rect -37945 8200 -37910 8235
rect -37900 8200 -37865 8235
rect -37855 8200 -37820 8235
rect -37810 8200 -37775 8235
rect -37765 8200 -37730 8235
rect -37720 8200 -37685 8235
rect -37675 8200 -37640 8235
rect -37630 8200 -37595 8235
rect -37585 8200 -37550 8235
rect -37540 8200 -37505 8235
rect -37495 8200 -37460 8235
rect -37450 8200 -37415 8235
rect -37405 8200 -37370 8235
rect -37360 8200 -37325 8235
rect -37315 8200 -37280 8235
rect -37270 8200 -37235 8235
rect -37225 8200 -37190 8235
rect -38755 8155 -38720 8190
rect -38710 8155 -38675 8190
rect -38665 8155 -38630 8190
rect -38620 8155 -38585 8190
rect -38575 8155 -38540 8190
rect -38530 8155 -38495 8190
rect -38485 8155 -38450 8190
rect -38440 8155 -38405 8190
rect -38395 8155 -38360 8190
rect -38350 8155 -38315 8190
rect -38305 8155 -38270 8190
rect -38260 8155 -38225 8190
rect -38215 8155 -38180 8190
rect -38170 8155 -38135 8190
rect -38125 8155 -38090 8190
rect -38080 8155 -38045 8190
rect -38035 8155 -38000 8190
rect -37990 8155 -37955 8190
rect -37945 8155 -37910 8190
rect -37900 8155 -37865 8190
rect -37855 8155 -37820 8190
rect -37810 8155 -37775 8190
rect -37765 8155 -37730 8190
rect -37720 8155 -37685 8190
rect -37675 8155 -37640 8190
rect -37630 8155 -37595 8190
rect -37585 8155 -37550 8190
rect -37540 8155 -37505 8190
rect -37495 8155 -37460 8190
rect -37450 8155 -37415 8190
rect -37405 8155 -37370 8190
rect -37360 8155 -37325 8190
rect -37315 8155 -37280 8190
rect -37270 8155 -37235 8190
rect -37225 8155 -37190 8190
rect -38755 8110 -38720 8145
rect -38710 8110 -38675 8145
rect -38665 8110 -38630 8145
rect -38620 8110 -38585 8145
rect -38575 8110 -38540 8145
rect -38530 8110 -38495 8145
rect -38485 8110 -38450 8145
rect -38440 8110 -38405 8145
rect -38395 8110 -38360 8145
rect -38350 8110 -38315 8145
rect -38305 8110 -38270 8145
rect -38260 8110 -38225 8145
rect -38215 8110 -38180 8145
rect -38170 8110 -38135 8145
rect -38125 8110 -38090 8145
rect -38080 8110 -38045 8145
rect -38035 8110 -38000 8145
rect -37990 8110 -37955 8145
rect -37945 8110 -37910 8145
rect -37900 8110 -37865 8145
rect -37855 8110 -37820 8145
rect -37810 8110 -37775 8145
rect -37765 8110 -37730 8145
rect -37720 8110 -37685 8145
rect -37675 8110 -37640 8145
rect -37630 8110 -37595 8145
rect -37585 8110 -37550 8145
rect -37540 8110 -37505 8145
rect -37495 8110 -37460 8145
rect -37450 8110 -37415 8145
rect -37405 8110 -37370 8145
rect -37360 8110 -37325 8145
rect -37315 8110 -37280 8145
rect -37270 8110 -37235 8145
rect -37225 8110 -37190 8145
rect -38755 8065 -38720 8100
rect -38710 8065 -38675 8100
rect -38665 8065 -38630 8100
rect -38620 8065 -38585 8100
rect -38575 8065 -38540 8100
rect -38530 8065 -38495 8100
rect -38485 8065 -38450 8100
rect -38440 8065 -38405 8100
rect -38395 8065 -38360 8100
rect -38350 8065 -38315 8100
rect -38305 8065 -38270 8100
rect -38260 8065 -38225 8100
rect -38215 8065 -38180 8100
rect -38170 8065 -38135 8100
rect -38125 8065 -38090 8100
rect -38080 8065 -38045 8100
rect -38035 8065 -38000 8100
rect -37990 8065 -37955 8100
rect -37945 8065 -37910 8100
rect -37900 8065 -37865 8100
rect -37855 8065 -37820 8100
rect -37810 8065 -37775 8100
rect -37765 8065 -37730 8100
rect -37720 8065 -37685 8100
rect -37675 8065 -37640 8100
rect -37630 8065 -37595 8100
rect -37585 8065 -37550 8100
rect -37540 8065 -37505 8100
rect -37495 8065 -37460 8100
rect -37450 8065 -37415 8100
rect -37405 8065 -37370 8100
rect -37360 8065 -37325 8100
rect -37315 8065 -37280 8100
rect -37270 8065 -37235 8100
rect -37225 8065 -37190 8100
rect -38755 7995 -38720 8030
rect -38710 7995 -38675 8030
rect -38665 7995 -38630 8030
rect -38620 7995 -38585 8030
rect -38575 7995 -38540 8030
rect -38530 7995 -38495 8030
rect -38485 7995 -38450 8030
rect -38440 7995 -38405 8030
rect -38395 7995 -38360 8030
rect -38350 7995 -38315 8030
rect -38305 7995 -38270 8030
rect -38260 7995 -38225 8030
rect -38215 7995 -38180 8030
rect -38170 7995 -38135 8030
rect -38125 7995 -38090 8030
rect -38080 7995 -38045 8030
rect -38035 7995 -38000 8030
rect -37990 7995 -37955 8030
rect -37945 7995 -37910 8030
rect -37900 7995 -37865 8030
rect -37855 7995 -37820 8030
rect -37810 7995 -37775 8030
rect -37765 7995 -37730 8030
rect -37720 7995 -37685 8030
rect -37675 7995 -37640 8030
rect -37630 7995 -37595 8030
rect -37585 7995 -37550 8030
rect -37540 7995 -37505 8030
rect -37495 7995 -37460 8030
rect -37450 7995 -37415 8030
rect -37405 7995 -37370 8030
rect -37360 7995 -37325 8030
rect -37315 7995 -37280 8030
rect -37270 7995 -37235 8030
rect -37225 7995 -37190 8030
rect -38755 7950 -38720 7985
rect -38710 7950 -38675 7985
rect -38665 7950 -38630 7985
rect -38620 7950 -38585 7985
rect -38575 7950 -38540 7985
rect -38530 7950 -38495 7985
rect -38485 7950 -38450 7985
rect -38440 7950 -38405 7985
rect -38395 7950 -38360 7985
rect -38350 7950 -38315 7985
rect -38305 7950 -38270 7985
rect -38260 7950 -38225 7985
rect -38215 7950 -38180 7985
rect -38170 7950 -38135 7985
rect -38125 7950 -38090 7985
rect -38080 7950 -38045 7985
rect -38035 7950 -38000 7985
rect -37990 7950 -37955 7985
rect -37945 7950 -37910 7985
rect -37900 7950 -37865 7985
rect -37855 7950 -37820 7985
rect -37810 7950 -37775 7985
rect -37765 7950 -37730 7985
rect -37720 7950 -37685 7985
rect -37675 7950 -37640 7985
rect -37630 7950 -37595 7985
rect -37585 7950 -37550 7985
rect -37540 7950 -37505 7985
rect -37495 7950 -37460 7985
rect -37450 7950 -37415 7985
rect -37405 7950 -37370 7985
rect -37360 7950 -37325 7985
rect -37315 7950 -37280 7985
rect -37270 7950 -37235 7985
rect -37225 7950 -37190 7985
rect -38755 7905 -38720 7940
rect -38710 7905 -38675 7940
rect -38665 7905 -38630 7940
rect -38620 7905 -38585 7940
rect -38575 7905 -38540 7940
rect -38530 7905 -38495 7940
rect -38485 7905 -38450 7940
rect -38440 7905 -38405 7940
rect -38395 7905 -38360 7940
rect -38350 7905 -38315 7940
rect -38305 7905 -38270 7940
rect -38260 7905 -38225 7940
rect -38215 7905 -38180 7940
rect -38170 7905 -38135 7940
rect -38125 7905 -38090 7940
rect -38080 7905 -38045 7940
rect -38035 7905 -38000 7940
rect -37990 7905 -37955 7940
rect -37945 7905 -37910 7940
rect -37900 7905 -37865 7940
rect -37855 7905 -37820 7940
rect -37810 7905 -37775 7940
rect -37765 7905 -37730 7940
rect -37720 7905 -37685 7940
rect -37675 7905 -37640 7940
rect -37630 7905 -37595 7940
rect -37585 7905 -37550 7940
rect -37540 7905 -37505 7940
rect -37495 7905 -37460 7940
rect -37450 7905 -37415 7940
rect -37405 7905 -37370 7940
rect -37360 7905 -37325 7940
rect -37315 7905 -37280 7940
rect -37270 7905 -37235 7940
rect -37225 7905 -37190 7940
rect -38755 7860 -38720 7895
rect -38710 7860 -38675 7895
rect -38665 7860 -38630 7895
rect -38620 7860 -38585 7895
rect -38575 7860 -38540 7895
rect -38530 7860 -38495 7895
rect -38485 7860 -38450 7895
rect -38440 7860 -38405 7895
rect -38395 7860 -38360 7895
rect -38350 7860 -38315 7895
rect -38305 7860 -38270 7895
rect -38260 7860 -38225 7895
rect -38215 7860 -38180 7895
rect -38170 7860 -38135 7895
rect -38125 7860 -38090 7895
rect -38080 7860 -38045 7895
rect -38035 7860 -38000 7895
rect -37990 7860 -37955 7895
rect -37945 7860 -37910 7895
rect -37900 7860 -37865 7895
rect -37855 7860 -37820 7895
rect -37810 7860 -37775 7895
rect -37765 7860 -37730 7895
rect -37720 7860 -37685 7895
rect -37675 7860 -37640 7895
rect -37630 7860 -37595 7895
rect -37585 7860 -37550 7895
rect -37540 7860 -37505 7895
rect -37495 7860 -37460 7895
rect -37450 7860 -37415 7895
rect -37405 7860 -37370 7895
rect -37360 7860 -37325 7895
rect -37315 7860 -37280 7895
rect -37270 7860 -37235 7895
rect -37225 7860 -37190 7895
rect -38755 7815 -38720 7850
rect -38710 7815 -38675 7850
rect -38665 7815 -38630 7850
rect -38620 7815 -38585 7850
rect -38575 7815 -38540 7850
rect -38530 7815 -38495 7850
rect -38485 7815 -38450 7850
rect -38440 7815 -38405 7850
rect -38395 7815 -38360 7850
rect -38350 7815 -38315 7850
rect -38305 7815 -38270 7850
rect -38260 7815 -38225 7850
rect -38215 7815 -38180 7850
rect -38170 7815 -38135 7850
rect -38125 7815 -38090 7850
rect -38080 7815 -38045 7850
rect -38035 7815 -38000 7850
rect -37990 7815 -37955 7850
rect -37945 7815 -37910 7850
rect -37900 7815 -37865 7850
rect -37855 7815 -37820 7850
rect -37810 7815 -37775 7850
rect -37765 7815 -37730 7850
rect -37720 7815 -37685 7850
rect -37675 7815 -37640 7850
rect -37630 7815 -37595 7850
rect -37585 7815 -37550 7850
rect -37540 7815 -37505 7850
rect -37495 7815 -37460 7850
rect -37450 7815 -37415 7850
rect -37405 7815 -37370 7850
rect -37360 7815 -37325 7850
rect -37315 7815 -37280 7850
rect -37270 7815 -37235 7850
rect -37225 7815 -37190 7850
rect -38755 7770 -38720 7805
rect -38710 7770 -38675 7805
rect -38665 7770 -38630 7805
rect -38620 7770 -38585 7805
rect -38575 7770 -38540 7805
rect -38530 7770 -38495 7805
rect -38485 7770 -38450 7805
rect -38440 7770 -38405 7805
rect -38395 7770 -38360 7805
rect -38350 7770 -38315 7805
rect -38305 7770 -38270 7805
rect -38260 7770 -38225 7805
rect -38215 7770 -38180 7805
rect -38170 7770 -38135 7805
rect -38125 7770 -38090 7805
rect -38080 7770 -38045 7805
rect -38035 7770 -38000 7805
rect -37990 7770 -37955 7805
rect -37945 7770 -37910 7805
rect -37900 7770 -37865 7805
rect -37855 7770 -37820 7805
rect -37810 7770 -37775 7805
rect -37765 7770 -37730 7805
rect -37720 7770 -37685 7805
rect -37675 7770 -37640 7805
rect -37630 7770 -37595 7805
rect -37585 7770 -37550 7805
rect -37540 7770 -37505 7805
rect -37495 7770 -37460 7805
rect -37450 7770 -37415 7805
rect -37405 7770 -37370 7805
rect -37360 7770 -37325 7805
rect -37315 7770 -37280 7805
rect -37270 7770 -37235 7805
rect -37225 7770 -37190 7805
rect -38755 7725 -38720 7760
rect -38710 7725 -38675 7760
rect -38665 7725 -38630 7760
rect -38620 7725 -38585 7760
rect -38575 7725 -38540 7760
rect -38530 7725 -38495 7760
rect -38485 7725 -38450 7760
rect -38440 7725 -38405 7760
rect -38395 7725 -38360 7760
rect -38350 7725 -38315 7760
rect -38305 7725 -38270 7760
rect -38260 7725 -38225 7760
rect -38215 7725 -38180 7760
rect -38170 7725 -38135 7760
rect -38125 7725 -38090 7760
rect -38080 7725 -38045 7760
rect -38035 7725 -38000 7760
rect -37990 7725 -37955 7760
rect -37945 7725 -37910 7760
rect -37900 7725 -37865 7760
rect -37855 7725 -37820 7760
rect -37810 7725 -37775 7760
rect -37765 7725 -37730 7760
rect -37720 7725 -37685 7760
rect -37675 7725 -37640 7760
rect -37630 7725 -37595 7760
rect -37585 7725 -37550 7760
rect -37540 7725 -37505 7760
rect -37495 7725 -37460 7760
rect -37450 7725 -37415 7760
rect -37405 7725 -37370 7760
rect -37360 7725 -37325 7760
rect -37315 7725 -37280 7760
rect -37270 7725 -37235 7760
rect -37225 7725 -37190 7760
rect -38755 7680 -38720 7715
rect -38710 7680 -38675 7715
rect -38665 7680 -38630 7715
rect -38620 7680 -38585 7715
rect -38575 7680 -38540 7715
rect -38530 7680 -38495 7715
rect -38485 7680 -38450 7715
rect -38440 7680 -38405 7715
rect -38395 7680 -38360 7715
rect -38350 7680 -38315 7715
rect -38305 7680 -38270 7715
rect -38260 7680 -38225 7715
rect -38215 7680 -38180 7715
rect -38170 7680 -38135 7715
rect -38125 7680 -38090 7715
rect -38080 7680 -38045 7715
rect -38035 7680 -38000 7715
rect -37990 7680 -37955 7715
rect -37945 7680 -37910 7715
rect -37900 7680 -37865 7715
rect -37855 7680 -37820 7715
rect -37810 7680 -37775 7715
rect -37765 7680 -37730 7715
rect -37720 7680 -37685 7715
rect -37675 7680 -37640 7715
rect -37630 7680 -37595 7715
rect -37585 7680 -37550 7715
rect -37540 7680 -37505 7715
rect -37495 7680 -37460 7715
rect -37450 7680 -37415 7715
rect -37405 7680 -37370 7715
rect -37360 7680 -37325 7715
rect -37315 7680 -37280 7715
rect -37270 7680 -37235 7715
rect -37225 7680 -37190 7715
rect -38755 7635 -38720 7670
rect -38710 7635 -38675 7670
rect -38665 7635 -38630 7670
rect -38620 7635 -38585 7670
rect -38575 7635 -38540 7670
rect -38530 7635 -38495 7670
rect -38485 7635 -38450 7670
rect -38440 7635 -38405 7670
rect -38395 7635 -38360 7670
rect -38350 7635 -38315 7670
rect -38305 7635 -38270 7670
rect -38260 7635 -38225 7670
rect -38215 7635 -38180 7670
rect -38170 7635 -38135 7670
rect -38125 7635 -38090 7670
rect -38080 7635 -38045 7670
rect -38035 7635 -38000 7670
rect -37990 7635 -37955 7670
rect -37945 7635 -37910 7670
rect -37900 7635 -37865 7670
rect -37855 7635 -37820 7670
rect -37810 7635 -37775 7670
rect -37765 7635 -37730 7670
rect -37720 7635 -37685 7670
rect -37675 7635 -37640 7670
rect -37630 7635 -37595 7670
rect -37585 7635 -37550 7670
rect -37540 7635 -37505 7670
rect -37495 7635 -37460 7670
rect -37450 7635 -37415 7670
rect -37405 7635 -37370 7670
rect -37360 7635 -37325 7670
rect -37315 7635 -37280 7670
rect -37270 7635 -37235 7670
rect -37225 7635 -37190 7670
rect -38755 7590 -38720 7625
rect -38710 7590 -38675 7625
rect -38665 7590 -38630 7625
rect -38620 7590 -38585 7625
rect -38575 7590 -38540 7625
rect -38530 7590 -38495 7625
rect -38485 7590 -38450 7625
rect -38440 7590 -38405 7625
rect -38395 7590 -38360 7625
rect -38350 7590 -38315 7625
rect -38305 7590 -38270 7625
rect -38260 7590 -38225 7625
rect -38215 7590 -38180 7625
rect -38170 7590 -38135 7625
rect -38125 7590 -38090 7625
rect -38080 7590 -38045 7625
rect -38035 7590 -38000 7625
rect -37990 7590 -37955 7625
rect -37945 7590 -37910 7625
rect -37900 7590 -37865 7625
rect -37855 7590 -37820 7625
rect -37810 7590 -37775 7625
rect -37765 7590 -37730 7625
rect -37720 7590 -37685 7625
rect -37675 7590 -37640 7625
rect -37630 7590 -37595 7625
rect -37585 7590 -37550 7625
rect -37540 7590 -37505 7625
rect -37495 7590 -37460 7625
rect -37450 7590 -37415 7625
rect -37405 7590 -37370 7625
rect -37360 7590 -37325 7625
rect -37315 7590 -37280 7625
rect -37270 7590 -37235 7625
rect -37225 7590 -37190 7625
rect -38755 7545 -38720 7580
rect -38710 7545 -38675 7580
rect -38665 7545 -38630 7580
rect -38620 7545 -38585 7580
rect -38575 7545 -38540 7580
rect -38530 7545 -38495 7580
rect -38485 7545 -38450 7580
rect -38440 7545 -38405 7580
rect -38395 7545 -38360 7580
rect -38350 7545 -38315 7580
rect -38305 7545 -38270 7580
rect -38260 7545 -38225 7580
rect -38215 7545 -38180 7580
rect -38170 7545 -38135 7580
rect -38125 7545 -38090 7580
rect -38080 7545 -38045 7580
rect -38035 7545 -38000 7580
rect -37990 7545 -37955 7580
rect -37945 7545 -37910 7580
rect -37900 7545 -37865 7580
rect -37855 7545 -37820 7580
rect -37810 7545 -37775 7580
rect -37765 7545 -37730 7580
rect -37720 7545 -37685 7580
rect -37675 7545 -37640 7580
rect -37630 7545 -37595 7580
rect -37585 7545 -37550 7580
rect -37540 7545 -37505 7580
rect -37495 7545 -37460 7580
rect -37450 7545 -37415 7580
rect -37405 7545 -37370 7580
rect -37360 7545 -37325 7580
rect -37315 7545 -37280 7580
rect -37270 7545 -37235 7580
rect -37225 7545 -37190 7580
rect -38755 7500 -38720 7535
rect -38710 7500 -38675 7535
rect -38665 7500 -38630 7535
rect -38620 7500 -38585 7535
rect -38575 7500 -38540 7535
rect -38530 7500 -38495 7535
rect -38485 7500 -38450 7535
rect -38440 7500 -38405 7535
rect -38395 7500 -38360 7535
rect -38350 7500 -38315 7535
rect -38305 7500 -38270 7535
rect -38260 7500 -38225 7535
rect -38215 7500 -38180 7535
rect -38170 7500 -38135 7535
rect -38125 7500 -38090 7535
rect -38080 7500 -38045 7535
rect -38035 7500 -38000 7535
rect -37990 7500 -37955 7535
rect -37945 7500 -37910 7535
rect -37900 7500 -37865 7535
rect -37855 7500 -37820 7535
rect -37810 7500 -37775 7535
rect -37765 7500 -37730 7535
rect -37720 7500 -37685 7535
rect -37675 7500 -37640 7535
rect -37630 7500 -37595 7535
rect -37585 7500 -37550 7535
rect -37540 7500 -37505 7535
rect -37495 7500 -37460 7535
rect -37450 7500 -37415 7535
rect -37405 7500 -37370 7535
rect -37360 7500 -37325 7535
rect -37315 7500 -37280 7535
rect -37270 7500 -37235 7535
rect -37225 7500 -37190 7535
rect -38755 7455 -38720 7490
rect -38710 7455 -38675 7490
rect -38665 7455 -38630 7490
rect -38620 7455 -38585 7490
rect -38575 7455 -38540 7490
rect -38530 7455 -38495 7490
rect -38485 7455 -38450 7490
rect -38440 7455 -38405 7490
rect -38395 7455 -38360 7490
rect -38350 7455 -38315 7490
rect -38305 7455 -38270 7490
rect -38260 7455 -38225 7490
rect -38215 7455 -38180 7490
rect -38170 7455 -38135 7490
rect -38125 7455 -38090 7490
rect -38080 7455 -38045 7490
rect -38035 7455 -38000 7490
rect -37990 7455 -37955 7490
rect -37945 7455 -37910 7490
rect -37900 7455 -37865 7490
rect -37855 7455 -37820 7490
rect -37810 7455 -37775 7490
rect -37765 7455 -37730 7490
rect -37720 7455 -37685 7490
rect -37675 7455 -37640 7490
rect -37630 7455 -37595 7490
rect -37585 7455 -37550 7490
rect -37540 7455 -37505 7490
rect -37495 7455 -37460 7490
rect -37450 7455 -37415 7490
rect -37405 7455 -37370 7490
rect -37360 7455 -37325 7490
rect -37315 7455 -37280 7490
rect -37270 7455 -37235 7490
rect -37225 7455 -37190 7490
rect -38755 7410 -38720 7445
rect -38710 7410 -38675 7445
rect -38665 7410 -38630 7445
rect -38620 7410 -38585 7445
rect -38575 7410 -38540 7445
rect -38530 7410 -38495 7445
rect -38485 7410 -38450 7445
rect -38440 7410 -38405 7445
rect -38395 7410 -38360 7445
rect -38350 7410 -38315 7445
rect -38305 7410 -38270 7445
rect -38260 7410 -38225 7445
rect -38215 7410 -38180 7445
rect -38170 7410 -38135 7445
rect -38125 7410 -38090 7445
rect -38080 7410 -38045 7445
rect -38035 7410 -38000 7445
rect -37990 7410 -37955 7445
rect -37945 7410 -37910 7445
rect -37900 7410 -37865 7445
rect -37855 7410 -37820 7445
rect -37810 7410 -37775 7445
rect -37765 7410 -37730 7445
rect -37720 7410 -37685 7445
rect -37675 7410 -37640 7445
rect -37630 7410 -37595 7445
rect -37585 7410 -37550 7445
rect -37540 7410 -37505 7445
rect -37495 7410 -37460 7445
rect -37450 7410 -37415 7445
rect -37405 7410 -37370 7445
rect -37360 7410 -37325 7445
rect -37315 7410 -37280 7445
rect -37270 7410 -37235 7445
rect -37225 7410 -37190 7445
rect -38755 7365 -38720 7400
rect -38710 7365 -38675 7400
rect -38665 7365 -38630 7400
rect -38620 7365 -38585 7400
rect -38575 7365 -38540 7400
rect -38530 7365 -38495 7400
rect -38485 7365 -38450 7400
rect -38440 7365 -38405 7400
rect -38395 7365 -38360 7400
rect -38350 7365 -38315 7400
rect -38305 7365 -38270 7400
rect -38260 7365 -38225 7400
rect -38215 7365 -38180 7400
rect -38170 7365 -38135 7400
rect -38125 7365 -38090 7400
rect -38080 7365 -38045 7400
rect -38035 7365 -38000 7400
rect -37990 7365 -37955 7400
rect -37945 7365 -37910 7400
rect -37900 7365 -37865 7400
rect -37855 7365 -37820 7400
rect -37810 7365 -37775 7400
rect -37765 7365 -37730 7400
rect -37720 7365 -37685 7400
rect -37675 7365 -37640 7400
rect -37630 7365 -37595 7400
rect -37585 7365 -37550 7400
rect -37540 7365 -37505 7400
rect -37495 7365 -37460 7400
rect -37450 7365 -37415 7400
rect -37405 7365 -37370 7400
rect -37360 7365 -37325 7400
rect -37315 7365 -37280 7400
rect -37270 7365 -37235 7400
rect -37225 7365 -37190 7400
rect -38755 7320 -38720 7355
rect -38710 7320 -38675 7355
rect -38665 7320 -38630 7355
rect -38620 7320 -38585 7355
rect -38575 7320 -38540 7355
rect -38530 7320 -38495 7355
rect -38485 7320 -38450 7355
rect -38440 7320 -38405 7355
rect -38395 7320 -38360 7355
rect -38350 7320 -38315 7355
rect -38305 7320 -38270 7355
rect -38260 7320 -38225 7355
rect -38215 7320 -38180 7355
rect -38170 7320 -38135 7355
rect -38125 7320 -38090 7355
rect -38080 7320 -38045 7355
rect -38035 7320 -38000 7355
rect -37990 7320 -37955 7355
rect -37945 7320 -37910 7355
rect -37900 7320 -37865 7355
rect -37855 7320 -37820 7355
rect -37810 7320 -37775 7355
rect -37765 7320 -37730 7355
rect -37720 7320 -37685 7355
rect -37675 7320 -37640 7355
rect -37630 7320 -37595 7355
rect -37585 7320 -37550 7355
rect -37540 7320 -37505 7355
rect -37495 7320 -37460 7355
rect -37450 7320 -37415 7355
rect -37405 7320 -37370 7355
rect -37360 7320 -37325 7355
rect -37315 7320 -37280 7355
rect -37270 7320 -37235 7355
rect -37225 7320 -37190 7355
rect -38755 7275 -38720 7310
rect -38710 7275 -38675 7310
rect -38665 7275 -38630 7310
rect -38620 7275 -38585 7310
rect -38575 7275 -38540 7310
rect -38530 7275 -38495 7310
rect -38485 7275 -38450 7310
rect -38440 7275 -38405 7310
rect -38395 7275 -38360 7310
rect -38350 7275 -38315 7310
rect -38305 7275 -38270 7310
rect -38260 7275 -38225 7310
rect -38215 7275 -38180 7310
rect -38170 7275 -38135 7310
rect -38125 7275 -38090 7310
rect -38080 7275 -38045 7310
rect -38035 7275 -38000 7310
rect -37990 7275 -37955 7310
rect -37945 7275 -37910 7310
rect -37900 7275 -37865 7310
rect -37855 7275 -37820 7310
rect -37810 7275 -37775 7310
rect -37765 7275 -37730 7310
rect -37720 7275 -37685 7310
rect -37675 7275 -37640 7310
rect -37630 7275 -37595 7310
rect -37585 7275 -37550 7310
rect -37540 7275 -37505 7310
rect -37495 7275 -37460 7310
rect -37450 7275 -37415 7310
rect -37405 7275 -37370 7310
rect -37360 7275 -37325 7310
rect -37315 7275 -37280 7310
rect -37270 7275 -37235 7310
rect -37225 7275 -37190 7310
rect -38755 7230 -38720 7265
rect -38710 7230 -38675 7265
rect -38665 7230 -38630 7265
rect -38620 7230 -38585 7265
rect -38575 7230 -38540 7265
rect -38530 7230 -38495 7265
rect -38485 7230 -38450 7265
rect -38440 7230 -38405 7265
rect -38395 7230 -38360 7265
rect -38350 7230 -38315 7265
rect -38305 7230 -38270 7265
rect -38260 7230 -38225 7265
rect -38215 7230 -38180 7265
rect -38170 7230 -38135 7265
rect -38125 7230 -38090 7265
rect -38080 7230 -38045 7265
rect -38035 7230 -38000 7265
rect -37990 7230 -37955 7265
rect -37945 7230 -37910 7265
rect -37900 7230 -37865 7265
rect -37855 7230 -37820 7265
rect -37810 7230 -37775 7265
rect -37765 7230 -37730 7265
rect -37720 7230 -37685 7265
rect -37675 7230 -37640 7265
rect -37630 7230 -37595 7265
rect -37585 7230 -37550 7265
rect -37540 7230 -37505 7265
rect -37495 7230 -37460 7265
rect -37450 7230 -37415 7265
rect -37405 7230 -37370 7265
rect -37360 7230 -37325 7265
rect -37315 7230 -37280 7265
rect -37270 7230 -37235 7265
rect -37225 7230 -37190 7265
rect -38755 7185 -38720 7220
rect -38710 7185 -38675 7220
rect -38665 7185 -38630 7220
rect -38620 7185 -38585 7220
rect -38575 7185 -38540 7220
rect -38530 7185 -38495 7220
rect -38485 7185 -38450 7220
rect -38440 7185 -38405 7220
rect -38395 7185 -38360 7220
rect -38350 7185 -38315 7220
rect -38305 7185 -38270 7220
rect -38260 7185 -38225 7220
rect -38215 7185 -38180 7220
rect -38170 7185 -38135 7220
rect -38125 7185 -38090 7220
rect -38080 7185 -38045 7220
rect -38035 7185 -38000 7220
rect -37990 7185 -37955 7220
rect -37945 7185 -37910 7220
rect -37900 7185 -37865 7220
rect -37855 7185 -37820 7220
rect -37810 7185 -37775 7220
rect -37765 7185 -37730 7220
rect -37720 7185 -37685 7220
rect -37675 7185 -37640 7220
rect -37630 7185 -37595 7220
rect -37585 7185 -37550 7220
rect -37540 7185 -37505 7220
rect -37495 7185 -37460 7220
rect -37450 7185 -37415 7220
rect -37405 7185 -37370 7220
rect -37360 7185 -37325 7220
rect -37315 7185 -37280 7220
rect -37270 7185 -37235 7220
rect -37225 7185 -37190 7220
rect -38755 7140 -38720 7175
rect -38710 7140 -38675 7175
rect -38665 7140 -38630 7175
rect -38620 7140 -38585 7175
rect -38575 7140 -38540 7175
rect -38530 7140 -38495 7175
rect -38485 7140 -38450 7175
rect -38440 7140 -38405 7175
rect -38395 7140 -38360 7175
rect -38350 7140 -38315 7175
rect -38305 7140 -38270 7175
rect -38260 7140 -38225 7175
rect -38215 7140 -38180 7175
rect -38170 7140 -38135 7175
rect -38125 7140 -38090 7175
rect -38080 7140 -38045 7175
rect -38035 7140 -38000 7175
rect -37990 7140 -37955 7175
rect -37945 7140 -37910 7175
rect -37900 7140 -37865 7175
rect -37855 7140 -37820 7175
rect -37810 7140 -37775 7175
rect -37765 7140 -37730 7175
rect -37720 7140 -37685 7175
rect -37675 7140 -37640 7175
rect -37630 7140 -37595 7175
rect -37585 7140 -37550 7175
rect -37540 7140 -37505 7175
rect -37495 7140 -37460 7175
rect -37450 7140 -37415 7175
rect -37405 7140 -37370 7175
rect -37360 7140 -37325 7175
rect -37315 7140 -37280 7175
rect -37270 7140 -37235 7175
rect -37225 7140 -37190 7175
rect -38755 7095 -38720 7130
rect -38710 7095 -38675 7130
rect -38665 7095 -38630 7130
rect -38620 7095 -38585 7130
rect -38575 7095 -38540 7130
rect -38530 7095 -38495 7130
rect -38485 7095 -38450 7130
rect -38440 7095 -38405 7130
rect -38395 7095 -38360 7130
rect -38350 7095 -38315 7130
rect -38305 7095 -38270 7130
rect -38260 7095 -38225 7130
rect -38215 7095 -38180 7130
rect -38170 7095 -38135 7130
rect -38125 7095 -38090 7130
rect -38080 7095 -38045 7130
rect -38035 7095 -38000 7130
rect -37990 7095 -37955 7130
rect -37945 7095 -37910 7130
rect -37900 7095 -37865 7130
rect -37855 7095 -37820 7130
rect -37810 7095 -37775 7130
rect -37765 7095 -37730 7130
rect -37720 7095 -37685 7130
rect -37675 7095 -37640 7130
rect -37630 7095 -37595 7130
rect -37585 7095 -37550 7130
rect -37540 7095 -37505 7130
rect -37495 7095 -37460 7130
rect -37450 7095 -37415 7130
rect -37405 7095 -37370 7130
rect -37360 7095 -37325 7130
rect -37315 7095 -37280 7130
rect -37270 7095 -37235 7130
rect -37225 7095 -37190 7130
rect -38755 7050 -38720 7085
rect -38710 7050 -38675 7085
rect -38665 7050 -38630 7085
rect -38620 7050 -38585 7085
rect -38575 7050 -38540 7085
rect -38530 7050 -38495 7085
rect -38485 7050 -38450 7085
rect -38440 7050 -38405 7085
rect -38395 7050 -38360 7085
rect -38350 7050 -38315 7085
rect -38305 7050 -38270 7085
rect -38260 7050 -38225 7085
rect -38215 7050 -38180 7085
rect -38170 7050 -38135 7085
rect -38125 7050 -38090 7085
rect -38080 7050 -38045 7085
rect -38035 7050 -38000 7085
rect -37990 7050 -37955 7085
rect -37945 7050 -37910 7085
rect -37900 7050 -37865 7085
rect -37855 7050 -37820 7085
rect -37810 7050 -37775 7085
rect -37765 7050 -37730 7085
rect -37720 7050 -37685 7085
rect -37675 7050 -37640 7085
rect -37630 7050 -37595 7085
rect -37585 7050 -37550 7085
rect -37540 7050 -37505 7085
rect -37495 7050 -37460 7085
rect -37450 7050 -37415 7085
rect -37405 7050 -37370 7085
rect -37360 7050 -37325 7085
rect -37315 7050 -37280 7085
rect -37270 7050 -37235 7085
rect -37225 7050 -37190 7085
rect -38755 7005 -38720 7040
rect -38710 7005 -38675 7040
rect -38665 7005 -38630 7040
rect -38620 7005 -38585 7040
rect -38575 7005 -38540 7040
rect -38530 7005 -38495 7040
rect -38485 7005 -38450 7040
rect -38440 7005 -38405 7040
rect -38395 7005 -38360 7040
rect -38350 7005 -38315 7040
rect -38305 7005 -38270 7040
rect -38260 7005 -38225 7040
rect -38215 7005 -38180 7040
rect -38170 7005 -38135 7040
rect -38125 7005 -38090 7040
rect -38080 7005 -38045 7040
rect -38035 7005 -38000 7040
rect -37990 7005 -37955 7040
rect -37945 7005 -37910 7040
rect -37900 7005 -37865 7040
rect -37855 7005 -37820 7040
rect -37810 7005 -37775 7040
rect -37765 7005 -37730 7040
rect -37720 7005 -37685 7040
rect -37675 7005 -37640 7040
rect -37630 7005 -37595 7040
rect -37585 7005 -37550 7040
rect -37540 7005 -37505 7040
rect -37495 7005 -37460 7040
rect -37450 7005 -37415 7040
rect -37405 7005 -37370 7040
rect -37360 7005 -37325 7040
rect -37315 7005 -37280 7040
rect -37270 7005 -37235 7040
rect -37225 7005 -37190 7040
rect -38755 6960 -38720 6995
rect -38710 6960 -38675 6995
rect -38665 6960 -38630 6995
rect -38620 6960 -38585 6995
rect -38575 6960 -38540 6995
rect -38530 6960 -38495 6995
rect -38485 6960 -38450 6995
rect -38440 6960 -38405 6995
rect -38395 6960 -38360 6995
rect -38350 6960 -38315 6995
rect -38305 6960 -38270 6995
rect -38260 6960 -38225 6995
rect -38215 6960 -38180 6995
rect -38170 6960 -38135 6995
rect -38125 6960 -38090 6995
rect -38080 6960 -38045 6995
rect -38035 6960 -38000 6995
rect -37990 6960 -37955 6995
rect -37945 6960 -37910 6995
rect -37900 6960 -37865 6995
rect -37855 6960 -37820 6995
rect -37810 6960 -37775 6995
rect -37765 6960 -37730 6995
rect -37720 6960 -37685 6995
rect -37675 6960 -37640 6995
rect -37630 6960 -37595 6995
rect -37585 6960 -37550 6995
rect -37540 6960 -37505 6995
rect -37495 6960 -37460 6995
rect -37450 6960 -37415 6995
rect -37405 6960 -37370 6995
rect -37360 6960 -37325 6995
rect -37315 6960 -37280 6995
rect -37270 6960 -37235 6995
rect -37225 6960 -37190 6995
rect -38755 6915 -38720 6950
rect -38710 6915 -38675 6950
rect -38665 6915 -38630 6950
rect -38620 6915 -38585 6950
rect -38575 6915 -38540 6950
rect -38530 6915 -38495 6950
rect -38485 6915 -38450 6950
rect -38440 6915 -38405 6950
rect -38395 6915 -38360 6950
rect -38350 6915 -38315 6950
rect -38305 6915 -38270 6950
rect -38260 6915 -38225 6950
rect -38215 6915 -38180 6950
rect -38170 6915 -38135 6950
rect -38125 6915 -38090 6950
rect -38080 6915 -38045 6950
rect -38035 6915 -38000 6950
rect -37990 6915 -37955 6950
rect -37945 6915 -37910 6950
rect -37900 6915 -37865 6950
rect -37855 6915 -37820 6950
rect -37810 6915 -37775 6950
rect -37765 6915 -37730 6950
rect -37720 6915 -37685 6950
rect -37675 6915 -37640 6950
rect -37630 6915 -37595 6950
rect -37585 6915 -37550 6950
rect -37540 6915 -37505 6950
rect -37495 6915 -37460 6950
rect -37450 6915 -37415 6950
rect -37405 6915 -37370 6950
rect -37360 6915 -37325 6950
rect -37315 6915 -37280 6950
rect -37270 6915 -37235 6950
rect -37225 6915 -37190 6950
rect -38755 6870 -38720 6905
rect -38710 6870 -38675 6905
rect -38665 6870 -38630 6905
rect -38620 6870 -38585 6905
rect -38575 6870 -38540 6905
rect -38530 6870 -38495 6905
rect -38485 6870 -38450 6905
rect -38440 6870 -38405 6905
rect -38395 6870 -38360 6905
rect -38350 6870 -38315 6905
rect -38305 6870 -38270 6905
rect -38260 6870 -38225 6905
rect -38215 6870 -38180 6905
rect -38170 6870 -38135 6905
rect -38125 6870 -38090 6905
rect -38080 6870 -38045 6905
rect -38035 6870 -38000 6905
rect -37990 6870 -37955 6905
rect -37945 6870 -37910 6905
rect -37900 6870 -37865 6905
rect -37855 6870 -37820 6905
rect -37810 6870 -37775 6905
rect -37765 6870 -37730 6905
rect -37720 6870 -37685 6905
rect -37675 6870 -37640 6905
rect -37630 6870 -37595 6905
rect -37585 6870 -37550 6905
rect -37540 6870 -37505 6905
rect -37495 6870 -37460 6905
rect -37450 6870 -37415 6905
rect -37405 6870 -37370 6905
rect -37360 6870 -37325 6905
rect -37315 6870 -37280 6905
rect -37270 6870 -37235 6905
rect -37225 6870 -37190 6905
rect -38755 6825 -38720 6860
rect -38710 6825 -38675 6860
rect -38665 6825 -38630 6860
rect -38620 6825 -38585 6860
rect -38575 6825 -38540 6860
rect -38530 6825 -38495 6860
rect -38485 6825 -38450 6860
rect -38440 6825 -38405 6860
rect -38395 6825 -38360 6860
rect -38350 6825 -38315 6860
rect -38305 6825 -38270 6860
rect -38260 6825 -38225 6860
rect -38215 6825 -38180 6860
rect -38170 6825 -38135 6860
rect -38125 6825 -38090 6860
rect -38080 6825 -38045 6860
rect -38035 6825 -38000 6860
rect -37990 6825 -37955 6860
rect -37945 6825 -37910 6860
rect -37900 6825 -37865 6860
rect -37855 6825 -37820 6860
rect -37810 6825 -37775 6860
rect -37765 6825 -37730 6860
rect -37720 6825 -37685 6860
rect -37675 6825 -37640 6860
rect -37630 6825 -37595 6860
rect -37585 6825 -37550 6860
rect -37540 6825 -37505 6860
rect -37495 6825 -37460 6860
rect -37450 6825 -37415 6860
rect -37405 6825 -37370 6860
rect -37360 6825 -37325 6860
rect -37315 6825 -37280 6860
rect -37270 6825 -37235 6860
rect -37225 6825 -37190 6860
rect -38755 6780 -38720 6815
rect -38710 6780 -38675 6815
rect -38665 6780 -38630 6815
rect -38620 6780 -38585 6815
rect -38575 6780 -38540 6815
rect -38530 6780 -38495 6815
rect -38485 6780 -38450 6815
rect -38440 6780 -38405 6815
rect -38395 6780 -38360 6815
rect -38350 6780 -38315 6815
rect -38305 6780 -38270 6815
rect -38260 6780 -38225 6815
rect -38215 6780 -38180 6815
rect -38170 6780 -38135 6815
rect -38125 6780 -38090 6815
rect -38080 6780 -38045 6815
rect -38035 6780 -38000 6815
rect -37990 6780 -37955 6815
rect -37945 6780 -37910 6815
rect -37900 6780 -37865 6815
rect -37855 6780 -37820 6815
rect -37810 6780 -37775 6815
rect -37765 6780 -37730 6815
rect -37720 6780 -37685 6815
rect -37675 6780 -37640 6815
rect -37630 6780 -37595 6815
rect -37585 6780 -37550 6815
rect -37540 6780 -37505 6815
rect -37495 6780 -37460 6815
rect -37450 6780 -37415 6815
rect -37405 6780 -37370 6815
rect -37360 6780 -37325 6815
rect -37315 6780 -37280 6815
rect -37270 6780 -37235 6815
rect -37225 6780 -37190 6815
rect -38755 6735 -38720 6770
rect -38710 6735 -38675 6770
rect -38665 6735 -38630 6770
rect -38620 6735 -38585 6770
rect -38575 6735 -38540 6770
rect -38530 6735 -38495 6770
rect -38485 6735 -38450 6770
rect -38440 6735 -38405 6770
rect -38395 6735 -38360 6770
rect -38350 6735 -38315 6770
rect -38305 6735 -38270 6770
rect -38260 6735 -38225 6770
rect -38215 6735 -38180 6770
rect -38170 6735 -38135 6770
rect -38125 6735 -38090 6770
rect -38080 6735 -38045 6770
rect -38035 6735 -38000 6770
rect -37990 6735 -37955 6770
rect -37945 6735 -37910 6770
rect -37900 6735 -37865 6770
rect -37855 6735 -37820 6770
rect -37810 6735 -37775 6770
rect -37765 6735 -37730 6770
rect -37720 6735 -37685 6770
rect -37675 6735 -37640 6770
rect -37630 6735 -37595 6770
rect -37585 6735 -37550 6770
rect -37540 6735 -37505 6770
rect -37495 6735 -37460 6770
rect -37450 6735 -37415 6770
rect -37405 6735 -37370 6770
rect -37360 6735 -37325 6770
rect -37315 6735 -37280 6770
rect -37270 6735 -37235 6770
rect -37225 6735 -37190 6770
rect -38755 6690 -38720 6725
rect -38710 6690 -38675 6725
rect -38665 6690 -38630 6725
rect -38620 6690 -38585 6725
rect -38575 6690 -38540 6725
rect -38530 6690 -38495 6725
rect -38485 6690 -38450 6725
rect -38440 6690 -38405 6725
rect -38395 6690 -38360 6725
rect -38350 6690 -38315 6725
rect -38305 6690 -38270 6725
rect -38260 6690 -38225 6725
rect -38215 6690 -38180 6725
rect -38170 6690 -38135 6725
rect -38125 6690 -38090 6725
rect -38080 6690 -38045 6725
rect -38035 6690 -38000 6725
rect -37990 6690 -37955 6725
rect -37945 6690 -37910 6725
rect -37900 6690 -37865 6725
rect -37855 6690 -37820 6725
rect -37810 6690 -37775 6725
rect -37765 6690 -37730 6725
rect -37720 6690 -37685 6725
rect -37675 6690 -37640 6725
rect -37630 6690 -37595 6725
rect -37585 6690 -37550 6725
rect -37540 6690 -37505 6725
rect -37495 6690 -37460 6725
rect -37450 6690 -37415 6725
rect -37405 6690 -37370 6725
rect -37360 6690 -37325 6725
rect -37315 6690 -37280 6725
rect -37270 6690 -37235 6725
rect -37225 6690 -37190 6725
rect -38755 6645 -38720 6680
rect -38710 6645 -38675 6680
rect -38665 6645 -38630 6680
rect -38620 6645 -38585 6680
rect -38575 6645 -38540 6680
rect -38530 6645 -38495 6680
rect -38485 6645 -38450 6680
rect -38440 6645 -38405 6680
rect -38395 6645 -38360 6680
rect -38350 6645 -38315 6680
rect -38305 6645 -38270 6680
rect -38260 6645 -38225 6680
rect -38215 6645 -38180 6680
rect -38170 6645 -38135 6680
rect -38125 6645 -38090 6680
rect -38080 6645 -38045 6680
rect -38035 6645 -38000 6680
rect -37990 6645 -37955 6680
rect -37945 6645 -37910 6680
rect -37900 6645 -37865 6680
rect -37855 6645 -37820 6680
rect -37810 6645 -37775 6680
rect -37765 6645 -37730 6680
rect -37720 6645 -37685 6680
rect -37675 6645 -37640 6680
rect -37630 6645 -37595 6680
rect -37585 6645 -37550 6680
rect -37540 6645 -37505 6680
rect -37495 6645 -37460 6680
rect -37450 6645 -37415 6680
rect -37405 6645 -37370 6680
rect -37360 6645 -37325 6680
rect -37315 6645 -37280 6680
rect -37270 6645 -37235 6680
rect -37225 6645 -37190 6680
rect -38755 6600 -38720 6635
rect -38710 6600 -38675 6635
rect -38665 6600 -38630 6635
rect -38620 6600 -38585 6635
rect -38575 6600 -38540 6635
rect -38530 6600 -38495 6635
rect -38485 6600 -38450 6635
rect -38440 6600 -38405 6635
rect -38395 6600 -38360 6635
rect -38350 6600 -38315 6635
rect -38305 6600 -38270 6635
rect -38260 6600 -38225 6635
rect -38215 6600 -38180 6635
rect -38170 6600 -38135 6635
rect -38125 6600 -38090 6635
rect -38080 6600 -38045 6635
rect -38035 6600 -38000 6635
rect -37990 6600 -37955 6635
rect -37945 6600 -37910 6635
rect -37900 6600 -37865 6635
rect -37855 6600 -37820 6635
rect -37810 6600 -37775 6635
rect -37765 6600 -37730 6635
rect -37720 6600 -37685 6635
rect -37675 6600 -37640 6635
rect -37630 6600 -37595 6635
rect -37585 6600 -37550 6635
rect -37540 6600 -37505 6635
rect -37495 6600 -37460 6635
rect -37450 6600 -37415 6635
rect -37405 6600 -37370 6635
rect -37360 6600 -37325 6635
rect -37315 6600 -37280 6635
rect -37270 6600 -37235 6635
rect -37225 6600 -37190 6635
rect -38755 6555 -38720 6590
rect -38710 6555 -38675 6590
rect -38665 6555 -38630 6590
rect -38620 6555 -38585 6590
rect -38575 6555 -38540 6590
rect -38530 6555 -38495 6590
rect -38485 6555 -38450 6590
rect -38440 6555 -38405 6590
rect -38395 6555 -38360 6590
rect -38350 6555 -38315 6590
rect -38305 6555 -38270 6590
rect -38260 6555 -38225 6590
rect -38215 6555 -38180 6590
rect -38170 6555 -38135 6590
rect -38125 6555 -38090 6590
rect -38080 6555 -38045 6590
rect -38035 6555 -38000 6590
rect -37990 6555 -37955 6590
rect -37945 6555 -37910 6590
rect -37900 6555 -37865 6590
rect -37855 6555 -37820 6590
rect -37810 6555 -37775 6590
rect -37765 6555 -37730 6590
rect -37720 6555 -37685 6590
rect -37675 6555 -37640 6590
rect -37630 6555 -37595 6590
rect -37585 6555 -37550 6590
rect -37540 6555 -37505 6590
rect -37495 6555 -37460 6590
rect -37450 6555 -37415 6590
rect -37405 6555 -37370 6590
rect -37360 6555 -37325 6590
rect -37315 6555 -37280 6590
rect -37270 6555 -37235 6590
rect -37225 6555 -37190 6590
rect -38755 6510 -38720 6545
rect -38710 6510 -38675 6545
rect -38665 6510 -38630 6545
rect -38620 6510 -38585 6545
rect -38575 6510 -38540 6545
rect -38530 6510 -38495 6545
rect -38485 6510 -38450 6545
rect -38440 6510 -38405 6545
rect -38395 6510 -38360 6545
rect -38350 6510 -38315 6545
rect -38305 6510 -38270 6545
rect -38260 6510 -38225 6545
rect -38215 6510 -38180 6545
rect -38170 6510 -38135 6545
rect -38125 6510 -38090 6545
rect -38080 6510 -38045 6545
rect -38035 6510 -38000 6545
rect -37990 6510 -37955 6545
rect -37945 6510 -37910 6545
rect -37900 6510 -37865 6545
rect -37855 6510 -37820 6545
rect -37810 6510 -37775 6545
rect -37765 6510 -37730 6545
rect -37720 6510 -37685 6545
rect -37675 6510 -37640 6545
rect -37630 6510 -37595 6545
rect -37585 6510 -37550 6545
rect -37540 6510 -37505 6545
rect -37495 6510 -37460 6545
rect -37450 6510 -37415 6545
rect -37405 6510 -37370 6545
rect -37360 6510 -37325 6545
rect -37315 6510 -37280 6545
rect -37270 6510 -37235 6545
rect -37225 6510 -37190 6545
rect -38755 6465 -38720 6500
rect -38710 6465 -38675 6500
rect -38665 6465 -38630 6500
rect -38620 6465 -38585 6500
rect -38575 6465 -38540 6500
rect -38530 6465 -38495 6500
rect -38485 6465 -38450 6500
rect -38440 6465 -38405 6500
rect -38395 6465 -38360 6500
rect -38350 6465 -38315 6500
rect -38305 6465 -38270 6500
rect -38260 6465 -38225 6500
rect -38215 6465 -38180 6500
rect -38170 6465 -38135 6500
rect -38125 6465 -38090 6500
rect -38080 6465 -38045 6500
rect -38035 6465 -38000 6500
rect -37990 6465 -37955 6500
rect -37945 6465 -37910 6500
rect -37900 6465 -37865 6500
rect -37855 6465 -37820 6500
rect -37810 6465 -37775 6500
rect -37765 6465 -37730 6500
rect -37720 6465 -37685 6500
rect -37675 6465 -37640 6500
rect -37630 6465 -37595 6500
rect -37585 6465 -37550 6500
rect -37540 6465 -37505 6500
rect -37495 6465 -37460 6500
rect -37450 6465 -37415 6500
rect -37405 6465 -37370 6500
rect -37360 6465 -37325 6500
rect -37315 6465 -37280 6500
rect -37270 6465 -37235 6500
rect -37225 6465 -37190 6500
rect -80 9635 -40 9640
rect -80 9605 -75 9635
rect -75 9605 -45 9635
rect -45 9605 -40 9635
rect -80 9600 -40 9605
rect -80 9570 -40 9575
rect -80 9540 -75 9570
rect -75 9540 -45 9570
rect -45 9540 -40 9570
rect -80 9535 -40 9540
rect -80 9500 -40 9505
rect -80 9470 -75 9500
rect -75 9470 -45 9500
rect -45 9470 -40 9500
rect -80 9465 -40 9470
rect -80 9430 -40 9435
rect -80 9400 -75 9430
rect -75 9400 -45 9430
rect -45 9400 -40 9430
rect -80 9395 -40 9400
rect -80 9360 -40 9365
rect -80 9330 -75 9360
rect -75 9330 -45 9360
rect -45 9330 -40 9360
rect -80 9325 -40 9330
rect -80 9295 -40 9300
rect -80 9265 -75 9295
rect -75 9265 -45 9295
rect -45 9265 -40 9295
rect -80 9260 -40 9265
rect -80 9235 -40 9240
rect -80 9205 -75 9235
rect -75 9205 -45 9235
rect -45 9205 -40 9235
rect -80 9200 -40 9205
rect -80 9170 -40 9175
rect -80 9140 -75 9170
rect -75 9140 -45 9170
rect -45 9140 -40 9170
rect -80 9135 -40 9140
rect -80 9100 -40 9105
rect -80 9070 -75 9100
rect -75 9070 -45 9100
rect -45 9070 -40 9100
rect -80 9065 -40 9070
rect -80 9030 -40 9035
rect -80 9000 -75 9030
rect -75 9000 -45 9030
rect -45 9000 -40 9030
rect -80 8995 -40 9000
rect -80 8960 -40 8965
rect -80 8930 -75 8960
rect -75 8930 -45 8960
rect -45 8930 -40 8960
rect -80 8925 -40 8930
rect -80 8895 -40 8900
rect -80 8865 -75 8895
rect -75 8865 -45 8895
rect -45 8865 -40 8895
rect -80 8860 -40 8865
rect -80 8835 -40 8840
rect -80 8805 -75 8835
rect -75 8805 -45 8835
rect -45 8805 -40 8835
rect -80 8800 -40 8805
rect -80 8770 -40 8775
rect -80 8740 -75 8770
rect -75 8740 -45 8770
rect -45 8740 -40 8770
rect -80 8735 -40 8740
rect -80 8700 -40 8705
rect -80 8670 -75 8700
rect -75 8670 -45 8700
rect -45 8670 -40 8700
rect -80 8665 -40 8670
rect -80 8630 -40 8635
rect -80 8600 -75 8630
rect -75 8600 -45 8630
rect -45 8600 -40 8630
rect -80 8595 -40 8600
rect -80 8560 -40 8565
rect -80 8530 -75 8560
rect -75 8530 -45 8560
rect -45 8530 -40 8560
rect -80 8525 -40 8530
rect -80 8495 -40 8500
rect -80 8465 -75 8495
rect -75 8465 -45 8495
rect -45 8465 -40 8495
rect -80 8460 -40 8465
rect -80 8435 -40 8440
rect -80 8405 -75 8435
rect -75 8405 -45 8435
rect -45 8405 -40 8435
rect -80 8400 -40 8405
rect -80 8370 -40 8375
rect -80 8340 -75 8370
rect -75 8340 -45 8370
rect -45 8340 -40 8370
rect -80 8335 -40 8340
rect -80 8300 -40 8305
rect -80 8270 -75 8300
rect -75 8270 -45 8300
rect -45 8270 -40 8300
rect -80 8265 -40 8270
rect -80 8230 -40 8235
rect -80 8200 -75 8230
rect -75 8200 -45 8230
rect -45 8200 -40 8230
rect -80 8195 -40 8200
rect -80 8160 -40 8165
rect -80 8130 -75 8160
rect -75 8130 -45 8160
rect -45 8130 -40 8160
rect -80 8125 -40 8130
rect -80 8095 -40 8100
rect -80 8065 -75 8095
rect -75 8065 -45 8095
rect -45 8065 -40 8095
rect -80 8060 -40 8065
rect -80 8035 -40 8040
rect -80 8005 -75 8035
rect -75 8005 -45 8035
rect -45 8005 -40 8035
rect -80 8000 -40 8005
rect -80 7970 -40 7975
rect -80 7940 -75 7970
rect -75 7940 -45 7970
rect -45 7940 -40 7970
rect -80 7935 -40 7940
rect -80 7900 -40 7905
rect -80 7870 -75 7900
rect -75 7870 -45 7900
rect -45 7870 -40 7900
rect -80 7865 -40 7870
rect -80 7830 -40 7835
rect -80 7800 -75 7830
rect -75 7800 -45 7830
rect -45 7800 -40 7830
rect -80 7795 -40 7800
rect -80 7760 -40 7765
rect -80 7730 -75 7760
rect -75 7730 -45 7760
rect -45 7730 -40 7760
rect -80 7725 -40 7730
rect -80 7695 -40 7700
rect -80 7665 -75 7695
rect -75 7665 -45 7695
rect -45 7665 -40 7695
rect -80 7660 -40 7665
rect -80 7635 -40 7640
rect -80 7605 -75 7635
rect -75 7605 -45 7635
rect -45 7605 -40 7635
rect -80 7600 -40 7605
rect -80 7570 -40 7575
rect -80 7540 -75 7570
rect -75 7540 -45 7570
rect -45 7540 -40 7570
rect -80 7535 -40 7540
rect -80 7500 -40 7505
rect -80 7470 -75 7500
rect -75 7470 -45 7500
rect -45 7470 -40 7500
rect -80 7465 -40 7470
rect -80 7430 -40 7435
rect -80 7400 -75 7430
rect -75 7400 -45 7430
rect -45 7400 -40 7430
rect -80 7395 -40 7400
rect -80 7360 -40 7365
rect -80 7330 -75 7360
rect -75 7330 -45 7360
rect -45 7330 -40 7360
rect -80 7325 -40 7330
rect -80 7295 -40 7300
rect -80 7265 -75 7295
rect -75 7265 -45 7295
rect -45 7265 -40 7295
rect -80 7260 -40 7265
rect -80 7235 -40 7240
rect -80 7205 -75 7235
rect -75 7205 -45 7235
rect -45 7205 -40 7235
rect -80 7200 -40 7205
rect -80 7170 -40 7175
rect -80 7140 -75 7170
rect -75 7140 -45 7170
rect -45 7140 -40 7170
rect -80 7135 -40 7140
rect -80 7100 -40 7105
rect -80 7070 -75 7100
rect -75 7070 -45 7100
rect -45 7070 -40 7100
rect -80 7065 -40 7070
rect -80 7030 -40 7035
rect -80 7000 -75 7030
rect -75 7000 -45 7030
rect -45 7000 -40 7030
rect -80 6995 -40 7000
rect -80 6960 -40 6965
rect -80 6930 -75 6960
rect -75 6930 -45 6960
rect -45 6930 -40 6960
rect -80 6925 -40 6930
rect -80 6895 -40 6900
rect -80 6865 -75 6895
rect -75 6865 -45 6895
rect -45 6865 -40 6895
rect -80 6860 -40 6865
rect -80 6835 -40 6840
rect -80 6805 -75 6835
rect -75 6805 -45 6835
rect -45 6805 -40 6835
rect -80 6800 -40 6805
rect -80 6770 -40 6775
rect -80 6740 -75 6770
rect -75 6740 -45 6770
rect -45 6740 -40 6770
rect -80 6735 -40 6740
rect -80 6700 -40 6705
rect -80 6670 -75 6700
rect -75 6670 -45 6700
rect -45 6670 -40 6700
rect -80 6665 -40 6670
rect -80 6630 -40 6635
rect -80 6600 -75 6630
rect -75 6600 -45 6630
rect -45 6600 -40 6630
rect -80 6595 -40 6600
rect -80 6560 -40 6565
rect -80 6530 -75 6560
rect -75 6530 -45 6560
rect -45 6530 -40 6560
rect -80 6525 -40 6530
rect -80 6495 -40 6500
rect -80 6465 -75 6495
rect -75 6465 -45 6495
rect -45 6465 -40 6495
rect -80 6460 -40 6465
rect 270 9635 310 9640
rect 270 9605 275 9635
rect 275 9605 305 9635
rect 305 9605 310 9635
rect 270 9600 310 9605
rect 270 9570 310 9575
rect 270 9540 275 9570
rect 275 9540 305 9570
rect 305 9540 310 9570
rect 270 9535 310 9540
rect 270 9500 310 9505
rect 270 9470 275 9500
rect 275 9470 305 9500
rect 305 9470 310 9500
rect 270 9465 310 9470
rect 270 9430 310 9435
rect 270 9400 275 9430
rect 275 9400 305 9430
rect 305 9400 310 9430
rect 270 9395 310 9400
rect 270 9360 310 9365
rect 270 9330 275 9360
rect 275 9330 305 9360
rect 305 9330 310 9360
rect 270 9325 310 9330
rect 270 9295 310 9300
rect 270 9265 275 9295
rect 275 9265 305 9295
rect 305 9265 310 9295
rect 270 9260 310 9265
rect 270 9235 310 9240
rect 270 9205 275 9235
rect 275 9205 305 9235
rect 305 9205 310 9235
rect 270 9200 310 9205
rect 270 9170 310 9175
rect 270 9140 275 9170
rect 275 9140 305 9170
rect 305 9140 310 9170
rect 270 9135 310 9140
rect 270 9100 310 9105
rect 270 9070 275 9100
rect 275 9070 305 9100
rect 305 9070 310 9100
rect 270 9065 310 9070
rect 270 9030 310 9035
rect 270 9000 275 9030
rect 275 9000 305 9030
rect 305 9000 310 9030
rect 270 8995 310 9000
rect 270 8960 310 8965
rect 270 8930 275 8960
rect 275 8930 305 8960
rect 305 8930 310 8960
rect 270 8925 310 8930
rect 270 8895 310 8900
rect 270 8865 275 8895
rect 275 8865 305 8895
rect 305 8865 310 8895
rect 270 8860 310 8865
rect 270 8835 310 8840
rect 270 8805 275 8835
rect 275 8805 305 8835
rect 305 8805 310 8835
rect 270 8800 310 8805
rect 270 8770 310 8775
rect 270 8740 275 8770
rect 275 8740 305 8770
rect 305 8740 310 8770
rect 270 8735 310 8740
rect 270 8700 310 8705
rect 270 8670 275 8700
rect 275 8670 305 8700
rect 305 8670 310 8700
rect 270 8665 310 8670
rect 270 8630 310 8635
rect 270 8600 275 8630
rect 275 8600 305 8630
rect 305 8600 310 8630
rect 270 8595 310 8600
rect 270 8560 310 8565
rect 270 8530 275 8560
rect 275 8530 305 8560
rect 305 8530 310 8560
rect 270 8525 310 8530
rect 270 8495 310 8500
rect 270 8465 275 8495
rect 275 8465 305 8495
rect 305 8465 310 8495
rect 270 8460 310 8465
rect 270 8435 310 8440
rect 270 8405 275 8435
rect 275 8405 305 8435
rect 305 8405 310 8435
rect 270 8400 310 8405
rect 270 8370 310 8375
rect 270 8340 275 8370
rect 275 8340 305 8370
rect 305 8340 310 8370
rect 270 8335 310 8340
rect 270 8300 310 8305
rect 270 8270 275 8300
rect 275 8270 305 8300
rect 305 8270 310 8300
rect 270 8265 310 8270
rect 270 8230 310 8235
rect 270 8200 275 8230
rect 275 8200 305 8230
rect 305 8200 310 8230
rect 270 8195 310 8200
rect 270 8160 310 8165
rect 270 8130 275 8160
rect 275 8130 305 8160
rect 305 8130 310 8160
rect 270 8125 310 8130
rect 270 8095 310 8100
rect 270 8065 275 8095
rect 275 8065 305 8095
rect 305 8065 310 8095
rect 270 8060 310 8065
rect 270 8035 310 8040
rect 270 8005 275 8035
rect 275 8005 305 8035
rect 305 8005 310 8035
rect 270 8000 310 8005
rect 270 7970 310 7975
rect 270 7940 275 7970
rect 275 7940 305 7970
rect 305 7940 310 7970
rect 270 7935 310 7940
rect 270 7900 310 7905
rect 270 7870 275 7900
rect 275 7870 305 7900
rect 305 7870 310 7900
rect 270 7865 310 7870
rect 270 7830 310 7835
rect 270 7800 275 7830
rect 275 7800 305 7830
rect 305 7800 310 7830
rect 270 7795 310 7800
rect 270 7760 310 7765
rect 270 7730 275 7760
rect 275 7730 305 7760
rect 305 7730 310 7760
rect 270 7725 310 7730
rect 270 7695 310 7700
rect 270 7665 275 7695
rect 275 7665 305 7695
rect 305 7665 310 7695
rect 270 7660 310 7665
rect 270 7635 310 7640
rect 270 7605 275 7635
rect 275 7605 305 7635
rect 305 7605 310 7635
rect 270 7600 310 7605
rect 270 7570 310 7575
rect 270 7540 275 7570
rect 275 7540 305 7570
rect 305 7540 310 7570
rect 270 7535 310 7540
rect 270 7500 310 7505
rect 270 7470 275 7500
rect 275 7470 305 7500
rect 305 7470 310 7500
rect 270 7465 310 7470
rect 270 7430 310 7435
rect 270 7400 275 7430
rect 275 7400 305 7430
rect 305 7400 310 7430
rect 270 7395 310 7400
rect 270 7360 310 7365
rect 270 7330 275 7360
rect 275 7330 305 7360
rect 305 7330 310 7360
rect 270 7325 310 7330
rect 270 7295 310 7300
rect 270 7265 275 7295
rect 275 7265 305 7295
rect 305 7265 310 7295
rect 270 7260 310 7265
rect 270 7235 310 7240
rect 270 7205 275 7235
rect 275 7205 305 7235
rect 305 7205 310 7235
rect 270 7200 310 7205
rect 270 7170 310 7175
rect 270 7140 275 7170
rect 275 7140 305 7170
rect 305 7140 310 7170
rect 270 7135 310 7140
rect 270 7100 310 7105
rect 270 7070 275 7100
rect 275 7070 305 7100
rect 305 7070 310 7100
rect 270 7065 310 7070
rect 270 7030 310 7035
rect 270 7000 275 7030
rect 275 7000 305 7030
rect 305 7000 310 7030
rect 270 6995 310 7000
rect 270 6960 310 6965
rect 270 6930 275 6960
rect 275 6930 305 6960
rect 305 6930 310 6960
rect 270 6925 310 6930
rect 270 6895 310 6900
rect 270 6865 275 6895
rect 275 6865 305 6895
rect 305 6865 310 6895
rect 270 6860 310 6865
rect 270 6835 310 6840
rect 270 6805 275 6835
rect 275 6805 305 6835
rect 305 6805 310 6835
rect 270 6800 310 6805
rect 270 6770 310 6775
rect 270 6740 275 6770
rect 275 6740 305 6770
rect 305 6740 310 6770
rect 270 6735 310 6740
rect 270 6700 310 6705
rect 270 6670 275 6700
rect 275 6670 305 6700
rect 305 6670 310 6700
rect 270 6665 310 6670
rect 270 6630 310 6635
rect 270 6600 275 6630
rect 275 6600 305 6630
rect 305 6600 310 6630
rect 270 6595 310 6600
rect 270 6560 310 6565
rect 270 6530 275 6560
rect 275 6530 305 6560
rect 305 6530 310 6560
rect 270 6525 310 6530
rect 270 6495 310 6500
rect 270 6465 275 6495
rect 275 6465 305 6495
rect 305 6465 310 6495
rect 270 6460 310 6465
rect 620 9635 660 9640
rect 620 9605 625 9635
rect 625 9605 655 9635
rect 655 9605 660 9635
rect 620 9600 660 9605
rect 620 9570 660 9575
rect 620 9540 625 9570
rect 625 9540 655 9570
rect 655 9540 660 9570
rect 620 9535 660 9540
rect 620 9500 660 9505
rect 620 9470 625 9500
rect 625 9470 655 9500
rect 655 9470 660 9500
rect 620 9465 660 9470
rect 620 9430 660 9435
rect 620 9400 625 9430
rect 625 9400 655 9430
rect 655 9400 660 9430
rect 620 9395 660 9400
rect 620 9360 660 9365
rect 620 9330 625 9360
rect 625 9330 655 9360
rect 655 9330 660 9360
rect 620 9325 660 9330
rect 620 9295 660 9300
rect 620 9265 625 9295
rect 625 9265 655 9295
rect 655 9265 660 9295
rect 620 9260 660 9265
rect 620 9235 660 9240
rect 620 9205 625 9235
rect 625 9205 655 9235
rect 655 9205 660 9235
rect 620 9200 660 9205
rect 620 9170 660 9175
rect 620 9140 625 9170
rect 625 9140 655 9170
rect 655 9140 660 9170
rect 620 9135 660 9140
rect 620 9100 660 9105
rect 620 9070 625 9100
rect 625 9070 655 9100
rect 655 9070 660 9100
rect 620 9065 660 9070
rect 620 9030 660 9035
rect 620 9000 625 9030
rect 625 9000 655 9030
rect 655 9000 660 9030
rect 620 8995 660 9000
rect 620 8960 660 8965
rect 620 8930 625 8960
rect 625 8930 655 8960
rect 655 8930 660 8960
rect 620 8925 660 8930
rect 620 8895 660 8900
rect 620 8865 625 8895
rect 625 8865 655 8895
rect 655 8865 660 8895
rect 620 8860 660 8865
rect 620 8835 660 8840
rect 620 8805 625 8835
rect 625 8805 655 8835
rect 655 8805 660 8835
rect 620 8800 660 8805
rect 620 8770 660 8775
rect 620 8740 625 8770
rect 625 8740 655 8770
rect 655 8740 660 8770
rect 620 8735 660 8740
rect 620 8700 660 8705
rect 620 8670 625 8700
rect 625 8670 655 8700
rect 655 8670 660 8700
rect 620 8665 660 8670
rect 620 8630 660 8635
rect 620 8600 625 8630
rect 625 8600 655 8630
rect 655 8600 660 8630
rect 620 8595 660 8600
rect 620 8560 660 8565
rect 620 8530 625 8560
rect 625 8530 655 8560
rect 655 8530 660 8560
rect 620 8525 660 8530
rect 620 8495 660 8500
rect 620 8465 625 8495
rect 625 8465 655 8495
rect 655 8465 660 8495
rect 620 8460 660 8465
rect 620 8435 660 8440
rect 620 8405 625 8435
rect 625 8405 655 8435
rect 655 8405 660 8435
rect 620 8400 660 8405
rect 620 8370 660 8375
rect 620 8340 625 8370
rect 625 8340 655 8370
rect 655 8340 660 8370
rect 620 8335 660 8340
rect 620 8300 660 8305
rect 620 8270 625 8300
rect 625 8270 655 8300
rect 655 8270 660 8300
rect 620 8265 660 8270
rect 620 8230 660 8235
rect 620 8200 625 8230
rect 625 8200 655 8230
rect 655 8200 660 8230
rect 620 8195 660 8200
rect 620 8160 660 8165
rect 620 8130 625 8160
rect 625 8130 655 8160
rect 655 8130 660 8160
rect 620 8125 660 8130
rect 620 8095 660 8100
rect 620 8065 625 8095
rect 625 8065 655 8095
rect 655 8065 660 8095
rect 620 8060 660 8065
rect 620 8035 660 8040
rect 620 8005 625 8035
rect 625 8005 655 8035
rect 655 8005 660 8035
rect 620 8000 660 8005
rect 620 7970 660 7975
rect 620 7940 625 7970
rect 625 7940 655 7970
rect 655 7940 660 7970
rect 620 7935 660 7940
rect 620 7900 660 7905
rect 620 7870 625 7900
rect 625 7870 655 7900
rect 655 7870 660 7900
rect 620 7865 660 7870
rect 620 7830 660 7835
rect 620 7800 625 7830
rect 625 7800 655 7830
rect 655 7800 660 7830
rect 620 7795 660 7800
rect 620 7760 660 7765
rect 620 7730 625 7760
rect 625 7730 655 7760
rect 655 7730 660 7760
rect 620 7725 660 7730
rect 620 7695 660 7700
rect 620 7665 625 7695
rect 625 7665 655 7695
rect 655 7665 660 7695
rect 620 7660 660 7665
rect 620 7635 660 7640
rect 620 7605 625 7635
rect 625 7605 655 7635
rect 655 7605 660 7635
rect 620 7600 660 7605
rect 620 7570 660 7575
rect 620 7540 625 7570
rect 625 7540 655 7570
rect 655 7540 660 7570
rect 620 7535 660 7540
rect 620 7500 660 7505
rect 620 7470 625 7500
rect 625 7470 655 7500
rect 655 7470 660 7500
rect 620 7465 660 7470
rect 620 7430 660 7435
rect 620 7400 625 7430
rect 625 7400 655 7430
rect 655 7400 660 7430
rect 620 7395 660 7400
rect 620 7360 660 7365
rect 620 7330 625 7360
rect 625 7330 655 7360
rect 655 7330 660 7360
rect 620 7325 660 7330
rect 620 7295 660 7300
rect 620 7265 625 7295
rect 625 7265 655 7295
rect 655 7265 660 7295
rect 620 7260 660 7265
rect 620 7235 660 7240
rect 620 7205 625 7235
rect 625 7205 655 7235
rect 655 7205 660 7235
rect 620 7200 660 7205
rect 620 7170 660 7175
rect 620 7140 625 7170
rect 625 7140 655 7170
rect 655 7140 660 7170
rect 620 7135 660 7140
rect 620 7100 660 7105
rect 620 7070 625 7100
rect 625 7070 655 7100
rect 655 7070 660 7100
rect 620 7065 660 7070
rect 620 7030 660 7035
rect 620 7000 625 7030
rect 625 7000 655 7030
rect 655 7000 660 7030
rect 620 6995 660 7000
rect 620 6960 660 6965
rect 620 6930 625 6960
rect 625 6930 655 6960
rect 655 6930 660 6960
rect 620 6925 660 6930
rect 620 6895 660 6900
rect 620 6865 625 6895
rect 625 6865 655 6895
rect 655 6865 660 6895
rect 620 6860 660 6865
rect 620 6835 660 6840
rect 620 6805 625 6835
rect 625 6805 655 6835
rect 655 6805 660 6835
rect 620 6800 660 6805
rect 620 6770 660 6775
rect 620 6740 625 6770
rect 625 6740 655 6770
rect 655 6740 660 6770
rect 620 6735 660 6740
rect 620 6700 660 6705
rect 620 6670 625 6700
rect 625 6670 655 6700
rect 655 6670 660 6700
rect 620 6665 660 6670
rect 620 6630 660 6635
rect 620 6600 625 6630
rect 625 6600 655 6630
rect 655 6600 660 6630
rect 620 6595 660 6600
rect 620 6560 660 6565
rect 620 6530 625 6560
rect 625 6530 655 6560
rect 655 6530 660 6560
rect 620 6525 660 6530
rect 620 6495 660 6500
rect 620 6465 625 6495
rect 625 6465 655 6495
rect 655 6465 660 6495
rect 620 6460 660 6465
rect 970 9635 1010 9640
rect 970 9605 975 9635
rect 975 9605 1005 9635
rect 1005 9605 1010 9635
rect 970 9600 1010 9605
rect 970 9570 1010 9575
rect 970 9540 975 9570
rect 975 9540 1005 9570
rect 1005 9540 1010 9570
rect 970 9535 1010 9540
rect 970 9500 1010 9505
rect 970 9470 975 9500
rect 975 9470 1005 9500
rect 1005 9470 1010 9500
rect 970 9465 1010 9470
rect 970 9430 1010 9435
rect 970 9400 975 9430
rect 975 9400 1005 9430
rect 1005 9400 1010 9430
rect 970 9395 1010 9400
rect 970 9360 1010 9365
rect 970 9330 975 9360
rect 975 9330 1005 9360
rect 1005 9330 1010 9360
rect 970 9325 1010 9330
rect 970 9295 1010 9300
rect 970 9265 975 9295
rect 975 9265 1005 9295
rect 1005 9265 1010 9295
rect 970 9260 1010 9265
rect 970 9235 1010 9240
rect 970 9205 975 9235
rect 975 9205 1005 9235
rect 1005 9205 1010 9235
rect 970 9200 1010 9205
rect 970 9170 1010 9175
rect 970 9140 975 9170
rect 975 9140 1005 9170
rect 1005 9140 1010 9170
rect 970 9135 1010 9140
rect 970 9100 1010 9105
rect 970 9070 975 9100
rect 975 9070 1005 9100
rect 1005 9070 1010 9100
rect 970 9065 1010 9070
rect 970 9030 1010 9035
rect 970 9000 975 9030
rect 975 9000 1005 9030
rect 1005 9000 1010 9030
rect 970 8995 1010 9000
rect 970 8960 1010 8965
rect 970 8930 975 8960
rect 975 8930 1005 8960
rect 1005 8930 1010 8960
rect 970 8925 1010 8930
rect 970 8895 1010 8900
rect 970 8865 975 8895
rect 975 8865 1005 8895
rect 1005 8865 1010 8895
rect 970 8860 1010 8865
rect 970 8835 1010 8840
rect 970 8805 975 8835
rect 975 8805 1005 8835
rect 1005 8805 1010 8835
rect 970 8800 1010 8805
rect 970 8770 1010 8775
rect 970 8740 975 8770
rect 975 8740 1005 8770
rect 1005 8740 1010 8770
rect 970 8735 1010 8740
rect 970 8700 1010 8705
rect 970 8670 975 8700
rect 975 8670 1005 8700
rect 1005 8670 1010 8700
rect 970 8665 1010 8670
rect 970 8630 1010 8635
rect 970 8600 975 8630
rect 975 8600 1005 8630
rect 1005 8600 1010 8630
rect 970 8595 1010 8600
rect 970 8560 1010 8565
rect 970 8530 975 8560
rect 975 8530 1005 8560
rect 1005 8530 1010 8560
rect 970 8525 1010 8530
rect 970 8495 1010 8500
rect 970 8465 975 8495
rect 975 8465 1005 8495
rect 1005 8465 1010 8495
rect 970 8460 1010 8465
rect 970 8435 1010 8440
rect 970 8405 975 8435
rect 975 8405 1005 8435
rect 1005 8405 1010 8435
rect 970 8400 1010 8405
rect 970 8370 1010 8375
rect 970 8340 975 8370
rect 975 8340 1005 8370
rect 1005 8340 1010 8370
rect 970 8335 1010 8340
rect 970 8300 1010 8305
rect 970 8270 975 8300
rect 975 8270 1005 8300
rect 1005 8270 1010 8300
rect 970 8265 1010 8270
rect 970 8230 1010 8235
rect 970 8200 975 8230
rect 975 8200 1005 8230
rect 1005 8200 1010 8230
rect 970 8195 1010 8200
rect 970 8160 1010 8165
rect 970 8130 975 8160
rect 975 8130 1005 8160
rect 1005 8130 1010 8160
rect 970 8125 1010 8130
rect 970 8095 1010 8100
rect 970 8065 975 8095
rect 975 8065 1005 8095
rect 1005 8065 1010 8095
rect 970 8060 1010 8065
rect 970 8035 1010 8040
rect 970 8005 975 8035
rect 975 8005 1005 8035
rect 1005 8005 1010 8035
rect 970 8000 1010 8005
rect 970 7970 1010 7975
rect 970 7940 975 7970
rect 975 7940 1005 7970
rect 1005 7940 1010 7970
rect 970 7935 1010 7940
rect 970 7900 1010 7905
rect 970 7870 975 7900
rect 975 7870 1005 7900
rect 1005 7870 1010 7900
rect 970 7865 1010 7870
rect 970 7830 1010 7835
rect 970 7800 975 7830
rect 975 7800 1005 7830
rect 1005 7800 1010 7830
rect 970 7795 1010 7800
rect 970 7760 1010 7765
rect 970 7730 975 7760
rect 975 7730 1005 7760
rect 1005 7730 1010 7760
rect 970 7725 1010 7730
rect 970 7695 1010 7700
rect 970 7665 975 7695
rect 975 7665 1005 7695
rect 1005 7665 1010 7695
rect 970 7660 1010 7665
rect 970 7635 1010 7640
rect 970 7605 975 7635
rect 975 7605 1005 7635
rect 1005 7605 1010 7635
rect 970 7600 1010 7605
rect 970 7570 1010 7575
rect 970 7540 975 7570
rect 975 7540 1005 7570
rect 1005 7540 1010 7570
rect 970 7535 1010 7540
rect 970 7500 1010 7505
rect 970 7470 975 7500
rect 975 7470 1005 7500
rect 1005 7470 1010 7500
rect 970 7465 1010 7470
rect 970 7430 1010 7435
rect 970 7400 975 7430
rect 975 7400 1005 7430
rect 1005 7400 1010 7430
rect 970 7395 1010 7400
rect 970 7360 1010 7365
rect 970 7330 975 7360
rect 975 7330 1005 7360
rect 1005 7330 1010 7360
rect 970 7325 1010 7330
rect 970 7295 1010 7300
rect 970 7265 975 7295
rect 975 7265 1005 7295
rect 1005 7265 1010 7295
rect 970 7260 1010 7265
rect 970 7235 1010 7240
rect 970 7205 975 7235
rect 975 7205 1005 7235
rect 1005 7205 1010 7235
rect 970 7200 1010 7205
rect 970 7170 1010 7175
rect 970 7140 975 7170
rect 975 7140 1005 7170
rect 1005 7140 1010 7170
rect 970 7135 1010 7140
rect 970 7100 1010 7105
rect 970 7070 975 7100
rect 975 7070 1005 7100
rect 1005 7070 1010 7100
rect 970 7065 1010 7070
rect 970 7030 1010 7035
rect 970 7000 975 7030
rect 975 7000 1005 7030
rect 1005 7000 1010 7030
rect 970 6995 1010 7000
rect 970 6960 1010 6965
rect 970 6930 975 6960
rect 975 6930 1005 6960
rect 1005 6930 1010 6960
rect 970 6925 1010 6930
rect 970 6895 1010 6900
rect 970 6865 975 6895
rect 975 6865 1005 6895
rect 1005 6865 1010 6895
rect 970 6860 1010 6865
rect 970 6835 1010 6840
rect 970 6805 975 6835
rect 975 6805 1005 6835
rect 1005 6805 1010 6835
rect 970 6800 1010 6805
rect 970 6770 1010 6775
rect 970 6740 975 6770
rect 975 6740 1005 6770
rect 1005 6740 1010 6770
rect 970 6735 1010 6740
rect 970 6700 1010 6705
rect 970 6670 975 6700
rect 975 6670 1005 6700
rect 1005 6670 1010 6700
rect 970 6665 1010 6670
rect 970 6630 1010 6635
rect 970 6600 975 6630
rect 975 6600 1005 6630
rect 1005 6600 1010 6630
rect 970 6595 1010 6600
rect 970 6560 1010 6565
rect 970 6530 975 6560
rect 975 6530 1005 6560
rect 1005 6530 1010 6560
rect 970 6525 1010 6530
rect 970 6495 1010 6500
rect 970 6465 975 6495
rect 975 6465 1005 6495
rect 1005 6465 1010 6495
rect 970 6460 1010 6465
rect 1670 9635 1710 9640
rect 1670 9605 1675 9635
rect 1675 9605 1705 9635
rect 1705 9605 1710 9635
rect 1670 9600 1710 9605
rect 1670 9570 1710 9575
rect 1670 9540 1675 9570
rect 1675 9540 1705 9570
rect 1705 9540 1710 9570
rect 1670 9535 1710 9540
rect 1670 9500 1710 9505
rect 1670 9470 1675 9500
rect 1675 9470 1705 9500
rect 1705 9470 1710 9500
rect 1670 9465 1710 9470
rect 1670 9430 1710 9435
rect 1670 9400 1675 9430
rect 1675 9400 1705 9430
rect 1705 9400 1710 9430
rect 1670 9395 1710 9400
rect 1670 9360 1710 9365
rect 1670 9330 1675 9360
rect 1675 9330 1705 9360
rect 1705 9330 1710 9360
rect 1670 9325 1710 9330
rect 1670 9295 1710 9300
rect 1670 9265 1675 9295
rect 1675 9265 1705 9295
rect 1705 9265 1710 9295
rect 1670 9260 1710 9265
rect 1670 9235 1710 9240
rect 1670 9205 1675 9235
rect 1675 9205 1705 9235
rect 1705 9205 1710 9235
rect 1670 9200 1710 9205
rect 1670 9170 1710 9175
rect 1670 9140 1675 9170
rect 1675 9140 1705 9170
rect 1705 9140 1710 9170
rect 1670 9135 1710 9140
rect 1670 9100 1710 9105
rect 1670 9070 1675 9100
rect 1675 9070 1705 9100
rect 1705 9070 1710 9100
rect 1670 9065 1710 9070
rect 1670 9030 1710 9035
rect 1670 9000 1675 9030
rect 1675 9000 1705 9030
rect 1705 9000 1710 9030
rect 1670 8995 1710 9000
rect 1670 8960 1710 8965
rect 1670 8930 1675 8960
rect 1675 8930 1705 8960
rect 1705 8930 1710 8960
rect 1670 8925 1710 8930
rect 1670 8895 1710 8900
rect 1670 8865 1675 8895
rect 1675 8865 1705 8895
rect 1705 8865 1710 8895
rect 1670 8860 1710 8865
rect 1670 8835 1710 8840
rect 1670 8805 1675 8835
rect 1675 8805 1705 8835
rect 1705 8805 1710 8835
rect 1670 8800 1710 8805
rect 1670 8770 1710 8775
rect 1670 8740 1675 8770
rect 1675 8740 1705 8770
rect 1705 8740 1710 8770
rect 1670 8735 1710 8740
rect 1670 8700 1710 8705
rect 1670 8670 1675 8700
rect 1675 8670 1705 8700
rect 1705 8670 1710 8700
rect 1670 8665 1710 8670
rect 1670 8630 1710 8635
rect 1670 8600 1675 8630
rect 1675 8600 1705 8630
rect 1705 8600 1710 8630
rect 1670 8595 1710 8600
rect 1670 8560 1710 8565
rect 1670 8530 1675 8560
rect 1675 8530 1705 8560
rect 1705 8530 1710 8560
rect 1670 8525 1710 8530
rect 1670 8495 1710 8500
rect 1670 8465 1675 8495
rect 1675 8465 1705 8495
rect 1705 8465 1710 8495
rect 1670 8460 1710 8465
rect 1670 8435 1710 8440
rect 1670 8405 1675 8435
rect 1675 8405 1705 8435
rect 1705 8405 1710 8435
rect 1670 8400 1710 8405
rect 1670 8370 1710 8375
rect 1670 8340 1675 8370
rect 1675 8340 1705 8370
rect 1705 8340 1710 8370
rect 1670 8335 1710 8340
rect 1670 8300 1710 8305
rect 1670 8270 1675 8300
rect 1675 8270 1705 8300
rect 1705 8270 1710 8300
rect 1670 8265 1710 8270
rect 1670 8230 1710 8235
rect 1670 8200 1675 8230
rect 1675 8200 1705 8230
rect 1705 8200 1710 8230
rect 1670 8195 1710 8200
rect 1670 8160 1710 8165
rect 1670 8130 1675 8160
rect 1675 8130 1705 8160
rect 1705 8130 1710 8160
rect 1670 8125 1710 8130
rect 1670 8095 1710 8100
rect 1670 8065 1675 8095
rect 1675 8065 1705 8095
rect 1705 8065 1710 8095
rect 1670 8060 1710 8065
rect 1670 8035 1710 8040
rect 1670 8005 1675 8035
rect 1675 8005 1705 8035
rect 1705 8005 1710 8035
rect 1670 8000 1710 8005
rect 1670 7970 1710 7975
rect 1670 7940 1675 7970
rect 1675 7940 1705 7970
rect 1705 7940 1710 7970
rect 1670 7935 1710 7940
rect 1670 7900 1710 7905
rect 1670 7870 1675 7900
rect 1675 7870 1705 7900
rect 1705 7870 1710 7900
rect 1670 7865 1710 7870
rect 1670 7830 1710 7835
rect 1670 7800 1675 7830
rect 1675 7800 1705 7830
rect 1705 7800 1710 7830
rect 1670 7795 1710 7800
rect 1670 7760 1710 7765
rect 1670 7730 1675 7760
rect 1675 7730 1705 7760
rect 1705 7730 1710 7760
rect 1670 7725 1710 7730
rect 1670 7695 1710 7700
rect 1670 7665 1675 7695
rect 1675 7665 1705 7695
rect 1705 7665 1710 7695
rect 1670 7660 1710 7665
rect 1670 7635 1710 7640
rect 1670 7605 1675 7635
rect 1675 7605 1705 7635
rect 1705 7605 1710 7635
rect 1670 7600 1710 7605
rect 1670 7570 1710 7575
rect 1670 7540 1675 7570
rect 1675 7540 1705 7570
rect 1705 7540 1710 7570
rect 1670 7535 1710 7540
rect 1670 7500 1710 7505
rect 1670 7470 1675 7500
rect 1675 7470 1705 7500
rect 1705 7470 1710 7500
rect 1670 7465 1710 7470
rect 1670 7430 1710 7435
rect 1670 7400 1675 7430
rect 1675 7400 1705 7430
rect 1705 7400 1710 7430
rect 1670 7395 1710 7400
rect 1670 7360 1710 7365
rect 1670 7330 1675 7360
rect 1675 7330 1705 7360
rect 1705 7330 1710 7360
rect 1670 7325 1710 7330
rect 1670 7295 1710 7300
rect 1670 7265 1675 7295
rect 1675 7265 1705 7295
rect 1705 7265 1710 7295
rect 1670 7260 1710 7265
rect 1670 7235 1710 7240
rect 1670 7205 1675 7235
rect 1675 7205 1705 7235
rect 1705 7205 1710 7235
rect 1670 7200 1710 7205
rect 1670 7170 1710 7175
rect 1670 7140 1675 7170
rect 1675 7140 1705 7170
rect 1705 7140 1710 7170
rect 1670 7135 1710 7140
rect 1670 7100 1710 7105
rect 1670 7070 1675 7100
rect 1675 7070 1705 7100
rect 1705 7070 1710 7100
rect 1670 7065 1710 7070
rect 1670 7030 1710 7035
rect 1670 7000 1675 7030
rect 1675 7000 1705 7030
rect 1705 7000 1710 7030
rect 1670 6995 1710 7000
rect 1670 6960 1710 6965
rect 1670 6930 1675 6960
rect 1675 6930 1705 6960
rect 1705 6930 1710 6960
rect 1670 6925 1710 6930
rect 1670 6895 1710 6900
rect 1670 6865 1675 6895
rect 1675 6865 1705 6895
rect 1705 6865 1710 6895
rect 1670 6860 1710 6865
rect 1670 6835 1710 6840
rect 1670 6805 1675 6835
rect 1675 6805 1705 6835
rect 1705 6805 1710 6835
rect 1670 6800 1710 6805
rect 1670 6770 1710 6775
rect 1670 6740 1675 6770
rect 1675 6740 1705 6770
rect 1705 6740 1710 6770
rect 1670 6735 1710 6740
rect 1670 6700 1710 6705
rect 1670 6670 1675 6700
rect 1675 6670 1705 6700
rect 1705 6670 1710 6700
rect 1670 6665 1710 6670
rect 1670 6630 1710 6635
rect 1670 6600 1675 6630
rect 1675 6600 1705 6630
rect 1705 6600 1710 6630
rect 1670 6595 1710 6600
rect 1670 6560 1710 6565
rect 1670 6530 1675 6560
rect 1675 6530 1705 6560
rect 1705 6530 1710 6560
rect 1670 6525 1710 6530
rect 1670 6495 1710 6500
rect 1670 6465 1675 6495
rect 1675 6465 1705 6495
rect 1705 6465 1710 6495
rect 1670 6460 1710 6465
rect 2245 9635 2285 9640
rect 2245 9605 2250 9635
rect 2250 9605 2280 9635
rect 2280 9605 2285 9635
rect 2245 9600 2285 9605
rect 2245 9570 2285 9575
rect 2245 9540 2250 9570
rect 2250 9540 2280 9570
rect 2280 9540 2285 9570
rect 2245 9535 2285 9540
rect 2245 9500 2285 9505
rect 2245 9470 2250 9500
rect 2250 9470 2280 9500
rect 2280 9470 2285 9500
rect 2245 9465 2285 9470
rect 2245 9430 2285 9435
rect 2245 9400 2250 9430
rect 2250 9400 2280 9430
rect 2280 9400 2285 9430
rect 2245 9395 2285 9400
rect 2245 9360 2285 9365
rect 2245 9330 2250 9360
rect 2250 9330 2280 9360
rect 2280 9330 2285 9360
rect 2245 9325 2285 9330
rect 2245 9295 2285 9300
rect 2245 9265 2250 9295
rect 2250 9265 2280 9295
rect 2280 9265 2285 9295
rect 2245 9260 2285 9265
rect 2245 9235 2285 9240
rect 2245 9205 2250 9235
rect 2250 9205 2280 9235
rect 2280 9205 2285 9235
rect 2245 9200 2285 9205
rect 2245 9170 2285 9175
rect 2245 9140 2250 9170
rect 2250 9140 2280 9170
rect 2280 9140 2285 9170
rect 2245 9135 2285 9140
rect 2245 9100 2285 9105
rect 2245 9070 2250 9100
rect 2250 9070 2280 9100
rect 2280 9070 2285 9100
rect 2245 9065 2285 9070
rect 2245 9030 2285 9035
rect 2245 9000 2250 9030
rect 2250 9000 2280 9030
rect 2280 9000 2285 9030
rect 2245 8995 2285 9000
rect 2245 8960 2285 8965
rect 2245 8930 2250 8960
rect 2250 8930 2280 8960
rect 2280 8930 2285 8960
rect 2245 8925 2285 8930
rect 2245 8895 2285 8900
rect 2245 8865 2250 8895
rect 2250 8865 2280 8895
rect 2280 8865 2285 8895
rect 2245 8860 2285 8865
rect 2245 8835 2285 8840
rect 2245 8805 2250 8835
rect 2250 8805 2280 8835
rect 2280 8805 2285 8835
rect 2245 8800 2285 8805
rect 2245 8770 2285 8775
rect 2245 8740 2250 8770
rect 2250 8740 2280 8770
rect 2280 8740 2285 8770
rect 2245 8735 2285 8740
rect 2245 8700 2285 8705
rect 2245 8670 2250 8700
rect 2250 8670 2280 8700
rect 2280 8670 2285 8700
rect 2245 8665 2285 8670
rect 2245 8630 2285 8635
rect 2245 8600 2250 8630
rect 2250 8600 2280 8630
rect 2280 8600 2285 8630
rect 2245 8595 2285 8600
rect 2245 8560 2285 8565
rect 2245 8530 2250 8560
rect 2250 8530 2280 8560
rect 2280 8530 2285 8560
rect 2245 8525 2285 8530
rect 2245 8495 2285 8500
rect 2245 8465 2250 8495
rect 2250 8465 2280 8495
rect 2280 8465 2285 8495
rect 2245 8460 2285 8465
rect 2245 8435 2285 8440
rect 2245 8405 2250 8435
rect 2250 8405 2280 8435
rect 2280 8405 2285 8435
rect 2245 8400 2285 8405
rect 2245 8370 2285 8375
rect 2245 8340 2250 8370
rect 2250 8340 2280 8370
rect 2280 8340 2285 8370
rect 2245 8335 2285 8340
rect 2245 8300 2285 8305
rect 2245 8270 2250 8300
rect 2250 8270 2280 8300
rect 2280 8270 2285 8300
rect 2245 8265 2285 8270
rect 2245 8230 2285 8235
rect 2245 8200 2250 8230
rect 2250 8200 2280 8230
rect 2280 8200 2285 8230
rect 2245 8195 2285 8200
rect 2245 8160 2285 8165
rect 2245 8130 2250 8160
rect 2250 8130 2280 8160
rect 2280 8130 2285 8160
rect 2245 8125 2285 8130
rect 2245 8095 2285 8100
rect 2245 8065 2250 8095
rect 2250 8065 2280 8095
rect 2280 8065 2285 8095
rect 2245 8060 2285 8065
rect 2245 8035 2285 8040
rect 2245 8005 2250 8035
rect 2250 8005 2280 8035
rect 2280 8005 2285 8035
rect 2245 8000 2285 8005
rect 2245 7970 2285 7975
rect 2245 7940 2250 7970
rect 2250 7940 2280 7970
rect 2280 7940 2285 7970
rect 2245 7935 2285 7940
rect 2245 7900 2285 7905
rect 2245 7870 2250 7900
rect 2250 7870 2280 7900
rect 2280 7870 2285 7900
rect 2245 7865 2285 7870
rect 2245 7830 2285 7835
rect 2245 7800 2250 7830
rect 2250 7800 2280 7830
rect 2280 7800 2285 7830
rect 2245 7795 2285 7800
rect 2245 7760 2285 7765
rect 2245 7730 2250 7760
rect 2250 7730 2280 7760
rect 2280 7730 2285 7760
rect 2245 7725 2285 7730
rect 2245 7695 2285 7700
rect 2245 7665 2250 7695
rect 2250 7665 2280 7695
rect 2280 7665 2285 7695
rect 2245 7660 2285 7665
rect 2245 7635 2285 7640
rect 2245 7605 2250 7635
rect 2250 7605 2280 7635
rect 2280 7605 2285 7635
rect 2245 7600 2285 7605
rect 2245 7570 2285 7575
rect 2245 7540 2250 7570
rect 2250 7540 2280 7570
rect 2280 7540 2285 7570
rect 2245 7535 2285 7540
rect 2245 7500 2285 7505
rect 2245 7470 2250 7500
rect 2250 7470 2280 7500
rect 2280 7470 2285 7500
rect 2245 7465 2285 7470
rect 2245 7430 2285 7435
rect 2245 7400 2250 7430
rect 2250 7400 2280 7430
rect 2280 7400 2285 7430
rect 2245 7395 2285 7400
rect 2245 7360 2285 7365
rect 2245 7330 2250 7360
rect 2250 7330 2280 7360
rect 2280 7330 2285 7360
rect 2245 7325 2285 7330
rect 2245 7295 2285 7300
rect 2245 7265 2250 7295
rect 2250 7265 2280 7295
rect 2280 7265 2285 7295
rect 2245 7260 2285 7265
rect 2245 7235 2285 7240
rect 2245 7205 2250 7235
rect 2250 7205 2280 7235
rect 2280 7205 2285 7235
rect 2245 7200 2285 7205
rect 2245 7170 2285 7175
rect 2245 7140 2250 7170
rect 2250 7140 2280 7170
rect 2280 7140 2285 7170
rect 2245 7135 2285 7140
rect 2245 7100 2285 7105
rect 2245 7070 2250 7100
rect 2250 7070 2280 7100
rect 2280 7070 2285 7100
rect 2245 7065 2285 7070
rect 2245 7030 2285 7035
rect 2245 7000 2250 7030
rect 2250 7000 2280 7030
rect 2280 7000 2285 7030
rect 2245 6995 2285 7000
rect 2245 6960 2285 6965
rect 2245 6930 2250 6960
rect 2250 6930 2280 6960
rect 2280 6930 2285 6960
rect 2245 6925 2285 6930
rect 2245 6895 2285 6900
rect 2245 6865 2250 6895
rect 2250 6865 2280 6895
rect 2280 6865 2285 6895
rect 2245 6860 2285 6865
rect 2245 6835 2285 6840
rect 2245 6805 2250 6835
rect 2250 6805 2280 6835
rect 2280 6805 2285 6835
rect 2245 6800 2285 6805
rect 2245 6770 2285 6775
rect 2245 6740 2250 6770
rect 2250 6740 2280 6770
rect 2280 6740 2285 6770
rect 2245 6735 2285 6740
rect 2245 6700 2285 6705
rect 2245 6670 2250 6700
rect 2250 6670 2280 6700
rect 2280 6670 2285 6700
rect 2245 6665 2285 6670
rect 2245 6630 2285 6635
rect 2245 6600 2250 6630
rect 2250 6600 2280 6630
rect 2280 6600 2285 6630
rect 2245 6595 2285 6600
rect 2245 6560 2285 6565
rect 2245 6530 2250 6560
rect 2250 6530 2280 6560
rect 2280 6530 2285 6560
rect 2245 6525 2285 6530
rect 2245 6495 2285 6500
rect 2245 6465 2250 6495
rect 2250 6465 2280 6495
rect 2280 6465 2285 6495
rect 2245 6460 2285 6465
rect 3175 9635 3215 9640
rect 3175 9605 3180 9635
rect 3180 9605 3210 9635
rect 3210 9605 3215 9635
rect 3175 9600 3215 9605
rect 3235 9635 3275 9640
rect 3235 9605 3240 9635
rect 3240 9605 3270 9635
rect 3270 9605 3275 9635
rect 3235 9600 3275 9605
rect 3175 9570 3215 9575
rect 3175 9540 3180 9570
rect 3180 9540 3210 9570
rect 3210 9540 3215 9570
rect 3175 9535 3215 9540
rect 3235 9570 3275 9575
rect 3235 9540 3240 9570
rect 3240 9540 3270 9570
rect 3270 9540 3275 9570
rect 3235 9535 3275 9540
rect 3175 9500 3215 9505
rect 3175 9470 3180 9500
rect 3180 9470 3210 9500
rect 3210 9470 3215 9500
rect 3175 9465 3215 9470
rect 3235 9500 3275 9505
rect 3235 9470 3240 9500
rect 3240 9470 3270 9500
rect 3270 9470 3275 9500
rect 3235 9465 3275 9470
rect 3175 9430 3215 9435
rect 3175 9400 3180 9430
rect 3180 9400 3210 9430
rect 3210 9400 3215 9430
rect 3175 9395 3215 9400
rect 3235 9430 3275 9435
rect 3235 9400 3240 9430
rect 3240 9400 3270 9430
rect 3270 9400 3275 9430
rect 3235 9395 3275 9400
rect 3175 9360 3215 9365
rect 3175 9330 3180 9360
rect 3180 9330 3210 9360
rect 3210 9330 3215 9360
rect 3175 9325 3215 9330
rect 3235 9360 3275 9365
rect 3235 9330 3240 9360
rect 3240 9330 3270 9360
rect 3270 9330 3275 9360
rect 3235 9325 3275 9330
rect 3175 9295 3215 9300
rect 3175 9265 3180 9295
rect 3180 9265 3210 9295
rect 3210 9265 3215 9295
rect 3175 9260 3215 9265
rect 3235 9295 3275 9300
rect 3235 9265 3240 9295
rect 3240 9265 3270 9295
rect 3270 9265 3275 9295
rect 3235 9260 3275 9265
rect 3175 9235 3215 9240
rect 3175 9205 3180 9235
rect 3180 9205 3210 9235
rect 3210 9205 3215 9235
rect 3175 9200 3215 9205
rect 3235 9235 3275 9240
rect 3235 9205 3240 9235
rect 3240 9205 3270 9235
rect 3270 9205 3275 9235
rect 3235 9200 3275 9205
rect 3175 9170 3215 9175
rect 3175 9140 3180 9170
rect 3180 9140 3210 9170
rect 3210 9140 3215 9170
rect 3175 9135 3215 9140
rect 3235 9170 3275 9175
rect 3235 9140 3240 9170
rect 3240 9140 3270 9170
rect 3270 9140 3275 9170
rect 3235 9135 3275 9140
rect 3175 9100 3215 9105
rect 3175 9070 3180 9100
rect 3180 9070 3210 9100
rect 3210 9070 3215 9100
rect 3175 9065 3215 9070
rect 3235 9100 3275 9105
rect 3235 9070 3240 9100
rect 3240 9070 3270 9100
rect 3270 9070 3275 9100
rect 3235 9065 3275 9070
rect 3175 9030 3215 9035
rect 3175 9000 3180 9030
rect 3180 9000 3210 9030
rect 3210 9000 3215 9030
rect 3175 8995 3215 9000
rect 3235 9030 3275 9035
rect 3235 9000 3240 9030
rect 3240 9000 3270 9030
rect 3270 9000 3275 9030
rect 3235 8995 3275 9000
rect 3175 8960 3215 8965
rect 3175 8930 3180 8960
rect 3180 8930 3210 8960
rect 3210 8930 3215 8960
rect 3175 8925 3215 8930
rect 3235 8960 3275 8965
rect 3235 8930 3240 8960
rect 3240 8930 3270 8960
rect 3270 8930 3275 8960
rect 3235 8925 3275 8930
rect 3175 8895 3215 8900
rect 3175 8865 3180 8895
rect 3180 8865 3210 8895
rect 3210 8865 3215 8895
rect 3175 8860 3215 8865
rect 3235 8895 3275 8900
rect 3235 8865 3240 8895
rect 3240 8865 3270 8895
rect 3270 8865 3275 8895
rect 3235 8860 3275 8865
rect 3175 8835 3215 8840
rect 3175 8805 3180 8835
rect 3180 8805 3210 8835
rect 3210 8805 3215 8835
rect 3175 8800 3215 8805
rect 3235 8835 3275 8840
rect 3235 8805 3240 8835
rect 3240 8805 3270 8835
rect 3270 8805 3275 8835
rect 3235 8800 3275 8805
rect 3175 8770 3215 8775
rect 3175 8740 3180 8770
rect 3180 8740 3210 8770
rect 3210 8740 3215 8770
rect 3175 8735 3215 8740
rect 3235 8770 3275 8775
rect 3235 8740 3240 8770
rect 3240 8740 3270 8770
rect 3270 8740 3275 8770
rect 3235 8735 3275 8740
rect 3175 8700 3215 8705
rect 3175 8670 3180 8700
rect 3180 8670 3210 8700
rect 3210 8670 3215 8700
rect 3175 8665 3215 8670
rect 3235 8700 3275 8705
rect 3235 8670 3240 8700
rect 3240 8670 3270 8700
rect 3270 8670 3275 8700
rect 3235 8665 3275 8670
rect 3175 8630 3215 8635
rect 3175 8600 3180 8630
rect 3180 8600 3210 8630
rect 3210 8600 3215 8630
rect 3175 8595 3215 8600
rect 3235 8630 3275 8635
rect 3235 8600 3240 8630
rect 3240 8600 3270 8630
rect 3270 8600 3275 8630
rect 3235 8595 3275 8600
rect 3175 8560 3215 8565
rect 3175 8530 3180 8560
rect 3180 8530 3210 8560
rect 3210 8530 3215 8560
rect 3175 8525 3215 8530
rect 3235 8560 3275 8565
rect 3235 8530 3240 8560
rect 3240 8530 3270 8560
rect 3270 8530 3275 8560
rect 3235 8525 3275 8530
rect 3175 8495 3215 8500
rect 3175 8465 3180 8495
rect 3180 8465 3210 8495
rect 3210 8465 3215 8495
rect 3175 8460 3215 8465
rect 3235 8495 3275 8500
rect 3235 8465 3240 8495
rect 3240 8465 3270 8495
rect 3270 8465 3275 8495
rect 3235 8460 3275 8465
rect 3175 8435 3215 8440
rect 3175 8405 3180 8435
rect 3180 8405 3210 8435
rect 3210 8405 3215 8435
rect 3175 8400 3215 8405
rect 3235 8435 3275 8440
rect 3235 8405 3240 8435
rect 3240 8405 3270 8435
rect 3270 8405 3275 8435
rect 3235 8400 3275 8405
rect 3175 8370 3215 8375
rect 3175 8340 3180 8370
rect 3180 8340 3210 8370
rect 3210 8340 3215 8370
rect 3175 8335 3215 8340
rect 3235 8370 3275 8375
rect 3235 8340 3240 8370
rect 3240 8340 3270 8370
rect 3270 8340 3275 8370
rect 3235 8335 3275 8340
rect 3175 8300 3215 8305
rect 3175 8270 3180 8300
rect 3180 8270 3210 8300
rect 3210 8270 3215 8300
rect 3175 8265 3215 8270
rect 3235 8300 3275 8305
rect 3235 8270 3240 8300
rect 3240 8270 3270 8300
rect 3270 8270 3275 8300
rect 3235 8265 3275 8270
rect 3175 8230 3215 8235
rect 3175 8200 3180 8230
rect 3180 8200 3210 8230
rect 3210 8200 3215 8230
rect 3175 8195 3215 8200
rect 3235 8230 3275 8235
rect 3235 8200 3240 8230
rect 3240 8200 3270 8230
rect 3270 8200 3275 8230
rect 3235 8195 3275 8200
rect 3175 8160 3215 8165
rect 3175 8130 3180 8160
rect 3180 8130 3210 8160
rect 3210 8130 3215 8160
rect 3175 8125 3215 8130
rect 3235 8160 3275 8165
rect 3235 8130 3240 8160
rect 3240 8130 3270 8160
rect 3270 8130 3275 8160
rect 3235 8125 3275 8130
rect 3175 8095 3215 8100
rect 3175 8065 3180 8095
rect 3180 8065 3210 8095
rect 3210 8065 3215 8095
rect 3175 8060 3215 8065
rect 3235 8095 3275 8100
rect 3235 8065 3240 8095
rect 3240 8065 3270 8095
rect 3270 8065 3275 8095
rect 3235 8060 3275 8065
rect 3175 8035 3215 8040
rect 3175 8005 3180 8035
rect 3180 8005 3210 8035
rect 3210 8005 3215 8035
rect 3175 8000 3215 8005
rect 3235 8035 3275 8040
rect 3235 8005 3240 8035
rect 3240 8005 3270 8035
rect 3270 8005 3275 8035
rect 3235 8000 3275 8005
rect 3175 7970 3215 7975
rect 3175 7940 3180 7970
rect 3180 7940 3210 7970
rect 3210 7940 3215 7970
rect 3175 7935 3215 7940
rect 3235 7970 3275 7975
rect 3235 7940 3240 7970
rect 3240 7940 3270 7970
rect 3270 7940 3275 7970
rect 3235 7935 3275 7940
rect 3175 7900 3215 7905
rect 3175 7870 3180 7900
rect 3180 7870 3210 7900
rect 3210 7870 3215 7900
rect 3175 7865 3215 7870
rect 3235 7900 3275 7905
rect 3235 7870 3240 7900
rect 3240 7870 3270 7900
rect 3270 7870 3275 7900
rect 3235 7865 3275 7870
rect 3175 7830 3215 7835
rect 3175 7800 3180 7830
rect 3180 7800 3210 7830
rect 3210 7800 3215 7830
rect 3175 7795 3215 7800
rect 3235 7830 3275 7835
rect 3235 7800 3240 7830
rect 3240 7800 3270 7830
rect 3270 7800 3275 7830
rect 3235 7795 3275 7800
rect 3175 7760 3215 7765
rect 3175 7730 3180 7760
rect 3180 7730 3210 7760
rect 3210 7730 3215 7760
rect 3175 7725 3215 7730
rect 3235 7760 3275 7765
rect 3235 7730 3240 7760
rect 3240 7730 3270 7760
rect 3270 7730 3275 7760
rect 3235 7725 3275 7730
rect 3175 7695 3215 7700
rect 3175 7665 3180 7695
rect 3180 7665 3210 7695
rect 3210 7665 3215 7695
rect 3175 7660 3215 7665
rect 3235 7695 3275 7700
rect 3235 7665 3240 7695
rect 3240 7665 3270 7695
rect 3270 7665 3275 7695
rect 3235 7660 3275 7665
rect 3175 7635 3215 7640
rect 3175 7605 3180 7635
rect 3180 7605 3210 7635
rect 3210 7605 3215 7635
rect 3175 7600 3215 7605
rect 3235 7635 3275 7640
rect 3235 7605 3240 7635
rect 3240 7605 3270 7635
rect 3270 7605 3275 7635
rect 3235 7600 3275 7605
rect 3175 7570 3215 7575
rect 3175 7540 3180 7570
rect 3180 7540 3210 7570
rect 3210 7540 3215 7570
rect 3175 7535 3215 7540
rect 3235 7570 3275 7575
rect 3235 7540 3240 7570
rect 3240 7540 3270 7570
rect 3270 7540 3275 7570
rect 3235 7535 3275 7540
rect 3175 7500 3215 7505
rect 3175 7470 3180 7500
rect 3180 7470 3210 7500
rect 3210 7470 3215 7500
rect 3175 7465 3215 7470
rect 3235 7500 3275 7505
rect 3235 7470 3240 7500
rect 3240 7470 3270 7500
rect 3270 7470 3275 7500
rect 3235 7465 3275 7470
rect 3175 7430 3215 7435
rect 3175 7400 3180 7430
rect 3180 7400 3210 7430
rect 3210 7400 3215 7430
rect 3175 7395 3215 7400
rect 3235 7430 3275 7435
rect 3235 7400 3240 7430
rect 3240 7400 3270 7430
rect 3270 7400 3275 7430
rect 3235 7395 3275 7400
rect 3175 7360 3215 7365
rect 3175 7330 3180 7360
rect 3180 7330 3210 7360
rect 3210 7330 3215 7360
rect 3175 7325 3215 7330
rect 3235 7360 3275 7365
rect 3235 7330 3240 7360
rect 3240 7330 3270 7360
rect 3270 7330 3275 7360
rect 3235 7325 3275 7330
rect 3175 7295 3215 7300
rect 3175 7265 3180 7295
rect 3180 7265 3210 7295
rect 3210 7265 3215 7295
rect 3175 7260 3215 7265
rect 3235 7295 3275 7300
rect 3235 7265 3240 7295
rect 3240 7265 3270 7295
rect 3270 7265 3275 7295
rect 3235 7260 3275 7265
rect 3175 7235 3215 7240
rect 3175 7205 3180 7235
rect 3180 7205 3210 7235
rect 3210 7205 3215 7235
rect 3175 7200 3215 7205
rect 3235 7235 3275 7240
rect 3235 7205 3240 7235
rect 3240 7205 3270 7235
rect 3270 7205 3275 7235
rect 3235 7200 3275 7205
rect 3175 7170 3215 7175
rect 3175 7140 3180 7170
rect 3180 7140 3210 7170
rect 3210 7140 3215 7170
rect 3175 7135 3215 7140
rect 3235 7170 3275 7175
rect 3235 7140 3240 7170
rect 3240 7140 3270 7170
rect 3270 7140 3275 7170
rect 3235 7135 3275 7140
rect 3175 7100 3215 7105
rect 3175 7070 3180 7100
rect 3180 7070 3210 7100
rect 3210 7070 3215 7100
rect 3175 7065 3215 7070
rect 3235 7100 3275 7105
rect 3235 7070 3240 7100
rect 3240 7070 3270 7100
rect 3270 7070 3275 7100
rect 3235 7065 3275 7070
rect 3175 7030 3215 7035
rect 3175 7000 3180 7030
rect 3180 7000 3210 7030
rect 3210 7000 3215 7030
rect 3175 6995 3215 7000
rect 3235 7030 3275 7035
rect 3235 7000 3240 7030
rect 3240 7000 3270 7030
rect 3270 7000 3275 7030
rect 3235 6995 3275 7000
rect 3175 6960 3215 6965
rect 3175 6930 3180 6960
rect 3180 6930 3210 6960
rect 3210 6930 3215 6960
rect 3175 6925 3215 6930
rect 3235 6960 3275 6965
rect 3235 6930 3240 6960
rect 3240 6930 3270 6960
rect 3270 6930 3275 6960
rect 3235 6925 3275 6930
rect 3175 6895 3215 6900
rect 3175 6865 3180 6895
rect 3180 6865 3210 6895
rect 3210 6865 3215 6895
rect 3175 6860 3215 6865
rect 3235 6895 3275 6900
rect 3235 6865 3240 6895
rect 3240 6865 3270 6895
rect 3270 6865 3275 6895
rect 3235 6860 3275 6865
rect 3175 6835 3215 6840
rect 3175 6805 3180 6835
rect 3180 6805 3210 6835
rect 3210 6805 3215 6835
rect 3175 6800 3215 6805
rect 3235 6835 3275 6840
rect 3235 6805 3240 6835
rect 3240 6805 3270 6835
rect 3270 6805 3275 6835
rect 3235 6800 3275 6805
rect 3175 6770 3215 6775
rect 3175 6740 3180 6770
rect 3180 6740 3210 6770
rect 3210 6740 3215 6770
rect 3175 6735 3215 6740
rect 3235 6770 3275 6775
rect 3235 6740 3240 6770
rect 3240 6740 3270 6770
rect 3270 6740 3275 6770
rect 3235 6735 3275 6740
rect 3175 6700 3215 6705
rect 3175 6670 3180 6700
rect 3180 6670 3210 6700
rect 3210 6670 3215 6700
rect 3175 6665 3215 6670
rect 3235 6700 3275 6705
rect 3235 6670 3240 6700
rect 3240 6670 3270 6700
rect 3270 6670 3275 6700
rect 3235 6665 3275 6670
rect 3175 6630 3215 6635
rect 3175 6600 3180 6630
rect 3180 6600 3210 6630
rect 3210 6600 3215 6630
rect 3175 6595 3215 6600
rect 3235 6630 3275 6635
rect 3235 6600 3240 6630
rect 3240 6600 3270 6630
rect 3270 6600 3275 6630
rect 3235 6595 3275 6600
rect 3175 6560 3215 6565
rect 3175 6530 3180 6560
rect 3180 6530 3210 6560
rect 3210 6530 3215 6560
rect 3175 6525 3215 6530
rect 3235 6560 3275 6565
rect 3235 6530 3240 6560
rect 3240 6530 3270 6560
rect 3270 6530 3275 6560
rect 3235 6525 3275 6530
rect 3175 6495 3215 6500
rect 3175 6465 3180 6495
rect 3180 6465 3210 6495
rect 3210 6465 3215 6495
rect 3175 6460 3215 6465
rect 3235 6495 3275 6500
rect 3235 6465 3240 6495
rect 3240 6465 3270 6495
rect 3270 6465 3275 6495
rect 3235 6460 3275 6465
rect 3345 9635 3385 9640
rect 3345 9605 3350 9635
rect 3350 9605 3380 9635
rect 3380 9605 3385 9635
rect 3345 9600 3385 9605
rect 3345 9570 3385 9575
rect 3345 9540 3350 9570
rect 3350 9540 3380 9570
rect 3380 9540 3385 9570
rect 3345 9535 3385 9540
rect 3345 9500 3385 9505
rect 3345 9470 3350 9500
rect 3350 9470 3380 9500
rect 3380 9470 3385 9500
rect 3345 9465 3385 9470
rect 3345 9430 3385 9435
rect 3345 9400 3350 9430
rect 3350 9400 3380 9430
rect 3380 9400 3385 9430
rect 3345 9395 3385 9400
rect 3345 9360 3385 9365
rect 3345 9330 3350 9360
rect 3350 9330 3380 9360
rect 3380 9330 3385 9360
rect 3345 9325 3385 9330
rect 3345 9295 3385 9300
rect 3345 9265 3350 9295
rect 3350 9265 3380 9295
rect 3380 9265 3385 9295
rect 3345 9260 3385 9265
rect 3345 9235 3385 9240
rect 3345 9205 3350 9235
rect 3350 9205 3380 9235
rect 3380 9205 3385 9235
rect 3345 9200 3385 9205
rect 3345 9170 3385 9175
rect 3345 9140 3350 9170
rect 3350 9140 3380 9170
rect 3380 9140 3385 9170
rect 3345 9135 3385 9140
rect 3345 9100 3385 9105
rect 3345 9070 3350 9100
rect 3350 9070 3380 9100
rect 3380 9070 3385 9100
rect 3345 9065 3385 9070
rect 3345 9030 3385 9035
rect 3345 9000 3350 9030
rect 3350 9000 3380 9030
rect 3380 9000 3385 9030
rect 3345 8995 3385 9000
rect 3345 8960 3385 8965
rect 3345 8930 3350 8960
rect 3350 8930 3380 8960
rect 3380 8930 3385 8960
rect 3345 8925 3385 8930
rect 3345 8895 3385 8900
rect 3345 8865 3350 8895
rect 3350 8865 3380 8895
rect 3380 8865 3385 8895
rect 3345 8860 3385 8865
rect 3345 8835 3385 8840
rect 3345 8805 3350 8835
rect 3350 8805 3380 8835
rect 3380 8805 3385 8835
rect 3345 8800 3385 8805
rect 3345 8770 3385 8775
rect 3345 8740 3350 8770
rect 3350 8740 3380 8770
rect 3380 8740 3385 8770
rect 3345 8735 3385 8740
rect 3345 8700 3385 8705
rect 3345 8670 3350 8700
rect 3350 8670 3380 8700
rect 3380 8670 3385 8700
rect 3345 8665 3385 8670
rect 3345 8630 3385 8635
rect 3345 8600 3350 8630
rect 3350 8600 3380 8630
rect 3380 8600 3385 8630
rect 3345 8595 3385 8600
rect 3345 8560 3385 8565
rect 3345 8530 3350 8560
rect 3350 8530 3380 8560
rect 3380 8530 3385 8560
rect 3345 8525 3385 8530
rect 3345 8495 3385 8500
rect 3345 8465 3350 8495
rect 3350 8465 3380 8495
rect 3380 8465 3385 8495
rect 3345 8460 3385 8465
rect 3345 8435 3385 8440
rect 3345 8405 3350 8435
rect 3350 8405 3380 8435
rect 3380 8405 3385 8435
rect 3345 8400 3385 8405
rect 3345 8370 3385 8375
rect 3345 8340 3350 8370
rect 3350 8340 3380 8370
rect 3380 8340 3385 8370
rect 3345 8335 3385 8340
rect 3345 8300 3385 8305
rect 3345 8270 3350 8300
rect 3350 8270 3380 8300
rect 3380 8270 3385 8300
rect 3345 8265 3385 8270
rect 3345 8230 3385 8235
rect 3345 8200 3350 8230
rect 3350 8200 3380 8230
rect 3380 8200 3385 8230
rect 3345 8195 3385 8200
rect 3345 8160 3385 8165
rect 3345 8130 3350 8160
rect 3350 8130 3380 8160
rect 3380 8130 3385 8160
rect 3345 8125 3385 8130
rect 3345 8095 3385 8100
rect 3345 8065 3350 8095
rect 3350 8065 3380 8095
rect 3380 8065 3385 8095
rect 3345 8060 3385 8065
rect 3345 8035 3385 8040
rect 3345 8005 3350 8035
rect 3350 8005 3380 8035
rect 3380 8005 3385 8035
rect 3345 8000 3385 8005
rect 3345 7970 3385 7975
rect 3345 7940 3350 7970
rect 3350 7940 3380 7970
rect 3380 7940 3385 7970
rect 3345 7935 3385 7940
rect 3345 7900 3385 7905
rect 3345 7870 3350 7900
rect 3350 7870 3380 7900
rect 3380 7870 3385 7900
rect 3345 7865 3385 7870
rect 3345 7830 3385 7835
rect 3345 7800 3350 7830
rect 3350 7800 3380 7830
rect 3380 7800 3385 7830
rect 3345 7795 3385 7800
rect 3345 7760 3385 7765
rect 3345 7730 3350 7760
rect 3350 7730 3380 7760
rect 3380 7730 3385 7760
rect 3345 7725 3385 7730
rect 3345 7695 3385 7700
rect 3345 7665 3350 7695
rect 3350 7665 3380 7695
rect 3380 7665 3385 7695
rect 3345 7660 3385 7665
rect 3345 7635 3385 7640
rect 3345 7605 3350 7635
rect 3350 7605 3380 7635
rect 3380 7605 3385 7635
rect 3345 7600 3385 7605
rect 3345 7570 3385 7575
rect 3345 7540 3350 7570
rect 3350 7540 3380 7570
rect 3380 7540 3385 7570
rect 3345 7535 3385 7540
rect 3345 7500 3385 7505
rect 3345 7470 3350 7500
rect 3350 7470 3380 7500
rect 3380 7470 3385 7500
rect 3345 7465 3385 7470
rect 3345 7430 3385 7435
rect 3345 7400 3350 7430
rect 3350 7400 3380 7430
rect 3380 7400 3385 7430
rect 3345 7395 3385 7400
rect 3345 7360 3385 7365
rect 3345 7330 3350 7360
rect 3350 7330 3380 7360
rect 3380 7330 3385 7360
rect 3345 7325 3385 7330
rect 3345 7295 3385 7300
rect 3345 7265 3350 7295
rect 3350 7265 3380 7295
rect 3380 7265 3385 7295
rect 3345 7260 3385 7265
rect 3345 7235 3385 7240
rect 3345 7205 3350 7235
rect 3350 7205 3380 7235
rect 3380 7205 3385 7235
rect 3345 7200 3385 7205
rect 3345 7170 3385 7175
rect 3345 7140 3350 7170
rect 3350 7140 3380 7170
rect 3380 7140 3385 7170
rect 3345 7135 3385 7140
rect 3345 7100 3385 7105
rect 3345 7070 3350 7100
rect 3350 7070 3380 7100
rect 3380 7070 3385 7100
rect 3345 7065 3385 7070
rect 3345 7030 3385 7035
rect 3345 7000 3350 7030
rect 3350 7000 3380 7030
rect 3380 7000 3385 7030
rect 3345 6995 3385 7000
rect 3345 6960 3385 6965
rect 3345 6930 3350 6960
rect 3350 6930 3380 6960
rect 3380 6930 3385 6960
rect 3345 6925 3385 6930
rect 3345 6895 3385 6900
rect 3345 6865 3350 6895
rect 3350 6865 3380 6895
rect 3380 6865 3385 6895
rect 3345 6860 3385 6865
rect 3345 6835 3385 6840
rect 3345 6805 3350 6835
rect 3350 6805 3380 6835
rect 3380 6805 3385 6835
rect 3345 6800 3385 6805
rect 3345 6770 3385 6775
rect 3345 6740 3350 6770
rect 3350 6740 3380 6770
rect 3380 6740 3385 6770
rect 3345 6735 3385 6740
rect 3345 6700 3385 6705
rect 3345 6670 3350 6700
rect 3350 6670 3380 6700
rect 3380 6670 3385 6700
rect 3345 6665 3385 6670
rect 3345 6630 3385 6635
rect 3345 6600 3350 6630
rect 3350 6600 3380 6630
rect 3380 6600 3385 6630
rect 3345 6595 3385 6600
rect 3345 6560 3385 6565
rect 3345 6530 3350 6560
rect 3350 6530 3380 6560
rect 3380 6530 3385 6560
rect 3345 6525 3385 6530
rect 3345 6495 3385 6500
rect 3345 6465 3350 6495
rect 3350 6465 3380 6495
rect 3380 6465 3385 6495
rect 3345 6460 3385 6465
rect 6700 9635 6740 9640
rect 6700 9605 6705 9635
rect 6705 9605 6735 9635
rect 6735 9605 6740 9635
rect 6700 9600 6740 9605
rect 6700 9570 6740 9575
rect 6700 9540 6705 9570
rect 6705 9540 6735 9570
rect 6735 9540 6740 9570
rect 6700 9535 6740 9540
rect 6700 9500 6740 9505
rect 6700 9470 6705 9500
rect 6705 9470 6735 9500
rect 6735 9470 6740 9500
rect 6700 9465 6740 9470
rect 6700 9430 6740 9435
rect 6700 9400 6705 9430
rect 6705 9400 6735 9430
rect 6735 9400 6740 9430
rect 6700 9395 6740 9400
rect 6700 9360 6740 9365
rect 6700 9330 6705 9360
rect 6705 9330 6735 9360
rect 6735 9330 6740 9360
rect 6700 9325 6740 9330
rect 6700 9295 6740 9300
rect 6700 9265 6705 9295
rect 6705 9265 6735 9295
rect 6735 9265 6740 9295
rect 6700 9260 6740 9265
rect 6700 9235 6740 9240
rect 6700 9205 6705 9235
rect 6705 9205 6735 9235
rect 6735 9205 6740 9235
rect 6700 9200 6740 9205
rect 6700 9170 6740 9175
rect 6700 9140 6705 9170
rect 6705 9140 6735 9170
rect 6735 9140 6740 9170
rect 6700 9135 6740 9140
rect 6700 9100 6740 9105
rect 6700 9070 6705 9100
rect 6705 9070 6735 9100
rect 6735 9070 6740 9100
rect 6700 9065 6740 9070
rect 6700 9030 6740 9035
rect 6700 9000 6705 9030
rect 6705 9000 6735 9030
rect 6735 9000 6740 9030
rect 6700 8995 6740 9000
rect 6700 8960 6740 8965
rect 6700 8930 6705 8960
rect 6705 8930 6735 8960
rect 6735 8930 6740 8960
rect 6700 8925 6740 8930
rect 6700 8895 6740 8900
rect 6700 8865 6705 8895
rect 6705 8865 6735 8895
rect 6735 8865 6740 8895
rect 6700 8860 6740 8865
rect 6700 8835 6740 8840
rect 6700 8805 6705 8835
rect 6705 8805 6735 8835
rect 6735 8805 6740 8835
rect 6700 8800 6740 8805
rect 6700 8770 6740 8775
rect 6700 8740 6705 8770
rect 6705 8740 6735 8770
rect 6735 8740 6740 8770
rect 6700 8735 6740 8740
rect 6700 8700 6740 8705
rect 6700 8670 6705 8700
rect 6705 8670 6735 8700
rect 6735 8670 6740 8700
rect 6700 8665 6740 8670
rect 6700 8630 6740 8635
rect 6700 8600 6705 8630
rect 6705 8600 6735 8630
rect 6735 8600 6740 8630
rect 6700 8595 6740 8600
rect 6700 8560 6740 8565
rect 6700 8530 6705 8560
rect 6705 8530 6735 8560
rect 6735 8530 6740 8560
rect 6700 8525 6740 8530
rect 6700 8495 6740 8500
rect 6700 8465 6705 8495
rect 6705 8465 6735 8495
rect 6735 8465 6740 8495
rect 6700 8460 6740 8465
rect 6700 8435 6740 8440
rect 6700 8405 6705 8435
rect 6705 8405 6735 8435
rect 6735 8405 6740 8435
rect 6700 8400 6740 8405
rect 6700 8370 6740 8375
rect 6700 8340 6705 8370
rect 6705 8340 6735 8370
rect 6735 8340 6740 8370
rect 6700 8335 6740 8340
rect 6700 8300 6740 8305
rect 6700 8270 6705 8300
rect 6705 8270 6735 8300
rect 6735 8270 6740 8300
rect 6700 8265 6740 8270
rect 6700 8230 6740 8235
rect 6700 8200 6705 8230
rect 6705 8200 6735 8230
rect 6735 8200 6740 8230
rect 6700 8195 6740 8200
rect 6700 8160 6740 8165
rect 6700 8130 6705 8160
rect 6705 8130 6735 8160
rect 6735 8130 6740 8160
rect 6700 8125 6740 8130
rect 6700 8095 6740 8100
rect 6700 8065 6705 8095
rect 6705 8065 6735 8095
rect 6735 8065 6740 8095
rect 6700 8060 6740 8065
rect 6700 8035 6740 8040
rect 6700 8005 6705 8035
rect 6705 8005 6735 8035
rect 6735 8005 6740 8035
rect 6700 8000 6740 8005
rect 6700 7970 6740 7975
rect 6700 7940 6705 7970
rect 6705 7940 6735 7970
rect 6735 7940 6740 7970
rect 6700 7935 6740 7940
rect 6700 7900 6740 7905
rect 6700 7870 6705 7900
rect 6705 7870 6735 7900
rect 6735 7870 6740 7900
rect 6700 7865 6740 7870
rect 6700 7830 6740 7835
rect 6700 7800 6705 7830
rect 6705 7800 6735 7830
rect 6735 7800 6740 7830
rect 6700 7795 6740 7800
rect 6700 7760 6740 7765
rect 6700 7730 6705 7760
rect 6705 7730 6735 7760
rect 6735 7730 6740 7760
rect 6700 7725 6740 7730
rect 6700 7695 6740 7700
rect 6700 7665 6705 7695
rect 6705 7665 6735 7695
rect 6735 7665 6740 7695
rect 6700 7660 6740 7665
rect 6700 7635 6740 7640
rect 6700 7605 6705 7635
rect 6705 7605 6735 7635
rect 6735 7605 6740 7635
rect 6700 7600 6740 7605
rect 6700 7570 6740 7575
rect 6700 7540 6705 7570
rect 6705 7540 6735 7570
rect 6735 7540 6740 7570
rect 6700 7535 6740 7540
rect 6700 7500 6740 7505
rect 6700 7470 6705 7500
rect 6705 7470 6735 7500
rect 6735 7470 6740 7500
rect 6700 7465 6740 7470
rect 6700 7430 6740 7435
rect 6700 7400 6705 7430
rect 6705 7400 6735 7430
rect 6735 7400 6740 7430
rect 6700 7395 6740 7400
rect 6700 7360 6740 7365
rect 6700 7330 6705 7360
rect 6705 7330 6735 7360
rect 6735 7330 6740 7360
rect 6700 7325 6740 7330
rect 6700 7295 6740 7300
rect 6700 7265 6705 7295
rect 6705 7265 6735 7295
rect 6735 7265 6740 7295
rect 6700 7260 6740 7265
rect 6700 7235 6740 7240
rect 6700 7205 6705 7235
rect 6705 7205 6735 7235
rect 6735 7205 6740 7235
rect 6700 7200 6740 7205
rect 6700 7170 6740 7175
rect 6700 7140 6705 7170
rect 6705 7140 6735 7170
rect 6735 7140 6740 7170
rect 6700 7135 6740 7140
rect 6700 7100 6740 7105
rect 6700 7070 6705 7100
rect 6705 7070 6735 7100
rect 6735 7070 6740 7100
rect 6700 7065 6740 7070
rect 6700 7030 6740 7035
rect 6700 7000 6705 7030
rect 6705 7000 6735 7030
rect 6735 7000 6740 7030
rect 6700 6995 6740 7000
rect 6700 6960 6740 6965
rect 6700 6930 6705 6960
rect 6705 6930 6735 6960
rect 6735 6930 6740 6960
rect 6700 6925 6740 6930
rect 6700 6895 6740 6900
rect 6700 6865 6705 6895
rect 6705 6865 6735 6895
rect 6735 6865 6740 6895
rect 6700 6860 6740 6865
rect 6700 6835 6740 6840
rect 6700 6805 6705 6835
rect 6705 6805 6735 6835
rect 6735 6805 6740 6835
rect 6700 6800 6740 6805
rect 6700 6770 6740 6775
rect 6700 6740 6705 6770
rect 6705 6740 6735 6770
rect 6735 6740 6740 6770
rect 6700 6735 6740 6740
rect 6700 6700 6740 6705
rect 6700 6670 6705 6700
rect 6705 6670 6735 6700
rect 6735 6670 6740 6700
rect 6700 6665 6740 6670
rect 6700 6630 6740 6635
rect 6700 6600 6705 6630
rect 6705 6600 6735 6630
rect 6735 6600 6740 6630
rect 6700 6595 6740 6600
rect 6700 6560 6740 6565
rect 6700 6530 6705 6560
rect 6705 6530 6735 6560
rect 6735 6530 6740 6560
rect 6700 6525 6740 6530
rect 6700 6495 6740 6500
rect 6700 6465 6705 6495
rect 6705 6465 6735 6495
rect 6735 6465 6740 6495
rect 6700 6460 6740 6465
rect 7270 9635 7310 9640
rect 7270 9605 7275 9635
rect 7275 9605 7305 9635
rect 7305 9605 7310 9635
rect 7270 9600 7310 9605
rect 7270 9570 7310 9575
rect 7270 9540 7275 9570
rect 7275 9540 7305 9570
rect 7305 9540 7310 9570
rect 7270 9535 7310 9540
rect 7270 9500 7310 9505
rect 7270 9470 7275 9500
rect 7275 9470 7305 9500
rect 7305 9470 7310 9500
rect 7270 9465 7310 9470
rect 7270 9430 7310 9435
rect 7270 9400 7275 9430
rect 7275 9400 7305 9430
rect 7305 9400 7310 9430
rect 7270 9395 7310 9400
rect 7270 9360 7310 9365
rect 7270 9330 7275 9360
rect 7275 9330 7305 9360
rect 7305 9330 7310 9360
rect 7270 9325 7310 9330
rect 7270 9295 7310 9300
rect 7270 9265 7275 9295
rect 7275 9265 7305 9295
rect 7305 9265 7310 9295
rect 7270 9260 7310 9265
rect 7270 9235 7310 9240
rect 7270 9205 7275 9235
rect 7275 9205 7305 9235
rect 7305 9205 7310 9235
rect 7270 9200 7310 9205
rect 7270 9170 7310 9175
rect 7270 9140 7275 9170
rect 7275 9140 7305 9170
rect 7305 9140 7310 9170
rect 7270 9135 7310 9140
rect 7270 9100 7310 9105
rect 7270 9070 7275 9100
rect 7275 9070 7305 9100
rect 7305 9070 7310 9100
rect 7270 9065 7310 9070
rect 7270 9030 7310 9035
rect 7270 9000 7275 9030
rect 7275 9000 7305 9030
rect 7305 9000 7310 9030
rect 7270 8995 7310 9000
rect 7270 8960 7310 8965
rect 7270 8930 7275 8960
rect 7275 8930 7305 8960
rect 7305 8930 7310 8960
rect 7270 8925 7310 8930
rect 7270 8895 7310 8900
rect 7270 8865 7275 8895
rect 7275 8865 7305 8895
rect 7305 8865 7310 8895
rect 7270 8860 7310 8865
rect 7270 8835 7310 8840
rect 7270 8805 7275 8835
rect 7275 8805 7305 8835
rect 7305 8805 7310 8835
rect 7270 8800 7310 8805
rect 7270 8770 7310 8775
rect 7270 8740 7275 8770
rect 7275 8740 7305 8770
rect 7305 8740 7310 8770
rect 7270 8735 7310 8740
rect 7270 8700 7310 8705
rect 7270 8670 7275 8700
rect 7275 8670 7305 8700
rect 7305 8670 7310 8700
rect 7270 8665 7310 8670
rect 7270 8630 7310 8635
rect 7270 8600 7275 8630
rect 7275 8600 7305 8630
rect 7305 8600 7310 8630
rect 7270 8595 7310 8600
rect 7270 8560 7310 8565
rect 7270 8530 7275 8560
rect 7275 8530 7305 8560
rect 7305 8530 7310 8560
rect 7270 8525 7310 8530
rect 7270 8495 7310 8500
rect 7270 8465 7275 8495
rect 7275 8465 7305 8495
rect 7305 8465 7310 8495
rect 7270 8460 7310 8465
rect 7270 8435 7310 8440
rect 7270 8405 7275 8435
rect 7275 8405 7305 8435
rect 7305 8405 7310 8435
rect 7270 8400 7310 8405
rect 7270 8370 7310 8375
rect 7270 8340 7275 8370
rect 7275 8340 7305 8370
rect 7305 8340 7310 8370
rect 7270 8335 7310 8340
rect 7270 8300 7310 8305
rect 7270 8270 7275 8300
rect 7275 8270 7305 8300
rect 7305 8270 7310 8300
rect 7270 8265 7310 8270
rect 7270 8230 7310 8235
rect 7270 8200 7275 8230
rect 7275 8200 7305 8230
rect 7305 8200 7310 8230
rect 7270 8195 7310 8200
rect 7270 8160 7310 8165
rect 7270 8130 7275 8160
rect 7275 8130 7305 8160
rect 7305 8130 7310 8160
rect 7270 8125 7310 8130
rect 7270 8095 7310 8100
rect 7270 8065 7275 8095
rect 7275 8065 7305 8095
rect 7305 8065 7310 8095
rect 7270 8060 7310 8065
rect 7270 8035 7310 8040
rect 7270 8005 7275 8035
rect 7275 8005 7305 8035
rect 7305 8005 7310 8035
rect 7270 8000 7310 8005
rect 7270 7970 7310 7975
rect 7270 7940 7275 7970
rect 7275 7940 7305 7970
rect 7305 7940 7310 7970
rect 7270 7935 7310 7940
rect 7270 7900 7310 7905
rect 7270 7870 7275 7900
rect 7275 7870 7305 7900
rect 7305 7870 7310 7900
rect 7270 7865 7310 7870
rect 7270 7830 7310 7835
rect 7270 7800 7275 7830
rect 7275 7800 7305 7830
rect 7305 7800 7310 7830
rect 7270 7795 7310 7800
rect 7270 7760 7310 7765
rect 7270 7730 7275 7760
rect 7275 7730 7305 7760
rect 7305 7730 7310 7760
rect 7270 7725 7310 7730
rect 7270 7695 7310 7700
rect 7270 7665 7275 7695
rect 7275 7665 7305 7695
rect 7305 7665 7310 7695
rect 7270 7660 7310 7665
rect 7270 7635 7310 7640
rect 7270 7605 7275 7635
rect 7275 7605 7305 7635
rect 7305 7605 7310 7635
rect 7270 7600 7310 7605
rect 7270 7570 7310 7575
rect 7270 7540 7275 7570
rect 7275 7540 7305 7570
rect 7305 7540 7310 7570
rect 7270 7535 7310 7540
rect 7270 7500 7310 7505
rect 7270 7470 7275 7500
rect 7275 7470 7305 7500
rect 7305 7470 7310 7500
rect 7270 7465 7310 7470
rect 7270 7430 7310 7435
rect 7270 7400 7275 7430
rect 7275 7400 7305 7430
rect 7305 7400 7310 7430
rect 7270 7395 7310 7400
rect 7270 7360 7310 7365
rect 7270 7330 7275 7360
rect 7275 7330 7305 7360
rect 7305 7330 7310 7360
rect 7270 7325 7310 7330
rect 7270 7295 7310 7300
rect 7270 7265 7275 7295
rect 7275 7265 7305 7295
rect 7305 7265 7310 7295
rect 7270 7260 7310 7265
rect 7270 7235 7310 7240
rect 7270 7205 7275 7235
rect 7275 7205 7305 7235
rect 7305 7205 7310 7235
rect 7270 7200 7310 7205
rect 7270 7170 7310 7175
rect 7270 7140 7275 7170
rect 7275 7140 7305 7170
rect 7305 7140 7310 7170
rect 7270 7135 7310 7140
rect 7270 7100 7310 7105
rect 7270 7070 7275 7100
rect 7275 7070 7305 7100
rect 7305 7070 7310 7100
rect 7270 7065 7310 7070
rect 7270 7030 7310 7035
rect 7270 7000 7275 7030
rect 7275 7000 7305 7030
rect 7305 7000 7310 7030
rect 7270 6995 7310 7000
rect 7270 6960 7310 6965
rect 7270 6930 7275 6960
rect 7275 6930 7305 6960
rect 7305 6930 7310 6960
rect 7270 6925 7310 6930
rect 7270 6895 7310 6900
rect 7270 6865 7275 6895
rect 7275 6865 7305 6895
rect 7305 6865 7310 6895
rect 7270 6860 7310 6865
rect 7270 6835 7310 6840
rect 7270 6805 7275 6835
rect 7275 6805 7305 6835
rect 7305 6805 7310 6835
rect 7270 6800 7310 6805
rect 7270 6770 7310 6775
rect 7270 6740 7275 6770
rect 7275 6740 7305 6770
rect 7305 6740 7310 6770
rect 7270 6735 7310 6740
rect 7270 6700 7310 6705
rect 7270 6670 7275 6700
rect 7275 6670 7305 6700
rect 7305 6670 7310 6700
rect 7270 6665 7310 6670
rect 7270 6630 7310 6635
rect 7270 6600 7275 6630
rect 7275 6600 7305 6630
rect 7305 6600 7310 6630
rect 7270 6595 7310 6600
rect 7270 6560 7310 6565
rect 7270 6530 7275 6560
rect 7275 6530 7305 6560
rect 7305 6530 7310 6560
rect 7270 6525 7310 6530
rect 7270 6495 7310 6500
rect 7270 6465 7275 6495
rect 7275 6465 7305 6495
rect 7305 6465 7310 6495
rect 7270 6460 7310 6465
rect 7970 9635 8010 9640
rect 7970 9605 7975 9635
rect 7975 9605 8005 9635
rect 8005 9605 8010 9635
rect 7970 9600 8010 9605
rect 7970 9570 8010 9575
rect 7970 9540 7975 9570
rect 7975 9540 8005 9570
rect 8005 9540 8010 9570
rect 7970 9535 8010 9540
rect 7970 9500 8010 9505
rect 7970 9470 7975 9500
rect 7975 9470 8005 9500
rect 8005 9470 8010 9500
rect 7970 9465 8010 9470
rect 7970 9430 8010 9435
rect 7970 9400 7975 9430
rect 7975 9400 8005 9430
rect 8005 9400 8010 9430
rect 7970 9395 8010 9400
rect 7970 9360 8010 9365
rect 7970 9330 7975 9360
rect 7975 9330 8005 9360
rect 8005 9330 8010 9360
rect 7970 9325 8010 9330
rect 7970 9295 8010 9300
rect 7970 9265 7975 9295
rect 7975 9265 8005 9295
rect 8005 9265 8010 9295
rect 7970 9260 8010 9265
rect 7970 9235 8010 9240
rect 7970 9205 7975 9235
rect 7975 9205 8005 9235
rect 8005 9205 8010 9235
rect 7970 9200 8010 9205
rect 7970 9170 8010 9175
rect 7970 9140 7975 9170
rect 7975 9140 8005 9170
rect 8005 9140 8010 9170
rect 7970 9135 8010 9140
rect 7970 9100 8010 9105
rect 7970 9070 7975 9100
rect 7975 9070 8005 9100
rect 8005 9070 8010 9100
rect 7970 9065 8010 9070
rect 7970 9030 8010 9035
rect 7970 9000 7975 9030
rect 7975 9000 8005 9030
rect 8005 9000 8010 9030
rect 7970 8995 8010 9000
rect 7970 8960 8010 8965
rect 7970 8930 7975 8960
rect 7975 8930 8005 8960
rect 8005 8930 8010 8960
rect 7970 8925 8010 8930
rect 7970 8895 8010 8900
rect 7970 8865 7975 8895
rect 7975 8865 8005 8895
rect 8005 8865 8010 8895
rect 7970 8860 8010 8865
rect 7970 8835 8010 8840
rect 7970 8805 7975 8835
rect 7975 8805 8005 8835
rect 8005 8805 8010 8835
rect 7970 8800 8010 8805
rect 7970 8770 8010 8775
rect 7970 8740 7975 8770
rect 7975 8740 8005 8770
rect 8005 8740 8010 8770
rect 7970 8735 8010 8740
rect 7970 8700 8010 8705
rect 7970 8670 7975 8700
rect 7975 8670 8005 8700
rect 8005 8670 8010 8700
rect 7970 8665 8010 8670
rect 7970 8630 8010 8635
rect 7970 8600 7975 8630
rect 7975 8600 8005 8630
rect 8005 8600 8010 8630
rect 7970 8595 8010 8600
rect 7970 8560 8010 8565
rect 7970 8530 7975 8560
rect 7975 8530 8005 8560
rect 8005 8530 8010 8560
rect 7970 8525 8010 8530
rect 7970 8495 8010 8500
rect 7970 8465 7975 8495
rect 7975 8465 8005 8495
rect 8005 8465 8010 8495
rect 7970 8460 8010 8465
rect 7970 8435 8010 8440
rect 7970 8405 7975 8435
rect 7975 8405 8005 8435
rect 8005 8405 8010 8435
rect 7970 8400 8010 8405
rect 7970 8370 8010 8375
rect 7970 8340 7975 8370
rect 7975 8340 8005 8370
rect 8005 8340 8010 8370
rect 7970 8335 8010 8340
rect 7970 8300 8010 8305
rect 7970 8270 7975 8300
rect 7975 8270 8005 8300
rect 8005 8270 8010 8300
rect 7970 8265 8010 8270
rect 7970 8230 8010 8235
rect 7970 8200 7975 8230
rect 7975 8200 8005 8230
rect 8005 8200 8010 8230
rect 7970 8195 8010 8200
rect 7970 8160 8010 8165
rect 7970 8130 7975 8160
rect 7975 8130 8005 8160
rect 8005 8130 8010 8160
rect 7970 8125 8010 8130
rect 7970 8095 8010 8100
rect 7970 8065 7975 8095
rect 7975 8065 8005 8095
rect 8005 8065 8010 8095
rect 7970 8060 8010 8065
rect 7970 8035 8010 8040
rect 7970 8005 7975 8035
rect 7975 8005 8005 8035
rect 8005 8005 8010 8035
rect 7970 8000 8010 8005
rect 7970 7970 8010 7975
rect 7970 7940 7975 7970
rect 7975 7940 8005 7970
rect 8005 7940 8010 7970
rect 7970 7935 8010 7940
rect 7970 7900 8010 7905
rect 7970 7870 7975 7900
rect 7975 7870 8005 7900
rect 8005 7870 8010 7900
rect 7970 7865 8010 7870
rect 7970 7830 8010 7835
rect 7970 7800 7975 7830
rect 7975 7800 8005 7830
rect 8005 7800 8010 7830
rect 7970 7795 8010 7800
rect 7970 7760 8010 7765
rect 7970 7730 7975 7760
rect 7975 7730 8005 7760
rect 8005 7730 8010 7760
rect 7970 7725 8010 7730
rect 7970 7695 8010 7700
rect 7970 7665 7975 7695
rect 7975 7665 8005 7695
rect 8005 7665 8010 7695
rect 7970 7660 8010 7665
rect 7970 7635 8010 7640
rect 7970 7605 7975 7635
rect 7975 7605 8005 7635
rect 8005 7605 8010 7635
rect 7970 7600 8010 7605
rect 7970 7570 8010 7575
rect 7970 7540 7975 7570
rect 7975 7540 8005 7570
rect 8005 7540 8010 7570
rect 7970 7535 8010 7540
rect 7970 7500 8010 7505
rect 7970 7470 7975 7500
rect 7975 7470 8005 7500
rect 8005 7470 8010 7500
rect 7970 7465 8010 7470
rect 7970 7430 8010 7435
rect 7970 7400 7975 7430
rect 7975 7400 8005 7430
rect 8005 7400 8010 7430
rect 7970 7395 8010 7400
rect 7970 7360 8010 7365
rect 7970 7330 7975 7360
rect 7975 7330 8005 7360
rect 8005 7330 8010 7360
rect 7970 7325 8010 7330
rect 7970 7295 8010 7300
rect 7970 7265 7975 7295
rect 7975 7265 8005 7295
rect 8005 7265 8010 7295
rect 7970 7260 8010 7265
rect 7970 7235 8010 7240
rect 7970 7205 7975 7235
rect 7975 7205 8005 7235
rect 8005 7205 8010 7235
rect 7970 7200 8010 7205
rect 7970 7170 8010 7175
rect 7970 7140 7975 7170
rect 7975 7140 8005 7170
rect 8005 7140 8010 7170
rect 7970 7135 8010 7140
rect 7970 7100 8010 7105
rect 7970 7070 7975 7100
rect 7975 7070 8005 7100
rect 8005 7070 8010 7100
rect 7970 7065 8010 7070
rect 7970 7030 8010 7035
rect 7970 7000 7975 7030
rect 7975 7000 8005 7030
rect 8005 7000 8010 7030
rect 7970 6995 8010 7000
rect 7970 6960 8010 6965
rect 7970 6930 7975 6960
rect 7975 6930 8005 6960
rect 8005 6930 8010 6960
rect 7970 6925 8010 6930
rect 7970 6895 8010 6900
rect 7970 6865 7975 6895
rect 7975 6865 8005 6895
rect 8005 6865 8010 6895
rect 7970 6860 8010 6865
rect 7970 6835 8010 6840
rect 7970 6805 7975 6835
rect 7975 6805 8005 6835
rect 8005 6805 8010 6835
rect 7970 6800 8010 6805
rect 7970 6770 8010 6775
rect 7970 6740 7975 6770
rect 7975 6740 8005 6770
rect 8005 6740 8010 6770
rect 7970 6735 8010 6740
rect 7970 6700 8010 6705
rect 7970 6670 7975 6700
rect 7975 6670 8005 6700
rect 8005 6670 8010 6700
rect 7970 6665 8010 6670
rect 7970 6630 8010 6635
rect 7970 6600 7975 6630
rect 7975 6600 8005 6630
rect 8005 6600 8010 6630
rect 7970 6595 8010 6600
rect 7970 6560 8010 6565
rect 7970 6530 7975 6560
rect 7975 6530 8005 6560
rect 8005 6530 8010 6560
rect 7970 6525 8010 6530
rect 7970 6495 8010 6500
rect 7970 6465 7975 6495
rect 7975 6465 8005 6495
rect 8005 6465 8010 6495
rect 7970 6460 8010 6465
rect 8320 9635 8360 9640
rect 8320 9605 8325 9635
rect 8325 9605 8355 9635
rect 8355 9605 8360 9635
rect 8320 9600 8360 9605
rect 8320 9570 8360 9575
rect 8320 9540 8325 9570
rect 8325 9540 8355 9570
rect 8355 9540 8360 9570
rect 8320 9535 8360 9540
rect 8320 9500 8360 9505
rect 8320 9470 8325 9500
rect 8325 9470 8355 9500
rect 8355 9470 8360 9500
rect 8320 9465 8360 9470
rect 8320 9430 8360 9435
rect 8320 9400 8325 9430
rect 8325 9400 8355 9430
rect 8355 9400 8360 9430
rect 8320 9395 8360 9400
rect 8320 9360 8360 9365
rect 8320 9330 8325 9360
rect 8325 9330 8355 9360
rect 8355 9330 8360 9360
rect 8320 9325 8360 9330
rect 8320 9295 8360 9300
rect 8320 9265 8325 9295
rect 8325 9265 8355 9295
rect 8355 9265 8360 9295
rect 8320 9260 8360 9265
rect 8320 9235 8360 9240
rect 8320 9205 8325 9235
rect 8325 9205 8355 9235
rect 8355 9205 8360 9235
rect 8320 9200 8360 9205
rect 8320 9170 8360 9175
rect 8320 9140 8325 9170
rect 8325 9140 8355 9170
rect 8355 9140 8360 9170
rect 8320 9135 8360 9140
rect 8320 9100 8360 9105
rect 8320 9070 8325 9100
rect 8325 9070 8355 9100
rect 8355 9070 8360 9100
rect 8320 9065 8360 9070
rect 8320 9030 8360 9035
rect 8320 9000 8325 9030
rect 8325 9000 8355 9030
rect 8355 9000 8360 9030
rect 8320 8995 8360 9000
rect 8320 8960 8360 8965
rect 8320 8930 8325 8960
rect 8325 8930 8355 8960
rect 8355 8930 8360 8960
rect 8320 8925 8360 8930
rect 8320 8895 8360 8900
rect 8320 8865 8325 8895
rect 8325 8865 8355 8895
rect 8355 8865 8360 8895
rect 8320 8860 8360 8865
rect 8320 8835 8360 8840
rect 8320 8805 8325 8835
rect 8325 8805 8355 8835
rect 8355 8805 8360 8835
rect 8320 8800 8360 8805
rect 8320 8770 8360 8775
rect 8320 8740 8325 8770
rect 8325 8740 8355 8770
rect 8355 8740 8360 8770
rect 8320 8735 8360 8740
rect 8320 8700 8360 8705
rect 8320 8670 8325 8700
rect 8325 8670 8355 8700
rect 8355 8670 8360 8700
rect 8320 8665 8360 8670
rect 8320 8630 8360 8635
rect 8320 8600 8325 8630
rect 8325 8600 8355 8630
rect 8355 8600 8360 8630
rect 8320 8595 8360 8600
rect 8320 8560 8360 8565
rect 8320 8530 8325 8560
rect 8325 8530 8355 8560
rect 8355 8530 8360 8560
rect 8320 8525 8360 8530
rect 8320 8495 8360 8500
rect 8320 8465 8325 8495
rect 8325 8465 8355 8495
rect 8355 8465 8360 8495
rect 8320 8460 8360 8465
rect 8320 8435 8360 8440
rect 8320 8405 8325 8435
rect 8325 8405 8355 8435
rect 8355 8405 8360 8435
rect 8320 8400 8360 8405
rect 8320 8370 8360 8375
rect 8320 8340 8325 8370
rect 8325 8340 8355 8370
rect 8355 8340 8360 8370
rect 8320 8335 8360 8340
rect 8320 8300 8360 8305
rect 8320 8270 8325 8300
rect 8325 8270 8355 8300
rect 8355 8270 8360 8300
rect 8320 8265 8360 8270
rect 8320 8230 8360 8235
rect 8320 8200 8325 8230
rect 8325 8200 8355 8230
rect 8355 8200 8360 8230
rect 8320 8195 8360 8200
rect 8320 8160 8360 8165
rect 8320 8130 8325 8160
rect 8325 8130 8355 8160
rect 8355 8130 8360 8160
rect 8320 8125 8360 8130
rect 8320 8095 8360 8100
rect 8320 8065 8325 8095
rect 8325 8065 8355 8095
rect 8355 8065 8360 8095
rect 8320 8060 8360 8065
rect 8320 8035 8360 8040
rect 8320 8005 8325 8035
rect 8325 8005 8355 8035
rect 8355 8005 8360 8035
rect 8320 8000 8360 8005
rect 8320 7970 8360 7975
rect 8320 7940 8325 7970
rect 8325 7940 8355 7970
rect 8355 7940 8360 7970
rect 8320 7935 8360 7940
rect 8320 7900 8360 7905
rect 8320 7870 8325 7900
rect 8325 7870 8355 7900
rect 8355 7870 8360 7900
rect 8320 7865 8360 7870
rect 8320 7830 8360 7835
rect 8320 7800 8325 7830
rect 8325 7800 8355 7830
rect 8355 7800 8360 7830
rect 8320 7795 8360 7800
rect 8320 7760 8360 7765
rect 8320 7730 8325 7760
rect 8325 7730 8355 7760
rect 8355 7730 8360 7760
rect 8320 7725 8360 7730
rect 8320 7695 8360 7700
rect 8320 7665 8325 7695
rect 8325 7665 8355 7695
rect 8355 7665 8360 7695
rect 8320 7660 8360 7665
rect 8320 7635 8360 7640
rect 8320 7605 8325 7635
rect 8325 7605 8355 7635
rect 8355 7605 8360 7635
rect 8320 7600 8360 7605
rect 8320 7570 8360 7575
rect 8320 7540 8325 7570
rect 8325 7540 8355 7570
rect 8355 7540 8360 7570
rect 8320 7535 8360 7540
rect 8320 7500 8360 7505
rect 8320 7470 8325 7500
rect 8325 7470 8355 7500
rect 8355 7470 8360 7500
rect 8320 7465 8360 7470
rect 8320 7430 8360 7435
rect 8320 7400 8325 7430
rect 8325 7400 8355 7430
rect 8355 7400 8360 7430
rect 8320 7395 8360 7400
rect 8320 7360 8360 7365
rect 8320 7330 8325 7360
rect 8325 7330 8355 7360
rect 8355 7330 8360 7360
rect 8320 7325 8360 7330
rect 8320 7295 8360 7300
rect 8320 7265 8325 7295
rect 8325 7265 8355 7295
rect 8355 7265 8360 7295
rect 8320 7260 8360 7265
rect 8320 7235 8360 7240
rect 8320 7205 8325 7235
rect 8325 7205 8355 7235
rect 8355 7205 8360 7235
rect 8320 7200 8360 7205
rect 8320 7170 8360 7175
rect 8320 7140 8325 7170
rect 8325 7140 8355 7170
rect 8355 7140 8360 7170
rect 8320 7135 8360 7140
rect 8320 7100 8360 7105
rect 8320 7070 8325 7100
rect 8325 7070 8355 7100
rect 8355 7070 8360 7100
rect 8320 7065 8360 7070
rect 8320 7030 8360 7035
rect 8320 7000 8325 7030
rect 8325 7000 8355 7030
rect 8355 7000 8360 7030
rect 8320 6995 8360 7000
rect 8320 6960 8360 6965
rect 8320 6930 8325 6960
rect 8325 6930 8355 6960
rect 8355 6930 8360 6960
rect 8320 6925 8360 6930
rect 8320 6895 8360 6900
rect 8320 6865 8325 6895
rect 8325 6865 8355 6895
rect 8355 6865 8360 6895
rect 8320 6860 8360 6865
rect 8320 6835 8360 6840
rect 8320 6805 8325 6835
rect 8325 6805 8355 6835
rect 8355 6805 8360 6835
rect 8320 6800 8360 6805
rect 8320 6770 8360 6775
rect 8320 6740 8325 6770
rect 8325 6740 8355 6770
rect 8355 6740 8360 6770
rect 8320 6735 8360 6740
rect 8320 6700 8360 6705
rect 8320 6670 8325 6700
rect 8325 6670 8355 6700
rect 8355 6670 8360 6700
rect 8320 6665 8360 6670
rect 8320 6630 8360 6635
rect 8320 6600 8325 6630
rect 8325 6600 8355 6630
rect 8355 6600 8360 6630
rect 8320 6595 8360 6600
rect 8320 6560 8360 6565
rect 8320 6530 8325 6560
rect 8325 6530 8355 6560
rect 8355 6530 8360 6560
rect 8320 6525 8360 6530
rect 8320 6495 8360 6500
rect 8320 6465 8325 6495
rect 8325 6465 8355 6495
rect 8355 6465 8360 6495
rect 8320 6460 8360 6465
rect 8670 9635 8710 9640
rect 8670 9605 8675 9635
rect 8675 9605 8705 9635
rect 8705 9605 8710 9635
rect 8670 9600 8710 9605
rect 8670 9570 8710 9575
rect 8670 9540 8675 9570
rect 8675 9540 8705 9570
rect 8705 9540 8710 9570
rect 8670 9535 8710 9540
rect 8670 9500 8710 9505
rect 8670 9470 8675 9500
rect 8675 9470 8705 9500
rect 8705 9470 8710 9500
rect 8670 9465 8710 9470
rect 8670 9430 8710 9435
rect 8670 9400 8675 9430
rect 8675 9400 8705 9430
rect 8705 9400 8710 9430
rect 8670 9395 8710 9400
rect 8670 9360 8710 9365
rect 8670 9330 8675 9360
rect 8675 9330 8705 9360
rect 8705 9330 8710 9360
rect 8670 9325 8710 9330
rect 8670 9295 8710 9300
rect 8670 9265 8675 9295
rect 8675 9265 8705 9295
rect 8705 9265 8710 9295
rect 8670 9260 8710 9265
rect 8670 9235 8710 9240
rect 8670 9205 8675 9235
rect 8675 9205 8705 9235
rect 8705 9205 8710 9235
rect 8670 9200 8710 9205
rect 8670 9170 8710 9175
rect 8670 9140 8675 9170
rect 8675 9140 8705 9170
rect 8705 9140 8710 9170
rect 8670 9135 8710 9140
rect 8670 9100 8710 9105
rect 8670 9070 8675 9100
rect 8675 9070 8705 9100
rect 8705 9070 8710 9100
rect 8670 9065 8710 9070
rect 8670 9030 8710 9035
rect 8670 9000 8675 9030
rect 8675 9000 8705 9030
rect 8705 9000 8710 9030
rect 8670 8995 8710 9000
rect 8670 8960 8710 8965
rect 8670 8930 8675 8960
rect 8675 8930 8705 8960
rect 8705 8930 8710 8960
rect 8670 8925 8710 8930
rect 8670 8895 8710 8900
rect 8670 8865 8675 8895
rect 8675 8865 8705 8895
rect 8705 8865 8710 8895
rect 8670 8860 8710 8865
rect 8670 8835 8710 8840
rect 8670 8805 8675 8835
rect 8675 8805 8705 8835
rect 8705 8805 8710 8835
rect 8670 8800 8710 8805
rect 8670 8770 8710 8775
rect 8670 8740 8675 8770
rect 8675 8740 8705 8770
rect 8705 8740 8710 8770
rect 8670 8735 8710 8740
rect 8670 8700 8710 8705
rect 8670 8670 8675 8700
rect 8675 8670 8705 8700
rect 8705 8670 8710 8700
rect 8670 8665 8710 8670
rect 8670 8630 8710 8635
rect 8670 8600 8675 8630
rect 8675 8600 8705 8630
rect 8705 8600 8710 8630
rect 8670 8595 8710 8600
rect 8670 8560 8710 8565
rect 8670 8530 8675 8560
rect 8675 8530 8705 8560
rect 8705 8530 8710 8560
rect 8670 8525 8710 8530
rect 8670 8495 8710 8500
rect 8670 8465 8675 8495
rect 8675 8465 8705 8495
rect 8705 8465 8710 8495
rect 8670 8460 8710 8465
rect 8670 8435 8710 8440
rect 8670 8405 8675 8435
rect 8675 8405 8705 8435
rect 8705 8405 8710 8435
rect 8670 8400 8710 8405
rect 8670 8370 8710 8375
rect 8670 8340 8675 8370
rect 8675 8340 8705 8370
rect 8705 8340 8710 8370
rect 8670 8335 8710 8340
rect 8670 8300 8710 8305
rect 8670 8270 8675 8300
rect 8675 8270 8705 8300
rect 8705 8270 8710 8300
rect 8670 8265 8710 8270
rect 8670 8230 8710 8235
rect 8670 8200 8675 8230
rect 8675 8200 8705 8230
rect 8705 8200 8710 8230
rect 8670 8195 8710 8200
rect 8670 8160 8710 8165
rect 8670 8130 8675 8160
rect 8675 8130 8705 8160
rect 8705 8130 8710 8160
rect 8670 8125 8710 8130
rect 8670 8095 8710 8100
rect 8670 8065 8675 8095
rect 8675 8065 8705 8095
rect 8705 8065 8710 8095
rect 8670 8060 8710 8065
rect 8670 8035 8710 8040
rect 8670 8005 8675 8035
rect 8675 8005 8705 8035
rect 8705 8005 8710 8035
rect 8670 8000 8710 8005
rect 8670 7970 8710 7975
rect 8670 7940 8675 7970
rect 8675 7940 8705 7970
rect 8705 7940 8710 7970
rect 8670 7935 8710 7940
rect 8670 7900 8710 7905
rect 8670 7870 8675 7900
rect 8675 7870 8705 7900
rect 8705 7870 8710 7900
rect 8670 7865 8710 7870
rect 8670 7830 8710 7835
rect 8670 7800 8675 7830
rect 8675 7800 8705 7830
rect 8705 7800 8710 7830
rect 8670 7795 8710 7800
rect 8670 7760 8710 7765
rect 8670 7730 8675 7760
rect 8675 7730 8705 7760
rect 8705 7730 8710 7760
rect 8670 7725 8710 7730
rect 8670 7695 8710 7700
rect 8670 7665 8675 7695
rect 8675 7665 8705 7695
rect 8705 7665 8710 7695
rect 8670 7660 8710 7665
rect 8670 7635 8710 7640
rect 8670 7605 8675 7635
rect 8675 7605 8705 7635
rect 8705 7605 8710 7635
rect 8670 7600 8710 7605
rect 8670 7570 8710 7575
rect 8670 7540 8675 7570
rect 8675 7540 8705 7570
rect 8705 7540 8710 7570
rect 8670 7535 8710 7540
rect 8670 7500 8710 7505
rect 8670 7470 8675 7500
rect 8675 7470 8705 7500
rect 8705 7470 8710 7500
rect 8670 7465 8710 7470
rect 8670 7430 8710 7435
rect 8670 7400 8675 7430
rect 8675 7400 8705 7430
rect 8705 7400 8710 7430
rect 8670 7395 8710 7400
rect 8670 7360 8710 7365
rect 8670 7330 8675 7360
rect 8675 7330 8705 7360
rect 8705 7330 8710 7360
rect 8670 7325 8710 7330
rect 8670 7295 8710 7300
rect 8670 7265 8675 7295
rect 8675 7265 8705 7295
rect 8705 7265 8710 7295
rect 8670 7260 8710 7265
rect 8670 7235 8710 7240
rect 8670 7205 8675 7235
rect 8675 7205 8705 7235
rect 8705 7205 8710 7235
rect 8670 7200 8710 7205
rect 8670 7170 8710 7175
rect 8670 7140 8675 7170
rect 8675 7140 8705 7170
rect 8705 7140 8710 7170
rect 8670 7135 8710 7140
rect 8670 7100 8710 7105
rect 8670 7070 8675 7100
rect 8675 7070 8705 7100
rect 8705 7070 8710 7100
rect 8670 7065 8710 7070
rect 8670 7030 8710 7035
rect 8670 7000 8675 7030
rect 8675 7000 8705 7030
rect 8705 7000 8710 7030
rect 8670 6995 8710 7000
rect 8670 6960 8710 6965
rect 8670 6930 8675 6960
rect 8675 6930 8705 6960
rect 8705 6930 8710 6960
rect 8670 6925 8710 6930
rect 8670 6895 8710 6900
rect 8670 6865 8675 6895
rect 8675 6865 8705 6895
rect 8705 6865 8710 6895
rect 8670 6860 8710 6865
rect 8670 6835 8710 6840
rect 8670 6805 8675 6835
rect 8675 6805 8705 6835
rect 8705 6805 8710 6835
rect 8670 6800 8710 6805
rect 8670 6770 8710 6775
rect 8670 6740 8675 6770
rect 8675 6740 8705 6770
rect 8705 6740 8710 6770
rect 8670 6735 8710 6740
rect 8670 6700 8710 6705
rect 8670 6670 8675 6700
rect 8675 6670 8705 6700
rect 8705 6670 8710 6700
rect 8670 6665 8710 6670
rect 8670 6630 8710 6635
rect 8670 6600 8675 6630
rect 8675 6600 8705 6630
rect 8705 6600 8710 6630
rect 8670 6595 8710 6600
rect 8670 6560 8710 6565
rect 8670 6530 8675 6560
rect 8675 6530 8705 6560
rect 8705 6530 8710 6560
rect 8670 6525 8710 6530
rect 8670 6495 8710 6500
rect 8670 6465 8675 6495
rect 8675 6465 8705 6495
rect 8705 6465 8710 6495
rect 8670 6460 8710 6465
rect 9020 9635 9060 9640
rect 9020 9605 9025 9635
rect 9025 9605 9055 9635
rect 9055 9605 9060 9635
rect 9020 9600 9060 9605
rect 9020 9570 9060 9575
rect 9020 9540 9025 9570
rect 9025 9540 9055 9570
rect 9055 9540 9060 9570
rect 9020 9535 9060 9540
rect 9020 9500 9060 9505
rect 9020 9470 9025 9500
rect 9025 9470 9055 9500
rect 9055 9470 9060 9500
rect 9020 9465 9060 9470
rect 9020 9430 9060 9435
rect 9020 9400 9025 9430
rect 9025 9400 9055 9430
rect 9055 9400 9060 9430
rect 9020 9395 9060 9400
rect 9020 9360 9060 9365
rect 9020 9330 9025 9360
rect 9025 9330 9055 9360
rect 9055 9330 9060 9360
rect 9020 9325 9060 9330
rect 9020 9295 9060 9300
rect 9020 9265 9025 9295
rect 9025 9265 9055 9295
rect 9055 9265 9060 9295
rect 9020 9260 9060 9265
rect 9020 9235 9060 9240
rect 9020 9205 9025 9235
rect 9025 9205 9055 9235
rect 9055 9205 9060 9235
rect 9020 9200 9060 9205
rect 9020 9170 9060 9175
rect 9020 9140 9025 9170
rect 9025 9140 9055 9170
rect 9055 9140 9060 9170
rect 9020 9135 9060 9140
rect 9020 9100 9060 9105
rect 9020 9070 9025 9100
rect 9025 9070 9055 9100
rect 9055 9070 9060 9100
rect 9020 9065 9060 9070
rect 9020 9030 9060 9035
rect 9020 9000 9025 9030
rect 9025 9000 9055 9030
rect 9055 9000 9060 9030
rect 9020 8995 9060 9000
rect 9020 8960 9060 8965
rect 9020 8930 9025 8960
rect 9025 8930 9055 8960
rect 9055 8930 9060 8960
rect 9020 8925 9060 8930
rect 9020 8895 9060 8900
rect 9020 8865 9025 8895
rect 9025 8865 9055 8895
rect 9055 8865 9060 8895
rect 9020 8860 9060 8865
rect 9020 8835 9060 8840
rect 9020 8805 9025 8835
rect 9025 8805 9055 8835
rect 9055 8805 9060 8835
rect 9020 8800 9060 8805
rect 9020 8770 9060 8775
rect 9020 8740 9025 8770
rect 9025 8740 9055 8770
rect 9055 8740 9060 8770
rect 9020 8735 9060 8740
rect 9020 8700 9060 8705
rect 9020 8670 9025 8700
rect 9025 8670 9055 8700
rect 9055 8670 9060 8700
rect 9020 8665 9060 8670
rect 9020 8630 9060 8635
rect 9020 8600 9025 8630
rect 9025 8600 9055 8630
rect 9055 8600 9060 8630
rect 9020 8595 9060 8600
rect 9020 8560 9060 8565
rect 9020 8530 9025 8560
rect 9025 8530 9055 8560
rect 9055 8530 9060 8560
rect 9020 8525 9060 8530
rect 9020 8495 9060 8500
rect 9020 8465 9025 8495
rect 9025 8465 9055 8495
rect 9055 8465 9060 8495
rect 9020 8460 9060 8465
rect 9020 8435 9060 8440
rect 9020 8405 9025 8435
rect 9025 8405 9055 8435
rect 9055 8405 9060 8435
rect 9020 8400 9060 8405
rect 9020 8370 9060 8375
rect 9020 8340 9025 8370
rect 9025 8340 9055 8370
rect 9055 8340 9060 8370
rect 9020 8335 9060 8340
rect 9020 8300 9060 8305
rect 9020 8270 9025 8300
rect 9025 8270 9055 8300
rect 9055 8270 9060 8300
rect 9020 8265 9060 8270
rect 9020 8230 9060 8235
rect 9020 8200 9025 8230
rect 9025 8200 9055 8230
rect 9055 8200 9060 8230
rect 9020 8195 9060 8200
rect 9020 8160 9060 8165
rect 9020 8130 9025 8160
rect 9025 8130 9055 8160
rect 9055 8130 9060 8160
rect 9020 8125 9060 8130
rect 9020 8095 9060 8100
rect 9020 8065 9025 8095
rect 9025 8065 9055 8095
rect 9055 8065 9060 8095
rect 9020 8060 9060 8065
rect 9020 8035 9060 8040
rect 9020 8005 9025 8035
rect 9025 8005 9055 8035
rect 9055 8005 9060 8035
rect 9020 8000 9060 8005
rect 9020 7970 9060 7975
rect 9020 7940 9025 7970
rect 9025 7940 9055 7970
rect 9055 7940 9060 7970
rect 9020 7935 9060 7940
rect 9020 7900 9060 7905
rect 9020 7870 9025 7900
rect 9025 7870 9055 7900
rect 9055 7870 9060 7900
rect 9020 7865 9060 7870
rect 9020 7830 9060 7835
rect 9020 7800 9025 7830
rect 9025 7800 9055 7830
rect 9055 7800 9060 7830
rect 9020 7795 9060 7800
rect 9020 7760 9060 7765
rect 9020 7730 9025 7760
rect 9025 7730 9055 7760
rect 9055 7730 9060 7760
rect 9020 7725 9060 7730
rect 9020 7695 9060 7700
rect 9020 7665 9025 7695
rect 9025 7665 9055 7695
rect 9055 7665 9060 7695
rect 9020 7660 9060 7665
rect 9020 7635 9060 7640
rect 9020 7605 9025 7635
rect 9025 7605 9055 7635
rect 9055 7605 9060 7635
rect 9020 7600 9060 7605
rect 9020 7570 9060 7575
rect 9020 7540 9025 7570
rect 9025 7540 9055 7570
rect 9055 7540 9060 7570
rect 9020 7535 9060 7540
rect 9020 7500 9060 7505
rect 9020 7470 9025 7500
rect 9025 7470 9055 7500
rect 9055 7470 9060 7500
rect 9020 7465 9060 7470
rect 9020 7430 9060 7435
rect 9020 7400 9025 7430
rect 9025 7400 9055 7430
rect 9055 7400 9060 7430
rect 9020 7395 9060 7400
rect 9020 7360 9060 7365
rect 9020 7330 9025 7360
rect 9025 7330 9055 7360
rect 9055 7330 9060 7360
rect 9020 7325 9060 7330
rect 9020 7295 9060 7300
rect 9020 7265 9025 7295
rect 9025 7265 9055 7295
rect 9055 7265 9060 7295
rect 9020 7260 9060 7265
rect 9020 7235 9060 7240
rect 9020 7205 9025 7235
rect 9025 7205 9055 7235
rect 9055 7205 9060 7235
rect 9020 7200 9060 7205
rect 9020 7170 9060 7175
rect 9020 7140 9025 7170
rect 9025 7140 9055 7170
rect 9055 7140 9060 7170
rect 9020 7135 9060 7140
rect 9020 7100 9060 7105
rect 9020 7070 9025 7100
rect 9025 7070 9055 7100
rect 9055 7070 9060 7100
rect 9020 7065 9060 7070
rect 9020 7030 9060 7035
rect 9020 7000 9025 7030
rect 9025 7000 9055 7030
rect 9055 7000 9060 7030
rect 9020 6995 9060 7000
rect 9020 6960 9060 6965
rect 9020 6930 9025 6960
rect 9025 6930 9055 6960
rect 9055 6930 9060 6960
rect 9020 6925 9060 6930
rect 9020 6895 9060 6900
rect 9020 6865 9025 6895
rect 9025 6865 9055 6895
rect 9055 6865 9060 6895
rect 9020 6860 9060 6865
rect 9020 6835 9060 6840
rect 9020 6805 9025 6835
rect 9025 6805 9055 6835
rect 9055 6805 9060 6835
rect 9020 6800 9060 6805
rect 9020 6770 9060 6775
rect 9020 6740 9025 6770
rect 9025 6740 9055 6770
rect 9055 6740 9060 6770
rect 9020 6735 9060 6740
rect 9020 6700 9060 6705
rect 9020 6670 9025 6700
rect 9025 6670 9055 6700
rect 9055 6670 9060 6700
rect 9020 6665 9060 6670
rect 9020 6630 9060 6635
rect 9020 6600 9025 6630
rect 9025 6600 9055 6630
rect 9055 6600 9060 6630
rect 9020 6595 9060 6600
rect 9020 6560 9060 6565
rect 9020 6530 9025 6560
rect 9025 6530 9055 6560
rect 9055 6530 9060 6560
rect 9020 6525 9060 6530
rect 9020 6495 9060 6500
rect 9020 6465 9025 6495
rect 9025 6465 9055 6495
rect 9055 6465 9060 6495
rect 9020 6460 9060 6465
rect 31305 7995 31340 8030
rect 31350 7995 31385 8030
rect 31395 7995 31430 8030
rect 31440 7995 31475 8030
rect 31485 7995 31520 8030
rect 31530 7995 31565 8030
rect 31575 7995 31610 8030
rect 31620 7995 31655 8030
rect 31665 7995 31700 8030
rect 31710 7995 31745 8030
rect 31755 7995 31790 8030
rect 31800 7995 31835 8030
rect 31845 7995 31880 8030
rect 31890 7995 31925 8030
rect 31935 7995 31970 8030
rect 31980 7995 32015 8030
rect 32025 7995 32060 8030
rect 32070 7995 32105 8030
rect 32115 7995 32150 8030
rect 32160 7995 32195 8030
rect 32205 7995 32240 8030
rect 32250 7995 32285 8030
rect 32295 7995 32330 8030
rect 32340 7995 32375 8030
rect 32385 7995 32420 8030
rect 32430 7995 32465 8030
rect 32475 7995 32510 8030
rect 32520 7995 32555 8030
rect 32565 7995 32600 8030
rect 32610 7995 32645 8030
rect 32655 7995 32690 8030
rect 32700 7995 32735 8030
rect 32745 7995 32780 8030
rect 32790 7995 32825 8030
rect 32835 7995 32870 8030
rect 31305 7950 31340 7985
rect 31350 7950 31385 7985
rect 31395 7950 31430 7985
rect 31440 7950 31475 7985
rect 31485 7950 31520 7985
rect 31530 7950 31565 7985
rect 31575 7950 31610 7985
rect 31620 7950 31655 7985
rect 31665 7950 31700 7985
rect 31710 7950 31745 7985
rect 31755 7950 31790 7985
rect 31800 7950 31835 7985
rect 31845 7950 31880 7985
rect 31890 7950 31925 7985
rect 31935 7950 31970 7985
rect 31980 7950 32015 7985
rect 32025 7950 32060 7985
rect 32070 7950 32105 7985
rect 32115 7950 32150 7985
rect 32160 7950 32195 7985
rect 32205 7950 32240 7985
rect 32250 7950 32285 7985
rect 32295 7950 32330 7985
rect 32340 7950 32375 7985
rect 32385 7950 32420 7985
rect 32430 7950 32465 7985
rect 32475 7950 32510 7985
rect 32520 7950 32555 7985
rect 32565 7950 32600 7985
rect 32610 7950 32645 7985
rect 32655 7950 32690 7985
rect 32700 7950 32735 7985
rect 32745 7950 32780 7985
rect 32790 7950 32825 7985
rect 32835 7950 32870 7985
rect 31305 7905 31340 7940
rect 31350 7905 31385 7940
rect 31395 7905 31430 7940
rect 31440 7905 31475 7940
rect 31485 7905 31520 7940
rect 31530 7905 31565 7940
rect 31575 7905 31610 7940
rect 31620 7905 31655 7940
rect 31665 7905 31700 7940
rect 31710 7905 31745 7940
rect 31755 7905 31790 7940
rect 31800 7905 31835 7940
rect 31845 7905 31880 7940
rect 31890 7905 31925 7940
rect 31935 7905 31970 7940
rect 31980 7905 32015 7940
rect 32025 7905 32060 7940
rect 32070 7905 32105 7940
rect 32115 7905 32150 7940
rect 32160 7905 32195 7940
rect 32205 7905 32240 7940
rect 32250 7905 32285 7940
rect 32295 7905 32330 7940
rect 32340 7905 32375 7940
rect 32385 7905 32420 7940
rect 32430 7905 32465 7940
rect 32475 7905 32510 7940
rect 32520 7905 32555 7940
rect 32565 7905 32600 7940
rect 32610 7905 32645 7940
rect 32655 7905 32690 7940
rect 32700 7905 32735 7940
rect 32745 7905 32780 7940
rect 32790 7905 32825 7940
rect 32835 7905 32870 7940
rect 31305 7860 31340 7895
rect 31350 7860 31385 7895
rect 31395 7860 31430 7895
rect 31440 7860 31475 7895
rect 31485 7860 31520 7895
rect 31530 7860 31565 7895
rect 31575 7860 31610 7895
rect 31620 7860 31655 7895
rect 31665 7860 31700 7895
rect 31710 7860 31745 7895
rect 31755 7860 31790 7895
rect 31800 7860 31835 7895
rect 31845 7860 31880 7895
rect 31890 7860 31925 7895
rect 31935 7860 31970 7895
rect 31980 7860 32015 7895
rect 32025 7860 32060 7895
rect 32070 7860 32105 7895
rect 32115 7860 32150 7895
rect 32160 7860 32195 7895
rect 32205 7860 32240 7895
rect 32250 7860 32285 7895
rect 32295 7860 32330 7895
rect 32340 7860 32375 7895
rect 32385 7860 32420 7895
rect 32430 7860 32465 7895
rect 32475 7860 32510 7895
rect 32520 7860 32555 7895
rect 32565 7860 32600 7895
rect 32610 7860 32645 7895
rect 32655 7860 32690 7895
rect 32700 7860 32735 7895
rect 32745 7860 32780 7895
rect 32790 7860 32825 7895
rect 32835 7860 32870 7895
rect 31305 7815 31340 7850
rect 31350 7815 31385 7850
rect 31395 7815 31430 7850
rect 31440 7815 31475 7850
rect 31485 7815 31520 7850
rect 31530 7815 31565 7850
rect 31575 7815 31610 7850
rect 31620 7815 31655 7850
rect 31665 7815 31700 7850
rect 31710 7815 31745 7850
rect 31755 7815 31790 7850
rect 31800 7815 31835 7850
rect 31845 7815 31880 7850
rect 31890 7815 31925 7850
rect 31935 7815 31970 7850
rect 31980 7815 32015 7850
rect 32025 7815 32060 7850
rect 32070 7815 32105 7850
rect 32115 7815 32150 7850
rect 32160 7815 32195 7850
rect 32205 7815 32240 7850
rect 32250 7815 32285 7850
rect 32295 7815 32330 7850
rect 32340 7815 32375 7850
rect 32385 7815 32420 7850
rect 32430 7815 32465 7850
rect 32475 7815 32510 7850
rect 32520 7815 32555 7850
rect 32565 7815 32600 7850
rect 32610 7815 32645 7850
rect 32655 7815 32690 7850
rect 32700 7815 32735 7850
rect 32745 7815 32780 7850
rect 32790 7815 32825 7850
rect 32835 7815 32870 7850
rect 31305 7770 31340 7805
rect 31350 7770 31385 7805
rect 31395 7770 31430 7805
rect 31440 7770 31475 7805
rect 31485 7770 31520 7805
rect 31530 7770 31565 7805
rect 31575 7770 31610 7805
rect 31620 7770 31655 7805
rect 31665 7770 31700 7805
rect 31710 7770 31745 7805
rect 31755 7770 31790 7805
rect 31800 7770 31835 7805
rect 31845 7770 31880 7805
rect 31890 7770 31925 7805
rect 31935 7770 31970 7805
rect 31980 7770 32015 7805
rect 32025 7770 32060 7805
rect 32070 7770 32105 7805
rect 32115 7770 32150 7805
rect 32160 7770 32195 7805
rect 32205 7770 32240 7805
rect 32250 7770 32285 7805
rect 32295 7770 32330 7805
rect 32340 7770 32375 7805
rect 32385 7770 32420 7805
rect 32430 7770 32465 7805
rect 32475 7770 32510 7805
rect 32520 7770 32555 7805
rect 32565 7770 32600 7805
rect 32610 7770 32645 7805
rect 32655 7770 32690 7805
rect 32700 7770 32735 7805
rect 32745 7770 32780 7805
rect 32790 7770 32825 7805
rect 32835 7770 32870 7805
rect 31305 7725 31340 7760
rect 31350 7725 31385 7760
rect 31395 7725 31430 7760
rect 31440 7725 31475 7760
rect 31485 7725 31520 7760
rect 31530 7725 31565 7760
rect 31575 7725 31610 7760
rect 31620 7725 31655 7760
rect 31665 7725 31700 7760
rect 31710 7725 31745 7760
rect 31755 7725 31790 7760
rect 31800 7725 31835 7760
rect 31845 7725 31880 7760
rect 31890 7725 31925 7760
rect 31935 7725 31970 7760
rect 31980 7725 32015 7760
rect 32025 7725 32060 7760
rect 32070 7725 32105 7760
rect 32115 7725 32150 7760
rect 32160 7725 32195 7760
rect 32205 7725 32240 7760
rect 32250 7725 32285 7760
rect 32295 7725 32330 7760
rect 32340 7725 32375 7760
rect 32385 7725 32420 7760
rect 32430 7725 32465 7760
rect 32475 7725 32510 7760
rect 32520 7725 32555 7760
rect 32565 7725 32600 7760
rect 32610 7725 32645 7760
rect 32655 7725 32690 7760
rect 32700 7725 32735 7760
rect 32745 7725 32780 7760
rect 32790 7725 32825 7760
rect 32835 7725 32870 7760
rect 31305 7680 31340 7715
rect 31350 7680 31385 7715
rect 31395 7680 31430 7715
rect 31440 7680 31475 7715
rect 31485 7680 31520 7715
rect 31530 7680 31565 7715
rect 31575 7680 31610 7715
rect 31620 7680 31655 7715
rect 31665 7680 31700 7715
rect 31710 7680 31745 7715
rect 31755 7680 31790 7715
rect 31800 7680 31835 7715
rect 31845 7680 31880 7715
rect 31890 7680 31925 7715
rect 31935 7680 31970 7715
rect 31980 7680 32015 7715
rect 32025 7680 32060 7715
rect 32070 7680 32105 7715
rect 32115 7680 32150 7715
rect 32160 7680 32195 7715
rect 32205 7680 32240 7715
rect 32250 7680 32285 7715
rect 32295 7680 32330 7715
rect 32340 7680 32375 7715
rect 32385 7680 32420 7715
rect 32430 7680 32465 7715
rect 32475 7680 32510 7715
rect 32520 7680 32555 7715
rect 32565 7680 32600 7715
rect 32610 7680 32645 7715
rect 32655 7680 32690 7715
rect 32700 7680 32735 7715
rect 32745 7680 32780 7715
rect 32790 7680 32825 7715
rect 32835 7680 32870 7715
rect 31305 7635 31340 7670
rect 31350 7635 31385 7670
rect 31395 7635 31430 7670
rect 31440 7635 31475 7670
rect 31485 7635 31520 7670
rect 31530 7635 31565 7670
rect 31575 7635 31610 7670
rect 31620 7635 31655 7670
rect 31665 7635 31700 7670
rect 31710 7635 31745 7670
rect 31755 7635 31790 7670
rect 31800 7635 31835 7670
rect 31845 7635 31880 7670
rect 31890 7635 31925 7670
rect 31935 7635 31970 7670
rect 31980 7635 32015 7670
rect 32025 7635 32060 7670
rect 32070 7635 32105 7670
rect 32115 7635 32150 7670
rect 32160 7635 32195 7670
rect 32205 7635 32240 7670
rect 32250 7635 32285 7670
rect 32295 7635 32330 7670
rect 32340 7635 32375 7670
rect 32385 7635 32420 7670
rect 32430 7635 32465 7670
rect 32475 7635 32510 7670
rect 32520 7635 32555 7670
rect 32565 7635 32600 7670
rect 32610 7635 32645 7670
rect 32655 7635 32690 7670
rect 32700 7635 32735 7670
rect 32745 7635 32780 7670
rect 32790 7635 32825 7670
rect 32835 7635 32870 7670
rect 31305 7590 31340 7625
rect 31350 7590 31385 7625
rect 31395 7590 31430 7625
rect 31440 7590 31475 7625
rect 31485 7590 31520 7625
rect 31530 7590 31565 7625
rect 31575 7590 31610 7625
rect 31620 7590 31655 7625
rect 31665 7590 31700 7625
rect 31710 7590 31745 7625
rect 31755 7590 31790 7625
rect 31800 7590 31835 7625
rect 31845 7590 31880 7625
rect 31890 7590 31925 7625
rect 31935 7590 31970 7625
rect 31980 7590 32015 7625
rect 32025 7590 32060 7625
rect 32070 7590 32105 7625
rect 32115 7590 32150 7625
rect 32160 7590 32195 7625
rect 32205 7590 32240 7625
rect 32250 7590 32285 7625
rect 32295 7590 32330 7625
rect 32340 7590 32375 7625
rect 32385 7590 32420 7625
rect 32430 7590 32465 7625
rect 32475 7590 32510 7625
rect 32520 7590 32555 7625
rect 32565 7590 32600 7625
rect 32610 7590 32645 7625
rect 32655 7590 32690 7625
rect 32700 7590 32735 7625
rect 32745 7590 32780 7625
rect 32790 7590 32825 7625
rect 32835 7590 32870 7625
rect 31305 7545 31340 7580
rect 31350 7545 31385 7580
rect 31395 7545 31430 7580
rect 31440 7545 31475 7580
rect 31485 7545 31520 7580
rect 31530 7545 31565 7580
rect 31575 7545 31610 7580
rect 31620 7545 31655 7580
rect 31665 7545 31700 7580
rect 31710 7545 31745 7580
rect 31755 7545 31790 7580
rect 31800 7545 31835 7580
rect 31845 7545 31880 7580
rect 31890 7545 31925 7580
rect 31935 7545 31970 7580
rect 31980 7545 32015 7580
rect 32025 7545 32060 7580
rect 32070 7545 32105 7580
rect 32115 7545 32150 7580
rect 32160 7545 32195 7580
rect 32205 7545 32240 7580
rect 32250 7545 32285 7580
rect 32295 7545 32330 7580
rect 32340 7545 32375 7580
rect 32385 7545 32420 7580
rect 32430 7545 32465 7580
rect 32475 7545 32510 7580
rect 32520 7545 32555 7580
rect 32565 7545 32600 7580
rect 32610 7545 32645 7580
rect 32655 7545 32690 7580
rect 32700 7545 32735 7580
rect 32745 7545 32780 7580
rect 32790 7545 32825 7580
rect 32835 7545 32870 7580
rect 31305 7500 31340 7535
rect 31350 7500 31385 7535
rect 31395 7500 31430 7535
rect 31440 7500 31475 7535
rect 31485 7500 31520 7535
rect 31530 7500 31565 7535
rect 31575 7500 31610 7535
rect 31620 7500 31655 7535
rect 31665 7500 31700 7535
rect 31710 7500 31745 7535
rect 31755 7500 31790 7535
rect 31800 7500 31835 7535
rect 31845 7500 31880 7535
rect 31890 7500 31925 7535
rect 31935 7500 31970 7535
rect 31980 7500 32015 7535
rect 32025 7500 32060 7535
rect 32070 7500 32105 7535
rect 32115 7500 32150 7535
rect 32160 7500 32195 7535
rect 32205 7500 32240 7535
rect 32250 7500 32285 7535
rect 32295 7500 32330 7535
rect 32340 7500 32375 7535
rect 32385 7500 32420 7535
rect 32430 7500 32465 7535
rect 32475 7500 32510 7535
rect 32520 7500 32555 7535
rect 32565 7500 32600 7535
rect 32610 7500 32645 7535
rect 32655 7500 32690 7535
rect 32700 7500 32735 7535
rect 32745 7500 32780 7535
rect 32790 7500 32825 7535
rect 32835 7500 32870 7535
rect 31305 7455 31340 7490
rect 31350 7455 31385 7490
rect 31395 7455 31430 7490
rect 31440 7455 31475 7490
rect 31485 7455 31520 7490
rect 31530 7455 31565 7490
rect 31575 7455 31610 7490
rect 31620 7455 31655 7490
rect 31665 7455 31700 7490
rect 31710 7455 31745 7490
rect 31755 7455 31790 7490
rect 31800 7455 31835 7490
rect 31845 7455 31880 7490
rect 31890 7455 31925 7490
rect 31935 7455 31970 7490
rect 31980 7455 32015 7490
rect 32025 7455 32060 7490
rect 32070 7455 32105 7490
rect 32115 7455 32150 7490
rect 32160 7455 32195 7490
rect 32205 7455 32240 7490
rect 32250 7455 32285 7490
rect 32295 7455 32330 7490
rect 32340 7455 32375 7490
rect 32385 7455 32420 7490
rect 32430 7455 32465 7490
rect 32475 7455 32510 7490
rect 32520 7455 32555 7490
rect 32565 7455 32600 7490
rect 32610 7455 32645 7490
rect 32655 7455 32690 7490
rect 32700 7455 32735 7490
rect 32745 7455 32780 7490
rect 32790 7455 32825 7490
rect 32835 7455 32870 7490
rect 31305 7410 31340 7445
rect 31350 7410 31385 7445
rect 31395 7410 31430 7445
rect 31440 7410 31475 7445
rect 31485 7410 31520 7445
rect 31530 7410 31565 7445
rect 31575 7410 31610 7445
rect 31620 7410 31655 7445
rect 31665 7410 31700 7445
rect 31710 7410 31745 7445
rect 31755 7410 31790 7445
rect 31800 7410 31835 7445
rect 31845 7410 31880 7445
rect 31890 7410 31925 7445
rect 31935 7410 31970 7445
rect 31980 7410 32015 7445
rect 32025 7410 32060 7445
rect 32070 7410 32105 7445
rect 32115 7410 32150 7445
rect 32160 7410 32195 7445
rect 32205 7410 32240 7445
rect 32250 7410 32285 7445
rect 32295 7410 32330 7445
rect 32340 7410 32375 7445
rect 32385 7410 32420 7445
rect 32430 7410 32465 7445
rect 32475 7410 32510 7445
rect 32520 7410 32555 7445
rect 32565 7410 32600 7445
rect 32610 7410 32645 7445
rect 32655 7410 32690 7445
rect 32700 7410 32735 7445
rect 32745 7410 32780 7445
rect 32790 7410 32825 7445
rect 32835 7410 32870 7445
rect 31305 7365 31340 7400
rect 31350 7365 31385 7400
rect 31395 7365 31430 7400
rect 31440 7365 31475 7400
rect 31485 7365 31520 7400
rect 31530 7365 31565 7400
rect 31575 7365 31610 7400
rect 31620 7365 31655 7400
rect 31665 7365 31700 7400
rect 31710 7365 31745 7400
rect 31755 7365 31790 7400
rect 31800 7365 31835 7400
rect 31845 7365 31880 7400
rect 31890 7365 31925 7400
rect 31935 7365 31970 7400
rect 31980 7365 32015 7400
rect 32025 7365 32060 7400
rect 32070 7365 32105 7400
rect 32115 7365 32150 7400
rect 32160 7365 32195 7400
rect 32205 7365 32240 7400
rect 32250 7365 32285 7400
rect 32295 7365 32330 7400
rect 32340 7365 32375 7400
rect 32385 7365 32420 7400
rect 32430 7365 32465 7400
rect 32475 7365 32510 7400
rect 32520 7365 32555 7400
rect 32565 7365 32600 7400
rect 32610 7365 32645 7400
rect 32655 7365 32690 7400
rect 32700 7365 32735 7400
rect 32745 7365 32780 7400
rect 32790 7365 32825 7400
rect 32835 7365 32870 7400
rect 31305 7320 31340 7355
rect 31350 7320 31385 7355
rect 31395 7320 31430 7355
rect 31440 7320 31475 7355
rect 31485 7320 31520 7355
rect 31530 7320 31565 7355
rect 31575 7320 31610 7355
rect 31620 7320 31655 7355
rect 31665 7320 31700 7355
rect 31710 7320 31745 7355
rect 31755 7320 31790 7355
rect 31800 7320 31835 7355
rect 31845 7320 31880 7355
rect 31890 7320 31925 7355
rect 31935 7320 31970 7355
rect 31980 7320 32015 7355
rect 32025 7320 32060 7355
rect 32070 7320 32105 7355
rect 32115 7320 32150 7355
rect 32160 7320 32195 7355
rect 32205 7320 32240 7355
rect 32250 7320 32285 7355
rect 32295 7320 32330 7355
rect 32340 7320 32375 7355
rect 32385 7320 32420 7355
rect 32430 7320 32465 7355
rect 32475 7320 32510 7355
rect 32520 7320 32555 7355
rect 32565 7320 32600 7355
rect 32610 7320 32645 7355
rect 32655 7320 32690 7355
rect 32700 7320 32735 7355
rect 32745 7320 32780 7355
rect 32790 7320 32825 7355
rect 32835 7320 32870 7355
rect 31305 7275 31340 7310
rect 31350 7275 31385 7310
rect 31395 7275 31430 7310
rect 31440 7275 31475 7310
rect 31485 7275 31520 7310
rect 31530 7275 31565 7310
rect 31575 7275 31610 7310
rect 31620 7275 31655 7310
rect 31665 7275 31700 7310
rect 31710 7275 31745 7310
rect 31755 7275 31790 7310
rect 31800 7275 31835 7310
rect 31845 7275 31880 7310
rect 31890 7275 31925 7310
rect 31935 7275 31970 7310
rect 31980 7275 32015 7310
rect 32025 7275 32060 7310
rect 32070 7275 32105 7310
rect 32115 7275 32150 7310
rect 32160 7275 32195 7310
rect 32205 7275 32240 7310
rect 32250 7275 32285 7310
rect 32295 7275 32330 7310
rect 32340 7275 32375 7310
rect 32385 7275 32420 7310
rect 32430 7275 32465 7310
rect 32475 7275 32510 7310
rect 32520 7275 32555 7310
rect 32565 7275 32600 7310
rect 32610 7275 32645 7310
rect 32655 7275 32690 7310
rect 32700 7275 32735 7310
rect 32745 7275 32780 7310
rect 32790 7275 32825 7310
rect 32835 7275 32870 7310
rect 31305 7230 31340 7265
rect 31350 7230 31385 7265
rect 31395 7230 31430 7265
rect 31440 7230 31475 7265
rect 31485 7230 31520 7265
rect 31530 7230 31565 7265
rect 31575 7230 31610 7265
rect 31620 7230 31655 7265
rect 31665 7230 31700 7265
rect 31710 7230 31745 7265
rect 31755 7230 31790 7265
rect 31800 7230 31835 7265
rect 31845 7230 31880 7265
rect 31890 7230 31925 7265
rect 31935 7230 31970 7265
rect 31980 7230 32015 7265
rect 32025 7230 32060 7265
rect 32070 7230 32105 7265
rect 32115 7230 32150 7265
rect 32160 7230 32195 7265
rect 32205 7230 32240 7265
rect 32250 7230 32285 7265
rect 32295 7230 32330 7265
rect 32340 7230 32375 7265
rect 32385 7230 32420 7265
rect 32430 7230 32465 7265
rect 32475 7230 32510 7265
rect 32520 7230 32555 7265
rect 32565 7230 32600 7265
rect 32610 7230 32645 7265
rect 32655 7230 32690 7265
rect 32700 7230 32735 7265
rect 32745 7230 32780 7265
rect 32790 7230 32825 7265
rect 32835 7230 32870 7265
rect 31305 7185 31340 7220
rect 31350 7185 31385 7220
rect 31395 7185 31430 7220
rect 31440 7185 31475 7220
rect 31485 7185 31520 7220
rect 31530 7185 31565 7220
rect 31575 7185 31610 7220
rect 31620 7185 31655 7220
rect 31665 7185 31700 7220
rect 31710 7185 31745 7220
rect 31755 7185 31790 7220
rect 31800 7185 31835 7220
rect 31845 7185 31880 7220
rect 31890 7185 31925 7220
rect 31935 7185 31970 7220
rect 31980 7185 32015 7220
rect 32025 7185 32060 7220
rect 32070 7185 32105 7220
rect 32115 7185 32150 7220
rect 32160 7185 32195 7220
rect 32205 7185 32240 7220
rect 32250 7185 32285 7220
rect 32295 7185 32330 7220
rect 32340 7185 32375 7220
rect 32385 7185 32420 7220
rect 32430 7185 32465 7220
rect 32475 7185 32510 7220
rect 32520 7185 32555 7220
rect 32565 7185 32600 7220
rect 32610 7185 32645 7220
rect 32655 7185 32690 7220
rect 32700 7185 32735 7220
rect 32745 7185 32780 7220
rect 32790 7185 32825 7220
rect 32835 7185 32870 7220
rect 31305 7140 31340 7175
rect 31350 7140 31385 7175
rect 31395 7140 31430 7175
rect 31440 7140 31475 7175
rect 31485 7140 31520 7175
rect 31530 7140 31565 7175
rect 31575 7140 31610 7175
rect 31620 7140 31655 7175
rect 31665 7140 31700 7175
rect 31710 7140 31745 7175
rect 31755 7140 31790 7175
rect 31800 7140 31835 7175
rect 31845 7140 31880 7175
rect 31890 7140 31925 7175
rect 31935 7140 31970 7175
rect 31980 7140 32015 7175
rect 32025 7140 32060 7175
rect 32070 7140 32105 7175
rect 32115 7140 32150 7175
rect 32160 7140 32195 7175
rect 32205 7140 32240 7175
rect 32250 7140 32285 7175
rect 32295 7140 32330 7175
rect 32340 7140 32375 7175
rect 32385 7140 32420 7175
rect 32430 7140 32465 7175
rect 32475 7140 32510 7175
rect 32520 7140 32555 7175
rect 32565 7140 32600 7175
rect 32610 7140 32645 7175
rect 32655 7140 32690 7175
rect 32700 7140 32735 7175
rect 32745 7140 32780 7175
rect 32790 7140 32825 7175
rect 32835 7140 32870 7175
rect 31305 7095 31340 7130
rect 31350 7095 31385 7130
rect 31395 7095 31430 7130
rect 31440 7095 31475 7130
rect 31485 7095 31520 7130
rect 31530 7095 31565 7130
rect 31575 7095 31610 7130
rect 31620 7095 31655 7130
rect 31665 7095 31700 7130
rect 31710 7095 31745 7130
rect 31755 7095 31790 7130
rect 31800 7095 31835 7130
rect 31845 7095 31880 7130
rect 31890 7095 31925 7130
rect 31935 7095 31970 7130
rect 31980 7095 32015 7130
rect 32025 7095 32060 7130
rect 32070 7095 32105 7130
rect 32115 7095 32150 7130
rect 32160 7095 32195 7130
rect 32205 7095 32240 7130
rect 32250 7095 32285 7130
rect 32295 7095 32330 7130
rect 32340 7095 32375 7130
rect 32385 7095 32420 7130
rect 32430 7095 32465 7130
rect 32475 7095 32510 7130
rect 32520 7095 32555 7130
rect 32565 7095 32600 7130
rect 32610 7095 32645 7130
rect 32655 7095 32690 7130
rect 32700 7095 32735 7130
rect 32745 7095 32780 7130
rect 32790 7095 32825 7130
rect 32835 7095 32870 7130
rect 31305 7050 31340 7085
rect 31350 7050 31385 7085
rect 31395 7050 31430 7085
rect 31440 7050 31475 7085
rect 31485 7050 31520 7085
rect 31530 7050 31565 7085
rect 31575 7050 31610 7085
rect 31620 7050 31655 7085
rect 31665 7050 31700 7085
rect 31710 7050 31745 7085
rect 31755 7050 31790 7085
rect 31800 7050 31835 7085
rect 31845 7050 31880 7085
rect 31890 7050 31925 7085
rect 31935 7050 31970 7085
rect 31980 7050 32015 7085
rect 32025 7050 32060 7085
rect 32070 7050 32105 7085
rect 32115 7050 32150 7085
rect 32160 7050 32195 7085
rect 32205 7050 32240 7085
rect 32250 7050 32285 7085
rect 32295 7050 32330 7085
rect 32340 7050 32375 7085
rect 32385 7050 32420 7085
rect 32430 7050 32465 7085
rect 32475 7050 32510 7085
rect 32520 7050 32555 7085
rect 32565 7050 32600 7085
rect 32610 7050 32645 7085
rect 32655 7050 32690 7085
rect 32700 7050 32735 7085
rect 32745 7050 32780 7085
rect 32790 7050 32825 7085
rect 32835 7050 32870 7085
rect 31305 7005 31340 7040
rect 31350 7005 31385 7040
rect 31395 7005 31430 7040
rect 31440 7005 31475 7040
rect 31485 7005 31520 7040
rect 31530 7005 31565 7040
rect 31575 7005 31610 7040
rect 31620 7005 31655 7040
rect 31665 7005 31700 7040
rect 31710 7005 31745 7040
rect 31755 7005 31790 7040
rect 31800 7005 31835 7040
rect 31845 7005 31880 7040
rect 31890 7005 31925 7040
rect 31935 7005 31970 7040
rect 31980 7005 32015 7040
rect 32025 7005 32060 7040
rect 32070 7005 32105 7040
rect 32115 7005 32150 7040
rect 32160 7005 32195 7040
rect 32205 7005 32240 7040
rect 32250 7005 32285 7040
rect 32295 7005 32330 7040
rect 32340 7005 32375 7040
rect 32385 7005 32420 7040
rect 32430 7005 32465 7040
rect 32475 7005 32510 7040
rect 32520 7005 32555 7040
rect 32565 7005 32600 7040
rect 32610 7005 32645 7040
rect 32655 7005 32690 7040
rect 32700 7005 32735 7040
rect 32745 7005 32780 7040
rect 32790 7005 32825 7040
rect 32835 7005 32870 7040
rect 31305 6960 31340 6995
rect 31350 6960 31385 6995
rect 31395 6960 31430 6995
rect 31440 6960 31475 6995
rect 31485 6960 31520 6995
rect 31530 6960 31565 6995
rect 31575 6960 31610 6995
rect 31620 6960 31655 6995
rect 31665 6960 31700 6995
rect 31710 6960 31745 6995
rect 31755 6960 31790 6995
rect 31800 6960 31835 6995
rect 31845 6960 31880 6995
rect 31890 6960 31925 6995
rect 31935 6960 31970 6995
rect 31980 6960 32015 6995
rect 32025 6960 32060 6995
rect 32070 6960 32105 6995
rect 32115 6960 32150 6995
rect 32160 6960 32195 6995
rect 32205 6960 32240 6995
rect 32250 6960 32285 6995
rect 32295 6960 32330 6995
rect 32340 6960 32375 6995
rect 32385 6960 32420 6995
rect 32430 6960 32465 6995
rect 32475 6960 32510 6995
rect 32520 6960 32555 6995
rect 32565 6960 32600 6995
rect 32610 6960 32645 6995
rect 32655 6960 32690 6995
rect 32700 6960 32735 6995
rect 32745 6960 32780 6995
rect 32790 6960 32825 6995
rect 32835 6960 32870 6995
rect 31305 6915 31340 6950
rect 31350 6915 31385 6950
rect 31395 6915 31430 6950
rect 31440 6915 31475 6950
rect 31485 6915 31520 6950
rect 31530 6915 31565 6950
rect 31575 6915 31610 6950
rect 31620 6915 31655 6950
rect 31665 6915 31700 6950
rect 31710 6915 31745 6950
rect 31755 6915 31790 6950
rect 31800 6915 31835 6950
rect 31845 6915 31880 6950
rect 31890 6915 31925 6950
rect 31935 6915 31970 6950
rect 31980 6915 32015 6950
rect 32025 6915 32060 6950
rect 32070 6915 32105 6950
rect 32115 6915 32150 6950
rect 32160 6915 32195 6950
rect 32205 6915 32240 6950
rect 32250 6915 32285 6950
rect 32295 6915 32330 6950
rect 32340 6915 32375 6950
rect 32385 6915 32420 6950
rect 32430 6915 32465 6950
rect 32475 6915 32510 6950
rect 32520 6915 32555 6950
rect 32565 6915 32600 6950
rect 32610 6915 32645 6950
rect 32655 6915 32690 6950
rect 32700 6915 32735 6950
rect 32745 6915 32780 6950
rect 32790 6915 32825 6950
rect 32835 6915 32870 6950
rect 31305 6870 31340 6905
rect 31350 6870 31385 6905
rect 31395 6870 31430 6905
rect 31440 6870 31475 6905
rect 31485 6870 31520 6905
rect 31530 6870 31565 6905
rect 31575 6870 31610 6905
rect 31620 6870 31655 6905
rect 31665 6870 31700 6905
rect 31710 6870 31745 6905
rect 31755 6870 31790 6905
rect 31800 6870 31835 6905
rect 31845 6870 31880 6905
rect 31890 6870 31925 6905
rect 31935 6870 31970 6905
rect 31980 6870 32015 6905
rect 32025 6870 32060 6905
rect 32070 6870 32105 6905
rect 32115 6870 32150 6905
rect 32160 6870 32195 6905
rect 32205 6870 32240 6905
rect 32250 6870 32285 6905
rect 32295 6870 32330 6905
rect 32340 6870 32375 6905
rect 32385 6870 32420 6905
rect 32430 6870 32465 6905
rect 32475 6870 32510 6905
rect 32520 6870 32555 6905
rect 32565 6870 32600 6905
rect 32610 6870 32645 6905
rect 32655 6870 32690 6905
rect 32700 6870 32735 6905
rect 32745 6870 32780 6905
rect 32790 6870 32825 6905
rect 32835 6870 32870 6905
rect 31305 6825 31340 6860
rect 31350 6825 31385 6860
rect 31395 6825 31430 6860
rect 31440 6825 31475 6860
rect 31485 6825 31520 6860
rect 31530 6825 31565 6860
rect 31575 6825 31610 6860
rect 31620 6825 31655 6860
rect 31665 6825 31700 6860
rect 31710 6825 31745 6860
rect 31755 6825 31790 6860
rect 31800 6825 31835 6860
rect 31845 6825 31880 6860
rect 31890 6825 31925 6860
rect 31935 6825 31970 6860
rect 31980 6825 32015 6860
rect 32025 6825 32060 6860
rect 32070 6825 32105 6860
rect 32115 6825 32150 6860
rect 32160 6825 32195 6860
rect 32205 6825 32240 6860
rect 32250 6825 32285 6860
rect 32295 6825 32330 6860
rect 32340 6825 32375 6860
rect 32385 6825 32420 6860
rect 32430 6825 32465 6860
rect 32475 6825 32510 6860
rect 32520 6825 32555 6860
rect 32565 6825 32600 6860
rect 32610 6825 32645 6860
rect 32655 6825 32690 6860
rect 32700 6825 32735 6860
rect 32745 6825 32780 6860
rect 32790 6825 32825 6860
rect 32835 6825 32870 6860
rect 31305 6780 31340 6815
rect 31350 6780 31385 6815
rect 31395 6780 31430 6815
rect 31440 6780 31475 6815
rect 31485 6780 31520 6815
rect 31530 6780 31565 6815
rect 31575 6780 31610 6815
rect 31620 6780 31655 6815
rect 31665 6780 31700 6815
rect 31710 6780 31745 6815
rect 31755 6780 31790 6815
rect 31800 6780 31835 6815
rect 31845 6780 31880 6815
rect 31890 6780 31925 6815
rect 31935 6780 31970 6815
rect 31980 6780 32015 6815
rect 32025 6780 32060 6815
rect 32070 6780 32105 6815
rect 32115 6780 32150 6815
rect 32160 6780 32195 6815
rect 32205 6780 32240 6815
rect 32250 6780 32285 6815
rect 32295 6780 32330 6815
rect 32340 6780 32375 6815
rect 32385 6780 32420 6815
rect 32430 6780 32465 6815
rect 32475 6780 32510 6815
rect 32520 6780 32555 6815
rect 32565 6780 32600 6815
rect 32610 6780 32645 6815
rect 32655 6780 32690 6815
rect 32700 6780 32735 6815
rect 32745 6780 32780 6815
rect 32790 6780 32825 6815
rect 32835 6780 32870 6815
rect 31305 6735 31340 6770
rect 31350 6735 31385 6770
rect 31395 6735 31430 6770
rect 31440 6735 31475 6770
rect 31485 6735 31520 6770
rect 31530 6735 31565 6770
rect 31575 6735 31610 6770
rect 31620 6735 31655 6770
rect 31665 6735 31700 6770
rect 31710 6735 31745 6770
rect 31755 6735 31790 6770
rect 31800 6735 31835 6770
rect 31845 6735 31880 6770
rect 31890 6735 31925 6770
rect 31935 6735 31970 6770
rect 31980 6735 32015 6770
rect 32025 6735 32060 6770
rect 32070 6735 32105 6770
rect 32115 6735 32150 6770
rect 32160 6735 32195 6770
rect 32205 6735 32240 6770
rect 32250 6735 32285 6770
rect 32295 6735 32330 6770
rect 32340 6735 32375 6770
rect 32385 6735 32420 6770
rect 32430 6735 32465 6770
rect 32475 6735 32510 6770
rect 32520 6735 32555 6770
rect 32565 6735 32600 6770
rect 32610 6735 32645 6770
rect 32655 6735 32690 6770
rect 32700 6735 32735 6770
rect 32745 6735 32780 6770
rect 32790 6735 32825 6770
rect 32835 6735 32870 6770
rect 31305 6690 31340 6725
rect 31350 6690 31385 6725
rect 31395 6690 31430 6725
rect 31440 6690 31475 6725
rect 31485 6690 31520 6725
rect 31530 6690 31565 6725
rect 31575 6690 31610 6725
rect 31620 6690 31655 6725
rect 31665 6690 31700 6725
rect 31710 6690 31745 6725
rect 31755 6690 31790 6725
rect 31800 6690 31835 6725
rect 31845 6690 31880 6725
rect 31890 6690 31925 6725
rect 31935 6690 31970 6725
rect 31980 6690 32015 6725
rect 32025 6690 32060 6725
rect 32070 6690 32105 6725
rect 32115 6690 32150 6725
rect 32160 6690 32195 6725
rect 32205 6690 32240 6725
rect 32250 6690 32285 6725
rect 32295 6690 32330 6725
rect 32340 6690 32375 6725
rect 32385 6690 32420 6725
rect 32430 6690 32465 6725
rect 32475 6690 32510 6725
rect 32520 6690 32555 6725
rect 32565 6690 32600 6725
rect 32610 6690 32645 6725
rect 32655 6690 32690 6725
rect 32700 6690 32735 6725
rect 32745 6690 32780 6725
rect 32790 6690 32825 6725
rect 32835 6690 32870 6725
rect 31305 6645 31340 6680
rect 31350 6645 31385 6680
rect 31395 6645 31430 6680
rect 31440 6645 31475 6680
rect 31485 6645 31520 6680
rect 31530 6645 31565 6680
rect 31575 6645 31610 6680
rect 31620 6645 31655 6680
rect 31665 6645 31700 6680
rect 31710 6645 31745 6680
rect 31755 6645 31790 6680
rect 31800 6645 31835 6680
rect 31845 6645 31880 6680
rect 31890 6645 31925 6680
rect 31935 6645 31970 6680
rect 31980 6645 32015 6680
rect 32025 6645 32060 6680
rect 32070 6645 32105 6680
rect 32115 6645 32150 6680
rect 32160 6645 32195 6680
rect 32205 6645 32240 6680
rect 32250 6645 32285 6680
rect 32295 6645 32330 6680
rect 32340 6645 32375 6680
rect 32385 6645 32420 6680
rect 32430 6645 32465 6680
rect 32475 6645 32510 6680
rect 32520 6645 32555 6680
rect 32565 6645 32600 6680
rect 32610 6645 32645 6680
rect 32655 6645 32690 6680
rect 32700 6645 32735 6680
rect 32745 6645 32780 6680
rect 32790 6645 32825 6680
rect 32835 6645 32870 6680
rect 31305 6600 31340 6635
rect 31350 6600 31385 6635
rect 31395 6600 31430 6635
rect 31440 6600 31475 6635
rect 31485 6600 31520 6635
rect 31530 6600 31565 6635
rect 31575 6600 31610 6635
rect 31620 6600 31655 6635
rect 31665 6600 31700 6635
rect 31710 6600 31745 6635
rect 31755 6600 31790 6635
rect 31800 6600 31835 6635
rect 31845 6600 31880 6635
rect 31890 6600 31925 6635
rect 31935 6600 31970 6635
rect 31980 6600 32015 6635
rect 32025 6600 32060 6635
rect 32070 6600 32105 6635
rect 32115 6600 32150 6635
rect 32160 6600 32195 6635
rect 32205 6600 32240 6635
rect 32250 6600 32285 6635
rect 32295 6600 32330 6635
rect 32340 6600 32375 6635
rect 32385 6600 32420 6635
rect 32430 6600 32465 6635
rect 32475 6600 32510 6635
rect 32520 6600 32555 6635
rect 32565 6600 32600 6635
rect 32610 6600 32645 6635
rect 32655 6600 32690 6635
rect 32700 6600 32735 6635
rect 32745 6600 32780 6635
rect 32790 6600 32825 6635
rect 32835 6600 32870 6635
rect 31305 6555 31340 6590
rect 31350 6555 31385 6590
rect 31395 6555 31430 6590
rect 31440 6555 31475 6590
rect 31485 6555 31520 6590
rect 31530 6555 31565 6590
rect 31575 6555 31610 6590
rect 31620 6555 31655 6590
rect 31665 6555 31700 6590
rect 31710 6555 31745 6590
rect 31755 6555 31790 6590
rect 31800 6555 31835 6590
rect 31845 6555 31880 6590
rect 31890 6555 31925 6590
rect 31935 6555 31970 6590
rect 31980 6555 32015 6590
rect 32025 6555 32060 6590
rect 32070 6555 32105 6590
rect 32115 6555 32150 6590
rect 32160 6555 32195 6590
rect 32205 6555 32240 6590
rect 32250 6555 32285 6590
rect 32295 6555 32330 6590
rect 32340 6555 32375 6590
rect 32385 6555 32420 6590
rect 32430 6555 32465 6590
rect 32475 6555 32510 6590
rect 32520 6555 32555 6590
rect 32565 6555 32600 6590
rect 32610 6555 32645 6590
rect 32655 6555 32690 6590
rect 32700 6555 32735 6590
rect 32745 6555 32780 6590
rect 32790 6555 32825 6590
rect 32835 6555 32870 6590
rect 31305 6510 31340 6545
rect 31350 6510 31385 6545
rect 31395 6510 31430 6545
rect 31440 6510 31475 6545
rect 31485 6510 31520 6545
rect 31530 6510 31565 6545
rect 31575 6510 31610 6545
rect 31620 6510 31655 6545
rect 31665 6510 31700 6545
rect 31710 6510 31745 6545
rect 31755 6510 31790 6545
rect 31800 6510 31835 6545
rect 31845 6510 31880 6545
rect 31890 6510 31925 6545
rect 31935 6510 31970 6545
rect 31980 6510 32015 6545
rect 32025 6510 32060 6545
rect 32070 6510 32105 6545
rect 32115 6510 32150 6545
rect 32160 6510 32195 6545
rect 32205 6510 32240 6545
rect 32250 6510 32285 6545
rect 32295 6510 32330 6545
rect 32340 6510 32375 6545
rect 32385 6510 32420 6545
rect 32430 6510 32465 6545
rect 32475 6510 32510 6545
rect 32520 6510 32555 6545
rect 32565 6510 32600 6545
rect 32610 6510 32645 6545
rect 32655 6510 32690 6545
rect 32700 6510 32735 6545
rect 32745 6510 32780 6545
rect 32790 6510 32825 6545
rect 32835 6510 32870 6545
rect 31305 6465 31340 6500
rect 31350 6465 31385 6500
rect 31395 6465 31430 6500
rect 31440 6465 31475 6500
rect 31485 6465 31520 6500
rect 31530 6465 31565 6500
rect 31575 6465 31610 6500
rect 31620 6465 31655 6500
rect 31665 6465 31700 6500
rect 31710 6465 31745 6500
rect 31755 6465 31790 6500
rect 31800 6465 31835 6500
rect 31845 6465 31880 6500
rect 31890 6465 31925 6500
rect 31935 6465 31970 6500
rect 31980 6465 32015 6500
rect 32025 6465 32060 6500
rect 32070 6465 32105 6500
rect 32115 6465 32150 6500
rect 32160 6465 32195 6500
rect 32205 6465 32240 6500
rect 32250 6465 32285 6500
rect 32295 6465 32330 6500
rect 32340 6465 32375 6500
rect 32385 6465 32420 6500
rect 32430 6465 32465 6500
rect 32475 6465 32510 6500
rect 32520 6465 32555 6500
rect 32565 6465 32600 6500
rect 32610 6465 32645 6500
rect 32655 6465 32690 6500
rect 32700 6465 32735 6500
rect 32745 6465 32780 6500
rect 32790 6465 32825 6500
rect 32835 6465 32870 6500
rect -80 -1305 -40 -1300
rect -80 -1335 -75 -1305
rect -75 -1335 -45 -1305
rect -45 -1335 -40 -1305
rect -80 -1340 -40 -1335
rect -80 -1370 -40 -1365
rect -80 -1400 -75 -1370
rect -75 -1400 -45 -1370
rect -45 -1400 -40 -1370
rect -80 -1405 -40 -1400
rect -80 -1440 -40 -1435
rect -80 -1470 -75 -1440
rect -75 -1470 -45 -1440
rect -45 -1470 -40 -1440
rect -80 -1475 -40 -1470
rect -80 -1510 -40 -1505
rect -80 -1540 -75 -1510
rect -75 -1540 -45 -1510
rect -45 -1540 -40 -1510
rect -80 -1545 -40 -1540
rect -80 -1580 -40 -1575
rect -80 -1610 -75 -1580
rect -75 -1610 -45 -1580
rect -45 -1610 -40 -1580
rect -80 -1615 -40 -1610
rect -80 -1645 -40 -1640
rect -80 -1675 -75 -1645
rect -75 -1675 -45 -1645
rect -45 -1675 -40 -1645
rect -80 -1680 -40 -1675
rect -80 -1705 -40 -1700
rect -80 -1735 -75 -1705
rect -75 -1735 -45 -1705
rect -45 -1735 -40 -1705
rect -80 -1740 -40 -1735
rect -80 -1770 -40 -1765
rect -80 -1800 -75 -1770
rect -75 -1800 -45 -1770
rect -45 -1800 -40 -1770
rect -80 -1805 -40 -1800
rect -80 -1840 -40 -1835
rect -80 -1870 -75 -1840
rect -75 -1870 -45 -1840
rect -45 -1870 -40 -1840
rect -80 -1875 -40 -1870
rect -80 -1910 -40 -1905
rect -80 -1940 -75 -1910
rect -75 -1940 -45 -1910
rect -45 -1940 -40 -1910
rect -80 -1945 -40 -1940
rect -80 -1980 -40 -1975
rect -80 -2010 -75 -1980
rect -75 -2010 -45 -1980
rect -45 -2010 -40 -1980
rect -80 -2015 -40 -2010
rect -80 -2045 -40 -2040
rect -80 -2075 -75 -2045
rect -75 -2075 -45 -2045
rect -45 -2075 -40 -2045
rect -80 -2080 -40 -2075
rect -80 -2105 -40 -2100
rect -80 -2135 -75 -2105
rect -75 -2135 -45 -2105
rect -45 -2135 -40 -2105
rect -80 -2140 -40 -2135
rect -80 -2170 -40 -2165
rect -80 -2200 -75 -2170
rect -75 -2200 -45 -2170
rect -45 -2200 -40 -2170
rect -80 -2205 -40 -2200
rect -80 -2240 -40 -2235
rect -80 -2270 -75 -2240
rect -75 -2270 -45 -2240
rect -45 -2270 -40 -2240
rect -80 -2275 -40 -2270
rect -80 -2310 -40 -2305
rect -80 -2340 -75 -2310
rect -75 -2340 -45 -2310
rect -45 -2340 -40 -2310
rect -80 -2345 -40 -2340
rect -80 -2380 -40 -2375
rect -80 -2410 -75 -2380
rect -75 -2410 -45 -2380
rect -45 -2410 -40 -2380
rect -80 -2415 -40 -2410
rect -80 -2445 -40 -2440
rect -80 -2475 -75 -2445
rect -75 -2475 -45 -2445
rect -45 -2475 -40 -2445
rect -80 -2480 -40 -2475
rect -80 -2505 -40 -2500
rect -80 -2535 -75 -2505
rect -75 -2535 -45 -2505
rect -45 -2535 -40 -2505
rect -80 -2540 -40 -2535
rect -80 -2570 -40 -2565
rect -80 -2600 -75 -2570
rect -75 -2600 -45 -2570
rect -45 -2600 -40 -2570
rect -80 -2605 -40 -2600
rect -80 -2640 -40 -2635
rect -80 -2670 -75 -2640
rect -75 -2670 -45 -2640
rect -45 -2670 -40 -2640
rect -80 -2675 -40 -2670
rect -80 -2710 -40 -2705
rect -80 -2740 -75 -2710
rect -75 -2740 -45 -2710
rect -45 -2740 -40 -2710
rect -80 -2745 -40 -2740
rect -80 -2780 -40 -2775
rect -80 -2810 -75 -2780
rect -75 -2810 -45 -2780
rect -45 -2810 -40 -2780
rect -80 -2815 -40 -2810
rect -80 -2845 -40 -2840
rect -80 -2875 -75 -2845
rect -75 -2875 -45 -2845
rect -45 -2875 -40 -2845
rect -80 -2880 -40 -2875
rect 270 -1305 310 -1300
rect 270 -1335 275 -1305
rect 275 -1335 305 -1305
rect 305 -1335 310 -1305
rect 270 -1340 310 -1335
rect 270 -1370 310 -1365
rect 270 -1400 275 -1370
rect 275 -1400 305 -1370
rect 305 -1400 310 -1370
rect 270 -1405 310 -1400
rect 270 -1440 310 -1435
rect 270 -1470 275 -1440
rect 275 -1470 305 -1440
rect 305 -1470 310 -1440
rect 270 -1475 310 -1470
rect 270 -1510 310 -1505
rect 270 -1540 275 -1510
rect 275 -1540 305 -1510
rect 305 -1540 310 -1510
rect 270 -1545 310 -1540
rect 270 -1580 310 -1575
rect 270 -1610 275 -1580
rect 275 -1610 305 -1580
rect 305 -1610 310 -1580
rect 270 -1615 310 -1610
rect 270 -1645 310 -1640
rect 270 -1675 275 -1645
rect 275 -1675 305 -1645
rect 305 -1675 310 -1645
rect 270 -1680 310 -1675
rect 270 -1705 310 -1700
rect 270 -1735 275 -1705
rect 275 -1735 305 -1705
rect 305 -1735 310 -1705
rect 270 -1740 310 -1735
rect 270 -1770 310 -1765
rect 270 -1800 275 -1770
rect 275 -1800 305 -1770
rect 305 -1800 310 -1770
rect 270 -1805 310 -1800
rect 270 -1840 310 -1835
rect 270 -1870 275 -1840
rect 275 -1870 305 -1840
rect 305 -1870 310 -1840
rect 270 -1875 310 -1870
rect 270 -1910 310 -1905
rect 270 -1940 275 -1910
rect 275 -1940 305 -1910
rect 305 -1940 310 -1910
rect 270 -1945 310 -1940
rect 270 -1980 310 -1975
rect 270 -2010 275 -1980
rect 275 -2010 305 -1980
rect 305 -2010 310 -1980
rect 270 -2015 310 -2010
rect 270 -2045 310 -2040
rect 270 -2075 275 -2045
rect 275 -2075 305 -2045
rect 305 -2075 310 -2045
rect 270 -2080 310 -2075
rect 270 -2105 310 -2100
rect 270 -2135 275 -2105
rect 275 -2135 305 -2105
rect 305 -2135 310 -2105
rect 270 -2140 310 -2135
rect 270 -2170 310 -2165
rect 270 -2200 275 -2170
rect 275 -2200 305 -2170
rect 305 -2200 310 -2170
rect 270 -2205 310 -2200
rect 270 -2240 310 -2235
rect 270 -2270 275 -2240
rect 275 -2270 305 -2240
rect 305 -2270 310 -2240
rect 270 -2275 310 -2270
rect 270 -2310 310 -2305
rect 270 -2340 275 -2310
rect 275 -2340 305 -2310
rect 305 -2340 310 -2310
rect 270 -2345 310 -2340
rect 270 -2380 310 -2375
rect 270 -2410 275 -2380
rect 275 -2410 305 -2380
rect 305 -2410 310 -2380
rect 270 -2415 310 -2410
rect 270 -2445 310 -2440
rect 270 -2475 275 -2445
rect 275 -2475 305 -2445
rect 305 -2475 310 -2445
rect 270 -2480 310 -2475
rect 270 -2505 310 -2500
rect 270 -2535 275 -2505
rect 275 -2535 305 -2505
rect 305 -2535 310 -2505
rect 270 -2540 310 -2535
rect 270 -2570 310 -2565
rect 270 -2600 275 -2570
rect 275 -2600 305 -2570
rect 305 -2600 310 -2570
rect 270 -2605 310 -2600
rect 270 -2640 310 -2635
rect 270 -2670 275 -2640
rect 275 -2670 305 -2640
rect 305 -2670 310 -2640
rect 270 -2675 310 -2670
rect 270 -2710 310 -2705
rect 270 -2740 275 -2710
rect 275 -2740 305 -2710
rect 305 -2740 310 -2710
rect 270 -2745 310 -2740
rect 270 -2780 310 -2775
rect 270 -2810 275 -2780
rect 275 -2810 305 -2780
rect 305 -2810 310 -2780
rect 270 -2815 310 -2810
rect 270 -2845 310 -2840
rect 270 -2875 275 -2845
rect 275 -2875 305 -2845
rect 305 -2875 310 -2845
rect 270 -2880 310 -2875
rect 620 -1305 660 -1300
rect 620 -1335 625 -1305
rect 625 -1335 655 -1305
rect 655 -1335 660 -1305
rect 620 -1340 660 -1335
rect 620 -1370 660 -1365
rect 620 -1400 625 -1370
rect 625 -1400 655 -1370
rect 655 -1400 660 -1370
rect 620 -1405 660 -1400
rect 620 -1440 660 -1435
rect 620 -1470 625 -1440
rect 625 -1470 655 -1440
rect 655 -1470 660 -1440
rect 620 -1475 660 -1470
rect 620 -1510 660 -1505
rect 620 -1540 625 -1510
rect 625 -1540 655 -1510
rect 655 -1540 660 -1510
rect 620 -1545 660 -1540
rect 620 -1580 660 -1575
rect 620 -1610 625 -1580
rect 625 -1610 655 -1580
rect 655 -1610 660 -1580
rect 620 -1615 660 -1610
rect 620 -1645 660 -1640
rect 620 -1675 625 -1645
rect 625 -1675 655 -1645
rect 655 -1675 660 -1645
rect 620 -1680 660 -1675
rect 620 -1705 660 -1700
rect 620 -1735 625 -1705
rect 625 -1735 655 -1705
rect 655 -1735 660 -1705
rect 620 -1740 660 -1735
rect 620 -1770 660 -1765
rect 620 -1800 625 -1770
rect 625 -1800 655 -1770
rect 655 -1800 660 -1770
rect 620 -1805 660 -1800
rect 620 -1840 660 -1835
rect 620 -1870 625 -1840
rect 625 -1870 655 -1840
rect 655 -1870 660 -1840
rect 620 -1875 660 -1870
rect 620 -1910 660 -1905
rect 620 -1940 625 -1910
rect 625 -1940 655 -1910
rect 655 -1940 660 -1910
rect 620 -1945 660 -1940
rect 620 -1980 660 -1975
rect 620 -2010 625 -1980
rect 625 -2010 655 -1980
rect 655 -2010 660 -1980
rect 620 -2015 660 -2010
rect 620 -2045 660 -2040
rect 620 -2075 625 -2045
rect 625 -2075 655 -2045
rect 655 -2075 660 -2045
rect 620 -2080 660 -2075
rect 620 -2105 660 -2100
rect 620 -2135 625 -2105
rect 625 -2135 655 -2105
rect 655 -2135 660 -2105
rect 620 -2140 660 -2135
rect 620 -2170 660 -2165
rect 620 -2200 625 -2170
rect 625 -2200 655 -2170
rect 655 -2200 660 -2170
rect 620 -2205 660 -2200
rect 620 -2240 660 -2235
rect 620 -2270 625 -2240
rect 625 -2270 655 -2240
rect 655 -2270 660 -2240
rect 620 -2275 660 -2270
rect 620 -2310 660 -2305
rect 620 -2340 625 -2310
rect 625 -2340 655 -2310
rect 655 -2340 660 -2310
rect 620 -2345 660 -2340
rect 620 -2380 660 -2375
rect 620 -2410 625 -2380
rect 625 -2410 655 -2380
rect 655 -2410 660 -2380
rect 620 -2415 660 -2410
rect 620 -2445 660 -2440
rect 620 -2475 625 -2445
rect 625 -2475 655 -2445
rect 655 -2475 660 -2445
rect 620 -2480 660 -2475
rect 620 -2505 660 -2500
rect 620 -2535 625 -2505
rect 625 -2535 655 -2505
rect 655 -2535 660 -2505
rect 620 -2540 660 -2535
rect 620 -2570 660 -2565
rect 620 -2600 625 -2570
rect 625 -2600 655 -2570
rect 655 -2600 660 -2570
rect 620 -2605 660 -2600
rect 620 -2640 660 -2635
rect 620 -2670 625 -2640
rect 625 -2670 655 -2640
rect 655 -2670 660 -2640
rect 620 -2675 660 -2670
rect 620 -2710 660 -2705
rect 620 -2740 625 -2710
rect 625 -2740 655 -2710
rect 655 -2740 660 -2710
rect 620 -2745 660 -2740
rect 620 -2780 660 -2775
rect 620 -2810 625 -2780
rect 625 -2810 655 -2780
rect 655 -2810 660 -2780
rect 620 -2815 660 -2810
rect 620 -2845 660 -2840
rect 620 -2875 625 -2845
rect 625 -2875 655 -2845
rect 655 -2875 660 -2845
rect 620 -2880 660 -2875
rect 970 -1305 1010 -1300
rect 970 -1335 975 -1305
rect 975 -1335 1005 -1305
rect 1005 -1335 1010 -1305
rect 970 -1340 1010 -1335
rect 970 -1370 1010 -1365
rect 970 -1400 975 -1370
rect 975 -1400 1005 -1370
rect 1005 -1400 1010 -1370
rect 970 -1405 1010 -1400
rect 970 -1440 1010 -1435
rect 970 -1470 975 -1440
rect 975 -1470 1005 -1440
rect 1005 -1470 1010 -1440
rect 970 -1475 1010 -1470
rect 970 -1510 1010 -1505
rect 970 -1540 975 -1510
rect 975 -1540 1005 -1510
rect 1005 -1540 1010 -1510
rect 970 -1545 1010 -1540
rect 970 -1580 1010 -1575
rect 970 -1610 975 -1580
rect 975 -1610 1005 -1580
rect 1005 -1610 1010 -1580
rect 970 -1615 1010 -1610
rect 970 -1645 1010 -1640
rect 970 -1675 975 -1645
rect 975 -1675 1005 -1645
rect 1005 -1675 1010 -1645
rect 970 -1680 1010 -1675
rect 970 -1705 1010 -1700
rect 970 -1735 975 -1705
rect 975 -1735 1005 -1705
rect 1005 -1735 1010 -1705
rect 970 -1740 1010 -1735
rect 970 -1770 1010 -1765
rect 970 -1800 975 -1770
rect 975 -1800 1005 -1770
rect 1005 -1800 1010 -1770
rect 970 -1805 1010 -1800
rect 970 -1840 1010 -1835
rect 970 -1870 975 -1840
rect 975 -1870 1005 -1840
rect 1005 -1870 1010 -1840
rect 970 -1875 1010 -1870
rect 970 -1910 1010 -1905
rect 970 -1940 975 -1910
rect 975 -1940 1005 -1910
rect 1005 -1940 1010 -1910
rect 970 -1945 1010 -1940
rect 970 -1980 1010 -1975
rect 970 -2010 975 -1980
rect 975 -2010 1005 -1980
rect 1005 -2010 1010 -1980
rect 970 -2015 1010 -2010
rect 970 -2045 1010 -2040
rect 970 -2075 975 -2045
rect 975 -2075 1005 -2045
rect 1005 -2075 1010 -2045
rect 970 -2080 1010 -2075
rect 970 -2105 1010 -2100
rect 970 -2135 975 -2105
rect 975 -2135 1005 -2105
rect 1005 -2135 1010 -2105
rect 970 -2140 1010 -2135
rect 970 -2170 1010 -2165
rect 970 -2200 975 -2170
rect 975 -2200 1005 -2170
rect 1005 -2200 1010 -2170
rect 970 -2205 1010 -2200
rect 970 -2240 1010 -2235
rect 970 -2270 975 -2240
rect 975 -2270 1005 -2240
rect 1005 -2270 1010 -2240
rect 970 -2275 1010 -2270
rect 970 -2310 1010 -2305
rect 970 -2340 975 -2310
rect 975 -2340 1005 -2310
rect 1005 -2340 1010 -2310
rect 970 -2345 1010 -2340
rect 970 -2380 1010 -2375
rect 970 -2410 975 -2380
rect 975 -2410 1005 -2380
rect 1005 -2410 1010 -2380
rect 970 -2415 1010 -2410
rect 970 -2445 1010 -2440
rect 970 -2475 975 -2445
rect 975 -2475 1005 -2445
rect 1005 -2475 1010 -2445
rect 970 -2480 1010 -2475
rect 970 -2505 1010 -2500
rect 970 -2535 975 -2505
rect 975 -2535 1005 -2505
rect 1005 -2535 1010 -2505
rect 970 -2540 1010 -2535
rect 970 -2570 1010 -2565
rect 970 -2600 975 -2570
rect 975 -2600 1005 -2570
rect 1005 -2600 1010 -2570
rect 970 -2605 1010 -2600
rect 970 -2640 1010 -2635
rect 970 -2670 975 -2640
rect 975 -2670 1005 -2640
rect 1005 -2670 1010 -2640
rect 970 -2675 1010 -2670
rect 970 -2710 1010 -2705
rect 970 -2740 975 -2710
rect 975 -2740 1005 -2710
rect 1005 -2740 1010 -2710
rect 970 -2745 1010 -2740
rect 970 -2780 1010 -2775
rect 970 -2810 975 -2780
rect 975 -2810 1005 -2780
rect 1005 -2810 1010 -2780
rect 970 -2815 1010 -2810
rect 970 -2845 1010 -2840
rect 970 -2875 975 -2845
rect 975 -2875 1005 -2845
rect 1005 -2875 1010 -2845
rect 970 -2880 1010 -2875
rect 1320 -1305 1360 -1300
rect 1320 -1335 1325 -1305
rect 1325 -1335 1355 -1305
rect 1355 -1335 1360 -1305
rect 1320 -1340 1360 -1335
rect 1320 -1370 1360 -1365
rect 1320 -1400 1325 -1370
rect 1325 -1400 1355 -1370
rect 1355 -1400 1360 -1370
rect 1320 -1405 1360 -1400
rect 1320 -1440 1360 -1435
rect 1320 -1470 1325 -1440
rect 1325 -1470 1355 -1440
rect 1355 -1470 1360 -1440
rect 1320 -1475 1360 -1470
rect 1320 -1510 1360 -1505
rect 1320 -1540 1325 -1510
rect 1325 -1540 1355 -1510
rect 1355 -1540 1360 -1510
rect 1320 -1545 1360 -1540
rect 1320 -1580 1360 -1575
rect 1320 -1610 1325 -1580
rect 1325 -1610 1355 -1580
rect 1355 -1610 1360 -1580
rect 1320 -1615 1360 -1610
rect 1320 -1645 1360 -1640
rect 1320 -1675 1325 -1645
rect 1325 -1675 1355 -1645
rect 1355 -1675 1360 -1645
rect 1320 -1680 1360 -1675
rect 1320 -1705 1360 -1700
rect 1320 -1735 1325 -1705
rect 1325 -1735 1355 -1705
rect 1355 -1735 1360 -1705
rect 1320 -1740 1360 -1735
rect 1320 -1770 1360 -1765
rect 1320 -1800 1325 -1770
rect 1325 -1800 1355 -1770
rect 1355 -1800 1360 -1770
rect 1320 -1805 1360 -1800
rect 1320 -1840 1360 -1835
rect 1320 -1870 1325 -1840
rect 1325 -1870 1355 -1840
rect 1355 -1870 1360 -1840
rect 1320 -1875 1360 -1870
rect 1320 -1910 1360 -1905
rect 1320 -1940 1325 -1910
rect 1325 -1940 1355 -1910
rect 1355 -1940 1360 -1910
rect 1320 -1945 1360 -1940
rect 1320 -1980 1360 -1975
rect 1320 -2010 1325 -1980
rect 1325 -2010 1355 -1980
rect 1355 -2010 1360 -1980
rect 1320 -2015 1360 -2010
rect 1320 -2045 1360 -2040
rect 1320 -2075 1325 -2045
rect 1325 -2075 1355 -2045
rect 1355 -2075 1360 -2045
rect 1320 -2080 1360 -2075
rect 1320 -2105 1360 -2100
rect 1320 -2135 1325 -2105
rect 1325 -2135 1355 -2105
rect 1355 -2135 1360 -2105
rect 1320 -2140 1360 -2135
rect 1320 -2170 1360 -2165
rect 1320 -2200 1325 -2170
rect 1325 -2200 1355 -2170
rect 1355 -2200 1360 -2170
rect 1320 -2205 1360 -2200
rect 1320 -2240 1360 -2235
rect 1320 -2270 1325 -2240
rect 1325 -2270 1355 -2240
rect 1355 -2270 1360 -2240
rect 1320 -2275 1360 -2270
rect 1320 -2310 1360 -2305
rect 1320 -2340 1325 -2310
rect 1325 -2340 1355 -2310
rect 1355 -2340 1360 -2310
rect 1320 -2345 1360 -2340
rect 1320 -2380 1360 -2375
rect 1320 -2410 1325 -2380
rect 1325 -2410 1355 -2380
rect 1355 -2410 1360 -2380
rect 1320 -2415 1360 -2410
rect 1320 -2445 1360 -2440
rect 1320 -2475 1325 -2445
rect 1325 -2475 1355 -2445
rect 1355 -2475 1360 -2445
rect 1320 -2480 1360 -2475
rect 1320 -2505 1360 -2500
rect 1320 -2535 1325 -2505
rect 1325 -2535 1355 -2505
rect 1355 -2535 1360 -2505
rect 1320 -2540 1360 -2535
rect 1320 -2570 1360 -2565
rect 1320 -2600 1325 -2570
rect 1325 -2600 1355 -2570
rect 1355 -2600 1360 -2570
rect 1320 -2605 1360 -2600
rect 1320 -2640 1360 -2635
rect 1320 -2670 1325 -2640
rect 1325 -2670 1355 -2640
rect 1355 -2670 1360 -2640
rect 1320 -2675 1360 -2670
rect 1320 -2710 1360 -2705
rect 1320 -2740 1325 -2710
rect 1325 -2740 1355 -2710
rect 1355 -2740 1360 -2710
rect 1320 -2745 1360 -2740
rect 1320 -2780 1360 -2775
rect 1320 -2810 1325 -2780
rect 1325 -2810 1355 -2780
rect 1355 -2810 1360 -2780
rect 1320 -2815 1360 -2810
rect 1320 -2845 1360 -2840
rect 1320 -2875 1325 -2845
rect 1325 -2875 1355 -2845
rect 1355 -2875 1360 -2845
rect 1320 -2880 1360 -2875
rect 1670 -1305 1710 -1300
rect 1670 -1335 1675 -1305
rect 1675 -1335 1705 -1305
rect 1705 -1335 1710 -1305
rect 1670 -1340 1710 -1335
rect 1670 -1370 1710 -1365
rect 1670 -1400 1675 -1370
rect 1675 -1400 1705 -1370
rect 1705 -1400 1710 -1370
rect 1670 -1405 1710 -1400
rect 1670 -1440 1710 -1435
rect 1670 -1470 1675 -1440
rect 1675 -1470 1705 -1440
rect 1705 -1470 1710 -1440
rect 1670 -1475 1710 -1470
rect 1670 -1510 1710 -1505
rect 1670 -1540 1675 -1510
rect 1675 -1540 1705 -1510
rect 1705 -1540 1710 -1510
rect 1670 -1545 1710 -1540
rect 1670 -1580 1710 -1575
rect 1670 -1610 1675 -1580
rect 1675 -1610 1705 -1580
rect 1705 -1610 1710 -1580
rect 1670 -1615 1710 -1610
rect 1670 -1645 1710 -1640
rect 1670 -1675 1675 -1645
rect 1675 -1675 1705 -1645
rect 1705 -1675 1710 -1645
rect 1670 -1680 1710 -1675
rect 1670 -1705 1710 -1700
rect 1670 -1735 1675 -1705
rect 1675 -1735 1705 -1705
rect 1705 -1735 1710 -1705
rect 1670 -1740 1710 -1735
rect 1670 -1770 1710 -1765
rect 1670 -1800 1675 -1770
rect 1675 -1800 1705 -1770
rect 1705 -1800 1710 -1770
rect 1670 -1805 1710 -1800
rect 1670 -1840 1710 -1835
rect 1670 -1870 1675 -1840
rect 1675 -1870 1705 -1840
rect 1705 -1870 1710 -1840
rect 1670 -1875 1710 -1870
rect 1670 -1910 1710 -1905
rect 1670 -1940 1675 -1910
rect 1675 -1940 1705 -1910
rect 1705 -1940 1710 -1910
rect 1670 -1945 1710 -1940
rect 1670 -1980 1710 -1975
rect 1670 -2010 1675 -1980
rect 1675 -2010 1705 -1980
rect 1705 -2010 1710 -1980
rect 1670 -2015 1710 -2010
rect 1670 -2045 1710 -2040
rect 1670 -2075 1675 -2045
rect 1675 -2075 1705 -2045
rect 1705 -2075 1710 -2045
rect 1670 -2080 1710 -2075
rect 1670 -2105 1710 -2100
rect 1670 -2135 1675 -2105
rect 1675 -2135 1705 -2105
rect 1705 -2135 1710 -2105
rect 1670 -2140 1710 -2135
rect 1670 -2170 1710 -2165
rect 1670 -2200 1675 -2170
rect 1675 -2200 1705 -2170
rect 1705 -2200 1710 -2170
rect 1670 -2205 1710 -2200
rect 1670 -2240 1710 -2235
rect 1670 -2270 1675 -2240
rect 1675 -2270 1705 -2240
rect 1705 -2270 1710 -2240
rect 1670 -2275 1710 -2270
rect 1670 -2310 1710 -2305
rect 1670 -2340 1675 -2310
rect 1675 -2340 1705 -2310
rect 1705 -2340 1710 -2310
rect 1670 -2345 1710 -2340
rect 1670 -2380 1710 -2375
rect 1670 -2410 1675 -2380
rect 1675 -2410 1705 -2380
rect 1705 -2410 1710 -2380
rect 1670 -2415 1710 -2410
rect 1670 -2445 1710 -2440
rect 1670 -2475 1675 -2445
rect 1675 -2475 1705 -2445
rect 1705 -2475 1710 -2445
rect 1670 -2480 1710 -2475
rect 1670 -2505 1710 -2500
rect 1670 -2535 1675 -2505
rect 1675 -2535 1705 -2505
rect 1705 -2535 1710 -2505
rect 1670 -2540 1710 -2535
rect 1670 -2570 1710 -2565
rect 1670 -2600 1675 -2570
rect 1675 -2600 1705 -2570
rect 1705 -2600 1710 -2570
rect 1670 -2605 1710 -2600
rect 1670 -2640 1710 -2635
rect 1670 -2670 1675 -2640
rect 1675 -2670 1705 -2640
rect 1705 -2670 1710 -2640
rect 1670 -2675 1710 -2670
rect 1670 -2710 1710 -2705
rect 1670 -2740 1675 -2710
rect 1675 -2740 1705 -2710
rect 1705 -2740 1710 -2710
rect 1670 -2745 1710 -2740
rect 1670 -2780 1710 -2775
rect 1670 -2810 1675 -2780
rect 1675 -2810 1705 -2780
rect 1705 -2810 1710 -2780
rect 1670 -2815 1710 -2810
rect 1670 -2845 1710 -2840
rect 1670 -2875 1675 -2845
rect 1675 -2875 1705 -2845
rect 1705 -2875 1710 -2845
rect 1670 -2880 1710 -2875
rect 2020 -1305 2060 -1300
rect 2020 -1335 2025 -1305
rect 2025 -1335 2055 -1305
rect 2055 -1335 2060 -1305
rect 2020 -1340 2060 -1335
rect 2020 -1370 2060 -1365
rect 2020 -1400 2025 -1370
rect 2025 -1400 2055 -1370
rect 2055 -1400 2060 -1370
rect 2020 -1405 2060 -1400
rect 2020 -1440 2060 -1435
rect 2020 -1470 2025 -1440
rect 2025 -1470 2055 -1440
rect 2055 -1470 2060 -1440
rect 2020 -1475 2060 -1470
rect 2020 -1510 2060 -1505
rect 2020 -1540 2025 -1510
rect 2025 -1540 2055 -1510
rect 2055 -1540 2060 -1510
rect 2020 -1545 2060 -1540
rect 2020 -1580 2060 -1575
rect 2020 -1610 2025 -1580
rect 2025 -1610 2055 -1580
rect 2055 -1610 2060 -1580
rect 2020 -1615 2060 -1610
rect 2020 -1645 2060 -1640
rect 2020 -1675 2025 -1645
rect 2025 -1675 2055 -1645
rect 2055 -1675 2060 -1645
rect 2020 -1680 2060 -1675
rect 2020 -1705 2060 -1700
rect 2020 -1735 2025 -1705
rect 2025 -1735 2055 -1705
rect 2055 -1735 2060 -1705
rect 2020 -1740 2060 -1735
rect 2020 -1770 2060 -1765
rect 2020 -1800 2025 -1770
rect 2025 -1800 2055 -1770
rect 2055 -1800 2060 -1770
rect 2020 -1805 2060 -1800
rect 2020 -1840 2060 -1835
rect 2020 -1870 2025 -1840
rect 2025 -1870 2055 -1840
rect 2055 -1870 2060 -1840
rect 2020 -1875 2060 -1870
rect 2020 -1910 2060 -1905
rect 2020 -1940 2025 -1910
rect 2025 -1940 2055 -1910
rect 2055 -1940 2060 -1910
rect 2020 -1945 2060 -1940
rect 2020 -1980 2060 -1975
rect 2020 -2010 2025 -1980
rect 2025 -2010 2055 -1980
rect 2055 -2010 2060 -1980
rect 2020 -2015 2060 -2010
rect 2020 -2045 2060 -2040
rect 2020 -2075 2025 -2045
rect 2025 -2075 2055 -2045
rect 2055 -2075 2060 -2045
rect 2020 -2080 2060 -2075
rect 2020 -2105 2060 -2100
rect 2020 -2135 2025 -2105
rect 2025 -2135 2055 -2105
rect 2055 -2135 2060 -2105
rect 2020 -2140 2060 -2135
rect 2020 -2170 2060 -2165
rect 2020 -2200 2025 -2170
rect 2025 -2200 2055 -2170
rect 2055 -2200 2060 -2170
rect 2020 -2205 2060 -2200
rect 2020 -2240 2060 -2235
rect 2020 -2270 2025 -2240
rect 2025 -2270 2055 -2240
rect 2055 -2270 2060 -2240
rect 2020 -2275 2060 -2270
rect 2020 -2310 2060 -2305
rect 2020 -2340 2025 -2310
rect 2025 -2340 2055 -2310
rect 2055 -2340 2060 -2310
rect 2020 -2345 2060 -2340
rect 2020 -2380 2060 -2375
rect 2020 -2410 2025 -2380
rect 2025 -2410 2055 -2380
rect 2055 -2410 2060 -2380
rect 2020 -2415 2060 -2410
rect 2020 -2445 2060 -2440
rect 2020 -2475 2025 -2445
rect 2025 -2475 2055 -2445
rect 2055 -2475 2060 -2445
rect 2020 -2480 2060 -2475
rect 2020 -2505 2060 -2500
rect 2020 -2535 2025 -2505
rect 2025 -2535 2055 -2505
rect 2055 -2535 2060 -2505
rect 2020 -2540 2060 -2535
rect 2020 -2570 2060 -2565
rect 2020 -2600 2025 -2570
rect 2025 -2600 2055 -2570
rect 2055 -2600 2060 -2570
rect 2020 -2605 2060 -2600
rect 2020 -2640 2060 -2635
rect 2020 -2670 2025 -2640
rect 2025 -2670 2055 -2640
rect 2055 -2670 2060 -2640
rect 2020 -2675 2060 -2670
rect 2020 -2710 2060 -2705
rect 2020 -2740 2025 -2710
rect 2025 -2740 2055 -2710
rect 2055 -2740 2060 -2710
rect 2020 -2745 2060 -2740
rect 2020 -2780 2060 -2775
rect 2020 -2810 2025 -2780
rect 2025 -2810 2055 -2780
rect 2055 -2810 2060 -2780
rect 2020 -2815 2060 -2810
rect 2020 -2845 2060 -2840
rect 2020 -2875 2025 -2845
rect 2025 -2875 2055 -2845
rect 2055 -2875 2060 -2845
rect 2020 -2880 2060 -2875
rect 2370 -1305 2410 -1300
rect 2370 -1335 2375 -1305
rect 2375 -1335 2405 -1305
rect 2405 -1335 2410 -1305
rect 2370 -1340 2410 -1335
rect 2370 -1370 2410 -1365
rect 2370 -1400 2375 -1370
rect 2375 -1400 2405 -1370
rect 2405 -1400 2410 -1370
rect 2370 -1405 2410 -1400
rect 2370 -1440 2410 -1435
rect 2370 -1470 2375 -1440
rect 2375 -1470 2405 -1440
rect 2405 -1470 2410 -1440
rect 2370 -1475 2410 -1470
rect 2370 -1510 2410 -1505
rect 2370 -1540 2375 -1510
rect 2375 -1540 2405 -1510
rect 2405 -1540 2410 -1510
rect 2370 -1545 2410 -1540
rect 2370 -1580 2410 -1575
rect 2370 -1610 2375 -1580
rect 2375 -1610 2405 -1580
rect 2405 -1610 2410 -1580
rect 2370 -1615 2410 -1610
rect 2370 -1645 2410 -1640
rect 2370 -1675 2375 -1645
rect 2375 -1675 2405 -1645
rect 2405 -1675 2410 -1645
rect 2370 -1680 2410 -1675
rect 2370 -1705 2410 -1700
rect 2370 -1735 2375 -1705
rect 2375 -1735 2405 -1705
rect 2405 -1735 2410 -1705
rect 2370 -1740 2410 -1735
rect 2370 -1770 2410 -1765
rect 2370 -1800 2375 -1770
rect 2375 -1800 2405 -1770
rect 2405 -1800 2410 -1770
rect 2370 -1805 2410 -1800
rect 2370 -1840 2410 -1835
rect 2370 -1870 2375 -1840
rect 2375 -1870 2405 -1840
rect 2405 -1870 2410 -1840
rect 2370 -1875 2410 -1870
rect 2370 -1910 2410 -1905
rect 2370 -1940 2375 -1910
rect 2375 -1940 2405 -1910
rect 2405 -1940 2410 -1910
rect 2370 -1945 2410 -1940
rect 2370 -1980 2410 -1975
rect 2370 -2010 2375 -1980
rect 2375 -2010 2405 -1980
rect 2405 -2010 2410 -1980
rect 2370 -2015 2410 -2010
rect 2370 -2045 2410 -2040
rect 2370 -2075 2375 -2045
rect 2375 -2075 2405 -2045
rect 2405 -2075 2410 -2045
rect 2370 -2080 2410 -2075
rect 2370 -2105 2410 -2100
rect 2370 -2135 2375 -2105
rect 2375 -2135 2405 -2105
rect 2405 -2135 2410 -2105
rect 2370 -2140 2410 -2135
rect 2370 -2170 2410 -2165
rect 2370 -2200 2375 -2170
rect 2375 -2200 2405 -2170
rect 2405 -2200 2410 -2170
rect 2370 -2205 2410 -2200
rect 2370 -2240 2410 -2235
rect 2370 -2270 2375 -2240
rect 2375 -2270 2405 -2240
rect 2405 -2270 2410 -2240
rect 2370 -2275 2410 -2270
rect 2370 -2310 2410 -2305
rect 2370 -2340 2375 -2310
rect 2375 -2340 2405 -2310
rect 2405 -2340 2410 -2310
rect 2370 -2345 2410 -2340
rect 2370 -2380 2410 -2375
rect 2370 -2410 2375 -2380
rect 2375 -2410 2405 -2380
rect 2405 -2410 2410 -2380
rect 2370 -2415 2410 -2410
rect 2370 -2445 2410 -2440
rect 2370 -2475 2375 -2445
rect 2375 -2475 2405 -2445
rect 2405 -2475 2410 -2445
rect 2370 -2480 2410 -2475
rect 2370 -2505 2410 -2500
rect 2370 -2535 2375 -2505
rect 2375 -2535 2405 -2505
rect 2405 -2535 2410 -2505
rect 2370 -2540 2410 -2535
rect 2370 -2570 2410 -2565
rect 2370 -2600 2375 -2570
rect 2375 -2600 2405 -2570
rect 2405 -2600 2410 -2570
rect 2370 -2605 2410 -2600
rect 2370 -2640 2410 -2635
rect 2370 -2670 2375 -2640
rect 2375 -2670 2405 -2640
rect 2405 -2670 2410 -2640
rect 2370 -2675 2410 -2670
rect 2370 -2710 2410 -2705
rect 2370 -2740 2375 -2710
rect 2375 -2740 2405 -2710
rect 2405 -2740 2410 -2710
rect 2370 -2745 2410 -2740
rect 2370 -2780 2410 -2775
rect 2370 -2810 2375 -2780
rect 2375 -2810 2405 -2780
rect 2405 -2810 2410 -2780
rect 2370 -2815 2410 -2810
rect 2370 -2845 2410 -2840
rect 2370 -2875 2375 -2845
rect 2375 -2875 2405 -2845
rect 2405 -2875 2410 -2845
rect 2370 -2880 2410 -2875
rect 2720 -1305 2760 -1300
rect 2720 -1335 2725 -1305
rect 2725 -1335 2755 -1305
rect 2755 -1335 2760 -1305
rect 2720 -1340 2760 -1335
rect 2720 -1370 2760 -1365
rect 2720 -1400 2725 -1370
rect 2725 -1400 2755 -1370
rect 2755 -1400 2760 -1370
rect 2720 -1405 2760 -1400
rect 2720 -1440 2760 -1435
rect 2720 -1470 2725 -1440
rect 2725 -1470 2755 -1440
rect 2755 -1470 2760 -1440
rect 2720 -1475 2760 -1470
rect 2720 -1510 2760 -1505
rect 2720 -1540 2725 -1510
rect 2725 -1540 2755 -1510
rect 2755 -1540 2760 -1510
rect 2720 -1545 2760 -1540
rect 2720 -1580 2760 -1575
rect 2720 -1610 2725 -1580
rect 2725 -1610 2755 -1580
rect 2755 -1610 2760 -1580
rect 2720 -1615 2760 -1610
rect 2720 -1645 2760 -1640
rect 2720 -1675 2725 -1645
rect 2725 -1675 2755 -1645
rect 2755 -1675 2760 -1645
rect 2720 -1680 2760 -1675
rect 2720 -1705 2760 -1700
rect 2720 -1735 2725 -1705
rect 2725 -1735 2755 -1705
rect 2755 -1735 2760 -1705
rect 2720 -1740 2760 -1735
rect 2720 -1770 2760 -1765
rect 2720 -1800 2725 -1770
rect 2725 -1800 2755 -1770
rect 2755 -1800 2760 -1770
rect 2720 -1805 2760 -1800
rect 2720 -1840 2760 -1835
rect 2720 -1870 2725 -1840
rect 2725 -1870 2755 -1840
rect 2755 -1870 2760 -1840
rect 2720 -1875 2760 -1870
rect 2720 -1910 2760 -1905
rect 2720 -1940 2725 -1910
rect 2725 -1940 2755 -1910
rect 2755 -1940 2760 -1910
rect 2720 -1945 2760 -1940
rect 2720 -1980 2760 -1975
rect 2720 -2010 2725 -1980
rect 2725 -2010 2755 -1980
rect 2755 -2010 2760 -1980
rect 2720 -2015 2760 -2010
rect 2720 -2045 2760 -2040
rect 2720 -2075 2725 -2045
rect 2725 -2075 2755 -2045
rect 2755 -2075 2760 -2045
rect 2720 -2080 2760 -2075
rect 2720 -2105 2760 -2100
rect 2720 -2135 2725 -2105
rect 2725 -2135 2755 -2105
rect 2755 -2135 2760 -2105
rect 2720 -2140 2760 -2135
rect 2720 -2170 2760 -2165
rect 2720 -2200 2725 -2170
rect 2725 -2200 2755 -2170
rect 2755 -2200 2760 -2170
rect 2720 -2205 2760 -2200
rect 2720 -2240 2760 -2235
rect 2720 -2270 2725 -2240
rect 2725 -2270 2755 -2240
rect 2755 -2270 2760 -2240
rect 2720 -2275 2760 -2270
rect 2720 -2310 2760 -2305
rect 2720 -2340 2725 -2310
rect 2725 -2340 2755 -2310
rect 2755 -2340 2760 -2310
rect 2720 -2345 2760 -2340
rect 2720 -2380 2760 -2375
rect 2720 -2410 2725 -2380
rect 2725 -2410 2755 -2380
rect 2755 -2410 2760 -2380
rect 2720 -2415 2760 -2410
rect 2720 -2445 2760 -2440
rect 2720 -2475 2725 -2445
rect 2725 -2475 2755 -2445
rect 2755 -2475 2760 -2445
rect 2720 -2480 2760 -2475
rect 2720 -2505 2760 -2500
rect 2720 -2535 2725 -2505
rect 2725 -2535 2755 -2505
rect 2755 -2535 2760 -2505
rect 2720 -2540 2760 -2535
rect 2720 -2570 2760 -2565
rect 2720 -2600 2725 -2570
rect 2725 -2600 2755 -2570
rect 2755 -2600 2760 -2570
rect 2720 -2605 2760 -2600
rect 2720 -2640 2760 -2635
rect 2720 -2670 2725 -2640
rect 2725 -2670 2755 -2640
rect 2755 -2670 2760 -2640
rect 2720 -2675 2760 -2670
rect 2720 -2710 2760 -2705
rect 2720 -2740 2725 -2710
rect 2725 -2740 2755 -2710
rect 2755 -2740 2760 -2710
rect 2720 -2745 2760 -2740
rect 2720 -2780 2760 -2775
rect 2720 -2810 2725 -2780
rect 2725 -2810 2755 -2780
rect 2755 -2810 2760 -2780
rect 2720 -2815 2760 -2810
rect 2720 -2845 2760 -2840
rect 2720 -2875 2725 -2845
rect 2725 -2875 2755 -2845
rect 2755 -2875 2760 -2845
rect 2720 -2880 2760 -2875
rect 3070 -1305 3110 -1300
rect 3070 -1335 3075 -1305
rect 3075 -1335 3105 -1305
rect 3105 -1335 3110 -1305
rect 3070 -1340 3110 -1335
rect 3070 -1370 3110 -1365
rect 3070 -1400 3075 -1370
rect 3075 -1400 3105 -1370
rect 3105 -1400 3110 -1370
rect 3070 -1405 3110 -1400
rect 3070 -1440 3110 -1435
rect 3070 -1470 3075 -1440
rect 3075 -1470 3105 -1440
rect 3105 -1470 3110 -1440
rect 3070 -1475 3110 -1470
rect 3070 -1510 3110 -1505
rect 3070 -1540 3075 -1510
rect 3075 -1540 3105 -1510
rect 3105 -1540 3110 -1510
rect 3070 -1545 3110 -1540
rect 3070 -1580 3110 -1575
rect 3070 -1610 3075 -1580
rect 3075 -1610 3105 -1580
rect 3105 -1610 3110 -1580
rect 3070 -1615 3110 -1610
rect 3070 -1645 3110 -1640
rect 3070 -1675 3075 -1645
rect 3075 -1675 3105 -1645
rect 3105 -1675 3110 -1645
rect 3070 -1680 3110 -1675
rect 3070 -1705 3110 -1700
rect 3070 -1735 3075 -1705
rect 3075 -1735 3105 -1705
rect 3105 -1735 3110 -1705
rect 3070 -1740 3110 -1735
rect 3070 -1770 3110 -1765
rect 3070 -1800 3075 -1770
rect 3075 -1800 3105 -1770
rect 3105 -1800 3110 -1770
rect 3070 -1805 3110 -1800
rect 3070 -1840 3110 -1835
rect 3070 -1870 3075 -1840
rect 3075 -1870 3105 -1840
rect 3105 -1870 3110 -1840
rect 3070 -1875 3110 -1870
rect 3070 -1910 3110 -1905
rect 3070 -1940 3075 -1910
rect 3075 -1940 3105 -1910
rect 3105 -1940 3110 -1910
rect 3070 -1945 3110 -1940
rect 3070 -1980 3110 -1975
rect 3070 -2010 3075 -1980
rect 3075 -2010 3105 -1980
rect 3105 -2010 3110 -1980
rect 3070 -2015 3110 -2010
rect 3070 -2045 3110 -2040
rect 3070 -2075 3075 -2045
rect 3075 -2075 3105 -2045
rect 3105 -2075 3110 -2045
rect 3070 -2080 3110 -2075
rect 3070 -2105 3110 -2100
rect 3070 -2135 3075 -2105
rect 3075 -2135 3105 -2105
rect 3105 -2135 3110 -2105
rect 3070 -2140 3110 -2135
rect 3070 -2170 3110 -2165
rect 3070 -2200 3075 -2170
rect 3075 -2200 3105 -2170
rect 3105 -2200 3110 -2170
rect 3070 -2205 3110 -2200
rect 3070 -2240 3110 -2235
rect 3070 -2270 3075 -2240
rect 3075 -2270 3105 -2240
rect 3105 -2270 3110 -2240
rect 3070 -2275 3110 -2270
rect 3070 -2310 3110 -2305
rect 3070 -2340 3075 -2310
rect 3075 -2340 3105 -2310
rect 3105 -2340 3110 -2310
rect 3070 -2345 3110 -2340
rect 3070 -2380 3110 -2375
rect 3070 -2410 3075 -2380
rect 3075 -2410 3105 -2380
rect 3105 -2410 3110 -2380
rect 3070 -2415 3110 -2410
rect 3070 -2445 3110 -2440
rect 3070 -2475 3075 -2445
rect 3075 -2475 3105 -2445
rect 3105 -2475 3110 -2445
rect 3070 -2480 3110 -2475
rect 3070 -2505 3110 -2500
rect 3070 -2535 3075 -2505
rect 3075 -2535 3105 -2505
rect 3105 -2535 3110 -2505
rect 3070 -2540 3110 -2535
rect 3070 -2570 3110 -2565
rect 3070 -2600 3075 -2570
rect 3075 -2600 3105 -2570
rect 3105 -2600 3110 -2570
rect 3070 -2605 3110 -2600
rect 3070 -2640 3110 -2635
rect 3070 -2670 3075 -2640
rect 3075 -2670 3105 -2640
rect 3105 -2670 3110 -2640
rect 3070 -2675 3110 -2670
rect 3070 -2710 3110 -2705
rect 3070 -2740 3075 -2710
rect 3075 -2740 3105 -2710
rect 3105 -2740 3110 -2710
rect 3070 -2745 3110 -2740
rect 3070 -2780 3110 -2775
rect 3070 -2810 3075 -2780
rect 3075 -2810 3105 -2780
rect 3105 -2810 3110 -2780
rect 3070 -2815 3110 -2810
rect 3070 -2845 3110 -2840
rect 3070 -2875 3075 -2845
rect 3075 -2875 3105 -2845
rect 3105 -2875 3110 -2845
rect 3070 -2880 3110 -2875
rect 3420 -1305 3460 -1300
rect 3420 -1335 3425 -1305
rect 3425 -1335 3455 -1305
rect 3455 -1335 3460 -1305
rect 3420 -1340 3460 -1335
rect 3420 -1370 3460 -1365
rect 3420 -1400 3425 -1370
rect 3425 -1400 3455 -1370
rect 3455 -1400 3460 -1370
rect 3420 -1405 3460 -1400
rect 3420 -1440 3460 -1435
rect 3420 -1470 3425 -1440
rect 3425 -1470 3455 -1440
rect 3455 -1470 3460 -1440
rect 3420 -1475 3460 -1470
rect 3420 -1510 3460 -1505
rect 3420 -1540 3425 -1510
rect 3425 -1540 3455 -1510
rect 3455 -1540 3460 -1510
rect 3420 -1545 3460 -1540
rect 3420 -1580 3460 -1575
rect 3420 -1610 3425 -1580
rect 3425 -1610 3455 -1580
rect 3455 -1610 3460 -1580
rect 3420 -1615 3460 -1610
rect 3420 -1645 3460 -1640
rect 3420 -1675 3425 -1645
rect 3425 -1675 3455 -1645
rect 3455 -1675 3460 -1645
rect 3420 -1680 3460 -1675
rect 3420 -1705 3460 -1700
rect 3420 -1735 3425 -1705
rect 3425 -1735 3455 -1705
rect 3455 -1735 3460 -1705
rect 3420 -1740 3460 -1735
rect 3420 -1770 3460 -1765
rect 3420 -1800 3425 -1770
rect 3425 -1800 3455 -1770
rect 3455 -1800 3460 -1770
rect 3420 -1805 3460 -1800
rect 3420 -1840 3460 -1835
rect 3420 -1870 3425 -1840
rect 3425 -1870 3455 -1840
rect 3455 -1870 3460 -1840
rect 3420 -1875 3460 -1870
rect 3420 -1910 3460 -1905
rect 3420 -1940 3425 -1910
rect 3425 -1940 3455 -1910
rect 3455 -1940 3460 -1910
rect 3420 -1945 3460 -1940
rect 3420 -1980 3460 -1975
rect 3420 -2010 3425 -1980
rect 3425 -2010 3455 -1980
rect 3455 -2010 3460 -1980
rect 3420 -2015 3460 -2010
rect 3420 -2045 3460 -2040
rect 3420 -2075 3425 -2045
rect 3425 -2075 3455 -2045
rect 3455 -2075 3460 -2045
rect 3420 -2080 3460 -2075
rect 3420 -2105 3460 -2100
rect 3420 -2135 3425 -2105
rect 3425 -2135 3455 -2105
rect 3455 -2135 3460 -2105
rect 3420 -2140 3460 -2135
rect 3420 -2170 3460 -2165
rect 3420 -2200 3425 -2170
rect 3425 -2200 3455 -2170
rect 3455 -2200 3460 -2170
rect 3420 -2205 3460 -2200
rect 3420 -2240 3460 -2235
rect 3420 -2270 3425 -2240
rect 3425 -2270 3455 -2240
rect 3455 -2270 3460 -2240
rect 3420 -2275 3460 -2270
rect 3420 -2310 3460 -2305
rect 3420 -2340 3425 -2310
rect 3425 -2340 3455 -2310
rect 3455 -2340 3460 -2310
rect 3420 -2345 3460 -2340
rect 3420 -2380 3460 -2375
rect 3420 -2410 3425 -2380
rect 3425 -2410 3455 -2380
rect 3455 -2410 3460 -2380
rect 3420 -2415 3460 -2410
rect 3420 -2445 3460 -2440
rect 3420 -2475 3425 -2445
rect 3425 -2475 3455 -2445
rect 3455 -2475 3460 -2445
rect 3420 -2480 3460 -2475
rect 3420 -2505 3460 -2500
rect 3420 -2535 3425 -2505
rect 3425 -2535 3455 -2505
rect 3455 -2535 3460 -2505
rect 3420 -2540 3460 -2535
rect 3420 -2570 3460 -2565
rect 3420 -2600 3425 -2570
rect 3425 -2600 3455 -2570
rect 3455 -2600 3460 -2570
rect 3420 -2605 3460 -2600
rect 3420 -2640 3460 -2635
rect 3420 -2670 3425 -2640
rect 3425 -2670 3455 -2640
rect 3455 -2670 3460 -2640
rect 3420 -2675 3460 -2670
rect 3420 -2710 3460 -2705
rect 3420 -2740 3425 -2710
rect 3425 -2740 3455 -2710
rect 3455 -2740 3460 -2710
rect 3420 -2745 3460 -2740
rect 3420 -2780 3460 -2775
rect 3420 -2810 3425 -2780
rect 3425 -2810 3455 -2780
rect 3455 -2810 3460 -2780
rect 3420 -2815 3460 -2810
rect 3420 -2845 3460 -2840
rect 3420 -2875 3425 -2845
rect 3425 -2875 3455 -2845
rect 3455 -2875 3460 -2845
rect 3420 -2880 3460 -2875
rect 3770 -1305 3810 -1300
rect 3770 -1335 3775 -1305
rect 3775 -1335 3805 -1305
rect 3805 -1335 3810 -1305
rect 3770 -1340 3810 -1335
rect 3770 -1370 3810 -1365
rect 3770 -1400 3775 -1370
rect 3775 -1400 3805 -1370
rect 3805 -1400 3810 -1370
rect 3770 -1405 3810 -1400
rect 3770 -1440 3810 -1435
rect 3770 -1470 3775 -1440
rect 3775 -1470 3805 -1440
rect 3805 -1470 3810 -1440
rect 3770 -1475 3810 -1470
rect 3770 -1510 3810 -1505
rect 3770 -1540 3775 -1510
rect 3775 -1540 3805 -1510
rect 3805 -1540 3810 -1510
rect 3770 -1545 3810 -1540
rect 3770 -1580 3810 -1575
rect 3770 -1610 3775 -1580
rect 3775 -1610 3805 -1580
rect 3805 -1610 3810 -1580
rect 3770 -1615 3810 -1610
rect 3770 -1645 3810 -1640
rect 3770 -1675 3775 -1645
rect 3775 -1675 3805 -1645
rect 3805 -1675 3810 -1645
rect 3770 -1680 3810 -1675
rect 3770 -1705 3810 -1700
rect 3770 -1735 3775 -1705
rect 3775 -1735 3805 -1705
rect 3805 -1735 3810 -1705
rect 3770 -1740 3810 -1735
rect 3770 -1770 3810 -1765
rect 3770 -1800 3775 -1770
rect 3775 -1800 3805 -1770
rect 3805 -1800 3810 -1770
rect 3770 -1805 3810 -1800
rect 3770 -1840 3810 -1835
rect 3770 -1870 3775 -1840
rect 3775 -1870 3805 -1840
rect 3805 -1870 3810 -1840
rect 3770 -1875 3810 -1870
rect 3770 -1910 3810 -1905
rect 3770 -1940 3775 -1910
rect 3775 -1940 3805 -1910
rect 3805 -1940 3810 -1910
rect 3770 -1945 3810 -1940
rect 3770 -1980 3810 -1975
rect 3770 -2010 3775 -1980
rect 3775 -2010 3805 -1980
rect 3805 -2010 3810 -1980
rect 3770 -2015 3810 -2010
rect 3770 -2045 3810 -2040
rect 3770 -2075 3775 -2045
rect 3775 -2075 3805 -2045
rect 3805 -2075 3810 -2045
rect 3770 -2080 3810 -2075
rect 3770 -2105 3810 -2100
rect 3770 -2135 3775 -2105
rect 3775 -2135 3805 -2105
rect 3805 -2135 3810 -2105
rect 3770 -2140 3810 -2135
rect 3770 -2170 3810 -2165
rect 3770 -2200 3775 -2170
rect 3775 -2200 3805 -2170
rect 3805 -2200 3810 -2170
rect 3770 -2205 3810 -2200
rect 3770 -2240 3810 -2235
rect 3770 -2270 3775 -2240
rect 3775 -2270 3805 -2240
rect 3805 -2270 3810 -2240
rect 3770 -2275 3810 -2270
rect 3770 -2310 3810 -2305
rect 3770 -2340 3775 -2310
rect 3775 -2340 3805 -2310
rect 3805 -2340 3810 -2310
rect 3770 -2345 3810 -2340
rect 3770 -2380 3810 -2375
rect 3770 -2410 3775 -2380
rect 3775 -2410 3805 -2380
rect 3805 -2410 3810 -2380
rect 3770 -2415 3810 -2410
rect 3770 -2445 3810 -2440
rect 3770 -2475 3775 -2445
rect 3775 -2475 3805 -2445
rect 3805 -2475 3810 -2445
rect 3770 -2480 3810 -2475
rect 3770 -2505 3810 -2500
rect 3770 -2535 3775 -2505
rect 3775 -2535 3805 -2505
rect 3805 -2535 3810 -2505
rect 3770 -2540 3810 -2535
rect 3770 -2570 3810 -2565
rect 3770 -2600 3775 -2570
rect 3775 -2600 3805 -2570
rect 3805 -2600 3810 -2570
rect 3770 -2605 3810 -2600
rect 3770 -2640 3810 -2635
rect 3770 -2670 3775 -2640
rect 3775 -2670 3805 -2640
rect 3805 -2670 3810 -2640
rect 3770 -2675 3810 -2670
rect 3770 -2710 3810 -2705
rect 3770 -2740 3775 -2710
rect 3775 -2740 3805 -2710
rect 3805 -2740 3810 -2710
rect 3770 -2745 3810 -2740
rect 3770 -2780 3810 -2775
rect 3770 -2810 3775 -2780
rect 3775 -2810 3805 -2780
rect 3805 -2810 3810 -2780
rect 3770 -2815 3810 -2810
rect 3770 -2845 3810 -2840
rect 3770 -2875 3775 -2845
rect 3775 -2875 3805 -2845
rect 3805 -2875 3810 -2845
rect 3770 -2880 3810 -2875
rect 4120 -1305 4160 -1300
rect 4120 -1335 4125 -1305
rect 4125 -1335 4155 -1305
rect 4155 -1335 4160 -1305
rect 4120 -1340 4160 -1335
rect 4120 -1370 4160 -1365
rect 4120 -1400 4125 -1370
rect 4125 -1400 4155 -1370
rect 4155 -1400 4160 -1370
rect 4120 -1405 4160 -1400
rect 4120 -1440 4160 -1435
rect 4120 -1470 4125 -1440
rect 4125 -1470 4155 -1440
rect 4155 -1470 4160 -1440
rect 4120 -1475 4160 -1470
rect 4120 -1510 4160 -1505
rect 4120 -1540 4125 -1510
rect 4125 -1540 4155 -1510
rect 4155 -1540 4160 -1510
rect 4120 -1545 4160 -1540
rect 4120 -1580 4160 -1575
rect 4120 -1610 4125 -1580
rect 4125 -1610 4155 -1580
rect 4155 -1610 4160 -1580
rect 4120 -1615 4160 -1610
rect 4120 -1645 4160 -1640
rect 4120 -1675 4125 -1645
rect 4125 -1675 4155 -1645
rect 4155 -1675 4160 -1645
rect 4120 -1680 4160 -1675
rect 4120 -1705 4160 -1700
rect 4120 -1735 4125 -1705
rect 4125 -1735 4155 -1705
rect 4155 -1735 4160 -1705
rect 4120 -1740 4160 -1735
rect 4120 -1770 4160 -1765
rect 4120 -1800 4125 -1770
rect 4125 -1800 4155 -1770
rect 4155 -1800 4160 -1770
rect 4120 -1805 4160 -1800
rect 4120 -1840 4160 -1835
rect 4120 -1870 4125 -1840
rect 4125 -1870 4155 -1840
rect 4155 -1870 4160 -1840
rect 4120 -1875 4160 -1870
rect 4120 -1910 4160 -1905
rect 4120 -1940 4125 -1910
rect 4125 -1940 4155 -1910
rect 4155 -1940 4160 -1910
rect 4120 -1945 4160 -1940
rect 4120 -1980 4160 -1975
rect 4120 -2010 4125 -1980
rect 4125 -2010 4155 -1980
rect 4155 -2010 4160 -1980
rect 4120 -2015 4160 -2010
rect 4120 -2045 4160 -2040
rect 4120 -2075 4125 -2045
rect 4125 -2075 4155 -2045
rect 4155 -2075 4160 -2045
rect 4120 -2080 4160 -2075
rect 4120 -2105 4160 -2100
rect 4120 -2135 4125 -2105
rect 4125 -2135 4155 -2105
rect 4155 -2135 4160 -2105
rect 4120 -2140 4160 -2135
rect 4120 -2170 4160 -2165
rect 4120 -2200 4125 -2170
rect 4125 -2200 4155 -2170
rect 4155 -2200 4160 -2170
rect 4120 -2205 4160 -2200
rect 4120 -2240 4160 -2235
rect 4120 -2270 4125 -2240
rect 4125 -2270 4155 -2240
rect 4155 -2270 4160 -2240
rect 4120 -2275 4160 -2270
rect 4120 -2310 4160 -2305
rect 4120 -2340 4125 -2310
rect 4125 -2340 4155 -2310
rect 4155 -2340 4160 -2310
rect 4120 -2345 4160 -2340
rect 4120 -2380 4160 -2375
rect 4120 -2410 4125 -2380
rect 4125 -2410 4155 -2380
rect 4155 -2410 4160 -2380
rect 4120 -2415 4160 -2410
rect 4120 -2445 4160 -2440
rect 4120 -2475 4125 -2445
rect 4125 -2475 4155 -2445
rect 4155 -2475 4160 -2445
rect 4120 -2480 4160 -2475
rect 4120 -2505 4160 -2500
rect 4120 -2535 4125 -2505
rect 4125 -2535 4155 -2505
rect 4155 -2535 4160 -2505
rect 4120 -2540 4160 -2535
rect 4120 -2570 4160 -2565
rect 4120 -2600 4125 -2570
rect 4125 -2600 4155 -2570
rect 4155 -2600 4160 -2570
rect 4120 -2605 4160 -2600
rect 4120 -2640 4160 -2635
rect 4120 -2670 4125 -2640
rect 4125 -2670 4155 -2640
rect 4155 -2670 4160 -2640
rect 4120 -2675 4160 -2670
rect 4120 -2710 4160 -2705
rect 4120 -2740 4125 -2710
rect 4125 -2740 4155 -2710
rect 4155 -2740 4160 -2710
rect 4120 -2745 4160 -2740
rect 4120 -2780 4160 -2775
rect 4120 -2810 4125 -2780
rect 4125 -2810 4155 -2780
rect 4155 -2810 4160 -2780
rect 4120 -2815 4160 -2810
rect 4120 -2845 4160 -2840
rect 4120 -2875 4125 -2845
rect 4125 -2875 4155 -2845
rect 4155 -2875 4160 -2845
rect 4120 -2880 4160 -2875
rect 4470 -1305 4510 -1300
rect 4470 -1335 4475 -1305
rect 4475 -1335 4505 -1305
rect 4505 -1335 4510 -1305
rect 4470 -1340 4510 -1335
rect 4470 -1370 4510 -1365
rect 4470 -1400 4475 -1370
rect 4475 -1400 4505 -1370
rect 4505 -1400 4510 -1370
rect 4470 -1405 4510 -1400
rect 4470 -1440 4510 -1435
rect 4470 -1470 4475 -1440
rect 4475 -1470 4505 -1440
rect 4505 -1470 4510 -1440
rect 4470 -1475 4510 -1470
rect 4470 -1510 4510 -1505
rect 4470 -1540 4475 -1510
rect 4475 -1540 4505 -1510
rect 4505 -1540 4510 -1510
rect 4470 -1545 4510 -1540
rect 4470 -1580 4510 -1575
rect 4470 -1610 4475 -1580
rect 4475 -1610 4505 -1580
rect 4505 -1610 4510 -1580
rect 4470 -1615 4510 -1610
rect 4470 -1645 4510 -1640
rect 4470 -1675 4475 -1645
rect 4475 -1675 4505 -1645
rect 4505 -1675 4510 -1645
rect 4470 -1680 4510 -1675
rect 4470 -1705 4510 -1700
rect 4470 -1735 4475 -1705
rect 4475 -1735 4505 -1705
rect 4505 -1735 4510 -1705
rect 4470 -1740 4510 -1735
rect 4470 -1770 4510 -1765
rect 4470 -1800 4475 -1770
rect 4475 -1800 4505 -1770
rect 4505 -1800 4510 -1770
rect 4470 -1805 4510 -1800
rect 4470 -1840 4510 -1835
rect 4470 -1870 4475 -1840
rect 4475 -1870 4505 -1840
rect 4505 -1870 4510 -1840
rect 4470 -1875 4510 -1870
rect 4470 -1910 4510 -1905
rect 4470 -1940 4475 -1910
rect 4475 -1940 4505 -1910
rect 4505 -1940 4510 -1910
rect 4470 -1945 4510 -1940
rect 4470 -1980 4510 -1975
rect 4470 -2010 4475 -1980
rect 4475 -2010 4505 -1980
rect 4505 -2010 4510 -1980
rect 4470 -2015 4510 -2010
rect 4470 -2045 4510 -2040
rect 4470 -2075 4475 -2045
rect 4475 -2075 4505 -2045
rect 4505 -2075 4510 -2045
rect 4470 -2080 4510 -2075
rect 4470 -2105 4510 -2100
rect 4470 -2135 4475 -2105
rect 4475 -2135 4505 -2105
rect 4505 -2135 4510 -2105
rect 4470 -2140 4510 -2135
rect 4470 -2170 4510 -2165
rect 4470 -2200 4475 -2170
rect 4475 -2200 4505 -2170
rect 4505 -2200 4510 -2170
rect 4470 -2205 4510 -2200
rect 4470 -2240 4510 -2235
rect 4470 -2270 4475 -2240
rect 4475 -2270 4505 -2240
rect 4505 -2270 4510 -2240
rect 4470 -2275 4510 -2270
rect 4470 -2310 4510 -2305
rect 4470 -2340 4475 -2310
rect 4475 -2340 4505 -2310
rect 4505 -2340 4510 -2310
rect 4470 -2345 4510 -2340
rect 4470 -2380 4510 -2375
rect 4470 -2410 4475 -2380
rect 4475 -2410 4505 -2380
rect 4505 -2410 4510 -2380
rect 4470 -2415 4510 -2410
rect 4470 -2445 4510 -2440
rect 4470 -2475 4475 -2445
rect 4475 -2475 4505 -2445
rect 4505 -2475 4510 -2445
rect 4470 -2480 4510 -2475
rect 4470 -2505 4510 -2500
rect 4470 -2535 4475 -2505
rect 4475 -2535 4505 -2505
rect 4505 -2535 4510 -2505
rect 4470 -2540 4510 -2535
rect 4470 -2570 4510 -2565
rect 4470 -2600 4475 -2570
rect 4475 -2600 4505 -2570
rect 4505 -2600 4510 -2570
rect 4470 -2605 4510 -2600
rect 4470 -2640 4510 -2635
rect 4470 -2670 4475 -2640
rect 4475 -2670 4505 -2640
rect 4505 -2670 4510 -2640
rect 4470 -2675 4510 -2670
rect 4470 -2710 4510 -2705
rect 4470 -2740 4475 -2710
rect 4475 -2740 4505 -2710
rect 4505 -2740 4510 -2710
rect 4470 -2745 4510 -2740
rect 4470 -2780 4510 -2775
rect 4470 -2810 4475 -2780
rect 4475 -2810 4505 -2780
rect 4505 -2810 4510 -2780
rect 4470 -2815 4510 -2810
rect 4470 -2845 4510 -2840
rect 4470 -2875 4475 -2845
rect 4475 -2875 4505 -2845
rect 4505 -2875 4510 -2845
rect 4470 -2880 4510 -2875
rect 4820 -1305 4860 -1300
rect 4820 -1335 4825 -1305
rect 4825 -1335 4855 -1305
rect 4855 -1335 4860 -1305
rect 4820 -1340 4860 -1335
rect 4820 -1370 4860 -1365
rect 4820 -1400 4825 -1370
rect 4825 -1400 4855 -1370
rect 4855 -1400 4860 -1370
rect 4820 -1405 4860 -1400
rect 4820 -1440 4860 -1435
rect 4820 -1470 4825 -1440
rect 4825 -1470 4855 -1440
rect 4855 -1470 4860 -1440
rect 4820 -1475 4860 -1470
rect 4820 -1510 4860 -1505
rect 4820 -1540 4825 -1510
rect 4825 -1540 4855 -1510
rect 4855 -1540 4860 -1510
rect 4820 -1545 4860 -1540
rect 4820 -1580 4860 -1575
rect 4820 -1610 4825 -1580
rect 4825 -1610 4855 -1580
rect 4855 -1610 4860 -1580
rect 4820 -1615 4860 -1610
rect 4820 -1645 4860 -1640
rect 4820 -1675 4825 -1645
rect 4825 -1675 4855 -1645
rect 4855 -1675 4860 -1645
rect 4820 -1680 4860 -1675
rect 4820 -1705 4860 -1700
rect 4820 -1735 4825 -1705
rect 4825 -1735 4855 -1705
rect 4855 -1735 4860 -1705
rect 4820 -1740 4860 -1735
rect 4820 -1770 4860 -1765
rect 4820 -1800 4825 -1770
rect 4825 -1800 4855 -1770
rect 4855 -1800 4860 -1770
rect 4820 -1805 4860 -1800
rect 4820 -1840 4860 -1835
rect 4820 -1870 4825 -1840
rect 4825 -1870 4855 -1840
rect 4855 -1870 4860 -1840
rect 4820 -1875 4860 -1870
rect 4820 -1910 4860 -1905
rect 4820 -1940 4825 -1910
rect 4825 -1940 4855 -1910
rect 4855 -1940 4860 -1910
rect 4820 -1945 4860 -1940
rect 4820 -1980 4860 -1975
rect 4820 -2010 4825 -1980
rect 4825 -2010 4855 -1980
rect 4855 -2010 4860 -1980
rect 4820 -2015 4860 -2010
rect 4820 -2045 4860 -2040
rect 4820 -2075 4825 -2045
rect 4825 -2075 4855 -2045
rect 4855 -2075 4860 -2045
rect 4820 -2080 4860 -2075
rect 4820 -2105 4860 -2100
rect 4820 -2135 4825 -2105
rect 4825 -2135 4855 -2105
rect 4855 -2135 4860 -2105
rect 4820 -2140 4860 -2135
rect 4820 -2170 4860 -2165
rect 4820 -2200 4825 -2170
rect 4825 -2200 4855 -2170
rect 4855 -2200 4860 -2170
rect 4820 -2205 4860 -2200
rect 4820 -2240 4860 -2235
rect 4820 -2270 4825 -2240
rect 4825 -2270 4855 -2240
rect 4855 -2270 4860 -2240
rect 4820 -2275 4860 -2270
rect 4820 -2310 4860 -2305
rect 4820 -2340 4825 -2310
rect 4825 -2340 4855 -2310
rect 4855 -2340 4860 -2310
rect 4820 -2345 4860 -2340
rect 4820 -2380 4860 -2375
rect 4820 -2410 4825 -2380
rect 4825 -2410 4855 -2380
rect 4855 -2410 4860 -2380
rect 4820 -2415 4860 -2410
rect 4820 -2445 4860 -2440
rect 4820 -2475 4825 -2445
rect 4825 -2475 4855 -2445
rect 4855 -2475 4860 -2445
rect 4820 -2480 4860 -2475
rect 4820 -2505 4860 -2500
rect 4820 -2535 4825 -2505
rect 4825 -2535 4855 -2505
rect 4855 -2535 4860 -2505
rect 4820 -2540 4860 -2535
rect 4820 -2570 4860 -2565
rect 4820 -2600 4825 -2570
rect 4825 -2600 4855 -2570
rect 4855 -2600 4860 -2570
rect 4820 -2605 4860 -2600
rect 4820 -2640 4860 -2635
rect 4820 -2670 4825 -2640
rect 4825 -2670 4855 -2640
rect 4855 -2670 4860 -2640
rect 4820 -2675 4860 -2670
rect 4820 -2710 4860 -2705
rect 4820 -2740 4825 -2710
rect 4825 -2740 4855 -2710
rect 4855 -2740 4860 -2710
rect 4820 -2745 4860 -2740
rect 4820 -2780 4860 -2775
rect 4820 -2810 4825 -2780
rect 4825 -2810 4855 -2780
rect 4855 -2810 4860 -2780
rect 4820 -2815 4860 -2810
rect 4820 -2845 4860 -2840
rect 4820 -2875 4825 -2845
rect 4825 -2875 4855 -2845
rect 4855 -2875 4860 -2845
rect 4820 -2880 4860 -2875
rect 5170 -1305 5210 -1300
rect 5170 -1335 5175 -1305
rect 5175 -1335 5205 -1305
rect 5205 -1335 5210 -1305
rect 5170 -1340 5210 -1335
rect 5170 -1370 5210 -1365
rect 5170 -1400 5175 -1370
rect 5175 -1400 5205 -1370
rect 5205 -1400 5210 -1370
rect 5170 -1405 5210 -1400
rect 5170 -1440 5210 -1435
rect 5170 -1470 5175 -1440
rect 5175 -1470 5205 -1440
rect 5205 -1470 5210 -1440
rect 5170 -1475 5210 -1470
rect 5170 -1510 5210 -1505
rect 5170 -1540 5175 -1510
rect 5175 -1540 5205 -1510
rect 5205 -1540 5210 -1510
rect 5170 -1545 5210 -1540
rect 5170 -1580 5210 -1575
rect 5170 -1610 5175 -1580
rect 5175 -1610 5205 -1580
rect 5205 -1610 5210 -1580
rect 5170 -1615 5210 -1610
rect 5170 -1645 5210 -1640
rect 5170 -1675 5175 -1645
rect 5175 -1675 5205 -1645
rect 5205 -1675 5210 -1645
rect 5170 -1680 5210 -1675
rect 5170 -1705 5210 -1700
rect 5170 -1735 5175 -1705
rect 5175 -1735 5205 -1705
rect 5205 -1735 5210 -1705
rect 5170 -1740 5210 -1735
rect 5170 -1770 5210 -1765
rect 5170 -1800 5175 -1770
rect 5175 -1800 5205 -1770
rect 5205 -1800 5210 -1770
rect 5170 -1805 5210 -1800
rect 5170 -1840 5210 -1835
rect 5170 -1870 5175 -1840
rect 5175 -1870 5205 -1840
rect 5205 -1870 5210 -1840
rect 5170 -1875 5210 -1870
rect 5170 -1910 5210 -1905
rect 5170 -1940 5175 -1910
rect 5175 -1940 5205 -1910
rect 5205 -1940 5210 -1910
rect 5170 -1945 5210 -1940
rect 5170 -1980 5210 -1975
rect 5170 -2010 5175 -1980
rect 5175 -2010 5205 -1980
rect 5205 -2010 5210 -1980
rect 5170 -2015 5210 -2010
rect 5170 -2045 5210 -2040
rect 5170 -2075 5175 -2045
rect 5175 -2075 5205 -2045
rect 5205 -2075 5210 -2045
rect 5170 -2080 5210 -2075
rect 5170 -2105 5210 -2100
rect 5170 -2135 5175 -2105
rect 5175 -2135 5205 -2105
rect 5205 -2135 5210 -2105
rect 5170 -2140 5210 -2135
rect 5170 -2170 5210 -2165
rect 5170 -2200 5175 -2170
rect 5175 -2200 5205 -2170
rect 5205 -2200 5210 -2170
rect 5170 -2205 5210 -2200
rect 5170 -2240 5210 -2235
rect 5170 -2270 5175 -2240
rect 5175 -2270 5205 -2240
rect 5205 -2270 5210 -2240
rect 5170 -2275 5210 -2270
rect 5170 -2310 5210 -2305
rect 5170 -2340 5175 -2310
rect 5175 -2340 5205 -2310
rect 5205 -2340 5210 -2310
rect 5170 -2345 5210 -2340
rect 5170 -2380 5210 -2375
rect 5170 -2410 5175 -2380
rect 5175 -2410 5205 -2380
rect 5205 -2410 5210 -2380
rect 5170 -2415 5210 -2410
rect 5170 -2445 5210 -2440
rect 5170 -2475 5175 -2445
rect 5175 -2475 5205 -2445
rect 5205 -2475 5210 -2445
rect 5170 -2480 5210 -2475
rect 5170 -2505 5210 -2500
rect 5170 -2535 5175 -2505
rect 5175 -2535 5205 -2505
rect 5205 -2535 5210 -2505
rect 5170 -2540 5210 -2535
rect 5170 -2570 5210 -2565
rect 5170 -2600 5175 -2570
rect 5175 -2600 5205 -2570
rect 5205 -2600 5210 -2570
rect 5170 -2605 5210 -2600
rect 5170 -2640 5210 -2635
rect 5170 -2670 5175 -2640
rect 5175 -2670 5205 -2640
rect 5205 -2670 5210 -2640
rect 5170 -2675 5210 -2670
rect 5170 -2710 5210 -2705
rect 5170 -2740 5175 -2710
rect 5175 -2740 5205 -2710
rect 5205 -2740 5210 -2710
rect 5170 -2745 5210 -2740
rect 5170 -2780 5210 -2775
rect 5170 -2810 5175 -2780
rect 5175 -2810 5205 -2780
rect 5205 -2810 5210 -2780
rect 5170 -2815 5210 -2810
rect 5170 -2845 5210 -2840
rect 5170 -2875 5175 -2845
rect 5175 -2875 5205 -2845
rect 5205 -2875 5210 -2845
rect 5170 -2880 5210 -2875
rect 5520 -1305 5560 -1300
rect 5520 -1335 5525 -1305
rect 5525 -1335 5555 -1305
rect 5555 -1335 5560 -1305
rect 5520 -1340 5560 -1335
rect 5520 -1370 5560 -1365
rect 5520 -1400 5525 -1370
rect 5525 -1400 5555 -1370
rect 5555 -1400 5560 -1370
rect 5520 -1405 5560 -1400
rect 5520 -1440 5560 -1435
rect 5520 -1470 5525 -1440
rect 5525 -1470 5555 -1440
rect 5555 -1470 5560 -1440
rect 5520 -1475 5560 -1470
rect 5520 -1510 5560 -1505
rect 5520 -1540 5525 -1510
rect 5525 -1540 5555 -1510
rect 5555 -1540 5560 -1510
rect 5520 -1545 5560 -1540
rect 5520 -1580 5560 -1575
rect 5520 -1610 5525 -1580
rect 5525 -1610 5555 -1580
rect 5555 -1610 5560 -1580
rect 5520 -1615 5560 -1610
rect 5520 -1645 5560 -1640
rect 5520 -1675 5525 -1645
rect 5525 -1675 5555 -1645
rect 5555 -1675 5560 -1645
rect 5520 -1680 5560 -1675
rect 5520 -1705 5560 -1700
rect 5520 -1735 5525 -1705
rect 5525 -1735 5555 -1705
rect 5555 -1735 5560 -1705
rect 5520 -1740 5560 -1735
rect 5520 -1770 5560 -1765
rect 5520 -1800 5525 -1770
rect 5525 -1800 5555 -1770
rect 5555 -1800 5560 -1770
rect 5520 -1805 5560 -1800
rect 5520 -1840 5560 -1835
rect 5520 -1870 5525 -1840
rect 5525 -1870 5555 -1840
rect 5555 -1870 5560 -1840
rect 5520 -1875 5560 -1870
rect 5520 -1910 5560 -1905
rect 5520 -1940 5525 -1910
rect 5525 -1940 5555 -1910
rect 5555 -1940 5560 -1910
rect 5520 -1945 5560 -1940
rect 5520 -1980 5560 -1975
rect 5520 -2010 5525 -1980
rect 5525 -2010 5555 -1980
rect 5555 -2010 5560 -1980
rect 5520 -2015 5560 -2010
rect 5520 -2045 5560 -2040
rect 5520 -2075 5525 -2045
rect 5525 -2075 5555 -2045
rect 5555 -2075 5560 -2045
rect 5520 -2080 5560 -2075
rect 5520 -2105 5560 -2100
rect 5520 -2135 5525 -2105
rect 5525 -2135 5555 -2105
rect 5555 -2135 5560 -2105
rect 5520 -2140 5560 -2135
rect 5520 -2170 5560 -2165
rect 5520 -2200 5525 -2170
rect 5525 -2200 5555 -2170
rect 5555 -2200 5560 -2170
rect 5520 -2205 5560 -2200
rect 5520 -2240 5560 -2235
rect 5520 -2270 5525 -2240
rect 5525 -2270 5555 -2240
rect 5555 -2270 5560 -2240
rect 5520 -2275 5560 -2270
rect 5520 -2310 5560 -2305
rect 5520 -2340 5525 -2310
rect 5525 -2340 5555 -2310
rect 5555 -2340 5560 -2310
rect 5520 -2345 5560 -2340
rect 5520 -2380 5560 -2375
rect 5520 -2410 5525 -2380
rect 5525 -2410 5555 -2380
rect 5555 -2410 5560 -2380
rect 5520 -2415 5560 -2410
rect 5520 -2445 5560 -2440
rect 5520 -2475 5525 -2445
rect 5525 -2475 5555 -2445
rect 5555 -2475 5560 -2445
rect 5520 -2480 5560 -2475
rect 5520 -2505 5560 -2500
rect 5520 -2535 5525 -2505
rect 5525 -2535 5555 -2505
rect 5555 -2535 5560 -2505
rect 5520 -2540 5560 -2535
rect 5520 -2570 5560 -2565
rect 5520 -2600 5525 -2570
rect 5525 -2600 5555 -2570
rect 5555 -2600 5560 -2570
rect 5520 -2605 5560 -2600
rect 5520 -2640 5560 -2635
rect 5520 -2670 5525 -2640
rect 5525 -2670 5555 -2640
rect 5555 -2670 5560 -2640
rect 5520 -2675 5560 -2670
rect 5520 -2710 5560 -2705
rect 5520 -2740 5525 -2710
rect 5525 -2740 5555 -2710
rect 5555 -2740 5560 -2710
rect 5520 -2745 5560 -2740
rect 5520 -2780 5560 -2775
rect 5520 -2810 5525 -2780
rect 5525 -2810 5555 -2780
rect 5555 -2810 5560 -2780
rect 5520 -2815 5560 -2810
rect 5520 -2845 5560 -2840
rect 5520 -2875 5525 -2845
rect 5525 -2875 5555 -2845
rect 5555 -2875 5560 -2845
rect 5520 -2880 5560 -2875
rect 5870 -1305 5910 -1300
rect 5870 -1335 5875 -1305
rect 5875 -1335 5905 -1305
rect 5905 -1335 5910 -1305
rect 5870 -1340 5910 -1335
rect 5870 -1370 5910 -1365
rect 5870 -1400 5875 -1370
rect 5875 -1400 5905 -1370
rect 5905 -1400 5910 -1370
rect 5870 -1405 5910 -1400
rect 5870 -1440 5910 -1435
rect 5870 -1470 5875 -1440
rect 5875 -1470 5905 -1440
rect 5905 -1470 5910 -1440
rect 5870 -1475 5910 -1470
rect 5870 -1510 5910 -1505
rect 5870 -1540 5875 -1510
rect 5875 -1540 5905 -1510
rect 5905 -1540 5910 -1510
rect 5870 -1545 5910 -1540
rect 5870 -1580 5910 -1575
rect 5870 -1610 5875 -1580
rect 5875 -1610 5905 -1580
rect 5905 -1610 5910 -1580
rect 5870 -1615 5910 -1610
rect 5870 -1645 5910 -1640
rect 5870 -1675 5875 -1645
rect 5875 -1675 5905 -1645
rect 5905 -1675 5910 -1645
rect 5870 -1680 5910 -1675
rect 5870 -1705 5910 -1700
rect 5870 -1735 5875 -1705
rect 5875 -1735 5905 -1705
rect 5905 -1735 5910 -1705
rect 5870 -1740 5910 -1735
rect 5870 -1770 5910 -1765
rect 5870 -1800 5875 -1770
rect 5875 -1800 5905 -1770
rect 5905 -1800 5910 -1770
rect 5870 -1805 5910 -1800
rect 5870 -1840 5910 -1835
rect 5870 -1870 5875 -1840
rect 5875 -1870 5905 -1840
rect 5905 -1870 5910 -1840
rect 5870 -1875 5910 -1870
rect 5870 -1910 5910 -1905
rect 5870 -1940 5875 -1910
rect 5875 -1940 5905 -1910
rect 5905 -1940 5910 -1910
rect 5870 -1945 5910 -1940
rect 5870 -1980 5910 -1975
rect 5870 -2010 5875 -1980
rect 5875 -2010 5905 -1980
rect 5905 -2010 5910 -1980
rect 5870 -2015 5910 -2010
rect 5870 -2045 5910 -2040
rect 5870 -2075 5875 -2045
rect 5875 -2075 5905 -2045
rect 5905 -2075 5910 -2045
rect 5870 -2080 5910 -2075
rect 5870 -2105 5910 -2100
rect 5870 -2135 5875 -2105
rect 5875 -2135 5905 -2105
rect 5905 -2135 5910 -2105
rect 5870 -2140 5910 -2135
rect 5870 -2170 5910 -2165
rect 5870 -2200 5875 -2170
rect 5875 -2200 5905 -2170
rect 5905 -2200 5910 -2170
rect 5870 -2205 5910 -2200
rect 5870 -2240 5910 -2235
rect 5870 -2270 5875 -2240
rect 5875 -2270 5905 -2240
rect 5905 -2270 5910 -2240
rect 5870 -2275 5910 -2270
rect 5870 -2310 5910 -2305
rect 5870 -2340 5875 -2310
rect 5875 -2340 5905 -2310
rect 5905 -2340 5910 -2310
rect 5870 -2345 5910 -2340
rect 5870 -2380 5910 -2375
rect 5870 -2410 5875 -2380
rect 5875 -2410 5905 -2380
rect 5905 -2410 5910 -2380
rect 5870 -2415 5910 -2410
rect 5870 -2445 5910 -2440
rect 5870 -2475 5875 -2445
rect 5875 -2475 5905 -2445
rect 5905 -2475 5910 -2445
rect 5870 -2480 5910 -2475
rect 5870 -2505 5910 -2500
rect 5870 -2535 5875 -2505
rect 5875 -2535 5905 -2505
rect 5905 -2535 5910 -2505
rect 5870 -2540 5910 -2535
rect 5870 -2570 5910 -2565
rect 5870 -2600 5875 -2570
rect 5875 -2600 5905 -2570
rect 5905 -2600 5910 -2570
rect 5870 -2605 5910 -2600
rect 5870 -2640 5910 -2635
rect 5870 -2670 5875 -2640
rect 5875 -2670 5905 -2640
rect 5905 -2670 5910 -2640
rect 5870 -2675 5910 -2670
rect 5870 -2710 5910 -2705
rect 5870 -2740 5875 -2710
rect 5875 -2740 5905 -2710
rect 5905 -2740 5910 -2710
rect 5870 -2745 5910 -2740
rect 5870 -2780 5910 -2775
rect 5870 -2810 5875 -2780
rect 5875 -2810 5905 -2780
rect 5905 -2810 5910 -2780
rect 5870 -2815 5910 -2810
rect 5870 -2845 5910 -2840
rect 5870 -2875 5875 -2845
rect 5875 -2875 5905 -2845
rect 5905 -2875 5910 -2845
rect 5870 -2880 5910 -2875
rect 6220 -1305 6260 -1300
rect 6220 -1335 6225 -1305
rect 6225 -1335 6255 -1305
rect 6255 -1335 6260 -1305
rect 6220 -1340 6260 -1335
rect 6220 -1370 6260 -1365
rect 6220 -1400 6225 -1370
rect 6225 -1400 6255 -1370
rect 6255 -1400 6260 -1370
rect 6220 -1405 6260 -1400
rect 6220 -1440 6260 -1435
rect 6220 -1470 6225 -1440
rect 6225 -1470 6255 -1440
rect 6255 -1470 6260 -1440
rect 6220 -1475 6260 -1470
rect 6220 -1510 6260 -1505
rect 6220 -1540 6225 -1510
rect 6225 -1540 6255 -1510
rect 6255 -1540 6260 -1510
rect 6220 -1545 6260 -1540
rect 6220 -1580 6260 -1575
rect 6220 -1610 6225 -1580
rect 6225 -1610 6255 -1580
rect 6255 -1610 6260 -1580
rect 6220 -1615 6260 -1610
rect 6220 -1645 6260 -1640
rect 6220 -1675 6225 -1645
rect 6225 -1675 6255 -1645
rect 6255 -1675 6260 -1645
rect 6220 -1680 6260 -1675
rect 6220 -1705 6260 -1700
rect 6220 -1735 6225 -1705
rect 6225 -1735 6255 -1705
rect 6255 -1735 6260 -1705
rect 6220 -1740 6260 -1735
rect 6220 -1770 6260 -1765
rect 6220 -1800 6225 -1770
rect 6225 -1800 6255 -1770
rect 6255 -1800 6260 -1770
rect 6220 -1805 6260 -1800
rect 6220 -1840 6260 -1835
rect 6220 -1870 6225 -1840
rect 6225 -1870 6255 -1840
rect 6255 -1870 6260 -1840
rect 6220 -1875 6260 -1870
rect 6220 -1910 6260 -1905
rect 6220 -1940 6225 -1910
rect 6225 -1940 6255 -1910
rect 6255 -1940 6260 -1910
rect 6220 -1945 6260 -1940
rect 6220 -1980 6260 -1975
rect 6220 -2010 6225 -1980
rect 6225 -2010 6255 -1980
rect 6255 -2010 6260 -1980
rect 6220 -2015 6260 -2010
rect 6220 -2045 6260 -2040
rect 6220 -2075 6225 -2045
rect 6225 -2075 6255 -2045
rect 6255 -2075 6260 -2045
rect 6220 -2080 6260 -2075
rect 6220 -2105 6260 -2100
rect 6220 -2135 6225 -2105
rect 6225 -2135 6255 -2105
rect 6255 -2135 6260 -2105
rect 6220 -2140 6260 -2135
rect 6220 -2170 6260 -2165
rect 6220 -2200 6225 -2170
rect 6225 -2200 6255 -2170
rect 6255 -2200 6260 -2170
rect 6220 -2205 6260 -2200
rect 6220 -2240 6260 -2235
rect 6220 -2270 6225 -2240
rect 6225 -2270 6255 -2240
rect 6255 -2270 6260 -2240
rect 6220 -2275 6260 -2270
rect 6220 -2310 6260 -2305
rect 6220 -2340 6225 -2310
rect 6225 -2340 6255 -2310
rect 6255 -2340 6260 -2310
rect 6220 -2345 6260 -2340
rect 6220 -2380 6260 -2375
rect 6220 -2410 6225 -2380
rect 6225 -2410 6255 -2380
rect 6255 -2410 6260 -2380
rect 6220 -2415 6260 -2410
rect 6220 -2445 6260 -2440
rect 6220 -2475 6225 -2445
rect 6225 -2475 6255 -2445
rect 6255 -2475 6260 -2445
rect 6220 -2480 6260 -2475
rect 6220 -2505 6260 -2500
rect 6220 -2535 6225 -2505
rect 6225 -2535 6255 -2505
rect 6255 -2535 6260 -2505
rect 6220 -2540 6260 -2535
rect 6220 -2570 6260 -2565
rect 6220 -2600 6225 -2570
rect 6225 -2600 6255 -2570
rect 6255 -2600 6260 -2570
rect 6220 -2605 6260 -2600
rect 6220 -2640 6260 -2635
rect 6220 -2670 6225 -2640
rect 6225 -2670 6255 -2640
rect 6255 -2670 6260 -2640
rect 6220 -2675 6260 -2670
rect 6220 -2710 6260 -2705
rect 6220 -2740 6225 -2710
rect 6225 -2740 6255 -2710
rect 6255 -2740 6260 -2710
rect 6220 -2745 6260 -2740
rect 6220 -2780 6260 -2775
rect 6220 -2810 6225 -2780
rect 6225 -2810 6255 -2780
rect 6255 -2810 6260 -2780
rect 6220 -2815 6260 -2810
rect 6220 -2845 6260 -2840
rect 6220 -2875 6225 -2845
rect 6225 -2875 6255 -2845
rect 6255 -2875 6260 -2845
rect 6220 -2880 6260 -2875
rect 6570 -1305 6610 -1300
rect 6570 -1335 6575 -1305
rect 6575 -1335 6605 -1305
rect 6605 -1335 6610 -1305
rect 6570 -1340 6610 -1335
rect 6570 -1370 6610 -1365
rect 6570 -1400 6575 -1370
rect 6575 -1400 6605 -1370
rect 6605 -1400 6610 -1370
rect 6570 -1405 6610 -1400
rect 6570 -1440 6610 -1435
rect 6570 -1470 6575 -1440
rect 6575 -1470 6605 -1440
rect 6605 -1470 6610 -1440
rect 6570 -1475 6610 -1470
rect 6570 -1510 6610 -1505
rect 6570 -1540 6575 -1510
rect 6575 -1540 6605 -1510
rect 6605 -1540 6610 -1510
rect 6570 -1545 6610 -1540
rect 6570 -1580 6610 -1575
rect 6570 -1610 6575 -1580
rect 6575 -1610 6605 -1580
rect 6605 -1610 6610 -1580
rect 6570 -1615 6610 -1610
rect 6570 -1645 6610 -1640
rect 6570 -1675 6575 -1645
rect 6575 -1675 6605 -1645
rect 6605 -1675 6610 -1645
rect 6570 -1680 6610 -1675
rect 6570 -1705 6610 -1700
rect 6570 -1735 6575 -1705
rect 6575 -1735 6605 -1705
rect 6605 -1735 6610 -1705
rect 6570 -1740 6610 -1735
rect 6570 -1770 6610 -1765
rect 6570 -1800 6575 -1770
rect 6575 -1800 6605 -1770
rect 6605 -1800 6610 -1770
rect 6570 -1805 6610 -1800
rect 6570 -1840 6610 -1835
rect 6570 -1870 6575 -1840
rect 6575 -1870 6605 -1840
rect 6605 -1870 6610 -1840
rect 6570 -1875 6610 -1870
rect 6570 -1910 6610 -1905
rect 6570 -1940 6575 -1910
rect 6575 -1940 6605 -1910
rect 6605 -1940 6610 -1910
rect 6570 -1945 6610 -1940
rect 6570 -1980 6610 -1975
rect 6570 -2010 6575 -1980
rect 6575 -2010 6605 -1980
rect 6605 -2010 6610 -1980
rect 6570 -2015 6610 -2010
rect 6570 -2045 6610 -2040
rect 6570 -2075 6575 -2045
rect 6575 -2075 6605 -2045
rect 6605 -2075 6610 -2045
rect 6570 -2080 6610 -2075
rect 6570 -2105 6610 -2100
rect 6570 -2135 6575 -2105
rect 6575 -2135 6605 -2105
rect 6605 -2135 6610 -2105
rect 6570 -2140 6610 -2135
rect 6570 -2170 6610 -2165
rect 6570 -2200 6575 -2170
rect 6575 -2200 6605 -2170
rect 6605 -2200 6610 -2170
rect 6570 -2205 6610 -2200
rect 6570 -2240 6610 -2235
rect 6570 -2270 6575 -2240
rect 6575 -2270 6605 -2240
rect 6605 -2270 6610 -2240
rect 6570 -2275 6610 -2270
rect 6570 -2310 6610 -2305
rect 6570 -2340 6575 -2310
rect 6575 -2340 6605 -2310
rect 6605 -2340 6610 -2310
rect 6570 -2345 6610 -2340
rect 6570 -2380 6610 -2375
rect 6570 -2410 6575 -2380
rect 6575 -2410 6605 -2380
rect 6605 -2410 6610 -2380
rect 6570 -2415 6610 -2410
rect 6570 -2445 6610 -2440
rect 6570 -2475 6575 -2445
rect 6575 -2475 6605 -2445
rect 6605 -2475 6610 -2445
rect 6570 -2480 6610 -2475
rect 6570 -2505 6610 -2500
rect 6570 -2535 6575 -2505
rect 6575 -2535 6605 -2505
rect 6605 -2535 6610 -2505
rect 6570 -2540 6610 -2535
rect 6570 -2570 6610 -2565
rect 6570 -2600 6575 -2570
rect 6575 -2600 6605 -2570
rect 6605 -2600 6610 -2570
rect 6570 -2605 6610 -2600
rect 6570 -2640 6610 -2635
rect 6570 -2670 6575 -2640
rect 6575 -2670 6605 -2640
rect 6605 -2670 6610 -2640
rect 6570 -2675 6610 -2670
rect 6570 -2710 6610 -2705
rect 6570 -2740 6575 -2710
rect 6575 -2740 6605 -2710
rect 6605 -2740 6610 -2710
rect 6570 -2745 6610 -2740
rect 6570 -2780 6610 -2775
rect 6570 -2810 6575 -2780
rect 6575 -2810 6605 -2780
rect 6605 -2810 6610 -2780
rect 6570 -2815 6610 -2810
rect 6570 -2845 6610 -2840
rect 6570 -2875 6575 -2845
rect 6575 -2875 6605 -2845
rect 6605 -2875 6610 -2845
rect 6570 -2880 6610 -2875
rect 6920 -1305 6960 -1300
rect 6920 -1335 6925 -1305
rect 6925 -1335 6955 -1305
rect 6955 -1335 6960 -1305
rect 6920 -1340 6960 -1335
rect 6920 -1370 6960 -1365
rect 6920 -1400 6925 -1370
rect 6925 -1400 6955 -1370
rect 6955 -1400 6960 -1370
rect 6920 -1405 6960 -1400
rect 6920 -1440 6960 -1435
rect 6920 -1470 6925 -1440
rect 6925 -1470 6955 -1440
rect 6955 -1470 6960 -1440
rect 6920 -1475 6960 -1470
rect 6920 -1510 6960 -1505
rect 6920 -1540 6925 -1510
rect 6925 -1540 6955 -1510
rect 6955 -1540 6960 -1510
rect 6920 -1545 6960 -1540
rect 6920 -1580 6960 -1575
rect 6920 -1610 6925 -1580
rect 6925 -1610 6955 -1580
rect 6955 -1610 6960 -1580
rect 6920 -1615 6960 -1610
rect 6920 -1645 6960 -1640
rect 6920 -1675 6925 -1645
rect 6925 -1675 6955 -1645
rect 6955 -1675 6960 -1645
rect 6920 -1680 6960 -1675
rect 6920 -1705 6960 -1700
rect 6920 -1735 6925 -1705
rect 6925 -1735 6955 -1705
rect 6955 -1735 6960 -1705
rect 6920 -1740 6960 -1735
rect 6920 -1770 6960 -1765
rect 6920 -1800 6925 -1770
rect 6925 -1800 6955 -1770
rect 6955 -1800 6960 -1770
rect 6920 -1805 6960 -1800
rect 6920 -1840 6960 -1835
rect 6920 -1870 6925 -1840
rect 6925 -1870 6955 -1840
rect 6955 -1870 6960 -1840
rect 6920 -1875 6960 -1870
rect 6920 -1910 6960 -1905
rect 6920 -1940 6925 -1910
rect 6925 -1940 6955 -1910
rect 6955 -1940 6960 -1910
rect 6920 -1945 6960 -1940
rect 6920 -1980 6960 -1975
rect 6920 -2010 6925 -1980
rect 6925 -2010 6955 -1980
rect 6955 -2010 6960 -1980
rect 6920 -2015 6960 -2010
rect 6920 -2045 6960 -2040
rect 6920 -2075 6925 -2045
rect 6925 -2075 6955 -2045
rect 6955 -2075 6960 -2045
rect 6920 -2080 6960 -2075
rect 6920 -2105 6960 -2100
rect 6920 -2135 6925 -2105
rect 6925 -2135 6955 -2105
rect 6955 -2135 6960 -2105
rect 6920 -2140 6960 -2135
rect 6920 -2170 6960 -2165
rect 6920 -2200 6925 -2170
rect 6925 -2200 6955 -2170
rect 6955 -2200 6960 -2170
rect 6920 -2205 6960 -2200
rect 6920 -2240 6960 -2235
rect 6920 -2270 6925 -2240
rect 6925 -2270 6955 -2240
rect 6955 -2270 6960 -2240
rect 6920 -2275 6960 -2270
rect 6920 -2310 6960 -2305
rect 6920 -2340 6925 -2310
rect 6925 -2340 6955 -2310
rect 6955 -2340 6960 -2310
rect 6920 -2345 6960 -2340
rect 6920 -2380 6960 -2375
rect 6920 -2410 6925 -2380
rect 6925 -2410 6955 -2380
rect 6955 -2410 6960 -2380
rect 6920 -2415 6960 -2410
rect 6920 -2445 6960 -2440
rect 6920 -2475 6925 -2445
rect 6925 -2475 6955 -2445
rect 6955 -2475 6960 -2445
rect 6920 -2480 6960 -2475
rect 6920 -2505 6960 -2500
rect 6920 -2535 6925 -2505
rect 6925 -2535 6955 -2505
rect 6955 -2535 6960 -2505
rect 6920 -2540 6960 -2535
rect 6920 -2570 6960 -2565
rect 6920 -2600 6925 -2570
rect 6925 -2600 6955 -2570
rect 6955 -2600 6960 -2570
rect 6920 -2605 6960 -2600
rect 6920 -2640 6960 -2635
rect 6920 -2670 6925 -2640
rect 6925 -2670 6955 -2640
rect 6955 -2670 6960 -2640
rect 6920 -2675 6960 -2670
rect 6920 -2710 6960 -2705
rect 6920 -2740 6925 -2710
rect 6925 -2740 6955 -2710
rect 6955 -2740 6960 -2710
rect 6920 -2745 6960 -2740
rect 6920 -2780 6960 -2775
rect 6920 -2810 6925 -2780
rect 6925 -2810 6955 -2780
rect 6955 -2810 6960 -2780
rect 6920 -2815 6960 -2810
rect 6920 -2845 6960 -2840
rect 6920 -2875 6925 -2845
rect 6925 -2875 6955 -2845
rect 6955 -2875 6960 -2845
rect 6920 -2880 6960 -2875
rect 7270 -1305 7310 -1300
rect 7270 -1335 7275 -1305
rect 7275 -1335 7305 -1305
rect 7305 -1335 7310 -1305
rect 7270 -1340 7310 -1335
rect 7270 -1370 7310 -1365
rect 7270 -1400 7275 -1370
rect 7275 -1400 7305 -1370
rect 7305 -1400 7310 -1370
rect 7270 -1405 7310 -1400
rect 7270 -1440 7310 -1435
rect 7270 -1470 7275 -1440
rect 7275 -1470 7305 -1440
rect 7305 -1470 7310 -1440
rect 7270 -1475 7310 -1470
rect 7270 -1510 7310 -1505
rect 7270 -1540 7275 -1510
rect 7275 -1540 7305 -1510
rect 7305 -1540 7310 -1510
rect 7270 -1545 7310 -1540
rect 7270 -1580 7310 -1575
rect 7270 -1610 7275 -1580
rect 7275 -1610 7305 -1580
rect 7305 -1610 7310 -1580
rect 7270 -1615 7310 -1610
rect 7270 -1645 7310 -1640
rect 7270 -1675 7275 -1645
rect 7275 -1675 7305 -1645
rect 7305 -1675 7310 -1645
rect 7270 -1680 7310 -1675
rect 7270 -1705 7310 -1700
rect 7270 -1735 7275 -1705
rect 7275 -1735 7305 -1705
rect 7305 -1735 7310 -1705
rect 7270 -1740 7310 -1735
rect 7270 -1770 7310 -1765
rect 7270 -1800 7275 -1770
rect 7275 -1800 7305 -1770
rect 7305 -1800 7310 -1770
rect 7270 -1805 7310 -1800
rect 7270 -1840 7310 -1835
rect 7270 -1870 7275 -1840
rect 7275 -1870 7305 -1840
rect 7305 -1870 7310 -1840
rect 7270 -1875 7310 -1870
rect 7270 -1910 7310 -1905
rect 7270 -1940 7275 -1910
rect 7275 -1940 7305 -1910
rect 7305 -1940 7310 -1910
rect 7270 -1945 7310 -1940
rect 7270 -1980 7310 -1975
rect 7270 -2010 7275 -1980
rect 7275 -2010 7305 -1980
rect 7305 -2010 7310 -1980
rect 7270 -2015 7310 -2010
rect 7270 -2045 7310 -2040
rect 7270 -2075 7275 -2045
rect 7275 -2075 7305 -2045
rect 7305 -2075 7310 -2045
rect 7270 -2080 7310 -2075
rect 7270 -2105 7310 -2100
rect 7270 -2135 7275 -2105
rect 7275 -2135 7305 -2105
rect 7305 -2135 7310 -2105
rect 7270 -2140 7310 -2135
rect 7270 -2170 7310 -2165
rect 7270 -2200 7275 -2170
rect 7275 -2200 7305 -2170
rect 7305 -2200 7310 -2170
rect 7270 -2205 7310 -2200
rect 7270 -2240 7310 -2235
rect 7270 -2270 7275 -2240
rect 7275 -2270 7305 -2240
rect 7305 -2270 7310 -2240
rect 7270 -2275 7310 -2270
rect 7270 -2310 7310 -2305
rect 7270 -2340 7275 -2310
rect 7275 -2340 7305 -2310
rect 7305 -2340 7310 -2310
rect 7270 -2345 7310 -2340
rect 7270 -2380 7310 -2375
rect 7270 -2410 7275 -2380
rect 7275 -2410 7305 -2380
rect 7305 -2410 7310 -2380
rect 7270 -2415 7310 -2410
rect 7270 -2445 7310 -2440
rect 7270 -2475 7275 -2445
rect 7275 -2475 7305 -2445
rect 7305 -2475 7310 -2445
rect 7270 -2480 7310 -2475
rect 7270 -2505 7310 -2500
rect 7270 -2535 7275 -2505
rect 7275 -2535 7305 -2505
rect 7305 -2535 7310 -2505
rect 7270 -2540 7310 -2535
rect 7270 -2570 7310 -2565
rect 7270 -2600 7275 -2570
rect 7275 -2600 7305 -2570
rect 7305 -2600 7310 -2570
rect 7270 -2605 7310 -2600
rect 7270 -2640 7310 -2635
rect 7270 -2670 7275 -2640
rect 7275 -2670 7305 -2640
rect 7305 -2670 7310 -2640
rect 7270 -2675 7310 -2670
rect 7270 -2710 7310 -2705
rect 7270 -2740 7275 -2710
rect 7275 -2740 7305 -2710
rect 7305 -2740 7310 -2710
rect 7270 -2745 7310 -2740
rect 7270 -2780 7310 -2775
rect 7270 -2810 7275 -2780
rect 7275 -2810 7305 -2780
rect 7305 -2810 7310 -2780
rect 7270 -2815 7310 -2810
rect 7270 -2845 7310 -2840
rect 7270 -2875 7275 -2845
rect 7275 -2875 7305 -2845
rect 7305 -2875 7310 -2845
rect 7270 -2880 7310 -2875
rect 7620 -1305 7660 -1300
rect 7620 -1335 7625 -1305
rect 7625 -1335 7655 -1305
rect 7655 -1335 7660 -1305
rect 7620 -1340 7660 -1335
rect 7620 -1370 7660 -1365
rect 7620 -1400 7625 -1370
rect 7625 -1400 7655 -1370
rect 7655 -1400 7660 -1370
rect 7620 -1405 7660 -1400
rect 7620 -1440 7660 -1435
rect 7620 -1470 7625 -1440
rect 7625 -1470 7655 -1440
rect 7655 -1470 7660 -1440
rect 7620 -1475 7660 -1470
rect 7620 -1510 7660 -1505
rect 7620 -1540 7625 -1510
rect 7625 -1540 7655 -1510
rect 7655 -1540 7660 -1510
rect 7620 -1545 7660 -1540
rect 7620 -1580 7660 -1575
rect 7620 -1610 7625 -1580
rect 7625 -1610 7655 -1580
rect 7655 -1610 7660 -1580
rect 7620 -1615 7660 -1610
rect 7620 -1645 7660 -1640
rect 7620 -1675 7625 -1645
rect 7625 -1675 7655 -1645
rect 7655 -1675 7660 -1645
rect 7620 -1680 7660 -1675
rect 7620 -1705 7660 -1700
rect 7620 -1735 7625 -1705
rect 7625 -1735 7655 -1705
rect 7655 -1735 7660 -1705
rect 7620 -1740 7660 -1735
rect 7620 -1770 7660 -1765
rect 7620 -1800 7625 -1770
rect 7625 -1800 7655 -1770
rect 7655 -1800 7660 -1770
rect 7620 -1805 7660 -1800
rect 7620 -1840 7660 -1835
rect 7620 -1870 7625 -1840
rect 7625 -1870 7655 -1840
rect 7655 -1870 7660 -1840
rect 7620 -1875 7660 -1870
rect 7620 -1910 7660 -1905
rect 7620 -1940 7625 -1910
rect 7625 -1940 7655 -1910
rect 7655 -1940 7660 -1910
rect 7620 -1945 7660 -1940
rect 7620 -1980 7660 -1975
rect 7620 -2010 7625 -1980
rect 7625 -2010 7655 -1980
rect 7655 -2010 7660 -1980
rect 7620 -2015 7660 -2010
rect 7620 -2045 7660 -2040
rect 7620 -2075 7625 -2045
rect 7625 -2075 7655 -2045
rect 7655 -2075 7660 -2045
rect 7620 -2080 7660 -2075
rect 7620 -2105 7660 -2100
rect 7620 -2135 7625 -2105
rect 7625 -2135 7655 -2105
rect 7655 -2135 7660 -2105
rect 7620 -2140 7660 -2135
rect 7620 -2170 7660 -2165
rect 7620 -2200 7625 -2170
rect 7625 -2200 7655 -2170
rect 7655 -2200 7660 -2170
rect 7620 -2205 7660 -2200
rect 7620 -2240 7660 -2235
rect 7620 -2270 7625 -2240
rect 7625 -2270 7655 -2240
rect 7655 -2270 7660 -2240
rect 7620 -2275 7660 -2270
rect 7620 -2310 7660 -2305
rect 7620 -2340 7625 -2310
rect 7625 -2340 7655 -2310
rect 7655 -2340 7660 -2310
rect 7620 -2345 7660 -2340
rect 7620 -2380 7660 -2375
rect 7620 -2410 7625 -2380
rect 7625 -2410 7655 -2380
rect 7655 -2410 7660 -2380
rect 7620 -2415 7660 -2410
rect 7620 -2445 7660 -2440
rect 7620 -2475 7625 -2445
rect 7625 -2475 7655 -2445
rect 7655 -2475 7660 -2445
rect 7620 -2480 7660 -2475
rect 7620 -2505 7660 -2500
rect 7620 -2535 7625 -2505
rect 7625 -2535 7655 -2505
rect 7655 -2535 7660 -2505
rect 7620 -2540 7660 -2535
rect 7620 -2570 7660 -2565
rect 7620 -2600 7625 -2570
rect 7625 -2600 7655 -2570
rect 7655 -2600 7660 -2570
rect 7620 -2605 7660 -2600
rect 7620 -2640 7660 -2635
rect 7620 -2670 7625 -2640
rect 7625 -2670 7655 -2640
rect 7655 -2670 7660 -2640
rect 7620 -2675 7660 -2670
rect 7620 -2710 7660 -2705
rect 7620 -2740 7625 -2710
rect 7625 -2740 7655 -2710
rect 7655 -2740 7660 -2710
rect 7620 -2745 7660 -2740
rect 7620 -2780 7660 -2775
rect 7620 -2810 7625 -2780
rect 7625 -2810 7655 -2780
rect 7655 -2810 7660 -2780
rect 7620 -2815 7660 -2810
rect 7620 -2845 7660 -2840
rect 7620 -2875 7625 -2845
rect 7625 -2875 7655 -2845
rect 7655 -2875 7660 -2845
rect 7620 -2880 7660 -2875
rect 7970 -1305 8010 -1300
rect 7970 -1335 7975 -1305
rect 7975 -1335 8005 -1305
rect 8005 -1335 8010 -1305
rect 7970 -1340 8010 -1335
rect 7970 -1370 8010 -1365
rect 7970 -1400 7975 -1370
rect 7975 -1400 8005 -1370
rect 8005 -1400 8010 -1370
rect 7970 -1405 8010 -1400
rect 7970 -1440 8010 -1435
rect 7970 -1470 7975 -1440
rect 7975 -1470 8005 -1440
rect 8005 -1470 8010 -1440
rect 7970 -1475 8010 -1470
rect 7970 -1510 8010 -1505
rect 7970 -1540 7975 -1510
rect 7975 -1540 8005 -1510
rect 8005 -1540 8010 -1510
rect 7970 -1545 8010 -1540
rect 7970 -1580 8010 -1575
rect 7970 -1610 7975 -1580
rect 7975 -1610 8005 -1580
rect 8005 -1610 8010 -1580
rect 7970 -1615 8010 -1610
rect 7970 -1645 8010 -1640
rect 7970 -1675 7975 -1645
rect 7975 -1675 8005 -1645
rect 8005 -1675 8010 -1645
rect 7970 -1680 8010 -1675
rect 7970 -1705 8010 -1700
rect 7970 -1735 7975 -1705
rect 7975 -1735 8005 -1705
rect 8005 -1735 8010 -1705
rect 7970 -1740 8010 -1735
rect 7970 -1770 8010 -1765
rect 7970 -1800 7975 -1770
rect 7975 -1800 8005 -1770
rect 8005 -1800 8010 -1770
rect 7970 -1805 8010 -1800
rect 7970 -1840 8010 -1835
rect 7970 -1870 7975 -1840
rect 7975 -1870 8005 -1840
rect 8005 -1870 8010 -1840
rect 7970 -1875 8010 -1870
rect 7970 -1910 8010 -1905
rect 7970 -1940 7975 -1910
rect 7975 -1940 8005 -1910
rect 8005 -1940 8010 -1910
rect 7970 -1945 8010 -1940
rect 7970 -1980 8010 -1975
rect 7970 -2010 7975 -1980
rect 7975 -2010 8005 -1980
rect 8005 -2010 8010 -1980
rect 7970 -2015 8010 -2010
rect 7970 -2045 8010 -2040
rect 7970 -2075 7975 -2045
rect 7975 -2075 8005 -2045
rect 8005 -2075 8010 -2045
rect 7970 -2080 8010 -2075
rect 7970 -2105 8010 -2100
rect 7970 -2135 7975 -2105
rect 7975 -2135 8005 -2105
rect 8005 -2135 8010 -2105
rect 7970 -2140 8010 -2135
rect 7970 -2170 8010 -2165
rect 7970 -2200 7975 -2170
rect 7975 -2200 8005 -2170
rect 8005 -2200 8010 -2170
rect 7970 -2205 8010 -2200
rect 7970 -2240 8010 -2235
rect 7970 -2270 7975 -2240
rect 7975 -2270 8005 -2240
rect 8005 -2270 8010 -2240
rect 7970 -2275 8010 -2270
rect 7970 -2310 8010 -2305
rect 7970 -2340 7975 -2310
rect 7975 -2340 8005 -2310
rect 8005 -2340 8010 -2310
rect 7970 -2345 8010 -2340
rect 7970 -2380 8010 -2375
rect 7970 -2410 7975 -2380
rect 7975 -2410 8005 -2380
rect 8005 -2410 8010 -2380
rect 7970 -2415 8010 -2410
rect 7970 -2445 8010 -2440
rect 7970 -2475 7975 -2445
rect 7975 -2475 8005 -2445
rect 8005 -2475 8010 -2445
rect 7970 -2480 8010 -2475
rect 7970 -2505 8010 -2500
rect 7970 -2535 7975 -2505
rect 7975 -2535 8005 -2505
rect 8005 -2535 8010 -2505
rect 7970 -2540 8010 -2535
rect 7970 -2570 8010 -2565
rect 7970 -2600 7975 -2570
rect 7975 -2600 8005 -2570
rect 8005 -2600 8010 -2570
rect 7970 -2605 8010 -2600
rect 7970 -2640 8010 -2635
rect 7970 -2670 7975 -2640
rect 7975 -2670 8005 -2640
rect 8005 -2670 8010 -2640
rect 7970 -2675 8010 -2670
rect 7970 -2710 8010 -2705
rect 7970 -2740 7975 -2710
rect 7975 -2740 8005 -2710
rect 8005 -2740 8010 -2710
rect 7970 -2745 8010 -2740
rect 7970 -2780 8010 -2775
rect 7970 -2810 7975 -2780
rect 7975 -2810 8005 -2780
rect 8005 -2810 8010 -2780
rect 7970 -2815 8010 -2810
rect 7970 -2845 8010 -2840
rect 7970 -2875 7975 -2845
rect 7975 -2875 8005 -2845
rect 8005 -2875 8010 -2845
rect 7970 -2880 8010 -2875
rect 8320 -1305 8360 -1300
rect 8320 -1335 8325 -1305
rect 8325 -1335 8355 -1305
rect 8355 -1335 8360 -1305
rect 8320 -1340 8360 -1335
rect 8320 -1370 8360 -1365
rect 8320 -1400 8325 -1370
rect 8325 -1400 8355 -1370
rect 8355 -1400 8360 -1370
rect 8320 -1405 8360 -1400
rect 8320 -1440 8360 -1435
rect 8320 -1470 8325 -1440
rect 8325 -1470 8355 -1440
rect 8355 -1470 8360 -1440
rect 8320 -1475 8360 -1470
rect 8320 -1510 8360 -1505
rect 8320 -1540 8325 -1510
rect 8325 -1540 8355 -1510
rect 8355 -1540 8360 -1510
rect 8320 -1545 8360 -1540
rect 8320 -1580 8360 -1575
rect 8320 -1610 8325 -1580
rect 8325 -1610 8355 -1580
rect 8355 -1610 8360 -1580
rect 8320 -1615 8360 -1610
rect 8320 -1645 8360 -1640
rect 8320 -1675 8325 -1645
rect 8325 -1675 8355 -1645
rect 8355 -1675 8360 -1645
rect 8320 -1680 8360 -1675
rect 8320 -1705 8360 -1700
rect 8320 -1735 8325 -1705
rect 8325 -1735 8355 -1705
rect 8355 -1735 8360 -1705
rect 8320 -1740 8360 -1735
rect 8320 -1770 8360 -1765
rect 8320 -1800 8325 -1770
rect 8325 -1800 8355 -1770
rect 8355 -1800 8360 -1770
rect 8320 -1805 8360 -1800
rect 8320 -1840 8360 -1835
rect 8320 -1870 8325 -1840
rect 8325 -1870 8355 -1840
rect 8355 -1870 8360 -1840
rect 8320 -1875 8360 -1870
rect 8320 -1910 8360 -1905
rect 8320 -1940 8325 -1910
rect 8325 -1940 8355 -1910
rect 8355 -1940 8360 -1910
rect 8320 -1945 8360 -1940
rect 8320 -1980 8360 -1975
rect 8320 -2010 8325 -1980
rect 8325 -2010 8355 -1980
rect 8355 -2010 8360 -1980
rect 8320 -2015 8360 -2010
rect 8320 -2045 8360 -2040
rect 8320 -2075 8325 -2045
rect 8325 -2075 8355 -2045
rect 8355 -2075 8360 -2045
rect 8320 -2080 8360 -2075
rect 8320 -2105 8360 -2100
rect 8320 -2135 8325 -2105
rect 8325 -2135 8355 -2105
rect 8355 -2135 8360 -2105
rect 8320 -2140 8360 -2135
rect 8320 -2170 8360 -2165
rect 8320 -2200 8325 -2170
rect 8325 -2200 8355 -2170
rect 8355 -2200 8360 -2170
rect 8320 -2205 8360 -2200
rect 8320 -2240 8360 -2235
rect 8320 -2270 8325 -2240
rect 8325 -2270 8355 -2240
rect 8355 -2270 8360 -2240
rect 8320 -2275 8360 -2270
rect 8320 -2310 8360 -2305
rect 8320 -2340 8325 -2310
rect 8325 -2340 8355 -2310
rect 8355 -2340 8360 -2310
rect 8320 -2345 8360 -2340
rect 8320 -2380 8360 -2375
rect 8320 -2410 8325 -2380
rect 8325 -2410 8355 -2380
rect 8355 -2410 8360 -2380
rect 8320 -2415 8360 -2410
rect 8320 -2445 8360 -2440
rect 8320 -2475 8325 -2445
rect 8325 -2475 8355 -2445
rect 8355 -2475 8360 -2445
rect 8320 -2480 8360 -2475
rect 8320 -2505 8360 -2500
rect 8320 -2535 8325 -2505
rect 8325 -2535 8355 -2505
rect 8355 -2535 8360 -2505
rect 8320 -2540 8360 -2535
rect 8320 -2570 8360 -2565
rect 8320 -2600 8325 -2570
rect 8325 -2600 8355 -2570
rect 8355 -2600 8360 -2570
rect 8320 -2605 8360 -2600
rect 8320 -2640 8360 -2635
rect 8320 -2670 8325 -2640
rect 8325 -2670 8355 -2640
rect 8355 -2670 8360 -2640
rect 8320 -2675 8360 -2670
rect 8320 -2710 8360 -2705
rect 8320 -2740 8325 -2710
rect 8325 -2740 8355 -2710
rect 8355 -2740 8360 -2710
rect 8320 -2745 8360 -2740
rect 8320 -2780 8360 -2775
rect 8320 -2810 8325 -2780
rect 8325 -2810 8355 -2780
rect 8355 -2810 8360 -2780
rect 8320 -2815 8360 -2810
rect 8320 -2845 8360 -2840
rect 8320 -2875 8325 -2845
rect 8325 -2875 8355 -2845
rect 8355 -2875 8360 -2845
rect 8320 -2880 8360 -2875
rect 31305 -1345 31340 -1310
rect 31350 -1345 31385 -1310
rect 31395 -1345 31430 -1310
rect 31440 -1345 31475 -1310
rect 31485 -1345 31520 -1310
rect 31530 -1345 31565 -1310
rect 31575 -1345 31610 -1310
rect 31620 -1345 31655 -1310
rect 31665 -1345 31700 -1310
rect 31710 -1345 31745 -1310
rect 31755 -1345 31790 -1310
rect 31800 -1345 31835 -1310
rect 31845 -1345 31880 -1310
rect 31890 -1345 31925 -1310
rect 31935 -1345 31970 -1310
rect 31980 -1345 32015 -1310
rect 32025 -1345 32060 -1310
rect 32070 -1345 32105 -1310
rect 32115 -1345 32150 -1310
rect 32160 -1345 32195 -1310
rect 32205 -1345 32240 -1310
rect 32250 -1345 32285 -1310
rect 32295 -1345 32330 -1310
rect 32340 -1345 32375 -1310
rect 32385 -1345 32420 -1310
rect 32430 -1345 32465 -1310
rect 32475 -1345 32510 -1310
rect 32520 -1345 32555 -1310
rect 32565 -1345 32600 -1310
rect 32610 -1345 32645 -1310
rect 32655 -1345 32690 -1310
rect 32700 -1345 32735 -1310
rect 32745 -1345 32780 -1310
rect 32790 -1345 32825 -1310
rect 32835 -1345 32870 -1310
rect 31305 -1390 31340 -1355
rect 31350 -1390 31385 -1355
rect 31395 -1390 31430 -1355
rect 31440 -1390 31475 -1355
rect 31485 -1390 31520 -1355
rect 31530 -1390 31565 -1355
rect 31575 -1390 31610 -1355
rect 31620 -1390 31655 -1355
rect 31665 -1390 31700 -1355
rect 31710 -1390 31745 -1355
rect 31755 -1390 31790 -1355
rect 31800 -1390 31835 -1355
rect 31845 -1390 31880 -1355
rect 31890 -1390 31925 -1355
rect 31935 -1390 31970 -1355
rect 31980 -1390 32015 -1355
rect 32025 -1390 32060 -1355
rect 32070 -1390 32105 -1355
rect 32115 -1390 32150 -1355
rect 32160 -1390 32195 -1355
rect 32205 -1390 32240 -1355
rect 32250 -1390 32285 -1355
rect 32295 -1390 32330 -1355
rect 32340 -1390 32375 -1355
rect 32385 -1390 32420 -1355
rect 32430 -1390 32465 -1355
rect 32475 -1390 32510 -1355
rect 32520 -1390 32555 -1355
rect 32565 -1390 32600 -1355
rect 32610 -1390 32645 -1355
rect 32655 -1390 32690 -1355
rect 32700 -1390 32735 -1355
rect 32745 -1390 32780 -1355
rect 32790 -1390 32825 -1355
rect 32835 -1390 32870 -1355
rect 31305 -1435 31340 -1400
rect 31350 -1435 31385 -1400
rect 31395 -1435 31430 -1400
rect 31440 -1435 31475 -1400
rect 31485 -1435 31520 -1400
rect 31530 -1435 31565 -1400
rect 31575 -1435 31610 -1400
rect 31620 -1435 31655 -1400
rect 31665 -1435 31700 -1400
rect 31710 -1435 31745 -1400
rect 31755 -1435 31790 -1400
rect 31800 -1435 31835 -1400
rect 31845 -1435 31880 -1400
rect 31890 -1435 31925 -1400
rect 31935 -1435 31970 -1400
rect 31980 -1435 32015 -1400
rect 32025 -1435 32060 -1400
rect 32070 -1435 32105 -1400
rect 32115 -1435 32150 -1400
rect 32160 -1435 32195 -1400
rect 32205 -1435 32240 -1400
rect 32250 -1435 32285 -1400
rect 32295 -1435 32330 -1400
rect 32340 -1435 32375 -1400
rect 32385 -1435 32420 -1400
rect 32430 -1435 32465 -1400
rect 32475 -1435 32510 -1400
rect 32520 -1435 32555 -1400
rect 32565 -1435 32600 -1400
rect 32610 -1435 32645 -1400
rect 32655 -1435 32690 -1400
rect 32700 -1435 32735 -1400
rect 32745 -1435 32780 -1400
rect 32790 -1435 32825 -1400
rect 32835 -1435 32870 -1400
rect 31305 -1480 31340 -1445
rect 31350 -1480 31385 -1445
rect 31395 -1480 31430 -1445
rect 31440 -1480 31475 -1445
rect 31485 -1480 31520 -1445
rect 31530 -1480 31565 -1445
rect 31575 -1480 31610 -1445
rect 31620 -1480 31655 -1445
rect 31665 -1480 31700 -1445
rect 31710 -1480 31745 -1445
rect 31755 -1480 31790 -1445
rect 31800 -1480 31835 -1445
rect 31845 -1480 31880 -1445
rect 31890 -1480 31925 -1445
rect 31935 -1480 31970 -1445
rect 31980 -1480 32015 -1445
rect 32025 -1480 32060 -1445
rect 32070 -1480 32105 -1445
rect 32115 -1480 32150 -1445
rect 32160 -1480 32195 -1445
rect 32205 -1480 32240 -1445
rect 32250 -1480 32285 -1445
rect 32295 -1480 32330 -1445
rect 32340 -1480 32375 -1445
rect 32385 -1480 32420 -1445
rect 32430 -1480 32465 -1445
rect 32475 -1480 32510 -1445
rect 32520 -1480 32555 -1445
rect 32565 -1480 32600 -1445
rect 32610 -1480 32645 -1445
rect 32655 -1480 32690 -1445
rect 32700 -1480 32735 -1445
rect 32745 -1480 32780 -1445
rect 32790 -1480 32825 -1445
rect 32835 -1480 32870 -1445
rect 31305 -1525 31340 -1490
rect 31350 -1525 31385 -1490
rect 31395 -1525 31430 -1490
rect 31440 -1525 31475 -1490
rect 31485 -1525 31520 -1490
rect 31530 -1525 31565 -1490
rect 31575 -1525 31610 -1490
rect 31620 -1525 31655 -1490
rect 31665 -1525 31700 -1490
rect 31710 -1525 31745 -1490
rect 31755 -1525 31790 -1490
rect 31800 -1525 31835 -1490
rect 31845 -1525 31880 -1490
rect 31890 -1525 31925 -1490
rect 31935 -1525 31970 -1490
rect 31980 -1525 32015 -1490
rect 32025 -1525 32060 -1490
rect 32070 -1525 32105 -1490
rect 32115 -1525 32150 -1490
rect 32160 -1525 32195 -1490
rect 32205 -1525 32240 -1490
rect 32250 -1525 32285 -1490
rect 32295 -1525 32330 -1490
rect 32340 -1525 32375 -1490
rect 32385 -1525 32420 -1490
rect 32430 -1525 32465 -1490
rect 32475 -1525 32510 -1490
rect 32520 -1525 32555 -1490
rect 32565 -1525 32600 -1490
rect 32610 -1525 32645 -1490
rect 32655 -1525 32690 -1490
rect 32700 -1525 32735 -1490
rect 32745 -1525 32780 -1490
rect 32790 -1525 32825 -1490
rect 32835 -1525 32870 -1490
rect 31305 -1570 31340 -1535
rect 31350 -1570 31385 -1535
rect 31395 -1570 31430 -1535
rect 31440 -1570 31475 -1535
rect 31485 -1570 31520 -1535
rect 31530 -1570 31565 -1535
rect 31575 -1570 31610 -1535
rect 31620 -1570 31655 -1535
rect 31665 -1570 31700 -1535
rect 31710 -1570 31745 -1535
rect 31755 -1570 31790 -1535
rect 31800 -1570 31835 -1535
rect 31845 -1570 31880 -1535
rect 31890 -1570 31925 -1535
rect 31935 -1570 31970 -1535
rect 31980 -1570 32015 -1535
rect 32025 -1570 32060 -1535
rect 32070 -1570 32105 -1535
rect 32115 -1570 32150 -1535
rect 32160 -1570 32195 -1535
rect 32205 -1570 32240 -1535
rect 32250 -1570 32285 -1535
rect 32295 -1570 32330 -1535
rect 32340 -1570 32375 -1535
rect 32385 -1570 32420 -1535
rect 32430 -1570 32465 -1535
rect 32475 -1570 32510 -1535
rect 32520 -1570 32555 -1535
rect 32565 -1570 32600 -1535
rect 32610 -1570 32645 -1535
rect 32655 -1570 32690 -1535
rect 32700 -1570 32735 -1535
rect 32745 -1570 32780 -1535
rect 32790 -1570 32825 -1535
rect 32835 -1570 32870 -1535
rect 31305 -1615 31340 -1580
rect 31350 -1615 31385 -1580
rect 31395 -1615 31430 -1580
rect 31440 -1615 31475 -1580
rect 31485 -1615 31520 -1580
rect 31530 -1615 31565 -1580
rect 31575 -1615 31610 -1580
rect 31620 -1615 31655 -1580
rect 31665 -1615 31700 -1580
rect 31710 -1615 31745 -1580
rect 31755 -1615 31790 -1580
rect 31800 -1615 31835 -1580
rect 31845 -1615 31880 -1580
rect 31890 -1615 31925 -1580
rect 31935 -1615 31970 -1580
rect 31980 -1615 32015 -1580
rect 32025 -1615 32060 -1580
rect 32070 -1615 32105 -1580
rect 32115 -1615 32150 -1580
rect 32160 -1615 32195 -1580
rect 32205 -1615 32240 -1580
rect 32250 -1615 32285 -1580
rect 32295 -1615 32330 -1580
rect 32340 -1615 32375 -1580
rect 32385 -1615 32420 -1580
rect 32430 -1615 32465 -1580
rect 32475 -1615 32510 -1580
rect 32520 -1615 32555 -1580
rect 32565 -1615 32600 -1580
rect 32610 -1615 32645 -1580
rect 32655 -1615 32690 -1580
rect 32700 -1615 32735 -1580
rect 32745 -1615 32780 -1580
rect 32790 -1615 32825 -1580
rect 32835 -1615 32870 -1580
rect 31305 -1660 31340 -1625
rect 31350 -1660 31385 -1625
rect 31395 -1660 31430 -1625
rect 31440 -1660 31475 -1625
rect 31485 -1660 31520 -1625
rect 31530 -1660 31565 -1625
rect 31575 -1660 31610 -1625
rect 31620 -1660 31655 -1625
rect 31665 -1660 31700 -1625
rect 31710 -1660 31745 -1625
rect 31755 -1660 31790 -1625
rect 31800 -1660 31835 -1625
rect 31845 -1660 31880 -1625
rect 31890 -1660 31925 -1625
rect 31935 -1660 31970 -1625
rect 31980 -1660 32015 -1625
rect 32025 -1660 32060 -1625
rect 32070 -1660 32105 -1625
rect 32115 -1660 32150 -1625
rect 32160 -1660 32195 -1625
rect 32205 -1660 32240 -1625
rect 32250 -1660 32285 -1625
rect 32295 -1660 32330 -1625
rect 32340 -1660 32375 -1625
rect 32385 -1660 32420 -1625
rect 32430 -1660 32465 -1625
rect 32475 -1660 32510 -1625
rect 32520 -1660 32555 -1625
rect 32565 -1660 32600 -1625
rect 32610 -1660 32645 -1625
rect 32655 -1660 32690 -1625
rect 32700 -1660 32735 -1625
rect 32745 -1660 32780 -1625
rect 32790 -1660 32825 -1625
rect 32835 -1660 32870 -1625
rect 31305 -1705 31340 -1670
rect 31350 -1705 31385 -1670
rect 31395 -1705 31430 -1670
rect 31440 -1705 31475 -1670
rect 31485 -1705 31520 -1670
rect 31530 -1705 31565 -1670
rect 31575 -1705 31610 -1670
rect 31620 -1705 31655 -1670
rect 31665 -1705 31700 -1670
rect 31710 -1705 31745 -1670
rect 31755 -1705 31790 -1670
rect 31800 -1705 31835 -1670
rect 31845 -1705 31880 -1670
rect 31890 -1705 31925 -1670
rect 31935 -1705 31970 -1670
rect 31980 -1705 32015 -1670
rect 32025 -1705 32060 -1670
rect 32070 -1705 32105 -1670
rect 32115 -1705 32150 -1670
rect 32160 -1705 32195 -1670
rect 32205 -1705 32240 -1670
rect 32250 -1705 32285 -1670
rect 32295 -1705 32330 -1670
rect 32340 -1705 32375 -1670
rect 32385 -1705 32420 -1670
rect 32430 -1705 32465 -1670
rect 32475 -1705 32510 -1670
rect 32520 -1705 32555 -1670
rect 32565 -1705 32600 -1670
rect 32610 -1705 32645 -1670
rect 32655 -1705 32690 -1670
rect 32700 -1705 32735 -1670
rect 32745 -1705 32780 -1670
rect 32790 -1705 32825 -1670
rect 32835 -1705 32870 -1670
rect 31305 -1750 31340 -1715
rect 31350 -1750 31385 -1715
rect 31395 -1750 31430 -1715
rect 31440 -1750 31475 -1715
rect 31485 -1750 31520 -1715
rect 31530 -1750 31565 -1715
rect 31575 -1750 31610 -1715
rect 31620 -1750 31655 -1715
rect 31665 -1750 31700 -1715
rect 31710 -1750 31745 -1715
rect 31755 -1750 31790 -1715
rect 31800 -1750 31835 -1715
rect 31845 -1750 31880 -1715
rect 31890 -1750 31925 -1715
rect 31935 -1750 31970 -1715
rect 31980 -1750 32015 -1715
rect 32025 -1750 32060 -1715
rect 32070 -1750 32105 -1715
rect 32115 -1750 32150 -1715
rect 32160 -1750 32195 -1715
rect 32205 -1750 32240 -1715
rect 32250 -1750 32285 -1715
rect 32295 -1750 32330 -1715
rect 32340 -1750 32375 -1715
rect 32385 -1750 32420 -1715
rect 32430 -1750 32465 -1715
rect 32475 -1750 32510 -1715
rect 32520 -1750 32555 -1715
rect 32565 -1750 32600 -1715
rect 32610 -1750 32645 -1715
rect 32655 -1750 32690 -1715
rect 32700 -1750 32735 -1715
rect 32745 -1750 32780 -1715
rect 32790 -1750 32825 -1715
rect 32835 -1750 32870 -1715
rect 31305 -1795 31340 -1760
rect 31350 -1795 31385 -1760
rect 31395 -1795 31430 -1760
rect 31440 -1795 31475 -1760
rect 31485 -1795 31520 -1760
rect 31530 -1795 31565 -1760
rect 31575 -1795 31610 -1760
rect 31620 -1795 31655 -1760
rect 31665 -1795 31700 -1760
rect 31710 -1795 31745 -1760
rect 31755 -1795 31790 -1760
rect 31800 -1795 31835 -1760
rect 31845 -1795 31880 -1760
rect 31890 -1795 31925 -1760
rect 31935 -1795 31970 -1760
rect 31980 -1795 32015 -1760
rect 32025 -1795 32060 -1760
rect 32070 -1795 32105 -1760
rect 32115 -1795 32150 -1760
rect 32160 -1795 32195 -1760
rect 32205 -1795 32240 -1760
rect 32250 -1795 32285 -1760
rect 32295 -1795 32330 -1760
rect 32340 -1795 32375 -1760
rect 32385 -1795 32420 -1760
rect 32430 -1795 32465 -1760
rect 32475 -1795 32510 -1760
rect 32520 -1795 32555 -1760
rect 32565 -1795 32600 -1760
rect 32610 -1795 32645 -1760
rect 32655 -1795 32690 -1760
rect 32700 -1795 32735 -1760
rect 32745 -1795 32780 -1760
rect 32790 -1795 32825 -1760
rect 32835 -1795 32870 -1760
rect 31305 -1840 31340 -1805
rect 31350 -1840 31385 -1805
rect 31395 -1840 31430 -1805
rect 31440 -1840 31475 -1805
rect 31485 -1840 31520 -1805
rect 31530 -1840 31565 -1805
rect 31575 -1840 31610 -1805
rect 31620 -1840 31655 -1805
rect 31665 -1840 31700 -1805
rect 31710 -1840 31745 -1805
rect 31755 -1840 31790 -1805
rect 31800 -1840 31835 -1805
rect 31845 -1840 31880 -1805
rect 31890 -1840 31925 -1805
rect 31935 -1840 31970 -1805
rect 31980 -1840 32015 -1805
rect 32025 -1840 32060 -1805
rect 32070 -1840 32105 -1805
rect 32115 -1840 32150 -1805
rect 32160 -1840 32195 -1805
rect 32205 -1840 32240 -1805
rect 32250 -1840 32285 -1805
rect 32295 -1840 32330 -1805
rect 32340 -1840 32375 -1805
rect 32385 -1840 32420 -1805
rect 32430 -1840 32465 -1805
rect 32475 -1840 32510 -1805
rect 32520 -1840 32555 -1805
rect 32565 -1840 32600 -1805
rect 32610 -1840 32645 -1805
rect 32655 -1840 32690 -1805
rect 32700 -1840 32735 -1805
rect 32745 -1840 32780 -1805
rect 32790 -1840 32825 -1805
rect 32835 -1840 32870 -1805
rect 31305 -1885 31340 -1850
rect 31350 -1885 31385 -1850
rect 31395 -1885 31430 -1850
rect 31440 -1885 31475 -1850
rect 31485 -1885 31520 -1850
rect 31530 -1885 31565 -1850
rect 31575 -1885 31610 -1850
rect 31620 -1885 31655 -1850
rect 31665 -1885 31700 -1850
rect 31710 -1885 31745 -1850
rect 31755 -1885 31790 -1850
rect 31800 -1885 31835 -1850
rect 31845 -1885 31880 -1850
rect 31890 -1885 31925 -1850
rect 31935 -1885 31970 -1850
rect 31980 -1885 32015 -1850
rect 32025 -1885 32060 -1850
rect 32070 -1885 32105 -1850
rect 32115 -1885 32150 -1850
rect 32160 -1885 32195 -1850
rect 32205 -1885 32240 -1850
rect 32250 -1885 32285 -1850
rect 32295 -1885 32330 -1850
rect 32340 -1885 32375 -1850
rect 32385 -1885 32420 -1850
rect 32430 -1885 32465 -1850
rect 32475 -1885 32510 -1850
rect 32520 -1885 32555 -1850
rect 32565 -1885 32600 -1850
rect 32610 -1885 32645 -1850
rect 32655 -1885 32690 -1850
rect 32700 -1885 32735 -1850
rect 32745 -1885 32780 -1850
rect 32790 -1885 32825 -1850
rect 32835 -1885 32870 -1850
rect 31305 -1930 31340 -1895
rect 31350 -1930 31385 -1895
rect 31395 -1930 31430 -1895
rect 31440 -1930 31475 -1895
rect 31485 -1930 31520 -1895
rect 31530 -1930 31565 -1895
rect 31575 -1930 31610 -1895
rect 31620 -1930 31655 -1895
rect 31665 -1930 31700 -1895
rect 31710 -1930 31745 -1895
rect 31755 -1930 31790 -1895
rect 31800 -1930 31835 -1895
rect 31845 -1930 31880 -1895
rect 31890 -1930 31925 -1895
rect 31935 -1930 31970 -1895
rect 31980 -1930 32015 -1895
rect 32025 -1930 32060 -1895
rect 32070 -1930 32105 -1895
rect 32115 -1930 32150 -1895
rect 32160 -1930 32195 -1895
rect 32205 -1930 32240 -1895
rect 32250 -1930 32285 -1895
rect 32295 -1930 32330 -1895
rect 32340 -1930 32375 -1895
rect 32385 -1930 32420 -1895
rect 32430 -1930 32465 -1895
rect 32475 -1930 32510 -1895
rect 32520 -1930 32555 -1895
rect 32565 -1930 32600 -1895
rect 32610 -1930 32645 -1895
rect 32655 -1930 32690 -1895
rect 32700 -1930 32735 -1895
rect 32745 -1930 32780 -1895
rect 32790 -1930 32825 -1895
rect 32835 -1930 32870 -1895
rect 31305 -1975 31340 -1940
rect 31350 -1975 31385 -1940
rect 31395 -1975 31430 -1940
rect 31440 -1975 31475 -1940
rect 31485 -1975 31520 -1940
rect 31530 -1975 31565 -1940
rect 31575 -1975 31610 -1940
rect 31620 -1975 31655 -1940
rect 31665 -1975 31700 -1940
rect 31710 -1975 31745 -1940
rect 31755 -1975 31790 -1940
rect 31800 -1975 31835 -1940
rect 31845 -1975 31880 -1940
rect 31890 -1975 31925 -1940
rect 31935 -1975 31970 -1940
rect 31980 -1975 32015 -1940
rect 32025 -1975 32060 -1940
rect 32070 -1975 32105 -1940
rect 32115 -1975 32150 -1940
rect 32160 -1975 32195 -1940
rect 32205 -1975 32240 -1940
rect 32250 -1975 32285 -1940
rect 32295 -1975 32330 -1940
rect 32340 -1975 32375 -1940
rect 32385 -1975 32420 -1940
rect 32430 -1975 32465 -1940
rect 32475 -1975 32510 -1940
rect 32520 -1975 32555 -1940
rect 32565 -1975 32600 -1940
rect 32610 -1975 32645 -1940
rect 32655 -1975 32690 -1940
rect 32700 -1975 32735 -1940
rect 32745 -1975 32780 -1940
rect 32790 -1975 32825 -1940
rect 32835 -1975 32870 -1940
rect 31305 -2020 31340 -1985
rect 31350 -2020 31385 -1985
rect 31395 -2020 31430 -1985
rect 31440 -2020 31475 -1985
rect 31485 -2020 31520 -1985
rect 31530 -2020 31565 -1985
rect 31575 -2020 31610 -1985
rect 31620 -2020 31655 -1985
rect 31665 -2020 31700 -1985
rect 31710 -2020 31745 -1985
rect 31755 -2020 31790 -1985
rect 31800 -2020 31835 -1985
rect 31845 -2020 31880 -1985
rect 31890 -2020 31925 -1985
rect 31935 -2020 31970 -1985
rect 31980 -2020 32015 -1985
rect 32025 -2020 32060 -1985
rect 32070 -2020 32105 -1985
rect 32115 -2020 32150 -1985
rect 32160 -2020 32195 -1985
rect 32205 -2020 32240 -1985
rect 32250 -2020 32285 -1985
rect 32295 -2020 32330 -1985
rect 32340 -2020 32375 -1985
rect 32385 -2020 32420 -1985
rect 32430 -2020 32465 -1985
rect 32475 -2020 32510 -1985
rect 32520 -2020 32555 -1985
rect 32565 -2020 32600 -1985
rect 32610 -2020 32645 -1985
rect 32655 -2020 32690 -1985
rect 32700 -2020 32735 -1985
rect 32745 -2020 32780 -1985
rect 32790 -2020 32825 -1985
rect 32835 -2020 32870 -1985
rect 31305 -2065 31340 -2030
rect 31350 -2065 31385 -2030
rect 31395 -2065 31430 -2030
rect 31440 -2065 31475 -2030
rect 31485 -2065 31520 -2030
rect 31530 -2065 31565 -2030
rect 31575 -2065 31610 -2030
rect 31620 -2065 31655 -2030
rect 31665 -2065 31700 -2030
rect 31710 -2065 31745 -2030
rect 31755 -2065 31790 -2030
rect 31800 -2065 31835 -2030
rect 31845 -2065 31880 -2030
rect 31890 -2065 31925 -2030
rect 31935 -2065 31970 -2030
rect 31980 -2065 32015 -2030
rect 32025 -2065 32060 -2030
rect 32070 -2065 32105 -2030
rect 32115 -2065 32150 -2030
rect 32160 -2065 32195 -2030
rect 32205 -2065 32240 -2030
rect 32250 -2065 32285 -2030
rect 32295 -2065 32330 -2030
rect 32340 -2065 32375 -2030
rect 32385 -2065 32420 -2030
rect 32430 -2065 32465 -2030
rect 32475 -2065 32510 -2030
rect 32520 -2065 32555 -2030
rect 32565 -2065 32600 -2030
rect 32610 -2065 32645 -2030
rect 32655 -2065 32690 -2030
rect 32700 -2065 32735 -2030
rect 32745 -2065 32780 -2030
rect 32790 -2065 32825 -2030
rect 32835 -2065 32870 -2030
rect 31305 -2110 31340 -2075
rect 31350 -2110 31385 -2075
rect 31395 -2110 31430 -2075
rect 31440 -2110 31475 -2075
rect 31485 -2110 31520 -2075
rect 31530 -2110 31565 -2075
rect 31575 -2110 31610 -2075
rect 31620 -2110 31655 -2075
rect 31665 -2110 31700 -2075
rect 31710 -2110 31745 -2075
rect 31755 -2110 31790 -2075
rect 31800 -2110 31835 -2075
rect 31845 -2110 31880 -2075
rect 31890 -2110 31925 -2075
rect 31935 -2110 31970 -2075
rect 31980 -2110 32015 -2075
rect 32025 -2110 32060 -2075
rect 32070 -2110 32105 -2075
rect 32115 -2110 32150 -2075
rect 32160 -2110 32195 -2075
rect 32205 -2110 32240 -2075
rect 32250 -2110 32285 -2075
rect 32295 -2110 32330 -2075
rect 32340 -2110 32375 -2075
rect 32385 -2110 32420 -2075
rect 32430 -2110 32465 -2075
rect 32475 -2110 32510 -2075
rect 32520 -2110 32555 -2075
rect 32565 -2110 32600 -2075
rect 32610 -2110 32645 -2075
rect 32655 -2110 32690 -2075
rect 32700 -2110 32735 -2075
rect 32745 -2110 32780 -2075
rect 32790 -2110 32825 -2075
rect 32835 -2110 32870 -2075
rect 31305 -2155 31340 -2120
rect 31350 -2155 31385 -2120
rect 31395 -2155 31430 -2120
rect 31440 -2155 31475 -2120
rect 31485 -2155 31520 -2120
rect 31530 -2155 31565 -2120
rect 31575 -2155 31610 -2120
rect 31620 -2155 31655 -2120
rect 31665 -2155 31700 -2120
rect 31710 -2155 31745 -2120
rect 31755 -2155 31790 -2120
rect 31800 -2155 31835 -2120
rect 31845 -2155 31880 -2120
rect 31890 -2155 31925 -2120
rect 31935 -2155 31970 -2120
rect 31980 -2155 32015 -2120
rect 32025 -2155 32060 -2120
rect 32070 -2155 32105 -2120
rect 32115 -2155 32150 -2120
rect 32160 -2155 32195 -2120
rect 32205 -2155 32240 -2120
rect 32250 -2155 32285 -2120
rect 32295 -2155 32330 -2120
rect 32340 -2155 32375 -2120
rect 32385 -2155 32420 -2120
rect 32430 -2155 32465 -2120
rect 32475 -2155 32510 -2120
rect 32520 -2155 32555 -2120
rect 32565 -2155 32600 -2120
rect 32610 -2155 32645 -2120
rect 32655 -2155 32690 -2120
rect 32700 -2155 32735 -2120
rect 32745 -2155 32780 -2120
rect 32790 -2155 32825 -2120
rect 32835 -2155 32870 -2120
rect 31305 -2200 31340 -2165
rect 31350 -2200 31385 -2165
rect 31395 -2200 31430 -2165
rect 31440 -2200 31475 -2165
rect 31485 -2200 31520 -2165
rect 31530 -2200 31565 -2165
rect 31575 -2200 31610 -2165
rect 31620 -2200 31655 -2165
rect 31665 -2200 31700 -2165
rect 31710 -2200 31745 -2165
rect 31755 -2200 31790 -2165
rect 31800 -2200 31835 -2165
rect 31845 -2200 31880 -2165
rect 31890 -2200 31925 -2165
rect 31935 -2200 31970 -2165
rect 31980 -2200 32015 -2165
rect 32025 -2200 32060 -2165
rect 32070 -2200 32105 -2165
rect 32115 -2200 32150 -2165
rect 32160 -2200 32195 -2165
rect 32205 -2200 32240 -2165
rect 32250 -2200 32285 -2165
rect 32295 -2200 32330 -2165
rect 32340 -2200 32375 -2165
rect 32385 -2200 32420 -2165
rect 32430 -2200 32465 -2165
rect 32475 -2200 32510 -2165
rect 32520 -2200 32555 -2165
rect 32565 -2200 32600 -2165
rect 32610 -2200 32645 -2165
rect 32655 -2200 32690 -2165
rect 32700 -2200 32735 -2165
rect 32745 -2200 32780 -2165
rect 32790 -2200 32825 -2165
rect 32835 -2200 32870 -2165
rect 31305 -2245 31340 -2210
rect 31350 -2245 31385 -2210
rect 31395 -2245 31430 -2210
rect 31440 -2245 31475 -2210
rect 31485 -2245 31520 -2210
rect 31530 -2245 31565 -2210
rect 31575 -2245 31610 -2210
rect 31620 -2245 31655 -2210
rect 31665 -2245 31700 -2210
rect 31710 -2245 31745 -2210
rect 31755 -2245 31790 -2210
rect 31800 -2245 31835 -2210
rect 31845 -2245 31880 -2210
rect 31890 -2245 31925 -2210
rect 31935 -2245 31970 -2210
rect 31980 -2245 32015 -2210
rect 32025 -2245 32060 -2210
rect 32070 -2245 32105 -2210
rect 32115 -2245 32150 -2210
rect 32160 -2245 32195 -2210
rect 32205 -2245 32240 -2210
rect 32250 -2245 32285 -2210
rect 32295 -2245 32330 -2210
rect 32340 -2245 32375 -2210
rect 32385 -2245 32420 -2210
rect 32430 -2245 32465 -2210
rect 32475 -2245 32510 -2210
rect 32520 -2245 32555 -2210
rect 32565 -2245 32600 -2210
rect 32610 -2245 32645 -2210
rect 32655 -2245 32690 -2210
rect 32700 -2245 32735 -2210
rect 32745 -2245 32780 -2210
rect 32790 -2245 32825 -2210
rect 32835 -2245 32870 -2210
rect 31305 -2290 31340 -2255
rect 31350 -2290 31385 -2255
rect 31395 -2290 31430 -2255
rect 31440 -2290 31475 -2255
rect 31485 -2290 31520 -2255
rect 31530 -2290 31565 -2255
rect 31575 -2290 31610 -2255
rect 31620 -2290 31655 -2255
rect 31665 -2290 31700 -2255
rect 31710 -2290 31745 -2255
rect 31755 -2290 31790 -2255
rect 31800 -2290 31835 -2255
rect 31845 -2290 31880 -2255
rect 31890 -2290 31925 -2255
rect 31935 -2290 31970 -2255
rect 31980 -2290 32015 -2255
rect 32025 -2290 32060 -2255
rect 32070 -2290 32105 -2255
rect 32115 -2290 32150 -2255
rect 32160 -2290 32195 -2255
rect 32205 -2290 32240 -2255
rect 32250 -2290 32285 -2255
rect 32295 -2290 32330 -2255
rect 32340 -2290 32375 -2255
rect 32385 -2290 32420 -2255
rect 32430 -2290 32465 -2255
rect 32475 -2290 32510 -2255
rect 32520 -2290 32555 -2255
rect 32565 -2290 32600 -2255
rect 32610 -2290 32645 -2255
rect 32655 -2290 32690 -2255
rect 32700 -2290 32735 -2255
rect 32745 -2290 32780 -2255
rect 32790 -2290 32825 -2255
rect 32835 -2290 32870 -2255
rect 31305 -2335 31340 -2300
rect 31350 -2335 31385 -2300
rect 31395 -2335 31430 -2300
rect 31440 -2335 31475 -2300
rect 31485 -2335 31520 -2300
rect 31530 -2335 31565 -2300
rect 31575 -2335 31610 -2300
rect 31620 -2335 31655 -2300
rect 31665 -2335 31700 -2300
rect 31710 -2335 31745 -2300
rect 31755 -2335 31790 -2300
rect 31800 -2335 31835 -2300
rect 31845 -2335 31880 -2300
rect 31890 -2335 31925 -2300
rect 31935 -2335 31970 -2300
rect 31980 -2335 32015 -2300
rect 32025 -2335 32060 -2300
rect 32070 -2335 32105 -2300
rect 32115 -2335 32150 -2300
rect 32160 -2335 32195 -2300
rect 32205 -2335 32240 -2300
rect 32250 -2335 32285 -2300
rect 32295 -2335 32330 -2300
rect 32340 -2335 32375 -2300
rect 32385 -2335 32420 -2300
rect 32430 -2335 32465 -2300
rect 32475 -2335 32510 -2300
rect 32520 -2335 32555 -2300
rect 32565 -2335 32600 -2300
rect 32610 -2335 32645 -2300
rect 32655 -2335 32690 -2300
rect 32700 -2335 32735 -2300
rect 32745 -2335 32780 -2300
rect 32790 -2335 32825 -2300
rect 32835 -2335 32870 -2300
rect 31305 -2380 31340 -2345
rect 31350 -2380 31385 -2345
rect 31395 -2380 31430 -2345
rect 31440 -2380 31475 -2345
rect 31485 -2380 31520 -2345
rect 31530 -2380 31565 -2345
rect 31575 -2380 31610 -2345
rect 31620 -2380 31655 -2345
rect 31665 -2380 31700 -2345
rect 31710 -2380 31745 -2345
rect 31755 -2380 31790 -2345
rect 31800 -2380 31835 -2345
rect 31845 -2380 31880 -2345
rect 31890 -2380 31925 -2345
rect 31935 -2380 31970 -2345
rect 31980 -2380 32015 -2345
rect 32025 -2380 32060 -2345
rect 32070 -2380 32105 -2345
rect 32115 -2380 32150 -2345
rect 32160 -2380 32195 -2345
rect 32205 -2380 32240 -2345
rect 32250 -2380 32285 -2345
rect 32295 -2380 32330 -2345
rect 32340 -2380 32375 -2345
rect 32385 -2380 32420 -2345
rect 32430 -2380 32465 -2345
rect 32475 -2380 32510 -2345
rect 32520 -2380 32555 -2345
rect 32565 -2380 32600 -2345
rect 32610 -2380 32645 -2345
rect 32655 -2380 32690 -2345
rect 32700 -2380 32735 -2345
rect 32745 -2380 32780 -2345
rect 32790 -2380 32825 -2345
rect 32835 -2380 32870 -2345
rect 31305 -2425 31340 -2390
rect 31350 -2425 31385 -2390
rect 31395 -2425 31430 -2390
rect 31440 -2425 31475 -2390
rect 31485 -2425 31520 -2390
rect 31530 -2425 31565 -2390
rect 31575 -2425 31610 -2390
rect 31620 -2425 31655 -2390
rect 31665 -2425 31700 -2390
rect 31710 -2425 31745 -2390
rect 31755 -2425 31790 -2390
rect 31800 -2425 31835 -2390
rect 31845 -2425 31880 -2390
rect 31890 -2425 31925 -2390
rect 31935 -2425 31970 -2390
rect 31980 -2425 32015 -2390
rect 32025 -2425 32060 -2390
rect 32070 -2425 32105 -2390
rect 32115 -2425 32150 -2390
rect 32160 -2425 32195 -2390
rect 32205 -2425 32240 -2390
rect 32250 -2425 32285 -2390
rect 32295 -2425 32330 -2390
rect 32340 -2425 32375 -2390
rect 32385 -2425 32420 -2390
rect 32430 -2425 32465 -2390
rect 32475 -2425 32510 -2390
rect 32520 -2425 32555 -2390
rect 32565 -2425 32600 -2390
rect 32610 -2425 32645 -2390
rect 32655 -2425 32690 -2390
rect 32700 -2425 32735 -2390
rect 32745 -2425 32780 -2390
rect 32790 -2425 32825 -2390
rect 32835 -2425 32870 -2390
rect 31305 -2470 31340 -2435
rect 31350 -2470 31385 -2435
rect 31395 -2470 31430 -2435
rect 31440 -2470 31475 -2435
rect 31485 -2470 31520 -2435
rect 31530 -2470 31565 -2435
rect 31575 -2470 31610 -2435
rect 31620 -2470 31655 -2435
rect 31665 -2470 31700 -2435
rect 31710 -2470 31745 -2435
rect 31755 -2470 31790 -2435
rect 31800 -2470 31835 -2435
rect 31845 -2470 31880 -2435
rect 31890 -2470 31925 -2435
rect 31935 -2470 31970 -2435
rect 31980 -2470 32015 -2435
rect 32025 -2470 32060 -2435
rect 32070 -2470 32105 -2435
rect 32115 -2470 32150 -2435
rect 32160 -2470 32195 -2435
rect 32205 -2470 32240 -2435
rect 32250 -2470 32285 -2435
rect 32295 -2470 32330 -2435
rect 32340 -2470 32375 -2435
rect 32385 -2470 32420 -2435
rect 32430 -2470 32465 -2435
rect 32475 -2470 32510 -2435
rect 32520 -2470 32555 -2435
rect 32565 -2470 32600 -2435
rect 32610 -2470 32645 -2435
rect 32655 -2470 32690 -2435
rect 32700 -2470 32735 -2435
rect 32745 -2470 32780 -2435
rect 32790 -2470 32825 -2435
rect 32835 -2470 32870 -2435
rect 31305 -2515 31340 -2480
rect 31350 -2515 31385 -2480
rect 31395 -2515 31430 -2480
rect 31440 -2515 31475 -2480
rect 31485 -2515 31520 -2480
rect 31530 -2515 31565 -2480
rect 31575 -2515 31610 -2480
rect 31620 -2515 31655 -2480
rect 31665 -2515 31700 -2480
rect 31710 -2515 31745 -2480
rect 31755 -2515 31790 -2480
rect 31800 -2515 31835 -2480
rect 31845 -2515 31880 -2480
rect 31890 -2515 31925 -2480
rect 31935 -2515 31970 -2480
rect 31980 -2515 32015 -2480
rect 32025 -2515 32060 -2480
rect 32070 -2515 32105 -2480
rect 32115 -2515 32150 -2480
rect 32160 -2515 32195 -2480
rect 32205 -2515 32240 -2480
rect 32250 -2515 32285 -2480
rect 32295 -2515 32330 -2480
rect 32340 -2515 32375 -2480
rect 32385 -2515 32420 -2480
rect 32430 -2515 32465 -2480
rect 32475 -2515 32510 -2480
rect 32520 -2515 32555 -2480
rect 32565 -2515 32600 -2480
rect 32610 -2515 32645 -2480
rect 32655 -2515 32690 -2480
rect 32700 -2515 32735 -2480
rect 32745 -2515 32780 -2480
rect 32790 -2515 32825 -2480
rect 32835 -2515 32870 -2480
rect 31305 -2560 31340 -2525
rect 31350 -2560 31385 -2525
rect 31395 -2560 31430 -2525
rect 31440 -2560 31475 -2525
rect 31485 -2560 31520 -2525
rect 31530 -2560 31565 -2525
rect 31575 -2560 31610 -2525
rect 31620 -2560 31655 -2525
rect 31665 -2560 31700 -2525
rect 31710 -2560 31745 -2525
rect 31755 -2560 31790 -2525
rect 31800 -2560 31835 -2525
rect 31845 -2560 31880 -2525
rect 31890 -2560 31925 -2525
rect 31935 -2560 31970 -2525
rect 31980 -2560 32015 -2525
rect 32025 -2560 32060 -2525
rect 32070 -2560 32105 -2525
rect 32115 -2560 32150 -2525
rect 32160 -2560 32195 -2525
rect 32205 -2560 32240 -2525
rect 32250 -2560 32285 -2525
rect 32295 -2560 32330 -2525
rect 32340 -2560 32375 -2525
rect 32385 -2560 32420 -2525
rect 32430 -2560 32465 -2525
rect 32475 -2560 32510 -2525
rect 32520 -2560 32555 -2525
rect 32565 -2560 32600 -2525
rect 32610 -2560 32645 -2525
rect 32655 -2560 32690 -2525
rect 32700 -2560 32735 -2525
rect 32745 -2560 32780 -2525
rect 32790 -2560 32825 -2525
rect 32835 -2560 32870 -2525
rect 31305 -2605 31340 -2570
rect 31350 -2605 31385 -2570
rect 31395 -2605 31430 -2570
rect 31440 -2605 31475 -2570
rect 31485 -2605 31520 -2570
rect 31530 -2605 31565 -2570
rect 31575 -2605 31610 -2570
rect 31620 -2605 31655 -2570
rect 31665 -2605 31700 -2570
rect 31710 -2605 31745 -2570
rect 31755 -2605 31790 -2570
rect 31800 -2605 31835 -2570
rect 31845 -2605 31880 -2570
rect 31890 -2605 31925 -2570
rect 31935 -2605 31970 -2570
rect 31980 -2605 32015 -2570
rect 32025 -2605 32060 -2570
rect 32070 -2605 32105 -2570
rect 32115 -2605 32150 -2570
rect 32160 -2605 32195 -2570
rect 32205 -2605 32240 -2570
rect 32250 -2605 32285 -2570
rect 32295 -2605 32330 -2570
rect 32340 -2605 32375 -2570
rect 32385 -2605 32420 -2570
rect 32430 -2605 32465 -2570
rect 32475 -2605 32510 -2570
rect 32520 -2605 32555 -2570
rect 32565 -2605 32600 -2570
rect 32610 -2605 32645 -2570
rect 32655 -2605 32690 -2570
rect 32700 -2605 32735 -2570
rect 32745 -2605 32780 -2570
rect 32790 -2605 32825 -2570
rect 32835 -2605 32870 -2570
rect 31305 -2650 31340 -2615
rect 31350 -2650 31385 -2615
rect 31395 -2650 31430 -2615
rect 31440 -2650 31475 -2615
rect 31485 -2650 31520 -2615
rect 31530 -2650 31565 -2615
rect 31575 -2650 31610 -2615
rect 31620 -2650 31655 -2615
rect 31665 -2650 31700 -2615
rect 31710 -2650 31745 -2615
rect 31755 -2650 31790 -2615
rect 31800 -2650 31835 -2615
rect 31845 -2650 31880 -2615
rect 31890 -2650 31925 -2615
rect 31935 -2650 31970 -2615
rect 31980 -2650 32015 -2615
rect 32025 -2650 32060 -2615
rect 32070 -2650 32105 -2615
rect 32115 -2650 32150 -2615
rect 32160 -2650 32195 -2615
rect 32205 -2650 32240 -2615
rect 32250 -2650 32285 -2615
rect 32295 -2650 32330 -2615
rect 32340 -2650 32375 -2615
rect 32385 -2650 32420 -2615
rect 32430 -2650 32465 -2615
rect 32475 -2650 32510 -2615
rect 32520 -2650 32555 -2615
rect 32565 -2650 32600 -2615
rect 32610 -2650 32645 -2615
rect 32655 -2650 32690 -2615
rect 32700 -2650 32735 -2615
rect 32745 -2650 32780 -2615
rect 32790 -2650 32825 -2615
rect 32835 -2650 32870 -2615
rect 31305 -2695 31340 -2660
rect 31350 -2695 31385 -2660
rect 31395 -2695 31430 -2660
rect 31440 -2695 31475 -2660
rect 31485 -2695 31520 -2660
rect 31530 -2695 31565 -2660
rect 31575 -2695 31610 -2660
rect 31620 -2695 31655 -2660
rect 31665 -2695 31700 -2660
rect 31710 -2695 31745 -2660
rect 31755 -2695 31790 -2660
rect 31800 -2695 31835 -2660
rect 31845 -2695 31880 -2660
rect 31890 -2695 31925 -2660
rect 31935 -2695 31970 -2660
rect 31980 -2695 32015 -2660
rect 32025 -2695 32060 -2660
rect 32070 -2695 32105 -2660
rect 32115 -2695 32150 -2660
rect 32160 -2695 32195 -2660
rect 32205 -2695 32240 -2660
rect 32250 -2695 32285 -2660
rect 32295 -2695 32330 -2660
rect 32340 -2695 32375 -2660
rect 32385 -2695 32420 -2660
rect 32430 -2695 32465 -2660
rect 32475 -2695 32510 -2660
rect 32520 -2695 32555 -2660
rect 32565 -2695 32600 -2660
rect 32610 -2695 32645 -2660
rect 32655 -2695 32690 -2660
rect 32700 -2695 32735 -2660
rect 32745 -2695 32780 -2660
rect 32790 -2695 32825 -2660
rect 32835 -2695 32870 -2660
rect 31305 -2740 31340 -2705
rect 31350 -2740 31385 -2705
rect 31395 -2740 31430 -2705
rect 31440 -2740 31475 -2705
rect 31485 -2740 31520 -2705
rect 31530 -2740 31565 -2705
rect 31575 -2740 31610 -2705
rect 31620 -2740 31655 -2705
rect 31665 -2740 31700 -2705
rect 31710 -2740 31745 -2705
rect 31755 -2740 31790 -2705
rect 31800 -2740 31835 -2705
rect 31845 -2740 31880 -2705
rect 31890 -2740 31925 -2705
rect 31935 -2740 31970 -2705
rect 31980 -2740 32015 -2705
rect 32025 -2740 32060 -2705
rect 32070 -2740 32105 -2705
rect 32115 -2740 32150 -2705
rect 32160 -2740 32195 -2705
rect 32205 -2740 32240 -2705
rect 32250 -2740 32285 -2705
rect 32295 -2740 32330 -2705
rect 32340 -2740 32375 -2705
rect 32385 -2740 32420 -2705
rect 32430 -2740 32465 -2705
rect 32475 -2740 32510 -2705
rect 32520 -2740 32555 -2705
rect 32565 -2740 32600 -2705
rect 32610 -2740 32645 -2705
rect 32655 -2740 32690 -2705
rect 32700 -2740 32735 -2705
rect 32745 -2740 32780 -2705
rect 32790 -2740 32825 -2705
rect 32835 -2740 32870 -2705
rect 31305 -2785 31340 -2750
rect 31350 -2785 31385 -2750
rect 31395 -2785 31430 -2750
rect 31440 -2785 31475 -2750
rect 31485 -2785 31520 -2750
rect 31530 -2785 31565 -2750
rect 31575 -2785 31610 -2750
rect 31620 -2785 31655 -2750
rect 31665 -2785 31700 -2750
rect 31710 -2785 31745 -2750
rect 31755 -2785 31790 -2750
rect 31800 -2785 31835 -2750
rect 31845 -2785 31880 -2750
rect 31890 -2785 31925 -2750
rect 31935 -2785 31970 -2750
rect 31980 -2785 32015 -2750
rect 32025 -2785 32060 -2750
rect 32070 -2785 32105 -2750
rect 32115 -2785 32150 -2750
rect 32160 -2785 32195 -2750
rect 32205 -2785 32240 -2750
rect 32250 -2785 32285 -2750
rect 32295 -2785 32330 -2750
rect 32340 -2785 32375 -2750
rect 32385 -2785 32420 -2750
rect 32430 -2785 32465 -2750
rect 32475 -2785 32510 -2750
rect 32520 -2785 32555 -2750
rect 32565 -2785 32600 -2750
rect 32610 -2785 32645 -2750
rect 32655 -2785 32690 -2750
rect 32700 -2785 32735 -2750
rect 32745 -2785 32780 -2750
rect 32790 -2785 32825 -2750
rect 32835 -2785 32870 -2750
rect 31305 -2830 31340 -2795
rect 31350 -2830 31385 -2795
rect 31395 -2830 31430 -2795
rect 31440 -2830 31475 -2795
rect 31485 -2830 31520 -2795
rect 31530 -2830 31565 -2795
rect 31575 -2830 31610 -2795
rect 31620 -2830 31655 -2795
rect 31665 -2830 31700 -2795
rect 31710 -2830 31745 -2795
rect 31755 -2830 31790 -2795
rect 31800 -2830 31835 -2795
rect 31845 -2830 31880 -2795
rect 31890 -2830 31925 -2795
rect 31935 -2830 31970 -2795
rect 31980 -2830 32015 -2795
rect 32025 -2830 32060 -2795
rect 32070 -2830 32105 -2795
rect 32115 -2830 32150 -2795
rect 32160 -2830 32195 -2795
rect 32205 -2830 32240 -2795
rect 32250 -2830 32285 -2795
rect 32295 -2830 32330 -2795
rect 32340 -2830 32375 -2795
rect 32385 -2830 32420 -2795
rect 32430 -2830 32465 -2795
rect 32475 -2830 32510 -2795
rect 32520 -2830 32555 -2795
rect 32565 -2830 32600 -2795
rect 32610 -2830 32645 -2795
rect 32655 -2830 32690 -2795
rect 32700 -2830 32735 -2795
rect 32745 -2830 32780 -2795
rect 32790 -2830 32825 -2795
rect 32835 -2830 32870 -2795
rect 31305 -2875 31340 -2840
rect 31350 -2875 31385 -2840
rect 31395 -2875 31430 -2840
rect 31440 -2875 31475 -2840
rect 31485 -2875 31520 -2840
rect 31530 -2875 31565 -2840
rect 31575 -2875 31610 -2840
rect 31620 -2875 31655 -2840
rect 31665 -2875 31700 -2840
rect 31710 -2875 31745 -2840
rect 31755 -2875 31790 -2840
rect 31800 -2875 31835 -2840
rect 31845 -2875 31880 -2840
rect 31890 -2875 31925 -2840
rect 31935 -2875 31970 -2840
rect 31980 -2875 32015 -2840
rect 32025 -2875 32060 -2840
rect 32070 -2875 32105 -2840
rect 32115 -2875 32150 -2840
rect 32160 -2875 32195 -2840
rect 32205 -2875 32240 -2840
rect 32250 -2875 32285 -2840
rect 32295 -2875 32330 -2840
rect 32340 -2875 32375 -2840
rect 32385 -2875 32420 -2840
rect 32430 -2875 32465 -2840
rect 32475 -2875 32510 -2840
rect 32520 -2875 32555 -2840
rect 32565 -2875 32600 -2840
rect 32610 -2875 32645 -2840
rect 32655 -2875 32690 -2840
rect 32700 -2875 32735 -2840
rect 32745 -2875 32780 -2840
rect 32790 -2875 32825 -2840
rect 32835 -2875 32870 -2840
<< metal4 >>
rect 2070 19315 32890 19325
rect 2070 19275 2110 19315
rect 2150 19275 6700 19315
rect 6740 19305 32890 19315
rect 6740 19275 31305 19305
rect 2070 19270 31305 19275
rect 31340 19270 31350 19305
rect 31385 19270 31395 19305
rect 31430 19270 31440 19305
rect 31475 19270 31485 19305
rect 31520 19270 31530 19305
rect 31565 19270 31575 19305
rect 31610 19270 31620 19305
rect 31655 19270 31665 19305
rect 31700 19270 31710 19305
rect 31745 19270 31755 19305
rect 31790 19270 31800 19305
rect 31835 19270 31845 19305
rect 31880 19270 31890 19305
rect 31925 19270 31935 19305
rect 31970 19270 31980 19305
rect 32015 19270 32025 19305
rect 32060 19270 32070 19305
rect 32105 19270 32115 19305
rect 32150 19270 32160 19305
rect 32195 19270 32205 19305
rect 32240 19270 32250 19305
rect 32285 19270 32295 19305
rect 32330 19270 32340 19305
rect 32375 19270 32385 19305
rect 32420 19270 32430 19305
rect 32465 19270 32475 19305
rect 32510 19270 32520 19305
rect 32555 19270 32565 19305
rect 32600 19270 32610 19305
rect 32645 19270 32655 19305
rect 32690 19270 32700 19305
rect 32735 19270 32745 19305
rect 32780 19270 32790 19305
rect 32825 19270 32835 19305
rect 32870 19270 32890 19305
rect 2070 19260 32890 19270
rect 2070 19250 31305 19260
rect 2070 19210 2110 19250
rect 2150 19210 6700 19250
rect 6740 19225 31305 19250
rect 31340 19225 31350 19260
rect 31385 19225 31395 19260
rect 31430 19225 31440 19260
rect 31475 19225 31485 19260
rect 31520 19225 31530 19260
rect 31565 19225 31575 19260
rect 31610 19225 31620 19260
rect 31655 19225 31665 19260
rect 31700 19225 31710 19260
rect 31745 19225 31755 19260
rect 31790 19225 31800 19260
rect 31835 19225 31845 19260
rect 31880 19225 31890 19260
rect 31925 19225 31935 19260
rect 31970 19225 31980 19260
rect 32015 19225 32025 19260
rect 32060 19225 32070 19260
rect 32105 19225 32115 19260
rect 32150 19225 32160 19260
rect 32195 19225 32205 19260
rect 32240 19225 32250 19260
rect 32285 19225 32295 19260
rect 32330 19225 32340 19260
rect 32375 19225 32385 19260
rect 32420 19225 32430 19260
rect 32465 19225 32475 19260
rect 32510 19225 32520 19260
rect 32555 19225 32565 19260
rect 32600 19225 32610 19260
rect 32645 19225 32655 19260
rect 32690 19225 32700 19260
rect 32735 19225 32745 19260
rect 32780 19225 32790 19260
rect 32825 19225 32835 19260
rect 32870 19225 32890 19260
rect 6740 19215 32890 19225
rect 6740 19210 31305 19215
rect 2070 19180 31305 19210
rect 31340 19180 31350 19215
rect 31385 19180 31395 19215
rect 31430 19180 31440 19215
rect 31475 19180 31485 19215
rect 31520 19180 31530 19215
rect 31565 19180 31575 19215
rect 31610 19180 31620 19215
rect 31655 19180 31665 19215
rect 31700 19180 31710 19215
rect 31745 19180 31755 19215
rect 31790 19180 31800 19215
rect 31835 19180 31845 19215
rect 31880 19180 31890 19215
rect 31925 19180 31935 19215
rect 31970 19180 31980 19215
rect 32015 19180 32025 19215
rect 32060 19180 32070 19215
rect 32105 19180 32115 19215
rect 32150 19180 32160 19215
rect 32195 19180 32205 19215
rect 32240 19180 32250 19215
rect 32285 19180 32295 19215
rect 32330 19180 32340 19215
rect 32375 19180 32385 19215
rect 32420 19180 32430 19215
rect 32465 19180 32475 19215
rect 32510 19180 32520 19215
rect 32555 19180 32565 19215
rect 32600 19180 32610 19215
rect 32645 19180 32655 19215
rect 32690 19180 32700 19215
rect 32735 19180 32745 19215
rect 32780 19180 32790 19215
rect 32825 19180 32835 19215
rect 32870 19180 32890 19215
rect 2070 19140 2110 19180
rect 2150 19140 6700 19180
rect 6740 19170 32890 19180
rect 6740 19140 31305 19170
rect 2070 19135 31305 19140
rect 31340 19135 31350 19170
rect 31385 19135 31395 19170
rect 31430 19135 31440 19170
rect 31475 19135 31485 19170
rect 31520 19135 31530 19170
rect 31565 19135 31575 19170
rect 31610 19135 31620 19170
rect 31655 19135 31665 19170
rect 31700 19135 31710 19170
rect 31745 19135 31755 19170
rect 31790 19135 31800 19170
rect 31835 19135 31845 19170
rect 31880 19135 31890 19170
rect 31925 19135 31935 19170
rect 31970 19135 31980 19170
rect 32015 19135 32025 19170
rect 32060 19135 32070 19170
rect 32105 19135 32115 19170
rect 32150 19135 32160 19170
rect 32195 19135 32205 19170
rect 32240 19135 32250 19170
rect 32285 19135 32295 19170
rect 32330 19135 32340 19170
rect 32375 19135 32385 19170
rect 32420 19135 32430 19170
rect 32465 19135 32475 19170
rect 32510 19135 32520 19170
rect 32555 19135 32565 19170
rect 32600 19135 32610 19170
rect 32645 19135 32655 19170
rect 32690 19135 32700 19170
rect 32735 19135 32745 19170
rect 32780 19135 32790 19170
rect 32825 19135 32835 19170
rect 32870 19135 32890 19170
rect 2070 19125 32890 19135
rect 2070 19110 31305 19125
rect 2070 19070 2110 19110
rect 2150 19070 6700 19110
rect 6740 19090 31305 19110
rect 31340 19090 31350 19125
rect 31385 19090 31395 19125
rect 31430 19090 31440 19125
rect 31475 19090 31485 19125
rect 31520 19090 31530 19125
rect 31565 19090 31575 19125
rect 31610 19090 31620 19125
rect 31655 19090 31665 19125
rect 31700 19090 31710 19125
rect 31745 19090 31755 19125
rect 31790 19090 31800 19125
rect 31835 19090 31845 19125
rect 31880 19090 31890 19125
rect 31925 19090 31935 19125
rect 31970 19090 31980 19125
rect 32015 19090 32025 19125
rect 32060 19090 32070 19125
rect 32105 19090 32115 19125
rect 32150 19090 32160 19125
rect 32195 19090 32205 19125
rect 32240 19090 32250 19125
rect 32285 19090 32295 19125
rect 32330 19090 32340 19125
rect 32375 19090 32385 19125
rect 32420 19090 32430 19125
rect 32465 19090 32475 19125
rect 32510 19090 32520 19125
rect 32555 19090 32565 19125
rect 32600 19090 32610 19125
rect 32645 19090 32655 19125
rect 32690 19090 32700 19125
rect 32735 19090 32745 19125
rect 32780 19090 32790 19125
rect 32825 19090 32835 19125
rect 32870 19090 32890 19125
rect 6740 19080 32890 19090
rect 6740 19070 31305 19080
rect 2070 19045 31305 19070
rect 31340 19045 31350 19080
rect 31385 19045 31395 19080
rect 31430 19045 31440 19080
rect 31475 19045 31485 19080
rect 31520 19045 31530 19080
rect 31565 19045 31575 19080
rect 31610 19045 31620 19080
rect 31655 19045 31665 19080
rect 31700 19045 31710 19080
rect 31745 19045 31755 19080
rect 31790 19045 31800 19080
rect 31835 19045 31845 19080
rect 31880 19045 31890 19080
rect 31925 19045 31935 19080
rect 31970 19045 31980 19080
rect 32015 19045 32025 19080
rect 32060 19045 32070 19080
rect 32105 19045 32115 19080
rect 32150 19045 32160 19080
rect 32195 19045 32205 19080
rect 32240 19045 32250 19080
rect 32285 19045 32295 19080
rect 32330 19045 32340 19080
rect 32375 19045 32385 19080
rect 32420 19045 32430 19080
rect 32465 19045 32475 19080
rect 32510 19045 32520 19080
rect 32555 19045 32565 19080
rect 32600 19045 32610 19080
rect 32645 19045 32655 19080
rect 32690 19045 32700 19080
rect 32735 19045 32745 19080
rect 32780 19045 32790 19080
rect 32825 19045 32835 19080
rect 32870 19045 32890 19080
rect 2070 19040 32890 19045
rect 2070 19000 2110 19040
rect 2150 19000 6700 19040
rect 6740 19035 32890 19040
rect 6740 19000 31305 19035
rect 31340 19000 31350 19035
rect 31385 19000 31395 19035
rect 31430 19000 31440 19035
rect 31475 19000 31485 19035
rect 31520 19000 31530 19035
rect 31565 19000 31575 19035
rect 31610 19000 31620 19035
rect 31655 19000 31665 19035
rect 31700 19000 31710 19035
rect 31745 19000 31755 19035
rect 31790 19000 31800 19035
rect 31835 19000 31845 19035
rect 31880 19000 31890 19035
rect 31925 19000 31935 19035
rect 31970 19000 31980 19035
rect 32015 19000 32025 19035
rect 32060 19000 32070 19035
rect 32105 19000 32115 19035
rect 32150 19000 32160 19035
rect 32195 19000 32205 19035
rect 32240 19000 32250 19035
rect 32285 19000 32295 19035
rect 32330 19000 32340 19035
rect 32375 19000 32385 19035
rect 32420 19000 32430 19035
rect 32465 19000 32475 19035
rect 32510 19000 32520 19035
rect 32555 19000 32565 19035
rect 32600 19000 32610 19035
rect 32645 19000 32655 19035
rect 32690 19000 32700 19035
rect 32735 19000 32745 19035
rect 32780 19000 32790 19035
rect 32825 19000 32835 19035
rect 32870 19000 32890 19035
rect 2070 18990 32890 19000
rect 2070 18975 31305 18990
rect 2070 18935 2110 18975
rect 2150 18935 6700 18975
rect 6740 18955 31305 18975
rect 31340 18955 31350 18990
rect 31385 18955 31395 18990
rect 31430 18955 31440 18990
rect 31475 18955 31485 18990
rect 31520 18955 31530 18990
rect 31565 18955 31575 18990
rect 31610 18955 31620 18990
rect 31655 18955 31665 18990
rect 31700 18955 31710 18990
rect 31745 18955 31755 18990
rect 31790 18955 31800 18990
rect 31835 18955 31845 18990
rect 31880 18955 31890 18990
rect 31925 18955 31935 18990
rect 31970 18955 31980 18990
rect 32015 18955 32025 18990
rect 32060 18955 32070 18990
rect 32105 18955 32115 18990
rect 32150 18955 32160 18990
rect 32195 18955 32205 18990
rect 32240 18955 32250 18990
rect 32285 18955 32295 18990
rect 32330 18955 32340 18990
rect 32375 18955 32385 18990
rect 32420 18955 32430 18990
rect 32465 18955 32475 18990
rect 32510 18955 32520 18990
rect 32555 18955 32565 18990
rect 32600 18955 32610 18990
rect 32645 18955 32655 18990
rect 32690 18955 32700 18990
rect 32735 18955 32745 18990
rect 32780 18955 32790 18990
rect 32825 18955 32835 18990
rect 32870 18955 32890 18990
rect 6740 18945 32890 18955
rect 6740 18935 31305 18945
rect 2070 18915 31305 18935
rect 2070 18875 2110 18915
rect 2150 18875 6700 18915
rect 6740 18910 31305 18915
rect 31340 18910 31350 18945
rect 31385 18910 31395 18945
rect 31430 18910 31440 18945
rect 31475 18910 31485 18945
rect 31520 18910 31530 18945
rect 31565 18910 31575 18945
rect 31610 18910 31620 18945
rect 31655 18910 31665 18945
rect 31700 18910 31710 18945
rect 31745 18910 31755 18945
rect 31790 18910 31800 18945
rect 31835 18910 31845 18945
rect 31880 18910 31890 18945
rect 31925 18910 31935 18945
rect 31970 18910 31980 18945
rect 32015 18910 32025 18945
rect 32060 18910 32070 18945
rect 32105 18910 32115 18945
rect 32150 18910 32160 18945
rect 32195 18910 32205 18945
rect 32240 18910 32250 18945
rect 32285 18910 32295 18945
rect 32330 18910 32340 18945
rect 32375 18910 32385 18945
rect 32420 18910 32430 18945
rect 32465 18910 32475 18945
rect 32510 18910 32520 18945
rect 32555 18910 32565 18945
rect 32600 18910 32610 18945
rect 32645 18910 32655 18945
rect 32690 18910 32700 18945
rect 32735 18910 32745 18945
rect 32780 18910 32790 18945
rect 32825 18910 32835 18945
rect 32870 18910 32890 18945
rect 6740 18900 32890 18910
rect 6740 18875 31305 18900
rect 2070 18865 31305 18875
rect 31340 18865 31350 18900
rect 31385 18865 31395 18900
rect 31430 18865 31440 18900
rect 31475 18865 31485 18900
rect 31520 18865 31530 18900
rect 31565 18865 31575 18900
rect 31610 18865 31620 18900
rect 31655 18865 31665 18900
rect 31700 18865 31710 18900
rect 31745 18865 31755 18900
rect 31790 18865 31800 18900
rect 31835 18865 31845 18900
rect 31880 18865 31890 18900
rect 31925 18865 31935 18900
rect 31970 18865 31980 18900
rect 32015 18865 32025 18900
rect 32060 18865 32070 18900
rect 32105 18865 32115 18900
rect 32150 18865 32160 18900
rect 32195 18865 32205 18900
rect 32240 18865 32250 18900
rect 32285 18865 32295 18900
rect 32330 18865 32340 18900
rect 32375 18865 32385 18900
rect 32420 18865 32430 18900
rect 32465 18865 32475 18900
rect 32510 18865 32520 18900
rect 32555 18865 32565 18900
rect 32600 18865 32610 18900
rect 32645 18865 32655 18900
rect 32690 18865 32700 18900
rect 32735 18865 32745 18900
rect 32780 18865 32790 18900
rect 32825 18865 32835 18900
rect 32870 18865 32890 18900
rect 2070 18855 32890 18865
rect 2070 18850 31305 18855
rect 2070 18810 2110 18850
rect 2150 18810 6700 18850
rect 6740 18820 31305 18850
rect 31340 18820 31350 18855
rect 31385 18820 31395 18855
rect 31430 18820 31440 18855
rect 31475 18820 31485 18855
rect 31520 18820 31530 18855
rect 31565 18820 31575 18855
rect 31610 18820 31620 18855
rect 31655 18820 31665 18855
rect 31700 18820 31710 18855
rect 31745 18820 31755 18855
rect 31790 18820 31800 18855
rect 31835 18820 31845 18855
rect 31880 18820 31890 18855
rect 31925 18820 31935 18855
rect 31970 18820 31980 18855
rect 32015 18820 32025 18855
rect 32060 18820 32070 18855
rect 32105 18820 32115 18855
rect 32150 18820 32160 18855
rect 32195 18820 32205 18855
rect 32240 18820 32250 18855
rect 32285 18820 32295 18855
rect 32330 18820 32340 18855
rect 32375 18820 32385 18855
rect 32420 18820 32430 18855
rect 32465 18820 32475 18855
rect 32510 18820 32520 18855
rect 32555 18820 32565 18855
rect 32600 18820 32610 18855
rect 32645 18820 32655 18855
rect 32690 18820 32700 18855
rect 32735 18820 32745 18855
rect 32780 18820 32790 18855
rect 32825 18820 32835 18855
rect 32870 18820 32890 18855
rect 6740 18810 32890 18820
rect 2070 18780 31305 18810
rect 2070 18740 2110 18780
rect 2150 18740 6700 18780
rect 6740 18775 31305 18780
rect 31340 18775 31350 18810
rect 31385 18775 31395 18810
rect 31430 18775 31440 18810
rect 31475 18775 31485 18810
rect 31520 18775 31530 18810
rect 31565 18775 31575 18810
rect 31610 18775 31620 18810
rect 31655 18775 31665 18810
rect 31700 18775 31710 18810
rect 31745 18775 31755 18810
rect 31790 18775 31800 18810
rect 31835 18775 31845 18810
rect 31880 18775 31890 18810
rect 31925 18775 31935 18810
rect 31970 18775 31980 18810
rect 32015 18775 32025 18810
rect 32060 18775 32070 18810
rect 32105 18775 32115 18810
rect 32150 18775 32160 18810
rect 32195 18775 32205 18810
rect 32240 18775 32250 18810
rect 32285 18775 32295 18810
rect 32330 18775 32340 18810
rect 32375 18775 32385 18810
rect 32420 18775 32430 18810
rect 32465 18775 32475 18810
rect 32510 18775 32520 18810
rect 32555 18775 32565 18810
rect 32600 18775 32610 18810
rect 32645 18775 32655 18810
rect 32690 18775 32700 18810
rect 32735 18775 32745 18810
rect 32780 18775 32790 18810
rect 32825 18775 32835 18810
rect 32870 18775 32890 18810
rect 6740 18765 32890 18775
rect 6740 18740 31305 18765
rect 2070 18730 31305 18740
rect 31340 18730 31350 18765
rect 31385 18730 31395 18765
rect 31430 18730 31440 18765
rect 31475 18730 31485 18765
rect 31520 18730 31530 18765
rect 31565 18730 31575 18765
rect 31610 18730 31620 18765
rect 31655 18730 31665 18765
rect 31700 18730 31710 18765
rect 31745 18730 31755 18765
rect 31790 18730 31800 18765
rect 31835 18730 31845 18765
rect 31880 18730 31890 18765
rect 31925 18730 31935 18765
rect 31970 18730 31980 18765
rect 32015 18730 32025 18765
rect 32060 18730 32070 18765
rect 32105 18730 32115 18765
rect 32150 18730 32160 18765
rect 32195 18730 32205 18765
rect 32240 18730 32250 18765
rect 32285 18730 32295 18765
rect 32330 18730 32340 18765
rect 32375 18730 32385 18765
rect 32420 18730 32430 18765
rect 32465 18730 32475 18765
rect 32510 18730 32520 18765
rect 32555 18730 32565 18765
rect 32600 18730 32610 18765
rect 32645 18730 32655 18765
rect 32690 18730 32700 18765
rect 32735 18730 32745 18765
rect 32780 18730 32790 18765
rect 32825 18730 32835 18765
rect 32870 18730 32890 18765
rect 2070 18720 32890 18730
rect 2070 18710 31305 18720
rect 2070 18670 2110 18710
rect 2150 18670 6700 18710
rect 6740 18685 31305 18710
rect 31340 18685 31350 18720
rect 31385 18685 31395 18720
rect 31430 18685 31440 18720
rect 31475 18685 31485 18720
rect 31520 18685 31530 18720
rect 31565 18685 31575 18720
rect 31610 18685 31620 18720
rect 31655 18685 31665 18720
rect 31700 18685 31710 18720
rect 31745 18685 31755 18720
rect 31790 18685 31800 18720
rect 31835 18685 31845 18720
rect 31880 18685 31890 18720
rect 31925 18685 31935 18720
rect 31970 18685 31980 18720
rect 32015 18685 32025 18720
rect 32060 18685 32070 18720
rect 32105 18685 32115 18720
rect 32150 18685 32160 18720
rect 32195 18685 32205 18720
rect 32240 18685 32250 18720
rect 32285 18685 32295 18720
rect 32330 18685 32340 18720
rect 32375 18685 32385 18720
rect 32420 18685 32430 18720
rect 32465 18685 32475 18720
rect 32510 18685 32520 18720
rect 32555 18685 32565 18720
rect 32600 18685 32610 18720
rect 32645 18685 32655 18720
rect 32690 18685 32700 18720
rect 32735 18685 32745 18720
rect 32780 18685 32790 18720
rect 32825 18685 32835 18720
rect 32870 18685 32890 18720
rect 6740 18675 32890 18685
rect 6740 18670 31305 18675
rect 2070 18640 31305 18670
rect 31340 18640 31350 18675
rect 31385 18640 31395 18675
rect 31430 18640 31440 18675
rect 31475 18640 31485 18675
rect 31520 18640 31530 18675
rect 31565 18640 31575 18675
rect 31610 18640 31620 18675
rect 31655 18640 31665 18675
rect 31700 18640 31710 18675
rect 31745 18640 31755 18675
rect 31790 18640 31800 18675
rect 31835 18640 31845 18675
rect 31880 18640 31890 18675
rect 31925 18640 31935 18675
rect 31970 18640 31980 18675
rect 32015 18640 32025 18675
rect 32060 18640 32070 18675
rect 32105 18640 32115 18675
rect 32150 18640 32160 18675
rect 32195 18640 32205 18675
rect 32240 18640 32250 18675
rect 32285 18640 32295 18675
rect 32330 18640 32340 18675
rect 32375 18640 32385 18675
rect 32420 18640 32430 18675
rect 32465 18640 32475 18675
rect 32510 18640 32520 18675
rect 32555 18640 32565 18675
rect 32600 18640 32610 18675
rect 32645 18640 32655 18675
rect 32690 18640 32700 18675
rect 32735 18640 32745 18675
rect 32780 18640 32790 18675
rect 32825 18640 32835 18675
rect 32870 18640 32890 18675
rect 2070 18600 2110 18640
rect 2150 18600 6700 18640
rect 6740 18630 32890 18640
rect 6740 18600 31305 18630
rect 2070 18595 31305 18600
rect 31340 18595 31350 18630
rect 31385 18595 31395 18630
rect 31430 18595 31440 18630
rect 31475 18595 31485 18630
rect 31520 18595 31530 18630
rect 31565 18595 31575 18630
rect 31610 18595 31620 18630
rect 31655 18595 31665 18630
rect 31700 18595 31710 18630
rect 31745 18595 31755 18630
rect 31790 18595 31800 18630
rect 31835 18595 31845 18630
rect 31880 18595 31890 18630
rect 31925 18595 31935 18630
rect 31970 18595 31980 18630
rect 32015 18595 32025 18630
rect 32060 18595 32070 18630
rect 32105 18595 32115 18630
rect 32150 18595 32160 18630
rect 32195 18595 32205 18630
rect 32240 18595 32250 18630
rect 32285 18595 32295 18630
rect 32330 18595 32340 18630
rect 32375 18595 32385 18630
rect 32420 18595 32430 18630
rect 32465 18595 32475 18630
rect 32510 18595 32520 18630
rect 32555 18595 32565 18630
rect 32600 18595 32610 18630
rect 32645 18595 32655 18630
rect 32690 18595 32700 18630
rect 32735 18595 32745 18630
rect 32780 18595 32790 18630
rect 32825 18595 32835 18630
rect 32870 18595 32890 18630
rect 2070 18585 32890 18595
rect 2070 18575 31305 18585
rect 2070 18535 2110 18575
rect 2150 18535 6700 18575
rect 6740 18550 31305 18575
rect 31340 18550 31350 18585
rect 31385 18550 31395 18585
rect 31430 18550 31440 18585
rect 31475 18550 31485 18585
rect 31520 18550 31530 18585
rect 31565 18550 31575 18585
rect 31610 18550 31620 18585
rect 31655 18550 31665 18585
rect 31700 18550 31710 18585
rect 31745 18550 31755 18585
rect 31790 18550 31800 18585
rect 31835 18550 31845 18585
rect 31880 18550 31890 18585
rect 31925 18550 31935 18585
rect 31970 18550 31980 18585
rect 32015 18550 32025 18585
rect 32060 18550 32070 18585
rect 32105 18550 32115 18585
rect 32150 18550 32160 18585
rect 32195 18550 32205 18585
rect 32240 18550 32250 18585
rect 32285 18550 32295 18585
rect 32330 18550 32340 18585
rect 32375 18550 32385 18585
rect 32420 18550 32430 18585
rect 32465 18550 32475 18585
rect 32510 18550 32520 18585
rect 32555 18550 32565 18585
rect 32600 18550 32610 18585
rect 32645 18550 32655 18585
rect 32690 18550 32700 18585
rect 32735 18550 32745 18585
rect 32780 18550 32790 18585
rect 32825 18550 32835 18585
rect 32870 18550 32890 18585
rect 6740 18540 32890 18550
rect 6740 18535 31305 18540
rect 2070 18515 31305 18535
rect 2070 18475 2110 18515
rect 2150 18475 6700 18515
rect 6740 18505 31305 18515
rect 31340 18505 31350 18540
rect 31385 18505 31395 18540
rect 31430 18505 31440 18540
rect 31475 18505 31485 18540
rect 31520 18505 31530 18540
rect 31565 18505 31575 18540
rect 31610 18505 31620 18540
rect 31655 18505 31665 18540
rect 31700 18505 31710 18540
rect 31745 18505 31755 18540
rect 31790 18505 31800 18540
rect 31835 18505 31845 18540
rect 31880 18505 31890 18540
rect 31925 18505 31935 18540
rect 31970 18505 31980 18540
rect 32015 18505 32025 18540
rect 32060 18505 32070 18540
rect 32105 18505 32115 18540
rect 32150 18505 32160 18540
rect 32195 18505 32205 18540
rect 32240 18505 32250 18540
rect 32285 18505 32295 18540
rect 32330 18505 32340 18540
rect 32375 18505 32385 18540
rect 32420 18505 32430 18540
rect 32465 18505 32475 18540
rect 32510 18505 32520 18540
rect 32555 18505 32565 18540
rect 32600 18505 32610 18540
rect 32645 18505 32655 18540
rect 32690 18505 32700 18540
rect 32735 18505 32745 18540
rect 32780 18505 32790 18540
rect 32825 18505 32835 18540
rect 32870 18505 32890 18540
rect 6740 18495 32890 18505
rect 6740 18475 31305 18495
rect 2070 18460 31305 18475
rect 31340 18460 31350 18495
rect 31385 18460 31395 18495
rect 31430 18460 31440 18495
rect 31475 18460 31485 18495
rect 31520 18460 31530 18495
rect 31565 18460 31575 18495
rect 31610 18460 31620 18495
rect 31655 18460 31665 18495
rect 31700 18460 31710 18495
rect 31745 18460 31755 18495
rect 31790 18460 31800 18495
rect 31835 18460 31845 18495
rect 31880 18460 31890 18495
rect 31925 18460 31935 18495
rect 31970 18460 31980 18495
rect 32015 18460 32025 18495
rect 32060 18460 32070 18495
rect 32105 18460 32115 18495
rect 32150 18460 32160 18495
rect 32195 18460 32205 18495
rect 32240 18460 32250 18495
rect 32285 18460 32295 18495
rect 32330 18460 32340 18495
rect 32375 18460 32385 18495
rect 32420 18460 32430 18495
rect 32465 18460 32475 18495
rect 32510 18460 32520 18495
rect 32555 18460 32565 18495
rect 32600 18460 32610 18495
rect 32645 18460 32655 18495
rect 32690 18460 32700 18495
rect 32735 18460 32745 18495
rect 32780 18460 32790 18495
rect 32825 18460 32835 18495
rect 32870 18460 32890 18495
rect 2070 18450 32890 18460
rect 2070 18410 2110 18450
rect 2150 18410 6700 18450
rect 6740 18415 31305 18450
rect 31340 18415 31350 18450
rect 31385 18415 31395 18450
rect 31430 18415 31440 18450
rect 31475 18415 31485 18450
rect 31520 18415 31530 18450
rect 31565 18415 31575 18450
rect 31610 18415 31620 18450
rect 31655 18415 31665 18450
rect 31700 18415 31710 18450
rect 31745 18415 31755 18450
rect 31790 18415 31800 18450
rect 31835 18415 31845 18450
rect 31880 18415 31890 18450
rect 31925 18415 31935 18450
rect 31970 18415 31980 18450
rect 32015 18415 32025 18450
rect 32060 18415 32070 18450
rect 32105 18415 32115 18450
rect 32150 18415 32160 18450
rect 32195 18415 32205 18450
rect 32240 18415 32250 18450
rect 32285 18415 32295 18450
rect 32330 18415 32340 18450
rect 32375 18415 32385 18450
rect 32420 18415 32430 18450
rect 32465 18415 32475 18450
rect 32510 18415 32520 18450
rect 32555 18415 32565 18450
rect 32600 18415 32610 18450
rect 32645 18415 32655 18450
rect 32690 18415 32700 18450
rect 32735 18415 32745 18450
rect 32780 18415 32790 18450
rect 32825 18415 32835 18450
rect 32870 18415 32890 18450
rect 6740 18410 32890 18415
rect 2070 18405 32890 18410
rect 2070 18380 31305 18405
rect 2070 18340 2110 18380
rect 2150 18340 6700 18380
rect 6740 18370 31305 18380
rect 31340 18370 31350 18405
rect 31385 18370 31395 18405
rect 31430 18370 31440 18405
rect 31475 18370 31485 18405
rect 31520 18370 31530 18405
rect 31565 18370 31575 18405
rect 31610 18370 31620 18405
rect 31655 18370 31665 18405
rect 31700 18370 31710 18405
rect 31745 18370 31755 18405
rect 31790 18370 31800 18405
rect 31835 18370 31845 18405
rect 31880 18370 31890 18405
rect 31925 18370 31935 18405
rect 31970 18370 31980 18405
rect 32015 18370 32025 18405
rect 32060 18370 32070 18405
rect 32105 18370 32115 18405
rect 32150 18370 32160 18405
rect 32195 18370 32205 18405
rect 32240 18370 32250 18405
rect 32285 18370 32295 18405
rect 32330 18370 32340 18405
rect 32375 18370 32385 18405
rect 32420 18370 32430 18405
rect 32465 18370 32475 18405
rect 32510 18370 32520 18405
rect 32555 18370 32565 18405
rect 32600 18370 32610 18405
rect 32645 18370 32655 18405
rect 32690 18370 32700 18405
rect 32735 18370 32745 18405
rect 32780 18370 32790 18405
rect 32825 18370 32835 18405
rect 32870 18370 32890 18405
rect 6740 18360 32890 18370
rect 6740 18340 31305 18360
rect 2070 18325 31305 18340
rect 31340 18325 31350 18360
rect 31385 18325 31395 18360
rect 31430 18325 31440 18360
rect 31475 18325 31485 18360
rect 31520 18325 31530 18360
rect 31565 18325 31575 18360
rect 31610 18325 31620 18360
rect 31655 18325 31665 18360
rect 31700 18325 31710 18360
rect 31745 18325 31755 18360
rect 31790 18325 31800 18360
rect 31835 18325 31845 18360
rect 31880 18325 31890 18360
rect 31925 18325 31935 18360
rect 31970 18325 31980 18360
rect 32015 18325 32025 18360
rect 32060 18325 32070 18360
rect 32105 18325 32115 18360
rect 32150 18325 32160 18360
rect 32195 18325 32205 18360
rect 32240 18325 32250 18360
rect 32285 18325 32295 18360
rect 32330 18325 32340 18360
rect 32375 18325 32385 18360
rect 32420 18325 32430 18360
rect 32465 18325 32475 18360
rect 32510 18325 32520 18360
rect 32555 18325 32565 18360
rect 32600 18325 32610 18360
rect 32645 18325 32655 18360
rect 32690 18325 32700 18360
rect 32735 18325 32745 18360
rect 32780 18325 32790 18360
rect 32825 18325 32835 18360
rect 32870 18325 32890 18360
rect 2070 18315 32890 18325
rect 2070 18310 31305 18315
rect 2070 18270 2110 18310
rect 2150 18270 6700 18310
rect 6740 18280 31305 18310
rect 31340 18280 31350 18315
rect 31385 18280 31395 18315
rect 31430 18280 31440 18315
rect 31475 18280 31485 18315
rect 31520 18280 31530 18315
rect 31565 18280 31575 18315
rect 31610 18280 31620 18315
rect 31655 18280 31665 18315
rect 31700 18280 31710 18315
rect 31745 18280 31755 18315
rect 31790 18280 31800 18315
rect 31835 18280 31845 18315
rect 31880 18280 31890 18315
rect 31925 18280 31935 18315
rect 31970 18280 31980 18315
rect 32015 18280 32025 18315
rect 32060 18280 32070 18315
rect 32105 18280 32115 18315
rect 32150 18280 32160 18315
rect 32195 18280 32205 18315
rect 32240 18280 32250 18315
rect 32285 18280 32295 18315
rect 32330 18280 32340 18315
rect 32375 18280 32385 18315
rect 32420 18280 32430 18315
rect 32465 18280 32475 18315
rect 32510 18280 32520 18315
rect 32555 18280 32565 18315
rect 32600 18280 32610 18315
rect 32645 18280 32655 18315
rect 32690 18280 32700 18315
rect 32735 18280 32745 18315
rect 32780 18280 32790 18315
rect 32825 18280 32835 18315
rect 32870 18280 32890 18315
rect 6740 18270 32890 18280
rect 2070 18240 31305 18270
rect 2070 18200 2110 18240
rect 2150 18200 6700 18240
rect 6740 18235 31305 18240
rect 31340 18235 31350 18270
rect 31385 18235 31395 18270
rect 31430 18235 31440 18270
rect 31475 18235 31485 18270
rect 31520 18235 31530 18270
rect 31565 18235 31575 18270
rect 31610 18235 31620 18270
rect 31655 18235 31665 18270
rect 31700 18235 31710 18270
rect 31745 18235 31755 18270
rect 31790 18235 31800 18270
rect 31835 18235 31845 18270
rect 31880 18235 31890 18270
rect 31925 18235 31935 18270
rect 31970 18235 31980 18270
rect 32015 18235 32025 18270
rect 32060 18235 32070 18270
rect 32105 18235 32115 18270
rect 32150 18235 32160 18270
rect 32195 18235 32205 18270
rect 32240 18235 32250 18270
rect 32285 18235 32295 18270
rect 32330 18235 32340 18270
rect 32375 18235 32385 18270
rect 32420 18235 32430 18270
rect 32465 18235 32475 18270
rect 32510 18235 32520 18270
rect 32555 18235 32565 18270
rect 32600 18235 32610 18270
rect 32645 18235 32655 18270
rect 32690 18235 32700 18270
rect 32735 18235 32745 18270
rect 32780 18235 32790 18270
rect 32825 18235 32835 18270
rect 32870 18235 32890 18270
rect 6740 18225 32890 18235
rect 6740 18200 31305 18225
rect 2070 18190 31305 18200
rect 31340 18190 31350 18225
rect 31385 18190 31395 18225
rect 31430 18190 31440 18225
rect 31475 18190 31485 18225
rect 31520 18190 31530 18225
rect 31565 18190 31575 18225
rect 31610 18190 31620 18225
rect 31655 18190 31665 18225
rect 31700 18190 31710 18225
rect 31745 18190 31755 18225
rect 31790 18190 31800 18225
rect 31835 18190 31845 18225
rect 31880 18190 31890 18225
rect 31925 18190 31935 18225
rect 31970 18190 31980 18225
rect 32015 18190 32025 18225
rect 32060 18190 32070 18225
rect 32105 18190 32115 18225
rect 32150 18190 32160 18225
rect 32195 18190 32205 18225
rect 32240 18190 32250 18225
rect 32285 18190 32295 18225
rect 32330 18190 32340 18225
rect 32375 18190 32385 18225
rect 32420 18190 32430 18225
rect 32465 18190 32475 18225
rect 32510 18190 32520 18225
rect 32555 18190 32565 18225
rect 32600 18190 32610 18225
rect 32645 18190 32655 18225
rect 32690 18190 32700 18225
rect 32735 18190 32745 18225
rect 32780 18190 32790 18225
rect 32825 18190 32835 18225
rect 32870 18190 32890 18225
rect 2070 18180 32890 18190
rect 2070 18175 31305 18180
rect 2070 18135 2110 18175
rect 2150 18135 6700 18175
rect 6740 18145 31305 18175
rect 31340 18145 31350 18180
rect 31385 18145 31395 18180
rect 31430 18145 31440 18180
rect 31475 18145 31485 18180
rect 31520 18145 31530 18180
rect 31565 18145 31575 18180
rect 31610 18145 31620 18180
rect 31655 18145 31665 18180
rect 31700 18145 31710 18180
rect 31745 18145 31755 18180
rect 31790 18145 31800 18180
rect 31835 18145 31845 18180
rect 31880 18145 31890 18180
rect 31925 18145 31935 18180
rect 31970 18145 31980 18180
rect 32015 18145 32025 18180
rect 32060 18145 32070 18180
rect 32105 18145 32115 18180
rect 32150 18145 32160 18180
rect 32195 18145 32205 18180
rect 32240 18145 32250 18180
rect 32285 18145 32295 18180
rect 32330 18145 32340 18180
rect 32375 18145 32385 18180
rect 32420 18145 32430 18180
rect 32465 18145 32475 18180
rect 32510 18145 32520 18180
rect 32555 18145 32565 18180
rect 32600 18145 32610 18180
rect 32645 18145 32655 18180
rect 32690 18145 32700 18180
rect 32735 18145 32745 18180
rect 32780 18145 32790 18180
rect 32825 18145 32835 18180
rect 32870 18145 32890 18180
rect 6740 18135 32890 18145
rect 2070 18115 31305 18135
rect 2070 18075 2110 18115
rect 2150 18075 6700 18115
rect 6740 18100 31305 18115
rect 31340 18100 31350 18135
rect 31385 18100 31395 18135
rect 31430 18100 31440 18135
rect 31475 18100 31485 18135
rect 31520 18100 31530 18135
rect 31565 18100 31575 18135
rect 31610 18100 31620 18135
rect 31655 18100 31665 18135
rect 31700 18100 31710 18135
rect 31745 18100 31755 18135
rect 31790 18100 31800 18135
rect 31835 18100 31845 18135
rect 31880 18100 31890 18135
rect 31925 18100 31935 18135
rect 31970 18100 31980 18135
rect 32015 18100 32025 18135
rect 32060 18100 32070 18135
rect 32105 18100 32115 18135
rect 32150 18100 32160 18135
rect 32195 18100 32205 18135
rect 32240 18100 32250 18135
rect 32285 18100 32295 18135
rect 32330 18100 32340 18135
rect 32375 18100 32385 18135
rect 32420 18100 32430 18135
rect 32465 18100 32475 18135
rect 32510 18100 32520 18135
rect 32555 18100 32565 18135
rect 32600 18100 32610 18135
rect 32645 18100 32655 18135
rect 32690 18100 32700 18135
rect 32735 18100 32745 18135
rect 32780 18100 32790 18135
rect 32825 18100 32835 18135
rect 32870 18100 32890 18135
rect 6740 18090 32890 18100
rect 6740 18075 31305 18090
rect 2070 18055 31305 18075
rect 31340 18055 31350 18090
rect 31385 18055 31395 18090
rect 31430 18055 31440 18090
rect 31475 18055 31485 18090
rect 31520 18055 31530 18090
rect 31565 18055 31575 18090
rect 31610 18055 31620 18090
rect 31655 18055 31665 18090
rect 31700 18055 31710 18090
rect 31745 18055 31755 18090
rect 31790 18055 31800 18090
rect 31835 18055 31845 18090
rect 31880 18055 31890 18090
rect 31925 18055 31935 18090
rect 31970 18055 31980 18090
rect 32015 18055 32025 18090
rect 32060 18055 32070 18090
rect 32105 18055 32115 18090
rect 32150 18055 32160 18090
rect 32195 18055 32205 18090
rect 32240 18055 32250 18090
rect 32285 18055 32295 18090
rect 32330 18055 32340 18090
rect 32375 18055 32385 18090
rect 32420 18055 32430 18090
rect 32465 18055 32475 18090
rect 32510 18055 32520 18090
rect 32555 18055 32565 18090
rect 32600 18055 32610 18090
rect 32645 18055 32655 18090
rect 32690 18055 32700 18090
rect 32735 18055 32745 18090
rect 32780 18055 32790 18090
rect 32825 18055 32835 18090
rect 32870 18055 32890 18090
rect 2070 18050 32890 18055
rect 2070 18010 2110 18050
rect 2150 18010 6700 18050
rect 6740 18045 32890 18050
rect 6740 18010 31305 18045
rect 31340 18010 31350 18045
rect 31385 18010 31395 18045
rect 31430 18010 31440 18045
rect 31475 18010 31485 18045
rect 31520 18010 31530 18045
rect 31565 18010 31575 18045
rect 31610 18010 31620 18045
rect 31655 18010 31665 18045
rect 31700 18010 31710 18045
rect 31745 18010 31755 18045
rect 31790 18010 31800 18045
rect 31835 18010 31845 18045
rect 31880 18010 31890 18045
rect 31925 18010 31935 18045
rect 31970 18010 31980 18045
rect 32015 18010 32025 18045
rect 32060 18010 32070 18045
rect 32105 18010 32115 18045
rect 32150 18010 32160 18045
rect 32195 18010 32205 18045
rect 32240 18010 32250 18045
rect 32285 18010 32295 18045
rect 32330 18010 32340 18045
rect 32375 18010 32385 18045
rect 32420 18010 32430 18045
rect 32465 18010 32475 18045
rect 32510 18010 32520 18045
rect 32555 18010 32565 18045
rect 32600 18010 32610 18045
rect 32645 18010 32655 18045
rect 32690 18010 32700 18045
rect 32735 18010 32745 18045
rect 32780 18010 32790 18045
rect 32825 18010 32835 18045
rect 32870 18010 32890 18045
rect 2070 18000 32890 18010
rect 2070 17980 31305 18000
rect 2070 17940 2110 17980
rect 2150 17940 6700 17980
rect 6740 17965 31305 17980
rect 31340 17965 31350 18000
rect 31385 17965 31395 18000
rect 31430 17965 31440 18000
rect 31475 17965 31485 18000
rect 31520 17965 31530 18000
rect 31565 17965 31575 18000
rect 31610 17965 31620 18000
rect 31655 17965 31665 18000
rect 31700 17965 31710 18000
rect 31745 17965 31755 18000
rect 31790 17965 31800 18000
rect 31835 17965 31845 18000
rect 31880 17965 31890 18000
rect 31925 17965 31935 18000
rect 31970 17965 31980 18000
rect 32015 17965 32025 18000
rect 32060 17965 32070 18000
rect 32105 17965 32115 18000
rect 32150 17965 32160 18000
rect 32195 17965 32205 18000
rect 32240 17965 32250 18000
rect 32285 17965 32295 18000
rect 32330 17965 32340 18000
rect 32375 17965 32385 18000
rect 32420 17965 32430 18000
rect 32465 17965 32475 18000
rect 32510 17965 32520 18000
rect 32555 17965 32565 18000
rect 32600 17965 32610 18000
rect 32645 17965 32655 18000
rect 32690 17965 32700 18000
rect 32735 17965 32745 18000
rect 32780 17965 32790 18000
rect 32825 17965 32835 18000
rect 32870 17965 32890 18000
rect 6740 17955 32890 17965
rect 6740 17940 31305 17955
rect 2070 17920 31305 17940
rect 31340 17920 31350 17955
rect 31385 17920 31395 17955
rect 31430 17920 31440 17955
rect 31475 17920 31485 17955
rect 31520 17920 31530 17955
rect 31565 17920 31575 17955
rect 31610 17920 31620 17955
rect 31655 17920 31665 17955
rect 31700 17920 31710 17955
rect 31745 17920 31755 17955
rect 31790 17920 31800 17955
rect 31835 17920 31845 17955
rect 31880 17920 31890 17955
rect 31925 17920 31935 17955
rect 31970 17920 31980 17955
rect 32015 17920 32025 17955
rect 32060 17920 32070 17955
rect 32105 17920 32115 17955
rect 32150 17920 32160 17955
rect 32195 17920 32205 17955
rect 32240 17920 32250 17955
rect 32285 17920 32295 17955
rect 32330 17920 32340 17955
rect 32375 17920 32385 17955
rect 32420 17920 32430 17955
rect 32465 17920 32475 17955
rect 32510 17920 32520 17955
rect 32555 17920 32565 17955
rect 32600 17920 32610 17955
rect 32645 17920 32655 17955
rect 32690 17920 32700 17955
rect 32735 17920 32745 17955
rect 32780 17920 32790 17955
rect 32825 17920 32835 17955
rect 32870 17920 32890 17955
rect 2070 17910 32890 17920
rect 2070 17870 2110 17910
rect 2150 17870 6700 17910
rect 6740 17875 31305 17910
rect 31340 17875 31350 17910
rect 31385 17875 31395 17910
rect 31430 17875 31440 17910
rect 31475 17875 31485 17910
rect 31520 17875 31530 17910
rect 31565 17875 31575 17910
rect 31610 17875 31620 17910
rect 31655 17875 31665 17910
rect 31700 17875 31710 17910
rect 31745 17875 31755 17910
rect 31790 17875 31800 17910
rect 31835 17875 31845 17910
rect 31880 17875 31890 17910
rect 31925 17875 31935 17910
rect 31970 17875 31980 17910
rect 32015 17875 32025 17910
rect 32060 17875 32070 17910
rect 32105 17875 32115 17910
rect 32150 17875 32160 17910
rect 32195 17875 32205 17910
rect 32240 17875 32250 17910
rect 32285 17875 32295 17910
rect 32330 17875 32340 17910
rect 32375 17875 32385 17910
rect 32420 17875 32430 17910
rect 32465 17875 32475 17910
rect 32510 17875 32520 17910
rect 32555 17875 32565 17910
rect 32600 17875 32610 17910
rect 32645 17875 32655 17910
rect 32690 17875 32700 17910
rect 32735 17875 32745 17910
rect 32780 17875 32790 17910
rect 32825 17875 32835 17910
rect 32870 17875 32890 17910
rect 6740 17870 32890 17875
rect 2070 17865 32890 17870
rect 2070 17840 31305 17865
rect 2070 17800 2110 17840
rect 2150 17800 6700 17840
rect 6740 17830 31305 17840
rect 31340 17830 31350 17865
rect 31385 17830 31395 17865
rect 31430 17830 31440 17865
rect 31475 17830 31485 17865
rect 31520 17830 31530 17865
rect 31565 17830 31575 17865
rect 31610 17830 31620 17865
rect 31655 17830 31665 17865
rect 31700 17830 31710 17865
rect 31745 17830 31755 17865
rect 31790 17830 31800 17865
rect 31835 17830 31845 17865
rect 31880 17830 31890 17865
rect 31925 17830 31935 17865
rect 31970 17830 31980 17865
rect 32015 17830 32025 17865
rect 32060 17830 32070 17865
rect 32105 17830 32115 17865
rect 32150 17830 32160 17865
rect 32195 17830 32205 17865
rect 32240 17830 32250 17865
rect 32285 17830 32295 17865
rect 32330 17830 32340 17865
rect 32375 17830 32385 17865
rect 32420 17830 32430 17865
rect 32465 17830 32475 17865
rect 32510 17830 32520 17865
rect 32555 17830 32565 17865
rect 32600 17830 32610 17865
rect 32645 17830 32655 17865
rect 32690 17830 32700 17865
rect 32735 17830 32745 17865
rect 32780 17830 32790 17865
rect 32825 17830 32835 17865
rect 32870 17830 32890 17865
rect 6740 17820 32890 17830
rect 6740 17800 31305 17820
rect 2070 17785 31305 17800
rect 31340 17785 31350 17820
rect 31385 17785 31395 17820
rect 31430 17785 31440 17820
rect 31475 17785 31485 17820
rect 31520 17785 31530 17820
rect 31565 17785 31575 17820
rect 31610 17785 31620 17820
rect 31655 17785 31665 17820
rect 31700 17785 31710 17820
rect 31745 17785 31755 17820
rect 31790 17785 31800 17820
rect 31835 17785 31845 17820
rect 31880 17785 31890 17820
rect 31925 17785 31935 17820
rect 31970 17785 31980 17820
rect 32015 17785 32025 17820
rect 32060 17785 32070 17820
rect 32105 17785 32115 17820
rect 32150 17785 32160 17820
rect 32195 17785 32205 17820
rect 32240 17785 32250 17820
rect 32285 17785 32295 17820
rect 32330 17785 32340 17820
rect 32375 17785 32385 17820
rect 32420 17785 32430 17820
rect 32465 17785 32475 17820
rect 32510 17785 32520 17820
rect 32555 17785 32565 17820
rect 32600 17785 32610 17820
rect 32645 17785 32655 17820
rect 32690 17785 32700 17820
rect 32735 17785 32745 17820
rect 32780 17785 32790 17820
rect 32825 17785 32835 17820
rect 32870 17785 32890 17820
rect 2070 17775 32890 17785
rect 2070 17735 2110 17775
rect 2150 17735 6700 17775
rect 6740 17740 31305 17775
rect 31340 17740 31350 17775
rect 31385 17740 31395 17775
rect 31430 17740 31440 17775
rect 31475 17740 31485 17775
rect 31520 17740 31530 17775
rect 31565 17740 31575 17775
rect 31610 17740 31620 17775
rect 31655 17740 31665 17775
rect 31700 17740 31710 17775
rect 31745 17740 31755 17775
rect 31790 17740 31800 17775
rect 31835 17740 31845 17775
rect 31880 17740 31890 17775
rect 31925 17740 31935 17775
rect 31970 17740 31980 17775
rect 32015 17740 32025 17775
rect 32060 17740 32070 17775
rect 32105 17740 32115 17775
rect 32150 17740 32160 17775
rect 32195 17740 32205 17775
rect 32240 17740 32250 17775
rect 32285 17740 32295 17775
rect 32330 17740 32340 17775
rect 32375 17740 32385 17775
rect 32420 17740 32430 17775
rect 32465 17740 32475 17775
rect 32510 17740 32520 17775
rect 32555 17740 32565 17775
rect 32600 17740 32610 17775
rect 32645 17740 32655 17775
rect 32690 17740 32700 17775
rect 32735 17740 32745 17775
rect 32780 17740 32790 17775
rect 32825 17740 32835 17775
rect 32870 17740 32890 17775
rect 6740 17735 32890 17740
rect 2070 17725 32890 17735
rect -38770 9640 9100 9650
rect -38770 9630 -80 9640
rect -38770 9595 -38755 9630
rect -38720 9595 -38710 9630
rect -38675 9595 -38665 9630
rect -38630 9595 -38620 9630
rect -38585 9595 -38575 9630
rect -38540 9595 -38530 9630
rect -38495 9595 -38485 9630
rect -38450 9595 -38440 9630
rect -38405 9595 -38395 9630
rect -38360 9595 -38350 9630
rect -38315 9595 -38305 9630
rect -38270 9595 -38260 9630
rect -38225 9595 -38215 9630
rect -38180 9595 -38170 9630
rect -38135 9595 -38125 9630
rect -38090 9595 -38080 9630
rect -38045 9595 -38035 9630
rect -38000 9595 -37990 9630
rect -37955 9595 -37945 9630
rect -37910 9595 -37900 9630
rect -37865 9595 -37855 9630
rect -37820 9595 -37810 9630
rect -37775 9595 -37765 9630
rect -37730 9595 -37720 9630
rect -37685 9595 -37675 9630
rect -37640 9595 -37630 9630
rect -37595 9595 -37585 9630
rect -37550 9595 -37540 9630
rect -37505 9595 -37495 9630
rect -37460 9595 -37450 9630
rect -37415 9595 -37405 9630
rect -37370 9595 -37360 9630
rect -37325 9595 -37315 9630
rect -37280 9595 -37270 9630
rect -37235 9595 -37225 9630
rect -37190 9600 -80 9630
rect -40 9600 270 9640
rect 310 9600 620 9640
rect 660 9600 970 9640
rect 1010 9600 1670 9640
rect 1710 9600 2245 9640
rect 2285 9600 3175 9640
rect 3215 9600 3235 9640
rect 3275 9600 3345 9640
rect 3385 9600 6700 9640
rect 6740 9600 7270 9640
rect 7310 9600 7970 9640
rect 8010 9600 8320 9640
rect 8360 9600 8670 9640
rect 8710 9600 9020 9640
rect 9060 9600 9100 9640
rect -37190 9595 9100 9600
rect -38770 9585 9100 9595
rect -38770 9550 -38755 9585
rect -38720 9550 -38710 9585
rect -38675 9550 -38665 9585
rect -38630 9550 -38620 9585
rect -38585 9550 -38575 9585
rect -38540 9550 -38530 9585
rect -38495 9550 -38485 9585
rect -38450 9550 -38440 9585
rect -38405 9550 -38395 9585
rect -38360 9550 -38350 9585
rect -38315 9550 -38305 9585
rect -38270 9550 -38260 9585
rect -38225 9550 -38215 9585
rect -38180 9550 -38170 9585
rect -38135 9550 -38125 9585
rect -38090 9550 -38080 9585
rect -38045 9550 -38035 9585
rect -38000 9550 -37990 9585
rect -37955 9550 -37945 9585
rect -37910 9550 -37900 9585
rect -37865 9550 -37855 9585
rect -37820 9550 -37810 9585
rect -37775 9550 -37765 9585
rect -37730 9550 -37720 9585
rect -37685 9550 -37675 9585
rect -37640 9550 -37630 9585
rect -37595 9550 -37585 9585
rect -37550 9550 -37540 9585
rect -37505 9550 -37495 9585
rect -37460 9550 -37450 9585
rect -37415 9550 -37405 9585
rect -37370 9550 -37360 9585
rect -37325 9550 -37315 9585
rect -37280 9550 -37270 9585
rect -37235 9550 -37225 9585
rect -37190 9575 9100 9585
rect -37190 9550 -80 9575
rect -38770 9540 -80 9550
rect -38770 9505 -38755 9540
rect -38720 9505 -38710 9540
rect -38675 9505 -38665 9540
rect -38630 9505 -38620 9540
rect -38585 9505 -38575 9540
rect -38540 9505 -38530 9540
rect -38495 9505 -38485 9540
rect -38450 9505 -38440 9540
rect -38405 9505 -38395 9540
rect -38360 9505 -38350 9540
rect -38315 9505 -38305 9540
rect -38270 9505 -38260 9540
rect -38225 9505 -38215 9540
rect -38180 9505 -38170 9540
rect -38135 9505 -38125 9540
rect -38090 9505 -38080 9540
rect -38045 9505 -38035 9540
rect -38000 9505 -37990 9540
rect -37955 9505 -37945 9540
rect -37910 9505 -37900 9540
rect -37865 9505 -37855 9540
rect -37820 9505 -37810 9540
rect -37775 9505 -37765 9540
rect -37730 9505 -37720 9540
rect -37685 9505 -37675 9540
rect -37640 9505 -37630 9540
rect -37595 9505 -37585 9540
rect -37550 9505 -37540 9540
rect -37505 9505 -37495 9540
rect -37460 9505 -37450 9540
rect -37415 9505 -37405 9540
rect -37370 9505 -37360 9540
rect -37325 9505 -37315 9540
rect -37280 9505 -37270 9540
rect -37235 9505 -37225 9540
rect -37190 9535 -80 9540
rect -40 9535 270 9575
rect 310 9535 620 9575
rect 660 9535 970 9575
rect 1010 9535 1670 9575
rect 1710 9535 2245 9575
rect 2285 9535 3175 9575
rect 3215 9535 3235 9575
rect 3275 9535 3345 9575
rect 3385 9535 6700 9575
rect 6740 9535 7270 9575
rect 7310 9535 7970 9575
rect 8010 9535 8320 9575
rect 8360 9535 8670 9575
rect 8710 9535 9020 9575
rect 9060 9535 9100 9575
rect -37190 9505 9100 9535
rect -38770 9495 -80 9505
rect -38770 9460 -38755 9495
rect -38720 9460 -38710 9495
rect -38675 9460 -38665 9495
rect -38630 9460 -38620 9495
rect -38585 9460 -38575 9495
rect -38540 9460 -38530 9495
rect -38495 9460 -38485 9495
rect -38450 9460 -38440 9495
rect -38405 9460 -38395 9495
rect -38360 9460 -38350 9495
rect -38315 9460 -38305 9495
rect -38270 9460 -38260 9495
rect -38225 9460 -38215 9495
rect -38180 9460 -38170 9495
rect -38135 9460 -38125 9495
rect -38090 9460 -38080 9495
rect -38045 9460 -38035 9495
rect -38000 9460 -37990 9495
rect -37955 9460 -37945 9495
rect -37910 9460 -37900 9495
rect -37865 9460 -37855 9495
rect -37820 9460 -37810 9495
rect -37775 9460 -37765 9495
rect -37730 9460 -37720 9495
rect -37685 9460 -37675 9495
rect -37640 9460 -37630 9495
rect -37595 9460 -37585 9495
rect -37550 9460 -37540 9495
rect -37505 9460 -37495 9495
rect -37460 9460 -37450 9495
rect -37415 9460 -37405 9495
rect -37370 9460 -37360 9495
rect -37325 9460 -37315 9495
rect -37280 9460 -37270 9495
rect -37235 9460 -37225 9495
rect -37190 9465 -80 9495
rect -40 9465 270 9505
rect 310 9465 620 9505
rect 660 9465 970 9505
rect 1010 9465 1670 9505
rect 1710 9465 2245 9505
rect 2285 9465 3175 9505
rect 3215 9465 3235 9505
rect 3275 9465 3345 9505
rect 3385 9465 6700 9505
rect 6740 9465 7270 9505
rect 7310 9465 7970 9505
rect 8010 9465 8320 9505
rect 8360 9465 8670 9505
rect 8710 9465 9020 9505
rect 9060 9465 9100 9505
rect -37190 9460 9100 9465
rect -38770 9450 9100 9460
rect -38770 9415 -38755 9450
rect -38720 9415 -38710 9450
rect -38675 9415 -38665 9450
rect -38630 9415 -38620 9450
rect -38585 9415 -38575 9450
rect -38540 9415 -38530 9450
rect -38495 9415 -38485 9450
rect -38450 9415 -38440 9450
rect -38405 9415 -38395 9450
rect -38360 9415 -38350 9450
rect -38315 9415 -38305 9450
rect -38270 9415 -38260 9450
rect -38225 9415 -38215 9450
rect -38180 9415 -38170 9450
rect -38135 9415 -38125 9450
rect -38090 9415 -38080 9450
rect -38045 9415 -38035 9450
rect -38000 9415 -37990 9450
rect -37955 9415 -37945 9450
rect -37910 9415 -37900 9450
rect -37865 9415 -37855 9450
rect -37820 9415 -37810 9450
rect -37775 9415 -37765 9450
rect -37730 9415 -37720 9450
rect -37685 9415 -37675 9450
rect -37640 9415 -37630 9450
rect -37595 9415 -37585 9450
rect -37550 9415 -37540 9450
rect -37505 9415 -37495 9450
rect -37460 9415 -37450 9450
rect -37415 9415 -37405 9450
rect -37370 9415 -37360 9450
rect -37325 9415 -37315 9450
rect -37280 9415 -37270 9450
rect -37235 9415 -37225 9450
rect -37190 9435 9100 9450
rect -37190 9415 -80 9435
rect -38770 9405 -80 9415
rect -38770 9370 -38755 9405
rect -38720 9370 -38710 9405
rect -38675 9370 -38665 9405
rect -38630 9370 -38620 9405
rect -38585 9370 -38575 9405
rect -38540 9370 -38530 9405
rect -38495 9370 -38485 9405
rect -38450 9370 -38440 9405
rect -38405 9370 -38395 9405
rect -38360 9370 -38350 9405
rect -38315 9370 -38305 9405
rect -38270 9370 -38260 9405
rect -38225 9370 -38215 9405
rect -38180 9370 -38170 9405
rect -38135 9370 -38125 9405
rect -38090 9370 -38080 9405
rect -38045 9370 -38035 9405
rect -38000 9370 -37990 9405
rect -37955 9370 -37945 9405
rect -37910 9370 -37900 9405
rect -37865 9370 -37855 9405
rect -37820 9370 -37810 9405
rect -37775 9370 -37765 9405
rect -37730 9370 -37720 9405
rect -37685 9370 -37675 9405
rect -37640 9370 -37630 9405
rect -37595 9370 -37585 9405
rect -37550 9370 -37540 9405
rect -37505 9370 -37495 9405
rect -37460 9370 -37450 9405
rect -37415 9370 -37405 9405
rect -37370 9370 -37360 9405
rect -37325 9370 -37315 9405
rect -37280 9370 -37270 9405
rect -37235 9370 -37225 9405
rect -37190 9395 -80 9405
rect -40 9395 270 9435
rect 310 9395 620 9435
rect 660 9395 970 9435
rect 1010 9395 1670 9435
rect 1710 9395 2245 9435
rect 2285 9395 3175 9435
rect 3215 9395 3235 9435
rect 3275 9395 3345 9435
rect 3385 9395 6700 9435
rect 6740 9395 7270 9435
rect 7310 9395 7970 9435
rect 8010 9395 8320 9435
rect 8360 9395 8670 9435
rect 8710 9395 9020 9435
rect 9060 9395 9100 9435
rect -37190 9370 9100 9395
rect -38770 9365 9100 9370
rect -38770 9360 -80 9365
rect -38770 9325 -38755 9360
rect -38720 9325 -38710 9360
rect -38675 9325 -38665 9360
rect -38630 9325 -38620 9360
rect -38585 9325 -38575 9360
rect -38540 9325 -38530 9360
rect -38495 9325 -38485 9360
rect -38450 9325 -38440 9360
rect -38405 9325 -38395 9360
rect -38360 9325 -38350 9360
rect -38315 9325 -38305 9360
rect -38270 9325 -38260 9360
rect -38225 9325 -38215 9360
rect -38180 9325 -38170 9360
rect -38135 9325 -38125 9360
rect -38090 9325 -38080 9360
rect -38045 9325 -38035 9360
rect -38000 9325 -37990 9360
rect -37955 9325 -37945 9360
rect -37910 9325 -37900 9360
rect -37865 9325 -37855 9360
rect -37820 9325 -37810 9360
rect -37775 9325 -37765 9360
rect -37730 9325 -37720 9360
rect -37685 9325 -37675 9360
rect -37640 9325 -37630 9360
rect -37595 9325 -37585 9360
rect -37550 9325 -37540 9360
rect -37505 9325 -37495 9360
rect -37460 9325 -37450 9360
rect -37415 9325 -37405 9360
rect -37370 9325 -37360 9360
rect -37325 9325 -37315 9360
rect -37280 9325 -37270 9360
rect -37235 9325 -37225 9360
rect -37190 9325 -80 9360
rect -40 9325 270 9365
rect 310 9325 620 9365
rect 660 9325 970 9365
rect 1010 9325 1670 9365
rect 1710 9325 2245 9365
rect 2285 9325 3175 9365
rect 3215 9325 3235 9365
rect 3275 9325 3345 9365
rect 3385 9325 6700 9365
rect 6740 9325 7270 9365
rect 7310 9325 7970 9365
rect 8010 9325 8320 9365
rect 8360 9325 8670 9365
rect 8710 9325 9020 9365
rect 9060 9325 9100 9365
rect -38770 9315 9100 9325
rect -38770 9280 -38755 9315
rect -38720 9280 -38710 9315
rect -38675 9280 -38665 9315
rect -38630 9280 -38620 9315
rect -38585 9280 -38575 9315
rect -38540 9280 -38530 9315
rect -38495 9280 -38485 9315
rect -38450 9280 -38440 9315
rect -38405 9280 -38395 9315
rect -38360 9280 -38350 9315
rect -38315 9280 -38305 9315
rect -38270 9280 -38260 9315
rect -38225 9280 -38215 9315
rect -38180 9280 -38170 9315
rect -38135 9280 -38125 9315
rect -38090 9280 -38080 9315
rect -38045 9280 -38035 9315
rect -38000 9280 -37990 9315
rect -37955 9280 -37945 9315
rect -37910 9280 -37900 9315
rect -37865 9280 -37855 9315
rect -37820 9280 -37810 9315
rect -37775 9280 -37765 9315
rect -37730 9280 -37720 9315
rect -37685 9280 -37675 9315
rect -37640 9280 -37630 9315
rect -37595 9280 -37585 9315
rect -37550 9280 -37540 9315
rect -37505 9280 -37495 9315
rect -37460 9280 -37450 9315
rect -37415 9280 -37405 9315
rect -37370 9280 -37360 9315
rect -37325 9280 -37315 9315
rect -37280 9280 -37270 9315
rect -37235 9280 -37225 9315
rect -37190 9300 9100 9315
rect -37190 9280 -80 9300
rect -38770 9270 -80 9280
rect -38770 9235 -38755 9270
rect -38720 9235 -38710 9270
rect -38675 9235 -38665 9270
rect -38630 9235 -38620 9270
rect -38585 9235 -38575 9270
rect -38540 9235 -38530 9270
rect -38495 9235 -38485 9270
rect -38450 9235 -38440 9270
rect -38405 9235 -38395 9270
rect -38360 9235 -38350 9270
rect -38315 9235 -38305 9270
rect -38270 9235 -38260 9270
rect -38225 9235 -38215 9270
rect -38180 9235 -38170 9270
rect -38135 9235 -38125 9270
rect -38090 9235 -38080 9270
rect -38045 9235 -38035 9270
rect -38000 9235 -37990 9270
rect -37955 9235 -37945 9270
rect -37910 9235 -37900 9270
rect -37865 9235 -37855 9270
rect -37820 9235 -37810 9270
rect -37775 9235 -37765 9270
rect -37730 9235 -37720 9270
rect -37685 9235 -37675 9270
rect -37640 9235 -37630 9270
rect -37595 9235 -37585 9270
rect -37550 9235 -37540 9270
rect -37505 9235 -37495 9270
rect -37460 9235 -37450 9270
rect -37415 9235 -37405 9270
rect -37370 9235 -37360 9270
rect -37325 9235 -37315 9270
rect -37280 9235 -37270 9270
rect -37235 9235 -37225 9270
rect -37190 9260 -80 9270
rect -40 9260 270 9300
rect 310 9260 620 9300
rect 660 9260 970 9300
rect 1010 9260 1670 9300
rect 1710 9260 2245 9300
rect 2285 9260 3175 9300
rect 3215 9260 3235 9300
rect 3275 9260 3345 9300
rect 3385 9260 6700 9300
rect 6740 9260 7270 9300
rect 7310 9260 7970 9300
rect 8010 9260 8320 9300
rect 8360 9260 8670 9300
rect 8710 9260 9020 9300
rect 9060 9260 9100 9300
rect -37190 9240 9100 9260
rect -37190 9235 -80 9240
rect -38770 9225 -80 9235
rect -38770 9190 -38755 9225
rect -38720 9190 -38710 9225
rect -38675 9190 -38665 9225
rect -38630 9190 -38620 9225
rect -38585 9190 -38575 9225
rect -38540 9190 -38530 9225
rect -38495 9190 -38485 9225
rect -38450 9190 -38440 9225
rect -38405 9190 -38395 9225
rect -38360 9190 -38350 9225
rect -38315 9190 -38305 9225
rect -38270 9190 -38260 9225
rect -38225 9190 -38215 9225
rect -38180 9190 -38170 9225
rect -38135 9190 -38125 9225
rect -38090 9190 -38080 9225
rect -38045 9190 -38035 9225
rect -38000 9190 -37990 9225
rect -37955 9190 -37945 9225
rect -37910 9190 -37900 9225
rect -37865 9190 -37855 9225
rect -37820 9190 -37810 9225
rect -37775 9190 -37765 9225
rect -37730 9190 -37720 9225
rect -37685 9190 -37675 9225
rect -37640 9190 -37630 9225
rect -37595 9190 -37585 9225
rect -37550 9190 -37540 9225
rect -37505 9190 -37495 9225
rect -37460 9190 -37450 9225
rect -37415 9190 -37405 9225
rect -37370 9190 -37360 9225
rect -37325 9190 -37315 9225
rect -37280 9190 -37270 9225
rect -37235 9190 -37225 9225
rect -37190 9200 -80 9225
rect -40 9200 270 9240
rect 310 9200 620 9240
rect 660 9200 970 9240
rect 1010 9200 1670 9240
rect 1710 9200 2245 9240
rect 2285 9200 3175 9240
rect 3215 9200 3235 9240
rect 3275 9200 3345 9240
rect 3385 9200 6700 9240
rect 6740 9200 7270 9240
rect 7310 9200 7970 9240
rect 8010 9200 8320 9240
rect 8360 9200 8670 9240
rect 8710 9200 9020 9240
rect 9060 9200 9100 9240
rect -37190 9190 9100 9200
rect -38770 9180 9100 9190
rect -38770 9145 -38755 9180
rect -38720 9145 -38710 9180
rect -38675 9145 -38665 9180
rect -38630 9145 -38620 9180
rect -38585 9145 -38575 9180
rect -38540 9145 -38530 9180
rect -38495 9145 -38485 9180
rect -38450 9145 -38440 9180
rect -38405 9145 -38395 9180
rect -38360 9145 -38350 9180
rect -38315 9145 -38305 9180
rect -38270 9145 -38260 9180
rect -38225 9145 -38215 9180
rect -38180 9145 -38170 9180
rect -38135 9145 -38125 9180
rect -38090 9145 -38080 9180
rect -38045 9145 -38035 9180
rect -38000 9145 -37990 9180
rect -37955 9145 -37945 9180
rect -37910 9145 -37900 9180
rect -37865 9145 -37855 9180
rect -37820 9145 -37810 9180
rect -37775 9145 -37765 9180
rect -37730 9145 -37720 9180
rect -37685 9145 -37675 9180
rect -37640 9145 -37630 9180
rect -37595 9145 -37585 9180
rect -37550 9145 -37540 9180
rect -37505 9145 -37495 9180
rect -37460 9145 -37450 9180
rect -37415 9145 -37405 9180
rect -37370 9145 -37360 9180
rect -37325 9145 -37315 9180
rect -37280 9145 -37270 9180
rect -37235 9145 -37225 9180
rect -37190 9175 9100 9180
rect -37190 9145 -80 9175
rect -38770 9135 -80 9145
rect -40 9135 270 9175
rect 310 9135 620 9175
rect 660 9135 970 9175
rect 1010 9135 1670 9175
rect 1710 9135 2245 9175
rect 2285 9135 3175 9175
rect 3215 9135 3235 9175
rect 3275 9135 3345 9175
rect 3385 9135 6700 9175
rect 6740 9135 7270 9175
rect 7310 9135 7970 9175
rect 8010 9135 8320 9175
rect 8360 9135 8670 9175
rect 8710 9135 9020 9175
rect 9060 9135 9100 9175
rect -38770 9100 -38755 9135
rect -38720 9100 -38710 9135
rect -38675 9100 -38665 9135
rect -38630 9100 -38620 9135
rect -38585 9100 -38575 9135
rect -38540 9100 -38530 9135
rect -38495 9100 -38485 9135
rect -38450 9100 -38440 9135
rect -38405 9100 -38395 9135
rect -38360 9100 -38350 9135
rect -38315 9100 -38305 9135
rect -38270 9100 -38260 9135
rect -38225 9100 -38215 9135
rect -38180 9100 -38170 9135
rect -38135 9100 -38125 9135
rect -38090 9100 -38080 9135
rect -38045 9100 -38035 9135
rect -38000 9100 -37990 9135
rect -37955 9100 -37945 9135
rect -37910 9100 -37900 9135
rect -37865 9100 -37855 9135
rect -37820 9100 -37810 9135
rect -37775 9100 -37765 9135
rect -37730 9100 -37720 9135
rect -37685 9100 -37675 9135
rect -37640 9100 -37630 9135
rect -37595 9100 -37585 9135
rect -37550 9100 -37540 9135
rect -37505 9100 -37495 9135
rect -37460 9100 -37450 9135
rect -37415 9100 -37405 9135
rect -37370 9100 -37360 9135
rect -37325 9100 -37315 9135
rect -37280 9100 -37270 9135
rect -37235 9100 -37225 9135
rect -37190 9105 9100 9135
rect -37190 9100 -80 9105
rect -38770 9090 -80 9100
rect -38770 9055 -38755 9090
rect -38720 9055 -38710 9090
rect -38675 9055 -38665 9090
rect -38630 9055 -38620 9090
rect -38585 9055 -38575 9090
rect -38540 9055 -38530 9090
rect -38495 9055 -38485 9090
rect -38450 9055 -38440 9090
rect -38405 9055 -38395 9090
rect -38360 9055 -38350 9090
rect -38315 9055 -38305 9090
rect -38270 9055 -38260 9090
rect -38225 9055 -38215 9090
rect -38180 9055 -38170 9090
rect -38135 9055 -38125 9090
rect -38090 9055 -38080 9090
rect -38045 9055 -38035 9090
rect -38000 9055 -37990 9090
rect -37955 9055 -37945 9090
rect -37910 9055 -37900 9090
rect -37865 9055 -37855 9090
rect -37820 9055 -37810 9090
rect -37775 9055 -37765 9090
rect -37730 9055 -37720 9090
rect -37685 9055 -37675 9090
rect -37640 9055 -37630 9090
rect -37595 9055 -37585 9090
rect -37550 9055 -37540 9090
rect -37505 9055 -37495 9090
rect -37460 9055 -37450 9090
rect -37415 9055 -37405 9090
rect -37370 9055 -37360 9090
rect -37325 9055 -37315 9090
rect -37280 9055 -37270 9090
rect -37235 9055 -37225 9090
rect -37190 9065 -80 9090
rect -40 9065 270 9105
rect 310 9065 620 9105
rect 660 9065 970 9105
rect 1010 9065 1670 9105
rect 1710 9065 2245 9105
rect 2285 9065 3175 9105
rect 3215 9065 3235 9105
rect 3275 9065 3345 9105
rect 3385 9065 6700 9105
rect 6740 9065 7270 9105
rect 7310 9065 7970 9105
rect 8010 9065 8320 9105
rect 8360 9065 8670 9105
rect 8710 9065 9020 9105
rect 9060 9065 9100 9105
rect -37190 9055 9100 9065
rect -38770 9045 9100 9055
rect -38770 9010 -38755 9045
rect -38720 9010 -38710 9045
rect -38675 9010 -38665 9045
rect -38630 9010 -38620 9045
rect -38585 9010 -38575 9045
rect -38540 9010 -38530 9045
rect -38495 9010 -38485 9045
rect -38450 9010 -38440 9045
rect -38405 9010 -38395 9045
rect -38360 9010 -38350 9045
rect -38315 9010 -38305 9045
rect -38270 9010 -38260 9045
rect -38225 9010 -38215 9045
rect -38180 9010 -38170 9045
rect -38135 9010 -38125 9045
rect -38090 9010 -38080 9045
rect -38045 9010 -38035 9045
rect -38000 9010 -37990 9045
rect -37955 9010 -37945 9045
rect -37910 9010 -37900 9045
rect -37865 9010 -37855 9045
rect -37820 9010 -37810 9045
rect -37775 9010 -37765 9045
rect -37730 9010 -37720 9045
rect -37685 9010 -37675 9045
rect -37640 9010 -37630 9045
rect -37595 9010 -37585 9045
rect -37550 9010 -37540 9045
rect -37505 9010 -37495 9045
rect -37460 9010 -37450 9045
rect -37415 9010 -37405 9045
rect -37370 9010 -37360 9045
rect -37325 9010 -37315 9045
rect -37280 9010 -37270 9045
rect -37235 9010 -37225 9045
rect -37190 9035 9100 9045
rect -37190 9010 -80 9035
rect -38770 9000 -80 9010
rect -38770 8965 -38755 9000
rect -38720 8965 -38710 9000
rect -38675 8965 -38665 9000
rect -38630 8965 -38620 9000
rect -38585 8965 -38575 9000
rect -38540 8965 -38530 9000
rect -38495 8965 -38485 9000
rect -38450 8965 -38440 9000
rect -38405 8965 -38395 9000
rect -38360 8965 -38350 9000
rect -38315 8965 -38305 9000
rect -38270 8965 -38260 9000
rect -38225 8965 -38215 9000
rect -38180 8965 -38170 9000
rect -38135 8965 -38125 9000
rect -38090 8965 -38080 9000
rect -38045 8965 -38035 9000
rect -38000 8965 -37990 9000
rect -37955 8965 -37945 9000
rect -37910 8965 -37900 9000
rect -37865 8965 -37855 9000
rect -37820 8965 -37810 9000
rect -37775 8965 -37765 9000
rect -37730 8965 -37720 9000
rect -37685 8965 -37675 9000
rect -37640 8965 -37630 9000
rect -37595 8965 -37585 9000
rect -37550 8965 -37540 9000
rect -37505 8965 -37495 9000
rect -37460 8965 -37450 9000
rect -37415 8965 -37405 9000
rect -37370 8965 -37360 9000
rect -37325 8965 -37315 9000
rect -37280 8965 -37270 9000
rect -37235 8965 -37225 9000
rect -37190 8995 -80 9000
rect -40 8995 270 9035
rect 310 8995 620 9035
rect 660 8995 970 9035
rect 1010 8995 1670 9035
rect 1710 8995 2245 9035
rect 2285 8995 3175 9035
rect 3215 8995 3235 9035
rect 3275 8995 3345 9035
rect 3385 8995 6700 9035
rect 6740 8995 7270 9035
rect 7310 8995 7970 9035
rect 8010 8995 8320 9035
rect 8360 8995 8670 9035
rect 8710 8995 9020 9035
rect 9060 8995 9100 9035
rect -37190 8965 9100 8995
rect -38770 8955 -80 8965
rect -38770 8920 -38755 8955
rect -38720 8920 -38710 8955
rect -38675 8920 -38665 8955
rect -38630 8920 -38620 8955
rect -38585 8920 -38575 8955
rect -38540 8920 -38530 8955
rect -38495 8920 -38485 8955
rect -38450 8920 -38440 8955
rect -38405 8920 -38395 8955
rect -38360 8920 -38350 8955
rect -38315 8920 -38305 8955
rect -38270 8920 -38260 8955
rect -38225 8920 -38215 8955
rect -38180 8920 -38170 8955
rect -38135 8920 -38125 8955
rect -38090 8920 -38080 8955
rect -38045 8920 -38035 8955
rect -38000 8920 -37990 8955
rect -37955 8920 -37945 8955
rect -37910 8920 -37900 8955
rect -37865 8920 -37855 8955
rect -37820 8920 -37810 8955
rect -37775 8920 -37765 8955
rect -37730 8920 -37720 8955
rect -37685 8920 -37675 8955
rect -37640 8920 -37630 8955
rect -37595 8920 -37585 8955
rect -37550 8920 -37540 8955
rect -37505 8920 -37495 8955
rect -37460 8920 -37450 8955
rect -37415 8920 -37405 8955
rect -37370 8920 -37360 8955
rect -37325 8920 -37315 8955
rect -37280 8920 -37270 8955
rect -37235 8920 -37225 8955
rect -37190 8925 -80 8955
rect -40 8925 270 8965
rect 310 8925 620 8965
rect 660 8925 970 8965
rect 1010 8925 1670 8965
rect 1710 8925 2245 8965
rect 2285 8925 3175 8965
rect 3215 8925 3235 8965
rect 3275 8925 3345 8965
rect 3385 8925 6700 8965
rect 6740 8925 7270 8965
rect 7310 8925 7970 8965
rect 8010 8925 8320 8965
rect 8360 8925 8670 8965
rect 8710 8925 9020 8965
rect 9060 8925 9100 8965
rect -37190 8920 9100 8925
rect -38770 8910 9100 8920
rect -38770 8875 -38755 8910
rect -38720 8875 -38710 8910
rect -38675 8875 -38665 8910
rect -38630 8875 -38620 8910
rect -38585 8875 -38575 8910
rect -38540 8875 -38530 8910
rect -38495 8875 -38485 8910
rect -38450 8875 -38440 8910
rect -38405 8875 -38395 8910
rect -38360 8875 -38350 8910
rect -38315 8875 -38305 8910
rect -38270 8875 -38260 8910
rect -38225 8875 -38215 8910
rect -38180 8875 -38170 8910
rect -38135 8875 -38125 8910
rect -38090 8875 -38080 8910
rect -38045 8875 -38035 8910
rect -38000 8875 -37990 8910
rect -37955 8875 -37945 8910
rect -37910 8875 -37900 8910
rect -37865 8875 -37855 8910
rect -37820 8875 -37810 8910
rect -37775 8875 -37765 8910
rect -37730 8875 -37720 8910
rect -37685 8875 -37675 8910
rect -37640 8875 -37630 8910
rect -37595 8875 -37585 8910
rect -37550 8875 -37540 8910
rect -37505 8875 -37495 8910
rect -37460 8875 -37450 8910
rect -37415 8875 -37405 8910
rect -37370 8875 -37360 8910
rect -37325 8875 -37315 8910
rect -37280 8875 -37270 8910
rect -37235 8875 -37225 8910
rect -37190 8900 9100 8910
rect -37190 8875 -80 8900
rect -38770 8865 -80 8875
rect -38770 8830 -38755 8865
rect -38720 8830 -38710 8865
rect -38675 8830 -38665 8865
rect -38630 8830 -38620 8865
rect -38585 8830 -38575 8865
rect -38540 8830 -38530 8865
rect -38495 8830 -38485 8865
rect -38450 8830 -38440 8865
rect -38405 8830 -38395 8865
rect -38360 8830 -38350 8865
rect -38315 8830 -38305 8865
rect -38270 8830 -38260 8865
rect -38225 8830 -38215 8865
rect -38180 8830 -38170 8865
rect -38135 8830 -38125 8865
rect -38090 8830 -38080 8865
rect -38045 8830 -38035 8865
rect -38000 8830 -37990 8865
rect -37955 8830 -37945 8865
rect -37910 8830 -37900 8865
rect -37865 8830 -37855 8865
rect -37820 8830 -37810 8865
rect -37775 8830 -37765 8865
rect -37730 8830 -37720 8865
rect -37685 8830 -37675 8865
rect -37640 8830 -37630 8865
rect -37595 8830 -37585 8865
rect -37550 8830 -37540 8865
rect -37505 8830 -37495 8865
rect -37460 8830 -37450 8865
rect -37415 8830 -37405 8865
rect -37370 8830 -37360 8865
rect -37325 8830 -37315 8865
rect -37280 8830 -37270 8865
rect -37235 8830 -37225 8865
rect -37190 8860 -80 8865
rect -40 8860 270 8900
rect 310 8860 620 8900
rect 660 8860 970 8900
rect 1010 8860 1670 8900
rect 1710 8860 2245 8900
rect 2285 8860 3175 8900
rect 3215 8860 3235 8900
rect 3275 8860 3345 8900
rect 3385 8860 6700 8900
rect 6740 8860 7270 8900
rect 7310 8860 7970 8900
rect 8010 8860 8320 8900
rect 8360 8860 8670 8900
rect 8710 8860 9020 8900
rect 9060 8860 9100 8900
rect -37190 8840 9100 8860
rect -37190 8830 -80 8840
rect -38770 8820 -80 8830
rect -38770 8785 -38755 8820
rect -38720 8785 -38710 8820
rect -38675 8785 -38665 8820
rect -38630 8785 -38620 8820
rect -38585 8785 -38575 8820
rect -38540 8785 -38530 8820
rect -38495 8785 -38485 8820
rect -38450 8785 -38440 8820
rect -38405 8785 -38395 8820
rect -38360 8785 -38350 8820
rect -38315 8785 -38305 8820
rect -38270 8785 -38260 8820
rect -38225 8785 -38215 8820
rect -38180 8785 -38170 8820
rect -38135 8785 -38125 8820
rect -38090 8785 -38080 8820
rect -38045 8785 -38035 8820
rect -38000 8785 -37990 8820
rect -37955 8785 -37945 8820
rect -37910 8785 -37900 8820
rect -37865 8785 -37855 8820
rect -37820 8785 -37810 8820
rect -37775 8785 -37765 8820
rect -37730 8785 -37720 8820
rect -37685 8785 -37675 8820
rect -37640 8785 -37630 8820
rect -37595 8785 -37585 8820
rect -37550 8785 -37540 8820
rect -37505 8785 -37495 8820
rect -37460 8785 -37450 8820
rect -37415 8785 -37405 8820
rect -37370 8785 -37360 8820
rect -37325 8785 -37315 8820
rect -37280 8785 -37270 8820
rect -37235 8785 -37225 8820
rect -37190 8800 -80 8820
rect -40 8800 270 8840
rect 310 8800 620 8840
rect 660 8800 970 8840
rect 1010 8800 1670 8840
rect 1710 8800 2245 8840
rect 2285 8800 3175 8840
rect 3215 8800 3235 8840
rect 3275 8800 3345 8840
rect 3385 8800 6700 8840
rect 6740 8800 7270 8840
rect 7310 8800 7970 8840
rect 8010 8800 8320 8840
rect 8360 8800 8670 8840
rect 8710 8800 9020 8840
rect 9060 8800 9100 8840
rect -37190 8785 9100 8800
rect -38770 8775 9100 8785
rect -38770 8740 -38755 8775
rect -38720 8740 -38710 8775
rect -38675 8740 -38665 8775
rect -38630 8740 -38620 8775
rect -38585 8740 -38575 8775
rect -38540 8740 -38530 8775
rect -38495 8740 -38485 8775
rect -38450 8740 -38440 8775
rect -38405 8740 -38395 8775
rect -38360 8740 -38350 8775
rect -38315 8740 -38305 8775
rect -38270 8740 -38260 8775
rect -38225 8740 -38215 8775
rect -38180 8740 -38170 8775
rect -38135 8740 -38125 8775
rect -38090 8740 -38080 8775
rect -38045 8740 -38035 8775
rect -38000 8740 -37990 8775
rect -37955 8740 -37945 8775
rect -37910 8740 -37900 8775
rect -37865 8740 -37855 8775
rect -37820 8740 -37810 8775
rect -37775 8740 -37765 8775
rect -37730 8740 -37720 8775
rect -37685 8740 -37675 8775
rect -37640 8740 -37630 8775
rect -37595 8740 -37585 8775
rect -37550 8740 -37540 8775
rect -37505 8740 -37495 8775
rect -37460 8740 -37450 8775
rect -37415 8740 -37405 8775
rect -37370 8740 -37360 8775
rect -37325 8740 -37315 8775
rect -37280 8740 -37270 8775
rect -37235 8740 -37225 8775
rect -37190 8740 -80 8775
rect -38770 8735 -80 8740
rect -40 8735 270 8775
rect 310 8735 620 8775
rect 660 8735 970 8775
rect 1010 8735 1670 8775
rect 1710 8735 2245 8775
rect 2285 8735 3175 8775
rect 3215 8735 3235 8775
rect 3275 8735 3345 8775
rect 3385 8735 6700 8775
rect 6740 8735 7270 8775
rect 7310 8735 7970 8775
rect 8010 8735 8320 8775
rect 8360 8735 8670 8775
rect 8710 8735 9020 8775
rect 9060 8735 9100 8775
rect -38770 8730 9100 8735
rect -38770 8695 -38755 8730
rect -38720 8695 -38710 8730
rect -38675 8695 -38665 8730
rect -38630 8695 -38620 8730
rect -38585 8695 -38575 8730
rect -38540 8695 -38530 8730
rect -38495 8695 -38485 8730
rect -38450 8695 -38440 8730
rect -38405 8695 -38395 8730
rect -38360 8695 -38350 8730
rect -38315 8695 -38305 8730
rect -38270 8695 -38260 8730
rect -38225 8695 -38215 8730
rect -38180 8695 -38170 8730
rect -38135 8695 -38125 8730
rect -38090 8695 -38080 8730
rect -38045 8695 -38035 8730
rect -38000 8695 -37990 8730
rect -37955 8695 -37945 8730
rect -37910 8695 -37900 8730
rect -37865 8695 -37855 8730
rect -37820 8695 -37810 8730
rect -37775 8695 -37765 8730
rect -37730 8695 -37720 8730
rect -37685 8695 -37675 8730
rect -37640 8695 -37630 8730
rect -37595 8695 -37585 8730
rect -37550 8695 -37540 8730
rect -37505 8695 -37495 8730
rect -37460 8695 -37450 8730
rect -37415 8695 -37405 8730
rect -37370 8695 -37360 8730
rect -37325 8695 -37315 8730
rect -37280 8695 -37270 8730
rect -37235 8695 -37225 8730
rect -37190 8705 9100 8730
rect -37190 8695 -80 8705
rect -38770 8685 -80 8695
rect -38770 8650 -38755 8685
rect -38720 8650 -38710 8685
rect -38675 8650 -38665 8685
rect -38630 8650 -38620 8685
rect -38585 8650 -38575 8685
rect -38540 8650 -38530 8685
rect -38495 8650 -38485 8685
rect -38450 8650 -38440 8685
rect -38405 8650 -38395 8685
rect -38360 8650 -38350 8685
rect -38315 8650 -38305 8685
rect -38270 8650 -38260 8685
rect -38225 8650 -38215 8685
rect -38180 8650 -38170 8685
rect -38135 8650 -38125 8685
rect -38090 8650 -38080 8685
rect -38045 8650 -38035 8685
rect -38000 8650 -37990 8685
rect -37955 8650 -37945 8685
rect -37910 8650 -37900 8685
rect -37865 8650 -37855 8685
rect -37820 8650 -37810 8685
rect -37775 8650 -37765 8685
rect -37730 8650 -37720 8685
rect -37685 8650 -37675 8685
rect -37640 8650 -37630 8685
rect -37595 8650 -37585 8685
rect -37550 8650 -37540 8685
rect -37505 8650 -37495 8685
rect -37460 8650 -37450 8685
rect -37415 8650 -37405 8685
rect -37370 8650 -37360 8685
rect -37325 8650 -37315 8685
rect -37280 8650 -37270 8685
rect -37235 8650 -37225 8685
rect -37190 8665 -80 8685
rect -40 8665 270 8705
rect 310 8665 620 8705
rect 660 8665 970 8705
rect 1010 8665 1670 8705
rect 1710 8665 2245 8705
rect 2285 8665 3175 8705
rect 3215 8665 3235 8705
rect 3275 8665 3345 8705
rect 3385 8665 6700 8705
rect 6740 8665 7270 8705
rect 7310 8665 7970 8705
rect 8010 8665 8320 8705
rect 8360 8665 8670 8705
rect 8710 8665 9020 8705
rect 9060 8665 9100 8705
rect -37190 8650 9100 8665
rect -38770 8640 9100 8650
rect -38770 8605 -38755 8640
rect -38720 8605 -38710 8640
rect -38675 8605 -38665 8640
rect -38630 8605 -38620 8640
rect -38585 8605 -38575 8640
rect -38540 8605 -38530 8640
rect -38495 8605 -38485 8640
rect -38450 8605 -38440 8640
rect -38405 8605 -38395 8640
rect -38360 8605 -38350 8640
rect -38315 8605 -38305 8640
rect -38270 8605 -38260 8640
rect -38225 8605 -38215 8640
rect -38180 8605 -38170 8640
rect -38135 8605 -38125 8640
rect -38090 8605 -38080 8640
rect -38045 8605 -38035 8640
rect -38000 8605 -37990 8640
rect -37955 8605 -37945 8640
rect -37910 8605 -37900 8640
rect -37865 8605 -37855 8640
rect -37820 8605 -37810 8640
rect -37775 8605 -37765 8640
rect -37730 8605 -37720 8640
rect -37685 8605 -37675 8640
rect -37640 8605 -37630 8640
rect -37595 8605 -37585 8640
rect -37550 8605 -37540 8640
rect -37505 8605 -37495 8640
rect -37460 8605 -37450 8640
rect -37415 8605 -37405 8640
rect -37370 8605 -37360 8640
rect -37325 8605 -37315 8640
rect -37280 8605 -37270 8640
rect -37235 8605 -37225 8640
rect -37190 8635 9100 8640
rect -37190 8605 -80 8635
rect -38770 8595 -80 8605
rect -40 8595 270 8635
rect 310 8595 620 8635
rect 660 8595 970 8635
rect 1010 8595 1670 8635
rect 1710 8595 2245 8635
rect 2285 8595 3175 8635
rect 3215 8595 3235 8635
rect 3275 8595 3345 8635
rect 3385 8595 6700 8635
rect 6740 8595 7270 8635
rect 7310 8595 7970 8635
rect 8010 8595 8320 8635
rect 8360 8595 8670 8635
rect 8710 8595 9020 8635
rect 9060 8595 9100 8635
rect -38770 8560 -38755 8595
rect -38720 8560 -38710 8595
rect -38675 8560 -38665 8595
rect -38630 8560 -38620 8595
rect -38585 8560 -38575 8595
rect -38540 8560 -38530 8595
rect -38495 8560 -38485 8595
rect -38450 8560 -38440 8595
rect -38405 8560 -38395 8595
rect -38360 8560 -38350 8595
rect -38315 8560 -38305 8595
rect -38270 8560 -38260 8595
rect -38225 8560 -38215 8595
rect -38180 8560 -38170 8595
rect -38135 8560 -38125 8595
rect -38090 8560 -38080 8595
rect -38045 8560 -38035 8595
rect -38000 8560 -37990 8595
rect -37955 8560 -37945 8595
rect -37910 8560 -37900 8595
rect -37865 8560 -37855 8595
rect -37820 8560 -37810 8595
rect -37775 8560 -37765 8595
rect -37730 8560 -37720 8595
rect -37685 8560 -37675 8595
rect -37640 8560 -37630 8595
rect -37595 8560 -37585 8595
rect -37550 8560 -37540 8595
rect -37505 8560 -37495 8595
rect -37460 8560 -37450 8595
rect -37415 8560 -37405 8595
rect -37370 8560 -37360 8595
rect -37325 8560 -37315 8595
rect -37280 8560 -37270 8595
rect -37235 8560 -37225 8595
rect -37190 8565 9100 8595
rect -37190 8560 -80 8565
rect -38770 8550 -80 8560
rect -38770 8515 -38755 8550
rect -38720 8515 -38710 8550
rect -38675 8515 -38665 8550
rect -38630 8515 -38620 8550
rect -38585 8515 -38575 8550
rect -38540 8515 -38530 8550
rect -38495 8515 -38485 8550
rect -38450 8515 -38440 8550
rect -38405 8515 -38395 8550
rect -38360 8515 -38350 8550
rect -38315 8515 -38305 8550
rect -38270 8515 -38260 8550
rect -38225 8515 -38215 8550
rect -38180 8515 -38170 8550
rect -38135 8515 -38125 8550
rect -38090 8515 -38080 8550
rect -38045 8515 -38035 8550
rect -38000 8515 -37990 8550
rect -37955 8515 -37945 8550
rect -37910 8515 -37900 8550
rect -37865 8515 -37855 8550
rect -37820 8515 -37810 8550
rect -37775 8515 -37765 8550
rect -37730 8515 -37720 8550
rect -37685 8515 -37675 8550
rect -37640 8515 -37630 8550
rect -37595 8515 -37585 8550
rect -37550 8515 -37540 8550
rect -37505 8515 -37495 8550
rect -37460 8515 -37450 8550
rect -37415 8515 -37405 8550
rect -37370 8515 -37360 8550
rect -37325 8515 -37315 8550
rect -37280 8515 -37270 8550
rect -37235 8515 -37225 8550
rect -37190 8525 -80 8550
rect -40 8525 270 8565
rect 310 8525 620 8565
rect 660 8525 970 8565
rect 1010 8525 1670 8565
rect 1710 8525 2245 8565
rect 2285 8525 3175 8565
rect 3215 8525 3235 8565
rect 3275 8525 3345 8565
rect 3385 8525 6700 8565
rect 6740 8525 7270 8565
rect 7310 8525 7970 8565
rect 8010 8525 8320 8565
rect 8360 8525 8670 8565
rect 8710 8525 9020 8565
rect 9060 8525 9100 8565
rect -37190 8515 9100 8525
rect -38770 8505 9100 8515
rect -38770 8470 -38755 8505
rect -38720 8470 -38710 8505
rect -38675 8470 -38665 8505
rect -38630 8470 -38620 8505
rect -38585 8470 -38575 8505
rect -38540 8470 -38530 8505
rect -38495 8470 -38485 8505
rect -38450 8470 -38440 8505
rect -38405 8470 -38395 8505
rect -38360 8470 -38350 8505
rect -38315 8470 -38305 8505
rect -38270 8470 -38260 8505
rect -38225 8470 -38215 8505
rect -38180 8470 -38170 8505
rect -38135 8470 -38125 8505
rect -38090 8470 -38080 8505
rect -38045 8470 -38035 8505
rect -38000 8470 -37990 8505
rect -37955 8470 -37945 8505
rect -37910 8470 -37900 8505
rect -37865 8470 -37855 8505
rect -37820 8470 -37810 8505
rect -37775 8470 -37765 8505
rect -37730 8470 -37720 8505
rect -37685 8470 -37675 8505
rect -37640 8470 -37630 8505
rect -37595 8470 -37585 8505
rect -37550 8470 -37540 8505
rect -37505 8470 -37495 8505
rect -37460 8470 -37450 8505
rect -37415 8470 -37405 8505
rect -37370 8470 -37360 8505
rect -37325 8470 -37315 8505
rect -37280 8470 -37270 8505
rect -37235 8470 -37225 8505
rect -37190 8500 9100 8505
rect -37190 8470 -80 8500
rect -38770 8460 -80 8470
rect -40 8460 270 8500
rect 310 8460 620 8500
rect 660 8460 970 8500
rect 1010 8460 1670 8500
rect 1710 8460 2245 8500
rect 2285 8460 3175 8500
rect 3215 8460 3235 8500
rect 3275 8460 3345 8500
rect 3385 8460 6700 8500
rect 6740 8460 7270 8500
rect 7310 8460 7970 8500
rect 8010 8460 8320 8500
rect 8360 8460 8670 8500
rect 8710 8460 9020 8500
rect 9060 8460 9100 8500
rect -38770 8425 -38755 8460
rect -38720 8425 -38710 8460
rect -38675 8425 -38665 8460
rect -38630 8425 -38620 8460
rect -38585 8425 -38575 8460
rect -38540 8425 -38530 8460
rect -38495 8425 -38485 8460
rect -38450 8425 -38440 8460
rect -38405 8425 -38395 8460
rect -38360 8425 -38350 8460
rect -38315 8425 -38305 8460
rect -38270 8425 -38260 8460
rect -38225 8425 -38215 8460
rect -38180 8425 -38170 8460
rect -38135 8425 -38125 8460
rect -38090 8425 -38080 8460
rect -38045 8425 -38035 8460
rect -38000 8425 -37990 8460
rect -37955 8425 -37945 8460
rect -37910 8425 -37900 8460
rect -37865 8425 -37855 8460
rect -37820 8425 -37810 8460
rect -37775 8425 -37765 8460
rect -37730 8425 -37720 8460
rect -37685 8425 -37675 8460
rect -37640 8425 -37630 8460
rect -37595 8425 -37585 8460
rect -37550 8425 -37540 8460
rect -37505 8425 -37495 8460
rect -37460 8425 -37450 8460
rect -37415 8425 -37405 8460
rect -37370 8425 -37360 8460
rect -37325 8425 -37315 8460
rect -37280 8425 -37270 8460
rect -37235 8425 -37225 8460
rect -37190 8440 9100 8460
rect -37190 8425 -80 8440
rect -38770 8415 -80 8425
rect -38770 8380 -38755 8415
rect -38720 8380 -38710 8415
rect -38675 8380 -38665 8415
rect -38630 8380 -38620 8415
rect -38585 8380 -38575 8415
rect -38540 8380 -38530 8415
rect -38495 8380 -38485 8415
rect -38450 8380 -38440 8415
rect -38405 8380 -38395 8415
rect -38360 8380 -38350 8415
rect -38315 8380 -38305 8415
rect -38270 8380 -38260 8415
rect -38225 8380 -38215 8415
rect -38180 8380 -38170 8415
rect -38135 8380 -38125 8415
rect -38090 8380 -38080 8415
rect -38045 8380 -38035 8415
rect -38000 8380 -37990 8415
rect -37955 8380 -37945 8415
rect -37910 8380 -37900 8415
rect -37865 8380 -37855 8415
rect -37820 8380 -37810 8415
rect -37775 8380 -37765 8415
rect -37730 8380 -37720 8415
rect -37685 8380 -37675 8415
rect -37640 8380 -37630 8415
rect -37595 8380 -37585 8415
rect -37550 8380 -37540 8415
rect -37505 8380 -37495 8415
rect -37460 8380 -37450 8415
rect -37415 8380 -37405 8415
rect -37370 8380 -37360 8415
rect -37325 8380 -37315 8415
rect -37280 8380 -37270 8415
rect -37235 8380 -37225 8415
rect -37190 8400 -80 8415
rect -40 8400 270 8440
rect 310 8400 620 8440
rect 660 8400 970 8440
rect 1010 8400 1670 8440
rect 1710 8400 2245 8440
rect 2285 8400 3175 8440
rect 3215 8400 3235 8440
rect 3275 8400 3345 8440
rect 3385 8400 6700 8440
rect 6740 8400 7270 8440
rect 7310 8400 7970 8440
rect 8010 8400 8320 8440
rect 8360 8400 8670 8440
rect 8710 8400 9020 8440
rect 9060 8400 9100 8440
rect -37190 8380 9100 8400
rect -38770 8375 9100 8380
rect -38770 8370 -80 8375
rect -38770 8335 -38755 8370
rect -38720 8335 -38710 8370
rect -38675 8335 -38665 8370
rect -38630 8335 -38620 8370
rect -38585 8335 -38575 8370
rect -38540 8335 -38530 8370
rect -38495 8335 -38485 8370
rect -38450 8335 -38440 8370
rect -38405 8335 -38395 8370
rect -38360 8335 -38350 8370
rect -38315 8335 -38305 8370
rect -38270 8335 -38260 8370
rect -38225 8335 -38215 8370
rect -38180 8335 -38170 8370
rect -38135 8335 -38125 8370
rect -38090 8335 -38080 8370
rect -38045 8335 -38035 8370
rect -38000 8335 -37990 8370
rect -37955 8335 -37945 8370
rect -37910 8335 -37900 8370
rect -37865 8335 -37855 8370
rect -37820 8335 -37810 8370
rect -37775 8335 -37765 8370
rect -37730 8335 -37720 8370
rect -37685 8335 -37675 8370
rect -37640 8335 -37630 8370
rect -37595 8335 -37585 8370
rect -37550 8335 -37540 8370
rect -37505 8335 -37495 8370
rect -37460 8335 -37450 8370
rect -37415 8335 -37405 8370
rect -37370 8335 -37360 8370
rect -37325 8335 -37315 8370
rect -37280 8335 -37270 8370
rect -37235 8335 -37225 8370
rect -37190 8335 -80 8370
rect -40 8335 270 8375
rect 310 8335 620 8375
rect 660 8335 970 8375
rect 1010 8335 1670 8375
rect 1710 8335 2245 8375
rect 2285 8335 3175 8375
rect 3215 8335 3235 8375
rect 3275 8335 3345 8375
rect 3385 8335 6700 8375
rect 6740 8335 7270 8375
rect 7310 8335 7970 8375
rect 8010 8335 8320 8375
rect 8360 8335 8670 8375
rect 8710 8335 9020 8375
rect 9060 8335 9100 8375
rect -38770 8325 9100 8335
rect -38770 8290 -38755 8325
rect -38720 8290 -38710 8325
rect -38675 8290 -38665 8325
rect -38630 8290 -38620 8325
rect -38585 8290 -38575 8325
rect -38540 8290 -38530 8325
rect -38495 8290 -38485 8325
rect -38450 8290 -38440 8325
rect -38405 8290 -38395 8325
rect -38360 8290 -38350 8325
rect -38315 8290 -38305 8325
rect -38270 8290 -38260 8325
rect -38225 8290 -38215 8325
rect -38180 8290 -38170 8325
rect -38135 8290 -38125 8325
rect -38090 8290 -38080 8325
rect -38045 8290 -38035 8325
rect -38000 8290 -37990 8325
rect -37955 8290 -37945 8325
rect -37910 8290 -37900 8325
rect -37865 8290 -37855 8325
rect -37820 8290 -37810 8325
rect -37775 8290 -37765 8325
rect -37730 8290 -37720 8325
rect -37685 8290 -37675 8325
rect -37640 8290 -37630 8325
rect -37595 8290 -37585 8325
rect -37550 8290 -37540 8325
rect -37505 8290 -37495 8325
rect -37460 8290 -37450 8325
rect -37415 8290 -37405 8325
rect -37370 8290 -37360 8325
rect -37325 8290 -37315 8325
rect -37280 8290 -37270 8325
rect -37235 8290 -37225 8325
rect -37190 8305 9100 8325
rect -37190 8290 -80 8305
rect -38770 8280 -80 8290
rect -38770 8245 -38755 8280
rect -38720 8245 -38710 8280
rect -38675 8245 -38665 8280
rect -38630 8245 -38620 8280
rect -38585 8245 -38575 8280
rect -38540 8245 -38530 8280
rect -38495 8245 -38485 8280
rect -38450 8245 -38440 8280
rect -38405 8245 -38395 8280
rect -38360 8245 -38350 8280
rect -38315 8245 -38305 8280
rect -38270 8245 -38260 8280
rect -38225 8245 -38215 8280
rect -38180 8245 -38170 8280
rect -38135 8245 -38125 8280
rect -38090 8245 -38080 8280
rect -38045 8245 -38035 8280
rect -38000 8245 -37990 8280
rect -37955 8245 -37945 8280
rect -37910 8245 -37900 8280
rect -37865 8245 -37855 8280
rect -37820 8245 -37810 8280
rect -37775 8245 -37765 8280
rect -37730 8245 -37720 8280
rect -37685 8245 -37675 8280
rect -37640 8245 -37630 8280
rect -37595 8245 -37585 8280
rect -37550 8245 -37540 8280
rect -37505 8245 -37495 8280
rect -37460 8245 -37450 8280
rect -37415 8245 -37405 8280
rect -37370 8245 -37360 8280
rect -37325 8245 -37315 8280
rect -37280 8245 -37270 8280
rect -37235 8245 -37225 8280
rect -37190 8265 -80 8280
rect -40 8265 270 8305
rect 310 8265 620 8305
rect 660 8265 970 8305
rect 1010 8265 1670 8305
rect 1710 8265 2245 8305
rect 2285 8265 3175 8305
rect 3215 8265 3235 8305
rect 3275 8265 3345 8305
rect 3385 8265 6700 8305
rect 6740 8265 7270 8305
rect 7310 8265 7970 8305
rect 8010 8265 8320 8305
rect 8360 8265 8670 8305
rect 8710 8265 9020 8305
rect 9060 8265 9100 8305
rect -37190 8245 9100 8265
rect -38770 8235 9100 8245
rect -38770 8200 -38755 8235
rect -38720 8200 -38710 8235
rect -38675 8200 -38665 8235
rect -38630 8200 -38620 8235
rect -38585 8200 -38575 8235
rect -38540 8200 -38530 8235
rect -38495 8200 -38485 8235
rect -38450 8200 -38440 8235
rect -38405 8200 -38395 8235
rect -38360 8200 -38350 8235
rect -38315 8200 -38305 8235
rect -38270 8200 -38260 8235
rect -38225 8200 -38215 8235
rect -38180 8200 -38170 8235
rect -38135 8200 -38125 8235
rect -38090 8200 -38080 8235
rect -38045 8200 -38035 8235
rect -38000 8200 -37990 8235
rect -37955 8200 -37945 8235
rect -37910 8200 -37900 8235
rect -37865 8200 -37855 8235
rect -37820 8200 -37810 8235
rect -37775 8200 -37765 8235
rect -37730 8200 -37720 8235
rect -37685 8200 -37675 8235
rect -37640 8200 -37630 8235
rect -37595 8200 -37585 8235
rect -37550 8200 -37540 8235
rect -37505 8200 -37495 8235
rect -37460 8200 -37450 8235
rect -37415 8200 -37405 8235
rect -37370 8200 -37360 8235
rect -37325 8200 -37315 8235
rect -37280 8200 -37270 8235
rect -37235 8200 -37225 8235
rect -37190 8200 -80 8235
rect -38770 8195 -80 8200
rect -40 8195 270 8235
rect 310 8195 620 8235
rect 660 8195 970 8235
rect 1010 8195 1670 8235
rect 1710 8195 2245 8235
rect 2285 8195 3175 8235
rect 3215 8195 3235 8235
rect 3275 8195 3345 8235
rect 3385 8195 6700 8235
rect 6740 8195 7270 8235
rect 7310 8195 7970 8235
rect 8010 8195 8320 8235
rect 8360 8195 8670 8235
rect 8710 8195 9020 8235
rect 9060 8195 9100 8235
rect -38770 8190 9100 8195
rect -38770 8155 -38755 8190
rect -38720 8155 -38710 8190
rect -38675 8155 -38665 8190
rect -38630 8155 -38620 8190
rect -38585 8155 -38575 8190
rect -38540 8155 -38530 8190
rect -38495 8155 -38485 8190
rect -38450 8155 -38440 8190
rect -38405 8155 -38395 8190
rect -38360 8155 -38350 8190
rect -38315 8155 -38305 8190
rect -38270 8155 -38260 8190
rect -38225 8155 -38215 8190
rect -38180 8155 -38170 8190
rect -38135 8155 -38125 8190
rect -38090 8155 -38080 8190
rect -38045 8155 -38035 8190
rect -38000 8155 -37990 8190
rect -37955 8155 -37945 8190
rect -37910 8155 -37900 8190
rect -37865 8155 -37855 8190
rect -37820 8155 -37810 8190
rect -37775 8155 -37765 8190
rect -37730 8155 -37720 8190
rect -37685 8155 -37675 8190
rect -37640 8155 -37630 8190
rect -37595 8155 -37585 8190
rect -37550 8155 -37540 8190
rect -37505 8155 -37495 8190
rect -37460 8155 -37450 8190
rect -37415 8155 -37405 8190
rect -37370 8155 -37360 8190
rect -37325 8155 -37315 8190
rect -37280 8155 -37270 8190
rect -37235 8155 -37225 8190
rect -37190 8165 9100 8190
rect -37190 8155 -80 8165
rect -38770 8145 -80 8155
rect -38770 8110 -38755 8145
rect -38720 8110 -38710 8145
rect -38675 8110 -38665 8145
rect -38630 8110 -38620 8145
rect -38585 8110 -38575 8145
rect -38540 8110 -38530 8145
rect -38495 8110 -38485 8145
rect -38450 8110 -38440 8145
rect -38405 8110 -38395 8145
rect -38360 8110 -38350 8145
rect -38315 8110 -38305 8145
rect -38270 8110 -38260 8145
rect -38225 8110 -38215 8145
rect -38180 8110 -38170 8145
rect -38135 8110 -38125 8145
rect -38090 8110 -38080 8145
rect -38045 8110 -38035 8145
rect -38000 8110 -37990 8145
rect -37955 8110 -37945 8145
rect -37910 8110 -37900 8145
rect -37865 8110 -37855 8145
rect -37820 8110 -37810 8145
rect -37775 8110 -37765 8145
rect -37730 8110 -37720 8145
rect -37685 8110 -37675 8145
rect -37640 8110 -37630 8145
rect -37595 8110 -37585 8145
rect -37550 8110 -37540 8145
rect -37505 8110 -37495 8145
rect -37460 8110 -37450 8145
rect -37415 8110 -37405 8145
rect -37370 8110 -37360 8145
rect -37325 8110 -37315 8145
rect -37280 8110 -37270 8145
rect -37235 8110 -37225 8145
rect -37190 8125 -80 8145
rect -40 8125 270 8165
rect 310 8125 620 8165
rect 660 8125 970 8165
rect 1010 8125 1670 8165
rect 1710 8125 2245 8165
rect 2285 8125 3175 8165
rect 3215 8125 3235 8165
rect 3275 8125 3345 8165
rect 3385 8125 6700 8165
rect 6740 8125 7270 8165
rect 7310 8125 7970 8165
rect 8010 8125 8320 8165
rect 8360 8125 8670 8165
rect 8710 8125 9020 8165
rect 9060 8125 9100 8165
rect -37190 8110 9100 8125
rect -38770 8100 9100 8110
rect -38770 8065 -38755 8100
rect -38720 8065 -38710 8100
rect -38675 8065 -38665 8100
rect -38630 8065 -38620 8100
rect -38585 8065 -38575 8100
rect -38540 8065 -38530 8100
rect -38495 8065 -38485 8100
rect -38450 8065 -38440 8100
rect -38405 8065 -38395 8100
rect -38360 8065 -38350 8100
rect -38315 8065 -38305 8100
rect -38270 8065 -38260 8100
rect -38225 8065 -38215 8100
rect -38180 8065 -38170 8100
rect -38135 8065 -38125 8100
rect -38090 8065 -38080 8100
rect -38045 8065 -38035 8100
rect -38000 8065 -37990 8100
rect -37955 8065 -37945 8100
rect -37910 8065 -37900 8100
rect -37865 8065 -37855 8100
rect -37820 8065 -37810 8100
rect -37775 8065 -37765 8100
rect -37730 8065 -37720 8100
rect -37685 8065 -37675 8100
rect -37640 8065 -37630 8100
rect -37595 8065 -37585 8100
rect -37550 8065 -37540 8100
rect -37505 8065 -37495 8100
rect -37460 8065 -37450 8100
rect -37415 8065 -37405 8100
rect -37370 8065 -37360 8100
rect -37325 8065 -37315 8100
rect -37280 8065 -37270 8100
rect -37235 8065 -37225 8100
rect -37190 8065 -80 8100
rect -38770 8060 -80 8065
rect -40 8060 270 8100
rect 310 8060 620 8100
rect 660 8060 970 8100
rect 1010 8060 1670 8100
rect 1710 8060 2245 8100
rect 2285 8060 3175 8100
rect 3215 8060 3235 8100
rect 3275 8060 3345 8100
rect 3385 8060 6700 8100
rect 6740 8060 7270 8100
rect 7310 8060 7970 8100
rect 8010 8060 8320 8100
rect 8360 8060 8670 8100
rect 8710 8060 9020 8100
rect 9060 8060 9100 8100
rect -38770 8040 9100 8060
rect -38770 8030 -80 8040
rect -38770 7995 -38755 8030
rect -38720 7995 -38710 8030
rect -38675 7995 -38665 8030
rect -38630 7995 -38620 8030
rect -38585 7995 -38575 8030
rect -38540 7995 -38530 8030
rect -38495 7995 -38485 8030
rect -38450 7995 -38440 8030
rect -38405 7995 -38395 8030
rect -38360 7995 -38350 8030
rect -38315 7995 -38305 8030
rect -38270 7995 -38260 8030
rect -38225 7995 -38215 8030
rect -38180 7995 -38170 8030
rect -38135 7995 -38125 8030
rect -38090 7995 -38080 8030
rect -38045 7995 -38035 8030
rect -38000 7995 -37990 8030
rect -37955 7995 -37945 8030
rect -37910 7995 -37900 8030
rect -37865 7995 -37855 8030
rect -37820 7995 -37810 8030
rect -37775 7995 -37765 8030
rect -37730 7995 -37720 8030
rect -37685 7995 -37675 8030
rect -37640 7995 -37630 8030
rect -37595 7995 -37585 8030
rect -37550 7995 -37540 8030
rect -37505 7995 -37495 8030
rect -37460 7995 -37450 8030
rect -37415 7995 -37405 8030
rect -37370 7995 -37360 8030
rect -37325 7995 -37315 8030
rect -37280 7995 -37270 8030
rect -37235 7995 -37225 8030
rect -37190 8000 -80 8030
rect -40 8000 270 8040
rect 310 8000 620 8040
rect 660 8000 970 8040
rect 1010 8000 1670 8040
rect 1710 8000 2245 8040
rect 2285 8000 3175 8040
rect 3215 8000 3235 8040
rect 3275 8000 3345 8040
rect 3385 8000 6700 8040
rect 6740 8000 7270 8040
rect 7310 8000 7970 8040
rect 8010 8000 8320 8040
rect 8360 8000 8670 8040
rect 8710 8000 9020 8040
rect 9060 8000 9100 8040
rect -37190 7995 9100 8000
rect -38770 7985 9100 7995
rect -38770 7950 -38755 7985
rect -38720 7950 -38710 7985
rect -38675 7950 -38665 7985
rect -38630 7950 -38620 7985
rect -38585 7950 -38575 7985
rect -38540 7950 -38530 7985
rect -38495 7950 -38485 7985
rect -38450 7950 -38440 7985
rect -38405 7950 -38395 7985
rect -38360 7950 -38350 7985
rect -38315 7950 -38305 7985
rect -38270 7950 -38260 7985
rect -38225 7950 -38215 7985
rect -38180 7950 -38170 7985
rect -38135 7950 -38125 7985
rect -38090 7950 -38080 7985
rect -38045 7950 -38035 7985
rect -38000 7950 -37990 7985
rect -37955 7950 -37945 7985
rect -37910 7950 -37900 7985
rect -37865 7950 -37855 7985
rect -37820 7950 -37810 7985
rect -37775 7950 -37765 7985
rect -37730 7950 -37720 7985
rect -37685 7950 -37675 7985
rect -37640 7950 -37630 7985
rect -37595 7950 -37585 7985
rect -37550 7950 -37540 7985
rect -37505 7950 -37495 7985
rect -37460 7950 -37450 7985
rect -37415 7950 -37405 7985
rect -37370 7950 -37360 7985
rect -37325 7950 -37315 7985
rect -37280 7950 -37270 7985
rect -37235 7950 -37225 7985
rect -37190 7975 9100 7985
rect -37190 7950 -80 7975
rect -38770 7940 -80 7950
rect -38770 7905 -38755 7940
rect -38720 7905 -38710 7940
rect -38675 7905 -38665 7940
rect -38630 7905 -38620 7940
rect -38585 7905 -38575 7940
rect -38540 7905 -38530 7940
rect -38495 7905 -38485 7940
rect -38450 7905 -38440 7940
rect -38405 7905 -38395 7940
rect -38360 7905 -38350 7940
rect -38315 7905 -38305 7940
rect -38270 7905 -38260 7940
rect -38225 7905 -38215 7940
rect -38180 7905 -38170 7940
rect -38135 7905 -38125 7940
rect -38090 7905 -38080 7940
rect -38045 7905 -38035 7940
rect -38000 7905 -37990 7940
rect -37955 7905 -37945 7940
rect -37910 7905 -37900 7940
rect -37865 7905 -37855 7940
rect -37820 7905 -37810 7940
rect -37775 7905 -37765 7940
rect -37730 7905 -37720 7940
rect -37685 7905 -37675 7940
rect -37640 7905 -37630 7940
rect -37595 7905 -37585 7940
rect -37550 7905 -37540 7940
rect -37505 7905 -37495 7940
rect -37460 7905 -37450 7940
rect -37415 7905 -37405 7940
rect -37370 7905 -37360 7940
rect -37325 7905 -37315 7940
rect -37280 7905 -37270 7940
rect -37235 7905 -37225 7940
rect -37190 7935 -80 7940
rect -40 7935 270 7975
rect 310 7935 620 7975
rect 660 7935 970 7975
rect 1010 7935 1670 7975
rect 1710 7935 2245 7975
rect 2285 7935 3175 7975
rect 3215 7935 3235 7975
rect 3275 7935 3345 7975
rect 3385 7935 6700 7975
rect 6740 7935 7270 7975
rect 7310 7935 7970 7975
rect 8010 7935 8320 7975
rect 8360 7935 8670 7975
rect 8710 7935 9020 7975
rect 9060 7935 9100 7975
rect -37190 7905 9100 7935
rect -38770 7895 -80 7905
rect -38770 7860 -38755 7895
rect -38720 7860 -38710 7895
rect -38675 7860 -38665 7895
rect -38630 7860 -38620 7895
rect -38585 7860 -38575 7895
rect -38540 7860 -38530 7895
rect -38495 7860 -38485 7895
rect -38450 7860 -38440 7895
rect -38405 7860 -38395 7895
rect -38360 7860 -38350 7895
rect -38315 7860 -38305 7895
rect -38270 7860 -38260 7895
rect -38225 7860 -38215 7895
rect -38180 7860 -38170 7895
rect -38135 7860 -38125 7895
rect -38090 7860 -38080 7895
rect -38045 7860 -38035 7895
rect -38000 7860 -37990 7895
rect -37955 7860 -37945 7895
rect -37910 7860 -37900 7895
rect -37865 7860 -37855 7895
rect -37820 7860 -37810 7895
rect -37775 7860 -37765 7895
rect -37730 7860 -37720 7895
rect -37685 7860 -37675 7895
rect -37640 7860 -37630 7895
rect -37595 7860 -37585 7895
rect -37550 7860 -37540 7895
rect -37505 7860 -37495 7895
rect -37460 7860 -37450 7895
rect -37415 7860 -37405 7895
rect -37370 7860 -37360 7895
rect -37325 7860 -37315 7895
rect -37280 7860 -37270 7895
rect -37235 7860 -37225 7895
rect -37190 7865 -80 7895
rect -40 7865 270 7905
rect 310 7865 620 7905
rect 660 7865 970 7905
rect 1010 7865 1670 7905
rect 1710 7865 2245 7905
rect 2285 7865 3175 7905
rect 3215 7865 3235 7905
rect 3275 7865 3345 7905
rect 3385 7865 6700 7905
rect 6740 7865 7270 7905
rect 7310 7865 7970 7905
rect 8010 7865 8320 7905
rect 8360 7865 8670 7905
rect 8710 7865 9020 7905
rect 9060 7865 9100 7905
rect -37190 7860 9100 7865
rect -38770 7850 9100 7860
rect -38770 7815 -38755 7850
rect -38720 7815 -38710 7850
rect -38675 7815 -38665 7850
rect -38630 7815 -38620 7850
rect -38585 7815 -38575 7850
rect -38540 7815 -38530 7850
rect -38495 7815 -38485 7850
rect -38450 7815 -38440 7850
rect -38405 7815 -38395 7850
rect -38360 7815 -38350 7850
rect -38315 7815 -38305 7850
rect -38270 7815 -38260 7850
rect -38225 7815 -38215 7850
rect -38180 7815 -38170 7850
rect -38135 7815 -38125 7850
rect -38090 7815 -38080 7850
rect -38045 7815 -38035 7850
rect -38000 7815 -37990 7850
rect -37955 7815 -37945 7850
rect -37910 7815 -37900 7850
rect -37865 7815 -37855 7850
rect -37820 7815 -37810 7850
rect -37775 7815 -37765 7850
rect -37730 7815 -37720 7850
rect -37685 7815 -37675 7850
rect -37640 7815 -37630 7850
rect -37595 7815 -37585 7850
rect -37550 7815 -37540 7850
rect -37505 7815 -37495 7850
rect -37460 7815 -37450 7850
rect -37415 7815 -37405 7850
rect -37370 7815 -37360 7850
rect -37325 7815 -37315 7850
rect -37280 7815 -37270 7850
rect -37235 7815 -37225 7850
rect -37190 7835 9100 7850
rect -37190 7815 -80 7835
rect -38770 7805 -80 7815
rect -38770 7770 -38755 7805
rect -38720 7770 -38710 7805
rect -38675 7770 -38665 7805
rect -38630 7770 -38620 7805
rect -38585 7770 -38575 7805
rect -38540 7770 -38530 7805
rect -38495 7770 -38485 7805
rect -38450 7770 -38440 7805
rect -38405 7770 -38395 7805
rect -38360 7770 -38350 7805
rect -38315 7770 -38305 7805
rect -38270 7770 -38260 7805
rect -38225 7770 -38215 7805
rect -38180 7770 -38170 7805
rect -38135 7770 -38125 7805
rect -38090 7770 -38080 7805
rect -38045 7770 -38035 7805
rect -38000 7770 -37990 7805
rect -37955 7770 -37945 7805
rect -37910 7770 -37900 7805
rect -37865 7770 -37855 7805
rect -37820 7770 -37810 7805
rect -37775 7770 -37765 7805
rect -37730 7770 -37720 7805
rect -37685 7770 -37675 7805
rect -37640 7770 -37630 7805
rect -37595 7770 -37585 7805
rect -37550 7770 -37540 7805
rect -37505 7770 -37495 7805
rect -37460 7770 -37450 7805
rect -37415 7770 -37405 7805
rect -37370 7770 -37360 7805
rect -37325 7770 -37315 7805
rect -37280 7770 -37270 7805
rect -37235 7770 -37225 7805
rect -37190 7795 -80 7805
rect -40 7795 270 7835
rect 310 7795 620 7835
rect 660 7795 970 7835
rect 1010 7795 1670 7835
rect 1710 7795 2245 7835
rect 2285 7795 3175 7835
rect 3215 7795 3235 7835
rect 3275 7795 3345 7835
rect 3385 7795 6700 7835
rect 6740 7795 7270 7835
rect 7310 7795 7970 7835
rect 8010 7795 8320 7835
rect 8360 7795 8670 7835
rect 8710 7795 9020 7835
rect 9060 7795 9100 7835
rect -37190 7770 9100 7795
rect -38770 7765 9100 7770
rect -38770 7760 -80 7765
rect -38770 7725 -38755 7760
rect -38720 7725 -38710 7760
rect -38675 7725 -38665 7760
rect -38630 7725 -38620 7760
rect -38585 7725 -38575 7760
rect -38540 7725 -38530 7760
rect -38495 7725 -38485 7760
rect -38450 7725 -38440 7760
rect -38405 7725 -38395 7760
rect -38360 7725 -38350 7760
rect -38315 7725 -38305 7760
rect -38270 7725 -38260 7760
rect -38225 7725 -38215 7760
rect -38180 7725 -38170 7760
rect -38135 7725 -38125 7760
rect -38090 7725 -38080 7760
rect -38045 7725 -38035 7760
rect -38000 7725 -37990 7760
rect -37955 7725 -37945 7760
rect -37910 7725 -37900 7760
rect -37865 7725 -37855 7760
rect -37820 7725 -37810 7760
rect -37775 7725 -37765 7760
rect -37730 7725 -37720 7760
rect -37685 7725 -37675 7760
rect -37640 7725 -37630 7760
rect -37595 7725 -37585 7760
rect -37550 7725 -37540 7760
rect -37505 7725 -37495 7760
rect -37460 7725 -37450 7760
rect -37415 7725 -37405 7760
rect -37370 7725 -37360 7760
rect -37325 7725 -37315 7760
rect -37280 7725 -37270 7760
rect -37235 7725 -37225 7760
rect -37190 7725 -80 7760
rect -40 7725 270 7765
rect 310 7725 620 7765
rect 660 7725 970 7765
rect 1010 7725 1670 7765
rect 1710 7725 2245 7765
rect 2285 7725 3175 7765
rect 3215 7725 3235 7765
rect 3275 7725 3345 7765
rect 3385 7725 6700 7765
rect 6740 7725 7270 7765
rect 7310 7725 7970 7765
rect 8010 7725 8320 7765
rect 8360 7725 8670 7765
rect 8710 7725 9020 7765
rect 9060 7725 9100 7765
rect -38770 7715 9100 7725
rect -38770 7680 -38755 7715
rect -38720 7680 -38710 7715
rect -38675 7680 -38665 7715
rect -38630 7680 -38620 7715
rect -38585 7680 -38575 7715
rect -38540 7680 -38530 7715
rect -38495 7680 -38485 7715
rect -38450 7680 -38440 7715
rect -38405 7680 -38395 7715
rect -38360 7680 -38350 7715
rect -38315 7680 -38305 7715
rect -38270 7680 -38260 7715
rect -38225 7680 -38215 7715
rect -38180 7680 -38170 7715
rect -38135 7680 -38125 7715
rect -38090 7680 -38080 7715
rect -38045 7680 -38035 7715
rect -38000 7680 -37990 7715
rect -37955 7680 -37945 7715
rect -37910 7680 -37900 7715
rect -37865 7680 -37855 7715
rect -37820 7680 -37810 7715
rect -37775 7680 -37765 7715
rect -37730 7680 -37720 7715
rect -37685 7680 -37675 7715
rect -37640 7680 -37630 7715
rect -37595 7680 -37585 7715
rect -37550 7680 -37540 7715
rect -37505 7680 -37495 7715
rect -37460 7680 -37450 7715
rect -37415 7680 -37405 7715
rect -37370 7680 -37360 7715
rect -37325 7680 -37315 7715
rect -37280 7680 -37270 7715
rect -37235 7680 -37225 7715
rect -37190 7700 9100 7715
rect -37190 7680 -80 7700
rect -38770 7670 -80 7680
rect -38770 7635 -38755 7670
rect -38720 7635 -38710 7670
rect -38675 7635 -38665 7670
rect -38630 7635 -38620 7670
rect -38585 7635 -38575 7670
rect -38540 7635 -38530 7670
rect -38495 7635 -38485 7670
rect -38450 7635 -38440 7670
rect -38405 7635 -38395 7670
rect -38360 7635 -38350 7670
rect -38315 7635 -38305 7670
rect -38270 7635 -38260 7670
rect -38225 7635 -38215 7670
rect -38180 7635 -38170 7670
rect -38135 7635 -38125 7670
rect -38090 7635 -38080 7670
rect -38045 7635 -38035 7670
rect -38000 7635 -37990 7670
rect -37955 7635 -37945 7670
rect -37910 7635 -37900 7670
rect -37865 7635 -37855 7670
rect -37820 7635 -37810 7670
rect -37775 7635 -37765 7670
rect -37730 7635 -37720 7670
rect -37685 7635 -37675 7670
rect -37640 7635 -37630 7670
rect -37595 7635 -37585 7670
rect -37550 7635 -37540 7670
rect -37505 7635 -37495 7670
rect -37460 7635 -37450 7670
rect -37415 7635 -37405 7670
rect -37370 7635 -37360 7670
rect -37325 7635 -37315 7670
rect -37280 7635 -37270 7670
rect -37235 7635 -37225 7670
rect -37190 7660 -80 7670
rect -40 7660 270 7700
rect 310 7660 620 7700
rect 660 7660 970 7700
rect 1010 7660 1670 7700
rect 1710 7660 2245 7700
rect 2285 7660 3175 7700
rect 3215 7660 3235 7700
rect 3275 7660 3345 7700
rect 3385 7660 6700 7700
rect 6740 7660 7270 7700
rect 7310 7660 7970 7700
rect 8010 7660 8320 7700
rect 8360 7660 8670 7700
rect 8710 7660 9020 7700
rect 9060 7660 9100 7700
rect -37190 7640 9100 7660
rect -37190 7635 -80 7640
rect -38770 7625 -80 7635
rect -38770 7590 -38755 7625
rect -38720 7590 -38710 7625
rect -38675 7590 -38665 7625
rect -38630 7590 -38620 7625
rect -38585 7590 -38575 7625
rect -38540 7590 -38530 7625
rect -38495 7590 -38485 7625
rect -38450 7590 -38440 7625
rect -38405 7590 -38395 7625
rect -38360 7590 -38350 7625
rect -38315 7590 -38305 7625
rect -38270 7590 -38260 7625
rect -38225 7590 -38215 7625
rect -38180 7590 -38170 7625
rect -38135 7590 -38125 7625
rect -38090 7590 -38080 7625
rect -38045 7590 -38035 7625
rect -38000 7590 -37990 7625
rect -37955 7590 -37945 7625
rect -37910 7590 -37900 7625
rect -37865 7590 -37855 7625
rect -37820 7590 -37810 7625
rect -37775 7590 -37765 7625
rect -37730 7590 -37720 7625
rect -37685 7590 -37675 7625
rect -37640 7590 -37630 7625
rect -37595 7590 -37585 7625
rect -37550 7590 -37540 7625
rect -37505 7590 -37495 7625
rect -37460 7590 -37450 7625
rect -37415 7590 -37405 7625
rect -37370 7590 -37360 7625
rect -37325 7590 -37315 7625
rect -37280 7590 -37270 7625
rect -37235 7590 -37225 7625
rect -37190 7600 -80 7625
rect -40 7600 270 7640
rect 310 7600 620 7640
rect 660 7600 970 7640
rect 1010 7600 1670 7640
rect 1710 7600 2245 7640
rect 2285 7600 3175 7640
rect 3215 7600 3235 7640
rect 3275 7600 3345 7640
rect 3385 7600 6700 7640
rect 6740 7600 7270 7640
rect 7310 7600 7970 7640
rect 8010 7600 8320 7640
rect 8360 7600 8670 7640
rect 8710 7600 9020 7640
rect 9060 7600 9100 7640
rect -37190 7590 9100 7600
rect -38770 7580 9100 7590
rect -38770 7545 -38755 7580
rect -38720 7545 -38710 7580
rect -38675 7545 -38665 7580
rect -38630 7545 -38620 7580
rect -38585 7545 -38575 7580
rect -38540 7545 -38530 7580
rect -38495 7545 -38485 7580
rect -38450 7545 -38440 7580
rect -38405 7545 -38395 7580
rect -38360 7545 -38350 7580
rect -38315 7545 -38305 7580
rect -38270 7545 -38260 7580
rect -38225 7545 -38215 7580
rect -38180 7545 -38170 7580
rect -38135 7545 -38125 7580
rect -38090 7545 -38080 7580
rect -38045 7545 -38035 7580
rect -38000 7545 -37990 7580
rect -37955 7545 -37945 7580
rect -37910 7545 -37900 7580
rect -37865 7545 -37855 7580
rect -37820 7545 -37810 7580
rect -37775 7545 -37765 7580
rect -37730 7545 -37720 7580
rect -37685 7545 -37675 7580
rect -37640 7545 -37630 7580
rect -37595 7545 -37585 7580
rect -37550 7545 -37540 7580
rect -37505 7545 -37495 7580
rect -37460 7545 -37450 7580
rect -37415 7545 -37405 7580
rect -37370 7545 -37360 7580
rect -37325 7545 -37315 7580
rect -37280 7545 -37270 7580
rect -37235 7545 -37225 7580
rect -37190 7575 9100 7580
rect -37190 7545 -80 7575
rect -38770 7535 -80 7545
rect -40 7535 270 7575
rect 310 7535 620 7575
rect 660 7535 970 7575
rect 1010 7535 1670 7575
rect 1710 7535 2245 7575
rect 2285 7535 3175 7575
rect 3215 7535 3235 7575
rect 3275 7535 3345 7575
rect 3385 7535 6700 7575
rect 6740 7535 7270 7575
rect 7310 7535 7970 7575
rect 8010 7535 8320 7575
rect 8360 7535 8670 7575
rect 8710 7535 9020 7575
rect 9060 7535 9100 7575
rect -38770 7500 -38755 7535
rect -38720 7500 -38710 7535
rect -38675 7500 -38665 7535
rect -38630 7500 -38620 7535
rect -38585 7500 -38575 7535
rect -38540 7500 -38530 7535
rect -38495 7500 -38485 7535
rect -38450 7500 -38440 7535
rect -38405 7500 -38395 7535
rect -38360 7500 -38350 7535
rect -38315 7500 -38305 7535
rect -38270 7500 -38260 7535
rect -38225 7500 -38215 7535
rect -38180 7500 -38170 7535
rect -38135 7500 -38125 7535
rect -38090 7500 -38080 7535
rect -38045 7500 -38035 7535
rect -38000 7500 -37990 7535
rect -37955 7500 -37945 7535
rect -37910 7500 -37900 7535
rect -37865 7500 -37855 7535
rect -37820 7500 -37810 7535
rect -37775 7500 -37765 7535
rect -37730 7500 -37720 7535
rect -37685 7500 -37675 7535
rect -37640 7500 -37630 7535
rect -37595 7500 -37585 7535
rect -37550 7500 -37540 7535
rect -37505 7500 -37495 7535
rect -37460 7500 -37450 7535
rect -37415 7500 -37405 7535
rect -37370 7500 -37360 7535
rect -37325 7500 -37315 7535
rect -37280 7500 -37270 7535
rect -37235 7500 -37225 7535
rect -37190 7505 9100 7535
rect -37190 7500 -80 7505
rect -38770 7490 -80 7500
rect -38770 7455 -38755 7490
rect -38720 7455 -38710 7490
rect -38675 7455 -38665 7490
rect -38630 7455 -38620 7490
rect -38585 7455 -38575 7490
rect -38540 7455 -38530 7490
rect -38495 7455 -38485 7490
rect -38450 7455 -38440 7490
rect -38405 7455 -38395 7490
rect -38360 7455 -38350 7490
rect -38315 7455 -38305 7490
rect -38270 7455 -38260 7490
rect -38225 7455 -38215 7490
rect -38180 7455 -38170 7490
rect -38135 7455 -38125 7490
rect -38090 7455 -38080 7490
rect -38045 7455 -38035 7490
rect -38000 7455 -37990 7490
rect -37955 7455 -37945 7490
rect -37910 7455 -37900 7490
rect -37865 7455 -37855 7490
rect -37820 7455 -37810 7490
rect -37775 7455 -37765 7490
rect -37730 7455 -37720 7490
rect -37685 7455 -37675 7490
rect -37640 7455 -37630 7490
rect -37595 7455 -37585 7490
rect -37550 7455 -37540 7490
rect -37505 7455 -37495 7490
rect -37460 7455 -37450 7490
rect -37415 7455 -37405 7490
rect -37370 7455 -37360 7490
rect -37325 7455 -37315 7490
rect -37280 7455 -37270 7490
rect -37235 7455 -37225 7490
rect -37190 7465 -80 7490
rect -40 7465 270 7505
rect 310 7465 620 7505
rect 660 7465 970 7505
rect 1010 7465 1670 7505
rect 1710 7465 2245 7505
rect 2285 7465 3175 7505
rect 3215 7465 3235 7505
rect 3275 7465 3345 7505
rect 3385 7465 6700 7505
rect 6740 7465 7270 7505
rect 7310 7465 7970 7505
rect 8010 7465 8320 7505
rect 8360 7465 8670 7505
rect 8710 7465 9020 7505
rect 9060 7465 9100 7505
rect -37190 7455 9100 7465
rect -38770 7445 9100 7455
rect -38770 7410 -38755 7445
rect -38720 7410 -38710 7445
rect -38675 7410 -38665 7445
rect -38630 7410 -38620 7445
rect -38585 7410 -38575 7445
rect -38540 7410 -38530 7445
rect -38495 7410 -38485 7445
rect -38450 7410 -38440 7445
rect -38405 7410 -38395 7445
rect -38360 7410 -38350 7445
rect -38315 7410 -38305 7445
rect -38270 7410 -38260 7445
rect -38225 7410 -38215 7445
rect -38180 7410 -38170 7445
rect -38135 7410 -38125 7445
rect -38090 7410 -38080 7445
rect -38045 7410 -38035 7445
rect -38000 7410 -37990 7445
rect -37955 7410 -37945 7445
rect -37910 7410 -37900 7445
rect -37865 7410 -37855 7445
rect -37820 7410 -37810 7445
rect -37775 7410 -37765 7445
rect -37730 7410 -37720 7445
rect -37685 7410 -37675 7445
rect -37640 7410 -37630 7445
rect -37595 7410 -37585 7445
rect -37550 7410 -37540 7445
rect -37505 7410 -37495 7445
rect -37460 7410 -37450 7445
rect -37415 7410 -37405 7445
rect -37370 7410 -37360 7445
rect -37325 7410 -37315 7445
rect -37280 7410 -37270 7445
rect -37235 7410 -37225 7445
rect -37190 7435 9100 7445
rect -37190 7410 -80 7435
rect -38770 7400 -80 7410
rect -38770 7365 -38755 7400
rect -38720 7365 -38710 7400
rect -38675 7365 -38665 7400
rect -38630 7365 -38620 7400
rect -38585 7365 -38575 7400
rect -38540 7365 -38530 7400
rect -38495 7365 -38485 7400
rect -38450 7365 -38440 7400
rect -38405 7365 -38395 7400
rect -38360 7365 -38350 7400
rect -38315 7365 -38305 7400
rect -38270 7365 -38260 7400
rect -38225 7365 -38215 7400
rect -38180 7365 -38170 7400
rect -38135 7365 -38125 7400
rect -38090 7365 -38080 7400
rect -38045 7365 -38035 7400
rect -38000 7365 -37990 7400
rect -37955 7365 -37945 7400
rect -37910 7365 -37900 7400
rect -37865 7365 -37855 7400
rect -37820 7365 -37810 7400
rect -37775 7365 -37765 7400
rect -37730 7365 -37720 7400
rect -37685 7365 -37675 7400
rect -37640 7365 -37630 7400
rect -37595 7365 -37585 7400
rect -37550 7365 -37540 7400
rect -37505 7365 -37495 7400
rect -37460 7365 -37450 7400
rect -37415 7365 -37405 7400
rect -37370 7365 -37360 7400
rect -37325 7365 -37315 7400
rect -37280 7365 -37270 7400
rect -37235 7365 -37225 7400
rect -37190 7395 -80 7400
rect -40 7395 270 7435
rect 310 7395 620 7435
rect 660 7395 970 7435
rect 1010 7395 1670 7435
rect 1710 7395 2245 7435
rect 2285 7395 3175 7435
rect 3215 7395 3235 7435
rect 3275 7395 3345 7435
rect 3385 7395 6700 7435
rect 6740 7395 7270 7435
rect 7310 7395 7970 7435
rect 8010 7395 8320 7435
rect 8360 7395 8670 7435
rect 8710 7395 9020 7435
rect 9060 7395 9100 7435
rect -37190 7365 9100 7395
rect -38770 7355 -80 7365
rect -38770 7320 -38755 7355
rect -38720 7320 -38710 7355
rect -38675 7320 -38665 7355
rect -38630 7320 -38620 7355
rect -38585 7320 -38575 7355
rect -38540 7320 -38530 7355
rect -38495 7320 -38485 7355
rect -38450 7320 -38440 7355
rect -38405 7320 -38395 7355
rect -38360 7320 -38350 7355
rect -38315 7320 -38305 7355
rect -38270 7320 -38260 7355
rect -38225 7320 -38215 7355
rect -38180 7320 -38170 7355
rect -38135 7320 -38125 7355
rect -38090 7320 -38080 7355
rect -38045 7320 -38035 7355
rect -38000 7320 -37990 7355
rect -37955 7320 -37945 7355
rect -37910 7320 -37900 7355
rect -37865 7320 -37855 7355
rect -37820 7320 -37810 7355
rect -37775 7320 -37765 7355
rect -37730 7320 -37720 7355
rect -37685 7320 -37675 7355
rect -37640 7320 -37630 7355
rect -37595 7320 -37585 7355
rect -37550 7320 -37540 7355
rect -37505 7320 -37495 7355
rect -37460 7320 -37450 7355
rect -37415 7320 -37405 7355
rect -37370 7320 -37360 7355
rect -37325 7320 -37315 7355
rect -37280 7320 -37270 7355
rect -37235 7320 -37225 7355
rect -37190 7325 -80 7355
rect -40 7325 270 7365
rect 310 7325 620 7365
rect 660 7325 970 7365
rect 1010 7325 1670 7365
rect 1710 7325 2245 7365
rect 2285 7325 3175 7365
rect 3215 7325 3235 7365
rect 3275 7325 3345 7365
rect 3385 7325 6700 7365
rect 6740 7325 7270 7365
rect 7310 7325 7970 7365
rect 8010 7325 8320 7365
rect 8360 7325 8670 7365
rect 8710 7325 9020 7365
rect 9060 7325 9100 7365
rect -37190 7320 9100 7325
rect -38770 7310 9100 7320
rect -38770 7275 -38755 7310
rect -38720 7275 -38710 7310
rect -38675 7275 -38665 7310
rect -38630 7275 -38620 7310
rect -38585 7275 -38575 7310
rect -38540 7275 -38530 7310
rect -38495 7275 -38485 7310
rect -38450 7275 -38440 7310
rect -38405 7275 -38395 7310
rect -38360 7275 -38350 7310
rect -38315 7275 -38305 7310
rect -38270 7275 -38260 7310
rect -38225 7275 -38215 7310
rect -38180 7275 -38170 7310
rect -38135 7275 -38125 7310
rect -38090 7275 -38080 7310
rect -38045 7275 -38035 7310
rect -38000 7275 -37990 7310
rect -37955 7275 -37945 7310
rect -37910 7275 -37900 7310
rect -37865 7275 -37855 7310
rect -37820 7275 -37810 7310
rect -37775 7275 -37765 7310
rect -37730 7275 -37720 7310
rect -37685 7275 -37675 7310
rect -37640 7275 -37630 7310
rect -37595 7275 -37585 7310
rect -37550 7275 -37540 7310
rect -37505 7275 -37495 7310
rect -37460 7275 -37450 7310
rect -37415 7275 -37405 7310
rect -37370 7275 -37360 7310
rect -37325 7275 -37315 7310
rect -37280 7275 -37270 7310
rect -37235 7275 -37225 7310
rect -37190 7300 9100 7310
rect -37190 7275 -80 7300
rect -38770 7265 -80 7275
rect -38770 7230 -38755 7265
rect -38720 7230 -38710 7265
rect -38675 7230 -38665 7265
rect -38630 7230 -38620 7265
rect -38585 7230 -38575 7265
rect -38540 7230 -38530 7265
rect -38495 7230 -38485 7265
rect -38450 7230 -38440 7265
rect -38405 7230 -38395 7265
rect -38360 7230 -38350 7265
rect -38315 7230 -38305 7265
rect -38270 7230 -38260 7265
rect -38225 7230 -38215 7265
rect -38180 7230 -38170 7265
rect -38135 7230 -38125 7265
rect -38090 7230 -38080 7265
rect -38045 7230 -38035 7265
rect -38000 7230 -37990 7265
rect -37955 7230 -37945 7265
rect -37910 7230 -37900 7265
rect -37865 7230 -37855 7265
rect -37820 7230 -37810 7265
rect -37775 7230 -37765 7265
rect -37730 7230 -37720 7265
rect -37685 7230 -37675 7265
rect -37640 7230 -37630 7265
rect -37595 7230 -37585 7265
rect -37550 7230 -37540 7265
rect -37505 7230 -37495 7265
rect -37460 7230 -37450 7265
rect -37415 7230 -37405 7265
rect -37370 7230 -37360 7265
rect -37325 7230 -37315 7265
rect -37280 7230 -37270 7265
rect -37235 7230 -37225 7265
rect -37190 7260 -80 7265
rect -40 7260 270 7300
rect 310 7260 620 7300
rect 660 7260 970 7300
rect 1010 7260 1670 7300
rect 1710 7260 2245 7300
rect 2285 7260 3175 7300
rect 3215 7260 3235 7300
rect 3275 7260 3345 7300
rect 3385 7260 6700 7300
rect 6740 7260 7270 7300
rect 7310 7260 7970 7300
rect 8010 7260 8320 7300
rect 8360 7260 8670 7300
rect 8710 7260 9020 7300
rect 9060 7260 9100 7300
rect -37190 7240 9100 7260
rect -37190 7230 -80 7240
rect -38770 7220 -80 7230
rect -38770 7185 -38755 7220
rect -38720 7185 -38710 7220
rect -38675 7185 -38665 7220
rect -38630 7185 -38620 7220
rect -38585 7185 -38575 7220
rect -38540 7185 -38530 7220
rect -38495 7185 -38485 7220
rect -38450 7185 -38440 7220
rect -38405 7185 -38395 7220
rect -38360 7185 -38350 7220
rect -38315 7185 -38305 7220
rect -38270 7185 -38260 7220
rect -38225 7185 -38215 7220
rect -38180 7185 -38170 7220
rect -38135 7185 -38125 7220
rect -38090 7185 -38080 7220
rect -38045 7185 -38035 7220
rect -38000 7185 -37990 7220
rect -37955 7185 -37945 7220
rect -37910 7185 -37900 7220
rect -37865 7185 -37855 7220
rect -37820 7185 -37810 7220
rect -37775 7185 -37765 7220
rect -37730 7185 -37720 7220
rect -37685 7185 -37675 7220
rect -37640 7185 -37630 7220
rect -37595 7185 -37585 7220
rect -37550 7185 -37540 7220
rect -37505 7185 -37495 7220
rect -37460 7185 -37450 7220
rect -37415 7185 -37405 7220
rect -37370 7185 -37360 7220
rect -37325 7185 -37315 7220
rect -37280 7185 -37270 7220
rect -37235 7185 -37225 7220
rect -37190 7200 -80 7220
rect -40 7200 270 7240
rect 310 7200 620 7240
rect 660 7200 970 7240
rect 1010 7200 1670 7240
rect 1710 7200 2245 7240
rect 2285 7200 3175 7240
rect 3215 7200 3235 7240
rect 3275 7200 3345 7240
rect 3385 7200 6700 7240
rect 6740 7200 7270 7240
rect 7310 7200 7970 7240
rect 8010 7200 8320 7240
rect 8360 7200 8670 7240
rect 8710 7200 9020 7240
rect 9060 7200 9100 7240
rect -37190 7185 9100 7200
rect -38770 7175 9100 7185
rect -38770 7140 -38755 7175
rect -38720 7140 -38710 7175
rect -38675 7140 -38665 7175
rect -38630 7140 -38620 7175
rect -38585 7140 -38575 7175
rect -38540 7140 -38530 7175
rect -38495 7140 -38485 7175
rect -38450 7140 -38440 7175
rect -38405 7140 -38395 7175
rect -38360 7140 -38350 7175
rect -38315 7140 -38305 7175
rect -38270 7140 -38260 7175
rect -38225 7140 -38215 7175
rect -38180 7140 -38170 7175
rect -38135 7140 -38125 7175
rect -38090 7140 -38080 7175
rect -38045 7140 -38035 7175
rect -38000 7140 -37990 7175
rect -37955 7140 -37945 7175
rect -37910 7140 -37900 7175
rect -37865 7140 -37855 7175
rect -37820 7140 -37810 7175
rect -37775 7140 -37765 7175
rect -37730 7140 -37720 7175
rect -37685 7140 -37675 7175
rect -37640 7140 -37630 7175
rect -37595 7140 -37585 7175
rect -37550 7140 -37540 7175
rect -37505 7140 -37495 7175
rect -37460 7140 -37450 7175
rect -37415 7140 -37405 7175
rect -37370 7140 -37360 7175
rect -37325 7140 -37315 7175
rect -37280 7140 -37270 7175
rect -37235 7140 -37225 7175
rect -37190 7140 -80 7175
rect -38770 7135 -80 7140
rect -40 7135 270 7175
rect 310 7135 620 7175
rect 660 7135 970 7175
rect 1010 7135 1670 7175
rect 1710 7135 2245 7175
rect 2285 7135 3175 7175
rect 3215 7135 3235 7175
rect 3275 7135 3345 7175
rect 3385 7135 6700 7175
rect 6740 7135 7270 7175
rect 7310 7135 7970 7175
rect 8010 7135 8320 7175
rect 8360 7135 8670 7175
rect 8710 7135 9020 7175
rect 9060 7135 9100 7175
rect -38770 7130 9100 7135
rect -38770 7095 -38755 7130
rect -38720 7095 -38710 7130
rect -38675 7095 -38665 7130
rect -38630 7095 -38620 7130
rect -38585 7095 -38575 7130
rect -38540 7095 -38530 7130
rect -38495 7095 -38485 7130
rect -38450 7095 -38440 7130
rect -38405 7095 -38395 7130
rect -38360 7095 -38350 7130
rect -38315 7095 -38305 7130
rect -38270 7095 -38260 7130
rect -38225 7095 -38215 7130
rect -38180 7095 -38170 7130
rect -38135 7095 -38125 7130
rect -38090 7095 -38080 7130
rect -38045 7095 -38035 7130
rect -38000 7095 -37990 7130
rect -37955 7095 -37945 7130
rect -37910 7095 -37900 7130
rect -37865 7095 -37855 7130
rect -37820 7095 -37810 7130
rect -37775 7095 -37765 7130
rect -37730 7095 -37720 7130
rect -37685 7095 -37675 7130
rect -37640 7095 -37630 7130
rect -37595 7095 -37585 7130
rect -37550 7095 -37540 7130
rect -37505 7095 -37495 7130
rect -37460 7095 -37450 7130
rect -37415 7095 -37405 7130
rect -37370 7095 -37360 7130
rect -37325 7095 -37315 7130
rect -37280 7095 -37270 7130
rect -37235 7095 -37225 7130
rect -37190 7105 9100 7130
rect -37190 7095 -80 7105
rect -38770 7085 -80 7095
rect -38770 7050 -38755 7085
rect -38720 7050 -38710 7085
rect -38675 7050 -38665 7085
rect -38630 7050 -38620 7085
rect -38585 7050 -38575 7085
rect -38540 7050 -38530 7085
rect -38495 7050 -38485 7085
rect -38450 7050 -38440 7085
rect -38405 7050 -38395 7085
rect -38360 7050 -38350 7085
rect -38315 7050 -38305 7085
rect -38270 7050 -38260 7085
rect -38225 7050 -38215 7085
rect -38180 7050 -38170 7085
rect -38135 7050 -38125 7085
rect -38090 7050 -38080 7085
rect -38045 7050 -38035 7085
rect -38000 7050 -37990 7085
rect -37955 7050 -37945 7085
rect -37910 7050 -37900 7085
rect -37865 7050 -37855 7085
rect -37820 7050 -37810 7085
rect -37775 7050 -37765 7085
rect -37730 7050 -37720 7085
rect -37685 7050 -37675 7085
rect -37640 7050 -37630 7085
rect -37595 7050 -37585 7085
rect -37550 7050 -37540 7085
rect -37505 7050 -37495 7085
rect -37460 7050 -37450 7085
rect -37415 7050 -37405 7085
rect -37370 7050 -37360 7085
rect -37325 7050 -37315 7085
rect -37280 7050 -37270 7085
rect -37235 7050 -37225 7085
rect -37190 7065 -80 7085
rect -40 7065 270 7105
rect 310 7065 620 7105
rect 660 7065 970 7105
rect 1010 7065 1670 7105
rect 1710 7065 2245 7105
rect 2285 7065 3175 7105
rect 3215 7065 3235 7105
rect 3275 7065 3345 7105
rect 3385 7065 6700 7105
rect 6740 7065 7270 7105
rect 7310 7065 7970 7105
rect 8010 7065 8320 7105
rect 8360 7065 8670 7105
rect 8710 7065 9020 7105
rect 9060 7065 9100 7105
rect -37190 7050 9100 7065
rect -38770 7040 9100 7050
rect -38770 7005 -38755 7040
rect -38720 7005 -38710 7040
rect -38675 7005 -38665 7040
rect -38630 7005 -38620 7040
rect -38585 7005 -38575 7040
rect -38540 7005 -38530 7040
rect -38495 7005 -38485 7040
rect -38450 7005 -38440 7040
rect -38405 7005 -38395 7040
rect -38360 7005 -38350 7040
rect -38315 7005 -38305 7040
rect -38270 7005 -38260 7040
rect -38225 7005 -38215 7040
rect -38180 7005 -38170 7040
rect -38135 7005 -38125 7040
rect -38090 7005 -38080 7040
rect -38045 7005 -38035 7040
rect -38000 7005 -37990 7040
rect -37955 7005 -37945 7040
rect -37910 7005 -37900 7040
rect -37865 7005 -37855 7040
rect -37820 7005 -37810 7040
rect -37775 7005 -37765 7040
rect -37730 7005 -37720 7040
rect -37685 7005 -37675 7040
rect -37640 7005 -37630 7040
rect -37595 7005 -37585 7040
rect -37550 7005 -37540 7040
rect -37505 7005 -37495 7040
rect -37460 7005 -37450 7040
rect -37415 7005 -37405 7040
rect -37370 7005 -37360 7040
rect -37325 7005 -37315 7040
rect -37280 7005 -37270 7040
rect -37235 7005 -37225 7040
rect -37190 7035 9100 7040
rect -37190 7005 -80 7035
rect -38770 6995 -80 7005
rect -40 6995 270 7035
rect 310 6995 620 7035
rect 660 6995 970 7035
rect 1010 6995 1670 7035
rect 1710 6995 2245 7035
rect 2285 6995 3175 7035
rect 3215 6995 3235 7035
rect 3275 6995 3345 7035
rect 3385 6995 6700 7035
rect 6740 6995 7270 7035
rect 7310 6995 7970 7035
rect 8010 6995 8320 7035
rect 8360 6995 8670 7035
rect 8710 6995 9020 7035
rect 9060 6995 9100 7035
rect -38770 6960 -38755 6995
rect -38720 6960 -38710 6995
rect -38675 6960 -38665 6995
rect -38630 6960 -38620 6995
rect -38585 6960 -38575 6995
rect -38540 6960 -38530 6995
rect -38495 6960 -38485 6995
rect -38450 6960 -38440 6995
rect -38405 6960 -38395 6995
rect -38360 6960 -38350 6995
rect -38315 6960 -38305 6995
rect -38270 6960 -38260 6995
rect -38225 6960 -38215 6995
rect -38180 6960 -38170 6995
rect -38135 6960 -38125 6995
rect -38090 6960 -38080 6995
rect -38045 6960 -38035 6995
rect -38000 6960 -37990 6995
rect -37955 6960 -37945 6995
rect -37910 6960 -37900 6995
rect -37865 6960 -37855 6995
rect -37820 6960 -37810 6995
rect -37775 6960 -37765 6995
rect -37730 6960 -37720 6995
rect -37685 6960 -37675 6995
rect -37640 6960 -37630 6995
rect -37595 6960 -37585 6995
rect -37550 6960 -37540 6995
rect -37505 6960 -37495 6995
rect -37460 6960 -37450 6995
rect -37415 6960 -37405 6995
rect -37370 6960 -37360 6995
rect -37325 6960 -37315 6995
rect -37280 6960 -37270 6995
rect -37235 6960 -37225 6995
rect -37190 6965 9100 6995
rect -37190 6960 -80 6965
rect -38770 6950 -80 6960
rect -38770 6915 -38755 6950
rect -38720 6915 -38710 6950
rect -38675 6915 -38665 6950
rect -38630 6915 -38620 6950
rect -38585 6915 -38575 6950
rect -38540 6915 -38530 6950
rect -38495 6915 -38485 6950
rect -38450 6915 -38440 6950
rect -38405 6915 -38395 6950
rect -38360 6915 -38350 6950
rect -38315 6915 -38305 6950
rect -38270 6915 -38260 6950
rect -38225 6915 -38215 6950
rect -38180 6915 -38170 6950
rect -38135 6915 -38125 6950
rect -38090 6915 -38080 6950
rect -38045 6915 -38035 6950
rect -38000 6915 -37990 6950
rect -37955 6915 -37945 6950
rect -37910 6915 -37900 6950
rect -37865 6915 -37855 6950
rect -37820 6915 -37810 6950
rect -37775 6915 -37765 6950
rect -37730 6915 -37720 6950
rect -37685 6915 -37675 6950
rect -37640 6915 -37630 6950
rect -37595 6915 -37585 6950
rect -37550 6915 -37540 6950
rect -37505 6915 -37495 6950
rect -37460 6915 -37450 6950
rect -37415 6915 -37405 6950
rect -37370 6915 -37360 6950
rect -37325 6915 -37315 6950
rect -37280 6915 -37270 6950
rect -37235 6915 -37225 6950
rect -37190 6925 -80 6950
rect -40 6925 270 6965
rect 310 6925 620 6965
rect 660 6925 970 6965
rect 1010 6925 1670 6965
rect 1710 6925 2245 6965
rect 2285 6925 3175 6965
rect 3215 6925 3235 6965
rect 3275 6925 3345 6965
rect 3385 6925 6700 6965
rect 6740 6925 7270 6965
rect 7310 6925 7970 6965
rect 8010 6925 8320 6965
rect 8360 6925 8670 6965
rect 8710 6925 9020 6965
rect 9060 6925 9100 6965
rect -37190 6915 9100 6925
rect -38770 6905 9100 6915
rect -38770 6870 -38755 6905
rect -38720 6870 -38710 6905
rect -38675 6870 -38665 6905
rect -38630 6870 -38620 6905
rect -38585 6870 -38575 6905
rect -38540 6870 -38530 6905
rect -38495 6870 -38485 6905
rect -38450 6870 -38440 6905
rect -38405 6870 -38395 6905
rect -38360 6870 -38350 6905
rect -38315 6870 -38305 6905
rect -38270 6870 -38260 6905
rect -38225 6870 -38215 6905
rect -38180 6870 -38170 6905
rect -38135 6870 -38125 6905
rect -38090 6870 -38080 6905
rect -38045 6870 -38035 6905
rect -38000 6870 -37990 6905
rect -37955 6870 -37945 6905
rect -37910 6870 -37900 6905
rect -37865 6870 -37855 6905
rect -37820 6870 -37810 6905
rect -37775 6870 -37765 6905
rect -37730 6870 -37720 6905
rect -37685 6870 -37675 6905
rect -37640 6870 -37630 6905
rect -37595 6870 -37585 6905
rect -37550 6870 -37540 6905
rect -37505 6870 -37495 6905
rect -37460 6870 -37450 6905
rect -37415 6870 -37405 6905
rect -37370 6870 -37360 6905
rect -37325 6870 -37315 6905
rect -37280 6870 -37270 6905
rect -37235 6870 -37225 6905
rect -37190 6900 9100 6905
rect -37190 6870 -80 6900
rect -38770 6860 -80 6870
rect -40 6860 270 6900
rect 310 6860 620 6900
rect 660 6860 970 6900
rect 1010 6860 1670 6900
rect 1710 6860 2245 6900
rect 2285 6860 3175 6900
rect 3215 6860 3235 6900
rect 3275 6860 3345 6900
rect 3385 6860 6700 6900
rect 6740 6860 7270 6900
rect 7310 6860 7970 6900
rect 8010 6860 8320 6900
rect 8360 6860 8670 6900
rect 8710 6860 9020 6900
rect 9060 6860 9100 6900
rect -38770 6825 -38755 6860
rect -38720 6825 -38710 6860
rect -38675 6825 -38665 6860
rect -38630 6825 -38620 6860
rect -38585 6825 -38575 6860
rect -38540 6825 -38530 6860
rect -38495 6825 -38485 6860
rect -38450 6825 -38440 6860
rect -38405 6825 -38395 6860
rect -38360 6825 -38350 6860
rect -38315 6825 -38305 6860
rect -38270 6825 -38260 6860
rect -38225 6825 -38215 6860
rect -38180 6825 -38170 6860
rect -38135 6825 -38125 6860
rect -38090 6825 -38080 6860
rect -38045 6825 -38035 6860
rect -38000 6825 -37990 6860
rect -37955 6825 -37945 6860
rect -37910 6825 -37900 6860
rect -37865 6825 -37855 6860
rect -37820 6825 -37810 6860
rect -37775 6825 -37765 6860
rect -37730 6825 -37720 6860
rect -37685 6825 -37675 6860
rect -37640 6825 -37630 6860
rect -37595 6825 -37585 6860
rect -37550 6825 -37540 6860
rect -37505 6825 -37495 6860
rect -37460 6825 -37450 6860
rect -37415 6825 -37405 6860
rect -37370 6825 -37360 6860
rect -37325 6825 -37315 6860
rect -37280 6825 -37270 6860
rect -37235 6825 -37225 6860
rect -37190 6840 9100 6860
rect -37190 6825 -80 6840
rect -38770 6815 -80 6825
rect -38770 6780 -38755 6815
rect -38720 6780 -38710 6815
rect -38675 6780 -38665 6815
rect -38630 6780 -38620 6815
rect -38585 6780 -38575 6815
rect -38540 6780 -38530 6815
rect -38495 6780 -38485 6815
rect -38450 6780 -38440 6815
rect -38405 6780 -38395 6815
rect -38360 6780 -38350 6815
rect -38315 6780 -38305 6815
rect -38270 6780 -38260 6815
rect -38225 6780 -38215 6815
rect -38180 6780 -38170 6815
rect -38135 6780 -38125 6815
rect -38090 6780 -38080 6815
rect -38045 6780 -38035 6815
rect -38000 6780 -37990 6815
rect -37955 6780 -37945 6815
rect -37910 6780 -37900 6815
rect -37865 6780 -37855 6815
rect -37820 6780 -37810 6815
rect -37775 6780 -37765 6815
rect -37730 6780 -37720 6815
rect -37685 6780 -37675 6815
rect -37640 6780 -37630 6815
rect -37595 6780 -37585 6815
rect -37550 6780 -37540 6815
rect -37505 6780 -37495 6815
rect -37460 6780 -37450 6815
rect -37415 6780 -37405 6815
rect -37370 6780 -37360 6815
rect -37325 6780 -37315 6815
rect -37280 6780 -37270 6815
rect -37235 6780 -37225 6815
rect -37190 6800 -80 6815
rect -40 6800 270 6840
rect 310 6800 620 6840
rect 660 6800 970 6840
rect 1010 6800 1670 6840
rect 1710 6800 2245 6840
rect 2285 6800 3175 6840
rect 3215 6800 3235 6840
rect 3275 6800 3345 6840
rect 3385 6800 6700 6840
rect 6740 6800 7270 6840
rect 7310 6800 7970 6840
rect 8010 6800 8320 6840
rect 8360 6800 8670 6840
rect 8710 6800 9020 6840
rect 9060 6800 9100 6840
rect -37190 6780 9100 6800
rect -38770 6775 9100 6780
rect -38770 6770 -80 6775
rect -38770 6735 -38755 6770
rect -38720 6735 -38710 6770
rect -38675 6735 -38665 6770
rect -38630 6735 -38620 6770
rect -38585 6735 -38575 6770
rect -38540 6735 -38530 6770
rect -38495 6735 -38485 6770
rect -38450 6735 -38440 6770
rect -38405 6735 -38395 6770
rect -38360 6735 -38350 6770
rect -38315 6735 -38305 6770
rect -38270 6735 -38260 6770
rect -38225 6735 -38215 6770
rect -38180 6735 -38170 6770
rect -38135 6735 -38125 6770
rect -38090 6735 -38080 6770
rect -38045 6735 -38035 6770
rect -38000 6735 -37990 6770
rect -37955 6735 -37945 6770
rect -37910 6735 -37900 6770
rect -37865 6735 -37855 6770
rect -37820 6735 -37810 6770
rect -37775 6735 -37765 6770
rect -37730 6735 -37720 6770
rect -37685 6735 -37675 6770
rect -37640 6735 -37630 6770
rect -37595 6735 -37585 6770
rect -37550 6735 -37540 6770
rect -37505 6735 -37495 6770
rect -37460 6735 -37450 6770
rect -37415 6735 -37405 6770
rect -37370 6735 -37360 6770
rect -37325 6735 -37315 6770
rect -37280 6735 -37270 6770
rect -37235 6735 -37225 6770
rect -37190 6735 -80 6770
rect -40 6735 270 6775
rect 310 6735 620 6775
rect 660 6735 970 6775
rect 1010 6735 1670 6775
rect 1710 6735 2245 6775
rect 2285 6735 3175 6775
rect 3215 6735 3235 6775
rect 3275 6735 3345 6775
rect 3385 6735 6700 6775
rect 6740 6735 7270 6775
rect 7310 6735 7970 6775
rect 8010 6735 8320 6775
rect 8360 6735 8670 6775
rect 8710 6735 9020 6775
rect 9060 6735 9100 6775
rect -38770 6725 9100 6735
rect -38770 6690 -38755 6725
rect -38720 6690 -38710 6725
rect -38675 6690 -38665 6725
rect -38630 6690 -38620 6725
rect -38585 6690 -38575 6725
rect -38540 6690 -38530 6725
rect -38495 6690 -38485 6725
rect -38450 6690 -38440 6725
rect -38405 6690 -38395 6725
rect -38360 6690 -38350 6725
rect -38315 6690 -38305 6725
rect -38270 6690 -38260 6725
rect -38225 6690 -38215 6725
rect -38180 6690 -38170 6725
rect -38135 6690 -38125 6725
rect -38090 6690 -38080 6725
rect -38045 6690 -38035 6725
rect -38000 6690 -37990 6725
rect -37955 6690 -37945 6725
rect -37910 6690 -37900 6725
rect -37865 6690 -37855 6725
rect -37820 6690 -37810 6725
rect -37775 6690 -37765 6725
rect -37730 6690 -37720 6725
rect -37685 6690 -37675 6725
rect -37640 6690 -37630 6725
rect -37595 6690 -37585 6725
rect -37550 6690 -37540 6725
rect -37505 6690 -37495 6725
rect -37460 6690 -37450 6725
rect -37415 6690 -37405 6725
rect -37370 6690 -37360 6725
rect -37325 6690 -37315 6725
rect -37280 6690 -37270 6725
rect -37235 6690 -37225 6725
rect -37190 6705 9100 6725
rect -37190 6690 -80 6705
rect -38770 6680 -80 6690
rect -38770 6645 -38755 6680
rect -38720 6645 -38710 6680
rect -38675 6645 -38665 6680
rect -38630 6645 -38620 6680
rect -38585 6645 -38575 6680
rect -38540 6645 -38530 6680
rect -38495 6645 -38485 6680
rect -38450 6645 -38440 6680
rect -38405 6645 -38395 6680
rect -38360 6645 -38350 6680
rect -38315 6645 -38305 6680
rect -38270 6645 -38260 6680
rect -38225 6645 -38215 6680
rect -38180 6645 -38170 6680
rect -38135 6645 -38125 6680
rect -38090 6645 -38080 6680
rect -38045 6645 -38035 6680
rect -38000 6645 -37990 6680
rect -37955 6645 -37945 6680
rect -37910 6645 -37900 6680
rect -37865 6645 -37855 6680
rect -37820 6645 -37810 6680
rect -37775 6645 -37765 6680
rect -37730 6645 -37720 6680
rect -37685 6645 -37675 6680
rect -37640 6645 -37630 6680
rect -37595 6645 -37585 6680
rect -37550 6645 -37540 6680
rect -37505 6645 -37495 6680
rect -37460 6645 -37450 6680
rect -37415 6645 -37405 6680
rect -37370 6645 -37360 6680
rect -37325 6645 -37315 6680
rect -37280 6645 -37270 6680
rect -37235 6645 -37225 6680
rect -37190 6665 -80 6680
rect -40 6665 270 6705
rect 310 6665 620 6705
rect 660 6665 970 6705
rect 1010 6665 1670 6705
rect 1710 6665 2245 6705
rect 2285 6665 3175 6705
rect 3215 6665 3235 6705
rect 3275 6665 3345 6705
rect 3385 6665 6700 6705
rect 6740 6665 7270 6705
rect 7310 6665 7970 6705
rect 8010 6665 8320 6705
rect 8360 6665 8670 6705
rect 8710 6665 9020 6705
rect 9060 6665 9100 6705
rect -37190 6645 9100 6665
rect -38770 6635 9100 6645
rect -38770 6600 -38755 6635
rect -38720 6600 -38710 6635
rect -38675 6600 -38665 6635
rect -38630 6600 -38620 6635
rect -38585 6600 -38575 6635
rect -38540 6600 -38530 6635
rect -38495 6600 -38485 6635
rect -38450 6600 -38440 6635
rect -38405 6600 -38395 6635
rect -38360 6600 -38350 6635
rect -38315 6600 -38305 6635
rect -38270 6600 -38260 6635
rect -38225 6600 -38215 6635
rect -38180 6600 -38170 6635
rect -38135 6600 -38125 6635
rect -38090 6600 -38080 6635
rect -38045 6600 -38035 6635
rect -38000 6600 -37990 6635
rect -37955 6600 -37945 6635
rect -37910 6600 -37900 6635
rect -37865 6600 -37855 6635
rect -37820 6600 -37810 6635
rect -37775 6600 -37765 6635
rect -37730 6600 -37720 6635
rect -37685 6600 -37675 6635
rect -37640 6600 -37630 6635
rect -37595 6600 -37585 6635
rect -37550 6600 -37540 6635
rect -37505 6600 -37495 6635
rect -37460 6600 -37450 6635
rect -37415 6600 -37405 6635
rect -37370 6600 -37360 6635
rect -37325 6600 -37315 6635
rect -37280 6600 -37270 6635
rect -37235 6600 -37225 6635
rect -37190 6600 -80 6635
rect -38770 6595 -80 6600
rect -40 6595 270 6635
rect 310 6595 620 6635
rect 660 6595 970 6635
rect 1010 6595 1670 6635
rect 1710 6595 2245 6635
rect 2285 6595 3175 6635
rect 3215 6595 3235 6635
rect 3275 6595 3345 6635
rect 3385 6595 6700 6635
rect 6740 6595 7270 6635
rect 7310 6595 7970 6635
rect 8010 6595 8320 6635
rect 8360 6595 8670 6635
rect 8710 6595 9020 6635
rect 9060 6595 9100 6635
rect -38770 6590 9100 6595
rect -38770 6555 -38755 6590
rect -38720 6555 -38710 6590
rect -38675 6555 -38665 6590
rect -38630 6555 -38620 6590
rect -38585 6555 -38575 6590
rect -38540 6555 -38530 6590
rect -38495 6555 -38485 6590
rect -38450 6555 -38440 6590
rect -38405 6555 -38395 6590
rect -38360 6555 -38350 6590
rect -38315 6555 -38305 6590
rect -38270 6555 -38260 6590
rect -38225 6555 -38215 6590
rect -38180 6555 -38170 6590
rect -38135 6555 -38125 6590
rect -38090 6555 -38080 6590
rect -38045 6555 -38035 6590
rect -38000 6555 -37990 6590
rect -37955 6555 -37945 6590
rect -37910 6555 -37900 6590
rect -37865 6555 -37855 6590
rect -37820 6555 -37810 6590
rect -37775 6555 -37765 6590
rect -37730 6555 -37720 6590
rect -37685 6555 -37675 6590
rect -37640 6555 -37630 6590
rect -37595 6555 -37585 6590
rect -37550 6555 -37540 6590
rect -37505 6555 -37495 6590
rect -37460 6555 -37450 6590
rect -37415 6555 -37405 6590
rect -37370 6555 -37360 6590
rect -37325 6555 -37315 6590
rect -37280 6555 -37270 6590
rect -37235 6555 -37225 6590
rect -37190 6565 9100 6590
rect -37190 6555 -80 6565
rect -38770 6545 -80 6555
rect -38770 6510 -38755 6545
rect -38720 6510 -38710 6545
rect -38675 6510 -38665 6545
rect -38630 6510 -38620 6545
rect -38585 6510 -38575 6545
rect -38540 6510 -38530 6545
rect -38495 6510 -38485 6545
rect -38450 6510 -38440 6545
rect -38405 6510 -38395 6545
rect -38360 6510 -38350 6545
rect -38315 6510 -38305 6545
rect -38270 6510 -38260 6545
rect -38225 6510 -38215 6545
rect -38180 6510 -38170 6545
rect -38135 6510 -38125 6545
rect -38090 6510 -38080 6545
rect -38045 6510 -38035 6545
rect -38000 6510 -37990 6545
rect -37955 6510 -37945 6545
rect -37910 6510 -37900 6545
rect -37865 6510 -37855 6545
rect -37820 6510 -37810 6545
rect -37775 6510 -37765 6545
rect -37730 6510 -37720 6545
rect -37685 6510 -37675 6545
rect -37640 6510 -37630 6545
rect -37595 6510 -37585 6545
rect -37550 6510 -37540 6545
rect -37505 6510 -37495 6545
rect -37460 6510 -37450 6545
rect -37415 6510 -37405 6545
rect -37370 6510 -37360 6545
rect -37325 6510 -37315 6545
rect -37280 6510 -37270 6545
rect -37235 6510 -37225 6545
rect -37190 6525 -80 6545
rect -40 6525 270 6565
rect 310 6525 620 6565
rect 660 6525 970 6565
rect 1010 6525 1670 6565
rect 1710 6525 2245 6565
rect 2285 6525 3175 6565
rect 3215 6525 3235 6565
rect 3275 6525 3345 6565
rect 3385 6525 6700 6565
rect 6740 6525 7270 6565
rect 7310 6525 7970 6565
rect 8010 6525 8320 6565
rect 8360 6525 8670 6565
rect 8710 6525 9020 6565
rect 9060 6525 9100 6565
rect -37190 6510 9100 6525
rect -38770 6500 9100 6510
rect -38770 6465 -38755 6500
rect -38720 6465 -38710 6500
rect -38675 6465 -38665 6500
rect -38630 6465 -38620 6500
rect -38585 6465 -38575 6500
rect -38540 6465 -38530 6500
rect -38495 6465 -38485 6500
rect -38450 6465 -38440 6500
rect -38405 6465 -38395 6500
rect -38360 6465 -38350 6500
rect -38315 6465 -38305 6500
rect -38270 6465 -38260 6500
rect -38225 6465 -38215 6500
rect -38180 6465 -38170 6500
rect -38135 6465 -38125 6500
rect -38090 6465 -38080 6500
rect -38045 6465 -38035 6500
rect -38000 6465 -37990 6500
rect -37955 6465 -37945 6500
rect -37910 6465 -37900 6500
rect -37865 6465 -37855 6500
rect -37820 6465 -37810 6500
rect -37775 6465 -37765 6500
rect -37730 6465 -37720 6500
rect -37685 6465 -37675 6500
rect -37640 6465 -37630 6500
rect -37595 6465 -37585 6500
rect -37550 6465 -37540 6500
rect -37505 6465 -37495 6500
rect -37460 6465 -37450 6500
rect -37415 6465 -37405 6500
rect -37370 6465 -37360 6500
rect -37325 6465 -37315 6500
rect -37280 6465 -37270 6500
rect -37235 6465 -37225 6500
rect -37190 6465 -80 6500
rect -38770 6460 -80 6465
rect -40 6460 270 6500
rect 310 6460 620 6500
rect 660 6460 970 6500
rect 1010 6460 1670 6500
rect 1710 6460 2245 6500
rect 2285 6460 3175 6500
rect 3215 6460 3235 6500
rect 3275 6460 3345 6500
rect 3385 6460 6700 6500
rect 6740 6460 7270 6500
rect 7310 6460 7970 6500
rect 8010 6460 8320 6500
rect 8360 6460 8670 6500
rect 8710 6460 9020 6500
rect 9060 6460 9100 6500
rect -38770 6450 9100 6460
rect 31290 8030 35620 8050
rect 31290 7995 31305 8030
rect 31340 7995 31350 8030
rect 31385 7995 31395 8030
rect 31430 7995 31440 8030
rect 31475 7995 31485 8030
rect 31520 7995 31530 8030
rect 31565 7995 31575 8030
rect 31610 7995 31620 8030
rect 31655 7995 31665 8030
rect 31700 7995 31710 8030
rect 31745 7995 31755 8030
rect 31790 7995 31800 8030
rect 31835 7995 31845 8030
rect 31880 7995 31890 8030
rect 31925 7995 31935 8030
rect 31970 7995 31980 8030
rect 32015 7995 32025 8030
rect 32060 7995 32070 8030
rect 32105 7995 32115 8030
rect 32150 7995 32160 8030
rect 32195 7995 32205 8030
rect 32240 7995 32250 8030
rect 32285 7995 32295 8030
rect 32330 7995 32340 8030
rect 32375 7995 32385 8030
rect 32420 7995 32430 8030
rect 32465 7995 32475 8030
rect 32510 7995 32520 8030
rect 32555 7995 32565 8030
rect 32600 7995 32610 8030
rect 32645 7995 32655 8030
rect 32690 7995 32700 8030
rect 32735 7995 32745 8030
rect 32780 7995 32790 8030
rect 32825 7995 32835 8030
rect 32870 7995 35620 8030
rect 31290 7985 35620 7995
rect 31290 7950 31305 7985
rect 31340 7950 31350 7985
rect 31385 7950 31395 7985
rect 31430 7950 31440 7985
rect 31475 7950 31485 7985
rect 31520 7950 31530 7985
rect 31565 7950 31575 7985
rect 31610 7950 31620 7985
rect 31655 7950 31665 7985
rect 31700 7950 31710 7985
rect 31745 7950 31755 7985
rect 31790 7950 31800 7985
rect 31835 7950 31845 7985
rect 31880 7950 31890 7985
rect 31925 7950 31935 7985
rect 31970 7950 31980 7985
rect 32015 7950 32025 7985
rect 32060 7950 32070 7985
rect 32105 7950 32115 7985
rect 32150 7950 32160 7985
rect 32195 7950 32205 7985
rect 32240 7950 32250 7985
rect 32285 7950 32295 7985
rect 32330 7950 32340 7985
rect 32375 7950 32385 7985
rect 32420 7950 32430 7985
rect 32465 7950 32475 7985
rect 32510 7950 32520 7985
rect 32555 7950 32565 7985
rect 32600 7950 32610 7985
rect 32645 7950 32655 7985
rect 32690 7950 32700 7985
rect 32735 7950 32745 7985
rect 32780 7950 32790 7985
rect 32825 7950 32835 7985
rect 32870 7950 35620 7985
rect 31290 7940 35620 7950
rect 31290 7905 31305 7940
rect 31340 7905 31350 7940
rect 31385 7905 31395 7940
rect 31430 7905 31440 7940
rect 31475 7905 31485 7940
rect 31520 7905 31530 7940
rect 31565 7905 31575 7940
rect 31610 7905 31620 7940
rect 31655 7905 31665 7940
rect 31700 7905 31710 7940
rect 31745 7905 31755 7940
rect 31790 7905 31800 7940
rect 31835 7905 31845 7940
rect 31880 7905 31890 7940
rect 31925 7905 31935 7940
rect 31970 7905 31980 7940
rect 32015 7905 32025 7940
rect 32060 7905 32070 7940
rect 32105 7905 32115 7940
rect 32150 7905 32160 7940
rect 32195 7905 32205 7940
rect 32240 7905 32250 7940
rect 32285 7905 32295 7940
rect 32330 7905 32340 7940
rect 32375 7905 32385 7940
rect 32420 7905 32430 7940
rect 32465 7905 32475 7940
rect 32510 7905 32520 7940
rect 32555 7905 32565 7940
rect 32600 7905 32610 7940
rect 32645 7905 32655 7940
rect 32690 7905 32700 7940
rect 32735 7905 32745 7940
rect 32780 7905 32790 7940
rect 32825 7905 32835 7940
rect 32870 7905 35620 7940
rect 31290 7895 35620 7905
rect 31290 7860 31305 7895
rect 31340 7860 31350 7895
rect 31385 7860 31395 7895
rect 31430 7860 31440 7895
rect 31475 7860 31485 7895
rect 31520 7860 31530 7895
rect 31565 7860 31575 7895
rect 31610 7860 31620 7895
rect 31655 7860 31665 7895
rect 31700 7860 31710 7895
rect 31745 7860 31755 7895
rect 31790 7860 31800 7895
rect 31835 7860 31845 7895
rect 31880 7860 31890 7895
rect 31925 7860 31935 7895
rect 31970 7860 31980 7895
rect 32015 7860 32025 7895
rect 32060 7860 32070 7895
rect 32105 7860 32115 7895
rect 32150 7860 32160 7895
rect 32195 7860 32205 7895
rect 32240 7860 32250 7895
rect 32285 7860 32295 7895
rect 32330 7860 32340 7895
rect 32375 7860 32385 7895
rect 32420 7860 32430 7895
rect 32465 7860 32475 7895
rect 32510 7860 32520 7895
rect 32555 7860 32565 7895
rect 32600 7860 32610 7895
rect 32645 7860 32655 7895
rect 32690 7860 32700 7895
rect 32735 7860 32745 7895
rect 32780 7860 32790 7895
rect 32825 7860 32835 7895
rect 32870 7860 35620 7895
rect 31290 7850 35620 7860
rect 31290 7815 31305 7850
rect 31340 7815 31350 7850
rect 31385 7815 31395 7850
rect 31430 7815 31440 7850
rect 31475 7815 31485 7850
rect 31520 7815 31530 7850
rect 31565 7815 31575 7850
rect 31610 7815 31620 7850
rect 31655 7815 31665 7850
rect 31700 7815 31710 7850
rect 31745 7815 31755 7850
rect 31790 7815 31800 7850
rect 31835 7815 31845 7850
rect 31880 7815 31890 7850
rect 31925 7815 31935 7850
rect 31970 7815 31980 7850
rect 32015 7815 32025 7850
rect 32060 7815 32070 7850
rect 32105 7815 32115 7850
rect 32150 7815 32160 7850
rect 32195 7815 32205 7850
rect 32240 7815 32250 7850
rect 32285 7815 32295 7850
rect 32330 7815 32340 7850
rect 32375 7815 32385 7850
rect 32420 7815 32430 7850
rect 32465 7815 32475 7850
rect 32510 7815 32520 7850
rect 32555 7815 32565 7850
rect 32600 7815 32610 7850
rect 32645 7815 32655 7850
rect 32690 7815 32700 7850
rect 32735 7815 32745 7850
rect 32780 7815 32790 7850
rect 32825 7815 32835 7850
rect 32870 7815 35620 7850
rect 31290 7805 35620 7815
rect 31290 7770 31305 7805
rect 31340 7770 31350 7805
rect 31385 7770 31395 7805
rect 31430 7770 31440 7805
rect 31475 7770 31485 7805
rect 31520 7770 31530 7805
rect 31565 7770 31575 7805
rect 31610 7770 31620 7805
rect 31655 7770 31665 7805
rect 31700 7770 31710 7805
rect 31745 7770 31755 7805
rect 31790 7770 31800 7805
rect 31835 7770 31845 7805
rect 31880 7770 31890 7805
rect 31925 7770 31935 7805
rect 31970 7770 31980 7805
rect 32015 7770 32025 7805
rect 32060 7770 32070 7805
rect 32105 7770 32115 7805
rect 32150 7770 32160 7805
rect 32195 7770 32205 7805
rect 32240 7770 32250 7805
rect 32285 7770 32295 7805
rect 32330 7770 32340 7805
rect 32375 7770 32385 7805
rect 32420 7770 32430 7805
rect 32465 7770 32475 7805
rect 32510 7770 32520 7805
rect 32555 7770 32565 7805
rect 32600 7770 32610 7805
rect 32645 7770 32655 7805
rect 32690 7770 32700 7805
rect 32735 7770 32745 7805
rect 32780 7770 32790 7805
rect 32825 7770 32835 7805
rect 32870 7770 35620 7805
rect 31290 7760 35620 7770
rect 31290 7725 31305 7760
rect 31340 7725 31350 7760
rect 31385 7725 31395 7760
rect 31430 7725 31440 7760
rect 31475 7725 31485 7760
rect 31520 7725 31530 7760
rect 31565 7725 31575 7760
rect 31610 7725 31620 7760
rect 31655 7725 31665 7760
rect 31700 7725 31710 7760
rect 31745 7725 31755 7760
rect 31790 7725 31800 7760
rect 31835 7725 31845 7760
rect 31880 7725 31890 7760
rect 31925 7725 31935 7760
rect 31970 7725 31980 7760
rect 32015 7725 32025 7760
rect 32060 7725 32070 7760
rect 32105 7725 32115 7760
rect 32150 7725 32160 7760
rect 32195 7725 32205 7760
rect 32240 7725 32250 7760
rect 32285 7725 32295 7760
rect 32330 7725 32340 7760
rect 32375 7725 32385 7760
rect 32420 7725 32430 7760
rect 32465 7725 32475 7760
rect 32510 7725 32520 7760
rect 32555 7725 32565 7760
rect 32600 7725 32610 7760
rect 32645 7725 32655 7760
rect 32690 7725 32700 7760
rect 32735 7725 32745 7760
rect 32780 7725 32790 7760
rect 32825 7725 32835 7760
rect 32870 7725 35620 7760
rect 31290 7715 35620 7725
rect 31290 7680 31305 7715
rect 31340 7680 31350 7715
rect 31385 7680 31395 7715
rect 31430 7680 31440 7715
rect 31475 7680 31485 7715
rect 31520 7680 31530 7715
rect 31565 7680 31575 7715
rect 31610 7680 31620 7715
rect 31655 7680 31665 7715
rect 31700 7680 31710 7715
rect 31745 7680 31755 7715
rect 31790 7680 31800 7715
rect 31835 7680 31845 7715
rect 31880 7680 31890 7715
rect 31925 7680 31935 7715
rect 31970 7680 31980 7715
rect 32015 7680 32025 7715
rect 32060 7680 32070 7715
rect 32105 7680 32115 7715
rect 32150 7680 32160 7715
rect 32195 7680 32205 7715
rect 32240 7680 32250 7715
rect 32285 7680 32295 7715
rect 32330 7680 32340 7715
rect 32375 7680 32385 7715
rect 32420 7680 32430 7715
rect 32465 7680 32475 7715
rect 32510 7680 32520 7715
rect 32555 7680 32565 7715
rect 32600 7680 32610 7715
rect 32645 7680 32655 7715
rect 32690 7680 32700 7715
rect 32735 7680 32745 7715
rect 32780 7680 32790 7715
rect 32825 7680 32835 7715
rect 32870 7680 35620 7715
rect 31290 7670 35620 7680
rect 31290 7635 31305 7670
rect 31340 7635 31350 7670
rect 31385 7635 31395 7670
rect 31430 7635 31440 7670
rect 31475 7635 31485 7670
rect 31520 7635 31530 7670
rect 31565 7635 31575 7670
rect 31610 7635 31620 7670
rect 31655 7635 31665 7670
rect 31700 7635 31710 7670
rect 31745 7635 31755 7670
rect 31790 7635 31800 7670
rect 31835 7635 31845 7670
rect 31880 7635 31890 7670
rect 31925 7635 31935 7670
rect 31970 7635 31980 7670
rect 32015 7635 32025 7670
rect 32060 7635 32070 7670
rect 32105 7635 32115 7670
rect 32150 7635 32160 7670
rect 32195 7635 32205 7670
rect 32240 7635 32250 7670
rect 32285 7635 32295 7670
rect 32330 7635 32340 7670
rect 32375 7635 32385 7670
rect 32420 7635 32430 7670
rect 32465 7635 32475 7670
rect 32510 7635 32520 7670
rect 32555 7635 32565 7670
rect 32600 7635 32610 7670
rect 32645 7635 32655 7670
rect 32690 7635 32700 7670
rect 32735 7635 32745 7670
rect 32780 7635 32790 7670
rect 32825 7635 32835 7670
rect 32870 7635 35620 7670
rect 31290 7625 35620 7635
rect 31290 7590 31305 7625
rect 31340 7590 31350 7625
rect 31385 7590 31395 7625
rect 31430 7590 31440 7625
rect 31475 7590 31485 7625
rect 31520 7590 31530 7625
rect 31565 7590 31575 7625
rect 31610 7590 31620 7625
rect 31655 7590 31665 7625
rect 31700 7590 31710 7625
rect 31745 7590 31755 7625
rect 31790 7590 31800 7625
rect 31835 7590 31845 7625
rect 31880 7590 31890 7625
rect 31925 7590 31935 7625
rect 31970 7590 31980 7625
rect 32015 7590 32025 7625
rect 32060 7590 32070 7625
rect 32105 7590 32115 7625
rect 32150 7590 32160 7625
rect 32195 7590 32205 7625
rect 32240 7590 32250 7625
rect 32285 7590 32295 7625
rect 32330 7590 32340 7625
rect 32375 7590 32385 7625
rect 32420 7590 32430 7625
rect 32465 7590 32475 7625
rect 32510 7590 32520 7625
rect 32555 7590 32565 7625
rect 32600 7590 32610 7625
rect 32645 7590 32655 7625
rect 32690 7590 32700 7625
rect 32735 7590 32745 7625
rect 32780 7590 32790 7625
rect 32825 7590 32835 7625
rect 32870 7590 35620 7625
rect 31290 7580 35620 7590
rect 31290 7545 31305 7580
rect 31340 7545 31350 7580
rect 31385 7545 31395 7580
rect 31430 7545 31440 7580
rect 31475 7545 31485 7580
rect 31520 7545 31530 7580
rect 31565 7545 31575 7580
rect 31610 7545 31620 7580
rect 31655 7545 31665 7580
rect 31700 7545 31710 7580
rect 31745 7545 31755 7580
rect 31790 7545 31800 7580
rect 31835 7545 31845 7580
rect 31880 7545 31890 7580
rect 31925 7545 31935 7580
rect 31970 7545 31980 7580
rect 32015 7545 32025 7580
rect 32060 7545 32070 7580
rect 32105 7545 32115 7580
rect 32150 7545 32160 7580
rect 32195 7545 32205 7580
rect 32240 7545 32250 7580
rect 32285 7545 32295 7580
rect 32330 7545 32340 7580
rect 32375 7545 32385 7580
rect 32420 7545 32430 7580
rect 32465 7545 32475 7580
rect 32510 7545 32520 7580
rect 32555 7545 32565 7580
rect 32600 7545 32610 7580
rect 32645 7545 32655 7580
rect 32690 7545 32700 7580
rect 32735 7545 32745 7580
rect 32780 7545 32790 7580
rect 32825 7545 32835 7580
rect 32870 7545 35620 7580
rect 31290 7535 35620 7545
rect 31290 7500 31305 7535
rect 31340 7500 31350 7535
rect 31385 7500 31395 7535
rect 31430 7500 31440 7535
rect 31475 7500 31485 7535
rect 31520 7500 31530 7535
rect 31565 7500 31575 7535
rect 31610 7500 31620 7535
rect 31655 7500 31665 7535
rect 31700 7500 31710 7535
rect 31745 7500 31755 7535
rect 31790 7500 31800 7535
rect 31835 7500 31845 7535
rect 31880 7500 31890 7535
rect 31925 7500 31935 7535
rect 31970 7500 31980 7535
rect 32015 7500 32025 7535
rect 32060 7500 32070 7535
rect 32105 7500 32115 7535
rect 32150 7500 32160 7535
rect 32195 7500 32205 7535
rect 32240 7500 32250 7535
rect 32285 7500 32295 7535
rect 32330 7500 32340 7535
rect 32375 7500 32385 7535
rect 32420 7500 32430 7535
rect 32465 7500 32475 7535
rect 32510 7500 32520 7535
rect 32555 7500 32565 7535
rect 32600 7500 32610 7535
rect 32645 7500 32655 7535
rect 32690 7500 32700 7535
rect 32735 7500 32745 7535
rect 32780 7500 32790 7535
rect 32825 7500 32835 7535
rect 32870 7500 35620 7535
rect 31290 7490 35620 7500
rect 31290 7455 31305 7490
rect 31340 7455 31350 7490
rect 31385 7455 31395 7490
rect 31430 7455 31440 7490
rect 31475 7455 31485 7490
rect 31520 7455 31530 7490
rect 31565 7455 31575 7490
rect 31610 7455 31620 7490
rect 31655 7455 31665 7490
rect 31700 7455 31710 7490
rect 31745 7455 31755 7490
rect 31790 7455 31800 7490
rect 31835 7455 31845 7490
rect 31880 7455 31890 7490
rect 31925 7455 31935 7490
rect 31970 7455 31980 7490
rect 32015 7455 32025 7490
rect 32060 7455 32070 7490
rect 32105 7455 32115 7490
rect 32150 7455 32160 7490
rect 32195 7455 32205 7490
rect 32240 7455 32250 7490
rect 32285 7455 32295 7490
rect 32330 7455 32340 7490
rect 32375 7455 32385 7490
rect 32420 7455 32430 7490
rect 32465 7455 32475 7490
rect 32510 7455 32520 7490
rect 32555 7455 32565 7490
rect 32600 7455 32610 7490
rect 32645 7455 32655 7490
rect 32690 7455 32700 7490
rect 32735 7455 32745 7490
rect 32780 7455 32790 7490
rect 32825 7455 32835 7490
rect 32870 7455 35620 7490
rect 31290 7445 35620 7455
rect 31290 7410 31305 7445
rect 31340 7410 31350 7445
rect 31385 7410 31395 7445
rect 31430 7410 31440 7445
rect 31475 7410 31485 7445
rect 31520 7410 31530 7445
rect 31565 7410 31575 7445
rect 31610 7410 31620 7445
rect 31655 7410 31665 7445
rect 31700 7410 31710 7445
rect 31745 7410 31755 7445
rect 31790 7410 31800 7445
rect 31835 7410 31845 7445
rect 31880 7410 31890 7445
rect 31925 7410 31935 7445
rect 31970 7410 31980 7445
rect 32015 7410 32025 7445
rect 32060 7410 32070 7445
rect 32105 7410 32115 7445
rect 32150 7410 32160 7445
rect 32195 7410 32205 7445
rect 32240 7410 32250 7445
rect 32285 7410 32295 7445
rect 32330 7410 32340 7445
rect 32375 7410 32385 7445
rect 32420 7410 32430 7445
rect 32465 7410 32475 7445
rect 32510 7410 32520 7445
rect 32555 7410 32565 7445
rect 32600 7410 32610 7445
rect 32645 7410 32655 7445
rect 32690 7410 32700 7445
rect 32735 7410 32745 7445
rect 32780 7410 32790 7445
rect 32825 7410 32835 7445
rect 32870 7410 35620 7445
rect 31290 7400 35620 7410
rect 31290 7365 31305 7400
rect 31340 7365 31350 7400
rect 31385 7365 31395 7400
rect 31430 7365 31440 7400
rect 31475 7365 31485 7400
rect 31520 7365 31530 7400
rect 31565 7365 31575 7400
rect 31610 7365 31620 7400
rect 31655 7365 31665 7400
rect 31700 7365 31710 7400
rect 31745 7365 31755 7400
rect 31790 7365 31800 7400
rect 31835 7365 31845 7400
rect 31880 7365 31890 7400
rect 31925 7365 31935 7400
rect 31970 7365 31980 7400
rect 32015 7365 32025 7400
rect 32060 7365 32070 7400
rect 32105 7365 32115 7400
rect 32150 7365 32160 7400
rect 32195 7365 32205 7400
rect 32240 7365 32250 7400
rect 32285 7365 32295 7400
rect 32330 7365 32340 7400
rect 32375 7365 32385 7400
rect 32420 7365 32430 7400
rect 32465 7365 32475 7400
rect 32510 7365 32520 7400
rect 32555 7365 32565 7400
rect 32600 7365 32610 7400
rect 32645 7365 32655 7400
rect 32690 7365 32700 7400
rect 32735 7365 32745 7400
rect 32780 7365 32790 7400
rect 32825 7365 32835 7400
rect 32870 7365 35620 7400
rect 31290 7355 35620 7365
rect 31290 7320 31305 7355
rect 31340 7320 31350 7355
rect 31385 7320 31395 7355
rect 31430 7320 31440 7355
rect 31475 7320 31485 7355
rect 31520 7320 31530 7355
rect 31565 7320 31575 7355
rect 31610 7320 31620 7355
rect 31655 7320 31665 7355
rect 31700 7320 31710 7355
rect 31745 7320 31755 7355
rect 31790 7320 31800 7355
rect 31835 7320 31845 7355
rect 31880 7320 31890 7355
rect 31925 7320 31935 7355
rect 31970 7320 31980 7355
rect 32015 7320 32025 7355
rect 32060 7320 32070 7355
rect 32105 7320 32115 7355
rect 32150 7320 32160 7355
rect 32195 7320 32205 7355
rect 32240 7320 32250 7355
rect 32285 7320 32295 7355
rect 32330 7320 32340 7355
rect 32375 7320 32385 7355
rect 32420 7320 32430 7355
rect 32465 7320 32475 7355
rect 32510 7320 32520 7355
rect 32555 7320 32565 7355
rect 32600 7320 32610 7355
rect 32645 7320 32655 7355
rect 32690 7320 32700 7355
rect 32735 7320 32745 7355
rect 32780 7320 32790 7355
rect 32825 7320 32835 7355
rect 32870 7320 35620 7355
rect 31290 7310 35620 7320
rect 31290 7275 31305 7310
rect 31340 7275 31350 7310
rect 31385 7275 31395 7310
rect 31430 7275 31440 7310
rect 31475 7275 31485 7310
rect 31520 7275 31530 7310
rect 31565 7275 31575 7310
rect 31610 7275 31620 7310
rect 31655 7275 31665 7310
rect 31700 7275 31710 7310
rect 31745 7275 31755 7310
rect 31790 7275 31800 7310
rect 31835 7275 31845 7310
rect 31880 7275 31890 7310
rect 31925 7275 31935 7310
rect 31970 7275 31980 7310
rect 32015 7275 32025 7310
rect 32060 7275 32070 7310
rect 32105 7275 32115 7310
rect 32150 7275 32160 7310
rect 32195 7275 32205 7310
rect 32240 7275 32250 7310
rect 32285 7275 32295 7310
rect 32330 7275 32340 7310
rect 32375 7275 32385 7310
rect 32420 7275 32430 7310
rect 32465 7275 32475 7310
rect 32510 7275 32520 7310
rect 32555 7275 32565 7310
rect 32600 7275 32610 7310
rect 32645 7275 32655 7310
rect 32690 7275 32700 7310
rect 32735 7275 32745 7310
rect 32780 7275 32790 7310
rect 32825 7275 32835 7310
rect 32870 7275 35620 7310
rect 31290 7265 35620 7275
rect 31290 7230 31305 7265
rect 31340 7230 31350 7265
rect 31385 7230 31395 7265
rect 31430 7230 31440 7265
rect 31475 7230 31485 7265
rect 31520 7230 31530 7265
rect 31565 7230 31575 7265
rect 31610 7230 31620 7265
rect 31655 7230 31665 7265
rect 31700 7230 31710 7265
rect 31745 7230 31755 7265
rect 31790 7230 31800 7265
rect 31835 7230 31845 7265
rect 31880 7230 31890 7265
rect 31925 7230 31935 7265
rect 31970 7230 31980 7265
rect 32015 7230 32025 7265
rect 32060 7230 32070 7265
rect 32105 7230 32115 7265
rect 32150 7230 32160 7265
rect 32195 7230 32205 7265
rect 32240 7230 32250 7265
rect 32285 7230 32295 7265
rect 32330 7230 32340 7265
rect 32375 7230 32385 7265
rect 32420 7230 32430 7265
rect 32465 7230 32475 7265
rect 32510 7230 32520 7265
rect 32555 7230 32565 7265
rect 32600 7230 32610 7265
rect 32645 7230 32655 7265
rect 32690 7230 32700 7265
rect 32735 7230 32745 7265
rect 32780 7230 32790 7265
rect 32825 7230 32835 7265
rect 32870 7230 35620 7265
rect 31290 7220 35620 7230
rect 31290 7185 31305 7220
rect 31340 7185 31350 7220
rect 31385 7185 31395 7220
rect 31430 7185 31440 7220
rect 31475 7185 31485 7220
rect 31520 7185 31530 7220
rect 31565 7185 31575 7220
rect 31610 7185 31620 7220
rect 31655 7185 31665 7220
rect 31700 7185 31710 7220
rect 31745 7185 31755 7220
rect 31790 7185 31800 7220
rect 31835 7185 31845 7220
rect 31880 7185 31890 7220
rect 31925 7185 31935 7220
rect 31970 7185 31980 7220
rect 32015 7185 32025 7220
rect 32060 7185 32070 7220
rect 32105 7185 32115 7220
rect 32150 7185 32160 7220
rect 32195 7185 32205 7220
rect 32240 7185 32250 7220
rect 32285 7185 32295 7220
rect 32330 7185 32340 7220
rect 32375 7185 32385 7220
rect 32420 7185 32430 7220
rect 32465 7185 32475 7220
rect 32510 7185 32520 7220
rect 32555 7185 32565 7220
rect 32600 7185 32610 7220
rect 32645 7185 32655 7220
rect 32690 7185 32700 7220
rect 32735 7185 32745 7220
rect 32780 7185 32790 7220
rect 32825 7185 32835 7220
rect 32870 7185 35620 7220
rect 31290 7175 35620 7185
rect 31290 7140 31305 7175
rect 31340 7140 31350 7175
rect 31385 7140 31395 7175
rect 31430 7140 31440 7175
rect 31475 7140 31485 7175
rect 31520 7140 31530 7175
rect 31565 7140 31575 7175
rect 31610 7140 31620 7175
rect 31655 7140 31665 7175
rect 31700 7140 31710 7175
rect 31745 7140 31755 7175
rect 31790 7140 31800 7175
rect 31835 7140 31845 7175
rect 31880 7140 31890 7175
rect 31925 7140 31935 7175
rect 31970 7140 31980 7175
rect 32015 7140 32025 7175
rect 32060 7140 32070 7175
rect 32105 7140 32115 7175
rect 32150 7140 32160 7175
rect 32195 7140 32205 7175
rect 32240 7140 32250 7175
rect 32285 7140 32295 7175
rect 32330 7140 32340 7175
rect 32375 7140 32385 7175
rect 32420 7140 32430 7175
rect 32465 7140 32475 7175
rect 32510 7140 32520 7175
rect 32555 7140 32565 7175
rect 32600 7140 32610 7175
rect 32645 7140 32655 7175
rect 32690 7140 32700 7175
rect 32735 7140 32745 7175
rect 32780 7140 32790 7175
rect 32825 7140 32835 7175
rect 32870 7140 35620 7175
rect 31290 7130 35620 7140
rect 31290 7095 31305 7130
rect 31340 7095 31350 7130
rect 31385 7095 31395 7130
rect 31430 7095 31440 7130
rect 31475 7095 31485 7130
rect 31520 7095 31530 7130
rect 31565 7095 31575 7130
rect 31610 7095 31620 7130
rect 31655 7095 31665 7130
rect 31700 7095 31710 7130
rect 31745 7095 31755 7130
rect 31790 7095 31800 7130
rect 31835 7095 31845 7130
rect 31880 7095 31890 7130
rect 31925 7095 31935 7130
rect 31970 7095 31980 7130
rect 32015 7095 32025 7130
rect 32060 7095 32070 7130
rect 32105 7095 32115 7130
rect 32150 7095 32160 7130
rect 32195 7095 32205 7130
rect 32240 7095 32250 7130
rect 32285 7095 32295 7130
rect 32330 7095 32340 7130
rect 32375 7095 32385 7130
rect 32420 7095 32430 7130
rect 32465 7095 32475 7130
rect 32510 7095 32520 7130
rect 32555 7095 32565 7130
rect 32600 7095 32610 7130
rect 32645 7095 32655 7130
rect 32690 7095 32700 7130
rect 32735 7095 32745 7130
rect 32780 7095 32790 7130
rect 32825 7095 32835 7130
rect 32870 7095 35620 7130
rect 31290 7085 35620 7095
rect 31290 7050 31305 7085
rect 31340 7050 31350 7085
rect 31385 7050 31395 7085
rect 31430 7050 31440 7085
rect 31475 7050 31485 7085
rect 31520 7050 31530 7085
rect 31565 7050 31575 7085
rect 31610 7050 31620 7085
rect 31655 7050 31665 7085
rect 31700 7050 31710 7085
rect 31745 7050 31755 7085
rect 31790 7050 31800 7085
rect 31835 7050 31845 7085
rect 31880 7050 31890 7085
rect 31925 7050 31935 7085
rect 31970 7050 31980 7085
rect 32015 7050 32025 7085
rect 32060 7050 32070 7085
rect 32105 7050 32115 7085
rect 32150 7050 32160 7085
rect 32195 7050 32205 7085
rect 32240 7050 32250 7085
rect 32285 7050 32295 7085
rect 32330 7050 32340 7085
rect 32375 7050 32385 7085
rect 32420 7050 32430 7085
rect 32465 7050 32475 7085
rect 32510 7050 32520 7085
rect 32555 7050 32565 7085
rect 32600 7050 32610 7085
rect 32645 7050 32655 7085
rect 32690 7050 32700 7085
rect 32735 7050 32745 7085
rect 32780 7050 32790 7085
rect 32825 7050 32835 7085
rect 32870 7050 35620 7085
rect 31290 7040 35620 7050
rect 31290 7005 31305 7040
rect 31340 7005 31350 7040
rect 31385 7005 31395 7040
rect 31430 7005 31440 7040
rect 31475 7005 31485 7040
rect 31520 7005 31530 7040
rect 31565 7005 31575 7040
rect 31610 7005 31620 7040
rect 31655 7005 31665 7040
rect 31700 7005 31710 7040
rect 31745 7005 31755 7040
rect 31790 7005 31800 7040
rect 31835 7005 31845 7040
rect 31880 7005 31890 7040
rect 31925 7005 31935 7040
rect 31970 7005 31980 7040
rect 32015 7005 32025 7040
rect 32060 7005 32070 7040
rect 32105 7005 32115 7040
rect 32150 7005 32160 7040
rect 32195 7005 32205 7040
rect 32240 7005 32250 7040
rect 32285 7005 32295 7040
rect 32330 7005 32340 7040
rect 32375 7005 32385 7040
rect 32420 7005 32430 7040
rect 32465 7005 32475 7040
rect 32510 7005 32520 7040
rect 32555 7005 32565 7040
rect 32600 7005 32610 7040
rect 32645 7005 32655 7040
rect 32690 7005 32700 7040
rect 32735 7005 32745 7040
rect 32780 7005 32790 7040
rect 32825 7005 32835 7040
rect 32870 7005 35620 7040
rect 31290 6995 35620 7005
rect 31290 6960 31305 6995
rect 31340 6960 31350 6995
rect 31385 6960 31395 6995
rect 31430 6960 31440 6995
rect 31475 6960 31485 6995
rect 31520 6960 31530 6995
rect 31565 6960 31575 6995
rect 31610 6960 31620 6995
rect 31655 6960 31665 6995
rect 31700 6960 31710 6995
rect 31745 6960 31755 6995
rect 31790 6960 31800 6995
rect 31835 6960 31845 6995
rect 31880 6960 31890 6995
rect 31925 6960 31935 6995
rect 31970 6960 31980 6995
rect 32015 6960 32025 6995
rect 32060 6960 32070 6995
rect 32105 6960 32115 6995
rect 32150 6960 32160 6995
rect 32195 6960 32205 6995
rect 32240 6960 32250 6995
rect 32285 6960 32295 6995
rect 32330 6960 32340 6995
rect 32375 6960 32385 6995
rect 32420 6960 32430 6995
rect 32465 6960 32475 6995
rect 32510 6960 32520 6995
rect 32555 6960 32565 6995
rect 32600 6960 32610 6995
rect 32645 6960 32655 6995
rect 32690 6960 32700 6995
rect 32735 6960 32745 6995
rect 32780 6960 32790 6995
rect 32825 6960 32835 6995
rect 32870 6960 35620 6995
rect 31290 6950 35620 6960
rect 31290 6915 31305 6950
rect 31340 6915 31350 6950
rect 31385 6915 31395 6950
rect 31430 6915 31440 6950
rect 31475 6915 31485 6950
rect 31520 6915 31530 6950
rect 31565 6915 31575 6950
rect 31610 6915 31620 6950
rect 31655 6915 31665 6950
rect 31700 6915 31710 6950
rect 31745 6915 31755 6950
rect 31790 6915 31800 6950
rect 31835 6915 31845 6950
rect 31880 6915 31890 6950
rect 31925 6915 31935 6950
rect 31970 6915 31980 6950
rect 32015 6915 32025 6950
rect 32060 6915 32070 6950
rect 32105 6915 32115 6950
rect 32150 6915 32160 6950
rect 32195 6915 32205 6950
rect 32240 6915 32250 6950
rect 32285 6915 32295 6950
rect 32330 6915 32340 6950
rect 32375 6915 32385 6950
rect 32420 6915 32430 6950
rect 32465 6915 32475 6950
rect 32510 6915 32520 6950
rect 32555 6915 32565 6950
rect 32600 6915 32610 6950
rect 32645 6915 32655 6950
rect 32690 6915 32700 6950
rect 32735 6915 32745 6950
rect 32780 6915 32790 6950
rect 32825 6915 32835 6950
rect 32870 6915 35620 6950
rect 31290 6905 35620 6915
rect 31290 6870 31305 6905
rect 31340 6870 31350 6905
rect 31385 6870 31395 6905
rect 31430 6870 31440 6905
rect 31475 6870 31485 6905
rect 31520 6870 31530 6905
rect 31565 6870 31575 6905
rect 31610 6870 31620 6905
rect 31655 6870 31665 6905
rect 31700 6870 31710 6905
rect 31745 6870 31755 6905
rect 31790 6870 31800 6905
rect 31835 6870 31845 6905
rect 31880 6870 31890 6905
rect 31925 6870 31935 6905
rect 31970 6870 31980 6905
rect 32015 6870 32025 6905
rect 32060 6870 32070 6905
rect 32105 6870 32115 6905
rect 32150 6870 32160 6905
rect 32195 6870 32205 6905
rect 32240 6870 32250 6905
rect 32285 6870 32295 6905
rect 32330 6870 32340 6905
rect 32375 6870 32385 6905
rect 32420 6870 32430 6905
rect 32465 6870 32475 6905
rect 32510 6870 32520 6905
rect 32555 6870 32565 6905
rect 32600 6870 32610 6905
rect 32645 6870 32655 6905
rect 32690 6870 32700 6905
rect 32735 6870 32745 6905
rect 32780 6870 32790 6905
rect 32825 6870 32835 6905
rect 32870 6870 35620 6905
rect 31290 6860 35620 6870
rect 31290 6825 31305 6860
rect 31340 6825 31350 6860
rect 31385 6825 31395 6860
rect 31430 6825 31440 6860
rect 31475 6825 31485 6860
rect 31520 6825 31530 6860
rect 31565 6825 31575 6860
rect 31610 6825 31620 6860
rect 31655 6825 31665 6860
rect 31700 6825 31710 6860
rect 31745 6825 31755 6860
rect 31790 6825 31800 6860
rect 31835 6825 31845 6860
rect 31880 6825 31890 6860
rect 31925 6825 31935 6860
rect 31970 6825 31980 6860
rect 32015 6825 32025 6860
rect 32060 6825 32070 6860
rect 32105 6825 32115 6860
rect 32150 6825 32160 6860
rect 32195 6825 32205 6860
rect 32240 6825 32250 6860
rect 32285 6825 32295 6860
rect 32330 6825 32340 6860
rect 32375 6825 32385 6860
rect 32420 6825 32430 6860
rect 32465 6825 32475 6860
rect 32510 6825 32520 6860
rect 32555 6825 32565 6860
rect 32600 6825 32610 6860
rect 32645 6825 32655 6860
rect 32690 6825 32700 6860
rect 32735 6825 32745 6860
rect 32780 6825 32790 6860
rect 32825 6825 32835 6860
rect 32870 6825 35620 6860
rect 31290 6815 35620 6825
rect 31290 6780 31305 6815
rect 31340 6780 31350 6815
rect 31385 6780 31395 6815
rect 31430 6780 31440 6815
rect 31475 6780 31485 6815
rect 31520 6780 31530 6815
rect 31565 6780 31575 6815
rect 31610 6780 31620 6815
rect 31655 6780 31665 6815
rect 31700 6780 31710 6815
rect 31745 6780 31755 6815
rect 31790 6780 31800 6815
rect 31835 6780 31845 6815
rect 31880 6780 31890 6815
rect 31925 6780 31935 6815
rect 31970 6780 31980 6815
rect 32015 6780 32025 6815
rect 32060 6780 32070 6815
rect 32105 6780 32115 6815
rect 32150 6780 32160 6815
rect 32195 6780 32205 6815
rect 32240 6780 32250 6815
rect 32285 6780 32295 6815
rect 32330 6780 32340 6815
rect 32375 6780 32385 6815
rect 32420 6780 32430 6815
rect 32465 6780 32475 6815
rect 32510 6780 32520 6815
rect 32555 6780 32565 6815
rect 32600 6780 32610 6815
rect 32645 6780 32655 6815
rect 32690 6780 32700 6815
rect 32735 6780 32745 6815
rect 32780 6780 32790 6815
rect 32825 6780 32835 6815
rect 32870 6780 35620 6815
rect 31290 6770 35620 6780
rect 31290 6735 31305 6770
rect 31340 6735 31350 6770
rect 31385 6735 31395 6770
rect 31430 6735 31440 6770
rect 31475 6735 31485 6770
rect 31520 6735 31530 6770
rect 31565 6735 31575 6770
rect 31610 6735 31620 6770
rect 31655 6735 31665 6770
rect 31700 6735 31710 6770
rect 31745 6735 31755 6770
rect 31790 6735 31800 6770
rect 31835 6735 31845 6770
rect 31880 6735 31890 6770
rect 31925 6735 31935 6770
rect 31970 6735 31980 6770
rect 32015 6735 32025 6770
rect 32060 6735 32070 6770
rect 32105 6735 32115 6770
rect 32150 6735 32160 6770
rect 32195 6735 32205 6770
rect 32240 6735 32250 6770
rect 32285 6735 32295 6770
rect 32330 6735 32340 6770
rect 32375 6735 32385 6770
rect 32420 6735 32430 6770
rect 32465 6735 32475 6770
rect 32510 6735 32520 6770
rect 32555 6735 32565 6770
rect 32600 6735 32610 6770
rect 32645 6735 32655 6770
rect 32690 6735 32700 6770
rect 32735 6735 32745 6770
rect 32780 6735 32790 6770
rect 32825 6735 32835 6770
rect 32870 6735 35620 6770
rect 31290 6725 35620 6735
rect 31290 6690 31305 6725
rect 31340 6690 31350 6725
rect 31385 6690 31395 6725
rect 31430 6690 31440 6725
rect 31475 6690 31485 6725
rect 31520 6690 31530 6725
rect 31565 6690 31575 6725
rect 31610 6690 31620 6725
rect 31655 6690 31665 6725
rect 31700 6690 31710 6725
rect 31745 6690 31755 6725
rect 31790 6690 31800 6725
rect 31835 6690 31845 6725
rect 31880 6690 31890 6725
rect 31925 6690 31935 6725
rect 31970 6690 31980 6725
rect 32015 6690 32025 6725
rect 32060 6690 32070 6725
rect 32105 6690 32115 6725
rect 32150 6690 32160 6725
rect 32195 6690 32205 6725
rect 32240 6690 32250 6725
rect 32285 6690 32295 6725
rect 32330 6690 32340 6725
rect 32375 6690 32385 6725
rect 32420 6690 32430 6725
rect 32465 6690 32475 6725
rect 32510 6690 32520 6725
rect 32555 6690 32565 6725
rect 32600 6690 32610 6725
rect 32645 6690 32655 6725
rect 32690 6690 32700 6725
rect 32735 6690 32745 6725
rect 32780 6690 32790 6725
rect 32825 6690 32835 6725
rect 32870 6690 35620 6725
rect 31290 6680 35620 6690
rect 31290 6645 31305 6680
rect 31340 6645 31350 6680
rect 31385 6645 31395 6680
rect 31430 6645 31440 6680
rect 31475 6645 31485 6680
rect 31520 6645 31530 6680
rect 31565 6645 31575 6680
rect 31610 6645 31620 6680
rect 31655 6645 31665 6680
rect 31700 6645 31710 6680
rect 31745 6645 31755 6680
rect 31790 6645 31800 6680
rect 31835 6645 31845 6680
rect 31880 6645 31890 6680
rect 31925 6645 31935 6680
rect 31970 6645 31980 6680
rect 32015 6645 32025 6680
rect 32060 6645 32070 6680
rect 32105 6645 32115 6680
rect 32150 6645 32160 6680
rect 32195 6645 32205 6680
rect 32240 6645 32250 6680
rect 32285 6645 32295 6680
rect 32330 6645 32340 6680
rect 32375 6645 32385 6680
rect 32420 6645 32430 6680
rect 32465 6645 32475 6680
rect 32510 6645 32520 6680
rect 32555 6645 32565 6680
rect 32600 6645 32610 6680
rect 32645 6645 32655 6680
rect 32690 6645 32700 6680
rect 32735 6645 32745 6680
rect 32780 6645 32790 6680
rect 32825 6645 32835 6680
rect 32870 6645 35620 6680
rect 31290 6635 35620 6645
rect 31290 6600 31305 6635
rect 31340 6600 31350 6635
rect 31385 6600 31395 6635
rect 31430 6600 31440 6635
rect 31475 6600 31485 6635
rect 31520 6600 31530 6635
rect 31565 6600 31575 6635
rect 31610 6600 31620 6635
rect 31655 6600 31665 6635
rect 31700 6600 31710 6635
rect 31745 6600 31755 6635
rect 31790 6600 31800 6635
rect 31835 6600 31845 6635
rect 31880 6600 31890 6635
rect 31925 6600 31935 6635
rect 31970 6600 31980 6635
rect 32015 6600 32025 6635
rect 32060 6600 32070 6635
rect 32105 6600 32115 6635
rect 32150 6600 32160 6635
rect 32195 6600 32205 6635
rect 32240 6600 32250 6635
rect 32285 6600 32295 6635
rect 32330 6600 32340 6635
rect 32375 6600 32385 6635
rect 32420 6600 32430 6635
rect 32465 6600 32475 6635
rect 32510 6600 32520 6635
rect 32555 6600 32565 6635
rect 32600 6600 32610 6635
rect 32645 6600 32655 6635
rect 32690 6600 32700 6635
rect 32735 6600 32745 6635
rect 32780 6600 32790 6635
rect 32825 6600 32835 6635
rect 32870 6600 35620 6635
rect 31290 6590 35620 6600
rect 31290 6555 31305 6590
rect 31340 6555 31350 6590
rect 31385 6555 31395 6590
rect 31430 6555 31440 6590
rect 31475 6555 31485 6590
rect 31520 6555 31530 6590
rect 31565 6555 31575 6590
rect 31610 6555 31620 6590
rect 31655 6555 31665 6590
rect 31700 6555 31710 6590
rect 31745 6555 31755 6590
rect 31790 6555 31800 6590
rect 31835 6555 31845 6590
rect 31880 6555 31890 6590
rect 31925 6555 31935 6590
rect 31970 6555 31980 6590
rect 32015 6555 32025 6590
rect 32060 6555 32070 6590
rect 32105 6555 32115 6590
rect 32150 6555 32160 6590
rect 32195 6555 32205 6590
rect 32240 6555 32250 6590
rect 32285 6555 32295 6590
rect 32330 6555 32340 6590
rect 32375 6555 32385 6590
rect 32420 6555 32430 6590
rect 32465 6555 32475 6590
rect 32510 6555 32520 6590
rect 32555 6555 32565 6590
rect 32600 6555 32610 6590
rect 32645 6555 32655 6590
rect 32690 6555 32700 6590
rect 32735 6555 32745 6590
rect 32780 6555 32790 6590
rect 32825 6555 32835 6590
rect 32870 6555 35620 6590
rect 31290 6545 35620 6555
rect 31290 6510 31305 6545
rect 31340 6510 31350 6545
rect 31385 6510 31395 6545
rect 31430 6510 31440 6545
rect 31475 6510 31485 6545
rect 31520 6510 31530 6545
rect 31565 6510 31575 6545
rect 31610 6510 31620 6545
rect 31655 6510 31665 6545
rect 31700 6510 31710 6545
rect 31745 6510 31755 6545
rect 31790 6510 31800 6545
rect 31835 6510 31845 6545
rect 31880 6510 31890 6545
rect 31925 6510 31935 6545
rect 31970 6510 31980 6545
rect 32015 6510 32025 6545
rect 32060 6510 32070 6545
rect 32105 6510 32115 6545
rect 32150 6510 32160 6545
rect 32195 6510 32205 6545
rect 32240 6510 32250 6545
rect 32285 6510 32295 6545
rect 32330 6510 32340 6545
rect 32375 6510 32385 6545
rect 32420 6510 32430 6545
rect 32465 6510 32475 6545
rect 32510 6510 32520 6545
rect 32555 6510 32565 6545
rect 32600 6510 32610 6545
rect 32645 6510 32655 6545
rect 32690 6510 32700 6545
rect 32735 6510 32745 6545
rect 32780 6510 32790 6545
rect 32825 6510 32835 6545
rect 32870 6510 35620 6545
rect 31290 6500 35620 6510
rect 31290 6465 31305 6500
rect 31340 6465 31350 6500
rect 31385 6465 31395 6500
rect 31430 6465 31440 6500
rect 31475 6465 31485 6500
rect 31520 6465 31530 6500
rect 31565 6465 31575 6500
rect 31610 6465 31620 6500
rect 31655 6465 31665 6500
rect 31700 6465 31710 6500
rect 31745 6465 31755 6500
rect 31790 6465 31800 6500
rect 31835 6465 31845 6500
rect 31880 6465 31890 6500
rect 31925 6465 31935 6500
rect 31970 6465 31980 6500
rect 32015 6465 32025 6500
rect 32060 6465 32070 6500
rect 32105 6465 32115 6500
rect 32150 6465 32160 6500
rect 32195 6465 32205 6500
rect 32240 6465 32250 6500
rect 32285 6465 32295 6500
rect 32330 6465 32340 6500
rect 32375 6465 32385 6500
rect 32420 6465 32430 6500
rect 32465 6465 32475 6500
rect 32510 6465 32520 6500
rect 32555 6465 32565 6500
rect 32600 6465 32610 6500
rect 32645 6465 32655 6500
rect 32690 6465 32700 6500
rect 32735 6465 32745 6500
rect 32780 6465 32790 6500
rect 32825 6465 32835 6500
rect 32870 6465 35620 6500
rect 31290 6450 35620 6465
rect -120 -1300 32890 -1290
rect -120 -1340 -80 -1300
rect -40 -1340 270 -1300
rect 310 -1340 620 -1300
rect 660 -1340 970 -1300
rect 1010 -1340 1320 -1300
rect 1360 -1340 1670 -1300
rect 1710 -1340 2020 -1300
rect 2060 -1340 2370 -1300
rect 2410 -1340 2720 -1300
rect 2760 -1340 3070 -1300
rect 3110 -1340 3420 -1300
rect 3460 -1340 3770 -1300
rect 3810 -1340 4120 -1300
rect 4160 -1340 4470 -1300
rect 4510 -1340 4820 -1300
rect 4860 -1340 5170 -1300
rect 5210 -1340 5520 -1300
rect 5560 -1340 5870 -1300
rect 5910 -1340 6220 -1300
rect 6260 -1340 6570 -1300
rect 6610 -1340 6920 -1300
rect 6960 -1340 7270 -1300
rect 7310 -1340 7620 -1300
rect 7660 -1340 7970 -1300
rect 8010 -1340 8320 -1300
rect 8360 -1310 32890 -1300
rect 8360 -1340 31305 -1310
rect -120 -1345 31305 -1340
rect 31340 -1345 31350 -1310
rect 31385 -1345 31395 -1310
rect 31430 -1345 31440 -1310
rect 31475 -1345 31485 -1310
rect 31520 -1345 31530 -1310
rect 31565 -1345 31575 -1310
rect 31610 -1345 31620 -1310
rect 31655 -1345 31665 -1310
rect 31700 -1345 31710 -1310
rect 31745 -1345 31755 -1310
rect 31790 -1345 31800 -1310
rect 31835 -1345 31845 -1310
rect 31880 -1345 31890 -1310
rect 31925 -1345 31935 -1310
rect 31970 -1345 31980 -1310
rect 32015 -1345 32025 -1310
rect 32060 -1345 32070 -1310
rect 32105 -1345 32115 -1310
rect 32150 -1345 32160 -1310
rect 32195 -1345 32205 -1310
rect 32240 -1345 32250 -1310
rect 32285 -1345 32295 -1310
rect 32330 -1345 32340 -1310
rect 32375 -1345 32385 -1310
rect 32420 -1345 32430 -1310
rect 32465 -1345 32475 -1310
rect 32510 -1345 32520 -1310
rect 32555 -1345 32565 -1310
rect 32600 -1345 32610 -1310
rect 32645 -1345 32655 -1310
rect 32690 -1345 32700 -1310
rect 32735 -1345 32745 -1310
rect 32780 -1345 32790 -1310
rect 32825 -1345 32835 -1310
rect 32870 -1345 32890 -1310
rect -120 -1355 32890 -1345
rect -120 -1365 31305 -1355
rect -120 -1405 -80 -1365
rect -40 -1405 270 -1365
rect 310 -1405 620 -1365
rect 660 -1405 970 -1365
rect 1010 -1405 1320 -1365
rect 1360 -1405 1670 -1365
rect 1710 -1405 2020 -1365
rect 2060 -1405 2370 -1365
rect 2410 -1405 2720 -1365
rect 2760 -1405 3070 -1365
rect 3110 -1405 3420 -1365
rect 3460 -1405 3770 -1365
rect 3810 -1405 4120 -1365
rect 4160 -1405 4470 -1365
rect 4510 -1405 4820 -1365
rect 4860 -1405 5170 -1365
rect 5210 -1405 5520 -1365
rect 5560 -1405 5870 -1365
rect 5910 -1405 6220 -1365
rect 6260 -1405 6570 -1365
rect 6610 -1405 6920 -1365
rect 6960 -1405 7270 -1365
rect 7310 -1405 7620 -1365
rect 7660 -1405 7970 -1365
rect 8010 -1405 8320 -1365
rect 8360 -1390 31305 -1365
rect 31340 -1390 31350 -1355
rect 31385 -1390 31395 -1355
rect 31430 -1390 31440 -1355
rect 31475 -1390 31485 -1355
rect 31520 -1390 31530 -1355
rect 31565 -1390 31575 -1355
rect 31610 -1390 31620 -1355
rect 31655 -1390 31665 -1355
rect 31700 -1390 31710 -1355
rect 31745 -1390 31755 -1355
rect 31790 -1390 31800 -1355
rect 31835 -1390 31845 -1355
rect 31880 -1390 31890 -1355
rect 31925 -1390 31935 -1355
rect 31970 -1390 31980 -1355
rect 32015 -1390 32025 -1355
rect 32060 -1390 32070 -1355
rect 32105 -1390 32115 -1355
rect 32150 -1390 32160 -1355
rect 32195 -1390 32205 -1355
rect 32240 -1390 32250 -1355
rect 32285 -1390 32295 -1355
rect 32330 -1390 32340 -1355
rect 32375 -1390 32385 -1355
rect 32420 -1390 32430 -1355
rect 32465 -1390 32475 -1355
rect 32510 -1390 32520 -1355
rect 32555 -1390 32565 -1355
rect 32600 -1390 32610 -1355
rect 32645 -1390 32655 -1355
rect 32690 -1390 32700 -1355
rect 32735 -1390 32745 -1355
rect 32780 -1390 32790 -1355
rect 32825 -1390 32835 -1355
rect 32870 -1390 32890 -1355
rect 8360 -1400 32890 -1390
rect 8360 -1405 31305 -1400
rect -120 -1435 31305 -1405
rect 31340 -1435 31350 -1400
rect 31385 -1435 31395 -1400
rect 31430 -1435 31440 -1400
rect 31475 -1435 31485 -1400
rect 31520 -1435 31530 -1400
rect 31565 -1435 31575 -1400
rect 31610 -1435 31620 -1400
rect 31655 -1435 31665 -1400
rect 31700 -1435 31710 -1400
rect 31745 -1435 31755 -1400
rect 31790 -1435 31800 -1400
rect 31835 -1435 31845 -1400
rect 31880 -1435 31890 -1400
rect 31925 -1435 31935 -1400
rect 31970 -1435 31980 -1400
rect 32015 -1435 32025 -1400
rect 32060 -1435 32070 -1400
rect 32105 -1435 32115 -1400
rect 32150 -1435 32160 -1400
rect 32195 -1435 32205 -1400
rect 32240 -1435 32250 -1400
rect 32285 -1435 32295 -1400
rect 32330 -1435 32340 -1400
rect 32375 -1435 32385 -1400
rect 32420 -1435 32430 -1400
rect 32465 -1435 32475 -1400
rect 32510 -1435 32520 -1400
rect 32555 -1435 32565 -1400
rect 32600 -1435 32610 -1400
rect 32645 -1435 32655 -1400
rect 32690 -1435 32700 -1400
rect 32735 -1435 32745 -1400
rect 32780 -1435 32790 -1400
rect 32825 -1435 32835 -1400
rect 32870 -1435 32890 -1400
rect -120 -1475 -80 -1435
rect -40 -1475 270 -1435
rect 310 -1475 620 -1435
rect 660 -1475 970 -1435
rect 1010 -1475 1320 -1435
rect 1360 -1475 1670 -1435
rect 1710 -1475 2020 -1435
rect 2060 -1475 2370 -1435
rect 2410 -1475 2720 -1435
rect 2760 -1475 3070 -1435
rect 3110 -1475 3420 -1435
rect 3460 -1475 3770 -1435
rect 3810 -1475 4120 -1435
rect 4160 -1475 4470 -1435
rect 4510 -1475 4820 -1435
rect 4860 -1475 5170 -1435
rect 5210 -1475 5520 -1435
rect 5560 -1475 5870 -1435
rect 5910 -1475 6220 -1435
rect 6260 -1475 6570 -1435
rect 6610 -1475 6920 -1435
rect 6960 -1475 7270 -1435
rect 7310 -1475 7620 -1435
rect 7660 -1475 7970 -1435
rect 8010 -1475 8320 -1435
rect 8360 -1445 32890 -1435
rect 8360 -1475 31305 -1445
rect -120 -1480 31305 -1475
rect 31340 -1480 31350 -1445
rect 31385 -1480 31395 -1445
rect 31430 -1480 31440 -1445
rect 31475 -1480 31485 -1445
rect 31520 -1480 31530 -1445
rect 31565 -1480 31575 -1445
rect 31610 -1480 31620 -1445
rect 31655 -1480 31665 -1445
rect 31700 -1480 31710 -1445
rect 31745 -1480 31755 -1445
rect 31790 -1480 31800 -1445
rect 31835 -1480 31845 -1445
rect 31880 -1480 31890 -1445
rect 31925 -1480 31935 -1445
rect 31970 -1480 31980 -1445
rect 32015 -1480 32025 -1445
rect 32060 -1480 32070 -1445
rect 32105 -1480 32115 -1445
rect 32150 -1480 32160 -1445
rect 32195 -1480 32205 -1445
rect 32240 -1480 32250 -1445
rect 32285 -1480 32295 -1445
rect 32330 -1480 32340 -1445
rect 32375 -1480 32385 -1445
rect 32420 -1480 32430 -1445
rect 32465 -1480 32475 -1445
rect 32510 -1480 32520 -1445
rect 32555 -1480 32565 -1445
rect 32600 -1480 32610 -1445
rect 32645 -1480 32655 -1445
rect 32690 -1480 32700 -1445
rect 32735 -1480 32745 -1445
rect 32780 -1480 32790 -1445
rect 32825 -1480 32835 -1445
rect 32870 -1480 32890 -1445
rect -120 -1490 32890 -1480
rect -120 -1505 31305 -1490
rect -120 -1545 -80 -1505
rect -40 -1545 270 -1505
rect 310 -1545 620 -1505
rect 660 -1545 970 -1505
rect 1010 -1545 1320 -1505
rect 1360 -1545 1670 -1505
rect 1710 -1545 2020 -1505
rect 2060 -1545 2370 -1505
rect 2410 -1545 2720 -1505
rect 2760 -1545 3070 -1505
rect 3110 -1545 3420 -1505
rect 3460 -1545 3770 -1505
rect 3810 -1545 4120 -1505
rect 4160 -1545 4470 -1505
rect 4510 -1545 4820 -1505
rect 4860 -1545 5170 -1505
rect 5210 -1545 5520 -1505
rect 5560 -1545 5870 -1505
rect 5910 -1545 6220 -1505
rect 6260 -1545 6570 -1505
rect 6610 -1545 6920 -1505
rect 6960 -1545 7270 -1505
rect 7310 -1545 7620 -1505
rect 7660 -1545 7970 -1505
rect 8010 -1545 8320 -1505
rect 8360 -1525 31305 -1505
rect 31340 -1525 31350 -1490
rect 31385 -1525 31395 -1490
rect 31430 -1525 31440 -1490
rect 31475 -1525 31485 -1490
rect 31520 -1525 31530 -1490
rect 31565 -1525 31575 -1490
rect 31610 -1525 31620 -1490
rect 31655 -1525 31665 -1490
rect 31700 -1525 31710 -1490
rect 31745 -1525 31755 -1490
rect 31790 -1525 31800 -1490
rect 31835 -1525 31845 -1490
rect 31880 -1525 31890 -1490
rect 31925 -1525 31935 -1490
rect 31970 -1525 31980 -1490
rect 32015 -1525 32025 -1490
rect 32060 -1525 32070 -1490
rect 32105 -1525 32115 -1490
rect 32150 -1525 32160 -1490
rect 32195 -1525 32205 -1490
rect 32240 -1525 32250 -1490
rect 32285 -1525 32295 -1490
rect 32330 -1525 32340 -1490
rect 32375 -1525 32385 -1490
rect 32420 -1525 32430 -1490
rect 32465 -1525 32475 -1490
rect 32510 -1525 32520 -1490
rect 32555 -1525 32565 -1490
rect 32600 -1525 32610 -1490
rect 32645 -1525 32655 -1490
rect 32690 -1525 32700 -1490
rect 32735 -1525 32745 -1490
rect 32780 -1525 32790 -1490
rect 32825 -1525 32835 -1490
rect 32870 -1525 32890 -1490
rect 8360 -1535 32890 -1525
rect 8360 -1545 31305 -1535
rect -120 -1570 31305 -1545
rect 31340 -1570 31350 -1535
rect 31385 -1570 31395 -1535
rect 31430 -1570 31440 -1535
rect 31475 -1570 31485 -1535
rect 31520 -1570 31530 -1535
rect 31565 -1570 31575 -1535
rect 31610 -1570 31620 -1535
rect 31655 -1570 31665 -1535
rect 31700 -1570 31710 -1535
rect 31745 -1570 31755 -1535
rect 31790 -1570 31800 -1535
rect 31835 -1570 31845 -1535
rect 31880 -1570 31890 -1535
rect 31925 -1570 31935 -1535
rect 31970 -1570 31980 -1535
rect 32015 -1570 32025 -1535
rect 32060 -1570 32070 -1535
rect 32105 -1570 32115 -1535
rect 32150 -1570 32160 -1535
rect 32195 -1570 32205 -1535
rect 32240 -1570 32250 -1535
rect 32285 -1570 32295 -1535
rect 32330 -1570 32340 -1535
rect 32375 -1570 32385 -1535
rect 32420 -1570 32430 -1535
rect 32465 -1570 32475 -1535
rect 32510 -1570 32520 -1535
rect 32555 -1570 32565 -1535
rect 32600 -1570 32610 -1535
rect 32645 -1570 32655 -1535
rect 32690 -1570 32700 -1535
rect 32735 -1570 32745 -1535
rect 32780 -1570 32790 -1535
rect 32825 -1570 32835 -1535
rect 32870 -1570 32890 -1535
rect -120 -1575 32890 -1570
rect -120 -1615 -80 -1575
rect -40 -1615 270 -1575
rect 310 -1615 620 -1575
rect 660 -1615 970 -1575
rect 1010 -1615 1320 -1575
rect 1360 -1615 1670 -1575
rect 1710 -1615 2020 -1575
rect 2060 -1615 2370 -1575
rect 2410 -1615 2720 -1575
rect 2760 -1615 3070 -1575
rect 3110 -1615 3420 -1575
rect 3460 -1615 3770 -1575
rect 3810 -1615 4120 -1575
rect 4160 -1615 4470 -1575
rect 4510 -1615 4820 -1575
rect 4860 -1615 5170 -1575
rect 5210 -1615 5520 -1575
rect 5560 -1615 5870 -1575
rect 5910 -1615 6220 -1575
rect 6260 -1615 6570 -1575
rect 6610 -1615 6920 -1575
rect 6960 -1615 7270 -1575
rect 7310 -1615 7620 -1575
rect 7660 -1615 7970 -1575
rect 8010 -1615 8320 -1575
rect 8360 -1580 32890 -1575
rect 8360 -1615 31305 -1580
rect 31340 -1615 31350 -1580
rect 31385 -1615 31395 -1580
rect 31430 -1615 31440 -1580
rect 31475 -1615 31485 -1580
rect 31520 -1615 31530 -1580
rect 31565 -1615 31575 -1580
rect 31610 -1615 31620 -1580
rect 31655 -1615 31665 -1580
rect 31700 -1615 31710 -1580
rect 31745 -1615 31755 -1580
rect 31790 -1615 31800 -1580
rect 31835 -1615 31845 -1580
rect 31880 -1615 31890 -1580
rect 31925 -1615 31935 -1580
rect 31970 -1615 31980 -1580
rect 32015 -1615 32025 -1580
rect 32060 -1615 32070 -1580
rect 32105 -1615 32115 -1580
rect 32150 -1615 32160 -1580
rect 32195 -1615 32205 -1580
rect 32240 -1615 32250 -1580
rect 32285 -1615 32295 -1580
rect 32330 -1615 32340 -1580
rect 32375 -1615 32385 -1580
rect 32420 -1615 32430 -1580
rect 32465 -1615 32475 -1580
rect 32510 -1615 32520 -1580
rect 32555 -1615 32565 -1580
rect 32600 -1615 32610 -1580
rect 32645 -1615 32655 -1580
rect 32690 -1615 32700 -1580
rect 32735 -1615 32745 -1580
rect 32780 -1615 32790 -1580
rect 32825 -1615 32835 -1580
rect 32870 -1615 32890 -1580
rect -120 -1625 32890 -1615
rect -120 -1640 31305 -1625
rect -120 -1680 -80 -1640
rect -40 -1680 270 -1640
rect 310 -1680 620 -1640
rect 660 -1680 970 -1640
rect 1010 -1680 1320 -1640
rect 1360 -1680 1670 -1640
rect 1710 -1680 2020 -1640
rect 2060 -1680 2370 -1640
rect 2410 -1680 2720 -1640
rect 2760 -1680 3070 -1640
rect 3110 -1680 3420 -1640
rect 3460 -1680 3770 -1640
rect 3810 -1680 4120 -1640
rect 4160 -1680 4470 -1640
rect 4510 -1680 4820 -1640
rect 4860 -1680 5170 -1640
rect 5210 -1680 5520 -1640
rect 5560 -1680 5870 -1640
rect 5910 -1680 6220 -1640
rect 6260 -1680 6570 -1640
rect 6610 -1680 6920 -1640
rect 6960 -1680 7270 -1640
rect 7310 -1680 7620 -1640
rect 7660 -1680 7970 -1640
rect 8010 -1680 8320 -1640
rect 8360 -1660 31305 -1640
rect 31340 -1660 31350 -1625
rect 31385 -1660 31395 -1625
rect 31430 -1660 31440 -1625
rect 31475 -1660 31485 -1625
rect 31520 -1660 31530 -1625
rect 31565 -1660 31575 -1625
rect 31610 -1660 31620 -1625
rect 31655 -1660 31665 -1625
rect 31700 -1660 31710 -1625
rect 31745 -1660 31755 -1625
rect 31790 -1660 31800 -1625
rect 31835 -1660 31845 -1625
rect 31880 -1660 31890 -1625
rect 31925 -1660 31935 -1625
rect 31970 -1660 31980 -1625
rect 32015 -1660 32025 -1625
rect 32060 -1660 32070 -1625
rect 32105 -1660 32115 -1625
rect 32150 -1660 32160 -1625
rect 32195 -1660 32205 -1625
rect 32240 -1660 32250 -1625
rect 32285 -1660 32295 -1625
rect 32330 -1660 32340 -1625
rect 32375 -1660 32385 -1625
rect 32420 -1660 32430 -1625
rect 32465 -1660 32475 -1625
rect 32510 -1660 32520 -1625
rect 32555 -1660 32565 -1625
rect 32600 -1660 32610 -1625
rect 32645 -1660 32655 -1625
rect 32690 -1660 32700 -1625
rect 32735 -1660 32745 -1625
rect 32780 -1660 32790 -1625
rect 32825 -1660 32835 -1625
rect 32870 -1660 32890 -1625
rect 8360 -1670 32890 -1660
rect 8360 -1680 31305 -1670
rect -120 -1700 31305 -1680
rect -120 -1740 -80 -1700
rect -40 -1740 270 -1700
rect 310 -1740 620 -1700
rect 660 -1740 970 -1700
rect 1010 -1740 1320 -1700
rect 1360 -1740 1670 -1700
rect 1710 -1740 2020 -1700
rect 2060 -1740 2370 -1700
rect 2410 -1740 2720 -1700
rect 2760 -1740 3070 -1700
rect 3110 -1740 3420 -1700
rect 3460 -1740 3770 -1700
rect 3810 -1740 4120 -1700
rect 4160 -1740 4470 -1700
rect 4510 -1740 4820 -1700
rect 4860 -1740 5170 -1700
rect 5210 -1740 5520 -1700
rect 5560 -1740 5870 -1700
rect 5910 -1740 6220 -1700
rect 6260 -1740 6570 -1700
rect 6610 -1740 6920 -1700
rect 6960 -1740 7270 -1700
rect 7310 -1740 7620 -1700
rect 7660 -1740 7970 -1700
rect 8010 -1740 8320 -1700
rect 8360 -1705 31305 -1700
rect 31340 -1705 31350 -1670
rect 31385 -1705 31395 -1670
rect 31430 -1705 31440 -1670
rect 31475 -1705 31485 -1670
rect 31520 -1705 31530 -1670
rect 31565 -1705 31575 -1670
rect 31610 -1705 31620 -1670
rect 31655 -1705 31665 -1670
rect 31700 -1705 31710 -1670
rect 31745 -1705 31755 -1670
rect 31790 -1705 31800 -1670
rect 31835 -1705 31845 -1670
rect 31880 -1705 31890 -1670
rect 31925 -1705 31935 -1670
rect 31970 -1705 31980 -1670
rect 32015 -1705 32025 -1670
rect 32060 -1705 32070 -1670
rect 32105 -1705 32115 -1670
rect 32150 -1705 32160 -1670
rect 32195 -1705 32205 -1670
rect 32240 -1705 32250 -1670
rect 32285 -1705 32295 -1670
rect 32330 -1705 32340 -1670
rect 32375 -1705 32385 -1670
rect 32420 -1705 32430 -1670
rect 32465 -1705 32475 -1670
rect 32510 -1705 32520 -1670
rect 32555 -1705 32565 -1670
rect 32600 -1705 32610 -1670
rect 32645 -1705 32655 -1670
rect 32690 -1705 32700 -1670
rect 32735 -1705 32745 -1670
rect 32780 -1705 32790 -1670
rect 32825 -1705 32835 -1670
rect 32870 -1705 32890 -1670
rect 8360 -1715 32890 -1705
rect 8360 -1740 31305 -1715
rect -120 -1750 31305 -1740
rect 31340 -1750 31350 -1715
rect 31385 -1750 31395 -1715
rect 31430 -1750 31440 -1715
rect 31475 -1750 31485 -1715
rect 31520 -1750 31530 -1715
rect 31565 -1750 31575 -1715
rect 31610 -1750 31620 -1715
rect 31655 -1750 31665 -1715
rect 31700 -1750 31710 -1715
rect 31745 -1750 31755 -1715
rect 31790 -1750 31800 -1715
rect 31835 -1750 31845 -1715
rect 31880 -1750 31890 -1715
rect 31925 -1750 31935 -1715
rect 31970 -1750 31980 -1715
rect 32015 -1750 32025 -1715
rect 32060 -1750 32070 -1715
rect 32105 -1750 32115 -1715
rect 32150 -1750 32160 -1715
rect 32195 -1750 32205 -1715
rect 32240 -1750 32250 -1715
rect 32285 -1750 32295 -1715
rect 32330 -1750 32340 -1715
rect 32375 -1750 32385 -1715
rect 32420 -1750 32430 -1715
rect 32465 -1750 32475 -1715
rect 32510 -1750 32520 -1715
rect 32555 -1750 32565 -1715
rect 32600 -1750 32610 -1715
rect 32645 -1750 32655 -1715
rect 32690 -1750 32700 -1715
rect 32735 -1750 32745 -1715
rect 32780 -1750 32790 -1715
rect 32825 -1750 32835 -1715
rect 32870 -1750 32890 -1715
rect -120 -1760 32890 -1750
rect -120 -1765 31305 -1760
rect -120 -1805 -80 -1765
rect -40 -1805 270 -1765
rect 310 -1805 620 -1765
rect 660 -1805 970 -1765
rect 1010 -1805 1320 -1765
rect 1360 -1805 1670 -1765
rect 1710 -1805 2020 -1765
rect 2060 -1805 2370 -1765
rect 2410 -1805 2720 -1765
rect 2760 -1805 3070 -1765
rect 3110 -1805 3420 -1765
rect 3460 -1805 3770 -1765
rect 3810 -1805 4120 -1765
rect 4160 -1805 4470 -1765
rect 4510 -1805 4820 -1765
rect 4860 -1805 5170 -1765
rect 5210 -1805 5520 -1765
rect 5560 -1805 5870 -1765
rect 5910 -1805 6220 -1765
rect 6260 -1805 6570 -1765
rect 6610 -1805 6920 -1765
rect 6960 -1805 7270 -1765
rect 7310 -1805 7620 -1765
rect 7660 -1805 7970 -1765
rect 8010 -1805 8320 -1765
rect 8360 -1795 31305 -1765
rect 31340 -1795 31350 -1760
rect 31385 -1795 31395 -1760
rect 31430 -1795 31440 -1760
rect 31475 -1795 31485 -1760
rect 31520 -1795 31530 -1760
rect 31565 -1795 31575 -1760
rect 31610 -1795 31620 -1760
rect 31655 -1795 31665 -1760
rect 31700 -1795 31710 -1760
rect 31745 -1795 31755 -1760
rect 31790 -1795 31800 -1760
rect 31835 -1795 31845 -1760
rect 31880 -1795 31890 -1760
rect 31925 -1795 31935 -1760
rect 31970 -1795 31980 -1760
rect 32015 -1795 32025 -1760
rect 32060 -1795 32070 -1760
rect 32105 -1795 32115 -1760
rect 32150 -1795 32160 -1760
rect 32195 -1795 32205 -1760
rect 32240 -1795 32250 -1760
rect 32285 -1795 32295 -1760
rect 32330 -1795 32340 -1760
rect 32375 -1795 32385 -1760
rect 32420 -1795 32430 -1760
rect 32465 -1795 32475 -1760
rect 32510 -1795 32520 -1760
rect 32555 -1795 32565 -1760
rect 32600 -1795 32610 -1760
rect 32645 -1795 32655 -1760
rect 32690 -1795 32700 -1760
rect 32735 -1795 32745 -1760
rect 32780 -1795 32790 -1760
rect 32825 -1795 32835 -1760
rect 32870 -1795 32890 -1760
rect 8360 -1805 32890 -1795
rect -120 -1835 31305 -1805
rect -120 -1875 -80 -1835
rect -40 -1875 270 -1835
rect 310 -1875 620 -1835
rect 660 -1875 970 -1835
rect 1010 -1875 1320 -1835
rect 1360 -1875 1670 -1835
rect 1710 -1875 2020 -1835
rect 2060 -1875 2370 -1835
rect 2410 -1875 2720 -1835
rect 2760 -1875 3070 -1835
rect 3110 -1875 3420 -1835
rect 3460 -1875 3770 -1835
rect 3810 -1875 4120 -1835
rect 4160 -1875 4470 -1835
rect 4510 -1875 4820 -1835
rect 4860 -1875 5170 -1835
rect 5210 -1875 5520 -1835
rect 5560 -1875 5870 -1835
rect 5910 -1875 6220 -1835
rect 6260 -1875 6570 -1835
rect 6610 -1875 6920 -1835
rect 6960 -1875 7270 -1835
rect 7310 -1875 7620 -1835
rect 7660 -1875 7970 -1835
rect 8010 -1875 8320 -1835
rect 8360 -1840 31305 -1835
rect 31340 -1840 31350 -1805
rect 31385 -1840 31395 -1805
rect 31430 -1840 31440 -1805
rect 31475 -1840 31485 -1805
rect 31520 -1840 31530 -1805
rect 31565 -1840 31575 -1805
rect 31610 -1840 31620 -1805
rect 31655 -1840 31665 -1805
rect 31700 -1840 31710 -1805
rect 31745 -1840 31755 -1805
rect 31790 -1840 31800 -1805
rect 31835 -1840 31845 -1805
rect 31880 -1840 31890 -1805
rect 31925 -1840 31935 -1805
rect 31970 -1840 31980 -1805
rect 32015 -1840 32025 -1805
rect 32060 -1840 32070 -1805
rect 32105 -1840 32115 -1805
rect 32150 -1840 32160 -1805
rect 32195 -1840 32205 -1805
rect 32240 -1840 32250 -1805
rect 32285 -1840 32295 -1805
rect 32330 -1840 32340 -1805
rect 32375 -1840 32385 -1805
rect 32420 -1840 32430 -1805
rect 32465 -1840 32475 -1805
rect 32510 -1840 32520 -1805
rect 32555 -1840 32565 -1805
rect 32600 -1840 32610 -1805
rect 32645 -1840 32655 -1805
rect 32690 -1840 32700 -1805
rect 32735 -1840 32745 -1805
rect 32780 -1840 32790 -1805
rect 32825 -1840 32835 -1805
rect 32870 -1840 32890 -1805
rect 8360 -1850 32890 -1840
rect 8360 -1875 31305 -1850
rect -120 -1885 31305 -1875
rect 31340 -1885 31350 -1850
rect 31385 -1885 31395 -1850
rect 31430 -1885 31440 -1850
rect 31475 -1885 31485 -1850
rect 31520 -1885 31530 -1850
rect 31565 -1885 31575 -1850
rect 31610 -1885 31620 -1850
rect 31655 -1885 31665 -1850
rect 31700 -1885 31710 -1850
rect 31745 -1885 31755 -1850
rect 31790 -1885 31800 -1850
rect 31835 -1885 31845 -1850
rect 31880 -1885 31890 -1850
rect 31925 -1885 31935 -1850
rect 31970 -1885 31980 -1850
rect 32015 -1885 32025 -1850
rect 32060 -1885 32070 -1850
rect 32105 -1885 32115 -1850
rect 32150 -1885 32160 -1850
rect 32195 -1885 32205 -1850
rect 32240 -1885 32250 -1850
rect 32285 -1885 32295 -1850
rect 32330 -1885 32340 -1850
rect 32375 -1885 32385 -1850
rect 32420 -1885 32430 -1850
rect 32465 -1885 32475 -1850
rect 32510 -1885 32520 -1850
rect 32555 -1885 32565 -1850
rect 32600 -1885 32610 -1850
rect 32645 -1885 32655 -1850
rect 32690 -1885 32700 -1850
rect 32735 -1885 32745 -1850
rect 32780 -1885 32790 -1850
rect 32825 -1885 32835 -1850
rect 32870 -1885 32890 -1850
rect -120 -1895 32890 -1885
rect -120 -1905 31305 -1895
rect -120 -1945 -80 -1905
rect -40 -1945 270 -1905
rect 310 -1945 620 -1905
rect 660 -1945 970 -1905
rect 1010 -1945 1320 -1905
rect 1360 -1945 1670 -1905
rect 1710 -1945 2020 -1905
rect 2060 -1945 2370 -1905
rect 2410 -1945 2720 -1905
rect 2760 -1945 3070 -1905
rect 3110 -1945 3420 -1905
rect 3460 -1945 3770 -1905
rect 3810 -1945 4120 -1905
rect 4160 -1945 4470 -1905
rect 4510 -1945 4820 -1905
rect 4860 -1945 5170 -1905
rect 5210 -1945 5520 -1905
rect 5560 -1945 5870 -1905
rect 5910 -1945 6220 -1905
rect 6260 -1945 6570 -1905
rect 6610 -1945 6920 -1905
rect 6960 -1945 7270 -1905
rect 7310 -1945 7620 -1905
rect 7660 -1945 7970 -1905
rect 8010 -1945 8320 -1905
rect 8360 -1930 31305 -1905
rect 31340 -1930 31350 -1895
rect 31385 -1930 31395 -1895
rect 31430 -1930 31440 -1895
rect 31475 -1930 31485 -1895
rect 31520 -1930 31530 -1895
rect 31565 -1930 31575 -1895
rect 31610 -1930 31620 -1895
rect 31655 -1930 31665 -1895
rect 31700 -1930 31710 -1895
rect 31745 -1930 31755 -1895
rect 31790 -1930 31800 -1895
rect 31835 -1930 31845 -1895
rect 31880 -1930 31890 -1895
rect 31925 -1930 31935 -1895
rect 31970 -1930 31980 -1895
rect 32015 -1930 32025 -1895
rect 32060 -1930 32070 -1895
rect 32105 -1930 32115 -1895
rect 32150 -1930 32160 -1895
rect 32195 -1930 32205 -1895
rect 32240 -1930 32250 -1895
rect 32285 -1930 32295 -1895
rect 32330 -1930 32340 -1895
rect 32375 -1930 32385 -1895
rect 32420 -1930 32430 -1895
rect 32465 -1930 32475 -1895
rect 32510 -1930 32520 -1895
rect 32555 -1930 32565 -1895
rect 32600 -1930 32610 -1895
rect 32645 -1930 32655 -1895
rect 32690 -1930 32700 -1895
rect 32735 -1930 32745 -1895
rect 32780 -1930 32790 -1895
rect 32825 -1930 32835 -1895
rect 32870 -1930 32890 -1895
rect 8360 -1940 32890 -1930
rect 8360 -1945 31305 -1940
rect -120 -1975 31305 -1945
rect 31340 -1975 31350 -1940
rect 31385 -1975 31395 -1940
rect 31430 -1975 31440 -1940
rect 31475 -1975 31485 -1940
rect 31520 -1975 31530 -1940
rect 31565 -1975 31575 -1940
rect 31610 -1975 31620 -1940
rect 31655 -1975 31665 -1940
rect 31700 -1975 31710 -1940
rect 31745 -1975 31755 -1940
rect 31790 -1975 31800 -1940
rect 31835 -1975 31845 -1940
rect 31880 -1975 31890 -1940
rect 31925 -1975 31935 -1940
rect 31970 -1975 31980 -1940
rect 32015 -1975 32025 -1940
rect 32060 -1975 32070 -1940
rect 32105 -1975 32115 -1940
rect 32150 -1975 32160 -1940
rect 32195 -1975 32205 -1940
rect 32240 -1975 32250 -1940
rect 32285 -1975 32295 -1940
rect 32330 -1975 32340 -1940
rect 32375 -1975 32385 -1940
rect 32420 -1975 32430 -1940
rect 32465 -1975 32475 -1940
rect 32510 -1975 32520 -1940
rect 32555 -1975 32565 -1940
rect 32600 -1975 32610 -1940
rect 32645 -1975 32655 -1940
rect 32690 -1975 32700 -1940
rect 32735 -1975 32745 -1940
rect 32780 -1975 32790 -1940
rect 32825 -1975 32835 -1940
rect 32870 -1975 32890 -1940
rect -120 -2015 -80 -1975
rect -40 -2015 270 -1975
rect 310 -2015 620 -1975
rect 660 -2015 970 -1975
rect 1010 -2015 1320 -1975
rect 1360 -2015 1670 -1975
rect 1710 -2015 2020 -1975
rect 2060 -2015 2370 -1975
rect 2410 -2015 2720 -1975
rect 2760 -2015 3070 -1975
rect 3110 -2015 3420 -1975
rect 3460 -2015 3770 -1975
rect 3810 -2015 4120 -1975
rect 4160 -2015 4470 -1975
rect 4510 -2015 4820 -1975
rect 4860 -2015 5170 -1975
rect 5210 -2015 5520 -1975
rect 5560 -2015 5870 -1975
rect 5910 -2015 6220 -1975
rect 6260 -2015 6570 -1975
rect 6610 -2015 6920 -1975
rect 6960 -2015 7270 -1975
rect 7310 -2015 7620 -1975
rect 7660 -2015 7970 -1975
rect 8010 -2015 8320 -1975
rect 8360 -1985 32890 -1975
rect 8360 -2015 31305 -1985
rect -120 -2020 31305 -2015
rect 31340 -2020 31350 -1985
rect 31385 -2020 31395 -1985
rect 31430 -2020 31440 -1985
rect 31475 -2020 31485 -1985
rect 31520 -2020 31530 -1985
rect 31565 -2020 31575 -1985
rect 31610 -2020 31620 -1985
rect 31655 -2020 31665 -1985
rect 31700 -2020 31710 -1985
rect 31745 -2020 31755 -1985
rect 31790 -2020 31800 -1985
rect 31835 -2020 31845 -1985
rect 31880 -2020 31890 -1985
rect 31925 -2020 31935 -1985
rect 31970 -2020 31980 -1985
rect 32015 -2020 32025 -1985
rect 32060 -2020 32070 -1985
rect 32105 -2020 32115 -1985
rect 32150 -2020 32160 -1985
rect 32195 -2020 32205 -1985
rect 32240 -2020 32250 -1985
rect 32285 -2020 32295 -1985
rect 32330 -2020 32340 -1985
rect 32375 -2020 32385 -1985
rect 32420 -2020 32430 -1985
rect 32465 -2020 32475 -1985
rect 32510 -2020 32520 -1985
rect 32555 -2020 32565 -1985
rect 32600 -2020 32610 -1985
rect 32645 -2020 32655 -1985
rect 32690 -2020 32700 -1985
rect 32735 -2020 32745 -1985
rect 32780 -2020 32790 -1985
rect 32825 -2020 32835 -1985
rect 32870 -2020 32890 -1985
rect -120 -2030 32890 -2020
rect -120 -2040 31305 -2030
rect -120 -2080 -80 -2040
rect -40 -2080 270 -2040
rect 310 -2080 620 -2040
rect 660 -2080 970 -2040
rect 1010 -2080 1320 -2040
rect 1360 -2080 1670 -2040
rect 1710 -2080 2020 -2040
rect 2060 -2080 2370 -2040
rect 2410 -2080 2720 -2040
rect 2760 -2080 3070 -2040
rect 3110 -2080 3420 -2040
rect 3460 -2080 3770 -2040
rect 3810 -2080 4120 -2040
rect 4160 -2080 4470 -2040
rect 4510 -2080 4820 -2040
rect 4860 -2080 5170 -2040
rect 5210 -2080 5520 -2040
rect 5560 -2080 5870 -2040
rect 5910 -2080 6220 -2040
rect 6260 -2080 6570 -2040
rect 6610 -2080 6920 -2040
rect 6960 -2080 7270 -2040
rect 7310 -2080 7620 -2040
rect 7660 -2080 7970 -2040
rect 8010 -2080 8320 -2040
rect 8360 -2065 31305 -2040
rect 31340 -2065 31350 -2030
rect 31385 -2065 31395 -2030
rect 31430 -2065 31440 -2030
rect 31475 -2065 31485 -2030
rect 31520 -2065 31530 -2030
rect 31565 -2065 31575 -2030
rect 31610 -2065 31620 -2030
rect 31655 -2065 31665 -2030
rect 31700 -2065 31710 -2030
rect 31745 -2065 31755 -2030
rect 31790 -2065 31800 -2030
rect 31835 -2065 31845 -2030
rect 31880 -2065 31890 -2030
rect 31925 -2065 31935 -2030
rect 31970 -2065 31980 -2030
rect 32015 -2065 32025 -2030
rect 32060 -2065 32070 -2030
rect 32105 -2065 32115 -2030
rect 32150 -2065 32160 -2030
rect 32195 -2065 32205 -2030
rect 32240 -2065 32250 -2030
rect 32285 -2065 32295 -2030
rect 32330 -2065 32340 -2030
rect 32375 -2065 32385 -2030
rect 32420 -2065 32430 -2030
rect 32465 -2065 32475 -2030
rect 32510 -2065 32520 -2030
rect 32555 -2065 32565 -2030
rect 32600 -2065 32610 -2030
rect 32645 -2065 32655 -2030
rect 32690 -2065 32700 -2030
rect 32735 -2065 32745 -2030
rect 32780 -2065 32790 -2030
rect 32825 -2065 32835 -2030
rect 32870 -2065 32890 -2030
rect 8360 -2075 32890 -2065
rect 8360 -2080 31305 -2075
rect -120 -2100 31305 -2080
rect -120 -2140 -80 -2100
rect -40 -2140 270 -2100
rect 310 -2140 620 -2100
rect 660 -2140 970 -2100
rect 1010 -2140 1320 -2100
rect 1360 -2140 1670 -2100
rect 1710 -2140 2020 -2100
rect 2060 -2140 2370 -2100
rect 2410 -2140 2720 -2100
rect 2760 -2140 3070 -2100
rect 3110 -2140 3420 -2100
rect 3460 -2140 3770 -2100
rect 3810 -2140 4120 -2100
rect 4160 -2140 4470 -2100
rect 4510 -2140 4820 -2100
rect 4860 -2140 5170 -2100
rect 5210 -2140 5520 -2100
rect 5560 -2140 5870 -2100
rect 5910 -2140 6220 -2100
rect 6260 -2140 6570 -2100
rect 6610 -2140 6920 -2100
rect 6960 -2140 7270 -2100
rect 7310 -2140 7620 -2100
rect 7660 -2140 7970 -2100
rect 8010 -2140 8320 -2100
rect 8360 -2110 31305 -2100
rect 31340 -2110 31350 -2075
rect 31385 -2110 31395 -2075
rect 31430 -2110 31440 -2075
rect 31475 -2110 31485 -2075
rect 31520 -2110 31530 -2075
rect 31565 -2110 31575 -2075
rect 31610 -2110 31620 -2075
rect 31655 -2110 31665 -2075
rect 31700 -2110 31710 -2075
rect 31745 -2110 31755 -2075
rect 31790 -2110 31800 -2075
rect 31835 -2110 31845 -2075
rect 31880 -2110 31890 -2075
rect 31925 -2110 31935 -2075
rect 31970 -2110 31980 -2075
rect 32015 -2110 32025 -2075
rect 32060 -2110 32070 -2075
rect 32105 -2110 32115 -2075
rect 32150 -2110 32160 -2075
rect 32195 -2110 32205 -2075
rect 32240 -2110 32250 -2075
rect 32285 -2110 32295 -2075
rect 32330 -2110 32340 -2075
rect 32375 -2110 32385 -2075
rect 32420 -2110 32430 -2075
rect 32465 -2110 32475 -2075
rect 32510 -2110 32520 -2075
rect 32555 -2110 32565 -2075
rect 32600 -2110 32610 -2075
rect 32645 -2110 32655 -2075
rect 32690 -2110 32700 -2075
rect 32735 -2110 32745 -2075
rect 32780 -2110 32790 -2075
rect 32825 -2110 32835 -2075
rect 32870 -2110 32890 -2075
rect 8360 -2120 32890 -2110
rect 8360 -2140 31305 -2120
rect -120 -2155 31305 -2140
rect 31340 -2155 31350 -2120
rect 31385 -2155 31395 -2120
rect 31430 -2155 31440 -2120
rect 31475 -2155 31485 -2120
rect 31520 -2155 31530 -2120
rect 31565 -2155 31575 -2120
rect 31610 -2155 31620 -2120
rect 31655 -2155 31665 -2120
rect 31700 -2155 31710 -2120
rect 31745 -2155 31755 -2120
rect 31790 -2155 31800 -2120
rect 31835 -2155 31845 -2120
rect 31880 -2155 31890 -2120
rect 31925 -2155 31935 -2120
rect 31970 -2155 31980 -2120
rect 32015 -2155 32025 -2120
rect 32060 -2155 32070 -2120
rect 32105 -2155 32115 -2120
rect 32150 -2155 32160 -2120
rect 32195 -2155 32205 -2120
rect 32240 -2155 32250 -2120
rect 32285 -2155 32295 -2120
rect 32330 -2155 32340 -2120
rect 32375 -2155 32385 -2120
rect 32420 -2155 32430 -2120
rect 32465 -2155 32475 -2120
rect 32510 -2155 32520 -2120
rect 32555 -2155 32565 -2120
rect 32600 -2155 32610 -2120
rect 32645 -2155 32655 -2120
rect 32690 -2155 32700 -2120
rect 32735 -2155 32745 -2120
rect 32780 -2155 32790 -2120
rect 32825 -2155 32835 -2120
rect 32870 -2155 32890 -2120
rect -120 -2165 32890 -2155
rect -120 -2205 -80 -2165
rect -40 -2205 270 -2165
rect 310 -2205 620 -2165
rect 660 -2205 970 -2165
rect 1010 -2205 1320 -2165
rect 1360 -2205 1670 -2165
rect 1710 -2205 2020 -2165
rect 2060 -2205 2370 -2165
rect 2410 -2205 2720 -2165
rect 2760 -2205 3070 -2165
rect 3110 -2205 3420 -2165
rect 3460 -2205 3770 -2165
rect 3810 -2205 4120 -2165
rect 4160 -2205 4470 -2165
rect 4510 -2205 4820 -2165
rect 4860 -2205 5170 -2165
rect 5210 -2205 5520 -2165
rect 5560 -2205 5870 -2165
rect 5910 -2205 6220 -2165
rect 6260 -2205 6570 -2165
rect 6610 -2205 6920 -2165
rect 6960 -2205 7270 -2165
rect 7310 -2205 7620 -2165
rect 7660 -2205 7970 -2165
rect 8010 -2205 8320 -2165
rect 8360 -2200 31305 -2165
rect 31340 -2200 31350 -2165
rect 31385 -2200 31395 -2165
rect 31430 -2200 31440 -2165
rect 31475 -2200 31485 -2165
rect 31520 -2200 31530 -2165
rect 31565 -2200 31575 -2165
rect 31610 -2200 31620 -2165
rect 31655 -2200 31665 -2165
rect 31700 -2200 31710 -2165
rect 31745 -2200 31755 -2165
rect 31790 -2200 31800 -2165
rect 31835 -2200 31845 -2165
rect 31880 -2200 31890 -2165
rect 31925 -2200 31935 -2165
rect 31970 -2200 31980 -2165
rect 32015 -2200 32025 -2165
rect 32060 -2200 32070 -2165
rect 32105 -2200 32115 -2165
rect 32150 -2200 32160 -2165
rect 32195 -2200 32205 -2165
rect 32240 -2200 32250 -2165
rect 32285 -2200 32295 -2165
rect 32330 -2200 32340 -2165
rect 32375 -2200 32385 -2165
rect 32420 -2200 32430 -2165
rect 32465 -2200 32475 -2165
rect 32510 -2200 32520 -2165
rect 32555 -2200 32565 -2165
rect 32600 -2200 32610 -2165
rect 32645 -2200 32655 -2165
rect 32690 -2200 32700 -2165
rect 32735 -2200 32745 -2165
rect 32780 -2200 32790 -2165
rect 32825 -2200 32835 -2165
rect 32870 -2200 32890 -2165
rect 8360 -2205 32890 -2200
rect -120 -2210 32890 -2205
rect -120 -2235 31305 -2210
rect -120 -2275 -80 -2235
rect -40 -2275 270 -2235
rect 310 -2275 620 -2235
rect 660 -2275 970 -2235
rect 1010 -2275 1320 -2235
rect 1360 -2275 1670 -2235
rect 1710 -2275 2020 -2235
rect 2060 -2275 2370 -2235
rect 2410 -2275 2720 -2235
rect 2760 -2275 3070 -2235
rect 3110 -2275 3420 -2235
rect 3460 -2275 3770 -2235
rect 3810 -2275 4120 -2235
rect 4160 -2275 4470 -2235
rect 4510 -2275 4820 -2235
rect 4860 -2275 5170 -2235
rect 5210 -2275 5520 -2235
rect 5560 -2275 5870 -2235
rect 5910 -2275 6220 -2235
rect 6260 -2275 6570 -2235
rect 6610 -2275 6920 -2235
rect 6960 -2275 7270 -2235
rect 7310 -2275 7620 -2235
rect 7660 -2275 7970 -2235
rect 8010 -2275 8320 -2235
rect 8360 -2245 31305 -2235
rect 31340 -2245 31350 -2210
rect 31385 -2245 31395 -2210
rect 31430 -2245 31440 -2210
rect 31475 -2245 31485 -2210
rect 31520 -2245 31530 -2210
rect 31565 -2245 31575 -2210
rect 31610 -2245 31620 -2210
rect 31655 -2245 31665 -2210
rect 31700 -2245 31710 -2210
rect 31745 -2245 31755 -2210
rect 31790 -2245 31800 -2210
rect 31835 -2245 31845 -2210
rect 31880 -2245 31890 -2210
rect 31925 -2245 31935 -2210
rect 31970 -2245 31980 -2210
rect 32015 -2245 32025 -2210
rect 32060 -2245 32070 -2210
rect 32105 -2245 32115 -2210
rect 32150 -2245 32160 -2210
rect 32195 -2245 32205 -2210
rect 32240 -2245 32250 -2210
rect 32285 -2245 32295 -2210
rect 32330 -2245 32340 -2210
rect 32375 -2245 32385 -2210
rect 32420 -2245 32430 -2210
rect 32465 -2245 32475 -2210
rect 32510 -2245 32520 -2210
rect 32555 -2245 32565 -2210
rect 32600 -2245 32610 -2210
rect 32645 -2245 32655 -2210
rect 32690 -2245 32700 -2210
rect 32735 -2245 32745 -2210
rect 32780 -2245 32790 -2210
rect 32825 -2245 32835 -2210
rect 32870 -2245 32890 -2210
rect 8360 -2255 32890 -2245
rect 8360 -2275 31305 -2255
rect -120 -2290 31305 -2275
rect 31340 -2290 31350 -2255
rect 31385 -2290 31395 -2255
rect 31430 -2290 31440 -2255
rect 31475 -2290 31485 -2255
rect 31520 -2290 31530 -2255
rect 31565 -2290 31575 -2255
rect 31610 -2290 31620 -2255
rect 31655 -2290 31665 -2255
rect 31700 -2290 31710 -2255
rect 31745 -2290 31755 -2255
rect 31790 -2290 31800 -2255
rect 31835 -2290 31845 -2255
rect 31880 -2290 31890 -2255
rect 31925 -2290 31935 -2255
rect 31970 -2290 31980 -2255
rect 32015 -2290 32025 -2255
rect 32060 -2290 32070 -2255
rect 32105 -2290 32115 -2255
rect 32150 -2290 32160 -2255
rect 32195 -2290 32205 -2255
rect 32240 -2290 32250 -2255
rect 32285 -2290 32295 -2255
rect 32330 -2290 32340 -2255
rect 32375 -2290 32385 -2255
rect 32420 -2290 32430 -2255
rect 32465 -2290 32475 -2255
rect 32510 -2290 32520 -2255
rect 32555 -2290 32565 -2255
rect 32600 -2290 32610 -2255
rect 32645 -2290 32655 -2255
rect 32690 -2290 32700 -2255
rect 32735 -2290 32745 -2255
rect 32780 -2290 32790 -2255
rect 32825 -2290 32835 -2255
rect 32870 -2290 32890 -2255
rect -120 -2300 32890 -2290
rect -120 -2305 31305 -2300
rect -120 -2345 -80 -2305
rect -40 -2345 270 -2305
rect 310 -2345 620 -2305
rect 660 -2345 970 -2305
rect 1010 -2345 1320 -2305
rect 1360 -2345 1670 -2305
rect 1710 -2345 2020 -2305
rect 2060 -2345 2370 -2305
rect 2410 -2345 2720 -2305
rect 2760 -2345 3070 -2305
rect 3110 -2345 3420 -2305
rect 3460 -2345 3770 -2305
rect 3810 -2345 4120 -2305
rect 4160 -2345 4470 -2305
rect 4510 -2345 4820 -2305
rect 4860 -2345 5170 -2305
rect 5210 -2345 5520 -2305
rect 5560 -2345 5870 -2305
rect 5910 -2345 6220 -2305
rect 6260 -2345 6570 -2305
rect 6610 -2345 6920 -2305
rect 6960 -2345 7270 -2305
rect 7310 -2345 7620 -2305
rect 7660 -2345 7970 -2305
rect 8010 -2345 8320 -2305
rect 8360 -2335 31305 -2305
rect 31340 -2335 31350 -2300
rect 31385 -2335 31395 -2300
rect 31430 -2335 31440 -2300
rect 31475 -2335 31485 -2300
rect 31520 -2335 31530 -2300
rect 31565 -2335 31575 -2300
rect 31610 -2335 31620 -2300
rect 31655 -2335 31665 -2300
rect 31700 -2335 31710 -2300
rect 31745 -2335 31755 -2300
rect 31790 -2335 31800 -2300
rect 31835 -2335 31845 -2300
rect 31880 -2335 31890 -2300
rect 31925 -2335 31935 -2300
rect 31970 -2335 31980 -2300
rect 32015 -2335 32025 -2300
rect 32060 -2335 32070 -2300
rect 32105 -2335 32115 -2300
rect 32150 -2335 32160 -2300
rect 32195 -2335 32205 -2300
rect 32240 -2335 32250 -2300
rect 32285 -2335 32295 -2300
rect 32330 -2335 32340 -2300
rect 32375 -2335 32385 -2300
rect 32420 -2335 32430 -2300
rect 32465 -2335 32475 -2300
rect 32510 -2335 32520 -2300
rect 32555 -2335 32565 -2300
rect 32600 -2335 32610 -2300
rect 32645 -2335 32655 -2300
rect 32690 -2335 32700 -2300
rect 32735 -2335 32745 -2300
rect 32780 -2335 32790 -2300
rect 32825 -2335 32835 -2300
rect 32870 -2335 32890 -2300
rect 8360 -2345 32890 -2335
rect -120 -2375 31305 -2345
rect -120 -2415 -80 -2375
rect -40 -2415 270 -2375
rect 310 -2415 620 -2375
rect 660 -2415 970 -2375
rect 1010 -2415 1320 -2375
rect 1360 -2415 1670 -2375
rect 1710 -2415 2020 -2375
rect 2060 -2415 2370 -2375
rect 2410 -2415 2720 -2375
rect 2760 -2415 3070 -2375
rect 3110 -2415 3420 -2375
rect 3460 -2415 3770 -2375
rect 3810 -2415 4120 -2375
rect 4160 -2415 4470 -2375
rect 4510 -2415 4820 -2375
rect 4860 -2415 5170 -2375
rect 5210 -2415 5520 -2375
rect 5560 -2415 5870 -2375
rect 5910 -2415 6220 -2375
rect 6260 -2415 6570 -2375
rect 6610 -2415 6920 -2375
rect 6960 -2415 7270 -2375
rect 7310 -2415 7620 -2375
rect 7660 -2415 7970 -2375
rect 8010 -2415 8320 -2375
rect 8360 -2380 31305 -2375
rect 31340 -2380 31350 -2345
rect 31385 -2380 31395 -2345
rect 31430 -2380 31440 -2345
rect 31475 -2380 31485 -2345
rect 31520 -2380 31530 -2345
rect 31565 -2380 31575 -2345
rect 31610 -2380 31620 -2345
rect 31655 -2380 31665 -2345
rect 31700 -2380 31710 -2345
rect 31745 -2380 31755 -2345
rect 31790 -2380 31800 -2345
rect 31835 -2380 31845 -2345
rect 31880 -2380 31890 -2345
rect 31925 -2380 31935 -2345
rect 31970 -2380 31980 -2345
rect 32015 -2380 32025 -2345
rect 32060 -2380 32070 -2345
rect 32105 -2380 32115 -2345
rect 32150 -2380 32160 -2345
rect 32195 -2380 32205 -2345
rect 32240 -2380 32250 -2345
rect 32285 -2380 32295 -2345
rect 32330 -2380 32340 -2345
rect 32375 -2380 32385 -2345
rect 32420 -2380 32430 -2345
rect 32465 -2380 32475 -2345
rect 32510 -2380 32520 -2345
rect 32555 -2380 32565 -2345
rect 32600 -2380 32610 -2345
rect 32645 -2380 32655 -2345
rect 32690 -2380 32700 -2345
rect 32735 -2380 32745 -2345
rect 32780 -2380 32790 -2345
rect 32825 -2380 32835 -2345
rect 32870 -2380 32890 -2345
rect 8360 -2390 32890 -2380
rect 8360 -2415 31305 -2390
rect -120 -2425 31305 -2415
rect 31340 -2425 31350 -2390
rect 31385 -2425 31395 -2390
rect 31430 -2425 31440 -2390
rect 31475 -2425 31485 -2390
rect 31520 -2425 31530 -2390
rect 31565 -2425 31575 -2390
rect 31610 -2425 31620 -2390
rect 31655 -2425 31665 -2390
rect 31700 -2425 31710 -2390
rect 31745 -2425 31755 -2390
rect 31790 -2425 31800 -2390
rect 31835 -2425 31845 -2390
rect 31880 -2425 31890 -2390
rect 31925 -2425 31935 -2390
rect 31970 -2425 31980 -2390
rect 32015 -2425 32025 -2390
rect 32060 -2425 32070 -2390
rect 32105 -2425 32115 -2390
rect 32150 -2425 32160 -2390
rect 32195 -2425 32205 -2390
rect 32240 -2425 32250 -2390
rect 32285 -2425 32295 -2390
rect 32330 -2425 32340 -2390
rect 32375 -2425 32385 -2390
rect 32420 -2425 32430 -2390
rect 32465 -2425 32475 -2390
rect 32510 -2425 32520 -2390
rect 32555 -2425 32565 -2390
rect 32600 -2425 32610 -2390
rect 32645 -2425 32655 -2390
rect 32690 -2425 32700 -2390
rect 32735 -2425 32745 -2390
rect 32780 -2425 32790 -2390
rect 32825 -2425 32835 -2390
rect 32870 -2425 32890 -2390
rect -120 -2435 32890 -2425
rect -120 -2440 31305 -2435
rect -120 -2480 -80 -2440
rect -40 -2480 270 -2440
rect 310 -2480 620 -2440
rect 660 -2480 970 -2440
rect 1010 -2480 1320 -2440
rect 1360 -2480 1670 -2440
rect 1710 -2480 2020 -2440
rect 2060 -2480 2370 -2440
rect 2410 -2480 2720 -2440
rect 2760 -2480 3070 -2440
rect 3110 -2480 3420 -2440
rect 3460 -2480 3770 -2440
rect 3810 -2480 4120 -2440
rect 4160 -2480 4470 -2440
rect 4510 -2480 4820 -2440
rect 4860 -2480 5170 -2440
rect 5210 -2480 5520 -2440
rect 5560 -2480 5870 -2440
rect 5910 -2480 6220 -2440
rect 6260 -2480 6570 -2440
rect 6610 -2480 6920 -2440
rect 6960 -2480 7270 -2440
rect 7310 -2480 7620 -2440
rect 7660 -2480 7970 -2440
rect 8010 -2480 8320 -2440
rect 8360 -2470 31305 -2440
rect 31340 -2470 31350 -2435
rect 31385 -2470 31395 -2435
rect 31430 -2470 31440 -2435
rect 31475 -2470 31485 -2435
rect 31520 -2470 31530 -2435
rect 31565 -2470 31575 -2435
rect 31610 -2470 31620 -2435
rect 31655 -2470 31665 -2435
rect 31700 -2470 31710 -2435
rect 31745 -2470 31755 -2435
rect 31790 -2470 31800 -2435
rect 31835 -2470 31845 -2435
rect 31880 -2470 31890 -2435
rect 31925 -2470 31935 -2435
rect 31970 -2470 31980 -2435
rect 32015 -2470 32025 -2435
rect 32060 -2470 32070 -2435
rect 32105 -2470 32115 -2435
rect 32150 -2470 32160 -2435
rect 32195 -2470 32205 -2435
rect 32240 -2470 32250 -2435
rect 32285 -2470 32295 -2435
rect 32330 -2470 32340 -2435
rect 32375 -2470 32385 -2435
rect 32420 -2470 32430 -2435
rect 32465 -2470 32475 -2435
rect 32510 -2470 32520 -2435
rect 32555 -2470 32565 -2435
rect 32600 -2470 32610 -2435
rect 32645 -2470 32655 -2435
rect 32690 -2470 32700 -2435
rect 32735 -2470 32745 -2435
rect 32780 -2470 32790 -2435
rect 32825 -2470 32835 -2435
rect 32870 -2470 32890 -2435
rect 8360 -2480 32890 -2470
rect -120 -2500 31305 -2480
rect -120 -2540 -80 -2500
rect -40 -2540 270 -2500
rect 310 -2540 620 -2500
rect 660 -2540 970 -2500
rect 1010 -2540 1320 -2500
rect 1360 -2540 1670 -2500
rect 1710 -2540 2020 -2500
rect 2060 -2540 2370 -2500
rect 2410 -2540 2720 -2500
rect 2760 -2540 3070 -2500
rect 3110 -2540 3420 -2500
rect 3460 -2540 3770 -2500
rect 3810 -2540 4120 -2500
rect 4160 -2540 4470 -2500
rect 4510 -2540 4820 -2500
rect 4860 -2540 5170 -2500
rect 5210 -2540 5520 -2500
rect 5560 -2540 5870 -2500
rect 5910 -2540 6220 -2500
rect 6260 -2540 6570 -2500
rect 6610 -2540 6920 -2500
rect 6960 -2540 7270 -2500
rect 7310 -2540 7620 -2500
rect 7660 -2540 7970 -2500
rect 8010 -2540 8320 -2500
rect 8360 -2515 31305 -2500
rect 31340 -2515 31350 -2480
rect 31385 -2515 31395 -2480
rect 31430 -2515 31440 -2480
rect 31475 -2515 31485 -2480
rect 31520 -2515 31530 -2480
rect 31565 -2515 31575 -2480
rect 31610 -2515 31620 -2480
rect 31655 -2515 31665 -2480
rect 31700 -2515 31710 -2480
rect 31745 -2515 31755 -2480
rect 31790 -2515 31800 -2480
rect 31835 -2515 31845 -2480
rect 31880 -2515 31890 -2480
rect 31925 -2515 31935 -2480
rect 31970 -2515 31980 -2480
rect 32015 -2515 32025 -2480
rect 32060 -2515 32070 -2480
rect 32105 -2515 32115 -2480
rect 32150 -2515 32160 -2480
rect 32195 -2515 32205 -2480
rect 32240 -2515 32250 -2480
rect 32285 -2515 32295 -2480
rect 32330 -2515 32340 -2480
rect 32375 -2515 32385 -2480
rect 32420 -2515 32430 -2480
rect 32465 -2515 32475 -2480
rect 32510 -2515 32520 -2480
rect 32555 -2515 32565 -2480
rect 32600 -2515 32610 -2480
rect 32645 -2515 32655 -2480
rect 32690 -2515 32700 -2480
rect 32735 -2515 32745 -2480
rect 32780 -2515 32790 -2480
rect 32825 -2515 32835 -2480
rect 32870 -2515 32890 -2480
rect 8360 -2525 32890 -2515
rect 8360 -2540 31305 -2525
rect -120 -2560 31305 -2540
rect 31340 -2560 31350 -2525
rect 31385 -2560 31395 -2525
rect 31430 -2560 31440 -2525
rect 31475 -2560 31485 -2525
rect 31520 -2560 31530 -2525
rect 31565 -2560 31575 -2525
rect 31610 -2560 31620 -2525
rect 31655 -2560 31665 -2525
rect 31700 -2560 31710 -2525
rect 31745 -2560 31755 -2525
rect 31790 -2560 31800 -2525
rect 31835 -2560 31845 -2525
rect 31880 -2560 31890 -2525
rect 31925 -2560 31935 -2525
rect 31970 -2560 31980 -2525
rect 32015 -2560 32025 -2525
rect 32060 -2560 32070 -2525
rect 32105 -2560 32115 -2525
rect 32150 -2560 32160 -2525
rect 32195 -2560 32205 -2525
rect 32240 -2560 32250 -2525
rect 32285 -2560 32295 -2525
rect 32330 -2560 32340 -2525
rect 32375 -2560 32385 -2525
rect 32420 -2560 32430 -2525
rect 32465 -2560 32475 -2525
rect 32510 -2560 32520 -2525
rect 32555 -2560 32565 -2525
rect 32600 -2560 32610 -2525
rect 32645 -2560 32655 -2525
rect 32690 -2560 32700 -2525
rect 32735 -2560 32745 -2525
rect 32780 -2560 32790 -2525
rect 32825 -2560 32835 -2525
rect 32870 -2560 32890 -2525
rect -120 -2565 32890 -2560
rect -120 -2605 -80 -2565
rect -40 -2605 270 -2565
rect 310 -2605 620 -2565
rect 660 -2605 970 -2565
rect 1010 -2605 1320 -2565
rect 1360 -2605 1670 -2565
rect 1710 -2605 2020 -2565
rect 2060 -2605 2370 -2565
rect 2410 -2605 2720 -2565
rect 2760 -2605 3070 -2565
rect 3110 -2605 3420 -2565
rect 3460 -2605 3770 -2565
rect 3810 -2605 4120 -2565
rect 4160 -2605 4470 -2565
rect 4510 -2605 4820 -2565
rect 4860 -2605 5170 -2565
rect 5210 -2605 5520 -2565
rect 5560 -2605 5870 -2565
rect 5910 -2605 6220 -2565
rect 6260 -2605 6570 -2565
rect 6610 -2605 6920 -2565
rect 6960 -2605 7270 -2565
rect 7310 -2605 7620 -2565
rect 7660 -2605 7970 -2565
rect 8010 -2605 8320 -2565
rect 8360 -2570 32890 -2565
rect 8360 -2605 31305 -2570
rect 31340 -2605 31350 -2570
rect 31385 -2605 31395 -2570
rect 31430 -2605 31440 -2570
rect 31475 -2605 31485 -2570
rect 31520 -2605 31530 -2570
rect 31565 -2605 31575 -2570
rect 31610 -2605 31620 -2570
rect 31655 -2605 31665 -2570
rect 31700 -2605 31710 -2570
rect 31745 -2605 31755 -2570
rect 31790 -2605 31800 -2570
rect 31835 -2605 31845 -2570
rect 31880 -2605 31890 -2570
rect 31925 -2605 31935 -2570
rect 31970 -2605 31980 -2570
rect 32015 -2605 32025 -2570
rect 32060 -2605 32070 -2570
rect 32105 -2605 32115 -2570
rect 32150 -2605 32160 -2570
rect 32195 -2605 32205 -2570
rect 32240 -2605 32250 -2570
rect 32285 -2605 32295 -2570
rect 32330 -2605 32340 -2570
rect 32375 -2605 32385 -2570
rect 32420 -2605 32430 -2570
rect 32465 -2605 32475 -2570
rect 32510 -2605 32520 -2570
rect 32555 -2605 32565 -2570
rect 32600 -2605 32610 -2570
rect 32645 -2605 32655 -2570
rect 32690 -2605 32700 -2570
rect 32735 -2605 32745 -2570
rect 32780 -2605 32790 -2570
rect 32825 -2605 32835 -2570
rect 32870 -2605 32890 -2570
rect -120 -2615 32890 -2605
rect -120 -2635 31305 -2615
rect -120 -2675 -80 -2635
rect -40 -2675 270 -2635
rect 310 -2675 620 -2635
rect 660 -2675 970 -2635
rect 1010 -2675 1320 -2635
rect 1360 -2675 1670 -2635
rect 1710 -2675 2020 -2635
rect 2060 -2675 2370 -2635
rect 2410 -2675 2720 -2635
rect 2760 -2675 3070 -2635
rect 3110 -2675 3420 -2635
rect 3460 -2675 3770 -2635
rect 3810 -2675 4120 -2635
rect 4160 -2675 4470 -2635
rect 4510 -2675 4820 -2635
rect 4860 -2675 5170 -2635
rect 5210 -2675 5520 -2635
rect 5560 -2675 5870 -2635
rect 5910 -2675 6220 -2635
rect 6260 -2675 6570 -2635
rect 6610 -2675 6920 -2635
rect 6960 -2675 7270 -2635
rect 7310 -2675 7620 -2635
rect 7660 -2675 7970 -2635
rect 8010 -2675 8320 -2635
rect 8360 -2650 31305 -2635
rect 31340 -2650 31350 -2615
rect 31385 -2650 31395 -2615
rect 31430 -2650 31440 -2615
rect 31475 -2650 31485 -2615
rect 31520 -2650 31530 -2615
rect 31565 -2650 31575 -2615
rect 31610 -2650 31620 -2615
rect 31655 -2650 31665 -2615
rect 31700 -2650 31710 -2615
rect 31745 -2650 31755 -2615
rect 31790 -2650 31800 -2615
rect 31835 -2650 31845 -2615
rect 31880 -2650 31890 -2615
rect 31925 -2650 31935 -2615
rect 31970 -2650 31980 -2615
rect 32015 -2650 32025 -2615
rect 32060 -2650 32070 -2615
rect 32105 -2650 32115 -2615
rect 32150 -2650 32160 -2615
rect 32195 -2650 32205 -2615
rect 32240 -2650 32250 -2615
rect 32285 -2650 32295 -2615
rect 32330 -2650 32340 -2615
rect 32375 -2650 32385 -2615
rect 32420 -2650 32430 -2615
rect 32465 -2650 32475 -2615
rect 32510 -2650 32520 -2615
rect 32555 -2650 32565 -2615
rect 32600 -2650 32610 -2615
rect 32645 -2650 32655 -2615
rect 32690 -2650 32700 -2615
rect 32735 -2650 32745 -2615
rect 32780 -2650 32790 -2615
rect 32825 -2650 32835 -2615
rect 32870 -2650 32890 -2615
rect 8360 -2660 32890 -2650
rect 8360 -2675 31305 -2660
rect -120 -2695 31305 -2675
rect 31340 -2695 31350 -2660
rect 31385 -2695 31395 -2660
rect 31430 -2695 31440 -2660
rect 31475 -2695 31485 -2660
rect 31520 -2695 31530 -2660
rect 31565 -2695 31575 -2660
rect 31610 -2695 31620 -2660
rect 31655 -2695 31665 -2660
rect 31700 -2695 31710 -2660
rect 31745 -2695 31755 -2660
rect 31790 -2695 31800 -2660
rect 31835 -2695 31845 -2660
rect 31880 -2695 31890 -2660
rect 31925 -2695 31935 -2660
rect 31970 -2695 31980 -2660
rect 32015 -2695 32025 -2660
rect 32060 -2695 32070 -2660
rect 32105 -2695 32115 -2660
rect 32150 -2695 32160 -2660
rect 32195 -2695 32205 -2660
rect 32240 -2695 32250 -2660
rect 32285 -2695 32295 -2660
rect 32330 -2695 32340 -2660
rect 32375 -2695 32385 -2660
rect 32420 -2695 32430 -2660
rect 32465 -2695 32475 -2660
rect 32510 -2695 32520 -2660
rect 32555 -2695 32565 -2660
rect 32600 -2695 32610 -2660
rect 32645 -2695 32655 -2660
rect 32690 -2695 32700 -2660
rect 32735 -2695 32745 -2660
rect 32780 -2695 32790 -2660
rect 32825 -2695 32835 -2660
rect 32870 -2695 32890 -2660
rect -120 -2705 32890 -2695
rect -120 -2745 -80 -2705
rect -40 -2745 270 -2705
rect 310 -2745 620 -2705
rect 660 -2745 970 -2705
rect 1010 -2745 1320 -2705
rect 1360 -2745 1670 -2705
rect 1710 -2745 2020 -2705
rect 2060 -2745 2370 -2705
rect 2410 -2745 2720 -2705
rect 2760 -2745 3070 -2705
rect 3110 -2745 3420 -2705
rect 3460 -2745 3770 -2705
rect 3810 -2745 4120 -2705
rect 4160 -2745 4470 -2705
rect 4510 -2745 4820 -2705
rect 4860 -2745 5170 -2705
rect 5210 -2745 5520 -2705
rect 5560 -2745 5870 -2705
rect 5910 -2745 6220 -2705
rect 6260 -2745 6570 -2705
rect 6610 -2745 6920 -2705
rect 6960 -2745 7270 -2705
rect 7310 -2745 7620 -2705
rect 7660 -2745 7970 -2705
rect 8010 -2745 8320 -2705
rect 8360 -2740 31305 -2705
rect 31340 -2740 31350 -2705
rect 31385 -2740 31395 -2705
rect 31430 -2740 31440 -2705
rect 31475 -2740 31485 -2705
rect 31520 -2740 31530 -2705
rect 31565 -2740 31575 -2705
rect 31610 -2740 31620 -2705
rect 31655 -2740 31665 -2705
rect 31700 -2740 31710 -2705
rect 31745 -2740 31755 -2705
rect 31790 -2740 31800 -2705
rect 31835 -2740 31845 -2705
rect 31880 -2740 31890 -2705
rect 31925 -2740 31935 -2705
rect 31970 -2740 31980 -2705
rect 32015 -2740 32025 -2705
rect 32060 -2740 32070 -2705
rect 32105 -2740 32115 -2705
rect 32150 -2740 32160 -2705
rect 32195 -2740 32205 -2705
rect 32240 -2740 32250 -2705
rect 32285 -2740 32295 -2705
rect 32330 -2740 32340 -2705
rect 32375 -2740 32385 -2705
rect 32420 -2740 32430 -2705
rect 32465 -2740 32475 -2705
rect 32510 -2740 32520 -2705
rect 32555 -2740 32565 -2705
rect 32600 -2740 32610 -2705
rect 32645 -2740 32655 -2705
rect 32690 -2740 32700 -2705
rect 32735 -2740 32745 -2705
rect 32780 -2740 32790 -2705
rect 32825 -2740 32835 -2705
rect 32870 -2740 32890 -2705
rect 8360 -2745 32890 -2740
rect -120 -2750 32890 -2745
rect -120 -2775 31305 -2750
rect -120 -2815 -80 -2775
rect -40 -2815 270 -2775
rect 310 -2815 620 -2775
rect 660 -2815 970 -2775
rect 1010 -2815 1320 -2775
rect 1360 -2815 1670 -2775
rect 1710 -2815 2020 -2775
rect 2060 -2815 2370 -2775
rect 2410 -2815 2720 -2775
rect 2760 -2815 3070 -2775
rect 3110 -2815 3420 -2775
rect 3460 -2815 3770 -2775
rect 3810 -2815 4120 -2775
rect 4160 -2815 4470 -2775
rect 4510 -2815 4820 -2775
rect 4860 -2815 5170 -2775
rect 5210 -2815 5520 -2775
rect 5560 -2815 5870 -2775
rect 5910 -2815 6220 -2775
rect 6260 -2815 6570 -2775
rect 6610 -2815 6920 -2775
rect 6960 -2815 7270 -2775
rect 7310 -2815 7620 -2775
rect 7660 -2815 7970 -2775
rect 8010 -2815 8320 -2775
rect 8360 -2785 31305 -2775
rect 31340 -2785 31350 -2750
rect 31385 -2785 31395 -2750
rect 31430 -2785 31440 -2750
rect 31475 -2785 31485 -2750
rect 31520 -2785 31530 -2750
rect 31565 -2785 31575 -2750
rect 31610 -2785 31620 -2750
rect 31655 -2785 31665 -2750
rect 31700 -2785 31710 -2750
rect 31745 -2785 31755 -2750
rect 31790 -2785 31800 -2750
rect 31835 -2785 31845 -2750
rect 31880 -2785 31890 -2750
rect 31925 -2785 31935 -2750
rect 31970 -2785 31980 -2750
rect 32015 -2785 32025 -2750
rect 32060 -2785 32070 -2750
rect 32105 -2785 32115 -2750
rect 32150 -2785 32160 -2750
rect 32195 -2785 32205 -2750
rect 32240 -2785 32250 -2750
rect 32285 -2785 32295 -2750
rect 32330 -2785 32340 -2750
rect 32375 -2785 32385 -2750
rect 32420 -2785 32430 -2750
rect 32465 -2785 32475 -2750
rect 32510 -2785 32520 -2750
rect 32555 -2785 32565 -2750
rect 32600 -2785 32610 -2750
rect 32645 -2785 32655 -2750
rect 32690 -2785 32700 -2750
rect 32735 -2785 32745 -2750
rect 32780 -2785 32790 -2750
rect 32825 -2785 32835 -2750
rect 32870 -2785 32890 -2750
rect 8360 -2795 32890 -2785
rect 8360 -2815 31305 -2795
rect -120 -2830 31305 -2815
rect 31340 -2830 31350 -2795
rect 31385 -2830 31395 -2795
rect 31430 -2830 31440 -2795
rect 31475 -2830 31485 -2795
rect 31520 -2830 31530 -2795
rect 31565 -2830 31575 -2795
rect 31610 -2830 31620 -2795
rect 31655 -2830 31665 -2795
rect 31700 -2830 31710 -2795
rect 31745 -2830 31755 -2795
rect 31790 -2830 31800 -2795
rect 31835 -2830 31845 -2795
rect 31880 -2830 31890 -2795
rect 31925 -2830 31935 -2795
rect 31970 -2830 31980 -2795
rect 32015 -2830 32025 -2795
rect 32060 -2830 32070 -2795
rect 32105 -2830 32115 -2795
rect 32150 -2830 32160 -2795
rect 32195 -2830 32205 -2795
rect 32240 -2830 32250 -2795
rect 32285 -2830 32295 -2795
rect 32330 -2830 32340 -2795
rect 32375 -2830 32385 -2795
rect 32420 -2830 32430 -2795
rect 32465 -2830 32475 -2795
rect 32510 -2830 32520 -2795
rect 32555 -2830 32565 -2795
rect 32600 -2830 32610 -2795
rect 32645 -2830 32655 -2795
rect 32690 -2830 32700 -2795
rect 32735 -2830 32745 -2795
rect 32780 -2830 32790 -2795
rect 32825 -2830 32835 -2795
rect 32870 -2830 32890 -2795
rect -120 -2840 32890 -2830
rect -120 -2880 -80 -2840
rect -40 -2880 270 -2840
rect 310 -2880 620 -2840
rect 660 -2880 970 -2840
rect 1010 -2880 1320 -2840
rect 1360 -2880 1670 -2840
rect 1710 -2880 2020 -2840
rect 2060 -2880 2370 -2840
rect 2410 -2880 2720 -2840
rect 2760 -2880 3070 -2840
rect 3110 -2880 3420 -2840
rect 3460 -2880 3770 -2840
rect 3810 -2880 4120 -2840
rect 4160 -2880 4470 -2840
rect 4510 -2880 4820 -2840
rect 4860 -2880 5170 -2840
rect 5210 -2880 5520 -2840
rect 5560 -2880 5870 -2840
rect 5910 -2880 6220 -2840
rect 6260 -2880 6570 -2840
rect 6610 -2880 6920 -2840
rect 6960 -2880 7270 -2840
rect 7310 -2880 7620 -2840
rect 7660 -2880 7970 -2840
rect 8010 -2880 8320 -2840
rect 8360 -2875 31305 -2840
rect 31340 -2875 31350 -2840
rect 31385 -2875 31395 -2840
rect 31430 -2875 31440 -2840
rect 31475 -2875 31485 -2840
rect 31520 -2875 31530 -2840
rect 31565 -2875 31575 -2840
rect 31610 -2875 31620 -2840
rect 31655 -2875 31665 -2840
rect 31700 -2875 31710 -2840
rect 31745 -2875 31755 -2840
rect 31790 -2875 31800 -2840
rect 31835 -2875 31845 -2840
rect 31880 -2875 31890 -2840
rect 31925 -2875 31935 -2840
rect 31970 -2875 31980 -2840
rect 32015 -2875 32025 -2840
rect 32060 -2875 32070 -2840
rect 32105 -2875 32115 -2840
rect 32150 -2875 32160 -2840
rect 32195 -2875 32205 -2840
rect 32240 -2875 32250 -2840
rect 32285 -2875 32295 -2840
rect 32330 -2875 32340 -2840
rect 32375 -2875 32385 -2840
rect 32420 -2875 32430 -2840
rect 32465 -2875 32475 -2840
rect 32510 -2875 32520 -2840
rect 32555 -2875 32565 -2840
rect 32600 -2875 32610 -2840
rect 32645 -2875 32655 -2840
rect 32690 -2875 32700 -2840
rect 32735 -2875 32745 -2840
rect 32780 -2875 32790 -2840
rect 32825 -2875 32835 -2840
rect 32870 -2875 32890 -2840
rect 8360 -2880 32890 -2875
rect -120 -2890 32890 -2880
use bgr_11  bgr_11_0
timestamp 1755893231
transform -1 0 22290 0 -1 11375
box 15640 -6260 19905 1640
use two_stage_opamp_dummy_magic_26  two_stage_opamp_dummy_magic_26_0
timestamp 1755896001
transform 1 0 -52410 0 1 100
box 52060 -1500 61740 6110
<< labels >>
flabel metal4 35620 6650 35620 6650 3 FreeSans 800 0 320 0 GNDA
port 2 e
flabel metal3 -37570 10155 -37570 10155 1 FreeSans 800 0 0 320 VDDA
port 1 n
flabel metal2 5375 2090 5375 2090 3 FreeSans 400 0 160 0 VIN-
port 6 e
flabel metal2 3605 2090 3605 2090 7 FreeSans 400 0 -160 0 VIN+
port 5 w
flabel metal2 6795 865 6795 865 5 FreeSans 800 0 0 -400 VOUT-
port 4 s
flabel metal2 2185 865 2185 865 5 FreeSans 800 0 0 -400 VOUT+
port 3 s
<< end >>
