magic
tech sky130A
timestamp 1749438161
<< nwell >>
rect 2545 1880 5285 2950
<< pwell >>
rect 16240 4340 16460 4403
rect 16570 4340 16970 4420
rect 17080 4335 17600 4395
rect 16250 4105 17500 4155
rect 16195 3800 16895 3850
rect 16935 3800 17635 3850
rect 15155 2985 15855 3585
rect 16220 3175 17580 3575
rect 17945 2985 18645 3585
rect 15155 2455 15855 2655
rect 16220 2495 17580 2895
rect 17945 2455 18645 2655
rect 15155 1965 15855 2265
rect 16275 1980 17525 2130
rect 17945 1965 18645 2265
rect -45 1685 130 1725
rect 3165 1615 3805 1665
rect 4205 1615 4845 1665
rect 2835 1205 3955 1455
rect 4055 1205 5175 1455
rect 2945 975 5065 1075
rect 15155 955 15795 1655
rect 16030 1515 16730 1665
rect 16770 1515 17030 1665
rect 17070 1515 17770 1665
rect 16205 935 17620 1185
rect 18005 955 18645 1655
rect 2995 780 5015 880
rect 16260 645 16530 745
rect 16880 700 17580 750
<< nmos >>
rect 16280 4340 16300 4403
rect 16340 4340 16360 4403
rect 16400 4340 16420 4403
rect 16610 4340 16630 4420
rect 16670 4340 16690 4420
rect 16730 4340 16750 4420
rect 16790 4340 16810 4420
rect 16850 4340 16870 4420
rect 16910 4340 16930 4420
rect 17120 4335 17140 4395
rect 17180 4335 17200 4395
rect 17240 4335 17260 4395
rect 17300 4335 17320 4395
rect 17360 4335 17380 4395
rect 17420 4335 17440 4395
rect 17480 4335 17500 4395
rect 17540 4335 17560 4395
rect 16290 4105 16305 4155
rect 16345 4105 16360 4155
rect 16400 4105 16415 4155
rect 16455 4105 16470 4155
rect 16510 4105 16525 4155
rect 16565 4105 16580 4155
rect 16620 4105 16635 4155
rect 16675 4105 16690 4155
rect 16730 4105 16745 4155
rect 16785 4105 16800 4155
rect 16840 4105 16855 4155
rect 16895 4105 16910 4155
rect 16950 4105 16965 4155
rect 17005 4105 17020 4155
rect 17060 4105 17075 4155
rect 17115 4105 17130 4155
rect 17170 4105 17185 4155
rect 17225 4105 17240 4155
rect 17280 4105 17295 4155
rect 17335 4105 17350 4155
rect 17390 4105 17405 4155
rect 17445 4105 17460 4155
rect 16235 3800 16250 3850
rect 16290 3800 16305 3850
rect 16345 3800 16360 3850
rect 16400 3800 16415 3850
rect 16455 3800 16470 3850
rect 16510 3800 16525 3850
rect 16565 3800 16580 3850
rect 16620 3800 16635 3850
rect 16675 3800 16690 3850
rect 16730 3800 16745 3850
rect 16785 3800 16800 3850
rect 16840 3800 16855 3850
rect 16975 3800 16990 3850
rect 17030 3800 17045 3850
rect 17085 3800 17100 3850
rect 17140 3800 17155 3850
rect 17195 3800 17210 3850
rect 17250 3800 17265 3850
rect 17305 3800 17320 3850
rect 17360 3800 17375 3850
rect 17415 3800 17430 3850
rect 17470 3800 17485 3850
rect 17525 3800 17540 3850
rect 17580 3800 17595 3850
rect 15195 2985 15210 3585
rect 15250 2985 15265 3585
rect 15305 2985 15320 3585
rect 15360 2985 15375 3585
rect 15415 2985 15430 3585
rect 15470 2985 15485 3585
rect 15525 2985 15540 3585
rect 15580 2985 15595 3585
rect 15635 2985 15650 3585
rect 15690 2985 15705 3585
rect 15745 2985 15760 3585
rect 15800 2985 15815 3585
rect 16260 3175 16280 3575
rect 16320 3175 16340 3575
rect 16380 3175 16400 3575
rect 16440 3175 16460 3575
rect 16500 3175 16520 3575
rect 16560 3175 16580 3575
rect 16620 3175 16640 3575
rect 16680 3175 16700 3575
rect 16740 3175 16760 3575
rect 16800 3175 16820 3575
rect 16860 3175 16880 3575
rect 16920 3175 16940 3575
rect 16980 3175 17000 3575
rect 17040 3175 17060 3575
rect 17100 3175 17120 3575
rect 17160 3175 17180 3575
rect 17220 3175 17240 3575
rect 17280 3175 17300 3575
rect 17340 3175 17360 3575
rect 17400 3175 17420 3575
rect 17460 3175 17480 3575
rect 17520 3175 17540 3575
rect 17985 2985 18000 3585
rect 18040 2985 18055 3585
rect 18095 2985 18110 3585
rect 18150 2985 18165 3585
rect 18205 2985 18220 3585
rect 18260 2985 18275 3585
rect 18315 2985 18330 3585
rect 18370 2985 18385 3585
rect 18425 2985 18440 3585
rect 18480 2985 18495 3585
rect 18535 2985 18550 3585
rect 18590 2985 18605 3585
rect 15195 2455 15210 2655
rect 15250 2455 15265 2655
rect 15305 2455 15320 2655
rect 15360 2455 15375 2655
rect 15415 2455 15430 2655
rect 15470 2455 15485 2655
rect 15525 2455 15540 2655
rect 15580 2455 15595 2655
rect 15635 2455 15650 2655
rect 15690 2455 15705 2655
rect 15745 2455 15760 2655
rect 15800 2455 15815 2655
rect 16260 2495 16280 2895
rect 16320 2495 16340 2895
rect 16380 2495 16400 2895
rect 16440 2495 16460 2895
rect 16500 2495 16520 2895
rect 16560 2495 16580 2895
rect 16620 2495 16640 2895
rect 16680 2495 16700 2895
rect 16740 2495 16760 2895
rect 16800 2495 16820 2895
rect 16860 2495 16880 2895
rect 16920 2495 16940 2895
rect 16980 2495 17000 2895
rect 17040 2495 17060 2895
rect 17100 2495 17120 2895
rect 17160 2495 17180 2895
rect 17220 2495 17240 2895
rect 17280 2495 17300 2895
rect 17340 2495 17360 2895
rect 17400 2495 17420 2895
rect 17460 2495 17480 2895
rect 17520 2495 17540 2895
rect 17985 2455 18000 2655
rect 18040 2455 18055 2655
rect 18095 2455 18110 2655
rect 18150 2455 18165 2655
rect 18205 2455 18220 2655
rect 18260 2455 18275 2655
rect 18315 2455 18330 2655
rect 18370 2455 18385 2655
rect 18425 2455 18440 2655
rect 18480 2455 18495 2655
rect 18535 2455 18550 2655
rect 18590 2455 18605 2655
rect 15195 1965 15210 2265
rect 15250 1965 15265 2265
rect 15305 1965 15320 2265
rect 15360 1965 15375 2265
rect 15415 1965 15430 2265
rect 15470 1965 15485 2265
rect 15525 1965 15540 2265
rect 15580 1965 15595 2265
rect 15635 1965 15650 2265
rect 15690 1965 15705 2265
rect 15745 1965 15760 2265
rect 15800 1965 15815 2265
rect 16315 1980 16330 2130
rect 16370 1980 16385 2130
rect 16425 1980 16440 2130
rect 16480 1980 16495 2130
rect 16535 1980 16550 2130
rect 16590 1980 16605 2130
rect 16645 1980 16660 2130
rect 16700 1980 16715 2130
rect 16755 1980 16770 2130
rect 16810 1980 16825 2130
rect 16865 1980 16880 2130
rect 16920 1980 16935 2130
rect 16975 1980 16990 2130
rect 17030 1980 17045 2130
rect 17085 1980 17100 2130
rect 17140 1980 17155 2130
rect 17195 1980 17210 2130
rect 17250 1980 17265 2130
rect 17305 1980 17320 2130
rect 17360 1980 17375 2130
rect 17415 1980 17430 2130
rect 17470 1980 17485 2130
rect 17985 1965 18000 2265
rect 18040 1965 18055 2265
rect 18095 1965 18110 2265
rect 18150 1965 18165 2265
rect 18205 1965 18220 2265
rect 18260 1965 18275 2265
rect 18315 1965 18330 2265
rect 18370 1965 18385 2265
rect 18425 1965 18440 2265
rect 18480 1965 18495 2265
rect 18535 1965 18550 2265
rect 18590 1965 18605 2265
rect 3205 1615 3225 1665
rect 3265 1615 3285 1665
rect 3325 1615 3345 1665
rect 3385 1615 3405 1665
rect 3445 1615 3465 1665
rect 3505 1615 3525 1665
rect 3565 1615 3585 1665
rect 3625 1615 3645 1665
rect 3685 1615 3705 1665
rect 3745 1615 3765 1665
rect 4245 1615 4265 1665
rect 4305 1615 4325 1665
rect 4365 1615 4385 1665
rect 4425 1615 4445 1665
rect 4485 1615 4505 1665
rect 4545 1615 4565 1665
rect 4605 1615 4625 1665
rect 4665 1615 4685 1665
rect 4725 1615 4745 1665
rect 4785 1615 4805 1665
rect 2875 1205 3375 1455
rect 3415 1205 3915 1455
rect 4095 1205 4595 1455
rect 4635 1205 5135 1455
rect 2985 975 3985 1075
rect 4025 975 5025 1075
rect 15195 955 15255 1655
rect 15295 955 15355 1655
rect 15395 955 15455 1655
rect 15495 955 15555 1655
rect 15595 955 15655 1655
rect 15695 955 15755 1655
rect 16070 1515 16085 1665
rect 16125 1515 16140 1665
rect 16180 1515 16195 1665
rect 16235 1515 16250 1665
rect 16290 1515 16305 1665
rect 16345 1515 16360 1665
rect 16400 1515 16415 1665
rect 16455 1515 16470 1665
rect 16510 1515 16525 1665
rect 16565 1515 16580 1665
rect 16620 1515 16635 1665
rect 16675 1515 16690 1665
rect 16810 1515 16825 1665
rect 16865 1515 16880 1665
rect 16920 1515 16935 1665
rect 16975 1515 16990 1665
rect 17110 1515 17125 1665
rect 17165 1515 17180 1665
rect 17220 1515 17235 1665
rect 17275 1515 17290 1665
rect 17330 1515 17345 1665
rect 17385 1515 17400 1665
rect 17440 1515 17455 1665
rect 17495 1515 17510 1665
rect 17550 1515 17565 1665
rect 17605 1515 17620 1665
rect 17660 1515 17675 1665
rect 17715 1515 17730 1665
rect 16245 935 16260 1185
rect 16300 935 16315 1185
rect 16355 935 16370 1185
rect 16410 935 16425 1185
rect 16465 935 16480 1185
rect 16520 935 16535 1185
rect 16575 935 16590 1185
rect 16630 935 16645 1185
rect 16685 935 16700 1185
rect 16740 935 16755 1185
rect 16795 935 16810 1185
rect 16850 935 16865 1185
rect 16905 935 16920 1185
rect 16960 935 16975 1185
rect 17015 935 17030 1185
rect 17070 935 17085 1185
rect 17125 935 17140 1185
rect 17180 935 17195 1185
rect 17235 935 17250 1185
rect 17290 935 17305 1185
rect 17345 935 17360 1185
rect 17400 935 17415 1185
rect 17455 935 17470 1185
rect 17510 935 17525 1185
rect 17565 935 17580 1185
rect 18045 955 18105 1655
rect 18145 955 18205 1655
rect 18245 955 18305 1655
rect 18345 955 18405 1655
rect 18445 955 18505 1655
rect 18545 955 18605 1655
rect 3035 780 3085 880
rect 3125 780 3175 880
rect 3215 780 3265 880
rect 3305 780 3355 880
rect 3395 780 3445 880
rect 3485 780 3535 880
rect 3575 780 3625 880
rect 3665 780 3715 880
rect 3755 780 3805 880
rect 3845 780 3895 880
rect 3935 780 3985 880
rect 4025 780 4075 880
rect 4115 780 4165 880
rect 4205 780 4255 880
rect 4295 780 4345 880
rect 4385 780 4435 880
rect 4475 780 4525 880
rect 4565 780 4615 880
rect 4655 780 4705 880
rect 4745 780 4795 880
rect 4835 780 4885 880
rect 4925 780 4975 880
rect 16300 645 16490 745
rect 16920 700 16935 750
rect 16975 700 16990 750
rect 17030 700 17045 750
rect 17085 700 17100 750
rect 17140 700 17155 750
rect 17195 700 17210 750
rect 17250 700 17265 750
rect 17305 700 17320 750
rect 17360 700 17375 750
rect 17415 700 17430 750
rect 17470 700 17485 750
rect 17525 700 17540 750
<< pmos >>
rect 3035 2830 3085 2930
rect 3125 2830 3175 2930
rect 3215 2830 3265 2930
rect 3305 2830 3355 2930
rect 3395 2830 3445 2930
rect 3485 2830 3535 2930
rect 3575 2830 3625 2930
rect 3665 2830 3715 2930
rect 3755 2830 3805 2930
rect 3845 2830 3895 2930
rect 3935 2830 3985 2930
rect 4025 2830 4075 2930
rect 4115 2830 4165 2930
rect 4205 2830 4255 2930
rect 4295 2830 4345 2930
rect 4385 2830 4435 2930
rect 4475 2830 4525 2930
rect 4565 2830 4615 2930
rect 4655 2830 4705 2930
rect 4745 2830 4795 2930
rect 4835 2830 4885 2930
rect 4925 2830 4975 2930
rect 3215 2400 3265 2700
rect 3305 2400 3355 2700
rect 3395 2400 3445 2700
rect 3485 2400 3535 2700
rect 3575 2400 3625 2700
rect 3665 2400 3715 2700
rect 3755 2400 3805 2700
rect 3845 2400 3895 2700
rect 3935 2400 3985 2700
rect 4025 2400 4075 2700
rect 4115 2400 4165 2700
rect 4205 2400 4255 2700
rect 4295 2400 4345 2700
rect 4385 2400 4435 2700
rect 4475 2400 4525 2700
rect 4565 2400 4615 2700
rect 4655 2400 4705 2700
rect 4745 2400 4795 2700
rect 2605 1900 2620 2000
rect 2660 1900 2675 2000
rect 2785 1900 2805 2000
rect 2845 1900 2865 2000
rect 2905 1900 2925 2000
rect 2965 1900 2985 2000
rect 3025 1900 3045 2000
rect 3085 1900 3105 2000
rect 3145 1900 3165 2000
rect 3205 1900 3225 2000
rect 3265 1900 3285 2000
rect 3325 1900 3345 2000
rect 3385 1900 3405 2000
rect 3445 1900 3465 2000
rect 3505 1900 3525 2000
rect 3565 1900 3585 2000
rect 3625 1900 3645 2000
rect 3685 1900 3705 2000
rect 3745 1900 3765 2000
rect 3805 1900 3825 2000
rect 3865 1900 3885 2000
rect 3925 1900 3945 2000
rect 4065 1900 4085 2000
rect 4125 1900 4145 2000
rect 4185 1900 4205 2000
rect 4245 1900 4265 2000
rect 4305 1900 4325 2000
rect 4365 1900 4385 2000
rect 4425 1900 4445 2000
rect 4485 1900 4505 2000
rect 4545 1900 4565 2000
rect 4605 1900 4625 2000
rect 4665 1900 4685 2000
rect 4725 1900 4745 2000
rect 4785 1900 4805 2000
rect 4845 1900 4865 2000
rect 4905 1900 4925 2000
rect 4965 1900 4985 2000
rect 5025 1900 5045 2000
rect 5085 1900 5105 2000
rect 5145 1900 5165 2000
rect 5205 1900 5225 2000
<< ndiff >>
rect 16240 4375 16280 4403
rect 16240 4355 16250 4375
rect 16270 4355 16280 4375
rect 16240 4340 16280 4355
rect 16300 4380 16340 4403
rect 16300 4360 16310 4380
rect 16330 4360 16340 4380
rect 16300 4340 16340 4360
rect 16360 4380 16400 4403
rect 16360 4360 16370 4380
rect 16390 4360 16400 4380
rect 16360 4340 16400 4360
rect 16420 4375 16460 4403
rect 16420 4355 16430 4375
rect 16450 4355 16460 4375
rect 16420 4340 16460 4355
rect 16570 4390 16610 4420
rect 16570 4370 16580 4390
rect 16600 4370 16610 4390
rect 16570 4340 16610 4370
rect 16630 4390 16670 4420
rect 16630 4370 16640 4390
rect 16660 4370 16670 4390
rect 16630 4340 16670 4370
rect 16690 4390 16730 4420
rect 16690 4370 16700 4390
rect 16720 4370 16730 4390
rect 16690 4340 16730 4370
rect 16750 4390 16790 4420
rect 16750 4370 16760 4390
rect 16780 4370 16790 4390
rect 16750 4340 16790 4370
rect 16810 4390 16850 4420
rect 16810 4370 16820 4390
rect 16840 4370 16850 4390
rect 16810 4340 16850 4370
rect 16870 4390 16910 4420
rect 16870 4370 16880 4390
rect 16900 4370 16910 4390
rect 16870 4340 16910 4370
rect 16930 4390 16970 4420
rect 16930 4370 16940 4390
rect 16960 4370 16970 4390
rect 16930 4340 16970 4370
rect 17080 4375 17120 4395
rect 17080 4355 17090 4375
rect 17110 4355 17120 4375
rect 17080 4335 17120 4355
rect 17140 4375 17180 4395
rect 17140 4355 17150 4375
rect 17170 4355 17180 4375
rect 17140 4335 17180 4355
rect 17200 4375 17240 4395
rect 17200 4355 17210 4375
rect 17230 4355 17240 4375
rect 17200 4335 17240 4355
rect 17260 4375 17300 4395
rect 17260 4355 17270 4375
rect 17290 4355 17300 4375
rect 17260 4335 17300 4355
rect 17320 4375 17360 4395
rect 17320 4355 17330 4375
rect 17350 4355 17360 4375
rect 17320 4335 17360 4355
rect 17380 4375 17420 4395
rect 17380 4355 17390 4375
rect 17410 4355 17420 4375
rect 17380 4335 17420 4355
rect 17440 4375 17480 4395
rect 17440 4355 17450 4375
rect 17470 4355 17480 4375
rect 17440 4335 17480 4355
rect 17500 4375 17540 4395
rect 17500 4355 17510 4375
rect 17530 4355 17540 4375
rect 17500 4335 17540 4355
rect 17560 4375 17600 4395
rect 17560 4355 17570 4375
rect 17590 4355 17600 4375
rect 17560 4335 17600 4355
rect 16250 4140 16290 4155
rect 16250 4120 16260 4140
rect 16280 4120 16290 4140
rect 16250 4105 16290 4120
rect 16305 4140 16345 4155
rect 16305 4120 16315 4140
rect 16335 4120 16345 4140
rect 16305 4105 16345 4120
rect 16360 4140 16400 4155
rect 16360 4120 16370 4140
rect 16390 4120 16400 4140
rect 16360 4105 16400 4120
rect 16415 4140 16455 4155
rect 16415 4120 16425 4140
rect 16445 4120 16455 4140
rect 16415 4105 16455 4120
rect 16470 4140 16510 4155
rect 16470 4120 16480 4140
rect 16500 4120 16510 4140
rect 16470 4105 16510 4120
rect 16525 4140 16565 4155
rect 16525 4120 16535 4140
rect 16555 4120 16565 4140
rect 16525 4105 16565 4120
rect 16580 4140 16620 4155
rect 16580 4120 16590 4140
rect 16610 4120 16620 4140
rect 16580 4105 16620 4120
rect 16635 4140 16675 4155
rect 16635 4120 16645 4140
rect 16665 4120 16675 4140
rect 16635 4105 16675 4120
rect 16690 4140 16730 4155
rect 16690 4120 16700 4140
rect 16720 4120 16730 4140
rect 16690 4105 16730 4120
rect 16745 4140 16785 4155
rect 16745 4120 16755 4140
rect 16775 4120 16785 4140
rect 16745 4105 16785 4120
rect 16800 4140 16840 4155
rect 16800 4120 16810 4140
rect 16830 4120 16840 4140
rect 16800 4105 16840 4120
rect 16855 4140 16895 4155
rect 16855 4120 16865 4140
rect 16885 4120 16895 4140
rect 16855 4105 16895 4120
rect 16910 4140 16950 4155
rect 16910 4120 16920 4140
rect 16940 4120 16950 4140
rect 16910 4105 16950 4120
rect 16965 4140 17005 4155
rect 16965 4120 16975 4140
rect 16995 4120 17005 4140
rect 16965 4105 17005 4120
rect 17020 4140 17060 4155
rect 17020 4120 17030 4140
rect 17050 4120 17060 4140
rect 17020 4105 17060 4120
rect 17075 4140 17115 4155
rect 17075 4120 17085 4140
rect 17105 4120 17115 4140
rect 17075 4105 17115 4120
rect 17130 4140 17170 4155
rect 17130 4120 17140 4140
rect 17160 4120 17170 4140
rect 17130 4105 17170 4120
rect 17185 4140 17225 4155
rect 17185 4120 17195 4140
rect 17215 4120 17225 4140
rect 17185 4105 17225 4120
rect 17240 4140 17280 4155
rect 17240 4120 17250 4140
rect 17270 4120 17280 4140
rect 17240 4105 17280 4120
rect 17295 4140 17335 4155
rect 17295 4120 17305 4140
rect 17325 4120 17335 4140
rect 17295 4105 17335 4120
rect 17350 4140 17390 4155
rect 17350 4120 17360 4140
rect 17380 4120 17390 4140
rect 17350 4105 17390 4120
rect 17405 4140 17445 4155
rect 17405 4120 17415 4140
rect 17435 4120 17445 4140
rect 17405 4105 17445 4120
rect 17460 4140 17500 4155
rect 17460 4120 17470 4140
rect 17490 4120 17500 4140
rect 17460 4105 17500 4120
rect 16195 3835 16235 3850
rect 16195 3815 16205 3835
rect 16225 3815 16235 3835
rect 16195 3800 16235 3815
rect 16250 3835 16290 3850
rect 16250 3815 16260 3835
rect 16280 3815 16290 3835
rect 16250 3800 16290 3815
rect 16305 3835 16345 3850
rect 16305 3815 16315 3835
rect 16335 3815 16345 3835
rect 16305 3800 16345 3815
rect 16360 3835 16400 3850
rect 16360 3815 16370 3835
rect 16390 3815 16400 3835
rect 16360 3800 16400 3815
rect 16415 3835 16455 3850
rect 16415 3815 16425 3835
rect 16445 3815 16455 3835
rect 16415 3800 16455 3815
rect 16470 3835 16510 3850
rect 16470 3815 16480 3835
rect 16500 3815 16510 3835
rect 16470 3800 16510 3815
rect 16525 3835 16565 3850
rect 16525 3815 16535 3835
rect 16555 3815 16565 3835
rect 16525 3800 16565 3815
rect 16580 3835 16620 3850
rect 16580 3815 16590 3835
rect 16610 3815 16620 3835
rect 16580 3800 16620 3815
rect 16635 3835 16675 3850
rect 16635 3815 16645 3835
rect 16665 3815 16675 3835
rect 16635 3800 16675 3815
rect 16690 3835 16730 3850
rect 16690 3815 16700 3835
rect 16720 3815 16730 3835
rect 16690 3800 16730 3815
rect 16745 3835 16785 3850
rect 16745 3815 16755 3835
rect 16775 3815 16785 3835
rect 16745 3800 16785 3815
rect 16800 3835 16840 3850
rect 16800 3815 16810 3835
rect 16830 3815 16840 3835
rect 16800 3800 16840 3815
rect 16855 3835 16895 3850
rect 16935 3835 16975 3850
rect 16855 3815 16865 3835
rect 16885 3815 16895 3835
rect 16935 3815 16945 3835
rect 16965 3815 16975 3835
rect 16855 3800 16895 3815
rect 16935 3800 16975 3815
rect 16990 3835 17030 3850
rect 16990 3815 17000 3835
rect 17020 3815 17030 3835
rect 16990 3800 17030 3815
rect 17045 3835 17085 3850
rect 17045 3815 17055 3835
rect 17075 3815 17085 3835
rect 17045 3800 17085 3815
rect 17100 3835 17140 3850
rect 17100 3815 17110 3835
rect 17130 3815 17140 3835
rect 17100 3800 17140 3815
rect 17155 3835 17195 3850
rect 17155 3815 17165 3835
rect 17185 3815 17195 3835
rect 17155 3800 17195 3815
rect 17210 3835 17250 3850
rect 17210 3815 17220 3835
rect 17240 3815 17250 3835
rect 17210 3800 17250 3815
rect 17265 3835 17305 3850
rect 17265 3815 17275 3835
rect 17295 3815 17305 3835
rect 17265 3800 17305 3815
rect 17320 3835 17360 3850
rect 17320 3815 17330 3835
rect 17350 3815 17360 3835
rect 17320 3800 17360 3815
rect 17375 3835 17415 3850
rect 17375 3815 17385 3835
rect 17405 3815 17415 3835
rect 17375 3800 17415 3815
rect 17430 3835 17470 3850
rect 17430 3815 17440 3835
rect 17460 3815 17470 3835
rect 17430 3800 17470 3815
rect 17485 3835 17525 3850
rect 17485 3815 17495 3835
rect 17515 3815 17525 3835
rect 17485 3800 17525 3815
rect 17540 3835 17580 3850
rect 17540 3815 17550 3835
rect 17570 3815 17580 3835
rect 17540 3800 17580 3815
rect 17595 3835 17635 3850
rect 17595 3815 17605 3835
rect 17625 3815 17635 3835
rect 17595 3800 17635 3815
rect 15155 3570 15195 3585
rect 15155 3550 15165 3570
rect 15185 3550 15195 3570
rect 15155 3520 15195 3550
rect 15155 3500 15165 3520
rect 15185 3500 15195 3520
rect 15155 3470 15195 3500
rect 15155 3450 15165 3470
rect 15185 3450 15195 3470
rect 15155 3420 15195 3450
rect 15155 3400 15165 3420
rect 15185 3400 15195 3420
rect 15155 3370 15195 3400
rect 15155 3350 15165 3370
rect 15185 3350 15195 3370
rect 15155 3320 15195 3350
rect 15155 3300 15165 3320
rect 15185 3300 15195 3320
rect 15155 3270 15195 3300
rect 15155 3250 15165 3270
rect 15185 3250 15195 3270
rect 15155 3220 15195 3250
rect 15155 3200 15165 3220
rect 15185 3200 15195 3220
rect 15155 3170 15195 3200
rect 15155 3150 15165 3170
rect 15185 3150 15195 3170
rect 15155 3120 15195 3150
rect 15155 3100 15165 3120
rect 15185 3100 15195 3120
rect 15155 3070 15195 3100
rect 15155 3050 15165 3070
rect 15185 3050 15195 3070
rect 15155 3020 15195 3050
rect 15155 3000 15165 3020
rect 15185 3000 15195 3020
rect 15155 2985 15195 3000
rect 15210 3570 15250 3585
rect 15210 3550 15220 3570
rect 15240 3550 15250 3570
rect 15210 3520 15250 3550
rect 15210 3500 15220 3520
rect 15240 3500 15250 3520
rect 15210 3470 15250 3500
rect 15210 3450 15220 3470
rect 15240 3450 15250 3470
rect 15210 3420 15250 3450
rect 15210 3400 15220 3420
rect 15240 3400 15250 3420
rect 15210 3370 15250 3400
rect 15210 3350 15220 3370
rect 15240 3350 15250 3370
rect 15210 3320 15250 3350
rect 15210 3300 15220 3320
rect 15240 3300 15250 3320
rect 15210 3270 15250 3300
rect 15210 3250 15220 3270
rect 15240 3250 15250 3270
rect 15210 3220 15250 3250
rect 15210 3200 15220 3220
rect 15240 3200 15250 3220
rect 15210 3170 15250 3200
rect 15210 3150 15220 3170
rect 15240 3150 15250 3170
rect 15210 3120 15250 3150
rect 15210 3100 15220 3120
rect 15240 3100 15250 3120
rect 15210 3070 15250 3100
rect 15210 3050 15220 3070
rect 15240 3050 15250 3070
rect 15210 3020 15250 3050
rect 15210 3000 15220 3020
rect 15240 3000 15250 3020
rect 15210 2985 15250 3000
rect 15265 3570 15305 3585
rect 15265 3550 15275 3570
rect 15295 3550 15305 3570
rect 15265 3520 15305 3550
rect 15265 3500 15275 3520
rect 15295 3500 15305 3520
rect 15265 3470 15305 3500
rect 15265 3450 15275 3470
rect 15295 3450 15305 3470
rect 15265 3420 15305 3450
rect 15265 3400 15275 3420
rect 15295 3400 15305 3420
rect 15265 3370 15305 3400
rect 15265 3350 15275 3370
rect 15295 3350 15305 3370
rect 15265 3320 15305 3350
rect 15265 3300 15275 3320
rect 15295 3300 15305 3320
rect 15265 3270 15305 3300
rect 15265 3250 15275 3270
rect 15295 3250 15305 3270
rect 15265 3220 15305 3250
rect 15265 3200 15275 3220
rect 15295 3200 15305 3220
rect 15265 3170 15305 3200
rect 15265 3150 15275 3170
rect 15295 3150 15305 3170
rect 15265 3120 15305 3150
rect 15265 3100 15275 3120
rect 15295 3100 15305 3120
rect 15265 3070 15305 3100
rect 15265 3050 15275 3070
rect 15295 3050 15305 3070
rect 15265 3020 15305 3050
rect 15265 3000 15275 3020
rect 15295 3000 15305 3020
rect 15265 2985 15305 3000
rect 15320 3570 15360 3585
rect 15320 3550 15330 3570
rect 15350 3550 15360 3570
rect 15320 3520 15360 3550
rect 15320 3500 15330 3520
rect 15350 3500 15360 3520
rect 15320 3470 15360 3500
rect 15320 3450 15330 3470
rect 15350 3450 15360 3470
rect 15320 3420 15360 3450
rect 15320 3400 15330 3420
rect 15350 3400 15360 3420
rect 15320 3370 15360 3400
rect 15320 3350 15330 3370
rect 15350 3350 15360 3370
rect 15320 3320 15360 3350
rect 15320 3300 15330 3320
rect 15350 3300 15360 3320
rect 15320 3270 15360 3300
rect 15320 3250 15330 3270
rect 15350 3250 15360 3270
rect 15320 3220 15360 3250
rect 15320 3200 15330 3220
rect 15350 3200 15360 3220
rect 15320 3170 15360 3200
rect 15320 3150 15330 3170
rect 15350 3150 15360 3170
rect 15320 3120 15360 3150
rect 15320 3100 15330 3120
rect 15350 3100 15360 3120
rect 15320 3070 15360 3100
rect 15320 3050 15330 3070
rect 15350 3050 15360 3070
rect 15320 3020 15360 3050
rect 15320 3000 15330 3020
rect 15350 3000 15360 3020
rect 15320 2985 15360 3000
rect 15375 3570 15415 3585
rect 15375 3550 15385 3570
rect 15405 3550 15415 3570
rect 15375 3520 15415 3550
rect 15375 3500 15385 3520
rect 15405 3500 15415 3520
rect 15375 3470 15415 3500
rect 15375 3450 15385 3470
rect 15405 3450 15415 3470
rect 15375 3420 15415 3450
rect 15375 3400 15385 3420
rect 15405 3400 15415 3420
rect 15375 3370 15415 3400
rect 15375 3350 15385 3370
rect 15405 3350 15415 3370
rect 15375 3320 15415 3350
rect 15375 3300 15385 3320
rect 15405 3300 15415 3320
rect 15375 3270 15415 3300
rect 15375 3250 15385 3270
rect 15405 3250 15415 3270
rect 15375 3220 15415 3250
rect 15375 3200 15385 3220
rect 15405 3200 15415 3220
rect 15375 3170 15415 3200
rect 15375 3150 15385 3170
rect 15405 3150 15415 3170
rect 15375 3120 15415 3150
rect 15375 3100 15385 3120
rect 15405 3100 15415 3120
rect 15375 3070 15415 3100
rect 15375 3050 15385 3070
rect 15405 3050 15415 3070
rect 15375 3020 15415 3050
rect 15375 3000 15385 3020
rect 15405 3000 15415 3020
rect 15375 2985 15415 3000
rect 15430 3570 15470 3585
rect 15430 3550 15440 3570
rect 15460 3550 15470 3570
rect 15430 3520 15470 3550
rect 15430 3500 15440 3520
rect 15460 3500 15470 3520
rect 15430 3470 15470 3500
rect 15430 3450 15440 3470
rect 15460 3450 15470 3470
rect 15430 3420 15470 3450
rect 15430 3400 15440 3420
rect 15460 3400 15470 3420
rect 15430 3370 15470 3400
rect 15430 3350 15440 3370
rect 15460 3350 15470 3370
rect 15430 3320 15470 3350
rect 15430 3300 15440 3320
rect 15460 3300 15470 3320
rect 15430 3270 15470 3300
rect 15430 3250 15440 3270
rect 15460 3250 15470 3270
rect 15430 3220 15470 3250
rect 15430 3200 15440 3220
rect 15460 3200 15470 3220
rect 15430 3170 15470 3200
rect 15430 3150 15440 3170
rect 15460 3150 15470 3170
rect 15430 3120 15470 3150
rect 15430 3100 15440 3120
rect 15460 3100 15470 3120
rect 15430 3070 15470 3100
rect 15430 3050 15440 3070
rect 15460 3050 15470 3070
rect 15430 3020 15470 3050
rect 15430 3000 15440 3020
rect 15460 3000 15470 3020
rect 15430 2985 15470 3000
rect 15485 3570 15525 3585
rect 15485 3550 15495 3570
rect 15515 3550 15525 3570
rect 15485 3520 15525 3550
rect 15485 3500 15495 3520
rect 15515 3500 15525 3520
rect 15485 3470 15525 3500
rect 15485 3450 15495 3470
rect 15515 3450 15525 3470
rect 15485 3420 15525 3450
rect 15485 3400 15495 3420
rect 15515 3400 15525 3420
rect 15485 3370 15525 3400
rect 15485 3350 15495 3370
rect 15515 3350 15525 3370
rect 15485 3320 15525 3350
rect 15485 3300 15495 3320
rect 15515 3300 15525 3320
rect 15485 3270 15525 3300
rect 15485 3250 15495 3270
rect 15515 3250 15525 3270
rect 15485 3220 15525 3250
rect 15485 3200 15495 3220
rect 15515 3200 15525 3220
rect 15485 3170 15525 3200
rect 15485 3150 15495 3170
rect 15515 3150 15525 3170
rect 15485 3120 15525 3150
rect 15485 3100 15495 3120
rect 15515 3100 15525 3120
rect 15485 3070 15525 3100
rect 15485 3050 15495 3070
rect 15515 3050 15525 3070
rect 15485 3020 15525 3050
rect 15485 3000 15495 3020
rect 15515 3000 15525 3020
rect 15485 2985 15525 3000
rect 15540 3570 15580 3585
rect 15540 3550 15550 3570
rect 15570 3550 15580 3570
rect 15540 3520 15580 3550
rect 15540 3500 15550 3520
rect 15570 3500 15580 3520
rect 15540 3470 15580 3500
rect 15540 3450 15550 3470
rect 15570 3450 15580 3470
rect 15540 3420 15580 3450
rect 15540 3400 15550 3420
rect 15570 3400 15580 3420
rect 15540 3370 15580 3400
rect 15540 3350 15550 3370
rect 15570 3350 15580 3370
rect 15540 3320 15580 3350
rect 15540 3300 15550 3320
rect 15570 3300 15580 3320
rect 15540 3270 15580 3300
rect 15540 3250 15550 3270
rect 15570 3250 15580 3270
rect 15540 3220 15580 3250
rect 15540 3200 15550 3220
rect 15570 3200 15580 3220
rect 15540 3170 15580 3200
rect 15540 3150 15550 3170
rect 15570 3150 15580 3170
rect 15540 3120 15580 3150
rect 15540 3100 15550 3120
rect 15570 3100 15580 3120
rect 15540 3070 15580 3100
rect 15540 3050 15550 3070
rect 15570 3050 15580 3070
rect 15540 3020 15580 3050
rect 15540 3000 15550 3020
rect 15570 3000 15580 3020
rect 15540 2985 15580 3000
rect 15595 3570 15635 3585
rect 15595 3550 15605 3570
rect 15625 3550 15635 3570
rect 15595 3520 15635 3550
rect 15595 3500 15605 3520
rect 15625 3500 15635 3520
rect 15595 3470 15635 3500
rect 15595 3450 15605 3470
rect 15625 3450 15635 3470
rect 15595 3420 15635 3450
rect 15595 3400 15605 3420
rect 15625 3400 15635 3420
rect 15595 3370 15635 3400
rect 15595 3350 15605 3370
rect 15625 3350 15635 3370
rect 15595 3320 15635 3350
rect 15595 3300 15605 3320
rect 15625 3300 15635 3320
rect 15595 3270 15635 3300
rect 15595 3250 15605 3270
rect 15625 3250 15635 3270
rect 15595 3220 15635 3250
rect 15595 3200 15605 3220
rect 15625 3200 15635 3220
rect 15595 3170 15635 3200
rect 15595 3150 15605 3170
rect 15625 3150 15635 3170
rect 15595 3120 15635 3150
rect 15595 3100 15605 3120
rect 15625 3100 15635 3120
rect 15595 3070 15635 3100
rect 15595 3050 15605 3070
rect 15625 3050 15635 3070
rect 15595 3020 15635 3050
rect 15595 3000 15605 3020
rect 15625 3000 15635 3020
rect 15595 2985 15635 3000
rect 15650 3570 15690 3585
rect 15650 3550 15660 3570
rect 15680 3550 15690 3570
rect 15650 3520 15690 3550
rect 15650 3500 15660 3520
rect 15680 3500 15690 3520
rect 15650 3470 15690 3500
rect 15650 3450 15660 3470
rect 15680 3450 15690 3470
rect 15650 3420 15690 3450
rect 15650 3400 15660 3420
rect 15680 3400 15690 3420
rect 15650 3370 15690 3400
rect 15650 3350 15660 3370
rect 15680 3350 15690 3370
rect 15650 3320 15690 3350
rect 15650 3300 15660 3320
rect 15680 3300 15690 3320
rect 15650 3270 15690 3300
rect 15650 3250 15660 3270
rect 15680 3250 15690 3270
rect 15650 3220 15690 3250
rect 15650 3200 15660 3220
rect 15680 3200 15690 3220
rect 15650 3170 15690 3200
rect 15650 3150 15660 3170
rect 15680 3150 15690 3170
rect 15650 3120 15690 3150
rect 15650 3100 15660 3120
rect 15680 3100 15690 3120
rect 15650 3070 15690 3100
rect 15650 3050 15660 3070
rect 15680 3050 15690 3070
rect 15650 3020 15690 3050
rect 15650 3000 15660 3020
rect 15680 3000 15690 3020
rect 15650 2985 15690 3000
rect 15705 3570 15745 3585
rect 15705 3550 15715 3570
rect 15735 3550 15745 3570
rect 15705 3520 15745 3550
rect 15705 3500 15715 3520
rect 15735 3500 15745 3520
rect 15705 3470 15745 3500
rect 15705 3450 15715 3470
rect 15735 3450 15745 3470
rect 15705 3420 15745 3450
rect 15705 3400 15715 3420
rect 15735 3400 15745 3420
rect 15705 3370 15745 3400
rect 15705 3350 15715 3370
rect 15735 3350 15745 3370
rect 15705 3320 15745 3350
rect 15705 3300 15715 3320
rect 15735 3300 15745 3320
rect 15705 3270 15745 3300
rect 15705 3250 15715 3270
rect 15735 3250 15745 3270
rect 15705 3220 15745 3250
rect 15705 3200 15715 3220
rect 15735 3200 15745 3220
rect 15705 3170 15745 3200
rect 15705 3150 15715 3170
rect 15735 3150 15745 3170
rect 15705 3120 15745 3150
rect 15705 3100 15715 3120
rect 15735 3100 15745 3120
rect 15705 3070 15745 3100
rect 15705 3050 15715 3070
rect 15735 3050 15745 3070
rect 15705 3020 15745 3050
rect 15705 3000 15715 3020
rect 15735 3000 15745 3020
rect 15705 2985 15745 3000
rect 15760 3570 15800 3585
rect 15760 3550 15770 3570
rect 15790 3550 15800 3570
rect 15760 3520 15800 3550
rect 15760 3500 15770 3520
rect 15790 3500 15800 3520
rect 15760 3470 15800 3500
rect 15760 3450 15770 3470
rect 15790 3450 15800 3470
rect 15760 3420 15800 3450
rect 15760 3400 15770 3420
rect 15790 3400 15800 3420
rect 15760 3370 15800 3400
rect 15760 3350 15770 3370
rect 15790 3350 15800 3370
rect 15760 3320 15800 3350
rect 15760 3300 15770 3320
rect 15790 3300 15800 3320
rect 15760 3270 15800 3300
rect 15760 3250 15770 3270
rect 15790 3250 15800 3270
rect 15760 3220 15800 3250
rect 15760 3200 15770 3220
rect 15790 3200 15800 3220
rect 15760 3170 15800 3200
rect 15760 3150 15770 3170
rect 15790 3150 15800 3170
rect 15760 3120 15800 3150
rect 15760 3100 15770 3120
rect 15790 3100 15800 3120
rect 15760 3070 15800 3100
rect 15760 3050 15770 3070
rect 15790 3050 15800 3070
rect 15760 3020 15800 3050
rect 15760 3000 15770 3020
rect 15790 3000 15800 3020
rect 15760 2985 15800 3000
rect 15815 3570 15855 3585
rect 15815 3550 15825 3570
rect 15845 3550 15855 3570
rect 15815 3520 15855 3550
rect 15815 3500 15825 3520
rect 15845 3500 15855 3520
rect 15815 3470 15855 3500
rect 15815 3450 15825 3470
rect 15845 3450 15855 3470
rect 15815 3420 15855 3450
rect 15815 3400 15825 3420
rect 15845 3400 15855 3420
rect 15815 3370 15855 3400
rect 15815 3350 15825 3370
rect 15845 3350 15855 3370
rect 15815 3320 15855 3350
rect 15815 3300 15825 3320
rect 15845 3300 15855 3320
rect 15815 3270 15855 3300
rect 15815 3250 15825 3270
rect 15845 3250 15855 3270
rect 15815 3220 15855 3250
rect 15815 3200 15825 3220
rect 15845 3200 15855 3220
rect 15815 3170 15855 3200
rect 16220 3560 16260 3575
rect 16220 3540 16230 3560
rect 16250 3540 16260 3560
rect 16220 3510 16260 3540
rect 16220 3490 16230 3510
rect 16250 3490 16260 3510
rect 16220 3460 16260 3490
rect 16220 3440 16230 3460
rect 16250 3440 16260 3460
rect 16220 3410 16260 3440
rect 16220 3390 16230 3410
rect 16250 3390 16260 3410
rect 16220 3360 16260 3390
rect 16220 3340 16230 3360
rect 16250 3340 16260 3360
rect 16220 3310 16260 3340
rect 16220 3290 16230 3310
rect 16250 3290 16260 3310
rect 16220 3260 16260 3290
rect 16220 3240 16230 3260
rect 16250 3240 16260 3260
rect 16220 3210 16260 3240
rect 16220 3190 16230 3210
rect 16250 3190 16260 3210
rect 16220 3175 16260 3190
rect 16280 3560 16320 3575
rect 16280 3540 16290 3560
rect 16310 3540 16320 3560
rect 16280 3510 16320 3540
rect 16280 3490 16290 3510
rect 16310 3490 16320 3510
rect 16280 3460 16320 3490
rect 16280 3440 16290 3460
rect 16310 3440 16320 3460
rect 16280 3410 16320 3440
rect 16280 3390 16290 3410
rect 16310 3390 16320 3410
rect 16280 3360 16320 3390
rect 16280 3340 16290 3360
rect 16310 3340 16320 3360
rect 16280 3310 16320 3340
rect 16280 3290 16290 3310
rect 16310 3290 16320 3310
rect 16280 3260 16320 3290
rect 16280 3240 16290 3260
rect 16310 3240 16320 3260
rect 16280 3210 16320 3240
rect 16280 3190 16290 3210
rect 16310 3190 16320 3210
rect 16280 3175 16320 3190
rect 16340 3560 16380 3575
rect 16340 3540 16350 3560
rect 16370 3540 16380 3560
rect 16340 3510 16380 3540
rect 16340 3490 16350 3510
rect 16370 3490 16380 3510
rect 16340 3460 16380 3490
rect 16340 3440 16350 3460
rect 16370 3440 16380 3460
rect 16340 3410 16380 3440
rect 16340 3390 16350 3410
rect 16370 3390 16380 3410
rect 16340 3360 16380 3390
rect 16340 3340 16350 3360
rect 16370 3340 16380 3360
rect 16340 3310 16380 3340
rect 16340 3290 16350 3310
rect 16370 3290 16380 3310
rect 16340 3260 16380 3290
rect 16340 3240 16350 3260
rect 16370 3240 16380 3260
rect 16340 3210 16380 3240
rect 16340 3190 16350 3210
rect 16370 3190 16380 3210
rect 16340 3175 16380 3190
rect 16400 3560 16440 3575
rect 16400 3540 16410 3560
rect 16430 3540 16440 3560
rect 16400 3510 16440 3540
rect 16400 3490 16410 3510
rect 16430 3490 16440 3510
rect 16400 3460 16440 3490
rect 16400 3440 16410 3460
rect 16430 3440 16440 3460
rect 16400 3410 16440 3440
rect 16400 3390 16410 3410
rect 16430 3390 16440 3410
rect 16400 3360 16440 3390
rect 16400 3340 16410 3360
rect 16430 3340 16440 3360
rect 16400 3310 16440 3340
rect 16400 3290 16410 3310
rect 16430 3290 16440 3310
rect 16400 3260 16440 3290
rect 16400 3240 16410 3260
rect 16430 3240 16440 3260
rect 16400 3210 16440 3240
rect 16400 3190 16410 3210
rect 16430 3190 16440 3210
rect 16400 3175 16440 3190
rect 16460 3560 16500 3575
rect 16460 3540 16470 3560
rect 16490 3540 16500 3560
rect 16460 3510 16500 3540
rect 16460 3490 16470 3510
rect 16490 3490 16500 3510
rect 16460 3460 16500 3490
rect 16460 3440 16470 3460
rect 16490 3440 16500 3460
rect 16460 3410 16500 3440
rect 16460 3390 16470 3410
rect 16490 3390 16500 3410
rect 16460 3360 16500 3390
rect 16460 3340 16470 3360
rect 16490 3340 16500 3360
rect 16460 3310 16500 3340
rect 16460 3290 16470 3310
rect 16490 3290 16500 3310
rect 16460 3260 16500 3290
rect 16460 3240 16470 3260
rect 16490 3240 16500 3260
rect 16460 3210 16500 3240
rect 16460 3190 16470 3210
rect 16490 3190 16500 3210
rect 16460 3175 16500 3190
rect 16520 3560 16560 3575
rect 16520 3540 16530 3560
rect 16550 3540 16560 3560
rect 16520 3510 16560 3540
rect 16520 3490 16530 3510
rect 16550 3490 16560 3510
rect 16520 3460 16560 3490
rect 16520 3440 16530 3460
rect 16550 3440 16560 3460
rect 16520 3410 16560 3440
rect 16520 3390 16530 3410
rect 16550 3390 16560 3410
rect 16520 3360 16560 3390
rect 16520 3340 16530 3360
rect 16550 3340 16560 3360
rect 16520 3310 16560 3340
rect 16520 3290 16530 3310
rect 16550 3290 16560 3310
rect 16520 3260 16560 3290
rect 16520 3240 16530 3260
rect 16550 3240 16560 3260
rect 16520 3210 16560 3240
rect 16520 3190 16530 3210
rect 16550 3190 16560 3210
rect 16520 3175 16560 3190
rect 16580 3560 16620 3575
rect 16580 3540 16590 3560
rect 16610 3540 16620 3560
rect 16580 3510 16620 3540
rect 16580 3490 16590 3510
rect 16610 3490 16620 3510
rect 16580 3460 16620 3490
rect 16580 3440 16590 3460
rect 16610 3440 16620 3460
rect 16580 3410 16620 3440
rect 16580 3390 16590 3410
rect 16610 3390 16620 3410
rect 16580 3360 16620 3390
rect 16580 3340 16590 3360
rect 16610 3340 16620 3360
rect 16580 3310 16620 3340
rect 16580 3290 16590 3310
rect 16610 3290 16620 3310
rect 16580 3260 16620 3290
rect 16580 3240 16590 3260
rect 16610 3240 16620 3260
rect 16580 3210 16620 3240
rect 16580 3190 16590 3210
rect 16610 3190 16620 3210
rect 16580 3175 16620 3190
rect 16640 3560 16680 3575
rect 16640 3540 16650 3560
rect 16670 3540 16680 3560
rect 16640 3510 16680 3540
rect 16640 3490 16650 3510
rect 16670 3490 16680 3510
rect 16640 3460 16680 3490
rect 16640 3440 16650 3460
rect 16670 3440 16680 3460
rect 16640 3410 16680 3440
rect 16640 3390 16650 3410
rect 16670 3390 16680 3410
rect 16640 3360 16680 3390
rect 16640 3340 16650 3360
rect 16670 3340 16680 3360
rect 16640 3310 16680 3340
rect 16640 3290 16650 3310
rect 16670 3290 16680 3310
rect 16640 3260 16680 3290
rect 16640 3240 16650 3260
rect 16670 3240 16680 3260
rect 16640 3210 16680 3240
rect 16640 3190 16650 3210
rect 16670 3190 16680 3210
rect 16640 3175 16680 3190
rect 16700 3560 16740 3575
rect 16700 3540 16710 3560
rect 16730 3540 16740 3560
rect 16700 3510 16740 3540
rect 16700 3490 16710 3510
rect 16730 3490 16740 3510
rect 16700 3460 16740 3490
rect 16700 3440 16710 3460
rect 16730 3440 16740 3460
rect 16700 3410 16740 3440
rect 16700 3390 16710 3410
rect 16730 3390 16740 3410
rect 16700 3360 16740 3390
rect 16700 3340 16710 3360
rect 16730 3340 16740 3360
rect 16700 3310 16740 3340
rect 16700 3290 16710 3310
rect 16730 3290 16740 3310
rect 16700 3260 16740 3290
rect 16700 3240 16710 3260
rect 16730 3240 16740 3260
rect 16700 3210 16740 3240
rect 16700 3190 16710 3210
rect 16730 3190 16740 3210
rect 16700 3175 16740 3190
rect 16760 3560 16800 3575
rect 16760 3540 16770 3560
rect 16790 3540 16800 3560
rect 16760 3510 16800 3540
rect 16760 3490 16770 3510
rect 16790 3490 16800 3510
rect 16760 3460 16800 3490
rect 16760 3440 16770 3460
rect 16790 3440 16800 3460
rect 16760 3410 16800 3440
rect 16760 3390 16770 3410
rect 16790 3390 16800 3410
rect 16760 3360 16800 3390
rect 16760 3340 16770 3360
rect 16790 3340 16800 3360
rect 16760 3310 16800 3340
rect 16760 3290 16770 3310
rect 16790 3290 16800 3310
rect 16760 3260 16800 3290
rect 16760 3240 16770 3260
rect 16790 3240 16800 3260
rect 16760 3210 16800 3240
rect 16760 3190 16770 3210
rect 16790 3190 16800 3210
rect 16760 3175 16800 3190
rect 16820 3560 16860 3575
rect 16820 3540 16830 3560
rect 16850 3540 16860 3560
rect 16820 3510 16860 3540
rect 16820 3490 16830 3510
rect 16850 3490 16860 3510
rect 16820 3460 16860 3490
rect 16820 3440 16830 3460
rect 16850 3440 16860 3460
rect 16820 3410 16860 3440
rect 16820 3390 16830 3410
rect 16850 3390 16860 3410
rect 16820 3360 16860 3390
rect 16820 3340 16830 3360
rect 16850 3340 16860 3360
rect 16820 3310 16860 3340
rect 16820 3290 16830 3310
rect 16850 3290 16860 3310
rect 16820 3260 16860 3290
rect 16820 3240 16830 3260
rect 16850 3240 16860 3260
rect 16820 3210 16860 3240
rect 16820 3190 16830 3210
rect 16850 3190 16860 3210
rect 16820 3175 16860 3190
rect 16880 3560 16920 3575
rect 16880 3540 16890 3560
rect 16910 3540 16920 3560
rect 16880 3510 16920 3540
rect 16880 3490 16890 3510
rect 16910 3490 16920 3510
rect 16880 3460 16920 3490
rect 16880 3440 16890 3460
rect 16910 3440 16920 3460
rect 16880 3410 16920 3440
rect 16880 3390 16890 3410
rect 16910 3390 16920 3410
rect 16880 3360 16920 3390
rect 16880 3340 16890 3360
rect 16910 3340 16920 3360
rect 16880 3310 16920 3340
rect 16880 3290 16890 3310
rect 16910 3290 16920 3310
rect 16880 3260 16920 3290
rect 16880 3240 16890 3260
rect 16910 3240 16920 3260
rect 16880 3210 16920 3240
rect 16880 3190 16890 3210
rect 16910 3190 16920 3210
rect 16880 3175 16920 3190
rect 16940 3560 16980 3575
rect 16940 3540 16950 3560
rect 16970 3540 16980 3560
rect 16940 3510 16980 3540
rect 16940 3490 16950 3510
rect 16970 3490 16980 3510
rect 16940 3460 16980 3490
rect 16940 3440 16950 3460
rect 16970 3440 16980 3460
rect 16940 3410 16980 3440
rect 16940 3390 16950 3410
rect 16970 3390 16980 3410
rect 16940 3360 16980 3390
rect 16940 3340 16950 3360
rect 16970 3340 16980 3360
rect 16940 3310 16980 3340
rect 16940 3290 16950 3310
rect 16970 3290 16980 3310
rect 16940 3260 16980 3290
rect 16940 3240 16950 3260
rect 16970 3240 16980 3260
rect 16940 3210 16980 3240
rect 16940 3190 16950 3210
rect 16970 3190 16980 3210
rect 16940 3175 16980 3190
rect 17000 3560 17040 3575
rect 17000 3540 17010 3560
rect 17030 3540 17040 3560
rect 17000 3510 17040 3540
rect 17000 3490 17010 3510
rect 17030 3490 17040 3510
rect 17000 3460 17040 3490
rect 17000 3440 17010 3460
rect 17030 3440 17040 3460
rect 17000 3410 17040 3440
rect 17000 3390 17010 3410
rect 17030 3390 17040 3410
rect 17000 3360 17040 3390
rect 17000 3340 17010 3360
rect 17030 3340 17040 3360
rect 17000 3310 17040 3340
rect 17000 3290 17010 3310
rect 17030 3290 17040 3310
rect 17000 3260 17040 3290
rect 17000 3240 17010 3260
rect 17030 3240 17040 3260
rect 17000 3210 17040 3240
rect 17000 3190 17010 3210
rect 17030 3190 17040 3210
rect 17000 3175 17040 3190
rect 17060 3560 17100 3575
rect 17060 3540 17070 3560
rect 17090 3540 17100 3560
rect 17060 3510 17100 3540
rect 17060 3490 17070 3510
rect 17090 3490 17100 3510
rect 17060 3460 17100 3490
rect 17060 3440 17070 3460
rect 17090 3440 17100 3460
rect 17060 3410 17100 3440
rect 17060 3390 17070 3410
rect 17090 3390 17100 3410
rect 17060 3360 17100 3390
rect 17060 3340 17070 3360
rect 17090 3340 17100 3360
rect 17060 3310 17100 3340
rect 17060 3290 17070 3310
rect 17090 3290 17100 3310
rect 17060 3260 17100 3290
rect 17060 3240 17070 3260
rect 17090 3240 17100 3260
rect 17060 3210 17100 3240
rect 17060 3190 17070 3210
rect 17090 3190 17100 3210
rect 17060 3175 17100 3190
rect 17120 3560 17160 3575
rect 17120 3540 17130 3560
rect 17150 3540 17160 3560
rect 17120 3510 17160 3540
rect 17120 3490 17130 3510
rect 17150 3490 17160 3510
rect 17120 3460 17160 3490
rect 17120 3440 17130 3460
rect 17150 3440 17160 3460
rect 17120 3410 17160 3440
rect 17120 3390 17130 3410
rect 17150 3390 17160 3410
rect 17120 3360 17160 3390
rect 17120 3340 17130 3360
rect 17150 3340 17160 3360
rect 17120 3310 17160 3340
rect 17120 3290 17130 3310
rect 17150 3290 17160 3310
rect 17120 3260 17160 3290
rect 17120 3240 17130 3260
rect 17150 3240 17160 3260
rect 17120 3210 17160 3240
rect 17120 3190 17130 3210
rect 17150 3190 17160 3210
rect 17120 3175 17160 3190
rect 17180 3560 17220 3575
rect 17180 3540 17190 3560
rect 17210 3540 17220 3560
rect 17180 3510 17220 3540
rect 17180 3490 17190 3510
rect 17210 3490 17220 3510
rect 17180 3460 17220 3490
rect 17180 3440 17190 3460
rect 17210 3440 17220 3460
rect 17180 3410 17220 3440
rect 17180 3390 17190 3410
rect 17210 3390 17220 3410
rect 17180 3360 17220 3390
rect 17180 3340 17190 3360
rect 17210 3340 17220 3360
rect 17180 3310 17220 3340
rect 17180 3290 17190 3310
rect 17210 3290 17220 3310
rect 17180 3260 17220 3290
rect 17180 3240 17190 3260
rect 17210 3240 17220 3260
rect 17180 3210 17220 3240
rect 17180 3190 17190 3210
rect 17210 3190 17220 3210
rect 17180 3175 17220 3190
rect 17240 3560 17280 3575
rect 17240 3540 17250 3560
rect 17270 3540 17280 3560
rect 17240 3510 17280 3540
rect 17240 3490 17250 3510
rect 17270 3490 17280 3510
rect 17240 3460 17280 3490
rect 17240 3440 17250 3460
rect 17270 3440 17280 3460
rect 17240 3410 17280 3440
rect 17240 3390 17250 3410
rect 17270 3390 17280 3410
rect 17240 3360 17280 3390
rect 17240 3340 17250 3360
rect 17270 3340 17280 3360
rect 17240 3310 17280 3340
rect 17240 3290 17250 3310
rect 17270 3290 17280 3310
rect 17240 3260 17280 3290
rect 17240 3240 17250 3260
rect 17270 3240 17280 3260
rect 17240 3210 17280 3240
rect 17240 3190 17250 3210
rect 17270 3190 17280 3210
rect 17240 3175 17280 3190
rect 17300 3560 17340 3575
rect 17300 3540 17310 3560
rect 17330 3540 17340 3560
rect 17300 3510 17340 3540
rect 17300 3490 17310 3510
rect 17330 3490 17340 3510
rect 17300 3460 17340 3490
rect 17300 3440 17310 3460
rect 17330 3440 17340 3460
rect 17300 3410 17340 3440
rect 17300 3390 17310 3410
rect 17330 3390 17340 3410
rect 17300 3360 17340 3390
rect 17300 3340 17310 3360
rect 17330 3340 17340 3360
rect 17300 3310 17340 3340
rect 17300 3290 17310 3310
rect 17330 3290 17340 3310
rect 17300 3260 17340 3290
rect 17300 3240 17310 3260
rect 17330 3240 17340 3260
rect 17300 3210 17340 3240
rect 17300 3190 17310 3210
rect 17330 3190 17340 3210
rect 17300 3175 17340 3190
rect 17360 3560 17400 3575
rect 17360 3540 17370 3560
rect 17390 3540 17400 3560
rect 17360 3510 17400 3540
rect 17360 3490 17370 3510
rect 17390 3490 17400 3510
rect 17360 3460 17400 3490
rect 17360 3440 17370 3460
rect 17390 3440 17400 3460
rect 17360 3410 17400 3440
rect 17360 3390 17370 3410
rect 17390 3390 17400 3410
rect 17360 3360 17400 3390
rect 17360 3340 17370 3360
rect 17390 3340 17400 3360
rect 17360 3310 17400 3340
rect 17360 3290 17370 3310
rect 17390 3290 17400 3310
rect 17360 3260 17400 3290
rect 17360 3240 17370 3260
rect 17390 3240 17400 3260
rect 17360 3210 17400 3240
rect 17360 3190 17370 3210
rect 17390 3190 17400 3210
rect 17360 3175 17400 3190
rect 17420 3560 17460 3575
rect 17420 3540 17430 3560
rect 17450 3540 17460 3560
rect 17420 3510 17460 3540
rect 17420 3490 17430 3510
rect 17450 3490 17460 3510
rect 17420 3460 17460 3490
rect 17420 3440 17430 3460
rect 17450 3440 17460 3460
rect 17420 3410 17460 3440
rect 17420 3390 17430 3410
rect 17450 3390 17460 3410
rect 17420 3360 17460 3390
rect 17420 3340 17430 3360
rect 17450 3340 17460 3360
rect 17420 3310 17460 3340
rect 17420 3290 17430 3310
rect 17450 3290 17460 3310
rect 17420 3260 17460 3290
rect 17420 3240 17430 3260
rect 17450 3240 17460 3260
rect 17420 3210 17460 3240
rect 17420 3190 17430 3210
rect 17450 3190 17460 3210
rect 17420 3175 17460 3190
rect 17480 3560 17520 3575
rect 17480 3540 17490 3560
rect 17510 3540 17520 3560
rect 17480 3510 17520 3540
rect 17480 3490 17490 3510
rect 17510 3490 17520 3510
rect 17480 3460 17520 3490
rect 17480 3440 17490 3460
rect 17510 3440 17520 3460
rect 17480 3410 17520 3440
rect 17480 3390 17490 3410
rect 17510 3390 17520 3410
rect 17480 3360 17520 3390
rect 17480 3340 17490 3360
rect 17510 3340 17520 3360
rect 17480 3310 17520 3340
rect 17480 3290 17490 3310
rect 17510 3290 17520 3310
rect 17480 3260 17520 3290
rect 17480 3240 17490 3260
rect 17510 3240 17520 3260
rect 17480 3210 17520 3240
rect 17480 3190 17490 3210
rect 17510 3190 17520 3210
rect 17480 3175 17520 3190
rect 17540 3560 17580 3575
rect 17540 3540 17550 3560
rect 17570 3540 17580 3560
rect 17540 3510 17580 3540
rect 17540 3490 17550 3510
rect 17570 3490 17580 3510
rect 17540 3460 17580 3490
rect 17540 3440 17550 3460
rect 17570 3440 17580 3460
rect 17540 3410 17580 3440
rect 17540 3390 17550 3410
rect 17570 3390 17580 3410
rect 17540 3360 17580 3390
rect 17540 3340 17550 3360
rect 17570 3340 17580 3360
rect 17540 3310 17580 3340
rect 17540 3290 17550 3310
rect 17570 3290 17580 3310
rect 17540 3260 17580 3290
rect 17540 3240 17550 3260
rect 17570 3240 17580 3260
rect 17540 3210 17580 3240
rect 17540 3190 17550 3210
rect 17570 3190 17580 3210
rect 17540 3175 17580 3190
rect 17945 3570 17985 3585
rect 17945 3550 17955 3570
rect 17975 3550 17985 3570
rect 17945 3520 17985 3550
rect 17945 3500 17955 3520
rect 17975 3500 17985 3520
rect 17945 3470 17985 3500
rect 17945 3450 17955 3470
rect 17975 3450 17985 3470
rect 17945 3420 17985 3450
rect 17945 3400 17955 3420
rect 17975 3400 17985 3420
rect 17945 3370 17985 3400
rect 17945 3350 17955 3370
rect 17975 3350 17985 3370
rect 17945 3320 17985 3350
rect 17945 3300 17955 3320
rect 17975 3300 17985 3320
rect 17945 3270 17985 3300
rect 17945 3250 17955 3270
rect 17975 3250 17985 3270
rect 17945 3220 17985 3250
rect 17945 3200 17955 3220
rect 17975 3200 17985 3220
rect 15815 3150 15825 3170
rect 15845 3150 15855 3170
rect 17945 3170 17985 3200
rect 17945 3150 17955 3170
rect 17975 3150 17985 3170
rect 15815 3120 15855 3150
rect 17945 3120 17985 3150
rect 15815 3100 15825 3120
rect 15845 3100 15855 3120
rect 15815 3070 15855 3100
rect 15815 3050 15825 3070
rect 15845 3050 15855 3070
rect 15815 3020 15855 3050
rect 15815 3000 15825 3020
rect 15845 3000 15855 3020
rect 15815 2985 15855 3000
rect 17945 3100 17955 3120
rect 17975 3100 17985 3120
rect 17945 3070 17985 3100
rect 17945 3050 17955 3070
rect 17975 3050 17985 3070
rect 17945 3020 17985 3050
rect 17945 3000 17955 3020
rect 17975 3000 17985 3020
rect 17945 2985 17985 3000
rect 18000 3570 18040 3585
rect 18000 3550 18010 3570
rect 18030 3550 18040 3570
rect 18000 3520 18040 3550
rect 18000 3500 18010 3520
rect 18030 3500 18040 3520
rect 18000 3470 18040 3500
rect 18000 3450 18010 3470
rect 18030 3450 18040 3470
rect 18000 3420 18040 3450
rect 18000 3400 18010 3420
rect 18030 3400 18040 3420
rect 18000 3370 18040 3400
rect 18000 3350 18010 3370
rect 18030 3350 18040 3370
rect 18000 3320 18040 3350
rect 18000 3300 18010 3320
rect 18030 3300 18040 3320
rect 18000 3270 18040 3300
rect 18000 3250 18010 3270
rect 18030 3250 18040 3270
rect 18000 3220 18040 3250
rect 18000 3200 18010 3220
rect 18030 3200 18040 3220
rect 18000 3170 18040 3200
rect 18000 3150 18010 3170
rect 18030 3150 18040 3170
rect 18000 3120 18040 3150
rect 18000 3100 18010 3120
rect 18030 3100 18040 3120
rect 18000 3070 18040 3100
rect 18000 3050 18010 3070
rect 18030 3050 18040 3070
rect 18000 3020 18040 3050
rect 18000 3000 18010 3020
rect 18030 3000 18040 3020
rect 18000 2985 18040 3000
rect 18055 3570 18095 3585
rect 18055 3550 18065 3570
rect 18085 3550 18095 3570
rect 18055 3520 18095 3550
rect 18055 3500 18065 3520
rect 18085 3500 18095 3520
rect 18055 3470 18095 3500
rect 18055 3450 18065 3470
rect 18085 3450 18095 3470
rect 18055 3420 18095 3450
rect 18055 3400 18065 3420
rect 18085 3400 18095 3420
rect 18055 3370 18095 3400
rect 18055 3350 18065 3370
rect 18085 3350 18095 3370
rect 18055 3320 18095 3350
rect 18055 3300 18065 3320
rect 18085 3300 18095 3320
rect 18055 3270 18095 3300
rect 18055 3250 18065 3270
rect 18085 3250 18095 3270
rect 18055 3220 18095 3250
rect 18055 3200 18065 3220
rect 18085 3200 18095 3220
rect 18055 3170 18095 3200
rect 18055 3150 18065 3170
rect 18085 3150 18095 3170
rect 18055 3120 18095 3150
rect 18055 3100 18065 3120
rect 18085 3100 18095 3120
rect 18055 3070 18095 3100
rect 18055 3050 18065 3070
rect 18085 3050 18095 3070
rect 18055 3020 18095 3050
rect 18055 3000 18065 3020
rect 18085 3000 18095 3020
rect 18055 2985 18095 3000
rect 18110 3570 18150 3585
rect 18110 3550 18120 3570
rect 18140 3550 18150 3570
rect 18110 3520 18150 3550
rect 18110 3500 18120 3520
rect 18140 3500 18150 3520
rect 18110 3470 18150 3500
rect 18110 3450 18120 3470
rect 18140 3450 18150 3470
rect 18110 3420 18150 3450
rect 18110 3400 18120 3420
rect 18140 3400 18150 3420
rect 18110 3370 18150 3400
rect 18110 3350 18120 3370
rect 18140 3350 18150 3370
rect 18110 3320 18150 3350
rect 18110 3300 18120 3320
rect 18140 3300 18150 3320
rect 18110 3270 18150 3300
rect 18110 3250 18120 3270
rect 18140 3250 18150 3270
rect 18110 3220 18150 3250
rect 18110 3200 18120 3220
rect 18140 3200 18150 3220
rect 18110 3170 18150 3200
rect 18110 3150 18120 3170
rect 18140 3150 18150 3170
rect 18110 3120 18150 3150
rect 18110 3100 18120 3120
rect 18140 3100 18150 3120
rect 18110 3070 18150 3100
rect 18110 3050 18120 3070
rect 18140 3050 18150 3070
rect 18110 3020 18150 3050
rect 18110 3000 18120 3020
rect 18140 3000 18150 3020
rect 18110 2985 18150 3000
rect 18165 3570 18205 3585
rect 18165 3550 18175 3570
rect 18195 3550 18205 3570
rect 18165 3520 18205 3550
rect 18165 3500 18175 3520
rect 18195 3500 18205 3520
rect 18165 3470 18205 3500
rect 18165 3450 18175 3470
rect 18195 3450 18205 3470
rect 18165 3420 18205 3450
rect 18165 3400 18175 3420
rect 18195 3400 18205 3420
rect 18165 3370 18205 3400
rect 18165 3350 18175 3370
rect 18195 3350 18205 3370
rect 18165 3320 18205 3350
rect 18165 3300 18175 3320
rect 18195 3300 18205 3320
rect 18165 3270 18205 3300
rect 18165 3250 18175 3270
rect 18195 3250 18205 3270
rect 18165 3220 18205 3250
rect 18165 3200 18175 3220
rect 18195 3200 18205 3220
rect 18165 3170 18205 3200
rect 18165 3150 18175 3170
rect 18195 3150 18205 3170
rect 18165 3120 18205 3150
rect 18165 3100 18175 3120
rect 18195 3100 18205 3120
rect 18165 3070 18205 3100
rect 18165 3050 18175 3070
rect 18195 3050 18205 3070
rect 18165 3020 18205 3050
rect 18165 3000 18175 3020
rect 18195 3000 18205 3020
rect 18165 2985 18205 3000
rect 18220 3570 18260 3585
rect 18220 3550 18230 3570
rect 18250 3550 18260 3570
rect 18220 3520 18260 3550
rect 18220 3500 18230 3520
rect 18250 3500 18260 3520
rect 18220 3470 18260 3500
rect 18220 3450 18230 3470
rect 18250 3450 18260 3470
rect 18220 3420 18260 3450
rect 18220 3400 18230 3420
rect 18250 3400 18260 3420
rect 18220 3370 18260 3400
rect 18220 3350 18230 3370
rect 18250 3350 18260 3370
rect 18220 3320 18260 3350
rect 18220 3300 18230 3320
rect 18250 3300 18260 3320
rect 18220 3270 18260 3300
rect 18220 3250 18230 3270
rect 18250 3250 18260 3270
rect 18220 3220 18260 3250
rect 18220 3200 18230 3220
rect 18250 3200 18260 3220
rect 18220 3170 18260 3200
rect 18220 3150 18230 3170
rect 18250 3150 18260 3170
rect 18220 3120 18260 3150
rect 18220 3100 18230 3120
rect 18250 3100 18260 3120
rect 18220 3070 18260 3100
rect 18220 3050 18230 3070
rect 18250 3050 18260 3070
rect 18220 3020 18260 3050
rect 18220 3000 18230 3020
rect 18250 3000 18260 3020
rect 18220 2985 18260 3000
rect 18275 3570 18315 3585
rect 18275 3550 18285 3570
rect 18305 3550 18315 3570
rect 18275 3520 18315 3550
rect 18275 3500 18285 3520
rect 18305 3500 18315 3520
rect 18275 3470 18315 3500
rect 18275 3450 18285 3470
rect 18305 3450 18315 3470
rect 18275 3420 18315 3450
rect 18275 3400 18285 3420
rect 18305 3400 18315 3420
rect 18275 3370 18315 3400
rect 18275 3350 18285 3370
rect 18305 3350 18315 3370
rect 18275 3320 18315 3350
rect 18275 3300 18285 3320
rect 18305 3300 18315 3320
rect 18275 3270 18315 3300
rect 18275 3250 18285 3270
rect 18305 3250 18315 3270
rect 18275 3220 18315 3250
rect 18275 3200 18285 3220
rect 18305 3200 18315 3220
rect 18275 3170 18315 3200
rect 18275 3150 18285 3170
rect 18305 3150 18315 3170
rect 18275 3120 18315 3150
rect 18275 3100 18285 3120
rect 18305 3100 18315 3120
rect 18275 3070 18315 3100
rect 18275 3050 18285 3070
rect 18305 3050 18315 3070
rect 18275 3020 18315 3050
rect 18275 3000 18285 3020
rect 18305 3000 18315 3020
rect 18275 2985 18315 3000
rect 18330 3570 18370 3585
rect 18330 3550 18340 3570
rect 18360 3550 18370 3570
rect 18330 3520 18370 3550
rect 18330 3500 18340 3520
rect 18360 3500 18370 3520
rect 18330 3470 18370 3500
rect 18330 3450 18340 3470
rect 18360 3450 18370 3470
rect 18330 3420 18370 3450
rect 18330 3400 18340 3420
rect 18360 3400 18370 3420
rect 18330 3370 18370 3400
rect 18330 3350 18340 3370
rect 18360 3350 18370 3370
rect 18330 3320 18370 3350
rect 18330 3300 18340 3320
rect 18360 3300 18370 3320
rect 18330 3270 18370 3300
rect 18330 3250 18340 3270
rect 18360 3250 18370 3270
rect 18330 3220 18370 3250
rect 18330 3200 18340 3220
rect 18360 3200 18370 3220
rect 18330 3170 18370 3200
rect 18330 3150 18340 3170
rect 18360 3150 18370 3170
rect 18330 3120 18370 3150
rect 18330 3100 18340 3120
rect 18360 3100 18370 3120
rect 18330 3070 18370 3100
rect 18330 3050 18340 3070
rect 18360 3050 18370 3070
rect 18330 3020 18370 3050
rect 18330 3000 18340 3020
rect 18360 3000 18370 3020
rect 18330 2985 18370 3000
rect 18385 3570 18425 3585
rect 18385 3550 18395 3570
rect 18415 3550 18425 3570
rect 18385 3520 18425 3550
rect 18385 3500 18395 3520
rect 18415 3500 18425 3520
rect 18385 3470 18425 3500
rect 18385 3450 18395 3470
rect 18415 3450 18425 3470
rect 18385 3420 18425 3450
rect 18385 3400 18395 3420
rect 18415 3400 18425 3420
rect 18385 3370 18425 3400
rect 18385 3350 18395 3370
rect 18415 3350 18425 3370
rect 18385 3320 18425 3350
rect 18385 3300 18395 3320
rect 18415 3300 18425 3320
rect 18385 3270 18425 3300
rect 18385 3250 18395 3270
rect 18415 3250 18425 3270
rect 18385 3220 18425 3250
rect 18385 3200 18395 3220
rect 18415 3200 18425 3220
rect 18385 3170 18425 3200
rect 18385 3150 18395 3170
rect 18415 3150 18425 3170
rect 18385 3120 18425 3150
rect 18385 3100 18395 3120
rect 18415 3100 18425 3120
rect 18385 3070 18425 3100
rect 18385 3050 18395 3070
rect 18415 3050 18425 3070
rect 18385 3020 18425 3050
rect 18385 3000 18395 3020
rect 18415 3000 18425 3020
rect 18385 2985 18425 3000
rect 18440 3570 18480 3585
rect 18440 3550 18450 3570
rect 18470 3550 18480 3570
rect 18440 3520 18480 3550
rect 18440 3500 18450 3520
rect 18470 3500 18480 3520
rect 18440 3470 18480 3500
rect 18440 3450 18450 3470
rect 18470 3450 18480 3470
rect 18440 3420 18480 3450
rect 18440 3400 18450 3420
rect 18470 3400 18480 3420
rect 18440 3370 18480 3400
rect 18440 3350 18450 3370
rect 18470 3350 18480 3370
rect 18440 3320 18480 3350
rect 18440 3300 18450 3320
rect 18470 3300 18480 3320
rect 18440 3270 18480 3300
rect 18440 3250 18450 3270
rect 18470 3250 18480 3270
rect 18440 3220 18480 3250
rect 18440 3200 18450 3220
rect 18470 3200 18480 3220
rect 18440 3170 18480 3200
rect 18440 3150 18450 3170
rect 18470 3150 18480 3170
rect 18440 3120 18480 3150
rect 18440 3100 18450 3120
rect 18470 3100 18480 3120
rect 18440 3070 18480 3100
rect 18440 3050 18450 3070
rect 18470 3050 18480 3070
rect 18440 3020 18480 3050
rect 18440 3000 18450 3020
rect 18470 3000 18480 3020
rect 18440 2985 18480 3000
rect 18495 3570 18535 3585
rect 18495 3550 18505 3570
rect 18525 3550 18535 3570
rect 18495 3520 18535 3550
rect 18495 3500 18505 3520
rect 18525 3500 18535 3520
rect 18495 3470 18535 3500
rect 18495 3450 18505 3470
rect 18525 3450 18535 3470
rect 18495 3420 18535 3450
rect 18495 3400 18505 3420
rect 18525 3400 18535 3420
rect 18495 3370 18535 3400
rect 18495 3350 18505 3370
rect 18525 3350 18535 3370
rect 18495 3320 18535 3350
rect 18495 3300 18505 3320
rect 18525 3300 18535 3320
rect 18495 3270 18535 3300
rect 18495 3250 18505 3270
rect 18525 3250 18535 3270
rect 18495 3220 18535 3250
rect 18495 3200 18505 3220
rect 18525 3200 18535 3220
rect 18495 3170 18535 3200
rect 18495 3150 18505 3170
rect 18525 3150 18535 3170
rect 18495 3120 18535 3150
rect 18495 3100 18505 3120
rect 18525 3100 18535 3120
rect 18495 3070 18535 3100
rect 18495 3050 18505 3070
rect 18525 3050 18535 3070
rect 18495 3020 18535 3050
rect 18495 3000 18505 3020
rect 18525 3000 18535 3020
rect 18495 2985 18535 3000
rect 18550 3570 18590 3585
rect 18550 3550 18560 3570
rect 18580 3550 18590 3570
rect 18550 3520 18590 3550
rect 18550 3500 18560 3520
rect 18580 3500 18590 3520
rect 18550 3470 18590 3500
rect 18550 3450 18560 3470
rect 18580 3450 18590 3470
rect 18550 3420 18590 3450
rect 18550 3400 18560 3420
rect 18580 3400 18590 3420
rect 18550 3370 18590 3400
rect 18550 3350 18560 3370
rect 18580 3350 18590 3370
rect 18550 3320 18590 3350
rect 18550 3300 18560 3320
rect 18580 3300 18590 3320
rect 18550 3270 18590 3300
rect 18550 3250 18560 3270
rect 18580 3250 18590 3270
rect 18550 3220 18590 3250
rect 18550 3200 18560 3220
rect 18580 3200 18590 3220
rect 18550 3170 18590 3200
rect 18550 3150 18560 3170
rect 18580 3150 18590 3170
rect 18550 3120 18590 3150
rect 18550 3100 18560 3120
rect 18580 3100 18590 3120
rect 18550 3070 18590 3100
rect 18550 3050 18560 3070
rect 18580 3050 18590 3070
rect 18550 3020 18590 3050
rect 18550 3000 18560 3020
rect 18580 3000 18590 3020
rect 18550 2985 18590 3000
rect 18605 3570 18645 3585
rect 18605 3550 18615 3570
rect 18635 3550 18645 3570
rect 18605 3520 18645 3550
rect 18605 3500 18615 3520
rect 18635 3500 18645 3520
rect 18605 3470 18645 3500
rect 18605 3450 18615 3470
rect 18635 3450 18645 3470
rect 18605 3420 18645 3450
rect 18605 3400 18615 3420
rect 18635 3400 18645 3420
rect 18605 3370 18645 3400
rect 18605 3350 18615 3370
rect 18635 3350 18645 3370
rect 18605 3320 18645 3350
rect 18605 3300 18615 3320
rect 18635 3300 18645 3320
rect 18605 3270 18645 3300
rect 18605 3250 18615 3270
rect 18635 3250 18645 3270
rect 18605 3220 18645 3250
rect 18605 3200 18615 3220
rect 18635 3200 18645 3220
rect 18605 3170 18645 3200
rect 18605 3150 18615 3170
rect 18635 3150 18645 3170
rect 18605 3120 18645 3150
rect 18605 3100 18615 3120
rect 18635 3100 18645 3120
rect 18605 3070 18645 3100
rect 18605 3050 18615 3070
rect 18635 3050 18645 3070
rect 18605 3020 18645 3050
rect 18605 3000 18615 3020
rect 18635 3000 18645 3020
rect 18605 2985 18645 3000
rect 16220 2880 16260 2895
rect 16220 2860 16230 2880
rect 16250 2860 16260 2880
rect 16220 2830 16260 2860
rect 16220 2810 16230 2830
rect 16250 2810 16260 2830
rect 16220 2780 16260 2810
rect 16220 2760 16230 2780
rect 16250 2760 16260 2780
rect 16220 2730 16260 2760
rect 16220 2710 16230 2730
rect 16250 2710 16260 2730
rect 16220 2680 16260 2710
rect 16220 2660 16230 2680
rect 16250 2660 16260 2680
rect 15155 2640 15195 2655
rect 15155 2620 15165 2640
rect 15185 2620 15195 2640
rect 15155 2590 15195 2620
rect 15155 2570 15165 2590
rect 15185 2570 15195 2590
rect 15155 2540 15195 2570
rect 15155 2520 15165 2540
rect 15185 2520 15195 2540
rect 15155 2490 15195 2520
rect 15155 2470 15165 2490
rect 15185 2470 15195 2490
rect 15155 2455 15195 2470
rect 15210 2640 15250 2655
rect 15210 2620 15220 2640
rect 15240 2620 15250 2640
rect 15210 2590 15250 2620
rect 15210 2570 15220 2590
rect 15240 2570 15250 2590
rect 15210 2540 15250 2570
rect 15210 2520 15220 2540
rect 15240 2520 15250 2540
rect 15210 2490 15250 2520
rect 15210 2470 15220 2490
rect 15240 2470 15250 2490
rect 15210 2455 15250 2470
rect 15265 2640 15305 2655
rect 15265 2620 15275 2640
rect 15295 2620 15305 2640
rect 15265 2590 15305 2620
rect 15265 2570 15275 2590
rect 15295 2570 15305 2590
rect 15265 2540 15305 2570
rect 15265 2520 15275 2540
rect 15295 2520 15305 2540
rect 15265 2490 15305 2520
rect 15265 2470 15275 2490
rect 15295 2470 15305 2490
rect 15265 2455 15305 2470
rect 15320 2640 15360 2655
rect 15320 2620 15330 2640
rect 15350 2620 15360 2640
rect 15320 2590 15360 2620
rect 15320 2570 15330 2590
rect 15350 2570 15360 2590
rect 15320 2540 15360 2570
rect 15320 2520 15330 2540
rect 15350 2520 15360 2540
rect 15320 2490 15360 2520
rect 15320 2470 15330 2490
rect 15350 2470 15360 2490
rect 15320 2455 15360 2470
rect 15375 2640 15415 2655
rect 15375 2620 15385 2640
rect 15405 2620 15415 2640
rect 15375 2590 15415 2620
rect 15375 2570 15385 2590
rect 15405 2570 15415 2590
rect 15375 2540 15415 2570
rect 15375 2520 15385 2540
rect 15405 2520 15415 2540
rect 15375 2490 15415 2520
rect 15375 2470 15385 2490
rect 15405 2470 15415 2490
rect 15375 2455 15415 2470
rect 15430 2640 15470 2655
rect 15430 2620 15440 2640
rect 15460 2620 15470 2640
rect 15430 2590 15470 2620
rect 15430 2570 15440 2590
rect 15460 2570 15470 2590
rect 15430 2540 15470 2570
rect 15430 2520 15440 2540
rect 15460 2520 15470 2540
rect 15430 2490 15470 2520
rect 15430 2470 15440 2490
rect 15460 2470 15470 2490
rect 15430 2455 15470 2470
rect 15485 2640 15525 2655
rect 15485 2620 15495 2640
rect 15515 2620 15525 2640
rect 15485 2590 15525 2620
rect 15485 2570 15495 2590
rect 15515 2570 15525 2590
rect 15485 2540 15525 2570
rect 15485 2520 15495 2540
rect 15515 2520 15525 2540
rect 15485 2490 15525 2520
rect 15485 2470 15495 2490
rect 15515 2470 15525 2490
rect 15485 2455 15525 2470
rect 15540 2640 15580 2655
rect 15540 2620 15550 2640
rect 15570 2620 15580 2640
rect 15540 2590 15580 2620
rect 15540 2570 15550 2590
rect 15570 2570 15580 2590
rect 15540 2540 15580 2570
rect 15540 2520 15550 2540
rect 15570 2520 15580 2540
rect 15540 2490 15580 2520
rect 15540 2470 15550 2490
rect 15570 2470 15580 2490
rect 15540 2455 15580 2470
rect 15595 2640 15635 2655
rect 15595 2620 15605 2640
rect 15625 2620 15635 2640
rect 15595 2590 15635 2620
rect 15595 2570 15605 2590
rect 15625 2570 15635 2590
rect 15595 2540 15635 2570
rect 15595 2520 15605 2540
rect 15625 2520 15635 2540
rect 15595 2490 15635 2520
rect 15595 2470 15605 2490
rect 15625 2470 15635 2490
rect 15595 2455 15635 2470
rect 15650 2640 15690 2655
rect 15650 2620 15660 2640
rect 15680 2620 15690 2640
rect 15650 2590 15690 2620
rect 15650 2570 15660 2590
rect 15680 2570 15690 2590
rect 15650 2540 15690 2570
rect 15650 2520 15660 2540
rect 15680 2520 15690 2540
rect 15650 2490 15690 2520
rect 15650 2470 15660 2490
rect 15680 2470 15690 2490
rect 15650 2455 15690 2470
rect 15705 2640 15745 2655
rect 15705 2620 15715 2640
rect 15735 2620 15745 2640
rect 15705 2590 15745 2620
rect 15705 2570 15715 2590
rect 15735 2570 15745 2590
rect 15705 2540 15745 2570
rect 15705 2520 15715 2540
rect 15735 2520 15745 2540
rect 15705 2490 15745 2520
rect 15705 2470 15715 2490
rect 15735 2470 15745 2490
rect 15705 2455 15745 2470
rect 15760 2640 15800 2655
rect 15760 2620 15770 2640
rect 15790 2620 15800 2640
rect 15760 2590 15800 2620
rect 15760 2570 15770 2590
rect 15790 2570 15800 2590
rect 15760 2540 15800 2570
rect 15760 2520 15770 2540
rect 15790 2520 15800 2540
rect 15760 2490 15800 2520
rect 15760 2470 15770 2490
rect 15790 2470 15800 2490
rect 15760 2455 15800 2470
rect 15815 2640 15855 2655
rect 15815 2620 15825 2640
rect 15845 2620 15855 2640
rect 15815 2590 15855 2620
rect 15815 2570 15825 2590
rect 15845 2570 15855 2590
rect 15815 2540 15855 2570
rect 15815 2520 15825 2540
rect 15845 2520 15855 2540
rect 15815 2490 15855 2520
rect 16220 2630 16260 2660
rect 16220 2610 16230 2630
rect 16250 2610 16260 2630
rect 16220 2580 16260 2610
rect 16220 2560 16230 2580
rect 16250 2560 16260 2580
rect 16220 2530 16260 2560
rect 16220 2510 16230 2530
rect 16250 2510 16260 2530
rect 16220 2495 16260 2510
rect 16280 2880 16320 2895
rect 16280 2860 16290 2880
rect 16310 2860 16320 2880
rect 16280 2830 16320 2860
rect 16280 2810 16290 2830
rect 16310 2810 16320 2830
rect 16280 2780 16320 2810
rect 16280 2760 16290 2780
rect 16310 2760 16320 2780
rect 16280 2730 16320 2760
rect 16280 2710 16290 2730
rect 16310 2710 16320 2730
rect 16280 2680 16320 2710
rect 16280 2660 16290 2680
rect 16310 2660 16320 2680
rect 16280 2630 16320 2660
rect 16280 2610 16290 2630
rect 16310 2610 16320 2630
rect 16280 2580 16320 2610
rect 16280 2560 16290 2580
rect 16310 2560 16320 2580
rect 16280 2530 16320 2560
rect 16280 2510 16290 2530
rect 16310 2510 16320 2530
rect 16280 2495 16320 2510
rect 16340 2880 16380 2895
rect 16340 2860 16350 2880
rect 16370 2860 16380 2880
rect 16340 2830 16380 2860
rect 16340 2810 16350 2830
rect 16370 2810 16380 2830
rect 16340 2780 16380 2810
rect 16340 2760 16350 2780
rect 16370 2760 16380 2780
rect 16340 2730 16380 2760
rect 16340 2710 16350 2730
rect 16370 2710 16380 2730
rect 16340 2680 16380 2710
rect 16340 2660 16350 2680
rect 16370 2660 16380 2680
rect 16340 2630 16380 2660
rect 16340 2610 16350 2630
rect 16370 2610 16380 2630
rect 16340 2580 16380 2610
rect 16340 2560 16350 2580
rect 16370 2560 16380 2580
rect 16340 2530 16380 2560
rect 16340 2510 16350 2530
rect 16370 2510 16380 2530
rect 16340 2495 16380 2510
rect 16400 2880 16440 2895
rect 16400 2860 16410 2880
rect 16430 2860 16440 2880
rect 16400 2830 16440 2860
rect 16400 2810 16410 2830
rect 16430 2810 16440 2830
rect 16400 2780 16440 2810
rect 16400 2760 16410 2780
rect 16430 2760 16440 2780
rect 16400 2730 16440 2760
rect 16400 2710 16410 2730
rect 16430 2710 16440 2730
rect 16400 2680 16440 2710
rect 16400 2660 16410 2680
rect 16430 2660 16440 2680
rect 16400 2630 16440 2660
rect 16400 2610 16410 2630
rect 16430 2610 16440 2630
rect 16400 2580 16440 2610
rect 16400 2560 16410 2580
rect 16430 2560 16440 2580
rect 16400 2530 16440 2560
rect 16400 2510 16410 2530
rect 16430 2510 16440 2530
rect 16400 2495 16440 2510
rect 16460 2880 16500 2895
rect 16460 2860 16470 2880
rect 16490 2860 16500 2880
rect 16460 2830 16500 2860
rect 16460 2810 16470 2830
rect 16490 2810 16500 2830
rect 16460 2780 16500 2810
rect 16460 2760 16470 2780
rect 16490 2760 16500 2780
rect 16460 2730 16500 2760
rect 16460 2710 16470 2730
rect 16490 2710 16500 2730
rect 16460 2680 16500 2710
rect 16460 2660 16470 2680
rect 16490 2660 16500 2680
rect 16460 2630 16500 2660
rect 16460 2610 16470 2630
rect 16490 2610 16500 2630
rect 16460 2580 16500 2610
rect 16460 2560 16470 2580
rect 16490 2560 16500 2580
rect 16460 2530 16500 2560
rect 16460 2510 16470 2530
rect 16490 2510 16500 2530
rect 16460 2495 16500 2510
rect 16520 2880 16560 2895
rect 16520 2860 16530 2880
rect 16550 2860 16560 2880
rect 16520 2830 16560 2860
rect 16520 2810 16530 2830
rect 16550 2810 16560 2830
rect 16520 2780 16560 2810
rect 16520 2760 16530 2780
rect 16550 2760 16560 2780
rect 16520 2730 16560 2760
rect 16520 2710 16530 2730
rect 16550 2710 16560 2730
rect 16520 2680 16560 2710
rect 16520 2660 16530 2680
rect 16550 2660 16560 2680
rect 16520 2630 16560 2660
rect 16520 2610 16530 2630
rect 16550 2610 16560 2630
rect 16520 2580 16560 2610
rect 16520 2560 16530 2580
rect 16550 2560 16560 2580
rect 16520 2530 16560 2560
rect 16520 2510 16530 2530
rect 16550 2510 16560 2530
rect 16520 2495 16560 2510
rect 16580 2880 16620 2895
rect 16580 2860 16590 2880
rect 16610 2860 16620 2880
rect 16580 2830 16620 2860
rect 16580 2810 16590 2830
rect 16610 2810 16620 2830
rect 16580 2780 16620 2810
rect 16580 2760 16590 2780
rect 16610 2760 16620 2780
rect 16580 2730 16620 2760
rect 16580 2710 16590 2730
rect 16610 2710 16620 2730
rect 16580 2680 16620 2710
rect 16580 2660 16590 2680
rect 16610 2660 16620 2680
rect 16580 2630 16620 2660
rect 16580 2610 16590 2630
rect 16610 2610 16620 2630
rect 16580 2580 16620 2610
rect 16580 2560 16590 2580
rect 16610 2560 16620 2580
rect 16580 2530 16620 2560
rect 16580 2510 16590 2530
rect 16610 2510 16620 2530
rect 16580 2495 16620 2510
rect 16640 2880 16680 2895
rect 16640 2860 16650 2880
rect 16670 2860 16680 2880
rect 16640 2830 16680 2860
rect 16640 2810 16650 2830
rect 16670 2810 16680 2830
rect 16640 2780 16680 2810
rect 16640 2760 16650 2780
rect 16670 2760 16680 2780
rect 16640 2730 16680 2760
rect 16640 2710 16650 2730
rect 16670 2710 16680 2730
rect 16640 2680 16680 2710
rect 16640 2660 16650 2680
rect 16670 2660 16680 2680
rect 16640 2630 16680 2660
rect 16640 2610 16650 2630
rect 16670 2610 16680 2630
rect 16640 2580 16680 2610
rect 16640 2560 16650 2580
rect 16670 2560 16680 2580
rect 16640 2530 16680 2560
rect 16640 2510 16650 2530
rect 16670 2510 16680 2530
rect 16640 2495 16680 2510
rect 16700 2880 16740 2895
rect 16700 2860 16710 2880
rect 16730 2860 16740 2880
rect 16700 2830 16740 2860
rect 16700 2810 16710 2830
rect 16730 2810 16740 2830
rect 16700 2780 16740 2810
rect 16700 2760 16710 2780
rect 16730 2760 16740 2780
rect 16700 2730 16740 2760
rect 16700 2710 16710 2730
rect 16730 2710 16740 2730
rect 16700 2680 16740 2710
rect 16700 2660 16710 2680
rect 16730 2660 16740 2680
rect 16700 2630 16740 2660
rect 16700 2610 16710 2630
rect 16730 2610 16740 2630
rect 16700 2580 16740 2610
rect 16700 2560 16710 2580
rect 16730 2560 16740 2580
rect 16700 2530 16740 2560
rect 16700 2510 16710 2530
rect 16730 2510 16740 2530
rect 16700 2495 16740 2510
rect 16760 2880 16800 2895
rect 16760 2860 16770 2880
rect 16790 2860 16800 2880
rect 16760 2830 16800 2860
rect 16760 2810 16770 2830
rect 16790 2810 16800 2830
rect 16760 2780 16800 2810
rect 16760 2760 16770 2780
rect 16790 2760 16800 2780
rect 16760 2730 16800 2760
rect 16760 2710 16770 2730
rect 16790 2710 16800 2730
rect 16760 2680 16800 2710
rect 16760 2660 16770 2680
rect 16790 2660 16800 2680
rect 16760 2630 16800 2660
rect 16760 2610 16770 2630
rect 16790 2610 16800 2630
rect 16760 2580 16800 2610
rect 16760 2560 16770 2580
rect 16790 2560 16800 2580
rect 16760 2530 16800 2560
rect 16760 2510 16770 2530
rect 16790 2510 16800 2530
rect 16760 2495 16800 2510
rect 16820 2880 16860 2895
rect 16820 2860 16830 2880
rect 16850 2860 16860 2880
rect 16820 2830 16860 2860
rect 16820 2810 16830 2830
rect 16850 2810 16860 2830
rect 16820 2780 16860 2810
rect 16820 2760 16830 2780
rect 16850 2760 16860 2780
rect 16820 2730 16860 2760
rect 16820 2710 16830 2730
rect 16850 2710 16860 2730
rect 16820 2680 16860 2710
rect 16820 2660 16830 2680
rect 16850 2660 16860 2680
rect 16820 2630 16860 2660
rect 16820 2610 16830 2630
rect 16850 2610 16860 2630
rect 16820 2580 16860 2610
rect 16820 2560 16830 2580
rect 16850 2560 16860 2580
rect 16820 2530 16860 2560
rect 16820 2510 16830 2530
rect 16850 2510 16860 2530
rect 16820 2495 16860 2510
rect 16880 2880 16920 2895
rect 16880 2860 16890 2880
rect 16910 2860 16920 2880
rect 16880 2830 16920 2860
rect 16880 2810 16890 2830
rect 16910 2810 16920 2830
rect 16880 2780 16920 2810
rect 16880 2760 16890 2780
rect 16910 2760 16920 2780
rect 16880 2730 16920 2760
rect 16880 2710 16890 2730
rect 16910 2710 16920 2730
rect 16880 2680 16920 2710
rect 16880 2660 16890 2680
rect 16910 2660 16920 2680
rect 16880 2630 16920 2660
rect 16880 2610 16890 2630
rect 16910 2610 16920 2630
rect 16880 2580 16920 2610
rect 16880 2560 16890 2580
rect 16910 2560 16920 2580
rect 16880 2530 16920 2560
rect 16880 2510 16890 2530
rect 16910 2510 16920 2530
rect 16880 2495 16920 2510
rect 16940 2880 16980 2895
rect 16940 2860 16950 2880
rect 16970 2860 16980 2880
rect 16940 2830 16980 2860
rect 16940 2810 16950 2830
rect 16970 2810 16980 2830
rect 16940 2780 16980 2810
rect 16940 2760 16950 2780
rect 16970 2760 16980 2780
rect 16940 2730 16980 2760
rect 16940 2710 16950 2730
rect 16970 2710 16980 2730
rect 16940 2680 16980 2710
rect 16940 2660 16950 2680
rect 16970 2660 16980 2680
rect 16940 2630 16980 2660
rect 16940 2610 16950 2630
rect 16970 2610 16980 2630
rect 16940 2580 16980 2610
rect 16940 2560 16950 2580
rect 16970 2560 16980 2580
rect 16940 2530 16980 2560
rect 16940 2510 16950 2530
rect 16970 2510 16980 2530
rect 16940 2495 16980 2510
rect 17000 2880 17040 2895
rect 17000 2860 17010 2880
rect 17030 2860 17040 2880
rect 17000 2830 17040 2860
rect 17000 2810 17010 2830
rect 17030 2810 17040 2830
rect 17000 2780 17040 2810
rect 17000 2760 17010 2780
rect 17030 2760 17040 2780
rect 17000 2730 17040 2760
rect 17000 2710 17010 2730
rect 17030 2710 17040 2730
rect 17000 2680 17040 2710
rect 17000 2660 17010 2680
rect 17030 2660 17040 2680
rect 17000 2630 17040 2660
rect 17000 2610 17010 2630
rect 17030 2610 17040 2630
rect 17000 2580 17040 2610
rect 17000 2560 17010 2580
rect 17030 2560 17040 2580
rect 17000 2530 17040 2560
rect 17000 2510 17010 2530
rect 17030 2510 17040 2530
rect 17000 2495 17040 2510
rect 17060 2880 17100 2895
rect 17060 2860 17070 2880
rect 17090 2860 17100 2880
rect 17060 2830 17100 2860
rect 17060 2810 17070 2830
rect 17090 2810 17100 2830
rect 17060 2780 17100 2810
rect 17060 2760 17070 2780
rect 17090 2760 17100 2780
rect 17060 2730 17100 2760
rect 17060 2710 17070 2730
rect 17090 2710 17100 2730
rect 17060 2680 17100 2710
rect 17060 2660 17070 2680
rect 17090 2660 17100 2680
rect 17060 2630 17100 2660
rect 17060 2610 17070 2630
rect 17090 2610 17100 2630
rect 17060 2580 17100 2610
rect 17060 2560 17070 2580
rect 17090 2560 17100 2580
rect 17060 2530 17100 2560
rect 17060 2510 17070 2530
rect 17090 2510 17100 2530
rect 17060 2495 17100 2510
rect 17120 2880 17160 2895
rect 17120 2860 17130 2880
rect 17150 2860 17160 2880
rect 17120 2830 17160 2860
rect 17120 2810 17130 2830
rect 17150 2810 17160 2830
rect 17120 2780 17160 2810
rect 17120 2760 17130 2780
rect 17150 2760 17160 2780
rect 17120 2730 17160 2760
rect 17120 2710 17130 2730
rect 17150 2710 17160 2730
rect 17120 2680 17160 2710
rect 17120 2660 17130 2680
rect 17150 2660 17160 2680
rect 17120 2630 17160 2660
rect 17120 2610 17130 2630
rect 17150 2610 17160 2630
rect 17120 2580 17160 2610
rect 17120 2560 17130 2580
rect 17150 2560 17160 2580
rect 17120 2530 17160 2560
rect 17120 2510 17130 2530
rect 17150 2510 17160 2530
rect 17120 2495 17160 2510
rect 17180 2880 17220 2895
rect 17180 2860 17190 2880
rect 17210 2860 17220 2880
rect 17180 2830 17220 2860
rect 17180 2810 17190 2830
rect 17210 2810 17220 2830
rect 17180 2780 17220 2810
rect 17180 2760 17190 2780
rect 17210 2760 17220 2780
rect 17180 2730 17220 2760
rect 17180 2710 17190 2730
rect 17210 2710 17220 2730
rect 17180 2680 17220 2710
rect 17180 2660 17190 2680
rect 17210 2660 17220 2680
rect 17180 2630 17220 2660
rect 17180 2610 17190 2630
rect 17210 2610 17220 2630
rect 17180 2580 17220 2610
rect 17180 2560 17190 2580
rect 17210 2560 17220 2580
rect 17180 2530 17220 2560
rect 17180 2510 17190 2530
rect 17210 2510 17220 2530
rect 17180 2495 17220 2510
rect 17240 2880 17280 2895
rect 17240 2860 17250 2880
rect 17270 2860 17280 2880
rect 17240 2830 17280 2860
rect 17240 2810 17250 2830
rect 17270 2810 17280 2830
rect 17240 2780 17280 2810
rect 17240 2760 17250 2780
rect 17270 2760 17280 2780
rect 17240 2730 17280 2760
rect 17240 2710 17250 2730
rect 17270 2710 17280 2730
rect 17240 2680 17280 2710
rect 17240 2660 17250 2680
rect 17270 2660 17280 2680
rect 17240 2630 17280 2660
rect 17240 2610 17250 2630
rect 17270 2610 17280 2630
rect 17240 2580 17280 2610
rect 17240 2560 17250 2580
rect 17270 2560 17280 2580
rect 17240 2530 17280 2560
rect 17240 2510 17250 2530
rect 17270 2510 17280 2530
rect 17240 2495 17280 2510
rect 17300 2880 17340 2895
rect 17300 2860 17310 2880
rect 17330 2860 17340 2880
rect 17300 2830 17340 2860
rect 17300 2810 17310 2830
rect 17330 2810 17340 2830
rect 17300 2780 17340 2810
rect 17300 2760 17310 2780
rect 17330 2760 17340 2780
rect 17300 2730 17340 2760
rect 17300 2710 17310 2730
rect 17330 2710 17340 2730
rect 17300 2680 17340 2710
rect 17300 2660 17310 2680
rect 17330 2660 17340 2680
rect 17300 2630 17340 2660
rect 17300 2610 17310 2630
rect 17330 2610 17340 2630
rect 17300 2580 17340 2610
rect 17300 2560 17310 2580
rect 17330 2560 17340 2580
rect 17300 2530 17340 2560
rect 17300 2510 17310 2530
rect 17330 2510 17340 2530
rect 17300 2495 17340 2510
rect 17360 2880 17400 2895
rect 17360 2860 17370 2880
rect 17390 2860 17400 2880
rect 17360 2830 17400 2860
rect 17360 2810 17370 2830
rect 17390 2810 17400 2830
rect 17360 2780 17400 2810
rect 17360 2760 17370 2780
rect 17390 2760 17400 2780
rect 17360 2730 17400 2760
rect 17360 2710 17370 2730
rect 17390 2710 17400 2730
rect 17360 2680 17400 2710
rect 17360 2660 17370 2680
rect 17390 2660 17400 2680
rect 17360 2630 17400 2660
rect 17360 2610 17370 2630
rect 17390 2610 17400 2630
rect 17360 2580 17400 2610
rect 17360 2560 17370 2580
rect 17390 2560 17400 2580
rect 17360 2530 17400 2560
rect 17360 2510 17370 2530
rect 17390 2510 17400 2530
rect 17360 2495 17400 2510
rect 17420 2880 17460 2895
rect 17420 2860 17430 2880
rect 17450 2860 17460 2880
rect 17420 2830 17460 2860
rect 17420 2810 17430 2830
rect 17450 2810 17460 2830
rect 17420 2780 17460 2810
rect 17420 2760 17430 2780
rect 17450 2760 17460 2780
rect 17420 2730 17460 2760
rect 17420 2710 17430 2730
rect 17450 2710 17460 2730
rect 17420 2680 17460 2710
rect 17420 2660 17430 2680
rect 17450 2660 17460 2680
rect 17420 2630 17460 2660
rect 17420 2610 17430 2630
rect 17450 2610 17460 2630
rect 17420 2580 17460 2610
rect 17420 2560 17430 2580
rect 17450 2560 17460 2580
rect 17420 2530 17460 2560
rect 17420 2510 17430 2530
rect 17450 2510 17460 2530
rect 17420 2495 17460 2510
rect 17480 2880 17520 2895
rect 17480 2860 17490 2880
rect 17510 2860 17520 2880
rect 17480 2830 17520 2860
rect 17480 2810 17490 2830
rect 17510 2810 17520 2830
rect 17480 2780 17520 2810
rect 17480 2760 17490 2780
rect 17510 2760 17520 2780
rect 17480 2730 17520 2760
rect 17480 2710 17490 2730
rect 17510 2710 17520 2730
rect 17480 2680 17520 2710
rect 17480 2660 17490 2680
rect 17510 2660 17520 2680
rect 17480 2630 17520 2660
rect 17480 2610 17490 2630
rect 17510 2610 17520 2630
rect 17480 2580 17520 2610
rect 17480 2560 17490 2580
rect 17510 2560 17520 2580
rect 17480 2530 17520 2560
rect 17480 2510 17490 2530
rect 17510 2510 17520 2530
rect 17480 2495 17520 2510
rect 17540 2880 17580 2895
rect 17540 2860 17550 2880
rect 17570 2860 17580 2880
rect 17540 2830 17580 2860
rect 17540 2810 17550 2830
rect 17570 2810 17580 2830
rect 17540 2780 17580 2810
rect 17540 2760 17550 2780
rect 17570 2760 17580 2780
rect 17540 2730 17580 2760
rect 17540 2710 17550 2730
rect 17570 2710 17580 2730
rect 17540 2680 17580 2710
rect 17540 2660 17550 2680
rect 17570 2660 17580 2680
rect 17540 2630 17580 2660
rect 17540 2610 17550 2630
rect 17570 2610 17580 2630
rect 17540 2580 17580 2610
rect 17540 2560 17550 2580
rect 17570 2560 17580 2580
rect 17540 2530 17580 2560
rect 17540 2510 17550 2530
rect 17570 2510 17580 2530
rect 17540 2495 17580 2510
rect 17945 2640 17985 2655
rect 17945 2620 17955 2640
rect 17975 2620 17985 2640
rect 17945 2590 17985 2620
rect 17945 2570 17955 2590
rect 17975 2570 17985 2590
rect 17945 2540 17985 2570
rect 17945 2520 17955 2540
rect 17975 2520 17985 2540
rect 15815 2470 15825 2490
rect 15845 2470 15855 2490
rect 17945 2490 17985 2520
rect 17945 2470 17955 2490
rect 17975 2470 17985 2490
rect 15815 2455 15855 2470
rect 17945 2455 17985 2470
rect 18000 2640 18040 2655
rect 18000 2620 18010 2640
rect 18030 2620 18040 2640
rect 18000 2590 18040 2620
rect 18000 2570 18010 2590
rect 18030 2570 18040 2590
rect 18000 2540 18040 2570
rect 18000 2520 18010 2540
rect 18030 2520 18040 2540
rect 18000 2490 18040 2520
rect 18000 2470 18010 2490
rect 18030 2470 18040 2490
rect 18000 2455 18040 2470
rect 18055 2640 18095 2655
rect 18055 2620 18065 2640
rect 18085 2620 18095 2640
rect 18055 2590 18095 2620
rect 18055 2570 18065 2590
rect 18085 2570 18095 2590
rect 18055 2540 18095 2570
rect 18055 2520 18065 2540
rect 18085 2520 18095 2540
rect 18055 2490 18095 2520
rect 18055 2470 18065 2490
rect 18085 2470 18095 2490
rect 18055 2455 18095 2470
rect 18110 2640 18150 2655
rect 18110 2620 18120 2640
rect 18140 2620 18150 2640
rect 18110 2590 18150 2620
rect 18110 2570 18120 2590
rect 18140 2570 18150 2590
rect 18110 2540 18150 2570
rect 18110 2520 18120 2540
rect 18140 2520 18150 2540
rect 18110 2490 18150 2520
rect 18110 2470 18120 2490
rect 18140 2470 18150 2490
rect 18110 2455 18150 2470
rect 18165 2640 18205 2655
rect 18165 2620 18175 2640
rect 18195 2620 18205 2640
rect 18165 2590 18205 2620
rect 18165 2570 18175 2590
rect 18195 2570 18205 2590
rect 18165 2540 18205 2570
rect 18165 2520 18175 2540
rect 18195 2520 18205 2540
rect 18165 2490 18205 2520
rect 18165 2470 18175 2490
rect 18195 2470 18205 2490
rect 18165 2455 18205 2470
rect 18220 2640 18260 2655
rect 18220 2620 18230 2640
rect 18250 2620 18260 2640
rect 18220 2590 18260 2620
rect 18220 2570 18230 2590
rect 18250 2570 18260 2590
rect 18220 2540 18260 2570
rect 18220 2520 18230 2540
rect 18250 2520 18260 2540
rect 18220 2490 18260 2520
rect 18220 2470 18230 2490
rect 18250 2470 18260 2490
rect 18220 2455 18260 2470
rect 18275 2640 18315 2655
rect 18275 2620 18285 2640
rect 18305 2620 18315 2640
rect 18275 2590 18315 2620
rect 18275 2570 18285 2590
rect 18305 2570 18315 2590
rect 18275 2540 18315 2570
rect 18275 2520 18285 2540
rect 18305 2520 18315 2540
rect 18275 2490 18315 2520
rect 18275 2470 18285 2490
rect 18305 2470 18315 2490
rect 18275 2455 18315 2470
rect 18330 2640 18370 2655
rect 18330 2620 18340 2640
rect 18360 2620 18370 2640
rect 18330 2590 18370 2620
rect 18330 2570 18340 2590
rect 18360 2570 18370 2590
rect 18330 2540 18370 2570
rect 18330 2520 18340 2540
rect 18360 2520 18370 2540
rect 18330 2490 18370 2520
rect 18330 2470 18340 2490
rect 18360 2470 18370 2490
rect 18330 2455 18370 2470
rect 18385 2640 18425 2655
rect 18385 2620 18395 2640
rect 18415 2620 18425 2640
rect 18385 2590 18425 2620
rect 18385 2570 18395 2590
rect 18415 2570 18425 2590
rect 18385 2540 18425 2570
rect 18385 2520 18395 2540
rect 18415 2520 18425 2540
rect 18385 2490 18425 2520
rect 18385 2470 18395 2490
rect 18415 2470 18425 2490
rect 18385 2455 18425 2470
rect 18440 2640 18480 2655
rect 18440 2620 18450 2640
rect 18470 2620 18480 2640
rect 18440 2590 18480 2620
rect 18440 2570 18450 2590
rect 18470 2570 18480 2590
rect 18440 2540 18480 2570
rect 18440 2520 18450 2540
rect 18470 2520 18480 2540
rect 18440 2490 18480 2520
rect 18440 2470 18450 2490
rect 18470 2470 18480 2490
rect 18440 2455 18480 2470
rect 18495 2640 18535 2655
rect 18495 2620 18505 2640
rect 18525 2620 18535 2640
rect 18495 2590 18535 2620
rect 18495 2570 18505 2590
rect 18525 2570 18535 2590
rect 18495 2540 18535 2570
rect 18495 2520 18505 2540
rect 18525 2520 18535 2540
rect 18495 2490 18535 2520
rect 18495 2470 18505 2490
rect 18525 2470 18535 2490
rect 18495 2455 18535 2470
rect 18550 2640 18590 2655
rect 18550 2620 18560 2640
rect 18580 2620 18590 2640
rect 18550 2590 18590 2620
rect 18550 2570 18560 2590
rect 18580 2570 18590 2590
rect 18550 2540 18590 2570
rect 18550 2520 18560 2540
rect 18580 2520 18590 2540
rect 18550 2490 18590 2520
rect 18550 2470 18560 2490
rect 18580 2470 18590 2490
rect 18550 2455 18590 2470
rect 18605 2640 18645 2655
rect 18605 2620 18615 2640
rect 18635 2620 18645 2640
rect 18605 2590 18645 2620
rect 18605 2570 18615 2590
rect 18635 2570 18645 2590
rect 18605 2540 18645 2570
rect 18605 2520 18615 2540
rect 18635 2520 18645 2540
rect 18605 2490 18645 2520
rect 18605 2470 18615 2490
rect 18635 2470 18645 2490
rect 18605 2455 18645 2470
rect 15155 2250 15195 2265
rect 15155 2230 15165 2250
rect 15185 2230 15195 2250
rect 15155 2200 15195 2230
rect 15155 2180 15165 2200
rect 15185 2180 15195 2200
rect 15155 2150 15195 2180
rect 15155 2130 15165 2150
rect 15185 2130 15195 2150
rect 15155 2100 15195 2130
rect 15155 2080 15165 2100
rect 15185 2080 15195 2100
rect 15155 2050 15195 2080
rect 15155 2030 15165 2050
rect 15185 2030 15195 2050
rect 15155 2000 15195 2030
rect 15155 1980 15165 2000
rect 15185 1980 15195 2000
rect 15155 1965 15195 1980
rect 15210 2250 15250 2265
rect 15210 2230 15220 2250
rect 15240 2230 15250 2250
rect 15210 2200 15250 2230
rect 15210 2180 15220 2200
rect 15240 2180 15250 2200
rect 15210 2150 15250 2180
rect 15210 2130 15220 2150
rect 15240 2130 15250 2150
rect 15210 2100 15250 2130
rect 15210 2080 15220 2100
rect 15240 2080 15250 2100
rect 15210 2050 15250 2080
rect 15210 2030 15220 2050
rect 15240 2030 15250 2050
rect 15210 2000 15250 2030
rect 15210 1980 15220 2000
rect 15240 1980 15250 2000
rect 15210 1965 15250 1980
rect 15265 2250 15305 2265
rect 15265 2230 15275 2250
rect 15295 2230 15305 2250
rect 15265 2200 15305 2230
rect 15265 2180 15275 2200
rect 15295 2180 15305 2200
rect 15265 2150 15305 2180
rect 15265 2130 15275 2150
rect 15295 2130 15305 2150
rect 15265 2100 15305 2130
rect 15265 2080 15275 2100
rect 15295 2080 15305 2100
rect 15265 2050 15305 2080
rect 15265 2030 15275 2050
rect 15295 2030 15305 2050
rect 15265 2000 15305 2030
rect 15265 1980 15275 2000
rect 15295 1980 15305 2000
rect 15265 1965 15305 1980
rect 15320 2250 15360 2265
rect 15320 2230 15330 2250
rect 15350 2230 15360 2250
rect 15320 2200 15360 2230
rect 15320 2180 15330 2200
rect 15350 2180 15360 2200
rect 15320 2150 15360 2180
rect 15320 2130 15330 2150
rect 15350 2130 15360 2150
rect 15320 2100 15360 2130
rect 15320 2080 15330 2100
rect 15350 2080 15360 2100
rect 15320 2050 15360 2080
rect 15320 2030 15330 2050
rect 15350 2030 15360 2050
rect 15320 2000 15360 2030
rect 15320 1980 15330 2000
rect 15350 1980 15360 2000
rect 15320 1965 15360 1980
rect 15375 2250 15415 2265
rect 15375 2230 15385 2250
rect 15405 2230 15415 2250
rect 15375 2200 15415 2230
rect 15375 2180 15385 2200
rect 15405 2180 15415 2200
rect 15375 2150 15415 2180
rect 15375 2130 15385 2150
rect 15405 2130 15415 2150
rect 15375 2100 15415 2130
rect 15375 2080 15385 2100
rect 15405 2080 15415 2100
rect 15375 2050 15415 2080
rect 15375 2030 15385 2050
rect 15405 2030 15415 2050
rect 15375 2000 15415 2030
rect 15375 1980 15385 2000
rect 15405 1980 15415 2000
rect 15375 1965 15415 1980
rect 15430 2250 15470 2265
rect 15430 2230 15440 2250
rect 15460 2230 15470 2250
rect 15430 2200 15470 2230
rect 15430 2180 15440 2200
rect 15460 2180 15470 2200
rect 15430 2150 15470 2180
rect 15430 2130 15440 2150
rect 15460 2130 15470 2150
rect 15430 2100 15470 2130
rect 15430 2080 15440 2100
rect 15460 2080 15470 2100
rect 15430 2050 15470 2080
rect 15430 2030 15440 2050
rect 15460 2030 15470 2050
rect 15430 2000 15470 2030
rect 15430 1980 15440 2000
rect 15460 1980 15470 2000
rect 15430 1965 15470 1980
rect 15485 2250 15525 2265
rect 15485 2230 15495 2250
rect 15515 2230 15525 2250
rect 15485 2200 15525 2230
rect 15485 2180 15495 2200
rect 15515 2180 15525 2200
rect 15485 2150 15525 2180
rect 15485 2130 15495 2150
rect 15515 2130 15525 2150
rect 15485 2100 15525 2130
rect 15485 2080 15495 2100
rect 15515 2080 15525 2100
rect 15485 2050 15525 2080
rect 15485 2030 15495 2050
rect 15515 2030 15525 2050
rect 15485 2000 15525 2030
rect 15485 1980 15495 2000
rect 15515 1980 15525 2000
rect 15485 1965 15525 1980
rect 15540 2250 15580 2265
rect 15540 2230 15550 2250
rect 15570 2230 15580 2250
rect 15540 2200 15580 2230
rect 15540 2180 15550 2200
rect 15570 2180 15580 2200
rect 15540 2150 15580 2180
rect 15540 2130 15550 2150
rect 15570 2130 15580 2150
rect 15540 2100 15580 2130
rect 15540 2080 15550 2100
rect 15570 2080 15580 2100
rect 15540 2050 15580 2080
rect 15540 2030 15550 2050
rect 15570 2030 15580 2050
rect 15540 2000 15580 2030
rect 15540 1980 15550 2000
rect 15570 1980 15580 2000
rect 15540 1965 15580 1980
rect 15595 2250 15635 2265
rect 15595 2230 15605 2250
rect 15625 2230 15635 2250
rect 15595 2200 15635 2230
rect 15595 2180 15605 2200
rect 15625 2180 15635 2200
rect 15595 2150 15635 2180
rect 15595 2130 15605 2150
rect 15625 2130 15635 2150
rect 15595 2100 15635 2130
rect 15595 2080 15605 2100
rect 15625 2080 15635 2100
rect 15595 2050 15635 2080
rect 15595 2030 15605 2050
rect 15625 2030 15635 2050
rect 15595 2000 15635 2030
rect 15595 1980 15605 2000
rect 15625 1980 15635 2000
rect 15595 1965 15635 1980
rect 15650 2250 15690 2265
rect 15650 2230 15660 2250
rect 15680 2230 15690 2250
rect 15650 2200 15690 2230
rect 15650 2180 15660 2200
rect 15680 2180 15690 2200
rect 15650 2150 15690 2180
rect 15650 2130 15660 2150
rect 15680 2130 15690 2150
rect 15650 2100 15690 2130
rect 15650 2080 15660 2100
rect 15680 2080 15690 2100
rect 15650 2050 15690 2080
rect 15650 2030 15660 2050
rect 15680 2030 15690 2050
rect 15650 2000 15690 2030
rect 15650 1980 15660 2000
rect 15680 1980 15690 2000
rect 15650 1965 15690 1980
rect 15705 2250 15745 2265
rect 15705 2230 15715 2250
rect 15735 2230 15745 2250
rect 15705 2200 15745 2230
rect 15705 2180 15715 2200
rect 15735 2180 15745 2200
rect 15705 2150 15745 2180
rect 15705 2130 15715 2150
rect 15735 2130 15745 2150
rect 15705 2100 15745 2130
rect 15705 2080 15715 2100
rect 15735 2080 15745 2100
rect 15705 2050 15745 2080
rect 15705 2030 15715 2050
rect 15735 2030 15745 2050
rect 15705 2000 15745 2030
rect 15705 1980 15715 2000
rect 15735 1980 15745 2000
rect 15705 1965 15745 1980
rect 15760 2250 15800 2265
rect 15760 2230 15770 2250
rect 15790 2230 15800 2250
rect 15760 2200 15800 2230
rect 15760 2180 15770 2200
rect 15790 2180 15800 2200
rect 15760 2150 15800 2180
rect 15760 2130 15770 2150
rect 15790 2130 15800 2150
rect 15760 2100 15800 2130
rect 15760 2080 15770 2100
rect 15790 2080 15800 2100
rect 15760 2050 15800 2080
rect 15760 2030 15770 2050
rect 15790 2030 15800 2050
rect 15760 2000 15800 2030
rect 15760 1980 15770 2000
rect 15790 1980 15800 2000
rect 15760 1965 15800 1980
rect 15815 2250 15855 2265
rect 15815 2230 15825 2250
rect 15845 2230 15855 2250
rect 15815 2200 15855 2230
rect 15815 2180 15825 2200
rect 15845 2180 15855 2200
rect 17945 2250 17985 2265
rect 17945 2230 17955 2250
rect 17975 2230 17985 2250
rect 17945 2200 17985 2230
rect 15815 2150 15855 2180
rect 17945 2180 17955 2200
rect 17975 2180 17985 2200
rect 15815 2130 15825 2150
rect 15845 2130 15855 2150
rect 17945 2150 17985 2180
rect 17945 2130 17955 2150
rect 17975 2130 17985 2150
rect 15815 2100 15855 2130
rect 15815 2080 15825 2100
rect 15845 2080 15855 2100
rect 15815 2050 15855 2080
rect 15815 2030 15825 2050
rect 15845 2030 15855 2050
rect 15815 2000 15855 2030
rect 15815 1980 15825 2000
rect 15845 1980 15855 2000
rect 16275 2115 16315 2130
rect 16275 2095 16285 2115
rect 16305 2095 16315 2115
rect 16275 2065 16315 2095
rect 16275 2045 16285 2065
rect 16305 2045 16315 2065
rect 16275 2015 16315 2045
rect 16275 1995 16285 2015
rect 16305 1995 16315 2015
rect 16275 1980 16315 1995
rect 16330 2115 16370 2130
rect 16330 2095 16340 2115
rect 16360 2095 16370 2115
rect 16330 2065 16370 2095
rect 16330 2045 16340 2065
rect 16360 2045 16370 2065
rect 16330 2015 16370 2045
rect 16330 1995 16340 2015
rect 16360 1995 16370 2015
rect 16330 1980 16370 1995
rect 16385 2115 16425 2130
rect 16385 2095 16395 2115
rect 16415 2095 16425 2115
rect 16385 2065 16425 2095
rect 16385 2045 16395 2065
rect 16415 2045 16425 2065
rect 16385 2015 16425 2045
rect 16385 1995 16395 2015
rect 16415 1995 16425 2015
rect 16385 1980 16425 1995
rect 16440 2115 16480 2130
rect 16440 2095 16450 2115
rect 16470 2095 16480 2115
rect 16440 2065 16480 2095
rect 16440 2045 16450 2065
rect 16470 2045 16480 2065
rect 16440 2015 16480 2045
rect 16440 1995 16450 2015
rect 16470 1995 16480 2015
rect 16440 1980 16480 1995
rect 16495 2115 16535 2130
rect 16495 2095 16505 2115
rect 16525 2095 16535 2115
rect 16495 2065 16535 2095
rect 16495 2045 16505 2065
rect 16525 2045 16535 2065
rect 16495 2015 16535 2045
rect 16495 1995 16505 2015
rect 16525 1995 16535 2015
rect 16495 1980 16535 1995
rect 16550 2115 16590 2130
rect 16550 2095 16560 2115
rect 16580 2095 16590 2115
rect 16550 2065 16590 2095
rect 16550 2045 16560 2065
rect 16580 2045 16590 2065
rect 16550 2015 16590 2045
rect 16550 1995 16560 2015
rect 16580 1995 16590 2015
rect 16550 1980 16590 1995
rect 16605 2115 16645 2130
rect 16605 2095 16615 2115
rect 16635 2095 16645 2115
rect 16605 2065 16645 2095
rect 16605 2045 16615 2065
rect 16635 2045 16645 2065
rect 16605 2015 16645 2045
rect 16605 1995 16615 2015
rect 16635 1995 16645 2015
rect 16605 1980 16645 1995
rect 16660 2115 16700 2130
rect 16660 2095 16670 2115
rect 16690 2095 16700 2115
rect 16660 2065 16700 2095
rect 16660 2045 16670 2065
rect 16690 2045 16700 2065
rect 16660 2015 16700 2045
rect 16660 1995 16670 2015
rect 16690 1995 16700 2015
rect 16660 1980 16700 1995
rect 16715 2115 16755 2130
rect 16715 2095 16725 2115
rect 16745 2095 16755 2115
rect 16715 2065 16755 2095
rect 16715 2045 16725 2065
rect 16745 2045 16755 2065
rect 16715 2015 16755 2045
rect 16715 1995 16725 2015
rect 16745 1995 16755 2015
rect 16715 1980 16755 1995
rect 16770 2115 16810 2130
rect 16770 2095 16780 2115
rect 16800 2095 16810 2115
rect 16770 2065 16810 2095
rect 16770 2045 16780 2065
rect 16800 2045 16810 2065
rect 16770 2015 16810 2045
rect 16770 1995 16780 2015
rect 16800 1995 16810 2015
rect 16770 1980 16810 1995
rect 16825 2115 16865 2130
rect 16825 2095 16835 2115
rect 16855 2095 16865 2115
rect 16825 2065 16865 2095
rect 16825 2045 16835 2065
rect 16855 2045 16865 2065
rect 16825 2015 16865 2045
rect 16825 1995 16835 2015
rect 16855 1995 16865 2015
rect 16825 1980 16865 1995
rect 16880 2115 16920 2130
rect 16880 2095 16890 2115
rect 16910 2095 16920 2115
rect 16880 2065 16920 2095
rect 16880 2045 16890 2065
rect 16910 2045 16920 2065
rect 16880 2015 16920 2045
rect 16880 1995 16890 2015
rect 16910 1995 16920 2015
rect 16880 1980 16920 1995
rect 16935 2115 16975 2130
rect 16935 2095 16945 2115
rect 16965 2095 16975 2115
rect 16935 2065 16975 2095
rect 16935 2045 16945 2065
rect 16965 2045 16975 2065
rect 16935 2015 16975 2045
rect 16935 1995 16945 2015
rect 16965 1995 16975 2015
rect 16935 1980 16975 1995
rect 16990 2115 17030 2130
rect 16990 2095 17000 2115
rect 17020 2095 17030 2115
rect 16990 2065 17030 2095
rect 16990 2045 17000 2065
rect 17020 2045 17030 2065
rect 16990 2015 17030 2045
rect 16990 1995 17000 2015
rect 17020 1995 17030 2015
rect 16990 1980 17030 1995
rect 17045 2115 17085 2130
rect 17045 2095 17055 2115
rect 17075 2095 17085 2115
rect 17045 2065 17085 2095
rect 17045 2045 17055 2065
rect 17075 2045 17085 2065
rect 17045 2015 17085 2045
rect 17045 1995 17055 2015
rect 17075 1995 17085 2015
rect 17045 1980 17085 1995
rect 17100 2115 17140 2130
rect 17100 2095 17110 2115
rect 17130 2095 17140 2115
rect 17100 2065 17140 2095
rect 17100 2045 17110 2065
rect 17130 2045 17140 2065
rect 17100 2015 17140 2045
rect 17100 1995 17110 2015
rect 17130 1995 17140 2015
rect 17100 1980 17140 1995
rect 17155 2115 17195 2130
rect 17155 2095 17165 2115
rect 17185 2095 17195 2115
rect 17155 2065 17195 2095
rect 17155 2045 17165 2065
rect 17185 2045 17195 2065
rect 17155 2015 17195 2045
rect 17155 1995 17165 2015
rect 17185 1995 17195 2015
rect 17155 1980 17195 1995
rect 17210 2115 17250 2130
rect 17210 2095 17220 2115
rect 17240 2095 17250 2115
rect 17210 2065 17250 2095
rect 17210 2045 17220 2065
rect 17240 2045 17250 2065
rect 17210 2015 17250 2045
rect 17210 1995 17220 2015
rect 17240 1995 17250 2015
rect 17210 1980 17250 1995
rect 17265 2115 17305 2130
rect 17265 2095 17275 2115
rect 17295 2095 17305 2115
rect 17265 2065 17305 2095
rect 17265 2045 17275 2065
rect 17295 2045 17305 2065
rect 17265 2015 17305 2045
rect 17265 1995 17275 2015
rect 17295 1995 17305 2015
rect 17265 1980 17305 1995
rect 17320 2115 17360 2130
rect 17320 2095 17330 2115
rect 17350 2095 17360 2115
rect 17320 2065 17360 2095
rect 17320 2045 17330 2065
rect 17350 2045 17360 2065
rect 17320 2015 17360 2045
rect 17320 1995 17330 2015
rect 17350 1995 17360 2015
rect 17320 1980 17360 1995
rect 17375 2115 17415 2130
rect 17375 2095 17385 2115
rect 17405 2095 17415 2115
rect 17375 2065 17415 2095
rect 17375 2045 17385 2065
rect 17405 2045 17415 2065
rect 17375 2015 17415 2045
rect 17375 1995 17385 2015
rect 17405 1995 17415 2015
rect 17375 1980 17415 1995
rect 17430 2115 17470 2130
rect 17430 2095 17440 2115
rect 17460 2095 17470 2115
rect 17430 2065 17470 2095
rect 17430 2045 17440 2065
rect 17460 2045 17470 2065
rect 17430 2015 17470 2045
rect 17430 1995 17440 2015
rect 17460 1995 17470 2015
rect 17430 1980 17470 1995
rect 17485 2115 17525 2130
rect 17485 2095 17495 2115
rect 17515 2095 17525 2115
rect 17485 2065 17525 2095
rect 17485 2045 17495 2065
rect 17515 2045 17525 2065
rect 17485 2015 17525 2045
rect 17485 1995 17495 2015
rect 17515 1995 17525 2015
rect 17485 1980 17525 1995
rect 17945 2100 17985 2130
rect 17945 2080 17955 2100
rect 17975 2080 17985 2100
rect 17945 2050 17985 2080
rect 17945 2030 17955 2050
rect 17975 2030 17985 2050
rect 17945 2000 17985 2030
rect 17945 1980 17955 2000
rect 17975 1980 17985 2000
rect 15815 1965 15855 1980
rect 17945 1965 17985 1980
rect 18000 2250 18040 2265
rect 18000 2230 18010 2250
rect 18030 2230 18040 2250
rect 18000 2200 18040 2230
rect 18000 2180 18010 2200
rect 18030 2180 18040 2200
rect 18000 2150 18040 2180
rect 18000 2130 18010 2150
rect 18030 2130 18040 2150
rect 18000 2100 18040 2130
rect 18000 2080 18010 2100
rect 18030 2080 18040 2100
rect 18000 2050 18040 2080
rect 18000 2030 18010 2050
rect 18030 2030 18040 2050
rect 18000 2000 18040 2030
rect 18000 1980 18010 2000
rect 18030 1980 18040 2000
rect 18000 1965 18040 1980
rect 18055 2250 18095 2265
rect 18055 2230 18065 2250
rect 18085 2230 18095 2250
rect 18055 2200 18095 2230
rect 18055 2180 18065 2200
rect 18085 2180 18095 2200
rect 18055 2150 18095 2180
rect 18055 2130 18065 2150
rect 18085 2130 18095 2150
rect 18055 2100 18095 2130
rect 18055 2080 18065 2100
rect 18085 2080 18095 2100
rect 18055 2050 18095 2080
rect 18055 2030 18065 2050
rect 18085 2030 18095 2050
rect 18055 2000 18095 2030
rect 18055 1980 18065 2000
rect 18085 1980 18095 2000
rect 18055 1965 18095 1980
rect 18110 2250 18150 2265
rect 18110 2230 18120 2250
rect 18140 2230 18150 2250
rect 18110 2200 18150 2230
rect 18110 2180 18120 2200
rect 18140 2180 18150 2200
rect 18110 2150 18150 2180
rect 18110 2130 18120 2150
rect 18140 2130 18150 2150
rect 18110 2100 18150 2130
rect 18110 2080 18120 2100
rect 18140 2080 18150 2100
rect 18110 2050 18150 2080
rect 18110 2030 18120 2050
rect 18140 2030 18150 2050
rect 18110 2000 18150 2030
rect 18110 1980 18120 2000
rect 18140 1980 18150 2000
rect 18110 1965 18150 1980
rect 18165 2250 18205 2265
rect 18165 2230 18175 2250
rect 18195 2230 18205 2250
rect 18165 2200 18205 2230
rect 18165 2180 18175 2200
rect 18195 2180 18205 2200
rect 18165 2150 18205 2180
rect 18165 2130 18175 2150
rect 18195 2130 18205 2150
rect 18165 2100 18205 2130
rect 18165 2080 18175 2100
rect 18195 2080 18205 2100
rect 18165 2050 18205 2080
rect 18165 2030 18175 2050
rect 18195 2030 18205 2050
rect 18165 2000 18205 2030
rect 18165 1980 18175 2000
rect 18195 1980 18205 2000
rect 18165 1965 18205 1980
rect 18220 2250 18260 2265
rect 18220 2230 18230 2250
rect 18250 2230 18260 2250
rect 18220 2200 18260 2230
rect 18220 2180 18230 2200
rect 18250 2180 18260 2200
rect 18220 2150 18260 2180
rect 18220 2130 18230 2150
rect 18250 2130 18260 2150
rect 18220 2100 18260 2130
rect 18220 2080 18230 2100
rect 18250 2080 18260 2100
rect 18220 2050 18260 2080
rect 18220 2030 18230 2050
rect 18250 2030 18260 2050
rect 18220 2000 18260 2030
rect 18220 1980 18230 2000
rect 18250 1980 18260 2000
rect 18220 1965 18260 1980
rect 18275 2250 18315 2265
rect 18275 2230 18285 2250
rect 18305 2230 18315 2250
rect 18275 2200 18315 2230
rect 18275 2180 18285 2200
rect 18305 2180 18315 2200
rect 18275 2150 18315 2180
rect 18275 2130 18285 2150
rect 18305 2130 18315 2150
rect 18275 2100 18315 2130
rect 18275 2080 18285 2100
rect 18305 2080 18315 2100
rect 18275 2050 18315 2080
rect 18275 2030 18285 2050
rect 18305 2030 18315 2050
rect 18275 2000 18315 2030
rect 18275 1980 18285 2000
rect 18305 1980 18315 2000
rect 18275 1965 18315 1980
rect 18330 2250 18370 2265
rect 18330 2230 18340 2250
rect 18360 2230 18370 2250
rect 18330 2200 18370 2230
rect 18330 2180 18340 2200
rect 18360 2180 18370 2200
rect 18330 2150 18370 2180
rect 18330 2130 18340 2150
rect 18360 2130 18370 2150
rect 18330 2100 18370 2130
rect 18330 2080 18340 2100
rect 18360 2080 18370 2100
rect 18330 2050 18370 2080
rect 18330 2030 18340 2050
rect 18360 2030 18370 2050
rect 18330 2000 18370 2030
rect 18330 1980 18340 2000
rect 18360 1980 18370 2000
rect 18330 1965 18370 1980
rect 18385 2250 18425 2265
rect 18385 2230 18395 2250
rect 18415 2230 18425 2250
rect 18385 2200 18425 2230
rect 18385 2180 18395 2200
rect 18415 2180 18425 2200
rect 18385 2150 18425 2180
rect 18385 2130 18395 2150
rect 18415 2130 18425 2150
rect 18385 2100 18425 2130
rect 18385 2080 18395 2100
rect 18415 2080 18425 2100
rect 18385 2050 18425 2080
rect 18385 2030 18395 2050
rect 18415 2030 18425 2050
rect 18385 2000 18425 2030
rect 18385 1980 18395 2000
rect 18415 1980 18425 2000
rect 18385 1965 18425 1980
rect 18440 2250 18480 2265
rect 18440 2230 18450 2250
rect 18470 2230 18480 2250
rect 18440 2200 18480 2230
rect 18440 2180 18450 2200
rect 18470 2180 18480 2200
rect 18440 2150 18480 2180
rect 18440 2130 18450 2150
rect 18470 2130 18480 2150
rect 18440 2100 18480 2130
rect 18440 2080 18450 2100
rect 18470 2080 18480 2100
rect 18440 2050 18480 2080
rect 18440 2030 18450 2050
rect 18470 2030 18480 2050
rect 18440 2000 18480 2030
rect 18440 1980 18450 2000
rect 18470 1980 18480 2000
rect 18440 1965 18480 1980
rect 18495 2250 18535 2265
rect 18495 2230 18505 2250
rect 18525 2230 18535 2250
rect 18495 2200 18535 2230
rect 18495 2180 18505 2200
rect 18525 2180 18535 2200
rect 18495 2150 18535 2180
rect 18495 2130 18505 2150
rect 18525 2130 18535 2150
rect 18495 2100 18535 2130
rect 18495 2080 18505 2100
rect 18525 2080 18535 2100
rect 18495 2050 18535 2080
rect 18495 2030 18505 2050
rect 18525 2030 18535 2050
rect 18495 2000 18535 2030
rect 18495 1980 18505 2000
rect 18525 1980 18535 2000
rect 18495 1965 18535 1980
rect 18550 2250 18590 2265
rect 18550 2230 18560 2250
rect 18580 2230 18590 2250
rect 18550 2200 18590 2230
rect 18550 2180 18560 2200
rect 18580 2180 18590 2200
rect 18550 2150 18590 2180
rect 18550 2130 18560 2150
rect 18580 2130 18590 2150
rect 18550 2100 18590 2130
rect 18550 2080 18560 2100
rect 18580 2080 18590 2100
rect 18550 2050 18590 2080
rect 18550 2030 18560 2050
rect 18580 2030 18590 2050
rect 18550 2000 18590 2030
rect 18550 1980 18560 2000
rect 18580 1980 18590 2000
rect 18550 1965 18590 1980
rect 18605 2250 18645 2265
rect 18605 2230 18615 2250
rect 18635 2230 18645 2250
rect 18605 2200 18645 2230
rect 18605 2180 18615 2200
rect 18635 2180 18645 2200
rect 18605 2150 18645 2180
rect 18605 2130 18615 2150
rect 18635 2130 18645 2150
rect 18605 2100 18645 2130
rect 18605 2080 18615 2100
rect 18635 2080 18645 2100
rect 18605 2050 18645 2080
rect 18605 2030 18615 2050
rect 18635 2030 18645 2050
rect 18605 2000 18645 2030
rect 18605 1980 18615 2000
rect 18635 1980 18645 2000
rect 18605 1965 18645 1980
rect 3165 1650 3205 1665
rect 3165 1630 3175 1650
rect 3195 1630 3205 1650
rect 3165 1615 3205 1630
rect 3225 1650 3265 1665
rect 3225 1630 3235 1650
rect 3255 1630 3265 1650
rect 3225 1615 3265 1630
rect 3285 1650 3325 1665
rect 3285 1630 3295 1650
rect 3315 1630 3325 1650
rect 3285 1615 3325 1630
rect 3345 1650 3385 1665
rect 3345 1630 3355 1650
rect 3375 1630 3385 1650
rect 3345 1615 3385 1630
rect 3405 1650 3445 1665
rect 3405 1630 3415 1650
rect 3435 1630 3445 1650
rect 3405 1615 3445 1630
rect 3465 1650 3505 1665
rect 3465 1630 3475 1650
rect 3495 1630 3505 1650
rect 3465 1615 3505 1630
rect 3525 1650 3565 1665
rect 3525 1630 3535 1650
rect 3555 1630 3565 1650
rect 3525 1615 3565 1630
rect 3585 1650 3625 1665
rect 3585 1630 3595 1650
rect 3615 1630 3625 1650
rect 3585 1615 3625 1630
rect 3645 1650 3685 1665
rect 3645 1630 3655 1650
rect 3675 1630 3685 1650
rect 3645 1615 3685 1630
rect 3705 1650 3745 1665
rect 3705 1630 3715 1650
rect 3735 1630 3745 1650
rect 3705 1615 3745 1630
rect 3765 1650 3805 1665
rect 3765 1630 3775 1650
rect 3795 1630 3805 1650
rect 3765 1615 3805 1630
rect 4205 1650 4245 1665
rect 4205 1630 4215 1650
rect 4235 1630 4245 1650
rect 4205 1615 4245 1630
rect 4265 1650 4305 1665
rect 4265 1630 4275 1650
rect 4295 1630 4305 1650
rect 4265 1615 4305 1630
rect 4325 1650 4365 1665
rect 4325 1630 4335 1650
rect 4355 1630 4365 1650
rect 4325 1615 4365 1630
rect 4385 1650 4425 1665
rect 4385 1630 4395 1650
rect 4415 1630 4425 1650
rect 4385 1615 4425 1630
rect 4445 1650 4485 1665
rect 4445 1630 4455 1650
rect 4475 1630 4485 1650
rect 4445 1615 4485 1630
rect 4505 1650 4545 1665
rect 4505 1630 4515 1650
rect 4535 1630 4545 1650
rect 4505 1615 4545 1630
rect 4565 1650 4605 1665
rect 4565 1630 4575 1650
rect 4595 1630 4605 1650
rect 4565 1615 4605 1630
rect 4625 1650 4665 1665
rect 4625 1630 4635 1650
rect 4655 1630 4665 1650
rect 4625 1615 4665 1630
rect 4685 1650 4725 1665
rect 4685 1630 4695 1650
rect 4715 1630 4725 1650
rect 4685 1615 4725 1630
rect 4745 1650 4785 1665
rect 4745 1630 4755 1650
rect 4775 1630 4785 1650
rect 4745 1615 4785 1630
rect 4805 1650 4845 1665
rect 4805 1630 4815 1650
rect 4835 1630 4845 1650
rect 4805 1615 4845 1630
rect 15155 1640 15195 1655
rect 15155 1620 15165 1640
rect 15185 1620 15195 1640
rect 2835 1440 2875 1455
rect 2835 1420 2845 1440
rect 2865 1420 2875 1440
rect 2835 1390 2875 1420
rect 2835 1370 2845 1390
rect 2865 1370 2875 1390
rect 2835 1340 2875 1370
rect 2835 1320 2845 1340
rect 2865 1320 2875 1340
rect 2835 1290 2875 1320
rect 2835 1270 2845 1290
rect 2865 1270 2875 1290
rect 2835 1240 2875 1270
rect 2835 1220 2845 1240
rect 2865 1220 2875 1240
rect 2835 1205 2875 1220
rect 3375 1440 3415 1455
rect 3375 1420 3385 1440
rect 3405 1420 3415 1440
rect 3375 1390 3415 1420
rect 3375 1370 3385 1390
rect 3405 1370 3415 1390
rect 3375 1340 3415 1370
rect 3375 1320 3385 1340
rect 3405 1320 3415 1340
rect 3375 1290 3415 1320
rect 3375 1270 3385 1290
rect 3405 1270 3415 1290
rect 3375 1240 3415 1270
rect 3375 1220 3385 1240
rect 3405 1220 3415 1240
rect 3375 1205 3415 1220
rect 3915 1440 3955 1455
rect 3915 1420 3925 1440
rect 3945 1420 3955 1440
rect 3915 1390 3955 1420
rect 3915 1370 3925 1390
rect 3945 1370 3955 1390
rect 3915 1340 3955 1370
rect 3915 1320 3925 1340
rect 3945 1320 3955 1340
rect 3915 1290 3955 1320
rect 3915 1270 3925 1290
rect 3945 1270 3955 1290
rect 3915 1240 3955 1270
rect 3915 1220 3925 1240
rect 3945 1220 3955 1240
rect 3915 1205 3955 1220
rect 4055 1440 4095 1455
rect 4055 1420 4065 1440
rect 4085 1420 4095 1440
rect 4055 1390 4095 1420
rect 4055 1370 4065 1390
rect 4085 1370 4095 1390
rect 4055 1340 4095 1370
rect 4055 1320 4065 1340
rect 4085 1320 4095 1340
rect 4055 1290 4095 1320
rect 4055 1270 4065 1290
rect 4085 1270 4095 1290
rect 4055 1240 4095 1270
rect 4055 1220 4065 1240
rect 4085 1220 4095 1240
rect 4055 1205 4095 1220
rect 4595 1440 4635 1455
rect 4595 1420 4605 1440
rect 4625 1420 4635 1440
rect 4595 1390 4635 1420
rect 4595 1370 4605 1390
rect 4625 1370 4635 1390
rect 4595 1340 4635 1370
rect 4595 1320 4605 1340
rect 4625 1320 4635 1340
rect 4595 1290 4635 1320
rect 4595 1270 4605 1290
rect 4625 1270 4635 1290
rect 4595 1240 4635 1270
rect 4595 1220 4605 1240
rect 4625 1220 4635 1240
rect 4595 1205 4635 1220
rect 5135 1440 5175 1455
rect 5135 1420 5145 1440
rect 5165 1420 5175 1440
rect 5135 1390 5175 1420
rect 5135 1370 5145 1390
rect 5165 1370 5175 1390
rect 5135 1340 5175 1370
rect 5135 1320 5145 1340
rect 5165 1320 5175 1340
rect 5135 1290 5175 1320
rect 5135 1270 5145 1290
rect 5165 1270 5175 1290
rect 5135 1240 5175 1270
rect 5135 1220 5145 1240
rect 5165 1220 5175 1240
rect 5135 1205 5175 1220
rect 2945 1060 2985 1075
rect 2945 1040 2955 1060
rect 2975 1040 2985 1060
rect 2945 1010 2985 1040
rect 2945 990 2955 1010
rect 2975 990 2985 1010
rect 2945 975 2985 990
rect 3985 1060 4025 1075
rect 3985 1040 3995 1060
rect 4015 1040 4025 1060
rect 3985 1010 4025 1040
rect 3985 990 3995 1010
rect 4015 990 4025 1010
rect 3985 975 4025 990
rect 5025 1060 5065 1075
rect 5025 1040 5035 1060
rect 5055 1040 5065 1060
rect 5025 1010 5065 1040
rect 5025 990 5035 1010
rect 5055 990 5065 1010
rect 5025 975 5065 990
rect 15155 1590 15195 1620
rect 15155 1570 15165 1590
rect 15185 1570 15195 1590
rect 15155 1540 15195 1570
rect 15155 1520 15165 1540
rect 15185 1520 15195 1540
rect 15155 1490 15195 1520
rect 15155 1470 15165 1490
rect 15185 1470 15195 1490
rect 15155 1440 15195 1470
rect 15155 1420 15165 1440
rect 15185 1420 15195 1440
rect 15155 1390 15195 1420
rect 15155 1370 15165 1390
rect 15185 1370 15195 1390
rect 15155 1340 15195 1370
rect 15155 1320 15165 1340
rect 15185 1320 15195 1340
rect 15155 1290 15195 1320
rect 15155 1270 15165 1290
rect 15185 1270 15195 1290
rect 15155 1240 15195 1270
rect 15155 1220 15165 1240
rect 15185 1220 15195 1240
rect 15155 1190 15195 1220
rect 15155 1170 15165 1190
rect 15185 1170 15195 1190
rect 15155 1140 15195 1170
rect 15155 1120 15165 1140
rect 15185 1120 15195 1140
rect 15155 1090 15195 1120
rect 15155 1070 15165 1090
rect 15185 1070 15195 1090
rect 15155 1040 15195 1070
rect 15155 1020 15165 1040
rect 15185 1020 15195 1040
rect 15155 990 15195 1020
rect 15155 970 15165 990
rect 15185 970 15195 990
rect 15155 955 15195 970
rect 15255 1640 15295 1655
rect 15255 1620 15265 1640
rect 15285 1620 15295 1640
rect 15255 1590 15295 1620
rect 15255 1570 15265 1590
rect 15285 1570 15295 1590
rect 15255 1540 15295 1570
rect 15255 1520 15265 1540
rect 15285 1520 15295 1540
rect 15255 1490 15295 1520
rect 15255 1470 15265 1490
rect 15285 1470 15295 1490
rect 15255 1440 15295 1470
rect 15255 1420 15265 1440
rect 15285 1420 15295 1440
rect 15255 1390 15295 1420
rect 15255 1370 15265 1390
rect 15285 1370 15295 1390
rect 15255 1340 15295 1370
rect 15255 1320 15265 1340
rect 15285 1320 15295 1340
rect 15255 1290 15295 1320
rect 15255 1270 15265 1290
rect 15285 1270 15295 1290
rect 15255 1240 15295 1270
rect 15255 1220 15265 1240
rect 15285 1220 15295 1240
rect 15255 1190 15295 1220
rect 15255 1170 15265 1190
rect 15285 1170 15295 1190
rect 15255 1140 15295 1170
rect 15255 1120 15265 1140
rect 15285 1120 15295 1140
rect 15255 1090 15295 1120
rect 15255 1070 15265 1090
rect 15285 1070 15295 1090
rect 15255 1040 15295 1070
rect 15255 1020 15265 1040
rect 15285 1020 15295 1040
rect 15255 990 15295 1020
rect 15255 970 15265 990
rect 15285 970 15295 990
rect 15255 955 15295 970
rect 15355 1640 15395 1655
rect 15355 1620 15365 1640
rect 15385 1620 15395 1640
rect 15355 1590 15395 1620
rect 15355 1570 15365 1590
rect 15385 1570 15395 1590
rect 15355 1540 15395 1570
rect 15355 1520 15365 1540
rect 15385 1520 15395 1540
rect 15355 1490 15395 1520
rect 15355 1470 15365 1490
rect 15385 1470 15395 1490
rect 15355 1440 15395 1470
rect 15355 1420 15365 1440
rect 15385 1420 15395 1440
rect 15355 1390 15395 1420
rect 15355 1370 15365 1390
rect 15385 1370 15395 1390
rect 15355 1340 15395 1370
rect 15355 1320 15365 1340
rect 15385 1320 15395 1340
rect 15355 1290 15395 1320
rect 15355 1270 15365 1290
rect 15385 1270 15395 1290
rect 15355 1240 15395 1270
rect 15355 1220 15365 1240
rect 15385 1220 15395 1240
rect 15355 1190 15395 1220
rect 15355 1170 15365 1190
rect 15385 1170 15395 1190
rect 15355 1140 15395 1170
rect 15355 1120 15365 1140
rect 15385 1120 15395 1140
rect 15355 1090 15395 1120
rect 15355 1070 15365 1090
rect 15385 1070 15395 1090
rect 15355 1040 15395 1070
rect 15355 1020 15365 1040
rect 15385 1020 15395 1040
rect 15355 990 15395 1020
rect 15355 970 15365 990
rect 15385 970 15395 990
rect 15355 955 15395 970
rect 15455 1640 15495 1655
rect 15455 1620 15465 1640
rect 15485 1620 15495 1640
rect 15455 1590 15495 1620
rect 15455 1570 15465 1590
rect 15485 1570 15495 1590
rect 15455 1540 15495 1570
rect 15455 1520 15465 1540
rect 15485 1520 15495 1540
rect 15455 1490 15495 1520
rect 15455 1470 15465 1490
rect 15485 1470 15495 1490
rect 15455 1440 15495 1470
rect 15455 1420 15465 1440
rect 15485 1420 15495 1440
rect 15455 1390 15495 1420
rect 15455 1370 15465 1390
rect 15485 1370 15495 1390
rect 15455 1340 15495 1370
rect 15455 1320 15465 1340
rect 15485 1320 15495 1340
rect 15455 1290 15495 1320
rect 15455 1270 15465 1290
rect 15485 1270 15495 1290
rect 15455 1240 15495 1270
rect 15455 1220 15465 1240
rect 15485 1220 15495 1240
rect 15455 1190 15495 1220
rect 15455 1170 15465 1190
rect 15485 1170 15495 1190
rect 15455 1140 15495 1170
rect 15455 1120 15465 1140
rect 15485 1120 15495 1140
rect 15455 1090 15495 1120
rect 15455 1070 15465 1090
rect 15485 1070 15495 1090
rect 15455 1040 15495 1070
rect 15455 1020 15465 1040
rect 15485 1020 15495 1040
rect 15455 990 15495 1020
rect 15455 970 15465 990
rect 15485 970 15495 990
rect 15455 955 15495 970
rect 15555 1640 15595 1655
rect 15555 1620 15565 1640
rect 15585 1620 15595 1640
rect 15555 1590 15595 1620
rect 15555 1570 15565 1590
rect 15585 1570 15595 1590
rect 15555 1540 15595 1570
rect 15555 1520 15565 1540
rect 15585 1520 15595 1540
rect 15555 1490 15595 1520
rect 15555 1470 15565 1490
rect 15585 1470 15595 1490
rect 15555 1440 15595 1470
rect 15555 1420 15565 1440
rect 15585 1420 15595 1440
rect 15555 1390 15595 1420
rect 15555 1370 15565 1390
rect 15585 1370 15595 1390
rect 15555 1340 15595 1370
rect 15555 1320 15565 1340
rect 15585 1320 15595 1340
rect 15555 1290 15595 1320
rect 15555 1270 15565 1290
rect 15585 1270 15595 1290
rect 15555 1240 15595 1270
rect 15555 1220 15565 1240
rect 15585 1220 15595 1240
rect 15555 1190 15595 1220
rect 15555 1170 15565 1190
rect 15585 1170 15595 1190
rect 15555 1140 15595 1170
rect 15555 1120 15565 1140
rect 15585 1120 15595 1140
rect 15555 1090 15595 1120
rect 15555 1070 15565 1090
rect 15585 1070 15595 1090
rect 15555 1040 15595 1070
rect 15555 1020 15565 1040
rect 15585 1020 15595 1040
rect 15555 990 15595 1020
rect 15555 970 15565 990
rect 15585 970 15595 990
rect 15555 955 15595 970
rect 15655 1640 15695 1655
rect 15655 1620 15665 1640
rect 15685 1620 15695 1640
rect 15655 1590 15695 1620
rect 15655 1570 15665 1590
rect 15685 1570 15695 1590
rect 15655 1540 15695 1570
rect 15655 1520 15665 1540
rect 15685 1520 15695 1540
rect 15655 1490 15695 1520
rect 15655 1470 15665 1490
rect 15685 1470 15695 1490
rect 15655 1440 15695 1470
rect 15655 1420 15665 1440
rect 15685 1420 15695 1440
rect 15655 1390 15695 1420
rect 15655 1370 15665 1390
rect 15685 1370 15695 1390
rect 15655 1340 15695 1370
rect 15655 1320 15665 1340
rect 15685 1320 15695 1340
rect 15655 1290 15695 1320
rect 15655 1270 15665 1290
rect 15685 1270 15695 1290
rect 15655 1240 15695 1270
rect 15655 1220 15665 1240
rect 15685 1220 15695 1240
rect 15655 1190 15695 1220
rect 15655 1170 15665 1190
rect 15685 1170 15695 1190
rect 15655 1140 15695 1170
rect 15655 1120 15665 1140
rect 15685 1120 15695 1140
rect 15655 1090 15695 1120
rect 15655 1070 15665 1090
rect 15685 1070 15695 1090
rect 15655 1040 15695 1070
rect 15655 1020 15665 1040
rect 15685 1020 15695 1040
rect 15655 990 15695 1020
rect 15655 970 15665 990
rect 15685 970 15695 990
rect 15655 955 15695 970
rect 15755 1640 15795 1655
rect 15755 1620 15765 1640
rect 15785 1620 15795 1640
rect 15755 1590 15795 1620
rect 15755 1570 15765 1590
rect 15785 1570 15795 1590
rect 15755 1540 15795 1570
rect 15755 1520 15765 1540
rect 15785 1520 15795 1540
rect 15755 1490 15795 1520
rect 16030 1650 16070 1665
rect 16030 1630 16040 1650
rect 16060 1630 16070 1650
rect 16030 1600 16070 1630
rect 16030 1580 16040 1600
rect 16060 1580 16070 1600
rect 16030 1550 16070 1580
rect 16030 1530 16040 1550
rect 16060 1530 16070 1550
rect 16030 1515 16070 1530
rect 16085 1650 16125 1665
rect 16085 1630 16095 1650
rect 16115 1630 16125 1650
rect 16085 1600 16125 1630
rect 16085 1580 16095 1600
rect 16115 1580 16125 1600
rect 16085 1550 16125 1580
rect 16085 1530 16095 1550
rect 16115 1530 16125 1550
rect 16085 1515 16125 1530
rect 16140 1650 16180 1665
rect 16140 1630 16150 1650
rect 16170 1630 16180 1650
rect 16140 1600 16180 1630
rect 16140 1580 16150 1600
rect 16170 1580 16180 1600
rect 16140 1550 16180 1580
rect 16140 1530 16150 1550
rect 16170 1530 16180 1550
rect 16140 1515 16180 1530
rect 16195 1650 16235 1665
rect 16195 1630 16205 1650
rect 16225 1630 16235 1650
rect 16195 1600 16235 1630
rect 16195 1580 16205 1600
rect 16225 1580 16235 1600
rect 16195 1550 16235 1580
rect 16195 1530 16205 1550
rect 16225 1530 16235 1550
rect 16195 1515 16235 1530
rect 16250 1650 16290 1665
rect 16250 1630 16260 1650
rect 16280 1630 16290 1650
rect 16250 1600 16290 1630
rect 16250 1580 16260 1600
rect 16280 1580 16290 1600
rect 16250 1550 16290 1580
rect 16250 1530 16260 1550
rect 16280 1530 16290 1550
rect 16250 1515 16290 1530
rect 16305 1650 16345 1665
rect 16305 1630 16315 1650
rect 16335 1630 16345 1650
rect 16305 1600 16345 1630
rect 16305 1580 16315 1600
rect 16335 1580 16345 1600
rect 16305 1550 16345 1580
rect 16305 1530 16315 1550
rect 16335 1530 16345 1550
rect 16305 1515 16345 1530
rect 16360 1650 16400 1665
rect 16360 1630 16370 1650
rect 16390 1630 16400 1650
rect 16360 1600 16400 1630
rect 16360 1580 16370 1600
rect 16390 1580 16400 1600
rect 16360 1550 16400 1580
rect 16360 1530 16370 1550
rect 16390 1530 16400 1550
rect 16360 1515 16400 1530
rect 16415 1650 16455 1665
rect 16415 1630 16425 1650
rect 16445 1630 16455 1650
rect 16415 1600 16455 1630
rect 16415 1580 16425 1600
rect 16445 1580 16455 1600
rect 16415 1550 16455 1580
rect 16415 1530 16425 1550
rect 16445 1530 16455 1550
rect 16415 1515 16455 1530
rect 16470 1650 16510 1665
rect 16470 1630 16480 1650
rect 16500 1630 16510 1650
rect 16470 1600 16510 1630
rect 16470 1580 16480 1600
rect 16500 1580 16510 1600
rect 16470 1550 16510 1580
rect 16470 1530 16480 1550
rect 16500 1530 16510 1550
rect 16470 1515 16510 1530
rect 16525 1650 16565 1665
rect 16525 1630 16535 1650
rect 16555 1630 16565 1650
rect 16525 1600 16565 1630
rect 16525 1580 16535 1600
rect 16555 1580 16565 1600
rect 16525 1550 16565 1580
rect 16525 1530 16535 1550
rect 16555 1530 16565 1550
rect 16525 1515 16565 1530
rect 16580 1650 16620 1665
rect 16580 1630 16590 1650
rect 16610 1630 16620 1650
rect 16580 1600 16620 1630
rect 16580 1580 16590 1600
rect 16610 1580 16620 1600
rect 16580 1550 16620 1580
rect 16580 1530 16590 1550
rect 16610 1530 16620 1550
rect 16580 1515 16620 1530
rect 16635 1650 16675 1665
rect 16635 1630 16645 1650
rect 16665 1630 16675 1650
rect 16635 1600 16675 1630
rect 16635 1580 16645 1600
rect 16665 1580 16675 1600
rect 16635 1550 16675 1580
rect 16635 1530 16645 1550
rect 16665 1530 16675 1550
rect 16635 1515 16675 1530
rect 16690 1650 16730 1665
rect 16770 1650 16810 1665
rect 16690 1630 16700 1650
rect 16720 1630 16730 1650
rect 16770 1630 16780 1650
rect 16800 1630 16810 1650
rect 16690 1600 16730 1630
rect 16770 1600 16810 1630
rect 16690 1580 16700 1600
rect 16720 1580 16730 1600
rect 16770 1580 16780 1600
rect 16800 1580 16810 1600
rect 16690 1550 16730 1580
rect 16770 1550 16810 1580
rect 16690 1530 16700 1550
rect 16720 1530 16730 1550
rect 16770 1530 16780 1550
rect 16800 1530 16810 1550
rect 16690 1515 16730 1530
rect 16770 1515 16810 1530
rect 16825 1650 16865 1665
rect 16825 1630 16835 1650
rect 16855 1630 16865 1650
rect 16825 1600 16865 1630
rect 16825 1580 16835 1600
rect 16855 1580 16865 1600
rect 16825 1550 16865 1580
rect 16825 1530 16835 1550
rect 16855 1530 16865 1550
rect 16825 1515 16865 1530
rect 16880 1650 16920 1665
rect 16880 1630 16890 1650
rect 16910 1630 16920 1650
rect 16880 1600 16920 1630
rect 16880 1580 16890 1600
rect 16910 1580 16920 1600
rect 16880 1550 16920 1580
rect 16880 1530 16890 1550
rect 16910 1530 16920 1550
rect 16880 1515 16920 1530
rect 16935 1650 16975 1665
rect 16935 1630 16945 1650
rect 16965 1630 16975 1650
rect 16935 1600 16975 1630
rect 16935 1580 16945 1600
rect 16965 1580 16975 1600
rect 16935 1550 16975 1580
rect 16935 1530 16945 1550
rect 16965 1530 16975 1550
rect 16935 1515 16975 1530
rect 16990 1650 17030 1665
rect 17070 1650 17110 1665
rect 16990 1630 17000 1650
rect 17020 1630 17030 1650
rect 17070 1630 17080 1650
rect 17100 1630 17110 1650
rect 16990 1600 17030 1630
rect 17070 1600 17110 1630
rect 16990 1580 17000 1600
rect 17020 1580 17030 1600
rect 17070 1580 17080 1600
rect 17100 1580 17110 1600
rect 16990 1550 17030 1580
rect 17070 1550 17110 1580
rect 16990 1530 17000 1550
rect 17020 1530 17030 1550
rect 17070 1530 17080 1550
rect 17100 1530 17110 1550
rect 16990 1515 17030 1530
rect 17070 1515 17110 1530
rect 17125 1650 17165 1665
rect 17125 1630 17135 1650
rect 17155 1630 17165 1650
rect 17125 1600 17165 1630
rect 17125 1580 17135 1600
rect 17155 1580 17165 1600
rect 17125 1550 17165 1580
rect 17125 1530 17135 1550
rect 17155 1530 17165 1550
rect 17125 1515 17165 1530
rect 17180 1650 17220 1665
rect 17180 1630 17190 1650
rect 17210 1630 17220 1650
rect 17180 1600 17220 1630
rect 17180 1580 17190 1600
rect 17210 1580 17220 1600
rect 17180 1550 17220 1580
rect 17180 1530 17190 1550
rect 17210 1530 17220 1550
rect 17180 1515 17220 1530
rect 17235 1650 17275 1665
rect 17235 1630 17245 1650
rect 17265 1630 17275 1650
rect 17235 1600 17275 1630
rect 17235 1580 17245 1600
rect 17265 1580 17275 1600
rect 17235 1550 17275 1580
rect 17235 1530 17245 1550
rect 17265 1530 17275 1550
rect 17235 1515 17275 1530
rect 17290 1650 17330 1665
rect 17290 1630 17300 1650
rect 17320 1630 17330 1650
rect 17290 1600 17330 1630
rect 17290 1580 17300 1600
rect 17320 1580 17330 1600
rect 17290 1550 17330 1580
rect 17290 1530 17300 1550
rect 17320 1530 17330 1550
rect 17290 1515 17330 1530
rect 17345 1650 17385 1665
rect 17345 1630 17355 1650
rect 17375 1630 17385 1650
rect 17345 1600 17385 1630
rect 17345 1580 17355 1600
rect 17375 1580 17385 1600
rect 17345 1550 17385 1580
rect 17345 1530 17355 1550
rect 17375 1530 17385 1550
rect 17345 1515 17385 1530
rect 17400 1650 17440 1665
rect 17400 1630 17410 1650
rect 17430 1630 17440 1650
rect 17400 1600 17440 1630
rect 17400 1580 17410 1600
rect 17430 1580 17440 1600
rect 17400 1550 17440 1580
rect 17400 1530 17410 1550
rect 17430 1530 17440 1550
rect 17400 1515 17440 1530
rect 17455 1650 17495 1665
rect 17455 1630 17465 1650
rect 17485 1630 17495 1650
rect 17455 1600 17495 1630
rect 17455 1580 17465 1600
rect 17485 1580 17495 1600
rect 17455 1550 17495 1580
rect 17455 1530 17465 1550
rect 17485 1530 17495 1550
rect 17455 1515 17495 1530
rect 17510 1650 17550 1665
rect 17510 1630 17520 1650
rect 17540 1630 17550 1650
rect 17510 1600 17550 1630
rect 17510 1580 17520 1600
rect 17540 1580 17550 1600
rect 17510 1550 17550 1580
rect 17510 1530 17520 1550
rect 17540 1530 17550 1550
rect 17510 1515 17550 1530
rect 17565 1650 17605 1665
rect 17565 1630 17575 1650
rect 17595 1630 17605 1650
rect 17565 1600 17605 1630
rect 17565 1580 17575 1600
rect 17595 1580 17605 1600
rect 17565 1550 17605 1580
rect 17565 1530 17575 1550
rect 17595 1530 17605 1550
rect 17565 1515 17605 1530
rect 17620 1650 17660 1665
rect 17620 1630 17630 1650
rect 17650 1630 17660 1650
rect 17620 1600 17660 1630
rect 17620 1580 17630 1600
rect 17650 1580 17660 1600
rect 17620 1550 17660 1580
rect 17620 1530 17630 1550
rect 17650 1530 17660 1550
rect 17620 1515 17660 1530
rect 17675 1650 17715 1665
rect 17675 1630 17685 1650
rect 17705 1630 17715 1650
rect 17675 1600 17715 1630
rect 17675 1580 17685 1600
rect 17705 1580 17715 1600
rect 17675 1550 17715 1580
rect 17675 1530 17685 1550
rect 17705 1530 17715 1550
rect 17675 1515 17715 1530
rect 17730 1650 17770 1665
rect 17730 1630 17740 1650
rect 17760 1630 17770 1650
rect 17730 1600 17770 1630
rect 17730 1580 17740 1600
rect 17760 1580 17770 1600
rect 17730 1550 17770 1580
rect 17730 1530 17740 1550
rect 17760 1530 17770 1550
rect 17730 1515 17770 1530
rect 18005 1640 18045 1655
rect 18005 1620 18015 1640
rect 18035 1620 18045 1640
rect 18005 1590 18045 1620
rect 18005 1570 18015 1590
rect 18035 1570 18045 1590
rect 18005 1540 18045 1570
rect 18005 1520 18015 1540
rect 18035 1520 18045 1540
rect 15755 1470 15765 1490
rect 15785 1470 15795 1490
rect 15755 1440 15795 1470
rect 18005 1490 18045 1520
rect 18005 1470 18015 1490
rect 18035 1470 18045 1490
rect 15755 1420 15765 1440
rect 15785 1420 15795 1440
rect 15755 1390 15795 1420
rect 15755 1370 15765 1390
rect 15785 1370 15795 1390
rect 15755 1340 15795 1370
rect 15755 1320 15765 1340
rect 15785 1320 15795 1340
rect 15755 1290 15795 1320
rect 15755 1270 15765 1290
rect 15785 1270 15795 1290
rect 15755 1240 15795 1270
rect 18005 1440 18045 1470
rect 18005 1420 18015 1440
rect 18035 1420 18045 1440
rect 18005 1390 18045 1420
rect 18005 1370 18015 1390
rect 18035 1370 18045 1390
rect 18005 1340 18045 1370
rect 18005 1320 18015 1340
rect 18035 1320 18045 1340
rect 18005 1290 18045 1320
rect 18005 1270 18015 1290
rect 18035 1270 18045 1290
rect 15755 1220 15765 1240
rect 15785 1220 15795 1240
rect 15755 1190 15795 1220
rect 15755 1170 15765 1190
rect 15785 1170 15795 1190
rect 18005 1240 18045 1270
rect 18005 1220 18015 1240
rect 18035 1220 18045 1240
rect 18005 1190 18045 1220
rect 15755 1140 15795 1170
rect 15755 1120 15765 1140
rect 15785 1120 15795 1140
rect 15755 1090 15795 1120
rect 15755 1070 15765 1090
rect 15785 1070 15795 1090
rect 15755 1040 15795 1070
rect 15755 1020 15765 1040
rect 15785 1020 15795 1040
rect 15755 990 15795 1020
rect 15755 970 15765 990
rect 15785 970 15795 990
rect 15755 955 15795 970
rect 16205 1170 16245 1185
rect 16205 1150 16215 1170
rect 16235 1150 16245 1170
rect 16205 1120 16245 1150
rect 16205 1100 16215 1120
rect 16235 1100 16245 1120
rect 16205 1070 16245 1100
rect 16205 1050 16215 1070
rect 16235 1050 16245 1070
rect 16205 1020 16245 1050
rect 16205 1000 16215 1020
rect 16235 1000 16245 1020
rect 16205 970 16245 1000
rect 16205 950 16215 970
rect 16235 950 16245 970
rect 16205 935 16245 950
rect 16260 1170 16300 1185
rect 16260 1150 16270 1170
rect 16290 1150 16300 1170
rect 16260 1120 16300 1150
rect 16260 1100 16270 1120
rect 16290 1100 16300 1120
rect 16260 1070 16300 1100
rect 16260 1050 16270 1070
rect 16290 1050 16300 1070
rect 16260 1020 16300 1050
rect 16260 1000 16270 1020
rect 16290 1000 16300 1020
rect 16260 970 16300 1000
rect 16260 950 16270 970
rect 16290 950 16300 970
rect 16260 935 16300 950
rect 16315 1170 16355 1185
rect 16315 1150 16325 1170
rect 16345 1150 16355 1170
rect 16315 1120 16355 1150
rect 16315 1100 16325 1120
rect 16345 1100 16355 1120
rect 16315 1070 16355 1100
rect 16315 1050 16325 1070
rect 16345 1050 16355 1070
rect 16315 1020 16355 1050
rect 16315 1000 16325 1020
rect 16345 1000 16355 1020
rect 16315 970 16355 1000
rect 16315 950 16325 970
rect 16345 950 16355 970
rect 16315 935 16355 950
rect 16370 1170 16410 1185
rect 16370 1150 16380 1170
rect 16400 1150 16410 1170
rect 16370 1120 16410 1150
rect 16370 1100 16380 1120
rect 16400 1100 16410 1120
rect 16370 1070 16410 1100
rect 16370 1050 16380 1070
rect 16400 1050 16410 1070
rect 16370 1020 16410 1050
rect 16370 1000 16380 1020
rect 16400 1000 16410 1020
rect 16370 970 16410 1000
rect 16370 950 16380 970
rect 16400 950 16410 970
rect 16370 935 16410 950
rect 16425 1170 16465 1185
rect 16425 1150 16435 1170
rect 16455 1150 16465 1170
rect 16425 1120 16465 1150
rect 16425 1100 16435 1120
rect 16455 1100 16465 1120
rect 16425 1070 16465 1100
rect 16425 1050 16435 1070
rect 16455 1050 16465 1070
rect 16425 1020 16465 1050
rect 16425 1000 16435 1020
rect 16455 1000 16465 1020
rect 16425 970 16465 1000
rect 16425 950 16435 970
rect 16455 950 16465 970
rect 16425 935 16465 950
rect 16480 1170 16520 1185
rect 16480 1150 16490 1170
rect 16510 1150 16520 1170
rect 16480 1120 16520 1150
rect 16480 1100 16490 1120
rect 16510 1100 16520 1120
rect 16480 1070 16520 1100
rect 16480 1050 16490 1070
rect 16510 1050 16520 1070
rect 16480 1020 16520 1050
rect 16480 1000 16490 1020
rect 16510 1000 16520 1020
rect 16480 970 16520 1000
rect 16480 950 16490 970
rect 16510 950 16520 970
rect 16480 935 16520 950
rect 16535 1170 16575 1185
rect 16535 1150 16545 1170
rect 16565 1150 16575 1170
rect 16535 1120 16575 1150
rect 16535 1100 16545 1120
rect 16565 1100 16575 1120
rect 16535 1070 16575 1100
rect 16535 1050 16545 1070
rect 16565 1050 16575 1070
rect 16535 1020 16575 1050
rect 16535 1000 16545 1020
rect 16565 1000 16575 1020
rect 16535 970 16575 1000
rect 16535 950 16545 970
rect 16565 950 16575 970
rect 16535 935 16575 950
rect 16590 1170 16630 1185
rect 16590 1150 16600 1170
rect 16620 1150 16630 1170
rect 16590 1120 16630 1150
rect 16590 1100 16600 1120
rect 16620 1100 16630 1120
rect 16590 1070 16630 1100
rect 16590 1050 16600 1070
rect 16620 1050 16630 1070
rect 16590 1020 16630 1050
rect 16590 1000 16600 1020
rect 16620 1000 16630 1020
rect 16590 970 16630 1000
rect 16590 950 16600 970
rect 16620 950 16630 970
rect 16590 935 16630 950
rect 16645 1170 16685 1185
rect 16645 1150 16655 1170
rect 16675 1150 16685 1170
rect 16645 1120 16685 1150
rect 16645 1100 16655 1120
rect 16675 1100 16685 1120
rect 16645 1070 16685 1100
rect 16645 1050 16655 1070
rect 16675 1050 16685 1070
rect 16645 1020 16685 1050
rect 16645 1000 16655 1020
rect 16675 1000 16685 1020
rect 16645 970 16685 1000
rect 16645 950 16655 970
rect 16675 950 16685 970
rect 16645 935 16685 950
rect 16700 1170 16740 1185
rect 16700 1150 16710 1170
rect 16730 1150 16740 1170
rect 16700 1120 16740 1150
rect 16700 1100 16710 1120
rect 16730 1100 16740 1120
rect 16700 1070 16740 1100
rect 16700 1050 16710 1070
rect 16730 1050 16740 1070
rect 16700 1020 16740 1050
rect 16700 1000 16710 1020
rect 16730 1000 16740 1020
rect 16700 970 16740 1000
rect 16700 950 16710 970
rect 16730 950 16740 970
rect 16700 935 16740 950
rect 16755 1170 16795 1185
rect 16755 1150 16765 1170
rect 16785 1150 16795 1170
rect 16755 1120 16795 1150
rect 16755 1100 16765 1120
rect 16785 1100 16795 1120
rect 16755 1070 16795 1100
rect 16755 1050 16765 1070
rect 16785 1050 16795 1070
rect 16755 1020 16795 1050
rect 16755 1000 16765 1020
rect 16785 1000 16795 1020
rect 16755 970 16795 1000
rect 16755 950 16765 970
rect 16785 950 16795 970
rect 16755 935 16795 950
rect 16810 1170 16850 1185
rect 16810 1150 16820 1170
rect 16840 1150 16850 1170
rect 16810 1120 16850 1150
rect 16810 1100 16820 1120
rect 16840 1100 16850 1120
rect 16810 1070 16850 1100
rect 16810 1050 16820 1070
rect 16840 1050 16850 1070
rect 16810 1020 16850 1050
rect 16810 1000 16820 1020
rect 16840 1000 16850 1020
rect 16810 970 16850 1000
rect 16810 950 16820 970
rect 16840 950 16850 970
rect 16810 935 16850 950
rect 16865 1170 16905 1185
rect 16865 1150 16875 1170
rect 16895 1150 16905 1170
rect 16865 1120 16905 1150
rect 16865 1100 16875 1120
rect 16895 1100 16905 1120
rect 16865 1070 16905 1100
rect 16865 1050 16875 1070
rect 16895 1050 16905 1070
rect 16865 1020 16905 1050
rect 16865 1000 16875 1020
rect 16895 1000 16905 1020
rect 16865 970 16905 1000
rect 16865 950 16875 970
rect 16895 950 16905 970
rect 16865 935 16905 950
rect 16920 1170 16960 1185
rect 16920 1150 16930 1170
rect 16950 1150 16960 1170
rect 16920 1120 16960 1150
rect 16920 1100 16930 1120
rect 16950 1100 16960 1120
rect 16920 1070 16960 1100
rect 16920 1050 16930 1070
rect 16950 1050 16960 1070
rect 16920 1020 16960 1050
rect 16920 1000 16930 1020
rect 16950 1000 16960 1020
rect 16920 970 16960 1000
rect 16920 950 16930 970
rect 16950 950 16960 970
rect 16920 935 16960 950
rect 16975 1170 17015 1185
rect 16975 1150 16985 1170
rect 17005 1150 17015 1170
rect 16975 1120 17015 1150
rect 16975 1100 16985 1120
rect 17005 1100 17015 1120
rect 16975 1070 17015 1100
rect 16975 1050 16985 1070
rect 17005 1050 17015 1070
rect 16975 1020 17015 1050
rect 16975 1000 16985 1020
rect 17005 1000 17015 1020
rect 16975 970 17015 1000
rect 16975 950 16985 970
rect 17005 950 17015 970
rect 16975 935 17015 950
rect 17030 1170 17070 1185
rect 17030 1150 17040 1170
rect 17060 1150 17070 1170
rect 17030 1120 17070 1150
rect 17030 1100 17040 1120
rect 17060 1100 17070 1120
rect 17030 1070 17070 1100
rect 17030 1050 17040 1070
rect 17060 1050 17070 1070
rect 17030 1020 17070 1050
rect 17030 1000 17040 1020
rect 17060 1000 17070 1020
rect 17030 970 17070 1000
rect 17030 950 17040 970
rect 17060 950 17070 970
rect 17030 935 17070 950
rect 17085 1170 17125 1185
rect 17085 1150 17095 1170
rect 17115 1150 17125 1170
rect 17085 1120 17125 1150
rect 17085 1100 17095 1120
rect 17115 1100 17125 1120
rect 17085 1070 17125 1100
rect 17085 1050 17095 1070
rect 17115 1050 17125 1070
rect 17085 1020 17125 1050
rect 17085 1000 17095 1020
rect 17115 1000 17125 1020
rect 17085 970 17125 1000
rect 17085 950 17095 970
rect 17115 950 17125 970
rect 17085 935 17125 950
rect 17140 1170 17180 1185
rect 17140 1150 17150 1170
rect 17170 1150 17180 1170
rect 17140 1120 17180 1150
rect 17140 1100 17150 1120
rect 17170 1100 17180 1120
rect 17140 1070 17180 1100
rect 17140 1050 17150 1070
rect 17170 1050 17180 1070
rect 17140 1020 17180 1050
rect 17140 1000 17150 1020
rect 17170 1000 17180 1020
rect 17140 970 17180 1000
rect 17140 950 17150 970
rect 17170 950 17180 970
rect 17140 935 17180 950
rect 17195 1170 17235 1185
rect 17195 1150 17205 1170
rect 17225 1150 17235 1170
rect 17195 1120 17235 1150
rect 17195 1100 17205 1120
rect 17225 1100 17235 1120
rect 17195 1070 17235 1100
rect 17195 1050 17205 1070
rect 17225 1050 17235 1070
rect 17195 1020 17235 1050
rect 17195 1000 17205 1020
rect 17225 1000 17235 1020
rect 17195 970 17235 1000
rect 17195 950 17205 970
rect 17225 950 17235 970
rect 17195 935 17235 950
rect 17250 1170 17290 1185
rect 17250 1150 17260 1170
rect 17280 1150 17290 1170
rect 17250 1120 17290 1150
rect 17250 1100 17260 1120
rect 17280 1100 17290 1120
rect 17250 1070 17290 1100
rect 17250 1050 17260 1070
rect 17280 1050 17290 1070
rect 17250 1020 17290 1050
rect 17250 1000 17260 1020
rect 17280 1000 17290 1020
rect 17250 970 17290 1000
rect 17250 950 17260 970
rect 17280 950 17290 970
rect 17250 935 17290 950
rect 17305 1170 17345 1185
rect 17305 1150 17315 1170
rect 17335 1150 17345 1170
rect 17305 1120 17345 1150
rect 17305 1100 17315 1120
rect 17335 1100 17345 1120
rect 17305 1070 17345 1100
rect 17305 1050 17315 1070
rect 17335 1050 17345 1070
rect 17305 1020 17345 1050
rect 17305 1000 17315 1020
rect 17335 1000 17345 1020
rect 17305 970 17345 1000
rect 17305 950 17315 970
rect 17335 950 17345 970
rect 17305 935 17345 950
rect 17360 1170 17400 1185
rect 17360 1150 17370 1170
rect 17390 1150 17400 1170
rect 17360 1120 17400 1150
rect 17360 1100 17370 1120
rect 17390 1100 17400 1120
rect 17360 1070 17400 1100
rect 17360 1050 17370 1070
rect 17390 1050 17400 1070
rect 17360 1020 17400 1050
rect 17360 1000 17370 1020
rect 17390 1000 17400 1020
rect 17360 970 17400 1000
rect 17360 950 17370 970
rect 17390 950 17400 970
rect 17360 935 17400 950
rect 17415 1170 17455 1185
rect 17415 1150 17425 1170
rect 17445 1150 17455 1170
rect 17415 1120 17455 1150
rect 17415 1100 17425 1120
rect 17445 1100 17455 1120
rect 17415 1070 17455 1100
rect 17415 1050 17425 1070
rect 17445 1050 17455 1070
rect 17415 1020 17455 1050
rect 17415 1000 17425 1020
rect 17445 1000 17455 1020
rect 17415 970 17455 1000
rect 17415 950 17425 970
rect 17445 950 17455 970
rect 17415 935 17455 950
rect 17470 1170 17510 1185
rect 17470 1150 17480 1170
rect 17500 1150 17510 1170
rect 17470 1120 17510 1150
rect 17470 1100 17480 1120
rect 17500 1100 17510 1120
rect 17470 1070 17510 1100
rect 17470 1050 17480 1070
rect 17500 1050 17510 1070
rect 17470 1020 17510 1050
rect 17470 1000 17480 1020
rect 17500 1000 17510 1020
rect 17470 970 17510 1000
rect 17470 950 17480 970
rect 17500 950 17510 970
rect 17470 935 17510 950
rect 17525 1170 17565 1185
rect 17525 1150 17535 1170
rect 17555 1150 17565 1170
rect 17525 1120 17565 1150
rect 17525 1100 17535 1120
rect 17555 1100 17565 1120
rect 17525 1070 17565 1100
rect 17525 1050 17535 1070
rect 17555 1050 17565 1070
rect 17525 1020 17565 1050
rect 17525 1000 17535 1020
rect 17555 1000 17565 1020
rect 17525 970 17565 1000
rect 17525 950 17535 970
rect 17555 950 17565 970
rect 17525 935 17565 950
rect 17580 1170 17620 1185
rect 17580 1150 17590 1170
rect 17610 1150 17620 1170
rect 17580 1120 17620 1150
rect 17580 1100 17590 1120
rect 17610 1100 17620 1120
rect 17580 1070 17620 1100
rect 17580 1050 17590 1070
rect 17610 1050 17620 1070
rect 17580 1020 17620 1050
rect 17580 1000 17590 1020
rect 17610 1000 17620 1020
rect 17580 970 17620 1000
rect 17580 950 17590 970
rect 17610 950 17620 970
rect 18005 1170 18015 1190
rect 18035 1170 18045 1190
rect 18005 1140 18045 1170
rect 18005 1120 18015 1140
rect 18035 1120 18045 1140
rect 18005 1090 18045 1120
rect 18005 1070 18015 1090
rect 18035 1070 18045 1090
rect 18005 1040 18045 1070
rect 18005 1020 18015 1040
rect 18035 1020 18045 1040
rect 18005 990 18045 1020
rect 18005 970 18015 990
rect 18035 970 18045 990
rect 18005 955 18045 970
rect 18105 1640 18145 1655
rect 18105 1620 18115 1640
rect 18135 1620 18145 1640
rect 18105 1590 18145 1620
rect 18105 1570 18115 1590
rect 18135 1570 18145 1590
rect 18105 1540 18145 1570
rect 18105 1520 18115 1540
rect 18135 1520 18145 1540
rect 18105 1490 18145 1520
rect 18105 1470 18115 1490
rect 18135 1470 18145 1490
rect 18105 1440 18145 1470
rect 18105 1420 18115 1440
rect 18135 1420 18145 1440
rect 18105 1390 18145 1420
rect 18105 1370 18115 1390
rect 18135 1370 18145 1390
rect 18105 1340 18145 1370
rect 18105 1320 18115 1340
rect 18135 1320 18145 1340
rect 18105 1290 18145 1320
rect 18105 1270 18115 1290
rect 18135 1270 18145 1290
rect 18105 1240 18145 1270
rect 18105 1220 18115 1240
rect 18135 1220 18145 1240
rect 18105 1190 18145 1220
rect 18105 1170 18115 1190
rect 18135 1170 18145 1190
rect 18105 1140 18145 1170
rect 18105 1120 18115 1140
rect 18135 1120 18145 1140
rect 18105 1090 18145 1120
rect 18105 1070 18115 1090
rect 18135 1070 18145 1090
rect 18105 1040 18145 1070
rect 18105 1020 18115 1040
rect 18135 1020 18145 1040
rect 18105 990 18145 1020
rect 18105 970 18115 990
rect 18135 970 18145 990
rect 18105 955 18145 970
rect 18205 1640 18245 1655
rect 18205 1620 18215 1640
rect 18235 1620 18245 1640
rect 18205 1590 18245 1620
rect 18205 1570 18215 1590
rect 18235 1570 18245 1590
rect 18205 1540 18245 1570
rect 18205 1520 18215 1540
rect 18235 1520 18245 1540
rect 18205 1490 18245 1520
rect 18205 1470 18215 1490
rect 18235 1470 18245 1490
rect 18205 1440 18245 1470
rect 18205 1420 18215 1440
rect 18235 1420 18245 1440
rect 18205 1390 18245 1420
rect 18205 1370 18215 1390
rect 18235 1370 18245 1390
rect 18205 1340 18245 1370
rect 18205 1320 18215 1340
rect 18235 1320 18245 1340
rect 18205 1290 18245 1320
rect 18205 1270 18215 1290
rect 18235 1270 18245 1290
rect 18205 1240 18245 1270
rect 18205 1220 18215 1240
rect 18235 1220 18245 1240
rect 18205 1190 18245 1220
rect 18205 1170 18215 1190
rect 18235 1170 18245 1190
rect 18205 1140 18245 1170
rect 18205 1120 18215 1140
rect 18235 1120 18245 1140
rect 18205 1090 18245 1120
rect 18205 1070 18215 1090
rect 18235 1070 18245 1090
rect 18205 1040 18245 1070
rect 18205 1020 18215 1040
rect 18235 1020 18245 1040
rect 18205 990 18245 1020
rect 18205 970 18215 990
rect 18235 970 18245 990
rect 18205 955 18245 970
rect 18305 1640 18345 1655
rect 18305 1620 18315 1640
rect 18335 1620 18345 1640
rect 18305 1590 18345 1620
rect 18305 1570 18315 1590
rect 18335 1570 18345 1590
rect 18305 1540 18345 1570
rect 18305 1520 18315 1540
rect 18335 1520 18345 1540
rect 18305 1490 18345 1520
rect 18305 1470 18315 1490
rect 18335 1470 18345 1490
rect 18305 1440 18345 1470
rect 18305 1420 18315 1440
rect 18335 1420 18345 1440
rect 18305 1390 18345 1420
rect 18305 1370 18315 1390
rect 18335 1370 18345 1390
rect 18305 1340 18345 1370
rect 18305 1320 18315 1340
rect 18335 1320 18345 1340
rect 18305 1290 18345 1320
rect 18305 1270 18315 1290
rect 18335 1270 18345 1290
rect 18305 1240 18345 1270
rect 18305 1220 18315 1240
rect 18335 1220 18345 1240
rect 18305 1190 18345 1220
rect 18305 1170 18315 1190
rect 18335 1170 18345 1190
rect 18305 1140 18345 1170
rect 18305 1120 18315 1140
rect 18335 1120 18345 1140
rect 18305 1090 18345 1120
rect 18305 1070 18315 1090
rect 18335 1070 18345 1090
rect 18305 1040 18345 1070
rect 18305 1020 18315 1040
rect 18335 1020 18345 1040
rect 18305 990 18345 1020
rect 18305 970 18315 990
rect 18335 970 18345 990
rect 18305 955 18345 970
rect 18405 1640 18445 1655
rect 18405 1620 18415 1640
rect 18435 1620 18445 1640
rect 18405 1590 18445 1620
rect 18405 1570 18415 1590
rect 18435 1570 18445 1590
rect 18405 1540 18445 1570
rect 18405 1520 18415 1540
rect 18435 1520 18445 1540
rect 18405 1490 18445 1520
rect 18405 1470 18415 1490
rect 18435 1470 18445 1490
rect 18405 1440 18445 1470
rect 18405 1420 18415 1440
rect 18435 1420 18445 1440
rect 18405 1390 18445 1420
rect 18405 1370 18415 1390
rect 18435 1370 18445 1390
rect 18405 1340 18445 1370
rect 18405 1320 18415 1340
rect 18435 1320 18445 1340
rect 18405 1290 18445 1320
rect 18405 1270 18415 1290
rect 18435 1270 18445 1290
rect 18405 1240 18445 1270
rect 18405 1220 18415 1240
rect 18435 1220 18445 1240
rect 18405 1190 18445 1220
rect 18405 1170 18415 1190
rect 18435 1170 18445 1190
rect 18405 1140 18445 1170
rect 18405 1120 18415 1140
rect 18435 1120 18445 1140
rect 18405 1090 18445 1120
rect 18405 1070 18415 1090
rect 18435 1070 18445 1090
rect 18405 1040 18445 1070
rect 18405 1020 18415 1040
rect 18435 1020 18445 1040
rect 18405 990 18445 1020
rect 18405 970 18415 990
rect 18435 970 18445 990
rect 18405 955 18445 970
rect 18505 1640 18545 1655
rect 18505 1620 18515 1640
rect 18535 1620 18545 1640
rect 18505 1590 18545 1620
rect 18505 1570 18515 1590
rect 18535 1570 18545 1590
rect 18505 1540 18545 1570
rect 18505 1520 18515 1540
rect 18535 1520 18545 1540
rect 18505 1490 18545 1520
rect 18505 1470 18515 1490
rect 18535 1470 18545 1490
rect 18505 1440 18545 1470
rect 18505 1420 18515 1440
rect 18535 1420 18545 1440
rect 18505 1390 18545 1420
rect 18505 1370 18515 1390
rect 18535 1370 18545 1390
rect 18505 1340 18545 1370
rect 18505 1320 18515 1340
rect 18535 1320 18545 1340
rect 18505 1290 18545 1320
rect 18505 1270 18515 1290
rect 18535 1270 18545 1290
rect 18505 1240 18545 1270
rect 18505 1220 18515 1240
rect 18535 1220 18545 1240
rect 18505 1190 18545 1220
rect 18505 1170 18515 1190
rect 18535 1170 18545 1190
rect 18505 1140 18545 1170
rect 18505 1120 18515 1140
rect 18535 1120 18545 1140
rect 18505 1090 18545 1120
rect 18505 1070 18515 1090
rect 18535 1070 18545 1090
rect 18505 1040 18545 1070
rect 18505 1020 18515 1040
rect 18535 1020 18545 1040
rect 18505 990 18545 1020
rect 18505 970 18515 990
rect 18535 970 18545 990
rect 18505 955 18545 970
rect 18605 1640 18645 1655
rect 18605 1620 18615 1640
rect 18635 1620 18645 1640
rect 18605 1590 18645 1620
rect 18605 1570 18615 1590
rect 18635 1570 18645 1590
rect 18605 1540 18645 1570
rect 18605 1520 18615 1540
rect 18635 1520 18645 1540
rect 18605 1490 18645 1520
rect 18605 1470 18615 1490
rect 18635 1470 18645 1490
rect 18605 1440 18645 1470
rect 18605 1420 18615 1440
rect 18635 1420 18645 1440
rect 18605 1390 18645 1420
rect 18605 1370 18615 1390
rect 18635 1370 18645 1390
rect 18605 1340 18645 1370
rect 18605 1320 18615 1340
rect 18635 1320 18645 1340
rect 18605 1290 18645 1320
rect 18605 1270 18615 1290
rect 18635 1270 18645 1290
rect 18605 1240 18645 1270
rect 18605 1220 18615 1240
rect 18635 1220 18645 1240
rect 18605 1190 18645 1220
rect 18605 1170 18615 1190
rect 18635 1170 18645 1190
rect 18605 1140 18645 1170
rect 18605 1120 18615 1140
rect 18635 1120 18645 1140
rect 18605 1090 18645 1120
rect 18605 1070 18615 1090
rect 18635 1070 18645 1090
rect 18605 1040 18645 1070
rect 18605 1020 18615 1040
rect 18635 1020 18645 1040
rect 18605 990 18645 1020
rect 18605 970 18615 990
rect 18635 970 18645 990
rect 18605 955 18645 970
rect 17580 935 17620 950
rect 2995 865 3035 880
rect 2995 845 3005 865
rect 3025 845 3035 865
rect 2995 815 3035 845
rect 2995 795 3005 815
rect 3025 795 3035 815
rect 2995 780 3035 795
rect 3085 865 3125 880
rect 3085 845 3095 865
rect 3115 845 3125 865
rect 3085 815 3125 845
rect 3085 795 3095 815
rect 3115 795 3125 815
rect 3085 780 3125 795
rect 3175 865 3215 880
rect 3175 845 3185 865
rect 3205 845 3215 865
rect 3175 815 3215 845
rect 3175 795 3185 815
rect 3205 795 3215 815
rect 3175 780 3215 795
rect 3265 865 3305 880
rect 3265 845 3275 865
rect 3295 845 3305 865
rect 3265 815 3305 845
rect 3265 795 3275 815
rect 3295 795 3305 815
rect 3265 780 3305 795
rect 3355 865 3395 880
rect 3355 845 3365 865
rect 3385 845 3395 865
rect 3355 815 3395 845
rect 3355 795 3365 815
rect 3385 795 3395 815
rect 3355 780 3395 795
rect 3445 865 3485 880
rect 3445 845 3455 865
rect 3475 845 3485 865
rect 3445 815 3485 845
rect 3445 795 3455 815
rect 3475 795 3485 815
rect 3445 780 3485 795
rect 3535 865 3575 880
rect 3535 845 3545 865
rect 3565 845 3575 865
rect 3535 815 3575 845
rect 3535 795 3545 815
rect 3565 795 3575 815
rect 3535 780 3575 795
rect 3625 865 3665 880
rect 3625 845 3635 865
rect 3655 845 3665 865
rect 3625 815 3665 845
rect 3625 795 3635 815
rect 3655 795 3665 815
rect 3625 780 3665 795
rect 3715 865 3755 880
rect 3715 845 3725 865
rect 3745 845 3755 865
rect 3715 815 3755 845
rect 3715 795 3725 815
rect 3745 795 3755 815
rect 3715 780 3755 795
rect 3805 865 3845 880
rect 3805 845 3815 865
rect 3835 845 3845 865
rect 3805 815 3845 845
rect 3805 795 3815 815
rect 3835 795 3845 815
rect 3805 780 3845 795
rect 3895 865 3935 880
rect 3895 845 3905 865
rect 3925 845 3935 865
rect 3895 815 3935 845
rect 3895 795 3905 815
rect 3925 795 3935 815
rect 3895 780 3935 795
rect 3985 865 4025 880
rect 3985 845 3995 865
rect 4015 845 4025 865
rect 3985 815 4025 845
rect 3985 795 3995 815
rect 4015 795 4025 815
rect 3985 780 4025 795
rect 4075 865 4115 880
rect 4075 845 4085 865
rect 4105 845 4115 865
rect 4075 815 4115 845
rect 4075 795 4085 815
rect 4105 795 4115 815
rect 4075 780 4115 795
rect 4165 865 4205 880
rect 4165 845 4175 865
rect 4195 845 4205 865
rect 4165 815 4205 845
rect 4165 795 4175 815
rect 4195 795 4205 815
rect 4165 780 4205 795
rect 4255 865 4295 880
rect 4255 845 4265 865
rect 4285 845 4295 865
rect 4255 815 4295 845
rect 4255 795 4265 815
rect 4285 795 4295 815
rect 4255 780 4295 795
rect 4345 865 4385 880
rect 4345 845 4355 865
rect 4375 845 4385 865
rect 4345 815 4385 845
rect 4345 795 4355 815
rect 4375 795 4385 815
rect 4345 780 4385 795
rect 4435 865 4475 880
rect 4435 845 4445 865
rect 4465 845 4475 865
rect 4435 815 4475 845
rect 4435 795 4445 815
rect 4465 795 4475 815
rect 4435 780 4475 795
rect 4525 865 4565 880
rect 4525 845 4535 865
rect 4555 845 4565 865
rect 4525 815 4565 845
rect 4525 795 4535 815
rect 4555 795 4565 815
rect 4525 780 4565 795
rect 4615 865 4655 880
rect 4615 845 4625 865
rect 4645 845 4655 865
rect 4615 815 4655 845
rect 4615 795 4625 815
rect 4645 795 4655 815
rect 4615 780 4655 795
rect 4705 865 4745 880
rect 4705 845 4715 865
rect 4735 845 4745 865
rect 4705 815 4745 845
rect 4705 795 4715 815
rect 4735 795 4745 815
rect 4705 780 4745 795
rect 4795 865 4835 880
rect 4795 845 4805 865
rect 4825 845 4835 865
rect 4795 815 4835 845
rect 4795 795 4805 815
rect 4825 795 4835 815
rect 4795 780 4835 795
rect 4885 865 4925 880
rect 4885 845 4895 865
rect 4915 845 4925 865
rect 4885 815 4925 845
rect 4885 795 4895 815
rect 4915 795 4925 815
rect 4885 780 4925 795
rect 4975 865 5015 880
rect 4975 845 4985 865
rect 5005 845 5015 865
rect 4975 815 5015 845
rect 4975 795 4985 815
rect 5005 795 5015 815
rect 4975 780 5015 795
rect 16260 730 16300 745
rect 16260 710 16270 730
rect 16290 710 16300 730
rect 16260 680 16300 710
rect 16260 660 16270 680
rect 16290 660 16300 680
rect 16260 645 16300 660
rect 16490 730 16530 745
rect 16490 710 16500 730
rect 16520 710 16530 730
rect 16490 680 16530 710
rect 16880 735 16920 750
rect 16880 715 16890 735
rect 16910 715 16920 735
rect 16880 700 16920 715
rect 16935 735 16975 750
rect 16935 715 16945 735
rect 16965 715 16975 735
rect 16935 700 16975 715
rect 16990 735 17030 750
rect 16990 715 17000 735
rect 17020 715 17030 735
rect 16990 700 17030 715
rect 17045 735 17085 750
rect 17045 715 17055 735
rect 17075 715 17085 735
rect 17045 700 17085 715
rect 17100 735 17140 750
rect 17100 715 17110 735
rect 17130 715 17140 735
rect 17100 700 17140 715
rect 17155 735 17195 750
rect 17155 715 17165 735
rect 17185 715 17195 735
rect 17155 700 17195 715
rect 17210 735 17250 750
rect 17210 715 17220 735
rect 17240 715 17250 735
rect 17210 700 17250 715
rect 17265 735 17305 750
rect 17265 715 17275 735
rect 17295 715 17305 735
rect 17265 700 17305 715
rect 17320 735 17360 750
rect 17320 715 17330 735
rect 17350 715 17360 735
rect 17320 700 17360 715
rect 17375 735 17415 750
rect 17375 715 17385 735
rect 17405 715 17415 735
rect 17375 700 17415 715
rect 17430 735 17470 750
rect 17430 715 17440 735
rect 17460 715 17470 735
rect 17430 700 17470 715
rect 17485 735 17525 750
rect 17485 715 17495 735
rect 17515 715 17525 735
rect 17485 700 17525 715
rect 17540 735 17580 750
rect 17540 715 17550 735
rect 17570 715 17580 735
rect 17540 700 17580 715
rect 16490 660 16500 680
rect 16520 660 16530 680
rect 16490 645 16530 660
<< pdiff >>
rect 2995 2915 3035 2930
rect 2995 2895 3005 2915
rect 3025 2895 3035 2915
rect 2995 2865 3035 2895
rect 2995 2845 3005 2865
rect 3025 2845 3035 2865
rect 2995 2830 3035 2845
rect 3085 2915 3125 2930
rect 3085 2895 3095 2915
rect 3115 2895 3125 2915
rect 3085 2865 3125 2895
rect 3085 2845 3095 2865
rect 3115 2845 3125 2865
rect 3085 2830 3125 2845
rect 3175 2915 3215 2930
rect 3175 2895 3185 2915
rect 3205 2895 3215 2915
rect 3175 2865 3215 2895
rect 3175 2845 3185 2865
rect 3205 2845 3215 2865
rect 3175 2830 3215 2845
rect 3265 2915 3305 2930
rect 3265 2895 3275 2915
rect 3295 2895 3305 2915
rect 3265 2865 3305 2895
rect 3265 2845 3275 2865
rect 3295 2845 3305 2865
rect 3265 2830 3305 2845
rect 3355 2915 3395 2930
rect 3355 2895 3365 2915
rect 3385 2895 3395 2915
rect 3355 2865 3395 2895
rect 3355 2845 3365 2865
rect 3385 2845 3395 2865
rect 3355 2830 3395 2845
rect 3445 2915 3485 2930
rect 3445 2895 3455 2915
rect 3475 2895 3485 2915
rect 3445 2865 3485 2895
rect 3445 2845 3455 2865
rect 3475 2845 3485 2865
rect 3445 2830 3485 2845
rect 3535 2915 3575 2930
rect 3535 2895 3545 2915
rect 3565 2895 3575 2915
rect 3535 2865 3575 2895
rect 3535 2845 3545 2865
rect 3565 2845 3575 2865
rect 3535 2830 3575 2845
rect 3625 2915 3665 2930
rect 3625 2895 3635 2915
rect 3655 2895 3665 2915
rect 3625 2865 3665 2895
rect 3625 2845 3635 2865
rect 3655 2845 3665 2865
rect 3625 2830 3665 2845
rect 3715 2915 3755 2930
rect 3715 2895 3725 2915
rect 3745 2895 3755 2915
rect 3715 2865 3755 2895
rect 3715 2845 3725 2865
rect 3745 2845 3755 2865
rect 3715 2830 3755 2845
rect 3805 2915 3845 2930
rect 3805 2895 3815 2915
rect 3835 2895 3845 2915
rect 3805 2865 3845 2895
rect 3805 2845 3815 2865
rect 3835 2845 3845 2865
rect 3805 2830 3845 2845
rect 3895 2915 3935 2930
rect 3895 2895 3905 2915
rect 3925 2895 3935 2915
rect 3895 2865 3935 2895
rect 3895 2845 3905 2865
rect 3925 2845 3935 2865
rect 3895 2830 3935 2845
rect 3985 2915 4025 2930
rect 3985 2895 3995 2915
rect 4015 2895 4025 2915
rect 3985 2865 4025 2895
rect 3985 2845 3995 2865
rect 4015 2845 4025 2865
rect 3985 2830 4025 2845
rect 4075 2915 4115 2930
rect 4075 2895 4085 2915
rect 4105 2895 4115 2915
rect 4075 2865 4115 2895
rect 4075 2845 4085 2865
rect 4105 2845 4115 2865
rect 4075 2830 4115 2845
rect 4165 2915 4205 2930
rect 4165 2895 4175 2915
rect 4195 2895 4205 2915
rect 4165 2865 4205 2895
rect 4165 2845 4175 2865
rect 4195 2845 4205 2865
rect 4165 2830 4205 2845
rect 4255 2915 4295 2930
rect 4255 2895 4265 2915
rect 4285 2895 4295 2915
rect 4255 2865 4295 2895
rect 4255 2845 4265 2865
rect 4285 2845 4295 2865
rect 4255 2830 4295 2845
rect 4345 2915 4385 2930
rect 4345 2895 4355 2915
rect 4375 2895 4385 2915
rect 4345 2865 4385 2895
rect 4345 2845 4355 2865
rect 4375 2845 4385 2865
rect 4345 2830 4385 2845
rect 4435 2915 4475 2930
rect 4435 2895 4445 2915
rect 4465 2895 4475 2915
rect 4435 2865 4475 2895
rect 4435 2845 4445 2865
rect 4465 2845 4475 2865
rect 4435 2830 4475 2845
rect 4525 2915 4565 2930
rect 4525 2895 4535 2915
rect 4555 2895 4565 2915
rect 4525 2865 4565 2895
rect 4525 2845 4535 2865
rect 4555 2845 4565 2865
rect 4525 2830 4565 2845
rect 4615 2915 4655 2930
rect 4615 2895 4625 2915
rect 4645 2895 4655 2915
rect 4615 2865 4655 2895
rect 4615 2845 4625 2865
rect 4645 2845 4655 2865
rect 4615 2830 4655 2845
rect 4705 2915 4745 2930
rect 4705 2895 4715 2915
rect 4735 2895 4745 2915
rect 4705 2865 4745 2895
rect 4705 2845 4715 2865
rect 4735 2845 4745 2865
rect 4705 2830 4745 2845
rect 4795 2915 4835 2930
rect 4795 2895 4805 2915
rect 4825 2895 4835 2915
rect 4795 2865 4835 2895
rect 4795 2845 4805 2865
rect 4825 2845 4835 2865
rect 4795 2830 4835 2845
rect 4885 2915 4925 2930
rect 4885 2895 4895 2915
rect 4915 2895 4925 2915
rect 4885 2865 4925 2895
rect 4885 2845 4895 2865
rect 4915 2845 4925 2865
rect 4885 2830 4925 2845
rect 4975 2915 5015 2930
rect 4975 2895 4985 2915
rect 5005 2895 5015 2915
rect 4975 2865 5015 2895
rect 4975 2845 4985 2865
rect 5005 2845 5015 2865
rect 4975 2830 5015 2845
rect 3175 2685 3215 2700
rect 3175 2665 3185 2685
rect 3205 2665 3215 2685
rect 3175 2635 3215 2665
rect 3175 2615 3185 2635
rect 3205 2615 3215 2635
rect 3175 2585 3215 2615
rect 3175 2565 3185 2585
rect 3205 2565 3215 2585
rect 3175 2535 3215 2565
rect 3175 2515 3185 2535
rect 3205 2515 3215 2535
rect 3175 2485 3215 2515
rect 3175 2465 3185 2485
rect 3205 2465 3215 2485
rect 3175 2435 3215 2465
rect 3175 2415 3185 2435
rect 3205 2415 3215 2435
rect 3175 2400 3215 2415
rect 3265 2685 3305 2700
rect 3265 2665 3275 2685
rect 3295 2665 3305 2685
rect 3265 2635 3305 2665
rect 3265 2615 3275 2635
rect 3295 2615 3305 2635
rect 3265 2585 3305 2615
rect 3265 2565 3275 2585
rect 3295 2565 3305 2585
rect 3265 2535 3305 2565
rect 3265 2515 3275 2535
rect 3295 2515 3305 2535
rect 3265 2485 3305 2515
rect 3265 2465 3275 2485
rect 3295 2465 3305 2485
rect 3265 2435 3305 2465
rect 3265 2415 3275 2435
rect 3295 2415 3305 2435
rect 3265 2400 3305 2415
rect 3355 2685 3395 2700
rect 3355 2665 3365 2685
rect 3385 2665 3395 2685
rect 3355 2635 3395 2665
rect 3355 2615 3365 2635
rect 3385 2615 3395 2635
rect 3355 2585 3395 2615
rect 3355 2565 3365 2585
rect 3385 2565 3395 2585
rect 3355 2535 3395 2565
rect 3355 2515 3365 2535
rect 3385 2515 3395 2535
rect 3355 2485 3395 2515
rect 3355 2465 3365 2485
rect 3385 2465 3395 2485
rect 3355 2435 3395 2465
rect 3355 2415 3365 2435
rect 3385 2415 3395 2435
rect 3355 2400 3395 2415
rect 3445 2685 3485 2700
rect 3445 2665 3455 2685
rect 3475 2665 3485 2685
rect 3445 2635 3485 2665
rect 3445 2615 3455 2635
rect 3475 2615 3485 2635
rect 3445 2585 3485 2615
rect 3445 2565 3455 2585
rect 3475 2565 3485 2585
rect 3445 2535 3485 2565
rect 3445 2515 3455 2535
rect 3475 2515 3485 2535
rect 3445 2485 3485 2515
rect 3445 2465 3455 2485
rect 3475 2465 3485 2485
rect 3445 2435 3485 2465
rect 3445 2415 3455 2435
rect 3475 2415 3485 2435
rect 3445 2400 3485 2415
rect 3535 2685 3575 2700
rect 3535 2665 3545 2685
rect 3565 2665 3575 2685
rect 3535 2635 3575 2665
rect 3535 2615 3545 2635
rect 3565 2615 3575 2635
rect 3535 2585 3575 2615
rect 3535 2565 3545 2585
rect 3565 2565 3575 2585
rect 3535 2535 3575 2565
rect 3535 2515 3545 2535
rect 3565 2515 3575 2535
rect 3535 2485 3575 2515
rect 3535 2465 3545 2485
rect 3565 2465 3575 2485
rect 3535 2435 3575 2465
rect 3535 2415 3545 2435
rect 3565 2415 3575 2435
rect 3535 2400 3575 2415
rect 3625 2685 3665 2700
rect 3625 2665 3635 2685
rect 3655 2665 3665 2685
rect 3625 2635 3665 2665
rect 3625 2615 3635 2635
rect 3655 2615 3665 2635
rect 3625 2585 3665 2615
rect 3625 2565 3635 2585
rect 3655 2565 3665 2585
rect 3625 2535 3665 2565
rect 3625 2515 3635 2535
rect 3655 2515 3665 2535
rect 3625 2485 3665 2515
rect 3625 2465 3635 2485
rect 3655 2465 3665 2485
rect 3625 2435 3665 2465
rect 3625 2415 3635 2435
rect 3655 2415 3665 2435
rect 3625 2400 3665 2415
rect 3715 2685 3755 2700
rect 3715 2665 3725 2685
rect 3745 2665 3755 2685
rect 3715 2635 3755 2665
rect 3715 2615 3725 2635
rect 3745 2615 3755 2635
rect 3715 2585 3755 2615
rect 3715 2565 3725 2585
rect 3745 2565 3755 2585
rect 3715 2535 3755 2565
rect 3715 2515 3725 2535
rect 3745 2515 3755 2535
rect 3715 2485 3755 2515
rect 3715 2465 3725 2485
rect 3745 2465 3755 2485
rect 3715 2435 3755 2465
rect 3715 2415 3725 2435
rect 3745 2415 3755 2435
rect 3715 2400 3755 2415
rect 3805 2685 3845 2700
rect 3805 2665 3815 2685
rect 3835 2665 3845 2685
rect 3805 2635 3845 2665
rect 3805 2615 3815 2635
rect 3835 2615 3845 2635
rect 3805 2585 3845 2615
rect 3805 2565 3815 2585
rect 3835 2565 3845 2585
rect 3805 2535 3845 2565
rect 3805 2515 3815 2535
rect 3835 2515 3845 2535
rect 3805 2485 3845 2515
rect 3805 2465 3815 2485
rect 3835 2465 3845 2485
rect 3805 2435 3845 2465
rect 3805 2415 3815 2435
rect 3835 2415 3845 2435
rect 3805 2400 3845 2415
rect 3895 2685 3935 2700
rect 3895 2665 3905 2685
rect 3925 2665 3935 2685
rect 3895 2635 3935 2665
rect 3895 2615 3905 2635
rect 3925 2615 3935 2635
rect 3895 2585 3935 2615
rect 3895 2565 3905 2585
rect 3925 2565 3935 2585
rect 3895 2535 3935 2565
rect 3895 2515 3905 2535
rect 3925 2515 3935 2535
rect 3895 2485 3935 2515
rect 3895 2465 3905 2485
rect 3925 2465 3935 2485
rect 3895 2435 3935 2465
rect 3895 2415 3905 2435
rect 3925 2415 3935 2435
rect 3895 2400 3935 2415
rect 3985 2685 4025 2700
rect 3985 2665 3995 2685
rect 4015 2665 4025 2685
rect 3985 2635 4025 2665
rect 3985 2615 3995 2635
rect 4015 2615 4025 2635
rect 3985 2585 4025 2615
rect 3985 2565 3995 2585
rect 4015 2565 4025 2585
rect 3985 2535 4025 2565
rect 3985 2515 3995 2535
rect 4015 2515 4025 2535
rect 3985 2485 4025 2515
rect 3985 2465 3995 2485
rect 4015 2465 4025 2485
rect 3985 2435 4025 2465
rect 3985 2415 3995 2435
rect 4015 2415 4025 2435
rect 3985 2400 4025 2415
rect 4075 2685 4115 2700
rect 4075 2665 4085 2685
rect 4105 2665 4115 2685
rect 4075 2635 4115 2665
rect 4075 2615 4085 2635
rect 4105 2615 4115 2635
rect 4075 2585 4115 2615
rect 4075 2565 4085 2585
rect 4105 2565 4115 2585
rect 4075 2535 4115 2565
rect 4075 2515 4085 2535
rect 4105 2515 4115 2535
rect 4075 2485 4115 2515
rect 4075 2465 4085 2485
rect 4105 2465 4115 2485
rect 4075 2435 4115 2465
rect 4075 2415 4085 2435
rect 4105 2415 4115 2435
rect 4075 2400 4115 2415
rect 4165 2685 4205 2700
rect 4165 2665 4175 2685
rect 4195 2665 4205 2685
rect 4165 2635 4205 2665
rect 4165 2615 4175 2635
rect 4195 2615 4205 2635
rect 4165 2585 4205 2615
rect 4165 2565 4175 2585
rect 4195 2565 4205 2585
rect 4165 2535 4205 2565
rect 4165 2515 4175 2535
rect 4195 2515 4205 2535
rect 4165 2485 4205 2515
rect 4165 2465 4175 2485
rect 4195 2465 4205 2485
rect 4165 2435 4205 2465
rect 4165 2415 4175 2435
rect 4195 2415 4205 2435
rect 4165 2400 4205 2415
rect 4255 2685 4295 2700
rect 4255 2665 4265 2685
rect 4285 2665 4295 2685
rect 4255 2635 4295 2665
rect 4255 2615 4265 2635
rect 4285 2615 4295 2635
rect 4255 2585 4295 2615
rect 4255 2565 4265 2585
rect 4285 2565 4295 2585
rect 4255 2535 4295 2565
rect 4255 2515 4265 2535
rect 4285 2515 4295 2535
rect 4255 2485 4295 2515
rect 4255 2465 4265 2485
rect 4285 2465 4295 2485
rect 4255 2435 4295 2465
rect 4255 2415 4265 2435
rect 4285 2415 4295 2435
rect 4255 2400 4295 2415
rect 4345 2685 4385 2700
rect 4345 2665 4355 2685
rect 4375 2665 4385 2685
rect 4345 2635 4385 2665
rect 4345 2615 4355 2635
rect 4375 2615 4385 2635
rect 4345 2585 4385 2615
rect 4345 2565 4355 2585
rect 4375 2565 4385 2585
rect 4345 2535 4385 2565
rect 4345 2515 4355 2535
rect 4375 2515 4385 2535
rect 4345 2485 4385 2515
rect 4345 2465 4355 2485
rect 4375 2465 4385 2485
rect 4345 2435 4385 2465
rect 4345 2415 4355 2435
rect 4375 2415 4385 2435
rect 4345 2400 4385 2415
rect 4435 2685 4475 2700
rect 4435 2665 4445 2685
rect 4465 2665 4475 2685
rect 4435 2635 4475 2665
rect 4435 2615 4445 2635
rect 4465 2615 4475 2635
rect 4435 2585 4475 2615
rect 4435 2565 4445 2585
rect 4465 2565 4475 2585
rect 4435 2535 4475 2565
rect 4435 2515 4445 2535
rect 4465 2515 4475 2535
rect 4435 2485 4475 2515
rect 4435 2465 4445 2485
rect 4465 2465 4475 2485
rect 4435 2435 4475 2465
rect 4435 2415 4445 2435
rect 4465 2415 4475 2435
rect 4435 2400 4475 2415
rect 4525 2685 4565 2700
rect 4525 2665 4535 2685
rect 4555 2665 4565 2685
rect 4525 2635 4565 2665
rect 4525 2615 4535 2635
rect 4555 2615 4565 2635
rect 4525 2585 4565 2615
rect 4525 2565 4535 2585
rect 4555 2565 4565 2585
rect 4525 2535 4565 2565
rect 4525 2515 4535 2535
rect 4555 2515 4565 2535
rect 4525 2485 4565 2515
rect 4525 2465 4535 2485
rect 4555 2465 4565 2485
rect 4525 2435 4565 2465
rect 4525 2415 4535 2435
rect 4555 2415 4565 2435
rect 4525 2400 4565 2415
rect 4615 2685 4655 2700
rect 4615 2665 4625 2685
rect 4645 2665 4655 2685
rect 4615 2635 4655 2665
rect 4615 2615 4625 2635
rect 4645 2615 4655 2635
rect 4615 2585 4655 2615
rect 4615 2565 4625 2585
rect 4645 2565 4655 2585
rect 4615 2535 4655 2565
rect 4615 2515 4625 2535
rect 4645 2515 4655 2535
rect 4615 2485 4655 2515
rect 4615 2465 4625 2485
rect 4645 2465 4655 2485
rect 4615 2435 4655 2465
rect 4615 2415 4625 2435
rect 4645 2415 4655 2435
rect 4615 2400 4655 2415
rect 4705 2685 4745 2700
rect 4705 2665 4715 2685
rect 4735 2665 4745 2685
rect 4705 2635 4745 2665
rect 4705 2615 4715 2635
rect 4735 2615 4745 2635
rect 4705 2585 4745 2615
rect 4705 2565 4715 2585
rect 4735 2565 4745 2585
rect 4705 2535 4745 2565
rect 4705 2515 4715 2535
rect 4735 2515 4745 2535
rect 4705 2485 4745 2515
rect 4705 2465 4715 2485
rect 4735 2465 4745 2485
rect 4705 2435 4745 2465
rect 4705 2415 4715 2435
rect 4735 2415 4745 2435
rect 4705 2400 4745 2415
rect 4795 2685 4835 2700
rect 4795 2665 4805 2685
rect 4825 2665 4835 2685
rect 4795 2635 4835 2665
rect 4795 2615 4805 2635
rect 4825 2615 4835 2635
rect 4795 2585 4835 2615
rect 4795 2565 4805 2585
rect 4825 2565 4835 2585
rect 4795 2535 4835 2565
rect 4795 2515 4805 2535
rect 4825 2515 4835 2535
rect 4795 2485 4835 2515
rect 4795 2465 4805 2485
rect 4825 2465 4835 2485
rect 4795 2435 4835 2465
rect 4795 2415 4805 2435
rect 4825 2415 4835 2435
rect 4795 2400 4835 2415
rect 2565 1985 2605 2000
rect 2565 1965 2575 1985
rect 2595 1965 2605 1985
rect 2565 1935 2605 1965
rect 2565 1915 2575 1935
rect 2595 1915 2605 1935
rect 2565 1900 2605 1915
rect 2620 1985 2660 2000
rect 2620 1965 2630 1985
rect 2650 1965 2660 1985
rect 2620 1935 2660 1965
rect 2620 1915 2630 1935
rect 2650 1915 2660 1935
rect 2620 1900 2660 1915
rect 2675 1985 2715 2000
rect 2675 1965 2685 1985
rect 2705 1965 2715 1985
rect 2675 1935 2715 1965
rect 2675 1915 2685 1935
rect 2705 1915 2715 1935
rect 2675 1900 2715 1915
rect 2745 1985 2785 2000
rect 2745 1965 2755 1985
rect 2775 1965 2785 1985
rect 2745 1935 2785 1965
rect 2745 1915 2755 1935
rect 2775 1915 2785 1935
rect 2745 1900 2785 1915
rect 2805 1985 2845 2000
rect 2805 1965 2815 1985
rect 2835 1965 2845 1985
rect 2805 1935 2845 1965
rect 2805 1915 2815 1935
rect 2835 1915 2845 1935
rect 2805 1900 2845 1915
rect 2865 1985 2905 2000
rect 2865 1965 2875 1985
rect 2895 1965 2905 1985
rect 2865 1935 2905 1965
rect 2865 1915 2875 1935
rect 2895 1915 2905 1935
rect 2865 1900 2905 1915
rect 2925 1985 2965 2000
rect 2925 1965 2935 1985
rect 2955 1965 2965 1985
rect 2925 1935 2965 1965
rect 2925 1915 2935 1935
rect 2955 1915 2965 1935
rect 2925 1900 2965 1915
rect 2985 1985 3025 2000
rect 2985 1965 2995 1985
rect 3015 1965 3025 1985
rect 2985 1935 3025 1965
rect 2985 1915 2995 1935
rect 3015 1915 3025 1935
rect 2985 1900 3025 1915
rect 3045 1985 3085 2000
rect 3045 1965 3055 1985
rect 3075 1965 3085 1985
rect 3045 1935 3085 1965
rect 3045 1915 3055 1935
rect 3075 1915 3085 1935
rect 3045 1900 3085 1915
rect 3105 1985 3145 2000
rect 3105 1965 3115 1985
rect 3135 1965 3145 1985
rect 3105 1935 3145 1965
rect 3105 1915 3115 1935
rect 3135 1915 3145 1935
rect 3105 1900 3145 1915
rect 3165 1985 3205 2000
rect 3165 1965 3175 1985
rect 3195 1965 3205 1985
rect 3165 1935 3205 1965
rect 3165 1915 3175 1935
rect 3195 1915 3205 1935
rect 3165 1900 3205 1915
rect 3225 1985 3265 2000
rect 3225 1965 3235 1985
rect 3255 1965 3265 1985
rect 3225 1935 3265 1965
rect 3225 1915 3235 1935
rect 3255 1915 3265 1935
rect 3225 1900 3265 1915
rect 3285 1985 3325 2000
rect 3285 1965 3295 1985
rect 3315 1965 3325 1985
rect 3285 1935 3325 1965
rect 3285 1915 3295 1935
rect 3315 1915 3325 1935
rect 3285 1900 3325 1915
rect 3345 1985 3385 2000
rect 3345 1965 3355 1985
rect 3375 1965 3385 1985
rect 3345 1935 3385 1965
rect 3345 1915 3355 1935
rect 3375 1915 3385 1935
rect 3345 1900 3385 1915
rect 3405 1985 3445 2000
rect 3405 1965 3415 1985
rect 3435 1965 3445 1985
rect 3405 1935 3445 1965
rect 3405 1915 3415 1935
rect 3435 1915 3445 1935
rect 3405 1900 3445 1915
rect 3465 1985 3505 2000
rect 3465 1965 3475 1985
rect 3495 1965 3505 1985
rect 3465 1935 3505 1965
rect 3465 1915 3475 1935
rect 3495 1915 3505 1935
rect 3465 1900 3505 1915
rect 3525 1985 3565 2000
rect 3525 1965 3535 1985
rect 3555 1965 3565 1985
rect 3525 1935 3565 1965
rect 3525 1915 3535 1935
rect 3555 1915 3565 1935
rect 3525 1900 3565 1915
rect 3585 1985 3625 2000
rect 3585 1965 3595 1985
rect 3615 1965 3625 1985
rect 3585 1935 3625 1965
rect 3585 1915 3595 1935
rect 3615 1915 3625 1935
rect 3585 1900 3625 1915
rect 3645 1985 3685 2000
rect 3645 1965 3655 1985
rect 3675 1965 3685 1985
rect 3645 1935 3685 1965
rect 3645 1915 3655 1935
rect 3675 1915 3685 1935
rect 3645 1900 3685 1915
rect 3705 1985 3745 2000
rect 3705 1965 3715 1985
rect 3735 1965 3745 1985
rect 3705 1935 3745 1965
rect 3705 1915 3715 1935
rect 3735 1915 3745 1935
rect 3705 1900 3745 1915
rect 3765 1985 3805 2000
rect 3765 1965 3775 1985
rect 3795 1965 3805 1985
rect 3765 1935 3805 1965
rect 3765 1915 3775 1935
rect 3795 1915 3805 1935
rect 3765 1900 3805 1915
rect 3825 1985 3865 2000
rect 3825 1965 3835 1985
rect 3855 1965 3865 1985
rect 3825 1935 3865 1965
rect 3825 1915 3835 1935
rect 3855 1915 3865 1935
rect 3825 1900 3865 1915
rect 3885 1985 3925 2000
rect 3885 1965 3895 1985
rect 3915 1965 3925 1985
rect 3885 1935 3925 1965
rect 3885 1915 3895 1935
rect 3915 1915 3925 1935
rect 3885 1900 3925 1915
rect 3945 1985 3985 2000
rect 4025 1985 4065 2000
rect 3945 1965 3955 1985
rect 3975 1965 3985 1985
rect 4025 1965 4035 1985
rect 4055 1965 4065 1985
rect 3945 1935 3985 1965
rect 4025 1935 4065 1965
rect 3945 1915 3955 1935
rect 3975 1915 3985 1935
rect 4025 1915 4035 1935
rect 4055 1915 4065 1935
rect 3945 1900 3985 1915
rect 4025 1900 4065 1915
rect 4085 1985 4125 2000
rect 4085 1965 4095 1985
rect 4115 1965 4125 1985
rect 4085 1935 4125 1965
rect 4085 1915 4095 1935
rect 4115 1915 4125 1935
rect 4085 1900 4125 1915
rect 4145 1985 4185 2000
rect 4145 1965 4155 1985
rect 4175 1965 4185 1985
rect 4145 1935 4185 1965
rect 4145 1915 4155 1935
rect 4175 1915 4185 1935
rect 4145 1900 4185 1915
rect 4205 1985 4245 2000
rect 4205 1965 4215 1985
rect 4235 1965 4245 1985
rect 4205 1935 4245 1965
rect 4205 1915 4215 1935
rect 4235 1915 4245 1935
rect 4205 1900 4245 1915
rect 4265 1985 4305 2000
rect 4265 1965 4275 1985
rect 4295 1965 4305 1985
rect 4265 1935 4305 1965
rect 4265 1915 4275 1935
rect 4295 1915 4305 1935
rect 4265 1900 4305 1915
rect 4325 1985 4365 2000
rect 4325 1965 4335 1985
rect 4355 1965 4365 1985
rect 4325 1935 4365 1965
rect 4325 1915 4335 1935
rect 4355 1915 4365 1935
rect 4325 1900 4365 1915
rect 4385 1985 4425 2000
rect 4385 1965 4395 1985
rect 4415 1965 4425 1985
rect 4385 1935 4425 1965
rect 4385 1915 4395 1935
rect 4415 1915 4425 1935
rect 4385 1900 4425 1915
rect 4445 1985 4485 2000
rect 4445 1965 4455 1985
rect 4475 1965 4485 1985
rect 4445 1935 4485 1965
rect 4445 1915 4455 1935
rect 4475 1915 4485 1935
rect 4445 1900 4485 1915
rect 4505 1985 4545 2000
rect 4505 1965 4515 1985
rect 4535 1965 4545 1985
rect 4505 1935 4545 1965
rect 4505 1915 4515 1935
rect 4535 1915 4545 1935
rect 4505 1900 4545 1915
rect 4565 1985 4605 2000
rect 4565 1965 4575 1985
rect 4595 1965 4605 1985
rect 4565 1935 4605 1965
rect 4565 1915 4575 1935
rect 4595 1915 4605 1935
rect 4565 1900 4605 1915
rect 4625 1985 4665 2000
rect 4625 1965 4635 1985
rect 4655 1965 4665 1985
rect 4625 1935 4665 1965
rect 4625 1915 4635 1935
rect 4655 1915 4665 1935
rect 4625 1900 4665 1915
rect 4685 1985 4725 2000
rect 4685 1965 4695 1985
rect 4715 1965 4725 1985
rect 4685 1935 4725 1965
rect 4685 1915 4695 1935
rect 4715 1915 4725 1935
rect 4685 1900 4725 1915
rect 4745 1985 4785 2000
rect 4745 1965 4755 1985
rect 4775 1965 4785 1985
rect 4745 1935 4785 1965
rect 4745 1915 4755 1935
rect 4775 1915 4785 1935
rect 4745 1900 4785 1915
rect 4805 1985 4845 2000
rect 4805 1965 4815 1985
rect 4835 1965 4845 1985
rect 4805 1935 4845 1965
rect 4805 1915 4815 1935
rect 4835 1915 4845 1935
rect 4805 1900 4845 1915
rect 4865 1985 4905 2000
rect 4865 1965 4875 1985
rect 4895 1965 4905 1985
rect 4865 1935 4905 1965
rect 4865 1915 4875 1935
rect 4895 1915 4905 1935
rect 4865 1900 4905 1915
rect 4925 1985 4965 2000
rect 4925 1965 4935 1985
rect 4955 1965 4965 1985
rect 4925 1935 4965 1965
rect 4925 1915 4935 1935
rect 4955 1915 4965 1935
rect 4925 1900 4965 1915
rect 4985 1985 5025 2000
rect 4985 1965 4995 1985
rect 5015 1965 5025 1985
rect 4985 1935 5025 1965
rect 4985 1915 4995 1935
rect 5015 1915 5025 1935
rect 4985 1900 5025 1915
rect 5045 1985 5085 2000
rect 5045 1965 5055 1985
rect 5075 1965 5085 1985
rect 5045 1935 5085 1965
rect 5045 1915 5055 1935
rect 5075 1915 5085 1935
rect 5045 1900 5085 1915
rect 5105 1985 5145 2000
rect 5105 1965 5115 1985
rect 5135 1965 5145 1985
rect 5105 1935 5145 1965
rect 5105 1915 5115 1935
rect 5135 1915 5145 1935
rect 5105 1900 5145 1915
rect 5165 1985 5205 2000
rect 5165 1965 5175 1985
rect 5195 1965 5205 1985
rect 5165 1935 5205 1965
rect 5165 1915 5175 1935
rect 5195 1915 5205 1935
rect 5165 1900 5205 1915
rect 5225 1985 5265 2000
rect 5225 1965 5235 1985
rect 5255 1965 5265 1985
rect 5225 1935 5265 1965
rect 5225 1915 5235 1935
rect 5255 1915 5265 1935
rect 5225 1900 5265 1915
<< ndiffc >>
rect 16250 4355 16270 4375
rect 16310 4360 16330 4380
rect 16370 4360 16390 4380
rect 16430 4355 16450 4375
rect 16580 4370 16600 4390
rect 16640 4370 16660 4390
rect 16700 4370 16720 4390
rect 16760 4370 16780 4390
rect 16820 4370 16840 4390
rect 16880 4370 16900 4390
rect 16940 4370 16960 4390
rect 17090 4355 17110 4375
rect 17150 4355 17170 4375
rect 17210 4355 17230 4375
rect 17270 4355 17290 4375
rect 17330 4355 17350 4375
rect 17390 4355 17410 4375
rect 17450 4355 17470 4375
rect 17510 4355 17530 4375
rect 17570 4355 17590 4375
rect 16260 4120 16280 4140
rect 16315 4120 16335 4140
rect 16370 4120 16390 4140
rect 16425 4120 16445 4140
rect 16480 4120 16500 4140
rect 16535 4120 16555 4140
rect 16590 4120 16610 4140
rect 16645 4120 16665 4140
rect 16700 4120 16720 4140
rect 16755 4120 16775 4140
rect 16810 4120 16830 4140
rect 16865 4120 16885 4140
rect 16920 4120 16940 4140
rect 16975 4120 16995 4140
rect 17030 4120 17050 4140
rect 17085 4120 17105 4140
rect 17140 4120 17160 4140
rect 17195 4120 17215 4140
rect 17250 4120 17270 4140
rect 17305 4120 17325 4140
rect 17360 4120 17380 4140
rect 17415 4120 17435 4140
rect 17470 4120 17490 4140
rect 16205 3815 16225 3835
rect 16260 3815 16280 3835
rect 16315 3815 16335 3835
rect 16370 3815 16390 3835
rect 16425 3815 16445 3835
rect 16480 3815 16500 3835
rect 16535 3815 16555 3835
rect 16590 3815 16610 3835
rect 16645 3815 16665 3835
rect 16700 3815 16720 3835
rect 16755 3815 16775 3835
rect 16810 3815 16830 3835
rect 16865 3815 16885 3835
rect 16945 3815 16965 3835
rect 17000 3815 17020 3835
rect 17055 3815 17075 3835
rect 17110 3815 17130 3835
rect 17165 3815 17185 3835
rect 17220 3815 17240 3835
rect 17275 3815 17295 3835
rect 17330 3815 17350 3835
rect 17385 3815 17405 3835
rect 17440 3815 17460 3835
rect 17495 3815 17515 3835
rect 17550 3815 17570 3835
rect 17605 3815 17625 3835
rect 15165 3550 15185 3570
rect 15165 3500 15185 3520
rect 15165 3450 15185 3470
rect 15165 3400 15185 3420
rect 15165 3350 15185 3370
rect 15165 3300 15185 3320
rect 15165 3250 15185 3270
rect 15165 3200 15185 3220
rect 15165 3150 15185 3170
rect 15165 3100 15185 3120
rect 15165 3050 15185 3070
rect 15165 3000 15185 3020
rect 15220 3550 15240 3570
rect 15220 3500 15240 3520
rect 15220 3450 15240 3470
rect 15220 3400 15240 3420
rect 15220 3350 15240 3370
rect 15220 3300 15240 3320
rect 15220 3250 15240 3270
rect 15220 3200 15240 3220
rect 15220 3150 15240 3170
rect 15220 3100 15240 3120
rect 15220 3050 15240 3070
rect 15220 3000 15240 3020
rect 15275 3550 15295 3570
rect 15275 3500 15295 3520
rect 15275 3450 15295 3470
rect 15275 3400 15295 3420
rect 15275 3350 15295 3370
rect 15275 3300 15295 3320
rect 15275 3250 15295 3270
rect 15275 3200 15295 3220
rect 15275 3150 15295 3170
rect 15275 3100 15295 3120
rect 15275 3050 15295 3070
rect 15275 3000 15295 3020
rect 15330 3550 15350 3570
rect 15330 3500 15350 3520
rect 15330 3450 15350 3470
rect 15330 3400 15350 3420
rect 15330 3350 15350 3370
rect 15330 3300 15350 3320
rect 15330 3250 15350 3270
rect 15330 3200 15350 3220
rect 15330 3150 15350 3170
rect 15330 3100 15350 3120
rect 15330 3050 15350 3070
rect 15330 3000 15350 3020
rect 15385 3550 15405 3570
rect 15385 3500 15405 3520
rect 15385 3450 15405 3470
rect 15385 3400 15405 3420
rect 15385 3350 15405 3370
rect 15385 3300 15405 3320
rect 15385 3250 15405 3270
rect 15385 3200 15405 3220
rect 15385 3150 15405 3170
rect 15385 3100 15405 3120
rect 15385 3050 15405 3070
rect 15385 3000 15405 3020
rect 15440 3550 15460 3570
rect 15440 3500 15460 3520
rect 15440 3450 15460 3470
rect 15440 3400 15460 3420
rect 15440 3350 15460 3370
rect 15440 3300 15460 3320
rect 15440 3250 15460 3270
rect 15440 3200 15460 3220
rect 15440 3150 15460 3170
rect 15440 3100 15460 3120
rect 15440 3050 15460 3070
rect 15440 3000 15460 3020
rect 15495 3550 15515 3570
rect 15495 3500 15515 3520
rect 15495 3450 15515 3470
rect 15495 3400 15515 3420
rect 15495 3350 15515 3370
rect 15495 3300 15515 3320
rect 15495 3250 15515 3270
rect 15495 3200 15515 3220
rect 15495 3150 15515 3170
rect 15495 3100 15515 3120
rect 15495 3050 15515 3070
rect 15495 3000 15515 3020
rect 15550 3550 15570 3570
rect 15550 3500 15570 3520
rect 15550 3450 15570 3470
rect 15550 3400 15570 3420
rect 15550 3350 15570 3370
rect 15550 3300 15570 3320
rect 15550 3250 15570 3270
rect 15550 3200 15570 3220
rect 15550 3150 15570 3170
rect 15550 3100 15570 3120
rect 15550 3050 15570 3070
rect 15550 3000 15570 3020
rect 15605 3550 15625 3570
rect 15605 3500 15625 3520
rect 15605 3450 15625 3470
rect 15605 3400 15625 3420
rect 15605 3350 15625 3370
rect 15605 3300 15625 3320
rect 15605 3250 15625 3270
rect 15605 3200 15625 3220
rect 15605 3150 15625 3170
rect 15605 3100 15625 3120
rect 15605 3050 15625 3070
rect 15605 3000 15625 3020
rect 15660 3550 15680 3570
rect 15660 3500 15680 3520
rect 15660 3450 15680 3470
rect 15660 3400 15680 3420
rect 15660 3350 15680 3370
rect 15660 3300 15680 3320
rect 15660 3250 15680 3270
rect 15660 3200 15680 3220
rect 15660 3150 15680 3170
rect 15660 3100 15680 3120
rect 15660 3050 15680 3070
rect 15660 3000 15680 3020
rect 15715 3550 15735 3570
rect 15715 3500 15735 3520
rect 15715 3450 15735 3470
rect 15715 3400 15735 3420
rect 15715 3350 15735 3370
rect 15715 3300 15735 3320
rect 15715 3250 15735 3270
rect 15715 3200 15735 3220
rect 15715 3150 15735 3170
rect 15715 3100 15735 3120
rect 15715 3050 15735 3070
rect 15715 3000 15735 3020
rect 15770 3550 15790 3570
rect 15770 3500 15790 3520
rect 15770 3450 15790 3470
rect 15770 3400 15790 3420
rect 15770 3350 15790 3370
rect 15770 3300 15790 3320
rect 15770 3250 15790 3270
rect 15770 3200 15790 3220
rect 15770 3150 15790 3170
rect 15770 3100 15790 3120
rect 15770 3050 15790 3070
rect 15770 3000 15790 3020
rect 15825 3550 15845 3570
rect 15825 3500 15845 3520
rect 15825 3450 15845 3470
rect 15825 3400 15845 3420
rect 15825 3350 15845 3370
rect 15825 3300 15845 3320
rect 15825 3250 15845 3270
rect 15825 3200 15845 3220
rect 16230 3540 16250 3560
rect 16230 3490 16250 3510
rect 16230 3440 16250 3460
rect 16230 3390 16250 3410
rect 16230 3340 16250 3360
rect 16230 3290 16250 3310
rect 16230 3240 16250 3260
rect 16230 3190 16250 3210
rect 16290 3540 16310 3560
rect 16290 3490 16310 3510
rect 16290 3440 16310 3460
rect 16290 3390 16310 3410
rect 16290 3340 16310 3360
rect 16290 3290 16310 3310
rect 16290 3240 16310 3260
rect 16290 3190 16310 3210
rect 16350 3540 16370 3560
rect 16350 3490 16370 3510
rect 16350 3440 16370 3460
rect 16350 3390 16370 3410
rect 16350 3340 16370 3360
rect 16350 3290 16370 3310
rect 16350 3240 16370 3260
rect 16350 3190 16370 3210
rect 16410 3540 16430 3560
rect 16410 3490 16430 3510
rect 16410 3440 16430 3460
rect 16410 3390 16430 3410
rect 16410 3340 16430 3360
rect 16410 3290 16430 3310
rect 16410 3240 16430 3260
rect 16410 3190 16430 3210
rect 16470 3540 16490 3560
rect 16470 3490 16490 3510
rect 16470 3440 16490 3460
rect 16470 3390 16490 3410
rect 16470 3340 16490 3360
rect 16470 3290 16490 3310
rect 16470 3240 16490 3260
rect 16470 3190 16490 3210
rect 16530 3540 16550 3560
rect 16530 3490 16550 3510
rect 16530 3440 16550 3460
rect 16530 3390 16550 3410
rect 16530 3340 16550 3360
rect 16530 3290 16550 3310
rect 16530 3240 16550 3260
rect 16530 3190 16550 3210
rect 16590 3540 16610 3560
rect 16590 3490 16610 3510
rect 16590 3440 16610 3460
rect 16590 3390 16610 3410
rect 16590 3340 16610 3360
rect 16590 3290 16610 3310
rect 16590 3240 16610 3260
rect 16590 3190 16610 3210
rect 16650 3540 16670 3560
rect 16650 3490 16670 3510
rect 16650 3440 16670 3460
rect 16650 3390 16670 3410
rect 16650 3340 16670 3360
rect 16650 3290 16670 3310
rect 16650 3240 16670 3260
rect 16650 3190 16670 3210
rect 16710 3540 16730 3560
rect 16710 3490 16730 3510
rect 16710 3440 16730 3460
rect 16710 3390 16730 3410
rect 16710 3340 16730 3360
rect 16710 3290 16730 3310
rect 16710 3240 16730 3260
rect 16710 3190 16730 3210
rect 16770 3540 16790 3560
rect 16770 3490 16790 3510
rect 16770 3440 16790 3460
rect 16770 3390 16790 3410
rect 16770 3340 16790 3360
rect 16770 3290 16790 3310
rect 16770 3240 16790 3260
rect 16770 3190 16790 3210
rect 16830 3540 16850 3560
rect 16830 3490 16850 3510
rect 16830 3440 16850 3460
rect 16830 3390 16850 3410
rect 16830 3340 16850 3360
rect 16830 3290 16850 3310
rect 16830 3240 16850 3260
rect 16830 3190 16850 3210
rect 16890 3540 16910 3560
rect 16890 3490 16910 3510
rect 16890 3440 16910 3460
rect 16890 3390 16910 3410
rect 16890 3340 16910 3360
rect 16890 3290 16910 3310
rect 16890 3240 16910 3260
rect 16890 3190 16910 3210
rect 16950 3540 16970 3560
rect 16950 3490 16970 3510
rect 16950 3440 16970 3460
rect 16950 3390 16970 3410
rect 16950 3340 16970 3360
rect 16950 3290 16970 3310
rect 16950 3240 16970 3260
rect 16950 3190 16970 3210
rect 17010 3540 17030 3560
rect 17010 3490 17030 3510
rect 17010 3440 17030 3460
rect 17010 3390 17030 3410
rect 17010 3340 17030 3360
rect 17010 3290 17030 3310
rect 17010 3240 17030 3260
rect 17010 3190 17030 3210
rect 17070 3540 17090 3560
rect 17070 3490 17090 3510
rect 17070 3440 17090 3460
rect 17070 3390 17090 3410
rect 17070 3340 17090 3360
rect 17070 3290 17090 3310
rect 17070 3240 17090 3260
rect 17070 3190 17090 3210
rect 17130 3540 17150 3560
rect 17130 3490 17150 3510
rect 17130 3440 17150 3460
rect 17130 3390 17150 3410
rect 17130 3340 17150 3360
rect 17130 3290 17150 3310
rect 17130 3240 17150 3260
rect 17130 3190 17150 3210
rect 17190 3540 17210 3560
rect 17190 3490 17210 3510
rect 17190 3440 17210 3460
rect 17190 3390 17210 3410
rect 17190 3340 17210 3360
rect 17190 3290 17210 3310
rect 17190 3240 17210 3260
rect 17190 3190 17210 3210
rect 17250 3540 17270 3560
rect 17250 3490 17270 3510
rect 17250 3440 17270 3460
rect 17250 3390 17270 3410
rect 17250 3340 17270 3360
rect 17250 3290 17270 3310
rect 17250 3240 17270 3260
rect 17250 3190 17270 3210
rect 17310 3540 17330 3560
rect 17310 3490 17330 3510
rect 17310 3440 17330 3460
rect 17310 3390 17330 3410
rect 17310 3340 17330 3360
rect 17310 3290 17330 3310
rect 17310 3240 17330 3260
rect 17310 3190 17330 3210
rect 17370 3540 17390 3560
rect 17370 3490 17390 3510
rect 17370 3440 17390 3460
rect 17370 3390 17390 3410
rect 17370 3340 17390 3360
rect 17370 3290 17390 3310
rect 17370 3240 17390 3260
rect 17370 3190 17390 3210
rect 17430 3540 17450 3560
rect 17430 3490 17450 3510
rect 17430 3440 17450 3460
rect 17430 3390 17450 3410
rect 17430 3340 17450 3360
rect 17430 3290 17450 3310
rect 17430 3240 17450 3260
rect 17430 3190 17450 3210
rect 17490 3540 17510 3560
rect 17490 3490 17510 3510
rect 17490 3440 17510 3460
rect 17490 3390 17510 3410
rect 17490 3340 17510 3360
rect 17490 3290 17510 3310
rect 17490 3240 17510 3260
rect 17490 3190 17510 3210
rect 17550 3540 17570 3560
rect 17550 3490 17570 3510
rect 17550 3440 17570 3460
rect 17550 3390 17570 3410
rect 17550 3340 17570 3360
rect 17550 3290 17570 3310
rect 17550 3240 17570 3260
rect 17550 3190 17570 3210
rect 17955 3550 17975 3570
rect 17955 3500 17975 3520
rect 17955 3450 17975 3470
rect 17955 3400 17975 3420
rect 17955 3350 17975 3370
rect 17955 3300 17975 3320
rect 17955 3250 17975 3270
rect 17955 3200 17975 3220
rect 15825 3150 15845 3170
rect 17955 3150 17975 3170
rect 15825 3100 15845 3120
rect 15825 3050 15845 3070
rect 15825 3000 15845 3020
rect 17955 3100 17975 3120
rect 17955 3050 17975 3070
rect 17955 3000 17975 3020
rect 18010 3550 18030 3570
rect 18010 3500 18030 3520
rect 18010 3450 18030 3470
rect 18010 3400 18030 3420
rect 18010 3350 18030 3370
rect 18010 3300 18030 3320
rect 18010 3250 18030 3270
rect 18010 3200 18030 3220
rect 18010 3150 18030 3170
rect 18010 3100 18030 3120
rect 18010 3050 18030 3070
rect 18010 3000 18030 3020
rect 18065 3550 18085 3570
rect 18065 3500 18085 3520
rect 18065 3450 18085 3470
rect 18065 3400 18085 3420
rect 18065 3350 18085 3370
rect 18065 3300 18085 3320
rect 18065 3250 18085 3270
rect 18065 3200 18085 3220
rect 18065 3150 18085 3170
rect 18065 3100 18085 3120
rect 18065 3050 18085 3070
rect 18065 3000 18085 3020
rect 18120 3550 18140 3570
rect 18120 3500 18140 3520
rect 18120 3450 18140 3470
rect 18120 3400 18140 3420
rect 18120 3350 18140 3370
rect 18120 3300 18140 3320
rect 18120 3250 18140 3270
rect 18120 3200 18140 3220
rect 18120 3150 18140 3170
rect 18120 3100 18140 3120
rect 18120 3050 18140 3070
rect 18120 3000 18140 3020
rect 18175 3550 18195 3570
rect 18175 3500 18195 3520
rect 18175 3450 18195 3470
rect 18175 3400 18195 3420
rect 18175 3350 18195 3370
rect 18175 3300 18195 3320
rect 18175 3250 18195 3270
rect 18175 3200 18195 3220
rect 18175 3150 18195 3170
rect 18175 3100 18195 3120
rect 18175 3050 18195 3070
rect 18175 3000 18195 3020
rect 18230 3550 18250 3570
rect 18230 3500 18250 3520
rect 18230 3450 18250 3470
rect 18230 3400 18250 3420
rect 18230 3350 18250 3370
rect 18230 3300 18250 3320
rect 18230 3250 18250 3270
rect 18230 3200 18250 3220
rect 18230 3150 18250 3170
rect 18230 3100 18250 3120
rect 18230 3050 18250 3070
rect 18230 3000 18250 3020
rect 18285 3550 18305 3570
rect 18285 3500 18305 3520
rect 18285 3450 18305 3470
rect 18285 3400 18305 3420
rect 18285 3350 18305 3370
rect 18285 3300 18305 3320
rect 18285 3250 18305 3270
rect 18285 3200 18305 3220
rect 18285 3150 18305 3170
rect 18285 3100 18305 3120
rect 18285 3050 18305 3070
rect 18285 3000 18305 3020
rect 18340 3550 18360 3570
rect 18340 3500 18360 3520
rect 18340 3450 18360 3470
rect 18340 3400 18360 3420
rect 18340 3350 18360 3370
rect 18340 3300 18360 3320
rect 18340 3250 18360 3270
rect 18340 3200 18360 3220
rect 18340 3150 18360 3170
rect 18340 3100 18360 3120
rect 18340 3050 18360 3070
rect 18340 3000 18360 3020
rect 18395 3550 18415 3570
rect 18395 3500 18415 3520
rect 18395 3450 18415 3470
rect 18395 3400 18415 3420
rect 18395 3350 18415 3370
rect 18395 3300 18415 3320
rect 18395 3250 18415 3270
rect 18395 3200 18415 3220
rect 18395 3150 18415 3170
rect 18395 3100 18415 3120
rect 18395 3050 18415 3070
rect 18395 3000 18415 3020
rect 18450 3550 18470 3570
rect 18450 3500 18470 3520
rect 18450 3450 18470 3470
rect 18450 3400 18470 3420
rect 18450 3350 18470 3370
rect 18450 3300 18470 3320
rect 18450 3250 18470 3270
rect 18450 3200 18470 3220
rect 18450 3150 18470 3170
rect 18450 3100 18470 3120
rect 18450 3050 18470 3070
rect 18450 3000 18470 3020
rect 18505 3550 18525 3570
rect 18505 3500 18525 3520
rect 18505 3450 18525 3470
rect 18505 3400 18525 3420
rect 18505 3350 18525 3370
rect 18505 3300 18525 3320
rect 18505 3250 18525 3270
rect 18505 3200 18525 3220
rect 18505 3150 18525 3170
rect 18505 3100 18525 3120
rect 18505 3050 18525 3070
rect 18505 3000 18525 3020
rect 18560 3550 18580 3570
rect 18560 3500 18580 3520
rect 18560 3450 18580 3470
rect 18560 3400 18580 3420
rect 18560 3350 18580 3370
rect 18560 3300 18580 3320
rect 18560 3250 18580 3270
rect 18560 3200 18580 3220
rect 18560 3150 18580 3170
rect 18560 3100 18580 3120
rect 18560 3050 18580 3070
rect 18560 3000 18580 3020
rect 18615 3550 18635 3570
rect 18615 3500 18635 3520
rect 18615 3450 18635 3470
rect 18615 3400 18635 3420
rect 18615 3350 18635 3370
rect 18615 3300 18635 3320
rect 18615 3250 18635 3270
rect 18615 3200 18635 3220
rect 18615 3150 18635 3170
rect 18615 3100 18635 3120
rect 18615 3050 18635 3070
rect 18615 3000 18635 3020
rect 16230 2860 16250 2880
rect 16230 2810 16250 2830
rect 16230 2760 16250 2780
rect 16230 2710 16250 2730
rect 16230 2660 16250 2680
rect 15165 2620 15185 2640
rect 15165 2570 15185 2590
rect 15165 2520 15185 2540
rect 15165 2470 15185 2490
rect 15220 2620 15240 2640
rect 15220 2570 15240 2590
rect 15220 2520 15240 2540
rect 15220 2470 15240 2490
rect 15275 2620 15295 2640
rect 15275 2570 15295 2590
rect 15275 2520 15295 2540
rect 15275 2470 15295 2490
rect 15330 2620 15350 2640
rect 15330 2570 15350 2590
rect 15330 2520 15350 2540
rect 15330 2470 15350 2490
rect 15385 2620 15405 2640
rect 15385 2570 15405 2590
rect 15385 2520 15405 2540
rect 15385 2470 15405 2490
rect 15440 2620 15460 2640
rect 15440 2570 15460 2590
rect 15440 2520 15460 2540
rect 15440 2470 15460 2490
rect 15495 2620 15515 2640
rect 15495 2570 15515 2590
rect 15495 2520 15515 2540
rect 15495 2470 15515 2490
rect 15550 2620 15570 2640
rect 15550 2570 15570 2590
rect 15550 2520 15570 2540
rect 15550 2470 15570 2490
rect 15605 2620 15625 2640
rect 15605 2570 15625 2590
rect 15605 2520 15625 2540
rect 15605 2470 15625 2490
rect 15660 2620 15680 2640
rect 15660 2570 15680 2590
rect 15660 2520 15680 2540
rect 15660 2470 15680 2490
rect 15715 2620 15735 2640
rect 15715 2570 15735 2590
rect 15715 2520 15735 2540
rect 15715 2470 15735 2490
rect 15770 2620 15790 2640
rect 15770 2570 15790 2590
rect 15770 2520 15790 2540
rect 15770 2470 15790 2490
rect 15825 2620 15845 2640
rect 15825 2570 15845 2590
rect 15825 2520 15845 2540
rect 16230 2610 16250 2630
rect 16230 2560 16250 2580
rect 16230 2510 16250 2530
rect 16290 2860 16310 2880
rect 16290 2810 16310 2830
rect 16290 2760 16310 2780
rect 16290 2710 16310 2730
rect 16290 2660 16310 2680
rect 16290 2610 16310 2630
rect 16290 2560 16310 2580
rect 16290 2510 16310 2530
rect 16350 2860 16370 2880
rect 16350 2810 16370 2830
rect 16350 2760 16370 2780
rect 16350 2710 16370 2730
rect 16350 2660 16370 2680
rect 16350 2610 16370 2630
rect 16350 2560 16370 2580
rect 16350 2510 16370 2530
rect 16410 2860 16430 2880
rect 16410 2810 16430 2830
rect 16410 2760 16430 2780
rect 16410 2710 16430 2730
rect 16410 2660 16430 2680
rect 16410 2610 16430 2630
rect 16410 2560 16430 2580
rect 16410 2510 16430 2530
rect 16470 2860 16490 2880
rect 16470 2810 16490 2830
rect 16470 2760 16490 2780
rect 16470 2710 16490 2730
rect 16470 2660 16490 2680
rect 16470 2610 16490 2630
rect 16470 2560 16490 2580
rect 16470 2510 16490 2530
rect 16530 2860 16550 2880
rect 16530 2810 16550 2830
rect 16530 2760 16550 2780
rect 16530 2710 16550 2730
rect 16530 2660 16550 2680
rect 16530 2610 16550 2630
rect 16530 2560 16550 2580
rect 16530 2510 16550 2530
rect 16590 2860 16610 2880
rect 16590 2810 16610 2830
rect 16590 2760 16610 2780
rect 16590 2710 16610 2730
rect 16590 2660 16610 2680
rect 16590 2610 16610 2630
rect 16590 2560 16610 2580
rect 16590 2510 16610 2530
rect 16650 2860 16670 2880
rect 16650 2810 16670 2830
rect 16650 2760 16670 2780
rect 16650 2710 16670 2730
rect 16650 2660 16670 2680
rect 16650 2610 16670 2630
rect 16650 2560 16670 2580
rect 16650 2510 16670 2530
rect 16710 2860 16730 2880
rect 16710 2810 16730 2830
rect 16710 2760 16730 2780
rect 16710 2710 16730 2730
rect 16710 2660 16730 2680
rect 16710 2610 16730 2630
rect 16710 2560 16730 2580
rect 16710 2510 16730 2530
rect 16770 2860 16790 2880
rect 16770 2810 16790 2830
rect 16770 2760 16790 2780
rect 16770 2710 16790 2730
rect 16770 2660 16790 2680
rect 16770 2610 16790 2630
rect 16770 2560 16790 2580
rect 16770 2510 16790 2530
rect 16830 2860 16850 2880
rect 16830 2810 16850 2830
rect 16830 2760 16850 2780
rect 16830 2710 16850 2730
rect 16830 2660 16850 2680
rect 16830 2610 16850 2630
rect 16830 2560 16850 2580
rect 16830 2510 16850 2530
rect 16890 2860 16910 2880
rect 16890 2810 16910 2830
rect 16890 2760 16910 2780
rect 16890 2710 16910 2730
rect 16890 2660 16910 2680
rect 16890 2610 16910 2630
rect 16890 2560 16910 2580
rect 16890 2510 16910 2530
rect 16950 2860 16970 2880
rect 16950 2810 16970 2830
rect 16950 2760 16970 2780
rect 16950 2710 16970 2730
rect 16950 2660 16970 2680
rect 16950 2610 16970 2630
rect 16950 2560 16970 2580
rect 16950 2510 16970 2530
rect 17010 2860 17030 2880
rect 17010 2810 17030 2830
rect 17010 2760 17030 2780
rect 17010 2710 17030 2730
rect 17010 2660 17030 2680
rect 17010 2610 17030 2630
rect 17010 2560 17030 2580
rect 17010 2510 17030 2530
rect 17070 2860 17090 2880
rect 17070 2810 17090 2830
rect 17070 2760 17090 2780
rect 17070 2710 17090 2730
rect 17070 2660 17090 2680
rect 17070 2610 17090 2630
rect 17070 2560 17090 2580
rect 17070 2510 17090 2530
rect 17130 2860 17150 2880
rect 17130 2810 17150 2830
rect 17130 2760 17150 2780
rect 17130 2710 17150 2730
rect 17130 2660 17150 2680
rect 17130 2610 17150 2630
rect 17130 2560 17150 2580
rect 17130 2510 17150 2530
rect 17190 2860 17210 2880
rect 17190 2810 17210 2830
rect 17190 2760 17210 2780
rect 17190 2710 17210 2730
rect 17190 2660 17210 2680
rect 17190 2610 17210 2630
rect 17190 2560 17210 2580
rect 17190 2510 17210 2530
rect 17250 2860 17270 2880
rect 17250 2810 17270 2830
rect 17250 2760 17270 2780
rect 17250 2710 17270 2730
rect 17250 2660 17270 2680
rect 17250 2610 17270 2630
rect 17250 2560 17270 2580
rect 17250 2510 17270 2530
rect 17310 2860 17330 2880
rect 17310 2810 17330 2830
rect 17310 2760 17330 2780
rect 17310 2710 17330 2730
rect 17310 2660 17330 2680
rect 17310 2610 17330 2630
rect 17310 2560 17330 2580
rect 17310 2510 17330 2530
rect 17370 2860 17390 2880
rect 17370 2810 17390 2830
rect 17370 2760 17390 2780
rect 17370 2710 17390 2730
rect 17370 2660 17390 2680
rect 17370 2610 17390 2630
rect 17370 2560 17390 2580
rect 17370 2510 17390 2530
rect 17430 2860 17450 2880
rect 17430 2810 17450 2830
rect 17430 2760 17450 2780
rect 17430 2710 17450 2730
rect 17430 2660 17450 2680
rect 17430 2610 17450 2630
rect 17430 2560 17450 2580
rect 17430 2510 17450 2530
rect 17490 2860 17510 2880
rect 17490 2810 17510 2830
rect 17490 2760 17510 2780
rect 17490 2710 17510 2730
rect 17490 2660 17510 2680
rect 17490 2610 17510 2630
rect 17490 2560 17510 2580
rect 17490 2510 17510 2530
rect 17550 2860 17570 2880
rect 17550 2810 17570 2830
rect 17550 2760 17570 2780
rect 17550 2710 17570 2730
rect 17550 2660 17570 2680
rect 17550 2610 17570 2630
rect 17550 2560 17570 2580
rect 17550 2510 17570 2530
rect 17955 2620 17975 2640
rect 17955 2570 17975 2590
rect 17955 2520 17975 2540
rect 15825 2470 15845 2490
rect 17955 2470 17975 2490
rect 18010 2620 18030 2640
rect 18010 2570 18030 2590
rect 18010 2520 18030 2540
rect 18010 2470 18030 2490
rect 18065 2620 18085 2640
rect 18065 2570 18085 2590
rect 18065 2520 18085 2540
rect 18065 2470 18085 2490
rect 18120 2620 18140 2640
rect 18120 2570 18140 2590
rect 18120 2520 18140 2540
rect 18120 2470 18140 2490
rect 18175 2620 18195 2640
rect 18175 2570 18195 2590
rect 18175 2520 18195 2540
rect 18175 2470 18195 2490
rect 18230 2620 18250 2640
rect 18230 2570 18250 2590
rect 18230 2520 18250 2540
rect 18230 2470 18250 2490
rect 18285 2620 18305 2640
rect 18285 2570 18305 2590
rect 18285 2520 18305 2540
rect 18285 2470 18305 2490
rect 18340 2620 18360 2640
rect 18340 2570 18360 2590
rect 18340 2520 18360 2540
rect 18340 2470 18360 2490
rect 18395 2620 18415 2640
rect 18395 2570 18415 2590
rect 18395 2520 18415 2540
rect 18395 2470 18415 2490
rect 18450 2620 18470 2640
rect 18450 2570 18470 2590
rect 18450 2520 18470 2540
rect 18450 2470 18470 2490
rect 18505 2620 18525 2640
rect 18505 2570 18525 2590
rect 18505 2520 18525 2540
rect 18505 2470 18525 2490
rect 18560 2620 18580 2640
rect 18560 2570 18580 2590
rect 18560 2520 18580 2540
rect 18560 2470 18580 2490
rect 18615 2620 18635 2640
rect 18615 2570 18635 2590
rect 18615 2520 18635 2540
rect 18615 2470 18635 2490
rect 15165 2230 15185 2250
rect 15165 2180 15185 2200
rect 15165 2130 15185 2150
rect 15165 2080 15185 2100
rect 15165 2030 15185 2050
rect 15165 1980 15185 2000
rect 15220 2230 15240 2250
rect 15220 2180 15240 2200
rect 15220 2130 15240 2150
rect 15220 2080 15240 2100
rect 15220 2030 15240 2050
rect 15220 1980 15240 2000
rect 15275 2230 15295 2250
rect 15275 2180 15295 2200
rect 15275 2130 15295 2150
rect 15275 2080 15295 2100
rect 15275 2030 15295 2050
rect 15275 1980 15295 2000
rect 15330 2230 15350 2250
rect 15330 2180 15350 2200
rect 15330 2130 15350 2150
rect 15330 2080 15350 2100
rect 15330 2030 15350 2050
rect 15330 1980 15350 2000
rect 15385 2230 15405 2250
rect 15385 2180 15405 2200
rect 15385 2130 15405 2150
rect 15385 2080 15405 2100
rect 15385 2030 15405 2050
rect 15385 1980 15405 2000
rect 15440 2230 15460 2250
rect 15440 2180 15460 2200
rect 15440 2130 15460 2150
rect 15440 2080 15460 2100
rect 15440 2030 15460 2050
rect 15440 1980 15460 2000
rect 15495 2230 15515 2250
rect 15495 2180 15515 2200
rect 15495 2130 15515 2150
rect 15495 2080 15515 2100
rect 15495 2030 15515 2050
rect 15495 1980 15515 2000
rect 15550 2230 15570 2250
rect 15550 2180 15570 2200
rect 15550 2130 15570 2150
rect 15550 2080 15570 2100
rect 15550 2030 15570 2050
rect 15550 1980 15570 2000
rect 15605 2230 15625 2250
rect 15605 2180 15625 2200
rect 15605 2130 15625 2150
rect 15605 2080 15625 2100
rect 15605 2030 15625 2050
rect 15605 1980 15625 2000
rect 15660 2230 15680 2250
rect 15660 2180 15680 2200
rect 15660 2130 15680 2150
rect 15660 2080 15680 2100
rect 15660 2030 15680 2050
rect 15660 1980 15680 2000
rect 15715 2230 15735 2250
rect 15715 2180 15735 2200
rect 15715 2130 15735 2150
rect 15715 2080 15735 2100
rect 15715 2030 15735 2050
rect 15715 1980 15735 2000
rect 15770 2230 15790 2250
rect 15770 2180 15790 2200
rect 15770 2130 15790 2150
rect 15770 2080 15790 2100
rect 15770 2030 15790 2050
rect 15770 1980 15790 2000
rect 15825 2230 15845 2250
rect 15825 2180 15845 2200
rect 17955 2230 17975 2250
rect 17955 2180 17975 2200
rect 15825 2130 15845 2150
rect 17955 2130 17975 2150
rect 15825 2080 15845 2100
rect 15825 2030 15845 2050
rect 15825 1980 15845 2000
rect 16285 2095 16305 2115
rect 16285 2045 16305 2065
rect 16285 1995 16305 2015
rect 16340 2095 16360 2115
rect 16340 2045 16360 2065
rect 16340 1995 16360 2015
rect 16395 2095 16415 2115
rect 16395 2045 16415 2065
rect 16395 1995 16415 2015
rect 16450 2095 16470 2115
rect 16450 2045 16470 2065
rect 16450 1995 16470 2015
rect 16505 2095 16525 2115
rect 16505 2045 16525 2065
rect 16505 1995 16525 2015
rect 16560 2095 16580 2115
rect 16560 2045 16580 2065
rect 16560 1995 16580 2015
rect 16615 2095 16635 2115
rect 16615 2045 16635 2065
rect 16615 1995 16635 2015
rect 16670 2095 16690 2115
rect 16670 2045 16690 2065
rect 16670 1995 16690 2015
rect 16725 2095 16745 2115
rect 16725 2045 16745 2065
rect 16725 1995 16745 2015
rect 16780 2095 16800 2115
rect 16780 2045 16800 2065
rect 16780 1995 16800 2015
rect 16835 2095 16855 2115
rect 16835 2045 16855 2065
rect 16835 1995 16855 2015
rect 16890 2095 16910 2115
rect 16890 2045 16910 2065
rect 16890 1995 16910 2015
rect 16945 2095 16965 2115
rect 16945 2045 16965 2065
rect 16945 1995 16965 2015
rect 17000 2095 17020 2115
rect 17000 2045 17020 2065
rect 17000 1995 17020 2015
rect 17055 2095 17075 2115
rect 17055 2045 17075 2065
rect 17055 1995 17075 2015
rect 17110 2095 17130 2115
rect 17110 2045 17130 2065
rect 17110 1995 17130 2015
rect 17165 2095 17185 2115
rect 17165 2045 17185 2065
rect 17165 1995 17185 2015
rect 17220 2095 17240 2115
rect 17220 2045 17240 2065
rect 17220 1995 17240 2015
rect 17275 2095 17295 2115
rect 17275 2045 17295 2065
rect 17275 1995 17295 2015
rect 17330 2095 17350 2115
rect 17330 2045 17350 2065
rect 17330 1995 17350 2015
rect 17385 2095 17405 2115
rect 17385 2045 17405 2065
rect 17385 1995 17405 2015
rect 17440 2095 17460 2115
rect 17440 2045 17460 2065
rect 17440 1995 17460 2015
rect 17495 2095 17515 2115
rect 17495 2045 17515 2065
rect 17495 1995 17515 2015
rect 17955 2080 17975 2100
rect 17955 2030 17975 2050
rect 17955 1980 17975 2000
rect 18010 2230 18030 2250
rect 18010 2180 18030 2200
rect 18010 2130 18030 2150
rect 18010 2080 18030 2100
rect 18010 2030 18030 2050
rect 18010 1980 18030 2000
rect 18065 2230 18085 2250
rect 18065 2180 18085 2200
rect 18065 2130 18085 2150
rect 18065 2080 18085 2100
rect 18065 2030 18085 2050
rect 18065 1980 18085 2000
rect 18120 2230 18140 2250
rect 18120 2180 18140 2200
rect 18120 2130 18140 2150
rect 18120 2080 18140 2100
rect 18120 2030 18140 2050
rect 18120 1980 18140 2000
rect 18175 2230 18195 2250
rect 18175 2180 18195 2200
rect 18175 2130 18195 2150
rect 18175 2080 18195 2100
rect 18175 2030 18195 2050
rect 18175 1980 18195 2000
rect 18230 2230 18250 2250
rect 18230 2180 18250 2200
rect 18230 2130 18250 2150
rect 18230 2080 18250 2100
rect 18230 2030 18250 2050
rect 18230 1980 18250 2000
rect 18285 2230 18305 2250
rect 18285 2180 18305 2200
rect 18285 2130 18305 2150
rect 18285 2080 18305 2100
rect 18285 2030 18305 2050
rect 18285 1980 18305 2000
rect 18340 2230 18360 2250
rect 18340 2180 18360 2200
rect 18340 2130 18360 2150
rect 18340 2080 18360 2100
rect 18340 2030 18360 2050
rect 18340 1980 18360 2000
rect 18395 2230 18415 2250
rect 18395 2180 18415 2200
rect 18395 2130 18415 2150
rect 18395 2080 18415 2100
rect 18395 2030 18415 2050
rect 18395 1980 18415 2000
rect 18450 2230 18470 2250
rect 18450 2180 18470 2200
rect 18450 2130 18470 2150
rect 18450 2080 18470 2100
rect 18450 2030 18470 2050
rect 18450 1980 18470 2000
rect 18505 2230 18525 2250
rect 18505 2180 18525 2200
rect 18505 2130 18525 2150
rect 18505 2080 18525 2100
rect 18505 2030 18525 2050
rect 18505 1980 18525 2000
rect 18560 2230 18580 2250
rect 18560 2180 18580 2200
rect 18560 2130 18580 2150
rect 18560 2080 18580 2100
rect 18560 2030 18580 2050
rect 18560 1980 18580 2000
rect 18615 2230 18635 2250
rect 18615 2180 18635 2200
rect 18615 2130 18635 2150
rect 18615 2080 18635 2100
rect 18615 2030 18635 2050
rect 18615 1980 18635 2000
rect 3175 1630 3195 1650
rect 3235 1630 3255 1650
rect 3295 1630 3315 1650
rect 3355 1630 3375 1650
rect 3415 1630 3435 1650
rect 3475 1630 3495 1650
rect 3535 1630 3555 1650
rect 3595 1630 3615 1650
rect 3655 1630 3675 1650
rect 3715 1630 3735 1650
rect 3775 1630 3795 1650
rect 4215 1630 4235 1650
rect 4275 1630 4295 1650
rect 4335 1630 4355 1650
rect 4395 1630 4415 1650
rect 4455 1630 4475 1650
rect 4515 1630 4535 1650
rect 4575 1630 4595 1650
rect 4635 1630 4655 1650
rect 4695 1630 4715 1650
rect 4755 1630 4775 1650
rect 4815 1630 4835 1650
rect 15165 1620 15185 1640
rect 2845 1420 2865 1440
rect 2845 1370 2865 1390
rect 2845 1320 2865 1340
rect 2845 1270 2865 1290
rect 2845 1220 2865 1240
rect 3385 1420 3405 1440
rect 3385 1370 3405 1390
rect 3385 1320 3405 1340
rect 3385 1270 3405 1290
rect 3385 1220 3405 1240
rect 3925 1420 3945 1440
rect 3925 1370 3945 1390
rect 3925 1320 3945 1340
rect 3925 1270 3945 1290
rect 3925 1220 3945 1240
rect 4065 1420 4085 1440
rect 4065 1370 4085 1390
rect 4065 1320 4085 1340
rect 4065 1270 4085 1290
rect 4065 1220 4085 1240
rect 4605 1420 4625 1440
rect 4605 1370 4625 1390
rect 4605 1320 4625 1340
rect 4605 1270 4625 1290
rect 4605 1220 4625 1240
rect 5145 1420 5165 1440
rect 5145 1370 5165 1390
rect 5145 1320 5165 1340
rect 5145 1270 5165 1290
rect 5145 1220 5165 1240
rect 2955 1040 2975 1060
rect 2955 990 2975 1010
rect 3995 1040 4015 1060
rect 3995 990 4015 1010
rect 5035 1040 5055 1060
rect 5035 990 5055 1010
rect 15165 1570 15185 1590
rect 15165 1520 15185 1540
rect 15165 1470 15185 1490
rect 15165 1420 15185 1440
rect 15165 1370 15185 1390
rect 15165 1320 15185 1340
rect 15165 1270 15185 1290
rect 15165 1220 15185 1240
rect 15165 1170 15185 1190
rect 15165 1120 15185 1140
rect 15165 1070 15185 1090
rect 15165 1020 15185 1040
rect 15165 970 15185 990
rect 15265 1620 15285 1640
rect 15265 1570 15285 1590
rect 15265 1520 15285 1540
rect 15265 1470 15285 1490
rect 15265 1420 15285 1440
rect 15265 1370 15285 1390
rect 15265 1320 15285 1340
rect 15265 1270 15285 1290
rect 15265 1220 15285 1240
rect 15265 1170 15285 1190
rect 15265 1120 15285 1140
rect 15265 1070 15285 1090
rect 15265 1020 15285 1040
rect 15265 970 15285 990
rect 15365 1620 15385 1640
rect 15365 1570 15385 1590
rect 15365 1520 15385 1540
rect 15365 1470 15385 1490
rect 15365 1420 15385 1440
rect 15365 1370 15385 1390
rect 15365 1320 15385 1340
rect 15365 1270 15385 1290
rect 15365 1220 15385 1240
rect 15365 1170 15385 1190
rect 15365 1120 15385 1140
rect 15365 1070 15385 1090
rect 15365 1020 15385 1040
rect 15365 970 15385 990
rect 15465 1620 15485 1640
rect 15465 1570 15485 1590
rect 15465 1520 15485 1540
rect 15465 1470 15485 1490
rect 15465 1420 15485 1440
rect 15465 1370 15485 1390
rect 15465 1320 15485 1340
rect 15465 1270 15485 1290
rect 15465 1220 15485 1240
rect 15465 1170 15485 1190
rect 15465 1120 15485 1140
rect 15465 1070 15485 1090
rect 15465 1020 15485 1040
rect 15465 970 15485 990
rect 15565 1620 15585 1640
rect 15565 1570 15585 1590
rect 15565 1520 15585 1540
rect 15565 1470 15585 1490
rect 15565 1420 15585 1440
rect 15565 1370 15585 1390
rect 15565 1320 15585 1340
rect 15565 1270 15585 1290
rect 15565 1220 15585 1240
rect 15565 1170 15585 1190
rect 15565 1120 15585 1140
rect 15565 1070 15585 1090
rect 15565 1020 15585 1040
rect 15565 970 15585 990
rect 15665 1620 15685 1640
rect 15665 1570 15685 1590
rect 15665 1520 15685 1540
rect 15665 1470 15685 1490
rect 15665 1420 15685 1440
rect 15665 1370 15685 1390
rect 15665 1320 15685 1340
rect 15665 1270 15685 1290
rect 15665 1220 15685 1240
rect 15665 1170 15685 1190
rect 15665 1120 15685 1140
rect 15665 1070 15685 1090
rect 15665 1020 15685 1040
rect 15665 970 15685 990
rect 15765 1620 15785 1640
rect 15765 1570 15785 1590
rect 15765 1520 15785 1540
rect 16040 1630 16060 1650
rect 16040 1580 16060 1600
rect 16040 1530 16060 1550
rect 16095 1630 16115 1650
rect 16095 1580 16115 1600
rect 16095 1530 16115 1550
rect 16150 1630 16170 1650
rect 16150 1580 16170 1600
rect 16150 1530 16170 1550
rect 16205 1630 16225 1650
rect 16205 1580 16225 1600
rect 16205 1530 16225 1550
rect 16260 1630 16280 1650
rect 16260 1580 16280 1600
rect 16260 1530 16280 1550
rect 16315 1630 16335 1650
rect 16315 1580 16335 1600
rect 16315 1530 16335 1550
rect 16370 1630 16390 1650
rect 16370 1580 16390 1600
rect 16370 1530 16390 1550
rect 16425 1630 16445 1650
rect 16425 1580 16445 1600
rect 16425 1530 16445 1550
rect 16480 1630 16500 1650
rect 16480 1580 16500 1600
rect 16480 1530 16500 1550
rect 16535 1630 16555 1650
rect 16535 1580 16555 1600
rect 16535 1530 16555 1550
rect 16590 1630 16610 1650
rect 16590 1580 16610 1600
rect 16590 1530 16610 1550
rect 16645 1630 16665 1650
rect 16645 1580 16665 1600
rect 16645 1530 16665 1550
rect 16700 1630 16720 1650
rect 16780 1630 16800 1650
rect 16700 1580 16720 1600
rect 16780 1580 16800 1600
rect 16700 1530 16720 1550
rect 16780 1530 16800 1550
rect 16835 1630 16855 1650
rect 16835 1580 16855 1600
rect 16835 1530 16855 1550
rect 16890 1630 16910 1650
rect 16890 1580 16910 1600
rect 16890 1530 16910 1550
rect 16945 1630 16965 1650
rect 16945 1580 16965 1600
rect 16945 1530 16965 1550
rect 17000 1630 17020 1650
rect 17080 1630 17100 1650
rect 17000 1580 17020 1600
rect 17080 1580 17100 1600
rect 17000 1530 17020 1550
rect 17080 1530 17100 1550
rect 17135 1630 17155 1650
rect 17135 1580 17155 1600
rect 17135 1530 17155 1550
rect 17190 1630 17210 1650
rect 17190 1580 17210 1600
rect 17190 1530 17210 1550
rect 17245 1630 17265 1650
rect 17245 1580 17265 1600
rect 17245 1530 17265 1550
rect 17300 1630 17320 1650
rect 17300 1580 17320 1600
rect 17300 1530 17320 1550
rect 17355 1630 17375 1650
rect 17355 1580 17375 1600
rect 17355 1530 17375 1550
rect 17410 1630 17430 1650
rect 17410 1580 17430 1600
rect 17410 1530 17430 1550
rect 17465 1630 17485 1650
rect 17465 1580 17485 1600
rect 17465 1530 17485 1550
rect 17520 1630 17540 1650
rect 17520 1580 17540 1600
rect 17520 1530 17540 1550
rect 17575 1630 17595 1650
rect 17575 1580 17595 1600
rect 17575 1530 17595 1550
rect 17630 1630 17650 1650
rect 17630 1580 17650 1600
rect 17630 1530 17650 1550
rect 17685 1630 17705 1650
rect 17685 1580 17705 1600
rect 17685 1530 17705 1550
rect 17740 1630 17760 1650
rect 17740 1580 17760 1600
rect 17740 1530 17760 1550
rect 18015 1620 18035 1640
rect 18015 1570 18035 1590
rect 18015 1520 18035 1540
rect 15765 1470 15785 1490
rect 18015 1470 18035 1490
rect 15765 1420 15785 1440
rect 15765 1370 15785 1390
rect 15765 1320 15785 1340
rect 15765 1270 15785 1290
rect 18015 1420 18035 1440
rect 18015 1370 18035 1390
rect 18015 1320 18035 1340
rect 18015 1270 18035 1290
rect 15765 1220 15785 1240
rect 15765 1170 15785 1190
rect 18015 1220 18035 1240
rect 15765 1120 15785 1140
rect 15765 1070 15785 1090
rect 15765 1020 15785 1040
rect 15765 970 15785 990
rect 16215 1150 16235 1170
rect 16215 1100 16235 1120
rect 16215 1050 16235 1070
rect 16215 1000 16235 1020
rect 16215 950 16235 970
rect 16270 1150 16290 1170
rect 16270 1100 16290 1120
rect 16270 1050 16290 1070
rect 16270 1000 16290 1020
rect 16270 950 16290 970
rect 16325 1150 16345 1170
rect 16325 1100 16345 1120
rect 16325 1050 16345 1070
rect 16325 1000 16345 1020
rect 16325 950 16345 970
rect 16380 1150 16400 1170
rect 16380 1100 16400 1120
rect 16380 1050 16400 1070
rect 16380 1000 16400 1020
rect 16380 950 16400 970
rect 16435 1150 16455 1170
rect 16435 1100 16455 1120
rect 16435 1050 16455 1070
rect 16435 1000 16455 1020
rect 16435 950 16455 970
rect 16490 1150 16510 1170
rect 16490 1100 16510 1120
rect 16490 1050 16510 1070
rect 16490 1000 16510 1020
rect 16490 950 16510 970
rect 16545 1150 16565 1170
rect 16545 1100 16565 1120
rect 16545 1050 16565 1070
rect 16545 1000 16565 1020
rect 16545 950 16565 970
rect 16600 1150 16620 1170
rect 16600 1100 16620 1120
rect 16600 1050 16620 1070
rect 16600 1000 16620 1020
rect 16600 950 16620 970
rect 16655 1150 16675 1170
rect 16655 1100 16675 1120
rect 16655 1050 16675 1070
rect 16655 1000 16675 1020
rect 16655 950 16675 970
rect 16710 1150 16730 1170
rect 16710 1100 16730 1120
rect 16710 1050 16730 1070
rect 16710 1000 16730 1020
rect 16710 950 16730 970
rect 16765 1150 16785 1170
rect 16765 1100 16785 1120
rect 16765 1050 16785 1070
rect 16765 1000 16785 1020
rect 16765 950 16785 970
rect 16820 1150 16840 1170
rect 16820 1100 16840 1120
rect 16820 1050 16840 1070
rect 16820 1000 16840 1020
rect 16820 950 16840 970
rect 16875 1150 16895 1170
rect 16875 1100 16895 1120
rect 16875 1050 16895 1070
rect 16875 1000 16895 1020
rect 16875 950 16895 970
rect 16930 1150 16950 1170
rect 16930 1100 16950 1120
rect 16930 1050 16950 1070
rect 16930 1000 16950 1020
rect 16930 950 16950 970
rect 16985 1150 17005 1170
rect 16985 1100 17005 1120
rect 16985 1050 17005 1070
rect 16985 1000 17005 1020
rect 16985 950 17005 970
rect 17040 1150 17060 1170
rect 17040 1100 17060 1120
rect 17040 1050 17060 1070
rect 17040 1000 17060 1020
rect 17040 950 17060 970
rect 17095 1150 17115 1170
rect 17095 1100 17115 1120
rect 17095 1050 17115 1070
rect 17095 1000 17115 1020
rect 17095 950 17115 970
rect 17150 1150 17170 1170
rect 17150 1100 17170 1120
rect 17150 1050 17170 1070
rect 17150 1000 17170 1020
rect 17150 950 17170 970
rect 17205 1150 17225 1170
rect 17205 1100 17225 1120
rect 17205 1050 17225 1070
rect 17205 1000 17225 1020
rect 17205 950 17225 970
rect 17260 1150 17280 1170
rect 17260 1100 17280 1120
rect 17260 1050 17280 1070
rect 17260 1000 17280 1020
rect 17260 950 17280 970
rect 17315 1150 17335 1170
rect 17315 1100 17335 1120
rect 17315 1050 17335 1070
rect 17315 1000 17335 1020
rect 17315 950 17335 970
rect 17370 1150 17390 1170
rect 17370 1100 17390 1120
rect 17370 1050 17390 1070
rect 17370 1000 17390 1020
rect 17370 950 17390 970
rect 17425 1150 17445 1170
rect 17425 1100 17445 1120
rect 17425 1050 17445 1070
rect 17425 1000 17445 1020
rect 17425 950 17445 970
rect 17480 1150 17500 1170
rect 17480 1100 17500 1120
rect 17480 1050 17500 1070
rect 17480 1000 17500 1020
rect 17480 950 17500 970
rect 17535 1150 17555 1170
rect 17535 1100 17555 1120
rect 17535 1050 17555 1070
rect 17535 1000 17555 1020
rect 17535 950 17555 970
rect 17590 1150 17610 1170
rect 17590 1100 17610 1120
rect 17590 1050 17610 1070
rect 17590 1000 17610 1020
rect 17590 950 17610 970
rect 18015 1170 18035 1190
rect 18015 1120 18035 1140
rect 18015 1070 18035 1090
rect 18015 1020 18035 1040
rect 18015 970 18035 990
rect 18115 1620 18135 1640
rect 18115 1570 18135 1590
rect 18115 1520 18135 1540
rect 18115 1470 18135 1490
rect 18115 1420 18135 1440
rect 18115 1370 18135 1390
rect 18115 1320 18135 1340
rect 18115 1270 18135 1290
rect 18115 1220 18135 1240
rect 18115 1170 18135 1190
rect 18115 1120 18135 1140
rect 18115 1070 18135 1090
rect 18115 1020 18135 1040
rect 18115 970 18135 990
rect 18215 1620 18235 1640
rect 18215 1570 18235 1590
rect 18215 1520 18235 1540
rect 18215 1470 18235 1490
rect 18215 1420 18235 1440
rect 18215 1370 18235 1390
rect 18215 1320 18235 1340
rect 18215 1270 18235 1290
rect 18215 1220 18235 1240
rect 18215 1170 18235 1190
rect 18215 1120 18235 1140
rect 18215 1070 18235 1090
rect 18215 1020 18235 1040
rect 18215 970 18235 990
rect 18315 1620 18335 1640
rect 18315 1570 18335 1590
rect 18315 1520 18335 1540
rect 18315 1470 18335 1490
rect 18315 1420 18335 1440
rect 18315 1370 18335 1390
rect 18315 1320 18335 1340
rect 18315 1270 18335 1290
rect 18315 1220 18335 1240
rect 18315 1170 18335 1190
rect 18315 1120 18335 1140
rect 18315 1070 18335 1090
rect 18315 1020 18335 1040
rect 18315 970 18335 990
rect 18415 1620 18435 1640
rect 18415 1570 18435 1590
rect 18415 1520 18435 1540
rect 18415 1470 18435 1490
rect 18415 1420 18435 1440
rect 18415 1370 18435 1390
rect 18415 1320 18435 1340
rect 18415 1270 18435 1290
rect 18415 1220 18435 1240
rect 18415 1170 18435 1190
rect 18415 1120 18435 1140
rect 18415 1070 18435 1090
rect 18415 1020 18435 1040
rect 18415 970 18435 990
rect 18515 1620 18535 1640
rect 18515 1570 18535 1590
rect 18515 1520 18535 1540
rect 18515 1470 18535 1490
rect 18515 1420 18535 1440
rect 18515 1370 18535 1390
rect 18515 1320 18535 1340
rect 18515 1270 18535 1290
rect 18515 1220 18535 1240
rect 18515 1170 18535 1190
rect 18515 1120 18535 1140
rect 18515 1070 18535 1090
rect 18515 1020 18535 1040
rect 18515 970 18535 990
rect 18615 1620 18635 1640
rect 18615 1570 18635 1590
rect 18615 1520 18635 1540
rect 18615 1470 18635 1490
rect 18615 1420 18635 1440
rect 18615 1370 18635 1390
rect 18615 1320 18635 1340
rect 18615 1270 18635 1290
rect 18615 1220 18635 1240
rect 18615 1170 18635 1190
rect 18615 1120 18635 1140
rect 18615 1070 18635 1090
rect 18615 1020 18635 1040
rect 18615 970 18635 990
rect 3005 845 3025 865
rect 3005 795 3025 815
rect 3095 845 3115 865
rect 3095 795 3115 815
rect 3185 845 3205 865
rect 3185 795 3205 815
rect 3275 845 3295 865
rect 3275 795 3295 815
rect 3365 845 3385 865
rect 3365 795 3385 815
rect 3455 845 3475 865
rect 3455 795 3475 815
rect 3545 845 3565 865
rect 3545 795 3565 815
rect 3635 845 3655 865
rect 3635 795 3655 815
rect 3725 845 3745 865
rect 3725 795 3745 815
rect 3815 845 3835 865
rect 3815 795 3835 815
rect 3905 845 3925 865
rect 3905 795 3925 815
rect 3995 845 4015 865
rect 3995 795 4015 815
rect 4085 845 4105 865
rect 4085 795 4105 815
rect 4175 845 4195 865
rect 4175 795 4195 815
rect 4265 845 4285 865
rect 4265 795 4285 815
rect 4355 845 4375 865
rect 4355 795 4375 815
rect 4445 845 4465 865
rect 4445 795 4465 815
rect 4535 845 4555 865
rect 4535 795 4555 815
rect 4625 845 4645 865
rect 4625 795 4645 815
rect 4715 845 4735 865
rect 4715 795 4735 815
rect 4805 845 4825 865
rect 4805 795 4825 815
rect 4895 845 4915 865
rect 4895 795 4915 815
rect 4985 845 5005 865
rect 4985 795 5005 815
rect 16270 710 16290 730
rect 16270 660 16290 680
rect 16500 710 16520 730
rect 16890 715 16910 735
rect 16945 715 16965 735
rect 17000 715 17020 735
rect 17055 715 17075 735
rect 17110 715 17130 735
rect 17165 715 17185 735
rect 17220 715 17240 735
rect 17275 715 17295 735
rect 17330 715 17350 735
rect 17385 715 17405 735
rect 17440 715 17460 735
rect 17495 715 17515 735
rect 17550 715 17570 735
rect 16500 660 16520 680
<< pdiffc >>
rect 3005 2895 3025 2915
rect 3005 2845 3025 2865
rect 3095 2895 3115 2915
rect 3095 2845 3115 2865
rect 3185 2895 3205 2915
rect 3185 2845 3205 2865
rect 3275 2895 3295 2915
rect 3275 2845 3295 2865
rect 3365 2895 3385 2915
rect 3365 2845 3385 2865
rect 3455 2895 3475 2915
rect 3455 2845 3475 2865
rect 3545 2895 3565 2915
rect 3545 2845 3565 2865
rect 3635 2895 3655 2915
rect 3635 2845 3655 2865
rect 3725 2895 3745 2915
rect 3725 2845 3745 2865
rect 3815 2895 3835 2915
rect 3815 2845 3835 2865
rect 3905 2895 3925 2915
rect 3905 2845 3925 2865
rect 3995 2895 4015 2915
rect 3995 2845 4015 2865
rect 4085 2895 4105 2915
rect 4085 2845 4105 2865
rect 4175 2895 4195 2915
rect 4175 2845 4195 2865
rect 4265 2895 4285 2915
rect 4265 2845 4285 2865
rect 4355 2895 4375 2915
rect 4355 2845 4375 2865
rect 4445 2895 4465 2915
rect 4445 2845 4465 2865
rect 4535 2895 4555 2915
rect 4535 2845 4555 2865
rect 4625 2895 4645 2915
rect 4625 2845 4645 2865
rect 4715 2895 4735 2915
rect 4715 2845 4735 2865
rect 4805 2895 4825 2915
rect 4805 2845 4825 2865
rect 4895 2895 4915 2915
rect 4895 2845 4915 2865
rect 4985 2895 5005 2915
rect 4985 2845 5005 2865
rect 3185 2665 3205 2685
rect 3185 2615 3205 2635
rect 3185 2565 3205 2585
rect 3185 2515 3205 2535
rect 3185 2465 3205 2485
rect 3185 2415 3205 2435
rect 3275 2665 3295 2685
rect 3275 2615 3295 2635
rect 3275 2565 3295 2585
rect 3275 2515 3295 2535
rect 3275 2465 3295 2485
rect 3275 2415 3295 2435
rect 3365 2665 3385 2685
rect 3365 2615 3385 2635
rect 3365 2565 3385 2585
rect 3365 2515 3385 2535
rect 3365 2465 3385 2485
rect 3365 2415 3385 2435
rect 3455 2665 3475 2685
rect 3455 2615 3475 2635
rect 3455 2565 3475 2585
rect 3455 2515 3475 2535
rect 3455 2465 3475 2485
rect 3455 2415 3475 2435
rect 3545 2665 3565 2685
rect 3545 2615 3565 2635
rect 3545 2565 3565 2585
rect 3545 2515 3565 2535
rect 3545 2465 3565 2485
rect 3545 2415 3565 2435
rect 3635 2665 3655 2685
rect 3635 2615 3655 2635
rect 3635 2565 3655 2585
rect 3635 2515 3655 2535
rect 3635 2465 3655 2485
rect 3635 2415 3655 2435
rect 3725 2665 3745 2685
rect 3725 2615 3745 2635
rect 3725 2565 3745 2585
rect 3725 2515 3745 2535
rect 3725 2465 3745 2485
rect 3725 2415 3745 2435
rect 3815 2665 3835 2685
rect 3815 2615 3835 2635
rect 3815 2565 3835 2585
rect 3815 2515 3835 2535
rect 3815 2465 3835 2485
rect 3815 2415 3835 2435
rect 3905 2665 3925 2685
rect 3905 2615 3925 2635
rect 3905 2565 3925 2585
rect 3905 2515 3925 2535
rect 3905 2465 3925 2485
rect 3905 2415 3925 2435
rect 3995 2665 4015 2685
rect 3995 2615 4015 2635
rect 3995 2565 4015 2585
rect 3995 2515 4015 2535
rect 3995 2465 4015 2485
rect 3995 2415 4015 2435
rect 4085 2665 4105 2685
rect 4085 2615 4105 2635
rect 4085 2565 4105 2585
rect 4085 2515 4105 2535
rect 4085 2465 4105 2485
rect 4085 2415 4105 2435
rect 4175 2665 4195 2685
rect 4175 2615 4195 2635
rect 4175 2565 4195 2585
rect 4175 2515 4195 2535
rect 4175 2465 4195 2485
rect 4175 2415 4195 2435
rect 4265 2665 4285 2685
rect 4265 2615 4285 2635
rect 4265 2565 4285 2585
rect 4265 2515 4285 2535
rect 4265 2465 4285 2485
rect 4265 2415 4285 2435
rect 4355 2665 4375 2685
rect 4355 2615 4375 2635
rect 4355 2565 4375 2585
rect 4355 2515 4375 2535
rect 4355 2465 4375 2485
rect 4355 2415 4375 2435
rect 4445 2665 4465 2685
rect 4445 2615 4465 2635
rect 4445 2565 4465 2585
rect 4445 2515 4465 2535
rect 4445 2465 4465 2485
rect 4445 2415 4465 2435
rect 4535 2665 4555 2685
rect 4535 2615 4555 2635
rect 4535 2565 4555 2585
rect 4535 2515 4555 2535
rect 4535 2465 4555 2485
rect 4535 2415 4555 2435
rect 4625 2665 4645 2685
rect 4625 2615 4645 2635
rect 4625 2565 4645 2585
rect 4625 2515 4645 2535
rect 4625 2465 4645 2485
rect 4625 2415 4645 2435
rect 4715 2665 4735 2685
rect 4715 2615 4735 2635
rect 4715 2565 4735 2585
rect 4715 2515 4735 2535
rect 4715 2465 4735 2485
rect 4715 2415 4735 2435
rect 4805 2665 4825 2685
rect 4805 2615 4825 2635
rect 4805 2565 4825 2585
rect 4805 2515 4825 2535
rect 4805 2465 4825 2485
rect 4805 2415 4825 2435
rect 2575 1965 2595 1985
rect 2575 1915 2595 1935
rect 2630 1965 2650 1985
rect 2630 1915 2650 1935
rect 2685 1965 2705 1985
rect 2685 1915 2705 1935
rect 2755 1965 2775 1985
rect 2755 1915 2775 1935
rect 2815 1965 2835 1985
rect 2815 1915 2835 1935
rect 2875 1965 2895 1985
rect 2875 1915 2895 1935
rect 2935 1965 2955 1985
rect 2935 1915 2955 1935
rect 2995 1965 3015 1985
rect 2995 1915 3015 1935
rect 3055 1965 3075 1985
rect 3055 1915 3075 1935
rect 3115 1965 3135 1985
rect 3115 1915 3135 1935
rect 3175 1965 3195 1985
rect 3175 1915 3195 1935
rect 3235 1965 3255 1985
rect 3235 1915 3255 1935
rect 3295 1965 3315 1985
rect 3295 1915 3315 1935
rect 3355 1965 3375 1985
rect 3355 1915 3375 1935
rect 3415 1965 3435 1985
rect 3415 1915 3435 1935
rect 3475 1965 3495 1985
rect 3475 1915 3495 1935
rect 3535 1965 3555 1985
rect 3535 1915 3555 1935
rect 3595 1965 3615 1985
rect 3595 1915 3615 1935
rect 3655 1965 3675 1985
rect 3655 1915 3675 1935
rect 3715 1965 3735 1985
rect 3715 1915 3735 1935
rect 3775 1965 3795 1985
rect 3775 1915 3795 1935
rect 3835 1965 3855 1985
rect 3835 1915 3855 1935
rect 3895 1965 3915 1985
rect 3895 1915 3915 1935
rect 3955 1965 3975 1985
rect 4035 1965 4055 1985
rect 3955 1915 3975 1935
rect 4035 1915 4055 1935
rect 4095 1965 4115 1985
rect 4095 1915 4115 1935
rect 4155 1965 4175 1985
rect 4155 1915 4175 1935
rect 4215 1965 4235 1985
rect 4215 1915 4235 1935
rect 4275 1965 4295 1985
rect 4275 1915 4295 1935
rect 4335 1965 4355 1985
rect 4335 1915 4355 1935
rect 4395 1965 4415 1985
rect 4395 1915 4415 1935
rect 4455 1965 4475 1985
rect 4455 1915 4475 1935
rect 4515 1965 4535 1985
rect 4515 1915 4535 1935
rect 4575 1965 4595 1985
rect 4575 1915 4595 1935
rect 4635 1965 4655 1985
rect 4635 1915 4655 1935
rect 4695 1965 4715 1985
rect 4695 1915 4715 1935
rect 4755 1965 4775 1985
rect 4755 1915 4775 1935
rect 4815 1965 4835 1985
rect 4815 1915 4835 1935
rect 4875 1965 4895 1985
rect 4875 1915 4895 1935
rect 4935 1965 4955 1985
rect 4935 1915 4955 1935
rect 4995 1965 5015 1985
rect 4995 1915 5015 1935
rect 5055 1965 5075 1985
rect 5055 1915 5075 1935
rect 5115 1965 5135 1985
rect 5115 1915 5135 1935
rect 5175 1965 5195 1985
rect 5175 1915 5195 1935
rect 5235 1965 5255 1985
rect 5235 1915 5255 1935
<< psubdiff >>
rect 16200 4375 16240 4403
rect 16200 4355 16210 4375
rect 16230 4355 16240 4375
rect 16200 4340 16240 4355
rect 16460 4375 16500 4403
rect 16460 4355 16470 4375
rect 16490 4355 16500 4375
rect 16460 4340 16500 4355
rect 16530 4390 16570 4420
rect 16530 4370 16540 4390
rect 16560 4370 16570 4390
rect 16530 4340 16570 4370
rect 16970 4390 17010 4420
rect 16970 4370 16980 4390
rect 17000 4370 17010 4390
rect 16970 4340 17010 4370
rect 17040 4375 17080 4395
rect 17040 4355 17050 4375
rect 17070 4355 17080 4375
rect 17040 4335 17080 4355
rect 17600 4375 17640 4395
rect 17600 4355 17610 4375
rect 17630 4355 17640 4375
rect 17600 4335 17640 4355
rect 16210 4140 16250 4155
rect 16210 4120 16220 4140
rect 16240 4120 16250 4140
rect 16210 4105 16250 4120
rect 17500 4140 17540 4155
rect 17500 4120 17510 4140
rect 17530 4120 17540 4140
rect 17500 4105 17540 4120
rect 16155 3835 16195 3850
rect 16155 3815 16165 3835
rect 16185 3815 16195 3835
rect 16155 3800 16195 3815
rect 16895 3835 16935 3850
rect 16895 3815 16905 3835
rect 16925 3815 16935 3835
rect 16895 3800 16935 3815
rect 17635 3835 17675 3850
rect 17635 3815 17645 3835
rect 17665 3815 17675 3835
rect 17635 3800 17675 3815
rect 15115 3570 15155 3585
rect 15115 3550 15125 3570
rect 15145 3550 15155 3570
rect 15115 3520 15155 3550
rect 15115 3500 15125 3520
rect 15145 3500 15155 3520
rect 15115 3470 15155 3500
rect 15115 3450 15125 3470
rect 15145 3450 15155 3470
rect 15115 3420 15155 3450
rect 15115 3400 15125 3420
rect 15145 3400 15155 3420
rect 15115 3370 15155 3400
rect 15115 3350 15125 3370
rect 15145 3350 15155 3370
rect 15115 3320 15155 3350
rect 15115 3300 15125 3320
rect 15145 3300 15155 3320
rect 15115 3270 15155 3300
rect 15115 3250 15125 3270
rect 15145 3250 15155 3270
rect 15115 3220 15155 3250
rect 15115 3200 15125 3220
rect 15145 3200 15155 3220
rect 15115 3170 15155 3200
rect 15115 3150 15125 3170
rect 15145 3150 15155 3170
rect 15115 3120 15155 3150
rect 15115 3100 15125 3120
rect 15145 3100 15155 3120
rect 15115 3070 15155 3100
rect 15115 3050 15125 3070
rect 15145 3050 15155 3070
rect 15115 3020 15155 3050
rect 15115 3000 15125 3020
rect 15145 3000 15155 3020
rect 15115 2985 15155 3000
rect 15855 3570 15895 3585
rect 15855 3550 15865 3570
rect 15885 3550 15895 3570
rect 15855 3520 15895 3550
rect 15855 3500 15865 3520
rect 15885 3500 15895 3520
rect 15855 3470 15895 3500
rect 15855 3450 15865 3470
rect 15885 3450 15895 3470
rect 15855 3420 15895 3450
rect 15855 3400 15865 3420
rect 15885 3400 15895 3420
rect 15855 3370 15895 3400
rect 15855 3350 15865 3370
rect 15885 3350 15895 3370
rect 15855 3320 15895 3350
rect 15855 3300 15865 3320
rect 15885 3300 15895 3320
rect 15855 3270 15895 3300
rect 15855 3250 15865 3270
rect 15885 3250 15895 3270
rect 15855 3220 15895 3250
rect 15855 3200 15865 3220
rect 15885 3200 15895 3220
rect 15855 3170 15895 3200
rect 16180 3560 16220 3575
rect 16180 3540 16190 3560
rect 16210 3540 16220 3560
rect 16180 3510 16220 3540
rect 16180 3490 16190 3510
rect 16210 3490 16220 3510
rect 16180 3460 16220 3490
rect 16180 3440 16190 3460
rect 16210 3440 16220 3460
rect 16180 3410 16220 3440
rect 16180 3390 16190 3410
rect 16210 3390 16220 3410
rect 16180 3360 16220 3390
rect 16180 3340 16190 3360
rect 16210 3340 16220 3360
rect 16180 3310 16220 3340
rect 16180 3290 16190 3310
rect 16210 3290 16220 3310
rect 16180 3260 16220 3290
rect 16180 3240 16190 3260
rect 16210 3240 16220 3260
rect 16180 3210 16220 3240
rect 16180 3190 16190 3210
rect 16210 3190 16220 3210
rect 16180 3175 16220 3190
rect 17580 3560 17620 3575
rect 17580 3540 17590 3560
rect 17610 3540 17620 3560
rect 17580 3510 17620 3540
rect 17580 3490 17590 3510
rect 17610 3490 17620 3510
rect 17580 3460 17620 3490
rect 17580 3440 17590 3460
rect 17610 3440 17620 3460
rect 17580 3410 17620 3440
rect 17580 3390 17590 3410
rect 17610 3390 17620 3410
rect 17580 3360 17620 3390
rect 17580 3340 17590 3360
rect 17610 3340 17620 3360
rect 17580 3310 17620 3340
rect 17580 3290 17590 3310
rect 17610 3290 17620 3310
rect 17580 3260 17620 3290
rect 17580 3240 17590 3260
rect 17610 3240 17620 3260
rect 17580 3210 17620 3240
rect 17580 3190 17590 3210
rect 17610 3190 17620 3210
rect 17580 3175 17620 3190
rect 17905 3570 17945 3585
rect 17905 3550 17915 3570
rect 17935 3550 17945 3570
rect 17905 3520 17945 3550
rect 17905 3500 17915 3520
rect 17935 3500 17945 3520
rect 17905 3470 17945 3500
rect 17905 3450 17915 3470
rect 17935 3450 17945 3470
rect 17905 3420 17945 3450
rect 17905 3400 17915 3420
rect 17935 3400 17945 3420
rect 17905 3370 17945 3400
rect 17905 3350 17915 3370
rect 17935 3350 17945 3370
rect 17905 3320 17945 3350
rect 17905 3300 17915 3320
rect 17935 3300 17945 3320
rect 17905 3270 17945 3300
rect 17905 3250 17915 3270
rect 17935 3250 17945 3270
rect 17905 3220 17945 3250
rect 17905 3200 17915 3220
rect 17935 3200 17945 3220
rect 15855 3150 15865 3170
rect 15885 3150 15895 3170
rect 17905 3170 17945 3200
rect 17905 3150 17915 3170
rect 17935 3150 17945 3170
rect 15855 3120 15895 3150
rect 17905 3120 17945 3150
rect 15855 3100 15865 3120
rect 15885 3100 15895 3120
rect 15855 3070 15895 3100
rect 15855 3050 15865 3070
rect 15885 3050 15895 3070
rect 15855 3020 15895 3050
rect 15855 3000 15865 3020
rect 15885 3000 15895 3020
rect 15855 2985 15895 3000
rect 17905 3100 17915 3120
rect 17935 3100 17945 3120
rect 17905 3070 17945 3100
rect 17905 3050 17915 3070
rect 17935 3050 17945 3070
rect 17905 3020 17945 3050
rect 17905 3000 17915 3020
rect 17935 3000 17945 3020
rect 17905 2985 17945 3000
rect 18645 3570 18685 3585
rect 18645 3550 18655 3570
rect 18675 3550 18685 3570
rect 18645 3520 18685 3550
rect 18645 3500 18655 3520
rect 18675 3500 18685 3520
rect 18645 3470 18685 3500
rect 18645 3450 18655 3470
rect 18675 3450 18685 3470
rect 18645 3420 18685 3450
rect 18645 3400 18655 3420
rect 18675 3400 18685 3420
rect 18645 3370 18685 3400
rect 18645 3350 18655 3370
rect 18675 3350 18685 3370
rect 18645 3320 18685 3350
rect 18645 3300 18655 3320
rect 18675 3300 18685 3320
rect 18645 3270 18685 3300
rect 18645 3250 18655 3270
rect 18675 3250 18685 3270
rect 18645 3220 18685 3250
rect 18645 3200 18655 3220
rect 18675 3200 18685 3220
rect 18645 3170 18685 3200
rect 18645 3150 18655 3170
rect 18675 3150 18685 3170
rect 18645 3120 18685 3150
rect 18645 3100 18655 3120
rect 18675 3100 18685 3120
rect 18645 3070 18685 3100
rect 18645 3050 18655 3070
rect 18675 3050 18685 3070
rect 18645 3020 18685 3050
rect 18645 3000 18655 3020
rect 18675 3000 18685 3020
rect 18645 2985 18685 3000
rect 905 2910 1125 2920
rect 905 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 905 2870 1125 2880
rect 16180 2880 16220 2895
rect 16180 2860 16190 2880
rect 16210 2860 16220 2880
rect 16180 2830 16220 2860
rect 16180 2810 16190 2830
rect 16210 2810 16220 2830
rect 16180 2780 16220 2810
rect 16180 2760 16190 2780
rect 16210 2760 16220 2780
rect 16180 2730 16220 2760
rect 16180 2710 16190 2730
rect 16210 2710 16220 2730
rect 16180 2680 16220 2710
rect 16180 2660 16190 2680
rect 16210 2660 16220 2680
rect 15115 2640 15155 2655
rect 15115 2620 15125 2640
rect 15145 2620 15155 2640
rect 15115 2590 15155 2620
rect 15115 2570 15125 2590
rect 15145 2570 15155 2590
rect 15115 2540 15155 2570
rect 15115 2520 15125 2540
rect 15145 2520 15155 2540
rect 15115 2490 15155 2520
rect 15115 2470 15125 2490
rect 15145 2470 15155 2490
rect 15115 2455 15155 2470
rect 15855 2640 15895 2655
rect 15855 2620 15865 2640
rect 15885 2620 15895 2640
rect 15855 2590 15895 2620
rect 15855 2570 15865 2590
rect 15885 2570 15895 2590
rect 15855 2540 15895 2570
rect 15855 2520 15865 2540
rect 15885 2520 15895 2540
rect 15855 2490 15895 2520
rect 16180 2630 16220 2660
rect 16180 2610 16190 2630
rect 16210 2610 16220 2630
rect 16180 2580 16220 2610
rect 16180 2560 16190 2580
rect 16210 2560 16220 2580
rect 16180 2530 16220 2560
rect 16180 2510 16190 2530
rect 16210 2510 16220 2530
rect 16180 2495 16220 2510
rect 17580 2880 17620 2895
rect 17580 2860 17590 2880
rect 17610 2860 17620 2880
rect 17580 2830 17620 2860
rect 17580 2810 17590 2830
rect 17610 2810 17620 2830
rect 17580 2780 17620 2810
rect 17580 2760 17590 2780
rect 17610 2760 17620 2780
rect 17580 2730 17620 2760
rect 17580 2710 17590 2730
rect 17610 2710 17620 2730
rect 17580 2680 17620 2710
rect 17580 2660 17590 2680
rect 17610 2660 17620 2680
rect 17580 2630 17620 2660
rect 17580 2610 17590 2630
rect 17610 2610 17620 2630
rect 17580 2580 17620 2610
rect 17580 2560 17590 2580
rect 17610 2560 17620 2580
rect 17580 2530 17620 2560
rect 17580 2510 17590 2530
rect 17610 2510 17620 2530
rect 17580 2495 17620 2510
rect 17905 2640 17945 2655
rect 17905 2620 17915 2640
rect 17935 2620 17945 2640
rect 17905 2590 17945 2620
rect 17905 2570 17915 2590
rect 17935 2570 17945 2590
rect 17905 2540 17945 2570
rect 17905 2520 17915 2540
rect 17935 2520 17945 2540
rect 15855 2470 15865 2490
rect 15885 2470 15895 2490
rect 17905 2490 17945 2520
rect 17905 2470 17915 2490
rect 17935 2470 17945 2490
rect 15855 2455 15895 2470
rect 17905 2455 17945 2470
rect 18645 2640 18685 2655
rect 18645 2620 18655 2640
rect 18675 2620 18685 2640
rect 18645 2590 18685 2620
rect 18645 2570 18655 2590
rect 18675 2570 18685 2590
rect 18645 2540 18685 2570
rect 18645 2520 18655 2540
rect 18675 2520 18685 2540
rect 18645 2490 18685 2520
rect 18645 2470 18655 2490
rect 18675 2470 18685 2490
rect 18645 2455 18685 2470
rect 15115 2250 15155 2265
rect 15115 2230 15125 2250
rect 15145 2230 15155 2250
rect 15115 2200 15155 2230
rect 15115 2180 15125 2200
rect 15145 2180 15155 2200
rect 15115 2150 15155 2180
rect 15115 2130 15125 2150
rect 15145 2130 15155 2150
rect 15115 2100 15155 2130
rect 15115 2080 15125 2100
rect 15145 2080 15155 2100
rect 15115 2050 15155 2080
rect 15115 2030 15125 2050
rect 15145 2030 15155 2050
rect 15115 2000 15155 2030
rect 15115 1980 15125 2000
rect 15145 1980 15155 2000
rect 15115 1965 15155 1980
rect 15855 2250 15895 2265
rect 15855 2230 15865 2250
rect 15885 2230 15895 2250
rect 15855 2200 15895 2230
rect 15855 2180 15865 2200
rect 15885 2180 15895 2200
rect 17905 2250 17945 2265
rect 17905 2230 17915 2250
rect 17935 2230 17945 2250
rect 17905 2200 17945 2230
rect 15855 2150 15895 2180
rect 17905 2180 17915 2200
rect 17935 2180 17945 2200
rect 15855 2130 15865 2150
rect 15885 2130 15895 2150
rect 17905 2150 17945 2180
rect 17905 2130 17915 2150
rect 17935 2130 17945 2150
rect 15855 2100 15895 2130
rect 15855 2080 15865 2100
rect 15885 2080 15895 2100
rect 15855 2050 15895 2080
rect 15855 2030 15865 2050
rect 15885 2030 15895 2050
rect 15855 2000 15895 2030
rect 15855 1980 15865 2000
rect 15885 1980 15895 2000
rect 16235 2115 16275 2130
rect 16235 2095 16245 2115
rect 16265 2095 16275 2115
rect 16235 2065 16275 2095
rect 16235 2045 16245 2065
rect 16265 2045 16275 2065
rect 16235 2015 16275 2045
rect 16235 1995 16245 2015
rect 16265 1995 16275 2015
rect 16235 1980 16275 1995
rect 17525 2115 17565 2130
rect 17525 2095 17535 2115
rect 17555 2095 17565 2115
rect 17525 2065 17565 2095
rect 17525 2045 17535 2065
rect 17555 2045 17565 2065
rect 17525 2015 17565 2045
rect 17525 1995 17535 2015
rect 17555 1995 17565 2015
rect 17525 1980 17565 1995
rect 17905 2100 17945 2130
rect 17905 2080 17915 2100
rect 17935 2080 17945 2100
rect 17905 2050 17945 2080
rect 17905 2030 17915 2050
rect 17935 2030 17945 2050
rect 17905 2000 17945 2030
rect 17905 1980 17915 2000
rect 17935 1980 17945 2000
rect 15855 1965 15895 1980
rect 17905 1965 17945 1980
rect 18645 2250 18685 2265
rect 18645 2230 18655 2250
rect 18675 2230 18685 2250
rect 18645 2200 18685 2230
rect 18645 2180 18655 2200
rect 18675 2180 18685 2200
rect 18645 2150 18685 2180
rect 18645 2130 18655 2150
rect 18675 2130 18685 2150
rect 18645 2100 18685 2130
rect 18645 2080 18655 2100
rect 18675 2080 18685 2100
rect 18645 2050 18685 2080
rect 18645 2030 18655 2050
rect 18675 2030 18685 2050
rect 18645 2000 18685 2030
rect 18645 1980 18655 2000
rect 18675 1980 18685 2000
rect 18645 1965 18685 1980
rect -50 1715 100 1730
rect -50 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 100 1715
rect -50 1680 100 1695
rect 3980 1650 4030 1665
rect 3980 1630 3995 1650
rect 4015 1630 4030 1650
rect 3980 1615 4030 1630
rect 15115 1640 15155 1655
rect 15115 1620 15125 1640
rect 15145 1620 15155 1640
rect 5065 1060 5105 1075
rect 5065 1040 5075 1060
rect 5095 1040 5105 1060
rect 5065 1010 5105 1040
rect 5065 990 5075 1010
rect 5095 990 5105 1010
rect 5065 975 5105 990
rect 15115 1590 15155 1620
rect 15115 1570 15125 1590
rect 15145 1570 15155 1590
rect 15115 1540 15155 1570
rect 15115 1520 15125 1540
rect 15145 1520 15155 1540
rect 15115 1490 15155 1520
rect 15115 1470 15125 1490
rect 15145 1470 15155 1490
rect 15115 1440 15155 1470
rect 15115 1420 15125 1440
rect 15145 1420 15155 1440
rect 15115 1390 15155 1420
rect 15115 1370 15125 1390
rect 15145 1370 15155 1390
rect 15115 1340 15155 1370
rect 15115 1320 15125 1340
rect 15145 1320 15155 1340
rect 15115 1290 15155 1320
rect 15115 1270 15125 1290
rect 15145 1270 15155 1290
rect 15115 1240 15155 1270
rect 15115 1220 15125 1240
rect 15145 1220 15155 1240
rect 15115 1190 15155 1220
rect 15115 1170 15125 1190
rect 15145 1170 15155 1190
rect 15115 1140 15155 1170
rect 15115 1120 15125 1140
rect 15145 1120 15155 1140
rect 15115 1090 15155 1120
rect 15115 1070 15125 1090
rect 15145 1070 15155 1090
rect 15115 1040 15155 1070
rect 15115 1020 15125 1040
rect 15145 1020 15155 1040
rect 15115 990 15155 1020
rect 15115 970 15125 990
rect 15145 970 15155 990
rect 15115 955 15155 970
rect 15795 1640 15835 1655
rect 15795 1620 15805 1640
rect 15825 1620 15835 1640
rect 15795 1590 15835 1620
rect 15795 1570 15805 1590
rect 15825 1570 15835 1590
rect 15795 1540 15835 1570
rect 15795 1520 15805 1540
rect 15825 1520 15835 1540
rect 15795 1490 15835 1520
rect 15990 1650 16030 1665
rect 15990 1630 16000 1650
rect 16020 1630 16030 1650
rect 15990 1600 16030 1630
rect 15990 1580 16000 1600
rect 16020 1580 16030 1600
rect 15990 1550 16030 1580
rect 15990 1530 16000 1550
rect 16020 1530 16030 1550
rect 15990 1515 16030 1530
rect 16730 1650 16770 1665
rect 16730 1630 16740 1650
rect 16760 1630 16770 1650
rect 16730 1600 16770 1630
rect 16730 1580 16740 1600
rect 16760 1580 16770 1600
rect 16730 1550 16770 1580
rect 16730 1530 16740 1550
rect 16760 1530 16770 1550
rect 16730 1515 16770 1530
rect 17030 1650 17070 1665
rect 17030 1630 17040 1650
rect 17060 1630 17070 1650
rect 17030 1600 17070 1630
rect 17030 1580 17040 1600
rect 17060 1580 17070 1600
rect 17030 1550 17070 1580
rect 17030 1530 17040 1550
rect 17060 1530 17070 1550
rect 17030 1515 17070 1530
rect 17770 1650 17810 1665
rect 17770 1630 17780 1650
rect 17800 1630 17810 1650
rect 17770 1600 17810 1630
rect 17770 1580 17780 1600
rect 17800 1580 17810 1600
rect 17770 1550 17810 1580
rect 17770 1530 17780 1550
rect 17800 1530 17810 1550
rect 17770 1515 17810 1530
rect 17965 1640 18005 1655
rect 17965 1620 17975 1640
rect 17995 1620 18005 1640
rect 17965 1590 18005 1620
rect 17965 1570 17975 1590
rect 17995 1570 18005 1590
rect 17965 1540 18005 1570
rect 17965 1520 17975 1540
rect 17995 1520 18005 1540
rect 15795 1470 15805 1490
rect 15825 1470 15835 1490
rect 15795 1440 15835 1470
rect 17965 1490 18005 1520
rect 17965 1470 17975 1490
rect 17995 1470 18005 1490
rect 15795 1420 15805 1440
rect 15825 1420 15835 1440
rect 15795 1390 15835 1420
rect 15795 1370 15805 1390
rect 15825 1370 15835 1390
rect 15795 1340 15835 1370
rect 15795 1320 15805 1340
rect 15825 1320 15835 1340
rect 15795 1290 15835 1320
rect 15795 1270 15805 1290
rect 15825 1270 15835 1290
rect 15795 1240 15835 1270
rect 17965 1440 18005 1470
rect 17965 1420 17975 1440
rect 17995 1420 18005 1440
rect 17965 1390 18005 1420
rect 17965 1370 17975 1390
rect 17995 1370 18005 1390
rect 17965 1340 18005 1370
rect 17965 1320 17975 1340
rect 17995 1320 18005 1340
rect 17965 1290 18005 1320
rect 17965 1270 17975 1290
rect 17995 1270 18005 1290
rect 15795 1220 15805 1240
rect 15825 1220 15835 1240
rect 15795 1190 15835 1220
rect 15795 1170 15805 1190
rect 15825 1170 15835 1190
rect 17965 1240 18005 1270
rect 17965 1220 17975 1240
rect 17995 1220 18005 1240
rect 17965 1190 18005 1220
rect 15795 1140 15835 1170
rect 15795 1120 15805 1140
rect 15825 1120 15835 1140
rect 15795 1090 15835 1120
rect 15795 1070 15805 1090
rect 15825 1070 15835 1090
rect 15795 1040 15835 1070
rect 15795 1020 15805 1040
rect 15825 1020 15835 1040
rect 15795 990 15835 1020
rect 15795 970 15805 990
rect 15825 970 15835 990
rect 15795 955 15835 970
rect 16165 1170 16205 1185
rect 16165 1150 16175 1170
rect 16195 1150 16205 1170
rect 16165 1120 16205 1150
rect 16165 1100 16175 1120
rect 16195 1100 16205 1120
rect 16165 1070 16205 1100
rect 16165 1050 16175 1070
rect 16195 1050 16205 1070
rect 16165 1020 16205 1050
rect 16165 1000 16175 1020
rect 16195 1000 16205 1020
rect 16165 970 16205 1000
rect 16165 950 16175 970
rect 16195 950 16205 970
rect 16165 935 16205 950
rect 17620 1170 17660 1185
rect 17620 1150 17630 1170
rect 17650 1150 17660 1170
rect 17620 1120 17660 1150
rect 17620 1100 17630 1120
rect 17650 1100 17660 1120
rect 17620 1070 17660 1100
rect 17620 1050 17630 1070
rect 17650 1050 17660 1070
rect 17620 1020 17660 1050
rect 17620 1000 17630 1020
rect 17650 1000 17660 1020
rect 17620 970 17660 1000
rect 17620 950 17630 970
rect 17650 950 17660 970
rect 17965 1170 17975 1190
rect 17995 1170 18005 1190
rect 17965 1140 18005 1170
rect 17965 1120 17975 1140
rect 17995 1120 18005 1140
rect 17965 1090 18005 1120
rect 17965 1070 17975 1090
rect 17995 1070 18005 1090
rect 17965 1040 18005 1070
rect 17965 1020 17975 1040
rect 17995 1020 18005 1040
rect 17965 990 18005 1020
rect 17965 970 17975 990
rect 17995 970 18005 990
rect 17965 955 18005 970
rect 18645 1640 18685 1655
rect 18645 1620 18655 1640
rect 18675 1620 18685 1640
rect 18645 1590 18685 1620
rect 18645 1570 18655 1590
rect 18675 1570 18685 1590
rect 18645 1540 18685 1570
rect 18645 1520 18655 1540
rect 18675 1520 18685 1540
rect 18645 1490 18685 1520
rect 18645 1470 18655 1490
rect 18675 1470 18685 1490
rect 18645 1440 18685 1470
rect 18645 1420 18655 1440
rect 18675 1420 18685 1440
rect 18645 1390 18685 1420
rect 18645 1370 18655 1390
rect 18675 1370 18685 1390
rect 18645 1340 18685 1370
rect 18645 1320 18655 1340
rect 18675 1320 18685 1340
rect 18645 1290 18685 1320
rect 18645 1270 18655 1290
rect 18675 1270 18685 1290
rect 18645 1240 18685 1270
rect 18645 1220 18655 1240
rect 18675 1220 18685 1240
rect 18645 1190 18685 1220
rect 18645 1170 18655 1190
rect 18675 1170 18685 1190
rect 18645 1140 18685 1170
rect 18645 1120 18655 1140
rect 18675 1120 18685 1140
rect 18645 1090 18685 1120
rect 18645 1070 18655 1090
rect 18675 1070 18685 1090
rect 18645 1040 18685 1070
rect 18645 1020 18655 1040
rect 18675 1020 18685 1040
rect 18645 990 18685 1020
rect 18645 970 18655 990
rect 18675 970 18685 990
rect 18645 955 18685 970
rect 17620 935 17660 950
rect 2955 865 2995 880
rect 2955 845 2965 865
rect 2985 845 2995 865
rect 2955 815 2995 845
rect 2955 795 2965 815
rect 2985 795 2995 815
rect 2955 780 2995 795
rect 5015 865 5055 880
rect 5015 845 5025 865
rect 5045 845 5055 865
rect 5015 815 5055 845
rect 5015 795 5025 815
rect 5045 795 5055 815
rect 5015 780 5055 795
rect 16840 735 16880 750
rect 16840 715 16850 735
rect 16870 715 16880 735
rect 16840 700 16880 715
rect 17580 735 17620 750
rect 17580 715 17590 735
rect 17610 715 17620 735
rect 17580 700 17620 715
<< nsubdiff >>
rect 2955 2915 2995 2930
rect 2955 2895 2965 2915
rect 2985 2895 2995 2915
rect 2955 2865 2995 2895
rect 2955 2845 2965 2865
rect 2985 2845 2995 2865
rect 2955 2830 2995 2845
rect 5015 2915 5055 2930
rect 5015 2895 5025 2915
rect 5045 2895 5055 2915
rect 5015 2865 5055 2895
rect 5015 2845 5025 2865
rect 5045 2845 5055 2865
rect 5015 2830 5055 2845
rect 3135 2685 3175 2700
rect 3135 2665 3145 2685
rect 3165 2665 3175 2685
rect 3135 2635 3175 2665
rect 3135 2615 3145 2635
rect 3165 2615 3175 2635
rect 3135 2585 3175 2615
rect 3135 2565 3145 2585
rect 3165 2565 3175 2585
rect 3135 2535 3175 2565
rect 3135 2515 3145 2535
rect 3165 2515 3175 2535
rect 3135 2485 3175 2515
rect 3135 2465 3145 2485
rect 3165 2465 3175 2485
rect 3135 2435 3175 2465
rect 3135 2415 3145 2435
rect 3165 2415 3175 2435
rect 3135 2400 3175 2415
rect 4835 2685 4875 2700
rect 4835 2665 4845 2685
rect 4865 2665 4875 2685
rect 4835 2635 4875 2665
rect 4835 2615 4845 2635
rect 4865 2615 4875 2635
rect 4835 2585 4875 2615
rect 4835 2565 4845 2585
rect 4865 2565 4875 2585
rect 4835 2535 4875 2565
rect 4835 2515 4845 2535
rect 4865 2515 4875 2535
rect 4835 2485 4875 2515
rect 4835 2465 4845 2485
rect 4865 2465 4875 2485
rect 4835 2435 4875 2465
rect 4835 2415 4845 2435
rect 4865 2415 4875 2435
rect 4835 2400 4875 2415
rect 3985 1985 4025 2000
rect 3985 1965 3995 1985
rect 4015 1965 4025 1985
rect 3985 1935 4025 1965
rect 3985 1915 3995 1935
rect 4015 1915 4025 1935
rect 3985 1900 4025 1915
<< psubdiffcont >>
rect 16210 4355 16230 4375
rect 16470 4355 16490 4375
rect 16540 4370 16560 4390
rect 16980 4370 17000 4390
rect 17050 4355 17070 4375
rect 17610 4355 17630 4375
rect 16220 4120 16240 4140
rect 17510 4120 17530 4140
rect 16165 3815 16185 3835
rect 16905 3815 16925 3835
rect 17645 3815 17665 3835
rect 15125 3550 15145 3570
rect 15125 3500 15145 3520
rect 15125 3450 15145 3470
rect 15125 3400 15145 3420
rect 15125 3350 15145 3370
rect 15125 3300 15145 3320
rect 15125 3250 15145 3270
rect 15125 3200 15145 3220
rect 15125 3150 15145 3170
rect 15125 3100 15145 3120
rect 15125 3050 15145 3070
rect 15125 3000 15145 3020
rect 15865 3550 15885 3570
rect 15865 3500 15885 3520
rect 15865 3450 15885 3470
rect 15865 3400 15885 3420
rect 15865 3350 15885 3370
rect 15865 3300 15885 3320
rect 15865 3250 15885 3270
rect 15865 3200 15885 3220
rect 16190 3540 16210 3560
rect 16190 3490 16210 3510
rect 16190 3440 16210 3460
rect 16190 3390 16210 3410
rect 16190 3340 16210 3360
rect 16190 3290 16210 3310
rect 16190 3240 16210 3260
rect 16190 3190 16210 3210
rect 17590 3540 17610 3560
rect 17590 3490 17610 3510
rect 17590 3440 17610 3460
rect 17590 3390 17610 3410
rect 17590 3340 17610 3360
rect 17590 3290 17610 3310
rect 17590 3240 17610 3260
rect 17590 3190 17610 3210
rect 17915 3550 17935 3570
rect 17915 3500 17935 3520
rect 17915 3450 17935 3470
rect 17915 3400 17935 3420
rect 17915 3350 17935 3370
rect 17915 3300 17935 3320
rect 17915 3250 17935 3270
rect 17915 3200 17935 3220
rect 15865 3150 15885 3170
rect 17915 3150 17935 3170
rect 15865 3100 15885 3120
rect 15865 3050 15885 3070
rect 15865 3000 15885 3020
rect 17915 3100 17935 3120
rect 17915 3050 17935 3070
rect 17915 3000 17935 3020
rect 18655 3550 18675 3570
rect 18655 3500 18675 3520
rect 18655 3450 18675 3470
rect 18655 3400 18675 3420
rect 18655 3350 18675 3370
rect 18655 3300 18675 3320
rect 18655 3250 18675 3270
rect 18655 3200 18675 3220
rect 18655 3150 18675 3170
rect 18655 3100 18675 3120
rect 18655 3050 18675 3070
rect 18655 3000 18675 3020
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 16190 2860 16210 2880
rect 16190 2810 16210 2830
rect 16190 2760 16210 2780
rect 16190 2710 16210 2730
rect 16190 2660 16210 2680
rect 15125 2620 15145 2640
rect 15125 2570 15145 2590
rect 15125 2520 15145 2540
rect 15125 2470 15145 2490
rect 15865 2620 15885 2640
rect 15865 2570 15885 2590
rect 15865 2520 15885 2540
rect 16190 2610 16210 2630
rect 16190 2560 16210 2580
rect 16190 2510 16210 2530
rect 17590 2860 17610 2880
rect 17590 2810 17610 2830
rect 17590 2760 17610 2780
rect 17590 2710 17610 2730
rect 17590 2660 17610 2680
rect 17590 2610 17610 2630
rect 17590 2560 17610 2580
rect 17590 2510 17610 2530
rect 17915 2620 17935 2640
rect 17915 2570 17935 2590
rect 17915 2520 17935 2540
rect 15865 2470 15885 2490
rect 17915 2470 17935 2490
rect 18655 2620 18675 2640
rect 18655 2570 18675 2590
rect 18655 2520 18675 2540
rect 18655 2470 18675 2490
rect 15125 2230 15145 2250
rect 15125 2180 15145 2200
rect 15125 2130 15145 2150
rect 15125 2080 15145 2100
rect 15125 2030 15145 2050
rect 15125 1980 15145 2000
rect 15865 2230 15885 2250
rect 15865 2180 15885 2200
rect 17915 2230 17935 2250
rect 17915 2180 17935 2200
rect 15865 2130 15885 2150
rect 17915 2130 17935 2150
rect 15865 2080 15885 2100
rect 15865 2030 15885 2050
rect 15865 1980 15885 2000
rect 16245 2095 16265 2115
rect 16245 2045 16265 2065
rect 16245 1995 16265 2015
rect 17535 2095 17555 2115
rect 17535 2045 17555 2065
rect 17535 1995 17555 2015
rect 17915 2080 17935 2100
rect 17915 2030 17935 2050
rect 17915 1980 17935 2000
rect 18655 2230 18675 2250
rect 18655 2180 18675 2200
rect 18655 2130 18675 2150
rect 18655 2080 18675 2100
rect 18655 2030 18675 2050
rect 18655 1980 18675 2000
rect -35 1695 -15 1715
rect 15 1695 35 1715
rect 65 1695 85 1715
rect 3995 1630 4015 1650
rect 15125 1620 15145 1640
rect 5075 1040 5095 1060
rect 5075 990 5095 1010
rect 15125 1570 15145 1590
rect 15125 1520 15145 1540
rect 15125 1470 15145 1490
rect 15125 1420 15145 1440
rect 15125 1370 15145 1390
rect 15125 1320 15145 1340
rect 15125 1270 15145 1290
rect 15125 1220 15145 1240
rect 15125 1170 15145 1190
rect 15125 1120 15145 1140
rect 15125 1070 15145 1090
rect 15125 1020 15145 1040
rect 15125 970 15145 990
rect 15805 1620 15825 1640
rect 15805 1570 15825 1590
rect 15805 1520 15825 1540
rect 16000 1630 16020 1650
rect 16000 1580 16020 1600
rect 16000 1530 16020 1550
rect 16740 1630 16760 1650
rect 16740 1580 16760 1600
rect 16740 1530 16760 1550
rect 17040 1630 17060 1650
rect 17040 1580 17060 1600
rect 17040 1530 17060 1550
rect 17780 1630 17800 1650
rect 17780 1580 17800 1600
rect 17780 1530 17800 1550
rect 17975 1620 17995 1640
rect 17975 1570 17995 1590
rect 17975 1520 17995 1540
rect 15805 1470 15825 1490
rect 17975 1470 17995 1490
rect 15805 1420 15825 1440
rect 15805 1370 15825 1390
rect 15805 1320 15825 1340
rect 15805 1270 15825 1290
rect 17975 1420 17995 1440
rect 17975 1370 17995 1390
rect 17975 1320 17995 1340
rect 17975 1270 17995 1290
rect 15805 1220 15825 1240
rect 15805 1170 15825 1190
rect 17975 1220 17995 1240
rect 15805 1120 15825 1140
rect 15805 1070 15825 1090
rect 15805 1020 15825 1040
rect 15805 970 15825 990
rect 16175 1150 16195 1170
rect 16175 1100 16195 1120
rect 16175 1050 16195 1070
rect 16175 1000 16195 1020
rect 16175 950 16195 970
rect 17630 1150 17650 1170
rect 17630 1100 17650 1120
rect 17630 1050 17650 1070
rect 17630 1000 17650 1020
rect 17630 950 17650 970
rect 17975 1170 17995 1190
rect 17975 1120 17995 1140
rect 17975 1070 17995 1090
rect 17975 1020 17995 1040
rect 17975 970 17995 990
rect 18655 1620 18675 1640
rect 18655 1570 18675 1590
rect 18655 1520 18675 1540
rect 18655 1470 18675 1490
rect 18655 1420 18675 1440
rect 18655 1370 18675 1390
rect 18655 1320 18675 1340
rect 18655 1270 18675 1290
rect 18655 1220 18675 1240
rect 18655 1170 18675 1190
rect 18655 1120 18675 1140
rect 18655 1070 18675 1090
rect 18655 1020 18675 1040
rect 18655 970 18675 990
rect 2965 845 2985 865
rect 2965 795 2985 815
rect 5025 845 5045 865
rect 5025 795 5045 815
rect 16850 715 16870 735
rect 17590 715 17610 735
<< nsubdiffcont >>
rect 2965 2895 2985 2915
rect 2965 2845 2985 2865
rect 5025 2895 5045 2915
rect 5025 2845 5045 2865
rect 3145 2665 3165 2685
rect 3145 2615 3165 2635
rect 3145 2565 3165 2585
rect 3145 2515 3165 2535
rect 3145 2465 3165 2485
rect 3145 2415 3165 2435
rect 4845 2665 4865 2685
rect 4845 2615 4865 2635
rect 4845 2565 4865 2585
rect 4845 2515 4865 2535
rect 4845 2465 4865 2485
rect 4845 2415 4865 2435
rect 3995 1965 4015 1985
rect 3995 1915 4015 1935
<< poly >>
rect 16632 4510 16668 4520
rect 16632 4490 16640 4510
rect 16660 4490 16668 4510
rect 16632 4480 16668 4490
rect 16752 4510 16788 4520
rect 16752 4490 16760 4510
rect 16780 4490 16788 4510
rect 16752 4480 16788 4490
rect 16872 4510 16908 4520
rect 16872 4490 16880 4510
rect 16900 4490 16908 4510
rect 16872 4480 16908 4490
rect 16570 4465 16610 4475
rect 16200 4450 16240 4460
rect 16200 4430 16210 4450
rect 16230 4430 16240 4450
rect 16460 4450 16500 4460
rect 16460 4430 16470 4450
rect 16490 4430 16500 4450
rect 16570 4445 16580 4465
rect 16600 4450 16610 4465
rect 16930 4465 16970 4475
rect 16930 4450 16940 4465
rect 16600 4445 16630 4450
rect 16570 4435 16630 4445
rect 16910 4445 16940 4450
rect 16960 4445 16970 4465
rect 16910 4435 16970 4445
rect 16200 4415 16300 4430
rect 16280 4403 16300 4415
rect 16340 4403 16360 4418
rect 16400 4415 16500 4430
rect 16610 4420 16630 4435
rect 16670 4420 16690 4435
rect 16730 4420 16750 4435
rect 16790 4420 16810 4435
rect 16850 4420 16870 4435
rect 16910 4420 16930 4435
rect 16400 4403 16420 4415
rect 17120 4395 17140 4410
rect 17180 4395 17200 4410
rect 17240 4395 17260 4410
rect 17300 4395 17320 4410
rect 17360 4395 17380 4410
rect 17420 4395 17440 4410
rect 17480 4395 17500 4410
rect 17540 4395 17560 4410
rect 16280 4325 16300 4340
rect 16340 4325 16360 4340
rect 16400 4325 16420 4340
rect 16610 4325 16630 4340
rect 16670 4330 16690 4340
rect 16730 4330 16750 4340
rect 16790 4330 16810 4340
rect 16850 4330 16870 4340
rect 16330 4315 16370 4325
rect 16670 4315 16870 4330
rect 16910 4325 16930 4340
rect 17120 4325 17140 4335
rect 17180 4325 17200 4335
rect 17240 4325 17260 4335
rect 17300 4325 17320 4335
rect 17360 4325 17380 4335
rect 17420 4325 17440 4335
rect 17480 4325 17500 4335
rect 17540 4325 17560 4335
rect 16330 4295 16340 4315
rect 16360 4295 16370 4315
rect 16330 4285 16370 4295
rect 16750 4310 16790 4315
rect 17120 4310 17560 4325
rect 16750 4290 16760 4310
rect 16780 4290 16790 4310
rect 16750 4280 16790 4290
rect 17203 4290 17211 4310
rect 17229 4290 17237 4310
rect 17203 4280 17237 4290
rect 16210 4200 16250 4210
rect 16210 4180 16220 4200
rect 16240 4180 16250 4200
rect 17500 4200 17540 4210
rect 17500 4180 17510 4200
rect 17530 4180 17540 4200
rect 16210 4165 16305 4180
rect 16290 4155 16305 4165
rect 16345 4155 16360 4170
rect 16400 4155 16415 4170
rect 16455 4155 16470 4170
rect 16510 4155 16525 4170
rect 16565 4155 16580 4170
rect 16620 4155 16635 4170
rect 16675 4155 16690 4170
rect 16730 4155 16745 4170
rect 16785 4155 16800 4170
rect 16840 4155 16855 4170
rect 16895 4155 16910 4170
rect 16950 4155 16965 4170
rect 17005 4155 17020 4170
rect 17060 4155 17075 4170
rect 17115 4155 17130 4170
rect 17170 4155 17185 4170
rect 17225 4155 17240 4170
rect 17280 4155 17295 4170
rect 17335 4155 17350 4170
rect 17390 4155 17405 4170
rect 17445 4165 17540 4180
rect 17445 4155 17460 4165
rect 16290 4090 16305 4105
rect 16345 4095 16360 4105
rect 16400 4095 16415 4105
rect 16455 4095 16470 4105
rect 16510 4095 16525 4105
rect 16565 4095 16580 4105
rect 16620 4095 16635 4105
rect 16675 4095 16690 4105
rect 16730 4095 16745 4105
rect 16785 4095 16800 4105
rect 16840 4095 16855 4105
rect 16895 4095 16910 4105
rect 16950 4095 16965 4105
rect 17005 4095 17020 4105
rect 17060 4095 17075 4105
rect 17115 4095 17130 4105
rect 17170 4095 17185 4105
rect 17225 4095 17240 4105
rect 17280 4095 17295 4105
rect 17335 4095 17350 4105
rect 17390 4095 17405 4105
rect 16345 4080 17405 4095
rect 17445 4090 17460 4105
rect 16362 4060 16370 4080
rect 16390 4060 16398 4080
rect 16362 4050 16398 4060
rect 16155 3895 16195 3905
rect 16155 3875 16165 3895
rect 16185 3875 16195 3895
rect 16271 3895 16303 3905
rect 16271 3875 16277 3895
rect 16294 3875 16303 3895
rect 16470 3895 16510 3905
rect 16470 3875 16480 3895
rect 16500 3875 16510 3895
rect 16690 3895 16730 3905
rect 16690 3875 16700 3895
rect 16720 3875 16730 3895
rect 16895 3895 16935 3905
rect 16895 3875 16905 3895
rect 16925 3875 16935 3895
rect 17011 3895 17043 3905
rect 17011 3875 17017 3895
rect 17034 3875 17043 3895
rect 17210 3895 17250 3905
rect 17210 3875 17220 3895
rect 17240 3875 17250 3895
rect 17430 3895 17470 3905
rect 17430 3875 17440 3895
rect 17460 3875 17470 3895
rect 17635 3895 17675 3905
rect 17635 3875 17645 3895
rect 17665 3875 17675 3895
rect 16155 3860 16250 3875
rect 16271 3865 16305 3875
rect 16235 3850 16250 3860
rect 16290 3850 16305 3865
rect 16345 3850 16360 3865
rect 16400 3850 16415 3865
rect 16455 3860 16525 3875
rect 16455 3850 16470 3860
rect 16510 3850 16525 3860
rect 16565 3850 16580 3865
rect 16620 3850 16635 3865
rect 16675 3860 16745 3875
rect 16675 3850 16690 3860
rect 16730 3850 16745 3860
rect 16785 3850 16800 3865
rect 16840 3860 16990 3875
rect 17011 3865 17045 3875
rect 16840 3850 16855 3860
rect 16975 3850 16990 3860
rect 17030 3850 17045 3865
rect 17085 3850 17100 3865
rect 17140 3850 17155 3865
rect 17195 3860 17265 3875
rect 17195 3850 17210 3860
rect 17250 3850 17265 3860
rect 17305 3850 17320 3865
rect 17360 3850 17375 3865
rect 17415 3860 17485 3875
rect 17415 3850 17430 3860
rect 17470 3850 17485 3860
rect 17525 3850 17540 3865
rect 17580 3860 17675 3875
rect 17580 3850 17595 3860
rect 16235 3785 16250 3800
rect 16290 3785 16305 3800
rect 16345 3790 16360 3800
rect 16400 3790 16415 3800
rect 16345 3785 16415 3790
rect 16455 3785 16470 3800
rect 16510 3785 16525 3800
rect 16565 3790 16580 3800
rect 16620 3790 16635 3800
rect 16565 3785 16635 3790
rect 16675 3785 16690 3800
rect 16730 3785 16745 3800
rect 16785 3785 16800 3800
rect 16840 3785 16855 3800
rect 16975 3785 16990 3800
rect 17030 3785 17045 3800
rect 17085 3790 17100 3800
rect 17140 3790 17155 3800
rect 17085 3785 17155 3790
rect 17195 3785 17210 3800
rect 17250 3785 17265 3800
rect 17305 3790 17320 3800
rect 17360 3790 17375 3800
rect 17305 3785 17375 3790
rect 17415 3785 17430 3800
rect 17470 3785 17485 3800
rect 17525 3785 17540 3800
rect 17580 3785 17595 3800
rect 16345 3775 16434 3785
rect 16565 3775 16654 3785
rect 16402 3755 16408 3775
rect 16425 3755 16434 3775
rect 16402 3745 16434 3755
rect 16622 3755 16628 3775
rect 16645 3755 16654 3775
rect 16622 3745 16654 3755
rect 16766 3775 16800 3785
rect 17085 3775 17174 3785
rect 17305 3775 17394 3785
rect 16766 3755 16775 3775
rect 16792 3755 16800 3775
rect 16766 3745 16800 3755
rect 17142 3755 17148 3775
rect 17165 3755 17174 3775
rect 17142 3745 17174 3755
rect 17362 3755 17368 3775
rect 17385 3755 17394 3775
rect 17362 3745 17394 3755
rect 17506 3775 17540 3785
rect 17506 3755 17515 3775
rect 17532 3755 17540 3775
rect 17506 3745 17540 3755
rect 16180 3620 16220 3630
rect 16180 3600 16190 3620
rect 16210 3600 16220 3620
rect 17580 3620 17620 3630
rect 17580 3600 17590 3620
rect 17610 3600 17620 3620
rect 15195 3585 15210 3600
rect 15250 3585 15265 3600
rect 15305 3585 15320 3600
rect 15360 3585 15375 3600
rect 15415 3585 15430 3600
rect 15470 3585 15485 3600
rect 15525 3585 15540 3600
rect 15580 3585 15595 3600
rect 15635 3585 15650 3600
rect 15690 3585 15705 3600
rect 15745 3585 15760 3600
rect 15800 3585 15815 3600
rect 16180 3585 16280 3600
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 3035 2930 3085 2945
rect 3125 2930 3175 2945
rect 3215 2930 3265 2945
rect 3305 2930 3355 2945
rect 3395 2930 3445 2945
rect 3485 2930 3535 2945
rect 3575 2930 3625 2945
rect 3665 2930 3715 2945
rect 3755 2930 3805 2945
rect 3845 2930 3895 2945
rect 3935 2930 3985 2945
rect 4025 2930 4075 2945
rect 4115 2930 4165 2945
rect 4205 2930 4255 2945
rect 4295 2930 4345 2945
rect 4385 2930 4435 2945
rect 4475 2930 4525 2945
rect 4565 2930 4615 2945
rect 4655 2930 4705 2945
rect 4745 2930 4795 2945
rect 4835 2930 4885 2945
rect 4925 2930 4975 2945
rect 16260 3575 16280 3585
rect 16320 3575 16340 3590
rect 16380 3575 16400 3590
rect 16440 3575 16460 3590
rect 16500 3575 16520 3590
rect 16560 3575 16580 3590
rect 16620 3575 16640 3590
rect 16680 3575 16700 3590
rect 16740 3575 16760 3590
rect 16800 3575 16820 3590
rect 16860 3575 16880 3590
rect 16920 3575 16940 3590
rect 16980 3575 17000 3590
rect 17040 3575 17060 3590
rect 17100 3575 17120 3590
rect 17160 3575 17180 3590
rect 17220 3575 17240 3590
rect 17280 3575 17300 3590
rect 17340 3575 17360 3590
rect 17400 3575 17420 3590
rect 17460 3575 17480 3590
rect 17520 3585 17620 3600
rect 17985 3585 18000 3600
rect 18040 3585 18055 3600
rect 18095 3585 18110 3600
rect 18150 3585 18165 3600
rect 18205 3585 18220 3600
rect 18260 3585 18275 3600
rect 18315 3585 18330 3600
rect 18370 3585 18385 3600
rect 18425 3585 18440 3600
rect 18480 3585 18495 3600
rect 18535 3585 18550 3600
rect 18590 3585 18605 3600
rect 17520 3575 17540 3585
rect 16260 3160 16280 3175
rect 16320 3165 16340 3175
rect 16380 3165 16400 3175
rect 16440 3165 16460 3175
rect 16500 3165 16520 3175
rect 16560 3165 16580 3175
rect 16620 3165 16640 3175
rect 16680 3165 16700 3175
rect 16740 3165 16760 3175
rect 16800 3165 16820 3175
rect 16860 3165 16880 3175
rect 16920 3165 16940 3175
rect 16980 3165 17000 3175
rect 17040 3165 17060 3175
rect 17100 3165 17120 3175
rect 17160 3165 17180 3175
rect 17220 3165 17240 3175
rect 17280 3165 17300 3175
rect 17340 3165 17360 3175
rect 17400 3165 17420 3175
rect 17460 3165 17480 3175
rect 16320 3150 17480 3165
rect 17520 3160 17540 3175
rect 16823 3130 16831 3150
rect 16849 3130 16857 3150
rect 16823 3120 16857 3130
rect 15195 2975 15210 2985
rect 15115 2960 15210 2975
rect 15250 2975 15265 2985
rect 15305 2975 15320 2985
rect 15360 2975 15375 2985
rect 15415 2975 15430 2985
rect 15470 2975 15485 2985
rect 15525 2975 15540 2985
rect 15580 2975 15595 2985
rect 15635 2975 15650 2985
rect 15690 2975 15705 2985
rect 15745 2975 15760 2985
rect 15250 2960 15760 2975
rect 15800 2975 15815 2985
rect 17985 2975 18000 2985
rect 15800 2960 15895 2975
rect 15115 2940 15125 2960
rect 15145 2940 15155 2960
rect 15115 2930 15155 2940
rect 15653 2940 15661 2960
rect 15679 2940 15687 2960
rect 15653 2930 15687 2940
rect 15855 2940 15865 2960
rect 15885 2940 15895 2960
rect 17905 2960 18000 2975
rect 18040 2975 18055 2985
rect 18095 2975 18110 2985
rect 18150 2975 18165 2985
rect 18205 2975 18220 2985
rect 18260 2975 18275 2985
rect 18315 2975 18330 2985
rect 18370 2975 18385 2985
rect 18425 2975 18440 2985
rect 18480 2975 18495 2985
rect 18535 2975 18550 2985
rect 18040 2960 18550 2975
rect 18590 2975 18605 2985
rect 18590 2960 18685 2975
rect 15855 2930 15895 2940
rect 16180 2940 16220 2950
rect 16180 2920 16190 2940
rect 16210 2920 16220 2940
rect 17580 2940 17620 2950
rect 17580 2920 17590 2940
rect 17610 2920 17620 2940
rect 17905 2940 17915 2960
rect 17935 2940 17945 2960
rect 17905 2930 17945 2940
rect 18113 2940 18121 2960
rect 18139 2940 18147 2960
rect 18113 2930 18147 2940
rect 18645 2940 18655 2960
rect 18675 2940 18685 2960
rect 18645 2930 18685 2940
rect 16180 2905 16280 2920
rect 16260 2895 16280 2905
rect 16320 2895 16340 2910
rect 16380 2895 16400 2910
rect 16440 2895 16460 2910
rect 16500 2895 16520 2910
rect 16560 2895 16580 2910
rect 16620 2895 16640 2910
rect 16680 2895 16700 2910
rect 16740 2895 16760 2910
rect 16800 2895 16820 2910
rect 16860 2895 16880 2910
rect 16920 2895 16940 2910
rect 16980 2895 17000 2910
rect 17040 2895 17060 2910
rect 17100 2895 17120 2910
rect 17160 2895 17180 2910
rect 17220 2895 17240 2910
rect 17280 2895 17300 2910
rect 17340 2895 17360 2910
rect 17400 2895 17420 2910
rect 17460 2895 17480 2910
rect 17520 2905 17620 2920
rect 17520 2895 17540 2905
rect 3035 2815 3085 2830
rect 2995 2805 3085 2815
rect 3125 2820 3175 2830
rect 3215 2820 3265 2830
rect 3305 2820 3355 2830
rect 3395 2820 3445 2830
rect 3485 2820 3535 2830
rect 3575 2820 3625 2830
rect 3665 2820 3715 2830
rect 3755 2820 3805 2830
rect 3845 2820 3895 2830
rect 3935 2820 3985 2830
rect 4025 2820 4075 2830
rect 4115 2820 4165 2830
rect 4205 2820 4255 2830
rect 4295 2820 4345 2830
rect 4385 2820 4435 2830
rect 4475 2820 4525 2830
rect 4565 2820 4615 2830
rect 4655 2820 4705 2830
rect 4745 2820 4795 2830
rect 4835 2820 4885 2830
rect 3125 2805 4885 2820
rect 4925 2815 4975 2830
rect 4925 2805 5015 2815
rect 2995 2785 3005 2805
rect 3025 2800 3085 2805
rect 4925 2800 4985 2805
rect 3025 2785 3035 2800
rect 2995 2775 3035 2785
rect 4975 2785 4985 2800
rect 5005 2785 5015 2805
rect 4975 2775 5015 2785
rect 3175 2745 3215 2755
rect 3175 2725 3185 2745
rect 3205 2730 3215 2745
rect 4795 2745 4835 2755
rect 4795 2730 4805 2745
rect 3205 2725 3265 2730
rect 3175 2715 3265 2725
rect 4745 2725 4805 2730
rect 4825 2725 4835 2745
rect 4745 2715 4835 2725
rect 3215 2700 3265 2715
rect 3305 2700 3355 2715
rect 3395 2700 3445 2715
rect 3485 2700 3535 2715
rect 3575 2700 3625 2715
rect 3665 2700 3715 2715
rect 3755 2700 3805 2715
rect 3845 2700 3895 2715
rect 3935 2700 3985 2715
rect 4025 2700 4075 2715
rect 4115 2700 4165 2715
rect 4205 2700 4255 2715
rect 4295 2700 4345 2715
rect 4385 2700 4435 2715
rect 4475 2700 4525 2715
rect 4565 2700 4615 2715
rect 4655 2700 4705 2715
rect 4745 2700 4795 2715
rect 15195 2655 15210 2670
rect 15250 2655 15265 2670
rect 15305 2655 15320 2670
rect 15360 2655 15375 2670
rect 15415 2655 15430 2670
rect 15470 2655 15485 2670
rect 15525 2655 15540 2670
rect 15580 2655 15595 2670
rect 15635 2655 15650 2670
rect 15690 2655 15705 2670
rect 15745 2655 15760 2670
rect 15800 2655 15815 2670
rect 3215 2385 3265 2400
rect 3305 2390 3355 2400
rect 3395 2390 3445 2400
rect 3485 2390 3535 2400
rect 3575 2390 3625 2400
rect 3665 2390 3715 2400
rect 3755 2390 3805 2400
rect 3845 2390 3895 2400
rect 3935 2390 3985 2400
rect 4025 2390 4075 2400
rect 4115 2390 4165 2400
rect 4205 2390 4255 2400
rect 4295 2390 4345 2400
rect 4385 2390 4435 2400
rect 4475 2390 4525 2400
rect 4565 2390 4615 2400
rect 4655 2390 4705 2400
rect 3305 2375 4705 2390
rect 4745 2385 4795 2400
rect 3355 2370 3395 2375
rect 3355 2350 3365 2370
rect 3385 2350 3395 2370
rect 3355 2340 3395 2350
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 2605 2000 2620 2015
rect 2660 2000 2675 2015
rect 2785 2000 2805 2015
rect 2845 2000 2865 2015
rect 2905 2000 2925 2015
rect 2965 2000 2985 2015
rect 3025 2000 3045 2015
rect 3085 2000 3105 2015
rect 3145 2000 3165 2015
rect 3205 2000 3225 2015
rect 3265 2000 3285 2015
rect 3325 2000 3345 2015
rect 3385 2000 3405 2015
rect 3445 2000 3465 2015
rect 3505 2000 3525 2015
rect 3565 2000 3585 2015
rect 3625 2000 3645 2015
rect 3685 2000 3705 2015
rect 3745 2000 3765 2015
rect 3805 2000 3825 2015
rect 3865 2000 3885 2015
rect 3925 2000 3945 2015
rect 4065 2000 4085 2015
rect 4125 2000 4145 2015
rect 4185 2000 4205 2015
rect 4245 2000 4265 2015
rect 4305 2000 4325 2015
rect 4365 2000 4385 2015
rect 4425 2000 4445 2015
rect 4485 2000 4505 2015
rect 4545 2000 4565 2015
rect 4605 2000 4625 2015
rect 4665 2000 4685 2015
rect 4725 2000 4745 2015
rect 4785 2000 4805 2015
rect 4845 2000 4865 2015
rect 4905 2000 4925 2015
rect 4965 2000 4985 2015
rect 5025 2000 5045 2015
rect 5085 2000 5105 2015
rect 5145 2000 5165 2015
rect 5205 2000 5225 2015
rect 17985 2655 18000 2670
rect 18040 2655 18055 2670
rect 18095 2655 18110 2670
rect 18150 2655 18165 2670
rect 18205 2655 18220 2670
rect 18260 2655 18275 2670
rect 18315 2655 18330 2670
rect 18370 2655 18385 2670
rect 18425 2655 18440 2670
rect 18480 2655 18495 2670
rect 18535 2655 18550 2670
rect 18590 2655 18605 2670
rect 16260 2480 16280 2495
rect 16320 2485 16340 2495
rect 16380 2485 16400 2495
rect 16440 2485 16460 2495
rect 16500 2485 16520 2495
rect 16560 2485 16580 2495
rect 16620 2485 16640 2495
rect 16680 2485 16700 2495
rect 16740 2485 16760 2495
rect 16800 2485 16820 2495
rect 16860 2485 16880 2495
rect 16920 2485 16940 2495
rect 16980 2485 17000 2495
rect 17040 2485 17060 2495
rect 17100 2485 17120 2495
rect 17160 2485 17180 2495
rect 17220 2485 17240 2495
rect 17280 2485 17300 2495
rect 17340 2485 17360 2495
rect 17400 2485 17420 2495
rect 17460 2485 17480 2495
rect 16320 2470 17480 2485
rect 17520 2480 17540 2495
rect 15195 2445 15210 2455
rect 15115 2430 15210 2445
rect 15250 2445 15265 2455
rect 15305 2445 15320 2455
rect 15360 2445 15375 2455
rect 15415 2445 15430 2455
rect 15470 2445 15485 2455
rect 15525 2445 15540 2455
rect 15580 2445 15595 2455
rect 15635 2445 15650 2455
rect 15690 2445 15705 2455
rect 15745 2445 15760 2455
rect 15250 2430 15760 2445
rect 15800 2445 15815 2455
rect 16823 2450 16831 2470
rect 16849 2450 16857 2470
rect 15800 2430 15895 2445
rect 16823 2440 16857 2450
rect 17985 2445 18000 2455
rect 15115 2410 15125 2430
rect 15145 2410 15155 2430
rect 15115 2400 15155 2410
rect 15745 2395 15760 2430
rect 15855 2410 15865 2430
rect 15885 2410 15895 2430
rect 15855 2400 15895 2410
rect 17905 2430 18000 2445
rect 18040 2445 18055 2455
rect 18095 2445 18110 2455
rect 18150 2445 18165 2455
rect 18205 2445 18220 2455
rect 18260 2445 18275 2455
rect 18315 2445 18330 2455
rect 18370 2445 18385 2455
rect 18425 2445 18440 2455
rect 18480 2445 18495 2455
rect 18535 2445 18550 2455
rect 18040 2430 18550 2445
rect 18590 2445 18605 2455
rect 18590 2430 18685 2445
rect 17905 2410 17915 2430
rect 17935 2410 17945 2430
rect 17905 2400 17945 2410
rect 15745 2385 15805 2395
rect 15745 2365 15775 2385
rect 15795 2365 15805 2385
rect 18040 2380 18055 2430
rect 18645 2410 18655 2430
rect 18675 2410 18685 2430
rect 18645 2400 18685 2410
rect 15745 2355 15805 2365
rect 18025 2370 18065 2380
rect 15115 2310 15155 2320
rect 15115 2290 15125 2310
rect 15145 2290 15155 2310
rect 15745 2290 15760 2355
rect 18025 2350 18035 2370
rect 18055 2350 18065 2370
rect 18025 2340 18065 2350
rect 15855 2310 15895 2320
rect 15855 2290 15865 2310
rect 15885 2290 15895 2310
rect 15115 2275 15210 2290
rect 15195 2265 15210 2275
rect 15250 2275 15760 2290
rect 15250 2265 15265 2275
rect 15305 2265 15320 2275
rect 15360 2265 15375 2275
rect 15415 2265 15430 2275
rect 15470 2265 15485 2275
rect 15525 2265 15540 2275
rect 15580 2265 15595 2275
rect 15635 2265 15650 2275
rect 15690 2265 15705 2275
rect 15745 2265 15760 2275
rect 15800 2275 15895 2290
rect 17905 2310 17945 2320
rect 17905 2290 17915 2310
rect 17935 2290 17945 2310
rect 18040 2290 18055 2340
rect 18645 2310 18685 2320
rect 18645 2290 18655 2310
rect 18675 2290 18685 2310
rect 17905 2275 18000 2290
rect 15800 2265 15815 2275
rect 17985 2265 18000 2275
rect 18040 2275 18550 2290
rect 18040 2265 18055 2275
rect 18095 2265 18110 2275
rect 18150 2265 18165 2275
rect 18205 2265 18220 2275
rect 18260 2265 18275 2275
rect 18315 2265 18330 2275
rect 18370 2265 18385 2275
rect 18425 2265 18440 2275
rect 18480 2265 18495 2275
rect 18535 2265 18550 2275
rect 18590 2275 18685 2290
rect 18590 2265 18605 2275
rect 16828 2175 16862 2185
rect 16828 2155 16836 2175
rect 16854 2155 16862 2175
rect 16315 2130 16330 2145
rect 16370 2140 17430 2155
rect 16370 2130 16385 2140
rect 16425 2130 16440 2140
rect 16480 2130 16495 2140
rect 16535 2130 16550 2140
rect 16590 2130 16605 2140
rect 16645 2130 16660 2140
rect 16700 2130 16715 2140
rect 16755 2130 16770 2140
rect 16810 2130 16825 2140
rect 16865 2130 16880 2140
rect 16920 2130 16935 2140
rect 16975 2130 16990 2140
rect 17030 2130 17045 2140
rect 17085 2130 17100 2140
rect 17140 2130 17155 2140
rect 17195 2130 17210 2140
rect 17250 2130 17265 2140
rect 17305 2130 17320 2140
rect 17360 2130 17375 2140
rect 17415 2130 17430 2140
rect 17470 2130 17485 2145
rect 16315 1970 16330 1980
rect 15195 1950 15210 1965
rect 15250 1950 15265 1965
rect 15305 1950 15320 1965
rect 15360 1950 15375 1965
rect 15415 1950 15430 1965
rect 15470 1950 15485 1965
rect 15525 1950 15540 1965
rect 15580 1950 15595 1965
rect 15635 1950 15650 1965
rect 15690 1950 15705 1965
rect 15745 1950 15760 1965
rect 15800 1950 15815 1965
rect 16235 1955 16330 1970
rect 16370 1965 16385 1980
rect 16425 1965 16440 1980
rect 16480 1965 16495 1980
rect 16535 1965 16550 1980
rect 16590 1965 16605 1980
rect 16645 1965 16660 1980
rect 16700 1965 16715 1980
rect 16755 1965 16770 1980
rect 16810 1965 16825 1980
rect 16865 1965 16880 1980
rect 16920 1965 16935 1980
rect 16975 1965 16990 1980
rect 17030 1965 17045 1980
rect 17085 1965 17100 1980
rect 17140 1965 17155 1980
rect 17195 1965 17210 1980
rect 17250 1965 17265 1980
rect 17305 1965 17320 1980
rect 17360 1965 17375 1980
rect 17415 1965 17430 1980
rect 17470 1970 17485 1980
rect 17470 1955 17565 1970
rect 16235 1935 16245 1955
rect 16265 1935 16275 1955
rect 16235 1925 16275 1935
rect 17525 1935 17535 1955
rect 17555 1935 17565 1955
rect 17985 1950 18000 1965
rect 18040 1950 18055 1965
rect 18095 1950 18110 1965
rect 18150 1950 18165 1965
rect 18205 1950 18220 1965
rect 18260 1950 18275 1965
rect 18315 1950 18330 1965
rect 18370 1950 18385 1965
rect 18425 1950 18440 1965
rect 18480 1950 18495 1965
rect 18535 1950 18550 1965
rect 18590 1950 18605 1965
rect 17525 1925 17565 1935
rect 2605 1890 2620 1900
rect 2660 1890 2675 1900
rect 2605 1875 2675 1890
rect 2785 1885 2805 1900
rect 2845 1885 2865 1900
rect 2905 1890 2925 1900
rect 2965 1890 2985 1900
rect 3025 1890 3045 1900
rect 3085 1890 3105 1900
rect 2765 1875 2805 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2765 1855 2775 1875
rect 2795 1855 2805 1875
rect 2765 1845 2805 1855
rect 2835 1875 2875 1885
rect 2905 1875 3105 1890
rect 3145 1890 3165 1900
rect 3205 1890 3225 1900
rect 3145 1875 3225 1890
rect 3265 1890 3285 1900
rect 3325 1890 3345 1900
rect 3385 1890 3405 1900
rect 3445 1890 3465 1900
rect 3265 1875 3465 1890
rect 3505 1890 3525 1900
rect 3565 1890 3585 1900
rect 3505 1875 3585 1890
rect 3625 1890 3645 1900
rect 3685 1890 3705 1900
rect 3745 1890 3765 1900
rect 3805 1890 3825 1900
rect 3625 1875 3825 1890
rect 3865 1885 3885 1900
rect 3925 1890 3945 1900
rect 4065 1890 4085 1900
rect 3855 1875 3895 1885
rect 3925 1875 4085 1890
rect 4125 1885 4145 1900
rect 4185 1890 4205 1900
rect 4245 1890 4265 1900
rect 4305 1890 4325 1900
rect 4365 1890 4385 1900
rect 4115 1875 4155 1885
rect 4185 1875 4385 1890
rect 4425 1890 4445 1900
rect 4485 1890 4505 1900
rect 4425 1875 4505 1890
rect 4545 1890 4565 1900
rect 4605 1890 4625 1900
rect 4665 1890 4685 1900
rect 4725 1890 4745 1900
rect 4545 1875 4745 1890
rect 4785 1890 4805 1900
rect 4845 1890 4865 1900
rect 4785 1875 4865 1890
rect 4905 1890 4925 1900
rect 4965 1890 4985 1900
rect 5025 1890 5045 1900
rect 5085 1890 5105 1900
rect 4905 1875 5105 1890
rect 5145 1885 5165 1900
rect 5205 1885 5225 1900
rect 5135 1875 5175 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1855 2935 1875
rect 2955 1855 2965 1875
rect 2925 1845 2965 1855
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1855 3295 1875
rect 3315 1855 3325 1875
rect 3285 1845 3325 1855
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1855 3655 1875
rect 3675 1855 3685 1875
rect 3645 1845 3685 1855
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 3985 1870 4025 1875
rect 3985 1850 3995 1870
rect 4015 1850 4025 1870
rect 3985 1840 4025 1850
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4325 1855 4335 1875
rect 4355 1855 4365 1875
rect 4325 1845 4365 1855
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4685 1855 4695 1875
rect 4715 1855 4725 1875
rect 4685 1845 4725 1855
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 5045 1855 5055 1875
rect 5075 1855 5085 1875
rect 5045 1845 5085 1855
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 5205 1875 5245 1885
rect 5205 1855 5215 1875
rect 5235 1855 5245 1875
rect 5205 1845 5245 1855
rect 3225 1755 3265 1765
rect 3225 1735 3235 1755
rect 3255 1735 3265 1755
rect 3225 1720 3265 1735
rect 4745 1755 4785 1765
rect 4745 1735 4755 1755
rect 4775 1735 4785 1755
rect 4745 1720 4785 1735
rect 3225 1705 3765 1720
rect 3205 1665 3225 1680
rect 3265 1665 3285 1705
rect 3325 1665 3345 1705
rect 3385 1665 3405 1680
rect 3445 1665 3465 1680
rect 3505 1665 3525 1705
rect 3565 1665 3585 1705
rect 3625 1665 3645 1680
rect 3685 1665 3705 1680
rect 3745 1665 3765 1705
rect 4245 1705 4785 1720
rect 16237 1710 16269 1720
rect 4245 1665 4265 1705
rect 4305 1665 4325 1680
rect 4365 1665 4385 1680
rect 4425 1665 4445 1705
rect 4485 1665 4505 1705
rect 4545 1665 4565 1680
rect 4605 1665 4625 1680
rect 4665 1665 4685 1705
rect 4725 1665 4745 1705
rect 15558 1700 15592 1710
rect 15558 1680 15566 1700
rect 15584 1680 15592 1700
rect 16237 1690 16243 1710
rect 16260 1690 16269 1710
rect 16457 1710 16489 1720
rect 16457 1690 16463 1710
rect 16480 1690 16489 1710
rect 16180 1680 16269 1690
rect 16400 1680 16489 1690
rect 16601 1710 16635 1720
rect 16601 1690 16610 1710
rect 16627 1690 16635 1710
rect 16867 1710 16899 1720
rect 16867 1695 16876 1710
rect 16601 1680 16635 1690
rect 16865 1690 16876 1695
rect 16893 1690 16899 1710
rect 17277 1710 17309 1720
rect 17277 1690 17283 1710
rect 17300 1690 17309 1710
rect 17497 1710 17529 1720
rect 17497 1690 17503 1710
rect 17520 1690 17529 1710
rect 16865 1680 16899 1690
rect 17220 1680 17309 1690
rect 17440 1680 17529 1690
rect 17641 1710 17675 1720
rect 17641 1690 17650 1710
rect 17667 1690 17675 1710
rect 17641 1680 17675 1690
rect 18208 1700 18242 1710
rect 18208 1680 18216 1700
rect 18234 1680 18242 1700
rect 4785 1665 4805 1680
rect 15195 1655 15255 1670
rect 15295 1665 15655 1680
rect 15295 1655 15355 1665
rect 15395 1655 15455 1665
rect 15495 1655 15555 1665
rect 15595 1655 15655 1665
rect 15695 1655 15755 1670
rect 16070 1665 16085 1680
rect 16125 1665 16140 1680
rect 16180 1675 16250 1680
rect 16180 1665 16195 1675
rect 16235 1665 16250 1675
rect 16290 1665 16305 1680
rect 16345 1665 16360 1680
rect 16400 1675 16470 1680
rect 16400 1665 16415 1675
rect 16455 1665 16470 1675
rect 16510 1665 16525 1680
rect 16565 1665 16580 1680
rect 16620 1665 16635 1680
rect 16675 1665 16690 1680
rect 16810 1665 16825 1680
rect 16865 1665 16880 1680
rect 16920 1665 16935 1680
rect 16975 1665 16990 1680
rect 17110 1665 17125 1680
rect 17165 1665 17180 1680
rect 17220 1675 17290 1680
rect 17220 1665 17235 1675
rect 17275 1665 17290 1675
rect 17330 1665 17345 1680
rect 17385 1665 17400 1680
rect 17440 1675 17510 1680
rect 17440 1665 17455 1675
rect 17495 1665 17510 1675
rect 17550 1665 17565 1680
rect 17605 1665 17620 1680
rect 17660 1665 17675 1680
rect 17715 1665 17730 1680
rect 3205 1600 3225 1615
rect 3265 1600 3285 1615
rect 3325 1600 3345 1615
rect 3165 1590 3225 1600
rect 3165 1570 3175 1590
rect 3195 1575 3225 1590
rect 3385 1575 3405 1615
rect 3445 1575 3465 1615
rect 3505 1600 3525 1615
rect 3565 1600 3585 1615
rect 3625 1575 3645 1615
rect 3685 1575 3705 1615
rect 3745 1600 3765 1615
rect 4245 1600 4265 1615
rect 3195 1570 3705 1575
rect 3165 1560 3705 1570
rect 4305 1575 4325 1615
rect 4365 1575 4385 1615
rect 4425 1600 4445 1615
rect 4485 1600 4505 1615
rect 4545 1575 4565 1615
rect 4605 1575 4625 1615
rect 4665 1600 4685 1615
rect 4725 1600 4745 1615
rect 4785 1600 4805 1615
rect 4785 1590 4845 1600
rect 4785 1575 4815 1590
rect 4305 1570 4815 1575
rect 4835 1570 4845 1590
rect 4305 1560 4845 1570
rect 2925 1495 2965 1505
rect 2925 1475 2935 1495
rect 2955 1475 2965 1495
rect 2925 1470 2965 1475
rect 3045 1495 3085 1505
rect 3045 1475 3055 1495
rect 3075 1475 3085 1495
rect 3045 1470 3085 1475
rect 3165 1495 3205 1505
rect 3165 1475 3175 1495
rect 3195 1475 3205 1495
rect 3165 1470 3205 1475
rect 3285 1495 3325 1505
rect 3285 1475 3295 1495
rect 3315 1475 3325 1495
rect 3285 1470 3325 1475
rect 3525 1495 3565 1505
rect 3525 1475 3535 1495
rect 3555 1475 3565 1495
rect 3525 1470 3565 1475
rect 3645 1495 3685 1505
rect 3645 1475 3655 1495
rect 3675 1475 3685 1495
rect 3645 1470 3685 1475
rect 3765 1495 3805 1505
rect 3765 1475 3775 1495
rect 3795 1475 3805 1495
rect 3765 1470 3805 1475
rect 4205 1495 4245 1505
rect 4205 1475 4215 1495
rect 4235 1475 4245 1495
rect 4205 1470 4245 1475
rect 4325 1495 4365 1505
rect 4325 1475 4335 1495
rect 4355 1475 4365 1495
rect 4325 1470 4365 1475
rect 4445 1495 4485 1505
rect 4445 1475 4455 1495
rect 4475 1475 4485 1495
rect 4445 1470 4485 1475
rect 4685 1495 4725 1505
rect 4685 1475 4695 1495
rect 4715 1475 4725 1495
rect 4685 1470 4725 1475
rect 4805 1495 4845 1505
rect 4805 1475 4815 1495
rect 4835 1475 4845 1495
rect 4805 1470 4845 1475
rect 4925 1495 4965 1505
rect 4925 1475 4935 1495
rect 4955 1475 4965 1495
rect 4925 1470 4965 1475
rect 5045 1495 5085 1505
rect 5045 1475 5055 1495
rect 5075 1475 5085 1495
rect 5045 1470 5085 1475
rect 2875 1455 3375 1470
rect 3415 1455 3915 1470
rect 4095 1455 4595 1470
rect 4635 1455 5135 1470
rect 2875 1190 3375 1205
rect 3415 1190 3915 1205
rect 4095 1190 4595 1205
rect 4635 1190 5135 1205
rect 3025 1120 3065 1130
rect 3025 1100 3035 1120
rect 3055 1100 3065 1120
rect 3025 1090 3065 1100
rect 3105 1120 3145 1130
rect 3105 1100 3115 1120
rect 3135 1100 3145 1120
rect 3105 1090 3145 1100
rect 3185 1120 3225 1130
rect 3185 1100 3195 1120
rect 3215 1100 3225 1120
rect 3185 1090 3225 1100
rect 3265 1120 3305 1130
rect 3265 1100 3275 1120
rect 3295 1100 3305 1120
rect 3265 1090 3305 1100
rect 3345 1120 3385 1130
rect 3345 1100 3355 1120
rect 3375 1100 3385 1120
rect 3345 1090 3385 1100
rect 3425 1120 3465 1130
rect 3425 1100 3435 1120
rect 3455 1100 3465 1120
rect 3425 1090 3465 1100
rect 3505 1120 3545 1130
rect 3505 1100 3515 1120
rect 3535 1100 3545 1120
rect 3505 1090 3545 1100
rect 3585 1120 3625 1130
rect 3585 1100 3595 1120
rect 3615 1100 3625 1120
rect 3585 1090 3625 1100
rect 3665 1120 3705 1130
rect 3665 1100 3675 1120
rect 3695 1100 3705 1120
rect 3665 1090 3705 1100
rect 3745 1120 3785 1130
rect 3745 1100 3755 1120
rect 3775 1100 3785 1120
rect 3745 1090 3785 1100
rect 3825 1120 3865 1130
rect 3825 1100 3835 1120
rect 3855 1100 3865 1120
rect 3825 1090 3865 1100
rect 3905 1120 3945 1130
rect 3905 1100 3915 1120
rect 3935 1100 3945 1120
rect 3905 1090 3945 1100
rect 4065 1120 4105 1130
rect 4065 1100 4075 1120
rect 4095 1100 4105 1120
rect 4065 1090 4105 1100
rect 4145 1120 4185 1130
rect 4145 1100 4155 1120
rect 4175 1100 4185 1120
rect 4145 1090 4185 1100
rect 4225 1120 4265 1130
rect 4225 1100 4235 1120
rect 4255 1100 4265 1120
rect 4225 1090 4265 1100
rect 4305 1120 4345 1130
rect 4305 1100 4315 1120
rect 4335 1100 4345 1120
rect 4305 1090 4345 1100
rect 4385 1120 4425 1130
rect 4385 1100 4395 1120
rect 4415 1100 4425 1120
rect 4385 1090 4425 1100
rect 4465 1120 4505 1130
rect 4465 1100 4475 1120
rect 4495 1100 4505 1120
rect 4465 1090 4505 1100
rect 4545 1120 4585 1130
rect 4545 1100 4555 1120
rect 4575 1100 4585 1120
rect 4545 1090 4585 1100
rect 4625 1120 4665 1130
rect 4625 1100 4635 1120
rect 4655 1100 4665 1120
rect 4625 1090 4665 1100
rect 4705 1120 4745 1130
rect 4705 1100 4715 1120
rect 4735 1100 4745 1120
rect 4705 1090 4745 1100
rect 4785 1120 4825 1130
rect 4785 1100 4795 1120
rect 4815 1100 4825 1120
rect 4785 1090 4825 1100
rect 4865 1120 4905 1130
rect 4865 1100 4875 1120
rect 4895 1100 4905 1120
rect 4865 1090 4905 1100
rect 4945 1120 4985 1130
rect 4945 1100 4955 1120
rect 4975 1100 4985 1120
rect 4945 1090 4985 1100
rect 2985 1075 3985 1090
rect 4025 1075 5025 1090
rect 2985 960 3985 975
rect 4025 960 5025 975
rect 2995 925 3035 935
rect 2995 905 3005 925
rect 3025 905 3035 925
rect 4975 925 5015 935
rect 4975 905 4985 925
rect 5005 905 5015 925
rect 18045 1655 18105 1670
rect 18145 1665 18505 1680
rect 18145 1655 18205 1665
rect 18245 1655 18305 1665
rect 18345 1655 18405 1665
rect 18445 1655 18505 1665
rect 18545 1655 18605 1670
rect 16070 1505 16085 1515
rect 15990 1490 16085 1505
rect 16125 1500 16140 1515
rect 16180 1500 16195 1515
rect 16235 1500 16250 1515
rect 16290 1505 16305 1515
rect 16345 1505 16360 1515
rect 16106 1490 16140 1500
rect 16290 1490 16360 1505
rect 16400 1500 16415 1515
rect 16455 1500 16470 1515
rect 16510 1505 16525 1515
rect 16565 1505 16580 1515
rect 16510 1490 16580 1505
rect 16620 1500 16635 1515
rect 16675 1505 16690 1515
rect 16810 1505 16825 1515
rect 16675 1490 16825 1505
rect 16865 1500 16880 1515
rect 16920 1500 16935 1515
rect 16975 1505 16990 1515
rect 17110 1505 17125 1515
rect 16920 1490 16954 1500
rect 16975 1490 17125 1505
rect 17165 1500 17180 1515
rect 17220 1500 17235 1515
rect 17275 1500 17290 1515
rect 17330 1505 17345 1515
rect 17385 1505 17400 1515
rect 17146 1490 17180 1500
rect 17330 1490 17400 1505
rect 17440 1500 17455 1515
rect 17495 1500 17510 1515
rect 17550 1505 17565 1515
rect 17605 1505 17620 1515
rect 17550 1490 17620 1505
rect 17660 1500 17675 1515
rect 17715 1505 17730 1515
rect 17715 1490 17810 1505
rect 15990 1470 16000 1490
rect 16020 1470 16030 1490
rect 15990 1460 16030 1470
rect 16106 1470 16112 1490
rect 16129 1470 16138 1490
rect 16106 1460 16138 1470
rect 16305 1470 16315 1490
rect 16335 1470 16345 1490
rect 16305 1460 16345 1470
rect 16525 1470 16535 1490
rect 16555 1470 16565 1490
rect 16525 1460 16565 1470
rect 16730 1470 16740 1490
rect 16760 1470 16770 1490
rect 16730 1460 16770 1470
rect 16922 1470 16928 1490
rect 16945 1470 16954 1490
rect 16922 1460 16954 1470
rect 17030 1470 17040 1490
rect 17060 1470 17070 1490
rect 17030 1460 17070 1470
rect 17146 1470 17152 1490
rect 17169 1470 17178 1490
rect 17146 1460 17178 1470
rect 17345 1470 17355 1490
rect 17375 1470 17385 1490
rect 17345 1460 17385 1470
rect 17565 1470 17575 1490
rect 17595 1470 17605 1490
rect 17565 1460 17605 1470
rect 17770 1470 17780 1490
rect 17800 1470 17810 1490
rect 17770 1460 17810 1470
rect 17595 1245 17635 1255
rect 17595 1240 17605 1245
rect 16815 1230 16845 1240
rect 16815 1210 16820 1230
rect 16840 1210 16845 1230
rect 17510 1225 17605 1240
rect 17625 1225 17635 1245
rect 16245 1185 16260 1200
rect 16300 1195 17360 1210
rect 16300 1185 16315 1195
rect 16355 1185 16370 1195
rect 16410 1185 16425 1195
rect 16465 1185 16480 1195
rect 16520 1185 16535 1195
rect 16575 1185 16590 1195
rect 16630 1185 16645 1195
rect 16685 1185 16700 1195
rect 16740 1185 16755 1195
rect 16795 1185 16810 1195
rect 16850 1185 16865 1195
rect 16905 1185 16920 1195
rect 16960 1185 16975 1195
rect 17015 1185 17030 1195
rect 17070 1185 17085 1195
rect 17125 1185 17140 1195
rect 17180 1185 17195 1195
rect 17235 1185 17250 1195
rect 17290 1185 17305 1195
rect 17345 1185 17360 1195
rect 17400 1195 17470 1210
rect 17400 1185 17415 1195
rect 17455 1185 17470 1195
rect 17510 1185 17525 1225
rect 17595 1215 17635 1225
rect 17565 1185 17580 1200
rect 15195 945 15255 955
rect 15115 930 15255 945
rect 15295 940 15355 955
rect 15395 940 15455 955
rect 15495 940 15555 955
rect 15595 940 15655 955
rect 15695 945 15755 955
rect 15695 930 15835 945
rect 18045 945 18105 955
rect 15115 910 15125 930
rect 15145 910 15155 930
rect 2995 890 3085 905
rect 3035 880 3085 890
rect 3125 890 4885 905
rect 3125 880 3175 890
rect 3215 880 3265 890
rect 3305 880 3355 890
rect 3395 880 3445 890
rect 3485 880 3535 890
rect 3575 880 3625 890
rect 3665 880 3715 890
rect 3755 880 3805 890
rect 3845 880 3895 890
rect 3935 880 3985 890
rect 4025 880 4075 890
rect 4115 880 4165 890
rect 4205 880 4255 890
rect 4295 880 4345 890
rect 4385 880 4435 890
rect 4475 880 4525 890
rect 4565 880 4615 890
rect 4655 880 4705 890
rect 4745 880 4795 890
rect 4835 880 4885 890
rect 4925 890 5015 905
rect 15115 900 15155 910
rect 15795 910 15805 930
rect 15825 910 15835 930
rect 16245 920 16260 935
rect 16300 920 16315 935
rect 16355 920 16370 935
rect 16410 920 16425 935
rect 16465 920 16480 935
rect 16520 920 16535 935
rect 16575 920 16590 935
rect 16630 920 16645 935
rect 16685 920 16700 935
rect 16740 920 16755 935
rect 16795 920 16810 935
rect 16850 920 16865 935
rect 16905 920 16920 935
rect 16960 920 16975 935
rect 17015 920 17030 935
rect 17070 920 17085 935
rect 17125 920 17140 935
rect 17180 920 17195 935
rect 17235 920 17250 935
rect 17290 920 17305 935
rect 17345 920 17360 935
rect 17400 920 17415 935
rect 17455 920 17470 935
rect 17510 920 17525 935
rect 17565 920 17580 935
rect 17965 930 18105 945
rect 18145 940 18205 955
rect 18245 940 18305 955
rect 18345 940 18405 955
rect 18445 940 18505 955
rect 18545 945 18605 955
rect 18545 930 18685 945
rect 15795 900 15835 910
rect 16165 910 16260 920
rect 16165 890 16175 910
rect 16195 905 16260 910
rect 17565 910 17660 920
rect 17565 905 17630 910
rect 16195 890 16205 905
rect 4925 880 4975 890
rect 16165 880 16205 890
rect 17620 890 17630 905
rect 17650 890 17660 910
rect 17965 910 17975 930
rect 17995 910 18005 930
rect 17965 900 18005 910
rect 18645 910 18655 930
rect 18675 910 18685 930
rect 18645 900 18685 910
rect 17620 880 17660 890
rect 16305 790 16345 800
rect 3035 765 3085 780
rect 3125 755 3175 780
rect 3215 765 3265 780
rect 3305 765 3355 780
rect 3395 765 3445 780
rect 3485 765 3535 780
rect 3575 765 3625 780
rect 3665 765 3715 780
rect 3755 765 3805 780
rect 3845 765 3895 780
rect 3935 765 3985 780
rect 4025 765 4075 780
rect 4115 765 4165 780
rect 4205 765 4255 780
rect 4295 765 4345 780
rect 4385 765 4435 780
rect 4475 765 4525 780
rect 4565 765 4615 780
rect 4655 765 4705 780
rect 4745 765 4795 780
rect 4835 765 4885 780
rect 4925 765 4975 780
rect 16305 770 16315 790
rect 16335 770 16345 790
rect 16305 760 16345 770
rect 16375 790 16415 800
rect 16375 770 16385 790
rect 16405 770 16415 790
rect 16375 760 16415 770
rect 16445 790 16485 800
rect 16445 770 16455 790
rect 16475 770 16485 790
rect 16935 795 16975 805
rect 16935 775 16945 795
rect 16965 775 16975 795
rect 17155 795 17195 805
rect 17155 775 17165 795
rect 17185 775 17195 795
rect 17375 795 17415 805
rect 17375 775 17385 795
rect 17405 775 17415 795
rect 16445 760 16485 770
rect 16920 760 17485 775
rect 3125 750 3140 755
rect 3130 735 3140 750
rect 3160 750 3175 755
rect 3160 735 3170 750
rect 16300 745 16490 760
rect 16920 750 16935 760
rect 16975 750 16990 760
rect 17030 750 17045 760
rect 17085 750 17100 760
rect 17140 750 17155 760
rect 17195 750 17210 760
rect 17250 750 17265 760
rect 17305 750 17320 760
rect 17360 750 17375 760
rect 17415 750 17430 760
rect 17470 750 17485 760
rect 17525 750 17540 765
rect 3130 725 3170 735
rect 16920 690 16935 700
rect 16840 675 16935 690
rect 16975 685 16990 700
rect 17030 685 17045 700
rect 17085 685 17100 700
rect 17140 685 17155 700
rect 17195 685 17210 700
rect 17250 685 17265 700
rect 17305 685 17320 700
rect 17360 685 17375 700
rect 17415 685 17430 700
rect 17470 685 17485 700
rect 17525 690 17540 700
rect 17525 675 17620 690
rect 16840 655 16850 675
rect 16870 655 16880 675
rect 16840 645 16880 655
rect 17580 655 17590 675
rect 17610 655 17620 675
rect 17580 645 17620 655
rect 16300 630 16490 645
<< polycont >>
rect 16640 4490 16660 4510
rect 16760 4490 16780 4510
rect 16880 4490 16900 4510
rect 16210 4430 16230 4450
rect 16470 4430 16490 4450
rect 16580 4445 16600 4465
rect 16940 4445 16960 4465
rect 16340 4295 16360 4315
rect 16760 4290 16780 4310
rect 17211 4290 17229 4310
rect 16220 4180 16240 4200
rect 17510 4180 17530 4200
rect 16370 4060 16390 4080
rect 16165 3875 16185 3895
rect 16277 3875 16294 3895
rect 16480 3875 16500 3895
rect 16700 3875 16720 3895
rect 16905 3875 16925 3895
rect 17017 3875 17034 3895
rect 17220 3875 17240 3895
rect 17440 3875 17460 3895
rect 17645 3875 17665 3895
rect 16408 3755 16425 3775
rect 16628 3755 16645 3775
rect 16775 3755 16792 3775
rect 17148 3755 17165 3775
rect 17368 3755 17385 3775
rect 17515 3755 17532 3775
rect 16190 3600 16210 3620
rect 17590 3600 17610 3620
rect 3145 2955 3165 2975
rect 4845 2955 4865 2975
rect 16831 3130 16849 3150
rect 15125 2940 15145 2960
rect 15661 2940 15679 2960
rect 15865 2940 15885 2960
rect 16190 2920 16210 2940
rect 17590 2920 17610 2940
rect 17915 2940 17935 2960
rect 18121 2940 18139 2960
rect 18655 2940 18675 2960
rect 3005 2785 3025 2805
rect 4985 2785 5005 2805
rect 3185 2725 3205 2745
rect 4805 2725 4825 2745
rect 3365 2350 3385 2370
rect 3895 2355 3915 2375
rect 16831 2450 16849 2470
rect 15125 2410 15145 2430
rect 15865 2410 15885 2430
rect 17915 2410 17935 2430
rect 15775 2365 15795 2385
rect 18655 2410 18675 2430
rect 15125 2290 15145 2310
rect 18035 2350 18055 2370
rect 15865 2290 15885 2310
rect 17915 2290 17935 2310
rect 18655 2290 18675 2310
rect 16836 2155 16854 2175
rect 16245 1935 16265 1955
rect 17535 1935 17555 1955
rect 2630 1855 2650 1875
rect 2775 1855 2795 1875
rect 2845 1855 2865 1875
rect 2935 1855 2955 1875
rect 3175 1855 3195 1875
rect 3295 1855 3315 1875
rect 3535 1855 3555 1875
rect 3655 1855 3675 1875
rect 3865 1855 3885 1875
rect 3995 1850 4015 1870
rect 4125 1855 4145 1875
rect 4335 1855 4355 1875
rect 4455 1855 4475 1875
rect 4695 1855 4715 1875
rect 4815 1855 4835 1875
rect 5055 1855 5075 1875
rect 5145 1855 5165 1875
rect 5215 1855 5235 1875
rect 3235 1735 3255 1755
rect 4755 1735 4775 1755
rect 15566 1680 15584 1700
rect 16243 1690 16260 1710
rect 16463 1690 16480 1710
rect 16610 1690 16627 1710
rect 16876 1690 16893 1710
rect 17283 1690 17300 1710
rect 17503 1690 17520 1710
rect 17650 1690 17667 1710
rect 18216 1680 18234 1700
rect 3175 1570 3195 1590
rect 4815 1570 4835 1590
rect 2935 1475 2955 1495
rect 3055 1475 3075 1495
rect 3175 1475 3195 1495
rect 3295 1475 3315 1495
rect 3535 1475 3555 1495
rect 3655 1475 3675 1495
rect 3775 1475 3795 1495
rect 4215 1475 4235 1495
rect 4335 1475 4355 1495
rect 4455 1475 4475 1495
rect 4695 1475 4715 1495
rect 4815 1475 4835 1495
rect 4935 1475 4955 1495
rect 5055 1475 5075 1495
rect 3035 1100 3055 1120
rect 3115 1100 3135 1120
rect 3195 1100 3215 1120
rect 3275 1100 3295 1120
rect 3355 1100 3375 1120
rect 3435 1100 3455 1120
rect 3515 1100 3535 1120
rect 3595 1100 3615 1120
rect 3675 1100 3695 1120
rect 3755 1100 3775 1120
rect 3835 1100 3855 1120
rect 3915 1100 3935 1120
rect 4075 1100 4095 1120
rect 4155 1100 4175 1120
rect 4235 1100 4255 1120
rect 4315 1100 4335 1120
rect 4395 1100 4415 1120
rect 4475 1100 4495 1120
rect 4555 1100 4575 1120
rect 4635 1100 4655 1120
rect 4715 1100 4735 1120
rect 4795 1100 4815 1120
rect 4875 1100 4895 1120
rect 4955 1100 4975 1120
rect 3005 905 3025 925
rect 4985 905 5005 925
rect 16000 1470 16020 1490
rect 16112 1470 16129 1490
rect 16315 1470 16335 1490
rect 16535 1470 16555 1490
rect 16740 1470 16760 1490
rect 16928 1470 16945 1490
rect 17040 1470 17060 1490
rect 17152 1470 17169 1490
rect 17355 1470 17375 1490
rect 17575 1470 17595 1490
rect 17780 1470 17800 1490
rect 16820 1210 16840 1230
rect 17605 1225 17625 1245
rect 15125 910 15145 930
rect 15805 910 15825 930
rect 16175 890 16195 910
rect 17630 890 17650 910
rect 17975 910 17995 930
rect 18655 910 18675 930
rect 16315 770 16335 790
rect 16385 770 16405 790
rect 16455 770 16475 790
rect 16945 775 16965 795
rect 17165 775 17185 795
rect 17385 775 17405 795
rect 3140 735 3160 755
rect 16850 655 16870 675
rect 17590 655 17610 675
<< xpolycontact >>
rect 14904 3300 15045 3520
rect 91 3170 311 3205
rect 925 3170 1145 3205
rect 1306 3165 1526 3200
rect 2110 3165 2330 3200
rect 91 3110 311 3145
rect 925 3110 1145 3145
rect 1306 3105 1526 3140
rect 2110 3105 2330 3140
rect 91 3030 311 3065
rect 895 3030 1115 3065
rect 1306 3045 1526 3080
rect 2110 3045 2330 3080
rect 91 2970 311 3005
rect 895 2970 1115 3005
rect 1306 2985 1526 3020
rect 2110 2985 2330 3020
rect 1306 2925 1526 2960
rect 2110 2925 2330 2960
rect 14904 2940 15045 3160
rect 18755 3300 18896 3520
rect 1306 2865 1526 2900
rect 2110 2865 2330 2900
rect 96 2820 315 2855
rect 504 2820 724 2855
rect 1306 2805 1526 2840
rect 1740 2805 1960 2840
rect 18755 2940 18896 3160
rect 96 2760 315 2795
rect 504 2760 724 2795
rect 14790 2405 14825 2625
rect 14790 2010 14825 2230
rect 14850 2405 14885 2625
rect 14850 2010 14885 2230
rect 14910 2405 14945 2625
rect 14910 2010 14945 2230
rect 14970 2405 15005 2625
rect 18795 2405 18830 2625
rect 14970 2010 15005 2230
rect 18795 2010 18830 2230
rect 18855 2405 18890 2625
rect 18855 2010 18890 2230
rect 18915 2405 18950 2625
rect 18915 2010 18950 2230
rect 18975 2405 19010 2625
rect 18975 2010 19010 2230
rect 14970 1385 15005 1605
rect 14970 910 15005 1130
rect 15030 1385 15065 1605
rect 15030 910 15065 1130
rect 18735 1385 18770 1605
rect 18735 910 18770 1130
rect 18795 1385 18830 1605
rect 18795 910 18830 1130
<< ppolyres >>
rect 14904 3160 15045 3300
rect 18755 3160 18896 3300
rect 315 2820 504 2855
rect 315 2760 504 2795
<< xpolyres >>
rect 311 3170 925 3205
rect 1526 3165 2110 3200
rect 311 3110 925 3145
rect 1526 3105 2110 3140
rect 311 3030 895 3065
rect 1526 3045 2110 3080
rect 311 2970 895 3005
rect 1526 2985 2110 3020
rect 1526 2925 2110 2960
rect 1526 2865 2110 2900
rect 1526 2805 1740 2840
rect 14790 2230 14825 2405
rect 14850 2230 14885 2405
rect 14910 2230 14945 2405
rect 14970 2230 15005 2405
rect 18795 2230 18830 2405
rect 18855 2230 18890 2405
rect 18915 2230 18950 2405
rect 18975 2230 19010 2405
rect 14970 1130 15005 1385
rect 15030 1130 15065 1385
rect 18735 1130 18770 1385
rect 18795 1130 18830 1385
<< locali >>
rect 16632 4510 16668 4520
rect 16632 4490 16640 4510
rect 16660 4490 16668 4510
rect 16632 4480 16668 4490
rect 16752 4510 16788 4520
rect 16752 4490 16760 4510
rect 16780 4490 16788 4510
rect 16752 4480 16788 4490
rect 16872 4510 16908 4520
rect 16872 4490 16880 4510
rect 16900 4490 16908 4510
rect 16872 4480 16908 4490
rect 16570 4465 16610 4475
rect 16200 4450 16240 4460
rect 16200 4430 16210 4450
rect 16230 4430 16240 4450
rect 16200 4420 16240 4430
rect 16460 4450 16500 4460
rect 16460 4430 16470 4450
rect 16490 4430 16500 4450
rect 16570 4445 16580 4465
rect 16600 4445 16610 4465
rect 16570 4435 16610 4445
rect 16460 4420 16500 4430
rect 16210 4398 16230 4420
rect 16470 4398 16490 4420
rect 16580 4415 16600 4435
rect 16640 4415 16660 4480
rect 16690 4465 16730 4475
rect 16690 4445 16700 4465
rect 16720 4445 16730 4465
rect 16690 4435 16730 4445
rect 16700 4415 16720 4435
rect 16760 4415 16780 4480
rect 16810 4465 16850 4475
rect 16810 4445 16820 4465
rect 16840 4445 16850 4465
rect 16810 4435 16850 4445
rect 16820 4415 16840 4435
rect 16880 4415 16900 4480
rect 16930 4465 16970 4475
rect 16930 4445 16940 4465
rect 16960 4445 16970 4465
rect 16930 4435 16970 4445
rect 17080 4440 17120 4450
rect 16940 4415 16960 4435
rect 17080 4420 17090 4440
rect 17110 4420 17120 4440
rect 16205 4375 16275 4398
rect 16205 4355 16210 4375
rect 16230 4355 16250 4375
rect 16270 4355 16275 4375
rect 16205 4345 16275 4355
rect 16305 4380 16335 4398
rect 16305 4360 16310 4380
rect 16330 4360 16335 4380
rect 16305 4345 16335 4360
rect 16365 4380 16395 4398
rect 16365 4360 16370 4380
rect 16390 4360 16395 4380
rect 16365 4345 16395 4360
rect 16425 4375 16495 4398
rect 16425 4355 16430 4375
rect 16450 4355 16470 4375
rect 16490 4355 16495 4375
rect 16425 4345 16495 4355
rect 16535 4390 16605 4415
rect 16535 4370 16540 4390
rect 16560 4370 16580 4390
rect 16600 4370 16605 4390
rect 16535 4345 16605 4370
rect 16635 4390 16665 4415
rect 16635 4370 16640 4390
rect 16660 4370 16665 4390
rect 16635 4345 16665 4370
rect 16695 4390 16725 4415
rect 16695 4370 16700 4390
rect 16720 4370 16725 4390
rect 16695 4345 16725 4370
rect 16755 4390 16785 4415
rect 16755 4370 16760 4390
rect 16780 4370 16785 4390
rect 16755 4345 16785 4370
rect 16815 4390 16845 4415
rect 16815 4370 16820 4390
rect 16840 4370 16845 4390
rect 16815 4345 16845 4370
rect 16875 4390 16905 4415
rect 16875 4370 16880 4390
rect 16900 4370 16905 4390
rect 16875 4345 16905 4370
rect 16935 4390 17005 4415
rect 17080 4410 17120 4420
rect 17200 4440 17240 4450
rect 17200 4420 17210 4440
rect 17230 4420 17240 4440
rect 17200 4410 17240 4420
rect 17320 4440 17360 4450
rect 17320 4420 17330 4440
rect 17350 4420 17360 4440
rect 17320 4410 17360 4420
rect 17440 4440 17480 4450
rect 17440 4420 17450 4440
rect 17470 4420 17480 4440
rect 17440 4410 17480 4420
rect 17560 4440 17600 4450
rect 17560 4420 17570 4440
rect 17590 4420 17600 4440
rect 17560 4410 17600 4420
rect 17090 4390 17110 4410
rect 17210 4390 17230 4410
rect 17330 4390 17350 4410
rect 17450 4390 17470 4410
rect 17570 4390 17590 4410
rect 16935 4370 16940 4390
rect 16960 4370 16980 4390
rect 17000 4370 17005 4390
rect 16935 4345 17005 4370
rect 17045 4375 17115 4390
rect 17045 4355 17050 4375
rect 17070 4355 17090 4375
rect 17110 4355 17115 4375
rect 16370 4325 16390 4345
rect 17045 4340 17115 4355
rect 17145 4375 17175 4390
rect 17145 4355 17150 4375
rect 17170 4355 17175 4375
rect 17145 4340 17175 4355
rect 17205 4375 17235 4390
rect 17205 4355 17210 4375
rect 17230 4355 17235 4375
rect 17205 4340 17235 4355
rect 17265 4375 17295 4390
rect 17265 4355 17270 4375
rect 17290 4355 17295 4375
rect 17265 4340 17295 4355
rect 17325 4375 17355 4390
rect 17325 4355 17330 4375
rect 17350 4355 17355 4375
rect 17325 4340 17355 4355
rect 17385 4375 17415 4390
rect 17385 4355 17390 4375
rect 17410 4355 17415 4375
rect 17385 4340 17415 4355
rect 17445 4375 17475 4390
rect 17445 4355 17450 4375
rect 17470 4355 17475 4375
rect 17445 4340 17475 4355
rect 17505 4375 17535 4390
rect 17505 4355 17510 4375
rect 17530 4355 17535 4375
rect 17505 4340 17535 4355
rect 17565 4375 17635 4390
rect 17565 4355 17570 4375
rect 17590 4355 17610 4375
rect 17630 4355 17635 4375
rect 17565 4340 17635 4355
rect 16330 4320 16390 4325
rect 17150 4320 17170 4340
rect 17270 4320 17290 4340
rect 17390 4320 17410 4340
rect 17510 4320 17530 4340
rect 16330 4295 16340 4320
rect 16360 4305 16390 4320
rect 16750 4310 16790 4320
rect 16360 4295 16370 4305
rect 16330 4285 16370 4295
rect 16750 4290 16760 4310
rect 16780 4290 16790 4310
rect 16750 4280 16790 4290
rect 17140 4310 17180 4320
rect 17140 4290 17150 4310
rect 17170 4290 17180 4310
rect 17140 4280 17180 4290
rect 17203 4310 17237 4320
rect 17203 4290 17211 4310
rect 17229 4290 17237 4310
rect 17203 4280 17237 4290
rect 17260 4310 17300 4320
rect 17260 4290 17270 4310
rect 17290 4290 17300 4310
rect 17260 4280 17300 4290
rect 17380 4310 17420 4320
rect 17380 4290 17390 4310
rect 17410 4290 17420 4310
rect 17380 4280 17420 4290
rect 17500 4310 17540 4320
rect 17500 4290 17510 4310
rect 17530 4290 17540 4310
rect 17500 4280 17540 4290
rect 16210 4200 16250 4210
rect 16210 4180 16220 4200
rect 16240 4180 16250 4200
rect 16210 4170 16250 4180
rect 16360 4200 16400 4210
rect 16360 4180 16370 4200
rect 16390 4180 16400 4200
rect 16360 4170 16400 4180
rect 16470 4200 16510 4210
rect 16470 4180 16480 4200
rect 16500 4180 16510 4200
rect 16470 4170 16510 4180
rect 16580 4200 16620 4210
rect 16580 4180 16590 4200
rect 16610 4180 16620 4200
rect 16580 4170 16620 4180
rect 16690 4200 16730 4210
rect 16690 4180 16700 4200
rect 16720 4180 16730 4200
rect 16690 4170 16730 4180
rect 16800 4200 16840 4210
rect 16800 4180 16810 4200
rect 16830 4180 16840 4200
rect 16800 4170 16840 4180
rect 16910 4200 16950 4210
rect 16910 4180 16920 4200
rect 16940 4180 16950 4200
rect 16910 4170 16950 4180
rect 17020 4200 17060 4210
rect 17020 4180 17030 4200
rect 17050 4180 17060 4200
rect 17020 4170 17060 4180
rect 17130 4200 17170 4210
rect 17130 4180 17140 4200
rect 17160 4180 17170 4200
rect 17130 4170 17170 4180
rect 17240 4200 17280 4210
rect 17240 4180 17250 4200
rect 17270 4180 17280 4200
rect 17240 4170 17280 4180
rect 17350 4200 17390 4210
rect 17350 4180 17360 4200
rect 17380 4180 17390 4200
rect 17350 4170 17390 4180
rect 17500 4200 17540 4210
rect 17500 4180 17510 4200
rect 17530 4180 17540 4200
rect 17500 4170 17540 4180
rect 16220 4150 16240 4170
rect 16370 4150 16390 4170
rect 16480 4150 16500 4170
rect 16590 4150 16610 4170
rect 16700 4150 16720 4170
rect 16810 4150 16830 4170
rect 16920 4150 16940 4170
rect 17030 4150 17050 4170
rect 17140 4150 17160 4170
rect 17250 4150 17270 4170
rect 17360 4150 17380 4170
rect 17510 4150 17530 4170
rect 16215 4140 16285 4150
rect 16215 4120 16220 4140
rect 16240 4120 16260 4140
rect 16280 4120 16285 4140
rect 16215 4110 16285 4120
rect 16310 4140 16340 4150
rect 16310 4120 16315 4140
rect 16335 4120 16340 4140
rect 16310 4110 16340 4120
rect 16365 4140 16395 4150
rect 16365 4120 16370 4140
rect 16390 4120 16395 4140
rect 16365 4110 16395 4120
rect 16420 4140 16450 4150
rect 16420 4120 16425 4140
rect 16445 4120 16450 4140
rect 16420 4110 16450 4120
rect 16475 4140 16505 4150
rect 16475 4120 16480 4140
rect 16500 4120 16505 4140
rect 16475 4110 16505 4120
rect 16530 4140 16560 4150
rect 16530 4120 16535 4140
rect 16555 4120 16560 4140
rect 16530 4110 16560 4120
rect 16585 4140 16615 4150
rect 16585 4120 16590 4140
rect 16610 4120 16615 4140
rect 16585 4110 16615 4120
rect 16640 4140 16670 4150
rect 16640 4120 16645 4140
rect 16665 4120 16670 4140
rect 16640 4110 16670 4120
rect 16695 4140 16725 4150
rect 16695 4120 16700 4140
rect 16720 4120 16725 4140
rect 16695 4110 16725 4120
rect 16750 4140 16780 4150
rect 16750 4120 16755 4140
rect 16775 4120 16780 4140
rect 16750 4110 16780 4120
rect 16805 4140 16835 4150
rect 16805 4120 16810 4140
rect 16830 4120 16835 4140
rect 16805 4110 16835 4120
rect 16860 4140 16890 4150
rect 16860 4120 16865 4140
rect 16885 4120 16890 4140
rect 16860 4110 16890 4120
rect 16915 4140 16945 4150
rect 16915 4120 16920 4140
rect 16940 4120 16945 4140
rect 16915 4110 16945 4120
rect 16970 4140 17000 4150
rect 16970 4120 16975 4140
rect 16995 4120 17000 4140
rect 16970 4110 17000 4120
rect 17025 4140 17055 4150
rect 17025 4120 17030 4140
rect 17050 4120 17055 4140
rect 17025 4110 17055 4120
rect 17080 4140 17110 4150
rect 17080 4120 17085 4140
rect 17105 4120 17110 4140
rect 17080 4110 17110 4120
rect 17135 4140 17165 4150
rect 17135 4120 17140 4140
rect 17160 4120 17165 4140
rect 17135 4110 17165 4120
rect 17190 4140 17220 4150
rect 17190 4120 17195 4140
rect 17215 4120 17220 4140
rect 17190 4110 17220 4120
rect 17245 4140 17275 4150
rect 17245 4120 17250 4140
rect 17270 4120 17275 4140
rect 17245 4110 17275 4120
rect 17300 4140 17330 4150
rect 17300 4120 17305 4140
rect 17325 4120 17330 4140
rect 17300 4110 17330 4120
rect 17355 4140 17385 4150
rect 17355 4120 17360 4140
rect 17380 4120 17385 4140
rect 17355 4110 17385 4120
rect 17410 4140 17440 4150
rect 17410 4120 17415 4140
rect 17435 4120 17440 4140
rect 17410 4110 17440 4120
rect 17465 4140 17535 4150
rect 17465 4120 17470 4140
rect 17490 4120 17510 4140
rect 17530 4120 17535 4140
rect 17465 4110 17535 4120
rect 16315 4090 16335 4110
rect 16425 4090 16445 4110
rect 16535 4090 16555 4110
rect 16645 4090 16665 4110
rect 16755 4090 16775 4110
rect 16865 4090 16885 4110
rect 16975 4090 16995 4110
rect 17085 4090 17105 4110
rect 17195 4090 17215 4110
rect 17305 4090 17325 4110
rect 17415 4090 17435 4110
rect 16305 4080 16345 4090
rect 16305 4060 16315 4080
rect 16335 4060 16345 4080
rect 16305 4050 16345 4060
rect 16362 4080 16398 4090
rect 16362 4060 16370 4080
rect 16390 4060 16398 4080
rect 16362 4050 16398 4060
rect 16415 4080 16455 4090
rect 16415 4060 16425 4080
rect 16445 4060 16455 4080
rect 16415 4050 16455 4060
rect 16525 4080 16565 4090
rect 16525 4060 16535 4080
rect 16555 4060 16565 4080
rect 16525 4050 16565 4060
rect 16635 4080 16675 4090
rect 16635 4060 16645 4080
rect 16665 4060 16675 4080
rect 16635 4050 16675 4060
rect 16745 4080 16785 4090
rect 16745 4060 16755 4080
rect 16775 4060 16785 4080
rect 16745 4050 16785 4060
rect 16855 4080 16895 4090
rect 16855 4060 16865 4080
rect 16885 4060 16895 4080
rect 16855 4050 16895 4060
rect 16965 4080 17005 4090
rect 16965 4060 16975 4080
rect 16995 4060 17005 4080
rect 16965 4050 17005 4060
rect 17075 4080 17115 4090
rect 17075 4060 17085 4080
rect 17105 4060 17115 4080
rect 17075 4050 17115 4060
rect 17185 4080 17225 4090
rect 17185 4060 17195 4080
rect 17215 4060 17225 4080
rect 17185 4050 17225 4060
rect 17295 4080 17335 4090
rect 17295 4060 17305 4080
rect 17325 4060 17335 4080
rect 17295 4050 17335 4060
rect 17405 4080 17445 4090
rect 17405 4060 17415 4080
rect 17435 4060 17445 4080
rect 17405 4050 17445 4060
rect 16415 3990 16455 4030
rect 16635 3990 16675 4030
rect 16855 3990 16895 4030
rect 17075 3990 17115 4030
rect 17295 3990 17335 4030
rect 16310 3955 16350 3965
rect 16310 3935 16320 3955
rect 16340 3935 16350 3955
rect 16310 3925 16350 3935
rect 16415 3955 16455 3965
rect 16415 3935 16425 3955
rect 16445 3935 16455 3955
rect 16415 3925 16455 3935
rect 16525 3955 16565 3965
rect 16525 3935 16535 3955
rect 16555 3935 16565 3955
rect 16525 3925 16565 3935
rect 16635 3955 16675 3965
rect 16635 3935 16645 3955
rect 16665 3935 16675 3955
rect 16635 3925 16675 3935
rect 16745 3955 16785 3965
rect 16745 3935 16755 3955
rect 16775 3935 16785 3955
rect 16745 3925 16785 3935
rect 17050 3955 17090 3965
rect 17050 3935 17060 3955
rect 17080 3935 17090 3955
rect 17050 3925 17090 3935
rect 17155 3955 17195 3965
rect 17155 3935 17165 3955
rect 17185 3935 17195 3955
rect 17155 3925 17195 3935
rect 17265 3955 17305 3965
rect 17265 3935 17275 3955
rect 17295 3935 17305 3955
rect 17265 3925 17305 3935
rect 17375 3955 17415 3965
rect 17375 3935 17385 3955
rect 17405 3935 17415 3955
rect 17375 3925 17415 3935
rect 17485 3955 17525 3965
rect 17485 3935 17495 3955
rect 17515 3935 17525 3955
rect 17485 3925 17525 3935
rect 16155 3895 16195 3905
rect 16155 3875 16165 3895
rect 16185 3875 16195 3895
rect 16155 3865 16195 3875
rect 16271 3895 16303 3905
rect 16271 3875 16277 3895
rect 16294 3875 16303 3895
rect 16271 3865 16303 3875
rect 16165 3845 16185 3865
rect 16320 3845 16340 3925
rect 16360 3895 16400 3905
rect 16360 3875 16370 3895
rect 16390 3875 16400 3895
rect 16360 3865 16400 3875
rect 16370 3845 16390 3865
rect 16425 3845 16445 3925
rect 16470 3895 16510 3905
rect 16470 3875 16480 3895
rect 16500 3875 16510 3895
rect 16470 3865 16510 3875
rect 16535 3845 16555 3925
rect 16645 3845 16665 3925
rect 16690 3895 16730 3905
rect 16690 3875 16700 3895
rect 16720 3875 16730 3895
rect 16690 3865 16730 3875
rect 16755 3845 16775 3925
rect 16800 3895 16840 3905
rect 16800 3875 16810 3895
rect 16830 3875 16840 3895
rect 16800 3865 16840 3875
rect 16895 3895 16935 3905
rect 16895 3875 16905 3895
rect 16925 3875 16935 3895
rect 16895 3865 16935 3875
rect 17011 3895 17043 3905
rect 17011 3875 17017 3895
rect 17034 3875 17043 3895
rect 17011 3865 17043 3875
rect 16810 3845 16830 3865
rect 16905 3845 16925 3865
rect 17060 3845 17080 3925
rect 17165 3845 17185 3925
rect 17210 3895 17250 3905
rect 17210 3875 17220 3895
rect 17240 3875 17250 3895
rect 17210 3865 17250 3875
rect 17275 3845 17295 3925
rect 17385 3845 17405 3925
rect 17430 3895 17470 3905
rect 17430 3875 17440 3895
rect 17460 3875 17470 3895
rect 17430 3865 17470 3875
rect 17495 3845 17515 3925
rect 17635 3895 17675 3905
rect 17635 3875 17645 3895
rect 17665 3875 17675 3895
rect 17635 3865 17675 3875
rect 17765 3870 17795 3900
rect 17645 3845 17665 3865
rect 16155 3835 16230 3845
rect 16155 3815 16165 3835
rect 16185 3815 16205 3835
rect 16225 3815 16230 3835
rect 16155 3805 16230 3815
rect 16255 3835 16285 3845
rect 16255 3815 16260 3835
rect 16280 3815 16285 3835
rect 16255 3805 16285 3815
rect 16310 3835 16340 3845
rect 16310 3815 16315 3835
rect 16335 3815 16340 3835
rect 16310 3805 16340 3815
rect 16365 3835 16395 3845
rect 16365 3815 16370 3835
rect 16390 3815 16395 3835
rect 16365 3805 16395 3815
rect 16420 3835 16450 3845
rect 16420 3815 16425 3835
rect 16445 3815 16450 3835
rect 16420 3805 16450 3815
rect 16475 3835 16505 3845
rect 16475 3815 16480 3835
rect 16500 3815 16505 3835
rect 16475 3805 16505 3815
rect 16530 3835 16560 3845
rect 16530 3815 16535 3835
rect 16555 3815 16560 3835
rect 16530 3805 16560 3815
rect 16585 3835 16615 3845
rect 16585 3815 16590 3835
rect 16610 3815 16615 3835
rect 16585 3805 16615 3815
rect 16640 3835 16670 3845
rect 16640 3815 16645 3835
rect 16665 3815 16670 3835
rect 16640 3805 16670 3815
rect 16695 3835 16725 3845
rect 16695 3815 16700 3835
rect 16720 3815 16725 3835
rect 16695 3805 16725 3815
rect 16750 3835 16780 3845
rect 16750 3815 16755 3835
rect 16775 3815 16780 3835
rect 16750 3805 16780 3815
rect 16805 3835 16835 3845
rect 16805 3815 16810 3835
rect 16830 3815 16835 3835
rect 16805 3805 16835 3815
rect 16860 3835 16970 3845
rect 16860 3815 16865 3835
rect 16885 3815 16905 3835
rect 16925 3815 16945 3835
rect 16965 3815 16970 3835
rect 16860 3805 16970 3815
rect 16995 3835 17025 3845
rect 16995 3815 17000 3835
rect 17020 3815 17025 3835
rect 16995 3805 17025 3815
rect 17050 3835 17080 3845
rect 17050 3815 17055 3835
rect 17075 3815 17080 3835
rect 17050 3805 17080 3815
rect 17105 3835 17135 3845
rect 17105 3815 17110 3835
rect 17130 3815 17135 3835
rect 17105 3805 17135 3815
rect 17160 3835 17190 3845
rect 17160 3815 17165 3835
rect 17185 3815 17190 3835
rect 17160 3805 17190 3815
rect 17215 3835 17245 3845
rect 17215 3815 17220 3835
rect 17240 3815 17245 3835
rect 17215 3805 17245 3815
rect 17270 3835 17300 3845
rect 17270 3815 17275 3835
rect 17295 3815 17300 3835
rect 17270 3805 17300 3815
rect 17325 3835 17355 3845
rect 17325 3815 17330 3835
rect 17350 3815 17355 3835
rect 17325 3805 17355 3815
rect 17380 3835 17410 3845
rect 17380 3815 17385 3835
rect 17405 3815 17410 3835
rect 17380 3805 17410 3815
rect 17435 3835 17465 3845
rect 17435 3815 17440 3835
rect 17460 3815 17465 3835
rect 17435 3805 17465 3815
rect 17490 3835 17520 3845
rect 17490 3815 17495 3835
rect 17515 3815 17520 3835
rect 17490 3805 17520 3815
rect 17545 3835 17575 3845
rect 17545 3815 17550 3835
rect 17570 3815 17575 3835
rect 17545 3805 17575 3815
rect 17600 3835 17675 3845
rect 17600 3815 17605 3835
rect 17625 3815 17645 3835
rect 17665 3815 17675 3835
rect 17600 3805 17675 3815
rect 16260 3725 16280 3805
rect 16365 3725 16385 3805
rect 16402 3775 16434 3785
rect 16402 3755 16408 3775
rect 16425 3755 16434 3775
rect 16402 3745 16434 3755
rect 16480 3725 16500 3805
rect 16585 3725 16605 3805
rect 16622 3775 16654 3785
rect 16622 3755 16628 3775
rect 16645 3755 16654 3775
rect 16622 3745 16654 3755
rect 16700 3725 16720 3805
rect 16766 3775 16798 3785
rect 16766 3755 16775 3775
rect 16792 3755 16798 3775
rect 16766 3745 16798 3755
rect 16815 3725 16835 3805
rect 17000 3735 17020 3805
rect 16990 3725 17030 3735
rect 16250 3715 16290 3725
rect 16250 3695 16260 3715
rect 16280 3695 16290 3715
rect 16250 3685 16290 3695
rect 16355 3715 16395 3725
rect 16355 3695 16365 3715
rect 16385 3695 16395 3715
rect 16355 3685 16395 3695
rect 16470 3715 16510 3725
rect 16470 3695 16480 3715
rect 16500 3695 16510 3715
rect 16470 3685 16510 3695
rect 16575 3715 16615 3725
rect 16575 3695 16585 3715
rect 16605 3695 16615 3715
rect 16575 3685 16615 3695
rect 16690 3715 16730 3725
rect 16690 3695 16700 3715
rect 16720 3695 16730 3715
rect 16690 3685 16730 3695
rect 16805 3715 16845 3725
rect 16805 3695 16815 3715
rect 16835 3695 16845 3715
rect 16990 3705 17000 3725
rect 17020 3705 17030 3725
rect 16990 3695 17030 3705
rect 16805 3685 16845 3695
rect 17105 3690 17125 3805
rect 17142 3775 17174 3785
rect 17142 3755 17148 3775
rect 17165 3755 17174 3775
rect 17142 3745 17174 3755
rect 17220 3735 17240 3805
rect 17210 3725 17250 3735
rect 17210 3705 17220 3725
rect 17240 3705 17250 3725
rect 17210 3695 17250 3705
rect 17325 3690 17345 3805
rect 17362 3775 17394 3785
rect 17362 3755 17368 3775
rect 17385 3755 17394 3775
rect 17362 3745 17394 3755
rect 17440 3735 17460 3805
rect 17506 3775 17538 3785
rect 17506 3755 17515 3775
rect 17532 3755 17538 3775
rect 17506 3745 17538 3755
rect 17430 3725 17470 3735
rect 17430 3705 17440 3725
rect 17460 3705 17470 3725
rect 17430 3695 17470 3705
rect 17555 3690 17575 3805
rect 17865 3700 17895 3730
rect 17095 3650 17135 3690
rect 17315 3650 17355 3690
rect 17545 3650 17585 3690
rect 17810 3655 17840 3685
rect 14960 3605 14990 3635
rect 15210 3630 15250 3640
rect 15210 3610 15220 3630
rect 15240 3610 15250 3630
rect 15210 3600 15250 3610
rect 15320 3630 15360 3640
rect 15320 3610 15330 3630
rect 15350 3610 15360 3630
rect 15320 3600 15360 3610
rect 15430 3630 15470 3640
rect 15430 3610 15440 3630
rect 15460 3610 15470 3630
rect 15430 3600 15470 3610
rect 15540 3630 15580 3640
rect 15540 3610 15550 3630
rect 15570 3610 15580 3630
rect 15540 3600 15580 3610
rect 15650 3630 15690 3640
rect 15650 3610 15660 3630
rect 15680 3610 15690 3630
rect 15650 3600 15690 3610
rect 15760 3630 15800 3640
rect 18000 3630 18040 3640
rect 15760 3610 15770 3630
rect 15790 3610 15800 3630
rect 15760 3600 15800 3610
rect 16180 3620 16220 3630
rect 16180 3600 16190 3620
rect 16210 3600 16220 3620
rect 15220 3580 15240 3600
rect 15330 3580 15350 3600
rect 15440 3580 15460 3600
rect 15550 3580 15570 3600
rect 15660 3580 15680 3600
rect 15770 3580 15790 3600
rect 16180 3590 16220 3600
rect 16340 3620 16380 3630
rect 16340 3600 16350 3620
rect 16370 3600 16380 3620
rect 16340 3590 16380 3600
rect 16460 3620 16500 3630
rect 16460 3600 16470 3620
rect 16490 3600 16500 3620
rect 16460 3590 16500 3600
rect 16580 3620 16620 3630
rect 16580 3600 16590 3620
rect 16610 3600 16620 3620
rect 16580 3590 16620 3600
rect 16700 3620 16740 3630
rect 16700 3600 16710 3620
rect 16730 3600 16740 3620
rect 16700 3590 16740 3600
rect 16820 3620 16860 3630
rect 16820 3600 16830 3620
rect 16850 3600 16860 3620
rect 16820 3590 16860 3600
rect 16940 3620 16980 3630
rect 16940 3600 16950 3620
rect 16970 3600 16980 3620
rect 16940 3590 16980 3600
rect 17060 3620 17100 3630
rect 17060 3600 17070 3620
rect 17090 3600 17100 3620
rect 17060 3590 17100 3600
rect 17180 3620 17220 3630
rect 17180 3600 17190 3620
rect 17210 3600 17220 3620
rect 17180 3590 17220 3600
rect 17300 3620 17340 3630
rect 17300 3600 17310 3620
rect 17330 3600 17340 3620
rect 17300 3590 17340 3600
rect 17420 3620 17460 3630
rect 17420 3600 17430 3620
rect 17450 3600 17460 3620
rect 17420 3590 17460 3600
rect 17580 3620 17620 3630
rect 17580 3600 17590 3620
rect 17610 3600 17620 3620
rect 18000 3610 18010 3630
rect 18030 3610 18040 3630
rect 18000 3600 18040 3610
rect 18110 3630 18150 3640
rect 18110 3610 18120 3630
rect 18140 3610 18150 3630
rect 18110 3600 18150 3610
rect 18220 3630 18260 3640
rect 18220 3610 18230 3630
rect 18250 3610 18260 3630
rect 18220 3600 18260 3610
rect 18330 3630 18370 3640
rect 18330 3610 18340 3630
rect 18360 3610 18370 3630
rect 18330 3600 18370 3610
rect 18440 3630 18480 3640
rect 18440 3610 18450 3630
rect 18470 3610 18480 3630
rect 18440 3600 18480 3610
rect 18550 3630 18590 3640
rect 18550 3610 18560 3630
rect 18580 3610 18590 3630
rect 18550 3600 18590 3610
rect 18810 3605 18840 3635
rect 17580 3590 17620 3600
rect 15120 3570 15190 3580
rect 1266 3495 1296 3525
rect 14904 3520 15045 3560
rect 4445 3465 4475 3495
rect -10 3415 20 3445
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 5145 3415 5175 3445
rect -55 3360 -25 3390
rect 2695 3360 2725 3390
rect 1210 3310 1240 3340
rect 3140 3310 3170 3340
rect 3395 3305 3425 3335
rect 5365 3305 5395 3335
rect 15120 3550 15125 3570
rect 15145 3550 15165 3570
rect 15185 3550 15190 3570
rect 15120 3520 15190 3550
rect 15120 3500 15125 3520
rect 15145 3500 15165 3520
rect 15185 3500 15190 3520
rect 15120 3470 15190 3500
rect 15120 3450 15125 3470
rect 15145 3450 15165 3470
rect 15185 3450 15190 3470
rect 15120 3420 15190 3450
rect 15120 3400 15125 3420
rect 15145 3400 15165 3420
rect 15185 3400 15190 3420
rect 15120 3370 15190 3400
rect 15120 3350 15125 3370
rect 15145 3350 15165 3370
rect 15185 3350 15190 3370
rect 15120 3320 15190 3350
rect 15120 3300 15125 3320
rect 15145 3300 15165 3320
rect 15185 3300 15190 3320
rect 1165 3255 1195 3285
rect 4890 3255 4920 3285
rect 5415 3255 5445 3285
rect 15120 3270 15190 3300
rect 15120 3250 15125 3270
rect 15145 3250 15165 3270
rect 15185 3250 15190 3270
rect 2740 3210 2770 3240
rect 15120 3220 15190 3250
rect 46 3200 91 3205
rect 46 3175 56 3200
rect 81 3175 91 3200
rect 46 3170 91 3175
rect 15120 3200 15125 3220
rect 15145 3200 15165 3220
rect 15185 3200 15190 3220
rect 1110 3145 1145 3170
rect 1261 3195 1306 3200
rect 1261 3170 1271 3195
rect 1296 3170 1306 3195
rect 1261 3165 1306 3170
rect 2330 3165 2370 3200
rect 46 3140 91 3145
rect 46 3115 56 3140
rect 81 3115 91 3140
rect 46 3110 91 3115
rect 1261 3135 1306 3140
rect 1261 3110 1271 3135
rect 1296 3110 1306 3135
rect 1261 3105 1306 3110
rect 1165 3070 1195 3100
rect 2295 3080 2330 3105
rect 46 3060 91 3065
rect 46 3035 56 3060
rect 81 3035 91 3060
rect 46 3030 91 3035
rect 1080 3005 1115 3030
rect 46 3000 91 3005
rect 46 2975 56 3000
rect 81 2975 91 3000
rect 46 2970 91 2975
rect 1266 3045 1306 3080
rect 910 2910 1120 2915
rect 910 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1120 2910
rect 910 2875 1120 2880
rect 1266 2900 1286 3045
rect 2350 3020 2370 3165
rect 2625 3155 2655 3185
rect 4445 3155 4475 3185
rect 15120 3170 15190 3200
rect 3140 3110 3170 3140
rect 4840 3110 4870 3140
rect 5320 3110 5350 3140
rect 3990 3050 4020 3080
rect 2330 2985 2370 3020
rect 3450 3005 3480 3035
rect 3810 3005 3840 3035
rect 4350 3005 4380 3035
rect 4710 3005 4740 3035
rect 1306 2960 1341 2985
rect 2330 2955 2375 2960
rect 2330 2930 2340 2955
rect 2365 2930 2375 2955
rect 2330 2925 2375 2930
rect 2430 2925 2460 2955
rect 2520 2945 2560 2985
rect 3080 2975 3120 2985
rect 3080 2955 3090 2975
rect 3110 2955 3120 2975
rect 3080 2945 3120 2955
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 3265 2975 3305 2985
rect 3265 2955 3275 2975
rect 3295 2955 3305 2975
rect 3265 2945 3305 2955
rect 3445 2975 3485 2985
rect 3445 2955 3455 2975
rect 3475 2955 3485 2975
rect 3445 2945 3485 2955
rect 3625 2975 3665 2985
rect 3625 2955 3635 2975
rect 3655 2955 3665 2975
rect 3625 2945 3665 2955
rect 3805 2975 3845 2985
rect 3805 2955 3815 2975
rect 3835 2955 3845 2975
rect 3805 2945 3845 2955
rect 3985 2975 4025 2985
rect 3985 2955 3995 2975
rect 4015 2955 4025 2975
rect 3985 2945 4025 2955
rect 4165 2975 4205 2985
rect 4165 2955 4175 2975
rect 4195 2955 4205 2975
rect 4165 2945 4205 2955
rect 4345 2975 4385 2985
rect 4345 2955 4355 2975
rect 4375 2955 4385 2975
rect 4345 2945 4385 2955
rect 4525 2975 4565 2985
rect 4525 2955 4535 2975
rect 4555 2955 4565 2975
rect 4525 2945 4565 2955
rect 4705 2975 4745 2985
rect 4705 2955 4715 2975
rect 4735 2955 4745 2975
rect 4705 2945 4745 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 4890 2975 4925 2985
rect 4890 2955 4895 2975
rect 4915 2955 4925 2975
rect 4890 2945 4925 2955
rect 3095 2925 3115 2945
rect 3275 2925 3295 2945
rect 3455 2925 3475 2945
rect 3635 2925 3655 2945
rect 3815 2925 3835 2945
rect 3995 2925 4015 2945
rect 4175 2925 4195 2945
rect 4355 2925 4375 2945
rect 4535 2925 4555 2945
rect 4715 2925 4735 2945
rect 4895 2925 4915 2945
rect 15120 3150 15125 3170
rect 15145 3150 15165 3170
rect 15185 3150 15190 3170
rect 15120 3120 15190 3150
rect 15120 3100 15125 3120
rect 15145 3100 15165 3120
rect 15185 3100 15190 3120
rect 15120 3070 15190 3100
rect 15120 3050 15125 3070
rect 15145 3050 15165 3070
rect 15185 3050 15190 3070
rect 15120 3020 15190 3050
rect 15120 3000 15125 3020
rect 15145 3000 15165 3020
rect 15185 3000 15190 3020
rect 15120 2990 15190 3000
rect 15215 3570 15245 3580
rect 15215 3550 15220 3570
rect 15240 3550 15245 3570
rect 15215 3520 15245 3550
rect 15215 3500 15220 3520
rect 15240 3500 15245 3520
rect 15215 3470 15245 3500
rect 15215 3450 15220 3470
rect 15240 3450 15245 3470
rect 15215 3420 15245 3450
rect 15215 3400 15220 3420
rect 15240 3400 15245 3420
rect 15215 3370 15245 3400
rect 15215 3350 15220 3370
rect 15240 3350 15245 3370
rect 15215 3320 15245 3350
rect 15215 3300 15220 3320
rect 15240 3300 15245 3320
rect 15215 3270 15245 3300
rect 15215 3250 15220 3270
rect 15240 3250 15245 3270
rect 15215 3220 15245 3250
rect 15215 3200 15220 3220
rect 15240 3200 15245 3220
rect 15215 3170 15245 3200
rect 15215 3150 15220 3170
rect 15240 3150 15245 3170
rect 15215 3120 15245 3150
rect 15215 3100 15220 3120
rect 15240 3100 15245 3120
rect 15215 3070 15245 3100
rect 15215 3050 15220 3070
rect 15240 3050 15245 3070
rect 15215 3020 15245 3050
rect 15215 3000 15220 3020
rect 15240 3000 15245 3020
rect 15215 2990 15245 3000
rect 15270 3570 15300 3580
rect 15270 3550 15275 3570
rect 15295 3550 15300 3570
rect 15270 3520 15300 3550
rect 15270 3500 15275 3520
rect 15295 3500 15300 3520
rect 15270 3470 15300 3500
rect 15270 3450 15275 3470
rect 15295 3450 15300 3470
rect 15270 3420 15300 3450
rect 15270 3400 15275 3420
rect 15295 3400 15300 3420
rect 15270 3370 15300 3400
rect 15270 3350 15275 3370
rect 15295 3350 15300 3370
rect 15270 3320 15300 3350
rect 15270 3300 15275 3320
rect 15295 3300 15300 3320
rect 15270 3270 15300 3300
rect 15270 3250 15275 3270
rect 15295 3250 15300 3270
rect 15270 3220 15300 3250
rect 15270 3200 15275 3220
rect 15295 3200 15300 3220
rect 15270 3170 15300 3200
rect 15270 3150 15275 3170
rect 15295 3150 15300 3170
rect 15270 3120 15300 3150
rect 15270 3100 15275 3120
rect 15295 3100 15300 3120
rect 15270 3070 15300 3100
rect 15270 3050 15275 3070
rect 15295 3050 15300 3070
rect 15270 3020 15300 3050
rect 15270 3000 15275 3020
rect 15295 3000 15300 3020
rect 15270 2990 15300 3000
rect 15325 3570 15355 3580
rect 15325 3550 15330 3570
rect 15350 3550 15355 3570
rect 15325 3520 15355 3550
rect 15325 3500 15330 3520
rect 15350 3500 15355 3520
rect 15325 3470 15355 3500
rect 15325 3450 15330 3470
rect 15350 3450 15355 3470
rect 15325 3420 15355 3450
rect 15325 3400 15330 3420
rect 15350 3400 15355 3420
rect 15325 3370 15355 3400
rect 15325 3350 15330 3370
rect 15350 3350 15355 3370
rect 15325 3320 15355 3350
rect 15325 3300 15330 3320
rect 15350 3300 15355 3320
rect 15325 3270 15355 3300
rect 15325 3250 15330 3270
rect 15350 3250 15355 3270
rect 15325 3220 15355 3250
rect 15325 3200 15330 3220
rect 15350 3200 15355 3220
rect 15325 3170 15355 3200
rect 15325 3150 15330 3170
rect 15350 3150 15355 3170
rect 15325 3120 15355 3150
rect 15325 3100 15330 3120
rect 15350 3100 15355 3120
rect 15325 3070 15355 3100
rect 15325 3050 15330 3070
rect 15350 3050 15355 3070
rect 15325 3020 15355 3050
rect 15325 3000 15330 3020
rect 15350 3000 15355 3020
rect 15325 2990 15355 3000
rect 15380 3570 15410 3580
rect 15380 3550 15385 3570
rect 15405 3550 15410 3570
rect 15380 3520 15410 3550
rect 15380 3500 15385 3520
rect 15405 3500 15410 3520
rect 15380 3470 15410 3500
rect 15380 3450 15385 3470
rect 15405 3450 15410 3470
rect 15380 3420 15410 3450
rect 15380 3400 15385 3420
rect 15405 3400 15410 3420
rect 15380 3370 15410 3400
rect 15380 3350 15385 3370
rect 15405 3350 15410 3370
rect 15380 3320 15410 3350
rect 15380 3300 15385 3320
rect 15405 3300 15410 3320
rect 15380 3270 15410 3300
rect 15380 3250 15385 3270
rect 15405 3250 15410 3270
rect 15380 3220 15410 3250
rect 15380 3200 15385 3220
rect 15405 3200 15410 3220
rect 15380 3170 15410 3200
rect 15380 3150 15385 3170
rect 15405 3150 15410 3170
rect 15380 3120 15410 3150
rect 15380 3100 15385 3120
rect 15405 3100 15410 3120
rect 15380 3070 15410 3100
rect 15380 3050 15385 3070
rect 15405 3050 15410 3070
rect 15380 3020 15410 3050
rect 15380 3000 15385 3020
rect 15405 3000 15410 3020
rect 15380 2990 15410 3000
rect 15435 3570 15465 3580
rect 15435 3550 15440 3570
rect 15460 3550 15465 3570
rect 15435 3520 15465 3550
rect 15435 3500 15440 3520
rect 15460 3500 15465 3520
rect 15435 3470 15465 3500
rect 15435 3450 15440 3470
rect 15460 3450 15465 3470
rect 15435 3420 15465 3450
rect 15435 3400 15440 3420
rect 15460 3400 15465 3420
rect 15435 3370 15465 3400
rect 15435 3350 15440 3370
rect 15460 3350 15465 3370
rect 15435 3320 15465 3350
rect 15435 3300 15440 3320
rect 15460 3300 15465 3320
rect 15435 3270 15465 3300
rect 15435 3250 15440 3270
rect 15460 3250 15465 3270
rect 15435 3220 15465 3250
rect 15435 3200 15440 3220
rect 15460 3200 15465 3220
rect 15435 3170 15465 3200
rect 15435 3150 15440 3170
rect 15460 3150 15465 3170
rect 15435 3120 15465 3150
rect 15435 3100 15440 3120
rect 15460 3100 15465 3120
rect 15435 3070 15465 3100
rect 15435 3050 15440 3070
rect 15460 3050 15465 3070
rect 15435 3020 15465 3050
rect 15435 3000 15440 3020
rect 15460 3000 15465 3020
rect 15435 2990 15465 3000
rect 15490 3570 15520 3580
rect 15490 3550 15495 3570
rect 15515 3550 15520 3570
rect 15490 3520 15520 3550
rect 15490 3500 15495 3520
rect 15515 3500 15520 3520
rect 15490 3470 15520 3500
rect 15490 3450 15495 3470
rect 15515 3450 15520 3470
rect 15490 3420 15520 3450
rect 15490 3400 15495 3420
rect 15515 3400 15520 3420
rect 15490 3370 15520 3400
rect 15490 3350 15495 3370
rect 15515 3350 15520 3370
rect 15490 3320 15520 3350
rect 15490 3300 15495 3320
rect 15515 3300 15520 3320
rect 15490 3270 15520 3300
rect 15490 3250 15495 3270
rect 15515 3250 15520 3270
rect 15490 3220 15520 3250
rect 15490 3200 15495 3220
rect 15515 3200 15520 3220
rect 15490 3170 15520 3200
rect 15490 3150 15495 3170
rect 15515 3150 15520 3170
rect 15490 3120 15520 3150
rect 15490 3100 15495 3120
rect 15515 3100 15520 3120
rect 15490 3070 15520 3100
rect 15490 3050 15495 3070
rect 15515 3050 15520 3070
rect 15490 3020 15520 3050
rect 15490 3000 15495 3020
rect 15515 3000 15520 3020
rect 15490 2990 15520 3000
rect 15545 3570 15575 3580
rect 15545 3550 15550 3570
rect 15570 3550 15575 3570
rect 15545 3520 15575 3550
rect 15545 3500 15550 3520
rect 15570 3500 15575 3520
rect 15545 3470 15575 3500
rect 15545 3450 15550 3470
rect 15570 3450 15575 3470
rect 15545 3420 15575 3450
rect 15545 3400 15550 3420
rect 15570 3400 15575 3420
rect 15545 3370 15575 3400
rect 15545 3350 15550 3370
rect 15570 3350 15575 3370
rect 15545 3320 15575 3350
rect 15545 3300 15550 3320
rect 15570 3300 15575 3320
rect 15545 3270 15575 3300
rect 15545 3250 15550 3270
rect 15570 3250 15575 3270
rect 15545 3220 15575 3250
rect 15545 3200 15550 3220
rect 15570 3200 15575 3220
rect 15545 3170 15575 3200
rect 15545 3150 15550 3170
rect 15570 3150 15575 3170
rect 15545 3120 15575 3150
rect 15545 3100 15550 3120
rect 15570 3100 15575 3120
rect 15545 3070 15575 3100
rect 15545 3050 15550 3070
rect 15570 3050 15575 3070
rect 15545 3020 15575 3050
rect 15545 3000 15550 3020
rect 15570 3000 15575 3020
rect 15545 2990 15575 3000
rect 15600 3570 15630 3580
rect 15600 3550 15605 3570
rect 15625 3550 15630 3570
rect 15600 3520 15630 3550
rect 15600 3500 15605 3520
rect 15625 3500 15630 3520
rect 15600 3470 15630 3500
rect 15600 3450 15605 3470
rect 15625 3450 15630 3470
rect 15600 3420 15630 3450
rect 15600 3400 15605 3420
rect 15625 3400 15630 3420
rect 15600 3370 15630 3400
rect 15600 3350 15605 3370
rect 15625 3350 15630 3370
rect 15600 3320 15630 3350
rect 15600 3300 15605 3320
rect 15625 3300 15630 3320
rect 15600 3270 15630 3300
rect 15600 3250 15605 3270
rect 15625 3250 15630 3270
rect 15600 3220 15630 3250
rect 15600 3200 15605 3220
rect 15625 3200 15630 3220
rect 15600 3170 15630 3200
rect 15600 3150 15605 3170
rect 15625 3150 15630 3170
rect 15600 3120 15630 3150
rect 15600 3100 15605 3120
rect 15625 3100 15630 3120
rect 15600 3070 15630 3100
rect 15600 3050 15605 3070
rect 15625 3050 15630 3070
rect 15600 3020 15630 3050
rect 15600 3000 15605 3020
rect 15625 3000 15630 3020
rect 15600 2990 15630 3000
rect 15655 3570 15685 3580
rect 15655 3550 15660 3570
rect 15680 3550 15685 3570
rect 15655 3520 15685 3550
rect 15655 3500 15660 3520
rect 15680 3500 15685 3520
rect 15655 3470 15685 3500
rect 15655 3450 15660 3470
rect 15680 3450 15685 3470
rect 15655 3420 15685 3450
rect 15655 3400 15660 3420
rect 15680 3400 15685 3420
rect 15655 3370 15685 3400
rect 15655 3350 15660 3370
rect 15680 3350 15685 3370
rect 15655 3320 15685 3350
rect 15655 3300 15660 3320
rect 15680 3300 15685 3320
rect 15655 3270 15685 3300
rect 15655 3250 15660 3270
rect 15680 3250 15685 3270
rect 15655 3220 15685 3250
rect 15655 3200 15660 3220
rect 15680 3200 15685 3220
rect 15655 3170 15685 3200
rect 15655 3150 15660 3170
rect 15680 3150 15685 3170
rect 15655 3120 15685 3150
rect 15655 3100 15660 3120
rect 15680 3100 15685 3120
rect 15655 3070 15685 3100
rect 15655 3050 15660 3070
rect 15680 3050 15685 3070
rect 15655 3020 15685 3050
rect 15655 3000 15660 3020
rect 15680 3000 15685 3020
rect 15655 2990 15685 3000
rect 15710 3570 15740 3580
rect 15710 3550 15715 3570
rect 15735 3550 15740 3570
rect 15710 3520 15740 3550
rect 15710 3500 15715 3520
rect 15735 3500 15740 3520
rect 15710 3470 15740 3500
rect 15710 3450 15715 3470
rect 15735 3450 15740 3470
rect 15710 3420 15740 3450
rect 15710 3400 15715 3420
rect 15735 3400 15740 3420
rect 15710 3370 15740 3400
rect 15710 3350 15715 3370
rect 15735 3350 15740 3370
rect 15710 3320 15740 3350
rect 15710 3300 15715 3320
rect 15735 3300 15740 3320
rect 15710 3270 15740 3300
rect 15710 3250 15715 3270
rect 15735 3250 15740 3270
rect 15710 3220 15740 3250
rect 15710 3200 15715 3220
rect 15735 3200 15740 3220
rect 15710 3170 15740 3200
rect 15710 3150 15715 3170
rect 15735 3150 15740 3170
rect 15710 3120 15740 3150
rect 15710 3100 15715 3120
rect 15735 3100 15740 3120
rect 15710 3070 15740 3100
rect 15710 3050 15715 3070
rect 15735 3050 15740 3070
rect 15710 3020 15740 3050
rect 15710 3000 15715 3020
rect 15735 3000 15740 3020
rect 15710 2990 15740 3000
rect 15765 3570 15795 3580
rect 15765 3550 15770 3570
rect 15790 3550 15795 3570
rect 15765 3520 15795 3550
rect 15765 3500 15770 3520
rect 15790 3500 15795 3520
rect 15765 3470 15795 3500
rect 15765 3450 15770 3470
rect 15790 3450 15795 3470
rect 15765 3420 15795 3450
rect 15765 3400 15770 3420
rect 15790 3400 15795 3420
rect 15765 3370 15795 3400
rect 15765 3350 15770 3370
rect 15790 3350 15795 3370
rect 15765 3320 15795 3350
rect 15765 3300 15770 3320
rect 15790 3300 15795 3320
rect 15765 3270 15795 3300
rect 15765 3250 15770 3270
rect 15790 3250 15795 3270
rect 15765 3220 15795 3250
rect 15765 3200 15770 3220
rect 15790 3200 15795 3220
rect 15765 3170 15795 3200
rect 15765 3150 15770 3170
rect 15790 3150 15795 3170
rect 15765 3120 15795 3150
rect 15765 3100 15770 3120
rect 15790 3100 15795 3120
rect 15765 3070 15795 3100
rect 15765 3050 15770 3070
rect 15790 3050 15795 3070
rect 15765 3020 15795 3050
rect 15765 3000 15770 3020
rect 15790 3000 15795 3020
rect 15765 2990 15795 3000
rect 15820 3570 15890 3580
rect 16190 3570 16210 3590
rect 16350 3570 16370 3590
rect 16470 3570 16490 3590
rect 16590 3570 16610 3590
rect 16710 3570 16730 3590
rect 16830 3570 16850 3590
rect 16950 3570 16970 3590
rect 17070 3570 17090 3590
rect 17190 3570 17210 3590
rect 17310 3570 17330 3590
rect 17430 3570 17450 3590
rect 17590 3570 17610 3590
rect 18010 3580 18030 3600
rect 18120 3580 18140 3600
rect 18230 3580 18250 3600
rect 18340 3580 18360 3600
rect 18450 3580 18470 3600
rect 18560 3580 18580 3600
rect 17910 3570 17980 3580
rect 15820 3550 15825 3570
rect 15845 3550 15865 3570
rect 15885 3550 15890 3570
rect 15820 3520 15890 3550
rect 15820 3500 15825 3520
rect 15845 3500 15865 3520
rect 15885 3500 15890 3520
rect 15820 3470 15890 3500
rect 15820 3450 15825 3470
rect 15845 3450 15865 3470
rect 15885 3450 15890 3470
rect 15820 3420 15890 3450
rect 15820 3400 15825 3420
rect 15845 3400 15865 3420
rect 15885 3400 15890 3420
rect 15820 3370 15890 3400
rect 15820 3350 15825 3370
rect 15845 3350 15865 3370
rect 15885 3350 15890 3370
rect 15820 3320 15890 3350
rect 15820 3300 15825 3320
rect 15845 3300 15865 3320
rect 15885 3300 15890 3320
rect 15820 3270 15890 3300
rect 15820 3250 15825 3270
rect 15845 3250 15865 3270
rect 15885 3250 15890 3270
rect 15820 3220 15890 3250
rect 15820 3200 15825 3220
rect 15845 3200 15865 3220
rect 15885 3200 15890 3220
rect 15820 3170 15890 3200
rect 16185 3560 16255 3570
rect 16185 3540 16190 3560
rect 16210 3540 16230 3560
rect 16250 3540 16255 3560
rect 16185 3510 16255 3540
rect 16185 3490 16190 3510
rect 16210 3490 16230 3510
rect 16250 3490 16255 3510
rect 16185 3460 16255 3490
rect 16185 3440 16190 3460
rect 16210 3440 16230 3460
rect 16250 3440 16255 3460
rect 16185 3410 16255 3440
rect 16185 3390 16190 3410
rect 16210 3390 16230 3410
rect 16250 3390 16255 3410
rect 16185 3360 16255 3390
rect 16185 3340 16190 3360
rect 16210 3340 16230 3360
rect 16250 3340 16255 3360
rect 16185 3310 16255 3340
rect 16185 3290 16190 3310
rect 16210 3290 16230 3310
rect 16250 3290 16255 3310
rect 16185 3260 16255 3290
rect 16185 3240 16190 3260
rect 16210 3240 16230 3260
rect 16250 3240 16255 3260
rect 16185 3210 16255 3240
rect 16185 3190 16190 3210
rect 16210 3190 16230 3210
rect 16250 3190 16255 3210
rect 16185 3180 16255 3190
rect 16285 3560 16315 3570
rect 16285 3540 16290 3560
rect 16310 3540 16315 3560
rect 16285 3510 16315 3540
rect 16285 3490 16290 3510
rect 16310 3490 16315 3510
rect 16285 3460 16315 3490
rect 16285 3440 16290 3460
rect 16310 3440 16315 3460
rect 16285 3410 16315 3440
rect 16285 3390 16290 3410
rect 16310 3390 16315 3410
rect 16285 3360 16315 3390
rect 16285 3340 16290 3360
rect 16310 3340 16315 3360
rect 16285 3310 16315 3340
rect 16285 3290 16290 3310
rect 16310 3290 16315 3310
rect 16285 3260 16315 3290
rect 16285 3240 16290 3260
rect 16310 3240 16315 3260
rect 16285 3210 16315 3240
rect 16285 3190 16290 3210
rect 16310 3190 16315 3210
rect 16285 3180 16315 3190
rect 16345 3560 16375 3570
rect 16345 3540 16350 3560
rect 16370 3540 16375 3560
rect 16345 3510 16375 3540
rect 16345 3490 16350 3510
rect 16370 3490 16375 3510
rect 16345 3460 16375 3490
rect 16345 3440 16350 3460
rect 16370 3440 16375 3460
rect 16345 3410 16375 3440
rect 16345 3390 16350 3410
rect 16370 3390 16375 3410
rect 16345 3360 16375 3390
rect 16345 3340 16350 3360
rect 16370 3340 16375 3360
rect 16345 3310 16375 3340
rect 16345 3290 16350 3310
rect 16370 3290 16375 3310
rect 16345 3260 16375 3290
rect 16345 3240 16350 3260
rect 16370 3240 16375 3260
rect 16345 3210 16375 3240
rect 16345 3190 16350 3210
rect 16370 3190 16375 3210
rect 16345 3180 16375 3190
rect 16405 3560 16435 3570
rect 16405 3540 16410 3560
rect 16430 3540 16435 3560
rect 16405 3510 16435 3540
rect 16405 3490 16410 3510
rect 16430 3490 16435 3510
rect 16405 3460 16435 3490
rect 16405 3440 16410 3460
rect 16430 3440 16435 3460
rect 16405 3410 16435 3440
rect 16405 3390 16410 3410
rect 16430 3390 16435 3410
rect 16405 3360 16435 3390
rect 16405 3340 16410 3360
rect 16430 3340 16435 3360
rect 16405 3310 16435 3340
rect 16405 3290 16410 3310
rect 16430 3290 16435 3310
rect 16405 3260 16435 3290
rect 16405 3240 16410 3260
rect 16430 3240 16435 3260
rect 16405 3210 16435 3240
rect 16405 3190 16410 3210
rect 16430 3190 16435 3210
rect 16405 3180 16435 3190
rect 16465 3560 16495 3570
rect 16465 3540 16470 3560
rect 16490 3540 16495 3560
rect 16465 3510 16495 3540
rect 16465 3490 16470 3510
rect 16490 3490 16495 3510
rect 16465 3460 16495 3490
rect 16465 3440 16470 3460
rect 16490 3440 16495 3460
rect 16465 3410 16495 3440
rect 16465 3390 16470 3410
rect 16490 3390 16495 3410
rect 16465 3360 16495 3390
rect 16465 3340 16470 3360
rect 16490 3340 16495 3360
rect 16465 3310 16495 3340
rect 16465 3290 16470 3310
rect 16490 3290 16495 3310
rect 16465 3260 16495 3290
rect 16465 3240 16470 3260
rect 16490 3240 16495 3260
rect 16465 3210 16495 3240
rect 16465 3190 16470 3210
rect 16490 3190 16495 3210
rect 16465 3180 16495 3190
rect 16525 3560 16555 3570
rect 16525 3540 16530 3560
rect 16550 3540 16555 3560
rect 16525 3510 16555 3540
rect 16525 3490 16530 3510
rect 16550 3490 16555 3510
rect 16525 3460 16555 3490
rect 16525 3440 16530 3460
rect 16550 3440 16555 3460
rect 16525 3410 16555 3440
rect 16525 3390 16530 3410
rect 16550 3390 16555 3410
rect 16525 3360 16555 3390
rect 16525 3340 16530 3360
rect 16550 3340 16555 3360
rect 16525 3310 16555 3340
rect 16525 3290 16530 3310
rect 16550 3290 16555 3310
rect 16525 3260 16555 3290
rect 16525 3240 16530 3260
rect 16550 3240 16555 3260
rect 16525 3210 16555 3240
rect 16525 3190 16530 3210
rect 16550 3190 16555 3210
rect 16525 3180 16555 3190
rect 16585 3560 16615 3570
rect 16585 3540 16590 3560
rect 16610 3540 16615 3560
rect 16585 3510 16615 3540
rect 16585 3490 16590 3510
rect 16610 3490 16615 3510
rect 16585 3460 16615 3490
rect 16585 3440 16590 3460
rect 16610 3440 16615 3460
rect 16585 3410 16615 3440
rect 16585 3390 16590 3410
rect 16610 3390 16615 3410
rect 16585 3360 16615 3390
rect 16585 3340 16590 3360
rect 16610 3340 16615 3360
rect 16585 3310 16615 3340
rect 16585 3290 16590 3310
rect 16610 3290 16615 3310
rect 16585 3260 16615 3290
rect 16585 3240 16590 3260
rect 16610 3240 16615 3260
rect 16585 3210 16615 3240
rect 16585 3190 16590 3210
rect 16610 3190 16615 3210
rect 16585 3180 16615 3190
rect 16645 3560 16675 3570
rect 16645 3540 16650 3560
rect 16670 3540 16675 3560
rect 16645 3510 16675 3540
rect 16645 3490 16650 3510
rect 16670 3490 16675 3510
rect 16645 3460 16675 3490
rect 16645 3440 16650 3460
rect 16670 3440 16675 3460
rect 16645 3410 16675 3440
rect 16645 3390 16650 3410
rect 16670 3390 16675 3410
rect 16645 3360 16675 3390
rect 16645 3340 16650 3360
rect 16670 3340 16675 3360
rect 16645 3310 16675 3340
rect 16645 3290 16650 3310
rect 16670 3290 16675 3310
rect 16645 3260 16675 3290
rect 16645 3240 16650 3260
rect 16670 3240 16675 3260
rect 16645 3210 16675 3240
rect 16645 3190 16650 3210
rect 16670 3190 16675 3210
rect 16645 3180 16675 3190
rect 16705 3560 16735 3570
rect 16705 3540 16710 3560
rect 16730 3540 16735 3560
rect 16705 3510 16735 3540
rect 16705 3490 16710 3510
rect 16730 3490 16735 3510
rect 16705 3460 16735 3490
rect 16705 3440 16710 3460
rect 16730 3440 16735 3460
rect 16705 3410 16735 3440
rect 16705 3390 16710 3410
rect 16730 3390 16735 3410
rect 16705 3360 16735 3390
rect 16705 3340 16710 3360
rect 16730 3340 16735 3360
rect 16705 3310 16735 3340
rect 16705 3290 16710 3310
rect 16730 3290 16735 3310
rect 16705 3260 16735 3290
rect 16705 3240 16710 3260
rect 16730 3240 16735 3260
rect 16705 3210 16735 3240
rect 16705 3190 16710 3210
rect 16730 3190 16735 3210
rect 16705 3180 16735 3190
rect 16765 3560 16795 3570
rect 16765 3540 16770 3560
rect 16790 3540 16795 3560
rect 16765 3510 16795 3540
rect 16765 3490 16770 3510
rect 16790 3490 16795 3510
rect 16765 3460 16795 3490
rect 16765 3440 16770 3460
rect 16790 3440 16795 3460
rect 16765 3410 16795 3440
rect 16765 3390 16770 3410
rect 16790 3390 16795 3410
rect 16765 3360 16795 3390
rect 16765 3340 16770 3360
rect 16790 3340 16795 3360
rect 16765 3310 16795 3340
rect 16765 3290 16770 3310
rect 16790 3290 16795 3310
rect 16765 3260 16795 3290
rect 16765 3240 16770 3260
rect 16790 3240 16795 3260
rect 16765 3210 16795 3240
rect 16765 3190 16770 3210
rect 16790 3190 16795 3210
rect 16765 3180 16795 3190
rect 16825 3560 16855 3570
rect 16825 3540 16830 3560
rect 16850 3540 16855 3560
rect 16825 3510 16855 3540
rect 16825 3490 16830 3510
rect 16850 3490 16855 3510
rect 16825 3460 16855 3490
rect 16825 3440 16830 3460
rect 16850 3440 16855 3460
rect 16825 3410 16855 3440
rect 16825 3390 16830 3410
rect 16850 3390 16855 3410
rect 16825 3360 16855 3390
rect 16825 3340 16830 3360
rect 16850 3340 16855 3360
rect 16825 3310 16855 3340
rect 16825 3290 16830 3310
rect 16850 3290 16855 3310
rect 16825 3260 16855 3290
rect 16825 3240 16830 3260
rect 16850 3240 16855 3260
rect 16825 3210 16855 3240
rect 16825 3190 16830 3210
rect 16850 3190 16855 3210
rect 16825 3180 16855 3190
rect 16885 3560 16915 3570
rect 16885 3540 16890 3560
rect 16910 3540 16915 3560
rect 16885 3510 16915 3540
rect 16885 3490 16890 3510
rect 16910 3490 16915 3510
rect 16885 3460 16915 3490
rect 16885 3440 16890 3460
rect 16910 3440 16915 3460
rect 16885 3410 16915 3440
rect 16885 3390 16890 3410
rect 16910 3390 16915 3410
rect 16885 3360 16915 3390
rect 16885 3340 16890 3360
rect 16910 3340 16915 3360
rect 16885 3310 16915 3340
rect 16885 3290 16890 3310
rect 16910 3290 16915 3310
rect 16885 3260 16915 3290
rect 16885 3240 16890 3260
rect 16910 3240 16915 3260
rect 16885 3210 16915 3240
rect 16885 3190 16890 3210
rect 16910 3190 16915 3210
rect 16885 3180 16915 3190
rect 16945 3560 16975 3570
rect 16945 3540 16950 3560
rect 16970 3540 16975 3560
rect 16945 3510 16975 3540
rect 16945 3490 16950 3510
rect 16970 3490 16975 3510
rect 16945 3460 16975 3490
rect 16945 3440 16950 3460
rect 16970 3440 16975 3460
rect 16945 3410 16975 3440
rect 16945 3390 16950 3410
rect 16970 3390 16975 3410
rect 16945 3360 16975 3390
rect 16945 3340 16950 3360
rect 16970 3340 16975 3360
rect 16945 3310 16975 3340
rect 16945 3290 16950 3310
rect 16970 3290 16975 3310
rect 16945 3260 16975 3290
rect 16945 3240 16950 3260
rect 16970 3240 16975 3260
rect 16945 3210 16975 3240
rect 16945 3190 16950 3210
rect 16970 3190 16975 3210
rect 16945 3180 16975 3190
rect 17005 3560 17035 3570
rect 17005 3540 17010 3560
rect 17030 3540 17035 3560
rect 17005 3510 17035 3540
rect 17005 3490 17010 3510
rect 17030 3490 17035 3510
rect 17005 3460 17035 3490
rect 17005 3440 17010 3460
rect 17030 3440 17035 3460
rect 17005 3410 17035 3440
rect 17005 3390 17010 3410
rect 17030 3390 17035 3410
rect 17005 3360 17035 3390
rect 17005 3340 17010 3360
rect 17030 3340 17035 3360
rect 17005 3310 17035 3340
rect 17005 3290 17010 3310
rect 17030 3290 17035 3310
rect 17005 3260 17035 3290
rect 17005 3240 17010 3260
rect 17030 3240 17035 3260
rect 17005 3210 17035 3240
rect 17005 3190 17010 3210
rect 17030 3190 17035 3210
rect 17005 3180 17035 3190
rect 17065 3560 17095 3570
rect 17065 3540 17070 3560
rect 17090 3540 17095 3560
rect 17065 3510 17095 3540
rect 17065 3490 17070 3510
rect 17090 3490 17095 3510
rect 17065 3460 17095 3490
rect 17065 3440 17070 3460
rect 17090 3440 17095 3460
rect 17065 3410 17095 3440
rect 17065 3390 17070 3410
rect 17090 3390 17095 3410
rect 17065 3360 17095 3390
rect 17065 3340 17070 3360
rect 17090 3340 17095 3360
rect 17065 3310 17095 3340
rect 17065 3290 17070 3310
rect 17090 3290 17095 3310
rect 17065 3260 17095 3290
rect 17065 3240 17070 3260
rect 17090 3240 17095 3260
rect 17065 3210 17095 3240
rect 17065 3190 17070 3210
rect 17090 3190 17095 3210
rect 17065 3180 17095 3190
rect 17125 3560 17155 3570
rect 17125 3540 17130 3560
rect 17150 3540 17155 3560
rect 17125 3510 17155 3540
rect 17125 3490 17130 3510
rect 17150 3490 17155 3510
rect 17125 3460 17155 3490
rect 17125 3440 17130 3460
rect 17150 3440 17155 3460
rect 17125 3410 17155 3440
rect 17125 3390 17130 3410
rect 17150 3390 17155 3410
rect 17125 3360 17155 3390
rect 17125 3340 17130 3360
rect 17150 3340 17155 3360
rect 17125 3310 17155 3340
rect 17125 3290 17130 3310
rect 17150 3290 17155 3310
rect 17125 3260 17155 3290
rect 17125 3240 17130 3260
rect 17150 3240 17155 3260
rect 17125 3210 17155 3240
rect 17125 3190 17130 3210
rect 17150 3190 17155 3210
rect 17125 3180 17155 3190
rect 17185 3560 17215 3570
rect 17185 3540 17190 3560
rect 17210 3540 17215 3560
rect 17185 3510 17215 3540
rect 17185 3490 17190 3510
rect 17210 3490 17215 3510
rect 17185 3460 17215 3490
rect 17185 3440 17190 3460
rect 17210 3440 17215 3460
rect 17185 3410 17215 3440
rect 17185 3390 17190 3410
rect 17210 3390 17215 3410
rect 17185 3360 17215 3390
rect 17185 3340 17190 3360
rect 17210 3340 17215 3360
rect 17185 3310 17215 3340
rect 17185 3290 17190 3310
rect 17210 3290 17215 3310
rect 17185 3260 17215 3290
rect 17185 3240 17190 3260
rect 17210 3240 17215 3260
rect 17185 3210 17215 3240
rect 17185 3190 17190 3210
rect 17210 3190 17215 3210
rect 17185 3180 17215 3190
rect 17245 3560 17275 3570
rect 17245 3540 17250 3560
rect 17270 3540 17275 3560
rect 17245 3510 17275 3540
rect 17245 3490 17250 3510
rect 17270 3490 17275 3510
rect 17245 3460 17275 3490
rect 17245 3440 17250 3460
rect 17270 3440 17275 3460
rect 17245 3410 17275 3440
rect 17245 3390 17250 3410
rect 17270 3390 17275 3410
rect 17245 3360 17275 3390
rect 17245 3340 17250 3360
rect 17270 3340 17275 3360
rect 17245 3310 17275 3340
rect 17245 3290 17250 3310
rect 17270 3290 17275 3310
rect 17245 3260 17275 3290
rect 17245 3240 17250 3260
rect 17270 3240 17275 3260
rect 17245 3210 17275 3240
rect 17245 3190 17250 3210
rect 17270 3190 17275 3210
rect 17245 3180 17275 3190
rect 17305 3560 17335 3570
rect 17305 3540 17310 3560
rect 17330 3540 17335 3560
rect 17305 3510 17335 3540
rect 17305 3490 17310 3510
rect 17330 3490 17335 3510
rect 17305 3460 17335 3490
rect 17305 3440 17310 3460
rect 17330 3440 17335 3460
rect 17305 3410 17335 3440
rect 17305 3390 17310 3410
rect 17330 3390 17335 3410
rect 17305 3360 17335 3390
rect 17305 3340 17310 3360
rect 17330 3340 17335 3360
rect 17305 3310 17335 3340
rect 17305 3290 17310 3310
rect 17330 3290 17335 3310
rect 17305 3260 17335 3290
rect 17305 3240 17310 3260
rect 17330 3240 17335 3260
rect 17305 3210 17335 3240
rect 17305 3190 17310 3210
rect 17330 3190 17335 3210
rect 17305 3180 17335 3190
rect 17365 3560 17395 3570
rect 17365 3540 17370 3560
rect 17390 3540 17395 3560
rect 17365 3510 17395 3540
rect 17365 3490 17370 3510
rect 17390 3490 17395 3510
rect 17365 3460 17395 3490
rect 17365 3440 17370 3460
rect 17390 3440 17395 3460
rect 17365 3410 17395 3440
rect 17365 3390 17370 3410
rect 17390 3390 17395 3410
rect 17365 3360 17395 3390
rect 17365 3340 17370 3360
rect 17390 3340 17395 3360
rect 17365 3310 17395 3340
rect 17365 3290 17370 3310
rect 17390 3290 17395 3310
rect 17365 3260 17395 3290
rect 17365 3240 17370 3260
rect 17390 3240 17395 3260
rect 17365 3210 17395 3240
rect 17365 3190 17370 3210
rect 17390 3190 17395 3210
rect 17365 3180 17395 3190
rect 17425 3560 17455 3570
rect 17425 3540 17430 3560
rect 17450 3540 17455 3560
rect 17425 3510 17455 3540
rect 17425 3490 17430 3510
rect 17450 3490 17455 3510
rect 17425 3460 17455 3490
rect 17425 3440 17430 3460
rect 17450 3440 17455 3460
rect 17425 3410 17455 3440
rect 17425 3390 17430 3410
rect 17450 3390 17455 3410
rect 17425 3360 17455 3390
rect 17425 3340 17430 3360
rect 17450 3340 17455 3360
rect 17425 3310 17455 3340
rect 17425 3290 17430 3310
rect 17450 3290 17455 3310
rect 17425 3260 17455 3290
rect 17425 3240 17430 3260
rect 17450 3240 17455 3260
rect 17425 3210 17455 3240
rect 17425 3190 17430 3210
rect 17450 3190 17455 3210
rect 17425 3180 17455 3190
rect 17485 3560 17515 3570
rect 17485 3540 17490 3560
rect 17510 3540 17515 3560
rect 17485 3510 17515 3540
rect 17485 3490 17490 3510
rect 17510 3490 17515 3510
rect 17485 3460 17515 3490
rect 17485 3440 17490 3460
rect 17510 3440 17515 3460
rect 17485 3410 17515 3440
rect 17485 3390 17490 3410
rect 17510 3390 17515 3410
rect 17485 3360 17515 3390
rect 17485 3340 17490 3360
rect 17510 3340 17515 3360
rect 17485 3310 17515 3340
rect 17485 3290 17490 3310
rect 17510 3290 17515 3310
rect 17485 3260 17515 3290
rect 17485 3240 17490 3260
rect 17510 3240 17515 3260
rect 17485 3210 17515 3240
rect 17485 3190 17490 3210
rect 17510 3190 17515 3210
rect 17485 3180 17515 3190
rect 17545 3560 17615 3570
rect 17545 3540 17550 3560
rect 17570 3540 17590 3560
rect 17610 3540 17615 3560
rect 17545 3510 17615 3540
rect 17545 3490 17550 3510
rect 17570 3490 17590 3510
rect 17610 3490 17615 3510
rect 17545 3460 17615 3490
rect 17545 3440 17550 3460
rect 17570 3440 17590 3460
rect 17610 3440 17615 3460
rect 17545 3410 17615 3440
rect 17545 3390 17550 3410
rect 17570 3390 17590 3410
rect 17610 3390 17615 3410
rect 17545 3360 17615 3390
rect 17545 3340 17550 3360
rect 17570 3340 17590 3360
rect 17610 3340 17615 3360
rect 17545 3310 17615 3340
rect 17545 3290 17550 3310
rect 17570 3290 17590 3310
rect 17610 3290 17615 3310
rect 17545 3260 17615 3290
rect 17545 3240 17550 3260
rect 17570 3240 17590 3260
rect 17610 3240 17615 3260
rect 17545 3210 17615 3240
rect 17545 3190 17550 3210
rect 17570 3190 17590 3210
rect 17610 3190 17615 3210
rect 17545 3180 17615 3190
rect 17910 3550 17915 3570
rect 17935 3550 17955 3570
rect 17975 3550 17980 3570
rect 17910 3520 17980 3550
rect 17910 3500 17915 3520
rect 17935 3500 17955 3520
rect 17975 3500 17980 3520
rect 17910 3470 17980 3500
rect 17910 3450 17915 3470
rect 17935 3450 17955 3470
rect 17975 3450 17980 3470
rect 17910 3420 17980 3450
rect 17910 3400 17915 3420
rect 17935 3400 17955 3420
rect 17975 3400 17980 3420
rect 17910 3370 17980 3400
rect 17910 3350 17915 3370
rect 17935 3350 17955 3370
rect 17975 3350 17980 3370
rect 17910 3320 17980 3350
rect 17910 3300 17915 3320
rect 17935 3300 17955 3320
rect 17975 3300 17980 3320
rect 17910 3270 17980 3300
rect 17910 3250 17915 3270
rect 17935 3250 17955 3270
rect 17975 3250 17980 3270
rect 17910 3220 17980 3250
rect 17910 3200 17915 3220
rect 17935 3200 17955 3220
rect 17975 3200 17980 3220
rect 15820 3150 15825 3170
rect 15845 3150 15865 3170
rect 15885 3150 15890 3170
rect 16290 3160 16310 3180
rect 16410 3160 16430 3180
rect 16530 3160 16550 3180
rect 16650 3160 16670 3180
rect 16770 3160 16790 3180
rect 16890 3160 16910 3180
rect 17010 3160 17030 3180
rect 17130 3160 17150 3180
rect 17250 3160 17270 3180
rect 17370 3160 17390 3180
rect 17490 3160 17510 3180
rect 17910 3170 17980 3200
rect 15820 3120 15890 3150
rect 16280 3150 16320 3160
rect 16280 3130 16290 3150
rect 16310 3130 16320 3150
rect 16280 3120 16320 3130
rect 16400 3150 16440 3160
rect 16400 3130 16410 3150
rect 16430 3130 16440 3150
rect 16400 3120 16440 3130
rect 16520 3150 16560 3160
rect 16520 3130 16530 3150
rect 16550 3130 16560 3150
rect 16520 3120 16560 3130
rect 16640 3150 16680 3160
rect 16640 3130 16650 3150
rect 16670 3130 16680 3150
rect 16640 3120 16680 3130
rect 16760 3150 16800 3160
rect 16760 3130 16770 3150
rect 16790 3130 16800 3150
rect 16760 3120 16800 3130
rect 16823 3150 16857 3160
rect 16823 3130 16831 3150
rect 16849 3130 16857 3150
rect 16823 3120 16857 3130
rect 16880 3150 16920 3160
rect 16880 3130 16890 3150
rect 16910 3130 16920 3150
rect 16880 3120 16920 3130
rect 17000 3150 17040 3160
rect 17000 3130 17010 3150
rect 17030 3130 17040 3150
rect 17000 3120 17040 3130
rect 17120 3150 17160 3160
rect 17120 3130 17130 3150
rect 17150 3130 17160 3150
rect 17120 3120 17160 3130
rect 17240 3150 17280 3160
rect 17240 3130 17250 3150
rect 17270 3130 17280 3150
rect 17240 3120 17280 3130
rect 17360 3150 17400 3160
rect 17360 3130 17370 3150
rect 17390 3130 17400 3150
rect 17360 3120 17400 3130
rect 17480 3150 17520 3160
rect 17480 3130 17490 3150
rect 17510 3130 17520 3150
rect 17480 3120 17520 3130
rect 17910 3150 17915 3170
rect 17935 3150 17955 3170
rect 17975 3150 17980 3170
rect 17910 3120 17980 3150
rect 15820 3100 15825 3120
rect 15845 3100 15865 3120
rect 15885 3100 15890 3120
rect 15820 3070 15890 3100
rect 15820 3050 15825 3070
rect 15845 3050 15865 3070
rect 15885 3050 15890 3070
rect 15820 3020 15890 3050
rect 15820 3000 15825 3020
rect 15845 3000 15865 3020
rect 15885 3000 15890 3020
rect 15820 2990 15890 3000
rect 17910 3100 17915 3120
rect 17935 3100 17955 3120
rect 17975 3100 17980 3120
rect 17910 3070 17980 3100
rect 17910 3050 17915 3070
rect 17935 3050 17955 3070
rect 17975 3050 17980 3070
rect 17910 3020 17980 3050
rect 17910 3000 17915 3020
rect 17935 3000 17955 3020
rect 17975 3000 17980 3020
rect 17910 2990 17980 3000
rect 18005 3570 18035 3580
rect 18005 3550 18010 3570
rect 18030 3550 18035 3570
rect 18005 3520 18035 3550
rect 18005 3500 18010 3520
rect 18030 3500 18035 3520
rect 18005 3470 18035 3500
rect 18005 3450 18010 3470
rect 18030 3450 18035 3470
rect 18005 3420 18035 3450
rect 18005 3400 18010 3420
rect 18030 3400 18035 3420
rect 18005 3370 18035 3400
rect 18005 3350 18010 3370
rect 18030 3350 18035 3370
rect 18005 3320 18035 3350
rect 18005 3300 18010 3320
rect 18030 3300 18035 3320
rect 18005 3270 18035 3300
rect 18005 3250 18010 3270
rect 18030 3250 18035 3270
rect 18005 3220 18035 3250
rect 18005 3200 18010 3220
rect 18030 3200 18035 3220
rect 18005 3170 18035 3200
rect 18005 3150 18010 3170
rect 18030 3150 18035 3170
rect 18005 3120 18035 3150
rect 18005 3100 18010 3120
rect 18030 3100 18035 3120
rect 18005 3070 18035 3100
rect 18005 3050 18010 3070
rect 18030 3050 18035 3070
rect 18005 3020 18035 3050
rect 18005 3000 18010 3020
rect 18030 3000 18035 3020
rect 18005 2990 18035 3000
rect 18060 3570 18090 3580
rect 18060 3550 18065 3570
rect 18085 3550 18090 3570
rect 18060 3520 18090 3550
rect 18060 3500 18065 3520
rect 18085 3500 18090 3520
rect 18060 3470 18090 3500
rect 18060 3450 18065 3470
rect 18085 3450 18090 3470
rect 18060 3420 18090 3450
rect 18060 3400 18065 3420
rect 18085 3400 18090 3420
rect 18060 3370 18090 3400
rect 18060 3350 18065 3370
rect 18085 3350 18090 3370
rect 18060 3320 18090 3350
rect 18060 3300 18065 3320
rect 18085 3300 18090 3320
rect 18060 3270 18090 3300
rect 18060 3250 18065 3270
rect 18085 3250 18090 3270
rect 18060 3220 18090 3250
rect 18060 3200 18065 3220
rect 18085 3200 18090 3220
rect 18060 3170 18090 3200
rect 18060 3150 18065 3170
rect 18085 3150 18090 3170
rect 18060 3120 18090 3150
rect 18060 3100 18065 3120
rect 18085 3100 18090 3120
rect 18060 3070 18090 3100
rect 18060 3050 18065 3070
rect 18085 3050 18090 3070
rect 18060 3020 18090 3050
rect 18060 3000 18065 3020
rect 18085 3000 18090 3020
rect 18060 2990 18090 3000
rect 18115 3570 18145 3580
rect 18115 3550 18120 3570
rect 18140 3550 18145 3570
rect 18115 3520 18145 3550
rect 18115 3500 18120 3520
rect 18140 3500 18145 3520
rect 18115 3470 18145 3500
rect 18115 3450 18120 3470
rect 18140 3450 18145 3470
rect 18115 3420 18145 3450
rect 18115 3400 18120 3420
rect 18140 3400 18145 3420
rect 18115 3370 18145 3400
rect 18115 3350 18120 3370
rect 18140 3350 18145 3370
rect 18115 3320 18145 3350
rect 18115 3300 18120 3320
rect 18140 3300 18145 3320
rect 18115 3270 18145 3300
rect 18115 3250 18120 3270
rect 18140 3250 18145 3270
rect 18115 3220 18145 3250
rect 18115 3200 18120 3220
rect 18140 3200 18145 3220
rect 18115 3170 18145 3200
rect 18115 3150 18120 3170
rect 18140 3150 18145 3170
rect 18115 3120 18145 3150
rect 18115 3100 18120 3120
rect 18140 3100 18145 3120
rect 18115 3070 18145 3100
rect 18115 3050 18120 3070
rect 18140 3050 18145 3070
rect 18115 3020 18145 3050
rect 18115 3000 18120 3020
rect 18140 3000 18145 3020
rect 18115 2990 18145 3000
rect 18170 3570 18200 3580
rect 18170 3550 18175 3570
rect 18195 3550 18200 3570
rect 18170 3520 18200 3550
rect 18170 3500 18175 3520
rect 18195 3500 18200 3520
rect 18170 3470 18200 3500
rect 18170 3450 18175 3470
rect 18195 3450 18200 3470
rect 18170 3420 18200 3450
rect 18170 3400 18175 3420
rect 18195 3400 18200 3420
rect 18170 3370 18200 3400
rect 18170 3350 18175 3370
rect 18195 3350 18200 3370
rect 18170 3320 18200 3350
rect 18170 3300 18175 3320
rect 18195 3300 18200 3320
rect 18170 3270 18200 3300
rect 18170 3250 18175 3270
rect 18195 3250 18200 3270
rect 18170 3220 18200 3250
rect 18170 3200 18175 3220
rect 18195 3200 18200 3220
rect 18170 3170 18200 3200
rect 18170 3150 18175 3170
rect 18195 3150 18200 3170
rect 18170 3120 18200 3150
rect 18170 3100 18175 3120
rect 18195 3100 18200 3120
rect 18170 3070 18200 3100
rect 18170 3050 18175 3070
rect 18195 3050 18200 3070
rect 18170 3020 18200 3050
rect 18170 3000 18175 3020
rect 18195 3000 18200 3020
rect 18170 2990 18200 3000
rect 18225 3570 18255 3580
rect 18225 3550 18230 3570
rect 18250 3550 18255 3570
rect 18225 3520 18255 3550
rect 18225 3500 18230 3520
rect 18250 3500 18255 3520
rect 18225 3470 18255 3500
rect 18225 3450 18230 3470
rect 18250 3450 18255 3470
rect 18225 3420 18255 3450
rect 18225 3400 18230 3420
rect 18250 3400 18255 3420
rect 18225 3370 18255 3400
rect 18225 3350 18230 3370
rect 18250 3350 18255 3370
rect 18225 3320 18255 3350
rect 18225 3300 18230 3320
rect 18250 3300 18255 3320
rect 18225 3270 18255 3300
rect 18225 3250 18230 3270
rect 18250 3250 18255 3270
rect 18225 3220 18255 3250
rect 18225 3200 18230 3220
rect 18250 3200 18255 3220
rect 18225 3170 18255 3200
rect 18225 3150 18230 3170
rect 18250 3150 18255 3170
rect 18225 3120 18255 3150
rect 18225 3100 18230 3120
rect 18250 3100 18255 3120
rect 18225 3070 18255 3100
rect 18225 3050 18230 3070
rect 18250 3050 18255 3070
rect 18225 3020 18255 3050
rect 18225 3000 18230 3020
rect 18250 3000 18255 3020
rect 18225 2990 18255 3000
rect 18280 3570 18310 3580
rect 18280 3550 18285 3570
rect 18305 3550 18310 3570
rect 18280 3520 18310 3550
rect 18280 3500 18285 3520
rect 18305 3500 18310 3520
rect 18280 3470 18310 3500
rect 18280 3450 18285 3470
rect 18305 3450 18310 3470
rect 18280 3420 18310 3450
rect 18280 3400 18285 3420
rect 18305 3400 18310 3420
rect 18280 3370 18310 3400
rect 18280 3350 18285 3370
rect 18305 3350 18310 3370
rect 18280 3320 18310 3350
rect 18280 3300 18285 3320
rect 18305 3300 18310 3320
rect 18280 3270 18310 3300
rect 18280 3250 18285 3270
rect 18305 3250 18310 3270
rect 18280 3220 18310 3250
rect 18280 3200 18285 3220
rect 18305 3200 18310 3220
rect 18280 3170 18310 3200
rect 18280 3150 18285 3170
rect 18305 3150 18310 3170
rect 18280 3120 18310 3150
rect 18280 3100 18285 3120
rect 18305 3100 18310 3120
rect 18280 3070 18310 3100
rect 18280 3050 18285 3070
rect 18305 3050 18310 3070
rect 18280 3020 18310 3050
rect 18280 3000 18285 3020
rect 18305 3000 18310 3020
rect 18280 2990 18310 3000
rect 18335 3570 18365 3580
rect 18335 3550 18340 3570
rect 18360 3550 18365 3570
rect 18335 3520 18365 3550
rect 18335 3500 18340 3520
rect 18360 3500 18365 3520
rect 18335 3470 18365 3500
rect 18335 3450 18340 3470
rect 18360 3450 18365 3470
rect 18335 3420 18365 3450
rect 18335 3400 18340 3420
rect 18360 3400 18365 3420
rect 18335 3370 18365 3400
rect 18335 3350 18340 3370
rect 18360 3350 18365 3370
rect 18335 3320 18365 3350
rect 18335 3300 18340 3320
rect 18360 3300 18365 3320
rect 18335 3270 18365 3300
rect 18335 3250 18340 3270
rect 18360 3250 18365 3270
rect 18335 3220 18365 3250
rect 18335 3200 18340 3220
rect 18360 3200 18365 3220
rect 18335 3170 18365 3200
rect 18335 3150 18340 3170
rect 18360 3150 18365 3170
rect 18335 3120 18365 3150
rect 18335 3100 18340 3120
rect 18360 3100 18365 3120
rect 18335 3070 18365 3100
rect 18335 3050 18340 3070
rect 18360 3050 18365 3070
rect 18335 3020 18365 3050
rect 18335 3000 18340 3020
rect 18360 3000 18365 3020
rect 18335 2990 18365 3000
rect 18390 3570 18420 3580
rect 18390 3550 18395 3570
rect 18415 3550 18420 3570
rect 18390 3520 18420 3550
rect 18390 3500 18395 3520
rect 18415 3500 18420 3520
rect 18390 3470 18420 3500
rect 18390 3450 18395 3470
rect 18415 3450 18420 3470
rect 18390 3420 18420 3450
rect 18390 3400 18395 3420
rect 18415 3400 18420 3420
rect 18390 3370 18420 3400
rect 18390 3350 18395 3370
rect 18415 3350 18420 3370
rect 18390 3320 18420 3350
rect 18390 3300 18395 3320
rect 18415 3300 18420 3320
rect 18390 3270 18420 3300
rect 18390 3250 18395 3270
rect 18415 3250 18420 3270
rect 18390 3220 18420 3250
rect 18390 3200 18395 3220
rect 18415 3200 18420 3220
rect 18390 3170 18420 3200
rect 18390 3150 18395 3170
rect 18415 3150 18420 3170
rect 18390 3120 18420 3150
rect 18390 3100 18395 3120
rect 18415 3100 18420 3120
rect 18390 3070 18420 3100
rect 18390 3050 18395 3070
rect 18415 3050 18420 3070
rect 18390 3020 18420 3050
rect 18390 3000 18395 3020
rect 18415 3000 18420 3020
rect 18390 2990 18420 3000
rect 18445 3570 18475 3580
rect 18445 3550 18450 3570
rect 18470 3550 18475 3570
rect 18445 3520 18475 3550
rect 18445 3500 18450 3520
rect 18470 3500 18475 3520
rect 18445 3470 18475 3500
rect 18445 3450 18450 3470
rect 18470 3450 18475 3470
rect 18445 3420 18475 3450
rect 18445 3400 18450 3420
rect 18470 3400 18475 3420
rect 18445 3370 18475 3400
rect 18445 3350 18450 3370
rect 18470 3350 18475 3370
rect 18445 3320 18475 3350
rect 18445 3300 18450 3320
rect 18470 3300 18475 3320
rect 18445 3270 18475 3300
rect 18445 3250 18450 3270
rect 18470 3250 18475 3270
rect 18445 3220 18475 3250
rect 18445 3200 18450 3220
rect 18470 3200 18475 3220
rect 18445 3170 18475 3200
rect 18445 3150 18450 3170
rect 18470 3150 18475 3170
rect 18445 3120 18475 3150
rect 18445 3100 18450 3120
rect 18470 3100 18475 3120
rect 18445 3070 18475 3100
rect 18445 3050 18450 3070
rect 18470 3050 18475 3070
rect 18445 3020 18475 3050
rect 18445 3000 18450 3020
rect 18470 3000 18475 3020
rect 18445 2990 18475 3000
rect 18500 3570 18530 3580
rect 18500 3550 18505 3570
rect 18525 3550 18530 3570
rect 18500 3520 18530 3550
rect 18500 3500 18505 3520
rect 18525 3500 18530 3520
rect 18500 3470 18530 3500
rect 18500 3450 18505 3470
rect 18525 3450 18530 3470
rect 18500 3420 18530 3450
rect 18500 3400 18505 3420
rect 18525 3400 18530 3420
rect 18500 3370 18530 3400
rect 18500 3350 18505 3370
rect 18525 3350 18530 3370
rect 18500 3320 18530 3350
rect 18500 3300 18505 3320
rect 18525 3300 18530 3320
rect 18500 3270 18530 3300
rect 18500 3250 18505 3270
rect 18525 3250 18530 3270
rect 18500 3220 18530 3250
rect 18500 3200 18505 3220
rect 18525 3200 18530 3220
rect 18500 3170 18530 3200
rect 18500 3150 18505 3170
rect 18525 3150 18530 3170
rect 18500 3120 18530 3150
rect 18500 3100 18505 3120
rect 18525 3100 18530 3120
rect 18500 3070 18530 3100
rect 18500 3050 18505 3070
rect 18525 3050 18530 3070
rect 18500 3020 18530 3050
rect 18500 3000 18505 3020
rect 18525 3000 18530 3020
rect 18500 2990 18530 3000
rect 18555 3570 18585 3580
rect 18555 3550 18560 3570
rect 18580 3550 18585 3570
rect 18555 3520 18585 3550
rect 18555 3500 18560 3520
rect 18580 3500 18585 3520
rect 18555 3470 18585 3500
rect 18555 3450 18560 3470
rect 18580 3450 18585 3470
rect 18555 3420 18585 3450
rect 18555 3400 18560 3420
rect 18580 3400 18585 3420
rect 18555 3370 18585 3400
rect 18555 3350 18560 3370
rect 18580 3350 18585 3370
rect 18555 3320 18585 3350
rect 18555 3300 18560 3320
rect 18580 3300 18585 3320
rect 18555 3270 18585 3300
rect 18555 3250 18560 3270
rect 18580 3250 18585 3270
rect 18555 3220 18585 3250
rect 18555 3200 18560 3220
rect 18580 3200 18585 3220
rect 18555 3170 18585 3200
rect 18555 3150 18560 3170
rect 18580 3150 18585 3170
rect 18555 3120 18585 3150
rect 18555 3100 18560 3120
rect 18580 3100 18585 3120
rect 18555 3070 18585 3100
rect 18555 3050 18560 3070
rect 18580 3050 18585 3070
rect 18555 3020 18585 3050
rect 18555 3000 18560 3020
rect 18580 3000 18585 3020
rect 18555 2990 18585 3000
rect 18610 3570 18680 3580
rect 18610 3550 18615 3570
rect 18635 3550 18655 3570
rect 18675 3550 18680 3570
rect 18610 3520 18680 3550
rect 18610 3500 18615 3520
rect 18635 3500 18655 3520
rect 18675 3500 18680 3520
rect 18610 3470 18680 3500
rect 18610 3450 18615 3470
rect 18635 3450 18655 3470
rect 18675 3450 18680 3470
rect 18610 3420 18680 3450
rect 18610 3400 18615 3420
rect 18635 3400 18655 3420
rect 18675 3400 18680 3420
rect 18610 3370 18680 3400
rect 18610 3350 18615 3370
rect 18635 3350 18655 3370
rect 18675 3350 18680 3370
rect 18610 3320 18680 3350
rect 18610 3300 18615 3320
rect 18635 3300 18655 3320
rect 18675 3300 18680 3320
rect 18755 3520 18896 3560
rect 18610 3270 18680 3300
rect 18610 3250 18615 3270
rect 18635 3250 18655 3270
rect 18675 3250 18680 3270
rect 18610 3220 18680 3250
rect 18610 3200 18615 3220
rect 18635 3200 18655 3220
rect 18675 3200 18680 3220
rect 18610 3170 18680 3200
rect 18610 3150 18615 3170
rect 18635 3150 18655 3170
rect 18675 3150 18680 3170
rect 18610 3120 18680 3150
rect 18610 3100 18615 3120
rect 18635 3100 18655 3120
rect 18675 3100 18680 3120
rect 18610 3070 18680 3100
rect 18610 3050 18615 3070
rect 18635 3050 18655 3070
rect 18675 3050 18680 3070
rect 18610 3020 18680 3050
rect 18610 3000 18615 3020
rect 18635 3000 18655 3020
rect 18675 3000 18680 3020
rect 18610 2990 18680 3000
rect 15125 2970 15145 2990
rect 15275 2970 15295 2990
rect 15385 2970 15405 2990
rect 15495 2970 15515 2990
rect 15605 2970 15625 2990
rect 15715 2970 15735 2990
rect 15865 2970 15885 2990
rect 17915 2970 17935 2990
rect 18065 2970 18085 2990
rect 18175 2970 18195 2990
rect 18285 2970 18305 2990
rect 18395 2970 18415 2990
rect 18505 2970 18525 2990
rect 18655 2970 18675 2990
rect 2960 2915 3030 2925
rect 1266 2865 1306 2900
rect 2330 2895 2375 2905
rect 2330 2870 2340 2895
rect 2365 2870 2375 2895
rect 2330 2860 2375 2870
rect 2960 2895 2965 2915
rect 2985 2895 3005 2915
rect 3025 2895 3030 2915
rect 2960 2865 3030 2895
rect -55 2825 -25 2855
rect 51 2850 96 2855
rect 51 2825 61 2850
rect 86 2825 96 2850
rect 51 2820 96 2825
rect 724 2850 769 2855
rect 724 2825 734 2850
rect 759 2825 769 2850
rect 724 2820 769 2825
rect 1210 2820 1240 2850
rect 2960 2845 2965 2865
rect 2985 2845 3005 2865
rect 3025 2845 3030 2865
rect 1261 2835 1306 2840
rect 1261 2810 1271 2835
rect 1296 2810 1306 2835
rect 1261 2805 1306 2810
rect 1960 2835 2005 2840
rect 1960 2810 1970 2835
rect 1995 2810 2005 2835
rect 1960 2805 2005 2810
rect 2330 2800 2370 2840
rect 2960 2835 3030 2845
rect 3090 2915 3120 2925
rect 3090 2895 3095 2915
rect 3115 2895 3120 2915
rect 3090 2865 3120 2895
rect 3090 2845 3095 2865
rect 3115 2845 3120 2865
rect 3090 2835 3120 2845
rect 3180 2915 3210 2925
rect 3180 2895 3185 2915
rect 3205 2895 3210 2915
rect 3180 2865 3210 2895
rect 3180 2845 3185 2865
rect 3205 2845 3210 2865
rect 3180 2835 3210 2845
rect 3270 2915 3300 2925
rect 3270 2895 3275 2915
rect 3295 2895 3300 2915
rect 3270 2865 3300 2895
rect 3270 2845 3275 2865
rect 3295 2845 3300 2865
rect 3270 2835 3300 2845
rect 3360 2915 3390 2925
rect 3360 2895 3365 2915
rect 3385 2895 3390 2915
rect 3360 2865 3390 2895
rect 3360 2845 3365 2865
rect 3385 2845 3390 2865
rect 3360 2835 3390 2845
rect 3450 2915 3480 2925
rect 3450 2895 3455 2915
rect 3475 2895 3480 2915
rect 3450 2865 3480 2895
rect 3450 2845 3455 2865
rect 3475 2845 3480 2865
rect 3450 2835 3480 2845
rect 3540 2915 3570 2925
rect 3540 2895 3545 2915
rect 3565 2895 3570 2915
rect 3540 2865 3570 2895
rect 3540 2845 3545 2865
rect 3565 2845 3570 2865
rect 3540 2835 3570 2845
rect 3630 2915 3660 2925
rect 3630 2895 3635 2915
rect 3655 2895 3660 2915
rect 3630 2865 3660 2895
rect 3630 2845 3635 2865
rect 3655 2845 3660 2865
rect 3630 2835 3660 2845
rect 3720 2915 3750 2925
rect 3720 2895 3725 2915
rect 3745 2895 3750 2915
rect 3720 2865 3750 2895
rect 3720 2845 3725 2865
rect 3745 2845 3750 2865
rect 3720 2835 3750 2845
rect 3810 2915 3840 2925
rect 3810 2895 3815 2915
rect 3835 2895 3840 2915
rect 3810 2865 3840 2895
rect 3810 2845 3815 2865
rect 3835 2845 3840 2865
rect 3810 2835 3840 2845
rect 3900 2915 3930 2925
rect 3900 2895 3905 2915
rect 3925 2895 3930 2915
rect 3900 2865 3930 2895
rect 3900 2845 3905 2865
rect 3925 2845 3930 2865
rect 3900 2835 3930 2845
rect 3990 2915 4020 2925
rect 3990 2895 3995 2915
rect 4015 2895 4020 2915
rect 3990 2865 4020 2895
rect 3990 2845 3995 2865
rect 4015 2845 4020 2865
rect 3990 2835 4020 2845
rect 4080 2915 4110 2925
rect 4080 2895 4085 2915
rect 4105 2895 4110 2915
rect 4080 2865 4110 2895
rect 4080 2845 4085 2865
rect 4105 2845 4110 2865
rect 4080 2835 4110 2845
rect 4170 2915 4200 2925
rect 4170 2895 4175 2915
rect 4195 2895 4200 2915
rect 4170 2865 4200 2895
rect 4170 2845 4175 2865
rect 4195 2845 4200 2865
rect 4170 2835 4200 2845
rect 4260 2915 4290 2925
rect 4260 2895 4265 2915
rect 4285 2895 4290 2915
rect 4260 2865 4290 2895
rect 4260 2845 4265 2865
rect 4285 2845 4290 2865
rect 4260 2835 4290 2845
rect 4350 2915 4380 2925
rect 4350 2895 4355 2915
rect 4375 2895 4380 2915
rect 4350 2865 4380 2895
rect 4350 2845 4355 2865
rect 4375 2845 4380 2865
rect 4350 2835 4380 2845
rect 4440 2915 4470 2925
rect 4440 2895 4445 2915
rect 4465 2895 4470 2915
rect 4440 2865 4470 2895
rect 4440 2845 4445 2865
rect 4465 2845 4470 2865
rect 4440 2835 4470 2845
rect 4530 2915 4560 2925
rect 4530 2895 4535 2915
rect 4555 2895 4560 2915
rect 4530 2865 4560 2895
rect 4530 2845 4535 2865
rect 4555 2845 4560 2865
rect 4530 2835 4560 2845
rect 4620 2915 4650 2925
rect 4620 2895 4625 2915
rect 4645 2895 4650 2915
rect 4620 2865 4650 2895
rect 4620 2845 4625 2865
rect 4645 2845 4650 2865
rect 4620 2835 4650 2845
rect 4710 2915 4740 2925
rect 4710 2895 4715 2915
rect 4735 2895 4740 2915
rect 4710 2865 4740 2895
rect 4710 2845 4715 2865
rect 4735 2845 4740 2865
rect 4710 2835 4740 2845
rect 4800 2915 4830 2925
rect 4800 2895 4805 2915
rect 4825 2895 4830 2915
rect 4800 2865 4830 2895
rect 4800 2845 4805 2865
rect 4825 2845 4830 2865
rect 4800 2835 4830 2845
rect 4890 2915 4920 2925
rect 4890 2895 4895 2915
rect 4915 2895 4920 2915
rect 4890 2865 4920 2895
rect 4890 2845 4895 2865
rect 4915 2845 4920 2865
rect 4890 2835 4920 2845
rect 4980 2915 5050 2925
rect 4980 2895 4985 2915
rect 5005 2895 5025 2915
rect 5045 2895 5050 2915
rect 14904 2900 15045 2940
rect 15115 2960 15155 2970
rect 15115 2940 15125 2960
rect 15145 2940 15155 2960
rect 15115 2930 15155 2940
rect 15265 2960 15305 2970
rect 15265 2940 15275 2960
rect 15295 2940 15305 2960
rect 15265 2930 15305 2940
rect 15375 2960 15415 2970
rect 15375 2940 15385 2960
rect 15405 2940 15415 2960
rect 15375 2930 15415 2940
rect 15485 2960 15525 2970
rect 15485 2940 15495 2960
rect 15515 2940 15525 2960
rect 15485 2930 15525 2940
rect 15595 2960 15635 2970
rect 15595 2940 15605 2960
rect 15625 2940 15635 2960
rect 15595 2930 15635 2940
rect 15653 2960 15687 2970
rect 15653 2940 15661 2960
rect 15679 2940 15687 2960
rect 15653 2930 15687 2940
rect 15705 2960 15745 2970
rect 15705 2940 15715 2960
rect 15735 2940 15745 2960
rect 15705 2930 15745 2940
rect 15855 2960 15895 2970
rect 15855 2940 15865 2960
rect 15885 2940 15895 2960
rect 17905 2960 17945 2970
rect 15855 2930 15895 2940
rect 16180 2940 16220 2950
rect 16180 2920 16190 2940
rect 16210 2920 16220 2940
rect 16180 2910 16220 2920
rect 16340 2940 16380 2950
rect 16340 2920 16350 2940
rect 16370 2920 16380 2940
rect 16340 2910 16380 2920
rect 16460 2940 16500 2950
rect 16460 2920 16470 2940
rect 16490 2920 16500 2940
rect 16460 2910 16500 2920
rect 16580 2940 16620 2950
rect 16580 2920 16590 2940
rect 16610 2920 16620 2940
rect 16580 2910 16620 2920
rect 16700 2940 16740 2950
rect 16700 2920 16710 2940
rect 16730 2920 16740 2940
rect 16700 2910 16740 2920
rect 16820 2940 16860 2950
rect 16820 2920 16830 2940
rect 16850 2920 16860 2940
rect 16820 2910 16860 2920
rect 16940 2940 16980 2950
rect 16940 2920 16950 2940
rect 16970 2920 16980 2940
rect 16940 2910 16980 2920
rect 17060 2940 17100 2950
rect 17060 2920 17070 2940
rect 17090 2920 17100 2940
rect 17060 2910 17100 2920
rect 17180 2940 17220 2950
rect 17180 2920 17190 2940
rect 17210 2920 17220 2940
rect 17180 2910 17220 2920
rect 17300 2940 17340 2950
rect 17300 2920 17310 2940
rect 17330 2920 17340 2940
rect 17300 2910 17340 2920
rect 17420 2940 17460 2950
rect 17420 2920 17430 2940
rect 17450 2920 17460 2940
rect 17420 2910 17460 2920
rect 17480 2910 17520 2950
rect 17580 2940 17620 2950
rect 17580 2920 17590 2940
rect 17610 2920 17620 2940
rect 17905 2940 17915 2960
rect 17935 2940 17945 2960
rect 17905 2930 17945 2940
rect 18055 2960 18095 2970
rect 18055 2940 18065 2960
rect 18085 2940 18095 2960
rect 18055 2930 18095 2940
rect 18113 2960 18147 2970
rect 18113 2940 18121 2960
rect 18139 2940 18147 2960
rect 18113 2930 18147 2940
rect 18165 2960 18205 2970
rect 18165 2940 18175 2960
rect 18195 2940 18205 2960
rect 18165 2930 18205 2940
rect 18275 2960 18315 2970
rect 18275 2940 18285 2960
rect 18305 2940 18315 2960
rect 18275 2930 18315 2940
rect 18385 2960 18425 2970
rect 18385 2940 18395 2960
rect 18415 2940 18425 2960
rect 18385 2930 18425 2940
rect 18495 2960 18535 2970
rect 18495 2940 18505 2960
rect 18525 2940 18535 2960
rect 18495 2930 18535 2940
rect 18645 2960 18685 2970
rect 18645 2940 18655 2960
rect 18675 2940 18685 2960
rect 18645 2930 18685 2940
rect 17580 2910 17620 2920
rect 4980 2865 5050 2895
rect 16190 2890 16210 2910
rect 16350 2890 16370 2910
rect 16470 2890 16490 2910
rect 16590 2890 16610 2910
rect 16710 2890 16730 2910
rect 16830 2890 16850 2910
rect 16950 2890 16970 2910
rect 17070 2890 17090 2910
rect 17190 2890 17210 2910
rect 17310 2890 17330 2910
rect 17430 2890 17450 2910
rect 17590 2890 17610 2910
rect 18755 2900 18896 2940
rect 4980 2845 4985 2865
rect 5005 2845 5025 2865
rect 5045 2845 5050 2865
rect 4980 2835 5050 2845
rect 16185 2880 16255 2890
rect 16185 2860 16190 2880
rect 16210 2860 16230 2880
rect 16250 2860 16255 2880
rect 3005 2815 3025 2835
rect 3185 2815 3205 2835
rect 3365 2815 3385 2835
rect 3545 2815 3565 2835
rect 3725 2815 3745 2835
rect 3905 2815 3925 2835
rect 4085 2815 4105 2835
rect 4265 2815 4285 2835
rect 4445 2815 4465 2835
rect 4625 2815 4645 2835
rect 4805 2815 4825 2835
rect 4985 2815 5005 2835
rect 16185 2830 16255 2860
rect 2995 2805 3035 2815
rect -10 2765 20 2795
rect 51 2790 96 2795
rect 51 2765 61 2790
rect 86 2765 96 2790
rect 51 2760 96 2765
rect 724 2790 769 2795
rect 724 2765 734 2790
rect 759 2765 769 2790
rect 724 2760 769 2765
rect 2620 2755 2660 2795
rect 2995 2785 3005 2805
rect 3025 2785 3035 2805
rect 2995 2775 3035 2785
rect 3175 2805 3215 2815
rect 3175 2785 3185 2805
rect 3205 2785 3215 2805
rect 3175 2775 3215 2785
rect 3355 2805 3395 2815
rect 3355 2785 3365 2805
rect 3385 2785 3395 2805
rect 3355 2775 3395 2785
rect 3535 2805 3575 2815
rect 3535 2785 3545 2805
rect 3565 2785 3575 2805
rect 3535 2775 3575 2785
rect 3715 2805 3755 2815
rect 3715 2785 3725 2805
rect 3745 2785 3755 2805
rect 3715 2775 3755 2785
rect 3895 2805 3935 2815
rect 3895 2785 3905 2805
rect 3925 2785 3935 2805
rect 3895 2775 3935 2785
rect 4075 2805 4115 2815
rect 4075 2785 4085 2805
rect 4105 2785 4115 2805
rect 4075 2775 4115 2785
rect 4255 2805 4295 2815
rect 4255 2785 4265 2805
rect 4285 2785 4295 2805
rect 4255 2775 4295 2785
rect 4435 2805 4475 2815
rect 4435 2785 4445 2805
rect 4465 2785 4475 2805
rect 4435 2775 4475 2785
rect 4615 2805 4655 2815
rect 4615 2785 4625 2805
rect 4645 2785 4655 2805
rect 4615 2775 4655 2785
rect 4795 2805 4835 2815
rect 4795 2785 4805 2805
rect 4825 2785 4835 2805
rect 4795 2775 4835 2785
rect 4975 2805 5015 2815
rect 4975 2785 4985 2805
rect 5005 2785 5015 2805
rect 4975 2775 5015 2785
rect 16185 2810 16190 2830
rect 16210 2810 16230 2830
rect 16250 2810 16255 2830
rect 16185 2780 16255 2810
rect 16185 2760 16190 2780
rect 16210 2760 16230 2780
rect 16250 2760 16255 2780
rect 1266 2715 1296 2745
rect 2150 2710 2190 2750
rect 3175 2745 3215 2755
rect 3175 2725 3185 2745
rect 3205 2725 3215 2745
rect 3175 2715 3215 2725
rect 3355 2745 3395 2755
rect 3355 2725 3365 2745
rect 3385 2725 3395 2745
rect 3355 2715 3395 2725
rect 3535 2745 3575 2755
rect 3535 2725 3545 2745
rect 3565 2725 3575 2745
rect 3535 2715 3575 2725
rect 3715 2745 3755 2755
rect 3715 2725 3725 2745
rect 3745 2725 3755 2745
rect 3715 2715 3755 2725
rect 3895 2745 3935 2755
rect 3895 2725 3905 2745
rect 3925 2725 3935 2745
rect 3895 2715 3935 2725
rect 4075 2745 4115 2755
rect 4075 2725 4085 2745
rect 4105 2725 4115 2745
rect 4075 2715 4115 2725
rect 4255 2745 4295 2755
rect 4255 2725 4265 2745
rect 4285 2725 4295 2745
rect 4255 2715 4295 2725
rect 4435 2745 4475 2755
rect 4435 2725 4445 2745
rect 4465 2725 4475 2745
rect 4435 2715 4475 2725
rect 4615 2745 4655 2755
rect 4615 2725 4625 2745
rect 4645 2725 4655 2745
rect 4615 2715 4655 2725
rect 4795 2745 4835 2755
rect 4795 2725 4805 2745
rect 4825 2725 4835 2745
rect 4795 2715 4835 2725
rect 16185 2730 16255 2760
rect 650 2055 775 2700
rect 1330 2055 1455 2700
rect 2010 2055 2135 2700
rect 3185 2695 3205 2715
rect 3365 2695 3385 2715
rect 3545 2695 3565 2715
rect 3725 2695 3745 2715
rect 3905 2695 3925 2715
rect 4085 2695 4105 2715
rect 4265 2695 4285 2715
rect 4445 2695 4465 2715
rect 4625 2695 4645 2715
rect 4805 2695 4825 2715
rect 16185 2710 16190 2730
rect 16210 2710 16230 2730
rect 16250 2710 16255 2730
rect 15210 2700 15250 2710
rect 3140 2685 3210 2695
rect 3140 2665 3145 2685
rect 3165 2665 3185 2685
rect 3205 2665 3210 2685
rect 3140 2635 3210 2665
rect 3140 2615 3145 2635
rect 3165 2615 3185 2635
rect 3205 2615 3210 2635
rect 3140 2585 3210 2615
rect 3140 2565 3145 2585
rect 3165 2565 3185 2585
rect 3205 2565 3210 2585
rect 3140 2535 3210 2565
rect 3140 2515 3145 2535
rect 3165 2515 3185 2535
rect 3205 2515 3210 2535
rect 3140 2485 3210 2515
rect 3140 2465 3145 2485
rect 3165 2465 3185 2485
rect 3205 2465 3210 2485
rect 3140 2435 3210 2465
rect 3140 2415 3145 2435
rect 3165 2415 3185 2435
rect 3205 2415 3210 2435
rect 3140 2405 3210 2415
rect 3270 2685 3300 2695
rect 3270 2665 3275 2685
rect 3295 2665 3300 2685
rect 3270 2635 3300 2665
rect 3270 2615 3275 2635
rect 3295 2615 3300 2635
rect 3270 2585 3300 2615
rect 3270 2565 3275 2585
rect 3295 2565 3300 2585
rect 3270 2535 3300 2565
rect 3270 2515 3275 2535
rect 3295 2515 3300 2535
rect 3270 2485 3300 2515
rect 3270 2465 3275 2485
rect 3295 2465 3300 2485
rect 3270 2435 3300 2465
rect 3270 2415 3275 2435
rect 3295 2415 3300 2435
rect 3270 2405 3300 2415
rect 3360 2685 3390 2695
rect 3360 2665 3365 2685
rect 3385 2665 3390 2685
rect 3360 2635 3390 2665
rect 3360 2615 3365 2635
rect 3385 2615 3390 2635
rect 3360 2585 3390 2615
rect 3360 2565 3365 2585
rect 3385 2565 3390 2585
rect 3360 2535 3390 2565
rect 3360 2515 3365 2535
rect 3385 2515 3390 2535
rect 3360 2485 3390 2515
rect 3360 2465 3365 2485
rect 3385 2465 3390 2485
rect 3360 2435 3390 2465
rect 3360 2415 3365 2435
rect 3385 2415 3390 2435
rect 3360 2405 3390 2415
rect 3450 2685 3480 2695
rect 3450 2665 3455 2685
rect 3475 2665 3480 2685
rect 3450 2635 3480 2665
rect 3450 2615 3455 2635
rect 3475 2615 3480 2635
rect 3450 2585 3480 2615
rect 3450 2565 3455 2585
rect 3475 2565 3480 2585
rect 3450 2535 3480 2565
rect 3450 2515 3455 2535
rect 3475 2515 3480 2535
rect 3450 2485 3480 2515
rect 3450 2465 3455 2485
rect 3475 2465 3480 2485
rect 3450 2435 3480 2465
rect 3450 2415 3455 2435
rect 3475 2415 3480 2435
rect 3450 2405 3480 2415
rect 3540 2685 3570 2695
rect 3540 2665 3545 2685
rect 3565 2665 3570 2685
rect 3540 2635 3570 2665
rect 3540 2615 3545 2635
rect 3565 2615 3570 2635
rect 3540 2585 3570 2615
rect 3540 2565 3545 2585
rect 3565 2565 3570 2585
rect 3540 2535 3570 2565
rect 3540 2515 3545 2535
rect 3565 2515 3570 2535
rect 3540 2485 3570 2515
rect 3540 2465 3545 2485
rect 3565 2465 3570 2485
rect 3540 2435 3570 2465
rect 3540 2415 3545 2435
rect 3565 2415 3570 2435
rect 3540 2405 3570 2415
rect 3630 2685 3660 2695
rect 3630 2665 3635 2685
rect 3655 2665 3660 2685
rect 3630 2635 3660 2665
rect 3630 2615 3635 2635
rect 3655 2615 3660 2635
rect 3630 2585 3660 2615
rect 3630 2565 3635 2585
rect 3655 2565 3660 2585
rect 3630 2535 3660 2565
rect 3630 2515 3635 2535
rect 3655 2515 3660 2535
rect 3630 2485 3660 2515
rect 3630 2465 3635 2485
rect 3655 2465 3660 2485
rect 3630 2435 3660 2465
rect 3630 2415 3635 2435
rect 3655 2415 3660 2435
rect 3630 2405 3660 2415
rect 3720 2685 3750 2695
rect 3720 2665 3725 2685
rect 3745 2665 3750 2685
rect 3720 2635 3750 2665
rect 3720 2615 3725 2635
rect 3745 2615 3750 2635
rect 3720 2585 3750 2615
rect 3720 2565 3725 2585
rect 3745 2565 3750 2585
rect 3720 2535 3750 2565
rect 3720 2515 3725 2535
rect 3745 2515 3750 2535
rect 3720 2485 3750 2515
rect 3720 2465 3725 2485
rect 3745 2465 3750 2485
rect 3720 2435 3750 2465
rect 3720 2415 3725 2435
rect 3745 2415 3750 2435
rect 3720 2405 3750 2415
rect 3810 2685 3840 2695
rect 3810 2665 3815 2685
rect 3835 2665 3840 2685
rect 3810 2635 3840 2665
rect 3810 2615 3815 2635
rect 3835 2615 3840 2635
rect 3810 2585 3840 2615
rect 3810 2565 3815 2585
rect 3835 2565 3840 2585
rect 3810 2535 3840 2565
rect 3810 2515 3815 2535
rect 3835 2515 3840 2535
rect 3810 2485 3840 2515
rect 3810 2465 3815 2485
rect 3835 2465 3840 2485
rect 3810 2435 3840 2465
rect 3810 2415 3815 2435
rect 3835 2415 3840 2435
rect 3810 2405 3840 2415
rect 3900 2685 3930 2695
rect 3900 2665 3905 2685
rect 3925 2665 3930 2685
rect 3900 2635 3930 2665
rect 3900 2615 3905 2635
rect 3925 2615 3930 2635
rect 3900 2585 3930 2615
rect 3900 2565 3905 2585
rect 3925 2565 3930 2585
rect 3900 2535 3930 2565
rect 3900 2515 3905 2535
rect 3925 2515 3930 2535
rect 3900 2485 3930 2515
rect 3900 2465 3905 2485
rect 3925 2465 3930 2485
rect 3900 2435 3930 2465
rect 3900 2415 3905 2435
rect 3925 2415 3930 2435
rect 3900 2405 3930 2415
rect 3990 2685 4020 2695
rect 3990 2665 3995 2685
rect 4015 2665 4020 2685
rect 3990 2635 4020 2665
rect 3990 2615 3995 2635
rect 4015 2615 4020 2635
rect 3990 2585 4020 2615
rect 3990 2565 3995 2585
rect 4015 2565 4020 2585
rect 3990 2535 4020 2565
rect 3990 2515 3995 2535
rect 4015 2515 4020 2535
rect 3990 2485 4020 2515
rect 3990 2465 3995 2485
rect 4015 2465 4020 2485
rect 3990 2435 4020 2465
rect 3990 2415 3995 2435
rect 4015 2415 4020 2435
rect 3990 2405 4020 2415
rect 4080 2685 4110 2695
rect 4080 2665 4085 2685
rect 4105 2665 4110 2685
rect 4080 2635 4110 2665
rect 4080 2615 4085 2635
rect 4105 2615 4110 2635
rect 4080 2585 4110 2615
rect 4080 2565 4085 2585
rect 4105 2565 4110 2585
rect 4080 2535 4110 2565
rect 4080 2515 4085 2535
rect 4105 2515 4110 2535
rect 4080 2485 4110 2515
rect 4080 2465 4085 2485
rect 4105 2465 4110 2485
rect 4080 2435 4110 2465
rect 4080 2415 4085 2435
rect 4105 2415 4110 2435
rect 4080 2405 4110 2415
rect 4170 2685 4200 2695
rect 4170 2665 4175 2685
rect 4195 2665 4200 2685
rect 4170 2635 4200 2665
rect 4170 2615 4175 2635
rect 4195 2615 4200 2635
rect 4170 2585 4200 2615
rect 4170 2565 4175 2585
rect 4195 2565 4200 2585
rect 4170 2535 4200 2565
rect 4170 2515 4175 2535
rect 4195 2515 4200 2535
rect 4170 2485 4200 2515
rect 4170 2465 4175 2485
rect 4195 2465 4200 2485
rect 4170 2435 4200 2465
rect 4170 2415 4175 2435
rect 4195 2415 4200 2435
rect 4170 2405 4200 2415
rect 4260 2685 4290 2695
rect 4260 2665 4265 2685
rect 4285 2665 4290 2685
rect 4260 2635 4290 2665
rect 4260 2615 4265 2635
rect 4285 2615 4290 2635
rect 4260 2585 4290 2615
rect 4260 2565 4265 2585
rect 4285 2565 4290 2585
rect 4260 2535 4290 2565
rect 4260 2515 4265 2535
rect 4285 2515 4290 2535
rect 4260 2485 4290 2515
rect 4260 2465 4265 2485
rect 4285 2465 4290 2485
rect 4260 2435 4290 2465
rect 4260 2415 4265 2435
rect 4285 2415 4290 2435
rect 4260 2405 4290 2415
rect 4350 2685 4380 2695
rect 4350 2665 4355 2685
rect 4375 2665 4380 2685
rect 4350 2635 4380 2665
rect 4350 2615 4355 2635
rect 4375 2615 4380 2635
rect 4350 2585 4380 2615
rect 4350 2565 4355 2585
rect 4375 2565 4380 2585
rect 4350 2535 4380 2565
rect 4350 2515 4355 2535
rect 4375 2515 4380 2535
rect 4350 2485 4380 2515
rect 4350 2465 4355 2485
rect 4375 2465 4380 2485
rect 4350 2435 4380 2465
rect 4350 2415 4355 2435
rect 4375 2415 4380 2435
rect 4350 2405 4380 2415
rect 4440 2685 4470 2695
rect 4440 2665 4445 2685
rect 4465 2665 4470 2685
rect 4440 2635 4470 2665
rect 4440 2615 4445 2635
rect 4465 2615 4470 2635
rect 4440 2585 4470 2615
rect 4440 2565 4445 2585
rect 4465 2565 4470 2585
rect 4440 2535 4470 2565
rect 4440 2515 4445 2535
rect 4465 2515 4470 2535
rect 4440 2485 4470 2515
rect 4440 2465 4445 2485
rect 4465 2465 4470 2485
rect 4440 2435 4470 2465
rect 4440 2415 4445 2435
rect 4465 2415 4470 2435
rect 4440 2405 4470 2415
rect 4530 2685 4560 2695
rect 4530 2665 4535 2685
rect 4555 2665 4560 2685
rect 4530 2635 4560 2665
rect 4530 2615 4535 2635
rect 4555 2615 4560 2635
rect 4530 2585 4560 2615
rect 4530 2565 4535 2585
rect 4555 2565 4560 2585
rect 4530 2535 4560 2565
rect 4530 2515 4535 2535
rect 4555 2515 4560 2535
rect 4530 2485 4560 2515
rect 4530 2465 4535 2485
rect 4555 2465 4560 2485
rect 4530 2435 4560 2465
rect 4530 2415 4535 2435
rect 4555 2415 4560 2435
rect 4530 2405 4560 2415
rect 4620 2685 4650 2695
rect 4620 2665 4625 2685
rect 4645 2665 4650 2685
rect 4620 2635 4650 2665
rect 4620 2615 4625 2635
rect 4645 2615 4650 2635
rect 4620 2585 4650 2615
rect 4620 2565 4625 2585
rect 4645 2565 4650 2585
rect 4620 2535 4650 2565
rect 4620 2515 4625 2535
rect 4645 2515 4650 2535
rect 4620 2485 4650 2515
rect 4620 2465 4625 2485
rect 4645 2465 4650 2485
rect 4620 2435 4650 2465
rect 4620 2415 4625 2435
rect 4645 2415 4650 2435
rect 4620 2405 4650 2415
rect 4710 2685 4740 2695
rect 4710 2665 4715 2685
rect 4735 2665 4740 2685
rect 4710 2635 4740 2665
rect 4710 2615 4715 2635
rect 4735 2615 4740 2635
rect 4710 2585 4740 2615
rect 4710 2565 4715 2585
rect 4735 2565 4740 2585
rect 4710 2535 4740 2565
rect 4710 2515 4715 2535
rect 4735 2515 4740 2535
rect 4710 2485 4740 2515
rect 4710 2465 4715 2485
rect 4735 2465 4740 2485
rect 4710 2435 4740 2465
rect 4710 2415 4715 2435
rect 4735 2415 4740 2435
rect 4710 2405 4740 2415
rect 4800 2685 4870 2695
rect 4800 2665 4805 2685
rect 4825 2665 4845 2685
rect 4865 2665 4870 2685
rect 15210 2680 15220 2700
rect 15240 2680 15250 2700
rect 15210 2670 15250 2680
rect 15320 2700 15360 2710
rect 15320 2680 15330 2700
rect 15350 2680 15360 2700
rect 15320 2670 15360 2680
rect 15430 2700 15470 2710
rect 15430 2680 15440 2700
rect 15460 2680 15470 2700
rect 15430 2670 15470 2680
rect 15540 2700 15580 2710
rect 15540 2680 15550 2700
rect 15570 2680 15580 2700
rect 15540 2670 15580 2680
rect 15650 2700 15690 2710
rect 15650 2680 15660 2700
rect 15680 2680 15690 2700
rect 15650 2670 15690 2680
rect 15760 2700 15800 2710
rect 15760 2680 15770 2700
rect 15790 2680 15800 2700
rect 15760 2670 15800 2680
rect 16185 2680 16255 2710
rect 4800 2635 4870 2665
rect 4800 2615 4805 2635
rect 4825 2615 4845 2635
rect 4865 2615 4870 2635
rect 4800 2585 4870 2615
rect 4800 2565 4805 2585
rect 4825 2565 4845 2585
rect 4865 2565 4870 2585
rect 4800 2535 4870 2565
rect 4800 2515 4805 2535
rect 4825 2515 4845 2535
rect 4865 2515 4870 2535
rect 4800 2485 4870 2515
rect 4800 2465 4805 2485
rect 4825 2465 4845 2485
rect 4865 2465 4870 2485
rect 4800 2435 4870 2465
rect 4800 2415 4805 2435
rect 4825 2415 4845 2435
rect 4865 2415 4870 2435
rect 4800 2405 4870 2415
rect 14790 2645 15005 2665
rect 15220 2650 15240 2670
rect 15330 2650 15350 2670
rect 15440 2650 15460 2670
rect 15550 2650 15570 2670
rect 15660 2650 15680 2670
rect 15770 2650 15790 2670
rect 16185 2660 16190 2680
rect 16210 2660 16230 2680
rect 16250 2660 16255 2680
rect 14790 2625 14825 2645
rect 14970 2625 15005 2645
rect 14885 2575 14910 2625
rect 15120 2640 15190 2650
rect 15120 2620 15125 2640
rect 15145 2620 15165 2640
rect 15185 2620 15190 2640
rect 15120 2590 15190 2620
rect 15120 2570 15125 2590
rect 15145 2570 15165 2590
rect 15185 2570 15190 2590
rect 15120 2540 15190 2570
rect 15120 2520 15125 2540
rect 15145 2520 15165 2540
rect 15185 2520 15190 2540
rect 15120 2490 15190 2520
rect 15120 2470 15125 2490
rect 15145 2470 15165 2490
rect 15185 2470 15190 2490
rect 15120 2460 15190 2470
rect 15215 2640 15245 2650
rect 15215 2620 15220 2640
rect 15240 2620 15245 2640
rect 15215 2590 15245 2620
rect 15215 2570 15220 2590
rect 15240 2570 15245 2590
rect 15215 2540 15245 2570
rect 15215 2520 15220 2540
rect 15240 2520 15245 2540
rect 15215 2490 15245 2520
rect 15215 2470 15220 2490
rect 15240 2470 15245 2490
rect 15215 2460 15245 2470
rect 15270 2640 15300 2650
rect 15270 2620 15275 2640
rect 15295 2620 15300 2640
rect 15270 2590 15300 2620
rect 15270 2570 15275 2590
rect 15295 2570 15300 2590
rect 15270 2540 15300 2570
rect 15270 2520 15275 2540
rect 15295 2520 15300 2540
rect 15270 2490 15300 2520
rect 15270 2470 15275 2490
rect 15295 2470 15300 2490
rect 15270 2460 15300 2470
rect 15325 2640 15355 2650
rect 15325 2620 15330 2640
rect 15350 2620 15355 2640
rect 15325 2590 15355 2620
rect 15325 2570 15330 2590
rect 15350 2570 15355 2590
rect 15325 2540 15355 2570
rect 15325 2520 15330 2540
rect 15350 2520 15355 2540
rect 15325 2490 15355 2520
rect 15325 2470 15330 2490
rect 15350 2470 15355 2490
rect 15325 2460 15355 2470
rect 15380 2640 15410 2650
rect 15380 2620 15385 2640
rect 15405 2620 15410 2640
rect 15380 2590 15410 2620
rect 15380 2570 15385 2590
rect 15405 2570 15410 2590
rect 15380 2540 15410 2570
rect 15380 2520 15385 2540
rect 15405 2520 15410 2540
rect 15380 2490 15410 2520
rect 15380 2470 15385 2490
rect 15405 2470 15410 2490
rect 15380 2460 15410 2470
rect 15435 2640 15465 2650
rect 15435 2620 15440 2640
rect 15460 2620 15465 2640
rect 15435 2590 15465 2620
rect 15435 2570 15440 2590
rect 15460 2570 15465 2590
rect 15435 2540 15465 2570
rect 15435 2520 15440 2540
rect 15460 2520 15465 2540
rect 15435 2490 15465 2520
rect 15435 2470 15440 2490
rect 15460 2470 15465 2490
rect 15435 2460 15465 2470
rect 15490 2640 15520 2650
rect 15490 2620 15495 2640
rect 15515 2620 15520 2640
rect 15490 2590 15520 2620
rect 15490 2570 15495 2590
rect 15515 2570 15520 2590
rect 15490 2540 15520 2570
rect 15490 2520 15495 2540
rect 15515 2520 15520 2540
rect 15490 2490 15520 2520
rect 15490 2470 15495 2490
rect 15515 2470 15520 2490
rect 15490 2460 15520 2470
rect 15545 2640 15575 2650
rect 15545 2620 15550 2640
rect 15570 2620 15575 2640
rect 15545 2590 15575 2620
rect 15545 2570 15550 2590
rect 15570 2570 15575 2590
rect 15545 2540 15575 2570
rect 15545 2520 15550 2540
rect 15570 2520 15575 2540
rect 15545 2490 15575 2520
rect 15545 2470 15550 2490
rect 15570 2470 15575 2490
rect 15545 2460 15575 2470
rect 15600 2640 15630 2650
rect 15600 2620 15605 2640
rect 15625 2620 15630 2640
rect 15600 2590 15630 2620
rect 15600 2570 15605 2590
rect 15625 2570 15630 2590
rect 15600 2540 15630 2570
rect 15600 2520 15605 2540
rect 15625 2520 15630 2540
rect 15600 2490 15630 2520
rect 15600 2470 15605 2490
rect 15625 2470 15630 2490
rect 15600 2460 15630 2470
rect 15655 2640 15685 2650
rect 15655 2620 15660 2640
rect 15680 2620 15685 2640
rect 15655 2590 15685 2620
rect 15655 2570 15660 2590
rect 15680 2570 15685 2590
rect 15655 2540 15685 2570
rect 15655 2520 15660 2540
rect 15680 2520 15685 2540
rect 15655 2490 15685 2520
rect 15655 2470 15660 2490
rect 15680 2470 15685 2490
rect 15655 2460 15685 2470
rect 15710 2640 15740 2650
rect 15710 2620 15715 2640
rect 15735 2620 15740 2640
rect 15710 2590 15740 2620
rect 15710 2570 15715 2590
rect 15735 2570 15740 2590
rect 15710 2540 15740 2570
rect 15710 2520 15715 2540
rect 15735 2520 15740 2540
rect 15710 2490 15740 2520
rect 15710 2470 15715 2490
rect 15735 2470 15740 2490
rect 15710 2460 15740 2470
rect 15765 2640 15795 2650
rect 15765 2620 15770 2640
rect 15790 2620 15795 2640
rect 15765 2590 15795 2620
rect 15765 2570 15770 2590
rect 15790 2570 15795 2590
rect 15765 2540 15795 2570
rect 15765 2520 15770 2540
rect 15790 2520 15795 2540
rect 15765 2490 15795 2520
rect 15765 2470 15770 2490
rect 15790 2470 15795 2490
rect 15765 2460 15795 2470
rect 15820 2640 15890 2650
rect 15820 2620 15825 2640
rect 15845 2620 15865 2640
rect 15885 2620 15890 2640
rect 15820 2590 15890 2620
rect 15820 2570 15825 2590
rect 15845 2570 15865 2590
rect 15885 2570 15890 2590
rect 15820 2540 15890 2570
rect 15820 2520 15825 2540
rect 15845 2520 15865 2540
rect 15885 2520 15890 2540
rect 15820 2490 15890 2520
rect 16185 2630 16255 2660
rect 16185 2610 16190 2630
rect 16210 2610 16230 2630
rect 16250 2610 16255 2630
rect 16185 2580 16255 2610
rect 16185 2560 16190 2580
rect 16210 2560 16230 2580
rect 16250 2560 16255 2580
rect 16185 2530 16255 2560
rect 16185 2510 16190 2530
rect 16210 2510 16230 2530
rect 16250 2510 16255 2530
rect 16185 2500 16255 2510
rect 16285 2880 16315 2890
rect 16285 2860 16290 2880
rect 16310 2860 16315 2880
rect 16285 2830 16315 2860
rect 16285 2810 16290 2830
rect 16310 2810 16315 2830
rect 16285 2780 16315 2810
rect 16285 2760 16290 2780
rect 16310 2760 16315 2780
rect 16285 2730 16315 2760
rect 16285 2710 16290 2730
rect 16310 2710 16315 2730
rect 16285 2680 16315 2710
rect 16285 2660 16290 2680
rect 16310 2660 16315 2680
rect 16285 2630 16315 2660
rect 16285 2610 16290 2630
rect 16310 2610 16315 2630
rect 16285 2580 16315 2610
rect 16285 2560 16290 2580
rect 16310 2560 16315 2580
rect 16285 2530 16315 2560
rect 16285 2510 16290 2530
rect 16310 2510 16315 2530
rect 16285 2500 16315 2510
rect 16345 2880 16375 2890
rect 16345 2860 16350 2880
rect 16370 2860 16375 2880
rect 16345 2830 16375 2860
rect 16345 2810 16350 2830
rect 16370 2810 16375 2830
rect 16345 2780 16375 2810
rect 16345 2760 16350 2780
rect 16370 2760 16375 2780
rect 16345 2730 16375 2760
rect 16345 2710 16350 2730
rect 16370 2710 16375 2730
rect 16345 2680 16375 2710
rect 16345 2660 16350 2680
rect 16370 2660 16375 2680
rect 16345 2630 16375 2660
rect 16345 2610 16350 2630
rect 16370 2610 16375 2630
rect 16345 2580 16375 2610
rect 16345 2560 16350 2580
rect 16370 2560 16375 2580
rect 16345 2530 16375 2560
rect 16345 2510 16350 2530
rect 16370 2510 16375 2530
rect 16345 2500 16375 2510
rect 16405 2880 16435 2890
rect 16405 2860 16410 2880
rect 16430 2860 16435 2880
rect 16405 2830 16435 2860
rect 16405 2810 16410 2830
rect 16430 2810 16435 2830
rect 16405 2780 16435 2810
rect 16405 2760 16410 2780
rect 16430 2760 16435 2780
rect 16405 2730 16435 2760
rect 16405 2710 16410 2730
rect 16430 2710 16435 2730
rect 16405 2680 16435 2710
rect 16405 2660 16410 2680
rect 16430 2660 16435 2680
rect 16405 2630 16435 2660
rect 16405 2610 16410 2630
rect 16430 2610 16435 2630
rect 16405 2580 16435 2610
rect 16405 2560 16410 2580
rect 16430 2560 16435 2580
rect 16405 2530 16435 2560
rect 16405 2510 16410 2530
rect 16430 2510 16435 2530
rect 16405 2500 16435 2510
rect 16465 2880 16495 2890
rect 16465 2860 16470 2880
rect 16490 2860 16495 2880
rect 16465 2830 16495 2860
rect 16465 2810 16470 2830
rect 16490 2810 16495 2830
rect 16465 2780 16495 2810
rect 16465 2760 16470 2780
rect 16490 2760 16495 2780
rect 16465 2730 16495 2760
rect 16465 2710 16470 2730
rect 16490 2710 16495 2730
rect 16465 2680 16495 2710
rect 16465 2660 16470 2680
rect 16490 2660 16495 2680
rect 16465 2630 16495 2660
rect 16465 2610 16470 2630
rect 16490 2610 16495 2630
rect 16465 2580 16495 2610
rect 16465 2560 16470 2580
rect 16490 2560 16495 2580
rect 16465 2530 16495 2560
rect 16465 2510 16470 2530
rect 16490 2510 16495 2530
rect 16465 2500 16495 2510
rect 16525 2880 16555 2890
rect 16525 2860 16530 2880
rect 16550 2860 16555 2880
rect 16525 2830 16555 2860
rect 16525 2810 16530 2830
rect 16550 2810 16555 2830
rect 16525 2780 16555 2810
rect 16525 2760 16530 2780
rect 16550 2760 16555 2780
rect 16525 2730 16555 2760
rect 16525 2710 16530 2730
rect 16550 2710 16555 2730
rect 16525 2680 16555 2710
rect 16525 2660 16530 2680
rect 16550 2660 16555 2680
rect 16525 2630 16555 2660
rect 16525 2610 16530 2630
rect 16550 2610 16555 2630
rect 16525 2580 16555 2610
rect 16525 2560 16530 2580
rect 16550 2560 16555 2580
rect 16525 2530 16555 2560
rect 16525 2510 16530 2530
rect 16550 2510 16555 2530
rect 16525 2500 16555 2510
rect 16585 2880 16615 2890
rect 16585 2860 16590 2880
rect 16610 2860 16615 2880
rect 16585 2830 16615 2860
rect 16585 2810 16590 2830
rect 16610 2810 16615 2830
rect 16585 2780 16615 2810
rect 16585 2760 16590 2780
rect 16610 2760 16615 2780
rect 16585 2730 16615 2760
rect 16585 2710 16590 2730
rect 16610 2710 16615 2730
rect 16585 2680 16615 2710
rect 16585 2660 16590 2680
rect 16610 2660 16615 2680
rect 16585 2630 16615 2660
rect 16585 2610 16590 2630
rect 16610 2610 16615 2630
rect 16585 2580 16615 2610
rect 16585 2560 16590 2580
rect 16610 2560 16615 2580
rect 16585 2530 16615 2560
rect 16585 2510 16590 2530
rect 16610 2510 16615 2530
rect 16585 2500 16615 2510
rect 16645 2880 16675 2890
rect 16645 2860 16650 2880
rect 16670 2860 16675 2880
rect 16645 2830 16675 2860
rect 16645 2810 16650 2830
rect 16670 2810 16675 2830
rect 16645 2780 16675 2810
rect 16645 2760 16650 2780
rect 16670 2760 16675 2780
rect 16645 2730 16675 2760
rect 16645 2710 16650 2730
rect 16670 2710 16675 2730
rect 16645 2680 16675 2710
rect 16645 2660 16650 2680
rect 16670 2660 16675 2680
rect 16645 2630 16675 2660
rect 16645 2610 16650 2630
rect 16670 2610 16675 2630
rect 16645 2580 16675 2610
rect 16645 2560 16650 2580
rect 16670 2560 16675 2580
rect 16645 2530 16675 2560
rect 16645 2510 16650 2530
rect 16670 2510 16675 2530
rect 16645 2500 16675 2510
rect 16705 2880 16735 2890
rect 16705 2860 16710 2880
rect 16730 2860 16735 2880
rect 16705 2830 16735 2860
rect 16705 2810 16710 2830
rect 16730 2810 16735 2830
rect 16705 2780 16735 2810
rect 16705 2760 16710 2780
rect 16730 2760 16735 2780
rect 16705 2730 16735 2760
rect 16705 2710 16710 2730
rect 16730 2710 16735 2730
rect 16705 2680 16735 2710
rect 16705 2660 16710 2680
rect 16730 2660 16735 2680
rect 16705 2630 16735 2660
rect 16705 2610 16710 2630
rect 16730 2610 16735 2630
rect 16705 2580 16735 2610
rect 16705 2560 16710 2580
rect 16730 2560 16735 2580
rect 16705 2530 16735 2560
rect 16705 2510 16710 2530
rect 16730 2510 16735 2530
rect 16705 2500 16735 2510
rect 16765 2880 16795 2890
rect 16765 2860 16770 2880
rect 16790 2860 16795 2880
rect 16765 2830 16795 2860
rect 16765 2810 16770 2830
rect 16790 2810 16795 2830
rect 16765 2780 16795 2810
rect 16765 2760 16770 2780
rect 16790 2760 16795 2780
rect 16765 2730 16795 2760
rect 16765 2710 16770 2730
rect 16790 2710 16795 2730
rect 16765 2680 16795 2710
rect 16765 2660 16770 2680
rect 16790 2660 16795 2680
rect 16765 2630 16795 2660
rect 16765 2610 16770 2630
rect 16790 2610 16795 2630
rect 16765 2580 16795 2610
rect 16765 2560 16770 2580
rect 16790 2560 16795 2580
rect 16765 2530 16795 2560
rect 16765 2510 16770 2530
rect 16790 2510 16795 2530
rect 16765 2500 16795 2510
rect 16825 2880 16855 2890
rect 16825 2860 16830 2880
rect 16850 2860 16855 2880
rect 16825 2830 16855 2860
rect 16825 2810 16830 2830
rect 16850 2810 16855 2830
rect 16825 2780 16855 2810
rect 16825 2760 16830 2780
rect 16850 2760 16855 2780
rect 16825 2730 16855 2760
rect 16825 2710 16830 2730
rect 16850 2710 16855 2730
rect 16825 2680 16855 2710
rect 16825 2660 16830 2680
rect 16850 2660 16855 2680
rect 16825 2630 16855 2660
rect 16825 2610 16830 2630
rect 16850 2610 16855 2630
rect 16825 2580 16855 2610
rect 16825 2560 16830 2580
rect 16850 2560 16855 2580
rect 16825 2530 16855 2560
rect 16825 2510 16830 2530
rect 16850 2510 16855 2530
rect 16825 2500 16855 2510
rect 16885 2880 16915 2890
rect 16885 2860 16890 2880
rect 16910 2860 16915 2880
rect 16885 2830 16915 2860
rect 16885 2810 16890 2830
rect 16910 2810 16915 2830
rect 16885 2780 16915 2810
rect 16885 2760 16890 2780
rect 16910 2760 16915 2780
rect 16885 2730 16915 2760
rect 16885 2710 16890 2730
rect 16910 2710 16915 2730
rect 16885 2680 16915 2710
rect 16885 2660 16890 2680
rect 16910 2660 16915 2680
rect 16885 2630 16915 2660
rect 16885 2610 16890 2630
rect 16910 2610 16915 2630
rect 16885 2580 16915 2610
rect 16885 2560 16890 2580
rect 16910 2560 16915 2580
rect 16885 2530 16915 2560
rect 16885 2510 16890 2530
rect 16910 2510 16915 2530
rect 16885 2500 16915 2510
rect 16945 2880 16975 2890
rect 16945 2860 16950 2880
rect 16970 2860 16975 2880
rect 16945 2830 16975 2860
rect 16945 2810 16950 2830
rect 16970 2810 16975 2830
rect 16945 2780 16975 2810
rect 16945 2760 16950 2780
rect 16970 2760 16975 2780
rect 16945 2730 16975 2760
rect 16945 2710 16950 2730
rect 16970 2710 16975 2730
rect 16945 2680 16975 2710
rect 16945 2660 16950 2680
rect 16970 2660 16975 2680
rect 16945 2630 16975 2660
rect 16945 2610 16950 2630
rect 16970 2610 16975 2630
rect 16945 2580 16975 2610
rect 16945 2560 16950 2580
rect 16970 2560 16975 2580
rect 16945 2530 16975 2560
rect 16945 2510 16950 2530
rect 16970 2510 16975 2530
rect 16945 2500 16975 2510
rect 17005 2880 17035 2890
rect 17005 2860 17010 2880
rect 17030 2860 17035 2880
rect 17005 2830 17035 2860
rect 17005 2810 17010 2830
rect 17030 2810 17035 2830
rect 17005 2780 17035 2810
rect 17005 2760 17010 2780
rect 17030 2760 17035 2780
rect 17005 2730 17035 2760
rect 17005 2710 17010 2730
rect 17030 2710 17035 2730
rect 17005 2680 17035 2710
rect 17005 2660 17010 2680
rect 17030 2660 17035 2680
rect 17005 2630 17035 2660
rect 17005 2610 17010 2630
rect 17030 2610 17035 2630
rect 17005 2580 17035 2610
rect 17005 2560 17010 2580
rect 17030 2560 17035 2580
rect 17005 2530 17035 2560
rect 17005 2510 17010 2530
rect 17030 2510 17035 2530
rect 17005 2500 17035 2510
rect 17065 2880 17095 2890
rect 17065 2860 17070 2880
rect 17090 2860 17095 2880
rect 17065 2830 17095 2860
rect 17065 2810 17070 2830
rect 17090 2810 17095 2830
rect 17065 2780 17095 2810
rect 17065 2760 17070 2780
rect 17090 2760 17095 2780
rect 17065 2730 17095 2760
rect 17065 2710 17070 2730
rect 17090 2710 17095 2730
rect 17065 2680 17095 2710
rect 17065 2660 17070 2680
rect 17090 2660 17095 2680
rect 17065 2630 17095 2660
rect 17065 2610 17070 2630
rect 17090 2610 17095 2630
rect 17065 2580 17095 2610
rect 17065 2560 17070 2580
rect 17090 2560 17095 2580
rect 17065 2530 17095 2560
rect 17065 2510 17070 2530
rect 17090 2510 17095 2530
rect 17065 2500 17095 2510
rect 17125 2880 17155 2890
rect 17125 2860 17130 2880
rect 17150 2860 17155 2880
rect 17125 2830 17155 2860
rect 17125 2810 17130 2830
rect 17150 2810 17155 2830
rect 17125 2780 17155 2810
rect 17125 2760 17130 2780
rect 17150 2760 17155 2780
rect 17125 2730 17155 2760
rect 17125 2710 17130 2730
rect 17150 2710 17155 2730
rect 17125 2680 17155 2710
rect 17125 2660 17130 2680
rect 17150 2660 17155 2680
rect 17125 2630 17155 2660
rect 17125 2610 17130 2630
rect 17150 2610 17155 2630
rect 17125 2580 17155 2610
rect 17125 2560 17130 2580
rect 17150 2560 17155 2580
rect 17125 2530 17155 2560
rect 17125 2510 17130 2530
rect 17150 2510 17155 2530
rect 17125 2500 17155 2510
rect 17185 2880 17215 2890
rect 17185 2860 17190 2880
rect 17210 2860 17215 2880
rect 17185 2830 17215 2860
rect 17185 2810 17190 2830
rect 17210 2810 17215 2830
rect 17185 2780 17215 2810
rect 17185 2760 17190 2780
rect 17210 2760 17215 2780
rect 17185 2730 17215 2760
rect 17185 2710 17190 2730
rect 17210 2710 17215 2730
rect 17185 2680 17215 2710
rect 17185 2660 17190 2680
rect 17210 2660 17215 2680
rect 17185 2630 17215 2660
rect 17185 2610 17190 2630
rect 17210 2610 17215 2630
rect 17185 2580 17215 2610
rect 17185 2560 17190 2580
rect 17210 2560 17215 2580
rect 17185 2530 17215 2560
rect 17185 2510 17190 2530
rect 17210 2510 17215 2530
rect 17185 2500 17215 2510
rect 17245 2880 17275 2890
rect 17245 2860 17250 2880
rect 17270 2860 17275 2880
rect 17245 2830 17275 2860
rect 17245 2810 17250 2830
rect 17270 2810 17275 2830
rect 17245 2780 17275 2810
rect 17245 2760 17250 2780
rect 17270 2760 17275 2780
rect 17245 2730 17275 2760
rect 17245 2710 17250 2730
rect 17270 2710 17275 2730
rect 17245 2680 17275 2710
rect 17245 2660 17250 2680
rect 17270 2660 17275 2680
rect 17245 2630 17275 2660
rect 17245 2610 17250 2630
rect 17270 2610 17275 2630
rect 17245 2580 17275 2610
rect 17245 2560 17250 2580
rect 17270 2560 17275 2580
rect 17245 2530 17275 2560
rect 17245 2510 17250 2530
rect 17270 2510 17275 2530
rect 17245 2500 17275 2510
rect 17305 2880 17335 2890
rect 17305 2860 17310 2880
rect 17330 2860 17335 2880
rect 17305 2830 17335 2860
rect 17305 2810 17310 2830
rect 17330 2810 17335 2830
rect 17305 2780 17335 2810
rect 17305 2760 17310 2780
rect 17330 2760 17335 2780
rect 17305 2730 17335 2760
rect 17305 2710 17310 2730
rect 17330 2710 17335 2730
rect 17305 2680 17335 2710
rect 17305 2660 17310 2680
rect 17330 2660 17335 2680
rect 17305 2630 17335 2660
rect 17305 2610 17310 2630
rect 17330 2610 17335 2630
rect 17305 2580 17335 2610
rect 17305 2560 17310 2580
rect 17330 2560 17335 2580
rect 17305 2530 17335 2560
rect 17305 2510 17310 2530
rect 17330 2510 17335 2530
rect 17305 2500 17335 2510
rect 17365 2880 17395 2890
rect 17365 2860 17370 2880
rect 17390 2860 17395 2880
rect 17365 2830 17395 2860
rect 17365 2810 17370 2830
rect 17390 2810 17395 2830
rect 17365 2780 17395 2810
rect 17365 2760 17370 2780
rect 17390 2760 17395 2780
rect 17365 2730 17395 2760
rect 17365 2710 17370 2730
rect 17390 2710 17395 2730
rect 17365 2680 17395 2710
rect 17365 2660 17370 2680
rect 17390 2660 17395 2680
rect 17365 2630 17395 2660
rect 17365 2610 17370 2630
rect 17390 2610 17395 2630
rect 17365 2580 17395 2610
rect 17365 2560 17370 2580
rect 17390 2560 17395 2580
rect 17365 2530 17395 2560
rect 17365 2510 17370 2530
rect 17390 2510 17395 2530
rect 17365 2500 17395 2510
rect 17425 2880 17455 2890
rect 17425 2860 17430 2880
rect 17450 2860 17455 2880
rect 17425 2830 17455 2860
rect 17425 2810 17430 2830
rect 17450 2810 17455 2830
rect 17425 2780 17455 2810
rect 17425 2760 17430 2780
rect 17450 2760 17455 2780
rect 17425 2730 17455 2760
rect 17425 2710 17430 2730
rect 17450 2710 17455 2730
rect 17425 2680 17455 2710
rect 17425 2660 17430 2680
rect 17450 2660 17455 2680
rect 17425 2630 17455 2660
rect 17425 2610 17430 2630
rect 17450 2610 17455 2630
rect 17425 2580 17455 2610
rect 17425 2560 17430 2580
rect 17450 2560 17455 2580
rect 17425 2530 17455 2560
rect 17425 2510 17430 2530
rect 17450 2510 17455 2530
rect 17425 2500 17455 2510
rect 17485 2880 17515 2890
rect 17485 2860 17490 2880
rect 17510 2860 17515 2880
rect 17485 2830 17515 2860
rect 17485 2810 17490 2830
rect 17510 2810 17515 2830
rect 17485 2780 17515 2810
rect 17485 2760 17490 2780
rect 17510 2760 17515 2780
rect 17485 2730 17515 2760
rect 17485 2710 17490 2730
rect 17510 2710 17515 2730
rect 17485 2680 17515 2710
rect 17485 2660 17490 2680
rect 17510 2660 17515 2680
rect 17485 2630 17515 2660
rect 17485 2610 17490 2630
rect 17510 2610 17515 2630
rect 17485 2580 17515 2610
rect 17485 2560 17490 2580
rect 17510 2560 17515 2580
rect 17485 2530 17515 2560
rect 17485 2510 17490 2530
rect 17510 2510 17515 2530
rect 17485 2500 17515 2510
rect 17545 2880 17615 2890
rect 17545 2860 17550 2880
rect 17570 2860 17590 2880
rect 17610 2860 17615 2880
rect 17545 2830 17615 2860
rect 17545 2810 17550 2830
rect 17570 2810 17590 2830
rect 17610 2810 17615 2830
rect 17545 2780 17615 2810
rect 17545 2760 17550 2780
rect 17570 2760 17590 2780
rect 17610 2760 17615 2780
rect 17545 2730 17615 2760
rect 17545 2710 17550 2730
rect 17570 2710 17590 2730
rect 17610 2710 17615 2730
rect 17545 2680 17615 2710
rect 17545 2660 17550 2680
rect 17570 2660 17590 2680
rect 17610 2660 17615 2680
rect 18000 2700 18040 2710
rect 18000 2680 18010 2700
rect 18030 2680 18040 2700
rect 18000 2670 18040 2680
rect 18110 2700 18150 2710
rect 18110 2680 18120 2700
rect 18140 2680 18150 2700
rect 18110 2670 18150 2680
rect 18220 2700 18260 2710
rect 18220 2680 18230 2700
rect 18250 2680 18260 2700
rect 18220 2670 18260 2680
rect 18330 2700 18370 2710
rect 18330 2680 18340 2700
rect 18360 2680 18370 2700
rect 18330 2670 18370 2680
rect 18440 2700 18480 2710
rect 18440 2680 18450 2700
rect 18470 2680 18480 2700
rect 18440 2670 18480 2680
rect 18550 2700 18590 2710
rect 18550 2680 18560 2700
rect 18580 2680 18590 2700
rect 18550 2670 18590 2680
rect 17545 2630 17615 2660
rect 18010 2650 18030 2670
rect 18120 2650 18140 2670
rect 18230 2650 18250 2670
rect 18340 2650 18360 2670
rect 18450 2650 18470 2670
rect 18560 2650 18580 2670
rect 17545 2610 17550 2630
rect 17570 2610 17590 2630
rect 17610 2610 17615 2630
rect 17545 2580 17615 2610
rect 17545 2560 17550 2580
rect 17570 2560 17590 2580
rect 17610 2560 17615 2580
rect 17545 2530 17615 2560
rect 17545 2510 17550 2530
rect 17570 2510 17590 2530
rect 17610 2510 17615 2530
rect 17545 2500 17615 2510
rect 17910 2640 17980 2650
rect 17910 2620 17915 2640
rect 17935 2620 17955 2640
rect 17975 2620 17980 2640
rect 17910 2590 17980 2620
rect 17910 2570 17915 2590
rect 17935 2570 17955 2590
rect 17975 2570 17980 2590
rect 17910 2540 17980 2570
rect 17910 2520 17915 2540
rect 17935 2520 17955 2540
rect 17975 2520 17980 2540
rect 15820 2470 15825 2490
rect 15845 2470 15865 2490
rect 15885 2470 15890 2490
rect 16290 2480 16310 2500
rect 16410 2480 16430 2500
rect 16530 2480 16550 2500
rect 16650 2480 16670 2500
rect 16770 2480 16790 2500
rect 16890 2480 16910 2500
rect 17010 2480 17030 2500
rect 17130 2480 17150 2500
rect 17250 2480 17270 2500
rect 17370 2480 17390 2500
rect 17490 2480 17510 2500
rect 17910 2490 17980 2520
rect 15820 2460 15890 2470
rect 16280 2470 16320 2480
rect 15125 2440 15145 2460
rect 15275 2440 15295 2460
rect 15385 2440 15405 2460
rect 15495 2440 15515 2460
rect 15605 2440 15625 2460
rect 15715 2440 15735 2460
rect 15865 2440 15885 2460
rect 16280 2450 16290 2470
rect 16310 2450 16320 2470
rect 16280 2440 16320 2450
rect 16400 2470 16440 2480
rect 16400 2450 16410 2470
rect 16430 2450 16440 2470
rect 16400 2440 16440 2450
rect 16520 2470 16560 2480
rect 16520 2450 16530 2470
rect 16550 2450 16560 2470
rect 16520 2440 16560 2450
rect 16640 2470 16680 2480
rect 16640 2450 16650 2470
rect 16670 2450 16680 2470
rect 16640 2440 16680 2450
rect 16760 2470 16800 2480
rect 16760 2450 16770 2470
rect 16790 2450 16800 2470
rect 16760 2440 16800 2450
rect 16823 2470 16857 2480
rect 16823 2450 16831 2470
rect 16849 2450 16857 2470
rect 16823 2440 16857 2450
rect 16880 2470 16920 2480
rect 16880 2450 16890 2470
rect 16910 2450 16920 2470
rect 16880 2440 16920 2450
rect 17000 2470 17040 2480
rect 17000 2450 17010 2470
rect 17030 2450 17040 2470
rect 17000 2440 17040 2450
rect 17120 2470 17160 2480
rect 17120 2450 17130 2470
rect 17150 2450 17160 2470
rect 17120 2440 17160 2450
rect 17240 2470 17280 2480
rect 17240 2450 17250 2470
rect 17270 2450 17280 2470
rect 17240 2440 17280 2450
rect 17360 2470 17400 2480
rect 17360 2450 17370 2470
rect 17390 2450 17400 2470
rect 17360 2440 17400 2450
rect 17480 2470 17520 2480
rect 17480 2450 17490 2470
rect 17510 2450 17520 2470
rect 17910 2470 17915 2490
rect 17935 2470 17955 2490
rect 17975 2470 17980 2490
rect 17910 2460 17980 2470
rect 18005 2640 18035 2650
rect 18005 2620 18010 2640
rect 18030 2620 18035 2640
rect 18005 2590 18035 2620
rect 18005 2570 18010 2590
rect 18030 2570 18035 2590
rect 18005 2540 18035 2570
rect 18005 2520 18010 2540
rect 18030 2520 18035 2540
rect 18005 2490 18035 2520
rect 18005 2470 18010 2490
rect 18030 2470 18035 2490
rect 18005 2460 18035 2470
rect 18060 2640 18090 2650
rect 18060 2620 18065 2640
rect 18085 2620 18090 2640
rect 18060 2590 18090 2620
rect 18060 2570 18065 2590
rect 18085 2570 18090 2590
rect 18060 2540 18090 2570
rect 18060 2520 18065 2540
rect 18085 2520 18090 2540
rect 18060 2490 18090 2520
rect 18060 2470 18065 2490
rect 18085 2470 18090 2490
rect 18060 2460 18090 2470
rect 18115 2640 18145 2650
rect 18115 2620 18120 2640
rect 18140 2620 18145 2640
rect 18115 2590 18145 2620
rect 18115 2570 18120 2590
rect 18140 2570 18145 2590
rect 18115 2540 18145 2570
rect 18115 2520 18120 2540
rect 18140 2520 18145 2540
rect 18115 2490 18145 2520
rect 18115 2470 18120 2490
rect 18140 2470 18145 2490
rect 18115 2460 18145 2470
rect 18170 2640 18200 2650
rect 18170 2620 18175 2640
rect 18195 2620 18200 2640
rect 18170 2590 18200 2620
rect 18170 2570 18175 2590
rect 18195 2570 18200 2590
rect 18170 2540 18200 2570
rect 18170 2520 18175 2540
rect 18195 2520 18200 2540
rect 18170 2490 18200 2520
rect 18170 2470 18175 2490
rect 18195 2470 18200 2490
rect 18170 2460 18200 2470
rect 18225 2640 18255 2650
rect 18225 2620 18230 2640
rect 18250 2620 18255 2640
rect 18225 2590 18255 2620
rect 18225 2570 18230 2590
rect 18250 2570 18255 2590
rect 18225 2540 18255 2570
rect 18225 2520 18230 2540
rect 18250 2520 18255 2540
rect 18225 2490 18255 2520
rect 18225 2470 18230 2490
rect 18250 2470 18255 2490
rect 18225 2460 18255 2470
rect 18280 2640 18310 2650
rect 18280 2620 18285 2640
rect 18305 2620 18310 2640
rect 18280 2590 18310 2620
rect 18280 2570 18285 2590
rect 18305 2570 18310 2590
rect 18280 2540 18310 2570
rect 18280 2520 18285 2540
rect 18305 2520 18310 2540
rect 18280 2490 18310 2520
rect 18280 2470 18285 2490
rect 18305 2470 18310 2490
rect 18280 2460 18310 2470
rect 18335 2640 18365 2650
rect 18335 2620 18340 2640
rect 18360 2620 18365 2640
rect 18335 2590 18365 2620
rect 18335 2570 18340 2590
rect 18360 2570 18365 2590
rect 18335 2540 18365 2570
rect 18335 2520 18340 2540
rect 18360 2520 18365 2540
rect 18335 2490 18365 2520
rect 18335 2470 18340 2490
rect 18360 2470 18365 2490
rect 18335 2460 18365 2470
rect 18390 2640 18420 2650
rect 18390 2620 18395 2640
rect 18415 2620 18420 2640
rect 18390 2590 18420 2620
rect 18390 2570 18395 2590
rect 18415 2570 18420 2590
rect 18390 2540 18420 2570
rect 18390 2520 18395 2540
rect 18415 2520 18420 2540
rect 18390 2490 18420 2520
rect 18390 2470 18395 2490
rect 18415 2470 18420 2490
rect 18390 2460 18420 2470
rect 18445 2640 18475 2650
rect 18445 2620 18450 2640
rect 18470 2620 18475 2640
rect 18445 2590 18475 2620
rect 18445 2570 18450 2590
rect 18470 2570 18475 2590
rect 18445 2540 18475 2570
rect 18445 2520 18450 2540
rect 18470 2520 18475 2540
rect 18445 2490 18475 2520
rect 18445 2470 18450 2490
rect 18470 2470 18475 2490
rect 18445 2460 18475 2470
rect 18500 2640 18530 2650
rect 18500 2620 18505 2640
rect 18525 2620 18530 2640
rect 18500 2590 18530 2620
rect 18500 2570 18505 2590
rect 18525 2570 18530 2590
rect 18500 2540 18530 2570
rect 18500 2520 18505 2540
rect 18525 2520 18530 2540
rect 18500 2490 18530 2520
rect 18500 2470 18505 2490
rect 18525 2470 18530 2490
rect 18500 2460 18530 2470
rect 18555 2640 18585 2650
rect 18555 2620 18560 2640
rect 18580 2620 18585 2640
rect 18555 2590 18585 2620
rect 18555 2570 18560 2590
rect 18580 2570 18585 2590
rect 18555 2540 18585 2570
rect 18555 2520 18560 2540
rect 18580 2520 18585 2540
rect 18555 2490 18585 2520
rect 18555 2470 18560 2490
rect 18580 2470 18585 2490
rect 18555 2460 18585 2470
rect 18610 2640 18680 2650
rect 18610 2620 18615 2640
rect 18635 2620 18655 2640
rect 18675 2620 18680 2640
rect 18610 2590 18680 2620
rect 18610 2570 18615 2590
rect 18635 2570 18655 2590
rect 18675 2570 18680 2590
rect 18610 2540 18680 2570
rect 18610 2520 18615 2540
rect 18635 2520 18655 2540
rect 18675 2520 18680 2540
rect 18610 2490 18680 2520
rect 18610 2470 18615 2490
rect 18635 2470 18655 2490
rect 18675 2470 18680 2490
rect 18610 2460 18680 2470
rect 18795 2645 19010 2665
rect 18795 2625 18830 2645
rect 18975 2625 19010 2645
rect 17480 2440 17520 2450
rect 17915 2440 17935 2460
rect 18065 2440 18085 2460
rect 18175 2440 18195 2460
rect 18285 2440 18305 2460
rect 18395 2440 18415 2460
rect 18505 2440 18525 2460
rect 18655 2440 18675 2460
rect 15115 2430 15155 2440
rect 15115 2410 15125 2430
rect 15145 2410 15155 2430
rect 3275 2385 3295 2405
rect 3455 2385 3475 2405
rect 3265 2375 3305 2385
rect 3265 2355 3275 2375
rect 3295 2355 3305 2375
rect 3265 2345 3305 2355
rect 3355 2370 3395 2380
rect 3355 2350 3365 2370
rect 3385 2350 3395 2370
rect 2625 2315 2655 2345
rect 3355 2340 3395 2350
rect 3445 2375 3485 2385
rect 3445 2355 3455 2375
rect 3475 2355 3485 2375
rect 3445 2345 3485 2355
rect 3635 2340 3655 2405
rect 3815 2385 3835 2405
rect 3995 2385 4015 2405
rect 4175 2385 4195 2405
rect 3805 2375 3845 2385
rect 3805 2355 3815 2375
rect 3835 2355 3845 2375
rect 3805 2345 3845 2355
rect 3885 2375 3925 2385
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 3985 2375 4025 2385
rect 3985 2355 3995 2375
rect 4015 2355 4025 2375
rect 3985 2345 4025 2355
rect 4165 2375 4205 2385
rect 4165 2355 4175 2375
rect 4195 2355 4205 2375
rect 4165 2345 4205 2355
rect 4355 2340 4375 2405
rect 4535 2385 4555 2405
rect 4715 2385 4735 2405
rect 15115 2400 15155 2410
rect 15265 2430 15305 2440
rect 15265 2410 15275 2430
rect 15295 2410 15305 2430
rect 15265 2400 15305 2410
rect 15375 2430 15415 2440
rect 15375 2410 15385 2430
rect 15405 2410 15415 2430
rect 15375 2400 15415 2410
rect 15485 2430 15525 2440
rect 15485 2410 15495 2430
rect 15515 2410 15525 2430
rect 15485 2400 15525 2410
rect 15595 2430 15635 2440
rect 15595 2410 15605 2430
rect 15625 2410 15635 2430
rect 15595 2400 15635 2410
rect 15705 2430 15745 2440
rect 15705 2410 15715 2430
rect 15735 2410 15745 2430
rect 15705 2400 15745 2410
rect 15855 2430 15895 2440
rect 15855 2410 15865 2430
rect 15885 2410 15895 2430
rect 15855 2400 15895 2410
rect 17905 2430 17945 2440
rect 17905 2410 17915 2430
rect 17935 2410 17945 2430
rect 17905 2400 17945 2410
rect 18055 2430 18095 2440
rect 18055 2410 18065 2430
rect 18085 2410 18095 2430
rect 18055 2400 18095 2410
rect 18165 2430 18205 2440
rect 18165 2410 18175 2430
rect 18195 2410 18205 2430
rect 18165 2400 18205 2410
rect 18275 2430 18315 2440
rect 18275 2410 18285 2430
rect 18305 2410 18315 2430
rect 18275 2400 18315 2410
rect 18385 2430 18425 2440
rect 18385 2410 18395 2430
rect 18415 2410 18425 2430
rect 18385 2400 18425 2410
rect 18495 2430 18535 2440
rect 18495 2410 18505 2430
rect 18525 2410 18535 2430
rect 18495 2400 18535 2410
rect 18645 2430 18685 2440
rect 18645 2410 18655 2430
rect 18675 2410 18685 2430
rect 18645 2400 18685 2410
rect 18890 2575 18915 2625
rect 15765 2385 15805 2395
rect 4525 2375 4565 2385
rect 4525 2355 4535 2375
rect 4555 2355 4565 2375
rect 4525 2345 4565 2355
rect 4705 2375 4745 2385
rect 4705 2355 4715 2375
rect 4735 2355 4745 2375
rect 15765 2365 15775 2385
rect 15795 2365 15805 2385
rect 15765 2355 15805 2365
rect 18025 2370 18065 2380
rect 4705 2345 4745 2355
rect 18025 2350 18035 2370
rect 18055 2350 18065 2370
rect 18025 2340 18065 2350
rect 3625 2330 3665 2340
rect 3625 2310 3635 2330
rect 3655 2310 3665 2330
rect 3625 2300 3665 2310
rect 4345 2330 4385 2340
rect 4345 2310 4355 2330
rect 4375 2310 4385 2330
rect 4345 2300 4385 2310
rect 15115 2310 15155 2320
rect 2740 2260 2770 2290
rect 3445 2285 3485 2295
rect 3445 2265 3455 2285
rect 3475 2265 3485 2285
rect 3445 2255 3485 2265
rect 4525 2285 4565 2295
rect 15115 2290 15125 2310
rect 15145 2290 15155 2310
rect 4525 2265 4535 2285
rect 4555 2265 4565 2285
rect 4525 2255 4565 2265
rect 5275 2260 5305 2290
rect 15115 2280 15155 2290
rect 15265 2310 15305 2320
rect 15265 2290 15275 2310
rect 15295 2290 15305 2310
rect 15265 2280 15305 2290
rect 15375 2310 15415 2320
rect 15375 2290 15385 2310
rect 15405 2290 15415 2310
rect 15375 2280 15415 2290
rect 15485 2310 15525 2320
rect 15485 2290 15495 2310
rect 15515 2290 15525 2310
rect 15485 2280 15525 2290
rect 15595 2310 15635 2320
rect 15595 2290 15605 2310
rect 15625 2290 15635 2310
rect 15595 2280 15635 2290
rect 15705 2310 15745 2320
rect 15705 2290 15715 2310
rect 15735 2290 15745 2310
rect 15705 2280 15745 2290
rect 15855 2310 15895 2320
rect 15855 2290 15865 2310
rect 15885 2290 15895 2310
rect 15855 2280 15895 2290
rect 17905 2310 17945 2320
rect 17905 2290 17915 2310
rect 17935 2290 17945 2310
rect 17905 2280 17945 2290
rect 18055 2310 18095 2320
rect 18055 2290 18065 2310
rect 18085 2290 18095 2310
rect 18055 2280 18095 2290
rect 18165 2310 18205 2320
rect 18165 2290 18175 2310
rect 18195 2290 18205 2310
rect 18165 2280 18205 2290
rect 18275 2310 18315 2320
rect 18275 2290 18285 2310
rect 18305 2290 18315 2310
rect 18275 2280 18315 2290
rect 18385 2310 18425 2320
rect 18385 2290 18395 2310
rect 18415 2290 18425 2310
rect 18385 2280 18425 2290
rect 18495 2310 18535 2320
rect 18495 2290 18505 2310
rect 18525 2290 18535 2310
rect 18495 2280 18535 2290
rect 18645 2310 18685 2320
rect 18645 2290 18655 2310
rect 18675 2290 18685 2310
rect 18645 2280 18685 2290
rect 15125 2260 15145 2280
rect 15275 2260 15295 2280
rect 15385 2260 15405 2280
rect 15495 2260 15515 2280
rect 15605 2260 15625 2280
rect 15715 2260 15735 2280
rect 15865 2260 15885 2280
rect 17915 2260 17935 2280
rect 18065 2260 18085 2280
rect 18175 2260 18195 2280
rect 18285 2260 18305 2280
rect 18395 2260 18415 2280
rect 18505 2260 18525 2280
rect 18655 2260 18675 2280
rect 15120 2250 15190 2260
rect 2430 2215 2460 2245
rect 3810 2215 3840 2245
rect 15120 2230 15125 2250
rect 15145 2230 15165 2250
rect 15185 2230 15190 2250
rect 2335 2170 2365 2200
rect 2385 2120 2415 2150
rect 3630 2120 3660 2150
rect 4090 2115 4120 2145
rect 5320 2115 5350 2145
rect 2745 2090 2785 2100
rect 2745 2070 2755 2090
rect 2775 2070 2785 2090
rect 2745 2060 2785 2070
rect 2865 2090 2905 2100
rect 2865 2070 2875 2090
rect 2895 2070 2905 2090
rect 2865 2060 2905 2070
rect 2985 2090 3025 2100
rect 2985 2070 2995 2090
rect 3015 2070 3025 2090
rect 2985 2060 3025 2070
rect 3105 2090 3145 2100
rect 3105 2070 3115 2090
rect 3135 2070 3145 2090
rect 3105 2060 3145 2070
rect 3225 2090 3265 2100
rect 3225 2070 3235 2090
rect 3255 2070 3265 2090
rect 3225 2060 3265 2070
rect 3345 2090 3385 2100
rect 3345 2070 3355 2090
rect 3375 2070 3385 2090
rect 3345 2060 3385 2070
rect 3465 2090 3505 2100
rect 3465 2070 3475 2090
rect 3495 2070 3505 2090
rect 3465 2060 3505 2070
rect 3585 2090 3625 2100
rect 3585 2070 3595 2090
rect 3615 2070 3625 2090
rect 3585 2060 3625 2070
rect 3705 2090 3745 2100
rect 3705 2070 3715 2090
rect 3735 2070 3745 2090
rect 3705 2060 3745 2070
rect 3825 2090 3865 2100
rect 3825 2070 3835 2090
rect 3855 2070 3865 2090
rect 3825 2060 3865 2070
rect 3985 2090 4025 2100
rect 3985 2070 3995 2090
rect 4015 2070 4025 2090
rect 3985 2060 4025 2070
rect 4145 2090 4185 2100
rect 4145 2070 4155 2090
rect 4175 2070 4185 2090
rect 4145 2060 4185 2070
rect 4265 2090 4305 2100
rect 4265 2070 4275 2090
rect 4295 2070 4305 2090
rect 4265 2060 4305 2070
rect 4385 2090 4425 2100
rect 4385 2070 4395 2090
rect 4415 2070 4425 2090
rect 4385 2060 4425 2070
rect 4505 2090 4545 2100
rect 4505 2070 4515 2090
rect 4535 2070 4545 2090
rect 4505 2060 4545 2070
rect 4625 2090 4665 2100
rect 4625 2070 4635 2090
rect 4655 2070 4665 2090
rect 4625 2060 4665 2070
rect 4745 2090 4785 2100
rect 4745 2070 4755 2090
rect 4775 2070 4785 2090
rect 4745 2060 4785 2070
rect 4865 2090 4905 2100
rect 4865 2070 4875 2090
rect 4895 2070 4905 2090
rect 4865 2060 4905 2070
rect 4985 2090 5025 2100
rect 4985 2070 4995 2090
rect 5015 2070 5025 2090
rect 4985 2060 5025 2070
rect 5105 2090 5145 2100
rect 5105 2070 5115 2090
rect 5135 2070 5145 2090
rect 5105 2060 5145 2070
rect 5225 2090 5265 2100
rect 5225 2070 5235 2090
rect 5255 2070 5265 2090
rect 5225 2060 5265 2070
rect 125 2015 2135 2055
rect 2620 2045 2660 2055
rect 2620 2025 2630 2045
rect 2650 2025 2660 2045
rect 2620 2015 2660 2025
rect -45 1715 130 1725
rect -45 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 130 1715
rect -45 1685 130 1695
rect 650 1375 775 2015
rect 1330 1375 1455 2015
rect 2010 1375 2135 2015
rect 2630 1995 2650 2015
rect 2755 1995 2775 2060
rect 2805 2045 2845 2055
rect 2805 2025 2815 2045
rect 2835 2025 2845 2045
rect 2805 2015 2845 2025
rect 2815 1995 2835 2015
rect 2875 1995 2895 2060
rect 2995 1995 3015 2060
rect 3115 1995 3135 2060
rect 3165 2045 3205 2055
rect 3165 2025 3175 2045
rect 3195 2025 3205 2045
rect 3165 2015 3205 2025
rect 3175 1995 3195 2015
rect 3235 1995 3255 2060
rect 3355 1995 3375 2060
rect 3475 1995 3495 2060
rect 3525 2045 3565 2055
rect 3525 2025 3535 2045
rect 3555 2025 3565 2045
rect 3525 2015 3565 2025
rect 3535 1995 3555 2015
rect 3595 1995 3615 2060
rect 3715 1995 3735 2060
rect 3835 1995 3855 2060
rect 3885 2045 3925 2055
rect 3885 2025 3895 2045
rect 3915 2025 3925 2045
rect 3885 2015 3925 2025
rect 3895 1995 3915 2015
rect 3995 1995 4015 2060
rect 4085 2045 4125 2055
rect 4085 2025 4095 2045
rect 4115 2025 4125 2045
rect 4085 2015 4125 2025
rect 4095 1995 4115 2015
rect 4155 1995 4175 2060
rect 4275 1995 4295 2060
rect 4395 1995 4415 2060
rect 4445 2045 4485 2055
rect 4445 2025 4455 2045
rect 4475 2025 4485 2045
rect 4445 2015 4485 2025
rect 4455 1995 4475 2015
rect 4515 1995 4535 2060
rect 4635 1995 4655 2060
rect 4755 1995 4775 2060
rect 4805 2045 4845 2055
rect 4805 2025 4815 2045
rect 4835 2025 4845 2045
rect 4805 2015 4845 2025
rect 4815 1995 4835 2015
rect 4875 1995 4895 2060
rect 4995 1995 5015 2060
rect 5115 1995 5135 2060
rect 5165 2045 5205 2055
rect 5165 2025 5175 2045
rect 5195 2025 5205 2045
rect 5165 2015 5205 2025
rect 5175 1995 5195 2015
rect 5235 1995 5255 2060
rect 14790 2000 14825 2010
rect 2570 1985 2600 1995
rect 2570 1965 2575 1985
rect 2595 1965 2600 1985
rect 2570 1935 2600 1965
rect 2570 1915 2575 1935
rect 2595 1915 2600 1935
rect 2570 1905 2600 1915
rect 2625 1985 2655 1995
rect 2625 1965 2630 1985
rect 2650 1965 2655 1985
rect 2625 1935 2655 1965
rect 2625 1915 2630 1935
rect 2650 1915 2655 1935
rect 2625 1905 2655 1915
rect 2680 1985 2710 1995
rect 2680 1965 2685 1985
rect 2705 1965 2710 1985
rect 2680 1935 2710 1965
rect 2680 1915 2685 1935
rect 2705 1915 2710 1935
rect 2680 1905 2710 1915
rect 2750 1985 2780 1995
rect 2750 1965 2755 1985
rect 2775 1965 2780 1985
rect 2750 1935 2780 1965
rect 2750 1915 2755 1935
rect 2775 1915 2780 1935
rect 2750 1905 2780 1915
rect 2810 1985 2840 1995
rect 2810 1965 2815 1985
rect 2835 1965 2840 1985
rect 2810 1935 2840 1965
rect 2810 1915 2815 1935
rect 2835 1915 2840 1935
rect 2810 1905 2840 1915
rect 2870 1985 2900 1995
rect 2870 1965 2875 1985
rect 2895 1965 2900 1985
rect 2870 1935 2900 1965
rect 2870 1915 2875 1935
rect 2895 1915 2900 1935
rect 2870 1905 2900 1915
rect 2930 1985 2960 1995
rect 2930 1965 2935 1985
rect 2955 1965 2960 1985
rect 2930 1935 2960 1965
rect 2930 1915 2935 1935
rect 2955 1915 2960 1935
rect 2930 1905 2960 1915
rect 2990 1985 3020 1995
rect 2990 1965 2995 1985
rect 3015 1965 3020 1985
rect 2990 1935 3020 1965
rect 2990 1915 2995 1935
rect 3015 1915 3020 1935
rect 2990 1905 3020 1915
rect 3050 1985 3080 1995
rect 3050 1965 3055 1985
rect 3075 1965 3080 1985
rect 3050 1935 3080 1965
rect 3050 1915 3055 1935
rect 3075 1915 3080 1935
rect 3050 1905 3080 1915
rect 3110 1985 3140 1995
rect 3110 1965 3115 1985
rect 3135 1965 3140 1985
rect 3110 1935 3140 1965
rect 3110 1915 3115 1935
rect 3135 1915 3140 1935
rect 3110 1905 3140 1915
rect 3170 1985 3200 1995
rect 3170 1965 3175 1985
rect 3195 1965 3200 1985
rect 3170 1935 3200 1965
rect 3170 1915 3175 1935
rect 3195 1915 3200 1935
rect 3170 1905 3200 1915
rect 3230 1985 3260 1995
rect 3230 1965 3235 1985
rect 3255 1965 3260 1985
rect 3230 1935 3260 1965
rect 3230 1915 3235 1935
rect 3255 1915 3260 1935
rect 3230 1905 3260 1915
rect 3290 1985 3320 1995
rect 3290 1965 3295 1985
rect 3315 1965 3320 1985
rect 3290 1935 3320 1965
rect 3290 1915 3295 1935
rect 3315 1915 3320 1935
rect 3290 1905 3320 1915
rect 3350 1985 3380 1995
rect 3350 1965 3355 1985
rect 3375 1965 3380 1985
rect 3350 1935 3380 1965
rect 3350 1915 3355 1935
rect 3375 1915 3380 1935
rect 3350 1905 3380 1915
rect 3410 1985 3440 1995
rect 3410 1965 3415 1985
rect 3435 1965 3440 1985
rect 3410 1935 3440 1965
rect 3410 1915 3415 1935
rect 3435 1915 3440 1935
rect 3410 1905 3440 1915
rect 3470 1985 3500 1995
rect 3470 1965 3475 1985
rect 3495 1965 3500 1985
rect 3470 1935 3500 1965
rect 3470 1915 3475 1935
rect 3495 1915 3500 1935
rect 3470 1905 3500 1915
rect 3530 1985 3560 1995
rect 3530 1965 3535 1985
rect 3555 1965 3560 1985
rect 3530 1935 3560 1965
rect 3530 1915 3535 1935
rect 3555 1915 3560 1935
rect 3530 1905 3560 1915
rect 3590 1985 3620 1995
rect 3590 1965 3595 1985
rect 3615 1965 3620 1985
rect 3590 1935 3620 1965
rect 3590 1915 3595 1935
rect 3615 1915 3620 1935
rect 3590 1905 3620 1915
rect 3650 1985 3680 1995
rect 3650 1965 3655 1985
rect 3675 1965 3680 1985
rect 3650 1935 3680 1965
rect 3650 1915 3655 1935
rect 3675 1915 3680 1935
rect 3650 1905 3680 1915
rect 3710 1985 3740 1995
rect 3710 1965 3715 1985
rect 3735 1965 3740 1985
rect 3710 1935 3740 1965
rect 3710 1915 3715 1935
rect 3735 1915 3740 1935
rect 3710 1905 3740 1915
rect 3770 1985 3800 1995
rect 3770 1965 3775 1985
rect 3795 1965 3800 1985
rect 3770 1935 3800 1965
rect 3770 1915 3775 1935
rect 3795 1915 3800 1935
rect 3770 1905 3800 1915
rect 3830 1985 3860 1995
rect 3830 1965 3835 1985
rect 3855 1965 3860 1985
rect 3830 1935 3860 1965
rect 3830 1915 3835 1935
rect 3855 1915 3860 1935
rect 3830 1905 3860 1915
rect 3890 1985 3920 1995
rect 3890 1965 3895 1985
rect 3915 1965 3920 1985
rect 3890 1935 3920 1965
rect 3890 1915 3895 1935
rect 3915 1915 3920 1935
rect 3890 1905 3920 1915
rect 3950 1985 4060 1995
rect 3950 1965 3955 1985
rect 3975 1965 3995 1985
rect 4015 1965 4035 1985
rect 4055 1965 4060 1985
rect 3950 1935 4060 1965
rect 3950 1915 3955 1935
rect 3975 1915 3995 1935
rect 4015 1915 4035 1935
rect 4055 1915 4060 1935
rect 3950 1905 4060 1915
rect 4090 1985 4120 1995
rect 4090 1965 4095 1985
rect 4115 1965 4120 1985
rect 4090 1935 4120 1965
rect 4090 1915 4095 1935
rect 4115 1915 4120 1935
rect 4090 1905 4120 1915
rect 4150 1985 4180 1995
rect 4150 1965 4155 1985
rect 4175 1965 4180 1985
rect 4150 1935 4180 1965
rect 4150 1915 4155 1935
rect 4175 1915 4180 1935
rect 4150 1905 4180 1915
rect 4210 1985 4240 1995
rect 4210 1965 4215 1985
rect 4235 1965 4240 1985
rect 4210 1935 4240 1965
rect 4210 1915 4215 1935
rect 4235 1915 4240 1935
rect 4210 1905 4240 1915
rect 4270 1985 4300 1995
rect 4270 1965 4275 1985
rect 4295 1965 4300 1985
rect 4270 1935 4300 1965
rect 4270 1915 4275 1935
rect 4295 1915 4300 1935
rect 4270 1905 4300 1915
rect 4330 1985 4360 1995
rect 4330 1965 4335 1985
rect 4355 1965 4360 1985
rect 4330 1935 4360 1965
rect 4330 1915 4335 1935
rect 4355 1915 4360 1935
rect 4330 1905 4360 1915
rect 4390 1985 4420 1995
rect 4390 1965 4395 1985
rect 4415 1965 4420 1985
rect 4390 1935 4420 1965
rect 4390 1915 4395 1935
rect 4415 1915 4420 1935
rect 4390 1905 4420 1915
rect 4450 1985 4480 1995
rect 4450 1965 4455 1985
rect 4475 1965 4480 1985
rect 4450 1935 4480 1965
rect 4450 1915 4455 1935
rect 4475 1915 4480 1935
rect 4450 1905 4480 1915
rect 4510 1985 4540 1995
rect 4510 1965 4515 1985
rect 4535 1965 4540 1985
rect 4510 1935 4540 1965
rect 4510 1915 4515 1935
rect 4535 1915 4540 1935
rect 4510 1905 4540 1915
rect 4570 1985 4600 1995
rect 4570 1965 4575 1985
rect 4595 1965 4600 1985
rect 4570 1935 4600 1965
rect 4570 1915 4575 1935
rect 4595 1915 4600 1935
rect 4570 1905 4600 1915
rect 4630 1985 4660 1995
rect 4630 1965 4635 1985
rect 4655 1965 4660 1985
rect 4630 1935 4660 1965
rect 4630 1915 4635 1935
rect 4655 1915 4660 1935
rect 4630 1905 4660 1915
rect 4690 1985 4720 1995
rect 4690 1965 4695 1985
rect 4715 1965 4720 1985
rect 4690 1935 4720 1965
rect 4690 1915 4695 1935
rect 4715 1915 4720 1935
rect 4690 1905 4720 1915
rect 4750 1985 4780 1995
rect 4750 1965 4755 1985
rect 4775 1965 4780 1985
rect 4750 1935 4780 1965
rect 4750 1915 4755 1935
rect 4775 1915 4780 1935
rect 4750 1905 4780 1915
rect 4810 1985 4840 1995
rect 4810 1965 4815 1985
rect 4835 1965 4840 1985
rect 4810 1935 4840 1965
rect 4810 1915 4815 1935
rect 4835 1915 4840 1935
rect 4810 1905 4840 1915
rect 4870 1985 4900 1995
rect 4870 1965 4875 1985
rect 4895 1965 4900 1985
rect 4870 1935 4900 1965
rect 4870 1915 4875 1935
rect 4895 1915 4900 1935
rect 4870 1905 4900 1915
rect 4930 1985 4960 1995
rect 4930 1965 4935 1985
rect 4955 1965 4960 1985
rect 4930 1935 4960 1965
rect 4930 1915 4935 1935
rect 4955 1915 4960 1935
rect 4930 1905 4960 1915
rect 4990 1985 5020 1995
rect 4990 1965 4995 1985
rect 5015 1965 5020 1985
rect 4990 1935 5020 1965
rect 4990 1915 4995 1935
rect 5015 1915 5020 1935
rect 4990 1905 5020 1915
rect 5050 1985 5080 1995
rect 5050 1965 5055 1985
rect 5075 1965 5080 1985
rect 5050 1935 5080 1965
rect 5050 1915 5055 1935
rect 5075 1915 5080 1935
rect 5050 1905 5080 1915
rect 5110 1985 5140 1995
rect 5110 1965 5115 1985
rect 5135 1965 5140 1985
rect 5110 1935 5140 1965
rect 5110 1915 5115 1935
rect 5135 1915 5140 1935
rect 5110 1905 5140 1915
rect 5170 1985 5200 1995
rect 5170 1965 5175 1985
rect 5195 1965 5200 1985
rect 5170 1935 5200 1965
rect 5170 1915 5175 1935
rect 5195 1915 5200 1935
rect 5170 1905 5200 1915
rect 5230 1985 5260 1995
rect 5230 1965 5235 1985
rect 5255 1965 5260 1985
rect 14790 1975 14795 2000
rect 14820 1975 14825 2000
rect 14790 1965 14825 1975
rect 14850 2000 14885 2010
rect 14850 1975 14855 2000
rect 14880 1975 14885 2000
rect 14850 1965 14885 1975
rect 14910 2000 14945 2010
rect 14910 1975 14915 2000
rect 14940 1975 14945 2000
rect 14910 1965 14945 1975
rect 14970 2000 15005 2010
rect 14970 1975 14975 2000
rect 15000 1975 15005 2000
rect 14970 1965 15005 1975
rect 15120 2200 15190 2230
rect 15120 2180 15125 2200
rect 15145 2180 15165 2200
rect 15185 2180 15190 2200
rect 15120 2150 15190 2180
rect 15120 2130 15125 2150
rect 15145 2130 15165 2150
rect 15185 2130 15190 2150
rect 15120 2100 15190 2130
rect 15120 2080 15125 2100
rect 15145 2080 15165 2100
rect 15185 2080 15190 2100
rect 15120 2050 15190 2080
rect 15120 2030 15125 2050
rect 15145 2030 15165 2050
rect 15185 2030 15190 2050
rect 15120 2000 15190 2030
rect 15120 1980 15125 2000
rect 15145 1980 15165 2000
rect 15185 1980 15190 2000
rect 15120 1970 15190 1980
rect 15215 2250 15245 2260
rect 15215 2230 15220 2250
rect 15240 2230 15245 2250
rect 15215 2200 15245 2230
rect 15215 2180 15220 2200
rect 15240 2180 15245 2200
rect 15215 2150 15245 2180
rect 15215 2130 15220 2150
rect 15240 2130 15245 2150
rect 15215 2100 15245 2130
rect 15215 2080 15220 2100
rect 15240 2080 15245 2100
rect 15215 2050 15245 2080
rect 15215 2030 15220 2050
rect 15240 2030 15245 2050
rect 15215 2000 15245 2030
rect 15215 1980 15220 2000
rect 15240 1980 15245 2000
rect 15215 1970 15245 1980
rect 15270 2250 15300 2260
rect 15270 2230 15275 2250
rect 15295 2230 15300 2250
rect 15270 2200 15300 2230
rect 15270 2180 15275 2200
rect 15295 2180 15300 2200
rect 15270 2150 15300 2180
rect 15270 2130 15275 2150
rect 15295 2130 15300 2150
rect 15270 2100 15300 2130
rect 15270 2080 15275 2100
rect 15295 2080 15300 2100
rect 15270 2050 15300 2080
rect 15270 2030 15275 2050
rect 15295 2030 15300 2050
rect 15270 2000 15300 2030
rect 15270 1980 15275 2000
rect 15295 1980 15300 2000
rect 15270 1970 15300 1980
rect 15325 2250 15355 2260
rect 15325 2230 15330 2250
rect 15350 2230 15355 2250
rect 15325 2200 15355 2230
rect 15325 2180 15330 2200
rect 15350 2180 15355 2200
rect 15325 2150 15355 2180
rect 15325 2130 15330 2150
rect 15350 2130 15355 2150
rect 15325 2100 15355 2130
rect 15325 2080 15330 2100
rect 15350 2080 15355 2100
rect 15325 2050 15355 2080
rect 15325 2030 15330 2050
rect 15350 2030 15355 2050
rect 15325 2000 15355 2030
rect 15325 1980 15330 2000
rect 15350 1980 15355 2000
rect 15325 1970 15355 1980
rect 15380 2250 15410 2260
rect 15380 2230 15385 2250
rect 15405 2230 15410 2250
rect 15380 2200 15410 2230
rect 15380 2180 15385 2200
rect 15405 2180 15410 2200
rect 15380 2150 15410 2180
rect 15380 2130 15385 2150
rect 15405 2130 15410 2150
rect 15380 2100 15410 2130
rect 15380 2080 15385 2100
rect 15405 2080 15410 2100
rect 15380 2050 15410 2080
rect 15380 2030 15385 2050
rect 15405 2030 15410 2050
rect 15380 2000 15410 2030
rect 15380 1980 15385 2000
rect 15405 1980 15410 2000
rect 15380 1970 15410 1980
rect 15435 2250 15465 2260
rect 15435 2230 15440 2250
rect 15460 2230 15465 2250
rect 15435 2200 15465 2230
rect 15435 2180 15440 2200
rect 15460 2180 15465 2200
rect 15435 2150 15465 2180
rect 15435 2130 15440 2150
rect 15460 2130 15465 2150
rect 15435 2100 15465 2130
rect 15435 2080 15440 2100
rect 15460 2080 15465 2100
rect 15435 2050 15465 2080
rect 15435 2030 15440 2050
rect 15460 2030 15465 2050
rect 15435 2000 15465 2030
rect 15435 1980 15440 2000
rect 15460 1980 15465 2000
rect 15435 1970 15465 1980
rect 15490 2250 15520 2260
rect 15490 2230 15495 2250
rect 15515 2230 15520 2250
rect 15490 2200 15520 2230
rect 15490 2180 15495 2200
rect 15515 2180 15520 2200
rect 15490 2150 15520 2180
rect 15490 2130 15495 2150
rect 15515 2130 15520 2150
rect 15490 2100 15520 2130
rect 15490 2080 15495 2100
rect 15515 2080 15520 2100
rect 15490 2050 15520 2080
rect 15490 2030 15495 2050
rect 15515 2030 15520 2050
rect 15490 2000 15520 2030
rect 15490 1980 15495 2000
rect 15515 1980 15520 2000
rect 15490 1970 15520 1980
rect 15545 2250 15575 2260
rect 15545 2230 15550 2250
rect 15570 2230 15575 2250
rect 15545 2200 15575 2230
rect 15545 2180 15550 2200
rect 15570 2180 15575 2200
rect 15545 2150 15575 2180
rect 15545 2130 15550 2150
rect 15570 2130 15575 2150
rect 15545 2100 15575 2130
rect 15545 2080 15550 2100
rect 15570 2080 15575 2100
rect 15545 2050 15575 2080
rect 15545 2030 15550 2050
rect 15570 2030 15575 2050
rect 15545 2000 15575 2030
rect 15545 1980 15550 2000
rect 15570 1980 15575 2000
rect 15545 1970 15575 1980
rect 15600 2250 15630 2260
rect 15600 2230 15605 2250
rect 15625 2230 15630 2250
rect 15600 2200 15630 2230
rect 15600 2180 15605 2200
rect 15625 2180 15630 2200
rect 15600 2150 15630 2180
rect 15600 2130 15605 2150
rect 15625 2130 15630 2150
rect 15600 2100 15630 2130
rect 15600 2080 15605 2100
rect 15625 2080 15630 2100
rect 15600 2050 15630 2080
rect 15600 2030 15605 2050
rect 15625 2030 15630 2050
rect 15600 2000 15630 2030
rect 15600 1980 15605 2000
rect 15625 1980 15630 2000
rect 15600 1970 15630 1980
rect 15655 2250 15685 2260
rect 15655 2230 15660 2250
rect 15680 2230 15685 2250
rect 15655 2200 15685 2230
rect 15655 2180 15660 2200
rect 15680 2180 15685 2200
rect 15655 2150 15685 2180
rect 15655 2130 15660 2150
rect 15680 2130 15685 2150
rect 15655 2100 15685 2130
rect 15655 2080 15660 2100
rect 15680 2080 15685 2100
rect 15655 2050 15685 2080
rect 15655 2030 15660 2050
rect 15680 2030 15685 2050
rect 15655 2000 15685 2030
rect 15655 1980 15660 2000
rect 15680 1980 15685 2000
rect 15655 1970 15685 1980
rect 15710 2250 15740 2260
rect 15710 2230 15715 2250
rect 15735 2230 15740 2250
rect 15710 2200 15740 2230
rect 15710 2180 15715 2200
rect 15735 2180 15740 2200
rect 15710 2150 15740 2180
rect 15710 2130 15715 2150
rect 15735 2130 15740 2150
rect 15710 2100 15740 2130
rect 15710 2080 15715 2100
rect 15735 2080 15740 2100
rect 15710 2050 15740 2080
rect 15710 2030 15715 2050
rect 15735 2030 15740 2050
rect 15710 2000 15740 2030
rect 15710 1980 15715 2000
rect 15735 1980 15740 2000
rect 15710 1970 15740 1980
rect 15765 2250 15795 2260
rect 15765 2230 15770 2250
rect 15790 2230 15795 2250
rect 15765 2200 15795 2230
rect 15765 2180 15770 2200
rect 15790 2180 15795 2200
rect 15765 2150 15795 2180
rect 15765 2130 15770 2150
rect 15790 2130 15795 2150
rect 15765 2100 15795 2130
rect 15765 2080 15770 2100
rect 15790 2080 15795 2100
rect 15765 2050 15795 2080
rect 15765 2030 15770 2050
rect 15790 2030 15795 2050
rect 15765 2000 15795 2030
rect 15765 1980 15770 2000
rect 15790 1980 15795 2000
rect 15765 1970 15795 1980
rect 15820 2250 15890 2260
rect 15820 2230 15825 2250
rect 15845 2230 15865 2250
rect 15885 2230 15890 2250
rect 15820 2200 15890 2230
rect 15820 2180 15825 2200
rect 15845 2180 15865 2200
rect 15885 2180 15890 2200
rect 17910 2250 17980 2260
rect 17910 2230 17915 2250
rect 17935 2230 17955 2250
rect 17975 2230 17980 2250
rect 17910 2200 17980 2230
rect 15820 2150 15890 2180
rect 15820 2130 15825 2150
rect 15845 2130 15865 2150
rect 15885 2130 15890 2150
rect 16330 2175 16370 2185
rect 16330 2155 16340 2175
rect 16360 2155 16370 2175
rect 16330 2145 16370 2155
rect 16440 2175 16480 2185
rect 16440 2155 16450 2175
rect 16470 2155 16480 2175
rect 16440 2145 16480 2155
rect 16550 2175 16590 2185
rect 16550 2155 16560 2175
rect 16580 2155 16590 2175
rect 16550 2145 16590 2155
rect 16660 2175 16700 2185
rect 16660 2155 16670 2175
rect 16690 2155 16700 2175
rect 16660 2145 16700 2155
rect 16770 2175 16810 2185
rect 16770 2155 16780 2175
rect 16800 2155 16810 2175
rect 16770 2145 16810 2155
rect 16828 2175 16862 2185
rect 16828 2155 16836 2175
rect 16854 2155 16862 2175
rect 16828 2145 16862 2155
rect 16880 2175 16920 2185
rect 16880 2155 16890 2175
rect 16910 2155 16920 2175
rect 16880 2145 16920 2155
rect 16990 2175 17030 2185
rect 16990 2155 17000 2175
rect 17020 2155 17030 2175
rect 16990 2145 17030 2155
rect 17100 2175 17140 2185
rect 17100 2155 17110 2175
rect 17130 2155 17140 2175
rect 17100 2145 17140 2155
rect 17210 2175 17250 2185
rect 17210 2155 17220 2175
rect 17240 2155 17250 2175
rect 17210 2145 17250 2155
rect 17320 2175 17360 2185
rect 17320 2155 17330 2175
rect 17350 2155 17360 2175
rect 17320 2145 17360 2155
rect 17430 2175 17470 2185
rect 17430 2155 17440 2175
rect 17460 2155 17470 2175
rect 17430 2145 17470 2155
rect 17910 2180 17915 2200
rect 17935 2180 17955 2200
rect 17975 2180 17980 2200
rect 17910 2150 17980 2180
rect 15820 2100 15890 2130
rect 16340 2125 16360 2145
rect 16450 2125 16470 2145
rect 16560 2125 16580 2145
rect 16670 2125 16690 2145
rect 16780 2125 16800 2145
rect 16890 2125 16910 2145
rect 17000 2125 17020 2145
rect 17110 2125 17130 2145
rect 17220 2125 17240 2145
rect 17330 2125 17350 2145
rect 17440 2125 17460 2145
rect 17910 2130 17915 2150
rect 17935 2130 17955 2150
rect 17975 2130 17980 2150
rect 15820 2080 15825 2100
rect 15845 2080 15865 2100
rect 15885 2080 15890 2100
rect 15820 2050 15890 2080
rect 15820 2030 15825 2050
rect 15845 2030 15865 2050
rect 15885 2030 15890 2050
rect 15820 2000 15890 2030
rect 15820 1980 15825 2000
rect 15845 1980 15865 2000
rect 15885 1980 15890 2000
rect 16240 2115 16310 2125
rect 16240 2095 16245 2115
rect 16265 2095 16285 2115
rect 16305 2095 16310 2115
rect 16240 2065 16310 2095
rect 16240 2045 16245 2065
rect 16265 2045 16285 2065
rect 16305 2045 16310 2065
rect 16240 2015 16310 2045
rect 16240 1995 16245 2015
rect 16265 1995 16285 2015
rect 16305 1995 16310 2015
rect 16240 1985 16310 1995
rect 16335 2115 16365 2125
rect 16335 2095 16340 2115
rect 16360 2095 16365 2115
rect 16335 2065 16365 2095
rect 16335 2045 16340 2065
rect 16360 2045 16365 2065
rect 16335 2015 16365 2045
rect 16335 1995 16340 2015
rect 16360 1995 16365 2015
rect 16335 1985 16365 1995
rect 16390 2115 16420 2125
rect 16390 2095 16395 2115
rect 16415 2095 16420 2115
rect 16390 2065 16420 2095
rect 16390 2045 16395 2065
rect 16415 2045 16420 2065
rect 16390 2015 16420 2045
rect 16390 1995 16395 2015
rect 16415 1995 16420 2015
rect 16390 1985 16420 1995
rect 16445 2115 16475 2125
rect 16445 2095 16450 2115
rect 16470 2095 16475 2115
rect 16445 2065 16475 2095
rect 16445 2045 16450 2065
rect 16470 2045 16475 2065
rect 16445 2015 16475 2045
rect 16445 1995 16450 2015
rect 16470 1995 16475 2015
rect 16445 1985 16475 1995
rect 16500 2115 16530 2125
rect 16500 2095 16505 2115
rect 16525 2095 16530 2115
rect 16500 2065 16530 2095
rect 16500 2045 16505 2065
rect 16525 2045 16530 2065
rect 16500 2015 16530 2045
rect 16500 1995 16505 2015
rect 16525 1995 16530 2015
rect 16500 1985 16530 1995
rect 16555 2115 16585 2125
rect 16555 2095 16560 2115
rect 16580 2095 16585 2115
rect 16555 2065 16585 2095
rect 16555 2045 16560 2065
rect 16580 2045 16585 2065
rect 16555 2015 16585 2045
rect 16555 1995 16560 2015
rect 16580 1995 16585 2015
rect 16555 1985 16585 1995
rect 16610 2115 16640 2125
rect 16610 2095 16615 2115
rect 16635 2095 16640 2115
rect 16610 2065 16640 2095
rect 16610 2045 16615 2065
rect 16635 2045 16640 2065
rect 16610 2015 16640 2045
rect 16610 1995 16615 2015
rect 16635 1995 16640 2015
rect 16610 1985 16640 1995
rect 16665 2115 16695 2125
rect 16665 2095 16670 2115
rect 16690 2095 16695 2115
rect 16665 2065 16695 2095
rect 16665 2045 16670 2065
rect 16690 2045 16695 2065
rect 16665 2015 16695 2045
rect 16665 1995 16670 2015
rect 16690 1995 16695 2015
rect 16665 1985 16695 1995
rect 16720 2115 16750 2125
rect 16720 2095 16725 2115
rect 16745 2095 16750 2115
rect 16720 2065 16750 2095
rect 16720 2045 16725 2065
rect 16745 2045 16750 2065
rect 16720 2015 16750 2045
rect 16720 1995 16725 2015
rect 16745 1995 16750 2015
rect 16720 1985 16750 1995
rect 16775 2115 16805 2125
rect 16775 2095 16780 2115
rect 16800 2095 16805 2115
rect 16775 2065 16805 2095
rect 16775 2045 16780 2065
rect 16800 2045 16805 2065
rect 16775 2015 16805 2045
rect 16775 1995 16780 2015
rect 16800 1995 16805 2015
rect 16775 1985 16805 1995
rect 16830 2115 16860 2125
rect 16830 2095 16835 2115
rect 16855 2095 16860 2115
rect 16830 2065 16860 2095
rect 16830 2045 16835 2065
rect 16855 2045 16860 2065
rect 16830 2015 16860 2045
rect 16830 1995 16835 2015
rect 16855 1995 16860 2015
rect 16830 1985 16860 1995
rect 16885 2115 16915 2125
rect 16885 2095 16890 2115
rect 16910 2095 16915 2115
rect 16885 2065 16915 2095
rect 16885 2045 16890 2065
rect 16910 2045 16915 2065
rect 16885 2015 16915 2045
rect 16885 1995 16890 2015
rect 16910 1995 16915 2015
rect 16885 1985 16915 1995
rect 16940 2115 16970 2125
rect 16940 2095 16945 2115
rect 16965 2095 16970 2115
rect 16940 2065 16970 2095
rect 16940 2045 16945 2065
rect 16965 2045 16970 2065
rect 16940 2015 16970 2045
rect 16940 1995 16945 2015
rect 16965 1995 16970 2015
rect 16940 1985 16970 1995
rect 16995 2115 17025 2125
rect 16995 2095 17000 2115
rect 17020 2095 17025 2115
rect 16995 2065 17025 2095
rect 16995 2045 17000 2065
rect 17020 2045 17025 2065
rect 16995 2015 17025 2045
rect 16995 1995 17000 2015
rect 17020 1995 17025 2015
rect 16995 1985 17025 1995
rect 17050 2115 17080 2125
rect 17050 2095 17055 2115
rect 17075 2095 17080 2115
rect 17050 2065 17080 2095
rect 17050 2045 17055 2065
rect 17075 2045 17080 2065
rect 17050 2015 17080 2045
rect 17050 1995 17055 2015
rect 17075 1995 17080 2015
rect 17050 1985 17080 1995
rect 17105 2115 17135 2125
rect 17105 2095 17110 2115
rect 17130 2095 17135 2115
rect 17105 2065 17135 2095
rect 17105 2045 17110 2065
rect 17130 2045 17135 2065
rect 17105 2015 17135 2045
rect 17105 1995 17110 2015
rect 17130 1995 17135 2015
rect 17105 1985 17135 1995
rect 17160 2115 17190 2125
rect 17160 2095 17165 2115
rect 17185 2095 17190 2115
rect 17160 2065 17190 2095
rect 17160 2045 17165 2065
rect 17185 2045 17190 2065
rect 17160 2015 17190 2045
rect 17160 1995 17165 2015
rect 17185 1995 17190 2015
rect 17160 1985 17190 1995
rect 17215 2115 17245 2125
rect 17215 2095 17220 2115
rect 17240 2095 17245 2115
rect 17215 2065 17245 2095
rect 17215 2045 17220 2065
rect 17240 2045 17245 2065
rect 17215 2015 17245 2045
rect 17215 1995 17220 2015
rect 17240 1995 17245 2015
rect 17215 1985 17245 1995
rect 17270 2115 17300 2125
rect 17270 2095 17275 2115
rect 17295 2095 17300 2115
rect 17270 2065 17300 2095
rect 17270 2045 17275 2065
rect 17295 2045 17300 2065
rect 17270 2015 17300 2045
rect 17270 1995 17275 2015
rect 17295 1995 17300 2015
rect 17270 1985 17300 1995
rect 17325 2115 17355 2125
rect 17325 2095 17330 2115
rect 17350 2095 17355 2115
rect 17325 2065 17355 2095
rect 17325 2045 17330 2065
rect 17350 2045 17355 2065
rect 17325 2015 17355 2045
rect 17325 1995 17330 2015
rect 17350 1995 17355 2015
rect 17325 1985 17355 1995
rect 17380 2115 17410 2125
rect 17380 2095 17385 2115
rect 17405 2095 17410 2115
rect 17380 2065 17410 2095
rect 17380 2045 17385 2065
rect 17405 2045 17410 2065
rect 17380 2015 17410 2045
rect 17380 1995 17385 2015
rect 17405 1995 17410 2015
rect 17380 1985 17410 1995
rect 17435 2115 17465 2125
rect 17435 2095 17440 2115
rect 17460 2095 17465 2115
rect 17435 2065 17465 2095
rect 17435 2045 17440 2065
rect 17460 2045 17465 2065
rect 17435 2015 17465 2045
rect 17435 1995 17440 2015
rect 17460 1995 17465 2015
rect 17435 1985 17465 1995
rect 17490 2115 17560 2125
rect 17490 2095 17495 2115
rect 17515 2095 17535 2115
rect 17555 2095 17560 2115
rect 17490 2065 17560 2095
rect 17490 2045 17495 2065
rect 17515 2045 17535 2065
rect 17555 2045 17560 2065
rect 17490 2015 17560 2045
rect 17490 1995 17495 2015
rect 17515 1995 17535 2015
rect 17555 1995 17560 2015
rect 17490 1985 17560 1995
rect 17910 2100 17980 2130
rect 17910 2080 17915 2100
rect 17935 2080 17955 2100
rect 17975 2080 17980 2100
rect 17910 2050 17980 2080
rect 17910 2030 17915 2050
rect 17935 2030 17955 2050
rect 17975 2030 17980 2050
rect 17910 2000 17980 2030
rect 15820 1970 15890 1980
rect 5230 1935 5260 1965
rect 15220 1950 15240 1970
rect 15330 1950 15350 1970
rect 15440 1950 15460 1970
rect 15550 1950 15570 1970
rect 15660 1950 15680 1970
rect 15770 1950 15790 1970
rect 16245 1965 16265 1985
rect 16395 1965 16415 1985
rect 16505 1965 16525 1985
rect 16615 1965 16635 1985
rect 16725 1965 16745 1985
rect 16835 1965 16855 1985
rect 16945 1965 16965 1985
rect 17055 1965 17075 1985
rect 17165 1965 17185 1985
rect 17275 1965 17295 1985
rect 17385 1965 17405 1985
rect 17535 1965 17555 1985
rect 17910 1980 17915 2000
rect 17935 1980 17955 2000
rect 17975 1980 17980 2000
rect 17910 1970 17980 1980
rect 18005 2250 18035 2260
rect 18005 2230 18010 2250
rect 18030 2230 18035 2250
rect 18005 2200 18035 2230
rect 18005 2180 18010 2200
rect 18030 2180 18035 2200
rect 18005 2150 18035 2180
rect 18005 2130 18010 2150
rect 18030 2130 18035 2150
rect 18005 2100 18035 2130
rect 18005 2080 18010 2100
rect 18030 2080 18035 2100
rect 18005 2050 18035 2080
rect 18005 2030 18010 2050
rect 18030 2030 18035 2050
rect 18005 2000 18035 2030
rect 18005 1980 18010 2000
rect 18030 1980 18035 2000
rect 18005 1970 18035 1980
rect 18060 2250 18090 2260
rect 18060 2230 18065 2250
rect 18085 2230 18090 2250
rect 18060 2200 18090 2230
rect 18060 2180 18065 2200
rect 18085 2180 18090 2200
rect 18060 2150 18090 2180
rect 18060 2130 18065 2150
rect 18085 2130 18090 2150
rect 18060 2100 18090 2130
rect 18060 2080 18065 2100
rect 18085 2080 18090 2100
rect 18060 2050 18090 2080
rect 18060 2030 18065 2050
rect 18085 2030 18090 2050
rect 18060 2000 18090 2030
rect 18060 1980 18065 2000
rect 18085 1980 18090 2000
rect 18060 1970 18090 1980
rect 18115 2250 18145 2260
rect 18115 2230 18120 2250
rect 18140 2230 18145 2250
rect 18115 2200 18145 2230
rect 18115 2180 18120 2200
rect 18140 2180 18145 2200
rect 18115 2150 18145 2180
rect 18115 2130 18120 2150
rect 18140 2130 18145 2150
rect 18115 2100 18145 2130
rect 18115 2080 18120 2100
rect 18140 2080 18145 2100
rect 18115 2050 18145 2080
rect 18115 2030 18120 2050
rect 18140 2030 18145 2050
rect 18115 2000 18145 2030
rect 18115 1980 18120 2000
rect 18140 1980 18145 2000
rect 18115 1970 18145 1980
rect 18170 2250 18200 2260
rect 18170 2230 18175 2250
rect 18195 2230 18200 2250
rect 18170 2200 18200 2230
rect 18170 2180 18175 2200
rect 18195 2180 18200 2200
rect 18170 2150 18200 2180
rect 18170 2130 18175 2150
rect 18195 2130 18200 2150
rect 18170 2100 18200 2130
rect 18170 2080 18175 2100
rect 18195 2080 18200 2100
rect 18170 2050 18200 2080
rect 18170 2030 18175 2050
rect 18195 2030 18200 2050
rect 18170 2000 18200 2030
rect 18170 1980 18175 2000
rect 18195 1980 18200 2000
rect 18170 1970 18200 1980
rect 18225 2250 18255 2260
rect 18225 2230 18230 2250
rect 18250 2230 18255 2250
rect 18225 2200 18255 2230
rect 18225 2180 18230 2200
rect 18250 2180 18255 2200
rect 18225 2150 18255 2180
rect 18225 2130 18230 2150
rect 18250 2130 18255 2150
rect 18225 2100 18255 2130
rect 18225 2080 18230 2100
rect 18250 2080 18255 2100
rect 18225 2050 18255 2080
rect 18225 2030 18230 2050
rect 18250 2030 18255 2050
rect 18225 2000 18255 2030
rect 18225 1980 18230 2000
rect 18250 1980 18255 2000
rect 18225 1970 18255 1980
rect 18280 2250 18310 2260
rect 18280 2230 18285 2250
rect 18305 2230 18310 2250
rect 18280 2200 18310 2230
rect 18280 2180 18285 2200
rect 18305 2180 18310 2200
rect 18280 2150 18310 2180
rect 18280 2130 18285 2150
rect 18305 2130 18310 2150
rect 18280 2100 18310 2130
rect 18280 2080 18285 2100
rect 18305 2080 18310 2100
rect 18280 2050 18310 2080
rect 18280 2030 18285 2050
rect 18305 2030 18310 2050
rect 18280 2000 18310 2030
rect 18280 1980 18285 2000
rect 18305 1980 18310 2000
rect 18280 1970 18310 1980
rect 18335 2250 18365 2260
rect 18335 2230 18340 2250
rect 18360 2230 18365 2250
rect 18335 2200 18365 2230
rect 18335 2180 18340 2200
rect 18360 2180 18365 2200
rect 18335 2150 18365 2180
rect 18335 2130 18340 2150
rect 18360 2130 18365 2150
rect 18335 2100 18365 2130
rect 18335 2080 18340 2100
rect 18360 2080 18365 2100
rect 18335 2050 18365 2080
rect 18335 2030 18340 2050
rect 18360 2030 18365 2050
rect 18335 2000 18365 2030
rect 18335 1980 18340 2000
rect 18360 1980 18365 2000
rect 18335 1970 18365 1980
rect 18390 2250 18420 2260
rect 18390 2230 18395 2250
rect 18415 2230 18420 2250
rect 18390 2200 18420 2230
rect 18390 2180 18395 2200
rect 18415 2180 18420 2200
rect 18390 2150 18420 2180
rect 18390 2130 18395 2150
rect 18415 2130 18420 2150
rect 18390 2100 18420 2130
rect 18390 2080 18395 2100
rect 18415 2080 18420 2100
rect 18390 2050 18420 2080
rect 18390 2030 18395 2050
rect 18415 2030 18420 2050
rect 18390 2000 18420 2030
rect 18390 1980 18395 2000
rect 18415 1980 18420 2000
rect 18390 1970 18420 1980
rect 18445 2250 18475 2260
rect 18445 2230 18450 2250
rect 18470 2230 18475 2250
rect 18445 2200 18475 2230
rect 18445 2180 18450 2200
rect 18470 2180 18475 2200
rect 18445 2150 18475 2180
rect 18445 2130 18450 2150
rect 18470 2130 18475 2150
rect 18445 2100 18475 2130
rect 18445 2080 18450 2100
rect 18470 2080 18475 2100
rect 18445 2050 18475 2080
rect 18445 2030 18450 2050
rect 18470 2030 18475 2050
rect 18445 2000 18475 2030
rect 18445 1980 18450 2000
rect 18470 1980 18475 2000
rect 18445 1970 18475 1980
rect 18500 2250 18530 2260
rect 18500 2230 18505 2250
rect 18525 2230 18530 2250
rect 18500 2200 18530 2230
rect 18500 2180 18505 2200
rect 18525 2180 18530 2200
rect 18500 2150 18530 2180
rect 18500 2130 18505 2150
rect 18525 2130 18530 2150
rect 18500 2100 18530 2130
rect 18500 2080 18505 2100
rect 18525 2080 18530 2100
rect 18500 2050 18530 2080
rect 18500 2030 18505 2050
rect 18525 2030 18530 2050
rect 18500 2000 18530 2030
rect 18500 1980 18505 2000
rect 18525 1980 18530 2000
rect 18500 1970 18530 1980
rect 18555 2250 18585 2260
rect 18555 2230 18560 2250
rect 18580 2230 18585 2250
rect 18555 2200 18585 2230
rect 18555 2180 18560 2200
rect 18580 2180 18585 2200
rect 18555 2150 18585 2180
rect 18555 2130 18560 2150
rect 18580 2130 18585 2150
rect 18555 2100 18585 2130
rect 18555 2080 18560 2100
rect 18580 2080 18585 2100
rect 18555 2050 18585 2080
rect 18555 2030 18560 2050
rect 18580 2030 18585 2050
rect 18555 2000 18585 2030
rect 18555 1980 18560 2000
rect 18580 1980 18585 2000
rect 18555 1970 18585 1980
rect 18610 2250 18680 2260
rect 18610 2230 18615 2250
rect 18635 2230 18655 2250
rect 18675 2230 18680 2250
rect 18610 2200 18680 2230
rect 18610 2180 18615 2200
rect 18635 2180 18655 2200
rect 18675 2180 18680 2200
rect 18610 2150 18680 2180
rect 18610 2130 18615 2150
rect 18635 2130 18655 2150
rect 18675 2130 18680 2150
rect 18610 2100 18680 2130
rect 18610 2080 18615 2100
rect 18635 2080 18655 2100
rect 18675 2080 18680 2100
rect 18610 2050 18680 2080
rect 18610 2030 18615 2050
rect 18635 2030 18655 2050
rect 18675 2030 18680 2050
rect 18610 2000 18680 2030
rect 18610 1980 18615 2000
rect 18635 1980 18655 2000
rect 18675 1980 18680 2000
rect 18610 1970 18680 1980
rect 18795 2000 18830 2010
rect 18795 1975 18800 2000
rect 18825 1975 18830 2000
rect 16235 1955 16275 1965
rect 5230 1915 5235 1935
rect 5255 1915 5260 1935
rect 5230 1905 5260 1915
rect 15210 1940 15250 1950
rect 15210 1920 15220 1940
rect 15238 1920 15250 1940
rect 15210 1910 15250 1920
rect 15320 1940 15360 1950
rect 15320 1920 15330 1940
rect 15348 1920 15360 1940
rect 15320 1910 15360 1920
rect 15430 1940 15470 1950
rect 15430 1920 15440 1940
rect 15458 1920 15470 1940
rect 15430 1910 15470 1920
rect 15540 1940 15580 1950
rect 15540 1920 15550 1940
rect 15568 1920 15580 1940
rect 15540 1910 15580 1920
rect 15650 1940 15690 1950
rect 15650 1920 15660 1940
rect 15678 1920 15690 1940
rect 15650 1910 15690 1920
rect 15760 1940 15800 1950
rect 15760 1920 15770 1940
rect 15788 1920 15800 1940
rect 16235 1935 16245 1955
rect 16265 1935 16275 1955
rect 16235 1925 16275 1935
rect 16385 1955 16425 1965
rect 16385 1935 16395 1955
rect 16415 1935 16425 1955
rect 16385 1925 16425 1935
rect 16495 1955 16535 1965
rect 16495 1935 16505 1955
rect 16525 1935 16535 1955
rect 16495 1925 16535 1935
rect 16605 1955 16645 1965
rect 16605 1935 16615 1955
rect 16635 1935 16645 1955
rect 16605 1925 16645 1935
rect 16715 1955 16755 1965
rect 16715 1935 16725 1955
rect 16745 1935 16755 1955
rect 16715 1925 16755 1935
rect 16825 1955 16865 1965
rect 16825 1935 16835 1955
rect 16855 1935 16865 1955
rect 16825 1925 16865 1935
rect 16935 1955 16975 1965
rect 16935 1935 16945 1955
rect 16965 1935 16975 1955
rect 16935 1925 16975 1935
rect 17045 1955 17085 1965
rect 17045 1935 17055 1955
rect 17075 1935 17085 1955
rect 17045 1925 17085 1935
rect 17155 1955 17195 1965
rect 17155 1935 17165 1955
rect 17185 1935 17195 1955
rect 17155 1925 17195 1935
rect 17265 1955 17305 1965
rect 17265 1935 17275 1955
rect 17295 1935 17305 1955
rect 17265 1925 17305 1935
rect 17375 1955 17415 1965
rect 17375 1935 17385 1955
rect 17405 1935 17415 1955
rect 17375 1925 17415 1935
rect 17525 1955 17565 1965
rect 17525 1935 17535 1955
rect 17555 1935 17565 1955
rect 18010 1950 18030 1970
rect 18120 1950 18140 1970
rect 18230 1950 18250 1970
rect 18340 1950 18360 1970
rect 18450 1950 18470 1970
rect 18560 1950 18580 1970
rect 18795 1965 18830 1975
rect 18855 2000 18890 2010
rect 18855 1975 18860 2000
rect 18885 1975 18890 2000
rect 18855 1965 18890 1975
rect 18915 2000 18950 2010
rect 18915 1975 18920 2000
rect 18945 1975 18950 2000
rect 18915 1965 18950 1975
rect 18975 2000 19010 2010
rect 18975 1975 18980 2000
rect 19005 1975 19010 2000
rect 18975 1965 19010 1975
rect 17525 1925 17565 1935
rect 18000 1940 18040 1950
rect 15760 1910 15800 1920
rect 18000 1920 18012 1940
rect 18030 1920 18040 1940
rect 18000 1910 18040 1920
rect 18110 1940 18150 1950
rect 18110 1920 18122 1940
rect 18140 1920 18150 1940
rect 18110 1910 18150 1920
rect 18220 1940 18260 1950
rect 18220 1920 18232 1940
rect 18250 1920 18260 1940
rect 18220 1910 18260 1920
rect 18330 1940 18370 1950
rect 18330 1920 18342 1940
rect 18360 1920 18370 1940
rect 18330 1910 18370 1920
rect 18440 1940 18480 1950
rect 18440 1920 18452 1940
rect 18470 1920 18480 1940
rect 18440 1910 18480 1920
rect 18550 1940 18590 1950
rect 18550 1920 18562 1940
rect 18580 1920 18590 1940
rect 18550 1910 18590 1920
rect 2575 1885 2595 1905
rect 2685 1885 2705 1905
rect 2755 1885 2775 1905
rect 2935 1885 2955 1905
rect 3055 1885 3075 1905
rect 3295 1885 3315 1905
rect 3415 1885 3435 1905
rect 3655 1885 3675 1905
rect 3775 1885 3795 1905
rect 2565 1875 2600 1885
rect 2565 1855 2575 1875
rect 2595 1855 2600 1875
rect 2565 1845 2600 1855
rect 2620 1875 2660 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2680 1875 2715 1885
rect 2680 1855 2685 1875
rect 2705 1855 2715 1875
rect 2680 1845 2715 1855
rect 2755 1875 2805 1885
rect 2755 1855 2775 1875
rect 2795 1855 2805 1875
rect 2755 1845 2805 1855
rect 2835 1875 2875 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1875 2965 1885
rect 2925 1855 2935 1875
rect 2955 1855 2965 1875
rect 2925 1845 2965 1855
rect 3045 1875 3085 1885
rect 3045 1855 3055 1875
rect 3075 1855 3085 1875
rect 3045 1845 3085 1855
rect 3165 1875 3205 1885
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1875 3325 1885
rect 3285 1855 3295 1875
rect 3315 1855 3325 1875
rect 3285 1845 3325 1855
rect 3405 1875 3445 1885
rect 3405 1855 3415 1875
rect 3435 1855 3445 1875
rect 3405 1845 3445 1855
rect 3525 1875 3565 1885
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1875 3685 1885
rect 3645 1855 3655 1875
rect 3675 1855 3685 1875
rect 3645 1845 3685 1855
rect 3765 1875 3805 1885
rect 3765 1855 3775 1875
rect 3795 1855 3805 1875
rect 3765 1845 3805 1855
rect 3855 1875 3895 1885
rect 3995 1880 4015 1905
rect 4215 1885 4235 1905
rect 4335 1885 4355 1905
rect 4575 1885 4595 1905
rect 4695 1885 4715 1905
rect 4935 1885 4955 1905
rect 5055 1885 5075 1905
rect 5235 1885 5255 1905
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 3985 1870 4025 1880
rect 3985 1850 3995 1870
rect 4015 1850 4025 1870
rect 3985 1840 4025 1850
rect 4115 1875 4155 1885
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4205 1875 4245 1885
rect 4205 1855 4215 1875
rect 4235 1855 4245 1875
rect 4205 1845 4245 1855
rect 4325 1875 4365 1885
rect 4325 1855 4335 1875
rect 4355 1855 4365 1875
rect 4325 1845 4365 1855
rect 4445 1875 4485 1885
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4565 1875 4605 1885
rect 4565 1855 4575 1875
rect 4595 1855 4605 1875
rect 4565 1845 4605 1855
rect 4685 1875 4725 1885
rect 4685 1855 4695 1875
rect 4715 1855 4725 1875
rect 4685 1845 4725 1855
rect 4805 1875 4845 1885
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 4925 1875 4965 1885
rect 4925 1855 4935 1875
rect 4955 1855 4965 1875
rect 4925 1845 4965 1855
rect 5045 1875 5085 1885
rect 5045 1855 5055 1875
rect 5075 1855 5085 1875
rect 5045 1845 5085 1855
rect 5135 1875 5175 1885
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 5205 1875 5255 1885
rect 5205 1855 5215 1875
rect 5235 1855 5255 1875
rect 5205 1845 5255 1855
rect 2475 1790 2505 1820
rect 2835 1785 2875 1825
rect 3045 1815 3085 1825
rect 3045 1795 3055 1815
rect 3075 1795 3085 1815
rect 3045 1785 3085 1795
rect 3165 1785 3205 1825
rect 3405 1815 3445 1825
rect 3405 1795 3415 1815
rect 3435 1795 3445 1815
rect 3405 1785 3445 1795
rect 3525 1785 3565 1825
rect 3765 1815 3805 1825
rect 3765 1795 3775 1815
rect 3795 1795 3805 1815
rect 3765 1785 3805 1795
rect 3855 1785 3895 1825
rect 4115 1785 4155 1825
rect 4205 1815 4245 1825
rect 4205 1795 4215 1815
rect 4235 1795 4245 1815
rect 4205 1785 4245 1795
rect 4445 1785 4485 1825
rect 4565 1815 4605 1825
rect 4565 1795 4575 1815
rect 4595 1795 4605 1815
rect 4565 1785 4605 1795
rect 4805 1785 4845 1825
rect 4925 1815 4965 1825
rect 4925 1795 4935 1815
rect 4955 1795 4965 1815
rect 4925 1785 4965 1795
rect 5135 1785 5175 1825
rect 5365 1790 5395 1820
rect 16190 1770 16230 1780
rect 2430 1730 2460 1760
rect 2570 1730 2600 1760
rect 2680 1730 2710 1760
rect 2805 1735 2835 1765
rect 3225 1755 3265 1765
rect 3225 1735 3235 1755
rect 3255 1735 3265 1755
rect 3225 1725 3265 1735
rect 3285 1755 3325 1765
rect 3285 1735 3295 1755
rect 3315 1735 3325 1755
rect 3285 1725 3325 1735
rect 3525 1755 3565 1765
rect 3525 1735 3535 1755
rect 3555 1735 3565 1755
rect 3525 1725 3565 1735
rect 3765 1755 3805 1765
rect 3765 1735 3775 1755
rect 3795 1735 3805 1755
rect 3765 1725 3805 1735
rect 4205 1755 4245 1765
rect 4205 1735 4215 1755
rect 4235 1735 4245 1755
rect 4205 1725 4245 1735
rect 4445 1755 4485 1765
rect 4445 1735 4455 1755
rect 4475 1735 4485 1755
rect 4445 1725 4485 1735
rect 4685 1755 4725 1765
rect 4685 1735 4695 1755
rect 4715 1735 4725 1755
rect 4685 1725 4725 1735
rect 4745 1755 4785 1765
rect 4745 1735 4755 1755
rect 4775 1735 4785 1755
rect 4745 1725 4785 1735
rect 5275 1730 5305 1760
rect 16085 1755 16125 1765
rect 16085 1735 16095 1755
rect 16115 1735 16125 1755
rect 16190 1750 16200 1770
rect 16220 1750 16230 1770
rect 16410 1770 16450 1780
rect 16190 1740 16230 1750
rect 16305 1755 16345 1765
rect 16085 1725 16125 1735
rect 3165 1710 3205 1720
rect 2805 1680 2835 1710
rect 3165 1690 3175 1710
rect 3195 1690 3205 1710
rect 3165 1680 3205 1690
rect 2385 1635 2415 1665
rect 2625 1635 2655 1665
rect 3175 1660 3195 1680
rect 3295 1660 3315 1725
rect 3405 1710 3445 1720
rect 3405 1690 3415 1710
rect 3435 1690 3445 1710
rect 3405 1680 3445 1690
rect 3415 1660 3435 1680
rect 3535 1660 3555 1725
rect 3645 1710 3685 1720
rect 3645 1690 3655 1710
rect 3675 1690 3685 1710
rect 3645 1680 3685 1690
rect 3655 1660 3675 1680
rect 3775 1660 3795 1725
rect 4215 1660 4235 1725
rect 4325 1710 4365 1720
rect 4325 1690 4335 1710
rect 4355 1690 4365 1710
rect 4325 1680 4365 1690
rect 4335 1660 4355 1680
rect 4455 1660 4475 1725
rect 4565 1710 4605 1720
rect 4565 1690 4575 1710
rect 4595 1690 4605 1710
rect 4565 1680 4605 1690
rect 4575 1660 4595 1680
rect 4695 1660 4715 1725
rect 4805 1710 4845 1720
rect 4805 1690 4815 1710
rect 4835 1690 4845 1710
rect 4805 1680 4845 1690
rect 15255 1700 15295 1710
rect 15255 1680 15265 1700
rect 15285 1680 15295 1700
rect 4815 1660 4835 1680
rect 15255 1670 15295 1680
rect 15455 1700 15495 1710
rect 15455 1680 15465 1700
rect 15485 1680 15495 1700
rect 15455 1670 15495 1680
rect 15558 1700 15592 1710
rect 15558 1680 15566 1700
rect 15584 1680 15592 1700
rect 15558 1670 15592 1680
rect 15655 1700 15695 1710
rect 15655 1680 15665 1700
rect 15685 1680 15695 1700
rect 15655 1670 15695 1680
rect 3170 1650 3200 1660
rect 3170 1630 3175 1650
rect 3195 1630 3200 1650
rect 3170 1620 3200 1630
rect 3230 1650 3260 1660
rect 3230 1630 3235 1650
rect 3255 1630 3260 1650
rect 3230 1620 3260 1630
rect 3290 1650 3320 1660
rect 3290 1630 3295 1650
rect 3315 1630 3320 1650
rect 3290 1620 3320 1630
rect 3350 1650 3380 1660
rect 3350 1630 3355 1650
rect 3375 1630 3380 1650
rect 3350 1620 3380 1630
rect 3410 1650 3440 1660
rect 3410 1630 3415 1650
rect 3435 1630 3440 1650
rect 3410 1620 3440 1630
rect 3470 1650 3500 1660
rect 3470 1630 3475 1650
rect 3495 1630 3500 1650
rect 3470 1620 3500 1630
rect 3530 1650 3560 1660
rect 3530 1630 3535 1650
rect 3555 1630 3560 1650
rect 3530 1620 3560 1630
rect 3590 1650 3620 1660
rect 3590 1630 3595 1650
rect 3615 1630 3620 1650
rect 3590 1620 3620 1630
rect 3650 1650 3680 1660
rect 3650 1630 3655 1650
rect 3675 1630 3680 1650
rect 3650 1620 3680 1630
rect 3710 1650 3740 1660
rect 3710 1630 3715 1650
rect 3735 1630 3740 1650
rect 3710 1620 3740 1630
rect 3770 1650 3800 1660
rect 3770 1630 3775 1650
rect 3795 1630 3800 1650
rect 3770 1620 3800 1630
rect 3985 1650 4025 1660
rect 3985 1630 3995 1650
rect 4015 1630 4025 1650
rect 3985 1620 4025 1630
rect 4210 1650 4240 1660
rect 4210 1630 4215 1650
rect 4235 1630 4240 1650
rect 4210 1620 4240 1630
rect 4270 1650 4300 1660
rect 4270 1630 4275 1650
rect 4295 1630 4300 1650
rect 4270 1620 4300 1630
rect 4330 1650 4360 1660
rect 4330 1630 4335 1650
rect 4355 1630 4360 1650
rect 4330 1620 4360 1630
rect 4390 1650 4420 1660
rect 4390 1630 4395 1650
rect 4415 1630 4420 1650
rect 4390 1620 4420 1630
rect 4450 1650 4480 1660
rect 4450 1630 4455 1650
rect 4475 1630 4480 1650
rect 4450 1620 4480 1630
rect 4510 1650 4540 1660
rect 4510 1630 4515 1650
rect 4535 1630 4540 1650
rect 4510 1620 4540 1630
rect 4570 1650 4600 1660
rect 4570 1630 4575 1650
rect 4595 1630 4600 1650
rect 4570 1620 4600 1630
rect 4630 1650 4660 1660
rect 4630 1630 4635 1650
rect 4655 1630 4660 1650
rect 4630 1620 4660 1630
rect 4690 1650 4720 1660
rect 4690 1630 4695 1650
rect 4715 1630 4720 1650
rect 4690 1620 4720 1630
rect 4750 1650 4780 1660
rect 4750 1630 4755 1650
rect 4775 1630 4780 1650
rect 4750 1620 4780 1630
rect 4810 1650 4840 1660
rect 15265 1650 15285 1670
rect 15465 1650 15485 1670
rect 15665 1650 15685 1670
rect 16095 1660 16115 1725
rect 16200 1660 16220 1740
rect 16305 1735 16315 1755
rect 16335 1735 16345 1755
rect 16410 1750 16420 1770
rect 16440 1750 16450 1770
rect 16640 1770 16680 1780
rect 16410 1740 16450 1750
rect 16525 1755 16565 1765
rect 16305 1725 16345 1735
rect 16237 1710 16269 1720
rect 16237 1690 16243 1710
rect 16260 1690 16269 1710
rect 16237 1680 16269 1690
rect 16315 1660 16335 1725
rect 16420 1660 16440 1740
rect 16525 1735 16535 1755
rect 16555 1735 16565 1755
rect 16640 1750 16650 1770
rect 16670 1750 16680 1770
rect 17230 1770 17270 1780
rect 16640 1740 16680 1750
rect 17125 1755 17165 1765
rect 16525 1725 16565 1735
rect 16457 1710 16489 1720
rect 16457 1690 16463 1710
rect 16480 1690 16489 1710
rect 16457 1680 16489 1690
rect 16535 1660 16555 1725
rect 16601 1710 16633 1720
rect 16601 1690 16610 1710
rect 16627 1690 16633 1710
rect 16601 1680 16633 1690
rect 16650 1660 16670 1740
rect 17125 1735 17135 1755
rect 17155 1735 17165 1755
rect 17230 1750 17240 1770
rect 17260 1750 17270 1770
rect 17450 1770 17490 1780
rect 17230 1740 17270 1750
rect 17345 1755 17385 1765
rect 17125 1725 17165 1735
rect 16820 1710 16850 1720
rect 16820 1690 16825 1710
rect 16845 1690 16850 1710
rect 16820 1680 16850 1690
rect 16867 1710 16899 1720
rect 16867 1690 16876 1710
rect 16893 1690 16899 1710
rect 16867 1680 16899 1690
rect 16950 1710 16980 1720
rect 16950 1690 16955 1710
rect 16975 1690 16980 1710
rect 16950 1680 16980 1690
rect 16830 1660 16850 1680
rect 16950 1660 16970 1680
rect 17135 1660 17155 1725
rect 17240 1660 17260 1740
rect 17345 1735 17355 1755
rect 17375 1735 17385 1755
rect 17450 1750 17460 1770
rect 17480 1750 17490 1770
rect 17680 1770 17720 1780
rect 17450 1740 17490 1750
rect 17565 1755 17605 1765
rect 17345 1725 17385 1735
rect 17277 1710 17309 1720
rect 17277 1690 17283 1710
rect 17300 1690 17309 1710
rect 17277 1680 17309 1690
rect 17355 1660 17375 1725
rect 17460 1660 17480 1740
rect 17565 1735 17575 1755
rect 17595 1735 17605 1755
rect 17680 1750 17690 1770
rect 17710 1750 17720 1770
rect 17680 1740 17720 1750
rect 17565 1725 17605 1735
rect 17497 1710 17529 1720
rect 17497 1690 17503 1710
rect 17520 1690 17529 1710
rect 17497 1680 17529 1690
rect 17575 1660 17595 1725
rect 17641 1710 17673 1720
rect 17641 1690 17650 1710
rect 17667 1690 17673 1710
rect 17641 1680 17673 1690
rect 17690 1660 17710 1740
rect 18105 1700 18145 1710
rect 18105 1680 18115 1700
rect 18135 1680 18145 1700
rect 18105 1670 18145 1680
rect 18208 1700 18242 1710
rect 18208 1680 18216 1700
rect 18234 1680 18242 1700
rect 18208 1670 18242 1680
rect 18305 1700 18345 1710
rect 18305 1680 18315 1700
rect 18335 1680 18345 1700
rect 18305 1670 18345 1680
rect 18505 1700 18545 1710
rect 18505 1680 18515 1700
rect 18535 1680 18545 1700
rect 18505 1670 18545 1680
rect 15990 1650 16065 1660
rect 4810 1630 4815 1650
rect 4835 1630 4840 1650
rect 4810 1620 4840 1630
rect 14970 1640 15005 1650
rect 2335 1565 2365 1595
rect 3165 1590 3205 1600
rect 3165 1570 3175 1590
rect 3195 1570 3205 1590
rect 3165 1560 3205 1570
rect 3235 1550 3255 1620
rect 3355 1550 3375 1620
rect 3475 1550 3495 1620
rect 3595 1550 3615 1620
rect 3715 1550 3735 1620
rect 4275 1550 4295 1620
rect 4395 1550 4415 1620
rect 4515 1550 4535 1620
rect 4635 1550 4655 1620
rect 4755 1550 4775 1620
rect 14970 1615 14975 1640
rect 15000 1615 15005 1640
rect 14970 1605 15005 1615
rect 4805 1590 4845 1600
rect 4805 1570 4815 1590
rect 4835 1570 4845 1590
rect 4805 1560 4845 1570
rect 5415 1565 5445 1595
rect 3225 1540 3265 1550
rect 3225 1520 3235 1540
rect 3255 1520 3265 1540
rect 3225 1510 3265 1520
rect 3345 1540 3385 1550
rect 3345 1520 3355 1540
rect 3375 1520 3385 1540
rect 3345 1510 3385 1520
rect 3465 1540 3505 1550
rect 3465 1520 3475 1540
rect 3495 1520 3505 1540
rect 3465 1510 3505 1520
rect 3585 1540 3625 1550
rect 3585 1520 3595 1540
rect 3615 1520 3625 1540
rect 3585 1510 3625 1520
rect 3705 1540 3745 1550
rect 3705 1520 3715 1540
rect 3735 1520 3745 1540
rect 3705 1510 3745 1520
rect 4265 1540 4305 1550
rect 4265 1520 4275 1540
rect 4295 1520 4305 1540
rect 4265 1510 4305 1520
rect 4385 1540 4425 1550
rect 4385 1520 4395 1540
rect 4415 1520 4425 1540
rect 4385 1510 4425 1520
rect 4505 1540 4545 1550
rect 4505 1520 4515 1540
rect 4535 1520 4545 1540
rect 4505 1510 4545 1520
rect 4625 1540 4665 1550
rect 4625 1520 4635 1540
rect 4655 1520 4665 1540
rect 4625 1510 4665 1520
rect 4745 1540 4785 1550
rect 4745 1520 4755 1540
rect 4775 1520 4785 1540
rect 4745 1510 4785 1520
rect 2925 1495 2965 1505
rect 2835 1480 2875 1490
rect 2835 1460 2845 1480
rect 2865 1460 2875 1480
rect 2925 1475 2935 1495
rect 2955 1475 2965 1495
rect 2925 1465 2965 1475
rect 3045 1495 3085 1505
rect 3045 1475 3055 1495
rect 3075 1475 3085 1495
rect 3045 1465 3085 1475
rect 3165 1495 3205 1505
rect 3165 1475 3175 1495
rect 3195 1475 3205 1495
rect 3165 1465 3205 1475
rect 3285 1495 3325 1505
rect 3285 1475 3295 1495
rect 3315 1475 3325 1495
rect 3285 1465 3325 1475
rect 3525 1495 3565 1505
rect 3525 1475 3535 1495
rect 3555 1475 3565 1495
rect 3525 1465 3565 1475
rect 3645 1495 3685 1505
rect 3645 1475 3655 1495
rect 3675 1475 3685 1495
rect 3645 1465 3685 1475
rect 3765 1495 3805 1505
rect 3765 1475 3775 1495
rect 3795 1475 3805 1495
rect 4205 1495 4245 1505
rect 3765 1465 3805 1475
rect 3915 1480 3955 1490
rect 2835 1450 2875 1460
rect 3915 1460 3925 1480
rect 3945 1460 3955 1480
rect 3915 1450 3955 1460
rect 4055 1480 4095 1490
rect 4055 1460 4065 1480
rect 4085 1460 4095 1480
rect 4205 1475 4215 1495
rect 4235 1475 4245 1495
rect 4205 1465 4245 1475
rect 4325 1495 4365 1505
rect 4325 1475 4335 1495
rect 4355 1475 4365 1495
rect 4325 1465 4365 1475
rect 4445 1495 4485 1505
rect 4445 1475 4455 1495
rect 4475 1475 4485 1495
rect 4445 1465 4485 1475
rect 4685 1495 4725 1505
rect 4685 1475 4695 1495
rect 4715 1475 4725 1495
rect 4685 1465 4725 1475
rect 4805 1495 4845 1505
rect 4805 1475 4815 1495
rect 4835 1475 4845 1495
rect 4805 1465 4845 1475
rect 4925 1495 4965 1505
rect 4925 1475 4935 1495
rect 4955 1475 4965 1495
rect 4925 1465 4965 1475
rect 5045 1495 5085 1505
rect 5045 1475 5055 1495
rect 5075 1475 5085 1495
rect 5045 1465 5085 1475
rect 5135 1480 5175 1490
rect 4055 1450 4095 1460
rect 5135 1460 5145 1480
rect 5165 1460 5175 1480
rect 5135 1450 5175 1460
rect 125 1335 2135 1375
rect 650 690 775 1335
rect 1330 690 1455 1335
rect 2010 695 2135 1335
rect 2840 1440 2870 1450
rect 2840 1420 2845 1440
rect 2865 1420 2870 1440
rect 2840 1390 2870 1420
rect 2840 1370 2845 1390
rect 2865 1370 2870 1390
rect 2840 1340 2870 1370
rect 2840 1320 2845 1340
rect 2865 1320 2870 1340
rect 2840 1290 2870 1320
rect 2840 1270 2845 1290
rect 2865 1270 2870 1290
rect 2840 1240 2870 1270
rect 2840 1220 2845 1240
rect 2865 1220 2870 1240
rect 2840 1210 2870 1220
rect 3380 1440 3410 1450
rect 3380 1420 3385 1440
rect 3405 1420 3410 1440
rect 3380 1390 3410 1420
rect 3380 1370 3385 1390
rect 3405 1370 3410 1390
rect 3380 1340 3410 1370
rect 3380 1320 3385 1340
rect 3405 1320 3410 1340
rect 3380 1290 3410 1320
rect 3380 1270 3385 1290
rect 3405 1270 3410 1290
rect 3380 1240 3410 1270
rect 3380 1220 3385 1240
rect 3405 1220 3410 1240
rect 3380 1210 3410 1220
rect 3920 1440 3950 1450
rect 3920 1420 3925 1440
rect 3945 1420 3950 1440
rect 3920 1390 3950 1420
rect 3920 1370 3925 1390
rect 3945 1370 3950 1390
rect 3920 1340 3950 1370
rect 3920 1320 3925 1340
rect 3945 1320 3950 1340
rect 3920 1290 3950 1320
rect 3920 1270 3925 1290
rect 3945 1270 3950 1290
rect 3920 1240 3950 1270
rect 3920 1220 3925 1240
rect 3945 1220 3950 1240
rect 3920 1210 3950 1220
rect 4060 1440 4090 1450
rect 4060 1420 4065 1440
rect 4085 1420 4090 1440
rect 4060 1390 4090 1420
rect 4060 1370 4065 1390
rect 4085 1370 4090 1390
rect 4060 1340 4090 1370
rect 4060 1320 4065 1340
rect 4085 1320 4090 1340
rect 4060 1290 4090 1320
rect 4060 1270 4065 1290
rect 4085 1270 4090 1290
rect 4060 1240 4090 1270
rect 4060 1220 4065 1240
rect 4085 1220 4090 1240
rect 4060 1210 4090 1220
rect 4600 1440 4630 1450
rect 4600 1420 4605 1440
rect 4625 1420 4630 1440
rect 4600 1390 4630 1420
rect 4600 1370 4605 1390
rect 4625 1370 4630 1390
rect 4600 1340 4630 1370
rect 4600 1320 4605 1340
rect 4625 1320 4630 1340
rect 4600 1290 4630 1320
rect 4600 1270 4605 1290
rect 4625 1270 4630 1290
rect 4600 1240 4630 1270
rect 4600 1220 4605 1240
rect 4625 1220 4630 1240
rect 4600 1210 4630 1220
rect 5140 1440 5170 1450
rect 5140 1420 5145 1440
rect 5165 1420 5170 1440
rect 5140 1390 5170 1420
rect 5140 1370 5145 1390
rect 5165 1370 5170 1390
rect 15030 1640 15065 1650
rect 15030 1615 15035 1640
rect 15060 1615 15065 1640
rect 15030 1605 15065 1615
rect 15120 1640 15190 1650
rect 15120 1620 15125 1640
rect 15145 1620 15165 1640
rect 15185 1620 15190 1640
rect 15120 1590 15190 1620
rect 15120 1570 15125 1590
rect 15145 1570 15165 1590
rect 15185 1570 15190 1590
rect 15120 1540 15190 1570
rect 15120 1520 15125 1540
rect 15145 1520 15165 1540
rect 15185 1520 15190 1540
rect 15120 1490 15190 1520
rect 15120 1470 15125 1490
rect 15145 1470 15165 1490
rect 15185 1470 15190 1490
rect 15120 1440 15190 1470
rect 15120 1420 15125 1440
rect 15145 1420 15165 1440
rect 15185 1420 15190 1440
rect 15120 1390 15190 1420
rect 5140 1340 5170 1370
rect 5140 1320 5145 1340
rect 5165 1320 5170 1340
rect 5140 1290 5170 1320
rect 5140 1270 5145 1290
rect 5165 1270 5170 1290
rect 5140 1240 5170 1270
rect 5140 1220 5145 1240
rect 5165 1220 5170 1240
rect 5140 1210 5170 1220
rect 15120 1370 15125 1390
rect 15145 1370 15165 1390
rect 15185 1370 15190 1390
rect 15120 1340 15190 1370
rect 15120 1320 15125 1340
rect 15145 1320 15165 1340
rect 15185 1320 15190 1340
rect 15120 1290 15190 1320
rect 15120 1270 15125 1290
rect 15145 1270 15165 1290
rect 15185 1270 15190 1290
rect 15120 1240 15190 1270
rect 15120 1220 15125 1240
rect 15145 1220 15165 1240
rect 15185 1220 15190 1240
rect 3385 1190 3405 1210
rect 4605 1190 4625 1210
rect 15120 1190 15190 1220
rect 3375 1180 3415 1190
rect 3375 1160 3385 1180
rect 3405 1160 3415 1180
rect 3375 1150 3415 1160
rect 3990 1155 4020 1185
rect 4595 1180 4635 1190
rect 4595 1160 4605 1180
rect 4625 1160 4635 1180
rect 4595 1150 4635 1160
rect 15120 1170 15125 1190
rect 15145 1170 15165 1190
rect 15185 1170 15190 1190
rect 15120 1140 15190 1170
rect 2945 1120 2985 1130
rect 2945 1100 2955 1120
rect 2975 1100 2985 1120
rect 2945 1090 2985 1100
rect 3025 1120 3065 1130
rect 3025 1100 3035 1120
rect 3055 1100 3065 1120
rect 3025 1090 3065 1100
rect 3105 1120 3145 1130
rect 3105 1100 3115 1120
rect 3135 1100 3145 1120
rect 3105 1090 3145 1100
rect 3185 1120 3225 1130
rect 3185 1100 3195 1120
rect 3215 1100 3225 1120
rect 3185 1090 3225 1100
rect 3265 1120 3305 1130
rect 3265 1100 3275 1120
rect 3295 1100 3305 1120
rect 3265 1090 3305 1100
rect 3345 1120 3385 1130
rect 3345 1100 3355 1120
rect 3375 1100 3385 1120
rect 3345 1090 3385 1100
rect 3425 1120 3465 1130
rect 3425 1100 3435 1120
rect 3455 1100 3465 1120
rect 3425 1090 3465 1100
rect 3505 1120 3545 1130
rect 3505 1100 3515 1120
rect 3535 1100 3545 1120
rect 3505 1090 3545 1100
rect 3585 1120 3625 1130
rect 3585 1100 3595 1120
rect 3615 1100 3625 1120
rect 3585 1090 3625 1100
rect 3665 1120 3705 1130
rect 3665 1100 3675 1120
rect 3695 1100 3705 1120
rect 3665 1090 3705 1100
rect 3745 1120 3785 1130
rect 3745 1100 3755 1120
rect 3775 1100 3785 1120
rect 3745 1090 3785 1100
rect 3825 1120 3865 1130
rect 3825 1100 3835 1120
rect 3855 1100 3865 1120
rect 3825 1090 3865 1100
rect 3905 1120 3945 1130
rect 3905 1100 3915 1120
rect 3935 1100 3945 1120
rect 3905 1090 3945 1100
rect 3985 1120 4025 1130
rect 3985 1100 3995 1120
rect 4015 1100 4025 1120
rect 3985 1090 4025 1100
rect 4065 1120 4105 1130
rect 4065 1100 4075 1120
rect 4095 1100 4105 1120
rect 4065 1090 4105 1100
rect 4145 1120 4185 1130
rect 4145 1100 4155 1120
rect 4175 1100 4185 1120
rect 4145 1090 4185 1100
rect 4225 1120 4265 1130
rect 4225 1100 4235 1120
rect 4255 1100 4265 1120
rect 4225 1090 4265 1100
rect 4305 1120 4345 1130
rect 4305 1100 4315 1120
rect 4335 1100 4345 1120
rect 4305 1090 4345 1100
rect 4385 1120 4425 1130
rect 4385 1100 4395 1120
rect 4415 1100 4425 1120
rect 4385 1090 4425 1100
rect 4465 1120 4505 1130
rect 4465 1100 4475 1120
rect 4495 1100 4505 1120
rect 4465 1090 4505 1100
rect 4545 1120 4585 1130
rect 4545 1100 4555 1120
rect 4575 1100 4585 1120
rect 4545 1090 4585 1100
rect 4625 1120 4665 1130
rect 4625 1100 4635 1120
rect 4655 1100 4665 1120
rect 4625 1090 4665 1100
rect 4705 1120 4745 1130
rect 4705 1100 4715 1120
rect 4735 1100 4745 1120
rect 4705 1090 4745 1100
rect 4785 1120 4825 1130
rect 4785 1100 4795 1120
rect 4815 1100 4825 1120
rect 4785 1090 4825 1100
rect 4865 1120 4905 1130
rect 4865 1100 4875 1120
rect 4895 1100 4905 1120
rect 4865 1090 4905 1100
rect 4945 1120 4985 1130
rect 4945 1100 4955 1120
rect 4975 1100 4985 1120
rect 4945 1090 4985 1100
rect 2955 1070 2975 1090
rect 3995 1070 4015 1090
rect 2950 1060 2980 1070
rect 2950 1045 2955 1060
rect 2935 1040 2955 1045
rect 2975 1040 2980 1060
rect 2625 1010 2655 1040
rect 2910 1035 2980 1040
rect 2910 1015 2915 1035
rect 2935 1015 2980 1035
rect 2910 1010 2980 1015
rect 2935 1005 2955 1010
rect 2950 990 2955 1005
rect 2975 990 2980 1010
rect 2950 980 2980 990
rect 3990 1060 4020 1070
rect 3990 1040 3995 1060
rect 4015 1040 4020 1060
rect 3990 1010 4020 1040
rect 3990 990 3995 1010
rect 4015 990 4020 1010
rect 3990 980 4020 990
rect 5030 1060 5100 1070
rect 5030 1040 5035 1060
rect 5055 1040 5075 1060
rect 5095 1045 5100 1060
rect 5095 1040 5150 1045
rect 5030 1035 5150 1040
rect 5030 1015 5120 1035
rect 5140 1015 5150 1035
rect 5030 1010 5150 1015
rect 5030 990 5035 1010
rect 5055 990 5075 1010
rect 5095 1005 5150 1010
rect 5095 990 5100 1005
rect 5030 980 5100 990
rect 2995 925 3035 935
rect 2995 905 3005 925
rect 3025 905 3035 925
rect 2995 895 3035 905
rect 3175 925 3215 935
rect 3175 905 3185 925
rect 3205 905 3215 925
rect 3175 895 3215 905
rect 3355 925 3395 935
rect 3355 905 3365 925
rect 3385 905 3395 925
rect 3355 895 3395 905
rect 3535 925 3575 935
rect 3535 905 3545 925
rect 3565 905 3575 925
rect 3535 895 3575 905
rect 3715 925 3755 935
rect 3715 905 3725 925
rect 3745 905 3755 925
rect 3715 895 3755 905
rect 3895 925 3935 935
rect 3895 905 3905 925
rect 3925 905 3935 925
rect 3895 895 3935 905
rect 4075 925 4115 935
rect 4075 905 4085 925
rect 4105 905 4115 925
rect 4075 895 4115 905
rect 4255 925 4295 935
rect 4255 905 4265 925
rect 4285 905 4295 925
rect 4255 895 4295 905
rect 4435 925 4475 935
rect 4435 905 4445 925
rect 4465 905 4475 925
rect 4435 895 4475 905
rect 4615 925 4655 935
rect 4615 905 4625 925
rect 4645 905 4655 925
rect 4615 895 4655 905
rect 4795 925 4835 935
rect 4795 905 4805 925
rect 4825 905 4835 925
rect 4795 895 4835 905
rect 4975 925 5015 935
rect 4975 905 4985 925
rect 5005 905 5015 925
rect 15005 910 15030 960
rect 15120 1120 15125 1140
rect 15145 1120 15165 1140
rect 15185 1120 15190 1140
rect 15120 1090 15190 1120
rect 15120 1070 15125 1090
rect 15145 1070 15165 1090
rect 15185 1070 15190 1090
rect 15120 1040 15190 1070
rect 15120 1020 15125 1040
rect 15145 1020 15165 1040
rect 15185 1020 15190 1040
rect 15120 990 15190 1020
rect 15120 970 15125 990
rect 15145 970 15165 990
rect 15185 970 15190 990
rect 15120 960 15190 970
rect 15260 1640 15290 1650
rect 15260 1620 15265 1640
rect 15285 1620 15290 1640
rect 15260 1590 15290 1620
rect 15260 1570 15265 1590
rect 15285 1570 15290 1590
rect 15260 1540 15290 1570
rect 15260 1520 15265 1540
rect 15285 1520 15290 1540
rect 15260 1490 15290 1520
rect 15260 1470 15265 1490
rect 15285 1470 15290 1490
rect 15260 1440 15290 1470
rect 15260 1420 15265 1440
rect 15285 1420 15290 1440
rect 15260 1390 15290 1420
rect 15260 1370 15265 1390
rect 15285 1370 15290 1390
rect 15260 1340 15290 1370
rect 15260 1320 15265 1340
rect 15285 1320 15290 1340
rect 15260 1290 15290 1320
rect 15260 1270 15265 1290
rect 15285 1270 15290 1290
rect 15260 1240 15290 1270
rect 15260 1220 15265 1240
rect 15285 1220 15290 1240
rect 15260 1190 15290 1220
rect 15260 1170 15265 1190
rect 15285 1170 15290 1190
rect 15260 1140 15290 1170
rect 15260 1120 15265 1140
rect 15285 1120 15290 1140
rect 15260 1090 15290 1120
rect 15260 1070 15265 1090
rect 15285 1070 15290 1090
rect 15260 1040 15290 1070
rect 15260 1020 15265 1040
rect 15285 1020 15290 1040
rect 15260 990 15290 1020
rect 15260 970 15265 990
rect 15285 970 15290 990
rect 15260 960 15290 970
rect 15360 1640 15390 1650
rect 15360 1620 15365 1640
rect 15385 1620 15390 1640
rect 15360 1590 15390 1620
rect 15360 1570 15365 1590
rect 15385 1570 15390 1590
rect 15360 1540 15390 1570
rect 15360 1520 15365 1540
rect 15385 1520 15390 1540
rect 15360 1490 15390 1520
rect 15360 1470 15365 1490
rect 15385 1470 15390 1490
rect 15360 1440 15390 1470
rect 15360 1420 15365 1440
rect 15385 1420 15390 1440
rect 15360 1390 15390 1420
rect 15360 1370 15365 1390
rect 15385 1370 15390 1390
rect 15360 1340 15390 1370
rect 15360 1320 15365 1340
rect 15385 1320 15390 1340
rect 15360 1290 15390 1320
rect 15360 1270 15365 1290
rect 15385 1270 15390 1290
rect 15360 1240 15390 1270
rect 15360 1220 15365 1240
rect 15385 1220 15390 1240
rect 15360 1190 15390 1220
rect 15360 1170 15365 1190
rect 15385 1170 15390 1190
rect 15360 1140 15390 1170
rect 15360 1120 15365 1140
rect 15385 1120 15390 1140
rect 15360 1090 15390 1120
rect 15360 1070 15365 1090
rect 15385 1070 15390 1090
rect 15360 1040 15390 1070
rect 15360 1020 15365 1040
rect 15385 1020 15390 1040
rect 15360 990 15390 1020
rect 15360 970 15365 990
rect 15385 970 15390 990
rect 15360 960 15390 970
rect 15460 1640 15490 1650
rect 15460 1620 15465 1640
rect 15485 1620 15490 1640
rect 15460 1590 15490 1620
rect 15460 1570 15465 1590
rect 15485 1570 15490 1590
rect 15460 1540 15490 1570
rect 15460 1520 15465 1540
rect 15485 1520 15490 1540
rect 15460 1490 15490 1520
rect 15460 1470 15465 1490
rect 15485 1470 15490 1490
rect 15460 1440 15490 1470
rect 15460 1420 15465 1440
rect 15485 1420 15490 1440
rect 15460 1390 15490 1420
rect 15460 1370 15465 1390
rect 15485 1370 15490 1390
rect 15460 1340 15490 1370
rect 15460 1320 15465 1340
rect 15485 1320 15490 1340
rect 15460 1290 15490 1320
rect 15460 1270 15465 1290
rect 15485 1270 15490 1290
rect 15460 1240 15490 1270
rect 15460 1220 15465 1240
rect 15485 1220 15490 1240
rect 15460 1190 15490 1220
rect 15460 1170 15465 1190
rect 15485 1170 15490 1190
rect 15460 1140 15490 1170
rect 15460 1120 15465 1140
rect 15485 1120 15490 1140
rect 15460 1090 15490 1120
rect 15460 1070 15465 1090
rect 15485 1070 15490 1090
rect 15460 1040 15490 1070
rect 15460 1020 15465 1040
rect 15485 1020 15490 1040
rect 15460 990 15490 1020
rect 15460 970 15465 990
rect 15485 970 15490 990
rect 15460 960 15490 970
rect 15560 1640 15590 1650
rect 15560 1620 15565 1640
rect 15585 1620 15590 1640
rect 15560 1590 15590 1620
rect 15560 1570 15565 1590
rect 15585 1570 15590 1590
rect 15560 1540 15590 1570
rect 15560 1520 15565 1540
rect 15585 1520 15590 1540
rect 15560 1490 15590 1520
rect 15560 1470 15565 1490
rect 15585 1470 15590 1490
rect 15560 1440 15590 1470
rect 15560 1420 15565 1440
rect 15585 1420 15590 1440
rect 15560 1390 15590 1420
rect 15560 1370 15565 1390
rect 15585 1370 15590 1390
rect 15560 1340 15590 1370
rect 15560 1320 15565 1340
rect 15585 1320 15590 1340
rect 15560 1290 15590 1320
rect 15560 1270 15565 1290
rect 15585 1270 15590 1290
rect 15560 1240 15590 1270
rect 15560 1220 15565 1240
rect 15585 1220 15590 1240
rect 15560 1190 15590 1220
rect 15560 1170 15565 1190
rect 15585 1170 15590 1190
rect 15560 1140 15590 1170
rect 15560 1120 15565 1140
rect 15585 1120 15590 1140
rect 15560 1090 15590 1120
rect 15560 1070 15565 1090
rect 15585 1070 15590 1090
rect 15560 1040 15590 1070
rect 15560 1020 15565 1040
rect 15585 1020 15590 1040
rect 15560 990 15590 1020
rect 15560 970 15565 990
rect 15585 970 15590 990
rect 15560 960 15590 970
rect 15660 1640 15690 1650
rect 15660 1620 15665 1640
rect 15685 1620 15690 1640
rect 15660 1590 15690 1620
rect 15660 1570 15665 1590
rect 15685 1570 15690 1590
rect 15660 1540 15690 1570
rect 15660 1520 15665 1540
rect 15685 1520 15690 1540
rect 15660 1490 15690 1520
rect 15660 1470 15665 1490
rect 15685 1470 15690 1490
rect 15660 1440 15690 1470
rect 15660 1420 15665 1440
rect 15685 1420 15690 1440
rect 15660 1390 15690 1420
rect 15660 1370 15665 1390
rect 15685 1370 15690 1390
rect 15660 1340 15690 1370
rect 15660 1320 15665 1340
rect 15685 1320 15690 1340
rect 15660 1290 15690 1320
rect 15660 1270 15665 1290
rect 15685 1270 15690 1290
rect 15660 1240 15690 1270
rect 15660 1220 15665 1240
rect 15685 1220 15690 1240
rect 15660 1190 15690 1220
rect 15660 1170 15665 1190
rect 15685 1170 15690 1190
rect 15660 1140 15690 1170
rect 15660 1120 15665 1140
rect 15685 1120 15690 1140
rect 15660 1090 15690 1120
rect 15660 1070 15665 1090
rect 15685 1070 15690 1090
rect 15660 1040 15690 1070
rect 15660 1020 15665 1040
rect 15685 1020 15690 1040
rect 15660 990 15690 1020
rect 15660 970 15665 990
rect 15685 970 15690 990
rect 15660 960 15690 970
rect 15760 1640 15830 1650
rect 15760 1620 15765 1640
rect 15785 1620 15805 1640
rect 15825 1620 15830 1640
rect 15760 1590 15830 1620
rect 15760 1570 15765 1590
rect 15785 1570 15805 1590
rect 15825 1570 15830 1590
rect 15760 1540 15830 1570
rect 15760 1520 15765 1540
rect 15785 1520 15805 1540
rect 15825 1520 15830 1540
rect 15990 1630 16000 1650
rect 16020 1630 16040 1650
rect 16060 1630 16065 1650
rect 15990 1600 16065 1630
rect 15990 1580 16000 1600
rect 16020 1580 16040 1600
rect 16060 1580 16065 1600
rect 15990 1550 16065 1580
rect 15990 1530 16000 1550
rect 16020 1530 16040 1550
rect 16060 1530 16065 1550
rect 15990 1520 16065 1530
rect 16090 1650 16120 1660
rect 16090 1630 16095 1650
rect 16115 1630 16120 1650
rect 16090 1600 16120 1630
rect 16090 1580 16095 1600
rect 16115 1580 16120 1600
rect 16090 1550 16120 1580
rect 16090 1530 16095 1550
rect 16115 1530 16120 1550
rect 16090 1520 16120 1530
rect 16145 1650 16175 1660
rect 16145 1630 16150 1650
rect 16170 1630 16175 1650
rect 16145 1600 16175 1630
rect 16145 1580 16150 1600
rect 16170 1580 16175 1600
rect 16145 1550 16175 1580
rect 16145 1530 16150 1550
rect 16170 1530 16175 1550
rect 16145 1520 16175 1530
rect 16200 1650 16230 1660
rect 16200 1630 16205 1650
rect 16225 1630 16230 1650
rect 16200 1600 16230 1630
rect 16200 1580 16205 1600
rect 16225 1580 16230 1600
rect 16200 1550 16230 1580
rect 16200 1530 16205 1550
rect 16225 1530 16230 1550
rect 16200 1520 16230 1530
rect 16255 1650 16285 1660
rect 16255 1630 16260 1650
rect 16280 1630 16285 1650
rect 16255 1600 16285 1630
rect 16255 1580 16260 1600
rect 16280 1580 16285 1600
rect 16255 1550 16285 1580
rect 16255 1530 16260 1550
rect 16280 1530 16285 1550
rect 16255 1520 16285 1530
rect 16310 1650 16340 1660
rect 16310 1630 16315 1650
rect 16335 1630 16340 1650
rect 16310 1600 16340 1630
rect 16310 1580 16315 1600
rect 16335 1580 16340 1600
rect 16310 1550 16340 1580
rect 16310 1530 16315 1550
rect 16335 1530 16340 1550
rect 16310 1520 16340 1530
rect 16365 1650 16395 1660
rect 16365 1630 16370 1650
rect 16390 1630 16395 1650
rect 16365 1600 16395 1630
rect 16365 1580 16370 1600
rect 16390 1580 16395 1600
rect 16365 1550 16395 1580
rect 16365 1530 16370 1550
rect 16390 1530 16395 1550
rect 16365 1520 16395 1530
rect 16420 1650 16450 1660
rect 16420 1630 16425 1650
rect 16445 1630 16450 1650
rect 16420 1600 16450 1630
rect 16420 1580 16425 1600
rect 16445 1580 16450 1600
rect 16420 1550 16450 1580
rect 16420 1530 16425 1550
rect 16445 1530 16450 1550
rect 16420 1520 16450 1530
rect 16475 1650 16505 1660
rect 16475 1630 16480 1650
rect 16500 1630 16505 1650
rect 16475 1600 16505 1630
rect 16475 1580 16480 1600
rect 16500 1580 16505 1600
rect 16475 1550 16505 1580
rect 16475 1530 16480 1550
rect 16500 1530 16505 1550
rect 16475 1520 16505 1530
rect 16530 1650 16560 1660
rect 16530 1630 16535 1650
rect 16555 1630 16560 1650
rect 16530 1600 16560 1630
rect 16530 1580 16535 1600
rect 16555 1580 16560 1600
rect 16530 1550 16560 1580
rect 16530 1530 16535 1550
rect 16555 1530 16560 1550
rect 16530 1520 16560 1530
rect 16585 1650 16615 1660
rect 16585 1630 16590 1650
rect 16610 1630 16615 1650
rect 16585 1600 16615 1630
rect 16585 1580 16590 1600
rect 16610 1580 16615 1600
rect 16585 1550 16615 1580
rect 16585 1530 16590 1550
rect 16610 1530 16615 1550
rect 16585 1520 16615 1530
rect 16640 1650 16670 1660
rect 16640 1630 16645 1650
rect 16665 1630 16670 1650
rect 16640 1600 16670 1630
rect 16640 1580 16645 1600
rect 16665 1580 16670 1600
rect 16640 1550 16670 1580
rect 16640 1530 16645 1550
rect 16665 1530 16670 1550
rect 16640 1520 16670 1530
rect 16695 1650 16805 1660
rect 16695 1630 16700 1650
rect 16720 1630 16740 1650
rect 16760 1630 16780 1650
rect 16800 1630 16805 1650
rect 16695 1600 16805 1630
rect 16695 1580 16700 1600
rect 16720 1580 16740 1600
rect 16760 1580 16780 1600
rect 16800 1580 16805 1600
rect 16695 1550 16805 1580
rect 16695 1530 16700 1550
rect 16720 1530 16740 1550
rect 16760 1530 16780 1550
rect 16800 1530 16805 1550
rect 16695 1520 16805 1530
rect 16830 1650 16860 1660
rect 16830 1630 16835 1650
rect 16855 1630 16860 1650
rect 16830 1600 16860 1630
rect 16830 1580 16835 1600
rect 16855 1580 16860 1600
rect 16830 1550 16860 1580
rect 16830 1530 16835 1550
rect 16855 1530 16860 1550
rect 16830 1520 16860 1530
rect 16885 1650 16915 1660
rect 16885 1630 16890 1650
rect 16910 1630 16915 1650
rect 16885 1600 16915 1630
rect 16885 1580 16890 1600
rect 16910 1580 16915 1600
rect 16885 1550 16915 1580
rect 16885 1530 16890 1550
rect 16910 1530 16915 1550
rect 16885 1520 16915 1530
rect 16940 1650 16970 1660
rect 16940 1630 16945 1650
rect 16965 1630 16970 1650
rect 16940 1600 16970 1630
rect 16940 1580 16945 1600
rect 16965 1580 16970 1600
rect 16940 1550 16970 1580
rect 16940 1530 16945 1550
rect 16965 1530 16970 1550
rect 16940 1520 16970 1530
rect 16995 1650 17105 1660
rect 16995 1630 17000 1650
rect 17020 1630 17040 1650
rect 17060 1630 17080 1650
rect 17100 1630 17105 1650
rect 16995 1600 17105 1630
rect 16995 1580 17000 1600
rect 17020 1580 17040 1600
rect 17060 1580 17080 1600
rect 17100 1580 17105 1600
rect 16995 1550 17105 1580
rect 16995 1530 17000 1550
rect 17020 1530 17040 1550
rect 17060 1530 17080 1550
rect 17100 1530 17105 1550
rect 16995 1520 17105 1530
rect 17130 1650 17160 1660
rect 17130 1630 17135 1650
rect 17155 1630 17160 1650
rect 17130 1600 17160 1630
rect 17130 1580 17135 1600
rect 17155 1580 17160 1600
rect 17130 1550 17160 1580
rect 17130 1530 17135 1550
rect 17155 1530 17160 1550
rect 17130 1520 17160 1530
rect 17185 1650 17215 1660
rect 17185 1630 17190 1650
rect 17210 1630 17215 1650
rect 17185 1600 17215 1630
rect 17185 1580 17190 1600
rect 17210 1580 17215 1600
rect 17185 1550 17215 1580
rect 17185 1530 17190 1550
rect 17210 1530 17215 1550
rect 17185 1520 17215 1530
rect 17240 1650 17270 1660
rect 17240 1630 17245 1650
rect 17265 1630 17270 1650
rect 17240 1600 17270 1630
rect 17240 1580 17245 1600
rect 17265 1580 17270 1600
rect 17240 1550 17270 1580
rect 17240 1530 17245 1550
rect 17265 1530 17270 1550
rect 17240 1520 17270 1530
rect 17295 1650 17325 1660
rect 17295 1630 17300 1650
rect 17320 1630 17325 1650
rect 17295 1600 17325 1630
rect 17295 1580 17300 1600
rect 17320 1580 17325 1600
rect 17295 1550 17325 1580
rect 17295 1530 17300 1550
rect 17320 1530 17325 1550
rect 17295 1520 17325 1530
rect 17350 1650 17380 1660
rect 17350 1630 17355 1650
rect 17375 1630 17380 1650
rect 17350 1600 17380 1630
rect 17350 1580 17355 1600
rect 17375 1580 17380 1600
rect 17350 1550 17380 1580
rect 17350 1530 17355 1550
rect 17375 1530 17380 1550
rect 17350 1520 17380 1530
rect 17405 1650 17435 1660
rect 17405 1630 17410 1650
rect 17430 1630 17435 1650
rect 17405 1600 17435 1630
rect 17405 1580 17410 1600
rect 17430 1580 17435 1600
rect 17405 1550 17435 1580
rect 17405 1530 17410 1550
rect 17430 1530 17435 1550
rect 17405 1520 17435 1530
rect 17460 1650 17490 1660
rect 17460 1630 17465 1650
rect 17485 1630 17490 1650
rect 17460 1600 17490 1630
rect 17460 1580 17465 1600
rect 17485 1580 17490 1600
rect 17460 1550 17490 1580
rect 17460 1530 17465 1550
rect 17485 1530 17490 1550
rect 17460 1520 17490 1530
rect 17515 1650 17545 1660
rect 17515 1630 17520 1650
rect 17540 1630 17545 1650
rect 17515 1600 17545 1630
rect 17515 1580 17520 1600
rect 17540 1580 17545 1600
rect 17515 1550 17545 1580
rect 17515 1530 17520 1550
rect 17540 1530 17545 1550
rect 17515 1520 17545 1530
rect 17570 1650 17600 1660
rect 17570 1630 17575 1650
rect 17595 1630 17600 1650
rect 17570 1600 17600 1630
rect 17570 1580 17575 1600
rect 17595 1580 17600 1600
rect 17570 1550 17600 1580
rect 17570 1530 17575 1550
rect 17595 1530 17600 1550
rect 17570 1520 17600 1530
rect 17625 1650 17655 1660
rect 17625 1630 17630 1650
rect 17650 1630 17655 1650
rect 17625 1600 17655 1630
rect 17625 1580 17630 1600
rect 17650 1580 17655 1600
rect 17625 1550 17655 1580
rect 17625 1530 17630 1550
rect 17650 1530 17655 1550
rect 17625 1520 17655 1530
rect 17680 1650 17710 1660
rect 17680 1630 17685 1650
rect 17705 1630 17710 1650
rect 17680 1600 17710 1630
rect 17680 1580 17685 1600
rect 17705 1580 17710 1600
rect 17680 1550 17710 1580
rect 17680 1530 17685 1550
rect 17705 1530 17710 1550
rect 17680 1520 17710 1530
rect 17735 1650 17810 1660
rect 18115 1650 18135 1670
rect 18315 1650 18335 1670
rect 18515 1650 18535 1670
rect 17735 1630 17740 1650
rect 17760 1630 17780 1650
rect 17800 1630 17810 1650
rect 17735 1600 17810 1630
rect 17735 1580 17740 1600
rect 17760 1580 17780 1600
rect 17800 1580 17810 1600
rect 17735 1550 17810 1580
rect 17735 1530 17740 1550
rect 17760 1530 17780 1550
rect 17800 1530 17810 1550
rect 17735 1520 17810 1530
rect 17970 1640 18040 1650
rect 17970 1620 17975 1640
rect 17995 1620 18015 1640
rect 18035 1620 18040 1640
rect 17970 1590 18040 1620
rect 17970 1570 17975 1590
rect 17995 1570 18015 1590
rect 18035 1570 18040 1590
rect 17970 1540 18040 1570
rect 17970 1520 17975 1540
rect 17995 1520 18015 1540
rect 18035 1520 18040 1540
rect 15760 1490 15830 1520
rect 16000 1500 16020 1520
rect 15760 1470 15765 1490
rect 15785 1470 15805 1490
rect 15825 1470 15830 1490
rect 15760 1440 15830 1470
rect 15990 1490 16030 1500
rect 15990 1470 16000 1490
rect 16020 1470 16030 1490
rect 15990 1460 16030 1470
rect 16106 1490 16138 1500
rect 16106 1470 16112 1490
rect 16129 1470 16138 1490
rect 16106 1460 16138 1470
rect 16155 1440 16175 1520
rect 16260 1440 16280 1520
rect 16305 1490 16345 1500
rect 16305 1470 16315 1490
rect 16335 1470 16345 1490
rect 16305 1460 16345 1470
rect 16370 1440 16390 1520
rect 16480 1440 16500 1520
rect 16525 1490 16565 1500
rect 16525 1470 16535 1490
rect 16555 1470 16565 1490
rect 16525 1460 16565 1470
rect 16590 1440 16610 1520
rect 16740 1500 16760 1520
rect 16830 1500 16850 1520
rect 16885 1500 16905 1520
rect 17040 1500 17060 1520
rect 16730 1490 16770 1500
rect 16730 1470 16740 1490
rect 16760 1470 16770 1490
rect 16730 1460 16770 1470
rect 16825 1490 16855 1500
rect 16825 1470 16830 1490
rect 16850 1470 16855 1490
rect 16825 1460 16855 1470
rect 16875 1490 16905 1500
rect 16875 1470 16880 1490
rect 16900 1470 16905 1490
rect 16875 1460 16905 1470
rect 16922 1490 16954 1500
rect 16922 1470 16928 1490
rect 16945 1470 16954 1490
rect 16922 1460 16954 1470
rect 17030 1490 17070 1500
rect 17030 1470 17040 1490
rect 17060 1470 17070 1490
rect 17030 1460 17070 1470
rect 17146 1490 17178 1500
rect 17146 1470 17152 1490
rect 17169 1470 17178 1490
rect 17146 1460 17178 1470
rect 17195 1440 17215 1520
rect 17300 1440 17320 1520
rect 17345 1490 17385 1500
rect 17345 1470 17355 1490
rect 17375 1470 17385 1490
rect 17345 1460 17385 1470
rect 17410 1440 17430 1520
rect 17520 1440 17540 1520
rect 17565 1490 17605 1500
rect 17565 1470 17575 1490
rect 17595 1470 17605 1490
rect 17565 1460 17605 1470
rect 17630 1440 17650 1520
rect 17780 1500 17800 1520
rect 17770 1490 17810 1500
rect 17770 1470 17780 1490
rect 17800 1470 17810 1490
rect 17770 1460 17810 1470
rect 17970 1490 18040 1520
rect 17970 1470 17975 1490
rect 17995 1470 18015 1490
rect 18035 1470 18040 1490
rect 17970 1440 18040 1470
rect 15760 1420 15765 1440
rect 15785 1420 15805 1440
rect 15825 1420 15830 1440
rect 15760 1390 15830 1420
rect 16145 1430 16185 1440
rect 16145 1410 16155 1430
rect 16175 1410 16185 1430
rect 16145 1400 16185 1410
rect 16250 1430 16290 1440
rect 16250 1410 16260 1430
rect 16280 1410 16290 1430
rect 16250 1400 16290 1410
rect 16360 1430 16400 1440
rect 16360 1410 16370 1430
rect 16390 1410 16400 1430
rect 16360 1400 16400 1410
rect 16470 1430 16510 1440
rect 16470 1410 16480 1430
rect 16500 1410 16510 1430
rect 16470 1400 16510 1410
rect 16580 1430 16620 1440
rect 16580 1410 16590 1430
rect 16610 1410 16620 1430
rect 16580 1400 16620 1410
rect 17185 1430 17225 1440
rect 17185 1410 17195 1430
rect 17215 1410 17225 1430
rect 17185 1400 17225 1410
rect 17290 1430 17330 1440
rect 17290 1410 17300 1430
rect 17320 1410 17330 1430
rect 17290 1400 17330 1410
rect 17400 1430 17440 1440
rect 17400 1410 17410 1430
rect 17430 1410 17440 1430
rect 17400 1400 17440 1410
rect 17510 1430 17550 1440
rect 17510 1410 17520 1430
rect 17540 1410 17550 1430
rect 17510 1400 17550 1410
rect 17620 1430 17660 1440
rect 17620 1410 17630 1430
rect 17650 1410 17660 1430
rect 17620 1400 17660 1410
rect 17970 1420 17975 1440
rect 17995 1420 18015 1440
rect 18035 1420 18040 1440
rect 15760 1370 15765 1390
rect 15785 1370 15805 1390
rect 15825 1370 15830 1390
rect 15760 1340 15830 1370
rect 17970 1390 18040 1420
rect 17970 1370 17975 1390
rect 17995 1370 18015 1390
rect 18035 1370 18040 1390
rect 15760 1320 15765 1340
rect 15785 1320 15805 1340
rect 15825 1320 15830 1340
rect 15760 1290 15830 1320
rect 16810 1310 16850 1350
rect 17970 1340 18040 1370
rect 17970 1320 17975 1340
rect 17995 1320 18015 1340
rect 18035 1320 18040 1340
rect 15760 1270 15765 1290
rect 15785 1270 15805 1290
rect 15825 1270 15830 1290
rect 15760 1240 15830 1270
rect 16315 1260 16355 1300
rect 16880 1260 16920 1300
rect 17970 1290 18040 1320
rect 17970 1270 17975 1290
rect 17995 1270 18015 1290
rect 18035 1270 18040 1290
rect 17595 1245 17635 1255
rect 15760 1220 15765 1240
rect 15785 1220 15805 1240
rect 15825 1220 15830 1240
rect 15760 1190 15830 1220
rect 16315 1230 16355 1240
rect 16315 1210 16325 1230
rect 16345 1210 16355 1230
rect 16315 1200 16355 1210
rect 16425 1230 16465 1240
rect 16425 1210 16435 1230
rect 16455 1210 16465 1230
rect 16425 1200 16465 1210
rect 16535 1230 16575 1240
rect 16535 1210 16545 1230
rect 16565 1210 16575 1230
rect 16535 1200 16575 1210
rect 16645 1230 16685 1240
rect 16645 1210 16655 1230
rect 16675 1210 16685 1230
rect 16645 1200 16685 1210
rect 16755 1230 16795 1240
rect 16755 1210 16765 1230
rect 16785 1210 16795 1230
rect 16755 1200 16795 1210
rect 16815 1230 16845 1240
rect 16815 1210 16820 1230
rect 16840 1210 16845 1230
rect 16815 1200 16845 1210
rect 16865 1230 16905 1240
rect 16865 1210 16875 1230
rect 16895 1210 16905 1230
rect 16865 1200 16905 1210
rect 16975 1230 17015 1240
rect 16975 1210 16985 1230
rect 17005 1210 17015 1230
rect 16975 1200 17015 1210
rect 17085 1230 17125 1240
rect 17085 1210 17095 1230
rect 17115 1210 17125 1230
rect 17085 1200 17125 1210
rect 17195 1230 17235 1240
rect 17195 1210 17205 1230
rect 17225 1210 17235 1230
rect 17195 1200 17235 1210
rect 17305 1230 17345 1240
rect 17305 1210 17315 1230
rect 17335 1210 17345 1230
rect 17305 1200 17345 1210
rect 17415 1230 17455 1240
rect 17415 1210 17425 1230
rect 17445 1210 17455 1230
rect 17415 1200 17455 1210
rect 17525 1230 17565 1240
rect 17525 1210 17535 1230
rect 17555 1210 17565 1230
rect 17595 1225 17605 1245
rect 17625 1225 17635 1245
rect 17595 1215 17635 1225
rect 17970 1240 18040 1270
rect 17970 1220 17975 1240
rect 17995 1220 18015 1240
rect 18035 1220 18040 1240
rect 17525 1200 17565 1210
rect 15760 1170 15765 1190
rect 15785 1170 15805 1190
rect 15825 1170 15830 1190
rect 16325 1180 16345 1200
rect 16435 1180 16455 1200
rect 16545 1180 16565 1200
rect 16655 1180 16675 1200
rect 16765 1180 16785 1200
rect 16875 1180 16895 1200
rect 16985 1180 17005 1200
rect 17095 1180 17115 1200
rect 17205 1180 17225 1200
rect 17315 1180 17335 1200
rect 17425 1180 17445 1200
rect 17535 1180 17555 1200
rect 17970 1190 18040 1220
rect 15760 1140 15830 1170
rect 15760 1120 15765 1140
rect 15785 1120 15805 1140
rect 15825 1120 15830 1140
rect 15760 1090 15830 1120
rect 15760 1070 15765 1090
rect 15785 1070 15805 1090
rect 15825 1070 15830 1090
rect 15760 1040 15830 1070
rect 15760 1020 15765 1040
rect 15785 1020 15805 1040
rect 15825 1020 15830 1040
rect 15760 990 15830 1020
rect 15760 970 15765 990
rect 15785 970 15805 990
rect 15825 970 15830 990
rect 15760 960 15830 970
rect 16170 1170 16240 1180
rect 16170 1150 16175 1170
rect 16195 1150 16215 1170
rect 16235 1150 16240 1170
rect 16170 1120 16240 1150
rect 16170 1100 16175 1120
rect 16195 1100 16215 1120
rect 16235 1100 16240 1120
rect 16170 1070 16240 1100
rect 16170 1050 16175 1070
rect 16195 1050 16215 1070
rect 16235 1050 16240 1070
rect 16170 1020 16240 1050
rect 16170 1000 16175 1020
rect 16195 1000 16215 1020
rect 16235 1000 16240 1020
rect 16170 970 16240 1000
rect 15125 940 15145 960
rect 15365 940 15385 960
rect 15565 940 15585 960
rect 15805 940 15825 960
rect 16170 950 16175 970
rect 16195 950 16215 970
rect 16235 950 16240 970
rect 16170 940 16240 950
rect 16265 1170 16295 1180
rect 16265 1150 16270 1170
rect 16290 1150 16295 1170
rect 16265 1120 16295 1150
rect 16265 1100 16270 1120
rect 16290 1100 16295 1120
rect 16265 1070 16295 1100
rect 16265 1050 16270 1070
rect 16290 1050 16295 1070
rect 16265 1020 16295 1050
rect 16265 1000 16270 1020
rect 16290 1000 16295 1020
rect 16265 970 16295 1000
rect 16265 950 16270 970
rect 16290 950 16295 970
rect 16265 940 16295 950
rect 16320 1170 16350 1180
rect 16320 1150 16325 1170
rect 16345 1150 16350 1170
rect 16320 1120 16350 1150
rect 16320 1100 16325 1120
rect 16345 1100 16350 1120
rect 16320 1070 16350 1100
rect 16320 1050 16325 1070
rect 16345 1050 16350 1070
rect 16320 1020 16350 1050
rect 16320 1000 16325 1020
rect 16345 1000 16350 1020
rect 16320 970 16350 1000
rect 16320 950 16325 970
rect 16345 950 16350 970
rect 16320 940 16350 950
rect 16375 1170 16405 1180
rect 16375 1150 16380 1170
rect 16400 1150 16405 1170
rect 16375 1120 16405 1150
rect 16375 1100 16380 1120
rect 16400 1100 16405 1120
rect 16375 1070 16405 1100
rect 16375 1050 16380 1070
rect 16400 1050 16405 1070
rect 16375 1020 16405 1050
rect 16375 1000 16380 1020
rect 16400 1000 16405 1020
rect 16375 970 16405 1000
rect 16375 950 16380 970
rect 16400 950 16405 970
rect 16375 940 16405 950
rect 16430 1170 16460 1180
rect 16430 1150 16435 1170
rect 16455 1150 16460 1170
rect 16430 1120 16460 1150
rect 16430 1100 16435 1120
rect 16455 1100 16460 1120
rect 16430 1070 16460 1100
rect 16430 1050 16435 1070
rect 16455 1050 16460 1070
rect 16430 1020 16460 1050
rect 16430 1000 16435 1020
rect 16455 1000 16460 1020
rect 16430 970 16460 1000
rect 16430 950 16435 970
rect 16455 950 16460 970
rect 16430 940 16460 950
rect 16485 1170 16515 1180
rect 16485 1150 16490 1170
rect 16510 1150 16515 1170
rect 16485 1120 16515 1150
rect 16485 1100 16490 1120
rect 16510 1100 16515 1120
rect 16485 1070 16515 1100
rect 16485 1050 16490 1070
rect 16510 1050 16515 1070
rect 16485 1020 16515 1050
rect 16485 1000 16490 1020
rect 16510 1000 16515 1020
rect 16485 970 16515 1000
rect 16485 950 16490 970
rect 16510 950 16515 970
rect 16485 940 16515 950
rect 16540 1170 16570 1180
rect 16540 1150 16545 1170
rect 16565 1150 16570 1170
rect 16540 1120 16570 1150
rect 16540 1100 16545 1120
rect 16565 1100 16570 1120
rect 16540 1070 16570 1100
rect 16540 1050 16545 1070
rect 16565 1050 16570 1070
rect 16540 1020 16570 1050
rect 16540 1000 16545 1020
rect 16565 1000 16570 1020
rect 16540 970 16570 1000
rect 16540 950 16545 970
rect 16565 950 16570 970
rect 16540 940 16570 950
rect 16595 1170 16625 1180
rect 16595 1150 16600 1170
rect 16620 1150 16625 1170
rect 16595 1120 16625 1150
rect 16595 1100 16600 1120
rect 16620 1100 16625 1120
rect 16595 1070 16625 1100
rect 16595 1050 16600 1070
rect 16620 1050 16625 1070
rect 16595 1020 16625 1050
rect 16595 1000 16600 1020
rect 16620 1000 16625 1020
rect 16595 970 16625 1000
rect 16595 950 16600 970
rect 16620 950 16625 970
rect 16595 940 16625 950
rect 16650 1170 16680 1180
rect 16650 1150 16655 1170
rect 16675 1150 16680 1170
rect 16650 1120 16680 1150
rect 16650 1100 16655 1120
rect 16675 1100 16680 1120
rect 16650 1070 16680 1100
rect 16650 1050 16655 1070
rect 16675 1050 16680 1070
rect 16650 1020 16680 1050
rect 16650 1000 16655 1020
rect 16675 1000 16680 1020
rect 16650 970 16680 1000
rect 16650 950 16655 970
rect 16675 950 16680 970
rect 16650 940 16680 950
rect 16705 1170 16735 1180
rect 16705 1150 16710 1170
rect 16730 1150 16735 1170
rect 16705 1120 16735 1150
rect 16705 1100 16710 1120
rect 16730 1100 16735 1120
rect 16705 1070 16735 1100
rect 16705 1050 16710 1070
rect 16730 1050 16735 1070
rect 16705 1020 16735 1050
rect 16705 1000 16710 1020
rect 16730 1000 16735 1020
rect 16705 970 16735 1000
rect 16705 950 16710 970
rect 16730 950 16735 970
rect 16705 940 16735 950
rect 16760 1170 16790 1180
rect 16760 1150 16765 1170
rect 16785 1150 16790 1170
rect 16760 1120 16790 1150
rect 16760 1100 16765 1120
rect 16785 1100 16790 1120
rect 16760 1070 16790 1100
rect 16760 1050 16765 1070
rect 16785 1050 16790 1070
rect 16760 1020 16790 1050
rect 16760 1000 16765 1020
rect 16785 1000 16790 1020
rect 16760 970 16790 1000
rect 16760 950 16765 970
rect 16785 950 16790 970
rect 16760 940 16790 950
rect 16815 1170 16845 1180
rect 16815 1150 16820 1170
rect 16840 1150 16845 1170
rect 16815 1120 16845 1150
rect 16815 1100 16820 1120
rect 16840 1100 16845 1120
rect 16815 1070 16845 1100
rect 16815 1050 16820 1070
rect 16840 1050 16845 1070
rect 16815 1020 16845 1050
rect 16815 1000 16820 1020
rect 16840 1000 16845 1020
rect 16815 970 16845 1000
rect 16815 950 16820 970
rect 16840 950 16845 970
rect 16815 940 16845 950
rect 16870 1170 16900 1180
rect 16870 1150 16875 1170
rect 16895 1150 16900 1170
rect 16870 1120 16900 1150
rect 16870 1100 16875 1120
rect 16895 1100 16900 1120
rect 16870 1070 16900 1100
rect 16870 1050 16875 1070
rect 16895 1050 16900 1070
rect 16870 1020 16900 1050
rect 16870 1000 16875 1020
rect 16895 1000 16900 1020
rect 16870 970 16900 1000
rect 16870 950 16875 970
rect 16895 950 16900 970
rect 16870 940 16900 950
rect 16925 1170 16955 1180
rect 16925 1150 16930 1170
rect 16950 1150 16955 1170
rect 16925 1120 16955 1150
rect 16925 1100 16930 1120
rect 16950 1100 16955 1120
rect 16925 1070 16955 1100
rect 16925 1050 16930 1070
rect 16950 1050 16955 1070
rect 16925 1020 16955 1050
rect 16925 1000 16930 1020
rect 16950 1000 16955 1020
rect 16925 970 16955 1000
rect 16925 950 16930 970
rect 16950 950 16955 970
rect 16925 940 16955 950
rect 16980 1170 17010 1180
rect 16980 1150 16985 1170
rect 17005 1150 17010 1170
rect 16980 1120 17010 1150
rect 16980 1100 16985 1120
rect 17005 1100 17010 1120
rect 16980 1070 17010 1100
rect 16980 1050 16985 1070
rect 17005 1050 17010 1070
rect 16980 1020 17010 1050
rect 16980 1000 16985 1020
rect 17005 1000 17010 1020
rect 16980 970 17010 1000
rect 16980 950 16985 970
rect 17005 950 17010 970
rect 16980 940 17010 950
rect 17035 1170 17065 1180
rect 17035 1150 17040 1170
rect 17060 1150 17065 1170
rect 17035 1120 17065 1150
rect 17035 1100 17040 1120
rect 17060 1100 17065 1120
rect 17035 1070 17065 1100
rect 17035 1050 17040 1070
rect 17060 1050 17065 1070
rect 17035 1020 17065 1050
rect 17035 1000 17040 1020
rect 17060 1000 17065 1020
rect 17035 970 17065 1000
rect 17035 950 17040 970
rect 17060 950 17065 970
rect 17035 940 17065 950
rect 17090 1170 17120 1180
rect 17090 1150 17095 1170
rect 17115 1150 17120 1170
rect 17090 1120 17120 1150
rect 17090 1100 17095 1120
rect 17115 1100 17120 1120
rect 17090 1070 17120 1100
rect 17090 1050 17095 1070
rect 17115 1050 17120 1070
rect 17090 1020 17120 1050
rect 17090 1000 17095 1020
rect 17115 1000 17120 1020
rect 17090 970 17120 1000
rect 17090 950 17095 970
rect 17115 950 17120 970
rect 17090 940 17120 950
rect 17145 1170 17175 1180
rect 17145 1150 17150 1170
rect 17170 1150 17175 1170
rect 17145 1120 17175 1150
rect 17145 1100 17150 1120
rect 17170 1100 17175 1120
rect 17145 1070 17175 1100
rect 17145 1050 17150 1070
rect 17170 1050 17175 1070
rect 17145 1020 17175 1050
rect 17145 1000 17150 1020
rect 17170 1000 17175 1020
rect 17145 970 17175 1000
rect 17145 950 17150 970
rect 17170 950 17175 970
rect 17145 940 17175 950
rect 17200 1170 17230 1180
rect 17200 1150 17205 1170
rect 17225 1150 17230 1170
rect 17200 1120 17230 1150
rect 17200 1100 17205 1120
rect 17225 1100 17230 1120
rect 17200 1070 17230 1100
rect 17200 1050 17205 1070
rect 17225 1050 17230 1070
rect 17200 1020 17230 1050
rect 17200 1000 17205 1020
rect 17225 1000 17230 1020
rect 17200 970 17230 1000
rect 17200 950 17205 970
rect 17225 950 17230 970
rect 17200 940 17230 950
rect 17255 1170 17285 1180
rect 17255 1150 17260 1170
rect 17280 1150 17285 1170
rect 17255 1120 17285 1150
rect 17255 1100 17260 1120
rect 17280 1100 17285 1120
rect 17255 1070 17285 1100
rect 17255 1050 17260 1070
rect 17280 1050 17285 1070
rect 17255 1020 17285 1050
rect 17255 1000 17260 1020
rect 17280 1000 17285 1020
rect 17255 970 17285 1000
rect 17255 950 17260 970
rect 17280 950 17285 970
rect 17255 940 17285 950
rect 17310 1170 17340 1180
rect 17310 1150 17315 1170
rect 17335 1150 17340 1170
rect 17310 1120 17340 1150
rect 17310 1100 17315 1120
rect 17335 1100 17340 1120
rect 17310 1070 17340 1100
rect 17310 1050 17315 1070
rect 17335 1050 17340 1070
rect 17310 1020 17340 1050
rect 17310 1000 17315 1020
rect 17335 1000 17340 1020
rect 17310 970 17340 1000
rect 17310 950 17315 970
rect 17335 950 17340 970
rect 17310 940 17340 950
rect 17365 1170 17395 1180
rect 17365 1150 17370 1170
rect 17390 1150 17395 1170
rect 17365 1120 17395 1150
rect 17365 1100 17370 1120
rect 17390 1100 17395 1120
rect 17365 1070 17395 1100
rect 17365 1050 17370 1070
rect 17390 1050 17395 1070
rect 17365 1020 17395 1050
rect 17365 1000 17370 1020
rect 17390 1000 17395 1020
rect 17365 970 17395 1000
rect 17365 950 17370 970
rect 17390 950 17395 970
rect 17365 940 17395 950
rect 17420 1170 17450 1180
rect 17420 1150 17425 1170
rect 17445 1150 17450 1170
rect 17420 1120 17450 1150
rect 17420 1100 17425 1120
rect 17445 1100 17450 1120
rect 17420 1070 17450 1100
rect 17420 1050 17425 1070
rect 17445 1050 17450 1070
rect 17420 1020 17450 1050
rect 17420 1000 17425 1020
rect 17445 1000 17450 1020
rect 17420 970 17450 1000
rect 17420 950 17425 970
rect 17445 950 17450 970
rect 17420 940 17450 950
rect 17475 1170 17505 1180
rect 17475 1150 17480 1170
rect 17500 1150 17505 1170
rect 17475 1120 17505 1150
rect 17475 1100 17480 1120
rect 17500 1100 17505 1120
rect 17475 1070 17505 1100
rect 17475 1050 17480 1070
rect 17500 1050 17505 1070
rect 17475 1020 17505 1050
rect 17475 1000 17480 1020
rect 17500 1000 17505 1020
rect 17475 970 17505 1000
rect 17475 950 17480 970
rect 17500 950 17505 970
rect 17475 940 17505 950
rect 17530 1170 17560 1180
rect 17530 1150 17535 1170
rect 17555 1150 17560 1170
rect 17530 1120 17560 1150
rect 17530 1100 17535 1120
rect 17555 1100 17560 1120
rect 17530 1070 17560 1100
rect 17530 1050 17535 1070
rect 17555 1050 17560 1070
rect 17530 1020 17560 1050
rect 17530 1000 17535 1020
rect 17555 1000 17560 1020
rect 17530 970 17560 1000
rect 17530 950 17535 970
rect 17555 950 17560 970
rect 17530 940 17560 950
rect 17585 1170 17655 1180
rect 17585 1150 17590 1170
rect 17610 1150 17630 1170
rect 17650 1150 17655 1170
rect 17585 1120 17655 1150
rect 17585 1100 17590 1120
rect 17610 1100 17630 1120
rect 17650 1100 17655 1120
rect 17585 1070 17655 1100
rect 17585 1050 17590 1070
rect 17610 1050 17630 1070
rect 17650 1050 17655 1070
rect 17585 1020 17655 1050
rect 17585 1000 17590 1020
rect 17610 1000 17630 1020
rect 17650 1000 17655 1020
rect 17585 970 17655 1000
rect 17585 950 17590 970
rect 17610 950 17630 970
rect 17650 950 17655 970
rect 17970 1170 17975 1190
rect 17995 1170 18015 1190
rect 18035 1170 18040 1190
rect 17970 1140 18040 1170
rect 17970 1120 17975 1140
rect 17995 1120 18015 1140
rect 18035 1120 18040 1140
rect 17970 1090 18040 1120
rect 17970 1070 17975 1090
rect 17995 1070 18015 1090
rect 18035 1070 18040 1090
rect 17970 1040 18040 1070
rect 17970 1020 17975 1040
rect 17995 1020 18015 1040
rect 18035 1020 18040 1040
rect 17970 990 18040 1020
rect 17970 970 17975 990
rect 17995 970 18015 990
rect 18035 970 18040 990
rect 17970 960 18040 970
rect 18110 1640 18140 1650
rect 18110 1620 18115 1640
rect 18135 1620 18140 1640
rect 18110 1590 18140 1620
rect 18110 1570 18115 1590
rect 18135 1570 18140 1590
rect 18110 1540 18140 1570
rect 18110 1520 18115 1540
rect 18135 1520 18140 1540
rect 18110 1490 18140 1520
rect 18110 1470 18115 1490
rect 18135 1470 18140 1490
rect 18110 1440 18140 1470
rect 18110 1420 18115 1440
rect 18135 1420 18140 1440
rect 18110 1390 18140 1420
rect 18110 1370 18115 1390
rect 18135 1370 18140 1390
rect 18110 1340 18140 1370
rect 18110 1320 18115 1340
rect 18135 1320 18140 1340
rect 18110 1290 18140 1320
rect 18110 1270 18115 1290
rect 18135 1270 18140 1290
rect 18110 1240 18140 1270
rect 18110 1220 18115 1240
rect 18135 1220 18140 1240
rect 18110 1190 18140 1220
rect 18110 1170 18115 1190
rect 18135 1170 18140 1190
rect 18110 1140 18140 1170
rect 18110 1120 18115 1140
rect 18135 1120 18140 1140
rect 18110 1090 18140 1120
rect 18110 1070 18115 1090
rect 18135 1070 18140 1090
rect 18110 1040 18140 1070
rect 18110 1020 18115 1040
rect 18135 1020 18140 1040
rect 18110 990 18140 1020
rect 18110 970 18115 990
rect 18135 970 18140 990
rect 18110 960 18140 970
rect 18210 1640 18240 1650
rect 18210 1620 18215 1640
rect 18235 1620 18240 1640
rect 18210 1590 18240 1620
rect 18210 1570 18215 1590
rect 18235 1570 18240 1590
rect 18210 1540 18240 1570
rect 18210 1520 18215 1540
rect 18235 1520 18240 1540
rect 18210 1490 18240 1520
rect 18210 1470 18215 1490
rect 18235 1470 18240 1490
rect 18210 1440 18240 1470
rect 18210 1420 18215 1440
rect 18235 1420 18240 1440
rect 18210 1390 18240 1420
rect 18210 1370 18215 1390
rect 18235 1370 18240 1390
rect 18210 1340 18240 1370
rect 18210 1320 18215 1340
rect 18235 1320 18240 1340
rect 18210 1290 18240 1320
rect 18210 1270 18215 1290
rect 18235 1270 18240 1290
rect 18210 1240 18240 1270
rect 18210 1220 18215 1240
rect 18235 1220 18240 1240
rect 18210 1190 18240 1220
rect 18210 1170 18215 1190
rect 18235 1170 18240 1190
rect 18210 1140 18240 1170
rect 18210 1120 18215 1140
rect 18235 1120 18240 1140
rect 18210 1090 18240 1120
rect 18210 1070 18215 1090
rect 18235 1070 18240 1090
rect 18210 1040 18240 1070
rect 18210 1020 18215 1040
rect 18235 1020 18240 1040
rect 18210 990 18240 1020
rect 18210 970 18215 990
rect 18235 970 18240 990
rect 18210 960 18240 970
rect 18310 1640 18340 1650
rect 18310 1620 18315 1640
rect 18335 1620 18340 1640
rect 18310 1590 18340 1620
rect 18310 1570 18315 1590
rect 18335 1570 18340 1590
rect 18310 1540 18340 1570
rect 18310 1520 18315 1540
rect 18335 1520 18340 1540
rect 18310 1490 18340 1520
rect 18310 1470 18315 1490
rect 18335 1470 18340 1490
rect 18310 1440 18340 1470
rect 18310 1420 18315 1440
rect 18335 1420 18340 1440
rect 18310 1390 18340 1420
rect 18310 1370 18315 1390
rect 18335 1370 18340 1390
rect 18310 1340 18340 1370
rect 18310 1320 18315 1340
rect 18335 1320 18340 1340
rect 18310 1290 18340 1320
rect 18310 1270 18315 1290
rect 18335 1270 18340 1290
rect 18310 1240 18340 1270
rect 18310 1220 18315 1240
rect 18335 1220 18340 1240
rect 18310 1190 18340 1220
rect 18310 1170 18315 1190
rect 18335 1170 18340 1190
rect 18310 1140 18340 1170
rect 18310 1120 18315 1140
rect 18335 1120 18340 1140
rect 18310 1090 18340 1120
rect 18310 1070 18315 1090
rect 18335 1070 18340 1090
rect 18310 1040 18340 1070
rect 18310 1020 18315 1040
rect 18335 1020 18340 1040
rect 18310 990 18340 1020
rect 18310 970 18315 990
rect 18335 970 18340 990
rect 18310 960 18340 970
rect 18410 1640 18440 1650
rect 18410 1620 18415 1640
rect 18435 1620 18440 1640
rect 18410 1590 18440 1620
rect 18410 1570 18415 1590
rect 18435 1570 18440 1590
rect 18410 1540 18440 1570
rect 18410 1520 18415 1540
rect 18435 1520 18440 1540
rect 18410 1490 18440 1520
rect 18410 1470 18415 1490
rect 18435 1470 18440 1490
rect 18410 1440 18440 1470
rect 18410 1420 18415 1440
rect 18435 1420 18440 1440
rect 18410 1390 18440 1420
rect 18410 1370 18415 1390
rect 18435 1370 18440 1390
rect 18410 1340 18440 1370
rect 18410 1320 18415 1340
rect 18435 1320 18440 1340
rect 18410 1290 18440 1320
rect 18410 1270 18415 1290
rect 18435 1270 18440 1290
rect 18410 1240 18440 1270
rect 18410 1220 18415 1240
rect 18435 1220 18440 1240
rect 18410 1190 18440 1220
rect 18410 1170 18415 1190
rect 18435 1170 18440 1190
rect 18410 1140 18440 1170
rect 18410 1120 18415 1140
rect 18435 1120 18440 1140
rect 18410 1090 18440 1120
rect 18410 1070 18415 1090
rect 18435 1070 18440 1090
rect 18410 1040 18440 1070
rect 18410 1020 18415 1040
rect 18435 1020 18440 1040
rect 18410 990 18440 1020
rect 18410 970 18415 990
rect 18435 970 18440 990
rect 18410 960 18440 970
rect 18510 1640 18540 1650
rect 18510 1620 18515 1640
rect 18535 1620 18540 1640
rect 18510 1590 18540 1620
rect 18510 1570 18515 1590
rect 18535 1570 18540 1590
rect 18510 1540 18540 1570
rect 18510 1520 18515 1540
rect 18535 1520 18540 1540
rect 18510 1490 18540 1520
rect 18510 1470 18515 1490
rect 18535 1470 18540 1490
rect 18510 1440 18540 1470
rect 18510 1420 18515 1440
rect 18535 1420 18540 1440
rect 18510 1390 18540 1420
rect 18510 1370 18515 1390
rect 18535 1370 18540 1390
rect 18510 1340 18540 1370
rect 18510 1320 18515 1340
rect 18535 1320 18540 1340
rect 18510 1290 18540 1320
rect 18510 1270 18515 1290
rect 18535 1270 18540 1290
rect 18510 1240 18540 1270
rect 18510 1220 18515 1240
rect 18535 1220 18540 1240
rect 18510 1190 18540 1220
rect 18510 1170 18515 1190
rect 18535 1170 18540 1190
rect 18510 1140 18540 1170
rect 18510 1120 18515 1140
rect 18535 1120 18540 1140
rect 18510 1090 18540 1120
rect 18510 1070 18515 1090
rect 18535 1070 18540 1090
rect 18510 1040 18540 1070
rect 18510 1020 18515 1040
rect 18535 1020 18540 1040
rect 18510 990 18540 1020
rect 18510 970 18515 990
rect 18535 970 18540 990
rect 18510 960 18540 970
rect 18610 1640 18680 1650
rect 18610 1620 18615 1640
rect 18635 1620 18655 1640
rect 18675 1620 18680 1640
rect 18610 1590 18680 1620
rect 18610 1570 18615 1590
rect 18635 1570 18655 1590
rect 18675 1570 18680 1590
rect 18610 1540 18680 1570
rect 18610 1520 18615 1540
rect 18635 1520 18655 1540
rect 18675 1520 18680 1540
rect 18610 1490 18680 1520
rect 18610 1470 18615 1490
rect 18635 1470 18655 1490
rect 18675 1470 18680 1490
rect 18610 1440 18680 1470
rect 18610 1420 18615 1440
rect 18635 1420 18655 1440
rect 18675 1420 18680 1440
rect 18610 1390 18680 1420
rect 18610 1370 18615 1390
rect 18635 1370 18655 1390
rect 18675 1370 18680 1390
rect 18735 1640 18770 1650
rect 18735 1615 18740 1640
rect 18765 1615 18770 1640
rect 18735 1605 18770 1615
rect 18795 1640 18830 1650
rect 18795 1615 18800 1640
rect 18825 1615 18830 1640
rect 18795 1605 18830 1615
rect 18610 1340 18680 1370
rect 18610 1320 18615 1340
rect 18635 1320 18655 1340
rect 18675 1320 18680 1340
rect 18610 1290 18680 1320
rect 18610 1270 18615 1290
rect 18635 1270 18655 1290
rect 18675 1270 18680 1290
rect 18610 1240 18680 1270
rect 18610 1220 18615 1240
rect 18635 1220 18655 1240
rect 18675 1220 18680 1240
rect 18610 1190 18680 1220
rect 18610 1170 18615 1190
rect 18635 1170 18655 1190
rect 18675 1170 18680 1190
rect 18610 1140 18680 1170
rect 18610 1120 18615 1140
rect 18635 1120 18655 1140
rect 18675 1120 18680 1140
rect 18610 1090 18680 1120
rect 18610 1070 18615 1090
rect 18635 1070 18655 1090
rect 18675 1070 18680 1090
rect 18610 1040 18680 1070
rect 18610 1020 18615 1040
rect 18635 1020 18655 1040
rect 18675 1020 18680 1040
rect 18610 990 18680 1020
rect 18610 970 18615 990
rect 18635 970 18655 990
rect 18675 970 18680 990
rect 18610 960 18680 970
rect 17585 940 17655 950
rect 17975 940 17995 960
rect 18215 940 18235 960
rect 18415 940 18435 960
rect 18655 940 18675 960
rect 15115 930 15155 940
rect 15115 910 15125 930
rect 15145 910 15155 930
rect 4975 895 5015 905
rect 15115 900 15155 910
rect 15355 930 15395 940
rect 15355 910 15365 930
rect 15385 910 15395 930
rect 15355 900 15395 910
rect 15555 930 15595 940
rect 15555 910 15565 930
rect 15585 910 15595 930
rect 15555 900 15595 910
rect 15795 930 15835 940
rect 15795 910 15805 930
rect 15825 910 15835 930
rect 16175 920 16195 940
rect 16270 920 16290 940
rect 16380 920 16400 940
rect 16490 920 16510 940
rect 16600 920 16620 940
rect 16710 920 16730 940
rect 16820 920 16840 940
rect 16930 920 16950 940
rect 17040 920 17060 940
rect 17150 920 17170 940
rect 17260 920 17280 940
rect 17370 920 17390 940
rect 17480 920 17500 940
rect 17630 920 17650 940
rect 17965 930 18005 940
rect 15795 900 15835 910
rect 16165 910 16205 920
rect 3005 875 3025 895
rect 3185 875 3205 895
rect 3365 875 3385 895
rect 3545 875 3565 895
rect 3725 875 3745 895
rect 3905 875 3925 895
rect 4085 875 4105 895
rect 4265 875 4285 895
rect 4445 875 4465 895
rect 4625 875 4645 895
rect 4805 875 4825 895
rect 4985 875 5005 895
rect 16165 890 16175 910
rect 16195 890 16205 910
rect 16165 880 16205 890
rect 16260 910 16300 920
rect 16260 890 16270 910
rect 16290 890 16300 910
rect 16260 880 16300 890
rect 16370 910 16410 920
rect 16370 890 16380 910
rect 16400 890 16410 910
rect 16370 880 16410 890
rect 16480 910 16520 920
rect 16480 890 16490 910
rect 16510 890 16520 910
rect 16480 880 16520 890
rect 16590 910 16630 920
rect 16590 890 16600 910
rect 16620 890 16630 910
rect 16590 880 16630 890
rect 16700 910 16740 920
rect 16700 890 16710 910
rect 16730 890 16740 910
rect 16700 880 16740 890
rect 16810 910 16850 920
rect 16810 890 16820 910
rect 16840 890 16850 910
rect 16810 880 16850 890
rect 16920 910 16960 920
rect 16920 890 16930 910
rect 16950 890 16960 910
rect 16920 880 16960 890
rect 17030 910 17070 920
rect 17030 890 17040 910
rect 17060 890 17070 910
rect 17030 880 17070 890
rect 17140 910 17180 920
rect 17140 890 17150 910
rect 17170 890 17180 910
rect 17140 880 17180 890
rect 17250 910 17290 920
rect 17250 890 17260 910
rect 17280 890 17290 910
rect 17250 880 17290 890
rect 17360 910 17400 920
rect 17360 890 17370 910
rect 17390 890 17400 910
rect 17360 880 17400 890
rect 17470 910 17510 920
rect 17470 890 17480 910
rect 17500 890 17510 910
rect 17470 880 17510 890
rect 17620 910 17660 920
rect 17620 890 17630 910
rect 17650 890 17660 910
rect 17965 910 17975 930
rect 17995 910 18005 930
rect 17965 900 18005 910
rect 18205 930 18245 940
rect 18205 910 18215 930
rect 18235 910 18245 930
rect 18205 900 18245 910
rect 18405 930 18445 940
rect 18405 910 18415 930
rect 18435 910 18445 930
rect 18405 900 18445 910
rect 18645 930 18685 940
rect 18645 910 18655 930
rect 18675 910 18685 930
rect 18770 910 18795 960
rect 18645 900 18685 910
rect 17620 880 17660 890
rect 2960 865 3030 875
rect 2960 845 2965 865
rect 2985 845 3005 865
rect 3025 845 3030 865
rect 2960 815 3030 845
rect 2960 795 2965 815
rect 2985 795 3005 815
rect 3025 795 3030 815
rect 2960 785 3030 795
rect 3090 865 3120 875
rect 3090 845 3095 865
rect 3115 845 3120 865
rect 3090 815 3120 845
rect 3090 795 3095 815
rect 3115 795 3120 815
rect 3090 785 3120 795
rect 3180 865 3210 875
rect 3180 845 3185 865
rect 3205 845 3210 865
rect 3180 815 3210 845
rect 3180 795 3185 815
rect 3205 795 3210 815
rect 3180 785 3210 795
rect 3270 865 3300 875
rect 3270 845 3275 865
rect 3295 845 3300 865
rect 3270 815 3300 845
rect 3270 795 3275 815
rect 3295 795 3300 815
rect 3270 785 3300 795
rect 3360 865 3390 875
rect 3360 845 3365 865
rect 3385 845 3390 865
rect 3360 815 3390 845
rect 3360 795 3365 815
rect 3385 795 3390 815
rect 3360 785 3390 795
rect 3450 865 3480 875
rect 3450 845 3455 865
rect 3475 845 3480 865
rect 3450 815 3480 845
rect 3450 795 3455 815
rect 3475 795 3480 815
rect 3450 785 3480 795
rect 3540 865 3570 875
rect 3540 845 3545 865
rect 3565 845 3570 865
rect 3540 815 3570 845
rect 3540 795 3545 815
rect 3565 795 3570 815
rect 3540 785 3570 795
rect 3630 865 3660 875
rect 3630 845 3635 865
rect 3655 845 3660 865
rect 3630 815 3660 845
rect 3630 795 3635 815
rect 3655 795 3660 815
rect 3630 785 3660 795
rect 3720 865 3750 875
rect 3720 845 3725 865
rect 3745 845 3750 865
rect 3720 815 3750 845
rect 3720 795 3725 815
rect 3745 795 3750 815
rect 3720 785 3750 795
rect 3810 865 3840 875
rect 3810 845 3815 865
rect 3835 845 3840 865
rect 3810 815 3840 845
rect 3810 795 3815 815
rect 3835 795 3840 815
rect 3810 785 3840 795
rect 3900 865 3930 875
rect 3900 845 3905 865
rect 3925 845 3930 865
rect 3900 815 3930 845
rect 3900 795 3905 815
rect 3925 795 3930 815
rect 3900 785 3930 795
rect 3990 865 4020 875
rect 3990 845 3995 865
rect 4015 845 4020 865
rect 3990 815 4020 845
rect 3990 795 3995 815
rect 4015 795 4020 815
rect 3990 785 4020 795
rect 4080 865 4110 875
rect 4080 845 4085 865
rect 4105 845 4110 865
rect 4080 815 4110 845
rect 4080 795 4085 815
rect 4105 795 4110 815
rect 4080 785 4110 795
rect 4170 865 4200 875
rect 4170 845 4175 865
rect 4195 845 4200 865
rect 4170 815 4200 845
rect 4170 795 4175 815
rect 4195 795 4200 815
rect 4170 785 4200 795
rect 4260 865 4290 875
rect 4260 845 4265 865
rect 4285 845 4290 865
rect 4260 815 4290 845
rect 4260 795 4265 815
rect 4285 795 4290 815
rect 4260 785 4290 795
rect 4350 865 4380 875
rect 4350 845 4355 865
rect 4375 845 4380 865
rect 4350 815 4380 845
rect 4350 795 4355 815
rect 4375 795 4380 815
rect 4350 785 4380 795
rect 4440 865 4470 875
rect 4440 845 4445 865
rect 4465 845 4470 865
rect 4440 815 4470 845
rect 4440 795 4445 815
rect 4465 795 4470 815
rect 4440 785 4470 795
rect 4530 865 4560 875
rect 4530 845 4535 865
rect 4555 845 4560 865
rect 4530 815 4560 845
rect 4530 795 4535 815
rect 4555 795 4560 815
rect 4530 785 4560 795
rect 4620 865 4650 875
rect 4620 845 4625 865
rect 4645 845 4650 865
rect 4620 815 4650 845
rect 4620 795 4625 815
rect 4645 795 4650 815
rect 4620 785 4650 795
rect 4710 865 4740 875
rect 4710 845 4715 865
rect 4735 845 4740 865
rect 4710 815 4740 845
rect 4710 795 4715 815
rect 4735 795 4740 815
rect 4710 785 4740 795
rect 4800 865 4830 875
rect 4800 845 4805 865
rect 4825 845 4830 865
rect 4800 815 4830 845
rect 4800 795 4805 815
rect 4825 795 4830 815
rect 4800 785 4830 795
rect 4890 865 4920 875
rect 4890 845 4895 865
rect 4915 845 4920 865
rect 4890 815 4920 845
rect 4890 795 4895 815
rect 4915 795 4920 815
rect 4890 785 4920 795
rect 4980 865 5050 875
rect 4980 845 4985 865
rect 5005 845 5025 865
rect 5045 845 5050 865
rect 4980 815 5050 845
rect 16010 825 16040 855
rect 16495 820 16535 860
rect 16940 830 16970 860
rect 17160 830 17190 860
rect 17380 830 17410 860
rect 17865 830 17895 860
rect 4980 795 4985 815
rect 5005 795 5025 815
rect 5045 795 5050 815
rect 4980 785 5050 795
rect 3095 765 3115 785
rect 3275 765 3295 785
rect 3455 765 3475 785
rect 3635 765 3655 785
rect 3815 765 3835 785
rect 3995 765 4015 785
rect 4175 765 4195 785
rect 4355 765 4375 785
rect 4535 765 4555 785
rect 4715 765 4735 785
rect 4895 765 4915 785
rect 15955 765 15985 795
rect 16305 790 16345 800
rect 16305 780 16315 790
rect 16275 770 16315 780
rect 16335 770 16345 790
rect 2525 730 2555 760
rect 3095 755 3170 765
rect 3095 745 3140 755
rect 3130 735 3140 745
rect 3160 735 3170 755
rect 3130 725 3170 735
rect 3265 755 3305 765
rect 3265 735 3275 755
rect 3295 735 3305 755
rect 3265 725 3305 735
rect 3445 755 3485 765
rect 3445 735 3455 755
rect 3475 735 3485 755
rect 3445 725 3485 735
rect 3625 755 3665 765
rect 3625 735 3635 755
rect 3655 735 3665 755
rect 3625 725 3665 735
rect 3805 755 3845 765
rect 3805 735 3815 755
rect 3835 735 3845 755
rect 3805 725 3845 735
rect 3985 755 4025 765
rect 3985 735 3995 755
rect 4015 735 4025 755
rect 3985 725 4025 735
rect 4165 755 4205 765
rect 4165 735 4175 755
rect 4195 735 4205 755
rect 4165 725 4205 735
rect 4345 755 4385 765
rect 4345 735 4355 755
rect 4375 735 4385 755
rect 4345 725 4385 735
rect 4525 755 4565 765
rect 4525 735 4535 755
rect 4555 735 4565 755
rect 4525 725 4565 735
rect 4705 755 4745 765
rect 4705 735 4715 755
rect 4735 735 4745 755
rect 4705 725 4745 735
rect 4885 755 4925 765
rect 4885 735 4895 755
rect 4915 735 4925 755
rect 16275 760 16345 770
rect 16375 790 16415 800
rect 16375 770 16385 790
rect 16405 770 16415 790
rect 16375 760 16415 770
rect 16445 790 16485 800
rect 16445 770 16455 790
rect 16475 770 16485 790
rect 16445 760 16485 770
rect 16275 740 16295 760
rect 16505 740 16525 820
rect 16935 795 16975 805
rect 16935 775 16945 795
rect 16965 775 16975 795
rect 16935 765 16975 775
rect 17045 795 17085 805
rect 17045 775 17055 795
rect 17075 775 17085 795
rect 17045 765 17085 775
rect 17155 795 17195 805
rect 17155 775 17165 795
rect 17185 775 17195 795
rect 17155 765 17195 775
rect 17265 795 17305 805
rect 17265 775 17275 795
rect 17295 775 17305 795
rect 17265 765 17305 775
rect 17375 795 17415 805
rect 17375 775 17385 795
rect 17405 775 17415 795
rect 17375 765 17415 775
rect 17485 795 17525 805
rect 17485 775 17495 795
rect 17515 775 17525 795
rect 17485 765 17525 775
rect 17810 770 17840 800
rect 16945 745 16965 765
rect 17055 745 17075 765
rect 17165 745 17185 765
rect 17275 745 17295 765
rect 17385 745 17405 765
rect 17495 745 17515 765
rect 4885 725 4925 735
rect 16265 730 16295 740
rect 16265 710 16270 730
rect 16290 710 16295 730
rect 3450 675 3480 705
rect 3810 675 3840 705
rect 4170 675 4200 705
rect 16265 680 16295 710
rect 16265 660 16270 680
rect 16290 660 16295 680
rect 16265 650 16295 660
rect 16495 730 16525 740
rect 16495 710 16500 730
rect 16520 710 16525 730
rect 16495 680 16525 710
rect 16845 735 16915 745
rect 16845 715 16850 735
rect 16870 715 16890 735
rect 16910 715 16915 735
rect 16845 705 16915 715
rect 16940 735 16970 745
rect 16940 715 16945 735
rect 16965 715 16970 735
rect 16940 705 16970 715
rect 16995 735 17025 745
rect 16995 715 17000 735
rect 17020 715 17025 735
rect 16995 705 17025 715
rect 17050 735 17080 745
rect 17050 715 17055 735
rect 17075 715 17080 735
rect 17050 705 17080 715
rect 17105 735 17135 745
rect 17105 715 17110 735
rect 17130 715 17135 735
rect 17105 705 17135 715
rect 17160 735 17190 745
rect 17160 715 17165 735
rect 17185 715 17190 735
rect 17160 705 17190 715
rect 17215 735 17245 745
rect 17215 715 17220 735
rect 17240 715 17245 735
rect 17215 705 17245 715
rect 17270 735 17300 745
rect 17270 715 17275 735
rect 17295 715 17300 735
rect 17270 705 17300 715
rect 17325 735 17355 745
rect 17325 715 17330 735
rect 17350 715 17355 735
rect 17325 705 17355 715
rect 17380 735 17410 745
rect 17380 715 17385 735
rect 17405 715 17410 735
rect 17380 705 17410 715
rect 17435 735 17465 745
rect 17435 715 17440 735
rect 17460 715 17465 735
rect 17435 705 17465 715
rect 17490 735 17520 745
rect 17490 715 17495 735
rect 17515 715 17520 735
rect 17490 705 17520 715
rect 17545 735 17615 745
rect 17545 715 17550 735
rect 17570 715 17590 735
rect 17610 715 17615 735
rect 17545 705 17615 715
rect 16850 685 16870 705
rect 17000 685 17020 705
rect 17110 685 17130 705
rect 17220 685 17240 705
rect 17330 685 17350 705
rect 17440 685 17460 705
rect 17590 685 17610 705
rect 16495 660 16500 680
rect 16520 660 16525 680
rect 16495 650 16525 660
rect 16840 675 16880 685
rect 16840 655 16850 675
rect 16870 655 16880 675
rect 16840 645 16880 655
rect 16990 675 17030 685
rect 16990 655 17000 675
rect 17020 655 17030 675
rect 16990 645 17030 655
rect 17100 675 17140 685
rect 17100 655 17110 675
rect 17130 655 17140 675
rect 17100 645 17140 655
rect 17210 675 17250 685
rect 17210 655 17220 675
rect 17240 655 17250 675
rect 17210 645 17250 655
rect 17320 675 17360 685
rect 17320 655 17330 675
rect 17350 655 17360 675
rect 17320 645 17360 655
rect 17430 675 17470 685
rect 17430 655 17440 675
rect 17460 655 17470 675
rect 17430 645 17470 655
rect 17580 675 17620 685
rect 17580 655 17590 675
rect 17610 655 17620 675
rect 17580 645 17620 655
<< viali >>
rect 16640 4490 16660 4510
rect 16760 4490 16780 4510
rect 16880 4490 16900 4510
rect 16210 4430 16230 4450
rect 16470 4430 16490 4450
rect 16580 4445 16600 4465
rect 16700 4445 16720 4465
rect 16820 4445 16840 4465
rect 16940 4445 16960 4465
rect 17090 4420 17110 4440
rect 17210 4420 17230 4440
rect 17330 4420 17350 4440
rect 17450 4420 17470 4440
rect 17570 4420 17590 4440
rect 16340 4315 16360 4320
rect 16340 4295 16360 4315
rect 16760 4290 16780 4310
rect 17150 4290 17170 4310
rect 17211 4290 17229 4310
rect 17270 4290 17290 4310
rect 17390 4290 17410 4310
rect 17510 4290 17530 4310
rect 16370 4180 16390 4200
rect 16480 4180 16500 4200
rect 16590 4180 16610 4200
rect 16700 4180 16720 4200
rect 16810 4180 16830 4200
rect 16920 4180 16940 4200
rect 17030 4180 17050 4200
rect 17140 4180 17160 4200
rect 17250 4180 17270 4200
rect 17360 4180 17380 4200
rect 16315 4060 16335 4080
rect 16370 4060 16390 4080
rect 16425 4060 16445 4080
rect 16535 4060 16555 4080
rect 16645 4060 16665 4080
rect 16755 4060 16775 4080
rect 16865 4060 16885 4080
rect 16975 4060 16995 4080
rect 17085 4060 17105 4080
rect 17195 4060 17215 4080
rect 17305 4060 17325 4080
rect 17415 4060 17435 4080
rect 16320 3935 16340 3955
rect 16425 3935 16445 3955
rect 16535 3935 16555 3955
rect 16645 3935 16665 3955
rect 16755 3935 16775 3955
rect 17060 3935 17080 3955
rect 17165 3935 17185 3955
rect 17275 3935 17295 3955
rect 17385 3935 17405 3955
rect 17495 3935 17515 3955
rect 16277 3875 16294 3895
rect 16370 3875 16390 3895
rect 16480 3875 16500 3895
rect 16700 3875 16720 3895
rect 16810 3875 16830 3895
rect 17017 3875 17034 3895
rect 17220 3875 17240 3895
rect 17440 3875 17460 3895
rect 16408 3755 16425 3775
rect 16628 3755 16645 3775
rect 16775 3755 16792 3775
rect 16260 3695 16280 3715
rect 16365 3695 16385 3715
rect 16480 3695 16500 3715
rect 16585 3695 16605 3715
rect 16700 3695 16720 3715
rect 16815 3695 16835 3715
rect 17000 3705 17020 3725
rect 17148 3755 17165 3775
rect 17220 3705 17240 3725
rect 17368 3755 17385 3775
rect 17515 3755 17532 3775
rect 17440 3705 17460 3725
rect 15220 3610 15240 3630
rect 15330 3610 15350 3630
rect 15440 3610 15460 3630
rect 15550 3610 15570 3630
rect 15660 3610 15680 3630
rect 15770 3610 15790 3630
rect 16350 3600 16370 3620
rect 16470 3600 16490 3620
rect 16590 3600 16610 3620
rect 16710 3600 16730 3620
rect 16830 3600 16850 3620
rect 16950 3600 16970 3620
rect 17070 3600 17090 3620
rect 17190 3600 17210 3620
rect 17310 3600 17330 3620
rect 17430 3600 17450 3620
rect 18010 3610 18030 3630
rect 18120 3610 18140 3630
rect 18230 3610 18250 3630
rect 18340 3610 18360 3630
rect 18450 3610 18470 3630
rect 18560 3610 18580 3630
rect 56 3175 81 3200
rect 1271 3170 1296 3195
rect 56 3115 81 3140
rect 1271 3110 1296 3135
rect 56 3035 81 3060
rect 56 2975 81 3000
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 2340 2930 2365 2955
rect 3090 2955 3110 2975
rect 3145 2955 3165 2975
rect 3275 2955 3295 2975
rect 3455 2955 3475 2975
rect 3635 2955 3655 2975
rect 3815 2955 3835 2975
rect 3995 2955 4015 2975
rect 4175 2955 4195 2975
rect 4355 2955 4375 2975
rect 4535 2955 4555 2975
rect 4715 2955 4735 2975
rect 4845 2955 4865 2975
rect 4895 2955 4915 2975
rect 16290 3130 16310 3150
rect 16410 3130 16430 3150
rect 16530 3130 16550 3150
rect 16650 3130 16670 3150
rect 16770 3130 16790 3150
rect 16831 3130 16849 3150
rect 16890 3130 16910 3150
rect 17010 3130 17030 3150
rect 17130 3130 17150 3150
rect 17250 3130 17270 3150
rect 17370 3130 17390 3150
rect 17490 3130 17510 3150
rect 2340 2870 2365 2895
rect 61 2825 86 2850
rect 734 2825 759 2850
rect 1271 2810 1296 2835
rect 1970 2810 1995 2835
rect 15275 2940 15295 2960
rect 15385 2940 15405 2960
rect 15495 2940 15515 2960
rect 15605 2940 15625 2960
rect 15661 2940 15679 2960
rect 15715 2940 15735 2960
rect 16350 2920 16370 2940
rect 16470 2920 16490 2940
rect 16590 2920 16610 2940
rect 16710 2920 16730 2940
rect 16830 2920 16850 2940
rect 16950 2920 16970 2940
rect 17070 2920 17090 2940
rect 17190 2920 17210 2940
rect 17310 2920 17330 2940
rect 17430 2920 17450 2940
rect 18065 2940 18085 2960
rect 18121 2940 18139 2960
rect 18175 2940 18195 2960
rect 18285 2940 18305 2960
rect 18395 2940 18415 2960
rect 18505 2940 18525 2960
rect 61 2765 86 2790
rect 734 2765 759 2790
rect 3005 2785 3025 2805
rect 3185 2785 3205 2805
rect 3365 2785 3385 2805
rect 3545 2785 3565 2805
rect 3725 2785 3745 2805
rect 3905 2785 3925 2805
rect 4085 2785 4105 2805
rect 4265 2785 4285 2805
rect 4445 2785 4465 2805
rect 4625 2785 4645 2805
rect 4805 2785 4825 2805
rect 4985 2785 5005 2805
rect 3185 2725 3205 2745
rect 3365 2725 3385 2745
rect 3545 2725 3565 2745
rect 3725 2725 3745 2745
rect 3905 2725 3925 2745
rect 4085 2725 4105 2745
rect 4265 2725 4285 2745
rect 4445 2725 4465 2745
rect 4625 2725 4645 2745
rect 4805 2725 4825 2745
rect 15220 2680 15240 2700
rect 15330 2680 15350 2700
rect 15440 2680 15460 2700
rect 15550 2680 15570 2700
rect 15660 2680 15680 2700
rect 15770 2680 15790 2700
rect 18010 2680 18030 2700
rect 18120 2680 18140 2700
rect 18230 2680 18250 2700
rect 18340 2680 18360 2700
rect 18450 2680 18470 2700
rect 18560 2680 18580 2700
rect 16290 2450 16310 2470
rect 16410 2450 16430 2470
rect 16530 2450 16550 2470
rect 16650 2450 16670 2470
rect 16770 2450 16790 2470
rect 16831 2450 16849 2470
rect 16890 2450 16910 2470
rect 17010 2450 17030 2470
rect 17130 2450 17150 2470
rect 17250 2450 17270 2470
rect 17370 2450 17390 2470
rect 17490 2450 17510 2470
rect 3275 2355 3295 2375
rect 3365 2350 3385 2370
rect 3455 2355 3475 2375
rect 3815 2355 3835 2375
rect 3895 2355 3915 2375
rect 3995 2355 4015 2375
rect 4175 2355 4195 2375
rect 15275 2410 15295 2430
rect 15385 2410 15405 2430
rect 15495 2410 15515 2430
rect 15605 2410 15625 2430
rect 15715 2410 15735 2430
rect 18065 2410 18085 2430
rect 18175 2410 18195 2430
rect 18285 2410 18305 2430
rect 18395 2410 18415 2430
rect 18505 2410 18525 2430
rect 4535 2355 4555 2375
rect 4715 2355 4735 2375
rect 15775 2365 15795 2385
rect 18035 2350 18055 2370
rect 3635 2310 3655 2330
rect 4355 2310 4375 2330
rect 3455 2265 3475 2285
rect 4535 2265 4555 2285
rect 15275 2290 15295 2310
rect 15385 2290 15405 2310
rect 15495 2290 15515 2310
rect 15605 2290 15625 2310
rect 15715 2290 15735 2310
rect 18065 2290 18085 2310
rect 18175 2290 18195 2310
rect 18285 2290 18305 2310
rect 18395 2290 18415 2310
rect 18505 2290 18525 2310
rect 2755 2070 2775 2090
rect 2875 2070 2895 2090
rect 2995 2070 3015 2090
rect 3115 2070 3135 2090
rect 3235 2070 3255 2090
rect 3355 2070 3375 2090
rect 3475 2070 3495 2090
rect 3595 2070 3615 2090
rect 3715 2070 3735 2090
rect 3835 2070 3855 2090
rect 3995 2070 4015 2090
rect 4155 2070 4175 2090
rect 4275 2070 4295 2090
rect 4395 2070 4415 2090
rect 4515 2070 4535 2090
rect 4635 2070 4655 2090
rect 4755 2070 4775 2090
rect 4875 2070 4895 2090
rect 4995 2070 5015 2090
rect 5115 2070 5135 2090
rect 5235 2070 5255 2090
rect 2630 2025 2650 2045
rect -35 1695 -15 1715
rect 2815 2025 2835 2045
rect 3175 2025 3195 2045
rect 3535 2025 3555 2045
rect 3895 2025 3915 2045
rect 4095 2025 4115 2045
rect 4455 2025 4475 2045
rect 4815 2025 4835 2045
rect 5175 2025 5195 2045
rect 14795 1975 14820 2000
rect 14855 1975 14880 2000
rect 14915 1975 14940 2000
rect 14975 1975 15000 2000
rect 16340 2155 16360 2175
rect 16450 2155 16470 2175
rect 16560 2155 16580 2175
rect 16670 2155 16690 2175
rect 16780 2155 16800 2175
rect 16836 2155 16854 2175
rect 16890 2155 16910 2175
rect 17000 2155 17020 2175
rect 17110 2155 17130 2175
rect 17220 2155 17240 2175
rect 17330 2155 17350 2175
rect 17440 2155 17460 2175
rect 18800 1975 18825 2000
rect 15220 1920 15238 1940
rect 15330 1920 15348 1940
rect 15440 1920 15458 1940
rect 15550 1920 15568 1940
rect 15660 1920 15678 1940
rect 15770 1920 15788 1940
rect 16395 1935 16415 1955
rect 16505 1935 16525 1955
rect 16615 1935 16635 1955
rect 16725 1935 16745 1955
rect 16835 1935 16855 1955
rect 16945 1935 16965 1955
rect 17055 1935 17075 1955
rect 17165 1935 17185 1955
rect 17275 1935 17295 1955
rect 17385 1935 17405 1955
rect 18860 1975 18885 2000
rect 18920 1975 18945 2000
rect 18980 1975 19005 2000
rect 18012 1920 18030 1940
rect 18122 1920 18140 1940
rect 18232 1920 18250 1940
rect 18342 1920 18360 1940
rect 18452 1920 18470 1940
rect 18562 1920 18580 1940
rect 2575 1855 2595 1875
rect 2630 1855 2650 1875
rect 2685 1855 2705 1875
rect 2845 1855 2865 1875
rect 2935 1855 2955 1875
rect 3055 1855 3075 1875
rect 3175 1855 3195 1875
rect 3295 1855 3315 1875
rect 3415 1855 3435 1875
rect 3535 1855 3555 1875
rect 3655 1855 3675 1875
rect 3775 1855 3795 1875
rect 3865 1855 3885 1875
rect 4125 1855 4145 1875
rect 4215 1855 4235 1875
rect 4335 1855 4355 1875
rect 4455 1855 4475 1875
rect 4575 1855 4595 1875
rect 4695 1855 4715 1875
rect 4815 1855 4835 1875
rect 4935 1855 4955 1875
rect 5055 1855 5075 1875
rect 5145 1855 5165 1875
rect 3055 1795 3075 1815
rect 3415 1795 3435 1815
rect 3775 1795 3795 1815
rect 4215 1795 4235 1815
rect 4575 1795 4595 1815
rect 4935 1795 4955 1815
rect 3235 1735 3255 1755
rect 3295 1735 3315 1755
rect 3535 1735 3555 1755
rect 3775 1735 3795 1755
rect 4215 1735 4235 1755
rect 4455 1735 4475 1755
rect 4695 1735 4715 1755
rect 4755 1735 4775 1755
rect 16095 1735 16115 1755
rect 16200 1750 16220 1770
rect 3175 1690 3195 1710
rect 3415 1690 3435 1710
rect 3655 1690 3675 1710
rect 4335 1690 4355 1710
rect 4575 1690 4595 1710
rect 4815 1690 4835 1710
rect 15265 1680 15285 1700
rect 15465 1680 15485 1700
rect 15566 1680 15584 1700
rect 15665 1680 15685 1700
rect 3995 1630 4015 1650
rect 16315 1735 16335 1755
rect 16420 1750 16440 1770
rect 16243 1690 16260 1710
rect 16535 1735 16555 1755
rect 16650 1750 16670 1770
rect 16463 1690 16480 1710
rect 16610 1690 16627 1710
rect 17135 1735 17155 1755
rect 17240 1750 17260 1770
rect 16825 1690 16845 1710
rect 16876 1690 16893 1710
rect 16955 1690 16975 1710
rect 17355 1735 17375 1755
rect 17460 1750 17480 1770
rect 17283 1690 17300 1710
rect 17575 1735 17595 1755
rect 17690 1750 17710 1770
rect 17503 1690 17520 1710
rect 17650 1690 17667 1710
rect 18115 1680 18135 1700
rect 18216 1680 18234 1700
rect 18315 1680 18335 1700
rect 18515 1680 18535 1700
rect 3175 1570 3195 1590
rect 14975 1615 15000 1640
rect 4815 1570 4835 1590
rect 3235 1520 3255 1540
rect 3355 1520 3375 1540
rect 3475 1520 3495 1540
rect 3595 1520 3615 1540
rect 3715 1520 3735 1540
rect 4275 1520 4295 1540
rect 4395 1520 4415 1540
rect 4515 1520 4535 1540
rect 4635 1520 4655 1540
rect 4755 1520 4775 1540
rect 2845 1460 2865 1480
rect 2935 1475 2955 1495
rect 3055 1475 3075 1495
rect 3175 1475 3195 1495
rect 3295 1475 3315 1495
rect 3535 1475 3555 1495
rect 3655 1475 3675 1495
rect 3775 1475 3795 1495
rect 3925 1460 3945 1480
rect 4065 1460 4085 1480
rect 4215 1475 4235 1495
rect 4335 1475 4355 1495
rect 4455 1475 4475 1495
rect 4695 1475 4715 1495
rect 4815 1475 4835 1495
rect 4935 1475 4955 1495
rect 5055 1475 5075 1495
rect 5145 1460 5165 1480
rect 15035 1615 15060 1640
rect 3385 1160 3405 1180
rect 4605 1160 4625 1180
rect 2955 1100 2975 1120
rect 3035 1100 3055 1120
rect 3115 1100 3135 1120
rect 3195 1100 3215 1120
rect 3275 1100 3295 1120
rect 3355 1100 3375 1120
rect 3435 1100 3455 1120
rect 3515 1100 3535 1120
rect 3595 1100 3615 1120
rect 3675 1100 3695 1120
rect 3755 1100 3775 1120
rect 3835 1100 3855 1120
rect 3915 1100 3935 1120
rect 3995 1100 4015 1120
rect 4075 1100 4095 1120
rect 4155 1100 4175 1120
rect 4235 1100 4255 1120
rect 4315 1100 4335 1120
rect 4395 1100 4415 1120
rect 4475 1100 4495 1120
rect 4555 1100 4575 1120
rect 4635 1100 4655 1120
rect 4715 1100 4735 1120
rect 4795 1100 4815 1120
rect 4875 1100 4895 1120
rect 4955 1100 4975 1120
rect 2915 1015 2935 1035
rect 5120 1015 5140 1035
rect 3005 905 3025 925
rect 3185 905 3205 925
rect 3365 905 3385 925
rect 3545 905 3565 925
rect 3725 905 3745 925
rect 3905 905 3925 925
rect 4085 905 4105 925
rect 4265 905 4285 925
rect 4445 905 4465 925
rect 4625 905 4645 925
rect 4805 905 4825 925
rect 4985 905 5005 925
rect 16112 1470 16129 1490
rect 16315 1470 16335 1490
rect 16535 1470 16555 1490
rect 16830 1470 16850 1490
rect 16880 1470 16900 1490
rect 16928 1470 16945 1490
rect 17152 1470 17169 1490
rect 17355 1470 17375 1490
rect 17575 1470 17595 1490
rect 16155 1410 16175 1430
rect 16260 1410 16280 1430
rect 16370 1410 16390 1430
rect 16480 1410 16500 1430
rect 16590 1410 16610 1430
rect 17195 1410 17215 1430
rect 17300 1410 17320 1430
rect 17410 1410 17430 1430
rect 17520 1410 17540 1430
rect 17630 1410 17650 1430
rect 16325 1210 16345 1230
rect 16435 1210 16455 1230
rect 16545 1210 16565 1230
rect 16655 1210 16675 1230
rect 16765 1210 16785 1230
rect 16820 1210 16840 1230
rect 16875 1210 16895 1230
rect 16985 1210 17005 1230
rect 17095 1210 17115 1230
rect 17205 1210 17225 1230
rect 17315 1210 17335 1230
rect 17425 1210 17445 1230
rect 17535 1210 17555 1230
rect 17605 1225 17625 1245
rect 18740 1615 18765 1640
rect 18800 1615 18825 1640
rect 15365 910 15385 930
rect 15565 910 15585 930
rect 16175 890 16195 910
rect 16270 890 16290 910
rect 16380 890 16400 910
rect 16490 890 16510 910
rect 16600 890 16620 910
rect 16710 890 16730 910
rect 16820 890 16840 910
rect 16930 890 16950 910
rect 17040 890 17060 910
rect 17150 890 17170 910
rect 17260 890 17280 910
rect 17370 890 17390 910
rect 17480 890 17500 910
rect 17630 890 17650 910
rect 18215 910 18235 930
rect 18415 910 18435 930
rect 16315 770 16335 790
rect 3140 735 3160 755
rect 3275 735 3295 755
rect 3455 735 3475 755
rect 3635 735 3655 755
rect 3815 735 3835 755
rect 3995 735 4015 755
rect 4175 735 4195 755
rect 4355 735 4375 755
rect 4535 735 4555 755
rect 4715 735 4735 755
rect 4895 735 4915 755
rect 16385 770 16405 790
rect 16455 770 16475 790
rect 16945 775 16965 795
rect 17055 775 17075 795
rect 17165 775 17185 795
rect 17275 775 17295 795
rect 17385 775 17405 795
rect 17495 775 17515 795
rect 17000 655 17020 675
rect 17110 655 17130 675
rect 17220 655 17240 675
rect 17330 655 17350 675
rect 17440 655 17460 675
<< metal1 >>
rect 16632 4515 16668 4520
rect 16632 4485 16635 4515
rect 16665 4485 16668 4515
rect 16632 4480 16668 4485
rect 16752 4515 16788 4520
rect 16752 4485 16755 4515
rect 16785 4485 16788 4515
rect 16752 4480 16788 4485
rect 16872 4515 16908 4520
rect 16872 4485 16875 4515
rect 16905 4485 16908 4515
rect 16872 4480 16908 4485
rect 17080 4515 17120 4520
rect 17080 4485 17085 4515
rect 17115 4485 17120 4515
rect 17080 4480 17120 4485
rect 16570 4470 16610 4475
rect 16200 4455 16240 4460
rect 16200 4425 16205 4455
rect 16235 4425 16240 4455
rect 16200 4420 16240 4425
rect 16460 4455 16500 4460
rect 16460 4425 16465 4455
rect 16495 4425 16500 4455
rect 16570 4440 16575 4470
rect 16605 4440 16610 4470
rect 16570 4435 16610 4440
rect 16690 4470 16730 4475
rect 16690 4440 16695 4470
rect 16725 4440 16730 4470
rect 16690 4435 16730 4440
rect 16810 4470 16850 4475
rect 16810 4440 16815 4470
rect 16845 4440 16850 4470
rect 16810 4435 16850 4440
rect 16930 4470 16970 4475
rect 16930 4440 16935 4470
rect 16965 4440 16970 4470
rect 17090 4450 17110 4480
rect 16930 4435 16970 4440
rect 17080 4445 17120 4450
rect 16460 4420 16500 4425
rect 17080 4415 17085 4445
rect 17115 4415 17120 4445
rect 17080 4410 17120 4415
rect 17200 4445 17240 4450
rect 17200 4415 17205 4445
rect 17235 4415 17240 4445
rect 17200 4410 17240 4415
rect 17320 4445 17360 4450
rect 17320 4415 17325 4445
rect 17355 4415 17360 4445
rect 17320 4410 17360 4415
rect 17440 4445 17480 4450
rect 17440 4415 17445 4445
rect 17475 4415 17480 4445
rect 17440 4410 17480 4415
rect 17560 4445 17600 4450
rect 17560 4415 17565 4445
rect 17595 4415 17600 4445
rect 17560 4410 17600 4415
rect 16330 4320 16370 4325
rect 16050 4315 16090 4320
rect 16050 4285 16055 4315
rect 16085 4285 16090 4315
rect 16330 4290 16335 4320
rect 16365 4290 16370 4320
rect 16330 4285 16370 4290
rect 16750 4315 16790 4320
rect 16750 4285 16755 4315
rect 16785 4285 16790 4315
rect 16050 4280 16090 4285
rect 14955 3635 14995 3640
rect 14955 3605 14960 3635
rect 14990 3605 14995 3635
rect 14955 3600 14995 3605
rect 15210 3635 15250 3640
rect 15210 3605 15215 3635
rect 15245 3605 15250 3635
rect 15210 3600 15250 3605
rect 15320 3635 15360 3640
rect 15320 3605 15325 3635
rect 15355 3605 15360 3635
rect 15320 3600 15360 3605
rect 15430 3635 15470 3640
rect 15430 3605 15435 3635
rect 15465 3605 15470 3635
rect 15430 3600 15470 3605
rect 15540 3635 15580 3640
rect 15540 3605 15545 3635
rect 15575 3605 15580 3635
rect 15540 3600 15580 3605
rect 15650 3635 15690 3640
rect 15650 3605 15655 3635
rect 15685 3605 15690 3635
rect 15650 3600 15690 3605
rect 15760 3635 15800 3640
rect 15760 3605 15765 3635
rect 15795 3605 15800 3635
rect 15760 3600 15800 3605
rect 14965 3560 14985 3600
rect 14904 3555 15045 3560
rect 1261 3525 1301 3530
rect 1261 3495 1266 3525
rect 1296 3495 1301 3525
rect 14904 3525 14910 3555
rect 14940 3525 14960 3555
rect 14990 3525 15010 3555
rect 15040 3525 15045 3555
rect 14904 3520 15045 3525
rect 1261 3490 1301 3495
rect 4440 3495 4480 3500
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3415 25 3445
rect -15 3410 25 3415
rect 940 3445 980 3450
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3360 -20 3390
rect -60 3355 -20 3360
rect -50 2860 -30 3355
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2825 -20 2855
rect -60 2820 -20 2825
rect -5 2800 15 3410
rect 1205 3340 1245 3345
rect 1205 3310 1210 3340
rect 1240 3310 1245 3340
rect 1205 3305 1245 3310
rect 1160 3285 1200 3290
rect 1160 3255 1165 3285
rect 1195 3255 1200 3285
rect 1160 3250 1200 3255
rect 46 3170 51 3205
rect 86 3170 91 3205
rect 46 3110 51 3145
rect 86 3110 91 3145
rect 1170 3105 1190 3250
rect 1160 3100 1200 3105
rect 1160 3070 1165 3100
rect 1195 3070 1200 3100
rect 1160 3065 1200 3070
rect 46 3030 51 3065
rect 86 3030 91 3065
rect 46 2970 51 3005
rect 86 2970 91 3005
rect 905 2910 1125 2920
rect 905 2880 920 2910
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 905 2870 1125 2880
rect 1215 2855 1235 3305
rect 1271 3200 1291 3490
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 1635 3445 1685 3455
rect 1635 3415 1645 3445
rect 1675 3415 1685 3445
rect 2470 3450 2510 3455
rect 2470 3420 2475 3450
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 1635 3405 1685 3415
rect 1261 3165 1266 3200
rect 1301 3165 1306 3200
rect 1271 3140 1291 3165
rect 1261 3105 1266 3140
rect 1301 3105 1306 3140
rect 2330 2925 2335 2960
rect 2370 2925 2375 2960
rect 2425 2955 2465 2960
rect 2425 2925 2430 2955
rect 2460 2925 2465 2955
rect 2425 2920 2465 2925
rect 2330 2900 2375 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 2330 2860 2375 2865
rect 51 2820 56 2855
rect 91 2820 96 2855
rect 724 2820 729 2855
rect 764 2820 769 2855
rect 1205 2850 1245 2855
rect 1205 2820 1210 2850
rect 1240 2820 1245 2850
rect 2340 2840 2360 2860
rect 1205 2815 1245 2820
rect 1261 2805 1266 2840
rect 1301 2805 1306 2840
rect 1960 2805 1965 2840
rect 2000 2805 2005 2840
rect 2330 2835 2370 2840
rect 2330 2805 2335 2835
rect 2365 2805 2370 2835
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2765 25 2795
rect -15 2760 25 2765
rect 51 2760 56 2795
rect 91 2760 96 2795
rect 724 2760 729 2795
rect 764 2760 769 2795
rect 1271 2750 1291 2805
rect 2330 2800 2370 2805
rect 1261 2745 1301 2750
rect 1261 2715 1266 2745
rect 1296 2715 1301 2745
rect 1261 2710 1301 2715
rect 2150 2745 2190 2750
rect 2150 2715 2155 2745
rect 2185 2715 2190 2745
rect 2150 2710 2190 2715
rect 275 2200 1985 2550
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1715 -70 1720
rect -45 1720 -5 1725
rect -45 1715 -40 1720
rect -75 1695 -40 1715
rect -75 1690 -70 1695
rect -110 1685 -70 1690
rect -45 1690 -40 1695
rect -10 1690 -5 1720
rect -45 1685 -5 1690
rect 275 1190 625 2200
rect 952 1710 1302 1870
rect 952 1680 1270 1710
rect 1297 1680 1302 1710
rect 952 1520 1302 1680
rect 1330 1190 1455 1345
rect 1635 1190 1985 2200
rect 2160 1190 2180 2710
rect 2340 2205 2360 2800
rect 2435 2250 2455 2920
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2215 2465 2245
rect 2425 2210 2465 2215
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2170 2370 2200
rect 2330 2165 2370 2170
rect 2340 1600 2360 2165
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2120 2420 2150
rect 2380 2115 2420 2120
rect 2390 1670 2410 2115
rect 2435 1765 2455 2210
rect 2480 1825 2500 3415
rect 2690 3390 2730 3395
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3135 3340 3175 3345
rect 3135 3310 3140 3340
rect 3170 3310 3175 3340
rect 3135 3305 3175 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3305 3435 3335
rect 2735 3240 2775 3245
rect 2735 3210 2740 3240
rect 2770 3210 2775 3240
rect 2735 3205 2775 3210
rect 2620 3185 2660 3190
rect 2620 3155 2625 3185
rect 2655 3155 2660 3185
rect 2620 3150 2660 3155
rect 2520 2980 2560 2985
rect 2520 2950 2525 2980
rect 2555 2950 2560 2980
rect 2520 2945 2560 2950
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1790 2510 1820
rect 2470 1785 2510 1790
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1730 2465 1760
rect 2425 1725 2465 1730
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1635 2420 1665
rect 2380 1630 2420 1635
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1565 2370 1595
rect 2330 1560 2370 1565
rect 275 840 2180 1190
rect 2530 765 2550 2945
rect 2630 2795 2650 3150
rect 2620 2790 2660 2795
rect 2620 2760 2625 2790
rect 2655 2760 2660 2790
rect 2620 2755 2660 2760
rect 2630 2350 2650 2755
rect 2620 2345 2660 2350
rect 2620 2315 2625 2345
rect 2655 2315 2660 2345
rect 2620 2310 2660 2315
rect 2630 2055 2650 2310
rect 2745 2295 2765 3205
rect 3145 3145 3165 3305
rect 3385 3295 3435 3305
rect 4450 3190 4470 3460
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3415 5185 3445
rect 5135 3405 5185 3415
rect 5360 3335 5400 3340
rect 5360 3305 5365 3335
rect 5395 3305 5400 3335
rect 5360 3300 5400 3305
rect 4885 3285 4925 3290
rect 4885 3255 4890 3285
rect 4920 3255 4925 3285
rect 4885 3250 4925 3255
rect 4440 3185 4480 3190
rect 4440 3155 4445 3185
rect 4475 3155 4480 3185
rect 4440 3150 4480 3155
rect 3135 3140 3175 3145
rect 3135 3110 3140 3140
rect 3170 3110 3175 3140
rect 3135 3105 3175 3110
rect 4835 3140 4875 3145
rect 4835 3110 4840 3140
rect 4870 3110 4875 3140
rect 4835 3105 4875 3110
rect 3145 2985 3165 3105
rect 3985 3080 4025 3085
rect 3985 3050 3990 3080
rect 4020 3050 4025 3080
rect 3985 3045 4025 3050
rect 3445 3035 3485 3040
rect 3445 3005 3450 3035
rect 3480 3005 3485 3035
rect 3445 3000 3485 3005
rect 3805 3035 3845 3040
rect 3805 3005 3810 3035
rect 3840 3005 3845 3035
rect 3805 3000 3845 3005
rect 3455 2985 3475 3000
rect 3815 2985 3835 3000
rect 3995 2985 4015 3045
rect 4345 3035 4385 3040
rect 4345 3005 4350 3035
rect 4380 3005 4385 3035
rect 4345 3000 4385 3005
rect 4705 3035 4745 3040
rect 4705 3005 4710 3035
rect 4740 3005 4745 3035
rect 4705 3000 4745 3005
rect 4355 2985 4375 3000
rect 4715 2985 4735 3000
rect 4845 2985 4865 3105
rect 4895 2985 4915 3250
rect 5315 3140 5355 3145
rect 5315 3110 5320 3140
rect 5350 3110 5355 3140
rect 5315 3105 5355 3110
rect 3080 2980 3120 2985
rect 3080 2950 3085 2980
rect 3115 2950 3120 2980
rect 3080 2945 3120 2950
rect 3140 2975 3175 2985
rect 3140 2955 3145 2975
rect 3165 2955 3175 2975
rect 3140 2945 3175 2955
rect 3265 2980 3305 2985
rect 3265 2950 3270 2980
rect 3300 2950 3305 2980
rect 3265 2945 3305 2950
rect 3445 2975 3485 2985
rect 3445 2955 3455 2975
rect 3475 2955 3485 2975
rect 3445 2945 3485 2955
rect 3625 2980 3665 2985
rect 3625 2950 3630 2980
rect 3660 2950 3665 2980
rect 3625 2945 3665 2950
rect 3805 2975 3845 2985
rect 3805 2955 3815 2975
rect 3835 2955 3845 2975
rect 3805 2945 3845 2955
rect 3985 2975 4025 2985
rect 3985 2955 3995 2975
rect 4015 2955 4025 2975
rect 3985 2945 4025 2955
rect 4165 2980 4205 2985
rect 4165 2950 4170 2980
rect 4200 2950 4205 2980
rect 4165 2945 4205 2950
rect 4345 2975 4385 2985
rect 4345 2955 4355 2975
rect 4375 2955 4385 2975
rect 4345 2945 4385 2955
rect 4525 2980 4565 2985
rect 4525 2950 4530 2980
rect 4560 2950 4565 2980
rect 4525 2945 4565 2950
rect 4705 2975 4745 2985
rect 4705 2955 4715 2975
rect 4735 2955 4745 2975
rect 4705 2945 4745 2955
rect 4835 2975 4870 2985
rect 4835 2955 4845 2975
rect 4865 2955 4870 2975
rect 4835 2945 4870 2955
rect 4890 2975 4925 2985
rect 4890 2955 4895 2975
rect 4915 2955 4925 2975
rect 4890 2945 4925 2955
rect 2995 2810 3035 2815
rect 2995 2780 3000 2810
rect 3030 2780 3035 2810
rect 2995 2775 3035 2780
rect 3175 2810 3215 2815
rect 3175 2780 3180 2810
rect 3210 2780 3215 2810
rect 3175 2775 3215 2780
rect 3355 2810 3395 2815
rect 3355 2780 3360 2810
rect 3390 2780 3395 2810
rect 3355 2775 3395 2780
rect 3535 2810 3575 2815
rect 3535 2780 3540 2810
rect 3570 2780 3575 2810
rect 3535 2775 3575 2780
rect 3715 2810 3755 2815
rect 3715 2780 3720 2810
rect 3750 2780 3755 2810
rect 3715 2775 3755 2780
rect 3895 2810 3935 2815
rect 3895 2780 3900 2810
rect 3930 2780 3935 2810
rect 3895 2775 3935 2780
rect 4075 2810 4115 2815
rect 4075 2780 4080 2810
rect 4110 2780 4115 2810
rect 4075 2775 4115 2780
rect 4255 2810 4295 2815
rect 4255 2780 4260 2810
rect 4290 2780 4295 2810
rect 4255 2775 4295 2780
rect 4435 2810 4475 2815
rect 4435 2780 4440 2810
rect 4470 2780 4475 2810
rect 4435 2775 4475 2780
rect 4615 2810 4655 2815
rect 4615 2780 4620 2810
rect 4650 2780 4655 2810
rect 4615 2775 4655 2780
rect 4795 2810 4835 2815
rect 4795 2780 4800 2810
rect 4830 2780 4835 2810
rect 4795 2775 4835 2780
rect 4975 2810 5015 2815
rect 4975 2780 4980 2810
rect 5010 2780 5015 2810
rect 4975 2775 5015 2780
rect 4805 2755 4825 2775
rect 3175 2750 3215 2755
rect 3175 2720 3180 2750
rect 3210 2720 3215 2750
rect 3175 2715 3215 2720
rect 3355 2750 3395 2755
rect 3355 2720 3360 2750
rect 3390 2720 3395 2750
rect 3355 2715 3395 2720
rect 3535 2750 3575 2755
rect 3535 2720 3540 2750
rect 3570 2720 3575 2750
rect 3535 2715 3575 2720
rect 3715 2750 3755 2755
rect 3715 2720 3720 2750
rect 3750 2720 3755 2750
rect 3715 2715 3755 2720
rect 3895 2750 3935 2755
rect 3895 2720 3900 2750
rect 3930 2720 3935 2750
rect 3895 2715 3935 2720
rect 4075 2750 4115 2755
rect 4075 2720 4080 2750
rect 4110 2720 4115 2750
rect 4075 2715 4115 2720
rect 4255 2750 4295 2755
rect 4255 2720 4260 2750
rect 4290 2720 4295 2750
rect 4255 2715 4295 2720
rect 4435 2750 4475 2755
rect 4435 2720 4440 2750
rect 4470 2720 4475 2750
rect 4435 2715 4475 2720
rect 4615 2750 4655 2755
rect 4615 2720 4620 2750
rect 4650 2720 4655 2750
rect 4615 2715 4655 2720
rect 4795 2750 4835 2755
rect 4795 2720 4800 2750
rect 4830 2720 4835 2750
rect 4795 2715 4835 2720
rect 3265 2375 3305 2385
rect 3265 2355 3275 2375
rect 3295 2355 3305 2375
rect 3265 2345 3305 2355
rect 3355 2375 3395 2380
rect 3355 2345 3360 2375
rect 3390 2345 3395 2375
rect 3445 2375 3485 2385
rect 3445 2355 3455 2375
rect 3475 2355 3485 2375
rect 3445 2345 3485 2355
rect 3805 2380 3845 2385
rect 3805 2350 3810 2380
rect 3840 2350 3845 2380
rect 3805 2345 3845 2350
rect 3885 2375 3925 2385
rect 3885 2355 3895 2375
rect 3915 2355 3925 2375
rect 3885 2345 3925 2355
rect 3985 2375 4025 2385
rect 3985 2355 3995 2375
rect 4015 2355 4025 2375
rect 3985 2345 4025 2355
rect 4165 2380 4205 2385
rect 4165 2350 4170 2380
rect 4200 2350 4205 2380
rect 4165 2345 4205 2350
rect 4525 2375 4565 2385
rect 4525 2355 4535 2375
rect 4555 2355 4565 2375
rect 4525 2345 4565 2355
rect 4705 2375 4745 2385
rect 4705 2355 4715 2375
rect 4735 2355 4745 2375
rect 4705 2345 4745 2355
rect 2735 2290 2775 2295
rect 2735 2260 2740 2290
rect 2770 2260 2775 2290
rect 2735 2255 2775 2260
rect 3275 2205 3295 2345
rect 3355 2340 3395 2345
rect 3455 2295 3475 2345
rect 3625 2335 3665 2340
rect 3625 2305 3630 2335
rect 3660 2305 3665 2335
rect 3625 2300 3665 2305
rect 3445 2290 3485 2295
rect 3445 2260 3450 2290
rect 3480 2260 3485 2290
rect 3445 2255 3485 2260
rect 3265 2200 3305 2205
rect 3265 2170 3270 2200
rect 3300 2170 3305 2200
rect 3265 2165 3305 2170
rect 3635 2155 3655 2300
rect 3815 2250 3835 2345
rect 3805 2245 3845 2250
rect 3805 2215 3810 2245
rect 3840 2215 3845 2245
rect 3805 2210 3845 2215
rect 3625 2150 3665 2155
rect 3625 2120 3630 2150
rect 3660 2120 3665 2150
rect 3625 2115 3665 2120
rect 2745 2095 2785 2100
rect 2745 2065 2750 2095
rect 2780 2065 2785 2095
rect 2745 2060 2785 2065
rect 2865 2095 2905 2100
rect 2865 2065 2870 2095
rect 2900 2065 2905 2095
rect 2865 2060 2905 2065
rect 2985 2095 3025 2100
rect 2985 2065 2990 2095
rect 3020 2065 3025 2095
rect 2985 2060 3025 2065
rect 3105 2095 3145 2100
rect 3105 2065 3110 2095
rect 3140 2065 3145 2095
rect 3105 2060 3145 2065
rect 3225 2095 3265 2100
rect 3225 2065 3230 2095
rect 3260 2065 3265 2095
rect 3225 2060 3265 2065
rect 3345 2095 3385 2100
rect 3345 2065 3350 2095
rect 3380 2065 3385 2095
rect 3345 2060 3385 2065
rect 3465 2095 3505 2100
rect 3465 2065 3470 2095
rect 3500 2065 3505 2095
rect 3465 2060 3505 2065
rect 3585 2095 3625 2100
rect 3585 2065 3590 2095
rect 3620 2065 3625 2095
rect 3585 2060 3625 2065
rect 3705 2095 3745 2100
rect 3705 2065 3710 2095
rect 3740 2065 3745 2095
rect 3705 2060 3745 2065
rect 3825 2095 3865 2100
rect 3825 2065 3830 2095
rect 3860 2065 3865 2095
rect 3825 2060 3865 2065
rect 3895 2055 3915 2345
rect 3995 2205 4015 2345
rect 4345 2335 4385 2340
rect 4345 2305 4350 2335
rect 4380 2305 4385 2335
rect 4345 2300 4385 2305
rect 4535 2295 4555 2345
rect 4525 2290 4565 2295
rect 4525 2260 4530 2290
rect 4560 2260 4565 2290
rect 4525 2255 4565 2260
rect 4715 2205 4735 2345
rect 5270 2290 5310 2295
rect 5270 2260 5275 2290
rect 5305 2260 5310 2290
rect 5270 2255 5310 2260
rect 3985 2200 4025 2205
rect 3985 2170 3990 2200
rect 4020 2170 4025 2200
rect 3985 2165 4025 2170
rect 4705 2200 4745 2205
rect 4705 2170 4710 2200
rect 4740 2170 4745 2200
rect 4705 2165 4745 2170
rect 4085 2145 4125 2150
rect 4085 2115 4090 2145
rect 4120 2115 4125 2145
rect 4085 2110 4125 2115
rect 3985 2095 4025 2100
rect 3985 2065 3990 2095
rect 4020 2065 4025 2095
rect 3985 2060 4025 2065
rect 4095 2055 4115 2110
rect 4145 2095 4185 2100
rect 4145 2065 4150 2095
rect 4180 2065 4185 2095
rect 4145 2060 4185 2065
rect 4265 2095 4305 2100
rect 4265 2065 4270 2095
rect 4300 2065 4305 2095
rect 4265 2060 4305 2065
rect 4385 2095 4425 2100
rect 4385 2065 4390 2095
rect 4420 2065 4425 2095
rect 4385 2060 4425 2065
rect 4505 2095 4545 2100
rect 4505 2065 4510 2095
rect 4540 2065 4545 2095
rect 4505 2060 4545 2065
rect 4625 2095 4665 2100
rect 4625 2065 4630 2095
rect 4660 2065 4665 2095
rect 4625 2060 4665 2065
rect 4745 2095 4785 2100
rect 4745 2065 4750 2095
rect 4780 2065 4785 2095
rect 4745 2060 4785 2065
rect 4865 2095 4905 2100
rect 4865 2065 4870 2095
rect 4900 2065 4905 2095
rect 4865 2060 4905 2065
rect 4985 2095 5025 2100
rect 4985 2065 4990 2095
rect 5020 2065 5025 2095
rect 4985 2060 5025 2065
rect 5105 2095 5145 2100
rect 5105 2065 5110 2095
rect 5140 2065 5145 2095
rect 5105 2060 5145 2065
rect 5225 2095 5265 2100
rect 5225 2065 5230 2095
rect 5260 2065 5265 2095
rect 5225 2060 5265 2065
rect 2620 2050 2660 2055
rect 2620 2020 2625 2050
rect 2655 2020 2660 2050
rect 2620 2015 2660 2020
rect 2805 2050 2845 2055
rect 2805 2020 2810 2050
rect 2840 2020 2845 2050
rect 2805 2015 2845 2020
rect 3165 2050 3205 2055
rect 3165 2020 3170 2050
rect 3200 2020 3205 2050
rect 3165 2015 3205 2020
rect 3525 2050 3565 2055
rect 3525 2020 3530 2050
rect 3560 2020 3565 2050
rect 3525 2015 3565 2020
rect 3885 2050 3925 2055
rect 3885 2020 3890 2050
rect 3920 2045 3925 2050
rect 4085 2050 4125 2055
rect 4085 2045 4090 2050
rect 3920 2020 3945 2045
rect 3885 2015 3945 2020
rect 2565 1875 2600 1885
rect 2565 1855 2575 1875
rect 2595 1855 2600 1875
rect 2565 1845 2600 1855
rect 2620 1875 2660 1885
rect 2620 1855 2630 1875
rect 2650 1855 2660 1875
rect 2620 1845 2660 1855
rect 2680 1875 2715 1885
rect 2680 1855 2685 1875
rect 2705 1855 2715 1875
rect 2680 1845 2715 1855
rect 2835 1875 2875 1885
rect 2835 1855 2845 1875
rect 2865 1855 2875 1875
rect 2835 1845 2875 1855
rect 2925 1880 2965 1885
rect 2925 1850 2930 1880
rect 2960 1850 2965 1880
rect 2925 1845 2965 1850
rect 3045 1875 3085 1885
rect 3045 1855 3055 1875
rect 3075 1855 3085 1875
rect 3045 1845 3085 1855
rect 3165 1875 3205 1885
rect 3165 1855 3175 1875
rect 3195 1855 3205 1875
rect 3165 1845 3205 1855
rect 3285 1880 3325 1885
rect 3285 1850 3290 1880
rect 3320 1850 3325 1880
rect 3285 1845 3325 1850
rect 3405 1875 3445 1885
rect 3405 1855 3415 1875
rect 3435 1855 3445 1875
rect 3405 1845 3445 1855
rect 3525 1875 3565 1885
rect 3525 1855 3535 1875
rect 3555 1855 3565 1875
rect 3525 1845 3565 1855
rect 3645 1880 3685 1885
rect 3645 1850 3650 1880
rect 3680 1850 3685 1880
rect 3645 1845 3685 1850
rect 3765 1875 3805 1885
rect 3765 1855 3775 1875
rect 3795 1855 3805 1875
rect 3765 1845 3805 1855
rect 3855 1875 3895 1885
rect 3855 1855 3865 1875
rect 3885 1855 3895 1875
rect 3855 1845 3895 1855
rect 2575 1765 2595 1845
rect 2565 1760 2605 1765
rect 2565 1730 2570 1760
rect 2600 1730 2605 1760
rect 2565 1725 2605 1730
rect 2630 1670 2650 1845
rect 2685 1765 2705 1845
rect 2845 1825 2865 1845
rect 3055 1825 3075 1845
rect 3175 1825 3195 1845
rect 2835 1820 2875 1825
rect 2835 1790 2840 1820
rect 2870 1790 2875 1820
rect 2835 1785 2875 1790
rect 3045 1820 3085 1825
rect 3045 1790 3050 1820
rect 3080 1790 3085 1820
rect 3045 1785 3085 1790
rect 3165 1820 3205 1825
rect 3165 1790 3170 1820
rect 3200 1790 3205 1820
rect 3165 1785 3205 1790
rect 2800 1765 2840 1770
rect 3295 1765 3315 1845
rect 3415 1825 3435 1845
rect 3535 1825 3555 1845
rect 3775 1825 3795 1845
rect 3865 1825 3885 1845
rect 3405 1820 3445 1825
rect 3405 1790 3410 1820
rect 3440 1790 3445 1820
rect 3405 1785 3445 1790
rect 3525 1820 3565 1825
rect 3525 1790 3530 1820
rect 3560 1790 3565 1820
rect 3525 1785 3565 1790
rect 3765 1820 3805 1825
rect 3765 1790 3770 1820
rect 3800 1790 3805 1820
rect 3765 1785 3805 1790
rect 3855 1820 3895 1825
rect 3855 1790 3860 1820
rect 3890 1790 3895 1820
rect 3855 1785 3895 1790
rect 2675 1760 2715 1765
rect 2675 1730 2680 1760
rect 2710 1730 2715 1760
rect 2800 1735 2805 1765
rect 2835 1735 2840 1765
rect 2800 1730 2840 1735
rect 3225 1760 3265 1765
rect 3225 1730 3230 1760
rect 3260 1730 3265 1760
rect 2675 1725 2715 1730
rect 2810 1715 2830 1730
rect 3225 1725 3265 1730
rect 3285 1760 3325 1765
rect 3285 1730 3290 1760
rect 3320 1730 3325 1760
rect 3285 1725 3325 1730
rect 3415 1720 3435 1785
rect 3525 1760 3565 1765
rect 3525 1730 3530 1760
rect 3560 1730 3565 1760
rect 3525 1725 3565 1730
rect 3765 1760 3805 1765
rect 3765 1730 3770 1760
rect 3800 1730 3805 1760
rect 3765 1725 3805 1730
rect 3165 1715 3205 1720
rect 2800 1710 2840 1715
rect 2800 1680 2805 1710
rect 2835 1680 2840 1710
rect 3165 1685 3170 1715
rect 3200 1685 3205 1715
rect 3165 1680 3205 1685
rect 3405 1715 3445 1720
rect 3405 1685 3410 1715
rect 3440 1685 3445 1715
rect 3405 1680 3445 1685
rect 3645 1715 3685 1720
rect 3645 1685 3650 1715
rect 3680 1685 3685 1715
rect 3645 1680 3685 1685
rect 2800 1675 2840 1680
rect 2620 1665 2660 1670
rect 2620 1635 2625 1665
rect 2655 1635 2660 1665
rect 2620 1630 2660 1635
rect 2630 1045 2650 1630
rect 3165 1595 3205 1600
rect 3165 1565 3170 1595
rect 3200 1565 3205 1595
rect 3165 1560 3205 1565
rect 2835 1545 2875 1550
rect 2835 1515 2840 1545
rect 2870 1515 2875 1545
rect 2835 1510 2875 1515
rect 3225 1545 3265 1550
rect 3225 1515 3230 1545
rect 3260 1515 3265 1545
rect 3225 1510 3265 1515
rect 3345 1545 3385 1550
rect 3345 1515 3350 1545
rect 3380 1515 3385 1545
rect 3345 1510 3385 1515
rect 3465 1545 3505 1550
rect 3465 1515 3470 1545
rect 3500 1515 3505 1545
rect 3465 1510 3505 1515
rect 3585 1545 3625 1550
rect 3585 1515 3590 1545
rect 3620 1515 3625 1545
rect 3585 1510 3625 1515
rect 3705 1545 3745 1550
rect 3705 1515 3710 1545
rect 3740 1515 3745 1545
rect 3705 1510 3745 1515
rect 2845 1490 2865 1510
rect 2925 1500 2965 1505
rect 2835 1480 2875 1490
rect 2835 1460 2845 1480
rect 2865 1460 2875 1480
rect 2925 1470 2930 1500
rect 2960 1470 2965 1500
rect 2925 1465 2965 1470
rect 3045 1500 3085 1505
rect 3045 1470 3050 1500
rect 3080 1470 3085 1500
rect 3045 1465 3085 1470
rect 3165 1500 3205 1505
rect 3165 1470 3170 1500
rect 3200 1470 3205 1500
rect 3165 1465 3205 1470
rect 3285 1500 3325 1505
rect 3285 1470 3290 1500
rect 3320 1470 3325 1500
rect 3285 1465 3325 1470
rect 3525 1500 3565 1505
rect 3525 1470 3530 1500
rect 3560 1470 3565 1500
rect 3525 1465 3565 1470
rect 3645 1500 3685 1505
rect 3645 1470 3650 1500
rect 3680 1470 3685 1500
rect 3645 1465 3685 1470
rect 3765 1500 3805 1505
rect 3765 1470 3770 1500
rect 3800 1470 3805 1500
rect 3925 1490 3945 2015
rect 4065 2020 4090 2045
rect 4120 2020 4125 2050
rect 4065 2015 4125 2020
rect 4445 2050 4485 2055
rect 4445 2020 4450 2050
rect 4480 2020 4485 2050
rect 4445 2015 4485 2020
rect 4805 2050 4845 2055
rect 4805 2020 4810 2050
rect 4840 2020 4845 2050
rect 4805 2015 4845 2020
rect 5165 2050 5205 2055
rect 5165 2020 5170 2050
rect 5200 2020 5205 2050
rect 5165 2015 5205 2020
rect 3985 1650 4025 1660
rect 3985 1630 3995 1650
rect 4015 1630 4025 1650
rect 3985 1620 4025 1630
rect 3765 1465 3805 1470
rect 3915 1480 3955 1490
rect 2835 1450 2875 1460
rect 3915 1460 3925 1480
rect 3945 1460 3955 1480
rect 3915 1450 3955 1460
rect 3995 1190 4015 1620
rect 4065 1490 4085 2015
rect 4115 1875 4155 1885
rect 4115 1855 4125 1875
rect 4145 1855 4155 1875
rect 4115 1845 4155 1855
rect 4205 1875 4245 1885
rect 4205 1855 4215 1875
rect 4235 1855 4245 1875
rect 4205 1845 4245 1855
rect 4325 1880 4365 1885
rect 4325 1850 4330 1880
rect 4360 1850 4365 1880
rect 4325 1845 4365 1850
rect 4445 1875 4485 1885
rect 4445 1855 4455 1875
rect 4475 1855 4485 1875
rect 4445 1845 4485 1855
rect 4565 1875 4605 1885
rect 4565 1855 4575 1875
rect 4595 1855 4605 1875
rect 4565 1845 4605 1855
rect 4685 1880 4725 1885
rect 4685 1850 4690 1880
rect 4720 1850 4725 1880
rect 4685 1845 4725 1850
rect 4805 1875 4845 1885
rect 4805 1855 4815 1875
rect 4835 1855 4845 1875
rect 4805 1845 4845 1855
rect 4925 1875 4965 1885
rect 4925 1855 4935 1875
rect 4955 1855 4965 1875
rect 4925 1845 4965 1855
rect 5045 1880 5085 1885
rect 5045 1850 5050 1880
rect 5080 1850 5085 1880
rect 5045 1845 5085 1850
rect 5135 1875 5175 1885
rect 5135 1855 5145 1875
rect 5165 1855 5175 1875
rect 5135 1845 5175 1855
rect 4125 1825 4145 1845
rect 4215 1825 4235 1845
rect 4455 1825 4475 1845
rect 4575 1825 4595 1845
rect 4115 1820 4155 1825
rect 4115 1790 4120 1820
rect 4150 1790 4155 1820
rect 4115 1785 4155 1790
rect 4205 1820 4245 1825
rect 4205 1790 4210 1820
rect 4240 1790 4245 1820
rect 4205 1785 4245 1790
rect 4445 1820 4485 1825
rect 4445 1790 4450 1820
rect 4480 1790 4485 1820
rect 4445 1785 4485 1790
rect 4565 1820 4605 1825
rect 4565 1790 4570 1820
rect 4600 1790 4605 1820
rect 4565 1785 4605 1790
rect 4205 1760 4245 1765
rect 4205 1730 4210 1760
rect 4240 1730 4245 1760
rect 4205 1725 4245 1730
rect 4445 1760 4485 1765
rect 4445 1730 4450 1760
rect 4480 1730 4485 1760
rect 4445 1725 4485 1730
rect 4575 1720 4595 1785
rect 4695 1765 4715 1845
rect 4815 1825 4835 1845
rect 4935 1825 4955 1845
rect 5145 1825 5165 1845
rect 4805 1820 4845 1825
rect 4805 1790 4810 1820
rect 4840 1790 4845 1820
rect 4805 1785 4845 1790
rect 4925 1820 4965 1825
rect 4925 1790 4930 1820
rect 4960 1790 4965 1820
rect 4925 1785 4965 1790
rect 5135 1820 5175 1825
rect 5135 1790 5140 1820
rect 5170 1790 5175 1820
rect 5135 1785 5175 1790
rect 5280 1765 5300 2255
rect 5325 2150 5345 3105
rect 5315 2145 5355 2150
rect 5315 2115 5320 2145
rect 5350 2115 5355 2145
rect 5315 2110 5355 2115
rect 5370 1825 5390 3300
rect 5410 3285 5450 3290
rect 5410 3255 5415 3285
rect 5445 3255 5450 3285
rect 5410 3250 5450 3255
rect 5360 1820 5400 1825
rect 5360 1790 5365 1820
rect 5395 1790 5400 1820
rect 5360 1785 5400 1790
rect 4685 1760 4725 1765
rect 4685 1730 4690 1760
rect 4720 1730 4725 1760
rect 4685 1725 4725 1730
rect 4745 1760 4785 1765
rect 4745 1730 4750 1760
rect 4780 1730 4785 1760
rect 4745 1725 4785 1730
rect 5270 1760 5310 1765
rect 5270 1730 5275 1760
rect 5305 1730 5310 1760
rect 5270 1725 5310 1730
rect 4325 1715 4365 1720
rect 4325 1685 4330 1715
rect 4360 1685 4365 1715
rect 4325 1680 4365 1685
rect 4565 1715 4605 1720
rect 4565 1685 4570 1715
rect 4600 1685 4605 1715
rect 4565 1680 4605 1685
rect 4805 1715 4845 1720
rect 4805 1685 4810 1715
rect 4840 1685 4845 1715
rect 4805 1680 4845 1685
rect 5420 1600 5440 3250
rect 16060 3160 16080 4280
rect 16340 4265 16360 4285
rect 16750 4280 16790 4285
rect 17140 4315 17180 4320
rect 17140 4285 17145 4315
rect 17175 4285 17180 4315
rect 17140 4280 17180 4285
rect 17203 4310 17237 4320
rect 17203 4290 17211 4310
rect 17229 4290 17237 4310
rect 17203 4280 17237 4290
rect 17260 4315 17300 4320
rect 17260 4285 17265 4315
rect 17295 4285 17300 4315
rect 17260 4280 17300 4285
rect 17380 4315 17420 4320
rect 17380 4285 17385 4315
rect 17415 4285 17420 4315
rect 17380 4280 17420 4285
rect 17500 4315 17540 4320
rect 17500 4285 17505 4315
rect 17535 4285 17540 4315
rect 17500 4280 17540 4285
rect 17210 4265 17230 4280
rect 16105 4260 16145 4265
rect 16105 4230 16110 4260
rect 16140 4230 16145 4260
rect 16105 4225 16145 4230
rect 16330 4260 16370 4265
rect 16330 4230 16335 4260
rect 16365 4230 16370 4260
rect 16330 4225 16370 4230
rect 17200 4260 17240 4265
rect 17200 4230 17205 4260
rect 17235 4230 17240 4260
rect 17200 4225 17240 4230
rect 16050 3155 16090 3160
rect 16050 3125 16055 3155
rect 16085 3125 16090 3155
rect 16050 3120 16090 3125
rect 15265 2965 15305 2970
rect 14904 2935 15045 2940
rect 14904 2905 14910 2935
rect 14940 2905 14960 2935
rect 14990 2905 15010 2935
rect 15040 2905 15045 2935
rect 15265 2935 15270 2965
rect 15300 2935 15305 2965
rect 15265 2930 15305 2935
rect 15375 2965 15415 2970
rect 15375 2935 15380 2965
rect 15410 2935 15415 2965
rect 15375 2930 15415 2935
rect 15485 2965 15525 2970
rect 15485 2935 15490 2965
rect 15520 2935 15525 2965
rect 15485 2930 15525 2935
rect 15595 2965 15635 2970
rect 15595 2935 15600 2965
rect 15630 2935 15635 2965
rect 15595 2930 15635 2935
rect 15653 2960 15687 2970
rect 15653 2940 15661 2960
rect 15679 2940 15687 2960
rect 15653 2930 15687 2940
rect 15705 2965 15745 2970
rect 15705 2935 15710 2965
rect 15740 2935 15745 2965
rect 15705 2930 15745 2935
rect 14904 2900 15045 2905
rect 14965 2885 14985 2900
rect 14955 2880 14995 2885
rect 14955 2850 14960 2880
rect 14990 2850 14995 2880
rect 14955 2845 14995 2850
rect 15385 2830 15405 2930
rect 15660 2885 15680 2930
rect 15650 2880 15690 2885
rect 15650 2850 15655 2880
rect 15685 2850 15690 2880
rect 15650 2845 15690 2850
rect 16000 2880 16040 2885
rect 16000 2850 16005 2880
rect 16035 2850 16040 2880
rect 16000 2845 16040 2850
rect 14515 2825 14555 2830
rect 14515 2795 14520 2825
rect 14550 2795 14555 2825
rect 14515 2790 14555 2795
rect 15375 2825 15415 2830
rect 15375 2795 15380 2825
rect 15410 2795 15415 2825
rect 15375 2790 15415 2795
rect 14525 2120 14545 2790
rect 15210 2705 15250 2710
rect 15210 2675 15215 2705
rect 15245 2675 15250 2705
rect 15210 2670 15250 2675
rect 15320 2705 15360 2710
rect 15320 2675 15325 2705
rect 15355 2675 15360 2705
rect 15320 2670 15360 2675
rect 15430 2705 15470 2710
rect 15430 2675 15435 2705
rect 15465 2675 15470 2705
rect 15430 2670 15470 2675
rect 15540 2705 15580 2710
rect 15540 2675 15545 2705
rect 15575 2675 15580 2705
rect 15540 2670 15580 2675
rect 15650 2705 15690 2710
rect 15650 2675 15655 2705
rect 15685 2675 15690 2705
rect 15650 2670 15690 2675
rect 15760 2705 15800 2710
rect 15760 2675 15765 2705
rect 15795 2675 15800 2705
rect 15760 2670 15800 2675
rect 15020 2435 15060 2440
rect 15020 2405 15025 2435
rect 15055 2405 15060 2435
rect 15020 2400 15060 2405
rect 15265 2435 15305 2440
rect 15265 2405 15270 2435
rect 15300 2405 15305 2435
rect 15265 2400 15305 2405
rect 15375 2435 15415 2440
rect 15375 2405 15380 2435
rect 15410 2405 15415 2435
rect 15375 2400 15415 2405
rect 15485 2435 15525 2440
rect 15485 2405 15490 2435
rect 15520 2405 15525 2435
rect 15485 2400 15525 2405
rect 15595 2435 15635 2440
rect 15595 2405 15600 2435
rect 15630 2405 15635 2435
rect 15595 2400 15635 2405
rect 15705 2435 15745 2440
rect 15705 2405 15710 2435
rect 15740 2405 15745 2435
rect 16010 2425 16030 2845
rect 16115 2480 16135 4225
rect 16360 4205 16400 4210
rect 16360 4175 16365 4205
rect 16395 4175 16400 4205
rect 16360 4170 16400 4175
rect 16470 4205 16510 4210
rect 16470 4175 16475 4205
rect 16505 4175 16510 4205
rect 16470 4170 16510 4175
rect 16580 4205 16620 4210
rect 16580 4175 16585 4205
rect 16615 4175 16620 4205
rect 16580 4170 16620 4175
rect 16690 4205 16730 4210
rect 16690 4175 16695 4205
rect 16725 4175 16730 4205
rect 16690 4170 16730 4175
rect 16800 4205 16840 4210
rect 16800 4175 16805 4205
rect 16835 4175 16840 4205
rect 16800 4170 16840 4175
rect 16910 4205 16950 4210
rect 16910 4175 16915 4205
rect 16945 4175 16950 4205
rect 16910 4170 16950 4175
rect 17020 4205 17060 4210
rect 17020 4175 17025 4205
rect 17055 4175 17060 4205
rect 17020 4170 17060 4175
rect 17130 4205 17170 4210
rect 17130 4175 17135 4205
rect 17165 4175 17170 4205
rect 17130 4170 17170 4175
rect 17240 4205 17280 4210
rect 17240 4175 17245 4205
rect 17275 4175 17280 4205
rect 17240 4170 17280 4175
rect 17350 4205 17390 4210
rect 17350 4175 17355 4205
rect 17385 4175 17390 4205
rect 17350 4170 17390 4175
rect 16305 4085 16345 4090
rect 16305 4055 16310 4085
rect 16340 4055 16345 4085
rect 16305 4050 16345 4055
rect 16362 4080 16398 4090
rect 16362 4060 16370 4080
rect 16390 4060 16398 4080
rect 16362 4050 16398 4060
rect 16415 4080 16455 4090
rect 16415 4060 16425 4080
rect 16445 4060 16455 4080
rect 16415 4050 16455 4060
rect 16525 4085 16565 4090
rect 16525 4055 16530 4085
rect 16560 4055 16565 4085
rect 16525 4050 16565 4055
rect 16635 4080 16675 4090
rect 16635 4060 16645 4080
rect 16665 4060 16675 4080
rect 16635 4050 16675 4060
rect 16745 4085 16785 4090
rect 16745 4055 16750 4085
rect 16780 4055 16785 4085
rect 16745 4050 16785 4055
rect 16855 4080 16895 4090
rect 16855 4060 16865 4080
rect 16885 4060 16895 4080
rect 16855 4050 16895 4060
rect 16965 4085 17005 4090
rect 16965 4055 16970 4085
rect 17000 4055 17005 4085
rect 16965 4050 17005 4055
rect 17075 4080 17115 4090
rect 17075 4060 17085 4080
rect 17105 4060 17115 4080
rect 17075 4050 17115 4060
rect 17185 4085 17225 4090
rect 17185 4055 17190 4085
rect 17220 4055 17225 4085
rect 17185 4050 17225 4055
rect 17295 4080 17335 4090
rect 17295 4060 17305 4080
rect 17325 4060 17335 4080
rect 17295 4050 17335 4060
rect 17405 4085 17445 4090
rect 17405 4055 17410 4085
rect 17440 4055 17445 4085
rect 17405 4050 17445 4055
rect 16310 3960 16350 3965
rect 16310 3930 16315 3960
rect 16345 3930 16350 3960
rect 16310 3925 16350 3930
rect 16370 3905 16390 4050
rect 16425 4030 16445 4050
rect 16645 4030 16665 4050
rect 16865 4030 16885 4050
rect 17085 4030 17105 4050
rect 17305 4030 17325 4050
rect 16415 4025 16455 4030
rect 16415 3995 16420 4025
rect 16450 3995 16455 4025
rect 16415 3990 16455 3995
rect 16635 4025 16675 4030
rect 16635 3995 16640 4025
rect 16670 3995 16675 4025
rect 16635 3990 16675 3995
rect 16855 4025 16895 4030
rect 16855 3995 16860 4025
rect 16890 3995 16895 4025
rect 16855 3990 16895 3995
rect 17075 4025 17115 4030
rect 17075 3995 17080 4025
rect 17110 3995 17115 4025
rect 17075 3990 17115 3995
rect 17295 4025 17335 4030
rect 17295 3995 17300 4025
rect 17330 3995 17335 4025
rect 17295 3990 17335 3995
rect 16425 3965 16445 3990
rect 17415 3965 17435 4050
rect 16415 3960 16455 3965
rect 16415 3930 16420 3960
rect 16450 3930 16455 3960
rect 16415 3925 16455 3930
rect 16525 3960 16565 3965
rect 16525 3930 16530 3960
rect 16560 3930 16565 3960
rect 16525 3925 16565 3930
rect 16635 3960 16675 3965
rect 16635 3930 16640 3960
rect 16670 3930 16675 3960
rect 16635 3925 16675 3930
rect 16745 3960 16785 3965
rect 16745 3930 16750 3960
rect 16780 3930 16785 3960
rect 16745 3925 16785 3930
rect 17050 3960 17090 3965
rect 17050 3930 17055 3960
rect 17085 3930 17090 3960
rect 17050 3925 17090 3930
rect 17155 3960 17195 3965
rect 17155 3930 17160 3960
rect 17190 3930 17195 3960
rect 17155 3925 17195 3930
rect 17265 3960 17305 3965
rect 17265 3930 17270 3960
rect 17300 3930 17305 3960
rect 17265 3925 17305 3930
rect 17375 3960 17435 3965
rect 17375 3930 17380 3960
rect 17410 3930 17435 3960
rect 17375 3925 17435 3930
rect 17485 3960 17525 3965
rect 17485 3930 17490 3960
rect 17520 3930 17525 3960
rect 17485 3925 17525 3930
rect 16271 3900 16303 3905
rect 16271 3870 16274 3900
rect 16300 3870 16303 3900
rect 16271 3865 16303 3870
rect 16360 3895 16400 3905
rect 16360 3875 16370 3895
rect 16390 3875 16400 3895
rect 16360 3865 16400 3875
rect 16470 3900 16510 3905
rect 16470 3870 16475 3900
rect 16505 3870 16510 3900
rect 16470 3865 16510 3870
rect 16690 3900 16730 3905
rect 16690 3870 16695 3900
rect 16725 3870 16730 3900
rect 16690 3865 16730 3870
rect 16800 3895 16840 3905
rect 16800 3875 16810 3895
rect 16830 3875 16840 3895
rect 16800 3865 16840 3875
rect 17011 3900 17043 3905
rect 17011 3870 17014 3900
rect 17040 3870 17043 3900
rect 17011 3865 17043 3870
rect 17210 3900 17250 3905
rect 17210 3870 17215 3900
rect 17245 3870 17250 3900
rect 17210 3865 17250 3870
rect 17430 3900 17470 3905
rect 17430 3870 17435 3900
rect 17465 3870 17470 3900
rect 17430 3865 17470 3870
rect 17760 3900 17800 3905
rect 17760 3870 17765 3900
rect 17795 3870 17800 3900
rect 17760 3865 17800 3870
rect 16402 3780 16434 3785
rect 16402 3750 16405 3780
rect 16431 3750 16434 3780
rect 16402 3745 16434 3750
rect 16622 3780 16654 3785
rect 16622 3750 16625 3780
rect 16651 3750 16654 3780
rect 16622 3745 16654 3750
rect 16766 3780 16798 3785
rect 16766 3750 16769 3780
rect 16795 3750 16798 3780
rect 16766 3745 16798 3750
rect 17142 3780 17174 3785
rect 17142 3750 17145 3780
rect 17171 3750 17174 3780
rect 17142 3745 17174 3750
rect 17362 3780 17394 3785
rect 17362 3750 17365 3780
rect 17391 3750 17394 3780
rect 17362 3745 17394 3750
rect 17506 3780 17538 3785
rect 17506 3750 17509 3780
rect 17535 3750 17538 3780
rect 17506 3745 17538 3750
rect 16990 3730 17030 3735
rect 16250 3720 16290 3725
rect 16250 3690 16255 3720
rect 16285 3690 16290 3720
rect 16250 3685 16290 3690
rect 16355 3720 16395 3725
rect 16355 3690 16360 3720
rect 16390 3690 16395 3720
rect 16355 3685 16395 3690
rect 16470 3720 16510 3725
rect 16470 3690 16475 3720
rect 16505 3690 16510 3720
rect 16470 3685 16510 3690
rect 16575 3720 16615 3725
rect 16575 3690 16580 3720
rect 16610 3690 16615 3720
rect 16575 3685 16615 3690
rect 16690 3720 16730 3725
rect 16690 3690 16695 3720
rect 16725 3690 16730 3720
rect 16690 3685 16730 3690
rect 16805 3720 16845 3725
rect 16805 3690 16810 3720
rect 16840 3690 16845 3720
rect 16990 3700 16995 3730
rect 17025 3700 17030 3730
rect 16990 3695 17030 3700
rect 17210 3730 17250 3735
rect 17210 3700 17215 3730
rect 17245 3700 17250 3730
rect 17210 3695 17250 3700
rect 17430 3730 17470 3735
rect 17430 3700 17435 3730
rect 17465 3700 17470 3730
rect 17430 3695 17470 3700
rect 16805 3685 16845 3690
rect 17095 3685 17135 3690
rect 17095 3655 17100 3685
rect 17130 3655 17135 3685
rect 17095 3650 17135 3655
rect 17315 3685 17355 3690
rect 17315 3655 17320 3685
rect 17350 3655 17355 3685
rect 17315 3650 17355 3655
rect 17545 3685 17585 3690
rect 17545 3655 17550 3685
rect 17580 3655 17585 3685
rect 17545 3650 17585 3655
rect 16340 3625 16380 3630
rect 16340 3595 16345 3625
rect 16375 3595 16380 3625
rect 16340 3590 16380 3595
rect 16460 3625 16500 3630
rect 16460 3595 16465 3625
rect 16495 3595 16500 3625
rect 16460 3590 16500 3595
rect 16580 3625 16620 3630
rect 16580 3595 16585 3625
rect 16615 3595 16620 3625
rect 16580 3590 16620 3595
rect 16700 3625 16740 3630
rect 16700 3595 16705 3625
rect 16735 3595 16740 3625
rect 16700 3590 16740 3595
rect 16820 3625 16860 3630
rect 16820 3595 16825 3625
rect 16855 3595 16860 3625
rect 16820 3590 16860 3595
rect 16940 3625 16980 3630
rect 16940 3595 16945 3625
rect 16975 3595 16980 3625
rect 16940 3590 16980 3595
rect 17060 3625 17100 3630
rect 17060 3595 17065 3625
rect 17095 3595 17100 3625
rect 17060 3590 17100 3595
rect 17180 3625 17220 3630
rect 17180 3595 17185 3625
rect 17215 3595 17220 3625
rect 17180 3590 17220 3595
rect 17300 3625 17340 3630
rect 17300 3595 17305 3625
rect 17335 3595 17340 3625
rect 17300 3590 17340 3595
rect 17420 3625 17460 3630
rect 17420 3595 17425 3625
rect 17455 3595 17460 3625
rect 17420 3590 17460 3595
rect 16280 3150 16320 3160
rect 16280 3130 16290 3150
rect 16310 3130 16320 3150
rect 16280 3120 16320 3130
rect 16400 3150 16440 3160
rect 16400 3130 16410 3150
rect 16430 3130 16440 3150
rect 16400 3120 16440 3130
rect 16520 3150 16560 3160
rect 16520 3130 16530 3150
rect 16550 3130 16560 3150
rect 16520 3120 16560 3130
rect 16640 3150 16680 3160
rect 16640 3130 16650 3150
rect 16670 3130 16680 3150
rect 16640 3120 16680 3130
rect 16760 3150 16800 3160
rect 16760 3130 16770 3150
rect 16790 3130 16800 3150
rect 16760 3120 16800 3130
rect 16823 3155 16857 3160
rect 16823 3125 16826 3155
rect 16854 3125 16857 3155
rect 16823 3120 16857 3125
rect 16880 3150 16920 3160
rect 16880 3130 16890 3150
rect 16910 3130 16920 3150
rect 16880 3120 16920 3130
rect 17000 3150 17040 3160
rect 17000 3130 17010 3150
rect 17030 3130 17040 3150
rect 17000 3120 17040 3130
rect 17120 3150 17160 3160
rect 17120 3130 17130 3150
rect 17150 3130 17160 3150
rect 17120 3120 17160 3130
rect 17240 3150 17280 3160
rect 17240 3130 17250 3150
rect 17270 3130 17280 3150
rect 17240 3120 17280 3130
rect 17360 3150 17400 3160
rect 17360 3130 17370 3150
rect 17390 3130 17400 3150
rect 17360 3120 17400 3130
rect 17480 3150 17520 3160
rect 17480 3130 17490 3150
rect 17510 3130 17520 3150
rect 17480 3120 17520 3130
rect 16290 3105 16310 3120
rect 16280 3100 16320 3105
rect 16280 3070 16285 3100
rect 16315 3070 16320 3100
rect 16280 3065 16320 3070
rect 16410 3060 16430 3120
rect 16530 3105 16550 3120
rect 16520 3100 16560 3105
rect 16520 3070 16525 3100
rect 16555 3070 16560 3100
rect 16520 3065 16560 3070
rect 16650 3060 16670 3120
rect 16770 3105 16790 3120
rect 16760 3100 16800 3105
rect 16760 3070 16765 3100
rect 16795 3070 16800 3100
rect 16760 3065 16800 3070
rect 16890 3060 16910 3120
rect 17010 3105 17030 3120
rect 17000 3100 17040 3105
rect 17000 3070 17005 3100
rect 17035 3070 17040 3100
rect 17000 3065 17040 3070
rect 17130 3060 17150 3120
rect 17250 3105 17270 3120
rect 17240 3100 17280 3105
rect 17240 3070 17245 3100
rect 17275 3070 17280 3100
rect 17240 3065 17280 3070
rect 17370 3060 17390 3120
rect 17490 3105 17510 3120
rect 17480 3100 17520 3105
rect 17480 3070 17485 3100
rect 17515 3070 17520 3100
rect 17480 3065 17520 3070
rect 16400 3055 16440 3060
rect 16400 3025 16405 3055
rect 16435 3025 16440 3055
rect 16400 3020 16440 3025
rect 16640 3055 16680 3060
rect 16640 3025 16645 3055
rect 16675 3025 16680 3055
rect 16640 3020 16680 3025
rect 16880 3055 16920 3060
rect 16880 3025 16885 3055
rect 16915 3025 16920 3055
rect 16880 3020 16920 3025
rect 17120 3055 17160 3060
rect 17120 3025 17125 3055
rect 17155 3025 17160 3055
rect 17120 3020 17160 3025
rect 17360 3055 17400 3060
rect 17360 3025 17365 3055
rect 17395 3025 17400 3055
rect 17360 3020 17400 3025
rect 16410 3005 16430 3020
rect 16340 3000 16380 3005
rect 16340 2970 16345 3000
rect 16375 2970 16380 3000
rect 16340 2965 16380 2970
rect 16400 3000 16440 3005
rect 16400 2970 16405 3000
rect 16435 2970 16440 3000
rect 16400 2965 16440 2970
rect 16580 3000 16620 3005
rect 16580 2970 16585 3000
rect 16615 2970 16620 3000
rect 16580 2965 16620 2970
rect 16820 3000 16860 3005
rect 16820 2970 16825 3000
rect 16855 2970 16860 3000
rect 16820 2965 16860 2970
rect 17060 3000 17100 3005
rect 17060 2970 17065 3000
rect 17095 2970 17100 3000
rect 17060 2965 17100 2970
rect 17300 3000 17340 3005
rect 17300 2970 17305 3000
rect 17335 2970 17340 3000
rect 17300 2965 17340 2970
rect 16350 2950 16370 2965
rect 16590 2950 16610 2965
rect 16830 2950 16850 2965
rect 17070 2950 17090 2965
rect 17310 2950 17330 2965
rect 17490 2950 17510 3065
rect 16340 2940 16380 2950
rect 16340 2920 16350 2940
rect 16370 2920 16380 2940
rect 16340 2910 16380 2920
rect 16460 2945 16500 2950
rect 16460 2915 16465 2945
rect 16495 2915 16500 2945
rect 16460 2910 16500 2915
rect 16580 2940 16620 2950
rect 16580 2920 16590 2940
rect 16610 2920 16620 2940
rect 16580 2910 16620 2920
rect 16700 2945 16740 2950
rect 16700 2915 16705 2945
rect 16735 2915 16740 2945
rect 16700 2910 16740 2915
rect 16820 2940 16860 2950
rect 16820 2920 16830 2940
rect 16850 2920 16860 2940
rect 16820 2910 16860 2920
rect 16940 2945 16980 2950
rect 16940 2915 16945 2945
rect 16975 2915 16980 2945
rect 16940 2910 16980 2915
rect 17060 2940 17100 2950
rect 17060 2920 17070 2940
rect 17090 2920 17100 2940
rect 17060 2910 17100 2920
rect 17180 2945 17220 2950
rect 17180 2915 17185 2945
rect 17215 2915 17220 2945
rect 17180 2910 17220 2915
rect 17300 2940 17340 2950
rect 17300 2920 17310 2940
rect 17330 2920 17340 2940
rect 17300 2910 17340 2920
rect 17420 2945 17460 2950
rect 17420 2915 17425 2945
rect 17455 2915 17460 2945
rect 17420 2910 17460 2915
rect 17480 2945 17520 2950
rect 17480 2915 17485 2945
rect 17515 2915 17520 2945
rect 17480 2910 17520 2915
rect 17690 2880 17730 2885
rect 17690 2850 17695 2880
rect 17725 2850 17730 2880
rect 17690 2845 17730 2850
rect 16105 2475 16145 2480
rect 16105 2445 16110 2475
rect 16140 2445 16145 2475
rect 16105 2440 16145 2445
rect 16280 2470 16320 2480
rect 16280 2450 16290 2470
rect 16310 2450 16320 2470
rect 16280 2440 16320 2450
rect 16400 2470 16440 2480
rect 16400 2450 16410 2470
rect 16430 2450 16440 2470
rect 16400 2440 16440 2450
rect 16520 2470 16560 2480
rect 16520 2450 16530 2470
rect 16550 2450 16560 2470
rect 16520 2440 16560 2450
rect 16640 2470 16680 2480
rect 16640 2450 16650 2470
rect 16670 2450 16680 2470
rect 16640 2440 16680 2450
rect 16760 2470 16800 2480
rect 16760 2450 16770 2470
rect 16790 2450 16800 2470
rect 16760 2440 16800 2450
rect 16823 2475 16857 2480
rect 16823 2445 16826 2475
rect 16854 2445 16857 2475
rect 16823 2440 16857 2445
rect 16880 2470 16920 2480
rect 16880 2450 16890 2470
rect 16910 2450 16920 2470
rect 16880 2440 16920 2450
rect 17000 2470 17040 2480
rect 17000 2450 17010 2470
rect 17030 2450 17040 2470
rect 17000 2440 17040 2450
rect 17120 2470 17160 2480
rect 17120 2450 17130 2470
rect 17150 2450 17160 2470
rect 17120 2440 17160 2450
rect 17240 2470 17280 2480
rect 17240 2450 17250 2470
rect 17270 2450 17280 2470
rect 17240 2440 17280 2450
rect 17360 2470 17400 2480
rect 17360 2450 17370 2470
rect 17390 2450 17400 2470
rect 17360 2440 17400 2450
rect 17480 2470 17520 2480
rect 17480 2450 17490 2470
rect 17510 2450 17520 2470
rect 17480 2440 17520 2450
rect 16290 2425 16310 2440
rect 15705 2400 15745 2405
rect 16000 2420 16040 2425
rect 14510 2110 14560 2120
rect 14510 2080 14520 2110
rect 14550 2080 14560 2110
rect 14510 2070 14560 2080
rect 14525 1710 14545 2070
rect 14790 2005 14825 2011
rect 14790 1965 14825 1970
rect 14850 2005 14885 2010
rect 14850 1965 14885 1970
rect 14910 2005 14945 2011
rect 14910 1965 14945 1970
rect 14970 2005 15005 2010
rect 15030 2005 15050 2400
rect 15765 2390 15805 2395
rect 15765 2360 15770 2390
rect 15800 2360 15805 2390
rect 16000 2390 16005 2420
rect 16035 2390 16040 2420
rect 16000 2385 16040 2390
rect 16280 2420 16320 2425
rect 16280 2390 16285 2420
rect 16315 2390 16320 2420
rect 16280 2385 16320 2390
rect 16410 2380 16430 2440
rect 16530 2425 16550 2440
rect 16520 2420 16560 2425
rect 16520 2390 16525 2420
rect 16555 2390 16560 2420
rect 16520 2385 16560 2390
rect 16650 2380 16670 2440
rect 16770 2425 16790 2440
rect 16760 2420 16800 2425
rect 16760 2390 16765 2420
rect 16795 2390 16800 2420
rect 16760 2385 16800 2390
rect 15765 2355 15805 2360
rect 16400 2375 16440 2380
rect 16400 2345 16405 2375
rect 16435 2345 16440 2375
rect 16400 2340 16440 2345
rect 16640 2375 16680 2380
rect 16640 2345 16645 2375
rect 16675 2345 16680 2375
rect 16640 2340 16680 2345
rect 16000 2325 16040 2330
rect 15065 2315 15105 2320
rect 15065 2285 15070 2315
rect 15100 2285 15105 2315
rect 15065 2280 15105 2285
rect 15265 2315 15305 2320
rect 15265 2285 15270 2315
rect 15300 2285 15305 2315
rect 15265 2280 15305 2285
rect 15375 2315 15415 2320
rect 15375 2285 15380 2315
rect 15410 2285 15415 2315
rect 15375 2280 15415 2285
rect 15485 2315 15525 2320
rect 15485 2285 15490 2315
rect 15520 2285 15525 2315
rect 15485 2280 15525 2285
rect 15595 2315 15635 2320
rect 15595 2285 15600 2315
rect 15630 2285 15635 2315
rect 15595 2280 15635 2285
rect 15705 2315 15745 2320
rect 15705 2285 15710 2315
rect 15740 2285 15745 2315
rect 16000 2295 16005 2325
rect 16035 2295 16040 2325
rect 16000 2290 16040 2295
rect 15705 2280 15745 2285
rect 14970 1965 15005 1970
rect 15020 2000 15060 2005
rect 15020 1970 15025 2000
rect 15055 1970 15060 2000
rect 15020 1965 15060 1970
rect 14800 1900 14820 1965
rect 14920 1950 14940 1965
rect 15075 1950 15095 2280
rect 15950 2180 15990 2185
rect 15950 2150 15955 2180
rect 15985 2150 15990 2180
rect 15950 2145 15990 2150
rect 14910 1945 14950 1950
rect 14910 1915 14915 1945
rect 14945 1915 14950 1945
rect 14910 1910 14950 1915
rect 15065 1945 15105 1950
rect 15065 1915 15070 1945
rect 15100 1915 15105 1945
rect 15065 1910 15105 1915
rect 15210 1945 15250 1950
rect 15210 1915 15215 1945
rect 15245 1915 15250 1945
rect 15210 1910 15250 1915
rect 15320 1945 15360 1950
rect 15320 1915 15325 1945
rect 15355 1915 15360 1945
rect 15320 1910 15360 1915
rect 15430 1945 15470 1950
rect 15430 1915 15435 1945
rect 15465 1915 15470 1945
rect 15430 1910 15470 1915
rect 15540 1945 15580 1950
rect 15540 1915 15545 1945
rect 15575 1915 15580 1945
rect 15540 1910 15580 1915
rect 15650 1945 15690 1950
rect 15650 1915 15655 1945
rect 15685 1915 15690 1945
rect 15650 1910 15690 1915
rect 15760 1945 15800 1950
rect 15760 1915 15765 1945
rect 15795 1915 15800 1945
rect 15760 1910 15800 1915
rect 14790 1895 14830 1900
rect 14790 1865 14795 1895
rect 14825 1865 14830 1895
rect 14790 1860 14830 1865
rect 14965 1760 15005 1765
rect 14965 1730 14970 1760
rect 15000 1730 15005 1760
rect 14965 1725 15005 1730
rect 15555 1760 15595 1765
rect 15555 1730 15560 1760
rect 15590 1730 15595 1760
rect 15555 1725 15595 1730
rect 15835 1760 15875 1765
rect 15835 1730 15840 1760
rect 15870 1730 15875 1760
rect 15835 1725 15875 1730
rect 14515 1705 14555 1710
rect 14515 1675 14520 1705
rect 14550 1675 14555 1705
rect 14515 1670 14555 1675
rect 14975 1650 14995 1725
rect 15565 1710 15585 1725
rect 15030 1705 15070 1710
rect 15030 1675 15035 1705
rect 15065 1675 15070 1705
rect 15030 1670 15070 1675
rect 15255 1705 15295 1710
rect 15255 1675 15260 1705
rect 15290 1675 15295 1705
rect 15255 1670 15295 1675
rect 15455 1705 15495 1710
rect 15455 1675 15460 1705
rect 15490 1675 15495 1705
rect 15455 1670 15495 1675
rect 15558 1700 15592 1710
rect 15558 1680 15566 1700
rect 15584 1680 15592 1700
rect 15558 1670 15592 1680
rect 15655 1705 15695 1710
rect 15655 1675 15660 1705
rect 15690 1675 15695 1705
rect 15655 1670 15695 1675
rect 15040 1650 15060 1670
rect 14970 1645 15005 1650
rect 14970 1605 15005 1610
rect 15030 1645 15065 1650
rect 15030 1605 15065 1610
rect 4805 1595 4845 1600
rect 4805 1565 4810 1595
rect 4840 1565 4845 1595
rect 4805 1560 4845 1565
rect 5410 1595 5450 1600
rect 5410 1565 5415 1595
rect 5445 1565 5450 1595
rect 5410 1560 5450 1565
rect 4265 1545 4305 1550
rect 4265 1515 4270 1545
rect 4300 1515 4305 1545
rect 4265 1510 4305 1515
rect 4385 1545 4425 1550
rect 4385 1515 4390 1545
rect 4420 1515 4425 1545
rect 4385 1510 4425 1515
rect 4505 1545 4545 1550
rect 4505 1515 4510 1545
rect 4540 1515 4545 1545
rect 4505 1510 4545 1515
rect 4625 1545 4665 1550
rect 4625 1515 4630 1545
rect 4660 1515 4665 1545
rect 4625 1510 4665 1515
rect 4745 1545 4785 1550
rect 4745 1515 4750 1545
rect 4780 1515 4785 1545
rect 4745 1510 4785 1515
rect 5135 1545 5175 1550
rect 5135 1515 5140 1545
rect 5170 1515 5175 1545
rect 5135 1510 5175 1515
rect 4205 1500 4245 1505
rect 4055 1480 4095 1490
rect 4055 1460 4065 1480
rect 4085 1460 4095 1480
rect 4205 1470 4210 1500
rect 4240 1470 4245 1500
rect 4205 1465 4245 1470
rect 4325 1500 4365 1505
rect 4325 1470 4330 1500
rect 4360 1470 4365 1500
rect 4325 1465 4365 1470
rect 4445 1500 4485 1505
rect 4445 1470 4450 1500
rect 4480 1470 4485 1500
rect 4445 1465 4485 1470
rect 4685 1500 4725 1505
rect 4685 1470 4690 1500
rect 4720 1470 4725 1500
rect 4685 1465 4725 1470
rect 4805 1500 4845 1505
rect 4805 1470 4810 1500
rect 4840 1470 4845 1500
rect 4805 1465 4845 1470
rect 4925 1500 4965 1505
rect 4925 1470 4930 1500
rect 4960 1470 4965 1500
rect 4925 1465 4965 1470
rect 5045 1500 5085 1505
rect 5045 1470 5050 1500
rect 5080 1470 5085 1500
rect 5145 1490 5165 1510
rect 5045 1465 5085 1470
rect 5135 1480 5175 1490
rect 4055 1450 4095 1460
rect 5135 1460 5145 1480
rect 5165 1460 5175 1480
rect 5135 1450 5175 1460
rect 15845 1395 15865 1725
rect 15835 1390 15875 1395
rect 15835 1360 15840 1390
rect 15870 1360 15875 1390
rect 15835 1355 15875 1360
rect 3375 1185 3415 1190
rect 3375 1155 3380 1185
rect 3410 1155 3415 1185
rect 3375 1150 3415 1155
rect 3985 1185 4025 1190
rect 3985 1155 3990 1185
rect 4020 1155 4025 1185
rect 3985 1150 4025 1155
rect 4595 1185 4635 1190
rect 4595 1155 4600 1185
rect 4630 1155 4635 1185
rect 4595 1150 4635 1155
rect 2945 1125 2985 1130
rect 2945 1095 2950 1125
rect 2980 1095 2985 1125
rect 2945 1090 2985 1095
rect 3025 1125 3065 1130
rect 3025 1095 3030 1125
rect 3060 1095 3065 1125
rect 3025 1090 3065 1095
rect 3105 1125 3145 1130
rect 3105 1095 3110 1125
rect 3140 1095 3145 1125
rect 3105 1090 3145 1095
rect 3185 1125 3225 1130
rect 3185 1095 3190 1125
rect 3220 1095 3225 1125
rect 3185 1090 3225 1095
rect 3265 1125 3305 1130
rect 3265 1095 3270 1125
rect 3300 1095 3305 1125
rect 3265 1090 3305 1095
rect 3345 1125 3385 1130
rect 3345 1095 3350 1125
rect 3380 1095 3385 1125
rect 3345 1090 3385 1095
rect 3425 1125 3465 1130
rect 3425 1095 3430 1125
rect 3460 1095 3465 1125
rect 3425 1090 3465 1095
rect 3505 1125 3545 1130
rect 3505 1095 3510 1125
rect 3540 1095 3545 1125
rect 3505 1090 3545 1095
rect 3585 1125 3625 1130
rect 3585 1095 3590 1125
rect 3620 1095 3625 1125
rect 3585 1090 3625 1095
rect 3665 1125 3705 1130
rect 3665 1095 3670 1125
rect 3700 1095 3705 1125
rect 3665 1090 3705 1095
rect 3745 1125 3785 1130
rect 3745 1095 3750 1125
rect 3780 1095 3785 1125
rect 3745 1090 3785 1095
rect 3825 1125 3865 1130
rect 3825 1095 3830 1125
rect 3860 1095 3865 1125
rect 3825 1090 3865 1095
rect 3905 1125 3945 1130
rect 3905 1095 3910 1125
rect 3940 1095 3945 1125
rect 3905 1090 3945 1095
rect 3985 1125 4025 1130
rect 3985 1095 3990 1125
rect 4020 1095 4025 1125
rect 3985 1090 4025 1095
rect 4065 1125 4105 1130
rect 4065 1095 4070 1125
rect 4100 1095 4105 1125
rect 4065 1090 4105 1095
rect 4145 1125 4185 1130
rect 4145 1095 4150 1125
rect 4180 1095 4185 1125
rect 4145 1090 4185 1095
rect 4225 1125 4265 1130
rect 4225 1095 4230 1125
rect 4260 1095 4265 1125
rect 4225 1090 4265 1095
rect 4305 1125 4345 1130
rect 4305 1095 4310 1125
rect 4340 1095 4345 1125
rect 4305 1090 4345 1095
rect 4385 1125 4425 1130
rect 4385 1095 4390 1125
rect 4420 1095 4425 1125
rect 4385 1090 4425 1095
rect 4465 1125 4505 1130
rect 4465 1095 4470 1125
rect 4500 1095 4505 1125
rect 4465 1090 4505 1095
rect 4545 1125 4585 1130
rect 4545 1095 4550 1125
rect 4580 1095 4585 1125
rect 4545 1090 4585 1095
rect 4625 1125 4665 1130
rect 4625 1095 4630 1125
rect 4660 1095 4665 1125
rect 4625 1090 4665 1095
rect 4705 1125 4745 1130
rect 4705 1095 4710 1125
rect 4740 1095 4745 1125
rect 4705 1090 4745 1095
rect 4785 1125 4825 1130
rect 4785 1095 4790 1125
rect 4820 1095 4825 1125
rect 4785 1090 4825 1095
rect 4865 1125 4905 1130
rect 4865 1095 4870 1125
rect 4900 1095 4905 1125
rect 4865 1090 4905 1095
rect 4945 1125 4985 1130
rect 4945 1095 4950 1125
rect 4980 1095 4985 1125
rect 4945 1090 4985 1095
rect 2620 1040 2660 1045
rect 2620 1010 2625 1040
rect 2655 1010 2660 1040
rect 2620 1005 2660 1010
rect 2905 1040 2945 1045
rect 2905 1010 2910 1040
rect 2940 1010 2945 1040
rect 2905 1005 2945 1010
rect 5110 1040 5150 1045
rect 5110 1010 5115 1040
rect 5145 1010 5150 1040
rect 5110 1005 5150 1010
rect 15355 935 15395 940
rect 2995 930 3035 935
rect 2995 900 3000 930
rect 3030 900 3035 930
rect 2995 895 3035 900
rect 3175 930 3215 935
rect 3175 900 3180 930
rect 3210 900 3215 930
rect 3175 895 3215 900
rect 3355 930 3395 935
rect 3355 900 3360 930
rect 3390 900 3395 930
rect 3355 895 3395 900
rect 3535 930 3575 935
rect 3535 900 3540 930
rect 3570 900 3575 930
rect 3535 895 3575 900
rect 3715 930 3755 935
rect 3715 900 3720 930
rect 3750 900 3755 930
rect 3715 895 3755 900
rect 3895 930 3935 935
rect 3895 900 3900 930
rect 3930 900 3935 930
rect 3895 895 3935 900
rect 4075 930 4115 935
rect 4075 900 4080 930
rect 4110 900 4115 930
rect 4075 895 4115 900
rect 4255 930 4295 935
rect 4255 900 4260 930
rect 4290 900 4295 930
rect 4255 895 4295 900
rect 4435 930 4475 935
rect 4435 900 4440 930
rect 4470 900 4475 930
rect 4435 895 4475 900
rect 4615 930 4655 935
rect 4615 900 4620 930
rect 4650 900 4655 930
rect 4615 895 4655 900
rect 4795 930 4835 935
rect 4795 900 4800 930
rect 4830 900 4835 930
rect 4795 895 4835 900
rect 4975 930 5015 935
rect 4975 900 4980 930
rect 5010 900 5015 930
rect 15355 905 15360 935
rect 15390 905 15395 935
rect 15355 900 15395 905
rect 15555 935 15595 940
rect 15555 905 15560 935
rect 15590 905 15595 935
rect 15555 900 15595 905
rect 4975 895 5015 900
rect 15960 800 15980 2145
rect 16010 1900 16030 2290
rect 16440 2280 16480 2285
rect 16440 2250 16445 2280
rect 16475 2250 16480 2280
rect 16440 2245 16480 2250
rect 16660 2280 16700 2285
rect 16660 2250 16665 2280
rect 16695 2250 16700 2280
rect 16660 2245 16700 2250
rect 16330 2235 16370 2240
rect 16330 2205 16335 2235
rect 16365 2205 16370 2235
rect 16330 2200 16370 2205
rect 16340 2185 16360 2200
rect 16450 2185 16470 2245
rect 16550 2235 16590 2240
rect 16550 2205 16555 2235
rect 16585 2205 16590 2235
rect 16550 2200 16590 2205
rect 16560 2185 16580 2200
rect 16670 2185 16690 2245
rect 16770 2240 16790 2385
rect 16890 2380 16910 2440
rect 17010 2425 17030 2440
rect 17000 2420 17040 2425
rect 17000 2390 17005 2420
rect 17035 2390 17040 2420
rect 17000 2385 17040 2390
rect 17130 2380 17150 2440
rect 17250 2425 17270 2440
rect 17240 2420 17280 2425
rect 17240 2390 17245 2420
rect 17275 2390 17280 2420
rect 17240 2385 17280 2390
rect 17370 2380 17390 2440
rect 17490 2425 17510 2440
rect 17480 2420 17520 2425
rect 17480 2390 17485 2420
rect 17515 2390 17520 2420
rect 17480 2385 17520 2390
rect 17700 2380 17720 2845
rect 16880 2375 16920 2380
rect 16880 2345 16885 2375
rect 16915 2345 16920 2375
rect 16880 2340 16920 2345
rect 17120 2375 17160 2380
rect 17120 2345 17125 2375
rect 17155 2345 17160 2375
rect 17120 2340 17160 2345
rect 17360 2375 17400 2380
rect 17360 2345 17365 2375
rect 17395 2345 17400 2375
rect 17360 2340 17400 2345
rect 17690 2375 17730 2380
rect 17690 2345 17695 2375
rect 17725 2345 17730 2375
rect 17690 2340 17730 2345
rect 17120 2285 17140 2340
rect 17770 2330 17790 3865
rect 17860 3730 17900 3735
rect 17860 3700 17865 3730
rect 17895 3700 17900 3730
rect 17860 3695 17900 3700
rect 17805 3685 17845 3690
rect 17805 3655 17810 3685
rect 17840 3655 17845 3685
rect 17805 3650 17845 3655
rect 17760 2325 17800 2330
rect 17760 2295 17765 2325
rect 17795 2295 17800 2325
rect 17760 2290 17800 2295
rect 16880 2280 16920 2285
rect 16880 2250 16885 2280
rect 16915 2250 16920 2280
rect 16880 2245 16920 2250
rect 17100 2280 17140 2285
rect 17100 2250 17105 2280
rect 17135 2250 17140 2280
rect 17100 2245 17140 2250
rect 17320 2280 17360 2285
rect 17320 2250 17325 2280
rect 17355 2250 17360 2280
rect 17320 2245 17360 2250
rect 16770 2235 16810 2240
rect 16770 2205 16775 2235
rect 16805 2205 16810 2235
rect 16770 2200 16810 2205
rect 16780 2185 16800 2200
rect 16890 2185 16910 2245
rect 16990 2235 17030 2240
rect 16990 2205 16995 2235
rect 17025 2205 17030 2235
rect 16990 2200 17030 2205
rect 17000 2185 17020 2200
rect 17110 2185 17130 2245
rect 17210 2235 17250 2240
rect 17210 2205 17215 2235
rect 17245 2205 17250 2235
rect 17210 2200 17250 2205
rect 17220 2185 17240 2200
rect 17330 2185 17350 2245
rect 17430 2235 17470 2240
rect 17430 2205 17435 2235
rect 17465 2205 17470 2235
rect 17430 2200 17470 2205
rect 17440 2185 17460 2200
rect 16330 2175 16370 2185
rect 16330 2155 16340 2175
rect 16360 2155 16370 2175
rect 16330 2145 16370 2155
rect 16440 2175 16480 2185
rect 16440 2155 16450 2175
rect 16470 2155 16480 2175
rect 16440 2145 16480 2155
rect 16550 2175 16590 2185
rect 16550 2155 16560 2175
rect 16580 2155 16590 2175
rect 16550 2145 16590 2155
rect 16660 2175 16700 2185
rect 16660 2155 16670 2175
rect 16690 2155 16700 2175
rect 16660 2145 16700 2155
rect 16770 2175 16810 2185
rect 16770 2155 16780 2175
rect 16800 2155 16810 2175
rect 16770 2145 16810 2155
rect 16828 2180 16862 2185
rect 16828 2150 16831 2180
rect 16859 2150 16862 2180
rect 16828 2145 16862 2150
rect 16880 2175 16920 2185
rect 16880 2155 16890 2175
rect 16910 2155 16920 2175
rect 16880 2145 16920 2155
rect 16990 2175 17030 2185
rect 16990 2155 17000 2175
rect 17020 2155 17030 2175
rect 16990 2145 17030 2155
rect 17100 2175 17140 2185
rect 17100 2155 17110 2175
rect 17130 2155 17140 2175
rect 17100 2145 17140 2155
rect 17210 2175 17250 2185
rect 17210 2155 17220 2175
rect 17240 2155 17250 2175
rect 17210 2145 17250 2155
rect 17320 2175 17360 2185
rect 17320 2155 17330 2175
rect 17350 2155 17360 2175
rect 17320 2145 17360 2155
rect 17430 2175 17470 2185
rect 17430 2155 17440 2175
rect 17460 2155 17470 2175
rect 17430 2145 17470 2155
rect 16385 1960 16425 1965
rect 16385 1930 16390 1960
rect 16420 1930 16425 1960
rect 16385 1925 16425 1930
rect 16495 1955 16535 1965
rect 16495 1935 16505 1955
rect 16525 1935 16535 1955
rect 16495 1925 16535 1935
rect 16605 1960 16645 1965
rect 16605 1930 16610 1960
rect 16640 1930 16645 1960
rect 16605 1925 16645 1930
rect 16715 1955 16755 1965
rect 16715 1935 16725 1955
rect 16745 1935 16755 1955
rect 16715 1925 16755 1935
rect 16825 1960 16865 1965
rect 16825 1930 16830 1960
rect 16860 1930 16865 1960
rect 16825 1925 16865 1930
rect 16935 1955 16975 1965
rect 16935 1935 16945 1955
rect 16965 1935 16975 1955
rect 16935 1925 16975 1935
rect 17045 1960 17085 1965
rect 17045 1930 17050 1960
rect 17080 1930 17085 1960
rect 17045 1925 17085 1930
rect 17155 1955 17195 1965
rect 17155 1935 17165 1955
rect 17185 1935 17195 1955
rect 17155 1925 17195 1935
rect 17245 1960 17305 1965
rect 17245 1930 17270 1960
rect 17300 1930 17305 1960
rect 17245 1925 17305 1930
rect 17375 1955 17415 1965
rect 17375 1935 17385 1955
rect 17405 1935 17415 1955
rect 17375 1925 17415 1935
rect 16505 1910 16525 1925
rect 16725 1910 16745 1925
rect 16945 1910 16965 1925
rect 17165 1910 17185 1925
rect 16495 1905 16555 1910
rect 16000 1895 16040 1900
rect 16000 1865 16005 1895
rect 16035 1865 16040 1895
rect 16495 1875 16500 1905
rect 16530 1875 16555 1905
rect 16495 1870 16555 1875
rect 16715 1905 16755 1910
rect 16715 1875 16720 1905
rect 16750 1875 16755 1905
rect 16715 1870 16755 1875
rect 16935 1905 16975 1910
rect 16935 1875 16940 1905
rect 16970 1875 16975 1905
rect 16935 1870 16975 1875
rect 17155 1905 17195 1910
rect 17155 1875 17160 1905
rect 17190 1875 17195 1905
rect 17155 1870 17195 1875
rect 16000 1860 16040 1865
rect 16190 1850 16230 1855
rect 16190 1820 16195 1850
rect 16225 1820 16230 1850
rect 16190 1815 16230 1820
rect 16410 1850 16450 1855
rect 16410 1820 16415 1850
rect 16445 1820 16450 1850
rect 16410 1815 16450 1820
rect 16200 1780 16220 1815
rect 16420 1780 16440 1815
rect 16190 1770 16230 1780
rect 16085 1760 16125 1765
rect 16085 1730 16090 1760
rect 16120 1730 16125 1760
rect 16190 1750 16200 1770
rect 16220 1750 16230 1770
rect 16410 1770 16450 1780
rect 16190 1740 16230 1750
rect 16305 1760 16345 1765
rect 16085 1725 16125 1730
rect 16305 1730 16310 1760
rect 16340 1730 16345 1760
rect 16410 1750 16420 1770
rect 16440 1750 16450 1770
rect 16535 1765 16555 1870
rect 17245 1855 17265 1925
rect 17385 1910 17405 1925
rect 17375 1905 17415 1910
rect 17375 1875 17380 1905
rect 17410 1875 17415 1905
rect 17770 1900 17790 2290
rect 17375 1870 17415 1875
rect 17760 1895 17800 1900
rect 17760 1865 17765 1895
rect 17795 1865 17800 1895
rect 17760 1860 17800 1865
rect 16640 1850 16680 1855
rect 16640 1820 16645 1850
rect 16675 1820 16680 1850
rect 16640 1815 16680 1820
rect 17230 1850 17270 1855
rect 17230 1820 17235 1850
rect 17265 1820 17270 1850
rect 17230 1815 17270 1820
rect 17450 1850 17490 1855
rect 17450 1820 17455 1850
rect 17485 1820 17490 1850
rect 17450 1815 17490 1820
rect 17680 1850 17720 1855
rect 17680 1820 17685 1850
rect 17715 1820 17720 1850
rect 17680 1815 17720 1820
rect 16650 1780 16670 1815
rect 16820 1805 16860 1810
rect 16640 1770 16680 1780
rect 16820 1775 16825 1805
rect 16855 1775 16860 1805
rect 16820 1770 16860 1775
rect 16940 1805 16980 1810
rect 16940 1775 16945 1805
rect 16975 1775 16980 1805
rect 17240 1780 17260 1815
rect 17460 1780 17480 1815
rect 17690 1780 17710 1815
rect 16940 1770 16980 1775
rect 17230 1770 17270 1780
rect 16410 1740 16450 1750
rect 16525 1760 16565 1765
rect 16305 1725 16345 1730
rect 16525 1730 16530 1760
rect 16560 1730 16565 1760
rect 16640 1750 16650 1770
rect 16670 1750 16680 1770
rect 16640 1740 16680 1750
rect 16525 1725 16565 1730
rect 16830 1720 16850 1770
rect 16950 1720 16970 1770
rect 17125 1760 17165 1765
rect 17125 1730 17130 1760
rect 17160 1730 17165 1760
rect 17230 1750 17240 1770
rect 17260 1750 17270 1770
rect 17450 1770 17490 1780
rect 17230 1740 17270 1750
rect 17345 1760 17385 1765
rect 17125 1725 17165 1730
rect 17345 1730 17350 1760
rect 17380 1730 17385 1760
rect 17450 1750 17460 1770
rect 17480 1750 17490 1770
rect 17680 1770 17720 1780
rect 17450 1740 17490 1750
rect 17565 1760 17605 1765
rect 17345 1725 17385 1730
rect 17565 1730 17570 1760
rect 17600 1730 17605 1760
rect 17680 1750 17690 1770
rect 17710 1750 17720 1770
rect 17680 1740 17720 1750
rect 17565 1725 17605 1730
rect 16237 1715 16269 1720
rect 16237 1685 16240 1715
rect 16266 1685 16269 1715
rect 16237 1680 16269 1685
rect 16457 1715 16489 1720
rect 16457 1685 16460 1715
rect 16486 1685 16489 1715
rect 16457 1680 16489 1685
rect 16601 1715 16633 1720
rect 16601 1685 16604 1715
rect 16630 1685 16633 1715
rect 16601 1680 16633 1685
rect 16820 1710 16850 1720
rect 16820 1690 16825 1710
rect 16845 1690 16850 1710
rect 16820 1680 16850 1690
rect 16867 1715 16899 1720
rect 16867 1685 16870 1715
rect 16896 1685 16899 1715
rect 16867 1680 16899 1685
rect 16950 1710 16980 1720
rect 16950 1690 16955 1710
rect 16975 1690 16980 1710
rect 16950 1680 16980 1690
rect 17277 1715 17309 1720
rect 17277 1685 17280 1715
rect 17306 1685 17309 1715
rect 17277 1680 17309 1685
rect 17497 1715 17529 1720
rect 17497 1685 17500 1715
rect 17526 1685 17529 1715
rect 17497 1680 17529 1685
rect 17641 1715 17673 1720
rect 17641 1685 17644 1715
rect 17670 1685 17673 1715
rect 17641 1680 17673 1685
rect 16106 1495 16138 1500
rect 16106 1465 16109 1495
rect 16135 1465 16138 1495
rect 16106 1460 16138 1465
rect 16305 1495 16345 1500
rect 16305 1465 16310 1495
rect 16340 1465 16345 1495
rect 16305 1460 16345 1465
rect 16525 1495 16565 1500
rect 16525 1465 16530 1495
rect 16560 1465 16565 1495
rect 16525 1460 16565 1465
rect 16825 1490 16855 1500
rect 16825 1470 16830 1490
rect 16850 1470 16855 1490
rect 16825 1460 16855 1470
rect 16875 1490 16905 1500
rect 16875 1470 16880 1490
rect 16900 1470 16905 1490
rect 16875 1460 16905 1470
rect 16922 1495 16954 1500
rect 16922 1465 16925 1495
rect 16951 1465 16954 1495
rect 16922 1460 16954 1465
rect 17146 1495 17178 1500
rect 17146 1465 17149 1495
rect 17175 1465 17178 1495
rect 17146 1460 17178 1465
rect 17345 1495 17385 1500
rect 17345 1465 17350 1495
rect 17380 1465 17385 1495
rect 17345 1460 17385 1465
rect 17565 1495 17605 1500
rect 17565 1465 17570 1495
rect 17600 1465 17605 1495
rect 17565 1460 17605 1465
rect 16145 1435 16185 1440
rect 16145 1405 16150 1435
rect 16180 1405 16185 1435
rect 16145 1400 16185 1405
rect 16250 1435 16290 1440
rect 16250 1405 16255 1435
rect 16285 1405 16290 1435
rect 16250 1400 16290 1405
rect 16360 1435 16400 1440
rect 16360 1405 16365 1435
rect 16395 1405 16400 1435
rect 16360 1400 16400 1405
rect 16470 1435 16510 1440
rect 16470 1405 16475 1435
rect 16505 1405 16510 1435
rect 16470 1400 16510 1405
rect 16580 1435 16620 1440
rect 16580 1405 16585 1435
rect 16615 1405 16620 1435
rect 16580 1400 16620 1405
rect 16830 1350 16850 1460
rect 16005 1345 16045 1350
rect 16005 1315 16010 1345
rect 16040 1315 16045 1345
rect 16005 1310 16045 1315
rect 16810 1345 16850 1350
rect 16810 1315 16815 1345
rect 16845 1315 16850 1345
rect 16810 1310 16850 1315
rect 16015 860 16035 1310
rect 16315 1295 16355 1300
rect 16315 1265 16320 1295
rect 16350 1265 16355 1295
rect 16315 1260 16355 1265
rect 16325 1240 16345 1260
rect 16820 1240 16840 1310
rect 16880 1300 16900 1460
rect 17185 1435 17225 1440
rect 17185 1405 17190 1435
rect 17220 1405 17225 1435
rect 17185 1400 17225 1405
rect 17290 1435 17330 1440
rect 17290 1405 17295 1435
rect 17325 1405 17330 1435
rect 17290 1400 17330 1405
rect 17400 1435 17440 1440
rect 17400 1405 17405 1435
rect 17435 1405 17440 1435
rect 17400 1400 17440 1405
rect 17510 1435 17550 1440
rect 17510 1405 17515 1435
rect 17545 1405 17550 1435
rect 17510 1400 17550 1405
rect 17620 1435 17660 1440
rect 17620 1405 17625 1435
rect 17655 1405 17660 1435
rect 17620 1400 17660 1405
rect 16880 1295 16920 1300
rect 16880 1265 16885 1295
rect 16915 1265 16920 1295
rect 16880 1260 16920 1265
rect 17815 1255 17835 3650
rect 17595 1250 17635 1255
rect 16315 1230 16355 1240
rect 16315 1210 16325 1230
rect 16345 1210 16355 1230
rect 16315 1200 16355 1210
rect 16425 1235 16465 1240
rect 16425 1205 16430 1235
rect 16460 1205 16465 1235
rect 16425 1200 16465 1205
rect 16535 1235 16575 1240
rect 16535 1205 16540 1235
rect 16570 1205 16575 1235
rect 16535 1200 16575 1205
rect 16645 1235 16685 1240
rect 16645 1205 16650 1235
rect 16680 1205 16685 1235
rect 16645 1200 16685 1205
rect 16755 1235 16795 1240
rect 16755 1205 16760 1235
rect 16790 1205 16795 1235
rect 16755 1200 16795 1205
rect 16815 1230 16845 1240
rect 16815 1210 16820 1230
rect 16840 1210 16845 1230
rect 16815 1200 16845 1210
rect 16865 1235 16905 1240
rect 16865 1205 16870 1235
rect 16900 1205 16905 1235
rect 16865 1200 16905 1205
rect 16975 1235 17015 1240
rect 16975 1205 16980 1235
rect 17010 1205 17015 1235
rect 16975 1200 17015 1205
rect 17085 1235 17125 1240
rect 17085 1205 17090 1235
rect 17120 1205 17125 1235
rect 17085 1200 17125 1205
rect 17195 1235 17235 1240
rect 17195 1205 17200 1235
rect 17230 1205 17235 1235
rect 17195 1200 17235 1205
rect 17305 1235 17345 1240
rect 17305 1205 17310 1235
rect 17340 1205 17345 1235
rect 17305 1200 17345 1205
rect 17415 1235 17455 1240
rect 17415 1205 17420 1235
rect 17450 1205 17455 1235
rect 17415 1200 17455 1205
rect 17525 1235 17565 1240
rect 17525 1205 17530 1235
rect 17560 1205 17565 1235
rect 17595 1220 17600 1250
rect 17630 1220 17635 1250
rect 17595 1215 17635 1220
rect 17805 1250 17845 1255
rect 17805 1220 17810 1250
rect 17840 1220 17845 1250
rect 17805 1215 17845 1220
rect 17525 1200 17565 1205
rect 16165 915 16205 920
rect 16165 885 16170 915
rect 16200 885 16205 915
rect 16165 880 16205 885
rect 16260 915 16300 920
rect 16260 885 16265 915
rect 16295 885 16300 915
rect 16260 880 16300 885
rect 16370 915 16410 920
rect 16370 885 16375 915
rect 16405 885 16410 915
rect 16370 880 16410 885
rect 16480 915 16520 920
rect 16480 885 16485 915
rect 16515 885 16520 915
rect 16480 880 16520 885
rect 16590 915 16630 920
rect 16590 885 16595 915
rect 16625 885 16630 915
rect 16590 880 16630 885
rect 16700 915 16740 920
rect 16700 885 16705 915
rect 16735 885 16740 915
rect 16700 880 16740 885
rect 16810 915 16850 920
rect 16810 885 16815 915
rect 16845 885 16850 915
rect 16810 880 16850 885
rect 16920 915 16960 920
rect 16920 885 16925 915
rect 16955 885 16960 915
rect 16920 880 16960 885
rect 17030 915 17070 920
rect 17030 885 17035 915
rect 17065 885 17070 915
rect 17030 880 17070 885
rect 17140 915 17180 920
rect 17140 885 17145 915
rect 17175 885 17180 915
rect 17140 880 17180 885
rect 17250 915 17290 920
rect 17250 885 17255 915
rect 17285 885 17290 915
rect 17250 880 17290 885
rect 17360 915 17400 920
rect 17360 885 17365 915
rect 17395 885 17400 915
rect 17360 880 17400 885
rect 17470 915 17510 920
rect 17470 885 17475 915
rect 17505 885 17510 915
rect 17470 880 17510 885
rect 17620 915 17660 920
rect 17620 885 17625 915
rect 17655 885 17660 915
rect 17620 880 17660 885
rect 16935 860 16975 865
rect 16005 855 16045 860
rect 16005 825 16010 855
rect 16040 825 16045 855
rect 16005 820 16045 825
rect 16495 855 16535 860
rect 16495 825 16500 855
rect 16530 825 16535 855
rect 16935 830 16940 860
rect 16970 830 16975 860
rect 16935 825 16975 830
rect 17155 860 17195 865
rect 17155 830 17160 860
rect 17190 830 17195 860
rect 17155 825 17195 830
rect 17375 860 17415 865
rect 17375 830 17380 860
rect 17410 830 17415 860
rect 17375 825 17415 830
rect 16495 820 16535 825
rect 16945 805 16965 825
rect 17165 805 17185 825
rect 17385 805 17405 825
rect 17815 805 17835 1215
rect 17870 865 17890 3695
rect 18000 3635 18040 3640
rect 18000 3605 18005 3635
rect 18035 3605 18040 3635
rect 18000 3600 18040 3605
rect 18110 3635 18150 3640
rect 18110 3605 18115 3635
rect 18145 3605 18150 3635
rect 18110 3600 18150 3605
rect 18220 3635 18260 3640
rect 18220 3605 18225 3635
rect 18255 3605 18260 3635
rect 18220 3600 18260 3605
rect 18330 3635 18370 3640
rect 18330 3605 18335 3635
rect 18365 3605 18370 3635
rect 18330 3600 18370 3605
rect 18440 3635 18480 3640
rect 18440 3605 18445 3635
rect 18475 3605 18480 3635
rect 18440 3600 18480 3605
rect 18550 3635 18590 3640
rect 18550 3605 18555 3635
rect 18585 3605 18590 3635
rect 18550 3600 18590 3605
rect 18805 3635 18845 3640
rect 18805 3605 18810 3635
rect 18840 3605 18845 3635
rect 18805 3600 18845 3605
rect 18815 3560 18835 3600
rect 18755 3555 18896 3560
rect 18755 3525 18760 3555
rect 18790 3525 18810 3555
rect 18840 3525 18860 3555
rect 18890 3525 18896 3555
rect 18755 3520 18896 3525
rect 18055 2965 18095 2970
rect 18055 2935 18060 2965
rect 18090 2935 18095 2965
rect 18055 2930 18095 2935
rect 18113 2960 18147 2970
rect 18113 2940 18121 2960
rect 18139 2940 18147 2960
rect 18113 2930 18147 2940
rect 18165 2965 18205 2970
rect 18165 2935 18170 2965
rect 18200 2935 18205 2965
rect 18165 2930 18205 2935
rect 18275 2965 18315 2970
rect 18275 2935 18280 2965
rect 18310 2935 18315 2965
rect 18275 2930 18315 2935
rect 18385 2965 18425 2970
rect 18385 2935 18390 2965
rect 18420 2935 18425 2965
rect 18385 2930 18425 2935
rect 18495 2965 18535 2970
rect 18495 2935 18500 2965
rect 18530 2935 18535 2965
rect 18495 2930 18535 2935
rect 18755 2935 18896 2940
rect 18120 2885 18140 2930
rect 18110 2880 18150 2885
rect 18110 2850 18115 2880
rect 18145 2850 18150 2880
rect 18110 2845 18150 2850
rect 18395 2830 18415 2930
rect 18755 2905 18760 2935
rect 18790 2905 18810 2935
rect 18840 2905 18860 2935
rect 18890 2905 18896 2935
rect 18755 2900 18896 2905
rect 18815 2885 18835 2900
rect 18805 2880 18845 2885
rect 18805 2850 18810 2880
rect 18840 2850 18845 2880
rect 18805 2845 18845 2850
rect 18385 2825 18425 2830
rect 18385 2795 18390 2825
rect 18420 2795 18425 2825
rect 18385 2790 18425 2795
rect 19245 2825 19285 2830
rect 19245 2795 19250 2825
rect 19280 2795 19285 2825
rect 19245 2790 19285 2795
rect 18000 2705 18040 2710
rect 18000 2675 18005 2705
rect 18035 2675 18040 2705
rect 18000 2670 18040 2675
rect 18110 2705 18150 2710
rect 18110 2675 18115 2705
rect 18145 2675 18150 2705
rect 18110 2670 18150 2675
rect 18220 2705 18260 2710
rect 18220 2675 18225 2705
rect 18255 2675 18260 2705
rect 18220 2670 18260 2675
rect 18330 2705 18370 2710
rect 18330 2675 18335 2705
rect 18365 2675 18370 2705
rect 18330 2670 18370 2675
rect 18440 2705 18480 2710
rect 18440 2675 18445 2705
rect 18475 2675 18480 2705
rect 18440 2670 18480 2675
rect 18550 2705 18590 2710
rect 18550 2675 18555 2705
rect 18585 2675 18590 2705
rect 18550 2670 18590 2675
rect 18055 2435 18095 2440
rect 18055 2405 18060 2435
rect 18090 2405 18095 2435
rect 18055 2400 18095 2405
rect 18165 2435 18205 2440
rect 18165 2405 18170 2435
rect 18200 2405 18205 2435
rect 18165 2400 18205 2405
rect 18275 2435 18315 2440
rect 18275 2405 18280 2435
rect 18310 2405 18315 2435
rect 18275 2400 18315 2405
rect 18385 2435 18425 2440
rect 18385 2405 18390 2435
rect 18420 2405 18425 2435
rect 18385 2400 18425 2405
rect 18495 2435 18535 2440
rect 18495 2405 18500 2435
rect 18530 2405 18535 2435
rect 18495 2400 18535 2405
rect 18740 2435 18780 2440
rect 18740 2405 18745 2435
rect 18775 2405 18780 2435
rect 18740 2400 18780 2405
rect 18025 2375 18065 2380
rect 18025 2345 18030 2375
rect 18060 2345 18065 2375
rect 18025 2340 18065 2345
rect 18055 2315 18095 2320
rect 18055 2285 18060 2315
rect 18090 2285 18095 2315
rect 18055 2280 18095 2285
rect 18165 2315 18205 2320
rect 18165 2285 18170 2315
rect 18200 2285 18205 2315
rect 18165 2280 18205 2285
rect 18275 2315 18315 2320
rect 18275 2285 18280 2315
rect 18310 2285 18315 2315
rect 18275 2280 18315 2285
rect 18385 2315 18425 2320
rect 18385 2285 18390 2315
rect 18420 2285 18425 2315
rect 18385 2280 18425 2285
rect 18495 2315 18535 2320
rect 18495 2285 18500 2315
rect 18530 2285 18535 2315
rect 18495 2280 18535 2285
rect 18695 2315 18735 2320
rect 18695 2285 18700 2315
rect 18730 2285 18735 2315
rect 18695 2280 18735 2285
rect 18705 1950 18725 2280
rect 18750 2005 18770 2400
rect 19255 2120 19275 2790
rect 19240 2110 19290 2120
rect 19240 2080 19250 2110
rect 19280 2080 19290 2110
rect 19240 2070 19290 2080
rect 18795 2005 18830 2010
rect 18740 2000 18780 2005
rect 18740 1970 18745 2000
rect 18775 1970 18780 2000
rect 18740 1965 18780 1970
rect 18795 1965 18830 1970
rect 18855 2005 18890 2011
rect 18855 1965 18890 1970
rect 18915 2005 18950 2010
rect 18915 1965 18950 1970
rect 18975 2005 19010 2011
rect 18975 1965 19010 1970
rect 18860 1950 18880 1965
rect 18000 1945 18040 1950
rect 18000 1915 18005 1945
rect 18035 1915 18040 1945
rect 18000 1910 18040 1915
rect 18110 1945 18150 1950
rect 18110 1915 18115 1945
rect 18145 1915 18150 1945
rect 18110 1910 18150 1915
rect 18220 1945 18260 1950
rect 18220 1915 18225 1945
rect 18255 1915 18260 1945
rect 18220 1910 18260 1915
rect 18330 1945 18370 1950
rect 18330 1915 18335 1945
rect 18365 1915 18370 1945
rect 18330 1910 18370 1915
rect 18440 1945 18480 1950
rect 18440 1915 18445 1945
rect 18475 1915 18480 1945
rect 18440 1910 18480 1915
rect 18550 1945 18590 1950
rect 18550 1915 18555 1945
rect 18585 1915 18590 1945
rect 18550 1910 18590 1915
rect 18695 1945 18735 1950
rect 18695 1915 18700 1945
rect 18730 1915 18735 1945
rect 18695 1910 18735 1915
rect 18850 1945 18890 1950
rect 18850 1915 18855 1945
rect 18885 1915 18890 1945
rect 18850 1910 18890 1915
rect 18980 1900 19000 1965
rect 18970 1895 19010 1900
rect 18970 1865 18975 1895
rect 19005 1865 19010 1895
rect 18970 1860 19010 1865
rect 17925 1760 17965 1765
rect 17925 1730 17930 1760
rect 17960 1730 17965 1760
rect 17925 1725 17965 1730
rect 18205 1760 18245 1765
rect 18205 1730 18210 1760
rect 18240 1730 18245 1760
rect 18205 1725 18245 1730
rect 18795 1760 18835 1765
rect 18795 1730 18800 1760
rect 18830 1730 18835 1760
rect 18795 1725 18835 1730
rect 17935 1395 17955 1725
rect 18215 1710 18235 1725
rect 18105 1705 18145 1710
rect 18105 1675 18110 1705
rect 18140 1675 18145 1705
rect 18105 1670 18145 1675
rect 18208 1700 18242 1710
rect 18208 1680 18216 1700
rect 18234 1680 18242 1700
rect 18208 1670 18242 1680
rect 18305 1705 18345 1710
rect 18305 1675 18310 1705
rect 18340 1675 18345 1705
rect 18305 1670 18345 1675
rect 18505 1705 18545 1710
rect 18505 1675 18510 1705
rect 18540 1675 18545 1705
rect 18505 1670 18545 1675
rect 18730 1705 18770 1710
rect 18730 1675 18735 1705
rect 18765 1675 18770 1705
rect 18730 1670 18770 1675
rect 18740 1650 18760 1670
rect 18805 1650 18825 1725
rect 19255 1710 19275 2070
rect 19245 1705 19285 1710
rect 19245 1675 19250 1705
rect 19280 1675 19285 1705
rect 19245 1670 19285 1675
rect 18735 1645 18770 1650
rect 18735 1605 18770 1610
rect 18795 1645 18830 1650
rect 18795 1605 18830 1610
rect 17925 1390 17965 1395
rect 17925 1360 17930 1390
rect 17960 1360 17965 1390
rect 17925 1355 17965 1360
rect 18205 935 18245 940
rect 18205 905 18210 935
rect 18240 905 18245 935
rect 18205 900 18245 905
rect 18405 935 18445 940
rect 18405 905 18410 935
rect 18440 905 18445 935
rect 18405 900 18445 905
rect 17860 860 17900 865
rect 17860 830 17865 860
rect 17895 830 17900 860
rect 17860 825 17900 830
rect 15950 795 15990 800
rect 15950 765 15955 795
rect 15985 765 15990 795
rect 2520 760 2560 765
rect 2520 730 2525 760
rect 2555 730 2560 760
rect 2520 725 2560 730
rect 3130 760 3170 765
rect 3130 730 3135 760
rect 3165 730 3170 760
rect 3130 725 3170 730
rect 3265 755 3305 765
rect 3265 735 3275 755
rect 3295 735 3305 755
rect 3265 725 3305 735
rect 3445 755 3485 765
rect 3445 735 3455 755
rect 3475 735 3485 755
rect 3445 725 3485 735
rect 3625 760 3665 765
rect 3625 730 3630 760
rect 3660 730 3665 760
rect 3625 725 3665 730
rect 3805 755 3845 765
rect 3805 735 3815 755
rect 3835 735 3845 755
rect 3805 725 3845 735
rect 3985 760 4025 765
rect 3985 730 3990 760
rect 4020 730 4025 760
rect 3985 725 4025 730
rect 4165 755 4205 765
rect 4165 735 4175 755
rect 4195 735 4205 755
rect 4165 725 4205 735
rect 4345 760 4385 765
rect 4345 730 4350 760
rect 4380 730 4385 760
rect 4345 725 4385 730
rect 4525 760 4565 765
rect 4525 730 4530 760
rect 4560 730 4565 760
rect 4525 725 4565 730
rect 4705 760 4745 765
rect 4705 730 4710 760
rect 4740 730 4745 760
rect 4705 725 4745 730
rect 4885 760 4925 765
rect 15950 760 15990 765
rect 16305 795 16345 800
rect 16305 765 16310 795
rect 16340 765 16345 795
rect 16305 760 16345 765
rect 16375 795 16415 800
rect 16375 765 16380 795
rect 16410 765 16415 795
rect 16375 760 16415 765
rect 16445 795 16485 800
rect 16445 765 16450 795
rect 16480 765 16485 795
rect 16935 795 16975 805
rect 16935 775 16945 795
rect 16965 775 16975 795
rect 16935 765 16975 775
rect 17045 800 17085 805
rect 17045 770 17050 800
rect 17080 770 17085 800
rect 17045 765 17085 770
rect 17155 795 17195 805
rect 17155 775 17165 795
rect 17185 775 17195 795
rect 17155 765 17195 775
rect 17265 800 17305 805
rect 17265 770 17270 800
rect 17300 770 17305 800
rect 17265 765 17305 770
rect 17375 795 17415 805
rect 17375 775 17385 795
rect 17405 775 17415 795
rect 17375 765 17415 775
rect 17485 800 17525 805
rect 17485 770 17490 800
rect 17520 770 17525 800
rect 17485 765 17525 770
rect 17805 800 17845 805
rect 17805 770 17810 800
rect 17840 770 17845 800
rect 17805 765 17845 770
rect 16445 760 16485 765
rect 4885 730 4890 760
rect 4920 730 4925 760
rect 4885 725 4925 730
rect 3275 295 3295 725
rect 3455 710 3475 725
rect 3815 710 3835 725
rect 3445 705 3485 710
rect 3445 675 3450 705
rect 3480 675 3485 705
rect 3445 670 3485 675
rect 3805 705 3845 710
rect 3805 675 3810 705
rect 3840 675 3845 705
rect 3805 670 3845 675
rect 3815 295 3835 670
rect 3995 295 4015 725
rect 4175 710 4195 725
rect 4165 705 4205 710
rect 4165 675 4170 705
rect 4200 675 4205 705
rect 4165 670 4205 675
rect 4715 295 4735 725
rect 16990 680 17030 685
rect 16990 650 16995 680
rect 17025 650 17030 680
rect 16990 645 17030 650
rect 17100 680 17140 685
rect 17100 650 17105 680
rect 17135 650 17140 680
rect 17100 645 17140 650
rect 17210 680 17250 685
rect 17210 650 17215 680
rect 17245 650 17250 680
rect 17210 645 17250 650
rect 17320 680 17360 685
rect 17320 650 17325 680
rect 17355 650 17360 680
rect 17320 645 17360 650
rect 17430 680 17470 685
rect 17430 650 17435 680
rect 17465 650 17470 680
rect 17430 645 17470 650
<< via1 >>
rect 16635 4510 16665 4515
rect 16635 4490 16640 4510
rect 16640 4490 16660 4510
rect 16660 4490 16665 4510
rect 16635 4485 16665 4490
rect 16755 4510 16785 4515
rect 16755 4490 16760 4510
rect 16760 4490 16780 4510
rect 16780 4490 16785 4510
rect 16755 4485 16785 4490
rect 16875 4510 16905 4515
rect 16875 4490 16880 4510
rect 16880 4490 16900 4510
rect 16900 4490 16905 4510
rect 16875 4485 16905 4490
rect 17085 4485 17115 4515
rect 16205 4450 16235 4455
rect 16205 4430 16210 4450
rect 16210 4430 16230 4450
rect 16230 4430 16235 4450
rect 16205 4425 16235 4430
rect 16465 4450 16495 4455
rect 16465 4430 16470 4450
rect 16470 4430 16490 4450
rect 16490 4430 16495 4450
rect 16465 4425 16495 4430
rect 16575 4465 16605 4470
rect 16575 4445 16580 4465
rect 16580 4445 16600 4465
rect 16600 4445 16605 4465
rect 16575 4440 16605 4445
rect 16695 4465 16725 4470
rect 16695 4445 16700 4465
rect 16700 4445 16720 4465
rect 16720 4445 16725 4465
rect 16695 4440 16725 4445
rect 16815 4465 16845 4470
rect 16815 4445 16820 4465
rect 16820 4445 16840 4465
rect 16840 4445 16845 4465
rect 16815 4440 16845 4445
rect 16935 4465 16965 4470
rect 16935 4445 16940 4465
rect 16940 4445 16960 4465
rect 16960 4445 16965 4465
rect 16935 4440 16965 4445
rect 17085 4440 17115 4445
rect 17085 4420 17090 4440
rect 17090 4420 17110 4440
rect 17110 4420 17115 4440
rect 17085 4415 17115 4420
rect 17205 4440 17235 4445
rect 17205 4420 17210 4440
rect 17210 4420 17230 4440
rect 17230 4420 17235 4440
rect 17205 4415 17235 4420
rect 17325 4440 17355 4445
rect 17325 4420 17330 4440
rect 17330 4420 17350 4440
rect 17350 4420 17355 4440
rect 17325 4415 17355 4420
rect 17445 4440 17475 4445
rect 17445 4420 17450 4440
rect 17450 4420 17470 4440
rect 17470 4420 17475 4440
rect 17445 4415 17475 4420
rect 17565 4440 17595 4445
rect 17565 4420 17570 4440
rect 17570 4420 17590 4440
rect 17590 4420 17595 4440
rect 17565 4415 17595 4420
rect 16055 4285 16085 4315
rect 16335 4295 16340 4320
rect 16340 4295 16360 4320
rect 16360 4295 16365 4320
rect 16335 4290 16365 4295
rect 16755 4310 16785 4315
rect 16755 4290 16760 4310
rect 16760 4290 16780 4310
rect 16780 4290 16785 4310
rect 16755 4285 16785 4290
rect 14960 3605 14990 3635
rect 15215 3630 15245 3635
rect 15215 3610 15220 3630
rect 15220 3610 15240 3630
rect 15240 3610 15245 3630
rect 15215 3605 15245 3610
rect 15325 3630 15355 3635
rect 15325 3610 15330 3630
rect 15330 3610 15350 3630
rect 15350 3610 15355 3630
rect 15325 3605 15355 3610
rect 15435 3630 15465 3635
rect 15435 3610 15440 3630
rect 15440 3610 15460 3630
rect 15460 3610 15465 3630
rect 15435 3605 15465 3610
rect 15545 3630 15575 3635
rect 15545 3610 15550 3630
rect 15550 3610 15570 3630
rect 15570 3610 15575 3630
rect 15545 3605 15575 3610
rect 15655 3630 15685 3635
rect 15655 3610 15660 3630
rect 15660 3610 15680 3630
rect 15680 3610 15685 3630
rect 15655 3605 15685 3610
rect 15765 3630 15795 3635
rect 15765 3610 15770 3630
rect 15770 3610 15790 3630
rect 15790 3610 15795 3630
rect 15765 3605 15795 3610
rect 1266 3495 1296 3525
rect 14910 3525 14940 3555
rect 14960 3525 14990 3555
rect 15010 3525 15040 3555
rect -10 3415 20 3445
rect 945 3415 975 3445
rect -55 3360 -25 3390
rect -55 2825 -25 2855
rect 1210 3310 1240 3340
rect 1165 3255 1195 3285
rect 51 3200 86 3205
rect 51 3175 56 3200
rect 56 3175 81 3200
rect 81 3175 86 3200
rect 51 3170 86 3175
rect 51 3140 86 3145
rect 51 3115 56 3140
rect 56 3115 81 3140
rect 81 3115 86 3140
rect 51 3110 86 3115
rect 1165 3070 1195 3100
rect 51 3060 86 3065
rect 51 3035 56 3060
rect 56 3035 81 3060
rect 81 3035 86 3060
rect 51 3030 86 3035
rect 51 3000 86 3005
rect 51 2975 56 3000
rect 56 2975 81 3000
rect 81 2975 86 3000
rect 51 2970 86 2975
rect 920 2880 950 2910
rect 1000 2880 1030 2910
rect 1080 2880 1110 2910
rect 4445 3465 4475 3495
rect 1645 3415 1675 3445
rect 2475 3420 2505 3450
rect 1266 3195 1301 3200
rect 1266 3170 1271 3195
rect 1271 3170 1296 3195
rect 1296 3170 1301 3195
rect 1266 3165 1301 3170
rect 1266 3135 1301 3140
rect 1266 3110 1271 3135
rect 1271 3110 1296 3135
rect 1296 3110 1301 3135
rect 1266 3105 1301 3110
rect 2335 2955 2370 2960
rect 2335 2930 2340 2955
rect 2340 2930 2365 2955
rect 2365 2930 2370 2955
rect 2335 2925 2370 2930
rect 2430 2925 2460 2955
rect 2335 2895 2370 2900
rect 2335 2870 2340 2895
rect 2340 2870 2365 2895
rect 2365 2870 2370 2895
rect 2335 2865 2370 2870
rect 56 2850 91 2855
rect 56 2825 61 2850
rect 61 2825 86 2850
rect 86 2825 91 2850
rect 56 2820 91 2825
rect 729 2850 764 2855
rect 729 2825 734 2850
rect 734 2825 759 2850
rect 759 2825 764 2850
rect 729 2820 764 2825
rect 1210 2820 1240 2850
rect 1266 2835 1301 2840
rect 1266 2810 1271 2835
rect 1271 2810 1296 2835
rect 1296 2810 1301 2835
rect 1266 2805 1301 2810
rect 1965 2835 2000 2840
rect 1965 2810 1970 2835
rect 1970 2810 1995 2835
rect 1995 2810 2000 2835
rect 1965 2805 2000 2810
rect 2335 2805 2365 2835
rect -10 2765 20 2795
rect 56 2790 91 2795
rect 56 2765 61 2790
rect 61 2765 86 2790
rect 86 2765 91 2790
rect 56 2760 91 2765
rect 729 2790 764 2795
rect 729 2765 734 2790
rect 734 2765 759 2790
rect 759 2765 764 2790
rect 729 2760 764 2765
rect 1266 2715 1296 2745
rect 2155 2715 2185 2745
rect -105 1690 -75 1720
rect -40 1715 -10 1720
rect -40 1695 -35 1715
rect -35 1695 -15 1715
rect -15 1695 -10 1715
rect -40 1690 -10 1695
rect 1270 1680 1297 1710
rect 2430 2215 2460 2245
rect 2335 2170 2365 2200
rect 2385 2120 2415 2150
rect 2695 3360 2725 3390
rect 3140 3310 3170 3340
rect 3395 3305 3425 3335
rect 2740 3210 2770 3240
rect 2625 3155 2655 3185
rect 2525 2950 2555 2980
rect 2475 1790 2505 1820
rect 2430 1730 2460 1760
rect 2385 1635 2415 1665
rect 2335 1565 2365 1595
rect 2625 2760 2655 2790
rect 2625 2315 2655 2345
rect 5145 3415 5175 3445
rect 5365 3305 5395 3335
rect 4890 3255 4920 3285
rect 4445 3155 4475 3185
rect 3140 3110 3170 3140
rect 4840 3110 4870 3140
rect 3990 3050 4020 3080
rect 3450 3005 3480 3035
rect 3810 3005 3840 3035
rect 4350 3005 4380 3035
rect 4710 3005 4740 3035
rect 5320 3110 5350 3140
rect 3085 2975 3115 2980
rect 3085 2955 3090 2975
rect 3090 2955 3110 2975
rect 3110 2955 3115 2975
rect 3085 2950 3115 2955
rect 3270 2975 3300 2980
rect 3270 2955 3275 2975
rect 3275 2955 3295 2975
rect 3295 2955 3300 2975
rect 3270 2950 3300 2955
rect 3630 2975 3660 2980
rect 3630 2955 3635 2975
rect 3635 2955 3655 2975
rect 3655 2955 3660 2975
rect 3630 2950 3660 2955
rect 4170 2975 4200 2980
rect 4170 2955 4175 2975
rect 4175 2955 4195 2975
rect 4195 2955 4200 2975
rect 4170 2950 4200 2955
rect 4530 2975 4560 2980
rect 4530 2955 4535 2975
rect 4535 2955 4555 2975
rect 4555 2955 4560 2975
rect 4530 2950 4560 2955
rect 3000 2805 3030 2810
rect 3000 2785 3005 2805
rect 3005 2785 3025 2805
rect 3025 2785 3030 2805
rect 3000 2780 3030 2785
rect 3180 2805 3210 2810
rect 3180 2785 3185 2805
rect 3185 2785 3205 2805
rect 3205 2785 3210 2805
rect 3180 2780 3210 2785
rect 3360 2805 3390 2810
rect 3360 2785 3365 2805
rect 3365 2785 3385 2805
rect 3385 2785 3390 2805
rect 3360 2780 3390 2785
rect 3540 2805 3570 2810
rect 3540 2785 3545 2805
rect 3545 2785 3565 2805
rect 3565 2785 3570 2805
rect 3540 2780 3570 2785
rect 3720 2805 3750 2810
rect 3720 2785 3725 2805
rect 3725 2785 3745 2805
rect 3745 2785 3750 2805
rect 3720 2780 3750 2785
rect 3900 2805 3930 2810
rect 3900 2785 3905 2805
rect 3905 2785 3925 2805
rect 3925 2785 3930 2805
rect 3900 2780 3930 2785
rect 4080 2805 4110 2810
rect 4080 2785 4085 2805
rect 4085 2785 4105 2805
rect 4105 2785 4110 2805
rect 4080 2780 4110 2785
rect 4260 2805 4290 2810
rect 4260 2785 4265 2805
rect 4265 2785 4285 2805
rect 4285 2785 4290 2805
rect 4260 2780 4290 2785
rect 4440 2805 4470 2810
rect 4440 2785 4445 2805
rect 4445 2785 4465 2805
rect 4465 2785 4470 2805
rect 4440 2780 4470 2785
rect 4620 2805 4650 2810
rect 4620 2785 4625 2805
rect 4625 2785 4645 2805
rect 4645 2785 4650 2805
rect 4620 2780 4650 2785
rect 4800 2805 4830 2810
rect 4800 2785 4805 2805
rect 4805 2785 4825 2805
rect 4825 2785 4830 2805
rect 4800 2780 4830 2785
rect 4980 2805 5010 2810
rect 4980 2785 4985 2805
rect 4985 2785 5005 2805
rect 5005 2785 5010 2805
rect 4980 2780 5010 2785
rect 3180 2745 3210 2750
rect 3180 2725 3185 2745
rect 3185 2725 3205 2745
rect 3205 2725 3210 2745
rect 3180 2720 3210 2725
rect 3360 2745 3390 2750
rect 3360 2725 3365 2745
rect 3365 2725 3385 2745
rect 3385 2725 3390 2745
rect 3360 2720 3390 2725
rect 3540 2745 3570 2750
rect 3540 2725 3545 2745
rect 3545 2725 3565 2745
rect 3565 2725 3570 2745
rect 3540 2720 3570 2725
rect 3720 2745 3750 2750
rect 3720 2725 3725 2745
rect 3725 2725 3745 2745
rect 3745 2725 3750 2745
rect 3720 2720 3750 2725
rect 3900 2745 3930 2750
rect 3900 2725 3905 2745
rect 3905 2725 3925 2745
rect 3925 2725 3930 2745
rect 3900 2720 3930 2725
rect 4080 2745 4110 2750
rect 4080 2725 4085 2745
rect 4085 2725 4105 2745
rect 4105 2725 4110 2745
rect 4080 2720 4110 2725
rect 4260 2745 4290 2750
rect 4260 2725 4265 2745
rect 4265 2725 4285 2745
rect 4285 2725 4290 2745
rect 4260 2720 4290 2725
rect 4440 2745 4470 2750
rect 4440 2725 4445 2745
rect 4445 2725 4465 2745
rect 4465 2725 4470 2745
rect 4440 2720 4470 2725
rect 4620 2745 4650 2750
rect 4620 2725 4625 2745
rect 4625 2725 4645 2745
rect 4645 2725 4650 2745
rect 4620 2720 4650 2725
rect 4800 2745 4830 2750
rect 4800 2725 4805 2745
rect 4805 2725 4825 2745
rect 4825 2725 4830 2745
rect 4800 2720 4830 2725
rect 3360 2370 3390 2375
rect 3360 2350 3365 2370
rect 3365 2350 3385 2370
rect 3385 2350 3390 2370
rect 3360 2345 3390 2350
rect 3810 2375 3840 2380
rect 3810 2355 3815 2375
rect 3815 2355 3835 2375
rect 3835 2355 3840 2375
rect 3810 2350 3840 2355
rect 4170 2375 4200 2380
rect 4170 2355 4175 2375
rect 4175 2355 4195 2375
rect 4195 2355 4200 2375
rect 4170 2350 4200 2355
rect 2740 2260 2770 2290
rect 3630 2330 3660 2335
rect 3630 2310 3635 2330
rect 3635 2310 3655 2330
rect 3655 2310 3660 2330
rect 3630 2305 3660 2310
rect 3450 2285 3480 2290
rect 3450 2265 3455 2285
rect 3455 2265 3475 2285
rect 3475 2265 3480 2285
rect 3450 2260 3480 2265
rect 3270 2170 3300 2200
rect 3810 2215 3840 2245
rect 3630 2120 3660 2150
rect 2750 2090 2780 2095
rect 2750 2070 2755 2090
rect 2755 2070 2775 2090
rect 2775 2070 2780 2090
rect 2750 2065 2780 2070
rect 2870 2090 2900 2095
rect 2870 2070 2875 2090
rect 2875 2070 2895 2090
rect 2895 2070 2900 2090
rect 2870 2065 2900 2070
rect 2990 2090 3020 2095
rect 2990 2070 2995 2090
rect 2995 2070 3015 2090
rect 3015 2070 3020 2090
rect 2990 2065 3020 2070
rect 3110 2090 3140 2095
rect 3110 2070 3115 2090
rect 3115 2070 3135 2090
rect 3135 2070 3140 2090
rect 3110 2065 3140 2070
rect 3230 2090 3260 2095
rect 3230 2070 3235 2090
rect 3235 2070 3255 2090
rect 3255 2070 3260 2090
rect 3230 2065 3260 2070
rect 3350 2090 3380 2095
rect 3350 2070 3355 2090
rect 3355 2070 3375 2090
rect 3375 2070 3380 2090
rect 3350 2065 3380 2070
rect 3470 2090 3500 2095
rect 3470 2070 3475 2090
rect 3475 2070 3495 2090
rect 3495 2070 3500 2090
rect 3470 2065 3500 2070
rect 3590 2090 3620 2095
rect 3590 2070 3595 2090
rect 3595 2070 3615 2090
rect 3615 2070 3620 2090
rect 3590 2065 3620 2070
rect 3710 2090 3740 2095
rect 3710 2070 3715 2090
rect 3715 2070 3735 2090
rect 3735 2070 3740 2090
rect 3710 2065 3740 2070
rect 3830 2090 3860 2095
rect 3830 2070 3835 2090
rect 3835 2070 3855 2090
rect 3855 2070 3860 2090
rect 3830 2065 3860 2070
rect 4350 2330 4380 2335
rect 4350 2310 4355 2330
rect 4355 2310 4375 2330
rect 4375 2310 4380 2330
rect 4350 2305 4380 2310
rect 4530 2285 4560 2290
rect 4530 2265 4535 2285
rect 4535 2265 4555 2285
rect 4555 2265 4560 2285
rect 4530 2260 4560 2265
rect 5275 2260 5305 2290
rect 3990 2170 4020 2200
rect 4710 2170 4740 2200
rect 4090 2115 4120 2145
rect 3990 2090 4020 2095
rect 3990 2070 3995 2090
rect 3995 2070 4015 2090
rect 4015 2070 4020 2090
rect 3990 2065 4020 2070
rect 4150 2090 4180 2095
rect 4150 2070 4155 2090
rect 4155 2070 4175 2090
rect 4175 2070 4180 2090
rect 4150 2065 4180 2070
rect 4270 2090 4300 2095
rect 4270 2070 4275 2090
rect 4275 2070 4295 2090
rect 4295 2070 4300 2090
rect 4270 2065 4300 2070
rect 4390 2090 4420 2095
rect 4390 2070 4395 2090
rect 4395 2070 4415 2090
rect 4415 2070 4420 2090
rect 4390 2065 4420 2070
rect 4510 2090 4540 2095
rect 4510 2070 4515 2090
rect 4515 2070 4535 2090
rect 4535 2070 4540 2090
rect 4510 2065 4540 2070
rect 4630 2090 4660 2095
rect 4630 2070 4635 2090
rect 4635 2070 4655 2090
rect 4655 2070 4660 2090
rect 4630 2065 4660 2070
rect 4750 2090 4780 2095
rect 4750 2070 4755 2090
rect 4755 2070 4775 2090
rect 4775 2070 4780 2090
rect 4750 2065 4780 2070
rect 4870 2090 4900 2095
rect 4870 2070 4875 2090
rect 4875 2070 4895 2090
rect 4895 2070 4900 2090
rect 4870 2065 4900 2070
rect 4990 2090 5020 2095
rect 4990 2070 4995 2090
rect 4995 2070 5015 2090
rect 5015 2070 5020 2090
rect 4990 2065 5020 2070
rect 5110 2090 5140 2095
rect 5110 2070 5115 2090
rect 5115 2070 5135 2090
rect 5135 2070 5140 2090
rect 5110 2065 5140 2070
rect 5230 2090 5260 2095
rect 5230 2070 5235 2090
rect 5235 2070 5255 2090
rect 5255 2070 5260 2090
rect 5230 2065 5260 2070
rect 2625 2045 2655 2050
rect 2625 2025 2630 2045
rect 2630 2025 2650 2045
rect 2650 2025 2655 2045
rect 2625 2020 2655 2025
rect 2810 2045 2840 2050
rect 2810 2025 2815 2045
rect 2815 2025 2835 2045
rect 2835 2025 2840 2045
rect 2810 2020 2840 2025
rect 3170 2045 3200 2050
rect 3170 2025 3175 2045
rect 3175 2025 3195 2045
rect 3195 2025 3200 2045
rect 3170 2020 3200 2025
rect 3530 2045 3560 2050
rect 3530 2025 3535 2045
rect 3535 2025 3555 2045
rect 3555 2025 3560 2045
rect 3530 2020 3560 2025
rect 3890 2045 3920 2050
rect 4090 2045 4120 2050
rect 3890 2025 3895 2045
rect 3895 2025 3915 2045
rect 3915 2025 3920 2045
rect 3890 2020 3920 2025
rect 2930 1875 2960 1880
rect 2930 1855 2935 1875
rect 2935 1855 2955 1875
rect 2955 1855 2960 1875
rect 2930 1850 2960 1855
rect 3290 1875 3320 1880
rect 3290 1855 3295 1875
rect 3295 1855 3315 1875
rect 3315 1855 3320 1875
rect 3290 1850 3320 1855
rect 3650 1875 3680 1880
rect 3650 1855 3655 1875
rect 3655 1855 3675 1875
rect 3675 1855 3680 1875
rect 3650 1850 3680 1855
rect 2570 1730 2600 1760
rect 2840 1790 2870 1820
rect 3050 1815 3080 1820
rect 3050 1795 3055 1815
rect 3055 1795 3075 1815
rect 3075 1795 3080 1815
rect 3050 1790 3080 1795
rect 3170 1790 3200 1820
rect 3410 1815 3440 1820
rect 3410 1795 3415 1815
rect 3415 1795 3435 1815
rect 3435 1795 3440 1815
rect 3410 1790 3440 1795
rect 3530 1790 3560 1820
rect 3770 1815 3800 1820
rect 3770 1795 3775 1815
rect 3775 1795 3795 1815
rect 3795 1795 3800 1815
rect 3770 1790 3800 1795
rect 3860 1790 3890 1820
rect 2680 1730 2710 1760
rect 2805 1735 2835 1765
rect 3230 1755 3260 1760
rect 3230 1735 3235 1755
rect 3235 1735 3255 1755
rect 3255 1735 3260 1755
rect 3230 1730 3260 1735
rect 3290 1755 3320 1760
rect 3290 1735 3295 1755
rect 3295 1735 3315 1755
rect 3315 1735 3320 1755
rect 3290 1730 3320 1735
rect 3530 1755 3560 1760
rect 3530 1735 3535 1755
rect 3535 1735 3555 1755
rect 3555 1735 3560 1755
rect 3530 1730 3560 1735
rect 3770 1755 3800 1760
rect 3770 1735 3775 1755
rect 3775 1735 3795 1755
rect 3795 1735 3800 1755
rect 3770 1730 3800 1735
rect 2805 1680 2835 1710
rect 3170 1710 3200 1715
rect 3170 1690 3175 1710
rect 3175 1690 3195 1710
rect 3195 1690 3200 1710
rect 3170 1685 3200 1690
rect 3410 1710 3440 1715
rect 3410 1690 3415 1710
rect 3415 1690 3435 1710
rect 3435 1690 3440 1710
rect 3410 1685 3440 1690
rect 3650 1710 3680 1715
rect 3650 1690 3655 1710
rect 3655 1690 3675 1710
rect 3675 1690 3680 1710
rect 3650 1685 3680 1690
rect 2625 1635 2655 1665
rect 3170 1590 3200 1595
rect 3170 1570 3175 1590
rect 3175 1570 3195 1590
rect 3195 1570 3200 1590
rect 3170 1565 3200 1570
rect 2840 1515 2870 1545
rect 3230 1540 3260 1545
rect 3230 1520 3235 1540
rect 3235 1520 3255 1540
rect 3255 1520 3260 1540
rect 3230 1515 3260 1520
rect 3350 1540 3380 1545
rect 3350 1520 3355 1540
rect 3355 1520 3375 1540
rect 3375 1520 3380 1540
rect 3350 1515 3380 1520
rect 3470 1540 3500 1545
rect 3470 1520 3475 1540
rect 3475 1520 3495 1540
rect 3495 1520 3500 1540
rect 3470 1515 3500 1520
rect 3590 1540 3620 1545
rect 3590 1520 3595 1540
rect 3595 1520 3615 1540
rect 3615 1520 3620 1540
rect 3590 1515 3620 1520
rect 3710 1540 3740 1545
rect 3710 1520 3715 1540
rect 3715 1520 3735 1540
rect 3735 1520 3740 1540
rect 3710 1515 3740 1520
rect 2930 1495 2960 1500
rect 2930 1475 2935 1495
rect 2935 1475 2955 1495
rect 2955 1475 2960 1495
rect 2930 1470 2960 1475
rect 3050 1495 3080 1500
rect 3050 1475 3055 1495
rect 3055 1475 3075 1495
rect 3075 1475 3080 1495
rect 3050 1470 3080 1475
rect 3170 1495 3200 1500
rect 3170 1475 3175 1495
rect 3175 1475 3195 1495
rect 3195 1475 3200 1495
rect 3170 1470 3200 1475
rect 3290 1495 3320 1500
rect 3290 1475 3295 1495
rect 3295 1475 3315 1495
rect 3315 1475 3320 1495
rect 3290 1470 3320 1475
rect 3530 1495 3560 1500
rect 3530 1475 3535 1495
rect 3535 1475 3555 1495
rect 3555 1475 3560 1495
rect 3530 1470 3560 1475
rect 3650 1495 3680 1500
rect 3650 1475 3655 1495
rect 3655 1475 3675 1495
rect 3675 1475 3680 1495
rect 3650 1470 3680 1475
rect 3770 1495 3800 1500
rect 3770 1475 3775 1495
rect 3775 1475 3795 1495
rect 3795 1475 3800 1495
rect 3770 1470 3800 1475
rect 4090 2025 4095 2045
rect 4095 2025 4115 2045
rect 4115 2025 4120 2045
rect 4090 2020 4120 2025
rect 4450 2045 4480 2050
rect 4450 2025 4455 2045
rect 4455 2025 4475 2045
rect 4475 2025 4480 2045
rect 4450 2020 4480 2025
rect 4810 2045 4840 2050
rect 4810 2025 4815 2045
rect 4815 2025 4835 2045
rect 4835 2025 4840 2045
rect 4810 2020 4840 2025
rect 5170 2045 5200 2050
rect 5170 2025 5175 2045
rect 5175 2025 5195 2045
rect 5195 2025 5200 2045
rect 5170 2020 5200 2025
rect 4330 1875 4360 1880
rect 4330 1855 4335 1875
rect 4335 1855 4355 1875
rect 4355 1855 4360 1875
rect 4330 1850 4360 1855
rect 4690 1875 4720 1880
rect 4690 1855 4695 1875
rect 4695 1855 4715 1875
rect 4715 1855 4720 1875
rect 4690 1850 4720 1855
rect 5050 1875 5080 1880
rect 5050 1855 5055 1875
rect 5055 1855 5075 1875
rect 5075 1855 5080 1875
rect 5050 1850 5080 1855
rect 4120 1790 4150 1820
rect 4210 1815 4240 1820
rect 4210 1795 4215 1815
rect 4215 1795 4235 1815
rect 4235 1795 4240 1815
rect 4210 1790 4240 1795
rect 4450 1790 4480 1820
rect 4570 1815 4600 1820
rect 4570 1795 4575 1815
rect 4575 1795 4595 1815
rect 4595 1795 4600 1815
rect 4570 1790 4600 1795
rect 4210 1755 4240 1760
rect 4210 1735 4215 1755
rect 4215 1735 4235 1755
rect 4235 1735 4240 1755
rect 4210 1730 4240 1735
rect 4450 1755 4480 1760
rect 4450 1735 4455 1755
rect 4455 1735 4475 1755
rect 4475 1735 4480 1755
rect 4450 1730 4480 1735
rect 4810 1790 4840 1820
rect 4930 1815 4960 1820
rect 4930 1795 4935 1815
rect 4935 1795 4955 1815
rect 4955 1795 4960 1815
rect 4930 1790 4960 1795
rect 5140 1790 5170 1820
rect 5320 2115 5350 2145
rect 5415 3255 5445 3285
rect 5365 1790 5395 1820
rect 4690 1755 4720 1760
rect 4690 1735 4695 1755
rect 4695 1735 4715 1755
rect 4715 1735 4720 1755
rect 4690 1730 4720 1735
rect 4750 1755 4780 1760
rect 4750 1735 4755 1755
rect 4755 1735 4775 1755
rect 4775 1735 4780 1755
rect 4750 1730 4780 1735
rect 5275 1730 5305 1760
rect 4330 1710 4360 1715
rect 4330 1690 4335 1710
rect 4335 1690 4355 1710
rect 4355 1690 4360 1710
rect 4330 1685 4360 1690
rect 4570 1710 4600 1715
rect 4570 1690 4575 1710
rect 4575 1690 4595 1710
rect 4595 1690 4600 1710
rect 4570 1685 4600 1690
rect 4810 1710 4840 1715
rect 4810 1690 4815 1710
rect 4815 1690 4835 1710
rect 4835 1690 4840 1710
rect 4810 1685 4840 1690
rect 17145 4310 17175 4315
rect 17145 4290 17150 4310
rect 17150 4290 17170 4310
rect 17170 4290 17175 4310
rect 17145 4285 17175 4290
rect 17265 4310 17295 4315
rect 17265 4290 17270 4310
rect 17270 4290 17290 4310
rect 17290 4290 17295 4310
rect 17265 4285 17295 4290
rect 17385 4310 17415 4315
rect 17385 4290 17390 4310
rect 17390 4290 17410 4310
rect 17410 4290 17415 4310
rect 17385 4285 17415 4290
rect 17505 4310 17535 4315
rect 17505 4290 17510 4310
rect 17510 4290 17530 4310
rect 17530 4290 17535 4310
rect 17505 4285 17535 4290
rect 16110 4230 16140 4260
rect 16335 4230 16365 4260
rect 17205 4230 17235 4260
rect 16055 3125 16085 3155
rect 14910 2905 14940 2935
rect 14960 2905 14990 2935
rect 15010 2905 15040 2935
rect 15270 2960 15300 2965
rect 15270 2940 15275 2960
rect 15275 2940 15295 2960
rect 15295 2940 15300 2960
rect 15270 2935 15300 2940
rect 15380 2960 15410 2965
rect 15380 2940 15385 2960
rect 15385 2940 15405 2960
rect 15405 2940 15410 2960
rect 15380 2935 15410 2940
rect 15490 2960 15520 2965
rect 15490 2940 15495 2960
rect 15495 2940 15515 2960
rect 15515 2940 15520 2960
rect 15490 2935 15520 2940
rect 15600 2960 15630 2965
rect 15600 2940 15605 2960
rect 15605 2940 15625 2960
rect 15625 2940 15630 2960
rect 15600 2935 15630 2940
rect 15710 2960 15740 2965
rect 15710 2940 15715 2960
rect 15715 2940 15735 2960
rect 15735 2940 15740 2960
rect 15710 2935 15740 2940
rect 14960 2850 14990 2880
rect 15655 2850 15685 2880
rect 16005 2850 16035 2880
rect 14520 2795 14550 2825
rect 15380 2795 15410 2825
rect 15215 2700 15245 2705
rect 15215 2680 15220 2700
rect 15220 2680 15240 2700
rect 15240 2680 15245 2700
rect 15215 2675 15245 2680
rect 15325 2700 15355 2705
rect 15325 2680 15330 2700
rect 15330 2680 15350 2700
rect 15350 2680 15355 2700
rect 15325 2675 15355 2680
rect 15435 2700 15465 2705
rect 15435 2680 15440 2700
rect 15440 2680 15460 2700
rect 15460 2680 15465 2700
rect 15435 2675 15465 2680
rect 15545 2700 15575 2705
rect 15545 2680 15550 2700
rect 15550 2680 15570 2700
rect 15570 2680 15575 2700
rect 15545 2675 15575 2680
rect 15655 2700 15685 2705
rect 15655 2680 15660 2700
rect 15660 2680 15680 2700
rect 15680 2680 15685 2700
rect 15655 2675 15685 2680
rect 15765 2700 15795 2705
rect 15765 2680 15770 2700
rect 15770 2680 15790 2700
rect 15790 2680 15795 2700
rect 15765 2675 15795 2680
rect 15025 2405 15055 2435
rect 15270 2430 15300 2435
rect 15270 2410 15275 2430
rect 15275 2410 15295 2430
rect 15295 2410 15300 2430
rect 15270 2405 15300 2410
rect 15380 2430 15410 2435
rect 15380 2410 15385 2430
rect 15385 2410 15405 2430
rect 15405 2410 15410 2430
rect 15380 2405 15410 2410
rect 15490 2430 15520 2435
rect 15490 2410 15495 2430
rect 15495 2410 15515 2430
rect 15515 2410 15520 2430
rect 15490 2405 15520 2410
rect 15600 2430 15630 2435
rect 15600 2410 15605 2430
rect 15605 2410 15625 2430
rect 15625 2410 15630 2430
rect 15600 2405 15630 2410
rect 15710 2430 15740 2435
rect 15710 2410 15715 2430
rect 15715 2410 15735 2430
rect 15735 2410 15740 2430
rect 15710 2405 15740 2410
rect 16365 4200 16395 4205
rect 16365 4180 16370 4200
rect 16370 4180 16390 4200
rect 16390 4180 16395 4200
rect 16365 4175 16395 4180
rect 16475 4200 16505 4205
rect 16475 4180 16480 4200
rect 16480 4180 16500 4200
rect 16500 4180 16505 4200
rect 16475 4175 16505 4180
rect 16585 4200 16615 4205
rect 16585 4180 16590 4200
rect 16590 4180 16610 4200
rect 16610 4180 16615 4200
rect 16585 4175 16615 4180
rect 16695 4200 16725 4205
rect 16695 4180 16700 4200
rect 16700 4180 16720 4200
rect 16720 4180 16725 4200
rect 16695 4175 16725 4180
rect 16805 4200 16835 4205
rect 16805 4180 16810 4200
rect 16810 4180 16830 4200
rect 16830 4180 16835 4200
rect 16805 4175 16835 4180
rect 16915 4200 16945 4205
rect 16915 4180 16920 4200
rect 16920 4180 16940 4200
rect 16940 4180 16945 4200
rect 16915 4175 16945 4180
rect 17025 4200 17055 4205
rect 17025 4180 17030 4200
rect 17030 4180 17050 4200
rect 17050 4180 17055 4200
rect 17025 4175 17055 4180
rect 17135 4200 17165 4205
rect 17135 4180 17140 4200
rect 17140 4180 17160 4200
rect 17160 4180 17165 4200
rect 17135 4175 17165 4180
rect 17245 4200 17275 4205
rect 17245 4180 17250 4200
rect 17250 4180 17270 4200
rect 17270 4180 17275 4200
rect 17245 4175 17275 4180
rect 17355 4200 17385 4205
rect 17355 4180 17360 4200
rect 17360 4180 17380 4200
rect 17380 4180 17385 4200
rect 17355 4175 17385 4180
rect 16310 4080 16340 4085
rect 16310 4060 16315 4080
rect 16315 4060 16335 4080
rect 16335 4060 16340 4080
rect 16310 4055 16340 4060
rect 16530 4080 16560 4085
rect 16530 4060 16535 4080
rect 16535 4060 16555 4080
rect 16555 4060 16560 4080
rect 16530 4055 16560 4060
rect 16750 4080 16780 4085
rect 16750 4060 16755 4080
rect 16755 4060 16775 4080
rect 16775 4060 16780 4080
rect 16750 4055 16780 4060
rect 16970 4080 17000 4085
rect 16970 4060 16975 4080
rect 16975 4060 16995 4080
rect 16995 4060 17000 4080
rect 16970 4055 17000 4060
rect 17190 4080 17220 4085
rect 17190 4060 17195 4080
rect 17195 4060 17215 4080
rect 17215 4060 17220 4080
rect 17190 4055 17220 4060
rect 17410 4080 17440 4085
rect 17410 4060 17415 4080
rect 17415 4060 17435 4080
rect 17435 4060 17440 4080
rect 17410 4055 17440 4060
rect 16315 3955 16345 3960
rect 16315 3935 16320 3955
rect 16320 3935 16340 3955
rect 16340 3935 16345 3955
rect 16315 3930 16345 3935
rect 16420 3995 16450 4025
rect 16640 3995 16670 4025
rect 16860 3995 16890 4025
rect 17080 3995 17110 4025
rect 17300 3995 17330 4025
rect 16420 3955 16450 3960
rect 16420 3935 16425 3955
rect 16425 3935 16445 3955
rect 16445 3935 16450 3955
rect 16420 3930 16450 3935
rect 16530 3955 16560 3960
rect 16530 3935 16535 3955
rect 16535 3935 16555 3955
rect 16555 3935 16560 3955
rect 16530 3930 16560 3935
rect 16640 3955 16670 3960
rect 16640 3935 16645 3955
rect 16645 3935 16665 3955
rect 16665 3935 16670 3955
rect 16640 3930 16670 3935
rect 16750 3955 16780 3960
rect 16750 3935 16755 3955
rect 16755 3935 16775 3955
rect 16775 3935 16780 3955
rect 16750 3930 16780 3935
rect 17055 3955 17085 3960
rect 17055 3935 17060 3955
rect 17060 3935 17080 3955
rect 17080 3935 17085 3955
rect 17055 3930 17085 3935
rect 17160 3955 17190 3960
rect 17160 3935 17165 3955
rect 17165 3935 17185 3955
rect 17185 3935 17190 3955
rect 17160 3930 17190 3935
rect 17270 3955 17300 3960
rect 17270 3935 17275 3955
rect 17275 3935 17295 3955
rect 17295 3935 17300 3955
rect 17270 3930 17300 3935
rect 17380 3955 17410 3960
rect 17380 3935 17385 3955
rect 17385 3935 17405 3955
rect 17405 3935 17410 3955
rect 17380 3930 17410 3935
rect 17490 3955 17520 3960
rect 17490 3935 17495 3955
rect 17495 3935 17515 3955
rect 17515 3935 17520 3955
rect 17490 3930 17520 3935
rect 16274 3895 16300 3900
rect 16274 3875 16277 3895
rect 16277 3875 16294 3895
rect 16294 3875 16300 3895
rect 16274 3870 16300 3875
rect 16475 3895 16505 3900
rect 16475 3875 16480 3895
rect 16480 3875 16500 3895
rect 16500 3875 16505 3895
rect 16475 3870 16505 3875
rect 16695 3895 16725 3900
rect 16695 3875 16700 3895
rect 16700 3875 16720 3895
rect 16720 3875 16725 3895
rect 16695 3870 16725 3875
rect 17014 3895 17040 3900
rect 17014 3875 17017 3895
rect 17017 3875 17034 3895
rect 17034 3875 17040 3895
rect 17014 3870 17040 3875
rect 17215 3895 17245 3900
rect 17215 3875 17220 3895
rect 17220 3875 17240 3895
rect 17240 3875 17245 3895
rect 17215 3870 17245 3875
rect 17435 3895 17465 3900
rect 17435 3875 17440 3895
rect 17440 3875 17460 3895
rect 17460 3875 17465 3895
rect 17435 3870 17465 3875
rect 17765 3870 17795 3900
rect 16405 3775 16431 3780
rect 16405 3755 16408 3775
rect 16408 3755 16425 3775
rect 16425 3755 16431 3775
rect 16405 3750 16431 3755
rect 16625 3775 16651 3780
rect 16625 3755 16628 3775
rect 16628 3755 16645 3775
rect 16645 3755 16651 3775
rect 16625 3750 16651 3755
rect 16769 3775 16795 3780
rect 16769 3755 16775 3775
rect 16775 3755 16792 3775
rect 16792 3755 16795 3775
rect 16769 3750 16795 3755
rect 17145 3775 17171 3780
rect 17145 3755 17148 3775
rect 17148 3755 17165 3775
rect 17165 3755 17171 3775
rect 17145 3750 17171 3755
rect 17365 3775 17391 3780
rect 17365 3755 17368 3775
rect 17368 3755 17385 3775
rect 17385 3755 17391 3775
rect 17365 3750 17391 3755
rect 17509 3775 17535 3780
rect 17509 3755 17515 3775
rect 17515 3755 17532 3775
rect 17532 3755 17535 3775
rect 17509 3750 17535 3755
rect 16255 3715 16285 3720
rect 16255 3695 16260 3715
rect 16260 3695 16280 3715
rect 16280 3695 16285 3715
rect 16255 3690 16285 3695
rect 16360 3715 16390 3720
rect 16360 3695 16365 3715
rect 16365 3695 16385 3715
rect 16385 3695 16390 3715
rect 16360 3690 16390 3695
rect 16475 3715 16505 3720
rect 16475 3695 16480 3715
rect 16480 3695 16500 3715
rect 16500 3695 16505 3715
rect 16475 3690 16505 3695
rect 16580 3715 16610 3720
rect 16580 3695 16585 3715
rect 16585 3695 16605 3715
rect 16605 3695 16610 3715
rect 16580 3690 16610 3695
rect 16695 3715 16725 3720
rect 16695 3695 16700 3715
rect 16700 3695 16720 3715
rect 16720 3695 16725 3715
rect 16695 3690 16725 3695
rect 16810 3715 16840 3720
rect 16810 3695 16815 3715
rect 16815 3695 16835 3715
rect 16835 3695 16840 3715
rect 16810 3690 16840 3695
rect 16995 3725 17025 3730
rect 16995 3705 17000 3725
rect 17000 3705 17020 3725
rect 17020 3705 17025 3725
rect 16995 3700 17025 3705
rect 17215 3725 17245 3730
rect 17215 3705 17220 3725
rect 17220 3705 17240 3725
rect 17240 3705 17245 3725
rect 17215 3700 17245 3705
rect 17435 3725 17465 3730
rect 17435 3705 17440 3725
rect 17440 3705 17460 3725
rect 17460 3705 17465 3725
rect 17435 3700 17465 3705
rect 17100 3655 17130 3685
rect 17320 3655 17350 3685
rect 17550 3655 17580 3685
rect 16345 3620 16375 3625
rect 16345 3600 16350 3620
rect 16350 3600 16370 3620
rect 16370 3600 16375 3620
rect 16345 3595 16375 3600
rect 16465 3620 16495 3625
rect 16465 3600 16470 3620
rect 16470 3600 16490 3620
rect 16490 3600 16495 3620
rect 16465 3595 16495 3600
rect 16585 3620 16615 3625
rect 16585 3600 16590 3620
rect 16590 3600 16610 3620
rect 16610 3600 16615 3620
rect 16585 3595 16615 3600
rect 16705 3620 16735 3625
rect 16705 3600 16710 3620
rect 16710 3600 16730 3620
rect 16730 3600 16735 3620
rect 16705 3595 16735 3600
rect 16825 3620 16855 3625
rect 16825 3600 16830 3620
rect 16830 3600 16850 3620
rect 16850 3600 16855 3620
rect 16825 3595 16855 3600
rect 16945 3620 16975 3625
rect 16945 3600 16950 3620
rect 16950 3600 16970 3620
rect 16970 3600 16975 3620
rect 16945 3595 16975 3600
rect 17065 3620 17095 3625
rect 17065 3600 17070 3620
rect 17070 3600 17090 3620
rect 17090 3600 17095 3620
rect 17065 3595 17095 3600
rect 17185 3620 17215 3625
rect 17185 3600 17190 3620
rect 17190 3600 17210 3620
rect 17210 3600 17215 3620
rect 17185 3595 17215 3600
rect 17305 3620 17335 3625
rect 17305 3600 17310 3620
rect 17310 3600 17330 3620
rect 17330 3600 17335 3620
rect 17305 3595 17335 3600
rect 17425 3620 17455 3625
rect 17425 3600 17430 3620
rect 17430 3600 17450 3620
rect 17450 3600 17455 3620
rect 17425 3595 17455 3600
rect 16826 3150 16854 3155
rect 16826 3130 16831 3150
rect 16831 3130 16849 3150
rect 16849 3130 16854 3150
rect 16826 3125 16854 3130
rect 16285 3070 16315 3100
rect 16525 3070 16555 3100
rect 16765 3070 16795 3100
rect 17005 3070 17035 3100
rect 17245 3070 17275 3100
rect 17485 3070 17515 3100
rect 16405 3025 16435 3055
rect 16645 3025 16675 3055
rect 16885 3025 16915 3055
rect 17125 3025 17155 3055
rect 17365 3025 17395 3055
rect 16345 2970 16375 3000
rect 16405 2970 16435 3000
rect 16585 2970 16615 3000
rect 16825 2970 16855 3000
rect 17065 2970 17095 3000
rect 17305 2970 17335 3000
rect 16465 2940 16495 2945
rect 16465 2920 16470 2940
rect 16470 2920 16490 2940
rect 16490 2920 16495 2940
rect 16465 2915 16495 2920
rect 16705 2940 16735 2945
rect 16705 2920 16710 2940
rect 16710 2920 16730 2940
rect 16730 2920 16735 2940
rect 16705 2915 16735 2920
rect 16945 2940 16975 2945
rect 16945 2920 16950 2940
rect 16950 2920 16970 2940
rect 16970 2920 16975 2940
rect 16945 2915 16975 2920
rect 17185 2940 17215 2945
rect 17185 2920 17190 2940
rect 17190 2920 17210 2940
rect 17210 2920 17215 2940
rect 17185 2915 17215 2920
rect 17425 2940 17455 2945
rect 17425 2920 17430 2940
rect 17430 2920 17450 2940
rect 17450 2920 17455 2940
rect 17425 2915 17455 2920
rect 17485 2915 17515 2945
rect 17695 2850 17725 2880
rect 16110 2445 16140 2475
rect 16826 2470 16854 2475
rect 16826 2450 16831 2470
rect 16831 2450 16849 2470
rect 16849 2450 16854 2470
rect 16826 2445 16854 2450
rect 14520 2080 14550 2110
rect 14790 2000 14825 2005
rect 14790 1975 14795 2000
rect 14795 1975 14820 2000
rect 14820 1975 14825 2000
rect 14790 1970 14825 1975
rect 14850 2000 14885 2005
rect 14850 1975 14855 2000
rect 14855 1975 14880 2000
rect 14880 1975 14885 2000
rect 14850 1970 14885 1975
rect 14910 2000 14945 2005
rect 14910 1975 14915 2000
rect 14915 1975 14940 2000
rect 14940 1975 14945 2000
rect 14910 1970 14945 1975
rect 15770 2385 15800 2390
rect 15770 2365 15775 2385
rect 15775 2365 15795 2385
rect 15795 2365 15800 2385
rect 15770 2360 15800 2365
rect 16005 2390 16035 2420
rect 16285 2390 16315 2420
rect 16525 2390 16555 2420
rect 16765 2390 16795 2420
rect 16405 2345 16435 2375
rect 16645 2345 16675 2375
rect 15070 2285 15100 2315
rect 15270 2310 15300 2315
rect 15270 2290 15275 2310
rect 15275 2290 15295 2310
rect 15295 2290 15300 2310
rect 15270 2285 15300 2290
rect 15380 2310 15410 2315
rect 15380 2290 15385 2310
rect 15385 2290 15405 2310
rect 15405 2290 15410 2310
rect 15380 2285 15410 2290
rect 15490 2310 15520 2315
rect 15490 2290 15495 2310
rect 15495 2290 15515 2310
rect 15515 2290 15520 2310
rect 15490 2285 15520 2290
rect 15600 2310 15630 2315
rect 15600 2290 15605 2310
rect 15605 2290 15625 2310
rect 15625 2290 15630 2310
rect 15600 2285 15630 2290
rect 15710 2310 15740 2315
rect 15710 2290 15715 2310
rect 15715 2290 15735 2310
rect 15735 2290 15740 2310
rect 15710 2285 15740 2290
rect 16005 2295 16035 2325
rect 14970 2000 15005 2005
rect 14970 1975 14975 2000
rect 14975 1975 15000 2000
rect 15000 1975 15005 2000
rect 14970 1970 15005 1975
rect 15025 1970 15055 2000
rect 15955 2150 15985 2180
rect 14915 1915 14945 1945
rect 15070 1915 15100 1945
rect 15215 1940 15245 1945
rect 15215 1920 15220 1940
rect 15220 1920 15238 1940
rect 15238 1920 15245 1940
rect 15215 1915 15245 1920
rect 15325 1940 15355 1945
rect 15325 1920 15330 1940
rect 15330 1920 15348 1940
rect 15348 1920 15355 1940
rect 15325 1915 15355 1920
rect 15435 1940 15465 1945
rect 15435 1920 15440 1940
rect 15440 1920 15458 1940
rect 15458 1920 15465 1940
rect 15435 1915 15465 1920
rect 15545 1940 15575 1945
rect 15545 1920 15550 1940
rect 15550 1920 15568 1940
rect 15568 1920 15575 1940
rect 15545 1915 15575 1920
rect 15655 1940 15685 1945
rect 15655 1920 15660 1940
rect 15660 1920 15678 1940
rect 15678 1920 15685 1940
rect 15655 1915 15685 1920
rect 15765 1940 15795 1945
rect 15765 1920 15770 1940
rect 15770 1920 15788 1940
rect 15788 1920 15795 1940
rect 15765 1915 15795 1920
rect 14795 1865 14825 1895
rect 14970 1730 15000 1760
rect 15560 1730 15590 1760
rect 15840 1730 15870 1760
rect 14520 1675 14550 1705
rect 15035 1675 15065 1705
rect 15260 1700 15290 1705
rect 15260 1680 15265 1700
rect 15265 1680 15285 1700
rect 15285 1680 15290 1700
rect 15260 1675 15290 1680
rect 15460 1700 15490 1705
rect 15460 1680 15465 1700
rect 15465 1680 15485 1700
rect 15485 1680 15490 1700
rect 15460 1675 15490 1680
rect 15660 1700 15690 1705
rect 15660 1680 15665 1700
rect 15665 1680 15685 1700
rect 15685 1680 15690 1700
rect 15660 1675 15690 1680
rect 14970 1640 15005 1645
rect 14970 1615 14975 1640
rect 14975 1615 15000 1640
rect 15000 1615 15005 1640
rect 14970 1610 15005 1615
rect 15030 1640 15065 1645
rect 15030 1615 15035 1640
rect 15035 1615 15060 1640
rect 15060 1615 15065 1640
rect 15030 1610 15065 1615
rect 4810 1590 4840 1595
rect 4810 1570 4815 1590
rect 4815 1570 4835 1590
rect 4835 1570 4840 1590
rect 4810 1565 4840 1570
rect 5415 1565 5445 1595
rect 4270 1540 4300 1545
rect 4270 1520 4275 1540
rect 4275 1520 4295 1540
rect 4295 1520 4300 1540
rect 4270 1515 4300 1520
rect 4390 1540 4420 1545
rect 4390 1520 4395 1540
rect 4395 1520 4415 1540
rect 4415 1520 4420 1540
rect 4390 1515 4420 1520
rect 4510 1540 4540 1545
rect 4510 1520 4515 1540
rect 4515 1520 4535 1540
rect 4535 1520 4540 1540
rect 4510 1515 4540 1520
rect 4630 1540 4660 1545
rect 4630 1520 4635 1540
rect 4635 1520 4655 1540
rect 4655 1520 4660 1540
rect 4630 1515 4660 1520
rect 4750 1540 4780 1545
rect 4750 1520 4755 1540
rect 4755 1520 4775 1540
rect 4775 1520 4780 1540
rect 4750 1515 4780 1520
rect 5140 1515 5170 1545
rect 4210 1495 4240 1500
rect 4210 1475 4215 1495
rect 4215 1475 4235 1495
rect 4235 1475 4240 1495
rect 4210 1470 4240 1475
rect 4330 1495 4360 1500
rect 4330 1475 4335 1495
rect 4335 1475 4355 1495
rect 4355 1475 4360 1495
rect 4330 1470 4360 1475
rect 4450 1495 4480 1500
rect 4450 1475 4455 1495
rect 4455 1475 4475 1495
rect 4475 1475 4480 1495
rect 4450 1470 4480 1475
rect 4690 1495 4720 1500
rect 4690 1475 4695 1495
rect 4695 1475 4715 1495
rect 4715 1475 4720 1495
rect 4690 1470 4720 1475
rect 4810 1495 4840 1500
rect 4810 1475 4815 1495
rect 4815 1475 4835 1495
rect 4835 1475 4840 1495
rect 4810 1470 4840 1475
rect 4930 1495 4960 1500
rect 4930 1475 4935 1495
rect 4935 1475 4955 1495
rect 4955 1475 4960 1495
rect 4930 1470 4960 1475
rect 5050 1495 5080 1500
rect 5050 1475 5055 1495
rect 5055 1475 5075 1495
rect 5075 1475 5080 1495
rect 5050 1470 5080 1475
rect 15840 1360 15870 1390
rect 3380 1180 3410 1185
rect 3380 1160 3385 1180
rect 3385 1160 3405 1180
rect 3405 1160 3410 1180
rect 3380 1155 3410 1160
rect 3990 1155 4020 1185
rect 4600 1180 4630 1185
rect 4600 1160 4605 1180
rect 4605 1160 4625 1180
rect 4625 1160 4630 1180
rect 4600 1155 4630 1160
rect 2950 1120 2980 1125
rect 2950 1100 2955 1120
rect 2955 1100 2975 1120
rect 2975 1100 2980 1120
rect 2950 1095 2980 1100
rect 3030 1120 3060 1125
rect 3030 1100 3035 1120
rect 3035 1100 3055 1120
rect 3055 1100 3060 1120
rect 3030 1095 3060 1100
rect 3110 1120 3140 1125
rect 3110 1100 3115 1120
rect 3115 1100 3135 1120
rect 3135 1100 3140 1120
rect 3110 1095 3140 1100
rect 3190 1120 3220 1125
rect 3190 1100 3195 1120
rect 3195 1100 3215 1120
rect 3215 1100 3220 1120
rect 3190 1095 3220 1100
rect 3270 1120 3300 1125
rect 3270 1100 3275 1120
rect 3275 1100 3295 1120
rect 3295 1100 3300 1120
rect 3270 1095 3300 1100
rect 3350 1120 3380 1125
rect 3350 1100 3355 1120
rect 3355 1100 3375 1120
rect 3375 1100 3380 1120
rect 3350 1095 3380 1100
rect 3430 1120 3460 1125
rect 3430 1100 3435 1120
rect 3435 1100 3455 1120
rect 3455 1100 3460 1120
rect 3430 1095 3460 1100
rect 3510 1120 3540 1125
rect 3510 1100 3515 1120
rect 3515 1100 3535 1120
rect 3535 1100 3540 1120
rect 3510 1095 3540 1100
rect 3590 1120 3620 1125
rect 3590 1100 3595 1120
rect 3595 1100 3615 1120
rect 3615 1100 3620 1120
rect 3590 1095 3620 1100
rect 3670 1120 3700 1125
rect 3670 1100 3675 1120
rect 3675 1100 3695 1120
rect 3695 1100 3700 1120
rect 3670 1095 3700 1100
rect 3750 1120 3780 1125
rect 3750 1100 3755 1120
rect 3755 1100 3775 1120
rect 3775 1100 3780 1120
rect 3750 1095 3780 1100
rect 3830 1120 3860 1125
rect 3830 1100 3835 1120
rect 3835 1100 3855 1120
rect 3855 1100 3860 1120
rect 3830 1095 3860 1100
rect 3910 1120 3940 1125
rect 3910 1100 3915 1120
rect 3915 1100 3935 1120
rect 3935 1100 3940 1120
rect 3910 1095 3940 1100
rect 3990 1120 4020 1125
rect 3990 1100 3995 1120
rect 3995 1100 4015 1120
rect 4015 1100 4020 1120
rect 3990 1095 4020 1100
rect 4070 1120 4100 1125
rect 4070 1100 4075 1120
rect 4075 1100 4095 1120
rect 4095 1100 4100 1120
rect 4070 1095 4100 1100
rect 4150 1120 4180 1125
rect 4150 1100 4155 1120
rect 4155 1100 4175 1120
rect 4175 1100 4180 1120
rect 4150 1095 4180 1100
rect 4230 1120 4260 1125
rect 4230 1100 4235 1120
rect 4235 1100 4255 1120
rect 4255 1100 4260 1120
rect 4230 1095 4260 1100
rect 4310 1120 4340 1125
rect 4310 1100 4315 1120
rect 4315 1100 4335 1120
rect 4335 1100 4340 1120
rect 4310 1095 4340 1100
rect 4390 1120 4420 1125
rect 4390 1100 4395 1120
rect 4395 1100 4415 1120
rect 4415 1100 4420 1120
rect 4390 1095 4420 1100
rect 4470 1120 4500 1125
rect 4470 1100 4475 1120
rect 4475 1100 4495 1120
rect 4495 1100 4500 1120
rect 4470 1095 4500 1100
rect 4550 1120 4580 1125
rect 4550 1100 4555 1120
rect 4555 1100 4575 1120
rect 4575 1100 4580 1120
rect 4550 1095 4580 1100
rect 4630 1120 4660 1125
rect 4630 1100 4635 1120
rect 4635 1100 4655 1120
rect 4655 1100 4660 1120
rect 4630 1095 4660 1100
rect 4710 1120 4740 1125
rect 4710 1100 4715 1120
rect 4715 1100 4735 1120
rect 4735 1100 4740 1120
rect 4710 1095 4740 1100
rect 4790 1120 4820 1125
rect 4790 1100 4795 1120
rect 4795 1100 4815 1120
rect 4815 1100 4820 1120
rect 4790 1095 4820 1100
rect 4870 1120 4900 1125
rect 4870 1100 4875 1120
rect 4875 1100 4895 1120
rect 4895 1100 4900 1120
rect 4870 1095 4900 1100
rect 4950 1120 4980 1125
rect 4950 1100 4955 1120
rect 4955 1100 4975 1120
rect 4975 1100 4980 1120
rect 4950 1095 4980 1100
rect 2625 1010 2655 1040
rect 2910 1035 2940 1040
rect 2910 1015 2915 1035
rect 2915 1015 2935 1035
rect 2935 1015 2940 1035
rect 2910 1010 2940 1015
rect 5115 1035 5145 1040
rect 5115 1015 5120 1035
rect 5120 1015 5140 1035
rect 5140 1015 5145 1035
rect 5115 1010 5145 1015
rect 3000 925 3030 930
rect 3000 905 3005 925
rect 3005 905 3025 925
rect 3025 905 3030 925
rect 3000 900 3030 905
rect 3180 925 3210 930
rect 3180 905 3185 925
rect 3185 905 3205 925
rect 3205 905 3210 925
rect 3180 900 3210 905
rect 3360 925 3390 930
rect 3360 905 3365 925
rect 3365 905 3385 925
rect 3385 905 3390 925
rect 3360 900 3390 905
rect 3540 925 3570 930
rect 3540 905 3545 925
rect 3545 905 3565 925
rect 3565 905 3570 925
rect 3540 900 3570 905
rect 3720 925 3750 930
rect 3720 905 3725 925
rect 3725 905 3745 925
rect 3745 905 3750 925
rect 3720 900 3750 905
rect 3900 925 3930 930
rect 3900 905 3905 925
rect 3905 905 3925 925
rect 3925 905 3930 925
rect 3900 900 3930 905
rect 4080 925 4110 930
rect 4080 905 4085 925
rect 4085 905 4105 925
rect 4105 905 4110 925
rect 4080 900 4110 905
rect 4260 925 4290 930
rect 4260 905 4265 925
rect 4265 905 4285 925
rect 4285 905 4290 925
rect 4260 900 4290 905
rect 4440 925 4470 930
rect 4440 905 4445 925
rect 4445 905 4465 925
rect 4465 905 4470 925
rect 4440 900 4470 905
rect 4620 925 4650 930
rect 4620 905 4625 925
rect 4625 905 4645 925
rect 4645 905 4650 925
rect 4620 900 4650 905
rect 4800 925 4830 930
rect 4800 905 4805 925
rect 4805 905 4825 925
rect 4825 905 4830 925
rect 4800 900 4830 905
rect 4980 925 5010 930
rect 4980 905 4985 925
rect 4985 905 5005 925
rect 5005 905 5010 925
rect 4980 900 5010 905
rect 15360 930 15390 935
rect 15360 910 15365 930
rect 15365 910 15385 930
rect 15385 910 15390 930
rect 15360 905 15390 910
rect 15560 930 15590 935
rect 15560 910 15565 930
rect 15565 910 15585 930
rect 15585 910 15590 930
rect 15560 905 15590 910
rect 16445 2250 16475 2280
rect 16665 2250 16695 2280
rect 16335 2205 16365 2235
rect 16555 2205 16585 2235
rect 17005 2390 17035 2420
rect 17245 2390 17275 2420
rect 17485 2390 17515 2420
rect 16885 2345 16915 2375
rect 17125 2345 17155 2375
rect 17365 2345 17395 2375
rect 17695 2345 17725 2375
rect 17865 3700 17895 3730
rect 17810 3655 17840 3685
rect 17765 2295 17795 2325
rect 16885 2250 16915 2280
rect 17105 2250 17135 2280
rect 17325 2250 17355 2280
rect 16775 2205 16805 2235
rect 16995 2205 17025 2235
rect 17215 2205 17245 2235
rect 17435 2205 17465 2235
rect 16831 2175 16859 2180
rect 16831 2155 16836 2175
rect 16836 2155 16854 2175
rect 16854 2155 16859 2175
rect 16831 2150 16859 2155
rect 16390 1955 16420 1960
rect 16390 1935 16395 1955
rect 16395 1935 16415 1955
rect 16415 1935 16420 1955
rect 16390 1930 16420 1935
rect 16610 1955 16640 1960
rect 16610 1935 16615 1955
rect 16615 1935 16635 1955
rect 16635 1935 16640 1955
rect 16610 1930 16640 1935
rect 16830 1955 16860 1960
rect 16830 1935 16835 1955
rect 16835 1935 16855 1955
rect 16855 1935 16860 1955
rect 16830 1930 16860 1935
rect 17050 1955 17080 1960
rect 17050 1935 17055 1955
rect 17055 1935 17075 1955
rect 17075 1935 17080 1955
rect 17050 1930 17080 1935
rect 17270 1955 17300 1960
rect 17270 1935 17275 1955
rect 17275 1935 17295 1955
rect 17295 1935 17300 1955
rect 17270 1930 17300 1935
rect 16005 1865 16035 1895
rect 16500 1875 16530 1905
rect 16720 1875 16750 1905
rect 16940 1875 16970 1905
rect 17160 1875 17190 1905
rect 16195 1820 16225 1850
rect 16415 1820 16445 1850
rect 16090 1755 16120 1760
rect 16090 1735 16095 1755
rect 16095 1735 16115 1755
rect 16115 1735 16120 1755
rect 16090 1730 16120 1735
rect 16310 1755 16340 1760
rect 16310 1735 16315 1755
rect 16315 1735 16335 1755
rect 16335 1735 16340 1755
rect 16310 1730 16340 1735
rect 17380 1875 17410 1905
rect 17765 1865 17795 1895
rect 16645 1820 16675 1850
rect 17235 1820 17265 1850
rect 17455 1820 17485 1850
rect 17685 1820 17715 1850
rect 16825 1775 16855 1805
rect 16945 1775 16975 1805
rect 16530 1755 16560 1760
rect 16530 1735 16535 1755
rect 16535 1735 16555 1755
rect 16555 1735 16560 1755
rect 16530 1730 16560 1735
rect 17130 1755 17160 1760
rect 17130 1735 17135 1755
rect 17135 1735 17155 1755
rect 17155 1735 17160 1755
rect 17130 1730 17160 1735
rect 17350 1755 17380 1760
rect 17350 1735 17355 1755
rect 17355 1735 17375 1755
rect 17375 1735 17380 1755
rect 17350 1730 17380 1735
rect 17570 1755 17600 1760
rect 17570 1735 17575 1755
rect 17575 1735 17595 1755
rect 17595 1735 17600 1755
rect 17570 1730 17600 1735
rect 16240 1710 16266 1715
rect 16240 1690 16243 1710
rect 16243 1690 16260 1710
rect 16260 1690 16266 1710
rect 16240 1685 16266 1690
rect 16460 1710 16486 1715
rect 16460 1690 16463 1710
rect 16463 1690 16480 1710
rect 16480 1690 16486 1710
rect 16460 1685 16486 1690
rect 16604 1710 16630 1715
rect 16604 1690 16610 1710
rect 16610 1690 16627 1710
rect 16627 1690 16630 1710
rect 16604 1685 16630 1690
rect 16870 1710 16896 1715
rect 16870 1690 16876 1710
rect 16876 1690 16893 1710
rect 16893 1690 16896 1710
rect 16870 1685 16896 1690
rect 17280 1710 17306 1715
rect 17280 1690 17283 1710
rect 17283 1690 17300 1710
rect 17300 1690 17306 1710
rect 17280 1685 17306 1690
rect 17500 1710 17526 1715
rect 17500 1690 17503 1710
rect 17503 1690 17520 1710
rect 17520 1690 17526 1710
rect 17500 1685 17526 1690
rect 17644 1710 17670 1715
rect 17644 1690 17650 1710
rect 17650 1690 17667 1710
rect 17667 1690 17670 1710
rect 17644 1685 17670 1690
rect 16109 1490 16135 1495
rect 16109 1470 16112 1490
rect 16112 1470 16129 1490
rect 16129 1470 16135 1490
rect 16109 1465 16135 1470
rect 16310 1490 16340 1495
rect 16310 1470 16315 1490
rect 16315 1470 16335 1490
rect 16335 1470 16340 1490
rect 16310 1465 16340 1470
rect 16530 1490 16560 1495
rect 16530 1470 16535 1490
rect 16535 1470 16555 1490
rect 16555 1470 16560 1490
rect 16530 1465 16560 1470
rect 16925 1490 16951 1495
rect 16925 1470 16928 1490
rect 16928 1470 16945 1490
rect 16945 1470 16951 1490
rect 16925 1465 16951 1470
rect 17149 1490 17175 1495
rect 17149 1470 17152 1490
rect 17152 1470 17169 1490
rect 17169 1470 17175 1490
rect 17149 1465 17175 1470
rect 17350 1490 17380 1495
rect 17350 1470 17355 1490
rect 17355 1470 17375 1490
rect 17375 1470 17380 1490
rect 17350 1465 17380 1470
rect 17570 1490 17600 1495
rect 17570 1470 17575 1490
rect 17575 1470 17595 1490
rect 17595 1470 17600 1490
rect 17570 1465 17600 1470
rect 16150 1430 16180 1435
rect 16150 1410 16155 1430
rect 16155 1410 16175 1430
rect 16175 1410 16180 1430
rect 16150 1405 16180 1410
rect 16255 1430 16285 1435
rect 16255 1410 16260 1430
rect 16260 1410 16280 1430
rect 16280 1410 16285 1430
rect 16255 1405 16285 1410
rect 16365 1430 16395 1435
rect 16365 1410 16370 1430
rect 16370 1410 16390 1430
rect 16390 1410 16395 1430
rect 16365 1405 16395 1410
rect 16475 1430 16505 1435
rect 16475 1410 16480 1430
rect 16480 1410 16500 1430
rect 16500 1410 16505 1430
rect 16475 1405 16505 1410
rect 16585 1430 16615 1435
rect 16585 1410 16590 1430
rect 16590 1410 16610 1430
rect 16610 1410 16615 1430
rect 16585 1405 16615 1410
rect 16010 1315 16040 1345
rect 16815 1315 16845 1345
rect 16320 1265 16350 1295
rect 17190 1430 17220 1435
rect 17190 1410 17195 1430
rect 17195 1410 17215 1430
rect 17215 1410 17220 1430
rect 17190 1405 17220 1410
rect 17295 1430 17325 1435
rect 17295 1410 17300 1430
rect 17300 1410 17320 1430
rect 17320 1410 17325 1430
rect 17295 1405 17325 1410
rect 17405 1430 17435 1435
rect 17405 1410 17410 1430
rect 17410 1410 17430 1430
rect 17430 1410 17435 1430
rect 17405 1405 17435 1410
rect 17515 1430 17545 1435
rect 17515 1410 17520 1430
rect 17520 1410 17540 1430
rect 17540 1410 17545 1430
rect 17515 1405 17545 1410
rect 17625 1430 17655 1435
rect 17625 1410 17630 1430
rect 17630 1410 17650 1430
rect 17650 1410 17655 1430
rect 17625 1405 17655 1410
rect 16885 1265 16915 1295
rect 16430 1230 16460 1235
rect 16430 1210 16435 1230
rect 16435 1210 16455 1230
rect 16455 1210 16460 1230
rect 16430 1205 16460 1210
rect 16540 1230 16570 1235
rect 16540 1210 16545 1230
rect 16545 1210 16565 1230
rect 16565 1210 16570 1230
rect 16540 1205 16570 1210
rect 16650 1230 16680 1235
rect 16650 1210 16655 1230
rect 16655 1210 16675 1230
rect 16675 1210 16680 1230
rect 16650 1205 16680 1210
rect 16760 1230 16790 1235
rect 16760 1210 16765 1230
rect 16765 1210 16785 1230
rect 16785 1210 16790 1230
rect 16760 1205 16790 1210
rect 16870 1230 16900 1235
rect 16870 1210 16875 1230
rect 16875 1210 16895 1230
rect 16895 1210 16900 1230
rect 16870 1205 16900 1210
rect 16980 1230 17010 1235
rect 16980 1210 16985 1230
rect 16985 1210 17005 1230
rect 17005 1210 17010 1230
rect 16980 1205 17010 1210
rect 17090 1230 17120 1235
rect 17090 1210 17095 1230
rect 17095 1210 17115 1230
rect 17115 1210 17120 1230
rect 17090 1205 17120 1210
rect 17200 1230 17230 1235
rect 17200 1210 17205 1230
rect 17205 1210 17225 1230
rect 17225 1210 17230 1230
rect 17200 1205 17230 1210
rect 17310 1230 17340 1235
rect 17310 1210 17315 1230
rect 17315 1210 17335 1230
rect 17335 1210 17340 1230
rect 17310 1205 17340 1210
rect 17420 1230 17450 1235
rect 17420 1210 17425 1230
rect 17425 1210 17445 1230
rect 17445 1210 17450 1230
rect 17420 1205 17450 1210
rect 17530 1230 17560 1235
rect 17530 1210 17535 1230
rect 17535 1210 17555 1230
rect 17555 1210 17560 1230
rect 17530 1205 17560 1210
rect 17600 1245 17630 1250
rect 17600 1225 17605 1245
rect 17605 1225 17625 1245
rect 17625 1225 17630 1245
rect 17600 1220 17630 1225
rect 17810 1220 17840 1250
rect 16170 910 16200 915
rect 16170 890 16175 910
rect 16175 890 16195 910
rect 16195 890 16200 910
rect 16170 885 16200 890
rect 16265 910 16295 915
rect 16265 890 16270 910
rect 16270 890 16290 910
rect 16290 890 16295 910
rect 16265 885 16295 890
rect 16375 910 16405 915
rect 16375 890 16380 910
rect 16380 890 16400 910
rect 16400 890 16405 910
rect 16375 885 16405 890
rect 16485 910 16515 915
rect 16485 890 16490 910
rect 16490 890 16510 910
rect 16510 890 16515 910
rect 16485 885 16515 890
rect 16595 910 16625 915
rect 16595 890 16600 910
rect 16600 890 16620 910
rect 16620 890 16625 910
rect 16595 885 16625 890
rect 16705 910 16735 915
rect 16705 890 16710 910
rect 16710 890 16730 910
rect 16730 890 16735 910
rect 16705 885 16735 890
rect 16815 910 16845 915
rect 16815 890 16820 910
rect 16820 890 16840 910
rect 16840 890 16845 910
rect 16815 885 16845 890
rect 16925 910 16955 915
rect 16925 890 16930 910
rect 16930 890 16950 910
rect 16950 890 16955 910
rect 16925 885 16955 890
rect 17035 910 17065 915
rect 17035 890 17040 910
rect 17040 890 17060 910
rect 17060 890 17065 910
rect 17035 885 17065 890
rect 17145 910 17175 915
rect 17145 890 17150 910
rect 17150 890 17170 910
rect 17170 890 17175 910
rect 17145 885 17175 890
rect 17255 910 17285 915
rect 17255 890 17260 910
rect 17260 890 17280 910
rect 17280 890 17285 910
rect 17255 885 17285 890
rect 17365 910 17395 915
rect 17365 890 17370 910
rect 17370 890 17390 910
rect 17390 890 17395 910
rect 17365 885 17395 890
rect 17475 910 17505 915
rect 17475 890 17480 910
rect 17480 890 17500 910
rect 17500 890 17505 910
rect 17475 885 17505 890
rect 17625 910 17655 915
rect 17625 890 17630 910
rect 17630 890 17650 910
rect 17650 890 17655 910
rect 17625 885 17655 890
rect 16010 825 16040 855
rect 16500 825 16530 855
rect 16940 830 16970 860
rect 17160 830 17190 860
rect 17380 830 17410 860
rect 18005 3630 18035 3635
rect 18005 3610 18010 3630
rect 18010 3610 18030 3630
rect 18030 3610 18035 3630
rect 18005 3605 18035 3610
rect 18115 3630 18145 3635
rect 18115 3610 18120 3630
rect 18120 3610 18140 3630
rect 18140 3610 18145 3630
rect 18115 3605 18145 3610
rect 18225 3630 18255 3635
rect 18225 3610 18230 3630
rect 18230 3610 18250 3630
rect 18250 3610 18255 3630
rect 18225 3605 18255 3610
rect 18335 3630 18365 3635
rect 18335 3610 18340 3630
rect 18340 3610 18360 3630
rect 18360 3610 18365 3630
rect 18335 3605 18365 3610
rect 18445 3630 18475 3635
rect 18445 3610 18450 3630
rect 18450 3610 18470 3630
rect 18470 3610 18475 3630
rect 18445 3605 18475 3610
rect 18555 3630 18585 3635
rect 18555 3610 18560 3630
rect 18560 3610 18580 3630
rect 18580 3610 18585 3630
rect 18555 3605 18585 3610
rect 18810 3605 18840 3635
rect 18760 3525 18790 3555
rect 18810 3525 18840 3555
rect 18860 3525 18890 3555
rect 18060 2960 18090 2965
rect 18060 2940 18065 2960
rect 18065 2940 18085 2960
rect 18085 2940 18090 2960
rect 18060 2935 18090 2940
rect 18170 2960 18200 2965
rect 18170 2940 18175 2960
rect 18175 2940 18195 2960
rect 18195 2940 18200 2960
rect 18170 2935 18200 2940
rect 18280 2960 18310 2965
rect 18280 2940 18285 2960
rect 18285 2940 18305 2960
rect 18305 2940 18310 2960
rect 18280 2935 18310 2940
rect 18390 2960 18420 2965
rect 18390 2940 18395 2960
rect 18395 2940 18415 2960
rect 18415 2940 18420 2960
rect 18390 2935 18420 2940
rect 18500 2960 18530 2965
rect 18500 2940 18505 2960
rect 18505 2940 18525 2960
rect 18525 2940 18530 2960
rect 18500 2935 18530 2940
rect 18115 2850 18145 2880
rect 18760 2905 18790 2935
rect 18810 2905 18840 2935
rect 18860 2905 18890 2935
rect 18810 2850 18840 2880
rect 18390 2795 18420 2825
rect 19250 2795 19280 2825
rect 18005 2700 18035 2705
rect 18005 2680 18010 2700
rect 18010 2680 18030 2700
rect 18030 2680 18035 2700
rect 18005 2675 18035 2680
rect 18115 2700 18145 2705
rect 18115 2680 18120 2700
rect 18120 2680 18140 2700
rect 18140 2680 18145 2700
rect 18115 2675 18145 2680
rect 18225 2700 18255 2705
rect 18225 2680 18230 2700
rect 18230 2680 18250 2700
rect 18250 2680 18255 2700
rect 18225 2675 18255 2680
rect 18335 2700 18365 2705
rect 18335 2680 18340 2700
rect 18340 2680 18360 2700
rect 18360 2680 18365 2700
rect 18335 2675 18365 2680
rect 18445 2700 18475 2705
rect 18445 2680 18450 2700
rect 18450 2680 18470 2700
rect 18470 2680 18475 2700
rect 18445 2675 18475 2680
rect 18555 2700 18585 2705
rect 18555 2680 18560 2700
rect 18560 2680 18580 2700
rect 18580 2680 18585 2700
rect 18555 2675 18585 2680
rect 18060 2430 18090 2435
rect 18060 2410 18065 2430
rect 18065 2410 18085 2430
rect 18085 2410 18090 2430
rect 18060 2405 18090 2410
rect 18170 2430 18200 2435
rect 18170 2410 18175 2430
rect 18175 2410 18195 2430
rect 18195 2410 18200 2430
rect 18170 2405 18200 2410
rect 18280 2430 18310 2435
rect 18280 2410 18285 2430
rect 18285 2410 18305 2430
rect 18305 2410 18310 2430
rect 18280 2405 18310 2410
rect 18390 2430 18420 2435
rect 18390 2410 18395 2430
rect 18395 2410 18415 2430
rect 18415 2410 18420 2430
rect 18390 2405 18420 2410
rect 18500 2430 18530 2435
rect 18500 2410 18505 2430
rect 18505 2410 18525 2430
rect 18525 2410 18530 2430
rect 18500 2405 18530 2410
rect 18745 2405 18775 2435
rect 18030 2370 18060 2375
rect 18030 2350 18035 2370
rect 18035 2350 18055 2370
rect 18055 2350 18060 2370
rect 18030 2345 18060 2350
rect 18060 2310 18090 2315
rect 18060 2290 18065 2310
rect 18065 2290 18085 2310
rect 18085 2290 18090 2310
rect 18060 2285 18090 2290
rect 18170 2310 18200 2315
rect 18170 2290 18175 2310
rect 18175 2290 18195 2310
rect 18195 2290 18200 2310
rect 18170 2285 18200 2290
rect 18280 2310 18310 2315
rect 18280 2290 18285 2310
rect 18285 2290 18305 2310
rect 18305 2290 18310 2310
rect 18280 2285 18310 2290
rect 18390 2310 18420 2315
rect 18390 2290 18395 2310
rect 18395 2290 18415 2310
rect 18415 2290 18420 2310
rect 18390 2285 18420 2290
rect 18500 2310 18530 2315
rect 18500 2290 18505 2310
rect 18505 2290 18525 2310
rect 18525 2290 18530 2310
rect 18500 2285 18530 2290
rect 18700 2285 18730 2315
rect 19250 2080 19280 2110
rect 18745 1970 18775 2000
rect 18795 2000 18830 2005
rect 18795 1975 18800 2000
rect 18800 1975 18825 2000
rect 18825 1975 18830 2000
rect 18795 1970 18830 1975
rect 18855 2000 18890 2005
rect 18855 1975 18860 2000
rect 18860 1975 18885 2000
rect 18885 1975 18890 2000
rect 18855 1970 18890 1975
rect 18915 2000 18950 2005
rect 18915 1975 18920 2000
rect 18920 1975 18945 2000
rect 18945 1975 18950 2000
rect 18915 1970 18950 1975
rect 18975 2000 19010 2005
rect 18975 1975 18980 2000
rect 18980 1975 19005 2000
rect 19005 1975 19010 2000
rect 18975 1970 19010 1975
rect 18005 1940 18035 1945
rect 18005 1920 18012 1940
rect 18012 1920 18030 1940
rect 18030 1920 18035 1940
rect 18005 1915 18035 1920
rect 18115 1940 18145 1945
rect 18115 1920 18122 1940
rect 18122 1920 18140 1940
rect 18140 1920 18145 1940
rect 18115 1915 18145 1920
rect 18225 1940 18255 1945
rect 18225 1920 18232 1940
rect 18232 1920 18250 1940
rect 18250 1920 18255 1940
rect 18225 1915 18255 1920
rect 18335 1940 18365 1945
rect 18335 1920 18342 1940
rect 18342 1920 18360 1940
rect 18360 1920 18365 1940
rect 18335 1915 18365 1920
rect 18445 1940 18475 1945
rect 18445 1920 18452 1940
rect 18452 1920 18470 1940
rect 18470 1920 18475 1940
rect 18445 1915 18475 1920
rect 18555 1940 18585 1945
rect 18555 1920 18562 1940
rect 18562 1920 18580 1940
rect 18580 1920 18585 1940
rect 18555 1915 18585 1920
rect 18700 1915 18730 1945
rect 18855 1915 18885 1945
rect 18975 1865 19005 1895
rect 17930 1730 17960 1760
rect 18210 1730 18240 1760
rect 18800 1730 18830 1760
rect 18110 1700 18140 1705
rect 18110 1680 18115 1700
rect 18115 1680 18135 1700
rect 18135 1680 18140 1700
rect 18110 1675 18140 1680
rect 18310 1700 18340 1705
rect 18310 1680 18315 1700
rect 18315 1680 18335 1700
rect 18335 1680 18340 1700
rect 18310 1675 18340 1680
rect 18510 1700 18540 1705
rect 18510 1680 18515 1700
rect 18515 1680 18535 1700
rect 18535 1680 18540 1700
rect 18510 1675 18540 1680
rect 18735 1675 18765 1705
rect 19250 1675 19280 1705
rect 18735 1640 18770 1645
rect 18735 1615 18740 1640
rect 18740 1615 18765 1640
rect 18765 1615 18770 1640
rect 18735 1610 18770 1615
rect 18795 1640 18830 1645
rect 18795 1615 18800 1640
rect 18800 1615 18825 1640
rect 18825 1615 18830 1640
rect 18795 1610 18830 1615
rect 17930 1360 17960 1390
rect 18210 930 18240 935
rect 18210 910 18215 930
rect 18215 910 18235 930
rect 18235 910 18240 930
rect 18210 905 18240 910
rect 18410 930 18440 935
rect 18410 910 18415 930
rect 18415 910 18435 930
rect 18435 910 18440 930
rect 18410 905 18440 910
rect 17865 830 17895 860
rect 15955 765 15985 795
rect 2525 730 2555 760
rect 3135 755 3165 760
rect 3135 735 3140 755
rect 3140 735 3160 755
rect 3160 735 3165 755
rect 3135 730 3165 735
rect 3630 755 3660 760
rect 3630 735 3635 755
rect 3635 735 3655 755
rect 3655 735 3660 755
rect 3630 730 3660 735
rect 3990 755 4020 760
rect 3990 735 3995 755
rect 3995 735 4015 755
rect 4015 735 4020 755
rect 3990 730 4020 735
rect 4350 755 4380 760
rect 4350 735 4355 755
rect 4355 735 4375 755
rect 4375 735 4380 755
rect 4350 730 4380 735
rect 4530 755 4560 760
rect 4530 735 4535 755
rect 4535 735 4555 755
rect 4555 735 4560 755
rect 4530 730 4560 735
rect 4710 755 4740 760
rect 4710 735 4715 755
rect 4715 735 4735 755
rect 4735 735 4740 755
rect 4710 730 4740 735
rect 16310 790 16340 795
rect 16310 770 16315 790
rect 16315 770 16335 790
rect 16335 770 16340 790
rect 16310 765 16340 770
rect 16380 790 16410 795
rect 16380 770 16385 790
rect 16385 770 16405 790
rect 16405 770 16410 790
rect 16380 765 16410 770
rect 16450 790 16480 795
rect 16450 770 16455 790
rect 16455 770 16475 790
rect 16475 770 16480 790
rect 16450 765 16480 770
rect 17050 795 17080 800
rect 17050 775 17055 795
rect 17055 775 17075 795
rect 17075 775 17080 795
rect 17050 770 17080 775
rect 17270 795 17300 800
rect 17270 775 17275 795
rect 17275 775 17295 795
rect 17295 775 17300 795
rect 17270 770 17300 775
rect 17490 795 17520 800
rect 17490 775 17495 795
rect 17495 775 17515 795
rect 17515 775 17520 795
rect 17490 770 17520 775
rect 17810 770 17840 800
rect 4890 755 4920 760
rect 4890 735 4895 755
rect 4895 735 4915 755
rect 4915 735 4920 755
rect 4890 730 4920 735
rect 3450 675 3480 705
rect 3810 675 3840 705
rect 4170 675 4200 705
rect 16995 675 17025 680
rect 16995 655 17000 675
rect 17000 655 17020 675
rect 17020 655 17025 675
rect 16995 650 17025 655
rect 17105 675 17135 680
rect 17105 655 17110 675
rect 17110 655 17130 675
rect 17130 655 17135 675
rect 17105 650 17135 655
rect 17215 675 17245 680
rect 17215 655 17220 675
rect 17220 655 17240 675
rect 17240 655 17245 675
rect 17215 650 17245 655
rect 17325 675 17355 680
rect 17325 655 17330 675
rect 17330 655 17350 675
rect 17350 655 17355 675
rect 17325 650 17355 655
rect 17435 675 17465 680
rect 17435 655 17440 675
rect 17440 655 17460 675
rect 17460 655 17465 675
rect 17435 650 17465 655
<< metal2 >>
rect -195 4990 -155 4995
rect -195 4960 -190 4990
rect -160 4960 -155 4990
rect -195 4955 -155 4960
rect 5550 4990 5590 4995
rect 5550 4960 5555 4990
rect 5585 4960 5590 4990
rect 5550 4955 5590 4960
rect 16632 4515 16668 4520
rect 16632 4485 16635 4515
rect 16665 4510 16668 4515
rect 16752 4515 16788 4520
rect 16752 4510 16755 4515
rect 16665 4490 16755 4510
rect 16665 4485 16668 4490
rect 16632 4480 16668 4485
rect 16752 4485 16755 4490
rect 16785 4510 16788 4515
rect 16872 4515 16908 4520
rect 16872 4510 16875 4515
rect 16785 4490 16875 4510
rect 16785 4485 16788 4490
rect 16752 4480 16788 4485
rect 16872 4485 16875 4490
rect 16905 4510 16908 4515
rect 17080 4515 17120 4520
rect 17080 4510 17085 4515
rect 16905 4490 17085 4510
rect 16905 4485 16908 4490
rect 16872 4480 16908 4485
rect 17080 4485 17085 4490
rect 17115 4485 17120 4515
rect 17080 4480 17120 4485
rect 16570 4470 16610 4475
rect 16570 4460 16575 4470
rect 16200 4455 16240 4460
rect 16200 4425 16205 4455
rect 16235 4425 16240 4455
rect 16200 4420 16240 4425
rect 16460 4455 16575 4460
rect 16460 4425 16465 4455
rect 16495 4440 16575 4455
rect 16605 4465 16610 4470
rect 16690 4470 16730 4475
rect 16690 4465 16695 4470
rect 16605 4445 16695 4465
rect 16605 4440 16610 4445
rect 16495 4425 16500 4440
rect 16570 4435 16610 4440
rect 16690 4440 16695 4445
rect 16725 4465 16730 4470
rect 16810 4470 16850 4475
rect 16810 4465 16815 4470
rect 16725 4445 16815 4465
rect 16725 4440 16730 4445
rect 16690 4435 16730 4440
rect 16810 4440 16815 4445
rect 16845 4465 16850 4470
rect 16930 4470 16970 4475
rect 16930 4465 16935 4470
rect 16845 4445 16935 4465
rect 16845 4440 16850 4445
rect 16810 4435 16850 4440
rect 16930 4440 16935 4445
rect 16965 4440 16970 4470
rect 16930 4435 16970 4440
rect 17080 4445 17120 4450
rect 16460 4420 16500 4425
rect 17080 4415 17085 4445
rect 17115 4440 17120 4445
rect 17200 4445 17240 4450
rect 17200 4440 17205 4445
rect 17115 4420 17205 4440
rect 17115 4415 17120 4420
rect 17080 4410 17120 4415
rect 17200 4415 17205 4420
rect 17235 4440 17240 4445
rect 17320 4445 17360 4450
rect 17320 4440 17325 4445
rect 17235 4420 17325 4440
rect 17235 4415 17240 4420
rect 17200 4410 17240 4415
rect 17320 4415 17325 4420
rect 17355 4440 17360 4445
rect 17440 4445 17480 4450
rect 17440 4440 17445 4445
rect 17355 4420 17445 4440
rect 17355 4415 17360 4420
rect 17320 4410 17360 4415
rect 17440 4415 17445 4420
rect 17475 4440 17480 4445
rect 17560 4445 17600 4450
rect 17560 4440 17565 4445
rect 17475 4420 17565 4440
rect 17475 4415 17480 4420
rect 17440 4410 17480 4415
rect 17560 4415 17565 4420
rect 17595 4415 17600 4445
rect 17560 4410 17600 4415
rect 16330 4320 16370 4325
rect 16050 4315 16090 4320
rect 16050 4285 16055 4315
rect 16085 4310 16090 4315
rect 16330 4310 16335 4320
rect 16085 4290 16335 4310
rect 16365 4310 16370 4320
rect 16750 4315 16790 4320
rect 16750 4310 16755 4315
rect 16365 4290 16755 4310
rect 16085 4285 16090 4290
rect 16330 4285 16370 4290
rect 16750 4285 16755 4290
rect 16785 4310 16790 4315
rect 17140 4315 17180 4320
rect 17140 4310 17145 4315
rect 16785 4290 17145 4310
rect 16785 4285 16790 4290
rect 16050 4280 16090 4285
rect 16750 4280 16790 4285
rect 17140 4285 17145 4290
rect 17175 4310 17180 4315
rect 17260 4315 17300 4320
rect 17260 4310 17265 4315
rect 17175 4290 17265 4310
rect 17175 4285 17180 4290
rect 17140 4280 17180 4285
rect 17260 4285 17265 4290
rect 17295 4310 17300 4315
rect 17380 4315 17420 4320
rect 17380 4310 17385 4315
rect 17295 4290 17385 4310
rect 17295 4285 17300 4290
rect 17260 4280 17300 4285
rect 17380 4285 17385 4290
rect 17415 4310 17420 4315
rect 17500 4315 17540 4320
rect 17500 4310 17505 4315
rect 17415 4290 17505 4310
rect 17415 4285 17420 4290
rect 17380 4280 17420 4285
rect 17500 4285 17505 4290
rect 17535 4285 17540 4315
rect 17500 4280 17540 4285
rect 16105 4260 16145 4265
rect 16105 4230 16110 4260
rect 16140 4255 16145 4260
rect 16330 4260 16370 4265
rect 16330 4255 16335 4260
rect 16140 4235 16335 4255
rect 16140 4230 16145 4235
rect 16105 4225 16145 4230
rect 16330 4230 16335 4235
rect 16365 4255 16370 4260
rect 17200 4260 17240 4265
rect 17200 4255 17205 4260
rect 16365 4235 17205 4255
rect 16365 4230 16370 4235
rect 16330 4225 16370 4230
rect 17200 4230 17205 4235
rect 17235 4230 17240 4260
rect 17200 4225 17240 4230
rect 16360 4205 16400 4210
rect 16360 4175 16365 4205
rect 16395 4200 16400 4205
rect 16470 4205 16510 4210
rect 16470 4200 16475 4205
rect 16395 4180 16475 4200
rect 16395 4175 16400 4180
rect 16360 4170 16400 4175
rect 16470 4175 16475 4180
rect 16505 4200 16510 4205
rect 16580 4205 16620 4210
rect 16580 4200 16585 4205
rect 16505 4180 16585 4200
rect 16505 4175 16510 4180
rect 16470 4170 16510 4175
rect 16580 4175 16585 4180
rect 16615 4200 16620 4205
rect 16690 4205 16730 4210
rect 16690 4200 16695 4205
rect 16615 4180 16695 4200
rect 16615 4175 16620 4180
rect 16580 4170 16620 4175
rect 16690 4175 16695 4180
rect 16725 4200 16730 4205
rect 16800 4205 16840 4210
rect 16800 4200 16805 4205
rect 16725 4180 16805 4200
rect 16725 4175 16730 4180
rect 16690 4170 16730 4175
rect 16800 4175 16805 4180
rect 16835 4200 16840 4205
rect 16910 4205 16950 4210
rect 16910 4200 16915 4205
rect 16835 4180 16915 4200
rect 16835 4175 16840 4180
rect 16800 4170 16840 4175
rect 16910 4175 16915 4180
rect 16945 4200 16950 4205
rect 17020 4205 17060 4210
rect 17020 4200 17025 4205
rect 16945 4180 17025 4200
rect 16945 4175 16950 4180
rect 16910 4170 16950 4175
rect 17020 4175 17025 4180
rect 17055 4200 17060 4205
rect 17130 4205 17170 4210
rect 17130 4200 17135 4205
rect 17055 4180 17135 4200
rect 17055 4175 17060 4180
rect 17020 4170 17060 4175
rect 17130 4175 17135 4180
rect 17165 4200 17170 4205
rect 17240 4205 17280 4210
rect 17240 4200 17245 4205
rect 17165 4180 17245 4200
rect 17165 4175 17170 4180
rect 17130 4170 17170 4175
rect 17240 4175 17245 4180
rect 17275 4200 17280 4205
rect 17350 4205 17390 4210
rect 17350 4200 17355 4205
rect 17275 4180 17355 4200
rect 17275 4175 17280 4180
rect 17240 4170 17280 4175
rect 17350 4175 17355 4180
rect 17385 4175 17390 4205
rect 17350 4170 17390 4175
rect 16305 4085 16345 4090
rect 16305 4055 16310 4085
rect 16340 4080 16345 4085
rect 16525 4085 16565 4090
rect 16525 4080 16530 4085
rect 16340 4060 16530 4080
rect 16340 4055 16345 4060
rect 16305 4050 16345 4055
rect 16525 4055 16530 4060
rect 16560 4080 16565 4085
rect 16745 4085 16785 4090
rect 16745 4080 16750 4085
rect 16560 4060 16750 4080
rect 16560 4055 16565 4060
rect 16525 4050 16565 4055
rect 16745 4055 16750 4060
rect 16780 4080 16785 4085
rect 16965 4085 17005 4090
rect 16965 4080 16970 4085
rect 16780 4060 16970 4080
rect 16780 4055 16785 4060
rect 16745 4050 16785 4055
rect 16965 4055 16970 4060
rect 17000 4080 17005 4085
rect 17185 4085 17225 4090
rect 17185 4080 17190 4085
rect 17000 4060 17190 4080
rect 17000 4055 17005 4060
rect 16965 4050 17005 4055
rect 17185 4055 17190 4060
rect 17220 4080 17225 4085
rect 17405 4085 17445 4090
rect 17405 4080 17410 4085
rect 17220 4060 17410 4080
rect 17220 4055 17225 4060
rect 17185 4050 17225 4055
rect 17405 4055 17410 4060
rect 17440 4055 17445 4085
rect 17405 4050 17445 4055
rect 16415 4025 16455 4030
rect 16415 3995 16420 4025
rect 16450 4020 16455 4025
rect 16635 4025 16675 4030
rect 16635 4020 16640 4025
rect 16450 4000 16640 4020
rect 16450 3995 16455 4000
rect 16415 3990 16455 3995
rect 16635 3995 16640 4000
rect 16670 4020 16675 4025
rect 16855 4025 16895 4030
rect 16855 4020 16860 4025
rect 16670 4000 16860 4020
rect 16670 3995 16675 4000
rect 16635 3990 16675 3995
rect 16855 3995 16860 4000
rect 16890 4020 16895 4025
rect 17075 4025 17115 4030
rect 17075 4020 17080 4025
rect 16890 4000 17080 4020
rect 16890 3995 16895 4000
rect 16855 3990 16895 3995
rect 17075 3995 17080 4000
rect 17110 4020 17115 4025
rect 17295 4025 17335 4030
rect 17295 4020 17300 4025
rect 17110 4000 17300 4020
rect 17110 3995 17115 4000
rect 17075 3990 17115 3995
rect 17295 3995 17300 4000
rect 17330 3995 17335 4025
rect 17295 3990 17335 3995
rect 16310 3960 16350 3965
rect 16310 3930 16315 3960
rect 16345 3955 16350 3960
rect 16415 3960 16455 3965
rect 16415 3955 16420 3960
rect 16345 3935 16420 3955
rect 16345 3930 16350 3935
rect 16310 3925 16350 3930
rect 16415 3930 16420 3935
rect 16450 3955 16455 3960
rect 16525 3960 16565 3965
rect 16525 3955 16530 3960
rect 16450 3935 16530 3955
rect 16450 3930 16455 3935
rect 16415 3925 16455 3930
rect 16525 3930 16530 3935
rect 16560 3955 16565 3960
rect 16635 3960 16675 3965
rect 16635 3955 16640 3960
rect 16560 3935 16640 3955
rect 16560 3930 16565 3935
rect 16525 3925 16565 3930
rect 16635 3930 16640 3935
rect 16670 3955 16675 3960
rect 16745 3960 16785 3965
rect 16745 3955 16750 3960
rect 16670 3935 16750 3955
rect 16670 3930 16675 3935
rect 16635 3925 16675 3930
rect 16745 3930 16750 3935
rect 16780 3930 16785 3960
rect 16745 3925 16785 3930
rect 17050 3960 17090 3965
rect 17050 3930 17055 3960
rect 17085 3955 17090 3960
rect 17155 3960 17195 3965
rect 17155 3955 17160 3960
rect 17085 3935 17160 3955
rect 17085 3930 17090 3935
rect 17050 3925 17090 3930
rect 17155 3930 17160 3935
rect 17190 3955 17195 3960
rect 17265 3960 17305 3965
rect 17265 3955 17270 3960
rect 17190 3935 17270 3955
rect 17190 3930 17195 3935
rect 17155 3925 17195 3930
rect 17265 3930 17270 3935
rect 17300 3955 17305 3960
rect 17375 3960 17415 3965
rect 17375 3955 17380 3960
rect 17300 3935 17380 3955
rect 17300 3930 17305 3935
rect 17265 3925 17305 3930
rect 17375 3930 17380 3935
rect 17410 3955 17415 3960
rect 17485 3960 17525 3965
rect 17485 3955 17490 3960
rect 17410 3935 17490 3955
rect 17410 3930 17415 3935
rect 17375 3925 17415 3930
rect 17485 3930 17490 3935
rect 17520 3930 17525 3960
rect 17485 3925 17525 3930
rect 16271 3900 16303 3905
rect 16271 3870 16274 3900
rect 16300 3895 16303 3900
rect 16470 3900 16510 3905
rect 16470 3895 16475 3900
rect 16300 3875 16475 3895
rect 16300 3870 16303 3875
rect 16271 3865 16303 3870
rect 16470 3870 16475 3875
rect 16505 3895 16510 3900
rect 16690 3900 16730 3905
rect 16690 3895 16695 3900
rect 16505 3875 16695 3895
rect 16505 3870 16510 3875
rect 16470 3865 16510 3870
rect 16690 3870 16695 3875
rect 16725 3895 16730 3900
rect 17011 3900 17043 3905
rect 17011 3895 17014 3900
rect 16725 3875 17014 3895
rect 16725 3870 16730 3875
rect 16690 3865 16730 3870
rect 17011 3870 17014 3875
rect 17040 3895 17043 3900
rect 17210 3900 17250 3905
rect 17210 3895 17215 3900
rect 17040 3875 17215 3895
rect 17040 3870 17043 3875
rect 17011 3865 17043 3870
rect 17210 3870 17215 3875
rect 17245 3895 17250 3900
rect 17430 3900 17470 3905
rect 17430 3895 17435 3900
rect 17245 3875 17435 3895
rect 17245 3870 17250 3875
rect 17210 3865 17250 3870
rect 17430 3870 17435 3875
rect 17465 3895 17470 3900
rect 17760 3900 17800 3905
rect 17760 3895 17765 3900
rect 17465 3875 17765 3895
rect 17465 3870 17470 3875
rect 17430 3865 17470 3870
rect 17760 3870 17765 3875
rect 17795 3870 17800 3900
rect 17760 3865 17800 3870
rect 16402 3780 16434 3785
rect 16402 3775 16405 3780
rect 15915 3755 16405 3775
rect 16402 3750 16405 3755
rect 16431 3775 16434 3780
rect 16622 3780 16654 3785
rect 16622 3775 16625 3780
rect 16431 3755 16625 3775
rect 16431 3750 16434 3755
rect 16402 3745 16434 3750
rect 16622 3750 16625 3755
rect 16651 3775 16654 3780
rect 16766 3780 16798 3785
rect 16766 3775 16769 3780
rect 16651 3755 16769 3775
rect 16651 3750 16654 3755
rect 16622 3745 16654 3750
rect 16766 3750 16769 3755
rect 16795 3775 16798 3780
rect 17142 3780 17174 3785
rect 17142 3775 17145 3780
rect 16795 3755 17145 3775
rect 16795 3750 16798 3755
rect 16766 3745 16798 3750
rect 17142 3750 17145 3755
rect 17171 3775 17174 3780
rect 17362 3780 17394 3785
rect 17362 3775 17365 3780
rect 17171 3755 17365 3775
rect 17171 3750 17174 3755
rect 17142 3745 17174 3750
rect 17362 3750 17365 3755
rect 17391 3775 17394 3780
rect 17506 3780 17538 3785
rect 17506 3775 17509 3780
rect 17391 3755 17509 3775
rect 17391 3750 17394 3755
rect 17362 3745 17394 3750
rect 17506 3750 17509 3755
rect 17535 3750 17538 3780
rect 17506 3745 17538 3750
rect 16990 3730 17030 3735
rect 16250 3720 16290 3725
rect 16250 3690 16255 3720
rect 16285 3715 16290 3720
rect 16355 3720 16395 3725
rect 16355 3715 16360 3720
rect 16285 3695 16360 3715
rect 16285 3690 16290 3695
rect 16250 3685 16290 3690
rect 16355 3690 16360 3695
rect 16390 3715 16395 3720
rect 16470 3720 16510 3725
rect 16470 3715 16475 3720
rect 16390 3695 16475 3715
rect 16390 3690 16395 3695
rect 16355 3685 16395 3690
rect 16470 3690 16475 3695
rect 16505 3715 16510 3720
rect 16575 3720 16615 3725
rect 16575 3715 16580 3720
rect 16505 3695 16580 3715
rect 16505 3690 16510 3695
rect 16470 3685 16510 3690
rect 16575 3690 16580 3695
rect 16610 3715 16615 3720
rect 16690 3720 16730 3725
rect 16690 3715 16695 3720
rect 16610 3695 16695 3715
rect 16610 3690 16615 3695
rect 16575 3685 16615 3690
rect 16690 3690 16695 3695
rect 16725 3715 16730 3720
rect 16805 3720 16845 3725
rect 16805 3715 16810 3720
rect 16725 3695 16810 3715
rect 16725 3690 16730 3695
rect 16690 3685 16730 3690
rect 16805 3690 16810 3695
rect 16840 3690 16845 3720
rect 16990 3700 16995 3730
rect 17025 3725 17030 3730
rect 17210 3730 17250 3735
rect 17210 3725 17215 3730
rect 17025 3705 17215 3725
rect 17025 3700 17030 3705
rect 16990 3695 17030 3700
rect 17210 3700 17215 3705
rect 17245 3725 17250 3730
rect 17430 3730 17470 3735
rect 17430 3725 17435 3730
rect 17245 3705 17435 3725
rect 17245 3700 17250 3705
rect 17210 3695 17250 3700
rect 17430 3700 17435 3705
rect 17465 3725 17470 3730
rect 17860 3730 17900 3735
rect 17860 3725 17865 3730
rect 17465 3705 17865 3725
rect 17465 3700 17470 3705
rect 17430 3695 17470 3700
rect 17860 3700 17865 3705
rect 17895 3700 17900 3730
rect 17860 3695 17900 3700
rect 16805 3685 16845 3690
rect 17095 3685 17135 3690
rect 17095 3655 17100 3685
rect 17130 3680 17135 3685
rect 17315 3685 17355 3690
rect 17315 3680 17320 3685
rect 17130 3660 17320 3680
rect 17130 3655 17135 3660
rect 17095 3650 17135 3655
rect 17315 3655 17320 3660
rect 17350 3680 17355 3685
rect 17545 3685 17585 3690
rect 17545 3680 17550 3685
rect 17350 3660 17550 3680
rect 17350 3655 17355 3660
rect 17315 3650 17355 3655
rect 17545 3655 17550 3660
rect 17580 3680 17585 3685
rect 17805 3685 17845 3690
rect 17805 3680 17810 3685
rect 17580 3660 17810 3680
rect 17580 3655 17585 3660
rect 17545 3650 17585 3655
rect 17805 3655 17810 3660
rect 17840 3655 17845 3685
rect 17805 3650 17845 3655
rect 14955 3635 14995 3640
rect 14955 3605 14960 3635
rect 14990 3605 14995 3635
rect 14955 3600 14995 3605
rect 15210 3635 15250 3640
rect 15210 3605 15215 3635
rect 15245 3630 15250 3635
rect 15320 3635 15360 3640
rect 15320 3630 15325 3635
rect 15245 3610 15325 3630
rect 15245 3605 15250 3610
rect 15210 3600 15250 3605
rect 15320 3605 15325 3610
rect 15355 3630 15360 3635
rect 15430 3635 15470 3640
rect 15430 3630 15435 3635
rect 15355 3610 15435 3630
rect 15355 3605 15360 3610
rect 15320 3600 15360 3605
rect 15430 3605 15435 3610
rect 15465 3630 15470 3635
rect 15540 3635 15580 3640
rect 15540 3630 15545 3635
rect 15465 3610 15545 3630
rect 15465 3605 15470 3610
rect 15430 3600 15470 3605
rect 15540 3605 15545 3610
rect 15575 3630 15580 3635
rect 15650 3635 15690 3640
rect 15650 3630 15655 3635
rect 15575 3610 15655 3630
rect 15575 3605 15580 3610
rect 15540 3600 15580 3605
rect 15650 3605 15655 3610
rect 15685 3630 15690 3635
rect 15760 3635 15800 3640
rect 15760 3630 15765 3635
rect 15685 3610 15765 3630
rect 15685 3605 15690 3610
rect 15650 3600 15690 3605
rect 15760 3605 15765 3610
rect 15795 3605 15800 3635
rect 18000 3635 18040 3640
rect 15760 3600 15800 3605
rect 16340 3625 16380 3630
rect 16340 3595 16345 3625
rect 16375 3620 16380 3625
rect 16460 3625 16500 3630
rect 16460 3620 16465 3625
rect 16375 3600 16465 3620
rect 16375 3595 16380 3600
rect 16340 3590 16380 3595
rect 16460 3595 16465 3600
rect 16495 3620 16500 3625
rect 16580 3625 16620 3630
rect 16580 3620 16585 3625
rect 16495 3600 16585 3620
rect 16495 3595 16500 3600
rect 16460 3590 16500 3595
rect 16580 3595 16585 3600
rect 16615 3620 16620 3625
rect 16700 3625 16740 3630
rect 16700 3620 16705 3625
rect 16615 3600 16705 3620
rect 16615 3595 16620 3600
rect 16580 3590 16620 3595
rect 16700 3595 16705 3600
rect 16735 3620 16740 3625
rect 16820 3625 16860 3630
rect 16820 3620 16825 3625
rect 16735 3600 16825 3620
rect 16735 3595 16740 3600
rect 16700 3590 16740 3595
rect 16820 3595 16825 3600
rect 16855 3620 16860 3625
rect 16940 3625 16980 3630
rect 16940 3620 16945 3625
rect 16855 3600 16945 3620
rect 16855 3595 16860 3600
rect 16820 3590 16860 3595
rect 16940 3595 16945 3600
rect 16975 3620 16980 3625
rect 17060 3625 17100 3630
rect 17060 3620 17065 3625
rect 16975 3600 17065 3620
rect 16975 3595 16980 3600
rect 16940 3590 16980 3595
rect 17060 3595 17065 3600
rect 17095 3620 17100 3625
rect 17180 3625 17220 3630
rect 17180 3620 17185 3625
rect 17095 3600 17185 3620
rect 17095 3595 17100 3600
rect 17060 3590 17100 3595
rect 17180 3595 17185 3600
rect 17215 3620 17220 3625
rect 17300 3625 17340 3630
rect 17300 3620 17305 3625
rect 17215 3600 17305 3620
rect 17215 3595 17220 3600
rect 17180 3590 17220 3595
rect 17300 3595 17305 3600
rect 17335 3620 17340 3625
rect 17420 3625 17460 3630
rect 17420 3620 17425 3625
rect 17335 3600 17425 3620
rect 17335 3595 17340 3600
rect 17300 3590 17340 3595
rect 17420 3595 17425 3600
rect 17455 3595 17460 3625
rect 18000 3605 18005 3635
rect 18035 3630 18040 3635
rect 18110 3635 18150 3640
rect 18110 3630 18115 3635
rect 18035 3610 18115 3630
rect 18035 3605 18040 3610
rect 18000 3600 18040 3605
rect 18110 3605 18115 3610
rect 18145 3630 18150 3635
rect 18220 3635 18260 3640
rect 18220 3630 18225 3635
rect 18145 3610 18225 3630
rect 18145 3605 18150 3610
rect 18110 3600 18150 3605
rect 18220 3605 18225 3610
rect 18255 3630 18260 3635
rect 18330 3635 18370 3640
rect 18330 3630 18335 3635
rect 18255 3610 18335 3630
rect 18255 3605 18260 3610
rect 18220 3600 18260 3605
rect 18330 3605 18335 3610
rect 18365 3630 18370 3635
rect 18440 3635 18480 3640
rect 18440 3630 18445 3635
rect 18365 3610 18445 3630
rect 18365 3605 18370 3610
rect 18330 3600 18370 3605
rect 18440 3605 18445 3610
rect 18475 3630 18480 3635
rect 18550 3635 18590 3640
rect 18550 3630 18555 3635
rect 18475 3610 18555 3630
rect 18475 3605 18480 3610
rect 18440 3600 18480 3605
rect 18550 3605 18555 3610
rect 18585 3605 18590 3635
rect 18550 3600 18590 3605
rect 18805 3635 18845 3640
rect 18805 3605 18810 3635
rect 18840 3605 18845 3635
rect 18805 3600 18845 3605
rect 17420 3590 17460 3595
rect 14904 3555 15045 3560
rect -110 3525 -70 3530
rect -110 3495 -105 3525
rect -75 3520 -70 3525
rect 1261 3525 1301 3530
rect 1261 3520 1266 3525
rect -75 3500 1266 3520
rect -75 3495 -70 3500
rect -110 3490 -70 3495
rect 1261 3495 1266 3500
rect 1296 3495 1301 3525
rect 14904 3525 14910 3555
rect 14940 3525 14960 3555
rect 14990 3525 15010 3555
rect 15040 3525 15045 3555
rect 14904 3520 15045 3525
rect 18755 3555 18896 3560
rect 18755 3525 18760 3555
rect 18790 3525 18810 3555
rect 18840 3525 18860 3555
rect 18890 3525 18896 3555
rect 18755 3520 18896 3525
rect 1261 3490 1301 3495
rect 4440 3495 4480 3500
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect -15 3445 25 3450
rect -15 3415 -10 3445
rect 20 3440 25 3445
rect 940 3445 980 3450
rect 940 3440 945 3445
rect 20 3420 945 3440
rect 20 3415 25 3420
rect -15 3410 25 3415
rect 940 3415 945 3420
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3445 1685 3455
rect 2470 3450 2510 3455
rect 2470 3445 2475 3450
rect 1635 3415 1645 3445
rect 1675 3425 2475 3445
rect 1675 3415 1685 3425
rect 2470 3420 2475 3425
rect 2505 3420 2510 3450
rect 2470 3415 2510 3420
rect 5135 3445 5185 3455
rect 5135 3415 5145 3445
rect 5175 3440 5185 3445
rect 5550 3445 5590 3450
rect 5550 3440 5555 3445
rect 5175 3420 5555 3440
rect 5175 3415 5185 3420
rect 1635 3405 1685 3415
rect 5135 3405 5185 3415
rect 5550 3415 5555 3420
rect 5585 3415 5590 3445
rect 5550 3410 5590 3415
rect -60 3390 -20 3395
rect -60 3360 -55 3390
rect -25 3385 -20 3390
rect 2690 3390 2730 3395
rect 2690 3385 2695 3390
rect -25 3365 2695 3385
rect -25 3360 -20 3365
rect -60 3355 -20 3360
rect 2690 3360 2695 3365
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 1205 3340 1245 3345
rect 1205 3310 1210 3340
rect 1240 3335 1245 3340
rect 3135 3340 3175 3345
rect 3135 3335 3140 3340
rect 1240 3315 3140 3335
rect 1240 3310 1245 3315
rect 1205 3305 1245 3310
rect 3135 3310 3140 3315
rect 3170 3310 3175 3340
rect 3135 3305 3175 3310
rect 3385 3335 3435 3345
rect 3385 3305 3395 3335
rect 3425 3330 3435 3335
rect 5360 3335 5400 3340
rect 5360 3330 5365 3335
rect 3425 3310 5365 3330
rect 3425 3305 3435 3310
rect 3385 3295 3435 3305
rect 5360 3305 5365 3310
rect 5395 3305 5400 3335
rect 5360 3300 5400 3305
rect 1160 3285 1200 3290
rect 1160 3255 1165 3285
rect 1195 3280 1200 3285
rect 4885 3285 4925 3290
rect 4885 3280 4890 3285
rect 1195 3260 4890 3280
rect 1195 3255 1200 3260
rect 1160 3250 1200 3255
rect 4885 3255 4890 3260
rect 4920 3280 4925 3285
rect 5410 3285 5450 3290
rect 5410 3280 5415 3285
rect 4920 3260 5415 3280
rect 4920 3255 4925 3260
rect 4885 3250 4925 3255
rect 5410 3255 5415 3260
rect 5445 3255 5450 3285
rect 5410 3250 5450 3255
rect 2735 3240 2775 3245
rect 2735 3235 2740 3240
rect 46 3215 2740 3235
rect 46 3205 91 3215
rect 2735 3210 2740 3215
rect 2770 3210 2775 3240
rect 2735 3205 2775 3210
rect 46 3170 51 3205
rect 86 3170 91 3205
rect 1261 3165 1266 3200
rect 1301 3165 1306 3200
rect 2620 3185 2660 3190
rect 2620 3155 2625 3185
rect 2655 3180 2660 3185
rect 4440 3185 4480 3190
rect 4440 3180 4445 3185
rect 2655 3160 4445 3180
rect 2655 3155 2660 3160
rect 2620 3150 2660 3155
rect 4440 3155 4445 3160
rect 4475 3155 4480 3185
rect 4440 3150 4480 3155
rect 16050 3155 16090 3160
rect -110 3140 -70 3145
rect -110 3110 -105 3140
rect -75 3135 -70 3140
rect 46 3135 51 3145
rect -75 3115 51 3135
rect -75 3110 -70 3115
rect 46 3110 51 3115
rect 86 3110 91 3145
rect 3135 3140 3175 3145
rect -110 3105 -70 3110
rect 1261 3105 1266 3140
rect 1301 3105 1306 3140
rect 3135 3110 3140 3140
rect 3170 3135 3175 3140
rect 4835 3140 4875 3145
rect 4835 3135 4840 3140
rect 3170 3115 4840 3135
rect 3170 3110 3175 3115
rect 3135 3105 3175 3110
rect 4835 3110 4840 3115
rect 4870 3135 4875 3140
rect 5315 3140 5355 3145
rect 5315 3135 5320 3140
rect 4870 3115 5320 3135
rect 4870 3110 4875 3115
rect 4835 3105 4875 3110
rect 5315 3110 5320 3115
rect 5350 3110 5355 3140
rect 16050 3125 16055 3155
rect 16085 3150 16090 3155
rect 16823 3155 16857 3160
rect 16823 3150 16826 3155
rect 16085 3130 16826 3150
rect 16085 3125 16090 3130
rect 16050 3120 16090 3125
rect 16823 3125 16826 3130
rect 16854 3125 16857 3155
rect 16823 3120 16857 3125
rect 5315 3105 5355 3110
rect 1160 3100 1200 3105
rect 1160 3095 1165 3100
rect 46 3075 1165 3095
rect 46 3065 91 3075
rect 1160 3070 1165 3075
rect 1195 3070 1200 3100
rect 16280 3100 16320 3105
rect 1160 3065 1200 3070
rect 3985 3080 4025 3085
rect 46 3030 51 3065
rect 86 3030 91 3065
rect 3985 3050 3990 3080
rect 4020 3075 4025 3080
rect 4020 3055 6100 3075
rect 16280 3070 16285 3100
rect 16315 3095 16320 3100
rect 16520 3100 16560 3105
rect 16520 3095 16525 3100
rect 16315 3075 16525 3095
rect 16315 3070 16320 3075
rect 16280 3065 16320 3070
rect 16520 3070 16525 3075
rect 16555 3095 16560 3100
rect 16760 3100 16800 3105
rect 16760 3095 16765 3100
rect 16555 3075 16765 3095
rect 16555 3070 16560 3075
rect 16520 3065 16560 3070
rect 16760 3070 16765 3075
rect 16795 3095 16800 3100
rect 17000 3100 17040 3105
rect 17000 3095 17005 3100
rect 16795 3075 17005 3095
rect 16795 3070 16800 3075
rect 16760 3065 16800 3070
rect 17000 3070 17005 3075
rect 17035 3095 17040 3100
rect 17240 3100 17280 3105
rect 17240 3095 17245 3100
rect 17035 3075 17245 3095
rect 17035 3070 17040 3075
rect 17000 3065 17040 3070
rect 17240 3070 17245 3075
rect 17275 3095 17280 3100
rect 17480 3100 17520 3105
rect 17480 3095 17485 3100
rect 17275 3075 17485 3095
rect 17275 3070 17280 3075
rect 17240 3065 17280 3070
rect 17480 3070 17485 3075
rect 17515 3070 17520 3100
rect 17480 3065 17520 3070
rect 16400 3055 16440 3060
rect 4020 3050 4025 3055
rect 3985 3045 4025 3050
rect 3445 3035 3485 3040
rect 3445 3005 3450 3035
rect 3480 3030 3485 3035
rect 3805 3035 3845 3040
rect 3805 3030 3810 3035
rect 3480 3010 3810 3030
rect 3480 3005 3485 3010
rect -110 3000 -70 3005
rect -110 2970 -105 3000
rect -75 2995 -70 3000
rect 46 2995 51 3005
rect -75 2975 51 2995
rect -75 2970 -70 2975
rect 46 2970 51 2975
rect 86 2970 91 3005
rect 3445 3000 3485 3005
rect 3805 3005 3810 3010
rect 3840 3030 3845 3035
rect 4345 3035 4385 3040
rect 4345 3030 4350 3035
rect 3840 3010 4350 3030
rect 3840 3005 3845 3010
rect 3805 3000 3845 3005
rect 4345 3005 4350 3010
rect 4380 3030 4385 3035
rect 4705 3035 4745 3040
rect 4705 3030 4710 3035
rect 4380 3010 4710 3030
rect 4380 3005 4385 3010
rect 4345 3000 4385 3005
rect 4705 3005 4710 3010
rect 4740 3030 4745 3035
rect 4740 3010 6100 3030
rect 16400 3025 16405 3055
rect 16435 3050 16440 3055
rect 16640 3055 16680 3060
rect 16640 3050 16645 3055
rect 16435 3030 16645 3050
rect 16435 3025 16440 3030
rect 16400 3020 16440 3025
rect 16640 3025 16645 3030
rect 16675 3050 16680 3055
rect 16880 3055 16920 3060
rect 16880 3050 16885 3055
rect 16675 3030 16885 3050
rect 16675 3025 16680 3030
rect 16640 3020 16680 3025
rect 16880 3025 16885 3030
rect 16915 3050 16920 3055
rect 17120 3055 17160 3060
rect 17120 3050 17125 3055
rect 16915 3030 17125 3050
rect 16915 3025 16920 3030
rect 16880 3020 16920 3025
rect 17120 3025 17125 3030
rect 17155 3050 17160 3055
rect 17360 3055 17400 3060
rect 17360 3050 17365 3055
rect 17155 3030 17365 3050
rect 17155 3025 17160 3030
rect 17120 3020 17160 3025
rect 17360 3025 17365 3030
rect 17395 3025 17400 3055
rect 17360 3020 17400 3025
rect 4740 3005 4745 3010
rect 4705 3000 4745 3005
rect 16340 3000 16380 3005
rect 2520 2980 2560 2985
rect -110 2965 -70 2970
rect 2330 2925 2335 2960
rect 2370 2950 2375 2960
rect 2425 2955 2465 2960
rect 2425 2950 2430 2955
rect 2370 2930 2430 2950
rect 2370 2925 2375 2930
rect 2425 2925 2430 2930
rect 2460 2925 2465 2955
rect 2520 2950 2525 2980
rect 2555 2975 2560 2980
rect 3080 2980 3120 2985
rect 3080 2975 3085 2980
rect 2555 2955 3085 2975
rect 2555 2950 2560 2955
rect 2520 2945 2560 2950
rect 3080 2950 3085 2955
rect 3115 2950 3120 2980
rect 3080 2945 3120 2950
rect 3265 2980 3305 2985
rect 3265 2950 3270 2980
rect 3300 2975 3305 2980
rect 3625 2980 3665 2985
rect 3625 2975 3630 2980
rect 3300 2955 3630 2975
rect 3300 2950 3305 2955
rect 3265 2945 3305 2950
rect 3625 2950 3630 2955
rect 3660 2975 3665 2980
rect 4165 2980 4205 2985
rect 4165 2975 4170 2980
rect 3660 2955 4170 2975
rect 3660 2950 3665 2955
rect 3625 2945 3665 2950
rect 4165 2950 4170 2955
rect 4200 2975 4205 2980
rect 4525 2980 4565 2985
rect 4525 2975 4530 2980
rect 4200 2955 4530 2975
rect 4200 2950 4205 2955
rect 4165 2945 4205 2950
rect 4525 2950 4530 2955
rect 4560 2975 4565 2980
rect 4560 2955 6100 2975
rect 16340 2970 16345 3000
rect 16375 2995 16380 3000
rect 16400 3000 16440 3005
rect 16400 2995 16405 3000
rect 16375 2975 16405 2995
rect 16375 2970 16380 2975
rect 15265 2965 15305 2970
rect 4560 2950 4565 2955
rect 4525 2945 4565 2950
rect 2425 2920 2465 2925
rect 14904 2935 15045 2940
rect -110 2910 -70 2915
rect -110 2880 -105 2910
rect -75 2905 -70 2910
rect 905 2910 1125 2920
rect 905 2905 920 2910
rect -75 2885 920 2905
rect -75 2880 -70 2885
rect -110 2875 -70 2880
rect 905 2880 920 2885
rect 950 2880 1000 2910
rect 1030 2880 1080 2910
rect 1110 2880 1125 2910
rect 14904 2905 14910 2935
rect 14940 2905 14960 2935
rect 14990 2905 15010 2935
rect 15040 2905 15045 2935
rect 15265 2935 15270 2965
rect 15300 2960 15305 2965
rect 15375 2965 15415 2970
rect 15375 2960 15380 2965
rect 15300 2940 15380 2960
rect 15300 2935 15305 2940
rect 15265 2930 15305 2935
rect 15375 2935 15380 2940
rect 15410 2960 15415 2965
rect 15485 2965 15525 2970
rect 15485 2960 15490 2965
rect 15410 2940 15490 2960
rect 15410 2935 15415 2940
rect 15375 2930 15415 2935
rect 15485 2935 15490 2940
rect 15520 2960 15525 2965
rect 15595 2965 15635 2970
rect 15595 2960 15600 2965
rect 15520 2940 15600 2960
rect 15520 2935 15525 2940
rect 15485 2930 15525 2935
rect 15595 2935 15600 2940
rect 15630 2960 15635 2965
rect 15705 2965 15745 2970
rect 16340 2965 16380 2970
rect 16400 2970 16405 2975
rect 16435 2995 16440 3000
rect 16580 3000 16620 3005
rect 16580 2995 16585 3000
rect 16435 2975 16585 2995
rect 16435 2970 16440 2975
rect 16400 2965 16440 2970
rect 16580 2970 16585 2975
rect 16615 2995 16620 3000
rect 16820 3000 16860 3005
rect 16820 2995 16825 3000
rect 16615 2975 16825 2995
rect 16615 2970 16620 2975
rect 16580 2965 16620 2970
rect 16820 2970 16825 2975
rect 16855 2995 16860 3000
rect 17060 3000 17100 3005
rect 17060 2995 17065 3000
rect 16855 2975 17065 2995
rect 16855 2970 16860 2975
rect 16820 2965 16860 2970
rect 17060 2970 17065 2975
rect 17095 2995 17100 3000
rect 17300 3000 17340 3005
rect 17300 2995 17305 3000
rect 17095 2975 17305 2995
rect 17095 2970 17100 2975
rect 17060 2965 17100 2970
rect 17300 2970 17305 2975
rect 17335 2970 17340 3000
rect 17300 2965 17340 2970
rect 18055 2965 18095 2970
rect 15705 2960 15710 2965
rect 15630 2940 15710 2960
rect 15630 2935 15635 2940
rect 15595 2930 15635 2935
rect 15705 2935 15710 2940
rect 15740 2935 15745 2965
rect 15705 2930 15745 2935
rect 16460 2945 16500 2950
rect 16460 2915 16465 2945
rect 16495 2940 16500 2945
rect 16700 2945 16740 2950
rect 16700 2940 16705 2945
rect 16495 2920 16705 2940
rect 16495 2915 16500 2920
rect 16460 2910 16500 2915
rect 16700 2915 16705 2920
rect 16735 2940 16740 2945
rect 16940 2945 16980 2950
rect 16940 2940 16945 2945
rect 16735 2920 16945 2940
rect 16735 2915 16740 2920
rect 16700 2910 16740 2915
rect 16940 2915 16945 2920
rect 16975 2940 16980 2945
rect 17180 2945 17220 2950
rect 17180 2940 17185 2945
rect 16975 2920 17185 2940
rect 16975 2915 16980 2920
rect 16940 2910 16980 2915
rect 17180 2915 17185 2920
rect 17215 2940 17220 2945
rect 17420 2945 17460 2950
rect 17420 2940 17425 2945
rect 17215 2920 17425 2940
rect 17215 2915 17220 2920
rect 17180 2910 17220 2915
rect 17420 2915 17425 2920
rect 17455 2940 17460 2945
rect 17480 2945 17520 2950
rect 17480 2940 17485 2945
rect 17455 2920 17485 2940
rect 17455 2915 17460 2920
rect 17420 2910 17460 2915
rect 17480 2915 17485 2920
rect 17515 2915 17520 2945
rect 18055 2935 18060 2965
rect 18090 2960 18095 2965
rect 18165 2965 18205 2970
rect 18165 2960 18170 2965
rect 18090 2940 18170 2960
rect 18090 2935 18095 2940
rect 18055 2930 18095 2935
rect 18165 2935 18170 2940
rect 18200 2960 18205 2965
rect 18275 2965 18315 2970
rect 18275 2960 18280 2965
rect 18200 2940 18280 2960
rect 18200 2935 18205 2940
rect 18165 2930 18205 2935
rect 18275 2935 18280 2940
rect 18310 2960 18315 2965
rect 18385 2965 18425 2970
rect 18385 2960 18390 2965
rect 18310 2940 18390 2960
rect 18310 2935 18315 2940
rect 18275 2930 18315 2935
rect 18385 2935 18390 2940
rect 18420 2960 18425 2965
rect 18495 2965 18535 2970
rect 18495 2960 18500 2965
rect 18420 2940 18500 2960
rect 18420 2935 18425 2940
rect 18385 2930 18425 2935
rect 18495 2935 18500 2940
rect 18530 2935 18535 2965
rect 18495 2930 18535 2935
rect 18755 2935 18896 2940
rect 17480 2910 17520 2915
rect 905 2870 1125 2880
rect 2330 2900 2375 2905
rect 14904 2900 15045 2905
rect 18755 2905 18760 2935
rect 18790 2905 18810 2935
rect 18840 2905 18860 2935
rect 18890 2905 18896 2935
rect 18755 2900 18896 2905
rect 2330 2865 2335 2900
rect 2370 2865 2375 2900
rect 2330 2860 2375 2865
rect 14955 2880 14995 2885
rect -60 2855 -20 2860
rect -60 2825 -55 2855
rect -25 2850 -20 2855
rect 51 2850 56 2855
rect -25 2830 56 2850
rect -25 2825 -20 2830
rect -60 2820 -20 2825
rect 51 2820 56 2830
rect 91 2820 96 2855
rect 724 2820 729 2855
rect 764 2845 769 2855
rect 1205 2850 1245 2855
rect 1205 2845 1210 2850
rect 764 2825 1210 2845
rect 764 2820 769 2825
rect 1205 2820 1210 2825
rect 1240 2820 1245 2850
rect 14955 2850 14960 2880
rect 14990 2875 14995 2880
rect 15650 2880 15690 2885
rect 15650 2875 15655 2880
rect 14990 2855 15655 2875
rect 14990 2850 14995 2855
rect 14955 2845 14995 2850
rect 15650 2850 15655 2855
rect 15685 2875 15690 2880
rect 16000 2880 16040 2885
rect 16000 2875 16005 2880
rect 15685 2855 16005 2875
rect 15685 2850 15690 2855
rect 15650 2845 15690 2850
rect 16000 2850 16005 2855
rect 16035 2850 16040 2880
rect 16000 2845 16040 2850
rect 17690 2880 17730 2885
rect 17690 2850 17695 2880
rect 17725 2875 17730 2880
rect 18110 2880 18150 2885
rect 18110 2875 18115 2880
rect 17725 2855 18115 2875
rect 17725 2850 17730 2855
rect 17690 2845 17730 2850
rect 18110 2850 18115 2855
rect 18145 2875 18150 2880
rect 18805 2880 18845 2885
rect 18805 2875 18810 2880
rect 18145 2855 18810 2875
rect 18145 2850 18150 2855
rect 18110 2845 18150 2850
rect 18805 2850 18810 2855
rect 18840 2850 18845 2880
rect 18805 2845 18845 2850
rect 1205 2815 1245 2820
rect 1261 2805 1266 2840
rect 1301 2805 1306 2840
rect 1960 2805 1965 2840
rect 2000 2830 2005 2840
rect 2330 2835 2370 2840
rect 2330 2830 2335 2835
rect 2000 2810 2335 2830
rect 2000 2805 2005 2810
rect 2330 2805 2335 2810
rect 2365 2805 2370 2835
rect 14515 2825 14555 2830
rect 2330 2800 2370 2805
rect 2995 2810 3035 2815
rect -15 2795 25 2800
rect -15 2765 -10 2795
rect 20 2785 25 2795
rect 51 2785 56 2795
rect 20 2765 56 2785
rect -15 2760 25 2765
rect 51 2760 56 2765
rect 91 2760 96 2795
rect 724 2760 729 2795
rect 764 2785 769 2795
rect 2620 2790 2660 2795
rect 2620 2785 2625 2790
rect 764 2765 2625 2785
rect 764 2760 769 2765
rect 2620 2760 2625 2765
rect 2655 2760 2660 2790
rect 2995 2780 3000 2810
rect 3030 2805 3035 2810
rect 3175 2810 3215 2815
rect 3175 2805 3180 2810
rect 3030 2785 3180 2805
rect 3030 2780 3035 2785
rect 2995 2775 3035 2780
rect 3175 2780 3180 2785
rect 3210 2805 3215 2810
rect 3355 2810 3395 2815
rect 3355 2805 3360 2810
rect 3210 2785 3360 2805
rect 3210 2780 3215 2785
rect 3175 2775 3215 2780
rect 3355 2780 3360 2785
rect 3390 2805 3395 2810
rect 3535 2810 3575 2815
rect 3535 2805 3540 2810
rect 3390 2785 3540 2805
rect 3390 2780 3395 2785
rect 3355 2775 3395 2780
rect 3535 2780 3540 2785
rect 3570 2805 3575 2810
rect 3715 2810 3755 2815
rect 3715 2805 3720 2810
rect 3570 2785 3720 2805
rect 3570 2780 3575 2785
rect 3535 2775 3575 2780
rect 3715 2780 3720 2785
rect 3750 2805 3755 2810
rect 3895 2810 3935 2815
rect 3895 2805 3900 2810
rect 3750 2785 3900 2805
rect 3750 2780 3755 2785
rect 3715 2775 3755 2780
rect 3895 2780 3900 2785
rect 3930 2805 3935 2810
rect 4075 2810 4115 2815
rect 4075 2805 4080 2810
rect 3930 2785 4080 2805
rect 3930 2780 3935 2785
rect 3895 2775 3935 2780
rect 4075 2780 4080 2785
rect 4110 2805 4115 2810
rect 4255 2810 4295 2815
rect 4255 2805 4260 2810
rect 4110 2785 4260 2805
rect 4110 2780 4115 2785
rect 4075 2775 4115 2780
rect 4255 2780 4260 2785
rect 4290 2805 4295 2810
rect 4435 2810 4475 2815
rect 4435 2805 4440 2810
rect 4290 2785 4440 2805
rect 4290 2780 4295 2785
rect 4255 2775 4295 2780
rect 4435 2780 4440 2785
rect 4470 2805 4475 2810
rect 4615 2810 4655 2815
rect 4615 2805 4620 2810
rect 4470 2785 4620 2805
rect 4470 2780 4475 2785
rect 4435 2775 4475 2780
rect 4615 2780 4620 2785
rect 4650 2805 4655 2810
rect 4795 2810 4835 2815
rect 4795 2805 4800 2810
rect 4650 2785 4800 2805
rect 4650 2780 4655 2785
rect 4615 2775 4655 2780
rect 4795 2780 4800 2785
rect 4830 2805 4835 2810
rect 4975 2810 5015 2815
rect 4975 2805 4980 2810
rect 4830 2785 4980 2805
rect 4830 2780 4835 2785
rect 4795 2775 4835 2780
rect 4975 2780 4980 2785
rect 5010 2805 5015 2810
rect 5550 2810 5590 2815
rect 5550 2805 5555 2810
rect 5010 2785 5555 2805
rect 5010 2780 5015 2785
rect 4975 2775 5015 2780
rect 5550 2780 5555 2785
rect 5585 2780 5590 2810
rect 14515 2795 14520 2825
rect 14550 2820 14555 2825
rect 15375 2825 15415 2830
rect 15375 2820 15380 2825
rect 14550 2800 15380 2820
rect 14550 2795 14555 2800
rect 14515 2790 14555 2795
rect 15375 2795 15380 2800
rect 15410 2795 15415 2825
rect 15375 2790 15415 2795
rect 18385 2825 18425 2830
rect 18385 2795 18390 2825
rect 18420 2820 18425 2825
rect 19245 2825 19285 2830
rect 19245 2820 19250 2825
rect 18420 2800 19250 2820
rect 18420 2795 18425 2800
rect 18385 2790 18425 2795
rect 19245 2795 19250 2800
rect 19280 2795 19285 2825
rect 19245 2790 19285 2795
rect 5550 2775 5590 2780
rect 2620 2755 2660 2760
rect 3175 2750 3215 2755
rect 1261 2745 1301 2750
rect 1261 2715 1266 2745
rect 1296 2740 1301 2745
rect 2150 2745 2190 2750
rect 2150 2740 2155 2745
rect 1296 2720 2155 2740
rect 1296 2715 1301 2720
rect 1261 2710 1301 2715
rect 2150 2715 2155 2720
rect 2185 2715 2190 2745
rect 3175 2720 3180 2750
rect 3210 2745 3215 2750
rect 3355 2750 3395 2755
rect 3355 2745 3360 2750
rect 3210 2725 3360 2745
rect 3210 2720 3215 2725
rect 3175 2715 3215 2720
rect 3355 2720 3360 2725
rect 3390 2745 3395 2750
rect 3535 2750 3575 2755
rect 3535 2745 3540 2750
rect 3390 2725 3540 2745
rect 3390 2720 3395 2725
rect 3355 2715 3395 2720
rect 3535 2720 3540 2725
rect 3570 2745 3575 2750
rect 3715 2750 3755 2755
rect 3715 2745 3720 2750
rect 3570 2725 3720 2745
rect 3570 2720 3575 2725
rect 3535 2715 3575 2720
rect 3715 2720 3720 2725
rect 3750 2745 3755 2750
rect 3895 2750 3935 2755
rect 3895 2745 3900 2750
rect 3750 2725 3900 2745
rect 3750 2720 3755 2725
rect 3715 2715 3755 2720
rect 3895 2720 3900 2725
rect 3930 2745 3935 2750
rect 4075 2750 4115 2755
rect 4075 2745 4080 2750
rect 3930 2725 4080 2745
rect 3930 2720 3935 2725
rect 3895 2715 3935 2720
rect 4075 2720 4080 2725
rect 4110 2745 4115 2750
rect 4255 2750 4295 2755
rect 4255 2745 4260 2750
rect 4110 2725 4260 2745
rect 4110 2720 4115 2725
rect 4075 2715 4115 2720
rect 4255 2720 4260 2725
rect 4290 2745 4295 2750
rect 4435 2750 4475 2755
rect 4435 2745 4440 2750
rect 4290 2725 4440 2745
rect 4290 2720 4295 2725
rect 4255 2715 4295 2720
rect 4435 2720 4440 2725
rect 4470 2745 4475 2750
rect 4615 2750 4655 2755
rect 4615 2745 4620 2750
rect 4470 2725 4620 2745
rect 4470 2720 4475 2725
rect 4435 2715 4475 2720
rect 4615 2720 4620 2725
rect 4650 2745 4655 2750
rect 4795 2750 4835 2755
rect 4795 2745 4800 2750
rect 4650 2725 4800 2745
rect 4650 2720 4655 2725
rect 4615 2715 4655 2720
rect 4795 2720 4800 2725
rect 4830 2720 4835 2750
rect 4795 2715 4835 2720
rect 2150 2710 2190 2715
rect 15210 2705 15250 2710
rect 15210 2675 15215 2705
rect 15245 2700 15250 2705
rect 15320 2705 15360 2710
rect 15320 2700 15325 2705
rect 15245 2680 15325 2700
rect 15245 2675 15250 2680
rect 15210 2670 15250 2675
rect 15320 2675 15325 2680
rect 15355 2700 15360 2705
rect 15430 2705 15470 2710
rect 15430 2700 15435 2705
rect 15355 2680 15435 2700
rect 15355 2675 15360 2680
rect 15320 2670 15360 2675
rect 15430 2675 15435 2680
rect 15465 2700 15470 2705
rect 15540 2705 15580 2710
rect 15540 2700 15545 2705
rect 15465 2680 15545 2700
rect 15465 2675 15470 2680
rect 15430 2670 15470 2675
rect 15540 2675 15545 2680
rect 15575 2700 15580 2705
rect 15650 2705 15690 2710
rect 15650 2700 15655 2705
rect 15575 2680 15655 2700
rect 15575 2675 15580 2680
rect 15540 2670 15580 2675
rect 15650 2675 15655 2680
rect 15685 2700 15690 2705
rect 15760 2705 15800 2710
rect 15760 2700 15765 2705
rect 15685 2680 15765 2700
rect 15685 2675 15690 2680
rect 15650 2670 15690 2675
rect 15760 2675 15765 2680
rect 15795 2675 15800 2705
rect 15760 2670 15800 2675
rect 18000 2705 18040 2710
rect 18000 2675 18005 2705
rect 18035 2700 18040 2705
rect 18110 2705 18150 2710
rect 18110 2700 18115 2705
rect 18035 2680 18115 2700
rect 18035 2675 18040 2680
rect 18000 2670 18040 2675
rect 18110 2675 18115 2680
rect 18145 2700 18150 2705
rect 18220 2705 18260 2710
rect 18220 2700 18225 2705
rect 18145 2680 18225 2700
rect 18145 2675 18150 2680
rect 18110 2670 18150 2675
rect 18220 2675 18225 2680
rect 18255 2700 18260 2705
rect 18330 2705 18370 2710
rect 18330 2700 18335 2705
rect 18255 2680 18335 2700
rect 18255 2675 18260 2680
rect 18220 2670 18260 2675
rect 18330 2675 18335 2680
rect 18365 2700 18370 2705
rect 18440 2705 18480 2710
rect 18440 2700 18445 2705
rect 18365 2680 18445 2700
rect 18365 2675 18370 2680
rect 18330 2670 18370 2675
rect 18440 2675 18445 2680
rect 18475 2700 18480 2705
rect 18550 2705 18590 2710
rect 18550 2700 18555 2705
rect 18475 2680 18555 2700
rect 18475 2675 18480 2680
rect 18440 2670 18480 2675
rect 18550 2675 18555 2680
rect 18585 2675 18590 2705
rect 18550 2670 18590 2675
rect 16105 2475 16145 2480
rect 16105 2445 16110 2475
rect 16140 2470 16145 2475
rect 16823 2475 16857 2480
rect 16823 2470 16826 2475
rect 16140 2450 16826 2470
rect 16140 2445 16145 2450
rect 16105 2440 16145 2445
rect 16823 2445 16826 2450
rect 16854 2445 16857 2475
rect 16823 2440 16857 2445
rect 15020 2435 15060 2440
rect 15020 2405 15025 2435
rect 15055 2430 15060 2435
rect 15265 2435 15305 2440
rect 15265 2430 15270 2435
rect 15055 2410 15270 2430
rect 15055 2405 15060 2410
rect 15020 2400 15060 2405
rect 15265 2405 15270 2410
rect 15300 2430 15305 2435
rect 15375 2435 15415 2440
rect 15375 2430 15380 2435
rect 15300 2410 15380 2430
rect 15300 2405 15305 2410
rect 15265 2400 15305 2405
rect 15375 2405 15380 2410
rect 15410 2430 15415 2435
rect 15485 2435 15525 2440
rect 15485 2430 15490 2435
rect 15410 2410 15490 2430
rect 15410 2405 15415 2410
rect 15375 2400 15415 2405
rect 15485 2405 15490 2410
rect 15520 2430 15525 2435
rect 15595 2435 15635 2440
rect 15595 2430 15600 2435
rect 15520 2410 15600 2430
rect 15520 2405 15525 2410
rect 15485 2400 15525 2405
rect 15595 2405 15600 2410
rect 15630 2430 15635 2435
rect 15705 2435 15745 2440
rect 15705 2430 15710 2435
rect 15630 2410 15710 2430
rect 15630 2405 15635 2410
rect 15595 2400 15635 2405
rect 15705 2405 15710 2410
rect 15740 2405 15745 2435
rect 18055 2435 18095 2440
rect 16000 2420 16040 2425
rect 16000 2415 16005 2420
rect 15705 2400 15745 2405
rect 15785 2395 16005 2415
rect 15765 2390 15805 2395
rect 3805 2380 3845 2385
rect 3355 2375 3395 2380
rect 2620 2345 2660 2350
rect 2620 2315 2625 2345
rect 2655 2340 2660 2345
rect 3355 2345 3360 2375
rect 3390 2345 3395 2375
rect 3805 2350 3810 2380
rect 3840 2375 3845 2380
rect 4165 2380 4205 2385
rect 4165 2375 4170 2380
rect 3840 2355 4170 2375
rect 3840 2350 3845 2355
rect 3805 2345 3845 2350
rect 4165 2350 4170 2355
rect 4200 2350 4205 2380
rect 15765 2360 15770 2390
rect 15800 2360 15805 2390
rect 16000 2390 16005 2395
rect 16035 2415 16040 2420
rect 16280 2420 16320 2425
rect 16280 2415 16285 2420
rect 16035 2395 16285 2415
rect 16035 2390 16040 2395
rect 16000 2385 16040 2390
rect 16280 2390 16285 2395
rect 16315 2415 16320 2420
rect 16520 2420 16560 2425
rect 16520 2415 16525 2420
rect 16315 2395 16525 2415
rect 16315 2390 16320 2395
rect 16280 2385 16320 2390
rect 16520 2390 16525 2395
rect 16555 2415 16560 2420
rect 16760 2420 16800 2425
rect 16760 2415 16765 2420
rect 16555 2395 16765 2415
rect 16555 2390 16560 2395
rect 16520 2385 16560 2390
rect 16760 2390 16765 2395
rect 16795 2415 16800 2420
rect 17000 2420 17040 2425
rect 17000 2415 17005 2420
rect 16795 2395 17005 2415
rect 16795 2390 16800 2395
rect 16760 2385 16800 2390
rect 17000 2390 17005 2395
rect 17035 2415 17040 2420
rect 17240 2420 17280 2425
rect 17240 2415 17245 2420
rect 17035 2395 17245 2415
rect 17035 2390 17040 2395
rect 17000 2385 17040 2390
rect 17240 2390 17245 2395
rect 17275 2415 17280 2420
rect 17480 2420 17520 2425
rect 17480 2415 17485 2420
rect 17275 2395 17485 2415
rect 17275 2390 17280 2395
rect 17240 2385 17280 2390
rect 17480 2390 17485 2395
rect 17515 2390 17520 2420
rect 18055 2405 18060 2435
rect 18090 2430 18095 2435
rect 18165 2435 18205 2440
rect 18165 2430 18170 2435
rect 18090 2410 18170 2430
rect 18090 2405 18095 2410
rect 18055 2400 18095 2405
rect 18165 2405 18170 2410
rect 18200 2430 18205 2435
rect 18275 2435 18315 2440
rect 18275 2430 18280 2435
rect 18200 2410 18280 2430
rect 18200 2405 18205 2410
rect 18165 2400 18205 2405
rect 18275 2405 18280 2410
rect 18310 2430 18315 2435
rect 18385 2435 18425 2440
rect 18385 2430 18390 2435
rect 18310 2410 18390 2430
rect 18310 2405 18315 2410
rect 18275 2400 18315 2405
rect 18385 2405 18390 2410
rect 18420 2430 18425 2435
rect 18495 2435 18535 2440
rect 18495 2430 18500 2435
rect 18420 2410 18500 2430
rect 18420 2405 18425 2410
rect 18385 2400 18425 2405
rect 18495 2405 18500 2410
rect 18530 2430 18535 2435
rect 18740 2435 18780 2440
rect 18740 2430 18745 2435
rect 18530 2410 18745 2430
rect 18530 2405 18535 2410
rect 18495 2400 18535 2405
rect 18740 2405 18745 2410
rect 18775 2405 18780 2435
rect 18740 2400 18780 2405
rect 17480 2385 17520 2390
rect 15765 2355 15805 2360
rect 16400 2375 16440 2380
rect 4165 2345 4205 2350
rect 16400 2345 16405 2375
rect 16435 2370 16440 2375
rect 16640 2375 16680 2380
rect 16640 2370 16645 2375
rect 16435 2350 16645 2370
rect 16435 2345 16440 2350
rect 3355 2340 3395 2345
rect 16400 2340 16440 2345
rect 16640 2345 16645 2350
rect 16675 2370 16680 2375
rect 16880 2375 16920 2380
rect 16880 2370 16885 2375
rect 16675 2350 16885 2370
rect 16675 2345 16680 2350
rect 16640 2340 16680 2345
rect 16880 2345 16885 2350
rect 16915 2370 16920 2375
rect 17120 2375 17160 2380
rect 17120 2370 17125 2375
rect 16915 2350 17125 2370
rect 16915 2345 16920 2350
rect 16880 2340 16920 2345
rect 17120 2345 17125 2350
rect 17155 2370 17160 2375
rect 17360 2375 17400 2380
rect 17360 2370 17365 2375
rect 17155 2350 17365 2370
rect 17155 2345 17160 2350
rect 17120 2340 17160 2345
rect 17360 2345 17365 2350
rect 17395 2370 17400 2375
rect 17690 2375 17730 2380
rect 17690 2370 17695 2375
rect 17395 2350 17695 2370
rect 17395 2345 17400 2350
rect 17360 2340 17400 2345
rect 17690 2345 17695 2350
rect 17725 2370 17730 2375
rect 18025 2375 18065 2380
rect 18025 2370 18030 2375
rect 17725 2350 18030 2370
rect 17725 2345 17730 2350
rect 17690 2340 17730 2345
rect 18025 2345 18030 2350
rect 18060 2345 18065 2375
rect 18025 2340 18065 2345
rect 2655 2320 3395 2340
rect 3625 2335 3665 2340
rect 2655 2315 2660 2320
rect 2620 2310 2660 2315
rect 3625 2305 3630 2335
rect 3660 2330 3665 2335
rect 4345 2335 4385 2340
rect 4345 2330 4350 2335
rect 3660 2310 4350 2330
rect 3660 2305 3665 2310
rect 3625 2300 3665 2305
rect 4345 2305 4350 2310
rect 4380 2305 4385 2335
rect 16000 2325 16040 2330
rect 4345 2300 4385 2305
rect 15065 2315 15105 2320
rect 2735 2290 2775 2295
rect 2735 2260 2740 2290
rect 2770 2285 2775 2290
rect 3445 2290 3485 2295
rect 3445 2285 3450 2290
rect 2770 2265 3450 2285
rect 2770 2260 2775 2265
rect 2735 2255 2775 2260
rect 3445 2260 3450 2265
rect 3480 2285 3485 2290
rect 4525 2290 4565 2295
rect 4525 2285 4530 2290
rect 3480 2265 4530 2285
rect 3480 2260 3485 2265
rect 3445 2255 3485 2260
rect 4525 2260 4530 2265
rect 4560 2285 4565 2290
rect 5270 2290 5310 2295
rect 5270 2285 5275 2290
rect 4560 2265 5275 2285
rect 4560 2260 4565 2265
rect 4525 2255 4565 2260
rect 5270 2260 5275 2265
rect 5305 2260 5310 2290
rect 15065 2285 15070 2315
rect 15100 2310 15105 2315
rect 15265 2315 15305 2320
rect 15265 2310 15270 2315
rect 15100 2290 15270 2310
rect 15100 2285 15105 2290
rect 15065 2280 15105 2285
rect 15265 2285 15270 2290
rect 15300 2310 15305 2315
rect 15375 2315 15415 2320
rect 15375 2310 15380 2315
rect 15300 2290 15380 2310
rect 15300 2285 15305 2290
rect 15265 2280 15305 2285
rect 15375 2285 15380 2290
rect 15410 2310 15415 2315
rect 15485 2315 15525 2320
rect 15485 2310 15490 2315
rect 15410 2290 15490 2310
rect 15410 2285 15415 2290
rect 15375 2280 15415 2285
rect 15485 2285 15490 2290
rect 15520 2310 15525 2315
rect 15595 2315 15635 2320
rect 15595 2310 15600 2315
rect 15520 2290 15600 2310
rect 15520 2285 15525 2290
rect 15485 2280 15525 2285
rect 15595 2285 15600 2290
rect 15630 2310 15635 2315
rect 15705 2315 15745 2320
rect 15705 2310 15710 2315
rect 15630 2290 15710 2310
rect 15630 2285 15635 2290
rect 15595 2280 15635 2285
rect 15705 2285 15710 2290
rect 15740 2285 15745 2315
rect 16000 2295 16005 2325
rect 16035 2320 16040 2325
rect 17760 2325 17800 2330
rect 17760 2320 17765 2325
rect 16035 2300 17765 2320
rect 16035 2295 16040 2300
rect 16000 2290 16040 2295
rect 17760 2295 17765 2300
rect 17795 2295 17800 2325
rect 17760 2290 17800 2295
rect 18055 2315 18095 2320
rect 18055 2285 18060 2315
rect 18090 2310 18095 2315
rect 18165 2315 18205 2320
rect 18165 2310 18170 2315
rect 18090 2290 18170 2310
rect 18090 2285 18095 2290
rect 15705 2280 15745 2285
rect 16440 2280 16480 2285
rect 5270 2255 5310 2260
rect 16440 2250 16445 2280
rect 16475 2275 16480 2280
rect 16660 2280 16700 2285
rect 16660 2275 16665 2280
rect 16475 2255 16665 2275
rect 16475 2250 16480 2255
rect 2425 2245 2465 2250
rect 2425 2215 2430 2245
rect 2460 2240 2465 2245
rect 3805 2245 3845 2250
rect 16440 2245 16480 2250
rect 16660 2250 16665 2255
rect 16695 2275 16700 2280
rect 16880 2280 16920 2285
rect 16880 2275 16885 2280
rect 16695 2255 16885 2275
rect 16695 2250 16700 2255
rect 16660 2245 16700 2250
rect 16880 2250 16885 2255
rect 16915 2275 16920 2280
rect 17100 2280 17140 2285
rect 17100 2275 17105 2280
rect 16915 2255 17105 2275
rect 16915 2250 16920 2255
rect 16880 2245 16920 2250
rect 17100 2250 17105 2255
rect 17135 2275 17140 2280
rect 17320 2280 17360 2285
rect 18055 2280 18095 2285
rect 18165 2285 18170 2290
rect 18200 2310 18205 2315
rect 18275 2315 18315 2320
rect 18275 2310 18280 2315
rect 18200 2290 18280 2310
rect 18200 2285 18205 2290
rect 18165 2280 18205 2285
rect 18275 2285 18280 2290
rect 18310 2310 18315 2315
rect 18385 2315 18425 2320
rect 18385 2310 18390 2315
rect 18310 2290 18390 2310
rect 18310 2285 18315 2290
rect 18275 2280 18315 2285
rect 18385 2285 18390 2290
rect 18420 2310 18425 2315
rect 18495 2315 18535 2320
rect 18495 2310 18500 2315
rect 18420 2290 18500 2310
rect 18420 2285 18425 2290
rect 18385 2280 18425 2285
rect 18495 2285 18500 2290
rect 18530 2310 18535 2315
rect 18695 2315 18735 2320
rect 18695 2310 18700 2315
rect 18530 2290 18700 2310
rect 18530 2285 18535 2290
rect 18495 2280 18535 2285
rect 18695 2285 18700 2290
rect 18730 2285 18735 2315
rect 18695 2280 18735 2285
rect 17320 2275 17325 2280
rect 17135 2255 17325 2275
rect 17135 2250 17140 2255
rect 17100 2245 17140 2250
rect 17320 2250 17325 2255
rect 17355 2250 17360 2280
rect 17320 2245 17360 2250
rect 3805 2240 3810 2245
rect 2460 2220 3810 2240
rect 2460 2215 2465 2220
rect 2425 2210 2465 2215
rect 3805 2215 3810 2220
rect 3840 2215 3845 2245
rect 3805 2210 3845 2215
rect 16330 2235 16370 2240
rect 16330 2205 16335 2235
rect 16365 2230 16370 2235
rect 16550 2235 16590 2240
rect 16550 2230 16555 2235
rect 16365 2210 16555 2230
rect 16365 2205 16370 2210
rect 2330 2200 2370 2205
rect 2330 2170 2335 2200
rect 2365 2195 2370 2200
rect 3265 2200 3305 2205
rect 3265 2195 3270 2200
rect 2365 2175 3270 2195
rect 2365 2170 2370 2175
rect 2330 2165 2370 2170
rect 3265 2170 3270 2175
rect 3300 2195 3305 2200
rect 3985 2200 4025 2205
rect 3985 2195 3990 2200
rect 3300 2175 3990 2195
rect 3300 2170 3305 2175
rect 3265 2165 3305 2170
rect 3985 2170 3990 2175
rect 4020 2195 4025 2200
rect 4705 2200 4745 2205
rect 16330 2200 16370 2205
rect 16550 2205 16555 2210
rect 16585 2230 16590 2235
rect 16770 2235 16810 2240
rect 16770 2230 16775 2235
rect 16585 2210 16775 2230
rect 16585 2205 16590 2210
rect 16550 2200 16590 2205
rect 16770 2205 16775 2210
rect 16805 2230 16810 2235
rect 16990 2235 17030 2240
rect 16990 2230 16995 2235
rect 16805 2210 16995 2230
rect 16805 2205 16810 2210
rect 16770 2200 16810 2205
rect 16990 2205 16995 2210
rect 17025 2230 17030 2235
rect 17210 2235 17250 2240
rect 17210 2230 17215 2235
rect 17025 2210 17215 2230
rect 17025 2205 17030 2210
rect 16990 2200 17030 2205
rect 17210 2205 17215 2210
rect 17245 2230 17250 2235
rect 17430 2235 17470 2240
rect 17430 2230 17435 2235
rect 17245 2210 17435 2230
rect 17245 2205 17250 2210
rect 17210 2200 17250 2205
rect 17430 2205 17435 2210
rect 17465 2205 17470 2235
rect 17430 2200 17470 2205
rect 4705 2195 4710 2200
rect 4020 2175 4710 2195
rect 4020 2170 4025 2175
rect 3985 2165 4025 2170
rect 4705 2170 4710 2175
rect 4740 2170 4745 2200
rect 4705 2165 4745 2170
rect 15950 2180 15990 2185
rect 2380 2150 2420 2155
rect 2380 2120 2385 2150
rect 2415 2145 2420 2150
rect 3625 2150 3665 2155
rect 15950 2150 15955 2180
rect 15985 2175 15990 2180
rect 16828 2180 16862 2185
rect 16828 2175 16831 2180
rect 15985 2155 16831 2175
rect 15985 2150 15990 2155
rect 3625 2145 3630 2150
rect 2415 2125 3630 2145
rect 2415 2120 2420 2125
rect 2380 2115 2420 2120
rect 3625 2120 3630 2125
rect 3660 2120 3665 2150
rect 3625 2115 3665 2120
rect 4085 2145 4125 2150
rect 4085 2115 4090 2145
rect 4120 2140 4125 2145
rect 5315 2145 5355 2150
rect 15950 2145 15990 2150
rect 16828 2150 16831 2155
rect 16859 2150 16862 2180
rect 16828 2145 16862 2150
rect 5315 2140 5320 2145
rect 4120 2120 5320 2140
rect 4120 2115 4125 2120
rect 4085 2110 4125 2115
rect 5315 2115 5320 2120
rect 5350 2115 5355 2145
rect 5315 2110 5355 2115
rect 14510 2110 14560 2120
rect 2745 2095 2785 2100
rect 2745 2065 2750 2095
rect 2780 2090 2785 2095
rect 2865 2095 2905 2100
rect 2865 2090 2870 2095
rect 2780 2070 2870 2090
rect 2780 2065 2785 2070
rect 2745 2060 2785 2065
rect 2865 2065 2870 2070
rect 2900 2090 2905 2095
rect 2985 2095 3025 2100
rect 2985 2090 2990 2095
rect 2900 2070 2990 2090
rect 2900 2065 2905 2070
rect 2865 2060 2905 2065
rect 2985 2065 2990 2070
rect 3020 2090 3025 2095
rect 3105 2095 3145 2100
rect 3105 2090 3110 2095
rect 3020 2070 3110 2090
rect 3020 2065 3025 2070
rect 2985 2060 3025 2065
rect 3105 2065 3110 2070
rect 3140 2090 3145 2095
rect 3225 2095 3265 2100
rect 3225 2090 3230 2095
rect 3140 2070 3230 2090
rect 3140 2065 3145 2070
rect 3105 2060 3145 2065
rect 3225 2065 3230 2070
rect 3260 2090 3265 2095
rect 3345 2095 3385 2100
rect 3345 2090 3350 2095
rect 3260 2070 3350 2090
rect 3260 2065 3265 2070
rect 3225 2060 3265 2065
rect 3345 2065 3350 2070
rect 3380 2090 3385 2095
rect 3465 2095 3505 2100
rect 3465 2090 3470 2095
rect 3380 2070 3470 2090
rect 3380 2065 3385 2070
rect 3345 2060 3385 2065
rect 3465 2065 3470 2070
rect 3500 2090 3505 2095
rect 3585 2095 3625 2100
rect 3585 2090 3590 2095
rect 3500 2070 3590 2090
rect 3500 2065 3505 2070
rect 3465 2060 3505 2065
rect 3585 2065 3590 2070
rect 3620 2090 3625 2095
rect 3705 2095 3745 2100
rect 3705 2090 3710 2095
rect 3620 2070 3710 2090
rect 3620 2065 3625 2070
rect 3585 2060 3625 2065
rect 3705 2065 3710 2070
rect 3740 2090 3745 2095
rect 3825 2095 3865 2100
rect 3825 2090 3830 2095
rect 3740 2070 3830 2090
rect 3740 2065 3745 2070
rect 3705 2060 3745 2065
rect 3825 2065 3830 2070
rect 3860 2090 3865 2095
rect 3985 2095 4025 2100
rect 3985 2090 3990 2095
rect 3860 2070 3990 2090
rect 3860 2065 3865 2070
rect 3825 2060 3865 2065
rect 3985 2065 3990 2070
rect 4020 2090 4025 2095
rect 4145 2095 4185 2100
rect 4145 2090 4150 2095
rect 4020 2070 4150 2090
rect 4020 2065 4025 2070
rect 3985 2060 4025 2065
rect 4145 2065 4150 2070
rect 4180 2090 4185 2095
rect 4265 2095 4305 2100
rect 4265 2090 4270 2095
rect 4180 2070 4270 2090
rect 4180 2065 4185 2070
rect 4145 2060 4185 2065
rect 4265 2065 4270 2070
rect 4300 2090 4305 2095
rect 4385 2095 4425 2100
rect 4385 2090 4390 2095
rect 4300 2070 4390 2090
rect 4300 2065 4305 2070
rect 4265 2060 4305 2065
rect 4385 2065 4390 2070
rect 4420 2090 4425 2095
rect 4505 2095 4545 2100
rect 4505 2090 4510 2095
rect 4420 2070 4510 2090
rect 4420 2065 4425 2070
rect 4385 2060 4425 2065
rect 4505 2065 4510 2070
rect 4540 2090 4545 2095
rect 4625 2095 4665 2100
rect 4625 2090 4630 2095
rect 4540 2070 4630 2090
rect 4540 2065 4545 2070
rect 4505 2060 4545 2065
rect 4625 2065 4630 2070
rect 4660 2090 4665 2095
rect 4745 2095 4785 2100
rect 4745 2090 4750 2095
rect 4660 2070 4750 2090
rect 4660 2065 4665 2070
rect 4625 2060 4665 2065
rect 4745 2065 4750 2070
rect 4780 2090 4785 2095
rect 4865 2095 4905 2100
rect 4865 2090 4870 2095
rect 4780 2070 4870 2090
rect 4780 2065 4785 2070
rect 4745 2060 4785 2065
rect 4865 2065 4870 2070
rect 4900 2090 4905 2095
rect 4985 2095 5025 2100
rect 4985 2090 4990 2095
rect 4900 2070 4990 2090
rect 4900 2065 4905 2070
rect 4865 2060 4905 2065
rect 4985 2065 4990 2070
rect 5020 2090 5025 2095
rect 5105 2095 5145 2100
rect 5105 2090 5110 2095
rect 5020 2070 5110 2090
rect 5020 2065 5025 2070
rect 4985 2060 5025 2065
rect 5105 2065 5110 2070
rect 5140 2090 5145 2095
rect 5225 2095 5265 2100
rect 5225 2090 5230 2095
rect 5140 2070 5230 2090
rect 5140 2065 5145 2070
rect 5105 2060 5145 2065
rect 5225 2065 5230 2070
rect 5260 2090 5265 2095
rect 5550 2095 5590 2100
rect 5550 2090 5555 2095
rect 5260 2070 5555 2090
rect 5260 2065 5265 2070
rect 5225 2060 5265 2065
rect 5550 2065 5555 2070
rect 5585 2065 5590 2095
rect 14510 2080 14520 2110
rect 14550 2080 14560 2110
rect 14510 2070 14560 2080
rect 19240 2110 19290 2120
rect 19240 2080 19250 2110
rect 19280 2080 19290 2110
rect 19240 2070 19290 2080
rect 5550 2060 5590 2065
rect 2620 2050 2660 2055
rect 2620 2020 2625 2050
rect 2655 2020 2660 2050
rect 2620 2015 2660 2020
rect 2805 2050 2845 2055
rect 2805 2020 2810 2050
rect 2840 2045 2845 2050
rect 3165 2050 3205 2055
rect 3165 2045 3170 2050
rect 2840 2025 3170 2045
rect 2840 2020 2845 2025
rect 2805 2015 2845 2020
rect 3165 2020 3170 2025
rect 3200 2045 3205 2050
rect 3525 2050 3565 2055
rect 3525 2045 3530 2050
rect 3200 2025 3530 2045
rect 3200 2020 3205 2025
rect 3165 2015 3205 2020
rect 3525 2020 3530 2025
rect 3560 2045 3565 2050
rect 3885 2050 3925 2055
rect 3885 2045 3890 2050
rect 3560 2025 3890 2045
rect 3560 2020 3565 2025
rect 3525 2015 3565 2020
rect 3885 2020 3890 2025
rect 3920 2020 3925 2050
rect 3885 2015 3925 2020
rect 4085 2050 4125 2055
rect 4085 2020 4090 2050
rect 4120 2045 4125 2050
rect 4445 2050 4485 2055
rect 4445 2045 4450 2050
rect 4120 2025 4450 2045
rect 4120 2020 4125 2025
rect 4085 2015 4125 2020
rect 4445 2020 4450 2025
rect 4480 2045 4485 2050
rect 4805 2050 4845 2055
rect 4805 2045 4810 2050
rect 4480 2025 4810 2045
rect 4480 2020 4485 2025
rect 4445 2015 4485 2020
rect 4805 2020 4810 2025
rect 4840 2045 4845 2050
rect 5165 2050 5205 2055
rect 5165 2045 5170 2050
rect 4840 2025 5170 2045
rect 4840 2020 4845 2025
rect 4805 2015 4845 2020
rect 5165 2020 5170 2025
rect 5200 2020 5205 2050
rect 5165 2015 5205 2020
rect 14790 2010 14825 2011
rect 14790 2005 14885 2010
rect 14825 1970 14850 2005
rect 14790 1965 14885 1970
rect 14910 2005 14945 2011
rect 14910 1965 14945 1970
rect 14970 2005 15005 2010
rect 18795 2005 18830 2010
rect 15020 2000 15060 2005
rect 15020 1995 15025 2000
rect 15005 1975 15025 1995
rect 14970 1965 15005 1970
rect 15020 1970 15025 1975
rect 15055 1970 15060 2000
rect 15020 1965 15060 1970
rect 18740 2000 18780 2005
rect 18740 1970 18745 2000
rect 18775 1995 18780 2000
rect 18775 1975 18795 1995
rect 18775 1970 18780 1975
rect 18740 1965 18780 1970
rect 18795 1965 18830 1970
rect 18855 2005 18890 2011
rect 18975 2010 19010 2011
rect 18855 1965 18890 1970
rect 18915 2005 19010 2010
rect 18950 1970 18975 2005
rect 18915 1965 19010 1970
rect 16385 1960 16425 1965
rect 14910 1945 14950 1950
rect 14910 1915 14915 1945
rect 14945 1940 14950 1945
rect 15065 1945 15105 1950
rect 15065 1940 15070 1945
rect 14945 1920 15070 1940
rect 14945 1915 14950 1920
rect 14910 1910 14950 1915
rect 15065 1915 15070 1920
rect 15100 1915 15105 1945
rect 15065 1910 15105 1915
rect 15210 1945 15250 1950
rect 15210 1915 15215 1945
rect 15245 1940 15250 1945
rect 15320 1945 15360 1950
rect 15320 1940 15325 1945
rect 15245 1920 15325 1940
rect 15245 1915 15250 1920
rect 15210 1910 15250 1915
rect 15320 1915 15325 1920
rect 15355 1940 15360 1945
rect 15430 1945 15470 1950
rect 15430 1940 15435 1945
rect 15355 1920 15435 1940
rect 15355 1915 15360 1920
rect 15320 1910 15360 1915
rect 15430 1915 15435 1920
rect 15465 1940 15470 1945
rect 15540 1945 15580 1950
rect 15540 1940 15545 1945
rect 15465 1920 15545 1940
rect 15465 1915 15470 1920
rect 15430 1910 15470 1915
rect 15540 1915 15545 1920
rect 15575 1940 15580 1945
rect 15650 1945 15690 1950
rect 15650 1940 15655 1945
rect 15575 1920 15655 1940
rect 15575 1915 15580 1920
rect 15540 1910 15580 1915
rect 15650 1915 15655 1920
rect 15685 1940 15690 1945
rect 15760 1945 15800 1950
rect 15760 1940 15765 1945
rect 15685 1920 15765 1940
rect 15685 1915 15690 1920
rect 15650 1910 15690 1915
rect 15760 1915 15765 1920
rect 15795 1915 15800 1945
rect 16385 1930 16390 1960
rect 16420 1955 16425 1960
rect 16605 1960 16645 1965
rect 16605 1955 16610 1960
rect 16420 1935 16610 1955
rect 16420 1930 16425 1935
rect 16385 1925 16425 1930
rect 16605 1930 16610 1935
rect 16640 1955 16645 1960
rect 16825 1960 16865 1965
rect 16825 1955 16830 1960
rect 16640 1935 16830 1955
rect 16640 1930 16645 1935
rect 16605 1925 16645 1930
rect 16825 1930 16830 1935
rect 16860 1955 16865 1960
rect 17045 1960 17085 1965
rect 17045 1955 17050 1960
rect 16860 1935 17050 1955
rect 16860 1930 16865 1935
rect 16825 1925 16865 1930
rect 17045 1930 17050 1935
rect 17080 1955 17085 1960
rect 17265 1960 17305 1965
rect 17265 1955 17270 1960
rect 17080 1935 17270 1955
rect 17080 1930 17085 1935
rect 17045 1925 17085 1930
rect 17265 1930 17270 1935
rect 17300 1930 17305 1960
rect 17265 1925 17305 1930
rect 18000 1945 18040 1950
rect 15760 1910 15800 1915
rect 18000 1915 18005 1945
rect 18035 1940 18040 1945
rect 18110 1945 18150 1950
rect 18110 1940 18115 1945
rect 18035 1920 18115 1940
rect 18035 1915 18040 1920
rect 18000 1910 18040 1915
rect 18110 1915 18115 1920
rect 18145 1940 18150 1945
rect 18220 1945 18260 1950
rect 18220 1940 18225 1945
rect 18145 1920 18225 1940
rect 18145 1915 18150 1920
rect 18110 1910 18150 1915
rect 18220 1915 18225 1920
rect 18255 1940 18260 1945
rect 18330 1945 18370 1950
rect 18330 1940 18335 1945
rect 18255 1920 18335 1940
rect 18255 1915 18260 1920
rect 18220 1910 18260 1915
rect 18330 1915 18335 1920
rect 18365 1940 18370 1945
rect 18440 1945 18480 1950
rect 18440 1940 18445 1945
rect 18365 1920 18445 1940
rect 18365 1915 18370 1920
rect 18330 1910 18370 1915
rect 18440 1915 18445 1920
rect 18475 1940 18480 1945
rect 18550 1945 18590 1950
rect 18550 1940 18555 1945
rect 18475 1920 18555 1940
rect 18475 1915 18480 1920
rect 18440 1910 18480 1915
rect 18550 1915 18555 1920
rect 18585 1915 18590 1945
rect 18550 1910 18590 1915
rect 18695 1945 18735 1950
rect 18695 1915 18700 1945
rect 18730 1940 18735 1945
rect 18850 1945 18890 1950
rect 18850 1940 18855 1945
rect 18730 1920 18855 1940
rect 18730 1915 18735 1920
rect 18695 1910 18735 1915
rect 18850 1915 18855 1920
rect 18885 1915 18890 1945
rect 18850 1910 18890 1915
rect 16495 1905 16535 1910
rect 14790 1895 14830 1900
rect 2925 1880 2965 1885
rect 2925 1850 2930 1880
rect 2960 1875 2965 1880
rect 3045 1875 3085 1885
rect 3285 1880 3325 1885
rect 3285 1875 3290 1880
rect 2960 1855 3290 1875
rect 2960 1850 2965 1855
rect 2925 1845 2965 1850
rect 3045 1845 3085 1855
rect 3285 1850 3290 1855
rect 3320 1875 3325 1880
rect 3405 1875 3445 1885
rect 3645 1880 3685 1885
rect 3645 1875 3650 1880
rect 3320 1855 3650 1875
rect 3320 1850 3325 1855
rect 3285 1845 3325 1850
rect 3405 1845 3445 1855
rect 3645 1850 3650 1855
rect 3680 1850 3685 1880
rect 3645 1845 3685 1850
rect 3765 1845 3805 1885
rect 4205 1845 4245 1885
rect 4325 1880 4365 1885
rect 4325 1850 4330 1880
rect 4360 1875 4365 1880
rect 4565 1875 4605 1885
rect 4685 1880 4725 1885
rect 4685 1875 4690 1880
rect 4360 1855 4690 1875
rect 4360 1850 4365 1855
rect 4325 1845 4365 1850
rect 4565 1845 4605 1855
rect 4685 1850 4690 1855
rect 4720 1875 4725 1880
rect 4925 1875 4965 1885
rect 5045 1880 5085 1885
rect 5045 1875 5050 1880
rect 4720 1855 5050 1875
rect 4720 1850 4725 1855
rect 4685 1845 4725 1850
rect 4925 1845 4965 1855
rect 5045 1850 5050 1855
rect 5080 1875 5085 1880
rect 5080 1855 5175 1875
rect 14790 1865 14795 1895
rect 14825 1890 14830 1895
rect 16000 1895 16040 1900
rect 16000 1890 16005 1895
rect 14825 1870 16005 1890
rect 14825 1865 14830 1870
rect 14790 1860 14830 1865
rect 16000 1865 16005 1870
rect 16035 1865 16040 1895
rect 16495 1875 16500 1905
rect 16530 1900 16535 1905
rect 16715 1905 16755 1910
rect 16715 1900 16720 1905
rect 16530 1880 16720 1900
rect 16530 1875 16535 1880
rect 16495 1870 16535 1875
rect 16715 1875 16720 1880
rect 16750 1900 16755 1905
rect 16935 1905 16975 1910
rect 16935 1900 16940 1905
rect 16750 1880 16940 1900
rect 16750 1875 16755 1880
rect 16715 1870 16755 1875
rect 16935 1875 16940 1880
rect 16970 1900 16975 1905
rect 17155 1905 17195 1910
rect 17155 1900 17160 1905
rect 16970 1880 17160 1900
rect 16970 1875 16975 1880
rect 16935 1870 16975 1875
rect 17155 1875 17160 1880
rect 17190 1900 17195 1905
rect 17375 1905 17415 1910
rect 17375 1900 17380 1905
rect 17190 1880 17380 1900
rect 17190 1875 17195 1880
rect 17155 1870 17195 1875
rect 17375 1875 17380 1880
rect 17410 1875 17415 1905
rect 17375 1870 17415 1875
rect 17760 1895 17800 1900
rect 16000 1860 16040 1865
rect 17760 1865 17765 1895
rect 17795 1890 17800 1895
rect 18970 1895 19010 1900
rect 18970 1890 18975 1895
rect 17795 1870 18975 1890
rect 17795 1865 17800 1870
rect 17760 1860 17800 1865
rect 18970 1865 18975 1870
rect 19005 1865 19010 1895
rect 18970 1860 19010 1865
rect 5080 1850 5085 1855
rect 5045 1845 5085 1850
rect 16190 1850 16230 1855
rect 2470 1820 2510 1825
rect 2470 1790 2475 1820
rect 2505 1815 2510 1820
rect 2835 1820 2875 1825
rect 2835 1815 2840 1820
rect 2505 1795 2840 1815
rect 2505 1790 2510 1795
rect 2470 1785 2510 1790
rect 2835 1790 2840 1795
rect 2870 1815 2875 1820
rect 3045 1820 3085 1825
rect 3045 1815 3050 1820
rect 2870 1795 3050 1815
rect 2870 1790 2875 1795
rect 2835 1785 2875 1790
rect 3045 1790 3050 1795
rect 3080 1815 3085 1820
rect 3165 1820 3205 1825
rect 3165 1815 3170 1820
rect 3080 1795 3170 1815
rect 3080 1790 3085 1795
rect 3045 1785 3085 1790
rect 3165 1790 3170 1795
rect 3200 1815 3205 1820
rect 3405 1820 3445 1825
rect 3405 1815 3410 1820
rect 3200 1795 3410 1815
rect 3200 1790 3205 1795
rect 3165 1785 3205 1790
rect 3405 1790 3410 1795
rect 3440 1815 3445 1820
rect 3525 1820 3565 1825
rect 3525 1815 3530 1820
rect 3440 1795 3530 1815
rect 3440 1790 3445 1795
rect 3405 1785 3445 1790
rect 3525 1790 3530 1795
rect 3560 1815 3565 1820
rect 3765 1820 3805 1825
rect 3765 1815 3770 1820
rect 3560 1795 3770 1815
rect 3560 1790 3565 1795
rect 3525 1785 3565 1790
rect 3765 1790 3770 1795
rect 3800 1815 3805 1820
rect 3855 1820 3895 1825
rect 3855 1815 3860 1820
rect 3800 1795 3860 1815
rect 3800 1790 3805 1795
rect 3765 1785 3805 1790
rect 3855 1790 3860 1795
rect 3890 1790 3895 1820
rect 3855 1785 3895 1790
rect 4115 1820 4155 1825
rect 4115 1790 4120 1820
rect 4150 1815 4155 1820
rect 4205 1820 4245 1825
rect 4205 1815 4210 1820
rect 4150 1795 4210 1815
rect 4150 1790 4155 1795
rect 4115 1785 4155 1790
rect 4205 1790 4210 1795
rect 4240 1815 4245 1820
rect 4445 1820 4485 1825
rect 4445 1815 4450 1820
rect 4240 1795 4450 1815
rect 4240 1790 4245 1795
rect 4205 1785 4245 1790
rect 4445 1790 4450 1795
rect 4480 1815 4485 1820
rect 4565 1820 4605 1825
rect 4565 1815 4570 1820
rect 4480 1795 4570 1815
rect 4480 1790 4485 1795
rect 4445 1785 4485 1790
rect 4565 1790 4570 1795
rect 4600 1815 4605 1820
rect 4805 1820 4845 1825
rect 4805 1815 4810 1820
rect 4600 1795 4810 1815
rect 4600 1790 4605 1795
rect 4565 1785 4605 1790
rect 4805 1790 4810 1795
rect 4840 1815 4845 1820
rect 4925 1820 4965 1825
rect 4925 1815 4930 1820
rect 4840 1795 4930 1815
rect 4840 1790 4845 1795
rect 4805 1785 4845 1790
rect 4925 1790 4930 1795
rect 4960 1815 4965 1820
rect 5135 1820 5175 1825
rect 5135 1815 5140 1820
rect 4960 1795 5140 1815
rect 4960 1790 4965 1795
rect 4925 1785 4965 1790
rect 5135 1790 5140 1795
rect 5170 1815 5175 1820
rect 5360 1820 5400 1825
rect 5360 1815 5365 1820
rect 5170 1795 5365 1815
rect 5170 1790 5175 1795
rect 5135 1785 5175 1790
rect 5360 1790 5365 1795
rect 5395 1790 5400 1820
rect 16190 1820 16195 1850
rect 16225 1845 16230 1850
rect 16410 1850 16450 1855
rect 16410 1845 16415 1850
rect 16225 1825 16415 1845
rect 16225 1820 16230 1825
rect 16190 1815 16230 1820
rect 16410 1820 16415 1825
rect 16445 1845 16450 1850
rect 16640 1850 16680 1855
rect 16640 1845 16645 1850
rect 16445 1825 16645 1845
rect 16445 1820 16450 1825
rect 16410 1815 16450 1820
rect 16640 1820 16645 1825
rect 16675 1845 16680 1850
rect 17230 1850 17270 1855
rect 17230 1845 17235 1850
rect 16675 1825 17235 1845
rect 16675 1820 16680 1825
rect 16640 1815 16680 1820
rect 17230 1820 17235 1825
rect 17265 1845 17270 1850
rect 17450 1850 17490 1855
rect 17450 1845 17455 1850
rect 17265 1825 17455 1845
rect 17265 1820 17270 1825
rect 17230 1815 17270 1820
rect 17450 1820 17455 1825
rect 17485 1845 17490 1850
rect 17680 1850 17720 1855
rect 17680 1845 17685 1850
rect 17485 1825 17685 1845
rect 17485 1820 17490 1825
rect 17450 1815 17490 1820
rect 17680 1820 17685 1825
rect 17715 1820 17720 1850
rect 17680 1815 17720 1820
rect 5360 1785 5400 1790
rect 16820 1805 16860 1810
rect 16820 1775 16825 1805
rect 16855 1800 16860 1805
rect 16940 1805 16980 1810
rect 16940 1800 16945 1805
rect 16855 1780 16945 1800
rect 16855 1775 16860 1780
rect 16820 1770 16860 1775
rect 16940 1775 16945 1780
rect 16975 1775 16980 1805
rect 16940 1770 16980 1775
rect 2800 1765 2840 1770
rect 2425 1760 2465 1765
rect 2425 1730 2430 1760
rect 2460 1755 2465 1760
rect 2565 1760 2605 1765
rect 2565 1755 2570 1760
rect 2460 1735 2570 1755
rect 2460 1730 2465 1735
rect 2425 1725 2465 1730
rect 2565 1730 2570 1735
rect 2600 1755 2605 1760
rect 2675 1760 2715 1765
rect 2675 1755 2680 1760
rect 2600 1735 2680 1755
rect 2600 1730 2605 1735
rect 2565 1725 2605 1730
rect 2675 1730 2680 1735
rect 2710 1755 2715 1760
rect 2800 1755 2805 1765
rect 2710 1735 2805 1755
rect 2835 1755 2840 1765
rect 3225 1760 3265 1765
rect 3225 1755 3230 1760
rect 2835 1735 3230 1755
rect 2710 1730 2715 1735
rect 2800 1730 2840 1735
rect 3225 1730 3230 1735
rect 3260 1730 3265 1760
rect 2675 1725 2715 1730
rect 3225 1725 3265 1730
rect 3285 1760 3325 1765
rect 3285 1730 3290 1760
rect 3320 1755 3325 1760
rect 3525 1760 3565 1765
rect 3525 1755 3530 1760
rect 3320 1735 3530 1755
rect 3320 1730 3325 1735
rect 3285 1725 3325 1730
rect 3525 1730 3530 1735
rect 3560 1755 3565 1760
rect 3765 1760 3805 1765
rect 3765 1755 3770 1760
rect 3560 1735 3770 1755
rect 3560 1730 3565 1735
rect 3525 1725 3565 1730
rect 3765 1730 3770 1735
rect 3800 1730 3805 1760
rect 3765 1725 3805 1730
rect 4205 1760 4245 1765
rect 4205 1730 4210 1760
rect 4240 1755 4245 1760
rect 4445 1760 4485 1765
rect 4445 1755 4450 1760
rect 4240 1735 4450 1755
rect 4240 1730 4245 1735
rect 4205 1725 4245 1730
rect 4445 1730 4450 1735
rect 4480 1755 4485 1760
rect 4685 1760 4725 1765
rect 4685 1755 4690 1760
rect 4480 1735 4690 1755
rect 4480 1730 4485 1735
rect 4445 1725 4485 1730
rect 4685 1730 4690 1735
rect 4720 1730 4725 1760
rect 4685 1725 4725 1730
rect 4745 1760 4785 1765
rect 4745 1730 4750 1760
rect 4780 1755 4785 1760
rect 5270 1760 5310 1765
rect 5270 1755 5275 1760
rect 4780 1735 5275 1755
rect 4780 1730 4785 1735
rect 4745 1725 4785 1730
rect 5270 1730 5275 1735
rect 5305 1755 5310 1760
rect 14965 1760 15005 1765
rect 5305 1735 6100 1755
rect 5305 1730 5310 1735
rect 5270 1725 5310 1730
rect 14965 1730 14970 1760
rect 15000 1755 15005 1760
rect 15555 1760 15595 1765
rect 15555 1755 15560 1760
rect 15000 1735 15560 1755
rect 15000 1730 15005 1735
rect 14965 1725 15005 1730
rect 15555 1730 15560 1735
rect 15590 1755 15595 1760
rect 15835 1760 15875 1765
rect 15835 1755 15840 1760
rect 15590 1735 15840 1755
rect 15590 1730 15595 1735
rect 15555 1725 15595 1730
rect 15835 1730 15840 1735
rect 15870 1730 15875 1760
rect 15835 1725 15875 1730
rect 16085 1760 16125 1765
rect 16085 1730 16090 1760
rect 16120 1755 16125 1760
rect 16305 1760 16345 1765
rect 16305 1755 16310 1760
rect 16120 1735 16310 1755
rect 16120 1730 16125 1735
rect 16085 1725 16125 1730
rect 16305 1730 16310 1735
rect 16340 1755 16345 1760
rect 16525 1760 16565 1765
rect 16525 1755 16530 1760
rect 16340 1735 16530 1755
rect 16340 1730 16345 1735
rect 16305 1725 16345 1730
rect 16525 1730 16530 1735
rect 16560 1755 16565 1760
rect 17125 1760 17165 1765
rect 17125 1755 17130 1760
rect 16560 1735 17130 1755
rect 16560 1730 16565 1735
rect 16525 1725 16565 1730
rect 17125 1730 17130 1735
rect 17160 1755 17165 1760
rect 17345 1760 17385 1765
rect 17345 1755 17350 1760
rect 17160 1735 17350 1755
rect 17160 1730 17165 1735
rect 17125 1725 17165 1730
rect 17345 1730 17350 1735
rect 17380 1755 17385 1760
rect 17565 1760 17605 1765
rect 17565 1755 17570 1760
rect 17380 1735 17570 1755
rect 17380 1730 17385 1735
rect 17345 1725 17385 1730
rect 17565 1730 17570 1735
rect 17600 1730 17605 1760
rect 17565 1725 17605 1730
rect 17925 1760 17965 1765
rect 17925 1730 17930 1760
rect 17960 1755 17965 1760
rect 18205 1760 18245 1765
rect 18205 1755 18210 1760
rect 17960 1735 18210 1755
rect 17960 1730 17965 1735
rect 17925 1725 17965 1730
rect 18205 1730 18210 1735
rect 18240 1755 18245 1760
rect 18795 1760 18835 1765
rect 18795 1755 18800 1760
rect 18240 1735 18800 1755
rect 18240 1730 18245 1735
rect 18205 1725 18245 1730
rect 18795 1730 18800 1735
rect 18830 1730 18835 1760
rect 18795 1725 18835 1730
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 1685 -70 1690
rect -45 1720 -5 1725
rect -45 1690 -40 1720
rect -10 1690 -5 1720
rect 3165 1715 3205 1720
rect -45 1685 -5 1690
rect 1262 1710 1302 1715
rect 1262 1680 1270 1710
rect 1297 1705 1302 1710
rect 2800 1710 2840 1715
rect 2800 1705 2805 1710
rect 1297 1685 2805 1705
rect 1297 1680 1302 1685
rect 1262 1675 1302 1680
rect 2800 1680 2805 1685
rect 2835 1680 2840 1710
rect 3165 1685 3170 1715
rect 3200 1710 3205 1715
rect 3405 1715 3445 1720
rect 3405 1710 3410 1715
rect 3200 1690 3410 1710
rect 3200 1685 3205 1690
rect 3165 1680 3205 1685
rect 3405 1685 3410 1690
rect 3440 1710 3445 1715
rect 3645 1715 3685 1720
rect 3645 1710 3650 1715
rect 3440 1690 3650 1710
rect 3440 1685 3445 1690
rect 3405 1680 3445 1685
rect 3645 1685 3650 1690
rect 3680 1685 3685 1715
rect 3645 1680 3685 1685
rect 4325 1715 4365 1720
rect 4325 1685 4330 1715
rect 4360 1710 4365 1715
rect 4565 1715 4605 1720
rect 4565 1710 4570 1715
rect 4360 1690 4570 1710
rect 4360 1685 4365 1690
rect 4325 1680 4365 1685
rect 4565 1685 4570 1690
rect 4600 1710 4605 1715
rect 4805 1715 4845 1720
rect 4805 1710 4810 1715
rect 4600 1690 4810 1710
rect 4600 1685 4605 1690
rect 4565 1680 4605 1685
rect 4805 1685 4810 1690
rect 4840 1685 4845 1715
rect 16237 1715 16269 1720
rect 16237 1710 16240 1715
rect 4805 1680 4845 1685
rect 14515 1705 14555 1710
rect 2800 1675 2840 1680
rect 14515 1675 14520 1705
rect 14550 1700 14555 1705
rect 15030 1705 15070 1710
rect 15030 1700 15035 1705
rect 14550 1680 15035 1700
rect 14550 1675 14555 1680
rect 14515 1670 14555 1675
rect 15030 1675 15035 1680
rect 15065 1700 15070 1705
rect 15255 1705 15295 1710
rect 15255 1700 15260 1705
rect 15065 1680 15260 1700
rect 15065 1675 15070 1680
rect 15030 1670 15070 1675
rect 15255 1675 15260 1680
rect 15290 1700 15295 1705
rect 15455 1705 15495 1710
rect 15455 1700 15460 1705
rect 15290 1680 15460 1700
rect 15290 1675 15295 1680
rect 15255 1670 15295 1675
rect 15455 1675 15460 1680
rect 15490 1700 15495 1705
rect 15655 1705 15695 1710
rect 15655 1700 15660 1705
rect 15490 1680 15660 1700
rect 15490 1675 15495 1680
rect 15455 1670 15495 1675
rect 15655 1675 15660 1680
rect 15690 1675 15695 1705
rect 15910 1690 16240 1710
rect 16237 1685 16240 1690
rect 16266 1710 16269 1715
rect 16457 1715 16489 1720
rect 16457 1710 16460 1715
rect 16266 1690 16460 1710
rect 16266 1685 16269 1690
rect 16237 1680 16269 1685
rect 16457 1685 16460 1690
rect 16486 1710 16489 1715
rect 16601 1715 16633 1720
rect 16601 1710 16604 1715
rect 16486 1690 16604 1710
rect 16486 1685 16489 1690
rect 16457 1680 16489 1685
rect 16601 1685 16604 1690
rect 16630 1710 16633 1715
rect 16867 1715 16899 1720
rect 16867 1710 16870 1715
rect 16630 1690 16870 1710
rect 16630 1685 16633 1690
rect 16601 1680 16633 1685
rect 16867 1685 16870 1690
rect 16896 1710 16899 1715
rect 17277 1715 17309 1720
rect 17277 1710 17280 1715
rect 16896 1690 17280 1710
rect 16896 1685 16899 1690
rect 16867 1680 16899 1685
rect 17277 1685 17280 1690
rect 17306 1710 17309 1715
rect 17497 1715 17529 1720
rect 17497 1710 17500 1715
rect 17306 1690 17500 1710
rect 17306 1685 17309 1690
rect 17277 1680 17309 1685
rect 17497 1685 17500 1690
rect 17526 1710 17529 1715
rect 17641 1715 17673 1720
rect 17641 1710 17644 1715
rect 17526 1690 17644 1710
rect 17526 1685 17529 1690
rect 17497 1680 17529 1685
rect 17641 1685 17644 1690
rect 17670 1685 17673 1715
rect 17641 1680 17673 1685
rect 18105 1705 18145 1710
rect 15655 1670 15695 1675
rect 18105 1675 18110 1705
rect 18140 1700 18145 1705
rect 18305 1705 18345 1710
rect 18305 1700 18310 1705
rect 18140 1680 18310 1700
rect 18140 1675 18145 1680
rect 18105 1670 18145 1675
rect 18305 1675 18310 1680
rect 18340 1700 18345 1705
rect 18505 1705 18545 1710
rect 18505 1700 18510 1705
rect 18340 1680 18510 1700
rect 18340 1675 18345 1680
rect 18305 1670 18345 1675
rect 18505 1675 18510 1680
rect 18540 1700 18545 1705
rect 18730 1705 18770 1710
rect 18730 1700 18735 1705
rect 18540 1680 18735 1700
rect 18540 1675 18545 1680
rect 18505 1670 18545 1675
rect 18730 1675 18735 1680
rect 18765 1700 18770 1705
rect 19245 1705 19285 1710
rect 19245 1700 19250 1705
rect 18765 1680 19250 1700
rect 18765 1675 18770 1680
rect 18730 1670 18770 1675
rect 19245 1675 19250 1680
rect 19280 1675 19285 1705
rect 19245 1670 19285 1675
rect 2380 1665 2420 1670
rect 2380 1635 2385 1665
rect 2415 1660 2420 1665
rect 2620 1665 2660 1670
rect 2620 1660 2625 1665
rect 2415 1640 2625 1660
rect 2415 1635 2420 1640
rect 2380 1630 2420 1635
rect 2620 1635 2625 1640
rect 2655 1635 2660 1665
rect 2620 1630 2660 1635
rect 14970 1645 15005 1650
rect 14970 1605 15005 1610
rect 15030 1645 15065 1650
rect 15030 1605 15065 1610
rect 18735 1645 18770 1650
rect 18735 1605 18770 1610
rect 18795 1645 18830 1650
rect 18795 1605 18830 1610
rect 2330 1595 2370 1600
rect 2330 1565 2335 1595
rect 2365 1590 2370 1595
rect 3165 1595 3205 1600
rect 3165 1590 3170 1595
rect 2365 1570 3170 1590
rect 2365 1565 2370 1570
rect 2330 1560 2370 1565
rect 3165 1565 3170 1570
rect 3200 1565 3205 1595
rect 3165 1560 3205 1565
rect 4805 1595 4845 1600
rect 4805 1565 4810 1595
rect 4840 1590 4845 1595
rect 5410 1595 5450 1600
rect 5410 1590 5415 1595
rect 4840 1570 5415 1590
rect 4840 1565 4845 1570
rect 4805 1560 4845 1565
rect 5410 1565 5415 1570
rect 5445 1565 5450 1595
rect 5410 1560 5450 1565
rect 2835 1545 2875 1550
rect 2835 1515 2840 1545
rect 2870 1540 2875 1545
rect 3225 1545 3265 1550
rect 3225 1540 3230 1545
rect 2870 1520 3230 1540
rect 2870 1515 2875 1520
rect 2835 1510 2875 1515
rect 3225 1515 3230 1520
rect 3260 1540 3265 1545
rect 3345 1545 3385 1550
rect 3345 1540 3350 1545
rect 3260 1520 3350 1540
rect 3260 1515 3265 1520
rect 3225 1510 3265 1515
rect 3345 1515 3350 1520
rect 3380 1540 3385 1545
rect 3465 1545 3505 1550
rect 3465 1540 3470 1545
rect 3380 1520 3470 1540
rect 3380 1515 3385 1520
rect 3345 1510 3385 1515
rect 3465 1515 3470 1520
rect 3500 1540 3505 1545
rect 3585 1545 3625 1550
rect 3585 1540 3590 1545
rect 3500 1520 3590 1540
rect 3500 1515 3505 1520
rect 3465 1510 3505 1515
rect 3585 1515 3590 1520
rect 3620 1540 3625 1545
rect 3705 1545 3745 1550
rect 3705 1540 3710 1545
rect 3620 1520 3710 1540
rect 3620 1515 3625 1520
rect 3585 1510 3625 1515
rect 3705 1515 3710 1520
rect 3740 1515 3745 1545
rect 3705 1510 3745 1515
rect 4265 1545 4305 1550
rect 4265 1515 4270 1545
rect 4300 1540 4305 1545
rect 4385 1545 4425 1550
rect 4385 1540 4390 1545
rect 4300 1520 4390 1540
rect 4300 1515 4305 1520
rect 4265 1510 4305 1515
rect 4385 1515 4390 1520
rect 4420 1540 4425 1545
rect 4505 1545 4545 1550
rect 4505 1540 4510 1545
rect 4420 1520 4510 1540
rect 4420 1515 4425 1520
rect 4385 1510 4425 1515
rect 4505 1515 4510 1520
rect 4540 1540 4545 1545
rect 4625 1545 4665 1550
rect 4625 1540 4630 1545
rect 4540 1520 4630 1540
rect 4540 1515 4545 1520
rect 4505 1510 4545 1515
rect 4625 1515 4630 1520
rect 4660 1540 4665 1545
rect 4745 1545 4785 1550
rect 4745 1540 4750 1545
rect 4660 1520 4750 1540
rect 4660 1515 4665 1520
rect 4625 1510 4665 1515
rect 4745 1515 4750 1520
rect 4780 1540 4785 1545
rect 5135 1545 5175 1550
rect 5135 1540 5140 1545
rect 4780 1520 5140 1540
rect 4780 1515 4785 1520
rect 4745 1510 4785 1515
rect 5135 1515 5140 1520
rect 5170 1515 5175 1545
rect 5135 1510 5175 1515
rect 2925 1500 2965 1505
rect 2925 1470 2930 1500
rect 2960 1495 2965 1500
rect 3045 1500 3085 1505
rect 3045 1495 3050 1500
rect 2960 1475 3050 1495
rect 2960 1470 2965 1475
rect 2925 1465 2965 1470
rect 3045 1470 3050 1475
rect 3080 1495 3085 1500
rect 3165 1500 3205 1505
rect 3165 1495 3170 1500
rect 3080 1475 3170 1495
rect 3080 1470 3085 1475
rect 3045 1465 3085 1470
rect 3165 1470 3170 1475
rect 3200 1495 3205 1500
rect 3285 1500 3325 1505
rect 3285 1495 3290 1500
rect 3200 1475 3290 1495
rect 3200 1470 3205 1475
rect 3165 1465 3205 1470
rect 3285 1470 3290 1475
rect 3320 1495 3325 1500
rect 3525 1500 3565 1505
rect 3525 1495 3530 1500
rect 3320 1475 3530 1495
rect 3320 1470 3325 1475
rect 3285 1465 3325 1470
rect 3525 1470 3530 1475
rect 3560 1495 3565 1500
rect 3645 1500 3685 1505
rect 3645 1495 3650 1500
rect 3560 1475 3650 1495
rect 3560 1470 3565 1475
rect 3525 1465 3565 1470
rect 3645 1470 3650 1475
rect 3680 1495 3685 1500
rect 3765 1500 3805 1505
rect 3765 1495 3770 1500
rect 3680 1475 3770 1495
rect 3680 1470 3685 1475
rect 3645 1465 3685 1470
rect 3765 1470 3770 1475
rect 3800 1495 3805 1500
rect 4205 1500 4245 1505
rect 4205 1495 4210 1500
rect 3800 1475 4210 1495
rect 3800 1470 3805 1475
rect 3765 1465 3805 1470
rect 4205 1470 4210 1475
rect 4240 1495 4245 1500
rect 4325 1500 4365 1505
rect 4325 1495 4330 1500
rect 4240 1475 4330 1495
rect 4240 1470 4245 1475
rect 4205 1465 4245 1470
rect 4325 1470 4330 1475
rect 4360 1495 4365 1500
rect 4445 1500 4485 1505
rect 4445 1495 4450 1500
rect 4360 1475 4450 1495
rect 4360 1470 4365 1475
rect 4325 1465 4365 1470
rect 4445 1470 4450 1475
rect 4480 1495 4485 1500
rect 4685 1500 4725 1505
rect 4685 1495 4690 1500
rect 4480 1475 4690 1495
rect 4480 1470 4485 1475
rect 4445 1465 4485 1470
rect 4685 1470 4690 1475
rect 4720 1495 4725 1500
rect 4805 1500 4845 1505
rect 4805 1495 4810 1500
rect 4720 1475 4810 1495
rect 4720 1470 4725 1475
rect 4685 1465 4725 1470
rect 4805 1470 4810 1475
rect 4840 1495 4845 1500
rect 4925 1500 4965 1505
rect 4925 1495 4930 1500
rect 4840 1475 4930 1495
rect 4840 1470 4845 1475
rect 4805 1465 4845 1470
rect 4925 1470 4930 1475
rect 4960 1495 4965 1500
rect 5045 1500 5085 1505
rect 5045 1495 5050 1500
rect 4960 1475 5050 1495
rect 4960 1470 4965 1475
rect 4925 1465 4965 1470
rect 5045 1470 5050 1475
rect 5080 1495 5085 1500
rect 5550 1500 5590 1505
rect 5550 1495 5555 1500
rect 5080 1475 5555 1495
rect 5080 1470 5085 1475
rect 5045 1465 5085 1470
rect 5550 1470 5555 1475
rect 5585 1470 5590 1500
rect 16106 1495 16138 1500
rect 16106 1490 16109 1495
rect 15905 1470 16109 1490
rect 5550 1465 5590 1470
rect 16106 1465 16109 1470
rect 16135 1490 16138 1495
rect 16305 1495 16345 1500
rect 16305 1490 16310 1495
rect 16135 1470 16310 1490
rect 16135 1465 16138 1470
rect 16106 1460 16138 1465
rect 16305 1465 16310 1470
rect 16340 1490 16345 1495
rect 16525 1495 16565 1500
rect 16525 1490 16530 1495
rect 16340 1470 16530 1490
rect 16340 1465 16345 1470
rect 16305 1460 16345 1465
rect 16525 1465 16530 1470
rect 16560 1490 16565 1495
rect 16922 1495 16954 1500
rect 16922 1490 16925 1495
rect 16560 1470 16925 1490
rect 16560 1465 16565 1470
rect 16525 1460 16565 1465
rect 16922 1465 16925 1470
rect 16951 1490 16954 1495
rect 17146 1495 17178 1500
rect 17146 1490 17149 1495
rect 16951 1470 17149 1490
rect 16951 1465 16954 1470
rect 16922 1460 16954 1465
rect 17146 1465 17149 1470
rect 17175 1490 17178 1495
rect 17345 1495 17385 1500
rect 17345 1490 17350 1495
rect 17175 1470 17350 1490
rect 17175 1465 17178 1470
rect 17146 1460 17178 1465
rect 17345 1465 17350 1470
rect 17380 1490 17385 1495
rect 17565 1495 17605 1500
rect 17565 1490 17570 1495
rect 17380 1470 17570 1490
rect 17380 1465 17385 1470
rect 17345 1460 17385 1465
rect 17565 1465 17570 1470
rect 17600 1465 17605 1495
rect 17565 1460 17605 1465
rect 16145 1435 16185 1440
rect 16145 1405 16150 1435
rect 16180 1430 16185 1435
rect 16250 1435 16290 1440
rect 16250 1430 16255 1435
rect 16180 1410 16255 1430
rect 16180 1405 16185 1410
rect 16145 1400 16185 1405
rect 16250 1405 16255 1410
rect 16285 1430 16290 1435
rect 16360 1435 16400 1440
rect 16360 1430 16365 1435
rect 16285 1410 16365 1430
rect 16285 1405 16290 1410
rect 16250 1400 16290 1405
rect 16360 1405 16365 1410
rect 16395 1430 16400 1435
rect 16470 1435 16510 1440
rect 16470 1430 16475 1435
rect 16395 1410 16475 1430
rect 16395 1405 16400 1410
rect 16360 1400 16400 1405
rect 16470 1405 16475 1410
rect 16505 1430 16510 1435
rect 16580 1435 16620 1440
rect 16580 1430 16585 1435
rect 16505 1410 16585 1430
rect 16505 1405 16510 1410
rect 16470 1400 16510 1405
rect 16580 1405 16585 1410
rect 16615 1430 16620 1435
rect 17185 1435 17225 1440
rect 17185 1430 17190 1435
rect 16615 1410 17190 1430
rect 16615 1405 16620 1410
rect 16580 1400 16620 1405
rect 17185 1405 17190 1410
rect 17220 1430 17225 1435
rect 17290 1435 17330 1440
rect 17290 1430 17295 1435
rect 17220 1410 17295 1430
rect 17220 1405 17225 1410
rect 17185 1400 17225 1405
rect 17290 1405 17295 1410
rect 17325 1430 17330 1435
rect 17400 1435 17440 1440
rect 17400 1430 17405 1435
rect 17325 1410 17405 1430
rect 17325 1405 17330 1410
rect 17290 1400 17330 1405
rect 17400 1405 17405 1410
rect 17435 1430 17440 1435
rect 17510 1435 17550 1440
rect 17510 1430 17515 1435
rect 17435 1410 17515 1430
rect 17435 1405 17440 1410
rect 17400 1400 17440 1405
rect 17510 1405 17515 1410
rect 17545 1430 17550 1435
rect 17620 1435 17660 1440
rect 17620 1430 17625 1435
rect 17545 1410 17625 1430
rect 17545 1405 17550 1410
rect 17510 1400 17550 1405
rect 17620 1405 17625 1410
rect 17655 1405 17660 1435
rect 17620 1400 17660 1405
rect 15835 1390 15875 1395
rect 15835 1360 15840 1390
rect 15870 1385 15875 1390
rect 17925 1390 17965 1395
rect 17925 1385 17930 1390
rect 15870 1365 17930 1385
rect 15870 1360 15875 1365
rect 15835 1355 15875 1360
rect 17925 1360 17930 1365
rect 17960 1360 17965 1390
rect 17925 1355 17965 1360
rect 16005 1345 16045 1350
rect 16005 1315 16010 1345
rect 16040 1340 16045 1345
rect 16810 1345 16850 1350
rect 16810 1340 16815 1345
rect 16040 1320 16815 1340
rect 16040 1315 16045 1320
rect 16005 1310 16045 1315
rect 16810 1315 16815 1320
rect 16845 1315 16850 1345
rect 16810 1310 16850 1315
rect 16315 1295 16355 1300
rect 16315 1265 16320 1295
rect 16350 1290 16355 1295
rect 16880 1295 16920 1300
rect 16880 1290 16885 1295
rect 16350 1270 16885 1290
rect 16350 1265 16355 1270
rect 16315 1260 16355 1265
rect 16880 1265 16885 1270
rect 16915 1265 16920 1295
rect 16880 1260 16920 1265
rect 17595 1250 17635 1255
rect 16425 1235 16465 1240
rect 16425 1205 16430 1235
rect 16460 1230 16465 1235
rect 16535 1235 16575 1240
rect 16535 1230 16540 1235
rect 16460 1210 16540 1230
rect 16460 1205 16465 1210
rect 16425 1200 16465 1205
rect 16535 1205 16540 1210
rect 16570 1230 16575 1235
rect 16645 1235 16685 1240
rect 16645 1230 16650 1235
rect 16570 1210 16650 1230
rect 16570 1205 16575 1210
rect 16535 1200 16575 1205
rect 16645 1205 16650 1210
rect 16680 1230 16685 1235
rect 16755 1235 16795 1240
rect 16755 1230 16760 1235
rect 16680 1210 16760 1230
rect 16680 1205 16685 1210
rect 16645 1200 16685 1205
rect 16755 1205 16760 1210
rect 16790 1230 16795 1235
rect 16865 1235 16905 1240
rect 16865 1230 16870 1235
rect 16790 1210 16870 1230
rect 16790 1205 16795 1210
rect 16755 1200 16795 1205
rect 16865 1205 16870 1210
rect 16900 1230 16905 1235
rect 16975 1235 17015 1240
rect 16975 1230 16980 1235
rect 16900 1210 16980 1230
rect 16900 1205 16905 1210
rect 16865 1200 16905 1205
rect 16975 1205 16980 1210
rect 17010 1230 17015 1235
rect 17085 1235 17125 1240
rect 17085 1230 17090 1235
rect 17010 1210 17090 1230
rect 17010 1205 17015 1210
rect 16975 1200 17015 1205
rect 17085 1205 17090 1210
rect 17120 1230 17125 1235
rect 17195 1235 17235 1240
rect 17195 1230 17200 1235
rect 17120 1210 17200 1230
rect 17120 1205 17125 1210
rect 17085 1200 17125 1205
rect 17195 1205 17200 1210
rect 17230 1230 17235 1235
rect 17305 1235 17345 1240
rect 17305 1230 17310 1235
rect 17230 1210 17310 1230
rect 17230 1205 17235 1210
rect 17195 1200 17235 1205
rect 17305 1205 17310 1210
rect 17340 1230 17345 1235
rect 17415 1235 17455 1240
rect 17415 1230 17420 1235
rect 17340 1210 17420 1230
rect 17340 1205 17345 1210
rect 17305 1200 17345 1205
rect 17415 1205 17420 1210
rect 17450 1230 17455 1235
rect 17525 1235 17565 1240
rect 17525 1230 17530 1235
rect 17450 1210 17530 1230
rect 17450 1205 17455 1210
rect 17415 1200 17455 1205
rect 17525 1205 17530 1210
rect 17560 1205 17565 1235
rect 17595 1220 17600 1250
rect 17630 1245 17635 1250
rect 17805 1250 17845 1255
rect 17805 1245 17810 1250
rect 17630 1225 17810 1245
rect 17630 1220 17635 1225
rect 17595 1215 17635 1220
rect 17805 1220 17810 1225
rect 17840 1220 17845 1250
rect 17805 1215 17845 1220
rect 17525 1200 17565 1205
rect 3375 1185 3415 1190
rect 3375 1155 3380 1185
rect 3410 1180 3415 1185
rect 3985 1185 4025 1190
rect 3985 1180 3990 1185
rect 3410 1160 3990 1180
rect 3410 1155 3415 1160
rect 3375 1150 3415 1155
rect 3985 1155 3990 1160
rect 4020 1180 4025 1185
rect 4595 1185 4635 1190
rect 4595 1180 4600 1185
rect 4020 1160 4600 1180
rect 4020 1155 4025 1160
rect 3985 1150 4025 1155
rect 4595 1155 4600 1160
rect 4630 1180 4635 1185
rect 5465 1185 5505 1190
rect 5465 1180 5470 1185
rect 4630 1160 5470 1180
rect 4630 1155 4635 1160
rect 4595 1150 4635 1155
rect 5465 1155 5470 1160
rect 5500 1155 5505 1185
rect 5465 1150 5505 1155
rect 2945 1125 2985 1130
rect 2945 1095 2950 1125
rect 2980 1120 2985 1125
rect 3025 1125 3065 1130
rect 3025 1120 3030 1125
rect 2980 1100 3030 1120
rect 2980 1095 2985 1100
rect 2945 1090 2985 1095
rect 3025 1095 3030 1100
rect 3060 1120 3065 1125
rect 3105 1125 3145 1130
rect 3105 1120 3110 1125
rect 3060 1100 3110 1120
rect 3060 1095 3065 1100
rect 3025 1090 3065 1095
rect 3105 1095 3110 1100
rect 3140 1120 3145 1125
rect 3185 1125 3225 1130
rect 3185 1120 3190 1125
rect 3140 1100 3190 1120
rect 3140 1095 3145 1100
rect 3105 1090 3145 1095
rect 3185 1095 3190 1100
rect 3220 1120 3225 1125
rect 3265 1125 3305 1130
rect 3265 1120 3270 1125
rect 3220 1100 3270 1120
rect 3220 1095 3225 1100
rect 3185 1090 3225 1095
rect 3265 1095 3270 1100
rect 3300 1120 3305 1125
rect 3345 1125 3385 1130
rect 3345 1120 3350 1125
rect 3300 1100 3350 1120
rect 3300 1095 3305 1100
rect 3265 1090 3305 1095
rect 3345 1095 3350 1100
rect 3380 1120 3385 1125
rect 3425 1125 3465 1130
rect 3425 1120 3430 1125
rect 3380 1100 3430 1120
rect 3380 1095 3385 1100
rect 3345 1090 3385 1095
rect 3425 1095 3430 1100
rect 3460 1120 3465 1125
rect 3505 1125 3545 1130
rect 3505 1120 3510 1125
rect 3460 1100 3510 1120
rect 3460 1095 3465 1100
rect 3425 1090 3465 1095
rect 3505 1095 3510 1100
rect 3540 1120 3545 1125
rect 3585 1125 3625 1130
rect 3585 1120 3590 1125
rect 3540 1100 3590 1120
rect 3540 1095 3545 1100
rect 3505 1090 3545 1095
rect 3585 1095 3590 1100
rect 3620 1120 3625 1125
rect 3665 1125 3705 1130
rect 3665 1120 3670 1125
rect 3620 1100 3670 1120
rect 3620 1095 3625 1100
rect 3585 1090 3625 1095
rect 3665 1095 3670 1100
rect 3700 1120 3705 1125
rect 3745 1125 3785 1130
rect 3745 1120 3750 1125
rect 3700 1100 3750 1120
rect 3700 1095 3705 1100
rect 3665 1090 3705 1095
rect 3745 1095 3750 1100
rect 3780 1120 3785 1125
rect 3825 1125 3865 1130
rect 3825 1120 3830 1125
rect 3780 1100 3830 1120
rect 3780 1095 3785 1100
rect 3745 1090 3785 1095
rect 3825 1095 3830 1100
rect 3860 1120 3865 1125
rect 3905 1125 3945 1130
rect 3905 1120 3910 1125
rect 3860 1100 3910 1120
rect 3860 1095 3865 1100
rect 3825 1090 3865 1095
rect 3905 1095 3910 1100
rect 3940 1095 3945 1125
rect 3905 1090 3945 1095
rect 3985 1125 4025 1130
rect 3985 1095 3990 1125
rect 4020 1120 4025 1125
rect 4065 1125 4105 1130
rect 4065 1120 4070 1125
rect 4020 1100 4070 1120
rect 4020 1095 4025 1100
rect 3985 1090 4025 1095
rect 4065 1095 4070 1100
rect 4100 1120 4105 1125
rect 4145 1125 4185 1130
rect 4145 1120 4150 1125
rect 4100 1100 4150 1120
rect 4100 1095 4105 1100
rect 4065 1090 4105 1095
rect 4145 1095 4150 1100
rect 4180 1120 4185 1125
rect 4225 1125 4265 1130
rect 4225 1120 4230 1125
rect 4180 1100 4230 1120
rect 4180 1095 4185 1100
rect 4145 1090 4185 1095
rect 4225 1095 4230 1100
rect 4260 1120 4265 1125
rect 4305 1125 4345 1130
rect 4305 1120 4310 1125
rect 4260 1100 4310 1120
rect 4260 1095 4265 1100
rect 4225 1090 4265 1095
rect 4305 1095 4310 1100
rect 4340 1120 4345 1125
rect 4385 1125 4425 1130
rect 4385 1120 4390 1125
rect 4340 1100 4390 1120
rect 4340 1095 4345 1100
rect 4305 1090 4345 1095
rect 4385 1095 4390 1100
rect 4420 1120 4425 1125
rect 4465 1125 4505 1130
rect 4465 1120 4470 1125
rect 4420 1100 4470 1120
rect 4420 1095 4425 1100
rect 4385 1090 4425 1095
rect 4465 1095 4470 1100
rect 4500 1120 4505 1125
rect 4545 1125 4585 1130
rect 4545 1120 4550 1125
rect 4500 1100 4550 1120
rect 4500 1095 4505 1100
rect 4465 1090 4505 1095
rect 4545 1095 4550 1100
rect 4580 1120 4585 1125
rect 4625 1125 4665 1130
rect 4625 1120 4630 1125
rect 4580 1100 4630 1120
rect 4580 1095 4585 1100
rect 4545 1090 4585 1095
rect 4625 1095 4630 1100
rect 4660 1120 4665 1125
rect 4705 1125 4745 1130
rect 4705 1120 4710 1125
rect 4660 1100 4710 1120
rect 4660 1095 4665 1100
rect 4625 1090 4665 1095
rect 4705 1095 4710 1100
rect 4740 1120 4745 1125
rect 4785 1125 4825 1130
rect 4785 1120 4790 1125
rect 4740 1100 4790 1120
rect 4740 1095 4745 1100
rect 4705 1090 4745 1095
rect 4785 1095 4790 1100
rect 4820 1120 4825 1125
rect 4865 1125 4905 1130
rect 4865 1120 4870 1125
rect 4820 1100 4870 1120
rect 4820 1095 4825 1100
rect 4785 1090 4825 1095
rect 4865 1095 4870 1100
rect 4900 1120 4905 1125
rect 4945 1125 4985 1130
rect 4945 1120 4950 1125
rect 4900 1100 4950 1120
rect 4900 1095 4905 1100
rect 4865 1090 4905 1095
rect 4945 1095 4950 1100
rect 4980 1095 4985 1125
rect 4945 1090 4985 1095
rect 2620 1040 2660 1045
rect 2620 1010 2625 1040
rect 2655 1035 2660 1040
rect 2905 1040 2945 1045
rect 2905 1035 2910 1040
rect 2655 1015 2910 1035
rect 2655 1010 2660 1015
rect 2620 1005 2660 1010
rect 2905 1010 2910 1015
rect 2940 1010 2945 1040
rect 2905 1005 2945 1010
rect 5110 1040 5150 1045
rect 5110 1010 5115 1040
rect 5145 1035 5150 1040
rect 5465 1040 5505 1045
rect 5465 1035 5470 1040
rect 5145 1015 5470 1035
rect 5145 1010 5150 1015
rect 5110 1005 5150 1010
rect 5465 1010 5470 1015
rect 5500 1010 5505 1040
rect 5465 1005 5505 1010
rect 15355 935 15395 940
rect 2995 930 3035 935
rect 2995 900 3000 930
rect 3030 925 3035 930
rect 3175 930 3215 935
rect 3175 925 3180 930
rect 3030 905 3180 925
rect 3030 900 3035 905
rect 2995 895 3035 900
rect 3175 900 3180 905
rect 3210 925 3215 930
rect 3355 930 3395 935
rect 3355 925 3360 930
rect 3210 905 3360 925
rect 3210 900 3215 905
rect 3175 895 3215 900
rect 3355 900 3360 905
rect 3390 925 3395 930
rect 3535 930 3575 935
rect 3535 925 3540 930
rect 3390 905 3540 925
rect 3390 900 3395 905
rect 3355 895 3395 900
rect 3535 900 3540 905
rect 3570 925 3575 930
rect 3715 930 3755 935
rect 3715 925 3720 930
rect 3570 905 3720 925
rect 3570 900 3575 905
rect 3535 895 3575 900
rect 3715 900 3720 905
rect 3750 925 3755 930
rect 3895 930 3935 935
rect 3895 925 3900 930
rect 3750 905 3900 925
rect 3750 900 3755 905
rect 3715 895 3755 900
rect 3895 900 3900 905
rect 3930 925 3935 930
rect 4075 930 4115 935
rect 4075 925 4080 930
rect 3930 905 4080 925
rect 3930 900 3935 905
rect 3895 895 3935 900
rect 4075 900 4080 905
rect 4110 925 4115 930
rect 4255 930 4295 935
rect 4255 925 4260 930
rect 4110 905 4260 925
rect 4110 900 4115 905
rect 4075 895 4115 900
rect 4255 900 4260 905
rect 4290 925 4295 930
rect 4435 930 4475 935
rect 4435 925 4440 930
rect 4290 905 4440 925
rect 4290 900 4295 905
rect 4255 895 4295 900
rect 4435 900 4440 905
rect 4470 925 4475 930
rect 4615 930 4655 935
rect 4615 925 4620 930
rect 4470 905 4620 925
rect 4470 900 4475 905
rect 4435 895 4475 900
rect 4615 900 4620 905
rect 4650 925 4655 930
rect 4795 930 4835 935
rect 4795 925 4800 930
rect 4650 905 4800 925
rect 4650 900 4655 905
rect 4615 895 4655 900
rect 4795 900 4800 905
rect 4830 925 4835 930
rect 4975 930 5015 935
rect 4975 925 4980 930
rect 4830 905 4980 925
rect 4830 900 4835 905
rect 4795 895 4835 900
rect 4975 900 4980 905
rect 5010 925 5015 930
rect 5465 930 5505 935
rect 5465 925 5470 930
rect 5010 905 5470 925
rect 5010 900 5015 905
rect 4975 895 5015 900
rect 5465 900 5470 905
rect 5500 900 5505 930
rect 15355 905 15360 935
rect 15390 930 15395 935
rect 15555 935 15595 940
rect 15555 930 15560 935
rect 15390 910 15560 930
rect 15390 905 15395 910
rect 15355 900 15395 905
rect 15555 905 15560 910
rect 15590 905 15595 935
rect 18205 935 18245 940
rect 15555 900 15595 905
rect 16165 915 16205 920
rect 5465 895 5505 900
rect 16165 885 16170 915
rect 16200 910 16205 915
rect 16260 915 16300 920
rect 16260 910 16265 915
rect 16200 890 16265 910
rect 16200 885 16205 890
rect 16165 880 16205 885
rect 16260 885 16265 890
rect 16295 910 16300 915
rect 16370 915 16410 920
rect 16370 910 16375 915
rect 16295 890 16375 910
rect 16295 885 16300 890
rect 16260 880 16300 885
rect 16370 885 16375 890
rect 16405 910 16410 915
rect 16480 915 16520 920
rect 16480 910 16485 915
rect 16405 890 16485 910
rect 16405 885 16410 890
rect 16370 880 16410 885
rect 16480 885 16485 890
rect 16515 910 16520 915
rect 16590 915 16630 920
rect 16590 910 16595 915
rect 16515 890 16595 910
rect 16515 885 16520 890
rect 16480 880 16520 885
rect 16590 885 16595 890
rect 16625 910 16630 915
rect 16700 915 16740 920
rect 16700 910 16705 915
rect 16625 890 16705 910
rect 16625 885 16630 890
rect 16590 880 16630 885
rect 16700 885 16705 890
rect 16735 910 16740 915
rect 16810 915 16850 920
rect 16810 910 16815 915
rect 16735 890 16815 910
rect 16735 885 16740 890
rect 16700 880 16740 885
rect 16810 885 16815 890
rect 16845 910 16850 915
rect 16920 915 16960 920
rect 16920 910 16925 915
rect 16845 890 16925 910
rect 16845 885 16850 890
rect 16810 880 16850 885
rect 16920 885 16925 890
rect 16955 910 16960 915
rect 17030 915 17070 920
rect 17030 910 17035 915
rect 16955 890 17035 910
rect 16955 885 16960 890
rect 16920 880 16960 885
rect 17030 885 17035 890
rect 17065 910 17070 915
rect 17140 915 17180 920
rect 17140 910 17145 915
rect 17065 890 17145 910
rect 17065 885 17070 890
rect 17030 880 17070 885
rect 17140 885 17145 890
rect 17175 910 17180 915
rect 17250 915 17290 920
rect 17250 910 17255 915
rect 17175 890 17255 910
rect 17175 885 17180 890
rect 17140 880 17180 885
rect 17250 885 17255 890
rect 17285 910 17290 915
rect 17360 915 17400 920
rect 17360 910 17365 915
rect 17285 890 17365 910
rect 17285 885 17290 890
rect 17250 880 17290 885
rect 17360 885 17365 890
rect 17395 910 17400 915
rect 17470 915 17510 920
rect 17470 910 17475 915
rect 17395 890 17475 910
rect 17395 885 17400 890
rect 17360 880 17400 885
rect 17470 885 17475 890
rect 17505 910 17510 915
rect 17620 915 17660 920
rect 17620 910 17625 915
rect 17505 890 17625 910
rect 17505 885 17510 890
rect 17470 880 17510 885
rect 17620 885 17625 890
rect 17655 885 17660 915
rect 18205 905 18210 935
rect 18240 930 18245 935
rect 18405 935 18445 940
rect 18405 930 18410 935
rect 18240 910 18410 930
rect 18240 905 18245 910
rect 18205 900 18245 905
rect 18405 905 18410 910
rect 18440 905 18445 935
rect 18405 900 18445 905
rect 17620 880 17660 885
rect 16935 860 16975 865
rect 16005 855 16045 860
rect 16005 825 16010 855
rect 16040 850 16045 855
rect 16495 855 16535 860
rect 16495 850 16500 855
rect 16040 830 16500 850
rect 16040 825 16045 830
rect 16005 820 16045 825
rect 16495 825 16500 830
rect 16530 825 16535 855
rect 16935 830 16940 860
rect 16970 855 16975 860
rect 17155 860 17195 865
rect 17155 855 17160 860
rect 16970 835 17160 855
rect 16970 830 16975 835
rect 16935 825 16975 830
rect 17155 830 17160 835
rect 17190 855 17195 860
rect 17375 860 17415 865
rect 17375 855 17380 860
rect 17190 835 17380 855
rect 17190 830 17195 835
rect 17155 825 17195 830
rect 17375 830 17380 835
rect 17410 855 17415 860
rect 17860 860 17900 865
rect 17860 855 17865 860
rect 17410 835 17865 855
rect 17410 830 17415 835
rect 17375 825 17415 830
rect 17860 830 17865 835
rect 17895 830 17900 860
rect 17860 825 17900 830
rect 16495 820 16535 825
rect 17045 800 17085 805
rect 15950 795 15990 800
rect 15950 765 15955 795
rect 15985 790 15990 795
rect 16305 795 16345 800
rect 16305 790 16310 795
rect 15985 770 16310 790
rect 15985 765 15990 770
rect 2520 760 2560 765
rect 2520 730 2525 760
rect 2555 755 2560 760
rect 3130 760 3170 765
rect 3130 755 3135 760
rect 2555 735 3135 755
rect 2555 730 2560 735
rect 2520 725 2560 730
rect 3130 730 3135 735
rect 3165 730 3170 760
rect 3130 725 3170 730
rect 3625 760 3665 765
rect 3625 730 3630 760
rect 3660 755 3665 760
rect 3985 760 4025 765
rect 3985 755 3990 760
rect 3660 735 3990 755
rect 3660 730 3665 735
rect 3625 725 3665 730
rect 3985 730 3990 735
rect 4020 755 4025 760
rect 4345 760 4385 765
rect 4345 755 4350 760
rect 4020 735 4350 755
rect 4020 730 4025 735
rect 3985 725 4025 730
rect 4345 730 4350 735
rect 4380 730 4385 760
rect 4345 725 4385 730
rect 4525 760 4565 765
rect 4525 730 4530 760
rect 4560 755 4565 760
rect 4705 760 4745 765
rect 4705 755 4710 760
rect 4560 735 4710 755
rect 4560 730 4565 735
rect 4525 725 4565 730
rect 4705 730 4710 735
rect 4740 755 4745 760
rect 4885 760 4925 765
rect 15950 760 15990 765
rect 16305 765 16310 770
rect 16340 790 16345 795
rect 16375 795 16415 800
rect 16375 790 16380 795
rect 16340 770 16380 790
rect 16340 765 16345 770
rect 16305 760 16345 765
rect 16375 765 16380 770
rect 16410 790 16415 795
rect 16445 795 16485 800
rect 16445 790 16450 795
rect 16410 770 16450 790
rect 16410 765 16415 770
rect 16375 760 16415 765
rect 16445 765 16450 770
rect 16480 765 16485 795
rect 17045 770 17050 800
rect 17080 795 17085 800
rect 17265 800 17305 805
rect 17265 795 17270 800
rect 17080 775 17270 795
rect 17080 770 17085 775
rect 17045 765 17085 770
rect 17265 770 17270 775
rect 17300 795 17305 800
rect 17485 800 17525 805
rect 17485 795 17490 800
rect 17300 775 17490 795
rect 17300 770 17305 775
rect 17265 765 17305 770
rect 17485 770 17490 775
rect 17520 795 17525 800
rect 17805 800 17845 805
rect 17805 795 17810 800
rect 17520 775 17810 795
rect 17520 770 17525 775
rect 17485 765 17525 770
rect 17805 770 17810 775
rect 17840 770 17845 800
rect 17805 765 17845 770
rect 16445 760 16485 765
rect 4885 755 4890 760
rect 4740 735 4890 755
rect 4740 730 4745 735
rect 4705 725 4745 730
rect 4885 730 4890 735
rect 4920 730 4925 760
rect 4885 725 4925 730
rect 3445 705 3485 710
rect 3445 675 3450 705
rect 3480 700 3485 705
rect 3805 705 3845 710
rect 3805 700 3810 705
rect 3480 680 3810 700
rect 3480 675 3485 680
rect 3445 670 3485 675
rect 3805 675 3810 680
rect 3840 700 3845 705
rect 4165 705 4205 710
rect 4165 700 4170 705
rect 3840 680 4170 700
rect 3840 675 3845 680
rect 3805 670 3845 675
rect 4165 675 4170 680
rect 4200 675 4205 705
rect 4165 670 4205 675
rect 16990 680 17030 685
rect 16990 650 16995 680
rect 17025 675 17030 680
rect 17100 680 17140 685
rect 17100 675 17105 680
rect 17025 655 17105 675
rect 17025 650 17030 655
rect 16990 645 17030 650
rect 17100 650 17105 655
rect 17135 675 17140 680
rect 17210 680 17250 685
rect 17210 675 17215 680
rect 17135 655 17215 675
rect 17135 650 17140 655
rect 17100 645 17140 650
rect 17210 650 17215 655
rect 17245 675 17250 680
rect 17320 680 17360 685
rect 17320 675 17325 680
rect 17245 655 17325 675
rect 17245 650 17250 655
rect 17210 645 17250 650
rect 17320 650 17325 655
rect 17355 675 17360 680
rect 17430 680 17470 685
rect 17430 675 17435 680
rect 17355 655 17435 675
rect 17355 650 17360 655
rect 17320 645 17360 650
rect 17430 650 17435 655
rect 17465 650 17470 680
rect 17430 645 17470 650
rect -195 575 -155 580
rect -195 545 -190 575
rect -160 545 -155 575
rect -195 540 -155 545
<< via2 >>
rect -190 4960 -160 4990
rect 5555 4960 5585 4990
rect 14960 3605 14990 3635
rect 18810 3605 18840 3635
rect -105 3495 -75 3525
rect 4445 3465 4475 3495
rect 945 3415 975 3445
rect 1645 3415 1675 3445
rect 5145 3415 5175 3445
rect 5555 3415 5585 3445
rect 2695 3360 2725 3390
rect 3395 3305 3425 3335
rect -105 3110 -75 3140
rect -105 2970 -75 3000
rect -105 2880 -75 2910
rect 5555 2780 5585 2810
rect 5555 2065 5585 2095
rect 14520 2080 14550 2110
rect 19250 2080 19280 2110
rect -105 1690 -75 1720
rect 5555 1470 5585 1500
rect 5470 1155 5500 1185
rect 5470 1010 5500 1040
rect 5470 900 5500 930
rect -190 545 -160 575
<< metal3 >>
rect 12760 5620 12990 5705
rect 13110 5620 13340 5705
rect 13460 5620 13690 5705
rect 12760 5570 13690 5620
rect 12760 5475 12990 5570
rect 13110 5475 13340 5570
rect 13460 5475 13690 5570
rect 13810 5475 14040 5705
rect 14160 5475 14390 5705
rect 14510 5475 14740 5705
rect 14860 5475 15090 5705
rect 15210 5475 15440 5705
rect 15560 5475 15790 5705
rect 15910 5475 16140 5705
rect 16260 5475 16490 5705
rect 16610 5475 16840 5705
rect 16960 5475 17190 5705
rect 17310 5475 17540 5705
rect 17660 5475 17890 5705
rect 18010 5475 18240 5705
rect 18360 5475 18590 5705
rect 18710 5475 18940 5705
rect 19060 5475 19290 5705
rect 19410 5475 19640 5705
rect 19760 5475 19990 5705
rect 20110 5620 20340 5705
rect 20460 5620 20690 5705
rect 20810 5620 21040 5705
rect 20110 5570 21040 5620
rect 20110 5475 20340 5570
rect 20460 5475 20690 5570
rect 20810 5475 21040 5570
rect 13550 5355 13600 5475
rect 13900 5355 13950 5475
rect 14250 5355 14300 5475
rect 14600 5355 14650 5475
rect 14950 5355 15000 5475
rect 15300 5355 15350 5475
rect 15650 5355 15700 5475
rect 16000 5355 16050 5475
rect 16350 5355 16400 5475
rect 16700 5355 16750 5475
rect 17050 5355 17100 5475
rect 17400 5355 17450 5475
rect 17750 5355 17800 5475
rect 18100 5355 18150 5475
rect 18450 5355 18500 5475
rect 18800 5355 18850 5475
rect 19150 5355 19200 5475
rect 19500 5355 19550 5475
rect 19850 5355 19900 5475
rect 20200 5355 20250 5475
rect 12760 5270 12990 5355
rect 13110 5270 13340 5355
rect 13460 5270 13690 5355
rect 13810 5270 14040 5355
rect 14160 5270 14390 5355
rect 14510 5270 14740 5355
rect 14860 5270 15090 5355
rect 15210 5270 15440 5355
rect 15560 5270 15790 5355
rect 15910 5270 16140 5355
rect 16260 5270 16490 5355
rect 16610 5270 16840 5355
rect 12760 5220 16840 5270
rect 12760 5125 12990 5220
rect 13110 5125 13340 5220
rect 13460 5125 13690 5220
rect 13810 5125 14040 5220
rect 14160 5125 14390 5220
rect 14510 5125 14740 5220
rect 14860 5125 15090 5220
rect 15210 5125 15440 5220
rect 15560 5125 15790 5220
rect 15910 5125 16140 5220
rect 16260 5125 16490 5220
rect 16610 5125 16840 5220
rect 16960 5270 17190 5355
rect 17310 5270 17540 5355
rect 17660 5270 17890 5355
rect 18010 5270 18240 5355
rect 18360 5270 18590 5355
rect 18710 5270 18940 5355
rect 19060 5270 19290 5355
rect 19410 5270 19640 5355
rect 19760 5270 19990 5355
rect 20110 5270 20340 5355
rect 20460 5270 20690 5355
rect 20810 5270 21040 5355
rect 16960 5220 21040 5270
rect 16960 5125 17190 5220
rect 17310 5125 17540 5220
rect 17660 5125 17890 5220
rect 18010 5125 18240 5220
rect 18360 5125 18590 5220
rect 18710 5125 18940 5220
rect 19060 5125 19290 5220
rect 19410 5125 19640 5220
rect 19760 5125 19990 5220
rect 20110 5125 20340 5220
rect 20460 5125 20690 5220
rect 20810 5125 21040 5220
rect 13550 5005 13600 5125
rect 14600 5005 14650 5125
rect 14950 5005 15000 5125
rect 15300 5005 15350 5125
rect 15650 5005 15700 5125
rect 16000 5005 16050 5125
rect 16350 5005 16400 5125
rect 16700 5005 16750 5125
rect 17050 5005 17100 5125
rect 17400 5005 17450 5125
rect 17750 5005 17800 5125
rect 18100 5005 18150 5125
rect 18450 5005 18500 5125
rect 18800 5005 18850 5125
rect 19150 5005 19200 5125
rect 20200 5005 20250 5125
rect -200 4995 -150 5000
rect -200 4955 -195 4995
rect -155 4955 -150 4995
rect -200 4950 -150 4955
rect 5545 4995 5595 5000
rect 5545 4955 5550 4995
rect 5590 4955 5595 4995
rect 5545 4950 5595 4955
rect -195 585 -155 4950
rect -115 4910 -65 4915
rect -115 4870 -110 4910
rect -70 4870 -65 4910
rect -115 4865 -65 4870
rect 5460 4910 5510 4915
rect 5460 4870 5465 4910
rect 5505 4870 5510 4910
rect 5460 4865 5510 4870
rect -110 3525 -70 4865
rect 145 4770 375 4855
rect 495 4770 725 4855
rect 845 4770 1075 4855
rect 1195 4770 1425 4855
rect 1545 4770 1775 4855
rect 145 4720 1775 4770
rect 145 4625 375 4720
rect 495 4625 725 4720
rect 845 4625 1075 4720
rect 1195 4625 1425 4720
rect 1545 4625 1775 4720
rect 1895 4770 2125 4855
rect 2245 4770 2475 4855
rect 2595 4770 2825 4855
rect 2945 4770 3175 4855
rect 3295 4770 3525 4855
rect 1895 4720 3525 4770
rect 1895 4625 2125 4720
rect 2245 4625 2475 4720
rect 2595 4625 2825 4720
rect 2945 4625 3175 4720
rect 3295 4625 3525 4720
rect 3645 4770 3875 4855
rect 3995 4770 4225 4855
rect 4345 4770 4575 4855
rect 4695 4770 4925 4855
rect 5045 4770 5275 4855
rect 3645 4720 5275 4770
rect 3645 4625 3875 4720
rect 3995 4625 4225 4720
rect 4345 4625 4575 4720
rect 4695 4625 4925 4720
rect 5045 4625 5275 4720
rect 935 4505 985 4625
rect 2685 4505 2735 4625
rect 4435 4505 4485 4625
rect 145 4420 375 4505
rect 495 4420 725 4505
rect 845 4420 1075 4505
rect 1195 4420 1425 4505
rect 1545 4420 1775 4505
rect 145 4370 1775 4420
rect 145 4275 375 4370
rect 495 4275 725 4370
rect 845 4275 1075 4370
rect 1195 4275 1425 4370
rect 1545 4275 1775 4370
rect 1895 4420 2125 4505
rect 2245 4420 2475 4505
rect 2595 4420 2825 4505
rect 2945 4420 3175 4505
rect 3295 4420 3525 4505
rect 1895 4370 3525 4420
rect 1895 4275 2125 4370
rect 2245 4275 2475 4370
rect 2595 4275 2825 4370
rect 2945 4275 3175 4370
rect 3295 4275 3525 4370
rect 3645 4420 3875 4505
rect 3995 4420 4225 4505
rect 4345 4420 4575 4505
rect 4695 4420 4925 4505
rect 5045 4420 5275 4505
rect 3645 4370 5275 4420
rect 3645 4275 3875 4370
rect 3995 4275 4225 4370
rect 4345 4275 4575 4370
rect 4695 4275 4925 4370
rect 5045 4275 5275 4370
rect 935 4155 985 4275
rect 2685 4155 2735 4275
rect 4435 4155 4485 4275
rect 145 4070 375 4155
rect 495 4070 725 4155
rect 845 4070 1075 4155
rect 1195 4070 1425 4155
rect 1545 4070 1775 4155
rect 145 4020 1775 4070
rect 145 3925 375 4020
rect 495 3925 725 4020
rect 845 3925 1075 4020
rect 1195 3925 1425 4020
rect 1545 3925 1775 4020
rect 1895 4070 2125 4155
rect 2245 4070 2475 4155
rect 2595 4070 2825 4155
rect 2945 4070 3175 4155
rect 3295 4070 3525 4155
rect 1895 4020 3525 4070
rect 1895 3925 2125 4020
rect 2245 3925 2475 4020
rect 2595 3925 2825 4020
rect 2945 3925 3175 4020
rect 3295 3925 3525 4020
rect 3645 4070 3875 4155
rect 3995 4070 4225 4155
rect 4345 4070 4575 4155
rect 4695 4070 4925 4155
rect 5045 4070 5275 4155
rect 3645 4020 5275 4070
rect 3645 3925 3875 4020
rect 3995 3925 4225 4020
rect 4345 3925 4575 4020
rect 4695 3925 4925 4020
rect 5045 3925 5275 4020
rect 935 3805 985 3925
rect 2685 3805 2735 3925
rect 4435 3805 4485 3925
rect 145 3720 375 3805
rect 495 3720 725 3805
rect 845 3720 1075 3805
rect 1195 3720 1425 3805
rect 1545 3720 1775 3805
rect 145 3670 1775 3720
rect 145 3575 375 3670
rect 495 3575 725 3670
rect 845 3575 1075 3670
rect 1195 3575 1425 3670
rect 1545 3575 1775 3670
rect 1895 3720 2125 3805
rect 2245 3720 2475 3805
rect 2595 3720 2825 3805
rect 2945 3720 3175 3805
rect 3295 3720 3525 3805
rect 1895 3670 3525 3720
rect 1895 3575 2125 3670
rect 2245 3575 2475 3670
rect 2595 3575 2825 3670
rect 2945 3575 3175 3670
rect 3295 3575 3525 3670
rect 3645 3720 3875 3805
rect 3995 3720 4225 3805
rect 4345 3720 4575 3805
rect 4695 3720 4925 3805
rect 5045 3720 5275 3805
rect 3645 3670 5275 3720
rect 3645 3575 3875 3670
rect 3995 3575 4225 3670
rect 4345 3575 4575 3670
rect 4695 3575 4925 3670
rect 5045 3575 5275 3670
rect -110 3495 -105 3525
rect -75 3495 -70 3525
rect -110 3140 -70 3495
rect 940 3445 980 3575
rect 940 3415 945 3445
rect 975 3415 980 3445
rect 940 3410 980 3415
rect 1635 3450 1685 3455
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 2690 3390 2730 3575
rect 4440 3495 4480 3575
rect 4440 3465 4445 3495
rect 4475 3465 4480 3495
rect 4440 3460 4480 3465
rect 5135 3450 5185 3455
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 2690 3360 2695 3390
rect 2725 3360 2730 3390
rect 2690 3355 2730 3360
rect 3385 3340 3435 3345
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect -110 3110 -105 3140
rect -75 3110 -70 3140
rect -110 3000 -70 3110
rect -110 2970 -105 3000
rect -75 2970 -70 3000
rect -110 2910 -70 2970
rect -110 2880 -105 2910
rect -75 2880 -70 2910
rect -110 1720 -70 2880
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 665 -70 1690
rect 5465 1185 5505 4865
rect 5465 1155 5470 1185
rect 5500 1155 5505 1185
rect 5465 1040 5505 1155
rect 5465 1010 5470 1040
rect 5500 1010 5505 1040
rect 5465 930 5505 1010
rect 5465 900 5470 930
rect 5500 900 5505 930
rect 5465 665 5505 900
rect 5550 3445 5590 4950
rect 12760 4920 12990 5005
rect 13110 4920 13340 5005
rect 13460 4920 13690 5005
rect 13810 4920 14040 5005
rect 14160 4920 14390 5005
rect 12760 4870 14390 4920
rect 12760 4775 12990 4870
rect 13110 4775 13340 4870
rect 13460 4775 13690 4870
rect 13810 4775 14040 4870
rect 14160 4775 14390 4870
rect 14510 4775 14740 5005
rect 14860 4775 15090 5005
rect 15210 4775 15440 5005
rect 15560 4775 15790 5005
rect 15910 4775 16140 5005
rect 16260 4775 16490 5005
rect 16610 4775 16840 5005
rect 16960 4775 17190 5005
rect 17310 4775 17540 5005
rect 17660 4775 17890 5005
rect 18010 4775 18240 5005
rect 18360 4775 18590 5005
rect 18710 4775 18940 5005
rect 19060 4775 19290 5005
rect 19410 4920 19640 5005
rect 19760 4920 19990 5005
rect 20110 4920 20340 5005
rect 20460 4920 20690 5005
rect 20810 4920 21040 5005
rect 19410 4870 21040 4920
rect 19410 4775 19640 4870
rect 19760 4775 19990 4870
rect 20110 4775 20340 4870
rect 20460 4775 20690 4870
rect 20810 4775 21040 4870
rect 13550 4655 13600 4775
rect 14600 4655 14650 4775
rect 14950 4655 15000 4775
rect 15300 4655 15350 4775
rect 15650 4655 15700 4775
rect 18100 4655 18150 4775
rect 18450 4655 18500 4775
rect 18800 4655 18850 4775
rect 19150 4655 19200 4775
rect 20200 4655 20250 4775
rect 12760 4570 12990 4655
rect 13110 4570 13340 4655
rect 13460 4570 13690 4655
rect 13810 4570 14040 4655
rect 14160 4570 14390 4655
rect 12760 4520 14390 4570
rect 12760 4425 12990 4520
rect 13110 4425 13340 4520
rect 13460 4425 13690 4520
rect 13810 4425 14040 4520
rect 14160 4425 14390 4520
rect 14510 4425 14740 4655
rect 14860 4425 15090 4655
rect 15210 4425 15440 4655
rect 15560 4425 15790 4655
rect 18010 4425 18240 4655
rect 18360 4425 18590 4655
rect 18710 4425 18940 4655
rect 19060 4425 19290 4655
rect 19410 4570 19640 4655
rect 19760 4570 19990 4655
rect 20110 4570 20340 4655
rect 20460 4570 20690 4655
rect 20810 4570 21040 4655
rect 19410 4520 21040 4570
rect 19410 4425 19640 4520
rect 19760 4425 19990 4520
rect 20110 4425 20340 4520
rect 20460 4425 20690 4520
rect 20810 4425 21040 4520
rect 13550 4305 13600 4425
rect 14600 4305 14650 4425
rect 14950 4305 15000 4425
rect 15300 4305 15350 4425
rect 15650 4305 15700 4425
rect 18100 4305 18150 4425
rect 18450 4305 18500 4425
rect 18800 4305 18850 4425
rect 19150 4305 19200 4425
rect 20200 4305 20250 4425
rect 12760 4220 12990 4305
rect 13110 4220 13340 4305
rect 13460 4220 13690 4305
rect 13810 4220 14040 4305
rect 14160 4220 14390 4305
rect 12760 4170 14390 4220
rect 12760 4075 12990 4170
rect 13110 4075 13340 4170
rect 13460 4075 13690 4170
rect 13810 4075 14040 4170
rect 14160 4075 14390 4170
rect 14510 4075 14740 4305
rect 14860 4075 15090 4305
rect 15210 4075 15440 4305
rect 15560 4075 15790 4305
rect 18010 4075 18240 4305
rect 18360 4075 18590 4305
rect 18710 4075 18940 4305
rect 19060 4075 19290 4305
rect 19410 4220 19640 4305
rect 19760 4220 19990 4305
rect 20110 4220 20340 4305
rect 20460 4220 20690 4305
rect 20810 4220 21040 4305
rect 19410 4170 21040 4220
rect 19410 4075 19640 4170
rect 19760 4075 19990 4170
rect 20110 4075 20340 4170
rect 20460 4075 20690 4170
rect 20810 4075 21040 4170
rect 13550 3955 13600 4075
rect 14600 3955 14650 4075
rect 14950 3955 15000 4075
rect 15300 3955 15350 4075
rect 15650 3955 15700 4075
rect 18100 3955 18150 4075
rect 18450 3955 18500 4075
rect 18800 3955 18850 4075
rect 19150 3955 19200 4075
rect 20200 3955 20250 4075
rect 12760 3870 12990 3955
rect 13110 3870 13340 3955
rect 13460 3870 13690 3955
rect 13810 3870 14040 3955
rect 14160 3870 14390 3955
rect 12760 3820 14390 3870
rect 12760 3725 12990 3820
rect 13110 3725 13340 3820
rect 13460 3725 13690 3820
rect 13810 3725 14040 3820
rect 14160 3725 14390 3820
rect 14510 3725 14740 3955
rect 14860 3725 15090 3955
rect 15210 3725 15440 3955
rect 15560 3725 15790 3955
rect 18010 3725 18240 3955
rect 18360 3725 18590 3955
rect 18710 3725 18940 3955
rect 19060 3725 19290 3955
rect 19410 3870 19640 3955
rect 19760 3870 19990 3955
rect 20110 3870 20340 3955
rect 20460 3870 20690 3955
rect 20810 3870 21040 3955
rect 19410 3820 21040 3870
rect 19410 3725 19640 3820
rect 19760 3725 19990 3820
rect 20110 3725 20340 3820
rect 20460 3725 20690 3820
rect 20810 3725 21040 3820
rect 13550 3605 13600 3725
rect 14955 3635 14995 3725
rect 14955 3605 14960 3635
rect 14990 3605 14995 3635
rect 5550 3415 5555 3445
rect 5585 3415 5590 3445
rect 5550 2810 5590 3415
rect 12760 3520 12990 3605
rect 13110 3520 13340 3605
rect 13460 3520 13690 3605
rect 13810 3520 14040 3605
rect 14160 3520 14390 3605
rect 14955 3600 14995 3605
rect 18805 3635 18845 3725
rect 18805 3605 18810 3635
rect 18840 3605 18845 3635
rect 20200 3605 20250 3725
rect 18805 3600 18845 3605
rect 12760 3470 14390 3520
rect 12760 3375 12990 3470
rect 13110 3375 13340 3470
rect 13460 3375 13690 3470
rect 13810 3375 14040 3470
rect 14160 3375 14390 3470
rect 19410 3520 19640 3605
rect 19760 3520 19990 3605
rect 20110 3520 20340 3605
rect 20460 3520 20690 3605
rect 20810 3520 21040 3605
rect 19410 3470 21040 3520
rect 19410 3375 19640 3470
rect 19760 3375 19990 3470
rect 20110 3375 20340 3470
rect 20460 3375 20690 3470
rect 20810 3375 21040 3470
rect 13550 3255 13600 3375
rect 20200 3255 20250 3375
rect 12760 3170 12990 3255
rect 13110 3170 13340 3255
rect 13460 3170 13690 3255
rect 13810 3170 14040 3255
rect 14160 3170 14390 3255
rect 12760 3120 14390 3170
rect 12760 3025 12990 3120
rect 13110 3025 13340 3120
rect 13460 3025 13690 3120
rect 13810 3025 14040 3120
rect 14160 3025 14390 3120
rect 19410 3170 19640 3255
rect 19760 3170 19990 3255
rect 20110 3170 20340 3255
rect 20460 3170 20690 3255
rect 20810 3170 21040 3255
rect 19410 3120 21040 3170
rect 19410 3025 19640 3120
rect 19760 3025 19990 3120
rect 20110 3025 20340 3120
rect 20460 3025 20690 3120
rect 20810 3025 21040 3120
rect 13550 2905 13600 3025
rect 20200 2905 20250 3025
rect 5550 2780 5555 2810
rect 5585 2780 5590 2810
rect 5550 2095 5590 2780
rect 12760 2820 12990 2905
rect 13110 2820 13340 2905
rect 13460 2820 13690 2905
rect 13810 2820 14040 2905
rect 14160 2820 14390 2905
rect 12760 2770 14390 2820
rect 12760 2675 12990 2770
rect 13110 2675 13340 2770
rect 13460 2675 13690 2770
rect 13810 2675 14040 2770
rect 14160 2675 14390 2770
rect 19410 2820 19640 2905
rect 19760 2820 19990 2905
rect 20110 2820 20340 2905
rect 20460 2820 20690 2905
rect 20810 2820 21040 2905
rect 19410 2770 21040 2820
rect 19410 2675 19640 2770
rect 19760 2675 19990 2770
rect 20110 2675 20340 2770
rect 20460 2675 20690 2770
rect 20810 2675 21040 2770
rect 13550 2555 13600 2675
rect 20200 2555 20250 2675
rect 12760 2470 12990 2555
rect 13110 2470 13340 2555
rect 13460 2470 13690 2555
rect 13810 2470 14040 2555
rect 14160 2470 14390 2555
rect 12760 2420 14390 2470
rect 12760 2325 12990 2420
rect 13110 2325 13340 2420
rect 13460 2325 13690 2420
rect 13810 2325 14040 2420
rect 14160 2325 14390 2420
rect 19410 2470 19640 2555
rect 19760 2470 19990 2555
rect 20110 2470 20340 2555
rect 20460 2470 20690 2555
rect 20810 2470 21040 2555
rect 19410 2420 21040 2470
rect 19410 2325 19640 2420
rect 19760 2325 19990 2420
rect 20110 2325 20340 2420
rect 20460 2325 20690 2420
rect 20810 2325 21040 2420
rect 13550 2205 13600 2325
rect 20200 2205 20250 2325
rect 5550 2065 5555 2095
rect 5585 2065 5590 2095
rect 5550 1500 5590 2065
rect 12760 2120 12990 2205
rect 13110 2120 13340 2205
rect 13460 2120 13690 2205
rect 13810 2120 14040 2205
rect 14160 2120 14390 2205
rect 19410 2120 19640 2205
rect 19760 2120 19990 2205
rect 20110 2120 20340 2205
rect 20460 2120 20690 2205
rect 20810 2120 21040 2205
rect 12760 2070 14390 2120
rect 14510 2115 14560 2120
rect 14510 2075 14515 2115
rect 14555 2075 14560 2115
rect 14510 2070 14560 2075
rect 19240 2115 19290 2120
rect 19240 2075 19245 2115
rect 19285 2075 19290 2115
rect 19240 2070 19290 2075
rect 19410 2070 21040 2120
rect 12760 1975 12990 2070
rect 13110 1975 13340 2070
rect 13460 1975 13690 2070
rect 13810 1975 14040 2070
rect 14160 1975 14390 2070
rect 19410 1975 19640 2070
rect 19760 1975 19990 2070
rect 20110 1975 20340 2070
rect 20460 1975 20690 2070
rect 20810 1975 21040 2070
rect 13550 1855 13600 1975
rect 20200 1855 20250 1975
rect 12760 1770 12990 1855
rect 13110 1770 13340 1855
rect 13460 1770 13690 1855
rect 13810 1770 14040 1855
rect 14160 1770 14390 1855
rect 12760 1720 14390 1770
rect 12760 1625 12990 1720
rect 13110 1625 13340 1720
rect 13460 1625 13690 1720
rect 13810 1625 14040 1720
rect 14160 1625 14390 1720
rect 19410 1770 19640 1855
rect 19760 1770 19990 1855
rect 20110 1770 20340 1855
rect 20460 1770 20690 1855
rect 20810 1770 21040 1855
rect 19410 1720 21040 1770
rect 19410 1625 19640 1720
rect 19760 1625 19990 1720
rect 20110 1625 20340 1720
rect 20460 1625 20690 1720
rect 20810 1625 21040 1720
rect 13550 1505 13600 1625
rect 20200 1505 20250 1625
rect 5550 1470 5555 1500
rect 5585 1470 5590 1500
rect -115 660 -65 665
rect -115 620 -110 660
rect -70 620 -65 660
rect -115 615 -65 620
rect 5460 660 5510 665
rect 5460 620 5465 660
rect 5505 620 5510 660
rect 5460 615 5510 620
rect 5550 585 5590 1470
rect 12760 1420 12990 1505
rect 13110 1420 13340 1505
rect 13460 1420 13690 1505
rect 13810 1420 14040 1505
rect 14160 1420 14390 1505
rect 12760 1370 14390 1420
rect 12760 1275 12990 1370
rect 13110 1275 13340 1370
rect 13460 1275 13690 1370
rect 13810 1275 14040 1370
rect 14160 1275 14390 1370
rect 19410 1420 19640 1505
rect 19760 1420 19990 1505
rect 20110 1420 20340 1505
rect 20460 1420 20690 1505
rect 20810 1420 21040 1505
rect 19410 1370 21040 1420
rect 19410 1275 19640 1370
rect 19760 1275 19990 1370
rect 20110 1275 20340 1370
rect 20460 1275 20690 1370
rect 20810 1275 21040 1370
rect 13550 1155 13600 1275
rect 20200 1155 20250 1275
rect 12760 1070 12990 1155
rect 13110 1070 13340 1155
rect 13460 1070 13690 1155
rect 13810 1070 14040 1155
rect 14160 1070 14390 1155
rect 12760 1020 14390 1070
rect 12760 925 12990 1020
rect 13110 925 13340 1020
rect 13460 925 13690 1020
rect 13810 925 14040 1020
rect 14160 925 14390 1020
rect 19410 1070 19640 1155
rect 19760 1070 19990 1155
rect 20110 1070 20340 1155
rect 20460 1070 20690 1155
rect 20810 1070 21040 1155
rect 19410 1020 21040 1070
rect 19410 925 19640 1020
rect 19760 925 19990 1020
rect 20110 925 20340 1020
rect 20460 925 20690 1020
rect 20810 925 21040 1020
rect 13550 805 13600 925
rect 20200 805 20250 925
rect 12760 720 12990 805
rect 13110 720 13340 805
rect 13460 720 13690 805
rect 13810 720 14040 805
rect 14160 720 14390 805
rect 12760 670 14390 720
rect -200 580 -150 585
rect -200 540 -195 580
rect -155 540 -150 580
rect -200 535 -150 540
rect 5545 580 5595 585
rect 5545 540 5550 580
rect 5590 540 5595 580
rect 12760 575 12990 670
rect 13110 575 13340 670
rect 13460 575 13690 670
rect 13810 575 14040 670
rect 14160 575 14390 670
rect 19410 720 19640 805
rect 19760 720 19990 805
rect 20110 720 20340 805
rect 20460 720 20690 805
rect 20810 720 21040 805
rect 19410 670 21040 720
rect 19410 575 19640 670
rect 19760 575 19990 670
rect 20110 575 20340 670
rect 20460 575 20690 670
rect 20810 575 21040 670
rect 5545 535 5595 540
rect 13550 455 13600 575
rect 20200 455 20250 575
rect 12760 370 12990 455
rect 13110 370 13340 455
rect 13460 370 13690 455
rect 12760 320 13690 370
rect 12760 225 12990 320
rect 13110 225 13340 320
rect 13460 225 13690 320
rect 13810 225 14040 455
rect 14160 225 14390 455
rect 14510 225 14740 455
rect 14860 225 15090 455
rect 15210 225 15440 455
rect 15560 225 15790 455
rect 15910 225 16140 455
rect 16260 225 16490 455
rect 16610 225 16840 455
rect 16960 225 17190 455
rect 17310 225 17540 455
rect 17660 225 17890 455
rect 18010 225 18240 455
rect 18360 225 18590 455
rect 18710 225 18940 455
rect 19060 225 19290 455
rect 19410 225 19640 455
rect 19760 225 19990 455
rect 20110 370 20340 455
rect 20460 370 20690 455
rect 20810 370 21040 455
rect 20110 320 21040 370
rect 20110 225 20340 320
rect 20460 225 20690 320
rect 20810 225 21040 320
rect 13550 105 13600 225
rect 13900 105 13950 225
rect 14250 105 14300 225
rect 14600 105 14650 225
rect 14950 105 15000 225
rect 15300 105 15350 225
rect 15650 105 15700 225
rect 16000 105 16050 225
rect 16350 105 16400 225
rect 16700 105 16750 225
rect 17050 105 17100 225
rect 17400 105 17450 225
rect 17750 105 17800 225
rect 18100 105 18150 225
rect 18450 105 18500 225
rect 18800 105 18850 225
rect 19150 105 19200 225
rect 19500 105 19550 225
rect 19850 105 19900 225
rect 20200 105 20250 225
rect 12760 20 12990 105
rect 13110 20 13340 105
rect 13460 20 13690 105
rect 13810 20 14040 105
rect 14160 20 14390 105
rect 14510 20 14740 105
rect 14860 20 15090 105
rect 15210 20 15440 105
rect 15560 20 15790 105
rect 15910 20 16140 105
rect 16260 20 16490 105
rect 16610 20 16840 105
rect 12760 -30 16840 20
rect 12760 -125 12990 -30
rect 13110 -125 13340 -30
rect 13460 -125 13690 -30
rect 13810 -125 14040 -30
rect 14160 -125 14390 -30
rect 14510 -125 14740 -30
rect 14860 -125 15090 -30
rect 15210 -125 15440 -30
rect 15560 -125 15790 -30
rect 15910 -125 16140 -30
rect 16260 -125 16490 -30
rect 16610 -125 16840 -30
rect 16960 20 17190 105
rect 17310 20 17540 105
rect 17660 20 17890 105
rect 18010 20 18240 105
rect 18360 20 18590 105
rect 18710 20 18940 105
rect 19060 20 19290 105
rect 19410 20 19640 105
rect 19760 20 19990 105
rect 20110 20 20340 105
rect 20460 20 20690 105
rect 20810 20 21040 105
rect 16960 -30 21040 20
rect 16960 -125 17190 -30
rect 17310 -125 17540 -30
rect 17660 -125 17890 -30
rect 18010 -125 18240 -30
rect 18360 -125 18590 -30
rect 18710 -125 18940 -30
rect 19060 -125 19290 -30
rect 19410 -125 19640 -30
rect 19760 -125 19990 -30
rect 20110 -125 20340 -30
rect 20460 -125 20690 -30
rect 20810 -125 21040 -30
rect 13550 -245 13600 -125
rect 13900 -245 13950 -125
rect 14250 -245 14300 -125
rect 14600 -245 14650 -125
rect 14950 -245 15000 -125
rect 15300 -245 15350 -125
rect 15650 -245 15700 -125
rect 16000 -245 16050 -125
rect 16350 -245 16400 -125
rect 16700 -245 16750 -125
rect 17050 -245 17100 -125
rect 17400 -245 17450 -125
rect 17750 -245 17800 -125
rect 18100 -245 18150 -125
rect 18450 -245 18500 -125
rect 18800 -245 18850 -125
rect 19150 -245 19200 -125
rect 19500 -245 19550 -125
rect 19850 -245 19900 -125
rect 20200 -245 20250 -125
rect 12760 -330 12990 -245
rect 13110 -330 13340 -245
rect 13460 -330 13690 -245
rect 12760 -380 13690 -330
rect 12760 -475 12990 -380
rect 13110 -475 13340 -380
rect 13460 -475 13690 -380
rect 13810 -475 14040 -245
rect 14160 -475 14390 -245
rect 14510 -475 14740 -245
rect 14860 -475 15090 -245
rect 15210 -475 15440 -245
rect 15560 -475 15790 -245
rect 15910 -475 16140 -245
rect 16260 -475 16490 -245
rect 16610 -475 16840 -245
rect 16960 -475 17190 -245
rect 17310 -475 17540 -245
rect 17660 -475 17890 -245
rect 18010 -475 18240 -245
rect 18360 -475 18590 -245
rect 18710 -475 18940 -245
rect 19060 -475 19290 -245
rect 19410 -475 19640 -245
rect 19760 -475 19990 -245
rect 20110 -330 20340 -245
rect 20460 -330 20690 -245
rect 20810 -330 21040 -245
rect 20110 -380 21040 -330
rect 20110 -475 20340 -380
rect 20460 -475 20690 -380
rect 20810 -475 21040 -380
<< via3 >>
rect -195 4990 -155 4995
rect -195 4960 -190 4990
rect -190 4960 -160 4990
rect -160 4960 -155 4990
rect -195 4955 -155 4960
rect 5550 4990 5590 4995
rect 5550 4960 5555 4990
rect 5555 4960 5585 4990
rect 5585 4960 5590 4990
rect 5550 4955 5590 4960
rect -110 4870 -70 4910
rect 5465 4870 5505 4910
rect 1640 3445 1680 3450
rect 1640 3415 1645 3445
rect 1645 3415 1675 3445
rect 1675 3415 1680 3445
rect 1640 3410 1680 3415
rect 5140 3445 5180 3450
rect 5140 3415 5145 3445
rect 5145 3415 5175 3445
rect 5175 3415 5180 3445
rect 5140 3410 5180 3415
rect 3390 3335 3430 3340
rect 3390 3305 3395 3335
rect 3395 3305 3425 3335
rect 3425 3305 3430 3335
rect 3390 3300 3430 3305
rect 14515 2110 14555 2115
rect 14515 2080 14520 2110
rect 14520 2080 14550 2110
rect 14550 2080 14555 2110
rect 14515 2075 14555 2080
rect 19245 2110 19285 2115
rect 19245 2080 19250 2110
rect 19250 2080 19280 2110
rect 19280 2080 19285 2110
rect 19245 2075 19285 2080
rect -110 620 -70 660
rect 5465 620 5505 660
rect -195 575 -155 580
rect -195 545 -190 575
rect -190 545 -160 575
rect -160 545 -155 575
rect -195 540 -155 545
rect 5550 540 5590 580
<< mimcap >>
rect 12775 5615 12975 5690
rect 12775 5575 12855 5615
rect 12895 5575 12975 5615
rect 12775 5490 12975 5575
rect 13125 5615 13325 5690
rect 13125 5575 13205 5615
rect 13245 5575 13325 5615
rect 13125 5490 13325 5575
rect 13475 5615 13675 5690
rect 13475 5575 13555 5615
rect 13595 5575 13675 5615
rect 13475 5490 13675 5575
rect 13825 5615 14025 5690
rect 13825 5575 13905 5615
rect 13945 5575 14025 5615
rect 13825 5490 14025 5575
rect 14175 5615 14375 5690
rect 14175 5575 14255 5615
rect 14295 5575 14375 5615
rect 14175 5490 14375 5575
rect 14525 5615 14725 5690
rect 14525 5575 14605 5615
rect 14645 5575 14725 5615
rect 14525 5490 14725 5575
rect 14875 5615 15075 5690
rect 14875 5575 14955 5615
rect 14995 5575 15075 5615
rect 14875 5490 15075 5575
rect 15225 5615 15425 5690
rect 15225 5575 15305 5615
rect 15345 5575 15425 5615
rect 15225 5490 15425 5575
rect 15575 5615 15775 5690
rect 15575 5575 15655 5615
rect 15695 5575 15775 5615
rect 15575 5490 15775 5575
rect 15925 5615 16125 5690
rect 15925 5575 16005 5615
rect 16045 5575 16125 5615
rect 15925 5490 16125 5575
rect 16275 5615 16475 5690
rect 16275 5575 16355 5615
rect 16395 5575 16475 5615
rect 16275 5490 16475 5575
rect 16625 5615 16825 5690
rect 16625 5575 16705 5615
rect 16745 5575 16825 5615
rect 16625 5490 16825 5575
rect 16975 5615 17175 5690
rect 16975 5575 17055 5615
rect 17095 5575 17175 5615
rect 16975 5490 17175 5575
rect 17325 5615 17525 5690
rect 17325 5575 17405 5615
rect 17445 5575 17525 5615
rect 17325 5490 17525 5575
rect 17675 5615 17875 5690
rect 17675 5575 17755 5615
rect 17795 5575 17875 5615
rect 17675 5490 17875 5575
rect 18025 5615 18225 5690
rect 18025 5575 18105 5615
rect 18145 5575 18225 5615
rect 18025 5490 18225 5575
rect 18375 5615 18575 5690
rect 18375 5575 18455 5615
rect 18495 5575 18575 5615
rect 18375 5490 18575 5575
rect 18725 5615 18925 5690
rect 18725 5575 18805 5615
rect 18845 5575 18925 5615
rect 18725 5490 18925 5575
rect 19075 5615 19275 5690
rect 19075 5575 19155 5615
rect 19195 5575 19275 5615
rect 19075 5490 19275 5575
rect 19425 5615 19625 5690
rect 19425 5575 19505 5615
rect 19545 5575 19625 5615
rect 19425 5490 19625 5575
rect 19775 5615 19975 5690
rect 19775 5575 19855 5615
rect 19895 5575 19975 5615
rect 19775 5490 19975 5575
rect 20125 5615 20325 5690
rect 20125 5575 20205 5615
rect 20245 5575 20325 5615
rect 20125 5490 20325 5575
rect 20475 5615 20675 5690
rect 20475 5575 20555 5615
rect 20595 5575 20675 5615
rect 20475 5490 20675 5575
rect 20825 5615 21025 5690
rect 20825 5575 20905 5615
rect 20945 5575 21025 5615
rect 20825 5490 21025 5575
rect 12775 5265 12975 5340
rect 12775 5225 12855 5265
rect 12895 5225 12975 5265
rect 12775 5140 12975 5225
rect 13125 5265 13325 5340
rect 13125 5225 13205 5265
rect 13245 5225 13325 5265
rect 13125 5140 13325 5225
rect 13475 5265 13675 5340
rect 13475 5225 13555 5265
rect 13595 5225 13675 5265
rect 13475 5140 13675 5225
rect 13825 5265 14025 5340
rect 13825 5225 13905 5265
rect 13945 5225 14025 5265
rect 13825 5140 14025 5225
rect 14175 5265 14375 5340
rect 14175 5225 14255 5265
rect 14295 5225 14375 5265
rect 14175 5140 14375 5225
rect 14525 5265 14725 5340
rect 14525 5225 14605 5265
rect 14645 5225 14725 5265
rect 14525 5140 14725 5225
rect 14875 5265 15075 5340
rect 14875 5225 14955 5265
rect 14995 5225 15075 5265
rect 14875 5140 15075 5225
rect 15225 5265 15425 5340
rect 15225 5225 15305 5265
rect 15345 5225 15425 5265
rect 15225 5140 15425 5225
rect 15575 5265 15775 5340
rect 15575 5225 15655 5265
rect 15695 5225 15775 5265
rect 15575 5140 15775 5225
rect 15925 5265 16125 5340
rect 15925 5225 16005 5265
rect 16045 5225 16125 5265
rect 15925 5140 16125 5225
rect 16275 5265 16475 5340
rect 16275 5225 16355 5265
rect 16395 5225 16475 5265
rect 16275 5140 16475 5225
rect 16625 5265 16825 5340
rect 16625 5225 16705 5265
rect 16745 5225 16825 5265
rect 16625 5140 16825 5225
rect 16975 5265 17175 5340
rect 16975 5225 17055 5265
rect 17095 5225 17175 5265
rect 16975 5140 17175 5225
rect 17325 5265 17525 5340
rect 17325 5225 17405 5265
rect 17445 5225 17525 5265
rect 17325 5140 17525 5225
rect 17675 5265 17875 5340
rect 17675 5225 17755 5265
rect 17795 5225 17875 5265
rect 17675 5140 17875 5225
rect 18025 5265 18225 5340
rect 18025 5225 18105 5265
rect 18145 5225 18225 5265
rect 18025 5140 18225 5225
rect 18375 5265 18575 5340
rect 18375 5225 18455 5265
rect 18495 5225 18575 5265
rect 18375 5140 18575 5225
rect 18725 5265 18925 5340
rect 18725 5225 18805 5265
rect 18845 5225 18925 5265
rect 18725 5140 18925 5225
rect 19075 5265 19275 5340
rect 19075 5225 19155 5265
rect 19195 5225 19275 5265
rect 19075 5140 19275 5225
rect 19425 5265 19625 5340
rect 19425 5225 19505 5265
rect 19545 5225 19625 5265
rect 19425 5140 19625 5225
rect 19775 5265 19975 5340
rect 19775 5225 19855 5265
rect 19895 5225 19975 5265
rect 19775 5140 19975 5225
rect 20125 5265 20325 5340
rect 20125 5225 20205 5265
rect 20245 5225 20325 5265
rect 20125 5140 20325 5225
rect 20475 5265 20675 5340
rect 20475 5225 20555 5265
rect 20595 5225 20675 5265
rect 20475 5140 20675 5225
rect 20825 5265 21025 5340
rect 20825 5225 20905 5265
rect 20945 5225 21025 5265
rect 20825 5140 21025 5225
rect 12775 4915 12975 4990
rect 12775 4875 12855 4915
rect 12895 4875 12975 4915
rect 160 4765 360 4840
rect 160 4725 240 4765
rect 280 4725 360 4765
rect 160 4640 360 4725
rect 510 4765 710 4840
rect 510 4725 590 4765
rect 630 4725 710 4765
rect 510 4640 710 4725
rect 860 4765 1060 4840
rect 860 4725 940 4765
rect 980 4725 1060 4765
rect 860 4640 1060 4725
rect 1210 4765 1410 4840
rect 1210 4725 1290 4765
rect 1330 4725 1410 4765
rect 1210 4640 1410 4725
rect 1560 4765 1760 4840
rect 1560 4725 1640 4765
rect 1680 4725 1760 4765
rect 1560 4640 1760 4725
rect 1910 4765 2110 4840
rect 1910 4725 1990 4765
rect 2030 4725 2110 4765
rect 1910 4640 2110 4725
rect 2260 4765 2460 4840
rect 2260 4725 2340 4765
rect 2380 4725 2460 4765
rect 2260 4640 2460 4725
rect 2610 4765 2810 4840
rect 2610 4725 2690 4765
rect 2730 4725 2810 4765
rect 2610 4640 2810 4725
rect 2960 4765 3160 4840
rect 2960 4725 3040 4765
rect 3080 4725 3160 4765
rect 2960 4640 3160 4725
rect 3310 4765 3510 4840
rect 3310 4725 3390 4765
rect 3430 4725 3510 4765
rect 3310 4640 3510 4725
rect 3660 4765 3860 4840
rect 3660 4725 3740 4765
rect 3780 4725 3860 4765
rect 3660 4640 3860 4725
rect 4010 4765 4210 4840
rect 4010 4725 4090 4765
rect 4130 4725 4210 4765
rect 4010 4640 4210 4725
rect 4360 4765 4560 4840
rect 4360 4725 4440 4765
rect 4480 4725 4560 4765
rect 4360 4640 4560 4725
rect 4710 4765 4910 4840
rect 4710 4725 4790 4765
rect 4830 4725 4910 4765
rect 4710 4640 4910 4725
rect 5060 4765 5260 4840
rect 12775 4790 12975 4875
rect 13125 4915 13325 4990
rect 13125 4875 13205 4915
rect 13245 4875 13325 4915
rect 13125 4790 13325 4875
rect 13475 4915 13675 4990
rect 13475 4875 13555 4915
rect 13595 4875 13675 4915
rect 13475 4790 13675 4875
rect 13825 4915 14025 4990
rect 13825 4875 13905 4915
rect 13945 4875 14025 4915
rect 13825 4790 14025 4875
rect 14175 4915 14375 4990
rect 14175 4875 14255 4915
rect 14295 4875 14375 4915
rect 14175 4790 14375 4875
rect 14525 4915 14725 4990
rect 14525 4875 14605 4915
rect 14645 4875 14725 4915
rect 14525 4790 14725 4875
rect 14875 4915 15075 4990
rect 14875 4875 14955 4915
rect 14995 4875 15075 4915
rect 14875 4790 15075 4875
rect 15225 4915 15425 4990
rect 15225 4875 15305 4915
rect 15345 4875 15425 4915
rect 15225 4790 15425 4875
rect 15575 4915 15775 4990
rect 15575 4875 15655 4915
rect 15695 4875 15775 4915
rect 15575 4790 15775 4875
rect 15925 4915 16125 4990
rect 15925 4875 16005 4915
rect 16045 4875 16125 4915
rect 15925 4790 16125 4875
rect 16275 4915 16475 4990
rect 16275 4875 16355 4915
rect 16395 4875 16475 4915
rect 16275 4790 16475 4875
rect 16625 4915 16825 4990
rect 16625 4875 16705 4915
rect 16745 4875 16825 4915
rect 16625 4790 16825 4875
rect 16975 4915 17175 4990
rect 16975 4875 17055 4915
rect 17095 4875 17175 4915
rect 16975 4790 17175 4875
rect 17325 4915 17525 4990
rect 17325 4875 17405 4915
rect 17445 4875 17525 4915
rect 17325 4790 17525 4875
rect 17675 4915 17875 4990
rect 17675 4875 17755 4915
rect 17795 4875 17875 4915
rect 17675 4790 17875 4875
rect 18025 4915 18225 4990
rect 18025 4875 18105 4915
rect 18145 4875 18225 4915
rect 18025 4790 18225 4875
rect 18375 4915 18575 4990
rect 18375 4875 18455 4915
rect 18495 4875 18575 4915
rect 18375 4790 18575 4875
rect 18725 4915 18925 4990
rect 18725 4875 18805 4915
rect 18845 4875 18925 4915
rect 18725 4790 18925 4875
rect 19075 4915 19275 4990
rect 19075 4875 19155 4915
rect 19195 4875 19275 4915
rect 19075 4790 19275 4875
rect 19425 4915 19625 4990
rect 19425 4875 19505 4915
rect 19545 4875 19625 4915
rect 19425 4790 19625 4875
rect 19775 4915 19975 4990
rect 19775 4875 19855 4915
rect 19895 4875 19975 4915
rect 19775 4790 19975 4875
rect 20125 4915 20325 4990
rect 20125 4875 20205 4915
rect 20245 4875 20325 4915
rect 20125 4790 20325 4875
rect 20475 4915 20675 4990
rect 20475 4875 20555 4915
rect 20595 4875 20675 4915
rect 20475 4790 20675 4875
rect 20825 4915 21025 4990
rect 20825 4875 20905 4915
rect 20945 4875 21025 4915
rect 20825 4790 21025 4875
rect 5060 4725 5140 4765
rect 5180 4725 5260 4765
rect 5060 4640 5260 4725
rect 12775 4565 12975 4640
rect 12775 4525 12855 4565
rect 12895 4525 12975 4565
rect 160 4415 360 4490
rect 160 4375 240 4415
rect 280 4375 360 4415
rect 160 4290 360 4375
rect 510 4415 710 4490
rect 510 4375 590 4415
rect 630 4375 710 4415
rect 510 4290 710 4375
rect 860 4415 1060 4490
rect 860 4375 940 4415
rect 980 4375 1060 4415
rect 860 4290 1060 4375
rect 1210 4415 1410 4490
rect 1210 4375 1290 4415
rect 1330 4375 1410 4415
rect 1210 4290 1410 4375
rect 1560 4415 1760 4490
rect 1560 4375 1640 4415
rect 1680 4375 1760 4415
rect 1560 4290 1760 4375
rect 1910 4415 2110 4490
rect 1910 4375 1990 4415
rect 2030 4375 2110 4415
rect 1910 4290 2110 4375
rect 2260 4415 2460 4490
rect 2260 4375 2340 4415
rect 2380 4375 2460 4415
rect 2260 4290 2460 4375
rect 2610 4415 2810 4490
rect 2610 4375 2690 4415
rect 2730 4375 2810 4415
rect 2610 4290 2810 4375
rect 2960 4415 3160 4490
rect 2960 4375 3040 4415
rect 3080 4375 3160 4415
rect 2960 4290 3160 4375
rect 3310 4415 3510 4490
rect 3310 4375 3390 4415
rect 3430 4375 3510 4415
rect 3310 4290 3510 4375
rect 3660 4415 3860 4490
rect 3660 4375 3740 4415
rect 3780 4375 3860 4415
rect 3660 4290 3860 4375
rect 4010 4415 4210 4490
rect 4010 4375 4090 4415
rect 4130 4375 4210 4415
rect 4010 4290 4210 4375
rect 4360 4415 4560 4490
rect 4360 4375 4440 4415
rect 4480 4375 4560 4415
rect 4360 4290 4560 4375
rect 4710 4415 4910 4490
rect 4710 4375 4790 4415
rect 4830 4375 4910 4415
rect 4710 4290 4910 4375
rect 5060 4415 5260 4490
rect 12775 4440 12975 4525
rect 13125 4565 13325 4640
rect 13125 4525 13205 4565
rect 13245 4525 13325 4565
rect 13125 4440 13325 4525
rect 13475 4565 13675 4640
rect 13475 4525 13555 4565
rect 13595 4525 13675 4565
rect 13475 4440 13675 4525
rect 13825 4565 14025 4640
rect 13825 4525 13905 4565
rect 13945 4525 14025 4565
rect 13825 4440 14025 4525
rect 14175 4565 14375 4640
rect 14175 4525 14255 4565
rect 14295 4525 14375 4565
rect 14175 4440 14375 4525
rect 14525 4565 14725 4640
rect 14525 4525 14605 4565
rect 14645 4525 14725 4565
rect 14525 4440 14725 4525
rect 14875 4565 15075 4640
rect 14875 4525 14955 4565
rect 14995 4525 15075 4565
rect 14875 4440 15075 4525
rect 15225 4565 15425 4640
rect 15225 4525 15305 4565
rect 15345 4525 15425 4565
rect 15225 4440 15425 4525
rect 15575 4565 15775 4640
rect 15575 4525 15655 4565
rect 15695 4525 15775 4565
rect 15575 4440 15775 4525
rect 18025 4565 18225 4640
rect 18025 4525 18105 4565
rect 18145 4525 18225 4565
rect 18025 4440 18225 4525
rect 18375 4565 18575 4640
rect 18375 4525 18455 4565
rect 18495 4525 18575 4565
rect 18375 4440 18575 4525
rect 18725 4565 18925 4640
rect 18725 4525 18805 4565
rect 18845 4525 18925 4565
rect 18725 4440 18925 4525
rect 19075 4565 19275 4640
rect 19075 4525 19155 4565
rect 19195 4525 19275 4565
rect 19075 4440 19275 4525
rect 19425 4565 19625 4640
rect 19425 4525 19505 4565
rect 19545 4525 19625 4565
rect 19425 4440 19625 4525
rect 19775 4565 19975 4640
rect 19775 4525 19855 4565
rect 19895 4525 19975 4565
rect 19775 4440 19975 4525
rect 20125 4565 20325 4640
rect 20125 4525 20205 4565
rect 20245 4525 20325 4565
rect 20125 4440 20325 4525
rect 20475 4565 20675 4640
rect 20475 4525 20555 4565
rect 20595 4525 20675 4565
rect 20475 4440 20675 4525
rect 20825 4565 21025 4640
rect 20825 4525 20905 4565
rect 20945 4525 21025 4565
rect 20825 4440 21025 4525
rect 5060 4375 5140 4415
rect 5180 4375 5260 4415
rect 5060 4290 5260 4375
rect 12775 4215 12975 4290
rect 12775 4175 12855 4215
rect 12895 4175 12975 4215
rect 160 4065 360 4140
rect 160 4025 240 4065
rect 280 4025 360 4065
rect 160 3940 360 4025
rect 510 4065 710 4140
rect 510 4025 590 4065
rect 630 4025 710 4065
rect 510 3940 710 4025
rect 860 4065 1060 4140
rect 860 4025 940 4065
rect 980 4025 1060 4065
rect 860 3940 1060 4025
rect 1210 4065 1410 4140
rect 1210 4025 1290 4065
rect 1330 4025 1410 4065
rect 1210 3940 1410 4025
rect 1560 4065 1760 4140
rect 1560 4025 1640 4065
rect 1680 4025 1760 4065
rect 1560 3940 1760 4025
rect 1910 4065 2110 4140
rect 1910 4025 1990 4065
rect 2030 4025 2110 4065
rect 1910 3940 2110 4025
rect 2260 4065 2460 4140
rect 2260 4025 2340 4065
rect 2380 4025 2460 4065
rect 2260 3940 2460 4025
rect 2610 4065 2810 4140
rect 2610 4025 2690 4065
rect 2730 4025 2810 4065
rect 2610 3940 2810 4025
rect 2960 4065 3160 4140
rect 2960 4025 3040 4065
rect 3080 4025 3160 4065
rect 2960 3940 3160 4025
rect 3310 4065 3510 4140
rect 3310 4025 3390 4065
rect 3430 4025 3510 4065
rect 3310 3940 3510 4025
rect 3660 4065 3860 4140
rect 3660 4025 3740 4065
rect 3780 4025 3860 4065
rect 3660 3940 3860 4025
rect 4010 4065 4210 4140
rect 4010 4025 4090 4065
rect 4130 4025 4210 4065
rect 4010 3940 4210 4025
rect 4360 4065 4560 4140
rect 4360 4025 4440 4065
rect 4480 4025 4560 4065
rect 4360 3940 4560 4025
rect 4710 4065 4910 4140
rect 4710 4025 4790 4065
rect 4830 4025 4910 4065
rect 4710 3940 4910 4025
rect 5060 4065 5260 4140
rect 12775 4090 12975 4175
rect 13125 4215 13325 4290
rect 13125 4175 13205 4215
rect 13245 4175 13325 4215
rect 13125 4090 13325 4175
rect 13475 4215 13675 4290
rect 13475 4175 13555 4215
rect 13595 4175 13675 4215
rect 13475 4090 13675 4175
rect 13825 4215 14025 4290
rect 13825 4175 13905 4215
rect 13945 4175 14025 4215
rect 13825 4090 14025 4175
rect 14175 4215 14375 4290
rect 14175 4175 14255 4215
rect 14295 4175 14375 4215
rect 14175 4090 14375 4175
rect 14525 4215 14725 4290
rect 14525 4175 14605 4215
rect 14645 4175 14725 4215
rect 14525 4090 14725 4175
rect 14875 4215 15075 4290
rect 14875 4175 14955 4215
rect 14995 4175 15075 4215
rect 14875 4090 15075 4175
rect 15225 4215 15425 4290
rect 15225 4175 15305 4215
rect 15345 4175 15425 4215
rect 15225 4090 15425 4175
rect 15575 4215 15775 4290
rect 15575 4175 15655 4215
rect 15695 4175 15775 4215
rect 15575 4090 15775 4175
rect 18025 4215 18225 4290
rect 18025 4175 18105 4215
rect 18145 4175 18225 4215
rect 18025 4090 18225 4175
rect 18375 4215 18575 4290
rect 18375 4175 18455 4215
rect 18495 4175 18575 4215
rect 18375 4090 18575 4175
rect 18725 4215 18925 4290
rect 18725 4175 18805 4215
rect 18845 4175 18925 4215
rect 18725 4090 18925 4175
rect 19075 4215 19275 4290
rect 19075 4175 19155 4215
rect 19195 4175 19275 4215
rect 19075 4090 19275 4175
rect 19425 4215 19625 4290
rect 19425 4175 19505 4215
rect 19545 4175 19625 4215
rect 19425 4090 19625 4175
rect 19775 4215 19975 4290
rect 19775 4175 19855 4215
rect 19895 4175 19975 4215
rect 19775 4090 19975 4175
rect 20125 4215 20325 4290
rect 20125 4175 20205 4215
rect 20245 4175 20325 4215
rect 20125 4090 20325 4175
rect 20475 4215 20675 4290
rect 20475 4175 20555 4215
rect 20595 4175 20675 4215
rect 20475 4090 20675 4175
rect 20825 4215 21025 4290
rect 20825 4175 20905 4215
rect 20945 4175 21025 4215
rect 20825 4090 21025 4175
rect 5060 4025 5140 4065
rect 5180 4025 5260 4065
rect 5060 3940 5260 4025
rect 12775 3865 12975 3940
rect 12775 3825 12855 3865
rect 12895 3825 12975 3865
rect 160 3715 360 3790
rect 160 3675 240 3715
rect 280 3675 360 3715
rect 160 3590 360 3675
rect 510 3715 710 3790
rect 510 3675 590 3715
rect 630 3675 710 3715
rect 510 3590 710 3675
rect 860 3715 1060 3790
rect 860 3675 940 3715
rect 980 3675 1060 3715
rect 860 3590 1060 3675
rect 1210 3715 1410 3790
rect 1210 3675 1290 3715
rect 1330 3675 1410 3715
rect 1210 3590 1410 3675
rect 1560 3715 1760 3790
rect 1560 3675 1640 3715
rect 1680 3675 1760 3715
rect 1560 3590 1760 3675
rect 1910 3715 2110 3790
rect 1910 3675 1990 3715
rect 2030 3675 2110 3715
rect 1910 3590 2110 3675
rect 2260 3715 2460 3790
rect 2260 3675 2340 3715
rect 2380 3675 2460 3715
rect 2260 3590 2460 3675
rect 2610 3715 2810 3790
rect 2610 3675 2690 3715
rect 2730 3675 2810 3715
rect 2610 3590 2810 3675
rect 2960 3715 3160 3790
rect 2960 3675 3040 3715
rect 3080 3675 3160 3715
rect 2960 3590 3160 3675
rect 3310 3715 3510 3790
rect 3310 3675 3390 3715
rect 3430 3675 3510 3715
rect 3310 3590 3510 3675
rect 3660 3715 3860 3790
rect 3660 3675 3740 3715
rect 3780 3675 3860 3715
rect 3660 3590 3860 3675
rect 4010 3715 4210 3790
rect 4010 3675 4090 3715
rect 4130 3675 4210 3715
rect 4010 3590 4210 3675
rect 4360 3715 4560 3790
rect 4360 3675 4440 3715
rect 4480 3675 4560 3715
rect 4360 3590 4560 3675
rect 4710 3715 4910 3790
rect 4710 3675 4790 3715
rect 4830 3675 4910 3715
rect 4710 3590 4910 3675
rect 5060 3715 5260 3790
rect 12775 3740 12975 3825
rect 13125 3865 13325 3940
rect 13125 3825 13205 3865
rect 13245 3825 13325 3865
rect 13125 3740 13325 3825
rect 13475 3865 13675 3940
rect 13475 3825 13555 3865
rect 13595 3825 13675 3865
rect 13475 3740 13675 3825
rect 13825 3865 14025 3940
rect 13825 3825 13905 3865
rect 13945 3825 14025 3865
rect 13825 3740 14025 3825
rect 14175 3865 14375 3940
rect 14175 3825 14255 3865
rect 14295 3825 14375 3865
rect 14175 3740 14375 3825
rect 14525 3865 14725 3940
rect 14525 3825 14605 3865
rect 14645 3825 14725 3865
rect 14525 3740 14725 3825
rect 14875 3865 15075 3940
rect 14875 3825 14955 3865
rect 14995 3825 15075 3865
rect 14875 3740 15075 3825
rect 15225 3865 15425 3940
rect 15225 3825 15305 3865
rect 15345 3825 15425 3865
rect 15225 3740 15425 3825
rect 15575 3865 15775 3940
rect 15575 3825 15655 3865
rect 15695 3825 15775 3865
rect 15575 3740 15775 3825
rect 18025 3865 18225 3940
rect 18025 3825 18105 3865
rect 18145 3825 18225 3865
rect 18025 3740 18225 3825
rect 18375 3865 18575 3940
rect 18375 3825 18455 3865
rect 18495 3825 18575 3865
rect 18375 3740 18575 3825
rect 18725 3865 18925 3940
rect 18725 3825 18805 3865
rect 18845 3825 18925 3865
rect 18725 3740 18925 3825
rect 19075 3865 19275 3940
rect 19075 3825 19155 3865
rect 19195 3825 19275 3865
rect 19075 3740 19275 3825
rect 19425 3865 19625 3940
rect 19425 3825 19505 3865
rect 19545 3825 19625 3865
rect 19425 3740 19625 3825
rect 19775 3865 19975 3940
rect 19775 3825 19855 3865
rect 19895 3825 19975 3865
rect 19775 3740 19975 3825
rect 20125 3865 20325 3940
rect 20125 3825 20205 3865
rect 20245 3825 20325 3865
rect 20125 3740 20325 3825
rect 20475 3865 20675 3940
rect 20475 3825 20555 3865
rect 20595 3825 20675 3865
rect 20475 3740 20675 3825
rect 20825 3865 21025 3940
rect 20825 3825 20905 3865
rect 20945 3825 21025 3865
rect 20825 3740 21025 3825
rect 5060 3675 5140 3715
rect 5180 3675 5260 3715
rect 5060 3590 5260 3675
rect 12775 3515 12975 3590
rect 12775 3475 12855 3515
rect 12895 3475 12975 3515
rect 12775 3390 12975 3475
rect 13125 3515 13325 3590
rect 13125 3475 13205 3515
rect 13245 3475 13325 3515
rect 13125 3390 13325 3475
rect 13475 3515 13675 3590
rect 13475 3475 13555 3515
rect 13595 3475 13675 3515
rect 13475 3390 13675 3475
rect 13825 3515 14025 3590
rect 13825 3475 13905 3515
rect 13945 3475 14025 3515
rect 13825 3390 14025 3475
rect 14175 3515 14375 3590
rect 14175 3475 14255 3515
rect 14295 3475 14375 3515
rect 14175 3390 14375 3475
rect 19425 3515 19625 3590
rect 19425 3475 19505 3515
rect 19545 3475 19625 3515
rect 19425 3390 19625 3475
rect 19775 3515 19975 3590
rect 19775 3475 19855 3515
rect 19895 3475 19975 3515
rect 19775 3390 19975 3475
rect 20125 3515 20325 3590
rect 20125 3475 20205 3515
rect 20245 3475 20325 3515
rect 20125 3390 20325 3475
rect 20475 3515 20675 3590
rect 20475 3475 20555 3515
rect 20595 3475 20675 3515
rect 20475 3390 20675 3475
rect 20825 3515 21025 3590
rect 20825 3475 20905 3515
rect 20945 3475 21025 3515
rect 20825 3390 21025 3475
rect 12775 3165 12975 3240
rect 12775 3125 12855 3165
rect 12895 3125 12975 3165
rect 12775 3040 12975 3125
rect 13125 3165 13325 3240
rect 13125 3125 13205 3165
rect 13245 3125 13325 3165
rect 13125 3040 13325 3125
rect 13475 3165 13675 3240
rect 13475 3125 13555 3165
rect 13595 3125 13675 3165
rect 13475 3040 13675 3125
rect 13825 3165 14025 3240
rect 13825 3125 13905 3165
rect 13945 3125 14025 3165
rect 13825 3040 14025 3125
rect 14175 3165 14375 3240
rect 14175 3125 14255 3165
rect 14295 3125 14375 3165
rect 14175 3040 14375 3125
rect 19425 3165 19625 3240
rect 19425 3125 19505 3165
rect 19545 3125 19625 3165
rect 19425 3040 19625 3125
rect 19775 3165 19975 3240
rect 19775 3125 19855 3165
rect 19895 3125 19975 3165
rect 19775 3040 19975 3125
rect 20125 3165 20325 3240
rect 20125 3125 20205 3165
rect 20245 3125 20325 3165
rect 20125 3040 20325 3125
rect 20475 3165 20675 3240
rect 20475 3125 20555 3165
rect 20595 3125 20675 3165
rect 20475 3040 20675 3125
rect 20825 3165 21025 3240
rect 20825 3125 20905 3165
rect 20945 3125 21025 3165
rect 20825 3040 21025 3125
rect 12775 2815 12975 2890
rect 12775 2775 12855 2815
rect 12895 2775 12975 2815
rect 12775 2690 12975 2775
rect 13125 2815 13325 2890
rect 13125 2775 13205 2815
rect 13245 2775 13325 2815
rect 13125 2690 13325 2775
rect 13475 2815 13675 2890
rect 13475 2775 13555 2815
rect 13595 2775 13675 2815
rect 13475 2690 13675 2775
rect 13825 2815 14025 2890
rect 13825 2775 13905 2815
rect 13945 2775 14025 2815
rect 13825 2690 14025 2775
rect 14175 2815 14375 2890
rect 14175 2775 14255 2815
rect 14295 2775 14375 2815
rect 14175 2690 14375 2775
rect 19425 2815 19625 2890
rect 19425 2775 19505 2815
rect 19545 2775 19625 2815
rect 19425 2690 19625 2775
rect 19775 2815 19975 2890
rect 19775 2775 19855 2815
rect 19895 2775 19975 2815
rect 19775 2690 19975 2775
rect 20125 2815 20325 2890
rect 20125 2775 20205 2815
rect 20245 2775 20325 2815
rect 20125 2690 20325 2775
rect 20475 2815 20675 2890
rect 20475 2775 20555 2815
rect 20595 2775 20675 2815
rect 20475 2690 20675 2775
rect 20825 2815 21025 2890
rect 20825 2775 20905 2815
rect 20945 2775 21025 2815
rect 20825 2690 21025 2775
rect 12775 2465 12975 2540
rect 12775 2425 12855 2465
rect 12895 2425 12975 2465
rect 12775 2340 12975 2425
rect 13125 2465 13325 2540
rect 13125 2425 13205 2465
rect 13245 2425 13325 2465
rect 13125 2340 13325 2425
rect 13475 2465 13675 2540
rect 13475 2425 13555 2465
rect 13595 2425 13675 2465
rect 13475 2340 13675 2425
rect 13825 2465 14025 2540
rect 13825 2425 13905 2465
rect 13945 2425 14025 2465
rect 13825 2340 14025 2425
rect 14175 2465 14375 2540
rect 14175 2425 14255 2465
rect 14295 2425 14375 2465
rect 14175 2340 14375 2425
rect 19425 2465 19625 2540
rect 19425 2425 19505 2465
rect 19545 2425 19625 2465
rect 19425 2340 19625 2425
rect 19775 2465 19975 2540
rect 19775 2425 19855 2465
rect 19895 2425 19975 2465
rect 19775 2340 19975 2425
rect 20125 2465 20325 2540
rect 20125 2425 20205 2465
rect 20245 2425 20325 2465
rect 20125 2340 20325 2425
rect 20475 2465 20675 2540
rect 20475 2425 20555 2465
rect 20595 2425 20675 2465
rect 20475 2340 20675 2425
rect 20825 2465 21025 2540
rect 20825 2425 20905 2465
rect 20945 2425 21025 2465
rect 20825 2340 21025 2425
rect 12775 2115 12975 2190
rect 12775 2075 12855 2115
rect 12895 2075 12975 2115
rect 12775 1990 12975 2075
rect 13125 2115 13325 2190
rect 13125 2075 13205 2115
rect 13245 2075 13325 2115
rect 13125 1990 13325 2075
rect 13475 2115 13675 2190
rect 13475 2075 13555 2115
rect 13595 2075 13675 2115
rect 13475 1990 13675 2075
rect 13825 2115 14025 2190
rect 13825 2075 13905 2115
rect 13945 2075 14025 2115
rect 13825 1990 14025 2075
rect 14175 2115 14375 2190
rect 14175 2075 14255 2115
rect 14295 2075 14375 2115
rect 14175 1990 14375 2075
rect 19425 2115 19625 2190
rect 19425 2075 19505 2115
rect 19545 2075 19625 2115
rect 19425 1990 19625 2075
rect 19775 2115 19975 2190
rect 19775 2075 19855 2115
rect 19895 2075 19975 2115
rect 19775 1990 19975 2075
rect 20125 2115 20325 2190
rect 20125 2075 20205 2115
rect 20245 2075 20325 2115
rect 20125 1990 20325 2075
rect 20475 2115 20675 2190
rect 20475 2075 20555 2115
rect 20595 2075 20675 2115
rect 20475 1990 20675 2075
rect 20825 2115 21025 2190
rect 20825 2075 20905 2115
rect 20945 2075 21025 2115
rect 20825 1990 21025 2075
rect 12775 1765 12975 1840
rect 12775 1725 12855 1765
rect 12895 1725 12975 1765
rect 12775 1640 12975 1725
rect 13125 1765 13325 1840
rect 13125 1725 13205 1765
rect 13245 1725 13325 1765
rect 13125 1640 13325 1725
rect 13475 1765 13675 1840
rect 13475 1725 13555 1765
rect 13595 1725 13675 1765
rect 13475 1640 13675 1725
rect 13825 1765 14025 1840
rect 13825 1725 13905 1765
rect 13945 1725 14025 1765
rect 13825 1640 14025 1725
rect 14175 1765 14375 1840
rect 14175 1725 14255 1765
rect 14295 1725 14375 1765
rect 14175 1640 14375 1725
rect 19425 1765 19625 1840
rect 19425 1725 19505 1765
rect 19545 1725 19625 1765
rect 19425 1640 19625 1725
rect 19775 1765 19975 1840
rect 19775 1725 19855 1765
rect 19895 1725 19975 1765
rect 19775 1640 19975 1725
rect 20125 1765 20325 1840
rect 20125 1725 20205 1765
rect 20245 1725 20325 1765
rect 20125 1640 20325 1725
rect 20475 1765 20675 1840
rect 20475 1725 20555 1765
rect 20595 1725 20675 1765
rect 20475 1640 20675 1725
rect 20825 1765 21025 1840
rect 20825 1725 20905 1765
rect 20945 1725 21025 1765
rect 20825 1640 21025 1725
rect 12775 1415 12975 1490
rect 12775 1375 12855 1415
rect 12895 1375 12975 1415
rect 12775 1290 12975 1375
rect 13125 1415 13325 1490
rect 13125 1375 13205 1415
rect 13245 1375 13325 1415
rect 13125 1290 13325 1375
rect 13475 1415 13675 1490
rect 13475 1375 13555 1415
rect 13595 1375 13675 1415
rect 13475 1290 13675 1375
rect 13825 1415 14025 1490
rect 13825 1375 13905 1415
rect 13945 1375 14025 1415
rect 13825 1290 14025 1375
rect 14175 1415 14375 1490
rect 14175 1375 14255 1415
rect 14295 1375 14375 1415
rect 14175 1290 14375 1375
rect 19425 1415 19625 1490
rect 19425 1375 19505 1415
rect 19545 1375 19625 1415
rect 19425 1290 19625 1375
rect 19775 1415 19975 1490
rect 19775 1375 19855 1415
rect 19895 1375 19975 1415
rect 19775 1290 19975 1375
rect 20125 1415 20325 1490
rect 20125 1375 20205 1415
rect 20245 1375 20325 1415
rect 20125 1290 20325 1375
rect 20475 1415 20675 1490
rect 20475 1375 20555 1415
rect 20595 1375 20675 1415
rect 20475 1290 20675 1375
rect 20825 1415 21025 1490
rect 20825 1375 20905 1415
rect 20945 1375 21025 1415
rect 20825 1290 21025 1375
rect 12775 1065 12975 1140
rect 12775 1025 12855 1065
rect 12895 1025 12975 1065
rect 12775 940 12975 1025
rect 13125 1065 13325 1140
rect 13125 1025 13205 1065
rect 13245 1025 13325 1065
rect 13125 940 13325 1025
rect 13475 1065 13675 1140
rect 13475 1025 13555 1065
rect 13595 1025 13675 1065
rect 13475 940 13675 1025
rect 13825 1065 14025 1140
rect 13825 1025 13905 1065
rect 13945 1025 14025 1065
rect 13825 940 14025 1025
rect 14175 1065 14375 1140
rect 14175 1025 14255 1065
rect 14295 1025 14375 1065
rect 14175 940 14375 1025
rect 19425 1065 19625 1140
rect 19425 1025 19505 1065
rect 19545 1025 19625 1065
rect 19425 940 19625 1025
rect 19775 1065 19975 1140
rect 19775 1025 19855 1065
rect 19895 1025 19975 1065
rect 19775 940 19975 1025
rect 20125 1065 20325 1140
rect 20125 1025 20205 1065
rect 20245 1025 20325 1065
rect 20125 940 20325 1025
rect 20475 1065 20675 1140
rect 20475 1025 20555 1065
rect 20595 1025 20675 1065
rect 20475 940 20675 1025
rect 20825 1065 21025 1140
rect 20825 1025 20905 1065
rect 20945 1025 21025 1065
rect 20825 940 21025 1025
rect 12775 715 12975 790
rect 12775 675 12855 715
rect 12895 675 12975 715
rect 12775 590 12975 675
rect 13125 715 13325 790
rect 13125 675 13205 715
rect 13245 675 13325 715
rect 13125 590 13325 675
rect 13475 715 13675 790
rect 13475 675 13555 715
rect 13595 675 13675 715
rect 13475 590 13675 675
rect 13825 715 14025 790
rect 13825 675 13905 715
rect 13945 675 14025 715
rect 13825 590 14025 675
rect 14175 715 14375 790
rect 14175 675 14255 715
rect 14295 675 14375 715
rect 14175 590 14375 675
rect 19425 715 19625 790
rect 19425 675 19505 715
rect 19545 675 19625 715
rect 19425 590 19625 675
rect 19775 715 19975 790
rect 19775 675 19855 715
rect 19895 675 19975 715
rect 19775 590 19975 675
rect 20125 715 20325 790
rect 20125 675 20205 715
rect 20245 675 20325 715
rect 20125 590 20325 675
rect 20475 715 20675 790
rect 20475 675 20555 715
rect 20595 675 20675 715
rect 20475 590 20675 675
rect 20825 715 21025 790
rect 20825 675 20905 715
rect 20945 675 21025 715
rect 20825 590 21025 675
rect 12775 365 12975 440
rect 12775 325 12855 365
rect 12895 325 12975 365
rect 12775 240 12975 325
rect 13125 365 13325 440
rect 13125 325 13205 365
rect 13245 325 13325 365
rect 13125 240 13325 325
rect 13475 365 13675 440
rect 13475 325 13555 365
rect 13595 325 13675 365
rect 13475 240 13675 325
rect 13825 365 14025 440
rect 13825 325 13905 365
rect 13945 325 14025 365
rect 13825 240 14025 325
rect 14175 365 14375 440
rect 14175 325 14255 365
rect 14295 325 14375 365
rect 14175 240 14375 325
rect 14525 365 14725 440
rect 14525 325 14605 365
rect 14645 325 14725 365
rect 14525 240 14725 325
rect 14875 365 15075 440
rect 14875 325 14955 365
rect 14995 325 15075 365
rect 14875 240 15075 325
rect 15225 365 15425 440
rect 15225 325 15305 365
rect 15345 325 15425 365
rect 15225 240 15425 325
rect 15575 365 15775 440
rect 15575 325 15655 365
rect 15695 325 15775 365
rect 15575 240 15775 325
rect 15925 365 16125 440
rect 15925 325 16005 365
rect 16045 325 16125 365
rect 15925 240 16125 325
rect 16275 365 16475 440
rect 16275 325 16355 365
rect 16395 325 16475 365
rect 16275 240 16475 325
rect 16625 365 16825 440
rect 16625 325 16705 365
rect 16745 325 16825 365
rect 16625 240 16825 325
rect 16975 365 17175 440
rect 16975 325 17055 365
rect 17095 325 17175 365
rect 16975 240 17175 325
rect 17325 365 17525 440
rect 17325 325 17405 365
rect 17445 325 17525 365
rect 17325 240 17525 325
rect 17675 365 17875 440
rect 17675 325 17755 365
rect 17795 325 17875 365
rect 17675 240 17875 325
rect 18025 365 18225 440
rect 18025 325 18105 365
rect 18145 325 18225 365
rect 18025 240 18225 325
rect 18375 365 18575 440
rect 18375 325 18455 365
rect 18495 325 18575 365
rect 18375 240 18575 325
rect 18725 365 18925 440
rect 18725 325 18805 365
rect 18845 325 18925 365
rect 18725 240 18925 325
rect 19075 365 19275 440
rect 19075 325 19155 365
rect 19195 325 19275 365
rect 19075 240 19275 325
rect 19425 365 19625 440
rect 19425 325 19505 365
rect 19545 325 19625 365
rect 19425 240 19625 325
rect 19775 365 19975 440
rect 19775 325 19855 365
rect 19895 325 19975 365
rect 19775 240 19975 325
rect 20125 365 20325 440
rect 20125 325 20205 365
rect 20245 325 20325 365
rect 20125 240 20325 325
rect 20475 365 20675 440
rect 20475 325 20555 365
rect 20595 325 20675 365
rect 20475 240 20675 325
rect 20825 365 21025 440
rect 20825 325 20905 365
rect 20945 325 21025 365
rect 20825 240 21025 325
rect 12775 15 12975 90
rect 12775 -25 12855 15
rect 12895 -25 12975 15
rect 12775 -110 12975 -25
rect 13125 15 13325 90
rect 13125 -25 13205 15
rect 13245 -25 13325 15
rect 13125 -110 13325 -25
rect 13475 15 13675 90
rect 13475 -25 13555 15
rect 13595 -25 13675 15
rect 13475 -110 13675 -25
rect 13825 15 14025 90
rect 13825 -25 13905 15
rect 13945 -25 14025 15
rect 13825 -110 14025 -25
rect 14175 15 14375 90
rect 14175 -25 14255 15
rect 14295 -25 14375 15
rect 14175 -110 14375 -25
rect 14525 15 14725 90
rect 14525 -25 14605 15
rect 14645 -25 14725 15
rect 14525 -110 14725 -25
rect 14875 15 15075 90
rect 14875 -25 14955 15
rect 14995 -25 15075 15
rect 14875 -110 15075 -25
rect 15225 15 15425 90
rect 15225 -25 15305 15
rect 15345 -25 15425 15
rect 15225 -110 15425 -25
rect 15575 15 15775 90
rect 15575 -25 15655 15
rect 15695 -25 15775 15
rect 15575 -110 15775 -25
rect 15925 15 16125 90
rect 15925 -25 16005 15
rect 16045 -25 16125 15
rect 15925 -110 16125 -25
rect 16275 15 16475 90
rect 16275 -25 16355 15
rect 16395 -25 16475 15
rect 16275 -110 16475 -25
rect 16625 15 16825 90
rect 16625 -25 16705 15
rect 16745 -25 16825 15
rect 16625 -110 16825 -25
rect 16975 15 17175 90
rect 16975 -25 17055 15
rect 17095 -25 17175 15
rect 16975 -110 17175 -25
rect 17325 15 17525 90
rect 17325 -25 17405 15
rect 17445 -25 17525 15
rect 17325 -110 17525 -25
rect 17675 15 17875 90
rect 17675 -25 17755 15
rect 17795 -25 17875 15
rect 17675 -110 17875 -25
rect 18025 15 18225 90
rect 18025 -25 18105 15
rect 18145 -25 18225 15
rect 18025 -110 18225 -25
rect 18375 15 18575 90
rect 18375 -25 18455 15
rect 18495 -25 18575 15
rect 18375 -110 18575 -25
rect 18725 15 18925 90
rect 18725 -25 18805 15
rect 18845 -25 18925 15
rect 18725 -110 18925 -25
rect 19075 15 19275 90
rect 19075 -25 19155 15
rect 19195 -25 19275 15
rect 19075 -110 19275 -25
rect 19425 15 19625 90
rect 19425 -25 19505 15
rect 19545 -25 19625 15
rect 19425 -110 19625 -25
rect 19775 15 19975 90
rect 19775 -25 19855 15
rect 19895 -25 19975 15
rect 19775 -110 19975 -25
rect 20125 15 20325 90
rect 20125 -25 20205 15
rect 20245 -25 20325 15
rect 20125 -110 20325 -25
rect 20475 15 20675 90
rect 20475 -25 20555 15
rect 20595 -25 20675 15
rect 20475 -110 20675 -25
rect 20825 15 21025 90
rect 20825 -25 20905 15
rect 20945 -25 21025 15
rect 20825 -110 21025 -25
rect 12775 -335 12975 -260
rect 12775 -375 12855 -335
rect 12895 -375 12975 -335
rect 12775 -460 12975 -375
rect 13125 -335 13325 -260
rect 13125 -375 13205 -335
rect 13245 -375 13325 -335
rect 13125 -460 13325 -375
rect 13475 -335 13675 -260
rect 13475 -375 13555 -335
rect 13595 -375 13675 -335
rect 13475 -460 13675 -375
rect 13825 -335 14025 -260
rect 13825 -375 13905 -335
rect 13945 -375 14025 -335
rect 13825 -460 14025 -375
rect 14175 -335 14375 -260
rect 14175 -375 14255 -335
rect 14295 -375 14375 -335
rect 14175 -460 14375 -375
rect 14525 -335 14725 -260
rect 14525 -375 14605 -335
rect 14645 -375 14725 -335
rect 14525 -460 14725 -375
rect 14875 -335 15075 -260
rect 14875 -375 14955 -335
rect 14995 -375 15075 -335
rect 14875 -460 15075 -375
rect 15225 -335 15425 -260
rect 15225 -375 15305 -335
rect 15345 -375 15425 -335
rect 15225 -460 15425 -375
rect 15575 -335 15775 -260
rect 15575 -375 15655 -335
rect 15695 -375 15775 -335
rect 15575 -460 15775 -375
rect 15925 -335 16125 -260
rect 15925 -375 16005 -335
rect 16045 -375 16125 -335
rect 15925 -460 16125 -375
rect 16275 -335 16475 -260
rect 16275 -375 16355 -335
rect 16395 -375 16475 -335
rect 16275 -460 16475 -375
rect 16625 -335 16825 -260
rect 16625 -375 16705 -335
rect 16745 -375 16825 -335
rect 16625 -460 16825 -375
rect 16975 -335 17175 -260
rect 16975 -375 17055 -335
rect 17095 -375 17175 -335
rect 16975 -460 17175 -375
rect 17325 -335 17525 -260
rect 17325 -375 17405 -335
rect 17445 -375 17525 -335
rect 17325 -460 17525 -375
rect 17675 -335 17875 -260
rect 17675 -375 17755 -335
rect 17795 -375 17875 -335
rect 17675 -460 17875 -375
rect 18025 -335 18225 -260
rect 18025 -375 18105 -335
rect 18145 -375 18225 -335
rect 18025 -460 18225 -375
rect 18375 -335 18575 -260
rect 18375 -375 18455 -335
rect 18495 -375 18575 -335
rect 18375 -460 18575 -375
rect 18725 -335 18925 -260
rect 18725 -375 18805 -335
rect 18845 -375 18925 -335
rect 18725 -460 18925 -375
rect 19075 -335 19275 -260
rect 19075 -375 19155 -335
rect 19195 -375 19275 -335
rect 19075 -460 19275 -375
rect 19425 -335 19625 -260
rect 19425 -375 19505 -335
rect 19545 -375 19625 -335
rect 19425 -460 19625 -375
rect 19775 -335 19975 -260
rect 19775 -375 19855 -335
rect 19895 -375 19975 -335
rect 19775 -460 19975 -375
rect 20125 -335 20325 -260
rect 20125 -375 20205 -335
rect 20245 -375 20325 -335
rect 20125 -460 20325 -375
rect 20475 -335 20675 -260
rect 20475 -375 20555 -335
rect 20595 -375 20675 -335
rect 20475 -460 20675 -375
rect 20825 -335 21025 -260
rect 20825 -375 20905 -335
rect 20945 -375 21025 -335
rect 20825 -460 21025 -375
<< mimcapcontact >>
rect 12855 5575 12895 5615
rect 13205 5575 13245 5615
rect 13555 5575 13595 5615
rect 13905 5575 13945 5615
rect 14255 5575 14295 5615
rect 14605 5575 14645 5615
rect 14955 5575 14995 5615
rect 15305 5575 15345 5615
rect 15655 5575 15695 5615
rect 16005 5575 16045 5615
rect 16355 5575 16395 5615
rect 16705 5575 16745 5615
rect 17055 5575 17095 5615
rect 17405 5575 17445 5615
rect 17755 5575 17795 5615
rect 18105 5575 18145 5615
rect 18455 5575 18495 5615
rect 18805 5575 18845 5615
rect 19155 5575 19195 5615
rect 19505 5575 19545 5615
rect 19855 5575 19895 5615
rect 20205 5575 20245 5615
rect 20555 5575 20595 5615
rect 20905 5575 20945 5615
rect 12855 5225 12895 5265
rect 13205 5225 13245 5265
rect 13555 5225 13595 5265
rect 13905 5225 13945 5265
rect 14255 5225 14295 5265
rect 14605 5225 14645 5265
rect 14955 5225 14995 5265
rect 15305 5225 15345 5265
rect 15655 5225 15695 5265
rect 16005 5225 16045 5265
rect 16355 5225 16395 5265
rect 16705 5225 16745 5265
rect 17055 5225 17095 5265
rect 17405 5225 17445 5265
rect 17755 5225 17795 5265
rect 18105 5225 18145 5265
rect 18455 5225 18495 5265
rect 18805 5225 18845 5265
rect 19155 5225 19195 5265
rect 19505 5225 19545 5265
rect 19855 5225 19895 5265
rect 20205 5225 20245 5265
rect 20555 5225 20595 5265
rect 20905 5225 20945 5265
rect 12855 4875 12895 4915
rect 240 4725 280 4765
rect 590 4725 630 4765
rect 940 4725 980 4765
rect 1290 4725 1330 4765
rect 1640 4725 1680 4765
rect 1990 4725 2030 4765
rect 2340 4725 2380 4765
rect 2690 4725 2730 4765
rect 3040 4725 3080 4765
rect 3390 4725 3430 4765
rect 3740 4725 3780 4765
rect 4090 4725 4130 4765
rect 4440 4725 4480 4765
rect 4790 4725 4830 4765
rect 13205 4875 13245 4915
rect 13555 4875 13595 4915
rect 13905 4875 13945 4915
rect 14255 4875 14295 4915
rect 14605 4875 14645 4915
rect 14955 4875 14995 4915
rect 15305 4875 15345 4915
rect 15655 4875 15695 4915
rect 16005 4875 16045 4915
rect 16355 4875 16395 4915
rect 16705 4875 16745 4915
rect 17055 4875 17095 4915
rect 17405 4875 17445 4915
rect 17755 4875 17795 4915
rect 18105 4875 18145 4915
rect 18455 4875 18495 4915
rect 18805 4875 18845 4915
rect 19155 4875 19195 4915
rect 19505 4875 19545 4915
rect 19855 4875 19895 4915
rect 20205 4875 20245 4915
rect 20555 4875 20595 4915
rect 20905 4875 20945 4915
rect 5140 4725 5180 4765
rect 12855 4525 12895 4565
rect 240 4375 280 4415
rect 590 4375 630 4415
rect 940 4375 980 4415
rect 1290 4375 1330 4415
rect 1640 4375 1680 4415
rect 1990 4375 2030 4415
rect 2340 4375 2380 4415
rect 2690 4375 2730 4415
rect 3040 4375 3080 4415
rect 3390 4375 3430 4415
rect 3740 4375 3780 4415
rect 4090 4375 4130 4415
rect 4440 4375 4480 4415
rect 4790 4375 4830 4415
rect 13205 4525 13245 4565
rect 13555 4525 13595 4565
rect 13905 4525 13945 4565
rect 14255 4525 14295 4565
rect 14605 4525 14645 4565
rect 14955 4525 14995 4565
rect 15305 4525 15345 4565
rect 15655 4525 15695 4565
rect 18105 4525 18145 4565
rect 18455 4525 18495 4565
rect 18805 4525 18845 4565
rect 19155 4525 19195 4565
rect 19505 4525 19545 4565
rect 19855 4525 19895 4565
rect 20205 4525 20245 4565
rect 20555 4525 20595 4565
rect 20905 4525 20945 4565
rect 5140 4375 5180 4415
rect 12855 4175 12895 4215
rect 240 4025 280 4065
rect 590 4025 630 4065
rect 940 4025 980 4065
rect 1290 4025 1330 4065
rect 1640 4025 1680 4065
rect 1990 4025 2030 4065
rect 2340 4025 2380 4065
rect 2690 4025 2730 4065
rect 3040 4025 3080 4065
rect 3390 4025 3430 4065
rect 3740 4025 3780 4065
rect 4090 4025 4130 4065
rect 4440 4025 4480 4065
rect 4790 4025 4830 4065
rect 13205 4175 13245 4215
rect 13555 4175 13595 4215
rect 13905 4175 13945 4215
rect 14255 4175 14295 4215
rect 14605 4175 14645 4215
rect 14955 4175 14995 4215
rect 15305 4175 15345 4215
rect 15655 4175 15695 4215
rect 18105 4175 18145 4215
rect 18455 4175 18495 4215
rect 18805 4175 18845 4215
rect 19155 4175 19195 4215
rect 19505 4175 19545 4215
rect 19855 4175 19895 4215
rect 20205 4175 20245 4215
rect 20555 4175 20595 4215
rect 20905 4175 20945 4215
rect 5140 4025 5180 4065
rect 12855 3825 12895 3865
rect 240 3675 280 3715
rect 590 3675 630 3715
rect 940 3675 980 3715
rect 1290 3675 1330 3715
rect 1640 3675 1680 3715
rect 1990 3675 2030 3715
rect 2340 3675 2380 3715
rect 2690 3675 2730 3715
rect 3040 3675 3080 3715
rect 3390 3675 3430 3715
rect 3740 3675 3780 3715
rect 4090 3675 4130 3715
rect 4440 3675 4480 3715
rect 4790 3675 4830 3715
rect 13205 3825 13245 3865
rect 13555 3825 13595 3865
rect 13905 3825 13945 3865
rect 14255 3825 14295 3865
rect 14605 3825 14645 3865
rect 14955 3825 14995 3865
rect 15305 3825 15345 3865
rect 15655 3825 15695 3865
rect 18105 3825 18145 3865
rect 18455 3825 18495 3865
rect 18805 3825 18845 3865
rect 19155 3825 19195 3865
rect 19505 3825 19545 3865
rect 19855 3825 19895 3865
rect 20205 3825 20245 3865
rect 20555 3825 20595 3865
rect 20905 3825 20945 3865
rect 5140 3675 5180 3715
rect 12855 3475 12895 3515
rect 13205 3475 13245 3515
rect 13555 3475 13595 3515
rect 13905 3475 13945 3515
rect 14255 3475 14295 3515
rect 19505 3475 19545 3515
rect 19855 3475 19895 3515
rect 20205 3475 20245 3515
rect 20555 3475 20595 3515
rect 20905 3475 20945 3515
rect 12855 3125 12895 3165
rect 13205 3125 13245 3165
rect 13555 3125 13595 3165
rect 13905 3125 13945 3165
rect 14255 3125 14295 3165
rect 19505 3125 19545 3165
rect 19855 3125 19895 3165
rect 20205 3125 20245 3165
rect 20555 3125 20595 3165
rect 20905 3125 20945 3165
rect 12855 2775 12895 2815
rect 13205 2775 13245 2815
rect 13555 2775 13595 2815
rect 13905 2775 13945 2815
rect 14255 2775 14295 2815
rect 19505 2775 19545 2815
rect 19855 2775 19895 2815
rect 20205 2775 20245 2815
rect 20555 2775 20595 2815
rect 20905 2775 20945 2815
rect 12855 2425 12895 2465
rect 13205 2425 13245 2465
rect 13555 2425 13595 2465
rect 13905 2425 13945 2465
rect 14255 2425 14295 2465
rect 19505 2425 19545 2465
rect 19855 2425 19895 2465
rect 20205 2425 20245 2465
rect 20555 2425 20595 2465
rect 20905 2425 20945 2465
rect 12855 2075 12895 2115
rect 13205 2075 13245 2115
rect 13555 2075 13595 2115
rect 13905 2075 13945 2115
rect 14255 2075 14295 2115
rect 19505 2075 19545 2115
rect 19855 2075 19895 2115
rect 20205 2075 20245 2115
rect 20555 2075 20595 2115
rect 20905 2075 20945 2115
rect 12855 1725 12895 1765
rect 13205 1725 13245 1765
rect 13555 1725 13595 1765
rect 13905 1725 13945 1765
rect 14255 1725 14295 1765
rect 19505 1725 19545 1765
rect 19855 1725 19895 1765
rect 20205 1725 20245 1765
rect 20555 1725 20595 1765
rect 20905 1725 20945 1765
rect 12855 1375 12895 1415
rect 13205 1375 13245 1415
rect 13555 1375 13595 1415
rect 13905 1375 13945 1415
rect 14255 1375 14295 1415
rect 19505 1375 19545 1415
rect 19855 1375 19895 1415
rect 20205 1375 20245 1415
rect 20555 1375 20595 1415
rect 20905 1375 20945 1415
rect 12855 1025 12895 1065
rect 13205 1025 13245 1065
rect 13555 1025 13595 1065
rect 13905 1025 13945 1065
rect 14255 1025 14295 1065
rect 19505 1025 19545 1065
rect 19855 1025 19895 1065
rect 20205 1025 20245 1065
rect 20555 1025 20595 1065
rect 20905 1025 20945 1065
rect 12855 675 12895 715
rect 13205 675 13245 715
rect 13555 675 13595 715
rect 13905 675 13945 715
rect 14255 675 14295 715
rect 19505 675 19545 715
rect 19855 675 19895 715
rect 20205 675 20245 715
rect 20555 675 20595 715
rect 20905 675 20945 715
rect 12855 325 12895 365
rect 13205 325 13245 365
rect 13555 325 13595 365
rect 13905 325 13945 365
rect 14255 325 14295 365
rect 14605 325 14645 365
rect 14955 325 14995 365
rect 15305 325 15345 365
rect 15655 325 15695 365
rect 16005 325 16045 365
rect 16355 325 16395 365
rect 16705 325 16745 365
rect 17055 325 17095 365
rect 17405 325 17445 365
rect 17755 325 17795 365
rect 18105 325 18145 365
rect 18455 325 18495 365
rect 18805 325 18845 365
rect 19155 325 19195 365
rect 19505 325 19545 365
rect 19855 325 19895 365
rect 20205 325 20245 365
rect 20555 325 20595 365
rect 20905 325 20945 365
rect 12855 -25 12895 15
rect 13205 -25 13245 15
rect 13555 -25 13595 15
rect 13905 -25 13945 15
rect 14255 -25 14295 15
rect 14605 -25 14645 15
rect 14955 -25 14995 15
rect 15305 -25 15345 15
rect 15655 -25 15695 15
rect 16005 -25 16045 15
rect 16355 -25 16395 15
rect 16705 -25 16745 15
rect 17055 -25 17095 15
rect 17405 -25 17445 15
rect 17755 -25 17795 15
rect 18105 -25 18145 15
rect 18455 -25 18495 15
rect 18805 -25 18845 15
rect 19155 -25 19195 15
rect 19505 -25 19545 15
rect 19855 -25 19895 15
rect 20205 -25 20245 15
rect 20555 -25 20595 15
rect 20905 -25 20945 15
rect 12855 -375 12895 -335
rect 13205 -375 13245 -335
rect 13555 -375 13595 -335
rect 13905 -375 13945 -335
rect 14255 -375 14295 -335
rect 14605 -375 14645 -335
rect 14955 -375 14995 -335
rect 15305 -375 15345 -335
rect 15655 -375 15695 -335
rect 16005 -375 16045 -335
rect 16355 -375 16395 -335
rect 16705 -375 16745 -335
rect 17055 -375 17095 -335
rect 17405 -375 17445 -335
rect 17755 -375 17795 -335
rect 18105 -375 18145 -335
rect 18455 -375 18495 -335
rect 18805 -375 18845 -335
rect 19155 -375 19195 -335
rect 19505 -375 19545 -335
rect 19855 -375 19895 -335
rect 20205 -375 20245 -335
rect 20555 -375 20595 -335
rect 20905 -375 20945 -335
<< metal4 >>
rect 12850 5615 13600 5620
rect 12850 5575 12855 5615
rect 12895 5575 13205 5615
rect 13245 5575 13555 5615
rect 13595 5575 13600 5615
rect 12850 5570 13600 5575
rect 13550 5270 13600 5570
rect 13900 5615 13950 5620
rect 13900 5575 13905 5615
rect 13945 5575 13950 5615
rect 13900 5270 13950 5575
rect 14250 5615 14300 5620
rect 14250 5575 14255 5615
rect 14295 5575 14300 5615
rect 14250 5270 14300 5575
rect 14600 5615 14650 5620
rect 14600 5575 14605 5615
rect 14645 5575 14650 5615
rect 14600 5270 14650 5575
rect 14950 5615 15000 5620
rect 14950 5575 14955 5615
rect 14995 5575 15000 5615
rect 14950 5270 15000 5575
rect 15300 5615 15350 5620
rect 15300 5575 15305 5615
rect 15345 5575 15350 5615
rect 15300 5270 15350 5575
rect 15650 5615 15700 5620
rect 15650 5575 15655 5615
rect 15695 5575 15700 5615
rect 15650 5270 15700 5575
rect 16000 5615 16050 5620
rect 16000 5575 16005 5615
rect 16045 5575 16050 5615
rect 16000 5270 16050 5575
rect 16350 5615 16400 5620
rect 16350 5575 16355 5615
rect 16395 5575 16400 5615
rect 16350 5270 16400 5575
rect 16700 5615 16750 5620
rect 16700 5575 16705 5615
rect 16745 5575 16750 5615
rect 16700 5270 16750 5575
rect 12850 5265 16750 5270
rect 12850 5225 12855 5265
rect 12895 5225 13205 5265
rect 13245 5225 13555 5265
rect 13595 5225 13905 5265
rect 13945 5225 14255 5265
rect 14295 5225 14605 5265
rect 14645 5225 14955 5265
rect 14995 5225 15305 5265
rect 15345 5225 15655 5265
rect 15695 5225 16005 5265
rect 16045 5225 16355 5265
rect 16395 5225 16705 5265
rect 16745 5225 16750 5265
rect 12850 5220 16750 5225
rect -200 4995 5595 5000
rect -200 4955 -195 4995
rect -155 4955 5550 4995
rect 5590 4955 5595 4995
rect -200 4950 5595 4955
rect 13550 4920 13600 5220
rect 12850 4915 14300 4920
rect -115 4910 5510 4915
rect -115 4870 -110 4910
rect -70 4870 5465 4910
rect 5505 4870 5510 4910
rect 12850 4875 12855 4915
rect 12895 4875 13205 4915
rect 13245 4875 13555 4915
rect 13595 4875 13905 4915
rect 13945 4875 14255 4915
rect 14295 4875 14300 4915
rect 12850 4870 14300 4875
rect 14600 4915 14650 5220
rect 14600 4875 14605 4915
rect 14645 4875 14650 4915
rect -115 4865 5510 4870
rect 235 4765 1685 4770
rect 235 4725 240 4765
rect 280 4725 590 4765
rect 630 4725 940 4765
rect 980 4725 1290 4765
rect 1330 4725 1640 4765
rect 1680 4725 1685 4765
rect 235 4720 1685 4725
rect 1985 4765 3435 4770
rect 1985 4725 1990 4765
rect 2030 4725 2340 4765
rect 2380 4725 2690 4765
rect 2730 4725 3040 4765
rect 3080 4725 3390 4765
rect 3430 4725 3435 4765
rect 1985 4720 3435 4725
rect 3735 4765 5185 4770
rect 3735 4725 3740 4765
rect 3780 4725 4090 4765
rect 4130 4725 4440 4765
rect 4480 4725 4790 4765
rect 4830 4725 5140 4765
rect 5180 4725 5185 4765
rect 3735 4720 5185 4725
rect 935 4420 985 4720
rect 2685 4420 2735 4720
rect 4435 4420 4485 4720
rect 13550 4570 13600 4870
rect 12850 4565 14300 4570
rect 12850 4525 12855 4565
rect 12895 4525 13205 4565
rect 13245 4525 13555 4565
rect 13595 4525 13905 4565
rect 13945 4525 14255 4565
rect 14295 4525 14300 4565
rect 12850 4520 14300 4525
rect 14600 4565 14650 4875
rect 14600 4525 14605 4565
rect 14645 4525 14650 4565
rect 235 4415 1685 4420
rect 235 4375 240 4415
rect 280 4375 590 4415
rect 630 4375 940 4415
rect 980 4375 1290 4415
rect 1330 4375 1640 4415
rect 1680 4375 1685 4415
rect 235 4370 1685 4375
rect 1985 4415 3435 4420
rect 1985 4375 1990 4415
rect 2030 4375 2340 4415
rect 2380 4375 2690 4415
rect 2730 4375 3040 4415
rect 3080 4375 3390 4415
rect 3430 4375 3435 4415
rect 1985 4370 3435 4375
rect 3735 4415 5185 4420
rect 3735 4375 3740 4415
rect 3780 4375 4090 4415
rect 4130 4375 4440 4415
rect 4480 4375 4790 4415
rect 4830 4375 5140 4415
rect 5180 4375 5185 4415
rect 3735 4370 5185 4375
rect 935 4070 985 4370
rect 2685 4070 2735 4370
rect 4435 4070 4485 4370
rect 13550 4220 13600 4520
rect 12850 4215 14300 4220
rect 12850 4175 12855 4215
rect 12895 4175 13205 4215
rect 13245 4175 13555 4215
rect 13595 4175 13905 4215
rect 13945 4175 14255 4215
rect 14295 4175 14300 4215
rect 12850 4170 14300 4175
rect 14600 4215 14650 4525
rect 14600 4175 14605 4215
rect 14645 4175 14650 4215
rect 235 4065 1685 4070
rect 235 4025 240 4065
rect 280 4025 590 4065
rect 630 4025 940 4065
rect 980 4025 1290 4065
rect 1330 4025 1640 4065
rect 1680 4025 1685 4065
rect 235 4020 1685 4025
rect 1985 4065 3435 4070
rect 1985 4025 1990 4065
rect 2030 4025 2340 4065
rect 2380 4025 2690 4065
rect 2730 4025 3040 4065
rect 3080 4025 3390 4065
rect 3430 4025 3435 4065
rect 1985 4020 3435 4025
rect 3735 4065 5185 4070
rect 3735 4025 3740 4065
rect 3780 4025 4090 4065
rect 4130 4025 4440 4065
rect 4480 4025 4790 4065
rect 4830 4025 5140 4065
rect 5180 4025 5185 4065
rect 3735 4020 5185 4025
rect 935 3720 985 4020
rect 2685 3720 2735 4020
rect 4435 3720 4485 4020
rect 13550 3870 13600 4170
rect 12850 3865 14300 3870
rect 12850 3825 12855 3865
rect 12895 3825 13205 3865
rect 13245 3825 13555 3865
rect 13595 3825 13905 3865
rect 13945 3825 14255 3865
rect 14295 3825 14300 3865
rect 12850 3820 14300 3825
rect 14600 3865 14650 4175
rect 14600 3825 14605 3865
rect 14645 3825 14650 3865
rect 14600 3820 14650 3825
rect 14950 4915 15000 5220
rect 14950 4875 14955 4915
rect 14995 4875 15000 4915
rect 14950 4565 15000 4875
rect 14950 4525 14955 4565
rect 14995 4525 15000 4565
rect 14950 4215 15000 4525
rect 14950 4175 14955 4215
rect 14995 4175 15000 4215
rect 14950 3865 15000 4175
rect 14950 3825 14955 3865
rect 14995 3825 15000 3865
rect 14950 3820 15000 3825
rect 15300 4915 15350 5220
rect 15300 4875 15305 4915
rect 15345 4875 15350 4915
rect 15300 4565 15350 4875
rect 15300 4525 15305 4565
rect 15345 4525 15350 4565
rect 15300 4215 15350 4525
rect 15300 4175 15305 4215
rect 15345 4175 15350 4215
rect 15300 3865 15350 4175
rect 15300 3825 15305 3865
rect 15345 3825 15350 3865
rect 15300 3820 15350 3825
rect 15650 4915 15700 5220
rect 15650 4875 15655 4915
rect 15695 4875 15700 4915
rect 15650 4565 15700 4875
rect 16000 4915 16050 5220
rect 16000 4875 16005 4915
rect 16045 4875 16050 4915
rect 16000 4870 16050 4875
rect 16350 4915 16400 5220
rect 16350 4875 16355 4915
rect 16395 4875 16400 4915
rect 16350 4870 16400 4875
rect 16700 4915 16750 5220
rect 16700 4875 16705 4915
rect 16745 4875 16750 4915
rect 16700 4870 16750 4875
rect 17050 5615 17100 5620
rect 17050 5575 17055 5615
rect 17095 5575 17100 5615
rect 17050 5270 17100 5575
rect 17400 5615 17450 5620
rect 17400 5575 17405 5615
rect 17445 5575 17450 5615
rect 17400 5270 17450 5575
rect 17750 5615 17800 5620
rect 17750 5575 17755 5615
rect 17795 5575 17800 5615
rect 17750 5270 17800 5575
rect 18100 5615 18150 5620
rect 18100 5575 18105 5615
rect 18145 5575 18150 5615
rect 18100 5270 18150 5575
rect 18450 5615 18500 5620
rect 18450 5575 18455 5615
rect 18495 5575 18500 5615
rect 18450 5270 18500 5575
rect 18800 5615 18850 5620
rect 18800 5575 18805 5615
rect 18845 5575 18850 5615
rect 18800 5270 18850 5575
rect 19150 5615 19200 5620
rect 19150 5575 19155 5615
rect 19195 5575 19200 5615
rect 19150 5270 19200 5575
rect 19500 5615 19550 5620
rect 19500 5575 19505 5615
rect 19545 5575 19550 5615
rect 19500 5270 19550 5575
rect 19850 5615 19900 5620
rect 19850 5575 19855 5615
rect 19895 5575 19900 5615
rect 19850 5270 19900 5575
rect 20200 5615 20950 5620
rect 20200 5575 20205 5615
rect 20245 5575 20555 5615
rect 20595 5575 20905 5615
rect 20945 5575 20950 5615
rect 20200 5570 20950 5575
rect 20200 5270 20250 5570
rect 17050 5265 20950 5270
rect 17050 5225 17055 5265
rect 17095 5225 17405 5265
rect 17445 5225 17755 5265
rect 17795 5225 18105 5265
rect 18145 5225 18455 5265
rect 18495 5225 18805 5265
rect 18845 5225 19155 5265
rect 19195 5225 19505 5265
rect 19545 5225 19855 5265
rect 19895 5225 20205 5265
rect 20245 5225 20555 5265
rect 20595 5225 20905 5265
rect 20945 5225 20950 5265
rect 17050 5220 20950 5225
rect 17050 4915 17100 5220
rect 17050 4875 17055 4915
rect 17095 4875 17100 4915
rect 17050 4870 17100 4875
rect 17400 4915 17450 5220
rect 17400 4875 17405 4915
rect 17445 4875 17450 4915
rect 17400 4870 17450 4875
rect 17750 4915 17800 5220
rect 17750 4875 17755 4915
rect 17795 4875 17800 4915
rect 17750 4870 17800 4875
rect 18100 4915 18150 5220
rect 18100 4875 18105 4915
rect 18145 4875 18150 4915
rect 15650 4525 15655 4565
rect 15695 4525 15700 4565
rect 15650 4215 15700 4525
rect 15650 4175 15655 4215
rect 15695 4175 15700 4215
rect 15650 3865 15700 4175
rect 15650 3825 15655 3865
rect 15695 3825 15700 3865
rect 15650 3820 15700 3825
rect 18100 4565 18150 4875
rect 18100 4525 18105 4565
rect 18145 4525 18150 4565
rect 18100 4215 18150 4525
rect 18100 4175 18105 4215
rect 18145 4175 18150 4215
rect 18100 3865 18150 4175
rect 18100 3825 18105 3865
rect 18145 3825 18150 3865
rect 18100 3820 18150 3825
rect 18450 4915 18500 5220
rect 18450 4875 18455 4915
rect 18495 4875 18500 4915
rect 18450 4565 18500 4875
rect 18450 4525 18455 4565
rect 18495 4525 18500 4565
rect 18450 4215 18500 4525
rect 18450 4175 18455 4215
rect 18495 4175 18500 4215
rect 18450 3865 18500 4175
rect 18450 3825 18455 3865
rect 18495 3825 18500 3865
rect 18450 3820 18500 3825
rect 18800 4915 18850 5220
rect 18800 4875 18805 4915
rect 18845 4875 18850 4915
rect 18800 4565 18850 4875
rect 18800 4525 18805 4565
rect 18845 4525 18850 4565
rect 18800 4215 18850 4525
rect 18800 4175 18805 4215
rect 18845 4175 18850 4215
rect 18800 3865 18850 4175
rect 18800 3825 18805 3865
rect 18845 3825 18850 3865
rect 18800 3820 18850 3825
rect 19150 4915 19200 5220
rect 20200 4920 20250 5220
rect 19150 4875 19155 4915
rect 19195 4875 19200 4915
rect 19150 4565 19200 4875
rect 19500 4915 20950 4920
rect 19500 4875 19505 4915
rect 19545 4875 19855 4915
rect 19895 4875 20205 4915
rect 20245 4875 20555 4915
rect 20595 4875 20905 4915
rect 20945 4875 20950 4915
rect 19500 4870 20950 4875
rect 20200 4570 20250 4870
rect 19150 4525 19155 4565
rect 19195 4525 19200 4565
rect 19150 4215 19200 4525
rect 19500 4565 20950 4570
rect 19500 4525 19505 4565
rect 19545 4525 19855 4565
rect 19895 4525 20205 4565
rect 20245 4525 20555 4565
rect 20595 4525 20905 4565
rect 20945 4525 20950 4565
rect 19500 4520 20950 4525
rect 20200 4220 20250 4520
rect 19150 4175 19155 4215
rect 19195 4175 19200 4215
rect 19150 3865 19200 4175
rect 19500 4215 20950 4220
rect 19500 4175 19505 4215
rect 19545 4175 19855 4215
rect 19895 4175 20205 4215
rect 20245 4175 20555 4215
rect 20595 4175 20905 4215
rect 20945 4175 20950 4215
rect 19500 4170 20950 4175
rect 20200 3870 20250 4170
rect 19150 3825 19155 3865
rect 19195 3825 19200 3865
rect 19150 3820 19200 3825
rect 19500 3865 20950 3870
rect 19500 3825 19505 3865
rect 19545 3825 19855 3865
rect 19895 3825 20205 3865
rect 20245 3825 20555 3865
rect 20595 3825 20905 3865
rect 20945 3825 20950 3865
rect 19500 3820 20950 3825
rect 235 3715 1685 3720
rect 235 3675 240 3715
rect 280 3675 590 3715
rect 630 3675 940 3715
rect 980 3675 1290 3715
rect 1330 3675 1640 3715
rect 1680 3675 1685 3715
rect 235 3670 1685 3675
rect 1985 3715 3435 3720
rect 1985 3675 1990 3715
rect 2030 3675 2340 3715
rect 2380 3675 2690 3715
rect 2730 3675 3040 3715
rect 3080 3675 3390 3715
rect 3430 3675 3435 3715
rect 1985 3670 3435 3675
rect 3735 3715 5185 3720
rect 3735 3675 3740 3715
rect 3780 3675 4090 3715
rect 4130 3675 4440 3715
rect 4480 3675 4790 3715
rect 4830 3675 5140 3715
rect 5180 3675 5185 3715
rect 3735 3670 5185 3675
rect 1635 3450 1685 3670
rect 1635 3410 1640 3450
rect 1680 3410 1685 3450
rect 1635 3405 1685 3410
rect 3385 3340 3435 3670
rect 5135 3450 5185 3670
rect 13550 3520 13600 3820
rect 20200 3520 20250 3820
rect 12850 3515 14300 3520
rect 12850 3475 12855 3515
rect 12895 3475 13205 3515
rect 13245 3475 13555 3515
rect 13595 3475 13905 3515
rect 13945 3475 14255 3515
rect 14295 3475 14300 3515
rect 12850 3470 14300 3475
rect 19500 3515 20950 3520
rect 19500 3475 19505 3515
rect 19545 3475 19855 3515
rect 19895 3475 20205 3515
rect 20245 3475 20555 3515
rect 20595 3475 20905 3515
rect 20945 3475 20950 3515
rect 19500 3470 20950 3475
rect 5135 3410 5140 3450
rect 5180 3410 5185 3450
rect 5135 3405 5185 3410
rect 3385 3300 3390 3340
rect 3430 3300 3435 3340
rect 3385 3295 3435 3300
rect 13550 3170 13600 3470
rect 20200 3170 20250 3470
rect 12850 3165 14300 3170
rect 12850 3125 12855 3165
rect 12895 3125 13205 3165
rect 13245 3125 13555 3165
rect 13595 3125 13905 3165
rect 13945 3125 14255 3165
rect 14295 3125 14300 3165
rect 12850 3120 14300 3125
rect 19500 3165 20950 3170
rect 19500 3125 19505 3165
rect 19545 3125 19855 3165
rect 19895 3125 20205 3165
rect 20245 3125 20555 3165
rect 20595 3125 20905 3165
rect 20945 3125 20950 3165
rect 19500 3120 20950 3125
rect 13550 2820 13600 3120
rect 20200 2820 20250 3120
rect 12850 2815 14300 2820
rect 12850 2775 12855 2815
rect 12895 2775 13205 2815
rect 13245 2775 13555 2815
rect 13595 2775 13905 2815
rect 13945 2775 14255 2815
rect 14295 2775 14300 2815
rect 12850 2770 14300 2775
rect 19500 2815 20950 2820
rect 19500 2775 19505 2815
rect 19545 2775 19855 2815
rect 19895 2775 20205 2815
rect 20245 2775 20555 2815
rect 20595 2775 20905 2815
rect 20945 2775 20950 2815
rect 19500 2770 20950 2775
rect 13550 2470 13600 2770
rect 20200 2470 20250 2770
rect 12850 2465 14300 2470
rect 12850 2425 12855 2465
rect 12895 2425 13205 2465
rect 13245 2425 13555 2465
rect 13595 2425 13905 2465
rect 13945 2425 14255 2465
rect 14295 2425 14300 2465
rect 12850 2420 14300 2425
rect 19500 2465 20950 2470
rect 19500 2425 19505 2465
rect 19545 2425 19855 2465
rect 19895 2425 20205 2465
rect 20245 2425 20555 2465
rect 20595 2425 20905 2465
rect 20945 2425 20950 2465
rect 19500 2420 20950 2425
rect 13550 2120 13600 2420
rect 20200 2120 20250 2420
rect 12850 2115 14560 2120
rect 12850 2075 12855 2115
rect 12895 2075 13205 2115
rect 13245 2075 13555 2115
rect 13595 2075 13905 2115
rect 13945 2075 14255 2115
rect 14295 2075 14515 2115
rect 14555 2075 14560 2115
rect 12850 2070 14560 2075
rect 19240 2115 20950 2120
rect 19240 2075 19245 2115
rect 19285 2075 19505 2115
rect 19545 2075 19855 2115
rect 19895 2075 20205 2115
rect 20245 2075 20555 2115
rect 20595 2075 20905 2115
rect 20945 2075 20950 2115
rect 19240 2070 20950 2075
rect 13550 1770 13600 2070
rect 20200 1770 20250 2070
rect 12850 1765 14300 1770
rect 12850 1725 12855 1765
rect 12895 1725 13205 1765
rect 13245 1725 13555 1765
rect 13595 1725 13905 1765
rect 13945 1725 14255 1765
rect 14295 1725 14300 1765
rect 12850 1720 14300 1725
rect 19500 1765 20950 1770
rect 19500 1725 19505 1765
rect 19545 1725 19855 1765
rect 19895 1725 20205 1765
rect 20245 1725 20555 1765
rect 20595 1725 20905 1765
rect 20945 1725 20950 1765
rect 19500 1720 20950 1725
rect 13550 1420 13600 1720
rect 20200 1420 20250 1720
rect 12850 1415 14300 1420
rect 12850 1375 12855 1415
rect 12895 1375 13205 1415
rect 13245 1375 13555 1415
rect 13595 1375 13905 1415
rect 13945 1375 14255 1415
rect 14295 1375 14300 1415
rect 12850 1370 14300 1375
rect 19500 1415 20950 1420
rect 19500 1375 19505 1415
rect 19545 1375 19855 1415
rect 19895 1375 20205 1415
rect 20245 1375 20555 1415
rect 20595 1375 20905 1415
rect 20945 1375 20950 1415
rect 19500 1370 20950 1375
rect 13550 1070 13600 1370
rect 20200 1070 20250 1370
rect 12850 1065 14300 1070
rect 12850 1025 12855 1065
rect 12895 1025 13205 1065
rect 13245 1025 13555 1065
rect 13595 1025 13905 1065
rect 13945 1025 14255 1065
rect 14295 1025 14300 1065
rect 12850 1020 14300 1025
rect 19500 1065 20950 1070
rect 19500 1025 19505 1065
rect 19545 1025 19855 1065
rect 19895 1025 20205 1065
rect 20245 1025 20555 1065
rect 20595 1025 20905 1065
rect 20945 1025 20950 1065
rect 19500 1020 20950 1025
rect 13550 720 13600 1020
rect 20200 720 20250 1020
rect 12850 715 14300 720
rect 12850 675 12855 715
rect 12895 675 13205 715
rect 13245 675 13555 715
rect 13595 675 13905 715
rect 13945 675 14255 715
rect 14295 675 14300 715
rect 12850 670 14300 675
rect 19500 715 20950 720
rect 19500 675 19505 715
rect 19545 675 19855 715
rect 19895 675 20205 715
rect 20245 675 20555 715
rect 20595 675 20905 715
rect 20945 675 20950 715
rect 19500 670 20950 675
rect -115 660 5510 665
rect -115 620 -110 660
rect -70 620 5465 660
rect 5505 620 5510 660
rect -115 615 5510 620
rect -200 580 5595 585
rect -200 540 -195 580
rect -155 540 5550 580
rect 5590 540 5595 580
rect -200 535 5595 540
rect 13550 370 13600 670
rect 20200 370 20250 670
rect 12850 365 13600 370
rect 12850 325 12855 365
rect 12895 325 13205 365
rect 13245 325 13555 365
rect 13595 325 13600 365
rect 12850 320 13600 325
rect 13550 20 13600 320
rect 13900 365 13950 370
rect 13900 325 13905 365
rect 13945 325 13950 365
rect 13900 20 13950 325
rect 14250 365 14300 370
rect 14250 325 14255 365
rect 14295 325 14300 365
rect 14250 20 14300 325
rect 14600 365 14650 370
rect 14600 325 14605 365
rect 14645 325 14650 365
rect 14600 20 14650 325
rect 14950 365 15000 370
rect 14950 325 14955 365
rect 14995 325 15000 365
rect 14950 20 15000 325
rect 15300 365 15350 370
rect 15300 325 15305 365
rect 15345 325 15350 365
rect 15300 20 15350 325
rect 15650 365 15700 370
rect 15650 325 15655 365
rect 15695 325 15700 365
rect 15650 20 15700 325
rect 16000 365 16050 370
rect 16000 325 16005 365
rect 16045 325 16050 365
rect 16000 20 16050 325
rect 16350 365 16400 370
rect 16350 325 16355 365
rect 16395 325 16400 365
rect 16350 20 16400 325
rect 16700 365 16750 370
rect 16700 325 16705 365
rect 16745 325 16750 365
rect 16700 20 16750 325
rect 12850 15 16750 20
rect 12850 -25 12855 15
rect 12895 -25 13205 15
rect 13245 -25 13555 15
rect 13595 -25 13905 15
rect 13945 -25 14255 15
rect 14295 -25 14605 15
rect 14645 -25 14955 15
rect 14995 -25 15305 15
rect 15345 -25 15655 15
rect 15695 -25 16005 15
rect 16045 -25 16355 15
rect 16395 -25 16705 15
rect 16745 -25 16750 15
rect 12850 -30 16750 -25
rect 13550 -330 13600 -30
rect 12850 -335 13600 -330
rect 12850 -375 12855 -335
rect 12895 -375 13205 -335
rect 13245 -375 13555 -335
rect 13595 -375 13600 -335
rect 12850 -380 13600 -375
rect 13900 -335 13950 -30
rect 13900 -375 13905 -335
rect 13945 -375 13950 -335
rect 13900 -380 13950 -375
rect 14250 -335 14300 -30
rect 14250 -375 14255 -335
rect 14295 -375 14300 -335
rect 14250 -380 14300 -375
rect 14600 -335 14650 -30
rect 14600 -375 14605 -335
rect 14645 -375 14650 -335
rect 14600 -380 14650 -375
rect 14950 -335 15000 -30
rect 14950 -375 14955 -335
rect 14995 -375 15000 -335
rect 14950 -380 15000 -375
rect 15300 -335 15350 -30
rect 15300 -375 15305 -335
rect 15345 -375 15350 -335
rect 15300 -380 15350 -375
rect 15650 -335 15700 -30
rect 15650 -375 15655 -335
rect 15695 -375 15700 -335
rect 15650 -380 15700 -375
rect 16000 -335 16050 -30
rect 16000 -375 16005 -335
rect 16045 -375 16050 -335
rect 16000 -380 16050 -375
rect 16350 -335 16400 -30
rect 16350 -375 16355 -335
rect 16395 -375 16400 -335
rect 16350 -380 16400 -375
rect 16700 -335 16750 -30
rect 16700 -375 16705 -335
rect 16745 -375 16750 -335
rect 16700 -380 16750 -375
rect 17050 365 17100 370
rect 17050 325 17055 365
rect 17095 325 17100 365
rect 17050 20 17100 325
rect 17400 365 17450 370
rect 17400 325 17405 365
rect 17445 325 17450 365
rect 17400 20 17450 325
rect 17750 365 17800 370
rect 17750 325 17755 365
rect 17795 325 17800 365
rect 17750 20 17800 325
rect 18100 365 18150 370
rect 18100 325 18105 365
rect 18145 325 18150 365
rect 18100 20 18150 325
rect 18450 365 18500 370
rect 18450 325 18455 365
rect 18495 325 18500 365
rect 18450 20 18500 325
rect 18800 365 18850 370
rect 18800 325 18805 365
rect 18845 325 18850 365
rect 18800 20 18850 325
rect 19150 365 19200 370
rect 19150 325 19155 365
rect 19195 325 19200 365
rect 19150 20 19200 325
rect 19500 365 19550 370
rect 19500 325 19505 365
rect 19545 325 19550 365
rect 19500 20 19550 325
rect 19850 365 19900 370
rect 19850 325 19855 365
rect 19895 325 19900 365
rect 19850 20 19900 325
rect 20200 365 20950 370
rect 20200 325 20205 365
rect 20245 325 20555 365
rect 20595 325 20905 365
rect 20945 325 20950 365
rect 20200 320 20950 325
rect 20200 20 20250 320
rect 17050 15 20950 20
rect 17050 -25 17055 15
rect 17095 -25 17405 15
rect 17445 -25 17755 15
rect 17795 -25 18105 15
rect 18145 -25 18455 15
rect 18495 -25 18805 15
rect 18845 -25 19155 15
rect 19195 -25 19505 15
rect 19545 -25 19855 15
rect 19895 -25 20205 15
rect 20245 -25 20555 15
rect 20595 -25 20905 15
rect 20945 -25 20950 15
rect 17050 -30 20950 -25
rect 17050 -335 17100 -30
rect 17050 -375 17055 -335
rect 17095 -375 17100 -335
rect 17050 -380 17100 -375
rect 17400 -335 17450 -30
rect 17400 -375 17405 -335
rect 17445 -375 17450 -335
rect 17400 -380 17450 -375
rect 17750 -335 17800 -30
rect 17750 -375 17755 -335
rect 17795 -375 17800 -335
rect 17750 -380 17800 -375
rect 18100 -335 18150 -30
rect 18100 -375 18105 -335
rect 18145 -375 18150 -335
rect 18100 -380 18150 -375
rect 18450 -335 18500 -30
rect 18450 -375 18455 -335
rect 18495 -375 18500 -335
rect 18450 -380 18500 -375
rect 18800 -335 18850 -30
rect 18800 -375 18805 -335
rect 18845 -375 18850 -335
rect 18800 -380 18850 -375
rect 19150 -335 19200 -30
rect 19150 -375 19155 -335
rect 19195 -375 19200 -335
rect 19150 -380 19200 -375
rect 19500 -335 19550 -30
rect 19500 -375 19505 -335
rect 19545 -375 19550 -335
rect 19500 -380 19550 -375
rect 19850 -335 19900 -30
rect 19850 -375 19855 -335
rect 19895 -375 19900 -335
rect 19850 -380 19900 -375
rect 20200 -330 20250 -30
rect 20200 -335 20950 -330
rect 20200 -375 20205 -335
rect 20245 -375 20555 -335
rect 20595 -375 20905 -335
rect 20945 -375 20950 -335
rect 20200 -380 20950 -375
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 795 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 795 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 795 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 115 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 115 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 115 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 1475 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_7
timestamp 1723858470
transform 1 0 1475 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8
timestamp 1723858470
transform 1 0 1475 0 1 1360
box 0 0 670 670
<< labels >>
flabel metal2 2950 1735 2950 1735 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 2955 1590 2955 1590 1 FreeSans 400 0 0 80 Vin+
flabel metal2 2945 1845 2945 1845 5 FreeSans 400 0 0 -40 V_mir1
flabel metal2 3745 1530 3745 1530 3 FreeSans 400 0 40 0 V_p1
flabel metal1 2650 1155 2650 1155 3 FreeSans 400 0 200 0 START_UP
flabel metal2 3785 1785 3785 1785 5 FreeSans 400 0 0 -40 1st_Vout1
flabel metal2 455 3440 455 3440 1 FreeSans 400 0 0 40 cap_res1
flabel metal3 2730 3375 2730 3375 3 FreeSans 400 0 40 0 cap_res2
flabel metal1 2550 845 2550 845 3 FreeSans 400 0 40 0 NFET_GATE_10uA
flabel metal2 5120 1590 5120 1590 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal2 4225 1785 4225 1785 5 FreeSans 400 0 0 -40 1st_Vout2
flabel metal2 5065 1845 5065 1845 5 FreeSans 400 0 0 -40 V_mir2
flabel metal2 4265 1530 4265 1530 7 FreeSans 400 0 -40 0 V_p2
flabel metal1 3275 350 3275 350 7 FreeSans 400 0 -400 0 CMFB_NFET_CUR_BIAS
port 8 w
flabel metal1 3825 295 3825 295 5 FreeSans 400 0 0 -200 VB2_CUR_BIAS
port 5 s
flabel metal1 4015 350 4015 350 3 FreeSans 400 0 200 0 ERR_AMP_CUR_BIAS
port 7 e
flabel metal1 4725 295 4725 295 5 FreeSans 400 0 0 -200 VB3_CUR_BIAS
port 6 s
flabel metal1 4985 1110 4985 1110 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal2 4115 3135 4115 3135 1 FreeSans 400 0 0 40 PFET_GATE_10uA
flabel metal2 6080 3075 6080 3075 1 FreeSans 400 0 0 200 VB1_CUR_BIAS
port 1 n
flabel metal2 6100 3020 6100 3020 3 FreeSans 400 0 200 0 TAIL_CUR_MIR_BIAS
port 9 e
flabel metal2 6080 2955 6080 2955 5 FreeSans 400 0 0 -200 CMFB_PFET_CUR_BIAS
port 10 s
flabel metal2 6100 1745 6100 1745 3 FreeSans 400 0 200 0 ERR_AMP_REF
port 3 e
flabel metal3 5590 4400 5590 4400 3 FreeSans 800 0 80 0 VDDA
port 4 e
flabel metal3 5505 4175 5505 4175 3 FreeSans 800 0 80 0 GNDA
port 2 e
flabel metal1 2180 1010 2180 1010 3 FreeSans 400 0 40 0 Vbe2
flabel poly 4635 2375 4635 2375 5 FreeSans 400 0 0 -40 V_TOP
<< end >>
