magic
tech sky130A
magscale 1 2
timestamp 1738562572
<< nwell >>
rect -30 520 3310 600
rect -460 350 3560 520
rect -460 -770 -290 350
rect -30 340 3560 350
rect -30 260 3310 340
rect -30 -720 3250 -716
rect -30 -740 3300 -720
rect -30 -770 3560 -740
rect -460 -920 3560 -770
rect -460 -950 3300 -920
rect -30 -1048 3300 -950
<< pwell >>
rect 10 40 3270 210
rect 770 0 990 40
rect 770 -50 870 0
rect 950 -50 990 0
rect 1790 20 1870 40
rect 1790 -190 1830 20
rect 770 -500 990 -410
rect 2730 -500 2990 -410
rect 10 -660 3260 -500
<< poly >>
rect 3300 620 3380 640
rect 3300 580 3320 620
rect 3360 580 3380 620
rect 3300 560 3380 580
rect 800 470 960 490
rect 800 460 900 470
rect 800 260 830 460
rect 880 430 900 460
rect 940 430 960 470
rect 880 410 960 430
rect 1790 290 1870 310
rect 1790 260 1810 290
rect 260 230 340 260
rect 750 230 830 260
rect 1730 250 1810 260
rect 1850 250 1870 290
rect 3300 260 3330 560
rect 1730 230 1870 250
rect 3240 230 3330 260
rect 3380 410 3460 430
rect 3380 370 3400 410
rect 3440 370 3460 410
rect 3380 350 3460 370
rect 310 -110 340 230
rect 1790 100 1820 230
rect 1790 80 1870 100
rect 1790 40 1810 80
rect 1850 40 1870 80
rect 1790 20 1870 40
rect 870 0 950 20
rect 870 -40 890 0
rect 930 -30 950 0
rect 2870 0 2950 20
rect 2870 -30 2890 0
rect 930 -40 2890 -30
rect 2930 -40 2950 0
rect 870 -60 2950 -40
rect 3380 -110 3410 350
rect 310 -130 3410 -110
rect 310 -140 1810 -130
rect 1790 -170 1810 -140
rect 1850 -140 3410 -130
rect 1850 -170 1870 -140
rect 1790 -190 1870 -170
rect 1400 -260 1480 -240
rect 1400 -290 1420 -260
rect 310 -300 1420 -290
rect 1460 -290 1480 -260
rect 1460 -300 3410 -290
rect 310 -320 3410 -300
rect 310 -688 340 -320
rect 870 -390 2950 -370
rect 870 -430 890 -390
rect 930 -400 2890 -390
rect 930 -430 950 -400
rect 870 -450 950 -430
rect 2870 -430 2890 -400
rect 2930 -430 2950 -390
rect 2870 -450 2950 -430
rect 260 -718 340 -688
rect 750 -718 830 -688
rect 3240 -690 3250 -688
rect 800 -918 830 -718
rect 3230 -720 3330 -690
rect 880 -890 960 -868
rect 880 -918 900 -890
rect 800 -930 900 -918
rect 940 -930 960 -890
rect 800 -948 960 -930
rect 3300 -1020 3330 -720
rect 3380 -810 3410 -320
rect 3380 -830 3460 -810
rect 3380 -870 3400 -830
rect 3440 -870 3460 -830
rect 3380 -890 3460 -870
rect 3300 -1040 3380 -1020
rect 3300 -1080 3320 -1040
rect 3360 -1080 3380 -1040
rect 3300 -1100 3380 -1080
<< polycont >>
rect 3320 580 3360 620
rect 900 430 940 470
rect 1810 250 1850 290
rect 3400 370 3440 410
rect 1810 40 1850 80
rect 890 -40 930 0
rect 2890 -40 2930 0
rect 1810 -170 1850 -130
rect 1420 -300 1460 -260
rect 890 -430 930 -390
rect 2890 -430 2930 -390
rect 900 -930 940 -890
rect 3400 -870 3440 -830
rect 3320 -1080 3360 -1040
<< locali >>
rect 410 620 3380 640
rect 410 600 3320 620
rect 410 340 450 600
rect 3300 580 3320 600
rect 3360 580 3380 620
rect 3300 560 3380 580
rect 880 470 1010 490
rect 880 430 900 470
rect 940 450 1010 470
rect 940 430 960 450
rect 1498 440 1510 480
rect 880 410 960 430
rect 3240 410 3630 430
rect 3240 390 3400 410
rect 3380 370 3400 390
rect 3440 390 3630 410
rect 3440 370 3460 390
rect 3380 350 3460 370
rect 260 300 450 340
rect 750 300 880 340
rect 410 260 450 300
rect 840 260 880 300
rect 1790 290 1870 310
rect -650 220 30 260
rect 410 220 520 260
rect 840 220 1010 260
rect 1240 220 1360 260
rect 910 20 950 220
rect 870 0 950 20
rect 870 -40 890 0
rect 930 -40 950 0
rect 870 -60 950 -40
rect 870 -390 950 -370
rect 870 -430 890 -390
rect 930 -430 950 -390
rect 870 -450 950 -430
rect 910 -678 950 -450
rect 1320 -678 1360 220
rect 1400 220 1502 260
rect 1730 220 1740 260
rect 1790 250 1810 290
rect 1850 250 1870 290
rect 1790 230 1870 250
rect 1960 220 2040 260
rect 2180 220 2530 260
rect 2670 220 2830 260
rect 1400 -240 1440 220
rect 1960 180 2000 220
rect 1730 140 2000 180
rect 1790 80 1870 100
rect 1790 40 1810 80
rect 1850 40 1870 80
rect 1790 20 1870 40
rect 1790 -110 1830 20
rect 1790 -130 1870 -110
rect 1790 -170 1810 -130
rect 1850 -170 1870 -130
rect 1790 -190 1870 -170
rect 1400 -260 1480 -240
rect 1400 -300 1420 -260
rect 1460 -300 1480 -260
rect 1400 -320 1480 -300
rect 2790 -678 2830 220
rect 2910 220 3010 260
rect 2910 20 2950 220
rect 2870 0 2950 20
rect 2870 -40 2890 0
rect 2930 -40 2950 0
rect 2870 -60 2950 -40
rect 2870 -390 2950 -370
rect 2870 -430 2890 -390
rect 2930 -430 2950 -390
rect 2870 -450 2950 -430
rect -650 -720 30 -680
rect 410 -718 520 -678
rect 840 -718 1010 -678
rect 1248 -718 1546 -678
rect 1692 -718 2040 -678
rect 2180 -718 2530 -678
rect 2670 -718 2830 -678
rect 2910 -670 2950 -450
rect 2910 -710 3010 -670
rect 3240 -718 3250 -678
rect 410 -758 450 -718
rect 840 -758 880 -718
rect 2670 -720 2790 -718
rect 260 -798 450 -758
rect 750 -798 880 -758
rect 410 -1058 450 -798
rect 3380 -830 3460 -810
rect 3380 -850 3400 -830
rect 880 -890 960 -868
rect 3240 -870 3400 -850
rect 3440 -850 3460 -830
rect 3440 -870 3630 -850
rect 3240 -890 3630 -870
rect 880 -930 900 -890
rect 940 -908 960 -890
rect 940 -930 1010 -908
rect 880 -948 1010 -930
rect 3300 -1040 3380 -1020
rect 3300 -1058 3320 -1040
rect 410 -1080 3320 -1058
rect 3360 -1080 3380 -1040
rect 410 -1098 3380 -1080
rect 1400 -1100 1480 -1098
rect 3300 -1100 3380 -1098
<< metal1 >>
rect -90 500 10 590
rect 280 500 510 590
rect 770 500 1000 590
rect 1260 500 1490 590
rect 1750 500 1980 590
rect 2240 500 2470 590
rect 2730 500 2990 590
rect -90 -960 -50 500
rect 10 -430 70 -20
rect 280 -50 500 40
rect 770 0 990 40
rect 770 -50 870 0
rect 950 -50 990 0
rect 1260 -50 1480 40
rect 1750 -50 1970 40
rect 2230 -60 3010 50
rect 2210 -410 2470 -400
rect 2730 -410 3010 -400
rect 280 -500 500 -410
rect 770 -500 990 -410
rect 1260 -500 1480 -410
rect 1750 -500 1970 -410
rect 2210 -500 3010 -410
rect 2210 -510 2480 -500
rect 2720 -510 3010 -500
rect -90 -1050 39 -960
rect 280 -1050 500 -960
rect 770 -1050 990 -960
rect 1260 -1050 1480 -960
rect 1750 -1050 1970 -960
rect 2240 -1050 2460 -960
rect 2730 -1050 2990 -960
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 2246 0 -1 -456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1723858470
transform -1 0 1756 0 -1 -456
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1723858470
transform 1 0 1970 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1723858470
transform 1 0 2460 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1723858470
transform -1 0 2736 0 -1 -456
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1480 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 286 0 -1 -456
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_1
timestamp 1723858470
transform -1 0 3266 0 -1 -456
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_2
timestamp 1723858470
transform -1 0 776 0 -1 -456
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_3
timestamp 1723858470
transform 1 0 990 0 -1 -456
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_4
timestamp 1723858470
transform -1 0 286 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_5
timestamp 1723858470
transform -1 0 776 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_6
timestamp 1723858470
transform 1 0 990 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  sky130_fd_sc_hd__nor2_1_7
timestamp 1723858470
transform -1 0 3266 0 1 0
box -38 -48 314 592
<< labels >>
flabel locali -650 240 -650 240 7 FreeSans 320 0 -160 0 F_REF
port 1 w
flabel locali -650 -700 -650 -700 7 FreeSans 320 0 -160 0 F_VCO
port 2 w
flabel locali 3630 -870 3630 -870 3 FreeSans 320 0 160 0 QB
port 4 e
flabel locali 3630 410 3630 410 3 FreeSans 320 0 160 0 QA
port 3 e
flabel metal1 -90 590 -90 590 7 FreeSans 320 0 -160 0 VDDA
port 5 w
flabel metal1 70 -230 70 -230 3 FreeSans 320 0 160 0 GNDA
port 6 e
<< end >>
