magic
tech sky130A
timestamp 1738032933
<< nwell >>
rect 1045 150 1935 2565
<< nmos >>
rect 1140 -175 1155 -75
rect 1295 -175 1310 -75
rect 1515 -175 1530 -75
rect 1670 -175 1685 -75
rect 1845 -175 1860 -75
rect 1615 -1320 1665 -320
rect 1815 -1320 1865 -320
<< pmos >>
rect 1115 510 1165 2510
rect 1315 510 1365 2510
rect 1140 175 1155 375
rect 1295 175 1310 375
rect 1515 175 1530 375
rect 1670 175 1685 375
rect 1845 175 1860 375
<< ndiff >>
rect 1090 -90 1140 -75
rect 1090 -160 1105 -90
rect 1125 -160 1140 -90
rect 1090 -175 1140 -160
rect 1155 -90 1205 -75
rect 1155 -160 1170 -90
rect 1190 -160 1205 -90
rect 1155 -175 1205 -160
rect 1245 -90 1295 -75
rect 1245 -160 1260 -90
rect 1280 -160 1295 -90
rect 1245 -175 1295 -160
rect 1310 -90 1360 -75
rect 1310 -160 1325 -90
rect 1345 -160 1360 -90
rect 1465 -90 1515 -75
rect 1310 -175 1360 -160
rect 1465 -160 1480 -90
rect 1500 -160 1515 -90
rect 1465 -175 1515 -160
rect 1530 -90 1580 -75
rect 1530 -160 1545 -90
rect 1565 -160 1580 -90
rect 1530 -175 1580 -160
rect 1620 -90 1670 -75
rect 1620 -160 1635 -90
rect 1655 -160 1670 -90
rect 1620 -175 1670 -160
rect 1685 -90 1735 -75
rect 1685 -160 1700 -90
rect 1720 -160 1735 -90
rect 1685 -175 1735 -160
rect 1795 -90 1845 -75
rect 1795 -160 1810 -90
rect 1830 -160 1845 -90
rect 1795 -175 1845 -160
rect 1860 -90 1910 -75
rect 1860 -160 1875 -90
rect 1895 -160 1910 -90
rect 1860 -175 1910 -160
rect 1565 -335 1615 -320
rect 1565 -1305 1580 -335
rect 1600 -1305 1615 -335
rect 1565 -1320 1615 -1305
rect 1665 -335 1715 -320
rect 1665 -1305 1680 -335
rect 1700 -1305 1715 -335
rect 1665 -1320 1715 -1305
rect 1765 -335 1815 -320
rect 1765 -1305 1780 -335
rect 1800 -1305 1815 -335
rect 1765 -1320 1815 -1305
rect 1865 -335 1915 -320
rect 1865 -1305 1880 -335
rect 1900 -1305 1915 -335
rect 1865 -1320 1915 -1305
<< pdiff >>
rect 1065 2495 1115 2510
rect 1065 525 1080 2495
rect 1100 525 1115 2495
rect 1065 510 1115 525
rect 1165 2495 1215 2510
rect 1165 525 1180 2495
rect 1200 525 1215 2495
rect 1165 510 1215 525
rect 1265 2495 1315 2510
rect 1265 525 1280 2495
rect 1300 525 1315 2495
rect 1265 510 1315 525
rect 1365 2495 1415 2510
rect 1365 525 1380 2495
rect 1400 525 1415 2495
rect 1365 510 1415 525
rect 1090 360 1140 375
rect 1090 190 1105 360
rect 1125 190 1140 360
rect 1090 175 1140 190
rect 1155 360 1205 375
rect 1155 190 1170 360
rect 1190 190 1205 360
rect 1155 175 1205 190
rect 1245 360 1295 375
rect 1245 190 1260 360
rect 1280 190 1295 360
rect 1245 175 1295 190
rect 1310 360 1360 375
rect 1310 190 1325 360
rect 1345 190 1360 360
rect 1310 175 1360 190
rect 1465 360 1515 375
rect 1465 190 1480 360
rect 1500 190 1515 360
rect 1465 175 1515 190
rect 1530 360 1580 375
rect 1530 190 1545 360
rect 1565 190 1580 360
rect 1530 175 1580 190
rect 1620 360 1670 375
rect 1620 190 1635 360
rect 1655 190 1670 360
rect 1620 175 1670 190
rect 1685 360 1735 375
rect 1685 190 1700 360
rect 1720 190 1735 360
rect 1685 175 1735 190
rect 1795 360 1845 375
rect 1795 190 1810 360
rect 1830 190 1845 360
rect 1795 175 1845 190
rect 1860 360 1910 375
rect 1860 190 1875 360
rect 1895 190 1910 360
rect 1860 175 1910 190
<< ndiffc >>
rect 1105 -160 1125 -90
rect 1170 -160 1190 -90
rect 1260 -160 1280 -90
rect 1325 -160 1345 -90
rect 1480 -160 1500 -90
rect 1545 -160 1565 -90
rect 1635 -160 1655 -90
rect 1700 -160 1720 -90
rect 1810 -160 1830 -90
rect 1875 -160 1895 -90
rect 1580 -1305 1600 -335
rect 1680 -1305 1700 -335
rect 1780 -1305 1800 -335
rect 1880 -1305 1900 -335
<< pdiffc >>
rect 1080 525 1100 2495
rect 1180 525 1200 2495
rect 1280 525 1300 2495
rect 1380 525 1400 2495
rect 1105 190 1125 360
rect 1170 190 1190 360
rect 1260 190 1280 360
rect 1325 190 1345 360
rect 1480 190 1500 360
rect 1545 190 1565 360
rect 1635 190 1655 360
rect 1700 190 1720 360
rect 1810 190 1830 360
rect 1875 190 1895 360
<< poly >>
rect 1115 2510 1165 2525
rect 1315 2510 1365 2525
rect 1115 500 1165 510
rect 1315 500 1365 510
rect 1115 480 1365 500
rect 1115 460 1130 480
rect 1150 475 1365 480
rect 1150 460 1165 475
rect 855 435 1070 450
rect 1115 445 1165 460
rect 1055 405 1070 435
rect 1055 390 1155 405
rect 1055 345 1070 390
rect 1140 375 1155 390
rect 1295 375 1310 390
rect 1515 375 1530 390
rect 1670 375 1685 390
rect 1845 375 1860 390
rect 625 330 1070 345
rect 625 -230 640 330
rect 1140 160 1155 175
rect 1295 85 1310 175
rect 1515 165 1530 175
rect 1670 165 1685 175
rect 1515 160 1685 165
rect 1845 160 1860 175
rect 1480 145 1685 160
rect 1805 145 1860 160
rect 1480 125 1495 145
rect 1515 125 1530 145
rect 1480 110 1530 125
rect 1805 125 1820 145
rect 1840 125 1860 145
rect 1805 110 1860 125
rect 1395 90 1445 105
rect 1395 85 1410 90
rect 1005 70 1410 85
rect 1430 70 1445 90
rect 1005 -35 1020 70
rect 1395 55 1445 70
rect 1325 10 1375 25
rect 1325 -10 1340 10
rect 1360 5 1375 10
rect 1360 -10 1860 5
rect 860 -50 1020 -35
rect 1105 -25 1155 -10
rect 1325 -25 1375 -10
rect 1105 -45 1120 -25
rect 1140 -45 1155 -25
rect 1105 -50 1155 -45
rect 1105 -60 1310 -50
rect 1140 -65 1310 -60
rect 1140 -75 1155 -65
rect 1295 -75 1310 -65
rect 1515 -75 1530 -60
rect 1670 -75 1685 -60
rect 1845 -75 1860 -10
rect 1400 -165 1450 -150
rect 1140 -190 1155 -175
rect 1295 -190 1310 -175
rect 1400 -185 1415 -165
rect 1435 -185 1450 -165
rect 1515 -185 1530 -175
rect 1400 -200 1530 -185
rect 1670 -230 1685 -175
rect 1845 -190 1860 -175
rect 625 -245 1685 -230
rect 1615 -320 1665 -305
rect 1815 -320 1865 -305
rect 1615 -1330 1665 -1320
rect 1815 -1330 1865 -1320
rect 1615 -1340 1865 -1330
rect 1615 -1350 1630 -1340
rect 1620 -1360 1630 -1350
rect 1650 -1350 1865 -1340
rect 1650 -1360 1660 -1350
rect 1620 -1370 1660 -1360
<< polycont >>
rect 1130 460 1150 480
rect 1495 125 1515 145
rect 1820 125 1840 145
rect 1410 70 1430 90
rect 1340 -10 1360 10
rect 1120 -45 1140 -25
rect 1415 -185 1435 -165
rect 1630 -1360 1650 -1340
<< xpolycontact >>
rect 2070 745 2105 965
rect 2070 410 2105 630
rect 2070 -230 2105 -10
rect 1020 -605 1240 -320
rect 1290 -605 1510 -320
rect 2070 -535 2105 -315
<< xpolyres >>
rect 2070 630 2105 745
rect 2070 -315 2105 -230
rect 1240 -605 1290 -320
<< locali >>
rect 1070 2495 1110 2505
rect 1070 525 1080 2495
rect 1100 525 1110 2495
rect 1070 515 1110 525
rect 1170 2495 1210 2505
rect 1170 525 1180 2495
rect 1200 525 1210 2495
rect 1170 515 1210 525
rect 1270 2495 1310 2505
rect 1270 525 1280 2495
rect 1300 525 1310 2495
rect 1270 515 1310 525
rect 1370 2495 1410 2505
rect 1370 525 1380 2495
rect 1400 525 1410 2495
rect 2125 1070 2165 1080
rect 2085 1050 2135 1070
rect 2155 1050 2165 1070
rect 2085 965 2105 1050
rect 2125 1040 2165 1050
rect 1370 515 1410 525
rect 1080 495 1100 515
rect 965 480 1165 495
rect 965 475 1130 480
rect 965 -320 985 475
rect 1115 460 1130 475
rect 1150 460 1165 480
rect 1115 445 1165 460
rect 1380 415 1400 515
rect 1170 395 1400 415
rect 1170 370 1190 395
rect 1260 370 1280 395
rect 1095 360 1135 370
rect 1095 190 1105 360
rect 1125 190 1135 360
rect 1095 180 1135 190
rect 1160 360 1200 370
rect 1160 190 1170 360
rect 1190 190 1200 360
rect 1160 180 1200 190
rect 1250 360 1290 370
rect 1250 190 1260 360
rect 1280 190 1290 360
rect 1250 180 1290 190
rect 1315 360 1355 370
rect 1315 190 1325 360
rect 1345 190 1355 360
rect 1315 180 1355 190
rect 1470 360 1510 370
rect 1470 190 1480 360
rect 1500 190 1510 360
rect 1470 180 1510 190
rect 1535 360 1575 370
rect 1535 190 1545 360
rect 1565 190 1575 360
rect 1535 180 1575 190
rect 1625 360 1665 370
rect 1625 190 1635 360
rect 1655 190 1665 360
rect 1625 180 1665 190
rect 1690 360 1730 370
rect 1690 190 1700 360
rect 1720 190 1730 360
rect 1690 180 1730 190
rect 1800 360 1840 370
rect 1800 190 1810 360
rect 1830 190 1840 360
rect 1800 180 1840 190
rect 1865 360 1905 370
rect 1865 190 1875 360
rect 1895 190 1905 360
rect 2085 240 2105 410
rect 1865 180 1905 190
rect 1975 220 2105 240
rect 2125 305 2165 315
rect 2125 285 2135 305
rect 2155 285 2165 305
rect 2125 275 2165 285
rect 1105 -10 1125 180
rect 1325 25 1345 180
rect 1480 160 1500 180
rect 1700 160 1720 180
rect 1480 145 1530 160
rect 1480 125 1495 145
rect 1515 125 1530 145
rect 1480 110 1530 125
rect 1700 145 1855 160
rect 1700 140 1820 145
rect 1395 90 1445 105
rect 1395 70 1410 90
rect 1430 70 1445 90
rect 1395 55 1445 70
rect 1325 10 1375 25
rect 1325 -10 1340 10
rect 1360 -10 1375 10
rect 1105 -25 1155 -10
rect 1105 -45 1120 -25
rect 1140 -45 1155 -25
rect 1105 -60 1155 -45
rect 1325 -25 1375 -10
rect 1105 -80 1125 -60
rect 1325 -80 1345 -25
rect 1095 -90 1135 -80
rect 1095 -160 1105 -90
rect 1125 -160 1135 -90
rect 1095 -170 1135 -160
rect 1160 -90 1200 -80
rect 1160 -160 1170 -90
rect 1190 -160 1200 -90
rect 1160 -170 1200 -160
rect 1250 -90 1290 -80
rect 1250 -160 1260 -90
rect 1280 -160 1290 -90
rect 1250 -170 1290 -160
rect 1315 -90 1355 -80
rect 1315 -160 1325 -90
rect 1345 -160 1355 -90
rect 1415 -150 1435 55
rect 1480 -80 1500 110
rect 1700 -80 1720 140
rect 1805 125 1820 140
rect 1840 125 1855 145
rect 1875 150 1895 180
rect 1975 150 1995 220
rect 1875 130 1995 150
rect 2125 185 2145 275
rect 2125 165 3055 185
rect 1805 110 1855 125
rect 2125 70 2145 165
rect 2125 60 2165 70
rect 2125 40 2135 60
rect 2155 40 2165 60
rect 1875 15 2105 35
rect 2125 30 2165 40
rect 1875 -80 1895 15
rect 2085 -10 2105 15
rect 1470 -90 1510 -80
rect 1315 -170 1355 -160
rect 1400 -165 1450 -150
rect 1400 -185 1415 -165
rect 1435 -185 1450 -165
rect 1470 -160 1480 -90
rect 1500 -160 1510 -90
rect 1470 -170 1510 -160
rect 1535 -90 1575 -80
rect 1535 -160 1545 -90
rect 1565 -160 1575 -90
rect 1535 -170 1575 -160
rect 1625 -90 1665 -80
rect 1625 -160 1635 -90
rect 1655 -160 1665 -90
rect 1625 -170 1665 -160
rect 1690 -90 1730 -80
rect 1690 -160 1700 -90
rect 1720 -160 1730 -90
rect 1690 -170 1730 -160
rect 1800 -90 1840 -80
rect 1800 -160 1810 -90
rect 1830 -160 1840 -90
rect 1800 -170 1840 -160
rect 1865 -90 1905 -80
rect 1865 -160 1875 -90
rect 1895 -160 1905 -90
rect 1865 -170 1905 -160
rect 1400 -200 1450 -185
rect 1545 -215 1565 -170
rect 1635 -215 1655 -170
rect 1545 -235 1800 -215
rect 1780 -270 1800 -235
rect 1780 -290 1900 -270
rect 965 -340 1020 -320
rect 1880 -325 1900 -290
rect 1570 -335 1610 -325
rect 1510 -1335 1530 -585
rect 1570 -1305 1580 -335
rect 1600 -1305 1610 -335
rect 1570 -1315 1610 -1305
rect 1670 -335 1710 -325
rect 1670 -1305 1680 -335
rect 1700 -1305 1710 -335
rect 1670 -1315 1710 -1305
rect 1770 -335 1810 -325
rect 1770 -1305 1780 -335
rect 1800 -1305 1810 -335
rect 1770 -1315 1810 -1305
rect 1870 -335 1910 -325
rect 1870 -1305 1880 -335
rect 1900 -1305 1910 -335
rect 2085 -705 2105 -535
rect 2125 -705 2165 -695
rect 2085 -725 2135 -705
rect 2155 -725 2165 -705
rect 2125 -735 2165 -725
rect 1870 -1315 1910 -1305
rect 1580 -1335 1600 -1315
rect 1620 -1335 1660 -1330
rect 1510 -1340 1665 -1335
rect 1510 -1355 1630 -1340
rect 1620 -1360 1630 -1355
rect 1650 -1355 1665 -1340
rect 1650 -1360 1660 -1355
rect 1620 -1370 1660 -1360
<< viali >>
rect 1180 525 1200 2495
rect 1280 525 1300 2495
rect 2135 1050 2155 1070
rect 1545 190 1565 360
rect 1635 190 1655 360
rect 1810 190 1830 360
rect 2135 285 2155 305
rect 1170 -160 1190 -90
rect 1260 -160 1280 -90
rect 2135 40 2155 60
rect 1810 -160 1830 -90
rect 1680 -1305 1700 -335
rect 1780 -1305 1800 -335
rect 2135 -725 2155 -705
<< metal1 >>
rect 1015 2495 1955 2565
rect 1015 525 1180 2495
rect 1200 525 1280 2495
rect 1300 525 1955 2495
rect 2125 1070 2165 1080
rect 2125 1050 2135 1070
rect 2155 1050 2165 1070
rect 2125 1040 2165 1050
rect 1015 360 1955 525
rect 1015 190 1545 360
rect 1565 190 1635 360
rect 1655 190 1810 360
rect 1830 190 1955 360
rect 2125 305 2165 315
rect 2125 285 2135 305
rect 2155 285 2165 305
rect 2125 275 2165 285
rect 1015 150 1955 190
rect 2125 60 2165 70
rect 2125 40 2135 60
rect 2155 40 2165 60
rect 2125 30 2165 40
rect 1015 -90 1955 -35
rect 1015 -160 1170 -90
rect 1190 -160 1260 -90
rect 1280 -160 1810 -90
rect 1830 -160 1955 -90
rect 1015 -335 1955 -160
rect 1015 -645 1680 -335
rect 1560 -1305 1680 -645
rect 1700 -1305 1780 -335
rect 1800 -645 1955 -335
rect 1800 -1305 1920 -645
rect 2125 -705 2165 -695
rect 2125 -725 2135 -705
rect 2155 -725 2165 -705
rect 2125 -735 2165 -725
rect 1560 -1375 1920 -1305
<< metal3 >>
rect 2125 1040 3010 1085
rect 2180 255 3010 1040
rect 2180 -695 3010 90
rect 2125 -740 3010 -695
<< mimcap >>
rect 2195 315 2995 1070
rect 2195 280 2205 315
rect 2240 280 2995 315
rect 2195 270 2995 280
rect 2195 65 2995 75
rect 2195 30 2205 65
rect 2240 30 2995 65
rect 2195 -725 2995 30
<< mimcapcontact >>
rect 2205 280 2240 315
rect 2205 30 2240 65
<< metal4 >>
rect 2125 315 2245 320
rect 2125 280 2205 315
rect 2240 280 2245 315
rect 2125 275 2245 280
rect 2125 65 2245 70
rect 2125 30 2205 65
rect 2240 30 2245 65
rect 2125 25 2245 30
<< labels >>
flabel locali 3055 170 3055 170 3 FreeSans 400 0 0 0 VOUT
flabel poly 860 -40 860 -40 7 FreeSans 400 0 0 0 VIN-
flabel metal1 1015 -260 1015 -260 7 FreeSans 400 0 0 0 GNDA
flabel poly 855 440 855 440 7 FreeSans 400 0 0 0 VIN+
flabel metal1 1015 795 1015 795 7 FreeSans 400 0 0 0 VDDA
<< end >>
