magic
tech sky130A
timestamp 1753588328
<< metal1 >>
rect 2950 6685 2990 6690
rect 2950 6655 2955 6685
rect 2985 6655 2990 6685
rect 2950 6650 2990 6655
rect 3030 6685 3070 6690
rect 3030 6655 3035 6685
rect 3065 6655 3070 6685
rect 6045 6685 6085 6690
rect 6045 6655 6050 6685
rect 6080 6655 6085 6685
rect 3030 6650 3070 6655
rect 2905 6580 2945 6585
rect 2905 6550 2910 6580
rect 2940 6550 2945 6580
rect 2905 6545 2945 6550
rect 2915 2710 2935 6545
rect 2960 2505 2980 6650
rect 3280 6525 3300 6650
rect 3400 6645 3440 6650
rect 3400 6615 3405 6645
rect 3435 6615 3440 6645
rect 3400 6610 3440 6615
rect 3270 6520 3310 6525
rect 3270 6490 3275 6520
rect 3305 6490 3310 6520
rect 3270 6485 3310 6490
rect 3555 6480 3575 6655
rect 3955 6645 3995 6650
rect 3955 6615 3960 6645
rect 3990 6615 3995 6645
rect 3955 6610 3995 6615
rect 3545 6475 3585 6480
rect 3545 6445 3550 6475
rect 3580 6445 3585 6475
rect 3545 6440 3585 6445
rect 3965 3360 3985 6610
rect 4340 6585 4360 6655
rect 4330 6580 4370 6585
rect 4330 6550 4335 6580
rect 4365 6550 4370 6580
rect 4330 6545 4370 6550
rect 4005 6475 4045 6480
rect 4005 6445 4010 6475
rect 4040 6445 4045 6475
rect 4005 6440 4045 6445
rect 3955 3355 3995 3360
rect 3955 3325 3960 3355
rect 3990 3325 3995 3355
rect 3955 3320 3995 3325
rect 4015 2790 4035 6440
rect 5085 5465 5105 6655
rect 5730 6585 5750 6655
rect 6045 6650 6085 6655
rect 6700 6685 6740 6690
rect 6700 6655 6705 6685
rect 6735 6655 6740 6685
rect 7020 6685 7060 6690
rect 7020 6655 7025 6685
rect 7055 6655 7060 6685
rect 6700 6650 6740 6655
rect 5720 6580 5760 6585
rect 5720 6550 5725 6580
rect 5755 6550 5760 6580
rect 5720 6545 5760 6550
rect 5375 6520 5415 6525
rect 5375 6490 5380 6520
rect 5410 6490 5415 6520
rect 5375 6485 5415 6490
rect 5075 5460 5115 5465
rect 5075 5430 5080 5460
rect 5110 5430 5115 5460
rect 5075 5425 5115 5430
rect 5385 5420 5405 6485
rect 5375 5415 5415 5420
rect 5375 5385 5380 5415
rect 5410 5385 5415 5415
rect 5375 5380 5415 5385
rect 5495 5415 5535 5420
rect 5495 5385 5500 5415
rect 5530 5385 5535 5415
rect 5495 5380 5535 5385
rect 5505 4805 5525 5380
rect 5495 4800 5535 4805
rect 5495 4770 5500 4800
rect 5530 4770 5535 4800
rect 5495 4765 5535 4770
rect 6055 3640 6075 6650
rect 6100 5460 6140 5465
rect 6100 5430 6105 5460
rect 6135 5430 6140 5460
rect 6785 5440 6805 6655
rect 7020 6650 7060 6655
rect 7100 6685 7140 6690
rect 7100 6655 7105 6685
rect 7135 6655 7140 6685
rect 7100 6650 7140 6655
rect 6100 5425 6140 5430
rect 6425 5435 6465 5440
rect 6045 3635 6085 3640
rect 4970 3630 5010 3635
rect 4970 3600 4975 3630
rect 5005 3600 5010 3630
rect 6045 3605 6050 3635
rect 6080 3605 6085 3635
rect 6045 3600 6085 3605
rect 4970 3595 5010 3600
rect 6110 2880 6130 5425
rect 6425 5405 6430 5435
rect 6460 5405 6465 5435
rect 6425 5400 6465 5405
rect 6775 5435 6815 5440
rect 6775 5405 6780 5435
rect 6810 5405 6815 5435
rect 6775 5400 6815 5405
rect 6435 4870 6455 5400
rect 6425 4865 6465 4870
rect 6425 4835 6430 4865
rect 6460 4835 6465 4865
rect 6425 4830 6465 4835
rect 5085 2875 5125 2880
rect 5085 2845 5090 2875
rect 5120 2845 5125 2875
rect 5085 2840 5125 2845
rect 6100 2875 6140 2880
rect 6100 2845 6105 2875
rect 6135 2845 6140 2875
rect 6100 2840 6140 2845
rect 5095 2410 5115 2840
rect 7110 2505 7130 6650
rect 7145 6580 7185 6585
rect 7145 6550 7150 6580
rect 7180 6550 7185 6580
rect 7145 6545 7185 6550
rect 7155 2710 7175 6545
rect 2440 1800 2480 1830
<< via1 >>
rect 2955 6655 2985 6685
rect 3035 6655 3065 6685
rect 6050 6655 6080 6685
rect 2910 6550 2940 6580
rect 3405 6615 3435 6645
rect 3275 6490 3305 6520
rect 3960 6615 3990 6645
rect 3550 6445 3580 6475
rect 4335 6550 4365 6580
rect 4010 6445 4040 6475
rect 3960 3325 3990 3355
rect 6705 6655 6735 6685
rect 7025 6655 7055 6685
rect 5725 6550 5755 6580
rect 5380 6490 5410 6520
rect 5080 5430 5110 5460
rect 5380 5385 5410 5415
rect 5500 5385 5530 5415
rect 5500 4770 5530 4800
rect 6105 5430 6135 5460
rect 7105 6655 7135 6685
rect 4975 3600 5005 3630
rect 6050 3605 6080 3635
rect 6430 5405 6460 5435
rect 6780 5405 6810 5435
rect 6430 4835 6460 4865
rect 5090 2845 5120 2875
rect 6105 2845 6135 2875
rect 7150 6550 7180 6580
<< metal2 >>
rect 2950 6685 2990 6690
rect 2950 6655 2955 6685
rect 2985 6680 2990 6685
rect 3030 6685 3070 6690
rect 3030 6680 3035 6685
rect 2985 6660 3035 6680
rect 2985 6655 2990 6660
rect 2950 6650 2990 6655
rect 3030 6655 3035 6660
rect 3065 6655 3070 6685
rect 3030 6650 3070 6655
rect 6045 6685 6085 6690
rect 6045 6655 6050 6685
rect 6080 6680 6085 6685
rect 6700 6685 6740 6690
rect 6700 6680 6705 6685
rect 6080 6660 6705 6680
rect 6080 6655 6085 6660
rect 6045 6650 6085 6655
rect 6700 6655 6705 6660
rect 6735 6655 6740 6685
rect 7020 6685 7060 6690
rect 7020 6680 7025 6685
rect 7010 6660 7025 6680
rect 6700 6650 6740 6655
rect 7020 6655 7025 6660
rect 7055 6680 7060 6685
rect 7100 6685 7140 6690
rect 7100 6680 7105 6685
rect 7055 6660 7105 6680
rect 7055 6655 7060 6660
rect 7020 6650 7060 6655
rect 7100 6655 7105 6660
rect 7135 6655 7140 6685
rect 7100 6650 7140 6655
rect 3400 6645 3440 6650
rect 3400 6615 3405 6645
rect 3435 6640 3440 6645
rect 3955 6645 3995 6650
rect 3955 6640 3960 6645
rect 3435 6620 3960 6640
rect 3435 6615 3440 6620
rect 3400 6610 3440 6615
rect 3955 6615 3960 6620
rect 3990 6615 3995 6645
rect 3955 6610 3995 6615
rect 2905 6580 2945 6585
rect 2905 6550 2910 6580
rect 2940 6575 2945 6580
rect 4330 6580 4370 6585
rect 4330 6575 4335 6580
rect 2940 6555 4335 6575
rect 2940 6550 2945 6555
rect 2905 6545 2945 6550
rect 4330 6550 4335 6555
rect 4365 6550 4370 6580
rect 4330 6545 4370 6550
rect 5720 6580 5760 6585
rect 5720 6550 5725 6580
rect 5755 6575 5760 6580
rect 7145 6580 7185 6585
rect 7145 6575 7150 6580
rect 5755 6555 7150 6575
rect 5755 6550 5760 6555
rect 5720 6545 5760 6550
rect 7145 6550 7150 6555
rect 7180 6550 7185 6580
rect 7145 6545 7185 6550
rect 3270 6520 3310 6525
rect 3270 6490 3275 6520
rect 3305 6515 3310 6520
rect 5375 6520 5415 6525
rect 5375 6515 5380 6520
rect 3305 6495 5380 6515
rect 3305 6490 3310 6495
rect 3270 6485 3310 6490
rect 5375 6490 5380 6495
rect 5410 6490 5415 6520
rect 5375 6485 5415 6490
rect 3545 6475 3585 6480
rect 3545 6445 3550 6475
rect 3580 6470 3585 6475
rect 4005 6475 4045 6480
rect 4005 6470 4010 6475
rect 3580 6450 4010 6470
rect 3580 6445 3585 6450
rect 3545 6440 3585 6445
rect 4005 6445 4010 6450
rect 4040 6445 4045 6475
rect 4005 6440 4045 6445
rect 5075 5460 5115 5465
rect 5075 5430 5080 5460
rect 5110 5455 5115 5460
rect 6100 5460 6140 5465
rect 6100 5455 6105 5460
rect 5110 5435 6105 5455
rect 5110 5430 5115 5435
rect 5075 5425 5115 5430
rect 6100 5430 6105 5435
rect 6135 5430 6140 5460
rect 6100 5425 6140 5430
rect 6425 5435 6465 5440
rect 5375 5415 5415 5420
rect 5375 5385 5380 5415
rect 5410 5410 5415 5415
rect 5495 5415 5535 5420
rect 5495 5410 5500 5415
rect 5410 5390 5500 5410
rect 5410 5385 5415 5390
rect 5375 5380 5415 5385
rect 5495 5385 5500 5390
rect 5530 5385 5535 5415
rect 6425 5405 6430 5435
rect 6460 5430 6465 5435
rect 6775 5435 6815 5440
rect 6775 5430 6780 5435
rect 6460 5410 6780 5430
rect 6460 5405 6465 5410
rect 6425 5400 6465 5405
rect 6775 5405 6780 5410
rect 6810 5405 6815 5435
rect 6775 5400 6815 5405
rect 5495 5380 5535 5385
rect 6425 4865 6465 4870
rect 6425 4860 6430 4865
rect 5750 4840 6430 4860
rect 6425 4835 6430 4840
rect 6460 4835 6465 4865
rect 6425 4830 6465 4835
rect 5495 4800 5535 4805
rect 5495 4770 5500 4800
rect 5530 4770 5535 4800
rect 5495 4765 5535 4770
rect 6045 3635 6085 3640
rect 4970 3630 5010 3635
rect 4970 3600 4975 3630
rect 5005 3625 5010 3630
rect 6045 3625 6050 3635
rect 5005 3605 6050 3625
rect 6080 3605 6085 3635
rect 5005 3600 5010 3605
rect 6045 3600 6085 3605
rect 4970 3595 5010 3600
rect 3955 3355 3995 3360
rect 3955 3325 3960 3355
rect 3990 3340 3995 3355
rect 3990 3325 4115 3340
rect 3955 3320 4115 3325
rect 5085 2875 5125 2880
rect 5085 2845 5090 2875
rect 5120 2870 5125 2875
rect 6100 2875 6140 2880
rect 6100 2870 6105 2875
rect 5120 2850 6105 2870
rect 5120 2845 5125 2850
rect 5085 2840 5125 2845
rect 6100 2845 6105 2850
rect 6135 2845 6140 2875
rect 6100 2840 6140 2845
rect 4160 2315 4180 2335
rect 5910 2315 5930 2335
rect 2440 1800 2480 1830
rect 2645 1785 2665 1805
rect 7380 1785 7400 1805
<< metal3 >>
rect 10185 14460 10235 14465
rect 10185 14420 10190 14460
rect 10230 14420 10235 14460
rect 10185 14415 10235 14420
rect 10190 50 10230 14415
rect 10405 14100 10635 14185
rect 10755 14100 10985 14185
rect 11105 14100 11335 14185
rect 11455 14100 11685 14185
rect 11805 14100 12035 14185
rect 10405 14050 12035 14100
rect 10405 13955 10635 14050
rect 10755 13955 10985 14050
rect 11105 13955 11335 14050
rect 11455 13955 11685 14050
rect 11805 13955 12035 14050
rect 11195 13835 11245 13955
rect 10405 13750 10635 13835
rect 10755 13750 10985 13835
rect 11105 13750 11335 13835
rect 11455 13750 11685 13835
rect 11805 13750 12035 13835
rect 10405 13700 12035 13750
rect 10405 13605 10635 13700
rect 10755 13605 10985 13700
rect 11105 13605 11335 13700
rect 11455 13605 11685 13700
rect 11805 13605 12035 13700
rect 11195 13485 11245 13605
rect 10405 13400 10635 13485
rect 10755 13400 10985 13485
rect 11105 13400 11335 13485
rect 11455 13400 11685 13485
rect 11805 13400 12035 13485
rect 10405 13350 12035 13400
rect 10405 13255 10635 13350
rect 10755 13255 10985 13350
rect 11105 13255 11335 13350
rect 11455 13255 11685 13350
rect 11805 13255 12035 13350
rect 11195 13135 11245 13255
rect 10405 13050 10635 13135
rect 10755 13050 10985 13135
rect 11105 13050 11335 13135
rect 11455 13050 11685 13135
rect 11805 13050 12035 13135
rect 10405 13000 12035 13050
rect 10405 12905 10635 13000
rect 10755 12905 10985 13000
rect 11105 12905 11335 13000
rect 11455 12905 11685 13000
rect 11805 12905 12035 13000
rect 11195 12785 11245 12905
rect 10405 12700 10635 12785
rect 10755 12700 10985 12785
rect 11105 12700 11335 12785
rect 11455 12700 11685 12785
rect 11805 12700 12035 12785
rect 10405 12650 12035 12700
rect 10405 12555 10635 12650
rect 10755 12555 10985 12650
rect 11105 12555 11335 12650
rect 11455 12555 11685 12650
rect 11805 12555 12035 12650
rect 11195 12435 11245 12555
rect 10405 12350 10635 12435
rect 10755 12350 10985 12435
rect 11105 12350 11335 12435
rect 11455 12350 11685 12435
rect 11805 12350 12035 12435
rect 10405 12300 12035 12350
rect 10405 12205 10635 12300
rect 10755 12205 10985 12300
rect 11105 12205 11335 12300
rect 11455 12205 11685 12300
rect 11805 12205 12035 12300
rect 11195 12085 11245 12205
rect 10405 12000 10635 12085
rect 10755 12000 10985 12085
rect 11105 12000 11335 12085
rect 11455 12000 11685 12085
rect 11805 12000 12035 12085
rect 10405 11950 12035 12000
rect 10405 11855 10635 11950
rect 10755 11855 10985 11950
rect 11105 11855 11335 11950
rect 11455 11855 11685 11950
rect 11805 11855 12035 11950
rect 11195 11735 11245 11855
rect 10405 11650 10635 11735
rect 10755 11650 10985 11735
rect 11105 11650 11335 11735
rect 11455 11650 11685 11735
rect 11805 11650 12035 11735
rect 10405 11600 12035 11650
rect 10405 11505 10635 11600
rect 10755 11505 10985 11600
rect 11105 11505 11335 11600
rect 11455 11505 11685 11600
rect 11805 11505 12035 11600
rect 11195 11385 11245 11505
rect 10405 11300 10635 11385
rect 10755 11300 10985 11385
rect 11105 11300 11335 11385
rect 11455 11300 11685 11385
rect 11805 11300 12035 11385
rect 10405 11250 12035 11300
rect 10405 11155 10635 11250
rect 10755 11155 10985 11250
rect 11105 11155 11335 11250
rect 11455 11155 11685 11250
rect 11805 11155 12035 11250
rect 11195 11035 11245 11155
rect 10405 10950 10635 11035
rect 10755 10950 10985 11035
rect 11105 10950 11335 11035
rect 11455 10950 11685 11035
rect 11805 10950 12035 11035
rect 10405 10900 12035 10950
rect 10405 10805 10635 10900
rect 10755 10805 10985 10900
rect 11105 10805 11335 10900
rect 11455 10805 11685 10900
rect 11805 10805 12035 10900
rect 11195 10685 11245 10805
rect 10405 10600 10635 10685
rect 10755 10600 10985 10685
rect 11105 10600 11335 10685
rect 11455 10600 11685 10685
rect 11805 10600 12035 10685
rect 10405 10550 12035 10600
rect 10405 10455 10635 10550
rect 10755 10455 10985 10550
rect 11105 10455 11335 10550
rect 11455 10455 11685 10550
rect 11805 10455 12035 10550
rect 11195 10335 11245 10455
rect 10405 10250 10635 10335
rect 10755 10250 10985 10335
rect 11105 10250 11335 10335
rect 11455 10250 11685 10335
rect 11805 10250 12035 10335
rect 10405 10200 12035 10250
rect 10405 10105 10635 10200
rect 10755 10105 10985 10200
rect 11105 10105 11335 10200
rect 11455 10105 11685 10200
rect 11805 10105 12035 10200
rect 11195 9985 11245 10105
rect 10405 9900 10635 9985
rect 10755 9900 10985 9985
rect 11105 9900 11335 9985
rect 11455 9900 11685 9985
rect 11805 9900 12035 9985
rect 10405 9850 12035 9900
rect 10405 9755 10635 9850
rect 10755 9755 10985 9850
rect 11105 9755 11335 9850
rect 11455 9755 11685 9850
rect 11805 9755 12035 9850
rect 11195 9635 11245 9755
rect 10405 9550 10635 9635
rect 10755 9550 10985 9635
rect 11105 9550 11335 9635
rect 11455 9550 11685 9635
rect 11805 9550 12035 9635
rect 10405 9500 12035 9550
rect 10405 9405 10635 9500
rect 10755 9405 10985 9500
rect 11105 9405 11335 9500
rect 11455 9405 11685 9500
rect 11805 9405 12035 9500
rect 11195 9285 11245 9405
rect 10405 9200 10635 9285
rect 10755 9200 10985 9285
rect 11105 9200 11335 9285
rect 11455 9200 11685 9285
rect 11805 9200 12035 9285
rect 10405 9150 12035 9200
rect 10405 9055 10635 9150
rect 10755 9055 10985 9150
rect 11105 9055 11335 9150
rect 11455 9055 11685 9150
rect 11805 9055 12035 9150
rect 11195 8935 11245 9055
rect 10405 8850 10635 8935
rect 10755 8850 10985 8935
rect 11105 8850 11335 8935
rect 11455 8850 11685 8935
rect 11805 8850 12035 8935
rect 10405 8800 12035 8850
rect 10405 8705 10635 8800
rect 10755 8705 10985 8800
rect 11105 8705 11335 8800
rect 11455 8705 11685 8800
rect 11805 8705 12035 8800
rect 11195 8585 11245 8705
rect 10405 8500 10635 8585
rect 10755 8500 10985 8585
rect 11105 8500 11335 8585
rect 11455 8500 11685 8585
rect 11805 8500 12035 8585
rect 10405 8450 12035 8500
rect 10405 8355 10635 8450
rect 10755 8355 10985 8450
rect 11105 8355 11335 8450
rect 11455 8355 11685 8450
rect 11805 8355 12035 8450
rect 11195 8235 11245 8355
rect 10405 8150 10635 8235
rect 10755 8150 10985 8235
rect 11105 8150 11335 8235
rect 11455 8150 11685 8235
rect 11805 8150 12035 8235
rect 10405 8100 12035 8150
rect 10405 8005 10635 8100
rect 10755 8005 10985 8100
rect 11105 8005 11335 8100
rect 11455 8005 11685 8100
rect 11805 8005 12035 8100
rect 11195 7885 11245 8005
rect 10405 7800 10635 7885
rect 10755 7800 10985 7885
rect 11105 7800 11335 7885
rect 11455 7800 11685 7885
rect 11805 7800 12035 7885
rect 10405 7750 12035 7800
rect 10405 7655 10635 7750
rect 10755 7655 10985 7750
rect 11105 7655 11335 7750
rect 11455 7655 11685 7750
rect 11805 7655 12035 7750
rect 11195 7535 11245 7655
rect 10405 7450 10635 7535
rect 10755 7450 10985 7535
rect 11105 7450 11335 7535
rect 11455 7450 11685 7535
rect 11805 7450 12035 7535
rect 10405 7400 12035 7450
rect 10405 7305 10635 7400
rect 10755 7305 10985 7400
rect 11105 7305 11335 7400
rect 11455 7305 11685 7400
rect 11805 7305 12035 7400
rect 11195 7185 11245 7305
rect 10405 7100 10635 7185
rect 10755 7100 10985 7185
rect 11105 7100 11335 7185
rect 11455 7100 11685 7185
rect 11805 7100 12035 7185
rect 10405 7050 12035 7100
rect 10405 6955 10635 7050
rect 10755 6955 10985 7050
rect 11105 6955 11335 7050
rect 11455 6955 11685 7050
rect 11805 6955 12035 7050
rect 11195 6835 11245 6955
rect 10405 6750 10635 6835
rect 10755 6750 10985 6835
rect 11105 6750 11335 6835
rect 11455 6750 11685 6835
rect 11805 6750 12035 6835
rect 10405 6700 12035 6750
rect 10405 6605 10635 6700
rect 10755 6605 10985 6700
rect 11105 6605 11335 6700
rect 11455 6605 11685 6700
rect 11805 6605 12035 6700
rect 11195 6485 11245 6605
rect 10405 6400 10635 6485
rect 10755 6400 10985 6485
rect 11105 6400 11335 6485
rect 11455 6400 11685 6485
rect 11805 6400 12035 6485
rect 10405 6350 12035 6400
rect 10405 6255 10635 6350
rect 10755 6255 10985 6350
rect 11105 6255 11335 6350
rect 11455 6255 11685 6350
rect 11805 6255 12035 6350
rect 11195 6135 11245 6255
rect 10405 6050 10635 6135
rect 10755 6050 10985 6135
rect 11105 6050 11335 6135
rect 11455 6050 11685 6135
rect 11805 6050 12035 6135
rect 10405 6000 12035 6050
rect 10405 5905 10635 6000
rect 10755 5905 10985 6000
rect 11105 5905 11335 6000
rect 11455 5905 11685 6000
rect 11805 5905 12035 6000
rect 11195 5785 11245 5905
rect 10405 5700 10635 5785
rect 10755 5700 10985 5785
rect 11105 5700 11335 5785
rect 11455 5700 11685 5785
rect 11805 5700 12035 5785
rect 10405 5650 12035 5700
rect 10405 5555 10635 5650
rect 10755 5555 10985 5650
rect 11105 5555 11335 5650
rect 11455 5555 11685 5650
rect 11805 5555 12035 5650
rect 11195 5435 11245 5555
rect 10405 5350 10635 5435
rect 10755 5350 10985 5435
rect 11105 5350 11335 5435
rect 11455 5350 11685 5435
rect 11805 5350 12035 5435
rect 10405 5300 12035 5350
rect 10405 5205 10635 5300
rect 10755 5205 10985 5300
rect 11105 5205 11335 5300
rect 11455 5205 11685 5300
rect 11805 5205 12035 5300
rect 11195 5085 11245 5205
rect 10405 5000 10635 5085
rect 10755 5000 10985 5085
rect 11105 5000 11335 5085
rect 11455 5000 11685 5085
rect 11805 5000 12035 5085
rect 10405 4950 12035 5000
rect 10405 4855 10635 4950
rect 10755 4855 10985 4950
rect 11105 4855 11335 4950
rect 11455 4855 11685 4950
rect 11805 4855 12035 4950
rect 11195 4735 11245 4855
rect 10405 4650 10635 4735
rect 10755 4650 10985 4735
rect 11105 4650 11335 4735
rect 11455 4650 11685 4735
rect 11805 4650 12035 4735
rect 10405 4600 12035 4650
rect 10405 4505 10635 4600
rect 10755 4505 10985 4600
rect 11105 4505 11335 4600
rect 11455 4505 11685 4600
rect 11805 4505 12035 4600
rect 11195 4385 11245 4505
rect 10405 4300 10635 4385
rect 10755 4300 10985 4385
rect 11105 4300 11335 4385
rect 11455 4300 11685 4385
rect 11805 4300 12035 4385
rect 10405 4250 12035 4300
rect 10405 4155 10635 4250
rect 10755 4155 10985 4250
rect 11105 4155 11335 4250
rect 11455 4155 11685 4250
rect 11805 4155 12035 4250
rect 11195 4035 11245 4155
rect 10405 3950 10635 4035
rect 10755 3950 10985 4035
rect 11105 3950 11335 4035
rect 11455 3950 11685 4035
rect 11805 3950 12035 4035
rect 10405 3900 12035 3950
rect 10405 3805 10635 3900
rect 10755 3805 10985 3900
rect 11105 3805 11335 3900
rect 11455 3805 11685 3900
rect 11805 3805 12035 3900
rect 11195 3685 11245 3805
rect 10405 3600 10635 3685
rect 10755 3600 10985 3685
rect 11105 3600 11335 3685
rect 11455 3600 11685 3685
rect 11805 3600 12035 3685
rect 10405 3550 12035 3600
rect 10405 3455 10635 3550
rect 10755 3455 10985 3550
rect 11105 3455 11335 3550
rect 11455 3455 11685 3550
rect 11805 3455 12035 3550
rect 11195 3335 11245 3455
rect 10405 3250 10635 3335
rect 10755 3250 10985 3335
rect 11105 3250 11335 3335
rect 11455 3250 11685 3335
rect 11805 3250 12035 3335
rect 10405 3200 12035 3250
rect 10405 3105 10635 3200
rect 10755 3105 10985 3200
rect 11105 3105 11335 3200
rect 11455 3105 11685 3200
rect 11805 3105 12035 3200
rect 11195 2985 11245 3105
rect 10405 2900 10635 2985
rect 10755 2900 10985 2985
rect 11105 2900 11335 2985
rect 11455 2900 11685 2985
rect 11805 2900 12035 2985
rect 10405 2850 12035 2900
rect 10405 2755 10635 2850
rect 10755 2755 10985 2850
rect 11105 2755 11335 2850
rect 11455 2755 11685 2850
rect 11805 2755 12035 2850
rect 11195 2635 11245 2755
rect 10405 2550 10635 2635
rect 10755 2550 10985 2635
rect 11105 2550 11335 2635
rect 11455 2550 11685 2635
rect 11805 2550 12035 2635
rect 10405 2500 12035 2550
rect 10405 2405 10635 2500
rect 10755 2405 10985 2500
rect 11105 2405 11335 2500
rect 11455 2405 11685 2500
rect 11805 2405 12035 2500
rect 11195 2285 11245 2405
rect 10405 2200 10635 2285
rect 10755 2200 10985 2285
rect 11105 2200 11335 2285
rect 11455 2200 11685 2285
rect 11805 2200 12035 2285
rect 10405 2150 12035 2200
rect 10405 2055 10635 2150
rect 10755 2055 10985 2150
rect 11105 2055 11335 2150
rect 11455 2055 11685 2150
rect 11805 2055 12035 2150
rect 11195 1935 11245 2055
rect 10405 1850 10635 1935
rect 10755 1850 10985 1935
rect 11105 1850 11335 1935
rect 11455 1850 11685 1935
rect 11805 1850 12035 1935
rect 10405 1800 12035 1850
rect 10405 1705 10635 1800
rect 10755 1705 10985 1800
rect 11105 1705 11335 1800
rect 11455 1705 11685 1800
rect 11805 1705 12035 1800
rect 11195 1585 11245 1705
rect 10405 1500 10635 1585
rect 10755 1500 10985 1585
rect 11105 1500 11335 1585
rect 11455 1500 11685 1585
rect 11805 1500 12035 1585
rect 10405 1450 12035 1500
rect 10405 1355 10635 1450
rect 10755 1355 10985 1450
rect 11105 1355 11335 1450
rect 11455 1355 11685 1450
rect 11805 1355 12035 1450
rect 11195 1235 11245 1355
rect 10405 1150 10635 1235
rect 10755 1150 10985 1235
rect 11105 1150 11335 1235
rect 11455 1150 11685 1235
rect 11805 1150 12035 1235
rect 10405 1100 12035 1150
rect 10405 1005 10635 1100
rect 10755 1005 10985 1100
rect 11105 1005 11335 1100
rect 11455 1005 11685 1100
rect 11805 1005 12035 1100
rect 11195 885 11245 1005
rect 10405 800 10635 885
rect 10755 800 10985 885
rect 11105 800 11335 885
rect 11455 800 11685 885
rect 11805 800 12035 885
rect 10405 750 12035 800
rect 10405 655 10635 750
rect 10755 655 10985 750
rect 11105 655 11335 750
rect 11455 655 11685 750
rect 11805 655 12035 750
rect 11195 535 11245 655
rect 10405 450 10635 535
rect 10755 450 10985 535
rect 11105 450 11335 535
rect 11455 450 11685 535
rect 11805 450 12035 535
rect 10405 400 12035 450
rect 10405 305 10635 400
rect 10755 305 10985 400
rect 11105 305 11335 400
rect 11455 305 11685 400
rect 11805 305 12035 400
rect 10185 45 10235 50
rect 10185 5 10190 45
rect 10230 5 10235 45
rect 10185 0 10235 5
<< via3 >>
rect 10190 14420 10230 14460
rect 10190 5 10230 45
<< mimcap >>
rect 10420 14095 10620 14170
rect 10420 14055 10500 14095
rect 10540 14055 10620 14095
rect 10420 13970 10620 14055
rect 10770 14095 10970 14170
rect 10770 14055 10850 14095
rect 10890 14055 10970 14095
rect 10770 13970 10970 14055
rect 11120 14095 11320 14170
rect 11120 14055 11200 14095
rect 11240 14055 11320 14095
rect 11120 13970 11320 14055
rect 11470 14095 11670 14170
rect 11470 14055 11550 14095
rect 11590 14055 11670 14095
rect 11470 13970 11670 14055
rect 11820 14095 12020 14170
rect 11820 14055 11900 14095
rect 11940 14055 12020 14095
rect 11820 13970 12020 14055
rect 10420 13745 10620 13820
rect 10420 13705 10500 13745
rect 10540 13705 10620 13745
rect 10420 13620 10620 13705
rect 10770 13745 10970 13820
rect 10770 13705 10850 13745
rect 10890 13705 10970 13745
rect 10770 13620 10970 13705
rect 11120 13745 11320 13820
rect 11120 13705 11200 13745
rect 11240 13705 11320 13745
rect 11120 13620 11320 13705
rect 11470 13745 11670 13820
rect 11470 13705 11550 13745
rect 11590 13705 11670 13745
rect 11470 13620 11670 13705
rect 11820 13745 12020 13820
rect 11820 13705 11900 13745
rect 11940 13705 12020 13745
rect 11820 13620 12020 13705
rect 10420 13395 10620 13470
rect 10420 13355 10500 13395
rect 10540 13355 10620 13395
rect 10420 13270 10620 13355
rect 10770 13395 10970 13470
rect 10770 13355 10850 13395
rect 10890 13355 10970 13395
rect 10770 13270 10970 13355
rect 11120 13395 11320 13470
rect 11120 13355 11200 13395
rect 11240 13355 11320 13395
rect 11120 13270 11320 13355
rect 11470 13395 11670 13470
rect 11470 13355 11550 13395
rect 11590 13355 11670 13395
rect 11470 13270 11670 13355
rect 11820 13395 12020 13470
rect 11820 13355 11900 13395
rect 11940 13355 12020 13395
rect 11820 13270 12020 13355
rect 10420 13045 10620 13120
rect 10420 13005 10500 13045
rect 10540 13005 10620 13045
rect 10420 12920 10620 13005
rect 10770 13045 10970 13120
rect 10770 13005 10850 13045
rect 10890 13005 10970 13045
rect 10770 12920 10970 13005
rect 11120 13045 11320 13120
rect 11120 13005 11200 13045
rect 11240 13005 11320 13045
rect 11120 12920 11320 13005
rect 11470 13045 11670 13120
rect 11470 13005 11550 13045
rect 11590 13005 11670 13045
rect 11470 12920 11670 13005
rect 11820 13045 12020 13120
rect 11820 13005 11900 13045
rect 11940 13005 12020 13045
rect 11820 12920 12020 13005
rect 10420 12695 10620 12770
rect 10420 12655 10500 12695
rect 10540 12655 10620 12695
rect 10420 12570 10620 12655
rect 10770 12695 10970 12770
rect 10770 12655 10850 12695
rect 10890 12655 10970 12695
rect 10770 12570 10970 12655
rect 11120 12695 11320 12770
rect 11120 12655 11200 12695
rect 11240 12655 11320 12695
rect 11120 12570 11320 12655
rect 11470 12695 11670 12770
rect 11470 12655 11550 12695
rect 11590 12655 11670 12695
rect 11470 12570 11670 12655
rect 11820 12695 12020 12770
rect 11820 12655 11900 12695
rect 11940 12655 12020 12695
rect 11820 12570 12020 12655
rect 10420 12345 10620 12420
rect 10420 12305 10500 12345
rect 10540 12305 10620 12345
rect 10420 12220 10620 12305
rect 10770 12345 10970 12420
rect 10770 12305 10850 12345
rect 10890 12305 10970 12345
rect 10770 12220 10970 12305
rect 11120 12345 11320 12420
rect 11120 12305 11200 12345
rect 11240 12305 11320 12345
rect 11120 12220 11320 12305
rect 11470 12345 11670 12420
rect 11470 12305 11550 12345
rect 11590 12305 11670 12345
rect 11470 12220 11670 12305
rect 11820 12345 12020 12420
rect 11820 12305 11900 12345
rect 11940 12305 12020 12345
rect 11820 12220 12020 12305
rect 10420 11995 10620 12070
rect 10420 11955 10500 11995
rect 10540 11955 10620 11995
rect 10420 11870 10620 11955
rect 10770 11995 10970 12070
rect 10770 11955 10850 11995
rect 10890 11955 10970 11995
rect 10770 11870 10970 11955
rect 11120 11995 11320 12070
rect 11120 11955 11200 11995
rect 11240 11955 11320 11995
rect 11120 11870 11320 11955
rect 11470 11995 11670 12070
rect 11470 11955 11550 11995
rect 11590 11955 11670 11995
rect 11470 11870 11670 11955
rect 11820 11995 12020 12070
rect 11820 11955 11900 11995
rect 11940 11955 12020 11995
rect 11820 11870 12020 11955
rect 10420 11645 10620 11720
rect 10420 11605 10500 11645
rect 10540 11605 10620 11645
rect 10420 11520 10620 11605
rect 10770 11645 10970 11720
rect 10770 11605 10850 11645
rect 10890 11605 10970 11645
rect 10770 11520 10970 11605
rect 11120 11645 11320 11720
rect 11120 11605 11200 11645
rect 11240 11605 11320 11645
rect 11120 11520 11320 11605
rect 11470 11645 11670 11720
rect 11470 11605 11550 11645
rect 11590 11605 11670 11645
rect 11470 11520 11670 11605
rect 11820 11645 12020 11720
rect 11820 11605 11900 11645
rect 11940 11605 12020 11645
rect 11820 11520 12020 11605
rect 10420 11295 10620 11370
rect 10420 11255 10500 11295
rect 10540 11255 10620 11295
rect 10420 11170 10620 11255
rect 10770 11295 10970 11370
rect 10770 11255 10850 11295
rect 10890 11255 10970 11295
rect 10770 11170 10970 11255
rect 11120 11295 11320 11370
rect 11120 11255 11200 11295
rect 11240 11255 11320 11295
rect 11120 11170 11320 11255
rect 11470 11295 11670 11370
rect 11470 11255 11550 11295
rect 11590 11255 11670 11295
rect 11470 11170 11670 11255
rect 11820 11295 12020 11370
rect 11820 11255 11900 11295
rect 11940 11255 12020 11295
rect 11820 11170 12020 11255
rect 10420 10945 10620 11020
rect 10420 10905 10500 10945
rect 10540 10905 10620 10945
rect 10420 10820 10620 10905
rect 10770 10945 10970 11020
rect 10770 10905 10850 10945
rect 10890 10905 10970 10945
rect 10770 10820 10970 10905
rect 11120 10945 11320 11020
rect 11120 10905 11200 10945
rect 11240 10905 11320 10945
rect 11120 10820 11320 10905
rect 11470 10945 11670 11020
rect 11470 10905 11550 10945
rect 11590 10905 11670 10945
rect 11470 10820 11670 10905
rect 11820 10945 12020 11020
rect 11820 10905 11900 10945
rect 11940 10905 12020 10945
rect 11820 10820 12020 10905
rect 10420 10595 10620 10670
rect 10420 10555 10500 10595
rect 10540 10555 10620 10595
rect 10420 10470 10620 10555
rect 10770 10595 10970 10670
rect 10770 10555 10850 10595
rect 10890 10555 10970 10595
rect 10770 10470 10970 10555
rect 11120 10595 11320 10670
rect 11120 10555 11200 10595
rect 11240 10555 11320 10595
rect 11120 10470 11320 10555
rect 11470 10595 11670 10670
rect 11470 10555 11550 10595
rect 11590 10555 11670 10595
rect 11470 10470 11670 10555
rect 11820 10595 12020 10670
rect 11820 10555 11900 10595
rect 11940 10555 12020 10595
rect 11820 10470 12020 10555
rect 10420 10245 10620 10320
rect 10420 10205 10500 10245
rect 10540 10205 10620 10245
rect 10420 10120 10620 10205
rect 10770 10245 10970 10320
rect 10770 10205 10850 10245
rect 10890 10205 10970 10245
rect 10770 10120 10970 10205
rect 11120 10245 11320 10320
rect 11120 10205 11200 10245
rect 11240 10205 11320 10245
rect 11120 10120 11320 10205
rect 11470 10245 11670 10320
rect 11470 10205 11550 10245
rect 11590 10205 11670 10245
rect 11470 10120 11670 10205
rect 11820 10245 12020 10320
rect 11820 10205 11900 10245
rect 11940 10205 12020 10245
rect 11820 10120 12020 10205
rect 10420 9895 10620 9970
rect 10420 9855 10500 9895
rect 10540 9855 10620 9895
rect 10420 9770 10620 9855
rect 10770 9895 10970 9970
rect 10770 9855 10850 9895
rect 10890 9855 10970 9895
rect 10770 9770 10970 9855
rect 11120 9895 11320 9970
rect 11120 9855 11200 9895
rect 11240 9855 11320 9895
rect 11120 9770 11320 9855
rect 11470 9895 11670 9970
rect 11470 9855 11550 9895
rect 11590 9855 11670 9895
rect 11470 9770 11670 9855
rect 11820 9895 12020 9970
rect 11820 9855 11900 9895
rect 11940 9855 12020 9895
rect 11820 9770 12020 9855
rect 10420 9545 10620 9620
rect 10420 9505 10500 9545
rect 10540 9505 10620 9545
rect 10420 9420 10620 9505
rect 10770 9545 10970 9620
rect 10770 9505 10850 9545
rect 10890 9505 10970 9545
rect 10770 9420 10970 9505
rect 11120 9545 11320 9620
rect 11120 9505 11200 9545
rect 11240 9505 11320 9545
rect 11120 9420 11320 9505
rect 11470 9545 11670 9620
rect 11470 9505 11550 9545
rect 11590 9505 11670 9545
rect 11470 9420 11670 9505
rect 11820 9545 12020 9620
rect 11820 9505 11900 9545
rect 11940 9505 12020 9545
rect 11820 9420 12020 9505
rect 10420 9195 10620 9270
rect 10420 9155 10500 9195
rect 10540 9155 10620 9195
rect 10420 9070 10620 9155
rect 10770 9195 10970 9270
rect 10770 9155 10850 9195
rect 10890 9155 10970 9195
rect 10770 9070 10970 9155
rect 11120 9195 11320 9270
rect 11120 9155 11200 9195
rect 11240 9155 11320 9195
rect 11120 9070 11320 9155
rect 11470 9195 11670 9270
rect 11470 9155 11550 9195
rect 11590 9155 11670 9195
rect 11470 9070 11670 9155
rect 11820 9195 12020 9270
rect 11820 9155 11900 9195
rect 11940 9155 12020 9195
rect 11820 9070 12020 9155
rect 10420 8845 10620 8920
rect 10420 8805 10500 8845
rect 10540 8805 10620 8845
rect 10420 8720 10620 8805
rect 10770 8845 10970 8920
rect 10770 8805 10850 8845
rect 10890 8805 10970 8845
rect 10770 8720 10970 8805
rect 11120 8845 11320 8920
rect 11120 8805 11200 8845
rect 11240 8805 11320 8845
rect 11120 8720 11320 8805
rect 11470 8845 11670 8920
rect 11470 8805 11550 8845
rect 11590 8805 11670 8845
rect 11470 8720 11670 8805
rect 11820 8845 12020 8920
rect 11820 8805 11900 8845
rect 11940 8805 12020 8845
rect 11820 8720 12020 8805
rect 10420 8495 10620 8570
rect 10420 8455 10500 8495
rect 10540 8455 10620 8495
rect 10420 8370 10620 8455
rect 10770 8495 10970 8570
rect 10770 8455 10850 8495
rect 10890 8455 10970 8495
rect 10770 8370 10970 8455
rect 11120 8495 11320 8570
rect 11120 8455 11200 8495
rect 11240 8455 11320 8495
rect 11120 8370 11320 8455
rect 11470 8495 11670 8570
rect 11470 8455 11550 8495
rect 11590 8455 11670 8495
rect 11470 8370 11670 8455
rect 11820 8495 12020 8570
rect 11820 8455 11900 8495
rect 11940 8455 12020 8495
rect 11820 8370 12020 8455
rect 10420 8145 10620 8220
rect 10420 8105 10500 8145
rect 10540 8105 10620 8145
rect 10420 8020 10620 8105
rect 10770 8145 10970 8220
rect 10770 8105 10850 8145
rect 10890 8105 10970 8145
rect 10770 8020 10970 8105
rect 11120 8145 11320 8220
rect 11120 8105 11200 8145
rect 11240 8105 11320 8145
rect 11120 8020 11320 8105
rect 11470 8145 11670 8220
rect 11470 8105 11550 8145
rect 11590 8105 11670 8145
rect 11470 8020 11670 8105
rect 11820 8145 12020 8220
rect 11820 8105 11900 8145
rect 11940 8105 12020 8145
rect 11820 8020 12020 8105
rect 10420 7795 10620 7870
rect 10420 7755 10500 7795
rect 10540 7755 10620 7795
rect 10420 7670 10620 7755
rect 10770 7795 10970 7870
rect 10770 7755 10850 7795
rect 10890 7755 10970 7795
rect 10770 7670 10970 7755
rect 11120 7795 11320 7870
rect 11120 7755 11200 7795
rect 11240 7755 11320 7795
rect 11120 7670 11320 7755
rect 11470 7795 11670 7870
rect 11470 7755 11550 7795
rect 11590 7755 11670 7795
rect 11470 7670 11670 7755
rect 11820 7795 12020 7870
rect 11820 7755 11900 7795
rect 11940 7755 12020 7795
rect 11820 7670 12020 7755
rect 10420 7445 10620 7520
rect 10420 7405 10500 7445
rect 10540 7405 10620 7445
rect 10420 7320 10620 7405
rect 10770 7445 10970 7520
rect 10770 7405 10850 7445
rect 10890 7405 10970 7445
rect 10770 7320 10970 7405
rect 11120 7445 11320 7520
rect 11120 7405 11200 7445
rect 11240 7405 11320 7445
rect 11120 7320 11320 7405
rect 11470 7445 11670 7520
rect 11470 7405 11550 7445
rect 11590 7405 11670 7445
rect 11470 7320 11670 7405
rect 11820 7445 12020 7520
rect 11820 7405 11900 7445
rect 11940 7405 12020 7445
rect 11820 7320 12020 7405
rect 10420 7095 10620 7170
rect 10420 7055 10500 7095
rect 10540 7055 10620 7095
rect 10420 6970 10620 7055
rect 10770 7095 10970 7170
rect 10770 7055 10850 7095
rect 10890 7055 10970 7095
rect 10770 6970 10970 7055
rect 11120 7095 11320 7170
rect 11120 7055 11200 7095
rect 11240 7055 11320 7095
rect 11120 6970 11320 7055
rect 11470 7095 11670 7170
rect 11470 7055 11550 7095
rect 11590 7055 11670 7095
rect 11470 6970 11670 7055
rect 11820 7095 12020 7170
rect 11820 7055 11900 7095
rect 11940 7055 12020 7095
rect 11820 6970 12020 7055
rect 10420 6745 10620 6820
rect 10420 6705 10500 6745
rect 10540 6705 10620 6745
rect 10420 6620 10620 6705
rect 10770 6745 10970 6820
rect 10770 6705 10850 6745
rect 10890 6705 10970 6745
rect 10770 6620 10970 6705
rect 11120 6745 11320 6820
rect 11120 6705 11200 6745
rect 11240 6705 11320 6745
rect 11120 6620 11320 6705
rect 11470 6745 11670 6820
rect 11470 6705 11550 6745
rect 11590 6705 11670 6745
rect 11470 6620 11670 6705
rect 11820 6745 12020 6820
rect 11820 6705 11900 6745
rect 11940 6705 12020 6745
rect 11820 6620 12020 6705
rect 10420 6395 10620 6470
rect 10420 6355 10500 6395
rect 10540 6355 10620 6395
rect 10420 6270 10620 6355
rect 10770 6395 10970 6470
rect 10770 6355 10850 6395
rect 10890 6355 10970 6395
rect 10770 6270 10970 6355
rect 11120 6395 11320 6470
rect 11120 6355 11200 6395
rect 11240 6355 11320 6395
rect 11120 6270 11320 6355
rect 11470 6395 11670 6470
rect 11470 6355 11550 6395
rect 11590 6355 11670 6395
rect 11470 6270 11670 6355
rect 11820 6395 12020 6470
rect 11820 6355 11900 6395
rect 11940 6355 12020 6395
rect 11820 6270 12020 6355
rect 10420 6045 10620 6120
rect 10420 6005 10500 6045
rect 10540 6005 10620 6045
rect 10420 5920 10620 6005
rect 10770 6045 10970 6120
rect 10770 6005 10850 6045
rect 10890 6005 10970 6045
rect 10770 5920 10970 6005
rect 11120 6045 11320 6120
rect 11120 6005 11200 6045
rect 11240 6005 11320 6045
rect 11120 5920 11320 6005
rect 11470 6045 11670 6120
rect 11470 6005 11550 6045
rect 11590 6005 11670 6045
rect 11470 5920 11670 6005
rect 11820 6045 12020 6120
rect 11820 6005 11900 6045
rect 11940 6005 12020 6045
rect 11820 5920 12020 6005
rect 10420 5695 10620 5770
rect 10420 5655 10500 5695
rect 10540 5655 10620 5695
rect 10420 5570 10620 5655
rect 10770 5695 10970 5770
rect 10770 5655 10850 5695
rect 10890 5655 10970 5695
rect 10770 5570 10970 5655
rect 11120 5695 11320 5770
rect 11120 5655 11200 5695
rect 11240 5655 11320 5695
rect 11120 5570 11320 5655
rect 11470 5695 11670 5770
rect 11470 5655 11550 5695
rect 11590 5655 11670 5695
rect 11470 5570 11670 5655
rect 11820 5695 12020 5770
rect 11820 5655 11900 5695
rect 11940 5655 12020 5695
rect 11820 5570 12020 5655
rect 10420 5345 10620 5420
rect 10420 5305 10500 5345
rect 10540 5305 10620 5345
rect 10420 5220 10620 5305
rect 10770 5345 10970 5420
rect 10770 5305 10850 5345
rect 10890 5305 10970 5345
rect 10770 5220 10970 5305
rect 11120 5345 11320 5420
rect 11120 5305 11200 5345
rect 11240 5305 11320 5345
rect 11120 5220 11320 5305
rect 11470 5345 11670 5420
rect 11470 5305 11550 5345
rect 11590 5305 11670 5345
rect 11470 5220 11670 5305
rect 11820 5345 12020 5420
rect 11820 5305 11900 5345
rect 11940 5305 12020 5345
rect 11820 5220 12020 5305
rect 10420 4995 10620 5070
rect 10420 4955 10500 4995
rect 10540 4955 10620 4995
rect 10420 4870 10620 4955
rect 10770 4995 10970 5070
rect 10770 4955 10850 4995
rect 10890 4955 10970 4995
rect 10770 4870 10970 4955
rect 11120 4995 11320 5070
rect 11120 4955 11200 4995
rect 11240 4955 11320 4995
rect 11120 4870 11320 4955
rect 11470 4995 11670 5070
rect 11470 4955 11550 4995
rect 11590 4955 11670 4995
rect 11470 4870 11670 4955
rect 11820 4995 12020 5070
rect 11820 4955 11900 4995
rect 11940 4955 12020 4995
rect 11820 4870 12020 4955
rect 10420 4645 10620 4720
rect 10420 4605 10500 4645
rect 10540 4605 10620 4645
rect 10420 4520 10620 4605
rect 10770 4645 10970 4720
rect 10770 4605 10850 4645
rect 10890 4605 10970 4645
rect 10770 4520 10970 4605
rect 11120 4645 11320 4720
rect 11120 4605 11200 4645
rect 11240 4605 11320 4645
rect 11120 4520 11320 4605
rect 11470 4645 11670 4720
rect 11470 4605 11550 4645
rect 11590 4605 11670 4645
rect 11470 4520 11670 4605
rect 11820 4645 12020 4720
rect 11820 4605 11900 4645
rect 11940 4605 12020 4645
rect 11820 4520 12020 4605
rect 10420 4295 10620 4370
rect 10420 4255 10500 4295
rect 10540 4255 10620 4295
rect 10420 4170 10620 4255
rect 10770 4295 10970 4370
rect 10770 4255 10850 4295
rect 10890 4255 10970 4295
rect 10770 4170 10970 4255
rect 11120 4295 11320 4370
rect 11120 4255 11200 4295
rect 11240 4255 11320 4295
rect 11120 4170 11320 4255
rect 11470 4295 11670 4370
rect 11470 4255 11550 4295
rect 11590 4255 11670 4295
rect 11470 4170 11670 4255
rect 11820 4295 12020 4370
rect 11820 4255 11900 4295
rect 11940 4255 12020 4295
rect 11820 4170 12020 4255
rect 10420 3945 10620 4020
rect 10420 3905 10500 3945
rect 10540 3905 10620 3945
rect 10420 3820 10620 3905
rect 10770 3945 10970 4020
rect 10770 3905 10850 3945
rect 10890 3905 10970 3945
rect 10770 3820 10970 3905
rect 11120 3945 11320 4020
rect 11120 3905 11200 3945
rect 11240 3905 11320 3945
rect 11120 3820 11320 3905
rect 11470 3945 11670 4020
rect 11470 3905 11550 3945
rect 11590 3905 11670 3945
rect 11470 3820 11670 3905
rect 11820 3945 12020 4020
rect 11820 3905 11900 3945
rect 11940 3905 12020 3945
rect 11820 3820 12020 3905
rect 10420 3595 10620 3670
rect 10420 3555 10500 3595
rect 10540 3555 10620 3595
rect 10420 3470 10620 3555
rect 10770 3595 10970 3670
rect 10770 3555 10850 3595
rect 10890 3555 10970 3595
rect 10770 3470 10970 3555
rect 11120 3595 11320 3670
rect 11120 3555 11200 3595
rect 11240 3555 11320 3595
rect 11120 3470 11320 3555
rect 11470 3595 11670 3670
rect 11470 3555 11550 3595
rect 11590 3555 11670 3595
rect 11470 3470 11670 3555
rect 11820 3595 12020 3670
rect 11820 3555 11900 3595
rect 11940 3555 12020 3595
rect 11820 3470 12020 3555
rect 10420 3245 10620 3320
rect 10420 3205 10500 3245
rect 10540 3205 10620 3245
rect 10420 3120 10620 3205
rect 10770 3245 10970 3320
rect 10770 3205 10850 3245
rect 10890 3205 10970 3245
rect 10770 3120 10970 3205
rect 11120 3245 11320 3320
rect 11120 3205 11200 3245
rect 11240 3205 11320 3245
rect 11120 3120 11320 3205
rect 11470 3245 11670 3320
rect 11470 3205 11550 3245
rect 11590 3205 11670 3245
rect 11470 3120 11670 3205
rect 11820 3245 12020 3320
rect 11820 3205 11900 3245
rect 11940 3205 12020 3245
rect 11820 3120 12020 3205
rect 10420 2895 10620 2970
rect 10420 2855 10500 2895
rect 10540 2855 10620 2895
rect 10420 2770 10620 2855
rect 10770 2895 10970 2970
rect 10770 2855 10850 2895
rect 10890 2855 10970 2895
rect 10770 2770 10970 2855
rect 11120 2895 11320 2970
rect 11120 2855 11200 2895
rect 11240 2855 11320 2895
rect 11120 2770 11320 2855
rect 11470 2895 11670 2970
rect 11470 2855 11550 2895
rect 11590 2855 11670 2895
rect 11470 2770 11670 2855
rect 11820 2895 12020 2970
rect 11820 2855 11900 2895
rect 11940 2855 12020 2895
rect 11820 2770 12020 2855
rect 10420 2545 10620 2620
rect 10420 2505 10500 2545
rect 10540 2505 10620 2545
rect 10420 2420 10620 2505
rect 10770 2545 10970 2620
rect 10770 2505 10850 2545
rect 10890 2505 10970 2545
rect 10770 2420 10970 2505
rect 11120 2545 11320 2620
rect 11120 2505 11200 2545
rect 11240 2505 11320 2545
rect 11120 2420 11320 2505
rect 11470 2545 11670 2620
rect 11470 2505 11550 2545
rect 11590 2505 11670 2545
rect 11470 2420 11670 2505
rect 11820 2545 12020 2620
rect 11820 2505 11900 2545
rect 11940 2505 12020 2545
rect 11820 2420 12020 2505
rect 10420 2195 10620 2270
rect 10420 2155 10500 2195
rect 10540 2155 10620 2195
rect 10420 2070 10620 2155
rect 10770 2195 10970 2270
rect 10770 2155 10850 2195
rect 10890 2155 10970 2195
rect 10770 2070 10970 2155
rect 11120 2195 11320 2270
rect 11120 2155 11200 2195
rect 11240 2155 11320 2195
rect 11120 2070 11320 2155
rect 11470 2195 11670 2270
rect 11470 2155 11550 2195
rect 11590 2155 11670 2195
rect 11470 2070 11670 2155
rect 11820 2195 12020 2270
rect 11820 2155 11900 2195
rect 11940 2155 12020 2195
rect 11820 2070 12020 2155
rect 10420 1845 10620 1920
rect 10420 1805 10500 1845
rect 10540 1805 10620 1845
rect 10420 1720 10620 1805
rect 10770 1845 10970 1920
rect 10770 1805 10850 1845
rect 10890 1805 10970 1845
rect 10770 1720 10970 1805
rect 11120 1845 11320 1920
rect 11120 1805 11200 1845
rect 11240 1805 11320 1845
rect 11120 1720 11320 1805
rect 11470 1845 11670 1920
rect 11470 1805 11550 1845
rect 11590 1805 11670 1845
rect 11470 1720 11670 1805
rect 11820 1845 12020 1920
rect 11820 1805 11900 1845
rect 11940 1805 12020 1845
rect 11820 1720 12020 1805
rect 10420 1495 10620 1570
rect 10420 1455 10500 1495
rect 10540 1455 10620 1495
rect 10420 1370 10620 1455
rect 10770 1495 10970 1570
rect 10770 1455 10850 1495
rect 10890 1455 10970 1495
rect 10770 1370 10970 1455
rect 11120 1495 11320 1570
rect 11120 1455 11200 1495
rect 11240 1455 11320 1495
rect 11120 1370 11320 1455
rect 11470 1495 11670 1570
rect 11470 1455 11550 1495
rect 11590 1455 11670 1495
rect 11470 1370 11670 1455
rect 11820 1495 12020 1570
rect 11820 1455 11900 1495
rect 11940 1455 12020 1495
rect 11820 1370 12020 1455
rect 10420 1145 10620 1220
rect 10420 1105 10500 1145
rect 10540 1105 10620 1145
rect 10420 1020 10620 1105
rect 10770 1145 10970 1220
rect 10770 1105 10850 1145
rect 10890 1105 10970 1145
rect 10770 1020 10970 1105
rect 11120 1145 11320 1220
rect 11120 1105 11200 1145
rect 11240 1105 11320 1145
rect 11120 1020 11320 1105
rect 11470 1145 11670 1220
rect 11470 1105 11550 1145
rect 11590 1105 11670 1145
rect 11470 1020 11670 1105
rect 11820 1145 12020 1220
rect 11820 1105 11900 1145
rect 11940 1105 12020 1145
rect 11820 1020 12020 1105
rect 10420 795 10620 870
rect 10420 755 10500 795
rect 10540 755 10620 795
rect 10420 670 10620 755
rect 10770 795 10970 870
rect 10770 755 10850 795
rect 10890 755 10970 795
rect 10770 670 10970 755
rect 11120 795 11320 870
rect 11120 755 11200 795
rect 11240 755 11320 795
rect 11120 670 11320 755
rect 11470 795 11670 870
rect 11470 755 11550 795
rect 11590 755 11670 795
rect 11470 670 11670 755
rect 11820 795 12020 870
rect 11820 755 11900 795
rect 11940 755 12020 795
rect 11820 670 12020 755
rect 10420 445 10620 520
rect 10420 405 10500 445
rect 10540 405 10620 445
rect 10420 320 10620 405
rect 10770 445 10970 520
rect 10770 405 10850 445
rect 10890 405 10970 445
rect 10770 320 10970 405
rect 11120 445 11320 520
rect 11120 405 11200 445
rect 11240 405 11320 445
rect 11120 320 11320 405
rect 11470 445 11670 520
rect 11470 405 11550 445
rect 11590 405 11670 445
rect 11470 320 11670 405
rect 11820 445 12020 520
rect 11820 405 11900 445
rect 11940 405 12020 445
rect 11820 320 12020 405
<< mimcapcontact >>
rect 10500 14055 10540 14095
rect 10850 14055 10890 14095
rect 11200 14055 11240 14095
rect 11550 14055 11590 14095
rect 11900 14055 11940 14095
rect 10500 13705 10540 13745
rect 10850 13705 10890 13745
rect 11200 13705 11240 13745
rect 11550 13705 11590 13745
rect 11900 13705 11940 13745
rect 10500 13355 10540 13395
rect 10850 13355 10890 13395
rect 11200 13355 11240 13395
rect 11550 13355 11590 13395
rect 11900 13355 11940 13395
rect 10500 13005 10540 13045
rect 10850 13005 10890 13045
rect 11200 13005 11240 13045
rect 11550 13005 11590 13045
rect 11900 13005 11940 13045
rect 10500 12655 10540 12695
rect 10850 12655 10890 12695
rect 11200 12655 11240 12695
rect 11550 12655 11590 12695
rect 11900 12655 11940 12695
rect 10500 12305 10540 12345
rect 10850 12305 10890 12345
rect 11200 12305 11240 12345
rect 11550 12305 11590 12345
rect 11900 12305 11940 12345
rect 10500 11955 10540 11995
rect 10850 11955 10890 11995
rect 11200 11955 11240 11995
rect 11550 11955 11590 11995
rect 11900 11955 11940 11995
rect 10500 11605 10540 11645
rect 10850 11605 10890 11645
rect 11200 11605 11240 11645
rect 11550 11605 11590 11645
rect 11900 11605 11940 11645
rect 10500 11255 10540 11295
rect 10850 11255 10890 11295
rect 11200 11255 11240 11295
rect 11550 11255 11590 11295
rect 11900 11255 11940 11295
rect 10500 10905 10540 10945
rect 10850 10905 10890 10945
rect 11200 10905 11240 10945
rect 11550 10905 11590 10945
rect 11900 10905 11940 10945
rect 10500 10555 10540 10595
rect 10850 10555 10890 10595
rect 11200 10555 11240 10595
rect 11550 10555 11590 10595
rect 11900 10555 11940 10595
rect 10500 10205 10540 10245
rect 10850 10205 10890 10245
rect 11200 10205 11240 10245
rect 11550 10205 11590 10245
rect 11900 10205 11940 10245
rect 10500 9855 10540 9895
rect 10850 9855 10890 9895
rect 11200 9855 11240 9895
rect 11550 9855 11590 9895
rect 11900 9855 11940 9895
rect 10500 9505 10540 9545
rect 10850 9505 10890 9545
rect 11200 9505 11240 9545
rect 11550 9505 11590 9545
rect 11900 9505 11940 9545
rect 10500 9155 10540 9195
rect 10850 9155 10890 9195
rect 11200 9155 11240 9195
rect 11550 9155 11590 9195
rect 11900 9155 11940 9195
rect 10500 8805 10540 8845
rect 10850 8805 10890 8845
rect 11200 8805 11240 8845
rect 11550 8805 11590 8845
rect 11900 8805 11940 8845
rect 10500 8455 10540 8495
rect 10850 8455 10890 8495
rect 11200 8455 11240 8495
rect 11550 8455 11590 8495
rect 11900 8455 11940 8495
rect 10500 8105 10540 8145
rect 10850 8105 10890 8145
rect 11200 8105 11240 8145
rect 11550 8105 11590 8145
rect 11900 8105 11940 8145
rect 10500 7755 10540 7795
rect 10850 7755 10890 7795
rect 11200 7755 11240 7795
rect 11550 7755 11590 7795
rect 11900 7755 11940 7795
rect 10500 7405 10540 7445
rect 10850 7405 10890 7445
rect 11200 7405 11240 7445
rect 11550 7405 11590 7445
rect 11900 7405 11940 7445
rect 10500 7055 10540 7095
rect 10850 7055 10890 7095
rect 11200 7055 11240 7095
rect 11550 7055 11590 7095
rect 11900 7055 11940 7095
rect 10500 6705 10540 6745
rect 10850 6705 10890 6745
rect 11200 6705 11240 6745
rect 11550 6705 11590 6745
rect 11900 6705 11940 6745
rect 10500 6355 10540 6395
rect 10850 6355 10890 6395
rect 11200 6355 11240 6395
rect 11550 6355 11590 6395
rect 11900 6355 11940 6395
rect 10500 6005 10540 6045
rect 10850 6005 10890 6045
rect 11200 6005 11240 6045
rect 11550 6005 11590 6045
rect 11900 6005 11940 6045
rect 10500 5655 10540 5695
rect 10850 5655 10890 5695
rect 11200 5655 11240 5695
rect 11550 5655 11590 5695
rect 11900 5655 11940 5695
rect 10500 5305 10540 5345
rect 10850 5305 10890 5345
rect 11200 5305 11240 5345
rect 11550 5305 11590 5345
rect 11900 5305 11940 5345
rect 10500 4955 10540 4995
rect 10850 4955 10890 4995
rect 11200 4955 11240 4995
rect 11550 4955 11590 4995
rect 11900 4955 11940 4995
rect 10500 4605 10540 4645
rect 10850 4605 10890 4645
rect 11200 4605 11240 4645
rect 11550 4605 11590 4645
rect 11900 4605 11940 4645
rect 10500 4255 10540 4295
rect 10850 4255 10890 4295
rect 11200 4255 11240 4295
rect 11550 4255 11590 4295
rect 11900 4255 11940 4295
rect 10500 3905 10540 3945
rect 10850 3905 10890 3945
rect 11200 3905 11240 3945
rect 11550 3905 11590 3945
rect 11900 3905 11940 3945
rect 10500 3555 10540 3595
rect 10850 3555 10890 3595
rect 11200 3555 11240 3595
rect 11550 3555 11590 3595
rect 11900 3555 11940 3595
rect 10500 3205 10540 3245
rect 10850 3205 10890 3245
rect 11200 3205 11240 3245
rect 11550 3205 11590 3245
rect 11900 3205 11940 3245
rect 10500 2855 10540 2895
rect 10850 2855 10890 2895
rect 11200 2855 11240 2895
rect 11550 2855 11590 2895
rect 11900 2855 11940 2895
rect 10500 2505 10540 2545
rect 10850 2505 10890 2545
rect 11200 2505 11240 2545
rect 11550 2505 11590 2545
rect 11900 2505 11940 2545
rect 10500 2155 10540 2195
rect 10850 2155 10890 2195
rect 11200 2155 11240 2195
rect 11550 2155 11590 2195
rect 11900 2155 11940 2195
rect 10500 1805 10540 1845
rect 10850 1805 10890 1845
rect 11200 1805 11240 1845
rect 11550 1805 11590 1845
rect 11900 1805 11940 1845
rect 10500 1455 10540 1495
rect 10850 1455 10890 1495
rect 11200 1455 11240 1495
rect 11550 1455 11590 1495
rect 11900 1455 11940 1495
rect 10500 1105 10540 1145
rect 10850 1105 10890 1145
rect 11200 1105 11240 1145
rect 11550 1105 11590 1145
rect 11900 1105 11940 1145
rect 10500 755 10540 795
rect 10850 755 10890 795
rect 11200 755 11240 795
rect 11550 755 11590 795
rect 11900 755 11940 795
rect 10500 405 10540 445
rect 10850 405 10890 445
rect 11200 405 11240 445
rect 11550 405 11590 445
rect 11900 405 11940 445
<< metal4 >>
rect 7255 14460 10235 14465
rect 7255 14420 10190 14460
rect 10230 14420 10235 14460
rect 7255 14415 10235 14420
rect 10495 14095 11945 14100
rect 10495 14055 10500 14095
rect 10540 14055 10850 14095
rect 10890 14055 11200 14095
rect 11240 14055 11550 14095
rect 11590 14055 11900 14095
rect 11940 14055 11945 14095
rect 10495 14050 11945 14055
rect 11195 13750 11245 14050
rect 10495 13745 11945 13750
rect 10495 13705 10500 13745
rect 10540 13705 10850 13745
rect 10890 13705 11200 13745
rect 11240 13705 11550 13745
rect 11590 13705 11900 13745
rect 11940 13705 11945 13745
rect 10495 13700 11945 13705
rect 11195 13400 11245 13700
rect 10495 13395 11945 13400
rect 10495 13355 10500 13395
rect 10540 13355 10850 13395
rect 10890 13355 11200 13395
rect 11240 13355 11550 13395
rect 11590 13355 11900 13395
rect 11940 13355 11945 13395
rect 10495 13350 11945 13355
rect 11195 13050 11245 13350
rect 10495 13045 11945 13050
rect 10495 13005 10500 13045
rect 10540 13005 10850 13045
rect 10890 13005 11200 13045
rect 11240 13005 11550 13045
rect 11590 13005 11900 13045
rect 11940 13005 11945 13045
rect 10495 13000 11945 13005
rect 11195 12700 11245 13000
rect 10495 12695 11945 12700
rect 10495 12655 10500 12695
rect 10540 12655 10850 12695
rect 10890 12655 11200 12695
rect 11240 12655 11550 12695
rect 11590 12655 11900 12695
rect 11940 12655 11945 12695
rect 10495 12650 11945 12655
rect 11195 12350 11245 12650
rect 10495 12345 11945 12350
rect 10495 12305 10500 12345
rect 10540 12305 10850 12345
rect 10890 12305 11200 12345
rect 11240 12305 11550 12345
rect 11590 12305 11900 12345
rect 11940 12305 11945 12345
rect 10495 12300 11945 12305
rect 11195 12000 11245 12300
rect 10495 11995 11945 12000
rect 10495 11955 10500 11995
rect 10540 11955 10850 11995
rect 10890 11955 11200 11995
rect 11240 11955 11550 11995
rect 11590 11955 11900 11995
rect 11940 11955 11945 11995
rect 10495 11950 11945 11955
rect 11195 11650 11245 11950
rect 10495 11645 11945 11650
rect 10495 11605 10500 11645
rect 10540 11605 10850 11645
rect 10890 11605 11200 11645
rect 11240 11605 11550 11645
rect 11590 11605 11900 11645
rect 11940 11605 11945 11645
rect 10495 11600 11945 11605
rect 11195 11300 11245 11600
rect 10495 11295 11945 11300
rect 10495 11255 10500 11295
rect 10540 11255 10850 11295
rect 10890 11255 11200 11295
rect 11240 11255 11550 11295
rect 11590 11255 11900 11295
rect 11940 11255 11945 11295
rect 10495 11250 11945 11255
rect 11195 10950 11245 11250
rect 10495 10945 11945 10950
rect 10495 10905 10500 10945
rect 10540 10905 10850 10945
rect 10890 10905 11200 10945
rect 11240 10905 11550 10945
rect 11590 10905 11900 10945
rect 11940 10905 11945 10945
rect 10495 10900 11945 10905
rect 11195 10600 11245 10900
rect 10495 10595 11945 10600
rect 10495 10555 10500 10595
rect 10540 10555 10850 10595
rect 10890 10555 11200 10595
rect 11240 10555 11550 10595
rect 11590 10555 11900 10595
rect 11940 10555 11945 10595
rect 10495 10550 11945 10555
rect 11195 10250 11245 10550
rect 10495 10245 11945 10250
rect 10495 10205 10500 10245
rect 10540 10205 10850 10245
rect 10890 10205 11200 10245
rect 11240 10205 11550 10245
rect 11590 10205 11900 10245
rect 11940 10205 11945 10245
rect 10495 10200 11945 10205
rect 11195 9900 11245 10200
rect 10495 9895 11945 9900
rect 10495 9855 10500 9895
rect 10540 9855 10850 9895
rect 10890 9855 11200 9895
rect 11240 9855 11550 9895
rect 11590 9855 11900 9895
rect 11940 9855 11945 9895
rect 10495 9850 11945 9855
rect 11195 9550 11245 9850
rect 10495 9545 11945 9550
rect 10495 9505 10500 9545
rect 10540 9505 10850 9545
rect 10890 9505 11200 9545
rect 11240 9505 11550 9545
rect 11590 9505 11900 9545
rect 11940 9505 11945 9545
rect 10495 9500 11945 9505
rect 11195 9200 11245 9500
rect 10495 9195 11945 9200
rect 10495 9155 10500 9195
rect 10540 9155 10850 9195
rect 10890 9155 11200 9195
rect 11240 9155 11550 9195
rect 11590 9155 11900 9195
rect 11940 9155 11945 9195
rect 10495 9150 11945 9155
rect 11195 8850 11245 9150
rect 10495 8845 11945 8850
rect 10495 8805 10500 8845
rect 10540 8805 10850 8845
rect 10890 8805 11200 8845
rect 11240 8805 11550 8845
rect 11590 8805 11900 8845
rect 11940 8805 11945 8845
rect 10495 8800 11945 8805
rect 11195 8500 11245 8800
rect 10495 8495 11945 8500
rect 10495 8455 10500 8495
rect 10540 8455 10850 8495
rect 10890 8455 11200 8495
rect 11240 8455 11550 8495
rect 11590 8455 11900 8495
rect 11940 8455 11945 8495
rect 10495 8450 11945 8455
rect 11195 8150 11245 8450
rect 10495 8145 11945 8150
rect 10495 8105 10500 8145
rect 10540 8105 10850 8145
rect 10890 8105 11200 8145
rect 11240 8105 11550 8145
rect 11590 8105 11900 8145
rect 11940 8105 11945 8145
rect 10495 8100 11945 8105
rect 11195 7800 11245 8100
rect 10495 7795 11945 7800
rect 10495 7755 10500 7795
rect 10540 7755 10850 7795
rect 10890 7755 11200 7795
rect 11240 7755 11550 7795
rect 11590 7755 11900 7795
rect 11940 7755 11945 7795
rect 10495 7750 11945 7755
rect 11195 7450 11245 7750
rect 10495 7445 11945 7450
rect 10495 7405 10500 7445
rect 10540 7405 10850 7445
rect 10890 7405 11200 7445
rect 11240 7405 11550 7445
rect 11590 7405 11900 7445
rect 11940 7405 11945 7445
rect 10495 7400 11945 7405
rect 11195 7100 11245 7400
rect 10495 7095 11945 7100
rect 10495 7055 10500 7095
rect 10540 7055 10850 7095
rect 10890 7055 11200 7095
rect 11240 7055 11550 7095
rect 11590 7055 11900 7095
rect 11940 7055 11945 7095
rect 10495 7050 11945 7055
rect 11195 6750 11245 7050
rect 540 6700 590 6750
rect 9690 6745 11945 6750
rect 9690 6705 10500 6745
rect 10540 6705 10850 6745
rect 10890 6705 11200 6745
rect 11240 6705 11550 6745
rect 11590 6705 11900 6745
rect 11940 6705 11945 6745
rect 9690 6700 11945 6705
rect 11195 6400 11245 6700
rect 10495 6395 11945 6400
rect 10495 6355 10500 6395
rect 10540 6355 10850 6395
rect 10890 6355 11200 6395
rect 11240 6355 11550 6395
rect 11590 6355 11900 6395
rect 11940 6355 11945 6395
rect 10495 6350 11945 6355
rect 11195 6050 11245 6350
rect 10495 6045 11945 6050
rect 10495 6005 10500 6045
rect 10540 6005 10850 6045
rect 10890 6005 11200 6045
rect 11240 6005 11550 6045
rect 11590 6005 11900 6045
rect 11940 6005 11945 6045
rect 10495 6000 11945 6005
rect 11195 5700 11245 6000
rect 10495 5695 11945 5700
rect 10495 5655 10500 5695
rect 10540 5655 10850 5695
rect 10890 5655 11200 5695
rect 11240 5655 11550 5695
rect 11590 5655 11900 5695
rect 11940 5655 11945 5695
rect 10495 5650 11945 5655
rect 11195 5350 11245 5650
rect 10495 5345 11945 5350
rect 10495 5305 10500 5345
rect 10540 5305 10850 5345
rect 10890 5305 11200 5345
rect 11240 5305 11550 5345
rect 11590 5305 11900 5345
rect 11940 5305 11945 5345
rect 10495 5300 11945 5305
rect 11195 5000 11245 5300
rect 10495 4995 11945 5000
rect 10495 4955 10500 4995
rect 10540 4955 10850 4995
rect 10890 4955 11200 4995
rect 11240 4955 11550 4995
rect 11590 4955 11900 4995
rect 11940 4955 11945 4995
rect 10495 4950 11945 4955
rect 11195 4650 11245 4950
rect 10495 4645 11945 4650
rect 10495 4605 10500 4645
rect 10540 4605 10850 4645
rect 10890 4605 11200 4645
rect 11240 4605 11550 4645
rect 11590 4605 11900 4645
rect 11940 4605 11945 4645
rect 10495 4600 11945 4605
rect 11195 4300 11245 4600
rect 10495 4295 11945 4300
rect 10495 4255 10500 4295
rect 10540 4255 10850 4295
rect 10890 4255 11200 4295
rect 11240 4255 11550 4295
rect 11590 4255 11900 4295
rect 11940 4255 11945 4295
rect 10495 4250 11945 4255
rect 11195 3950 11245 4250
rect 10495 3945 11945 3950
rect 10495 3905 10500 3945
rect 10540 3905 10850 3945
rect 10890 3905 11200 3945
rect 11240 3905 11550 3945
rect 11590 3905 11900 3945
rect 11940 3905 11945 3945
rect 10495 3900 11945 3905
rect 11195 3600 11245 3900
rect 10495 3595 11945 3600
rect 10495 3555 10500 3595
rect 10540 3555 10850 3595
rect 10890 3555 11200 3595
rect 11240 3555 11550 3595
rect 11590 3555 11900 3595
rect 11940 3555 11945 3595
rect 10495 3550 11945 3555
rect 11195 3250 11245 3550
rect 10495 3245 11945 3250
rect 10495 3205 10500 3245
rect 10540 3205 10850 3245
rect 10890 3205 11200 3245
rect 11240 3205 11550 3245
rect 11590 3205 11900 3245
rect 11940 3205 11945 3245
rect 10495 3200 11945 3205
rect 11195 2900 11245 3200
rect 10495 2895 11945 2900
rect 10495 2855 10500 2895
rect 10540 2855 10850 2895
rect 10890 2855 11200 2895
rect 11240 2855 11550 2895
rect 11590 2855 11900 2895
rect 11940 2855 11945 2895
rect 10495 2850 11945 2855
rect 11195 2550 11245 2850
rect 10495 2545 11945 2550
rect 10495 2505 10500 2545
rect 10540 2505 10850 2545
rect 10890 2505 11200 2545
rect 11240 2505 11550 2545
rect 11590 2505 11900 2545
rect 11940 2505 11945 2545
rect 10495 2500 11945 2505
rect 11195 2200 11245 2500
rect 10495 2195 11945 2200
rect 10495 2155 10500 2195
rect 10540 2155 10850 2195
rect 10890 2155 11200 2195
rect 11240 2155 11550 2195
rect 11590 2155 11900 2195
rect 11940 2155 11945 2195
rect 10495 2150 11945 2155
rect 11195 1850 11245 2150
rect 10495 1845 11945 1850
rect 10495 1805 10500 1845
rect 10540 1805 10850 1845
rect 10890 1805 11200 1845
rect 11240 1805 11550 1845
rect 11590 1805 11900 1845
rect 11940 1805 11945 1845
rect 10495 1800 11945 1805
rect 11195 1500 11245 1800
rect 10495 1495 11945 1500
rect 10495 1455 10500 1495
rect 10540 1455 10850 1495
rect 10890 1455 11200 1495
rect 11240 1455 11550 1495
rect 11590 1455 11900 1495
rect 11940 1455 11945 1495
rect 10495 1450 11945 1455
rect 11195 1150 11245 1450
rect 10495 1145 11945 1150
rect 10495 1105 10500 1145
rect 10540 1105 10850 1145
rect 10890 1105 11200 1145
rect 11240 1105 11550 1145
rect 11590 1105 11900 1145
rect 11940 1105 11945 1145
rect 10495 1100 11945 1105
rect 11195 800 11245 1100
rect 10495 795 11945 800
rect 10495 755 10500 795
rect 10540 755 10850 795
rect 10890 755 11200 795
rect 11240 755 11550 795
rect 11590 755 11900 795
rect 11940 755 11945 795
rect 10495 750 11945 755
rect 11195 450 11245 750
rect 10495 445 11945 450
rect 10495 405 10500 445
rect 10540 405 10850 445
rect 10890 405 11200 445
rect 11240 405 11550 445
rect 11590 405 11900 445
rect 11940 405 11945 445
rect 10495 400 11945 405
rect 540 0 590 50
rect 9685 45 10235 50
rect 9685 5 10190 45
rect 10230 5 10235 45
rect 9685 0 10235 5
use bgr  bgr_0
timestamp 1752419158
transform -1 0 22845 0 -1 8250
box 15505 -6295 20095 1600
use two_stage_opamp_dummy_magic_21  two_stage_opamp_dummy_magic_21_0
timestamp 1752828052
transform 1 0 -51855 0 1 555
box 51855 -555 61545 6195
<< labels >>
flabel metal4 565 0 565 0 5 FreeSans 800 0 0 -320 GNDA
port 2 s
flabel metal2 4160 2325 4160 2325 7 FreeSans 800 0 -320 0 VIN+
port 5 w
flabel metal2 5930 2325 5930 2325 3 FreeSans 800 0 320 0 VIN-
port 6 e
flabel metal2 2655 1785 2655 1785 5 FreeSans 800 0 0 -320 VOUT+
port 3 s
flabel metal2 7390 1785 7390 1785 5 FreeSans 800 0 0 -320 VOUT-
port 4 s
flabel metal4 565 6750 565 6750 1 FreeSans 800 0 0 320 VDDA
port 1 n
<< end >>
