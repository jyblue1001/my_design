magic
tech sky130A
timestamp 1727625507
use sky130_fd_sc_hd__and2_0  sky130_fd_sc_hd__and2_0_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 0 0 1 0
box -19 -24 249 296
<< end >>
