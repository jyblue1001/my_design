* PEX produced on Sun Feb 16 02:11:13 PM CET 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from pfd_5.ext - technology: sky130A

.subckt pfd_5 F_REF F_VCO VDDA GNDA UP_input DOWN_input I_IN
X0 a_n150_n6120.t1 F_REF.t0 VDDA.t34 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X1 UP.t1 UP_PFD_b.t2 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X2 a_n150_n6880.t1 F_VCO.t0 VDDA.t37 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X3 DOWN_b.t1 GNDA.t60 DOWN_PFD_b.t3 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X4 DOWN_input.t2 DOWN_b.t2 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X5 E.t1 E_b.t3 a_750_n6120.t1 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X6 F.t0 F_b.t3 a_750_n6880.t1 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X7 GNDA.t1 QB.t3 QB_b.t2 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X8 QA.t1 QA_b.t3 GNDA.t28 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X9 E_b.t0 E.t3 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X10 GNDA.t26 a_2410_n7330.t2 a_2080_n7330.t1 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X11 E.t0 QA_b.t4 GNDA.t40 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X12 DOWN_input.t0 DOWN.t2 I_IN.t0 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X13 a_370_n6120.t0 QA_b.t5 QA.t0 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X14 a_1270_n6120.t1 E.t4 E_b.t1 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X15 a_370_n6880.t0 QB_b.t3 QB.t0 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X16 a_1270_n6880.t1 F.t3 F_b.t0 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X17 DOWN.t1 DOWN_b.t3 GNDA.t43 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X18 GNDA.t38 F.t4 QB.t2 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X19 GNDA.t23 Reset.t2 F_b.t2 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X20 a_750_n6120.t0 QA_b.t6 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X21 a_750_n6880.t0 QB_b.t4 VDDA.t16 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X22 DOWN_b.t0 VDDA.t41 DOWN_PFD_b.t2 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X23 UP_PFD_b.t0 QA.t3 GNDA.t17 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X24 QB_b.t0 F_VCO.t1 GNDA.t45 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X25 before_Reset.t0 QA.t4 a_1710_n5500.t0 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X26 VDDA.t20 a_2080_n7330.t2 a_1750_n7330.t0 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X27 GNDA.t15 F_b.t4 F.t1 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X28 GNDA.t13 QA.t5 QA_b.t1 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X29 before_Reset.t1 QA.t6 VDDA.t26 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X30 UP_PFD_b.t1 QA.t7 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X31 VDDA.t30 a_1750_n7330.t2 Reset.t1 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X32 DOWN_PFD_b.t1 QB.t4 VDDA.t31 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X33 UP_input.t0 UP.t2 VDDA.t22 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X34 QA_b.t0 QA.t8 a_n150_n6120.t0 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X35 QB_b.t1 QB.t5 a_n150_n6880.t0 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X36 a_2150_n6120.t1 before_Reset.t3 GNDA.t52 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X37 a_2410_n7330.t0 a_2150_n6120.t2 GNDA.t54 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X38 QB.t1 QB_b.t5 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X39 F_b.t1 F.t5 GNDA.t21 GNDA.t20 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X40 UP_input.t1 UP.t3 opamp_out.t0 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X41 UP_b.t1 UP.t4 GNDA.t56 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X42 GNDA.t32 Reset.t3 E_b.t2 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X43 a_1710_n5500.t1 QB.t6 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X44 GNDA.t9 E.t5 QA.t2 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X45 VDDA.t12 a_2410_n7330.t3 a_2080_n7330.t0 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X46 F.t2 QB_b.t6 GNDA.t34 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X47 a_2150_n6120.t0 before_Reset.t4 VDDA.t36 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X48 a_2410_n7330.t1 a_2150_n6120.t3 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X49 QA_b.t2 F_REF.t1 GNDA.t47 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X50 UP.t0 UP_PFD_b.t3 GNDA.t50 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X51 UP_input.t2 UP_b.t2 opamp_out.t1 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X52 DOWN_input.t1 DOWN_b.t4 I_IN.t1 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X53 GNDA.t19 a_2080_n7330.t3 a_1750_n7330.t1 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X54 UP_b.t0 UP.t5 VDDA.t38 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X55 DOWN.t0 DOWN_b.t5 VDDA.t7 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X56 GNDA.t3 E_b.t4 E.t2 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X57 VDDA.t8 E.t6 a_370_n6120.t1 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X58 VDDA.t1 Reset.t4 a_1270_n6120.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X59 VDDA.t15 QB.t7 before_Reset.t2 VDDA.t14 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X60 VDDA.t3 F.t6 a_370_n6880.t1 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X61 VDDA.t32 Reset.t5 a_1270_n6880.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X62 GNDA.t30 a_1750_n7330.t3 Reset.t0 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X63 DOWN_PFD_b.t0 QB.t8 GNDA.t11 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
R0 F_REF.n0 F_REF.t0 514.134
R1 F_REF.n0 F_REF.t1 273.134
R2 F_REF F_REF.n0 216.9
R3 VDDA.n196 VDDA.n188 831.25
R4 VDDA.n191 VDDA.n190 831.25
R5 VDDA.n185 VDDA.n177 831.25
R6 VDDA.n180 VDDA.n179 831.25
R7 VDDA.n189 VDDA.n188 585
R8 VDDA.n193 VDDA.n191 585
R9 VDDA.n120 VDDA.n115 585
R10 VDDA.n115 VDDA.n34 585
R11 VDDA.n94 VDDA.n40 585
R12 VDDA.n89 VDDA.n40 585
R13 VDDA.n66 VDDA.n60 585
R14 VDDA.n61 VDDA.n60 585
R15 VDDA.n72 VDDA.n46 585
R16 VDDA.n76 VDDA.n46 585
R17 VDDA.n178 VDDA.n177 585
R18 VDDA.n182 VDDA.n180 585
R19 VDDA.n124 VDDA.n35 585
R20 VDDA.n109 VDDA.n35 585
R21 VDDA.n57 VDDA.n51 585
R22 VDDA.n52 VDDA.n51 585
R23 VDDA.n195 VDDA.t10 465.079
R24 VDDA.t10 VDDA.n194 465.079
R25 VDDA.n184 VDDA.t16 465.079
R26 VDDA.t16 VDDA.n183 465.079
R27 VDDA.n105 VDDA.t12 464.281
R28 VDDA.n102 VDDA.t12 464.281
R29 VDDA.t34 VDDA.n169 464.281
R30 VDDA.n170 VDDA.t34 464.281
R31 VDDA.n212 VDDA.t1 464.281
R32 VDDA.t1 VDDA.n211 464.281
R33 VDDA.n226 VDDA.t36 464.281
R34 VDDA.t36 VDDA.n22 464.281
R35 VDDA.n142 VDDA.t40 464.281
R36 VDDA.t40 VDDA.n141 464.281
R37 VDDA.t37 VDDA.n161 464.281
R38 VDDA.n162 VDDA.t37 464.281
R39 VDDA.t32 VDDA.n201 464.281
R40 VDDA.n202 VDDA.t32 464.281
R41 VDDA.t30 VDDA.n216 464.281
R42 VDDA.n217 VDDA.t30 464.281
R43 VDDA.n151 VDDA.t20 464.281
R44 VDDA.t20 VDDA.n150 464.281
R45 VDDA.n83 VDDA.t41 415.336
R46 VDDA.t5 VDDA.t4 314.113
R47 VDDA.t17 VDDA.t18 314.113
R48 VDDA.n118 VDDA.n115 290.733
R49 VDDA.n92 VDDA.n40 290.733
R50 VDDA.n64 VDDA.n60 290.733
R51 VDDA.n70 VDDA.n46 290.733
R52 VDDA.n110 VDDA.n35 290.733
R53 VDDA.n55 VDDA.n51 290.733
R54 VDDA.n169 VDDA.n158 243.698
R55 VDDA.n213 VDDA.n212 243.698
R56 VDDA.n227 VDDA.n226 243.698
R57 VDDA.n143 VDDA.n142 243.698
R58 VDDA.n162 VDDA.n159 243.698
R59 VDDA.n202 VDDA.n199 243.698
R60 VDDA.n217 VDDA.n155 243.698
R61 VDDA.n150 VDDA.n145 243.698
R62 VDDA.n197 VDDA.n196 238.367
R63 VDDA.n190 VDDA.n157 238.367
R64 VDDA.n156 VDDA.n13 238.367
R65 VDDA.n230 VDDA.n229 238.367
R66 VDDA.n138 VDDA.n24 238.367
R67 VDDA.n166 VDDA.n2 238.367
R68 VDDA.n186 VDDA.n185 238.367
R69 VDDA.n206 VDDA.n14 238.367
R70 VDDA.n221 VDDA.n18 238.367
R71 VDDA.n153 VDDA.n152 238.367
R72 VDDA.n179 VDDA.n175 238.367
R73 VDDA.n173 VDDA.n1 238.367
R74 VDDA.n121 VDDA.n120 230.308
R75 VDDA.n97 VDDA.n34 230.308
R76 VDDA.n95 VDDA.n94 230.308
R77 VDDA.n89 VDDA.n38 230.308
R78 VDDA.n67 VDDA.n66 230.308
R79 VDDA.n61 VDDA.n48 230.308
R80 VDDA.n73 VDDA.n72 230.308
R81 VDDA.n76 VDDA.n75 230.308
R82 VDDA.n124 VDDA.n123 230.308
R83 VDDA.n58 VDDA.n57 230.308
R84 VDDA.n52 VDDA.n49 230.308
R85 VDDA.n113 VDDA.n109 230.308
R86 VDDA.n239 VDDA.n17 226.888
R87 VDDA.t13 VDDA.t6 222.178
R88 VDDA.n102 VDDA.n99 190.333
R89 VDDA.n56 VDDA.n50 185
R90 VDDA.n54 VDDA.n53 185
R91 VDDA.n37 VDDA.n36 185
R92 VDDA.n112 VDDA.n111 185
R93 VDDA.n147 VDDA.n146 185
R94 VDDA.n149 VDDA.n148 185
R95 VDDA.n220 VDDA.n219 185
R96 VDDA.n218 VDDA.n215 185
R97 VDDA.n205 VDDA.n204 185
R98 VDDA.n203 VDDA.n200 185
R99 VDDA.n178 VDDA.n176 185
R100 VDDA.n182 VDDA.n181 185
R101 VDDA.n165 VDDA.n164 185
R102 VDDA.n163 VDDA.n160 185
R103 VDDA.n71 VDDA.n69 185
R104 VDDA.n47 VDDA.n45 185
R105 VDDA.n65 VDDA.n59 185
R106 VDDA.n63 VDDA.n62 185
R107 VDDA.n93 VDDA.n39 185
R108 VDDA.n91 VDDA.n90 185
R109 VDDA.n119 VDDA.n114 185
R110 VDDA.n117 VDDA.n116 185
R111 VDDA.n26 VDDA.n25 185
R112 VDDA.n140 VDDA.n139 185
R113 VDDA.n225 VDDA.n223 185
R114 VDDA.n224 VDDA.n23 185
R115 VDDA.n208 VDDA.n207 185
R116 VDDA.n210 VDDA.n209 185
R117 VDDA.n189 VDDA.n187 185
R118 VDDA.n193 VDDA.n192 185
R119 VDDA.n168 VDDA.n167 185
R120 VDDA.n172 VDDA.n171 185
R121 VDDA.n107 VDDA.n106 185
R122 VDDA.n108 VDDA.n107 185
R123 VDDA.n104 VDDA.n100 185
R124 VDDA.n103 VDDA.n101 185
R125 VDDA.n108 VDDA.n99 185
R126 VDDA.n74 VDDA.t13 172.38
R127 VDDA.n68 VDDA.t23 172.38
R128 VDDA.t27 VDDA.n96 172.38
R129 VDDA.n172 VDDA.n167 150
R130 VDDA.n192 VDDA.n187 150
R131 VDDA.n209 VDDA.n207 150
R132 VDDA.n223 VDDA.n23 150
R133 VDDA.n139 VDDA.n25 150
R134 VDDA.n165 VDDA.n160 150
R135 VDDA.n181 VDDA.n176 150
R136 VDDA.n205 VDDA.n200 150
R137 VDDA.n220 VDDA.n215 150
R138 VDDA.n148 VDDA.n146 150
R139 VDDA.n107 VDDA.n100 150
R140 VDDA.n101 VDDA.n99 150
R141 VDDA.t14 VDDA.n214 149.395
R142 VDDA.n122 VDDA.n108 145.565
R143 VDDA.n74 VDDA.t21 126.412
R144 VDDA.t6 VDDA.n68 126.412
R145 VDDA.n96 VDDA.t23 126.412
R146 VDDA.n122 VDDA.t27 126.412
R147 VDDA.t8 VDDA.n188 123.126
R148 VDDA.n191 VDDA.t8 123.126
R149 VDDA.t3 VDDA.n177 123.126
R150 VDDA.n180 VDDA.t3 123.126
R151 VDDA.n116 VDDA.n114 120.001
R152 VDDA.n90 VDDA.n39 120.001
R153 VDDA.n62 VDDA.n59 120.001
R154 VDDA.n69 VDDA.n47 120.001
R155 VDDA.n112 VDDA.n37 120.001
R156 VDDA.n53 VDDA.n50 120.001
R157 VDDA.n214 VDDA.t0 103.427
R158 VDDA.t9 VDDA.n198 103.427
R159 VDDA.n198 VDDA.t2 103.427
R160 VDDA.t33 VDDA.n174 103.427
R161 VDDA.t0 VDDA.t5 84.2747
R162 VDDA.t4 VDDA.t9 84.2747
R163 VDDA.t2 VDDA.t17 84.2747
R164 VDDA.t18 VDDA.t33 84.2747
R165 VDDA.n154 VDDA.n144 76.6134
R166 VDDA.n228 VDDA.n222 76.6134
R167 VDDA.n108 VDDA.t39 72.7828
R168 VDDA.n144 VDDA.t11 72.7828
R169 VDDA.t35 VDDA.n154 72.7828
R170 VDDA.n228 VDDA.t19 72.7828
R171 VDDA.n222 VDDA.t25 72.7828
R172 VDDA.n68 VDDA.n58 69.8479
R173 VDDA.n68 VDDA.n49 69.8479
R174 VDDA.n123 VDDA.n122 69.8479
R175 VDDA.n122 VDDA.n113 69.8479
R176 VDDA.n74 VDDA.n73 69.8479
R177 VDDA.n75 VDDA.n74 69.8479
R178 VDDA.n68 VDDA.n67 69.8479
R179 VDDA.n68 VDDA.n48 69.8479
R180 VDDA.n96 VDDA.n95 69.8479
R181 VDDA.n96 VDDA.n38 69.8479
R182 VDDA.n122 VDDA.n121 69.8479
R183 VDDA.n122 VDDA.n97 69.8479
R184 VDDA.n77 VDDA.n76 66.3886
R185 VDDA.n154 VDDA.n153 65.8183
R186 VDDA.n154 VDDA.n145 65.8183
R187 VDDA.n222 VDDA.n221 65.8183
R188 VDDA.n222 VDDA.n155 65.8183
R189 VDDA.n214 VDDA.n206 65.8183
R190 VDDA.n214 VDDA.n199 65.8183
R191 VDDA.n198 VDDA.n186 65.8183
R192 VDDA.n198 VDDA.n175 65.8183
R193 VDDA.n174 VDDA.n166 65.8183
R194 VDDA.n174 VDDA.n159 65.8183
R195 VDDA.n144 VDDA.n143 65.8183
R196 VDDA.n144 VDDA.n24 65.8183
R197 VDDA.n228 VDDA.n227 65.8183
R198 VDDA.n229 VDDA.n228 65.8183
R199 VDDA.n214 VDDA.n213 65.8183
R200 VDDA.n214 VDDA.n156 65.8183
R201 VDDA.n198 VDDA.n197 65.8183
R202 VDDA.n198 VDDA.n157 65.8183
R203 VDDA.n174 VDDA.n158 65.8183
R204 VDDA.n174 VDDA.n173 65.8183
R205 VDDA.n108 VDDA.n98 65.8183
R206 VDDA.n273 VDDA.n1 58.0576
R207 VDDA.n245 VDDA.n13 58.0576
R208 VDDA.n231 VDDA.n230 58.0576
R209 VDDA.n138 VDDA.n137 58.0576
R210 VDDA.n273 VDDA.n2 58.0576
R211 VDDA.n245 VDDA.n14 58.0576
R212 VDDA.n237 VDDA.n18 58.0576
R213 VDDA.n152 VDDA.n21 58.0576
R214 VDDA.n106 VDDA.n27 58.0576
R215 VDDA.n125 VDDA.n34 57.2449
R216 VDDA.n89 VDDA.n88 57.2449
R217 VDDA.n61 VDDA.n44 57.2449
R218 VDDA.n125 VDDA.n124 57.2449
R219 VDDA.n57 VDDA.n44 57.2449
R220 VDDA.n260 VDDA.n7 54.4005
R221 VDDA.n258 VDDA.n7 54.4005
R222 VDDA.n258 VDDA.n8 54.4005
R223 VDDA.n260 VDDA.n8 54.4005
R224 VDDA.t29 VDDA.t14 53.6295
R225 VDDA.n167 VDDA.n158 53.3664
R226 VDDA.n173 VDDA.n172 53.3664
R227 VDDA.n160 VDDA.n159 53.3664
R228 VDDA.n181 VDDA.n175 53.3664
R229 VDDA.n200 VDDA.n199 53.3664
R230 VDDA.n153 VDDA.n146 53.3664
R231 VDDA.n148 VDDA.n145 53.3664
R232 VDDA.n221 VDDA.n220 53.3664
R233 VDDA.n215 VDDA.n155 53.3664
R234 VDDA.n206 VDDA.n205 53.3664
R235 VDDA.n186 VDDA.n176 53.3664
R236 VDDA.n166 VDDA.n165 53.3664
R237 VDDA.n143 VDDA.n25 53.3664
R238 VDDA.n139 VDDA.n24 53.3664
R239 VDDA.n227 VDDA.n223 53.3664
R240 VDDA.n229 VDDA.n23 53.3664
R241 VDDA.n213 VDDA.n207 53.3664
R242 VDDA.n209 VDDA.n156 53.3664
R243 VDDA.n197 VDDA.n187 53.3664
R244 VDDA.n192 VDDA.n157 53.3664
R245 VDDA.n100 VDDA.n98 53.3664
R246 VDDA.n101 VDDA.n98 53.3664
R247 VDDA.n113 VDDA.n112 45.3071
R248 VDDA.n53 VDDA.n49 45.3071
R249 VDDA.n58 VDDA.n50 45.3071
R250 VDDA.n123 VDDA.n37 45.3071
R251 VDDA.n73 VDDA.n69 45.3071
R252 VDDA.n75 VDDA.n47 45.3071
R253 VDDA.n67 VDDA.n59 45.3071
R254 VDDA.n62 VDDA.n48 45.3071
R255 VDDA.n95 VDDA.n39 45.3071
R256 VDDA.n90 VDDA.n38 45.3071
R257 VDDA.n121 VDDA.n114 45.3071
R258 VDDA.n116 VDDA.n97 45.3071
R259 VDDA.n274 VDDA.n273 34.9005
R260 VDDA.n80 VDDA.n79 32.0005
R261 VDDA.n81 VDDA.n80 32.0005
R262 VDDA.n81 VDDA.n41 32.0005
R263 VDDA.n87 VDDA.n42 32.0005
R264 VDDA.n42 VDDA.n33 32.0005
R265 VDDA.n126 VDDA.n33 32.0005
R266 VDDA.n130 VDDA.n31 32.0005
R267 VDDA.n131 VDDA.n130 32.0005
R268 VDDA.n132 VDDA.n131 32.0005
R269 VDDA.n136 VDDA.n29 32.0005
R270 VDDA.n29 VDDA.n28 32.0005
R271 VDDA.n236 VDDA.n19 32.0005
R272 VDDA.n240 VDDA.n15 32.0005
R273 VDDA.n244 VDDA.n15 32.0005
R274 VDDA.n247 VDDA.n246 32.0005
R275 VDDA.n247 VDDA.n11 32.0005
R276 VDDA.n251 VDDA.n11 32.0005
R277 VDDA.n252 VDDA.n251 32.0005
R278 VDDA.n253 VDDA.n252 32.0005
R279 VDDA.n253 VDDA.n9 32.0005
R280 VDDA.n257 VDDA.n9 32.0005
R281 VDDA.n261 VDDA.n5 32.0005
R282 VDDA.n265 VDDA.n5 32.0005
R283 VDDA.n266 VDDA.n265 32.0005
R284 VDDA.n267 VDDA.n266 32.0005
R285 VDDA.n267 VDDA.n3 32.0005
R286 VDDA.n271 VDDA.n3 32.0005
R287 VDDA.n272 VDDA.n271 32.0005
R288 VDDA.t39 VDDA.t11 30.6457
R289 VDDA.t19 VDDA.t35 30.6457
R290 VDDA.t25 VDDA.t29 30.6457
R291 VDDA.n77 VDDA.n44 29.8986
R292 VDDA.n231 VDDA.n19 25.6005
R293 VDDA.n237 VDDA.n236 25.6005
R294 VDDA.n245 VDDA.n244 25.6005
R295 VDDA.n259 VDDA.n258 25.6005
R296 VDDA.n260 VDDA.n259 25.6005
R297 VDDA.n115 VDDA.t28 24.6255
R298 VDDA.n40 VDDA.t24 24.6255
R299 VDDA.n60 VDDA.t38 24.6255
R300 VDDA.n46 VDDA.t22 24.6255
R301 VDDA.n35 VDDA.t31 24.6255
R302 VDDA.n51 VDDA.t7 24.6255
R303 VDDA.n137 VDDA.n27 22.4005
R304 VDDA.n17 VDDA.t26 19.7005
R305 VDDA.n17 VDDA.t15 19.7005
R306 VDDA.n88 VDDA.n41 19.2005
R307 VDDA.n240 VDDA.n239 19.2005
R308 VDDA.n126 VDDA.n125 16.0005
R309 VDDA.n125 VDDA.n31 16.0005
R310 VDDA.n28 VDDA.n21 16.0005
R311 VDDA.n232 VDDA.n21 16.0005
R312 VDDA.n88 VDDA.n87 12.8005
R313 VDDA.n239 VDDA.n238 12.8005
R314 VDDA.n79 VDDA.n44 9.6005
R315 VDDA.n79 VDDA.n78 9.3005
R316 VDDA.n80 VDDA.n43 9.3005
R317 VDDA.n82 VDDA.n81 9.3005
R318 VDDA.n84 VDDA.n41 9.3005
R319 VDDA.n87 VDDA.n86 9.3005
R320 VDDA.n85 VDDA.n42 9.3005
R321 VDDA.n33 VDDA.n32 9.3005
R322 VDDA.n127 VDDA.n126 9.3005
R323 VDDA.n128 VDDA.n31 9.3005
R324 VDDA.n130 VDDA.n129 9.3005
R325 VDDA.n131 VDDA.n30 9.3005
R326 VDDA.n133 VDDA.n132 9.3005
R327 VDDA.n136 VDDA.n135 9.3005
R328 VDDA.n134 VDDA.n29 9.3005
R329 VDDA.n28 VDDA.n20 9.3005
R330 VDDA.n233 VDDA.n232 9.3005
R331 VDDA.n234 VDDA.n19 9.3005
R332 VDDA.n236 VDDA.n235 9.3005
R333 VDDA.n238 VDDA.n16 9.3005
R334 VDDA.n241 VDDA.n240 9.3005
R335 VDDA.n242 VDDA.n15 9.3005
R336 VDDA.n244 VDDA.n243 9.3005
R337 VDDA.n246 VDDA.n12 9.3005
R338 VDDA.n248 VDDA.n247 9.3005
R339 VDDA.n249 VDDA.n11 9.3005
R340 VDDA.n251 VDDA.n250 9.3005
R341 VDDA.n252 VDDA.n10 9.3005
R342 VDDA.n254 VDDA.n253 9.3005
R343 VDDA.n255 VDDA.n9 9.3005
R344 VDDA.n257 VDDA.n256 9.3005
R345 VDDA.n259 VDDA.n6 9.3005
R346 VDDA.n262 VDDA.n261 9.3005
R347 VDDA.n263 VDDA.n5 9.3005
R348 VDDA.n265 VDDA.n264 9.3005
R349 VDDA.n266 VDDA.n4 9.3005
R350 VDDA.n268 VDDA.n267 9.3005
R351 VDDA.n269 VDDA.n3 9.3005
R352 VDDA.n271 VDDA.n270 9.3005
R353 VDDA.n272 VDDA.n0 9.3005
R354 VDDA.n171 VDDA.n168 9.14336
R355 VDDA.n210 VDDA.n208 9.14336
R356 VDDA.n225 VDDA.n224 9.14336
R357 VDDA.n140 VDDA.n26 9.14336
R358 VDDA.n164 VDDA.n163 9.14336
R359 VDDA.n204 VDDA.n203 9.14336
R360 VDDA.n219 VDDA.n218 9.14336
R361 VDDA.n149 VDDA.n147 9.14336
R362 VDDA.n104 VDDA.n103 9.14336
R363 VDDA.n120 VDDA.n119 7.11161
R364 VDDA.n117 VDDA.n34 7.11161
R365 VDDA.n94 VDDA.n93 7.11161
R366 VDDA.n91 VDDA.n89 7.11161
R367 VDDA.n66 VDDA.n65 7.11161
R368 VDDA.n63 VDDA.n61 7.11161
R369 VDDA.n72 VDDA.n71 7.11161
R370 VDDA.n76 VDDA.n45 7.11161
R371 VDDA.n124 VDDA.n36 7.11161
R372 VDDA.n111 VDDA.n109 7.11161
R373 VDDA.n57 VDDA.n56 7.11161
R374 VDDA.n54 VDDA.n52 7.11161
R375 VDDA.n132 VDDA.n27 6.4005
R376 VDDA.n232 VDDA.n231 6.4005
R377 VDDA.n238 VDDA.n237 6.4005
R378 VDDA.n246 VDDA.n245 6.4005
R379 VDDA.n258 VDDA.n257 6.4005
R380 VDDA.n261 VDDA.n260 6.4005
R381 VDDA.n273 VDDA.n272 6.4005
R382 VDDA.n193 VDDA.n189 5.81868
R383 VDDA.n182 VDDA.n178 5.81868
R384 VDDA.n106 VDDA.n105 5.33286
R385 VDDA.n170 VDDA.n1 5.33286
R386 VDDA.n211 VDDA.n13 5.33286
R387 VDDA.n230 VDDA.n22 5.33286
R388 VDDA.n141 VDDA.n138 5.33286
R389 VDDA.n161 VDDA.n2 5.33286
R390 VDDA.n201 VDDA.n14 5.33286
R391 VDDA.n216 VDDA.n18 5.33286
R392 VDDA.n152 VDDA.n151 5.33286
R393 VDDA.n169 VDDA.n168 3.75335
R394 VDDA.n171 VDDA.n170 3.75335
R395 VDDA.n212 VDDA.n208 3.75335
R396 VDDA.n211 VDDA.n210 3.75335
R397 VDDA.n226 VDDA.n225 3.75335
R398 VDDA.n224 VDDA.n22 3.75335
R399 VDDA.n142 VDDA.n26 3.75335
R400 VDDA.n141 VDDA.n140 3.75335
R401 VDDA.n164 VDDA.n161 3.75335
R402 VDDA.n163 VDDA.n162 3.75335
R403 VDDA.n204 VDDA.n201 3.75335
R404 VDDA.n203 VDDA.n202 3.75335
R405 VDDA.n219 VDDA.n216 3.75335
R406 VDDA.n218 VDDA.n217 3.75335
R407 VDDA.n151 VDDA.n147 3.75335
R408 VDDA.n150 VDDA.n149 3.75335
R409 VDDA.n105 VDDA.n104 3.75335
R410 VDDA.n103 VDDA.n102 3.75335
R411 VDDA.n119 VDDA.n118 3.53508
R412 VDDA.n118 VDDA.n117 3.53508
R413 VDDA.n93 VDDA.n92 3.53508
R414 VDDA.n92 VDDA.n91 3.53508
R415 VDDA.n65 VDDA.n64 3.53508
R416 VDDA.n64 VDDA.n63 3.53508
R417 VDDA.n71 VDDA.n70 3.53508
R418 VDDA.n70 VDDA.n45 3.53508
R419 VDDA.n110 VDDA.n36 3.53508
R420 VDDA.n111 VDDA.n110 3.53508
R421 VDDA.n56 VDDA.n55 3.53508
R422 VDDA.n55 VDDA.n54 3.53508
R423 VDDA.n196 VDDA.n195 3.40194
R424 VDDA.n194 VDDA.n190 3.40194
R425 VDDA.n185 VDDA.n184 3.40194
R426 VDDA.n183 VDDA.n179 3.40194
R427 VDDA.n137 VDDA.n136 3.2005
R428 VDDA.n195 VDDA.n189 2.39444
R429 VDDA.n194 VDDA.n193 2.39444
R430 VDDA.n184 VDDA.n178 2.39444
R431 VDDA.n183 VDDA.n182 2.39444
R432 VDDA.n190 VDDA.n7 2.32777
R433 VDDA.n185 VDDA.n8 2.32777
R434 VDDA.n78 VDDA.n77 0.1943
R435 VDDA.n78 VDDA.n43 0.15675
R436 VDDA.n82 VDDA.n43 0.15675
R437 VDDA.n86 VDDA.n84 0.15675
R438 VDDA.n86 VDDA.n85 0.15675
R439 VDDA.n85 VDDA.n32 0.15675
R440 VDDA.n127 VDDA.n32 0.15675
R441 VDDA.n128 VDDA.n127 0.15675
R442 VDDA.n129 VDDA.n128 0.15675
R443 VDDA.n129 VDDA.n30 0.15675
R444 VDDA.n133 VDDA.n30 0.15675
R445 VDDA.n135 VDDA.n133 0.15675
R446 VDDA.n135 VDDA.n134 0.15675
R447 VDDA.n134 VDDA.n20 0.15675
R448 VDDA.n233 VDDA.n20 0.15675
R449 VDDA.n234 VDDA.n233 0.15675
R450 VDDA.n235 VDDA.n234 0.15675
R451 VDDA.n235 VDDA.n16 0.15675
R452 VDDA.n241 VDDA.n16 0.15675
R453 VDDA.n242 VDDA.n241 0.15675
R454 VDDA.n243 VDDA.n242 0.15675
R455 VDDA.n243 VDDA.n12 0.15675
R456 VDDA.n248 VDDA.n12 0.15675
R457 VDDA.n249 VDDA.n248 0.15675
R458 VDDA.n250 VDDA.n249 0.15675
R459 VDDA.n250 VDDA.n10 0.15675
R460 VDDA.n254 VDDA.n10 0.15675
R461 VDDA.n255 VDDA.n254 0.15675
R462 VDDA.n256 VDDA.n255 0.15675
R463 VDDA.n256 VDDA.n6 0.15675
R464 VDDA.n262 VDDA.n6 0.15675
R465 VDDA.n263 VDDA.n262 0.15675
R466 VDDA.n264 VDDA.n263 0.15675
R467 VDDA.n264 VDDA.n4 0.15675
R468 VDDA.n268 VDDA.n4 0.15675
R469 VDDA.n269 VDDA.n268 0.15675
R470 VDDA.n270 VDDA.n269 0.15675
R471 VDDA.n270 VDDA.n0 0.15675
R472 VDDA.n274 VDDA.n0 0.15675
R473 VDDA.n84 VDDA.n83 0.1255
R474 VDDA VDDA.n274 0.1255
R475 VDDA.n83 VDDA.n82 0.03175
R476 a_n150_n6120.t0 a_n150_n6120.t1 39.4005
R477 UP_PFD_b.n0 UP_PFD_b.t2 441.834
R478 UP_PFD_b.n0 UP_PFD_b.t3 313.3
R479 UP_PFD_b.n1 UP_PFD_b.n0 235.201
R480 UP_PFD_b.t1 UP_PFD_b.n1 219.528
R481 UP_PFD_b.n1 UP_PFD_b.t0 167.935
R482 UP.n0 UP.t2 1205
R483 UP.n2 UP.t5 522.168
R484 UP.n1 UP.n0 441.834
R485 UP.n3 UP.n2 235.201
R486 UP.t1 UP.n3 229.127
R487 UP.n1 UP.t4 217.905
R488 UP.n0 UP.t3 208.868
R489 UP.n3 UP.t0 158.335
R490 UP.n2 UP.n1 15.063
R491 F_VCO.n0 F_VCO.t0 514.134
R492 F_VCO.n0 F_VCO.t1 273.134
R493 F_VCO F_VCO.n0 216.9
R494 a_n150_n6880.t0 a_n150_n6880.t1 39.4005
R495 GNDA.n149 GNDA.n148 21560
R496 GNDA.t4 GNDA.t2 3006.67
R497 GNDA.t27 GNDA.t12 3006.67
R498 GNDA.t20 GNDA.t14 3006.67
R499 GNDA.t35 GNDA.t0 3006.67
R500 GNDA.t48 GNDA.t10 2860
R501 GNDA.n73 GNDA.t53 2163.33
R502 GNDA.t55 GNDA.t57 2126.67
R503 GNDA.t41 GNDA.t42 2126.67
R504 GNDA.t29 GNDA.n152 1943.33
R505 GNDA.n76 GNDA.t49 1723.33
R506 GNDA.n75 GNDA.t16 1723.33
R507 GNDA.n31 GNDA.t41 1650
R508 GNDA.n30 GNDA.t48 1650
R509 GNDA.t51 GNDA.n109 1430
R510 GNDA.t24 GNDA.n110 1430
R511 GNDA.n114 GNDA.t58 1430
R512 GNDA.t25 GNDA.n154 1430
R513 GNDA.t18 GNDA.n153 1430
R514 GNDA.n155 GNDA.n52 1393.33
R515 GNDA.n31 GNDA.t6 1210
R516 GNDA.t42 GNDA.n30 1210
R517 GNDA.n52 GNDA.t10 1210
R518 GNDA.n76 GNDA.t55 1136.67
R519 GNDA.t49 GNDA.n75 1136.67
R520 GNDA.t16 GNDA.n73 1136.67
R521 GNDA.n109 GNDA.t53 990
R522 GNDA.n110 GNDA.t51 990
R523 GNDA.n114 GNDA.t31 990
R524 GNDA.t39 GNDA.n113 990
R525 GNDA.n113 GNDA.t8 990
R526 GNDA.n148 GNDA.t46 990
R527 GNDA.n155 GNDA.t25 990
R528 GNDA.n154 GNDA.t18 990
R529 GNDA.n153 GNDA.t29 990
R530 GNDA.n152 GNDA.t22 990
R531 GNDA.t33 GNDA.n151 990
R532 GNDA.n151 GNDA.t37 990
R533 GNDA.t44 GNDA.n149 990
R534 GNDA.t58 GNDA.t24 806.668
R535 GNDA.t31 GNDA.t4 806.668
R536 GNDA.t2 GNDA.t39 806.668
R537 GNDA.t8 GNDA.t27 806.668
R538 GNDA.t12 GNDA.t46 806.668
R539 GNDA.t22 GNDA.t20 806.668
R540 GNDA.t14 GNDA.t33 806.668
R541 GNDA.t37 GNDA.t35 806.668
R542 GNDA.t0 GNDA.t44 806.668
R543 GNDA.n110 GNDA.t52 715.004
R544 GNDA.n151 GNDA.n150 585.003
R545 GNDA.n113 GNDA.n112 585.003
R546 GNDA.n115 GNDA.n114 585.001
R547 GNDA.n109 GNDA.n108 585.001
R548 GNDA.n77 GNDA.n76 585.001
R549 GNDA.n75 GNDA.n74 585.001
R550 GNDA.n73 GNDA.n72 585.001
R551 GNDA.n148 GNDA.n147 585.001
R552 GNDA.n32 GNDA.n31 585.001
R553 GNDA.n30 GNDA.n29 585.001
R554 GNDA.n52 GNDA.n51 585.001
R555 GNDA.n156 GNDA.n155 585.001
R556 GNDA.n154 GNDA.n19 585.001
R557 GNDA.n153 GNDA.n16 585.001
R558 GNDA.n152 GNDA.n13 585.001
R559 GNDA.n149 GNDA.n2 585.001
R560 GNDA.n40 GNDA.t60 566.966
R561 GNDA.n3 GNDA.t1 198.058
R562 GNDA.n197 GNDA.t36 198.058
R563 GNDA.n185 GNDA.t15 198.058
R564 GNDA.n11 GNDA.t21 198.058
R565 GNDA.n141 GNDA.t13 198.058
R566 GNDA.n55 GNDA.t28 198.058
R567 GNDA.n127 GNDA.t3 198.058
R568 GNDA.n122 GNDA.t5 198.058
R569 GNDA.n94 GNDA.t59 198.058
R570 GNDA.n7 GNDA.t38 130.713
R571 GNDA.n13 GNDA.t23 130.001
R572 GNDA.n16 GNDA.t30 130.001
R573 GNDA.n19 GNDA.t19 130.001
R574 GNDA.n156 GNDA.t26 130.001
R575 GNDA.n147 GNDA.t47 130.001
R576 GNDA.n115 GNDA.t32 130.001
R577 GNDA.n108 GNDA.t54 130.001
R578 GNDA.n2 GNDA.t45 130.001
R579 GNDA.n8 GNDA.t34 130.001
R580 GNDA.n111 GNDA.t40 130.001
R581 GNDA.n57 GNDA.t9 130.001
R582 GNDA.n51 GNDA.t11 122.501
R583 GNDA.n29 GNDA.t43 122.501
R584 GNDA.n32 GNDA.t7 122.501
R585 GNDA.n72 GNDA.t17 122.501
R586 GNDA.n74 GNDA.t50 122.501
R587 GNDA.n77 GNDA.t56 122.501
R588 GNDA.n78 GNDA.n77 70.8139
R589 GNDA.n33 GNDA.n32 68.1246
R590 GNDA.n177 GNDA.n13 60.29
R591 GNDA.n170 GNDA.n16 60.29
R592 GNDA.n164 GNDA.n19 60.29
R593 GNDA.n157 GNDA.n156 60.29
R594 GNDA.n147 GNDA.n146 60.29
R595 GNDA.n116 GNDA.n115 60.29
R596 GNDA.n108 GNDA.n107 60.29
R597 GNDA.n205 GNDA.n2 60.29
R598 GNDA.n72 GNDA.n68 59.5478
R599 GNDA.n74 GNDA.n71 59.5478
R600 GNDA.n51 GNDA.n50 58.9809
R601 GNDA.n29 GNDA.n28 58.9809
R602 GNDA.n190 GNDA.n8 54.4005
R603 GNDA.n192 GNDA.n7 54.4005
R604 GNDA.n133 GNDA.n57 54.4005
R605 GNDA.n111 GNDA.n58 54.4005
R606 GNDA.n146 GNDA.n0 33.0991
R607 GNDA.n206 GNDA.n205 33.0991
R608 GNDA.n81 GNDA.n70 32.0005
R609 GNDA.n82 GNDA.n81 32.0005
R610 GNDA.n83 GNDA.n82 32.0005
R611 GNDA.n87 GNDA.n86 32.0005
R612 GNDA.n88 GNDA.n87 32.0005
R613 GNDA.n88 GNDA.n65 32.0005
R614 GNDA.n106 GNDA.n66 32.0005
R615 GNDA.n102 GNDA.n66 32.0005
R616 GNDA.n102 GNDA.n101 32.0005
R617 GNDA.n101 GNDA.n100 32.0005
R618 GNDA.n100 GNDA.n92 32.0005
R619 GNDA.n96 GNDA.n92 32.0005
R620 GNDA.n96 GNDA.n95 32.0005
R621 GNDA.n117 GNDA.n64 32.0005
R622 GNDA.n121 GNDA.n62 32.0005
R623 GNDA.n122 GNDA.n121 32.0005
R624 GNDA.n123 GNDA.n122 32.0005
R625 GNDA.n123 GNDA.n60 32.0005
R626 GNDA.n127 GNDA.n60 32.0005
R627 GNDA.n128 GNDA.n127 32.0005
R628 GNDA.n129 GNDA.n128 32.0005
R629 GNDA.n135 GNDA.n134 32.0005
R630 GNDA.n135 GNDA.n55 32.0005
R631 GNDA.n139 GNDA.n55 32.0005
R632 GNDA.n140 GNDA.n139 32.0005
R633 GNDA.n141 GNDA.n140 32.0005
R634 GNDA.n141 GNDA.n53 32.0005
R635 GNDA.n145 GNDA.n53 32.0005
R636 GNDA.n36 GNDA.n35 32.0005
R637 GNDA.n37 GNDA.n36 32.0005
R638 GNDA.n37 GNDA.n26 32.0005
R639 GNDA.n42 GNDA.n26 32.0005
R640 GNDA.n43 GNDA.n42 32.0005
R641 GNDA.n44 GNDA.n43 32.0005
R642 GNDA.n44 GNDA.n23 32.0005
R643 GNDA.n49 GNDA.n24 32.0005
R644 GNDA.n24 GNDA.n22 32.0005
R645 GNDA.n158 GNDA.n22 32.0005
R646 GNDA.n162 GNDA.n20 32.0005
R647 GNDA.n163 GNDA.n162 32.0005
R648 GNDA.n165 GNDA.n17 32.0005
R649 GNDA.n169 GNDA.n17 32.0005
R650 GNDA.n172 GNDA.n171 32.0005
R651 GNDA.n172 GNDA.n14 32.0005
R652 GNDA.n176 GNDA.n14 32.0005
R653 GNDA.n179 GNDA.n178 32.0005
R654 GNDA.n179 GNDA.n11 32.0005
R655 GNDA.n183 GNDA.n11 32.0005
R656 GNDA.n184 GNDA.n183 32.0005
R657 GNDA.n185 GNDA.n184 32.0005
R658 GNDA.n185 GNDA.n9 32.0005
R659 GNDA.n189 GNDA.n9 32.0005
R660 GNDA.n193 GNDA.n5 32.0005
R661 GNDA.n197 GNDA.n5 32.0005
R662 GNDA.n198 GNDA.n197 32.0005
R663 GNDA.n199 GNDA.n198 32.0005
R664 GNDA.n199 GNDA.n3 32.0005
R665 GNDA.n203 GNDA.n3 32.0005
R666 GNDA.n204 GNDA.n203 32.0005
R667 GNDA.n33 GNDA.n28 29.8986
R668 GNDA.n107 GNDA.n65 28.8005
R669 GNDA.n78 GNDA.n71 26.6601
R670 GNDA.n117 GNDA.n116 25.6005
R671 GNDA.n132 GNDA.n58 25.6005
R672 GNDA.n133 GNDA.n132 25.6005
R673 GNDA.n157 GNDA.n20 25.6005
R674 GNDA.n170 GNDA.n169 25.6005
R675 GNDA.n177 GNDA.n176 25.6005
R676 GNDA.n191 GNDA.n190 25.6005
R677 GNDA.n192 GNDA.n191 22.4005
R678 GNDA.n95 GNDA.n94 19.2005
R679 GNDA.n83 GNDA.n68 16.0005
R680 GNDA.n86 GNDA.n68 16.0005
R681 GNDA.n50 GNDA.n23 16.0005
R682 GNDA.n50 GNDA.n49 16.0005
R683 GNDA.n164 GNDA.n163 16.0005
R684 GNDA.n165 GNDA.n164 16.0005
R685 GNDA.n71 GNDA.n70 12.8005
R686 GNDA.n94 GNDA.n64 12.8005
R687 GNDA GNDA.n0 12.7806
R688 GNDA GNDA.n206 11.8876
R689 GNDA.n35 GNDA.n28 9.6005
R690 GNDA.n193 GNDA.n192 9.6005
R691 GNDA.n79 GNDA.n70 9.3005
R692 GNDA.n81 GNDA.n80 9.3005
R693 GNDA.n82 GNDA.n69 9.3005
R694 GNDA.n84 GNDA.n83 9.3005
R695 GNDA.n86 GNDA.n85 9.3005
R696 GNDA.n87 GNDA.n67 9.3005
R697 GNDA.n89 GNDA.n88 9.3005
R698 GNDA.n90 GNDA.n65 9.3005
R699 GNDA.n106 GNDA.n105 9.3005
R700 GNDA.n104 GNDA.n66 9.3005
R701 GNDA.n103 GNDA.n102 9.3005
R702 GNDA.n101 GNDA.n91 9.3005
R703 GNDA.n100 GNDA.n99 9.3005
R704 GNDA.n98 GNDA.n92 9.3005
R705 GNDA.n97 GNDA.n96 9.3005
R706 GNDA.n95 GNDA.n93 9.3005
R707 GNDA.n64 GNDA.n63 9.3005
R708 GNDA.n118 GNDA.n117 9.3005
R709 GNDA.n119 GNDA.n62 9.3005
R710 GNDA.n121 GNDA.n120 9.3005
R711 GNDA.n122 GNDA.n61 9.3005
R712 GNDA.n124 GNDA.n123 9.3005
R713 GNDA.n125 GNDA.n60 9.3005
R714 GNDA.n127 GNDA.n126 9.3005
R715 GNDA.n128 GNDA.n59 9.3005
R716 GNDA.n130 GNDA.n129 9.3005
R717 GNDA.n132 GNDA.n131 9.3005
R718 GNDA.n134 GNDA.n56 9.3005
R719 GNDA.n136 GNDA.n135 9.3005
R720 GNDA.n137 GNDA.n55 9.3005
R721 GNDA.n139 GNDA.n138 9.3005
R722 GNDA.n140 GNDA.n54 9.3005
R723 GNDA.n142 GNDA.n141 9.3005
R724 GNDA.n143 GNDA.n53 9.3005
R725 GNDA.n145 GNDA.n144 9.3005
R726 GNDA.n35 GNDA.n34 9.3005
R727 GNDA.n36 GNDA.n27 9.3005
R728 GNDA.n38 GNDA.n37 9.3005
R729 GNDA.n39 GNDA.n26 9.3005
R730 GNDA.n42 GNDA.n41 9.3005
R731 GNDA.n43 GNDA.n25 9.3005
R732 GNDA.n45 GNDA.n44 9.3005
R733 GNDA.n46 GNDA.n23 9.3005
R734 GNDA.n49 GNDA.n48 9.3005
R735 GNDA.n47 GNDA.n24 9.3005
R736 GNDA.n22 GNDA.n21 9.3005
R737 GNDA.n159 GNDA.n158 9.3005
R738 GNDA.n160 GNDA.n20 9.3005
R739 GNDA.n162 GNDA.n161 9.3005
R740 GNDA.n163 GNDA.n18 9.3005
R741 GNDA.n166 GNDA.n165 9.3005
R742 GNDA.n167 GNDA.n17 9.3005
R743 GNDA.n169 GNDA.n168 9.3005
R744 GNDA.n171 GNDA.n15 9.3005
R745 GNDA.n173 GNDA.n172 9.3005
R746 GNDA.n174 GNDA.n14 9.3005
R747 GNDA.n176 GNDA.n175 9.3005
R748 GNDA.n178 GNDA.n12 9.3005
R749 GNDA.n180 GNDA.n179 9.3005
R750 GNDA.n181 GNDA.n11 9.3005
R751 GNDA.n183 GNDA.n182 9.3005
R752 GNDA.n184 GNDA.n10 9.3005
R753 GNDA.n186 GNDA.n185 9.3005
R754 GNDA.n187 GNDA.n9 9.3005
R755 GNDA.n189 GNDA.n188 9.3005
R756 GNDA.n191 GNDA.n6 9.3005
R757 GNDA.n194 GNDA.n193 9.3005
R758 GNDA.n195 GNDA.n5 9.3005
R759 GNDA.n197 GNDA.n196 9.3005
R760 GNDA.n198 GNDA.n4 9.3005
R761 GNDA.n200 GNDA.n199 9.3005
R762 GNDA.n201 GNDA.n3 9.3005
R763 GNDA.n203 GNDA.n202 9.3005
R764 GNDA.n204 GNDA.n1 9.3005
R765 GNDA.n116 GNDA.n62 6.4005
R766 GNDA.n129 GNDA.n58 6.4005
R767 GNDA.n134 GNDA.n133 6.4005
R768 GNDA.n146 GNDA.n145 6.4005
R769 GNDA.n158 GNDA.n157 6.4005
R770 GNDA.n171 GNDA.n170 6.4005
R771 GNDA.n178 GNDA.n177 6.4005
R772 GNDA.n190 GNDA.n189 6.4005
R773 GNDA.n205 GNDA.n204 6.4005
R774 GNDA.n150 GNDA.n8 5.68939
R775 GNDA.n112 GNDA.n111 5.68939
R776 GNDA.n112 GNDA.n57 5.68939
R777 GNDA.n150 GNDA.n7 4.97828
R778 GNDA.n107 GNDA.n106 3.2005
R779 GNDA.n79 GNDA.n78 0.232799
R780 GNDA.n34 GNDA.n33 0.1943
R781 GNDA.n144 GNDA.n0 0.193881
R782 GNDA.n206 GNDA.n1 0.193881
R783 GNDA.n80 GNDA.n79 0.15675
R784 GNDA.n80 GNDA.n69 0.15675
R785 GNDA.n84 GNDA.n69 0.15675
R786 GNDA.n85 GNDA.n84 0.15675
R787 GNDA.n85 GNDA.n67 0.15675
R788 GNDA.n89 GNDA.n67 0.15675
R789 GNDA.n90 GNDA.n89 0.15675
R790 GNDA.n105 GNDA.n90 0.15675
R791 GNDA.n105 GNDA.n104 0.15675
R792 GNDA.n104 GNDA.n103 0.15675
R793 GNDA.n103 GNDA.n91 0.15675
R794 GNDA.n99 GNDA.n91 0.15675
R795 GNDA.n99 GNDA.n98 0.15675
R796 GNDA.n98 GNDA.n97 0.15675
R797 GNDA.n97 GNDA.n93 0.15675
R798 GNDA.n93 GNDA.n63 0.15675
R799 GNDA.n118 GNDA.n63 0.15675
R800 GNDA.n119 GNDA.n118 0.15675
R801 GNDA.n120 GNDA.n119 0.15675
R802 GNDA.n120 GNDA.n61 0.15675
R803 GNDA.n124 GNDA.n61 0.15675
R804 GNDA.n125 GNDA.n124 0.15675
R805 GNDA.n126 GNDA.n125 0.15675
R806 GNDA.n126 GNDA.n59 0.15675
R807 GNDA.n130 GNDA.n59 0.15675
R808 GNDA.n131 GNDA.n130 0.15675
R809 GNDA.n131 GNDA.n56 0.15675
R810 GNDA.n136 GNDA.n56 0.15675
R811 GNDA.n137 GNDA.n136 0.15675
R812 GNDA.n138 GNDA.n137 0.15675
R813 GNDA.n138 GNDA.n54 0.15675
R814 GNDA.n142 GNDA.n54 0.15675
R815 GNDA.n143 GNDA.n142 0.15675
R816 GNDA.n144 GNDA.n143 0.15675
R817 GNDA.n34 GNDA.n27 0.15675
R818 GNDA.n38 GNDA.n27 0.15675
R819 GNDA.n39 GNDA.n38 0.15675
R820 GNDA.n41 GNDA.n25 0.15675
R821 GNDA.n45 GNDA.n25 0.15675
R822 GNDA.n46 GNDA.n45 0.15675
R823 GNDA.n48 GNDA.n46 0.15675
R824 GNDA.n48 GNDA.n47 0.15675
R825 GNDA.n47 GNDA.n21 0.15675
R826 GNDA.n159 GNDA.n21 0.15675
R827 GNDA.n160 GNDA.n159 0.15675
R828 GNDA.n161 GNDA.n160 0.15675
R829 GNDA.n161 GNDA.n18 0.15675
R830 GNDA.n166 GNDA.n18 0.15675
R831 GNDA.n167 GNDA.n166 0.15675
R832 GNDA.n168 GNDA.n167 0.15675
R833 GNDA.n168 GNDA.n15 0.15675
R834 GNDA.n173 GNDA.n15 0.15675
R835 GNDA.n174 GNDA.n173 0.15675
R836 GNDA.n175 GNDA.n174 0.15675
R837 GNDA.n175 GNDA.n12 0.15675
R838 GNDA.n180 GNDA.n12 0.15675
R839 GNDA.n181 GNDA.n180 0.15675
R840 GNDA.n182 GNDA.n181 0.15675
R841 GNDA.n182 GNDA.n10 0.15675
R842 GNDA.n186 GNDA.n10 0.15675
R843 GNDA.n187 GNDA.n186 0.15675
R844 GNDA.n188 GNDA.n187 0.15675
R845 GNDA.n188 GNDA.n6 0.15675
R846 GNDA.n194 GNDA.n6 0.15675
R847 GNDA.n195 GNDA.n194 0.15675
R848 GNDA.n196 GNDA.n195 0.15675
R849 GNDA.n196 GNDA.n4 0.15675
R850 GNDA.n200 GNDA.n4 0.15675
R851 GNDA.n201 GNDA.n200 0.15675
R852 GNDA.n202 GNDA.n201 0.15675
R853 GNDA.n202 GNDA.n1 0.15675
R854 GNDA.n41 GNDA.n40 0.09425
R855 GNDA.n40 GNDA.n39 0.063
R856 DOWN_PFD_b.t1 DOWN_PFD_b.n1 203.528
R857 DOWN_PFD_b.n0 DOWN_PFD_b.t3 203.528
R858 DOWN_PFD_b.n1 DOWN_PFD_b.t0 183.935
R859 DOWN_PFD_b.n0 DOWN_PFD_b.t2 183.935
R860 DOWN_PFD_b.n1 DOWN_PFD_b.n0 83.2005
R861 DOWN_b.n0 DOWN_b.t2 1028.27
R862 DOWN_b.n2 DOWN_b.n1 569.734
R863 DOWN_b.n1 DOWN_b.n0 465.933
R864 DOWN_b.n1 DOWN_b.t3 401.668
R865 DOWN_b.n0 DOWN_b.t4 385.601
R866 DOWN_b.n1 DOWN_b.t5 385.601
R867 DOWN_b.t1 DOWN_b.n2 211.847
R868 DOWN_b.n2 DOWN_b.t0 173.055
R869 DOWN_input.n0 DOWN_input.t1 229.127
R870 DOWN_input.n0 DOWN_input.t0 158.335
R871 DOWN_input.n2 DOWN_input.t2 158.335
R872 DOWN_input.n2 DOWN_input.n0 124.8
R873 DOWN_input DOWN_input.n2 6.4005
R874 DOWN_input.n2 DOWN_input.n1 6.4005
R875 E_b.n0 E_b.t3 517.347
R876 E_b.n2 E_b.n0 417.574
R877 E_b.n2 E_b.n1 244.716
R878 E_b.n0 E_b.t4 228.148
R879 E_b.t1 E_b.n2 221.411
R880 E_b.n1 E_b.t2 24.0005
R881 E_b.n1 E_b.t0 24.0005
R882 a_750_n6120.t0 a_750_n6120.t1 39.4005
R883 E.n4 E.n0 1319.38
R884 E.n0 E.t4 562.333
R885 E.n2 E.t6 388.813
R886 E.n2 E.t5 356.68
R887 E.n3 E.n2 232
R888 E.n0 E.t3 224.934
R889 E.t1 E.n4 221.411
R890 E.n3 E.n1 157.278
R891 E.n4 E.n3 90.64
R892 E.n1 E.t2 24.0005
R893 E.n1 E.t0 24.0005
R894 F_b.n0 F_b.t3 517.347
R895 F_b.n2 F_b.n0 417.574
R896 F_b.n2 F_b.n1 244.716
R897 F_b.n0 F_b.t4 228.148
R898 F_b.t0 F_b.n2 221.411
R899 F_b.n1 F_b.t2 24.0005
R900 F_b.n1 F_b.t1 24.0005
R901 a_750_n6880.t0 a_750_n6880.t1 39.4005
R902 F.n4 F.n0 1319.38
R903 F.n0 F.t3 562.333
R904 F.n2 F.t6 388.813
R905 F.n2 F.t4 356.68
R906 F.n3 F.n2 232
R907 F.n0 F.t5 224.934
R908 F.t0 F.n4 221.411
R909 F.n3 F.n1 157.278
R910 F.n4 F.n3 90.64
R911 F.n1 F.t1 24.0005
R912 F.n1 F.t2 24.0005
R913 QB.t7 QB.t6 835.467
R914 QB.n2 QB.t7 561.913
R915 QB.n3 QB.t5 517.347
R916 QB.n1 QB.t4 514.134
R917 QB.n2 QB.n1 455.5
R918 QB.n4 QB.n3 363.2
R919 QB.n1 QB.t8 273.134
R920 QB.n5 QB.n0 244.716
R921 QB.n3 QB.t3 228.148
R922 QB.t0 QB.n5 221.411
R923 QB.n5 QB.n4 54.3734
R924 QB.n4 QB.n2 32.6567
R925 QB.n0 QB.t2 24.0005
R926 QB.n0 QB.t1 24.0005
R927 QB_b.t5 QB_b.t6 1188.93
R928 QB_b QB_b.n2 899.734
R929 QB_b.t6 QB_b.t4 835.467
R930 QB_b.n2 QB_b.t3 562.333
R931 QB_b QB_b.n1 419.647
R932 QB_b.n1 QB_b.n0 247.917
R933 QB_b.n2 QB_b.t5 224.934
R934 QB_b.n1 QB_b.t1 221.411
R935 QB_b.n0 QB_b.t2 24.0005
R936 QB_b.n0 QB_b.t0 24.0005
R937 QA_b.t3 QA_b.t4 1188.93
R938 QA_b QA_b.n2 837.38
R939 QA_b.t4 QA_b.t6 835.467
R940 QA_b.n0 QA_b.t5 562.333
R941 QA_b QA_b.n0 482
R942 QA_b.n2 QA_b.n1 247.917
R943 QA_b.n0 QA_b.t3 224.934
R944 QA_b.n2 QA_b.t0 221.411
R945 QA_b.n1 QA_b.t1 24.0005
R946 QA_b.n1 QA_b.t2 24.0005
R947 QA.t4 QA.t6 835.467
R948 QA.n2 QA.t8 517.347
R949 QA.n0 QA.t7 465.933
R950 QA.n1 QA.n0 454.062
R951 QA.n1 QA.t4 394.267
R952 QA.n0 QA.t3 321.334
R953 QA.n4 QA.n3 244.715
R954 QA.n2 QA.t5 228.148
R955 QA.n4 QA.t0 221.411
R956 QA.n5 QA.n2 216
R957 QA.n5 QA.n4 201.573
R958 QA QA.n5 60.8005
R959 QA QA.n1 55.9005
R960 QA.n3 QA.t2 24.0005
R961 QA.n3 QA.t1 24.0005
R962 a_2410_n7330.t1 a_2410_n7330.n2 500.086
R963 a_2410_n7330.n0 a_2410_n7330.t3 465.933
R964 a_2410_n7330.t1 a_2410_n7330.n2 461.389
R965 a_2410_n7330.n1 a_2410_n7330.n0 392.586
R966 a_2410_n7330.n0 a_2410_n7330.t2 321.334
R967 a_2410_n7330.n1 a_2410_n7330.t0 177.577
R968 a_2410_n7330.n2 a_2410_n7330.n1 48.3899
R969 a_2080_n7330.t0 a_2080_n7330.n2 500.086
R970 a_2080_n7330.n1 a_2080_n7330.n0 473.334
R971 a_2080_n7330.n0 a_2080_n7330.t2 465.933
R972 a_2080_n7330.t0 a_2080_n7330.n2 461.389
R973 a_2080_n7330.n0 a_2080_n7330.t3 321.334
R974 a_2080_n7330.n1 a_2080_n7330.t1 177.577
R975 a_2080_n7330.n2 a_2080_n7330.n1 48.3898
R976 DOWN.n0 DOWN.t2 605.311
R977 DOWN.t0 DOWN.n0 240.327
R978 DOWN.n0 DOWN.t1 148.736
R979 I_IN I_IN.t1 241.928
R980 I_IN I_IN.t0 158.335
R981 a_370_n6120.t0 a_370_n6120.t1 39.4005
R982 a_1270_n6120.t0 a_1270_n6120.t1 39.4005
R983 a_370_n6880.t0 a_370_n6880.t1 39.4005
R984 a_1270_n6880.t0 a_1270_n6880.t1 39.4005
R985 Reset.n1 Reset.t4 562.333
R986 Reset.n2 Reset.n1 480.45
R987 Reset.n0 Reset.t5 417.733
R988 Reset.n0 Reset.t2 369.534
R989 Reset.n3 Reset.n2 328.733
R990 Reset.t1 Reset.n3 288.37
R991 Reset.n1 Reset.t3 224.934
R992 Reset.n3 Reset.t0 177.577
R993 Reset.n2 Reset.n0 176.733
R994 a_1710_n5500.t0 a_1710_n5500.t1 48.0005
R995 before_Reset.t1 before_Reset.n3 500.086
R996 before_Reset.n1 before_Reset.n0 478.134
R997 before_Reset.n0 before_Reset.t4 465.933
R998 before_Reset.t1 before_Reset.n3 461.389
R999 before_Reset.n2 before_Reset.t2 337.649
R1000 before_Reset.n0 before_Reset.t3 321.334
R1001 before_Reset.n1 before_Reset.t0 187.941
R1002 before_Reset.n3 before_Reset.n2 40.0699
R1003 before_Reset.n2 before_Reset.n1 16.0005
R1004 a_1750_n7330.t0 a_1750_n7330.n2 500.086
R1005 a_1750_n7330.n1 a_1750_n7330.n0 473.334
R1006 a_1750_n7330.n0 a_1750_n7330.t2 465.933
R1007 a_1750_n7330.t0 a_1750_n7330.n2 461.389
R1008 a_1750_n7330.n0 a_1750_n7330.t3 321.334
R1009 a_1750_n7330.n1 a_1750_n7330.t1 177.577
R1010 a_1750_n7330.n2 a_1750_n7330.n1 48.3898
R1011 UP_input.n0 UP_input.t2 241.928
R1012 UP_input.n2 UP_input.t0 241.928
R1013 UP_input.n0 UP_input.t1 145.536
R1014 UP_input.n2 UP_input.n0 124.8
R1015 UP_input UP_input.n2 6.4005
R1016 UP_input.n2 UP_input.n1 6.4005
R1017 a_2150_n6120.t0 a_2150_n6120.n2 500.086
R1018 a_2150_n6120.n1 a_2150_n6120.n0 473.334
R1019 a_2150_n6120.n0 a_2150_n6120.t3 465.933
R1020 a_2150_n6120.t0 a_2150_n6120.n2 461.389
R1021 a_2150_n6120.n0 a_2150_n6120.t2 321.334
R1022 a_2150_n6120.n1 a_2150_n6120.t1 177.577
R1023 a_2150_n6120.n2 a_2150_n6120.n1 48.3899
R1024 opamp_out.t1 opamp_out.t0 400.264
R1025 UP_b.n0 UP_b.t2 778.601
R1026 UP_b.t0 UP_b.n0 209.928
R1027 UP_b.n0 UP_b.t1 177.536
C0 DOWN_input I_IN 0.243956f
C1 I_IN VDDA 0.051398f
C2 UP_input VDDA 0.353708f
C3 DOWN_input VDDA 0.152386f
C4 QA_b VDDA 0.521329f
C5 F_VCO VDDA 0.085127f
C6 QA VDDA 0.542812f
C7 QA_b QA 0.422773f
C8 F_REF VDDA 0.085173f
C9 QA_b F_REF 0.026369f
C10 QB_b VDDA 0.513239f
C11 QA F_REF 0.056f
C12 QB_b F_VCO 0.026369f
C13 DOWN_input GNDA 0.389223f
C14 I_IN GNDA 0.049563f
C15 F_VCO GNDA 0.236218f
C16 UP_input GNDA 0.315799f
C17 F_REF GNDA 0.236218f
C18 VDDA GNDA 19.844099f
C19 QB_b GNDA 1.06416f
C20 QA GNDA 3.0346f
C21 QA_b GNDA 1.05211f
C22 QB.t2 GNDA 0.025496f
C23 QB.t1 GNDA 0.025496f
C24 QB.n0 GNDA 0.136139f
C25 QB.t4 GNDA 0.063104f
C26 QB.t8 GNDA 0.02964f
C27 QB.n1 GNDA 0.091471f
C28 QB.t6 GNDA 0.063104f
C29 QB.t7 GNDA 0.096881f
C30 QB.n2 GNDA 1.18281f
C31 QB.t5 GNDA 0.063727f
C32 QB.t3 GNDA 0.027943f
C33 QB.n3 GNDA 0.160969f
C34 QB.n4 GNDA 0.257153f
C35 QB.n5 GNDA 0.24187f
C36 QB.t0 GNDA 0.134194f
C37 VDDA.t11 GNDA 0.023511f
C38 VDDA.t23 GNDA 0.067921f
C39 VDDA.t21 GNDA 0.082725f
C40 VDDA.n68 GNDA 0.067921f
C41 VDDA.t6 GNDA 0.079242f
C42 VDDA.t13 GNDA 0.089691f
C43 VDDA.n74 GNDA 0.067921f
C44 VDDA.n77 GNDA 0.029108f
C45 VDDA.n83 GNDA 0.021634f
C46 VDDA.n96 GNDA 0.067921f
C47 VDDA.t27 GNDA 0.067921f
C48 VDDA.t39 GNDA 0.023511f
C49 VDDA.n108 GNDA 0.049635f
C50 VDDA.n122 GNDA 0.061826f
C51 VDDA.n144 GNDA 0.033961f
C52 VDDA.n154 GNDA 0.033961f
C53 VDDA.t35 GNDA 0.023511f
C54 VDDA.t19 GNDA 0.023511f
C55 VDDA.n174 GNDA 0.051376f
C56 VDDA.t33 GNDA 0.042668f
C57 VDDA.t18 GNDA 0.090562f
C58 VDDA.t17 GNDA 0.090562f
C59 VDDA.t2 GNDA 0.042668f
C60 VDDA.n198 GNDA 0.047022f
C61 VDDA.t9 GNDA 0.042668f
C62 VDDA.t4 GNDA 0.090562f
C63 VDDA.t5 GNDA 0.090562f
C64 VDDA.t0 GNDA 0.042668f
C65 VDDA.n214 GNDA 0.057472f
C66 VDDA.t14 GNDA 0.046152f
C67 VDDA.t29 GNDA 0.019157f
C68 VDDA.t25 GNDA 0.023511f
C69 VDDA.n222 GNDA 0.033961f
C70 VDDA.n228 GNDA 0.033961f
.ends

