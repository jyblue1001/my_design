* PEX produced on Mon Aug 25 12:40:01 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_opamp_dummy_magic_20.ext - technology: sky130A

.subckt bgr_opamp_dummy_magic_20 VDDA GNDA VOUT+ VOUT- VIN+ VIN-
X0 VDDA.t211 bgr_11_0.1st_Vout_2.t7 bgr_11_0.PFET_GATE_10uA.t8 VDDA.t210 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X1 two_stage_opamp_dummy_magic_29_0.VD4.t31 two_stage_opamp_dummy_magic_29_0.Vb3.t8 VDDA.t53 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t16 two_stage_opamp_dummy_magic_29_0.X.t25 GNDA.t177 VDDA.t106 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X3 VDDA.t168 two_stage_opamp_dummy_magic_29_0.Y.t25 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t10 GNDA.t121 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X4 GNDA.t65 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t12 two_stage_opamp_dummy_magic_29_0.V_source.t39 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X5 GNDA.t276 GNDA.t274 two_stage_opamp_dummy_magic_29_0.Vb2.t9 GNDA.t275 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X6 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t12 two_stage_opamp_dummy_magic_29_0.X.t26 VDDA.t51 GNDA.t176 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X7 GNDA.t4 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t13 two_stage_opamp_dummy_magic_29_0.V_source.t38 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X8 VOUT-.t19 two_stage_opamp_dummy_magic_29_0.cap_res_X.t142 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 VOUT-.t20 two_stage_opamp_dummy_magic_29_0.cap_res_X.t141 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X10 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t3 two_stage_opamp_dummy_magic_29_0.Y.t0 GNDA.t16 sky130_fd_pr__res_high_po_1p41 l=1.41
X11 VOUT+.t19 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X12 two_stage_opamp_dummy_magic_29_0.VD4.t37 two_stage_opamp_dummy_magic_29_0.VD4.t35 two_stage_opamp_dummy_magic_29_0.Y.t21 two_stage_opamp_dummy_magic_29_0.VD4.t36 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X13 VDDA.t366 VDDA.t364 VOUT-.t6 VDDA.t365 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X14 VDDA.t140 bgr_11_0.V_TOP.t14 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t3 VDDA.t139 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X15 two_stage_opamp_dummy_magic_29_0.VD2.t17 two_stage_opamp_dummy_magic_29_0.Vb1.t12 two_stage_opamp_dummy_magic_29_0.Y.t16 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X16 VOUT-.t21 two_stage_opamp_dummy_magic_29_0.cap_res_X.t140 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X17 VOUT+.t20 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X18 bgr_11_0.1st_Vout_1.t7 bgr_11_0.cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X19 two_stage_opamp_dummy_magic_29_0.VD3.t19 two_stage_opamp_dummy_magic_29_0.Vb2.t11 two_stage_opamp_dummy_magic_29_0.X.t8 two_stage_opamp_dummy_magic_29_0.VD3.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X20 two_stage_opamp_dummy_magic_29_0.Vb2.t1 bgr_11_0.NFET_GATE_10uA.t5 GNDA.t37 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X21 bgr_11_0.V_TOP.t15 VDDA.t141 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 GNDA.t71 bgr_11_0.NFET_GATE_10uA.t6 two_stage_opamp_dummy_magic_29_0.Vb2.t2 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X23 two_stage_opamp_dummy_magic_29_0.VD4.t30 two_stage_opamp_dummy_magic_29_0.Vb3.t9 VDDA.t55 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X24 VDDA.t363 VDDA.t360 VDDA.t362 VDDA.t361 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0 ps=0 w=1.8 l=0.2
X25 bgr_11_0.START_UP_NFET1.t0 bgr_11_0.START_UP_NFET1 GNDA.t15 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X26 bgr_11_0.1st_Vout_1.t6 bgr_11_0.V_mir1.t13 VDDA.t414 VDDA.t413 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X27 two_stage_opamp_dummy_magic_29_0.VD3.t21 VDDA.t357 VDDA.t359 VDDA.t358 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X28 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t9 two_stage_opamp_dummy_magic_29_0.Y.t26 GNDA.t69 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X29 VOUT+.t21 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 a_3230_6968.t1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t10 GNDA.t135 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X31 VOUT-.t22 two_stage_opamp_dummy_magic_29_0.cap_res_X.t139 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 two_stage_opamp_dummy_magic_29_0.VD2.t3 VIN+.t0 two_stage_opamp_dummy_magic_29_0.V_source.t7 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X33 VOUT-.t23 two_stage_opamp_dummy_magic_29_0.cap_res_X.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 bgr_11_0.V_TOP.t16 VDDA.t387 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X35 two_stage_opamp_dummy_magic_29_0.V_source.t37 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t14 GNDA.t6 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X36 VOUT+.t22 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t140 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X37 VDDA.t118 two_stage_opamp_dummy_magic_29_0.Y.t27 VOUT+.t10 VDDA.t117 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X38 VOUT-.t24 two_stage_opamp_dummy_magic_29_0.cap_res_X.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 GNDA.t273 GNDA.t272 two_stage_opamp_dummy_magic_29_0.Vb1.t11 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X40 two_stage_opamp_dummy_magic_29_0.VD3.t17 two_stage_opamp_dummy_magic_29_0.Vb2.t12 two_stage_opamp_dummy_magic_29_0.X.t6 two_stage_opamp_dummy_magic_29_0.VD3.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X41 VOUT+.t23 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t141 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X42 VOUT+.t24 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X43 a_6350_30238.t0 bgr_11_0.Vin+.t5 GNDA.t84 sky130_fd_pr__res_xhigh_po_0p35 l=6
X44 bgr_11_0.V_TOP.t17 VDDA.t388 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 two_stage_opamp_dummy_magic_29_0.V_err_gate.t2 bgr_11_0.NFET_GATE_10uA.t7 GNDA.t291 GNDA.t290 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X46 VOUT-.t25 two_stage_opamp_dummy_magic_29_0.cap_res_X.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 VDDA.t171 a_6540_22450.t11 a_6540_22450.t12 VDDA.t170 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X48 two_stage_opamp_dummy_magic_29_0.VD3.t31 two_stage_opamp_dummy_magic_29_0.Vb3.t10 VDDA.t90 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X49 VDDA.t385 bgr_11_0.V_mir1.t10 bgr_11_0.V_mir1.t11 VDDA.t384 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X50 VOUT-.t26 two_stage_opamp_dummy_magic_29_0.cap_res_X.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 two_stage_opamp_dummy_magic_29_0.err_amp_out.t1 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t5 GNDA.t126 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X52 GNDA.t271 GNDA.t269 VOUT-.t18 GNDA.t270 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X53 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t14 bgr_11_0.PFET_GATE_10uA.t10 VDDA.t249 VDDA.t248 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X54 GNDA.t68 two_stage_opamp_dummy_magic_29_0.Y.t28 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t8 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X55 VDDA.t247 bgr_11_0.PFET_GATE_10uA.t11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t13 VDDA.t246 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X56 two_stage_opamp_dummy_magic_29_0.VD4.t21 VDDA.t354 VDDA.t356 VDDA.t355 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X57 VOUT-.t27 two_stage_opamp_dummy_magic_29_0.cap_res_X.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X58 bgr_11_0.V_TOP.t18 VDDA.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 bgr_11_0.cap_res1.t0 bgr_11_0.V_TOP.t0 GNDA.t13 sky130_fd_pr__res_high_po_0p35 l=2.05
X60 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t15 two_stage_opamp_dummy_magic_29_0.X.t27 GNDA.t175 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X61 VOUT+.t25 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X62 two_stage_opamp_dummy_magic_29_0.V_source.t5 two_stage_opamp_dummy_magic_29_0.Vb1.t13 two_stage_opamp_dummy_magic_29_0.Vb1_2.t0 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.6 ps=3.8 w=1.5 l=3
X63 VOUT-.t28 two_stage_opamp_dummy_magic_29_0.cap_res_X.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X64 two_stage_opamp_dummy_magic_29_0.VD1.t11 two_stage_opamp_dummy_magic_29_0.Vb1.t14 two_stage_opamp_dummy_magic_29_0.X.t13 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X65 VOUT+.t26 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X66 GNDA.t57 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t15 two_stage_opamp_dummy_magic_29_0.V_source.t36 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X67 VOUT-.t29 two_stage_opamp_dummy_magic_29_0.cap_res_X.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X68 VOUT-.t30 two_stage_opamp_dummy_magic_29_0.cap_res_X.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X69 VOUT+.t27 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X70 VDDA.t85 two_stage_opamp_dummy_magic_29_0.X.t28 VOUT-.t16 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X71 bgr_11_0.V_TOP.t19 VDDA.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X72 bgr_11_0.1st_Vout_2.t8 bgr_11_0.cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X73 VDDA.t373 two_stage_opamp_dummy_magic_29_0.X.t29 VOUT-.t15 VDDA.t372 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X74 two_stage_opamp_dummy_magic_29_0.VD2.t16 two_stage_opamp_dummy_magic_29_0.Vb1.t15 two_stage_opamp_dummy_magic_29_0.Y.t15 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X75 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t1 a_3830_3166.t1 GNDA.t284 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X76 GNDA.t186 GNDA.t258 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X77 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t9 VDDA.t351 VDDA.t353 VDDA.t352 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X78 VOUT-.t31 two_stage_opamp_dummy_magic_29_0.cap_res_X.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X79 two_stage_opamp_dummy_magic_29_0.VD1.t10 two_stage_opamp_dummy_magic_29_0.Vb1.t16 two_stage_opamp_dummy_magic_29_0.X.t11 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X80 VOUT-.t32 two_stage_opamp_dummy_magic_29_0.cap_res_X.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X81 VDDA.t209 bgr_11_0.1st_Vout_2.t9 bgr_11_0.PFET_GATE_10uA.t7 VDDA.t208 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X82 two_stage_opamp_dummy_magic_29_0.VD1.t1 VIN-.t0 two_stage_opamp_dummy_magic_29_0.V_source.t4 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X83 VOUT-.t33 two_stage_opamp_dummy_magic_29_0.cap_res_X.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X84 VOUT+.t28 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t138 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X85 bgr_11_0.1st_Vout_2.t10 bgr_11_0.cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X86 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t9 bgr_11_0.PFET_GATE_10uA.t12 VDDA.t245 VDDA.t244 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X87 VOUT-.t34 two_stage_opamp_dummy_magic_29_0.cap_res_X.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 VOUT-.t35 two_stage_opamp_dummy_magic_29_0.cap_res_X.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X89 VOUT+.t29 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t139 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X90 two_stage_opamp_dummy_magic_29_0.VD3.t15 two_stage_opamp_dummy_magic_29_0.Vb2.t13 two_stage_opamp_dummy_magic_29_0.X.t7 two_stage_opamp_dummy_magic_29_0.VD3.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 bgr_11_0.Vin+.t0 GNDA.t42 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X92 two_stage_opamp_dummy_magic_29_0.VD2.t20 GNDA.t267 GNDA.t268 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X93 VOUT-.t36 two_stage_opamp_dummy_magic_29_0.cap_res_X.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X94 bgr_11_0.1st_Vout_1.t8 bgr_11_0.cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 GNDA.t266 GNDA.t265 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t11 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X96 two_stage_opamp_dummy_magic_29_0.VD1.t0 VIN-.t1 two_stage_opamp_dummy_magic_29_0.V_source.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X97 bgr_11_0.1st_Vout_2.t11 bgr_11_0.cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 two_stage_opamp_dummy_magic_29_0.VD4.t11 two_stage_opamp_dummy_magic_29_0.Vb2.t14 two_stage_opamp_dummy_magic_29_0.Y.t9 two_stage_opamp_dummy_magic_29_0.VD4.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X99 VDDA.t115 two_stage_opamp_dummy_magic_29_0.Y.t29 VOUT+.t9 VDDA.t114 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X100 VOUT-.t37 two_stage_opamp_dummy_magic_29_0.cap_res_X.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 two_stage_opamp_dummy_magic_29_0.Vb1_2.t4 two_stage_opamp_dummy_magic_29_0.Vb1.t4 two_stage_opamp_dummy_magic_29_0.Vb1.t5 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X102 VDDA.t8 two_stage_opamp_dummy_magic_29_0.Y.t30 VOUT+.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X103 bgr_11_0.V_TOP.t20 VDDA.t159 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 VDDA.t243 bgr_11_0.PFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t4 VDDA.t242 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X105 VOUT+.t30 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X106 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t6 VDDA.t348 VDDA.t350 VDDA.t349 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X107 VOUT+.t31 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X108 VDDA.t193 a_6540_22450.t13 bgr_11_0.1st_Vout_2.t3 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X109 VDDA.t161 bgr_11_0.V_TOP.t21 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t2 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X110 VOUT+.t32 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X111 VOUT-.t38 two_stage_opamp_dummy_magic_29_0.cap_res_X.t123 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X112 VOUT-.t39 two_stage_opamp_dummy_magic_29_0.cap_res_X.t122 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X113 VOUT-.t40 two_stage_opamp_dummy_magic_29_0.cap_res_X.t121 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X114 VOUT-.t41 two_stage_opamp_dummy_magic_29_0.cap_res_X.t120 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 VDDA.t9 two_stage_opamp_dummy_magic_29_0.Y.t31 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t9 GNDA.t12 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X116 VOUT-.t42 two_stage_opamp_dummy_magic_29_0.cap_res_X.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X117 VOUT-.t17 GNDA.t262 GNDA.t264 GNDA.t263 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X118 two_stage_opamp_dummy_magic_29_0.VD4.t13 two_stage_opamp_dummy_magic_29_0.Vb2.t15 two_stage_opamp_dummy_magic_29_0.Y.t10 two_stage_opamp_dummy_magic_29_0.VD4.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X119 VOUT+.t33 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X120 VOUT+.t34 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X121 two_stage_opamp_dummy_magic_29_0.VD1.t9 two_stage_opamp_dummy_magic_29_0.Vb1.t17 two_stage_opamp_dummy_magic_29_0.X.t15 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X122 bgr_11_0.1st_Vout_2.t12 bgr_11_0.cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X123 VOUT+.t35 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t119 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X124 GNDA.t58 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t16 two_stage_opamp_dummy_magic_29_0.V_source.t35 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X125 bgr_11_0.V_TOP.t22 VDDA.t418 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X126 VOUT-.t43 two_stage_opamp_dummy_magic_29_0.cap_res_X.t118 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X127 VOUT+.t36 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X128 VDDA.t155 two_stage_opamp_dummy_magic_29_0.X.t30 VOUT-.t14 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X129 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t5 VDDA.t345 VDDA.t347 VDDA.t346 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X130 VOUT-.t44 two_stage_opamp_dummy_magic_29_0.cap_res_X.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X131 VOUT+.t37 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X132 two_stage_opamp_dummy_magic_29_0.VD2.t15 two_stage_opamp_dummy_magic_29_0.Vb1.t18 two_stage_opamp_dummy_magic_29_0.Y.t11 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X133 VOUT-.t45 two_stage_opamp_dummy_magic_29_0.cap_res_X.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X134 two_stage_opamp_dummy_magic_29_0.VD1.t8 two_stage_opamp_dummy_magic_29_0.Vb1.t19 two_stage_opamp_dummy_magic_29_0.X.t5 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X135 VOUT-.t46 two_stage_opamp_dummy_magic_29_0.cap_res_X.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X136 VOUT-.t3 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t2 GNDA.t128 GNDA.t127 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X137 GNDA.t261 GNDA.t259 GNDA.t261 GNDA.t260 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0 ps=0 w=2.5 l=0.15
X138 GNDA.t278 bgr_11_0.NFET_GATE_10uA.t8 two_stage_opamp_dummy_magic_29_0.Vb3.t6 GNDA.t277 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X139 VOUT-.t47 two_stage_opamp_dummy_magic_29_0.cap_res_X.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X140 VDDA.t390 a_6540_22450.t9 a_6540_22450.t10 VDDA.t389 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X141 a_3110_6968.t1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t11 GNDA.t75 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X142 VOUT+.t38 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X143 bgr_11_0.START_UP.t3 bgr_11_0.V_TOP.t23 VDDA.t420 VDDA.t419 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X144 VOUT+.t39 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 two_stage_opamp_dummy_magic_29_0.VD1.t20 VIN-.t2 two_stage_opamp_dummy_magic_29_0.V_source.t20 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X146 VOUT+.t40 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X147 a_11420_30238.t1 bgr_11_0.Vin-.t6 GNDA.t92 sky130_fd_pr__res_xhigh_po_0p35 l=6
X148 bgr_11_0.V_TOP.t12 VDDA.t342 VDDA.t344 VDDA.t343 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.45 ps=2.9 w=1 l=0.15
X149 GNDA.t91 a_11950_28880.t1 GNDA.t90 sky130_fd_pr__res_xhigh_po_0p35 l=4
X150 two_stage_opamp_dummy_magic_29_0.VD3.t13 two_stage_opamp_dummy_magic_29_0.Vb2.t16 two_stage_opamp_dummy_magic_29_0.X.t21 two_stage_opamp_dummy_magic_29_0.VD3.t12 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X151 bgr_11_0.V_TOP.t24 VDDA.t369 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 VDDA.t0 two_stage_opamp_dummy_magic_29_0.X.t31 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t11 GNDA.t174 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X153 VOUT-.t48 two_stage_opamp_dummy_magic_29_0.cap_res_X.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X154 VOUT+.t41 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X155 VOUT+.t42 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X156 bgr_11_0.Vin+.t4 bgr_11_0.V_TOP.t25 VDDA.t371 VDDA.t370 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X157 VDDA.t341 VDDA.t339 two_stage_opamp_dummy_magic_29_0.Vb2_2.t3 VDDA.t340 sky130_fd_pr__pfet_01v8 ad=0.72 pd=4.4 as=0.36 ps=2.2 w=1.8 l=0.2
X158 two_stage_opamp_dummy_magic_29_0.VD4.t19 two_stage_opamp_dummy_magic_29_0.Vb2.t17 two_stage_opamp_dummy_magic_29_0.Y.t19 two_stage_opamp_dummy_magic_29_0.VD4.t18 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X159 two_stage_opamp_dummy_magic_29_0.VD1.t18 VIN-.t3 two_stage_opamp_dummy_magic_29_0.V_source.t18 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X160 VOUT-.t49 two_stage_opamp_dummy_magic_29_0.cap_res_X.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X161 VDDA.t173 bgr_11_0.V_mir1.t14 bgr_11_0.1st_Vout_1.t5 VDDA.t172 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X162 two_stage_opamp_dummy_magic_29_0.V_err_gate.t4 VDDA.t336 VDDA.t338 VDDA.t337 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X163 VDDA.t65 two_stage_opamp_dummy_magic_29_0.Y.t32 VOUT+.t7 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X164 VOUT-.t50 two_stage_opamp_dummy_magic_29_0.cap_res_X.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X165 VOUT+.t43 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 two_stage_opamp_dummy_magic_29_0.V_err_gate.t5 two_stage_opamp_dummy_magic_29_0.V_tot.t4 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t1 VDDA.t407 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X167 VOUT-.t51 two_stage_opamp_dummy_magic_29_0.cap_res_X.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X168 VOUT-.t52 two_stage_opamp_dummy_magic_29_0.cap_res_X.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X169 VOUT-.t53 two_stage_opamp_dummy_magic_29_0.cap_res_X.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X170 VOUT+.t44 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X171 bgr_11_0.1st_Vout_2.t13 bgr_11_0.cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 VDDA.t335 VDDA.t332 VDDA.t334 VDDA.t333 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.15
X173 VDDA.t331 VDDA.t328 VDDA.t330 VDDA.t329 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X174 two_stage_opamp_dummy_magic_29_0.V_err_p.t3 two_stage_opamp_dummy_magic_29_0.V_err_gate.t6 VDDA.t189 VDDA.t188 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X175 VOUT+.t45 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X176 VOUT+.t46 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t126 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X177 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t3 VDDA.t325 VDDA.t327 VDDA.t326 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X178 VOUT+.t47 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X179 VOUT-.t54 two_stage_opamp_dummy_magic_29_0.cap_res_X.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X180 VDDA.t241 bgr_11_0.PFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t8 VDDA.t240 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X181 GNDA.t257 GNDA.t256 two_stage_opamp_dummy_magic_29_0.VD1.t15 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X182 VOUT+.t48 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X183 GNDA.t50 two_stage_opamp_dummy_magic_29_0.Y.t33 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t7 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X184 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t14 bgr_11_0.NFET_GATE_10uA.t9 GNDA.t289 GNDA.t288 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X185 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t6 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t4 two_stage_opamp_dummy_magic_29_0.Vb3.t7 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t5 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X186 VDDA.t410 two_stage_opamp_dummy_magic_29_0.Y.t34 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t8 GNDA.t285 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X187 VOUT-.t55 two_stage_opamp_dummy_magic_29_0.cap_res_X.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X188 two_stage_opamp_dummy_magic_29_0.Vb2.t10 bgr_11_0.NFET_GATE_10uA.t10 GNDA.t287 GNDA.t286 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X189 VDDA.t402 bgr_11_0.V_TOP.t26 bgr_11_0.Vin-.t3 VDDA.t401 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X190 VOUT+.t49 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X191 GNDA.t101 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t17 two_stage_opamp_dummy_magic_29_0.V_p_mir.t2 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X192 VDDA.t324 VDDA.t322 bgr_11_0.V_TOP.t11 VDDA.t323 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X193 VDDA.t321 VDDA.t319 two_stage_opamp_dummy_magic_29_0.VD3.t20 VDDA.t320 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X194 GNDA.t255 GNDA.t254 two_stage_opamp_dummy_magic_29_0.VD2.t19 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X195 VOUT-.t56 two_stage_opamp_dummy_magic_29_0.cap_res_X.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X196 GNDA.t186 GNDA.t243 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X197 GNDA.t102 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t18 two_stage_opamp_dummy_magic_29_0.V_source.t34 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X198 VOUT+.t12 a_3830_3166.t0 GNDA.t82 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X199 VOUT+.t50 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X200 two_stage_opamp_dummy_magic_29_0.VD4.t29 two_stage_opamp_dummy_magic_29_0.Vb3.t11 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X201 VOUT-.t57 two_stage_opamp_dummy_magic_29_0.cap_res_X.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 VOUT-.t58 two_stage_opamp_dummy_magic_29_0.cap_res_X.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X203 VDDA.t105 two_stage_opamp_dummy_magic_29_0.X.t32 VOUT-.t13 VDDA.t104 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X204 bgr_11_0.1st_Vout_1.t9 bgr_11_0.cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X205 VOUT+.t51 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X206 GNDA.t218 GNDA.t242 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X207 VDDA.t137 bgr_11_0.1st_Vout_1.t10 bgr_11_0.V_TOP.t3 VDDA.t136 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X208 VOUT+.t52 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 bgr_11_0.START_UP.t5 bgr_11_0.START_UP.t4 bgr_11_0.START_UP_NFET1.t0 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X210 VOUT+.t53 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X211 GNDA.t64 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t0 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t1 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X212 two_stage_opamp_dummy_magic_29_0.VD1.t7 two_stage_opamp_dummy_magic_29_0.Vb1.t20 two_stage_opamp_dummy_magic_29_0.X.t14 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X213 VOUT-.t59 two_stage_opamp_dummy_magic_29_0.cap_res_X.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X214 two_stage_opamp_dummy_magic_29_0.V_source.t3 two_stage_opamp_dummy_magic_29_0.err_amp_out.t4 GNDA.t40 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X215 bgr_11_0.NFET_GATE_10uA.t1 bgr_11_0.NFET_GATE_10uA.t0 GNDA.t104 GNDA.t103 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X216 VOUT+.t54 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 VDDA.t404 bgr_11_0.V_TOP.t27 bgr_11_0.Vin+.t3 VDDA.t403 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X218 VOUT+.t55 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 VOUT+.t56 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 GNDA.t173 two_stage_opamp_dummy_magic_29_0.X.t33 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t14 VDDA.t156 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X221 bgr_11_0.1st_Vout_1.t11 bgr_11_0.cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 VOUT-.t60 two_stage_opamp_dummy_magic_29_0.cap_res_X.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X223 VDDA.t367 two_stage_opamp_dummy_magic_29_0.X.t34 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t10 GNDA.t172 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X224 VDDA.t318 VDDA.t316 two_stage_opamp_dummy_magic_29_0.VD4.t20 VDDA.t317 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X225 two_stage_opamp_dummy_magic_29_0.X.t22 two_stage_opamp_dummy_magic_29_0.Vb1.t21 two_stage_opamp_dummy_magic_29_0.VD1.t6 GNDA.t178 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X226 VOUT+.t57 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X227 VOUT+.t58 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X228 VDDA.t386 two_stage_opamp_dummy_magic_29_0.X.t35 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t9 GNDA.t171 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X229 VOUT-.t61 two_stage_opamp_dummy_magic_29_0.cap_res_X.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X230 bgr_11_0.V_TOP.t28 VDDA.t415 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X231 VOUT+.t59 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X232 GNDA.t186 GNDA.t251 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X233 VDDA.t181 bgr_11_0.V_mir1.t8 bgr_11_0.V_mir1.t9 VDDA.t180 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X234 two_stage_opamp_dummy_magic_29_0.VD1.t14 GNDA.t252 GNDA.t253 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X235 GNDA.t250 GNDA.t247 GNDA.t249 GNDA.t248 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X236 VDDA.t315 VDDA.t313 bgr_11_0.NFET_GATE_10uA.t3 VDDA.t314 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X237 bgr_11_0.1st_Vout_1.t12 bgr_11_0.cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X238 VDDA.t412 two_stage_opamp_dummy_magic_29_0.Y.t35 VOUT+.t6 VDDA.t411 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X239 VOUT+.t60 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X240 VOUT+.t61 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X241 VOUT+.t62 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X242 VOUT+.t63 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X243 two_stage_opamp_dummy_magic_29_0.Y.t24 two_stage_opamp_dummy_magic_29_0.Vb1.t22 two_stage_opamp_dummy_magic_29_0.VD2.t14 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X244 VDDA.t177 bgr_11_0.1st_Vout_1.t13 bgr_11_0.V_TOP.t7 VDDA.t176 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X245 bgr_11_0.Vin+.t2 bgr_11_0.V_TOP.t29 VDDA.t417 VDDA.t416 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X246 GNDA.t72 two_stage_opamp_dummy_magic_29_0.Y.t36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t6 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X247 VOUT-.t62 two_stage_opamp_dummy_magic_29_0.cap_res_X.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X248 VDDA.t368 GNDA.t244 GNDA.t246 GNDA.t245 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X249 bgr_11_0.V_TOP.t30 VDDA.t152 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X250 bgr_11_0.PFET_GATE_10uA.t6 bgr_11_0.1st_Vout_2.t14 VDDA.t207 VDDA.t206 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X251 VDDA.t2 two_stage_opamp_dummy_magic_29_0.Vb3.t12 two_stage_opamp_dummy_magic_29_0.VD3.t30 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X252 VDDA.t126 two_stage_opamp_dummy_magic_29_0.Y.t37 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t7 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X253 VOUT+.t64 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X254 GNDA.t241 GNDA.t238 GNDA.t240 GNDA.t239 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0 ps=0 w=2.5 l=0.15
X255 VOUT-.t63 two_stage_opamp_dummy_magic_29_0.cap_res_X.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X256 two_stage_opamp_dummy_magic_29_0.Vb2.t6 bgr_11_0.NFET_GATE_10uA.t11 GNDA.t96 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X257 two_stage_opamp_dummy_magic_29_0.V_source.t40 VIN+.t1 two_stage_opamp_dummy_magic_29_0.VD2.t21 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X258 VOUT-.t64 two_stage_opamp_dummy_magic_29_0.cap_res_X.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X259 VOUT+.t65 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t97 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X260 GNDA.t48 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t19 two_stage_opamp_dummy_magic_29_0.V_source.t33 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X261 bgr_11_0.1st_Vout_1.t14 bgr_11_0.cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X262 two_stage_opamp_dummy_magic_29_0.Vb1.t3 two_stage_opamp_dummy_magic_29_0.Vb1.t2 two_stage_opamp_dummy_magic_29_0.Vb1_2.t3 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X263 VOUT-.t65 two_stage_opamp_dummy_magic_29_0.cap_res_X.t96 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X264 VDDA.t396 bgr_11_0.V_mir1.t6 bgr_11_0.V_mir1.t7 VDDA.t395 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X265 VOUT+.t11 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t3 GNDA.t81 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X266 VOUT+.t5 two_stage_opamp_dummy_magic_29_0.Y.t38 VDDA.t87 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X267 bgr_11_0.V_TOP.t31 VDDA.t153 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X268 VOUT-.t66 two_stage_opamp_dummy_magic_29_0.cap_res_X.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X269 VDDA.t102 two_stage_opamp_dummy_magic_29_0.X.t36 VOUT-.t12 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X270 VDDA.t205 bgr_11_0.1st_Vout_2.t15 bgr_11_0.PFET_GATE_10uA.t5 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X271 GNDA.t20 a_11300_28630.t0 GNDA.t19 sky130_fd_pr__res_xhigh_po_0p35 l=6
X272 GNDA.t94 bgr_11_0.NFET_GATE_10uA.t12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t12 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X273 two_stage_opamp_dummy_magic_29_0.Vb2.t8 GNDA.t235 GNDA.t237 GNDA.t236 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X274 two_stage_opamp_dummy_magic_29_0.Vb2_2.t2 two_stage_opamp_dummy_magic_29_0.Vb2.t4 two_stage_opamp_dummy_magic_29_0.Vb2.t5 two_stage_opamp_dummy_magic_29_0.Vb2_2.t1 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X275 GNDA.t170 two_stage_opamp_dummy_magic_29_0.X.t37 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t13 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X276 VOUT-.t67 two_stage_opamp_dummy_magic_29_0.cap_res_X.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X277 bgr_11_0.1st_Vout_2.t16 bgr_11_0.cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X278 bgr_11_0.V_TOP.t32 VDDA.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X279 GNDA.t169 two_stage_opamp_dummy_magic_29_0.X.t38 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t12 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X280 VOUT+.t66 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t116 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X281 VDDA.t73 two_stage_opamp_dummy_magic_29_0.X.t39 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t8 GNDA.t168 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X282 VOUT+.t67 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t117 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X283 bgr_11_0.V_p_1.t2 bgr_11_0.Vin+.t6 bgr_11_0.1st_Vout_1.t3 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X284 VOUT+.t68 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t136 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X285 VDDA.t383 a_6540_22450.t14 bgr_11_0.1st_Vout_2.t4 VDDA.t382 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X286 bgr_11_0.1st_Vout_1.t15 bgr_11_0.cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X287 VOUT+.t69 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t137 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X288 two_stage_opamp_dummy_magic_29_0.Y.t5 two_stage_opamp_dummy_magic_29_0.Vb1.t23 two_stage_opamp_dummy_magic_29_0.VD2.t13 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X289 VOUT-.t68 two_stage_opamp_dummy_magic_29_0.cap_res_X.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X290 bgr_11_0.1st_Vout_2.t17 bgr_11_0.cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X291 two_stage_opamp_dummy_magic_29_0.X.t20 two_stage_opamp_dummy_magic_29_0.Vb2.t18 two_stage_opamp_dummy_magic_29_0.VD3.t11 two_stage_opamp_dummy_magic_29_0.VD3.t10 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X292 two_stage_opamp_dummy_magic_29_0.Y.t8 two_stage_opamp_dummy_magic_29_0.Vb1.t24 two_stage_opamp_dummy_magic_29_0.VD2.t12 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X293 GNDA.t234 GNDA.t231 GNDA.t233 GNDA.t232 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0 ps=0 w=1 l=0.15
X294 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t3 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t0 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t2 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t1 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0 ps=0 w=3.5 l=0.2
X295 VOUT-.t69 two_stage_opamp_dummy_magic_29_0.cap_res_X.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X296 two_stage_opamp_dummy_magic_29_0.VD4.t17 two_stage_opamp_dummy_magic_29_0.Vb2.t19 two_stage_opamp_dummy_magic_29_0.Y.t18 two_stage_opamp_dummy_magic_29_0.VD4.t16 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X297 VOUT-.t70 two_stage_opamp_dummy_magic_29_0.cap_res_X.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X298 VOUT-.t71 two_stage_opamp_dummy_magic_29_0.cap_res_X.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X299 VOUT+.t70 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X300 bgr_11_0.1st_Vout_1.t16 bgr_11_0.cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X301 a_5700_30088.t0 a_5820_28824.t0 GNDA.t2 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X302 VDDA.t61 two_stage_opamp_dummy_magic_29_0.Vb3.t13 two_stage_opamp_dummy_magic_29_0.VD3.t29 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X303 VOUT-.t72 two_stage_opamp_dummy_magic_29_0.cap_res_X.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X304 VOUT-.t73 two_stage_opamp_dummy_magic_29_0.cap_res_X.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X305 bgr_11_0.1st_Vout_2.t18 bgr_11_0.cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X306 VDDA.t239 bgr_11_0.PFET_GATE_10uA.t15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t12 VDDA.t238 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X307 GNDA.t151 VDDA.t310 VDDA.t312 VDDA.t311 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X308 VOUT+.t71 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X309 VOUT-.t74 two_stage_opamp_dummy_magic_29_0.cap_res_X.t87 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X310 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t16 VDDA.t307 VDDA.t309 VDDA.t308 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X311 GNDA.t60 two_stage_opamp_dummy_magic_29_0.Y.t39 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t5 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X312 VOUT-.t75 two_stage_opamp_dummy_magic_29_0.cap_res_X.t86 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X313 a_6540_22450.t8 a_6540_22450.t7 VDDA.t13 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X314 VDDA.t381 two_stage_opamp_dummy_magic_29_0.Vb3.t14 two_stage_opamp_dummy_magic_29_0.VD4.t28 VDDA.t380 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X315 VDDA.t74 two_stage_opamp_dummy_magic_29_0.Y.t40 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t6 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X316 bgr_11_0.1st_Vout_1.t17 bgr_11_0.cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X317 two_stage_opamp_dummy_magic_29_0.V_source.t9 VIN+.t2 two_stage_opamp_dummy_magic_29_0.VD2.t5 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X318 bgr_11_0.1st_Vout_2.t19 bgr_11_0.cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X319 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t10 GNDA.t229 GNDA.t230 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X320 GNDA.t49 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t20 two_stage_opamp_dummy_magic_29_0.V_source.t32 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X321 VOUT+.t72 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X322 GNDA.t186 GNDA.t228 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X323 VOUT+.t73 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X324 VOUT-.t76 two_stage_opamp_dummy_magic_29_0.cap_res_X.t85 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X325 VOUT-.t77 two_stage_opamp_dummy_magic_29_0.cap_res_X.t84 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X326 VOUT-.t78 two_stage_opamp_dummy_magic_29_0.cap_res_X.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X327 bgr_11_0.1st_Vout_2.t20 bgr_11_0.cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X328 VOUT+.t74 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X329 VOUT+.t75 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X330 VOUT-.t79 two_stage_opamp_dummy_magic_29_0.cap_res_X.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X331 VOUT-.t80 two_stage_opamp_dummy_magic_29_0.cap_res_X.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X332 VDDA.t92 two_stage_opamp_dummy_magic_29_0.Vb3.t15 two_stage_opamp_dummy_magic_29_0.VD4.t27 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X333 bgr_11_0.START_UP.t2 bgr_11_0.V_TOP.t33 VDDA.t131 VDDA.t130 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X334 GNDA.t167 two_stage_opamp_dummy_magic_29_0.X.t40 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t11 VDDA.t186 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X335 VDDA.t306 VDDA.t304 VDDA.t306 VDDA.t305 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0 ps=0 w=1 l=0.15
X336 VOUT+.t76 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t114 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X337 bgr_11_0.1st_Vout_1.t18 bgr_11_0.cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X338 VDDA.t80 bgr_11_0.V_mir1.t15 bgr_11_0.1st_Vout_1.t2 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X339 VDDA.t237 bgr_11_0.PFET_GATE_10uA.t16 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t7 VDDA.t236 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X340 two_stage_opamp_dummy_magic_29_0.Vb2_2.t0 two_stage_opamp_dummy_magic_29_0.Vb2.t20 VDDA.t195 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.36 pd=2.2 as=0.36 ps=2.2 w=1.8 l=0.2
X341 VDDA.t94 two_stage_opamp_dummy_magic_29_0.Vb3.t16 two_stage_opamp_dummy_magic_29_0.VD3.t28 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X342 GNDA.t227 GNDA.t225 VDDA.t81 GNDA.t226 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X343 bgr_11_0.cap_res2.t0 bgr_11_0.PFET_GATE_10uA.t0 GNDA.t18 sky130_fd_pr__res_high_po_0p35 l=2.05
X344 bgr_11_0.V_TOP.t34 VDDA.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X345 VOUT-.t0 a_13940_3166.t0 GNDA.t9 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X346 two_stage_opamp_dummy_magic_29_0.V_source.t31 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t21 GNDA.t44 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X347 VDDA.t107 two_stage_opamp_dummy_magic_29_0.X.t41 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t7 GNDA.t166 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X348 GNDA.t137 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t4 VOUT+.t13 GNDA.t136 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X349 VOUT-.t81 two_stage_opamp_dummy_magic_29_0.cap_res_X.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X350 two_stage_opamp_dummy_magic_29_0.V_source.t30 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t22 GNDA.t45 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X351 VOUT+.t77 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t115 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X352 GNDA.t186 GNDA.t224 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X353 VOUT+.t78 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X354 two_stage_opamp_dummy_magic_29_0.Y.t14 two_stage_opamp_dummy_magic_29_0.Vb1.t25 two_stage_opamp_dummy_magic_29_0.VD2.t11 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X355 VOUT-.t82 two_stage_opamp_dummy_magic_29_0.cap_res_X.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X356 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t3 bgr_11_0.PFET_GATE_10uA.t17 VDDA.t235 VDDA.t234 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X357 two_stage_opamp_dummy_magic_29_0.X.t19 two_stage_opamp_dummy_magic_29_0.Vb2.t21 two_stage_opamp_dummy_magic_29_0.VD3.t9 two_stage_opamp_dummy_magic_29_0.VD3.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X358 VOUT-.t83 two_stage_opamp_dummy_magic_29_0.cap_res_X.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X359 VOUT-.t84 two_stage_opamp_dummy_magic_29_0.cap_res_X.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X360 VOUT-.t85 two_stage_opamp_dummy_magic_29_0.cap_res_X.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X361 VOUT+.t79 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X362 VOUT+.t80 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X363 a_6350_30238.t1 a_6470_28630.t1 GNDA.t84 sky130_fd_pr__res_xhigh_po_0p35 l=6
X364 VOUT+.t81 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X365 VOUT+.t82 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t90 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X366 bgr_11_0.1st_Vout_2.t0 a_6540_22450.t15 VDDA.t21 VDDA.t20 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X367 VDDA.t41 bgr_11_0.1st_Vout_1.t19 bgr_11_0.V_TOP.t1 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X368 VDDA.t375 two_stage_opamp_dummy_magic_29_0.Vb3.t17 two_stage_opamp_dummy_magic_29_0.VD3.t27 VDDA.t374 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X369 VOUT-.t86 two_stage_opamp_dummy_magic_29_0.cap_res_X.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X370 GNDA.t55 two_stage_opamp_dummy_magic_29_0.Y.t41 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t4 VDDA.t75 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X371 VOUT+.t83 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t91 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X372 VDDA.t50 bgr_11_0.V_mir1.t16 bgr_11_0.1st_Vout_1.t0 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X373 VDDA.t96 two_stage_opamp_dummy_magic_29_0.Vb3.t18 two_stage_opamp_dummy_magic_29_0.VD4.t26 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X374 two_stage_opamp_dummy_magic_29_0.V_source.t2 VIN+.t3 two_stage_opamp_dummy_magic_29_0.VD2.t1 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X375 a_14420_6968.t1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t14 GNDA.t283 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X376 VOUT-.t87 two_stage_opamp_dummy_magic_29_0.cap_res_X.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X377 bgr_11_0.V_TOP.t35 VDDA.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X378 VOUT-.t88 two_stage_opamp_dummy_magic_29_0.cap_res_X.t73 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X379 GNDA.t98 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t23 two_stage_opamp_dummy_magic_29_0.V_source.t29 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X380 VOUT+.t4 two_stage_opamp_dummy_magic_29_0.Y.t42 VDDA.t4 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X381 VOUT+.t84 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X382 VOUT-.t89 two_stage_opamp_dummy_magic_29_0.cap_res_X.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X383 VOUT+.t85 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X384 GNDA.t218 GNDA.t217 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X385 a_12070_30088.t0 a_11950_28880.t0 GNDA.t1 sky130_fd_pr__res_xhigh_po_0p35 l=4
X386 VOUT+.t86 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t112 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X387 VOUT+.t87 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t113 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X388 VDDA.t32 bgr_11_0.V_TOP.t36 bgr_11_0.Vin+.t1 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X389 VOUT+.t88 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t134 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X390 VOUT-.t90 two_stage_opamp_dummy_magic_29_0.cap_res_X.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X391 GNDA.t223 GNDA.t221 two_stage_opamp_dummy_magic_29_0.Vb3.t2 GNDA.t222 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X392 VDDA.t39 two_stage_opamp_dummy_magic_29_0.Vb3.t19 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t10 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X393 GNDA.t220 GNDA.t219 two_stage_opamp_dummy_magic_29_0.err_amp_out.t3 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X394 VDDA.t303 VDDA.t301 GNDA.t157 VDDA.t302 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X395 bgr_11_0.V_TOP.t6 bgr_11_0.START_UP.t6 bgr_11_0.Vin-.t5 VDDA.t169 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X396 GNDA.t165 two_stage_opamp_dummy_magic_29_0.X.t42 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t10 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X397 VOUT+.t89 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t135 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X398 a_6540_22450.t6 a_6540_22450.t5 VDDA.t78 VDDA.t77 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X399 VOUT-.t91 two_stage_opamp_dummy_magic_29_0.cap_res_X.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X400 VOUT+.t90 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X401 bgr_11_0.1st_Vout_1.t20 bgr_11_0.cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X402 VDDA.t300 VDDA.t298 bgr_11_0.V_TOP.t10 VDDA.t299 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X403 VOUT-.t92 two_stage_opamp_dummy_magic_29_0.cap_res_X.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X404 VOUT+.t91 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X405 VDDA.t124 GNDA.t214 GNDA.t216 GNDA.t215 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.15
X406 VOUT-.t93 two_stage_opamp_dummy_magic_29_0.cap_res_X.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X407 VOUT-.t94 two_stage_opamp_dummy_magic_29_0.cap_res_X.t67 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X408 two_stage_opamp_dummy_magic_29_0.V_source.t28 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t24 GNDA.t99 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X409 two_stage_opamp_dummy_magic_29_0.X.t2 two_stage_opamp_dummy_magic_29_0.Vb2.t22 two_stage_opamp_dummy_magic_29_0.VD3.t7 two_stage_opamp_dummy_magic_29_0.VD3.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X410 VOUT-.t95 two_stage_opamp_dummy_magic_29_0.cap_res_X.t66 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X411 VOUT+.t92 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X412 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t1 bgr_11_0.V_TOP.t37 VDDA.t34 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X413 VOUT-.t96 two_stage_opamp_dummy_magic_29_0.cap_res_X.t65 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X414 VOUT+.t93 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X415 VOUT+.t94 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X416 VOUT+.t95 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X417 VOUT+.t96 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t110 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X418 VOUT-.t97 two_stage_opamp_dummy_magic_29_0.cap_res_X.t64 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X419 VOUT-.t11 two_stage_opamp_dummy_magic_29_0.X.t43 VDDA.t36 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X420 VOUT+.t97 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t111 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X421 VOUT+.t98 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X422 VOUT+.t99 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X423 VOUT-.t4 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t5 GNDA.t139 GNDA.t138 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X424 two_stage_opamp_dummy_magic_29_0.Y.t3 two_stage_opamp_dummy_magic_29_0.Vb2.t23 two_stage_opamp_dummy_magic_29_0.VD4.t5 two_stage_opamp_dummy_magic_29_0.VD4.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X425 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t3 two_stage_opamp_dummy_magic_29_0.V_err_gate.t7 VDDA.t17 VDDA.t16 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X426 two_stage_opamp_dummy_magic_29_0.Y.t13 two_stage_opamp_dummy_magic_29_0.Vb1.t26 two_stage_opamp_dummy_magic_29_0.VD2.t10 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X427 VOUT-.t98 two_stage_opamp_dummy_magic_29_0.cap_res_X.t63 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X428 VDDA.t297 VDDA.t295 two_stage_opamp_dummy_magic_29_0.Vb1.t9 VDDA.t296 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X429 VDDA.t233 bgr_11_0.PFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t6 VDDA.t232 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X430 VDDA.t294 VDDA.t292 two_stage_opamp_dummy_magic_29_0.err_amp_out.t2 VDDA.t293 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X431 VDDA.t175 two_stage_opamp_dummy_magic_29_0.V_err_gate.t8 two_stage_opamp_dummy_magic_29_0.V_err_p.t2 VDDA.t174 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X432 VOUT+.t100 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X433 bgr_11_0.PFET_GATE_10uA.t4 bgr_11_0.1st_Vout_2.t21 VDDA.t203 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X434 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t5 bgr_11_0.PFET_GATE_10uA.t19 VDDA.t231 VDDA.t230 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X435 VOUT+.t101 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X436 two_stage_opamp_dummy_magic_29_0.V_source.t19 VIN-.t4 two_stage_opamp_dummy_magic_29_0.VD1.t19 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X437 VOUT+.t102 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t88 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X438 bgr_11_0.1st_Vout_1.t21 bgr_11_0.cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X439 VOUT-.t99 two_stage_opamp_dummy_magic_29_0.cap_res_X.t62 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X440 VOUT+.t103 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t89 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X441 VOUT+.t104 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t108 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X442 VOUT-.t100 two_stage_opamp_dummy_magic_29_0.cap_res_X.t61 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X443 VOUT+.t105 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t109 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X444 GNDA.t111 bgr_11_0.NFET_GATE_10uA.t13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t1 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X445 VDDA.t120 bgr_11_0.V_TOP.t38 bgr_11_0.START_UP.t1 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X446 two_stage_opamp_dummy_magic_29_0.V_source.t11 VIN+.t4 two_stage_opamp_dummy_magic_29_0.VD2.t7 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X447 bgr_11_0.Vin-.t2 bgr_11_0.V_TOP.t39 VDDA.t122 VDDA.t121 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X448 bgr_11_0.1st_Vout_1.t22 bgr_11_0.cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X449 two_stage_opamp_dummy_magic_29_0.Y.t2 two_stage_opamp_dummy_magic_29_0.Vb2.t24 two_stage_opamp_dummy_magic_29_0.VD4.t3 two_stage_opamp_dummy_magic_29_0.VD4.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X450 two_stage_opamp_dummy_magic_29_0.V_source.t16 VIN-.t5 two_stage_opamp_dummy_magic_29_0.VD1.t16 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X451 VOUT+.t106 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t132 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X452 VOUT-.t101 two_stage_opamp_dummy_magic_29_0.cap_res_X.t60 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X453 VOUT+.t3 two_stage_opamp_dummy_magic_29_0.Y.t43 VDDA.t6 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X454 VOUT+.t107 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t133 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X455 VOUT+.t108 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X456 VOUT+.t109 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X457 two_stage_opamp_dummy_magic_29_0.Vb1.t1 two_stage_opamp_dummy_magic_29_0.Vb1.t0 two_stage_opamp_dummy_magic_29_0.Vb1_2.t2 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X458 VOUT-.t102 two_stage_opamp_dummy_magic_29_0.cap_res_X.t59 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X459 two_stage_opamp_dummy_magic_29_0.X.t23 two_stage_opamp_dummy_magic_29_0.VD3.t35 two_stage_opamp_dummy_magic_29_0.VD3.t37 two_stage_opamp_dummy_magic_29_0.VD3.t36 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X460 VDDA.t59 two_stage_opamp_dummy_magic_29_0.Vb3.t20 two_stage_opamp_dummy_magic_29_0.VD4.t25 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X461 VOUT-.t103 two_stage_opamp_dummy_magic_29_0.cap_res_X.t58 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X462 VOUT+.t110 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t80 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X463 GNDA.t156 VDDA.t421 bgr_11_0.V_TOP.t13 GNDA.t155 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X464 bgr_11_0.1st_Vout_1.t23 bgr_11_0.cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X465 VOUT-.t104 two_stage_opamp_dummy_magic_29_0.cap_res_X.t57 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X466 VOUT+.t111 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t81 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X467 GNDA.t114 bgr_11_0.NFET_GATE_10uA.t14 two_stage_opamp_dummy_magic_29_0.V_err_gate.t1 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X468 bgr_11_0.V_TOP.t40 VDDA.t82 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X469 VOUT-.t105 two_stage_opamp_dummy_magic_29_0.cap_res_X.t56 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X470 bgr_11_0.1st_Vout_2.t6 a_6540_22450.t16 VDDA.t406 VDDA.t405 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X471 VOUT-.t106 two_stage_opamp_dummy_magic_29_0.cap_res_X.t55 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X472 GNDA.t154 VDDA.t289 VDDA.t291 VDDA.t290 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X473 VOUT+.t112 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t106 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X474 VOUT+.t113 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t107 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X475 two_stage_opamp_dummy_magic_29_0.X.t10 two_stage_opamp_dummy_magic_29_0.Vb1.t27 two_stage_opamp_dummy_magic_29_0.VD1.t5 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X476 VOUT+.t114 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t130 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X477 bgr_11_0.V_p_1.t1 VDDA.t422 GNDA.t153 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X478 two_stage_opamp_dummy_magic_29_0.X.t1 two_stage_opamp_dummy_magic_29_0.Vb2.t25 two_stage_opamp_dummy_magic_29_0.VD3.t5 two_stage_opamp_dummy_magic_29_0.VD3.t4 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X479 VOUT+.t115 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t131 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X480 two_stage_opamp_dummy_magic_29_0.V_source.t27 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t25 GNDA.t118 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X481 bgr_11_0.NFET_GATE_10uA.t2 bgr_11_0.PFET_GATE_10uA.t20 VDDA.t229 VDDA.t228 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X482 VOUT-.t10 two_stage_opamp_dummy_magic_29_0.X.t44 VDDA.t112 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X483 two_stage_opamp_dummy_magic_29_0.Vb3.t5 bgr_11_0.NFET_GATE_10uA.t15 GNDA.t130 GNDA.t129 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X484 bgr_11_0.1st_Vout_2.t22 bgr_11_0.cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X485 VDDA.t26 two_stage_opamp_dummy_magic_29_0.Vb3.t21 two_stage_opamp_dummy_magic_29_0.VD3.t26 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X486 two_stage_opamp_dummy_magic_29_0.Y.t6 two_stage_opamp_dummy_magic_29_0.Vb2.t26 two_stage_opamp_dummy_magic_29_0.VD4.t7 two_stage_opamp_dummy_magic_29_0.VD4.t6 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X487 VOUT-.t9 two_stage_opamp_dummy_magic_29_0.X.t45 VDDA.t392 VDDA.t391 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X488 bgr_11_0.V_mir1.t5 bgr_11_0.V_mir1.t4 VDDA.t166 VDDA.t165 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X489 two_stage_opamp_dummy_magic_29_0.Y.t23 GNDA.t211 GNDA.t213 GNDA.t212 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X490 bgr_11_0.1st_Vout_2.t5 bgr_11_0.V_CUR_REF_REG.t3 bgr_11_0.V_p_2.t1 GNDA.t280 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X491 two_stage_opamp_dummy_magic_29_0.X.t4 two_stage_opamp_dummy_magic_29_0.Vb1.t28 two_stage_opamp_dummy_magic_29_0.VD1.t4 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X492 bgr_11_0.1st_Vout_1.t24 bgr_11_0.cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X493 VOUT-.t107 two_stage_opamp_dummy_magic_29_0.cap_res_X.t54 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X494 VOUT+.t116 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X495 two_stage_opamp_dummy_magic_29_0.V_source.t15 VIN-.t6 two_stage_opamp_dummy_magic_29_0.VD1.t13 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X496 VOUT-.t108 two_stage_opamp_dummy_magic_29_0.cap_res_X.t53 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X497 VOUT+.t117 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X498 bgr_11_0.1st_Vout_2.t23 bgr_11_0.cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X499 a_14540_6968.t1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t0 GNDA.t83 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X500 VOUT+.t118 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t104 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X501 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t0 bgr_11_0.NFET_GATE_10uA.t16 GNDA.t25 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X502 GNDA.t120 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t26 two_stage_opamp_dummy_magic_29_0.V_source.t26 GNDA.t119 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X503 GNDA.t209 GNDA.t207 VDDA.t69 GNDA.t208 sky130_fd_pr__nfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.15
X504 VOUT-.t109 two_stage_opamp_dummy_magic_29_0.cap_res_X.t52 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X505 GNDA.t186 GNDA.t210 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X506 GNDA.t132 bgr_11_0.NFET_GATE_10uA.t17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t2 GNDA.t131 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X507 two_stage_opamp_dummy_magic_29_0.V_source.t10 VIN+.t5 two_stage_opamp_dummy_magic_29_0.VD2.t6 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X508 VOUT+.t119 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t105 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X509 VOUT-.t110 two_stage_opamp_dummy_magic_29_0.cap_res_X.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X510 two_stage_opamp_dummy_magic_29_0.Vb1.t10 GNDA.t205 GNDA.t206 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X511 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t1 VIN-.t7 two_stage_opamp_dummy_magic_29_0.V_p_mir.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X512 two_stage_opamp_dummy_magic_29_0.V_source.t21 VIN-.t8 two_stage_opamp_dummy_magic_29_0.VD1.t21 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X513 bgr_11_0.1st_Vout_2.t24 bgr_11_0.cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X514 GNDA.t23 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t6 VOUT-.t1 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X515 VOUT+.t16 VDDA.t286 VDDA.t288 VDDA.t287 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X516 VOUT+.t2 two_stage_opamp_dummy_magic_29_0.Y.t44 VDDA.t148 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X517 VOUT+.t120 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t124 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X518 VOUT-.t111 two_stage_opamp_dummy_magic_29_0.cap_res_X.t50 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X519 VDDA.t98 two_stage_opamp_dummy_magic_29_0.Vb3.t22 two_stage_opamp_dummy_magic_29_0.VD4.t24 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X520 VOUT+.t121 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t125 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X521 VOUT-.t112 two_stage_opamp_dummy_magic_29_0.cap_res_X.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X522 bgr_11_0.1st_Vout_1.t25 bgr_11_0.cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X523 GNDA.t11 bgr_11_0.NFET_GATE_10uA.t18 two_stage_opamp_dummy_magic_29_0.Vb2.t0 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X524 bgr_11_0.1st_Vout_2.t25 bgr_11_0.cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X525 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t0 bgr_11_0.NFET_GATE_10uA.t19 GNDA.t62 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X526 bgr_11_0.PFET_GATE_10uA.t9 bgr_11_0.1st_Vout_2.t26 VDDA.t201 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X527 VOUT+.t122 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X528 VOUT+.t123 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X529 bgr_11_0.1st_Vout_1.t26 bgr_11_0.cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X530 VOUT-.t113 two_stage_opamp_dummy_magic_29_0.cap_res_X.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X531 VOUT-.t114 two_stage_opamp_dummy_magic_29_0.cap_res_X.t47 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X532 GNDA.t34 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t7 VOUT-.t2 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X533 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t5 two_stage_opamp_dummy_magic_29_0.Y.t45 VDDA.t149 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X534 VOUT-.t115 two_stage_opamp_dummy_magic_29_0.cap_res_X.t46 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X535 bgr_11_0.1st_Vout_2.t27 bgr_11_0.cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X536 GNDA.t186 GNDA.t185 bgr_11_0.Vin-.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X537 two_stage_opamp_dummy_magic_29_0.X.t9 two_stage_opamp_dummy_magic_29_0.Vb1.t29 two_stage_opamp_dummy_magic_29_0.VD1.t3 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X538 two_stage_opamp_dummy_magic_29_0.V_source.t25 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t27 GNDA.t122 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X539 VOUT-.t116 two_stage_opamp_dummy_magic_29_0.cap_res_X.t45 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X540 a_3110_6968.t0 two_stage_opamp_dummy_magic_29_0.V_tot.t0 GNDA.t17 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X541 VOUT-.t117 two_stage_opamp_dummy_magic_29_0.cap_res_X.t44 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X542 bgr_11_0.1st_Vout_2.t1 a_6540_22450.t17 VDDA.t57 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X543 VOUT-.t8 two_stage_opamp_dummy_magic_29_0.X.t46 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X544 VOUT-.t118 two_stage_opamp_dummy_magic_29_0.cap_res_X.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X545 bgr_11_0.1st_Vout_1.t27 bgr_11_0.cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X546 bgr_11_0.V_TOP.t2 bgr_11_0.1st_Vout_1.t28 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X547 VOUT-.t119 two_stage_opamp_dummy_magic_29_0.cap_res_X.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X548 VOUT-.t120 two_stage_opamp_dummy_magic_29_0.cap_res_X.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X549 VOUT+.t124 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t42 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X550 VOUT+.t125 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t43 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X551 two_stage_opamp_dummy_magic_29_0.X.t3 two_stage_opamp_dummy_magic_29_0.Vb1.t30 two_stage_opamp_dummy_magic_29_0.VD1.t2 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X552 VOUT-.t121 two_stage_opamp_dummy_magic_29_0.cap_res_X.t40 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X553 bgr_11_0.1st_Vout_1.t1 bgr_11_0.V_mir1.t17 VDDA.t68 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X554 GNDA.t134 two_stage_opamp_dummy_magic_29_0.err_amp_out.t5 two_stage_opamp_dummy_magic_29_0.V_source.t13 GNDA.t133 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X555 VDDA.t282 VDDA.t280 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t15 VDDA.t281 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X556 VOUT+.t126 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t100 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X557 bgr_11_0.PFET_GATE_10uA.t1 VDDA.t423 GNDA.t149 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X558 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t11 bgr_11_0.PFET_GATE_10uA.t21 VDDA.t227 VDDA.t226 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X559 two_stage_opamp_dummy_magic_29_0.Y.t7 two_stage_opamp_dummy_magic_29_0.Vb2.t27 two_stage_opamp_dummy_magic_29_0.VD4.t9 two_stage_opamp_dummy_magic_29_0.VD4.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X560 VDDA.t285 VDDA.t283 GNDA.t150 VDDA.t284 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X561 VOUT+.t127 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t101 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X562 GNDA.t204 GNDA.t202 two_stage_opamp_dummy_magic_29_0.X.t12 GNDA.t203 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X563 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t6 two_stage_opamp_dummy_magic_29_0.X.t47 VDDA.t394 GNDA.t164 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X564 bgr_11_0.V_TOP.t41 VDDA.t83 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X565 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t5 two_stage_opamp_dummy_magic_29_0.X.t48 VDDA.t135 GNDA.t163 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X566 VDDA.t279 VDDA.t277 bgr_11_0.PFET_GATE_10uA.t3 VDDA.t278 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X567 VDDA.t71 bgr_11_0.V_TOP.t42 bgr_11_0.START_UP.t0 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X568 two_stage_opamp_dummy_magic_29_0.V_source.t17 VIN-.t9 two_stage_opamp_dummy_magic_29_0.VD1.t17 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X569 VOUT-.t122 two_stage_opamp_dummy_magic_29_0.cap_res_X.t39 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X570 VOUT+.t1 two_stage_opamp_dummy_magic_29_0.Y.t46 VDDA.t109 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X571 VOUT+.t128 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X572 GNDA.t201 GNDA.t200 two_stage_opamp_dummy_magic_29_0.Y.t22 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.8 as=0.3 ps=1.9 w=1.5 l=0.15
X573 VOUT-.t123 two_stage_opamp_dummy_magic_29_0.cap_res_X.t38 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X574 VOUT-.t124 two_stage_opamp_dummy_magic_29_0.cap_res_X.t37 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X575 VOUT+.t129 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X576 a_6540_22450.t4 a_6540_22450.t3 VDDA.t158 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X577 bgr_11_0.V_TOP.t43 VDDA.t72 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X578 VOUT-.t125 two_stage_opamp_dummy_magic_29_0.cap_res_X.t36 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X579 VOUT+.t130 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X580 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t3 two_stage_opamp_dummy_magic_29_0.Y.t47 GNDA.t67 VDDA.t110 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X581 two_stage_opamp_dummy_magic_29_0.VD1.t12 VIN-.t10 two_stage_opamp_dummy_magic_29_0.V_source.t14 GNDA.t178 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X582 a_11420_30238.t0 a_11300_28630.t1 GNDA.t79 sky130_fd_pr__res_xhigh_po_0p35 l=6
X583 two_stage_opamp_dummy_magic_29_0.Vb2_2.t9 two_stage_opamp_dummy_magic_29_0.Vb2_2.t7 two_stage_opamp_dummy_magic_29_0.Vb2_2.t9 two_stage_opamp_dummy_magic_29_0.Vb2_2.t8 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X584 two_stage_opamp_dummy_magic_29_0.cap_res_X.t143 two_stage_opamp_dummy_magic_29_0.X.t24 GNDA.t282 sky130_fd_pr__res_high_po_1p41 l=1.41
X585 VOUT-.t126 two_stage_opamp_dummy_magic_29_0.cap_res_X.t35 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X586 two_stage_opamp_dummy_magic_29_0.X.t0 two_stage_opamp_dummy_magic_29_0.Vb2.t28 two_stage_opamp_dummy_magic_29_0.VD3.t3 two_stage_opamp_dummy_magic_29_0.VD3.t2 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X587 VDDA.t225 bgr_11_0.PFET_GATE_10uA.t22 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t4 VDDA.t224 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X588 VOUT-.t127 two_stage_opamp_dummy_magic_29_0.cap_res_X.t34 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X589 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t3 bgr_11_0.PFET_GATE_10uA.t23 VDDA.t223 VDDA.t222 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X590 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t4 two_stage_opamp_dummy_magic_29_0.Y.t48 VDDA.t145 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X591 bgr_11_0.V_TOP.t44 VDDA.t142 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X592 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t3 two_stage_opamp_dummy_magic_29_0.Y.t49 VDDA.t146 GNDA.t86 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X593 VOUT-.t128 two_stage_opamp_dummy_magic_29_0.cap_res_X.t33 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X594 two_stage_opamp_dummy_magic_29_0.V_p_mir.t1 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t28 GNDA.t124 GNDA.t123 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X595 two_stage_opamp_dummy_magic_29_0.Y.t20 two_stage_opamp_dummy_magic_29_0.VD4.t32 two_stage_opamp_dummy_magic_29_0.VD4.t34 two_stage_opamp_dummy_magic_29_0.VD4.t33 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X596 two_stage_opamp_dummy_magic_29_0.VD2.t18 VIN+.t6 two_stage_opamp_dummy_magic_29_0.V_source.t12 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X597 VOUT-.t129 two_stage_opamp_dummy_magic_29_0.cap_res_X.t32 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X598 VOUT+.t131 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X599 two_stage_opamp_dummy_magic_29_0.V_source.t24 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t29 GNDA.t29 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X600 bgr_11_0.1st_Vout_1.t4 bgr_11_0.V_mir1.t18 VDDA.t164 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X601 VOUT-.t130 two_stage_opamp_dummy_magic_29_0.cap_res_X.t31 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X602 VDDA.t276 VDDA.t274 VOUT+.t15 VDDA.t275 sky130_fd_pr__pfet_01v8 ad=2.4 pd=12.8 as=1.2 ps=6.4 w=6 l=0.15
X603 VOUT+.t132 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t70 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X604 bgr_11_0.V_mir1.t12 bgr_11_0.Vin-.t8 bgr_11_0.V_p_1.t0 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.2
X605 VOUT-.t131 two_stage_opamp_dummy_magic_29_0.cap_res_X.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X606 VOUT+.t133 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t71 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X607 VOUT+.t134 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X608 VOUT+.t135 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t49 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X609 VOUT+.t136 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t94 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X610 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t2 bgr_11_0.PFET_GATE_10uA.t24 VDDA.t221 VDDA.t220 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X611 VOUT-.t7 two_stage_opamp_dummy_magic_29_0.X.t49 VDDA.t409 VDDA.t408 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=1.2 ps=6.4 w=6 l=0.15
X612 VOUT+.t137 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t95 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X613 VDDA.t219 bgr_11_0.PFET_GATE_10uA.t25 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t1 VDDA.t218 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X614 VDDA.t273 VDDA.t271 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t5 VDDA.t272 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X615 two_stage_opamp_dummy_magic_29_0.VD3.t34 two_stage_opamp_dummy_magic_29_0.VD3.t32 two_stage_opamp_dummy_magic_29_0.X.t16 two_stage_opamp_dummy_magic_29_0.VD3.t33 sky130_fd_pr__pfet_01v8 ad=1.4 pd=7.8 as=0.7 ps=3.9 w=3.5 l=0.2
X616 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t4 GNDA.t198 GNDA.t199 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.15
X617 two_stage_opamp_dummy_magic_29_0.X.t17 GNDA.t196 GNDA.t197 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.6 ps=3.8 w=1.5 l=0.15
X618 two_stage_opamp_dummy_magic_29_0.Vb3.t0 two_stage_opamp_dummy_magic_29_0.Vb2.t29 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t8 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t7 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X619 VOUT-.t132 two_stage_opamp_dummy_magic_29_0.cap_res_X.t29 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X620 a_14540_6968.t0 two_stage_opamp_dummy_magic_29_0.V_tot.t1 GNDA.t53 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X621 VOUT+.t138 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X622 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t0 bgr_11_0.V_TOP.t45 VDDA.t144 VDDA.t143 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X623 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t9 two_stage_opamp_dummy_magic_29_0.X.t50 GNDA.t162 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X624 VOUT-.t133 two_stage_opamp_dummy_magic_29_0.cap_res_X.t28 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X625 bgr_11_0.V_TOP.t46 VDDA.t127 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X626 GNDA.t52 a_5820_28824.t1 GNDA.t51 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X627 two_stage_opamp_dummy_magic_29_0.Y.t17 two_stage_opamp_dummy_magic_29_0.Vb2.t30 two_stage_opamp_dummy_magic_29_0.VD4.t15 two_stage_opamp_dummy_magic_29_0.VD4.t14 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X628 bgr_11_0.V_TOP.t4 bgr_11_0.1st_Vout_1.t29 VDDA.t151 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X629 two_stage_opamp_dummy_magic_29_0.VD3.t25 two_stage_opamp_dummy_magic_29_0.Vb3.t23 VDDA.t379 VDDA.t378 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X630 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t8 two_stage_opamp_dummy_magic_29_0.X.t51 GNDA.t161 VDDA.t187 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X631 GNDA.t145 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t8 VOUT+.t14 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X632 VOUT-.t134 two_stage_opamp_dummy_magic_29_0.cap_res_X.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X633 VOUT-.t135 two_stage_opamp_dummy_magic_29_0.cap_res_X.t26 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X634 VOUT-.t136 two_stage_opamp_dummy_magic_29_0.cap_res_X.t25 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X635 VOUT+.t139 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t79 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X636 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t4 two_stage_opamp_dummy_magic_29_0.X.t52 VDDA.t46 GNDA.t160 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X637 VOUT-.t137 two_stage_opamp_dummy_magic_29_0.cap_res_X.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X638 VOUT+.t140 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X639 two_stage_opamp_dummy_magic_29_0.VD4.t23 two_stage_opamp_dummy_magic_29_0.Vb3.t24 VDDA.t199 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X640 VOUT-.t138 two_stage_opamp_dummy_magic_29_0.cap_res_X.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X641 bgr_11_0.V_TOP.t8 bgr_11_0.1st_Vout_1.t30 VDDA.t191 VDDA.t190 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X642 bgr_11_0.1st_Vout_2.t28 bgr_11_0.cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X643 two_stage_opamp_dummy_magic_29_0.VD2.t9 two_stage_opamp_dummy_magic_29_0.Vb1.t31 two_stage_opamp_dummy_magic_29_0.Y.t12 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X644 VOUT-.t139 two_stage_opamp_dummy_magic_29_0.cap_res_X.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X645 VOUT+.t141 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X646 VDDA.t270 VDDA.t268 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t4 VDDA.t269 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X647 VOUT+.t142 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t76 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X648 two_stage_opamp_dummy_magic_29_0.Vb3.t4 bgr_11_0.NFET_GATE_10uA.t20 GNDA.t106 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X649 GNDA.t195 GNDA.t193 VOUT+.t18 GNDA.t194 sky130_fd_pr__nfet_01v8 ad=2.8 pd=14.8 as=1.4 ps=7.4 w=7 l=0.6
X650 VOUT+.t143 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t77 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X651 VOUT-.t140 two_stage_opamp_dummy_magic_29_0.cap_res_X.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X652 bgr_11_0.1st_Vout_1.t31 bgr_11_0.cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X653 VOUT-.t141 two_stage_opamp_dummy_magic_29_0.cap_res_X.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X654 VOUT+.t144 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X655 VOUT+.t145 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X656 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t2 two_stage_opamp_dummy_magic_29_0.Y.t50 GNDA.t140 VDDA.t182 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X657 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t1 two_stage_opamp_dummy_magic_29_0.Y.t51 GNDA.t141 VDDA.t183 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X658 VOUT-.t142 two_stage_opamp_dummy_magic_29_0.cap_res_X.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X659 VOUT+.t146 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X660 bgr_11_0.Vin-.t4 bgr_11_0.START_UP.t7 bgr_11_0.V_TOP.t5 VDDA.t162 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X661 two_stage_opamp_dummy_magic_29_0.VD4.t22 two_stage_opamp_dummy_magic_29_0.Vb3.t25 VDDA.t63 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X662 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t2 two_stage_opamp_dummy_magic_29_0.Y.t52 VDDA.t184 GNDA.t142 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X663 two_stage_opamp_dummy_magic_29_0.VD2.t4 VIN+.t7 two_stage_opamp_dummy_magic_29_0.V_source.t8 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X664 VOUT+.t147 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X665 VOUT-.t143 two_stage_opamp_dummy_magic_29_0.cap_res_X.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X666 VOUT+.t148 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t98 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X667 VOUT+.t149 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t99 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X668 VOUT-.t144 two_stage_opamp_dummy_magic_29_0.cap_res_X.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X669 bgr_11_0.V_mir1.t3 bgr_11_0.V_mir1.t2 VDDA.t19 VDDA.t18 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X670 two_stage_opamp_dummy_magic_29_0.VD3.t24 two_stage_opamp_dummy_magic_29_0.Vb3.t26 VDDA.t377 VDDA.t376 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X671 a_3230_6968.t0 two_stage_opamp_dummy_magic_29_0.V_tot.t3 GNDA.t109 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X672 two_stage_opamp_dummy_magic_29_0.VD2.t0 VIN+.t8 two_stage_opamp_dummy_magic_29_0.V_source.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X673 two_stage_opamp_dummy_magic_29_0.V_p_mir.t3 VIN+.t9 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X674 two_stage_opamp_dummy_magic_29_0.V_source.t23 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t30 GNDA.t30 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X675 two_stage_opamp_dummy_magic_29_0.Vb1_2.t1 two_stage_opamp_dummy_magic_29_0.Vb1.t6 two_stage_opamp_dummy_magic_29_0.Vb1.t7 GNDA.t47 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X676 bgr_11_0.V_p_2.t0 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t7 a_6540_22450.t0 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=1 ps=5.8 w=2.5 l=0.2
X677 bgr_11_0.V_TOP.t9 VDDA.t265 VDDA.t267 VDDA.t266 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X678 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t0 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t8 two_stage_opamp_dummy_magic_29_0.V_err_gate.t0 VDDA.t22 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X679 bgr_11_0.V_TOP.t47 VDDA.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X680 VDDA.t264 VDDA.t262 two_stage_opamp_dummy_magic_29_0.V_err_gate.t3 VDDA.t263 sky130_fd_pr__pfet_01v8 ad=1 pd=5.8 as=0.5 ps=2.9 w=2.5 l=0.15
X681 VOUT-.t5 VDDA.t259 VDDA.t261 VDDA.t260 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.4 as=2.4 ps=12.8 w=6 l=0.15
X682 VOUT-.t145 two_stage_opamp_dummy_magic_29_0.cap_res_X.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X683 VDDA.t398 bgr_11_0.V_TOP.t48 bgr_11_0.Vin-.t1 VDDA.t397 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X684 VDDA.t133 two_stage_opamp_dummy_magic_29_0.V_err_gate.t9 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t2 VDDA.t132 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X685 VOUT+.t150 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X686 VOUT+.t151 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X687 VOUT-.t146 two_stage_opamp_dummy_magic_29_0.cap_res_X.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X688 VOUT+.t152 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t68 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X689 two_stage_opamp_dummy_magic_29_0.Vb1.t8 bgr_11_0.PFET_GATE_10uA.t26 VDDA.t217 VDDA.t216 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X690 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t2 bgr_11_0.PFET_GATE_10uA.t27 VDDA.t215 VDDA.t214 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X691 two_stage_opamp_dummy_magic_29_0.err_amp_out.t0 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t9 two_stage_opamp_dummy_magic_29_0.V_err_p.t0 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X692 two_stage_opamp_dummy_magic_29_0.V_err_p.t1 two_stage_opamp_dummy_magic_29_0.V_tot.t5 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t2 VDDA.t138 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X693 VOUT-.t147 two_stage_opamp_dummy_magic_29_0.cap_res_X.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X694 VOUT-.t148 two_stage_opamp_dummy_magic_29_0.cap_res_X.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X695 GNDA.t108 a_6470_28630.t0 GNDA.t84 sky130_fd_pr__res_xhigh_po_0p35 l=6
X696 VOUT-.t149 two_stage_opamp_dummy_magic_29_0.cap_res_X.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X697 GNDA.t192 GNDA.t190 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t13 GNDA.t191 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X698 VDDA.t100 a_6540_22450.t18 bgr_11_0.1st_Vout_2.t2 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X699 two_stage_opamp_dummy_magic_29_0.VD3.t23 two_stage_opamp_dummy_magic_29_0.Vb3.t27 VDDA.t197 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X700 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t7 two_stage_opamp_dummy_magic_29_0.X.t53 GNDA.t159 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X701 VOUT+.t153 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t69 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X702 bgr_11_0.1st_Vout_2.t29 bgr_11_0.cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X703 VOUT+.t154 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t142 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X704 VOUT+.t155 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t143 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X705 GNDA.t116 bgr_11_0.NFET_GATE_10uA.t21 two_stage_opamp_dummy_magic_29_0.Vb2.t7 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X706 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t13 GNDA.t187 GNDA.t189 GNDA.t188 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X707 GNDA.t147 VDDA.t424 bgr_11_0.V_p_2.t2 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X708 bgr_11_0.V_mir1.t1 bgr_11_0.V_mir1.t0 VDDA.t11 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X709 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t3 two_stage_opamp_dummy_magic_29_0.X.t54 VDDA.t393 GNDA.t158 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X710 VOUT+.t156 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t92 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X711 bgr_11_0.PFET_GATE_10uA.t2 VDDA.t256 VDDA.t258 VDDA.t257 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X712 VOUT+.t157 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t93 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X713 two_stage_opamp_dummy_magic_29_0.VD2.t8 two_stage_opamp_dummy_magic_29_0.Vb1.t32 two_stage_opamp_dummy_magic_29_0.Y.t4 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X714 VOUT-.t150 two_stage_opamp_dummy_magic_29_0.cap_res_X.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X715 two_stage_opamp_dummy_magic_29_0.Vb2.t3 two_stage_opamp_dummy_magic_29_0.Vb2_2.t4 two_stage_opamp_dummy_magic_29_0.Vb2_2.t6 two_stage_opamp_dummy_magic_29_0.Vb2_2.t5 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=1.4 ps=7.8 w=3.5 l=0.2
X716 a_12070_30088.t1 bgr_11_0.V_CUR_REF_REG.t2 GNDA.t279 sky130_fd_pr__res_xhigh_po_0p35 l=4
X717 VOUT-.t151 two_stage_opamp_dummy_magic_29_0.cap_res_X.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X718 VOUT-.t152 two_stage_opamp_dummy_magic_29_0.cap_res_X.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X719 bgr_11_0.1st_Vout_2.t30 bgr_11_0.cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X720 GNDA.t184 GNDA.t182 bgr_11_0.NFET_GATE_10uA.t4 GNDA.t183 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X721 bgr_11_0.Vin-.t0 bgr_11_0.V_TOP.t49 VDDA.t400 VDDA.t399 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X722 VOUT+.t17 GNDA.t179 GNDA.t181 GNDA.t180 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=2.8 ps=14.8 w=7 l=0.6
X723 VDDA.t255 VDDA.t253 VDDA.t255 VDDA.t254 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0 ps=0 w=3.5 l=0.2
X724 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t0 two_stage_opamp_dummy_magic_29_0.Y.t53 GNDA.t143 VDDA.t185 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X725 VOUT+.t158 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t102 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X726 VOUT-.t153 two_stage_opamp_dummy_magic_29_0.cap_res_X.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X727 VOUT-.t154 two_stage_opamp_dummy_magic_29_0.cap_res_X.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X728 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t0 a_13940_3166.t1 GNDA.t66 sky130_fd_pr__res_xhigh_po_0p35 l=2.63
X729 VDDA.t179 a_6540_22450.t1 a_6540_22450.t2 VDDA.t178 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X730 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t1 two_stage_opamp_dummy_magic_29_0.Y.t54 VDDA.t167 GNDA.t117 sky130_fd_pr__nfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.15
X731 two_stage_opamp_dummy_magic_29_0.VD2.t2 VIN+.t10 two_stage_opamp_dummy_magic_29_0.V_source.t6 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.3 pd=1.9 as=0.3 ps=1.9 w=1.5 l=0.15
X732 VOUT-.t155 two_stage_opamp_dummy_magic_29_0.cap_res_X.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X733 bgr_11_0.1st_Vout_2.t31 bgr_11_0.cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X734 VOUT-.t156 two_stage_opamp_dummy_magic_29_0.cap_res_X.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X735 two_stage_opamp_dummy_magic_29_0.V_source.t22 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t31 GNDA.t35 GNDA.t3 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.9 as=0.5 ps=2.9 w=2.5 l=0.15
X736 VOUT+.t159 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t103 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X737 bgr_11_0.V_CUR_REF_REG.t1 VDDA.t250 VDDA.t252 VDDA.t251 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X738 VOUT+.t160 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t128 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X739 two_stage_opamp_dummy_magic_29_0.Vb3.t1 bgr_11_0.NFET_GATE_10uA.t22 GNDA.t27 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X740 VDDA.t213 bgr_11_0.PFET_GATE_10uA.t28 bgr_11_0.V_CUR_REF_REG.t0 VDDA.t212 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X741 two_stage_opamp_dummy_magic_29_0.VD3.t1 two_stage_opamp_dummy_magic_29_0.Vb2.t31 two_stage_opamp_dummy_magic_29_0.X.t18 two_stage_opamp_dummy_magic_29_0.VD3.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X742 GNDA.t89 bgr_11_0.NFET_GATE_10uA.t23 two_stage_opamp_dummy_magic_29_0.Vb3.t3 GNDA.t88 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X743 VOUT-.t157 two_stage_opamp_dummy_magic_29_0.cap_res_X.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X744 bgr_11_0.1st_Vout_1.t32 bgr_11_0.cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X745 VOUT-.t158 two_stage_opamp_dummy_magic_29_0.cap_res_X.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X746 VOUT-.t159 two_stage_opamp_dummy_magic_29_0.cap_res_X.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X747 VOUT+.t0 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t9 GNDA.t8 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=1.4 pd=7.4 as=1.4 ps=7.4 w=7 l=0.6
X748 VOUT+.t161 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t129 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X749 a_14420_6968.t0 two_stage_opamp_dummy_magic_29_0.V_tot.t2 GNDA.t107 sky130_fd_pr__res_xhigh_po_0p35 l=1.75
X750 VOUT-.t160 two_stage_opamp_dummy_magic_29_0.cap_res_X.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X751 a_5700_30088.t1 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t6 GNDA.t281 sky130_fd_pr__res_xhigh_po_0p35 l=4.28
X752 two_stage_opamp_dummy_magic_29_0.VD3.t22 two_stage_opamp_dummy_magic_29_0.Vb3.t28 VDDA.t30 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X753 two_stage_opamp_dummy_magic_29_0.VD4.t1 two_stage_opamp_dummy_magic_29_0.Vb2.t32 two_stage_opamp_dummy_magic_29_0.Y.t1 two_stage_opamp_dummy_magic_29_0.VD4.t0 sky130_fd_pr__pfet_01v8 ad=0.7 pd=3.9 as=0.7 ps=3.9 w=3.5 l=0.2
X754 bgr_11_0.1st_Vout_2.t32 bgr_11_0.cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X755 VOUT-.t161 two_stage_opamp_dummy_magic_29_0.cap_res_X.t0 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
R0 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.t15 362.341
R1 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.t14 355.094
R2 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n10 302.183
R3 bgr_11_0.1st_Vout_2.n7 bgr_11_0.1st_Vout_2.n6 302.183
R4 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n5 297.683
R5 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t26 194.809
R6 bgr_11_0.1st_Vout_2.n11 bgr_11_0.1st_Vout_2.t9 194.809
R7 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t21 194.809
R8 bgr_11_0.1st_Vout_2.n8 bgr_11_0.1st_Vout_2.t7 194.809
R9 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n11 166.03
R10 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n8 166.03
R11 bgr_11_0.1st_Vout_2.t5 bgr_11_0.1st_Vout_2.n12 49.5021
R12 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t4 39.4005
R13 bgr_11_0.1st_Vout_2.n10 bgr_11_0.1st_Vout_2.t6 39.4005
R14 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t2 39.4005
R15 bgr_11_0.1st_Vout_2.n6 bgr_11_0.1st_Vout_2.t0 39.4005
R16 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t3 39.4005
R17 bgr_11_0.1st_Vout_2.n5 bgr_11_0.1st_Vout_2.t1 39.4005
R18 bgr_11_0.1st_Vout_2.n9 bgr_11_0.1st_Vout_2.n0 35.7185
R19 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t32 4.8295
R20 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t12 4.8295
R21 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t13 4.8295
R22 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t19 4.8295
R23 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t30 4.8295
R24 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t11 4.8295
R25 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t23 4.8295
R26 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t28 4.8295
R27 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t8 4.8295
R28 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t27 4.5005
R29 bgr_11_0.1st_Vout_2.n1 bgr_11_0.1st_Vout_2.t20 4.5005
R30 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t31 4.5005
R31 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t25 4.5005
R32 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t24 4.5005
R33 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.t18 4.5005
R34 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t17 4.5005
R35 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t10 4.5005
R36 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t29 4.5005
R37 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t22 4.5005
R38 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.t16 4.5005
R39 bgr_11_0.1st_Vout_2.n12 bgr_11_0.1st_Vout_2.n3 4.5005
R40 bgr_11_0.1st_Vout_2.n4 bgr_11_0.1st_Vout_2.n9 2.90725
R41 bgr_11_0.1st_Vout_2.n0 bgr_11_0.1st_Vout_2.n2 2.2095
R42 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n4 1.1255
R43 bgr_11_0.1st_Vout_2.n3 bgr_11_0.1st_Vout_2.n7 1.1255
R44 bgr_11_0.1st_Vout_2.n2 bgr_11_0.1st_Vout_2.n1 0.8935
R45 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.t26 614.04
R46 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.n0 510.991
R47 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n25 509.226
R48 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t22 369.534
R49 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t27 369.534
R50 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.t11 369.534
R51 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.t10 369.534
R52 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.t25 369.534
R53 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t24 369.534
R54 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.n11 301.933
R55 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n9 301.933
R56 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.n7 301.933
R57 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.n5 301.933
R58 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t20 249.034
R59 bgr_11_0.PFET_GATE_10uA.n0 bgr_11_0.PFET_GATE_10uA.t28 249.034
R60 bgr_11_0.PFET_GATE_10uA.n22 bgr_11_0.PFET_GATE_10uA.t12 192.8
R61 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.t16 192.8
R62 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.t23 192.8
R63 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.t14 192.8
R64 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.t19 192.8
R65 bgr_11_0.PFET_GATE_10uA.n19 bgr_11_0.PFET_GATE_10uA.t18 192.8
R66 bgr_11_0.PFET_GATE_10uA.n16 bgr_11_0.PFET_GATE_10uA.t21 192.8
R67 bgr_11_0.PFET_GATE_10uA.n15 bgr_11_0.PFET_GATE_10uA.t15 192.8
R68 bgr_11_0.PFET_GATE_10uA.n2 bgr_11_0.PFET_GATE_10uA.t17 192.8
R69 bgr_11_0.PFET_GATE_10uA.n1 bgr_11_0.PFET_GATE_10uA.t13 192.8
R70 bgr_11_0.PFET_GATE_10uA.n21 bgr_11_0.PFET_GATE_10uA.n20 176.733
R71 bgr_11_0.PFET_GATE_10uA.n20 bgr_11_0.PFET_GATE_10uA.n19 176.733
R72 bgr_11_0.PFET_GATE_10uA.n23 bgr_11_0.PFET_GATE_10uA.n22 176.733
R73 bgr_11_0.PFET_GATE_10uA.n24 bgr_11_0.PFET_GATE_10uA.n23 176.733
R74 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.n17 166.343
R75 bgr_11_0.PFET_GATE_10uA.n4 bgr_11_0.PFET_GATE_10uA.n3 166.343
R76 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.t0 119.118
R77 bgr_11_0.PFET_GATE_10uA.n6 bgr_11_0.PFET_GATE_10uA.t1 104.474
R78 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n16 56.2338
R79 bgr_11_0.PFET_GATE_10uA.n17 bgr_11_0.PFET_GATE_10uA.n15 56.2338
R80 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.n2 56.2338
R81 bgr_11_0.PFET_GATE_10uA.n3 bgr_11_0.PFET_GATE_10uA.n1 56.2338
R82 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n21 56.2338
R83 bgr_11_0.PFET_GATE_10uA.n25 bgr_11_0.PFET_GATE_10uA.n24 56.2338
R84 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t5 39.4005
R85 bgr_11_0.PFET_GATE_10uA.n11 bgr_11_0.PFET_GATE_10uA.t2 39.4005
R86 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t7 39.4005
R87 bgr_11_0.PFET_GATE_10uA.n9 bgr_11_0.PFET_GATE_10uA.t9 39.4005
R88 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.t8 39.4005
R89 bgr_11_0.PFET_GATE_10uA.n7 bgr_11_0.PFET_GATE_10uA.t4 39.4005
R90 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.t3 39.4005
R91 bgr_11_0.PFET_GATE_10uA.n5 bgr_11_0.PFET_GATE_10uA.t6 39.4005
R92 bgr_11_0.PFET_GATE_10uA.n18 bgr_11_0.PFET_GATE_10uA.n14 10.3755
R93 bgr_11_0.PFET_GATE_10uA.n13 bgr_11_0.PFET_GATE_10uA.n12 6.15675
R94 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n4 2.28175
R95 bgr_11_0.PFET_GATE_10uA bgr_11_0.PFET_GATE_10uA.n18 2.28175
R96 bgr_11_0.PFET_GATE_10uA.n14 bgr_11_0.PFET_GATE_10uA.n13 1.54738
R97 bgr_11_0.PFET_GATE_10uA.n8 bgr_11_0.PFET_GATE_10uA.n6 1.1255
R98 bgr_11_0.PFET_GATE_10uA.n10 bgr_11_0.PFET_GATE_10uA.n8 1.1255
R99 bgr_11_0.PFET_GATE_10uA.n12 bgr_11_0.PFET_GATE_10uA.n10 1.1255
R100 VDDA.n296 VDDA.n281 2100
R101 VDDA.n294 VDDA.n281 2070
R102 VDDA.n296 VDDA.n282 1830
R103 VDDA.n294 VDDA.n282 1800
R104 VDDA.n872 VDDA.t274 1231.74
R105 VDDA.n875 VDDA.t286 1231.74
R106 VDDA.n737 VDDA.t364 1231.74
R107 VDDA.n740 VDDA.t259 1231.74
R108 VDDA.n754 VDDA.t292 858.933
R109 VDDA.n799 VDDA.t336 858.933
R110 VDDA.n794 VDDA.t262 858.933
R111 VDDA.n188 VDDA.t325 858.933
R112 VDDA.t279 VDDA.n425 708.125
R113 VDDA.n448 VDDA.t279 708.125
R114 VDDA.n445 VDDA.t258 708.125
R115 VDDA.t258 VDDA.n426 708.125
R116 VDDA.t324 VDDA.n405 708.125
R117 VDDA.n458 VDDA.t324 708.125
R118 VDDA.n455 VDDA.t267 708.125
R119 VDDA.t267 VDDA.n406 708.125
R120 VDDA.t343 VDDA.n535 676.966
R121 VDDA.n765 VDDA.t253 661.375
R122 VDDA.n768 VDDA.t351 661.375
R123 VDDA.n816 VDDA.t316 661.375
R124 VDDA.n813 VDDA.t354 661.375
R125 VDDA.n202 VDDA.t319 661.375
R126 VDDA.n205 VDDA.t357 661.375
R127 VDDA.n447 VDDA.t278 657.76
R128 VDDA.n457 VDDA.t323 657.76
R129 VDDA.t281 VDDA.n565 648.726
R130 VDDA.n566 VDDA.t308 648.726
R131 VDDA.t272 VDDA.n552 648.726
R132 VDDA.n553 VDDA.t349 648.726
R133 VDDA.n536 VDDA.t299 643.038
R134 VDDA.n562 VDDA.t329 642.992
R135 VDDA.t305 VDDA.n561 642.992
R136 VDDA.n549 VDDA.t251 642.992
R137 VDDA.t314 VDDA.n548 642.992
R138 VDDA.n305 VDDA.t332 605.143
R139 VDDA.n285 VDDA.t295 589.076
R140 VDDA.n234 VDDA.t283 589.076
R141 VDDA.n237 VDDA.t289 589.076
R142 VDDA.n852 VDDA.t301 589.076
R143 VDDA.n849 VDDA.t310 589.076
R144 VDDA.n487 VDDA.n485 587.407
R145 VDDA.n491 VDDA.n488 587.407
R146 VDDA.n517 VDDA.n516 587.407
R147 VDDA.n512 VDDA.n478 587.407
R148 VDDA.n516 VDDA.n515 585
R149 VDDA.n514 VDDA.n512 585
R150 VDDA.n498 VDDA.n487 585
R151 VDDA.n495 VDDA.n488 585
R152 VDDA.t257 VDDA.n446 540.818
R153 VDDA.t266 VDDA.n456 540.818
R154 VDDA.t335 VDDA.n302 461.389
R155 VDDA.n303 VDDA.t335 461.389
R156 VDDA.n290 VDDA.t297 461.389
R157 VDDA.t297 VDDA.n289 461.389
R158 VDDA.n781 VDDA.t339 456.526
R159 VDDA.n778 VDDA.t360 456.526
R160 VDDA.n555 VDDA.t304 441.2
R161 VDDA.n563 VDDA.t328 441.2
R162 VDDA.n546 VDDA.t313 441.2
R163 VDDA.n550 VDDA.t250 441.2
R164 VDDA.n564 VDDA.t280 418.368
R165 VDDA.n567 VDDA.t307 418.368
R166 VDDA.n551 VDDA.t271 418.368
R167 VDDA.n554 VDDA.t348 418.368
R168 VDDA.n537 VDDA.t298 413.084
R169 VDDA.n534 VDDA.t342 413.084
R170 VDDA.t278 VDDA.t206 407.144
R171 VDDA.t206 VDDA.t99 407.144
R172 VDDA.t99 VDDA.t20 407.144
R173 VDDA.t20 VDDA.t170 407.144
R174 VDDA.t170 VDDA.t12 407.144
R175 VDDA.t12 VDDA.t210 407.144
R176 VDDA.t210 VDDA.t202 407.144
R177 VDDA.t202 VDDA.t192 407.144
R178 VDDA.t192 VDDA.t56 407.144
R179 VDDA.t56 VDDA.t178 407.144
R180 VDDA.t178 VDDA.t77 407.144
R181 VDDA.t77 VDDA.t208 407.144
R182 VDDA.t208 VDDA.t200 407.144
R183 VDDA.t200 VDDA.t382 407.144
R184 VDDA.t382 VDDA.t405 407.144
R185 VDDA.t405 VDDA.t389 407.144
R186 VDDA.t389 VDDA.t157 407.144
R187 VDDA.t157 VDDA.t204 407.144
R188 VDDA.t204 VDDA.t257 407.144
R189 VDDA.t323 VDDA.t150 407.144
R190 VDDA.t150 VDDA.t384 407.144
R191 VDDA.t384 VDDA.t165 407.144
R192 VDDA.t165 VDDA.t172 407.144
R193 VDDA.t172 VDDA.t163 407.144
R194 VDDA.t163 VDDA.t40 407.144
R195 VDDA.t40 VDDA.t47 407.144
R196 VDDA.t47 VDDA.t180 407.144
R197 VDDA.t180 VDDA.t18 407.144
R198 VDDA.t18 VDDA.t79 407.144
R199 VDDA.t79 VDDA.t413 407.144
R200 VDDA.t413 VDDA.t136 407.144
R201 VDDA.t136 VDDA.t190 407.144
R202 VDDA.t190 VDDA.t395 407.144
R203 VDDA.t395 VDDA.t10 407.144
R204 VDDA.t10 VDDA.t49 407.144
R205 VDDA.t49 VDDA.t67 407.144
R206 VDDA.t67 VDDA.t176 407.144
R207 VDDA.t176 VDDA.t266 407.144
R208 VDDA.n780 VDDA.t340 397.784
R209 VDDA.t361 VDDA.n779 397.784
R210 VDDA.t248 VDDA.t281 373.214
R211 VDDA.t238 VDDA.t248 373.214
R212 VDDA.t226 VDDA.t238 373.214
R213 VDDA.t246 VDDA.t226 373.214
R214 VDDA.t308 VDDA.t246 373.214
R215 VDDA.t224 VDDA.t305 373.214
R216 VDDA.t244 VDDA.t224 373.214
R217 VDDA.t236 VDDA.t244 373.214
R218 VDDA.t222 VDDA.t236 373.214
R219 VDDA.t240 VDDA.t222 373.214
R220 VDDA.t230 VDDA.t240 373.214
R221 VDDA.t232 VDDA.t230 373.214
R222 VDDA.t214 VDDA.t232 373.214
R223 VDDA.t329 VDDA.t214 373.214
R224 VDDA.t220 VDDA.t272 373.214
R225 VDDA.t242 VDDA.t220 373.214
R226 VDDA.t234 VDDA.t242 373.214
R227 VDDA.t218 VDDA.t234 373.214
R228 VDDA.t349 VDDA.t218 373.214
R229 VDDA.t228 VDDA.t314 373.214
R230 VDDA.t212 VDDA.t228 373.214
R231 VDDA.t251 VDDA.t212 373.214
R232 VDDA.t299 VDDA.t169 373.214
R233 VDDA.t169 VDDA.t162 373.214
R234 VDDA.t162 VDDA.t343 373.214
R235 VDDA.n450 VDDA.t277 370.168
R236 VDDA.n443 VDDA.t256 370.168
R237 VDDA.n460 VDDA.t322 370.168
R238 VDDA.n453 VDDA.t265 370.168
R239 VDDA.n469 VDDA.t268 360.868
R240 VDDA.n523 VDDA.t345 360.868
R241 VDDA.n562 VDDA.t331 354.154
R242 VDDA.n561 VDDA.t306 354.154
R243 VDDA.n549 VDDA.t252 354.154
R244 VDDA.n548 VDDA.t315 354.154
R245 VDDA.n536 VDDA.t300 354.063
R246 VDDA.n535 VDDA.t344 347.224
R247 VDDA.t284 VDDA.n235 343.882
R248 VDDA.n236 VDDA.t290 343.882
R249 VDDA.n851 VDDA.t302 343.882
R250 VDDA.t311 VDDA.n850 343.882
R251 VDDA.n574 VDDA.n560 336.341
R252 VDDA.n575 VDDA.n559 336.341
R253 VDDA.n576 VDDA.n558 336.341
R254 VDDA.n577 VDDA.n557 336.341
R255 VDDA.n578 VDDA.n556 336.341
R256 VDDA.n587 VDDA.n547 336.341
R257 VDDA.n565 VDDA.t282 331.901
R258 VDDA.n566 VDDA.t309 331.901
R259 VDDA.n552 VDDA.t273 331.901
R260 VDDA.n553 VDDA.t350 331.901
R261 VDDA.n442 VDDA.n441 299.231
R262 VDDA.n440 VDDA.n439 299.231
R263 VDDA.n438 VDDA.n437 299.231
R264 VDDA.n436 VDDA.n435 299.231
R265 VDDA.n434 VDDA.n433 299.231
R266 VDDA.n432 VDDA.n431 299.231
R267 VDDA.n430 VDDA.n429 299.231
R268 VDDA.n428 VDDA.n427 299.231
R269 VDDA.n424 VDDA.n423 299.231
R270 VDDA.n422 VDDA.n421 299.231
R271 VDDA.n420 VDDA.n419 299.231
R272 VDDA.n418 VDDA.n417 299.231
R273 VDDA.n416 VDDA.n415 299.231
R274 VDDA.n414 VDDA.n413 299.231
R275 VDDA.n412 VDDA.n411 299.231
R276 VDDA.n410 VDDA.n409 299.231
R277 VDDA.n408 VDDA.n407 299.231
R278 VDDA.n404 VDDA.n403 299.231
R279 VDDA.n569 VDDA.n568 299.053
R280 VDDA.n571 VDDA.n570 299.053
R281 VDDA.n582 VDDA.n581 299.053
R282 VDDA.n584 VDDA.n583 299.053
R283 VDDA.n753 VDDA.t293 282.788
R284 VDDA.n798 VDDA.t337 282.788
R285 VDDA.t296 VDDA.n294 279.298
R286 VDDA.n296 VDDA.t333 279.298
R287 VDDA.t340 VDDA.t194 259.091
R288 VDDA.t194 VDDA.t361 259.091
R289 VDDA.t33 VDDA.t269 251.471
R290 VDDA.t119 VDDA.t33 251.471
R291 VDDA.t419 VDDA.t119 251.471
R292 VDDA.t397 VDDA.t419 251.471
R293 VDDA.t121 VDDA.t397 251.471
R294 VDDA.t403 VDDA.t121 251.471
R295 VDDA.t416 VDDA.t403 251.471
R296 VDDA.t139 VDDA.t416 251.471
R297 VDDA.t143 VDDA.t139 251.471
R298 VDDA.t31 VDDA.t143 251.471
R299 VDDA.t370 VDDA.t31 251.471
R300 VDDA.t401 VDDA.t370 251.471
R301 VDDA.t399 VDDA.t401 251.471
R302 VDDA.t70 VDDA.t399 251.471
R303 VDDA.t130 VDDA.t70 251.471
R304 VDDA.t160 VDDA.t130 251.471
R305 VDDA.t346 VDDA.t160 251.471
R306 VDDA.n519 VDDA.n518 238.367
R307 VDDA.n446 VDDA.n445 238.367
R308 VDDA.n446 VDDA.n426 238.367
R309 VDDA.n456 VDDA.n455 238.367
R310 VDDA.n456 VDDA.n406 238.367
R311 VDDA.t269 VDDA.n503 237.5
R312 VDDA.n520 VDDA.t346 237.5
R313 VDDA.n187 VDDA.n186 222.524
R314 VDDA.n757 VDDA.n756 222.524
R315 VDDA.n797 VDDA.t326 221.121
R316 VDDA.t263 VDDA.n797 221.121
R317 VDDA.t156 VDDA.t284 217.708
R318 VDDA.t187 VDDA.t156 217.708
R319 VDDA.t45 VDDA.t187 217.708
R320 VDDA.t123 VDDA.t45 217.708
R321 VDDA.t37 VDDA.t123 217.708
R322 VDDA.t134 VDDA.t37 217.708
R323 VDDA.t186 VDDA.t134 217.708
R324 VDDA.t106 VDDA.t186 217.708
R325 VDDA.t76 VDDA.t106 217.708
R326 VDDA.t103 VDDA.t76 217.708
R327 VDDA.t290 VDDA.t103 217.708
R328 VDDA.t302 VDDA.t113 217.708
R329 VDDA.t113 VDDA.t183 217.708
R330 VDDA.t183 VDDA.t88 217.708
R331 VDDA.t88 VDDA.t185 217.708
R332 VDDA.t185 VDDA.t75 217.708
R333 VDDA.t75 VDDA.t116 217.708
R334 VDDA.t116 VDDA.t66 217.708
R335 VDDA.t66 VDDA.t110 217.708
R336 VDDA.t110 VDDA.t125 217.708
R337 VDDA.t125 VDDA.t182 217.708
R338 VDDA.t182 VDDA.t311 217.708
R339 VDDA.t254 VDDA.n766 213.131
R340 VDDA.n767 VDDA.t352 213.131
R341 VDDA.n815 VDDA.t317 213.131
R342 VDDA.t355 VDDA.n814 213.131
R343 VDDA.t320 VDDA.n203 213.131
R344 VDDA.n204 VDDA.t358 213.131
R345 VDDA.n297 VDDA.n280 195.201
R346 VDDA.n293 VDDA.n280 192
R347 VDDA.n508 VDDA.n506 185
R348 VDDA.n515 VDDA.n505 185
R349 VDDA.n520 VDDA.n505 185
R350 VDDA.n514 VDDA.n513 185
R351 VDDA.n511 VDDA.n480 185
R352 VDDA.n522 VDDA.n521 185
R353 VDDA.n521 VDDA.n520 185
R354 VDDA.n502 VDDA.n501 185
R355 VDDA.n503 VDDA.n502 185
R356 VDDA.n499 VDDA.n484 185
R357 VDDA.n498 VDDA.n497 185
R358 VDDA.n496 VDDA.n495 185
R359 VDDA.n490 VDDA.n489 185
R360 VDDA.n492 VDDA.n483 185
R361 VDDA.n503 VDDA.n483 185
R362 VDDA.t293 VDDA.t42 180.173
R363 VDDA.t42 VDDA.t188 180.173
R364 VDDA.t188 VDDA.t174 180.173
R365 VDDA.t174 VDDA.t138 180.173
R366 VDDA.t138 VDDA.t326 180.173
R367 VDDA.t407 VDDA.t263 180.173
R368 VDDA.t16 VDDA.t407 180.173
R369 VDDA.t132 VDDA.t16 180.173
R370 VDDA.t22 VDDA.t132 180.173
R371 VDDA.t337 VDDA.t22 180.173
R372 VDDA.n780 VDDA.t341 168.139
R373 VDDA.n779 VDDA.t363 168.139
R374 VDDA.n298 VDDA.n297 163.201
R375 VDDA.n293 VDDA.n292 163.201
R376 VDDA.n777 VDDA.n776 150.643
R377 VDDA.n276 VDDA.n275 150.558
R378 VDDA.n506 VDDA.n505 150
R379 VDDA.n513 VDDA.n505 150
R380 VDDA.n521 VDDA.n480 150
R381 VDDA.n502 VDDA.n484 150
R382 VDDA.n497 VDDA.n496 150
R383 VDDA.n489 VDDA.n483 150
R384 VDDA.t38 VDDA.t254 146.155
R385 VDDA.t352 VDDA.t38 146.155
R386 VDDA.t317 VDDA.t62 146.155
R387 VDDA.t62 VDDA.t91 146.155
R388 VDDA.t91 VDDA.t54 146.155
R389 VDDA.t54 VDDA.t58 146.155
R390 VDDA.t58 VDDA.t198 146.155
R391 VDDA.t198 VDDA.t380 146.155
R392 VDDA.t380 VDDA.t52 146.155
R393 VDDA.t52 VDDA.t97 146.155
R394 VDDA.t97 VDDA.t27 146.155
R395 VDDA.t27 VDDA.t95 146.155
R396 VDDA.t95 VDDA.t355 146.155
R397 VDDA.t378 VDDA.t320 146.155
R398 VDDA.t60 VDDA.t378 146.155
R399 VDDA.t29 VDDA.t60 146.155
R400 VDDA.t1 VDDA.t29 146.155
R401 VDDA.t196 VDDA.t1 146.155
R402 VDDA.t374 VDDA.t196 146.155
R403 VDDA.t89 VDDA.t374 146.155
R404 VDDA.t25 VDDA.t89 146.155
R405 VDDA.t376 VDDA.t25 146.155
R406 VDDA.t93 VDDA.t376 146.155
R407 VDDA.t358 VDDA.t93 146.155
R408 VDDA.n524 VDDA.n477 141.712
R409 VDDA.n525 VDDA.n476 141.712
R410 VDDA.n526 VDDA.n475 141.712
R411 VDDA.n527 VDDA.n474 141.712
R412 VDDA.n528 VDDA.n473 141.712
R413 VDDA.n529 VDDA.n472 141.712
R414 VDDA.n530 VDDA.n471 141.712
R415 VDDA.n531 VDDA.n470 141.712
R416 VDDA.n235 VDDA.t285 136.701
R417 VDDA.n236 VDDA.t291 136.701
R418 VDDA.n851 VDDA.t303 136.701
R419 VDDA.n850 VDDA.t312 136.701
R420 VDDA.t270 VDDA.n487 123.126
R421 VDDA.n488 VDDA.t270 123.126
R422 VDDA.n516 VDDA.t347 123.126
R423 VDDA.n512 VDDA.t347 123.126
R424 VDDA.t275 VDDA.n873 122.829
R425 VDDA.n874 VDDA.t287 122.829
R426 VDDA.t365 VDDA.n738 122.829
R427 VDDA.n739 VDDA.t260 122.829
R428 VDDA.t333 VDDA.t216 117.416
R429 VDDA.n753 VDDA.t294 113.26
R430 VDDA.n798 VDDA.t338 113.26
R431 VDDA.n796 VDDA.t264 113.26
R432 VDDA.n796 VDDA.t327 113.26
R433 VDDA.n295 VDDA.t296 112.079
R434 VDDA.n297 VDDA.n296 92.5005
R435 VDDA.n282 VDDA.n280 92.5005
R436 VDDA.n295 VDDA.n282 92.5005
R437 VDDA.n294 VDDA.n293 92.5005
R438 VDDA.n281 VDDA.n279 92.5005
R439 VDDA.n295 VDDA.n281 92.5005
R440 VDDA.n799 VDDA.n798 82.7434
R441 VDDA.n754 VDDA.n753 82.7434
R442 VDDA.t86 VDDA.t275 81.6411
R443 VDDA.t7 VDDA.t86 81.6411
R444 VDDA.t147 VDDA.t7 81.6411
R445 VDDA.t64 VDDA.t147 81.6411
R446 VDDA.t108 VDDA.t64 81.6411
R447 VDDA.t411 VDDA.t108 81.6411
R448 VDDA.t3 VDDA.t411 81.6411
R449 VDDA.t117 VDDA.t3 81.6411
R450 VDDA.t5 VDDA.t117 81.6411
R451 VDDA.t114 VDDA.t5 81.6411
R452 VDDA.t287 VDDA.t114 81.6411
R453 VDDA.t35 VDDA.t365 81.6411
R454 VDDA.t372 VDDA.t35 81.6411
R455 VDDA.t391 VDDA.t372 81.6411
R456 VDDA.t84 VDDA.t391 81.6411
R457 VDDA.t111 VDDA.t84 81.6411
R458 VDDA.t154 VDDA.t111 81.6411
R459 VDDA.t23 VDDA.t154 81.6411
R460 VDDA.t104 VDDA.t23 81.6411
R461 VDDA.t408 VDDA.t104 81.6411
R462 VDDA.t101 VDDA.t408 81.6411
R463 VDDA.t260 VDDA.t101 81.6411
R464 VDDA.n766 VDDA.t255 76.2576
R465 VDDA.n767 VDDA.t353 76.2576
R466 VDDA.n815 VDDA.t318 76.2576
R467 VDDA.n814 VDDA.t356 76.2576
R468 VDDA.n203 VDDA.t321 76.2576
R469 VDDA.n204 VDDA.t359 76.2576
R470 VDDA.n812 VDDA.n811 71.388
R471 VDDA.n810 VDDA.n809 71.388
R472 VDDA.n808 VDDA.n807 71.388
R473 VDDA.n806 VDDA.n805 71.388
R474 VDDA.n804 VDDA.n803 71.388
R475 VDDA.n193 VDDA.n192 71.388
R476 VDDA.n195 VDDA.n194 71.388
R477 VDDA.n197 VDDA.n196 71.388
R478 VDDA.n199 VDDA.n198 71.388
R479 VDDA.n201 VDDA.n200 71.388
R480 VDDA.n764 VDDA.n763 68.4557
R481 VDDA.n520 VDDA.n519 65.8183
R482 VDDA.n520 VDDA.n504 65.8183
R483 VDDA.n503 VDDA.n481 65.8183
R484 VDDA.n503 VDDA.n482 65.8183
R485 VDDA.n797 VDDA.n796 61.6672
R486 VDDA.n795 VDDA.n794 60.8005
R487 VDDA.n795 VDDA.n188 60.8005
R488 VDDA.n394 VDDA.t421 58.8005
R489 VDDA.n393 VDDA.t423 58.8005
R490 VDDA.n513 VDDA.n504 53.3664
R491 VDDA.n519 VDDA.n506 53.3664
R492 VDDA.n504 VDDA.n480 53.3664
R493 VDDA.n484 VDDA.n481 53.3664
R494 VDDA.n496 VDDA.n482 53.3664
R495 VDDA.n497 VDDA.n481 53.3664
R496 VDDA.n489 VDDA.n482 53.3664
R497 VDDA.n393 VDDA.t424 49.1638
R498 VDDA.n395 VDDA.t422 48.5162
R499 VDDA.n298 VDDA.n279 48.0005
R500 VDDA.n292 VDDA.n279 44.8005
R501 VDDA.n873 VDDA.t276 40.9789
R502 VDDA.n874 VDDA.t288 40.9789
R503 VDDA.n738 VDDA.t366 40.9789
R504 VDDA.n739 VDDA.t261 40.9789
R505 VDDA.n560 VDDA.t215 39.4005
R506 VDDA.n560 VDDA.t330 39.4005
R507 VDDA.n559 VDDA.t231 39.4005
R508 VDDA.n559 VDDA.t233 39.4005
R509 VDDA.n558 VDDA.t223 39.4005
R510 VDDA.n558 VDDA.t241 39.4005
R511 VDDA.n557 VDDA.t245 39.4005
R512 VDDA.n557 VDDA.t237 39.4005
R513 VDDA.t306 VDDA.n556 39.4005
R514 VDDA.n556 VDDA.t225 39.4005
R515 VDDA.n547 VDDA.t229 39.4005
R516 VDDA.n547 VDDA.t213 39.4005
R517 VDDA.n568 VDDA.t227 39.4005
R518 VDDA.n568 VDDA.t247 39.4005
R519 VDDA.n570 VDDA.t249 39.4005
R520 VDDA.n570 VDDA.t239 39.4005
R521 VDDA.n581 VDDA.t235 39.4005
R522 VDDA.n581 VDDA.t219 39.4005
R523 VDDA.n583 VDDA.t221 39.4005
R524 VDDA.n583 VDDA.t243 39.4005
R525 VDDA.n441 VDDA.t158 39.4005
R526 VDDA.n441 VDDA.t205 39.4005
R527 VDDA.n439 VDDA.t406 39.4005
R528 VDDA.n439 VDDA.t390 39.4005
R529 VDDA.n437 VDDA.t201 39.4005
R530 VDDA.n437 VDDA.t383 39.4005
R531 VDDA.n435 VDDA.t78 39.4005
R532 VDDA.n435 VDDA.t209 39.4005
R533 VDDA.n433 VDDA.t57 39.4005
R534 VDDA.n433 VDDA.t179 39.4005
R535 VDDA.n431 VDDA.t203 39.4005
R536 VDDA.n431 VDDA.t193 39.4005
R537 VDDA.n429 VDDA.t13 39.4005
R538 VDDA.n429 VDDA.t211 39.4005
R539 VDDA.n427 VDDA.t21 39.4005
R540 VDDA.n427 VDDA.t171 39.4005
R541 VDDA.n423 VDDA.t207 39.4005
R542 VDDA.n423 VDDA.t100 39.4005
R543 VDDA.n421 VDDA.t68 39.4005
R544 VDDA.n421 VDDA.t177 39.4005
R545 VDDA.n419 VDDA.t11 39.4005
R546 VDDA.n419 VDDA.t50 39.4005
R547 VDDA.n417 VDDA.t191 39.4005
R548 VDDA.n417 VDDA.t396 39.4005
R549 VDDA.n415 VDDA.t414 39.4005
R550 VDDA.n415 VDDA.t137 39.4005
R551 VDDA.n413 VDDA.t19 39.4005
R552 VDDA.n413 VDDA.t80 39.4005
R553 VDDA.n411 VDDA.t48 39.4005
R554 VDDA.n411 VDDA.t181 39.4005
R555 VDDA.n409 VDDA.t164 39.4005
R556 VDDA.n409 VDDA.t41 39.4005
R557 VDDA.n407 VDDA.t166 39.4005
R558 VDDA.n407 VDDA.t173 39.4005
R559 VDDA.n403 VDDA.t151 39.4005
R560 VDDA.n403 VDDA.t385 39.4005
R561 VDDA.n181 VDDA.n180 38.2695
R562 VDDA.n864 VDDA.n863 38.2695
R563 VDDA.n866 VDDA.n865 38.2695
R564 VDDA.n868 VDDA.n867 38.2695
R565 VDDA.n870 VDDA.n869 38.2695
R566 VDDA.n246 VDDA.n245 38.2695
R567 VDDA.n729 VDDA.n728 38.2695
R568 VDDA.n731 VDDA.n730 38.2695
R569 VDDA.n733 VDDA.n732 38.2695
R570 VDDA.n735 VDDA.n734 38.2695
R571 VDDA.n220 VDDA.n218 26.8887
R572 VDDA.n834 VDDA.n832 26.8887
R573 VDDA.n228 VDDA.n227 26.7741
R574 VDDA.n226 VDDA.n225 26.7741
R575 VDDA.n224 VDDA.n223 26.7741
R576 VDDA.n222 VDDA.n221 26.7741
R577 VDDA.n220 VDDA.n219 26.7741
R578 VDDA.n834 VDDA.n833 26.7741
R579 VDDA.n836 VDDA.n835 26.7741
R580 VDDA.n838 VDDA.n837 26.7741
R581 VDDA.n840 VDDA.n839 26.7741
R582 VDDA.n842 VDDA.n841 26.7741
R583 VDDA.n563 VDDA.n562 24.9931
R584 VDDA.n561 VDDA.n555 24.9931
R585 VDDA.n550 VDDA.n549 24.9931
R586 VDDA.n548 VDDA.n546 24.9931
R587 VDDA.n48 VDDA.t141 24.1029
R588 VDDA.n537 VDDA.n536 22.9536
R589 VDDA.n523 VDDA.n522 22.8576
R590 VDDA.n492 VDDA.n469 22.8576
R591 VDDA.n776 VDDA.t195 21.8894
R592 VDDA.n776 VDDA.t362 21.8894
R593 VDDA.n302 VDDA.n299 21.6365
R594 VDDA.n304 VDDA.n303 21.6365
R595 VDDA.n291 VDDA.n290 21.6365
R596 VDDA.n289 VDDA.n286 21.6365
R597 VDDA.n301 VDDA.n278 21.3338
R598 VDDA.n288 VDDA.n284 21.3338
R599 VDDA.n535 VDDA.n534 20.4312
R600 VDDA.n275 VDDA.t217 19.7005
R601 VDDA.n275 VDDA.t334 19.7005
R602 VDDA.n186 VDDA.t17 15.7605
R603 VDDA.n186 VDDA.t133 15.7605
R604 VDDA.n756 VDDA.t189 15.7605
R605 VDDA.n756 VDDA.t175 15.7605
R606 VDDA.n796 VDDA.n795 13.9641
R607 VDDA.n477 VDDA.t131 13.1338
R608 VDDA.n477 VDDA.t161 13.1338
R609 VDDA.n476 VDDA.t400 13.1338
R610 VDDA.n476 VDDA.t71 13.1338
R611 VDDA.n475 VDDA.t371 13.1338
R612 VDDA.n475 VDDA.t402 13.1338
R613 VDDA.n474 VDDA.t144 13.1338
R614 VDDA.n474 VDDA.t32 13.1338
R615 VDDA.n473 VDDA.t417 13.1338
R616 VDDA.n473 VDDA.t140 13.1338
R617 VDDA.n472 VDDA.t122 13.1338
R618 VDDA.n472 VDDA.t404 13.1338
R619 VDDA.n471 VDDA.t420 13.1338
R620 VDDA.n471 VDDA.t398 13.1338
R621 VDDA.n470 VDDA.t34 13.1338
R622 VDDA.n470 VDDA.t120 13.1338
R623 VDDA.n534 VDDA.n533 11.37
R624 VDDA.n538 VDDA.n537 11.37
R625 VDDA.t255 VDDA.n764 11.2576
R626 VDDA.n764 VDDA.t39 11.2576
R627 VDDA.n811 VDDA.t28 11.2576
R628 VDDA.n811 VDDA.t96 11.2576
R629 VDDA.n809 VDDA.t53 11.2576
R630 VDDA.n809 VDDA.t98 11.2576
R631 VDDA.n807 VDDA.t199 11.2576
R632 VDDA.n807 VDDA.t381 11.2576
R633 VDDA.n805 VDDA.t55 11.2576
R634 VDDA.n805 VDDA.t59 11.2576
R635 VDDA.n803 VDDA.t63 11.2576
R636 VDDA.n803 VDDA.t92 11.2576
R637 VDDA.n192 VDDA.t377 11.2576
R638 VDDA.n192 VDDA.t94 11.2576
R639 VDDA.n194 VDDA.t90 11.2576
R640 VDDA.n194 VDDA.t26 11.2576
R641 VDDA.n196 VDDA.t197 11.2576
R642 VDDA.n196 VDDA.t375 11.2576
R643 VDDA.n198 VDDA.t30 11.2576
R644 VDDA.n198 VDDA.t2 11.2576
R645 VDDA.n200 VDDA.t379 11.2576
R646 VDDA.n200 VDDA.t61 11.2576
R647 VDDA.n524 VDDA.n523 11.0575
R648 VDDA.n579 VDDA.n555 10.87
R649 VDDA.n588 VDDA.n546 10.87
R650 VDDA.n586 VDDA.n550 10.87
R651 VDDA.n573 VDDA.n563 10.87
R652 VDDA.n532 VDDA.n469 10.87
R653 VDDA.n755 VDDA.n754 10.8696
R654 VDDA.n800 VDDA.n799 10.869
R655 VDDA.n292 VDDA.n291 9.8005
R656 VDDA.n299 VDDA.n298 9.8005
R657 VDDA.n501 VDDA.n500 9.50883
R658 VDDA.n493 VDDA.n492 9.50883
R659 VDDA.n518 VDDA.n507 9.50883
R660 VDDA.n522 VDDA.n479 9.50883
R661 VDDA.n449 VDDA.n425 9.50883
R662 VDDA.n459 VDDA.n405 9.50883
R663 VDDA.n288 VDDA.n287 9.3005
R664 VDDA.n284 VDDA.n283 9.3005
R665 VDDA.n278 VDDA.n277 9.3005
R666 VDDA.n301 VDDA.n300 9.3005
R667 VDDA.n511 VDDA.n479 9.3005
R668 VDDA.n514 VDDA.n510 9.3005
R669 VDDA.n515 VDDA.n509 9.3005
R670 VDDA.n508 VDDA.n507 9.3005
R671 VDDA.n493 VDDA.n490 9.3005
R672 VDDA.n495 VDDA.n494 9.3005
R673 VDDA.n498 VDDA.n486 9.3005
R674 VDDA.n500 VDDA.n499 9.3005
R675 VDDA.n449 VDDA.n448 9.3005
R676 VDDA.n459 VDDA.n458 9.3005
R677 VDDA.n794 VDDA.n793 9.3005
R678 VDDA.n793 VDDA.n188 9.3005
R679 VDDA.n515 VDDA.n508 9.14336
R680 VDDA.n515 VDDA.n514 9.14336
R681 VDDA.n514 VDDA.n511 9.14336
R682 VDDA.n499 VDDA.n498 9.14336
R683 VDDA.n498 VDDA.n495 9.14336
R684 VDDA.n495 VDDA.n490 9.14336
R685 VDDA.n302 VDDA.n301 8.68224
R686 VDDA.n303 VDDA.n278 8.68224
R687 VDDA.n290 VDDA.n284 8.68224
R688 VDDA.n289 VDDA.n288 8.68224
R689 VDDA.n227 VDDA.t51 8.0005
R690 VDDA.n227 VDDA.t124 8.0005
R691 VDDA.n225 VDDA.t393 8.0005
R692 VDDA.n225 VDDA.t107 8.0005
R693 VDDA.n223 VDDA.t46 8.0005
R694 VDDA.n223 VDDA.t73 8.0005
R695 VDDA.n221 VDDA.t394 8.0005
R696 VDDA.n221 VDDA.t367 8.0005
R697 VDDA.n219 VDDA.t135 8.0005
R698 VDDA.n219 VDDA.t386 8.0005
R699 VDDA.n218 VDDA.t69 8.0005
R700 VDDA.n218 VDDA.t0 8.0005
R701 VDDA.n832 VDDA.t145 8.0005
R702 VDDA.n832 VDDA.t368 8.0005
R703 VDDA.n833 VDDA.t149 8.0005
R704 VDDA.n833 VDDA.t410 8.0005
R705 VDDA.n835 VDDA.t167 8.0005
R706 VDDA.n835 VDDA.t9 8.0005
R707 VDDA.n837 VDDA.t184 8.0005
R708 VDDA.n837 VDDA.t74 8.0005
R709 VDDA.n839 VDDA.t146 8.0005
R710 VDDA.n839 VDDA.t126 8.0005
R711 VDDA.n841 VDDA.t81 8.0005
R712 VDDA.n841 VDDA.t168 8.0005
R713 VDDA.n180 VDDA.t6 6.56717
R714 VDDA.n180 VDDA.t115 6.56717
R715 VDDA.n863 VDDA.t4 6.56717
R716 VDDA.n863 VDDA.t118 6.56717
R717 VDDA.n865 VDDA.t109 6.56717
R718 VDDA.n865 VDDA.t412 6.56717
R719 VDDA.n867 VDDA.t148 6.56717
R720 VDDA.n867 VDDA.t65 6.56717
R721 VDDA.n869 VDDA.t87 6.56717
R722 VDDA.n869 VDDA.t8 6.56717
R723 VDDA.n245 VDDA.t409 6.56717
R724 VDDA.n245 VDDA.t102 6.56717
R725 VDDA.n728 VDDA.t24 6.56717
R726 VDDA.n728 VDDA.t105 6.56717
R727 VDDA.n730 VDDA.t112 6.56717
R728 VDDA.n730 VDDA.t155 6.56717
R729 VDDA.n732 VDDA.t392 6.56717
R730 VDDA.n732 VDDA.t85 6.56717
R731 VDDA.n734 VDDA.t36 6.56717
R732 VDDA.n734 VDDA.t373 6.56717
R733 VDDA.t216 VDDA.n295 5.33758
R734 VDDA.n518 VDDA.n517 5.33286
R735 VDDA.n522 VDDA.n478 5.33286
R736 VDDA.n501 VDDA.n485 5.33286
R737 VDDA.n492 VDDA.n491 5.33286
R738 VDDA.n567 VDDA.n566 4.98383
R739 VDDA.n565 VDDA.n564 4.98383
R740 VDDA.n554 VDDA.n553 4.98383
R741 VDDA.n552 VDDA.n551 4.98383
R742 VDDA.n813 VDDA.n812 4.8755
R743 VDDA.n202 VDDA.n201 4.8755
R744 VDDA.n308 VDDA.n307 4.5005
R745 VDDA.n309 VDDA.n274 4.5005
R746 VDDA.n313 VDDA.n310 4.5005
R747 VDDA.n314 VDDA.n273 4.5005
R748 VDDA.n318 VDDA.n317 4.5005
R749 VDDA.n319 VDDA.n272 4.5005
R750 VDDA.n323 VDDA.n320 4.5005
R751 VDDA.n324 VDDA.n271 4.5005
R752 VDDA.n328 VDDA.n327 4.5005
R753 VDDA.n329 VDDA.n270 4.5005
R754 VDDA.n333 VDDA.n330 4.5005
R755 VDDA.n334 VDDA.n269 4.5005
R756 VDDA.n338 VDDA.n337 4.5005
R757 VDDA.n339 VDDA.n268 4.5005
R758 VDDA.n343 VDDA.n340 4.5005
R759 VDDA.n344 VDDA.n267 4.5005
R760 VDDA.n348 VDDA.n347 4.5005
R761 VDDA.n349 VDDA.n266 4.5005
R762 VDDA.n353 VDDA.n350 4.5005
R763 VDDA.n354 VDDA.n265 4.5005
R764 VDDA.n358 VDDA.n357 4.5005
R765 VDDA.n48 VDDA.n47 4.5005
R766 VDDA.n49 VDDA.n41 4.5005
R767 VDDA.n53 VDDA.n50 4.5005
R768 VDDA.n54 VDDA.n40 4.5005
R769 VDDA.n58 VDDA.n57 4.5005
R770 VDDA.n59 VDDA.n39 4.5005
R771 VDDA.n63 VDDA.n60 4.5005
R772 VDDA.n64 VDDA.n38 4.5005
R773 VDDA.n68 VDDA.n67 4.5005
R774 VDDA.n69 VDDA.n37 4.5005
R775 VDDA.n73 VDDA.n70 4.5005
R776 VDDA.n74 VDDA.n36 4.5005
R777 VDDA.n78 VDDA.n77 4.5005
R778 VDDA.n79 VDDA.n35 4.5005
R779 VDDA.n83 VDDA.n80 4.5005
R780 VDDA.n84 VDDA.n34 4.5005
R781 VDDA.n88 VDDA.n87 4.5005
R782 VDDA.n89 VDDA.n33 4.5005
R783 VDDA.n93 VDDA.n90 4.5005
R784 VDDA.n94 VDDA.n32 4.5005
R785 VDDA.n98 VDDA.n97 4.5005
R786 VDDA.n399 VDDA.n398 4.5005
R787 VDDA.n465 VDDA.n464 4.5005
R788 VDDA.n542 VDDA.n541 4.5005
R789 VDDA.n592 VDDA.n591 4.5005
R790 VDDA.n595 VDDA.n384 4.5005
R791 VDDA.n598 VDDA.n596 4.5005
R792 VDDA.n599 VDDA.n383 4.5005
R793 VDDA.n603 VDDA.n602 4.5005
R794 VDDA.n604 VDDA.n382 4.5005
R795 VDDA.n608 VDDA.n605 4.5005
R796 VDDA.n609 VDDA.n381 4.5005
R797 VDDA.n613 VDDA.n612 4.5005
R798 VDDA.n614 VDDA.n380 4.5005
R799 VDDA.n618 VDDA.n615 4.5005
R800 VDDA.n619 VDDA.n379 4.5005
R801 VDDA.n623 VDDA.n622 4.5005
R802 VDDA.n624 VDDA.n378 4.5005
R803 VDDA.n628 VDDA.n625 4.5005
R804 VDDA.n629 VDDA.n377 4.5005
R805 VDDA.n633 VDDA.n632 4.5005
R806 VDDA.n634 VDDA.n376 4.5005
R807 VDDA.n638 VDDA.n635 4.5005
R808 VDDA.n639 VDDA.n375 4.5005
R809 VDDA.n643 VDDA.n642 4.5005
R810 VDDA.n786 VDDA.n760 4.5005
R811 VDDA.n771 VDDA.n762 4.5005
R812 VDDA.n137 VDDA.n136 4.5005
R813 VDDA.n138 VDDA.n131 4.5005
R814 VDDA.n142 VDDA.n141 4.5005
R815 VDDA.n143 VDDA.n128 4.5005
R816 VDDA.n145 VDDA.n144 4.5005
R817 VDDA.n146 VDDA.n127 4.5005
R818 VDDA.n150 VDDA.n149 4.5005
R819 VDDA.n151 VDDA.n124 4.5005
R820 VDDA.n153 VDDA.n152 4.5005
R821 VDDA.n154 VDDA.n123 4.5005
R822 VDDA.n158 VDDA.n157 4.5005
R823 VDDA.n159 VDDA.n120 4.5005
R824 VDDA.n161 VDDA.n160 4.5005
R825 VDDA.n162 VDDA.n119 4.5005
R826 VDDA.n166 VDDA.n165 4.5005
R827 VDDA.n167 VDDA.n116 4.5005
R828 VDDA.n169 VDDA.n168 4.5005
R829 VDDA.n170 VDDA.n115 4.5005
R830 VDDA.n174 VDDA.n173 4.5005
R831 VDDA.n175 VDDA.n114 4.5005
R832 VDDA.n883 VDDA.n882 4.5005
R833 VDDA.n877 VDDA.n177 4.5005
R834 VDDA.n879 VDDA.n878 4.5005
R835 VDDA.n878 VDDA.n877 4.5005
R836 VDDA.n817 VDDA.n816 4.5005
R837 VDDA.n823 VDDA.n183 4.5005
R838 VDDA.n826 VDDA.n825 4.5005
R839 VDDA.n829 VDDA.n828 4.5005
R840 VDDA.n821 VDDA.n801 4.5005
R841 VDDA.n822 VDDA.n185 4.5005
R842 VDDA.n822 VDDA.n821 4.5005
R843 VDDA.n790 VDDA.n758 4.5005
R844 VDDA.n793 VDDA.n792 4.5005
R845 VDDA.n206 VDDA.n205 4.5005
R846 VDDA.n207 VDDA.n191 4.5005
R847 VDDA.n214 VDDA.n213 4.5005
R848 VDDA.n217 VDDA.n216 4.5005
R849 VDDA.n742 VDDA.n209 4.5005
R850 VDDA.n744 VDDA.n743 4.5005
R851 VDDA.n743 VDDA.n742 4.5005
R852 VDDA.n722 VDDA.n248 4.5005
R853 VDDA.n714 VDDA.n659 4.5005
R854 VDDA.n713 VDDA.n660 4.5005
R855 VDDA.n710 VDDA.n661 4.5005
R856 VDDA.n709 VDDA.n662 4.5005
R857 VDDA.n706 VDDA.n663 4.5005
R858 VDDA.n705 VDDA.n664 4.5005
R859 VDDA.n702 VDDA.n665 4.5005
R860 VDDA.n701 VDDA.n666 4.5005
R861 VDDA.n698 VDDA.n667 4.5005
R862 VDDA.n697 VDDA.n668 4.5005
R863 VDDA.n694 VDDA.n669 4.5005
R864 VDDA.n693 VDDA.n670 4.5005
R865 VDDA.n690 VDDA.n671 4.5005
R866 VDDA.n689 VDDA.n672 4.5005
R867 VDDA.n686 VDDA.n673 4.5005
R868 VDDA.n685 VDDA.n674 4.5005
R869 VDDA.n682 VDDA.n675 4.5005
R870 VDDA.n681 VDDA.n676 4.5005
R871 VDDA.n678 VDDA.n677 4.5005
R872 VDDA.n250 VDDA.n249 4.5005
R873 VDDA.n721 VDDA.n720 4.5005
R874 VDDA.n448 VDDA.n447 4.48641
R875 VDDA.n447 VDDA.n425 4.48641
R876 VDDA.n458 VDDA.n457 4.48641
R877 VDDA.n457 VDDA.n405 4.48641
R878 VDDA.n517 VDDA.n508 3.75335
R879 VDDA.n511 VDDA.n478 3.75335
R880 VDDA.n499 VDDA.n485 3.75335
R881 VDDA.n491 VDDA.n490 3.75335
R882 VDDA.n135 VDDA.n112 3.50398
R883 VDDA.n717 VDDA.n657 3.50398
R884 VDDA.n360 VDDA.n359 3.48392
R885 VDDA.n100 VDDA.n99 3.48334
R886 VDDA.n645 VDDA.n644 3.48334
R887 VDDA.n307 VDDA.n262 3.43627
R888 VDDA.n47 VDDA.n29 3.43627
R889 VDDA.n444 VDDA.n443 3.41464
R890 VDDA.n454 VDDA.n453 3.41464
R891 VDDA.n264 VDDA.n263 3.4105
R892 VDDA.n357 VDDA.n356 3.4105
R893 VDDA.n355 VDDA.n354 3.4105
R894 VDDA.n353 VDDA.n352 3.4105
R895 VDDA.n351 VDDA.n266 3.4105
R896 VDDA.n347 VDDA.n346 3.4105
R897 VDDA.n345 VDDA.n344 3.4105
R898 VDDA.n343 VDDA.n342 3.4105
R899 VDDA.n341 VDDA.n268 3.4105
R900 VDDA.n337 VDDA.n336 3.4105
R901 VDDA.n335 VDDA.n334 3.4105
R902 VDDA.n333 VDDA.n332 3.4105
R903 VDDA.n331 VDDA.n270 3.4105
R904 VDDA.n327 VDDA.n326 3.4105
R905 VDDA.n325 VDDA.n324 3.4105
R906 VDDA.n323 VDDA.n322 3.4105
R907 VDDA.n321 VDDA.n272 3.4105
R908 VDDA.n317 VDDA.n316 3.4105
R909 VDDA.n315 VDDA.n314 3.4105
R910 VDDA.n313 VDDA.n312 3.4105
R911 VDDA.n311 VDDA.n274 3.4105
R912 VDDA.n31 VDDA.n30 3.4105
R913 VDDA.n97 VDDA.n96 3.4105
R914 VDDA.n95 VDDA.n94 3.4105
R915 VDDA.n93 VDDA.n92 3.4105
R916 VDDA.n91 VDDA.n33 3.4105
R917 VDDA.n87 VDDA.n86 3.4105
R918 VDDA.n85 VDDA.n84 3.4105
R919 VDDA.n83 VDDA.n82 3.4105
R920 VDDA.n81 VDDA.n35 3.4105
R921 VDDA.n77 VDDA.n76 3.4105
R922 VDDA.n75 VDDA.n74 3.4105
R923 VDDA.n73 VDDA.n72 3.4105
R924 VDDA.n71 VDDA.n37 3.4105
R925 VDDA.n67 VDDA.n66 3.4105
R926 VDDA.n65 VDDA.n64 3.4105
R927 VDDA.n63 VDDA.n62 3.4105
R928 VDDA.n61 VDDA.n39 3.4105
R929 VDDA.n57 VDDA.n56 3.4105
R930 VDDA.n55 VDDA.n54 3.4105
R931 VDDA.n53 VDDA.n52 3.4105
R932 VDDA.n51 VDDA.n41 3.4105
R933 VDDA.n374 VDDA.n373 3.4105
R934 VDDA.n642 VDDA.n641 3.4105
R935 VDDA.n640 VDDA.n639 3.4105
R936 VDDA.n638 VDDA.n637 3.4105
R937 VDDA.n636 VDDA.n376 3.4105
R938 VDDA.n632 VDDA.n631 3.4105
R939 VDDA.n630 VDDA.n629 3.4105
R940 VDDA.n628 VDDA.n627 3.4105
R941 VDDA.n626 VDDA.n378 3.4105
R942 VDDA.n622 VDDA.n621 3.4105
R943 VDDA.n620 VDDA.n619 3.4105
R944 VDDA.n618 VDDA.n617 3.4105
R945 VDDA.n616 VDDA.n380 3.4105
R946 VDDA.n612 VDDA.n611 3.4105
R947 VDDA.n610 VDDA.n609 3.4105
R948 VDDA.n608 VDDA.n607 3.4105
R949 VDDA.n606 VDDA.n382 3.4105
R950 VDDA.n602 VDDA.n601 3.4105
R951 VDDA.n600 VDDA.n599 3.4105
R952 VDDA.n598 VDDA.n597 3.4105
R953 VDDA.n114 VDDA.n113 3.4105
R954 VDDA.n173 VDDA.n172 3.4105
R955 VDDA.n171 VDDA.n170 3.4105
R956 VDDA.n169 VDDA.n118 3.4105
R957 VDDA.n117 VDDA.n116 3.4105
R958 VDDA.n165 VDDA.n164 3.4105
R959 VDDA.n163 VDDA.n162 3.4105
R960 VDDA.n161 VDDA.n122 3.4105
R961 VDDA.n121 VDDA.n120 3.4105
R962 VDDA.n157 VDDA.n156 3.4105
R963 VDDA.n155 VDDA.n154 3.4105
R964 VDDA.n153 VDDA.n126 3.4105
R965 VDDA.n125 VDDA.n124 3.4105
R966 VDDA.n149 VDDA.n148 3.4105
R967 VDDA.n147 VDDA.n146 3.4105
R968 VDDA.n145 VDDA.n130 3.4105
R969 VDDA.n129 VDDA.n128 3.4105
R970 VDDA.n141 VDDA.n140 3.4105
R971 VDDA.n139 VDDA.n138 3.4105
R972 VDDA.n137 VDDA.n134 3.4105
R973 VDDA.n133 VDDA.n132 3.4105
R974 VDDA.n884 VDDA.n883 3.4105
R975 VDDA.n251 VDDA.n250 3.4105
R976 VDDA.n679 VDDA.n678 3.4105
R977 VDDA.n681 VDDA.n680 3.4105
R978 VDDA.n683 VDDA.n682 3.4105
R979 VDDA.n685 VDDA.n684 3.4105
R980 VDDA.n687 VDDA.n686 3.4105
R981 VDDA.n689 VDDA.n688 3.4105
R982 VDDA.n691 VDDA.n690 3.4105
R983 VDDA.n693 VDDA.n692 3.4105
R984 VDDA.n695 VDDA.n694 3.4105
R985 VDDA.n697 VDDA.n696 3.4105
R986 VDDA.n699 VDDA.n698 3.4105
R987 VDDA.n701 VDDA.n700 3.4105
R988 VDDA.n703 VDDA.n702 3.4105
R989 VDDA.n705 VDDA.n704 3.4105
R990 VDDA.n707 VDDA.n706 3.4105
R991 VDDA.n709 VDDA.n708 3.4105
R992 VDDA.n711 VDDA.n710 3.4105
R993 VDDA.n713 VDDA.n712 3.4105
R994 VDDA.n715 VDDA.n714 3.4105
R995 VDDA.n716 VDDA.n658 3.4105
R996 VDDA.n720 VDDA.n719 3.4105
R997 VDDA.n719 VDDA.n718 3.4105
R998 VDDA.n646 VDDA.n645 3.4105
R999 VDDA.n885 VDDA.n884 3.4105
R1000 VDDA.n101 VDDA.n100 3.4105
R1001 VDDA.n361 VDDA.n360 3.4105
R1002 VDDA.n1000 VDDA.n17 3.4105
R1003 VDDA.n1000 VDDA.n16 3.4105
R1004 VDDA.n1000 VDDA.n18 3.4105
R1005 VDDA.n1000 VDDA.n999 3.4105
R1006 VDDA.n999 VDDA.n904 3.4105
R1007 VDDA.n901 VDDA.n16 3.4105
R1008 VDDA.n969 VDDA.n901 3.4105
R1009 VDDA.n966 VDDA.n901 3.4105
R1010 VDDA.n971 VDDA.n901 3.4105
R1011 VDDA.n965 VDDA.n901 3.4105
R1012 VDDA.n973 VDDA.n901 3.4105
R1013 VDDA.n964 VDDA.n901 3.4105
R1014 VDDA.n975 VDDA.n901 3.4105
R1015 VDDA.n963 VDDA.n901 3.4105
R1016 VDDA.n977 VDDA.n901 3.4105
R1017 VDDA.n962 VDDA.n901 3.4105
R1018 VDDA.n979 VDDA.n901 3.4105
R1019 VDDA.n961 VDDA.n901 3.4105
R1020 VDDA.n981 VDDA.n901 3.4105
R1021 VDDA.n960 VDDA.n901 3.4105
R1022 VDDA.n983 VDDA.n901 3.4105
R1023 VDDA.n959 VDDA.n901 3.4105
R1024 VDDA.n985 VDDA.n901 3.4105
R1025 VDDA.n958 VDDA.n901 3.4105
R1026 VDDA.n987 VDDA.n901 3.4105
R1027 VDDA.n957 VDDA.n901 3.4105
R1028 VDDA.n989 VDDA.n901 3.4105
R1029 VDDA.n956 VDDA.n901 3.4105
R1030 VDDA.n991 VDDA.n901 3.4105
R1031 VDDA.n955 VDDA.n901 3.4105
R1032 VDDA.n993 VDDA.n901 3.4105
R1033 VDDA.n954 VDDA.n901 3.4105
R1034 VDDA.n995 VDDA.n901 3.4105
R1035 VDDA.n953 VDDA.n901 3.4105
R1036 VDDA.n997 VDDA.n901 3.4105
R1037 VDDA.n952 VDDA.n901 3.4105
R1038 VDDA.n901 VDDA.n18 3.4105
R1039 VDDA.n999 VDDA.n901 3.4105
R1040 VDDA.n907 VDDA.n16 3.4105
R1041 VDDA.n969 VDDA.n907 3.4105
R1042 VDDA.n966 VDDA.n907 3.4105
R1043 VDDA.n971 VDDA.n907 3.4105
R1044 VDDA.n965 VDDA.n907 3.4105
R1045 VDDA.n973 VDDA.n907 3.4105
R1046 VDDA.n964 VDDA.n907 3.4105
R1047 VDDA.n975 VDDA.n907 3.4105
R1048 VDDA.n963 VDDA.n907 3.4105
R1049 VDDA.n977 VDDA.n907 3.4105
R1050 VDDA.n962 VDDA.n907 3.4105
R1051 VDDA.n979 VDDA.n907 3.4105
R1052 VDDA.n961 VDDA.n907 3.4105
R1053 VDDA.n981 VDDA.n907 3.4105
R1054 VDDA.n960 VDDA.n907 3.4105
R1055 VDDA.n983 VDDA.n907 3.4105
R1056 VDDA.n959 VDDA.n907 3.4105
R1057 VDDA.n985 VDDA.n907 3.4105
R1058 VDDA.n958 VDDA.n907 3.4105
R1059 VDDA.n987 VDDA.n907 3.4105
R1060 VDDA.n957 VDDA.n907 3.4105
R1061 VDDA.n989 VDDA.n907 3.4105
R1062 VDDA.n956 VDDA.n907 3.4105
R1063 VDDA.n991 VDDA.n907 3.4105
R1064 VDDA.n955 VDDA.n907 3.4105
R1065 VDDA.n993 VDDA.n907 3.4105
R1066 VDDA.n954 VDDA.n907 3.4105
R1067 VDDA.n995 VDDA.n907 3.4105
R1068 VDDA.n953 VDDA.n907 3.4105
R1069 VDDA.n997 VDDA.n907 3.4105
R1070 VDDA.n952 VDDA.n907 3.4105
R1071 VDDA.n907 VDDA.n18 3.4105
R1072 VDDA.n999 VDDA.n907 3.4105
R1073 VDDA.n900 VDDA.n16 3.4105
R1074 VDDA.n969 VDDA.n900 3.4105
R1075 VDDA.n966 VDDA.n900 3.4105
R1076 VDDA.n971 VDDA.n900 3.4105
R1077 VDDA.n965 VDDA.n900 3.4105
R1078 VDDA.n973 VDDA.n900 3.4105
R1079 VDDA.n964 VDDA.n900 3.4105
R1080 VDDA.n975 VDDA.n900 3.4105
R1081 VDDA.n963 VDDA.n900 3.4105
R1082 VDDA.n977 VDDA.n900 3.4105
R1083 VDDA.n962 VDDA.n900 3.4105
R1084 VDDA.n979 VDDA.n900 3.4105
R1085 VDDA.n961 VDDA.n900 3.4105
R1086 VDDA.n981 VDDA.n900 3.4105
R1087 VDDA.n960 VDDA.n900 3.4105
R1088 VDDA.n983 VDDA.n900 3.4105
R1089 VDDA.n959 VDDA.n900 3.4105
R1090 VDDA.n985 VDDA.n900 3.4105
R1091 VDDA.n958 VDDA.n900 3.4105
R1092 VDDA.n987 VDDA.n900 3.4105
R1093 VDDA.n957 VDDA.n900 3.4105
R1094 VDDA.n989 VDDA.n900 3.4105
R1095 VDDA.n956 VDDA.n900 3.4105
R1096 VDDA.n991 VDDA.n900 3.4105
R1097 VDDA.n955 VDDA.n900 3.4105
R1098 VDDA.n993 VDDA.n900 3.4105
R1099 VDDA.n954 VDDA.n900 3.4105
R1100 VDDA.n995 VDDA.n900 3.4105
R1101 VDDA.n953 VDDA.n900 3.4105
R1102 VDDA.n997 VDDA.n900 3.4105
R1103 VDDA.n952 VDDA.n900 3.4105
R1104 VDDA.n900 VDDA.n18 3.4105
R1105 VDDA.n999 VDDA.n900 3.4105
R1106 VDDA.n910 VDDA.n16 3.4105
R1107 VDDA.n969 VDDA.n910 3.4105
R1108 VDDA.n966 VDDA.n910 3.4105
R1109 VDDA.n971 VDDA.n910 3.4105
R1110 VDDA.n965 VDDA.n910 3.4105
R1111 VDDA.n973 VDDA.n910 3.4105
R1112 VDDA.n964 VDDA.n910 3.4105
R1113 VDDA.n975 VDDA.n910 3.4105
R1114 VDDA.n963 VDDA.n910 3.4105
R1115 VDDA.n977 VDDA.n910 3.4105
R1116 VDDA.n962 VDDA.n910 3.4105
R1117 VDDA.n979 VDDA.n910 3.4105
R1118 VDDA.n961 VDDA.n910 3.4105
R1119 VDDA.n981 VDDA.n910 3.4105
R1120 VDDA.n960 VDDA.n910 3.4105
R1121 VDDA.n983 VDDA.n910 3.4105
R1122 VDDA.n959 VDDA.n910 3.4105
R1123 VDDA.n985 VDDA.n910 3.4105
R1124 VDDA.n958 VDDA.n910 3.4105
R1125 VDDA.n987 VDDA.n910 3.4105
R1126 VDDA.n957 VDDA.n910 3.4105
R1127 VDDA.n989 VDDA.n910 3.4105
R1128 VDDA.n956 VDDA.n910 3.4105
R1129 VDDA.n991 VDDA.n910 3.4105
R1130 VDDA.n955 VDDA.n910 3.4105
R1131 VDDA.n993 VDDA.n910 3.4105
R1132 VDDA.n954 VDDA.n910 3.4105
R1133 VDDA.n995 VDDA.n910 3.4105
R1134 VDDA.n953 VDDA.n910 3.4105
R1135 VDDA.n997 VDDA.n910 3.4105
R1136 VDDA.n952 VDDA.n910 3.4105
R1137 VDDA.n910 VDDA.n18 3.4105
R1138 VDDA.n999 VDDA.n910 3.4105
R1139 VDDA.n899 VDDA.n16 3.4105
R1140 VDDA.n969 VDDA.n899 3.4105
R1141 VDDA.n966 VDDA.n899 3.4105
R1142 VDDA.n971 VDDA.n899 3.4105
R1143 VDDA.n965 VDDA.n899 3.4105
R1144 VDDA.n973 VDDA.n899 3.4105
R1145 VDDA.n964 VDDA.n899 3.4105
R1146 VDDA.n975 VDDA.n899 3.4105
R1147 VDDA.n963 VDDA.n899 3.4105
R1148 VDDA.n977 VDDA.n899 3.4105
R1149 VDDA.n962 VDDA.n899 3.4105
R1150 VDDA.n979 VDDA.n899 3.4105
R1151 VDDA.n961 VDDA.n899 3.4105
R1152 VDDA.n981 VDDA.n899 3.4105
R1153 VDDA.n960 VDDA.n899 3.4105
R1154 VDDA.n983 VDDA.n899 3.4105
R1155 VDDA.n959 VDDA.n899 3.4105
R1156 VDDA.n985 VDDA.n899 3.4105
R1157 VDDA.n958 VDDA.n899 3.4105
R1158 VDDA.n987 VDDA.n899 3.4105
R1159 VDDA.n957 VDDA.n899 3.4105
R1160 VDDA.n989 VDDA.n899 3.4105
R1161 VDDA.n956 VDDA.n899 3.4105
R1162 VDDA.n991 VDDA.n899 3.4105
R1163 VDDA.n955 VDDA.n899 3.4105
R1164 VDDA.n993 VDDA.n899 3.4105
R1165 VDDA.n954 VDDA.n899 3.4105
R1166 VDDA.n995 VDDA.n899 3.4105
R1167 VDDA.n953 VDDA.n899 3.4105
R1168 VDDA.n997 VDDA.n899 3.4105
R1169 VDDA.n952 VDDA.n899 3.4105
R1170 VDDA.n899 VDDA.n18 3.4105
R1171 VDDA.n999 VDDA.n899 3.4105
R1172 VDDA.n913 VDDA.n16 3.4105
R1173 VDDA.n969 VDDA.n913 3.4105
R1174 VDDA.n966 VDDA.n913 3.4105
R1175 VDDA.n971 VDDA.n913 3.4105
R1176 VDDA.n965 VDDA.n913 3.4105
R1177 VDDA.n973 VDDA.n913 3.4105
R1178 VDDA.n964 VDDA.n913 3.4105
R1179 VDDA.n975 VDDA.n913 3.4105
R1180 VDDA.n963 VDDA.n913 3.4105
R1181 VDDA.n977 VDDA.n913 3.4105
R1182 VDDA.n962 VDDA.n913 3.4105
R1183 VDDA.n979 VDDA.n913 3.4105
R1184 VDDA.n961 VDDA.n913 3.4105
R1185 VDDA.n981 VDDA.n913 3.4105
R1186 VDDA.n960 VDDA.n913 3.4105
R1187 VDDA.n983 VDDA.n913 3.4105
R1188 VDDA.n959 VDDA.n913 3.4105
R1189 VDDA.n985 VDDA.n913 3.4105
R1190 VDDA.n958 VDDA.n913 3.4105
R1191 VDDA.n987 VDDA.n913 3.4105
R1192 VDDA.n957 VDDA.n913 3.4105
R1193 VDDA.n989 VDDA.n913 3.4105
R1194 VDDA.n956 VDDA.n913 3.4105
R1195 VDDA.n991 VDDA.n913 3.4105
R1196 VDDA.n955 VDDA.n913 3.4105
R1197 VDDA.n993 VDDA.n913 3.4105
R1198 VDDA.n954 VDDA.n913 3.4105
R1199 VDDA.n995 VDDA.n913 3.4105
R1200 VDDA.n953 VDDA.n913 3.4105
R1201 VDDA.n997 VDDA.n913 3.4105
R1202 VDDA.n952 VDDA.n913 3.4105
R1203 VDDA.n913 VDDA.n18 3.4105
R1204 VDDA.n999 VDDA.n913 3.4105
R1205 VDDA.n898 VDDA.n16 3.4105
R1206 VDDA.n969 VDDA.n898 3.4105
R1207 VDDA.n966 VDDA.n898 3.4105
R1208 VDDA.n971 VDDA.n898 3.4105
R1209 VDDA.n965 VDDA.n898 3.4105
R1210 VDDA.n973 VDDA.n898 3.4105
R1211 VDDA.n964 VDDA.n898 3.4105
R1212 VDDA.n975 VDDA.n898 3.4105
R1213 VDDA.n963 VDDA.n898 3.4105
R1214 VDDA.n977 VDDA.n898 3.4105
R1215 VDDA.n962 VDDA.n898 3.4105
R1216 VDDA.n979 VDDA.n898 3.4105
R1217 VDDA.n961 VDDA.n898 3.4105
R1218 VDDA.n981 VDDA.n898 3.4105
R1219 VDDA.n960 VDDA.n898 3.4105
R1220 VDDA.n983 VDDA.n898 3.4105
R1221 VDDA.n959 VDDA.n898 3.4105
R1222 VDDA.n985 VDDA.n898 3.4105
R1223 VDDA.n958 VDDA.n898 3.4105
R1224 VDDA.n987 VDDA.n898 3.4105
R1225 VDDA.n957 VDDA.n898 3.4105
R1226 VDDA.n989 VDDA.n898 3.4105
R1227 VDDA.n956 VDDA.n898 3.4105
R1228 VDDA.n991 VDDA.n898 3.4105
R1229 VDDA.n955 VDDA.n898 3.4105
R1230 VDDA.n993 VDDA.n898 3.4105
R1231 VDDA.n954 VDDA.n898 3.4105
R1232 VDDA.n995 VDDA.n898 3.4105
R1233 VDDA.n953 VDDA.n898 3.4105
R1234 VDDA.n997 VDDA.n898 3.4105
R1235 VDDA.n952 VDDA.n898 3.4105
R1236 VDDA.n898 VDDA.n18 3.4105
R1237 VDDA.n999 VDDA.n898 3.4105
R1238 VDDA.n916 VDDA.n16 3.4105
R1239 VDDA.n969 VDDA.n916 3.4105
R1240 VDDA.n966 VDDA.n916 3.4105
R1241 VDDA.n971 VDDA.n916 3.4105
R1242 VDDA.n965 VDDA.n916 3.4105
R1243 VDDA.n973 VDDA.n916 3.4105
R1244 VDDA.n964 VDDA.n916 3.4105
R1245 VDDA.n975 VDDA.n916 3.4105
R1246 VDDA.n963 VDDA.n916 3.4105
R1247 VDDA.n977 VDDA.n916 3.4105
R1248 VDDA.n962 VDDA.n916 3.4105
R1249 VDDA.n979 VDDA.n916 3.4105
R1250 VDDA.n961 VDDA.n916 3.4105
R1251 VDDA.n981 VDDA.n916 3.4105
R1252 VDDA.n960 VDDA.n916 3.4105
R1253 VDDA.n983 VDDA.n916 3.4105
R1254 VDDA.n959 VDDA.n916 3.4105
R1255 VDDA.n985 VDDA.n916 3.4105
R1256 VDDA.n958 VDDA.n916 3.4105
R1257 VDDA.n987 VDDA.n916 3.4105
R1258 VDDA.n957 VDDA.n916 3.4105
R1259 VDDA.n989 VDDA.n916 3.4105
R1260 VDDA.n956 VDDA.n916 3.4105
R1261 VDDA.n991 VDDA.n916 3.4105
R1262 VDDA.n955 VDDA.n916 3.4105
R1263 VDDA.n993 VDDA.n916 3.4105
R1264 VDDA.n954 VDDA.n916 3.4105
R1265 VDDA.n995 VDDA.n916 3.4105
R1266 VDDA.n953 VDDA.n916 3.4105
R1267 VDDA.n997 VDDA.n916 3.4105
R1268 VDDA.n952 VDDA.n916 3.4105
R1269 VDDA.n916 VDDA.n18 3.4105
R1270 VDDA.n999 VDDA.n916 3.4105
R1271 VDDA.n897 VDDA.n16 3.4105
R1272 VDDA.n969 VDDA.n897 3.4105
R1273 VDDA.n966 VDDA.n897 3.4105
R1274 VDDA.n971 VDDA.n897 3.4105
R1275 VDDA.n965 VDDA.n897 3.4105
R1276 VDDA.n973 VDDA.n897 3.4105
R1277 VDDA.n964 VDDA.n897 3.4105
R1278 VDDA.n975 VDDA.n897 3.4105
R1279 VDDA.n963 VDDA.n897 3.4105
R1280 VDDA.n977 VDDA.n897 3.4105
R1281 VDDA.n962 VDDA.n897 3.4105
R1282 VDDA.n979 VDDA.n897 3.4105
R1283 VDDA.n961 VDDA.n897 3.4105
R1284 VDDA.n981 VDDA.n897 3.4105
R1285 VDDA.n960 VDDA.n897 3.4105
R1286 VDDA.n983 VDDA.n897 3.4105
R1287 VDDA.n959 VDDA.n897 3.4105
R1288 VDDA.n985 VDDA.n897 3.4105
R1289 VDDA.n958 VDDA.n897 3.4105
R1290 VDDA.n987 VDDA.n897 3.4105
R1291 VDDA.n957 VDDA.n897 3.4105
R1292 VDDA.n989 VDDA.n897 3.4105
R1293 VDDA.n956 VDDA.n897 3.4105
R1294 VDDA.n991 VDDA.n897 3.4105
R1295 VDDA.n955 VDDA.n897 3.4105
R1296 VDDA.n993 VDDA.n897 3.4105
R1297 VDDA.n954 VDDA.n897 3.4105
R1298 VDDA.n995 VDDA.n897 3.4105
R1299 VDDA.n953 VDDA.n897 3.4105
R1300 VDDA.n997 VDDA.n897 3.4105
R1301 VDDA.n952 VDDA.n897 3.4105
R1302 VDDA.n897 VDDA.n18 3.4105
R1303 VDDA.n999 VDDA.n897 3.4105
R1304 VDDA.n919 VDDA.n16 3.4105
R1305 VDDA.n969 VDDA.n919 3.4105
R1306 VDDA.n966 VDDA.n919 3.4105
R1307 VDDA.n971 VDDA.n919 3.4105
R1308 VDDA.n965 VDDA.n919 3.4105
R1309 VDDA.n973 VDDA.n919 3.4105
R1310 VDDA.n964 VDDA.n919 3.4105
R1311 VDDA.n975 VDDA.n919 3.4105
R1312 VDDA.n963 VDDA.n919 3.4105
R1313 VDDA.n977 VDDA.n919 3.4105
R1314 VDDA.n962 VDDA.n919 3.4105
R1315 VDDA.n979 VDDA.n919 3.4105
R1316 VDDA.n961 VDDA.n919 3.4105
R1317 VDDA.n981 VDDA.n919 3.4105
R1318 VDDA.n960 VDDA.n919 3.4105
R1319 VDDA.n983 VDDA.n919 3.4105
R1320 VDDA.n959 VDDA.n919 3.4105
R1321 VDDA.n985 VDDA.n919 3.4105
R1322 VDDA.n958 VDDA.n919 3.4105
R1323 VDDA.n987 VDDA.n919 3.4105
R1324 VDDA.n957 VDDA.n919 3.4105
R1325 VDDA.n989 VDDA.n919 3.4105
R1326 VDDA.n956 VDDA.n919 3.4105
R1327 VDDA.n991 VDDA.n919 3.4105
R1328 VDDA.n955 VDDA.n919 3.4105
R1329 VDDA.n993 VDDA.n919 3.4105
R1330 VDDA.n954 VDDA.n919 3.4105
R1331 VDDA.n995 VDDA.n919 3.4105
R1332 VDDA.n953 VDDA.n919 3.4105
R1333 VDDA.n997 VDDA.n919 3.4105
R1334 VDDA.n952 VDDA.n919 3.4105
R1335 VDDA.n919 VDDA.n18 3.4105
R1336 VDDA.n999 VDDA.n919 3.4105
R1337 VDDA.n896 VDDA.n16 3.4105
R1338 VDDA.n969 VDDA.n896 3.4105
R1339 VDDA.n966 VDDA.n896 3.4105
R1340 VDDA.n971 VDDA.n896 3.4105
R1341 VDDA.n965 VDDA.n896 3.4105
R1342 VDDA.n973 VDDA.n896 3.4105
R1343 VDDA.n964 VDDA.n896 3.4105
R1344 VDDA.n975 VDDA.n896 3.4105
R1345 VDDA.n963 VDDA.n896 3.4105
R1346 VDDA.n977 VDDA.n896 3.4105
R1347 VDDA.n962 VDDA.n896 3.4105
R1348 VDDA.n979 VDDA.n896 3.4105
R1349 VDDA.n961 VDDA.n896 3.4105
R1350 VDDA.n981 VDDA.n896 3.4105
R1351 VDDA.n960 VDDA.n896 3.4105
R1352 VDDA.n983 VDDA.n896 3.4105
R1353 VDDA.n959 VDDA.n896 3.4105
R1354 VDDA.n985 VDDA.n896 3.4105
R1355 VDDA.n958 VDDA.n896 3.4105
R1356 VDDA.n987 VDDA.n896 3.4105
R1357 VDDA.n957 VDDA.n896 3.4105
R1358 VDDA.n989 VDDA.n896 3.4105
R1359 VDDA.n956 VDDA.n896 3.4105
R1360 VDDA.n991 VDDA.n896 3.4105
R1361 VDDA.n955 VDDA.n896 3.4105
R1362 VDDA.n993 VDDA.n896 3.4105
R1363 VDDA.n954 VDDA.n896 3.4105
R1364 VDDA.n995 VDDA.n896 3.4105
R1365 VDDA.n953 VDDA.n896 3.4105
R1366 VDDA.n997 VDDA.n896 3.4105
R1367 VDDA.n952 VDDA.n896 3.4105
R1368 VDDA.n896 VDDA.n18 3.4105
R1369 VDDA.n999 VDDA.n896 3.4105
R1370 VDDA.n922 VDDA.n16 3.4105
R1371 VDDA.n969 VDDA.n922 3.4105
R1372 VDDA.n966 VDDA.n922 3.4105
R1373 VDDA.n971 VDDA.n922 3.4105
R1374 VDDA.n965 VDDA.n922 3.4105
R1375 VDDA.n973 VDDA.n922 3.4105
R1376 VDDA.n964 VDDA.n922 3.4105
R1377 VDDA.n975 VDDA.n922 3.4105
R1378 VDDA.n963 VDDA.n922 3.4105
R1379 VDDA.n977 VDDA.n922 3.4105
R1380 VDDA.n962 VDDA.n922 3.4105
R1381 VDDA.n979 VDDA.n922 3.4105
R1382 VDDA.n961 VDDA.n922 3.4105
R1383 VDDA.n981 VDDA.n922 3.4105
R1384 VDDA.n960 VDDA.n922 3.4105
R1385 VDDA.n983 VDDA.n922 3.4105
R1386 VDDA.n959 VDDA.n922 3.4105
R1387 VDDA.n985 VDDA.n922 3.4105
R1388 VDDA.n958 VDDA.n922 3.4105
R1389 VDDA.n987 VDDA.n922 3.4105
R1390 VDDA.n957 VDDA.n922 3.4105
R1391 VDDA.n989 VDDA.n922 3.4105
R1392 VDDA.n956 VDDA.n922 3.4105
R1393 VDDA.n991 VDDA.n922 3.4105
R1394 VDDA.n955 VDDA.n922 3.4105
R1395 VDDA.n993 VDDA.n922 3.4105
R1396 VDDA.n954 VDDA.n922 3.4105
R1397 VDDA.n995 VDDA.n922 3.4105
R1398 VDDA.n953 VDDA.n922 3.4105
R1399 VDDA.n997 VDDA.n922 3.4105
R1400 VDDA.n952 VDDA.n922 3.4105
R1401 VDDA.n922 VDDA.n18 3.4105
R1402 VDDA.n999 VDDA.n922 3.4105
R1403 VDDA.n895 VDDA.n16 3.4105
R1404 VDDA.n969 VDDA.n895 3.4105
R1405 VDDA.n966 VDDA.n895 3.4105
R1406 VDDA.n971 VDDA.n895 3.4105
R1407 VDDA.n965 VDDA.n895 3.4105
R1408 VDDA.n973 VDDA.n895 3.4105
R1409 VDDA.n964 VDDA.n895 3.4105
R1410 VDDA.n975 VDDA.n895 3.4105
R1411 VDDA.n963 VDDA.n895 3.4105
R1412 VDDA.n977 VDDA.n895 3.4105
R1413 VDDA.n962 VDDA.n895 3.4105
R1414 VDDA.n979 VDDA.n895 3.4105
R1415 VDDA.n961 VDDA.n895 3.4105
R1416 VDDA.n981 VDDA.n895 3.4105
R1417 VDDA.n960 VDDA.n895 3.4105
R1418 VDDA.n983 VDDA.n895 3.4105
R1419 VDDA.n959 VDDA.n895 3.4105
R1420 VDDA.n985 VDDA.n895 3.4105
R1421 VDDA.n958 VDDA.n895 3.4105
R1422 VDDA.n987 VDDA.n895 3.4105
R1423 VDDA.n957 VDDA.n895 3.4105
R1424 VDDA.n989 VDDA.n895 3.4105
R1425 VDDA.n956 VDDA.n895 3.4105
R1426 VDDA.n991 VDDA.n895 3.4105
R1427 VDDA.n955 VDDA.n895 3.4105
R1428 VDDA.n993 VDDA.n895 3.4105
R1429 VDDA.n954 VDDA.n895 3.4105
R1430 VDDA.n995 VDDA.n895 3.4105
R1431 VDDA.n953 VDDA.n895 3.4105
R1432 VDDA.n997 VDDA.n895 3.4105
R1433 VDDA.n952 VDDA.n895 3.4105
R1434 VDDA.n895 VDDA.n18 3.4105
R1435 VDDA.n999 VDDA.n895 3.4105
R1436 VDDA.n925 VDDA.n16 3.4105
R1437 VDDA.n969 VDDA.n925 3.4105
R1438 VDDA.n966 VDDA.n925 3.4105
R1439 VDDA.n971 VDDA.n925 3.4105
R1440 VDDA.n965 VDDA.n925 3.4105
R1441 VDDA.n973 VDDA.n925 3.4105
R1442 VDDA.n964 VDDA.n925 3.4105
R1443 VDDA.n975 VDDA.n925 3.4105
R1444 VDDA.n963 VDDA.n925 3.4105
R1445 VDDA.n977 VDDA.n925 3.4105
R1446 VDDA.n962 VDDA.n925 3.4105
R1447 VDDA.n979 VDDA.n925 3.4105
R1448 VDDA.n961 VDDA.n925 3.4105
R1449 VDDA.n981 VDDA.n925 3.4105
R1450 VDDA.n960 VDDA.n925 3.4105
R1451 VDDA.n983 VDDA.n925 3.4105
R1452 VDDA.n959 VDDA.n925 3.4105
R1453 VDDA.n985 VDDA.n925 3.4105
R1454 VDDA.n958 VDDA.n925 3.4105
R1455 VDDA.n987 VDDA.n925 3.4105
R1456 VDDA.n957 VDDA.n925 3.4105
R1457 VDDA.n989 VDDA.n925 3.4105
R1458 VDDA.n956 VDDA.n925 3.4105
R1459 VDDA.n991 VDDA.n925 3.4105
R1460 VDDA.n955 VDDA.n925 3.4105
R1461 VDDA.n993 VDDA.n925 3.4105
R1462 VDDA.n954 VDDA.n925 3.4105
R1463 VDDA.n995 VDDA.n925 3.4105
R1464 VDDA.n953 VDDA.n925 3.4105
R1465 VDDA.n997 VDDA.n925 3.4105
R1466 VDDA.n952 VDDA.n925 3.4105
R1467 VDDA.n925 VDDA.n18 3.4105
R1468 VDDA.n999 VDDA.n925 3.4105
R1469 VDDA.n894 VDDA.n16 3.4105
R1470 VDDA.n969 VDDA.n894 3.4105
R1471 VDDA.n966 VDDA.n894 3.4105
R1472 VDDA.n971 VDDA.n894 3.4105
R1473 VDDA.n965 VDDA.n894 3.4105
R1474 VDDA.n973 VDDA.n894 3.4105
R1475 VDDA.n964 VDDA.n894 3.4105
R1476 VDDA.n975 VDDA.n894 3.4105
R1477 VDDA.n963 VDDA.n894 3.4105
R1478 VDDA.n977 VDDA.n894 3.4105
R1479 VDDA.n962 VDDA.n894 3.4105
R1480 VDDA.n979 VDDA.n894 3.4105
R1481 VDDA.n961 VDDA.n894 3.4105
R1482 VDDA.n981 VDDA.n894 3.4105
R1483 VDDA.n960 VDDA.n894 3.4105
R1484 VDDA.n983 VDDA.n894 3.4105
R1485 VDDA.n959 VDDA.n894 3.4105
R1486 VDDA.n985 VDDA.n894 3.4105
R1487 VDDA.n958 VDDA.n894 3.4105
R1488 VDDA.n987 VDDA.n894 3.4105
R1489 VDDA.n957 VDDA.n894 3.4105
R1490 VDDA.n989 VDDA.n894 3.4105
R1491 VDDA.n956 VDDA.n894 3.4105
R1492 VDDA.n991 VDDA.n894 3.4105
R1493 VDDA.n955 VDDA.n894 3.4105
R1494 VDDA.n993 VDDA.n894 3.4105
R1495 VDDA.n954 VDDA.n894 3.4105
R1496 VDDA.n995 VDDA.n894 3.4105
R1497 VDDA.n953 VDDA.n894 3.4105
R1498 VDDA.n997 VDDA.n894 3.4105
R1499 VDDA.n952 VDDA.n894 3.4105
R1500 VDDA.n894 VDDA.n18 3.4105
R1501 VDDA.n999 VDDA.n894 3.4105
R1502 VDDA.n928 VDDA.n16 3.4105
R1503 VDDA.n969 VDDA.n928 3.4105
R1504 VDDA.n966 VDDA.n928 3.4105
R1505 VDDA.n971 VDDA.n928 3.4105
R1506 VDDA.n965 VDDA.n928 3.4105
R1507 VDDA.n973 VDDA.n928 3.4105
R1508 VDDA.n964 VDDA.n928 3.4105
R1509 VDDA.n975 VDDA.n928 3.4105
R1510 VDDA.n963 VDDA.n928 3.4105
R1511 VDDA.n977 VDDA.n928 3.4105
R1512 VDDA.n962 VDDA.n928 3.4105
R1513 VDDA.n979 VDDA.n928 3.4105
R1514 VDDA.n961 VDDA.n928 3.4105
R1515 VDDA.n981 VDDA.n928 3.4105
R1516 VDDA.n960 VDDA.n928 3.4105
R1517 VDDA.n983 VDDA.n928 3.4105
R1518 VDDA.n959 VDDA.n928 3.4105
R1519 VDDA.n985 VDDA.n928 3.4105
R1520 VDDA.n958 VDDA.n928 3.4105
R1521 VDDA.n987 VDDA.n928 3.4105
R1522 VDDA.n957 VDDA.n928 3.4105
R1523 VDDA.n989 VDDA.n928 3.4105
R1524 VDDA.n956 VDDA.n928 3.4105
R1525 VDDA.n991 VDDA.n928 3.4105
R1526 VDDA.n955 VDDA.n928 3.4105
R1527 VDDA.n993 VDDA.n928 3.4105
R1528 VDDA.n954 VDDA.n928 3.4105
R1529 VDDA.n995 VDDA.n928 3.4105
R1530 VDDA.n953 VDDA.n928 3.4105
R1531 VDDA.n997 VDDA.n928 3.4105
R1532 VDDA.n952 VDDA.n928 3.4105
R1533 VDDA.n928 VDDA.n18 3.4105
R1534 VDDA.n999 VDDA.n928 3.4105
R1535 VDDA.n893 VDDA.n16 3.4105
R1536 VDDA.n969 VDDA.n893 3.4105
R1537 VDDA.n966 VDDA.n893 3.4105
R1538 VDDA.n971 VDDA.n893 3.4105
R1539 VDDA.n965 VDDA.n893 3.4105
R1540 VDDA.n973 VDDA.n893 3.4105
R1541 VDDA.n964 VDDA.n893 3.4105
R1542 VDDA.n975 VDDA.n893 3.4105
R1543 VDDA.n963 VDDA.n893 3.4105
R1544 VDDA.n977 VDDA.n893 3.4105
R1545 VDDA.n962 VDDA.n893 3.4105
R1546 VDDA.n979 VDDA.n893 3.4105
R1547 VDDA.n961 VDDA.n893 3.4105
R1548 VDDA.n981 VDDA.n893 3.4105
R1549 VDDA.n960 VDDA.n893 3.4105
R1550 VDDA.n983 VDDA.n893 3.4105
R1551 VDDA.n959 VDDA.n893 3.4105
R1552 VDDA.n985 VDDA.n893 3.4105
R1553 VDDA.n958 VDDA.n893 3.4105
R1554 VDDA.n987 VDDA.n893 3.4105
R1555 VDDA.n957 VDDA.n893 3.4105
R1556 VDDA.n989 VDDA.n893 3.4105
R1557 VDDA.n956 VDDA.n893 3.4105
R1558 VDDA.n991 VDDA.n893 3.4105
R1559 VDDA.n955 VDDA.n893 3.4105
R1560 VDDA.n993 VDDA.n893 3.4105
R1561 VDDA.n954 VDDA.n893 3.4105
R1562 VDDA.n995 VDDA.n893 3.4105
R1563 VDDA.n953 VDDA.n893 3.4105
R1564 VDDA.n997 VDDA.n893 3.4105
R1565 VDDA.n952 VDDA.n893 3.4105
R1566 VDDA.n893 VDDA.n18 3.4105
R1567 VDDA.n999 VDDA.n893 3.4105
R1568 VDDA.n931 VDDA.n16 3.4105
R1569 VDDA.n969 VDDA.n931 3.4105
R1570 VDDA.n966 VDDA.n931 3.4105
R1571 VDDA.n971 VDDA.n931 3.4105
R1572 VDDA.n965 VDDA.n931 3.4105
R1573 VDDA.n973 VDDA.n931 3.4105
R1574 VDDA.n964 VDDA.n931 3.4105
R1575 VDDA.n975 VDDA.n931 3.4105
R1576 VDDA.n963 VDDA.n931 3.4105
R1577 VDDA.n977 VDDA.n931 3.4105
R1578 VDDA.n962 VDDA.n931 3.4105
R1579 VDDA.n979 VDDA.n931 3.4105
R1580 VDDA.n961 VDDA.n931 3.4105
R1581 VDDA.n981 VDDA.n931 3.4105
R1582 VDDA.n960 VDDA.n931 3.4105
R1583 VDDA.n983 VDDA.n931 3.4105
R1584 VDDA.n959 VDDA.n931 3.4105
R1585 VDDA.n985 VDDA.n931 3.4105
R1586 VDDA.n958 VDDA.n931 3.4105
R1587 VDDA.n987 VDDA.n931 3.4105
R1588 VDDA.n957 VDDA.n931 3.4105
R1589 VDDA.n989 VDDA.n931 3.4105
R1590 VDDA.n956 VDDA.n931 3.4105
R1591 VDDA.n991 VDDA.n931 3.4105
R1592 VDDA.n955 VDDA.n931 3.4105
R1593 VDDA.n993 VDDA.n931 3.4105
R1594 VDDA.n954 VDDA.n931 3.4105
R1595 VDDA.n995 VDDA.n931 3.4105
R1596 VDDA.n953 VDDA.n931 3.4105
R1597 VDDA.n997 VDDA.n931 3.4105
R1598 VDDA.n952 VDDA.n931 3.4105
R1599 VDDA.n931 VDDA.n18 3.4105
R1600 VDDA.n999 VDDA.n931 3.4105
R1601 VDDA.n892 VDDA.n16 3.4105
R1602 VDDA.n969 VDDA.n892 3.4105
R1603 VDDA.n966 VDDA.n892 3.4105
R1604 VDDA.n971 VDDA.n892 3.4105
R1605 VDDA.n965 VDDA.n892 3.4105
R1606 VDDA.n973 VDDA.n892 3.4105
R1607 VDDA.n964 VDDA.n892 3.4105
R1608 VDDA.n975 VDDA.n892 3.4105
R1609 VDDA.n963 VDDA.n892 3.4105
R1610 VDDA.n977 VDDA.n892 3.4105
R1611 VDDA.n962 VDDA.n892 3.4105
R1612 VDDA.n979 VDDA.n892 3.4105
R1613 VDDA.n961 VDDA.n892 3.4105
R1614 VDDA.n981 VDDA.n892 3.4105
R1615 VDDA.n960 VDDA.n892 3.4105
R1616 VDDA.n983 VDDA.n892 3.4105
R1617 VDDA.n959 VDDA.n892 3.4105
R1618 VDDA.n985 VDDA.n892 3.4105
R1619 VDDA.n958 VDDA.n892 3.4105
R1620 VDDA.n987 VDDA.n892 3.4105
R1621 VDDA.n957 VDDA.n892 3.4105
R1622 VDDA.n989 VDDA.n892 3.4105
R1623 VDDA.n956 VDDA.n892 3.4105
R1624 VDDA.n991 VDDA.n892 3.4105
R1625 VDDA.n955 VDDA.n892 3.4105
R1626 VDDA.n993 VDDA.n892 3.4105
R1627 VDDA.n954 VDDA.n892 3.4105
R1628 VDDA.n995 VDDA.n892 3.4105
R1629 VDDA.n953 VDDA.n892 3.4105
R1630 VDDA.n997 VDDA.n892 3.4105
R1631 VDDA.n952 VDDA.n892 3.4105
R1632 VDDA.n892 VDDA.n18 3.4105
R1633 VDDA.n999 VDDA.n892 3.4105
R1634 VDDA.n934 VDDA.n16 3.4105
R1635 VDDA.n969 VDDA.n934 3.4105
R1636 VDDA.n966 VDDA.n934 3.4105
R1637 VDDA.n971 VDDA.n934 3.4105
R1638 VDDA.n965 VDDA.n934 3.4105
R1639 VDDA.n973 VDDA.n934 3.4105
R1640 VDDA.n964 VDDA.n934 3.4105
R1641 VDDA.n975 VDDA.n934 3.4105
R1642 VDDA.n963 VDDA.n934 3.4105
R1643 VDDA.n977 VDDA.n934 3.4105
R1644 VDDA.n962 VDDA.n934 3.4105
R1645 VDDA.n979 VDDA.n934 3.4105
R1646 VDDA.n961 VDDA.n934 3.4105
R1647 VDDA.n981 VDDA.n934 3.4105
R1648 VDDA.n960 VDDA.n934 3.4105
R1649 VDDA.n983 VDDA.n934 3.4105
R1650 VDDA.n959 VDDA.n934 3.4105
R1651 VDDA.n985 VDDA.n934 3.4105
R1652 VDDA.n958 VDDA.n934 3.4105
R1653 VDDA.n987 VDDA.n934 3.4105
R1654 VDDA.n957 VDDA.n934 3.4105
R1655 VDDA.n989 VDDA.n934 3.4105
R1656 VDDA.n956 VDDA.n934 3.4105
R1657 VDDA.n991 VDDA.n934 3.4105
R1658 VDDA.n955 VDDA.n934 3.4105
R1659 VDDA.n993 VDDA.n934 3.4105
R1660 VDDA.n954 VDDA.n934 3.4105
R1661 VDDA.n995 VDDA.n934 3.4105
R1662 VDDA.n953 VDDA.n934 3.4105
R1663 VDDA.n997 VDDA.n934 3.4105
R1664 VDDA.n952 VDDA.n934 3.4105
R1665 VDDA.n934 VDDA.n18 3.4105
R1666 VDDA.n999 VDDA.n934 3.4105
R1667 VDDA.n891 VDDA.n16 3.4105
R1668 VDDA.n969 VDDA.n891 3.4105
R1669 VDDA.n966 VDDA.n891 3.4105
R1670 VDDA.n971 VDDA.n891 3.4105
R1671 VDDA.n965 VDDA.n891 3.4105
R1672 VDDA.n973 VDDA.n891 3.4105
R1673 VDDA.n964 VDDA.n891 3.4105
R1674 VDDA.n975 VDDA.n891 3.4105
R1675 VDDA.n963 VDDA.n891 3.4105
R1676 VDDA.n977 VDDA.n891 3.4105
R1677 VDDA.n962 VDDA.n891 3.4105
R1678 VDDA.n979 VDDA.n891 3.4105
R1679 VDDA.n961 VDDA.n891 3.4105
R1680 VDDA.n981 VDDA.n891 3.4105
R1681 VDDA.n960 VDDA.n891 3.4105
R1682 VDDA.n983 VDDA.n891 3.4105
R1683 VDDA.n959 VDDA.n891 3.4105
R1684 VDDA.n985 VDDA.n891 3.4105
R1685 VDDA.n958 VDDA.n891 3.4105
R1686 VDDA.n987 VDDA.n891 3.4105
R1687 VDDA.n957 VDDA.n891 3.4105
R1688 VDDA.n989 VDDA.n891 3.4105
R1689 VDDA.n956 VDDA.n891 3.4105
R1690 VDDA.n991 VDDA.n891 3.4105
R1691 VDDA.n955 VDDA.n891 3.4105
R1692 VDDA.n993 VDDA.n891 3.4105
R1693 VDDA.n954 VDDA.n891 3.4105
R1694 VDDA.n995 VDDA.n891 3.4105
R1695 VDDA.n953 VDDA.n891 3.4105
R1696 VDDA.n997 VDDA.n891 3.4105
R1697 VDDA.n952 VDDA.n891 3.4105
R1698 VDDA.n891 VDDA.n18 3.4105
R1699 VDDA.n999 VDDA.n891 3.4105
R1700 VDDA.n937 VDDA.n16 3.4105
R1701 VDDA.n969 VDDA.n937 3.4105
R1702 VDDA.n966 VDDA.n937 3.4105
R1703 VDDA.n971 VDDA.n937 3.4105
R1704 VDDA.n965 VDDA.n937 3.4105
R1705 VDDA.n973 VDDA.n937 3.4105
R1706 VDDA.n964 VDDA.n937 3.4105
R1707 VDDA.n975 VDDA.n937 3.4105
R1708 VDDA.n963 VDDA.n937 3.4105
R1709 VDDA.n977 VDDA.n937 3.4105
R1710 VDDA.n962 VDDA.n937 3.4105
R1711 VDDA.n979 VDDA.n937 3.4105
R1712 VDDA.n961 VDDA.n937 3.4105
R1713 VDDA.n981 VDDA.n937 3.4105
R1714 VDDA.n960 VDDA.n937 3.4105
R1715 VDDA.n983 VDDA.n937 3.4105
R1716 VDDA.n959 VDDA.n937 3.4105
R1717 VDDA.n985 VDDA.n937 3.4105
R1718 VDDA.n958 VDDA.n937 3.4105
R1719 VDDA.n987 VDDA.n937 3.4105
R1720 VDDA.n957 VDDA.n937 3.4105
R1721 VDDA.n989 VDDA.n937 3.4105
R1722 VDDA.n956 VDDA.n937 3.4105
R1723 VDDA.n991 VDDA.n937 3.4105
R1724 VDDA.n955 VDDA.n937 3.4105
R1725 VDDA.n993 VDDA.n937 3.4105
R1726 VDDA.n954 VDDA.n937 3.4105
R1727 VDDA.n995 VDDA.n937 3.4105
R1728 VDDA.n953 VDDA.n937 3.4105
R1729 VDDA.n997 VDDA.n937 3.4105
R1730 VDDA.n952 VDDA.n937 3.4105
R1731 VDDA.n937 VDDA.n18 3.4105
R1732 VDDA.n999 VDDA.n937 3.4105
R1733 VDDA.n890 VDDA.n16 3.4105
R1734 VDDA.n969 VDDA.n890 3.4105
R1735 VDDA.n966 VDDA.n890 3.4105
R1736 VDDA.n971 VDDA.n890 3.4105
R1737 VDDA.n965 VDDA.n890 3.4105
R1738 VDDA.n973 VDDA.n890 3.4105
R1739 VDDA.n964 VDDA.n890 3.4105
R1740 VDDA.n975 VDDA.n890 3.4105
R1741 VDDA.n963 VDDA.n890 3.4105
R1742 VDDA.n977 VDDA.n890 3.4105
R1743 VDDA.n962 VDDA.n890 3.4105
R1744 VDDA.n979 VDDA.n890 3.4105
R1745 VDDA.n961 VDDA.n890 3.4105
R1746 VDDA.n981 VDDA.n890 3.4105
R1747 VDDA.n960 VDDA.n890 3.4105
R1748 VDDA.n983 VDDA.n890 3.4105
R1749 VDDA.n959 VDDA.n890 3.4105
R1750 VDDA.n985 VDDA.n890 3.4105
R1751 VDDA.n958 VDDA.n890 3.4105
R1752 VDDA.n987 VDDA.n890 3.4105
R1753 VDDA.n957 VDDA.n890 3.4105
R1754 VDDA.n989 VDDA.n890 3.4105
R1755 VDDA.n956 VDDA.n890 3.4105
R1756 VDDA.n991 VDDA.n890 3.4105
R1757 VDDA.n955 VDDA.n890 3.4105
R1758 VDDA.n993 VDDA.n890 3.4105
R1759 VDDA.n954 VDDA.n890 3.4105
R1760 VDDA.n995 VDDA.n890 3.4105
R1761 VDDA.n953 VDDA.n890 3.4105
R1762 VDDA.n997 VDDA.n890 3.4105
R1763 VDDA.n952 VDDA.n890 3.4105
R1764 VDDA.n890 VDDA.n18 3.4105
R1765 VDDA.n999 VDDA.n890 3.4105
R1766 VDDA.n940 VDDA.n16 3.4105
R1767 VDDA.n969 VDDA.n940 3.4105
R1768 VDDA.n966 VDDA.n940 3.4105
R1769 VDDA.n971 VDDA.n940 3.4105
R1770 VDDA.n965 VDDA.n940 3.4105
R1771 VDDA.n973 VDDA.n940 3.4105
R1772 VDDA.n964 VDDA.n940 3.4105
R1773 VDDA.n975 VDDA.n940 3.4105
R1774 VDDA.n963 VDDA.n940 3.4105
R1775 VDDA.n977 VDDA.n940 3.4105
R1776 VDDA.n962 VDDA.n940 3.4105
R1777 VDDA.n979 VDDA.n940 3.4105
R1778 VDDA.n961 VDDA.n940 3.4105
R1779 VDDA.n981 VDDA.n940 3.4105
R1780 VDDA.n960 VDDA.n940 3.4105
R1781 VDDA.n983 VDDA.n940 3.4105
R1782 VDDA.n959 VDDA.n940 3.4105
R1783 VDDA.n985 VDDA.n940 3.4105
R1784 VDDA.n958 VDDA.n940 3.4105
R1785 VDDA.n987 VDDA.n940 3.4105
R1786 VDDA.n957 VDDA.n940 3.4105
R1787 VDDA.n989 VDDA.n940 3.4105
R1788 VDDA.n956 VDDA.n940 3.4105
R1789 VDDA.n991 VDDA.n940 3.4105
R1790 VDDA.n955 VDDA.n940 3.4105
R1791 VDDA.n993 VDDA.n940 3.4105
R1792 VDDA.n954 VDDA.n940 3.4105
R1793 VDDA.n995 VDDA.n940 3.4105
R1794 VDDA.n953 VDDA.n940 3.4105
R1795 VDDA.n997 VDDA.n940 3.4105
R1796 VDDA.n952 VDDA.n940 3.4105
R1797 VDDA.n940 VDDA.n18 3.4105
R1798 VDDA.n999 VDDA.n940 3.4105
R1799 VDDA.n889 VDDA.n16 3.4105
R1800 VDDA.n969 VDDA.n889 3.4105
R1801 VDDA.n966 VDDA.n889 3.4105
R1802 VDDA.n971 VDDA.n889 3.4105
R1803 VDDA.n965 VDDA.n889 3.4105
R1804 VDDA.n973 VDDA.n889 3.4105
R1805 VDDA.n964 VDDA.n889 3.4105
R1806 VDDA.n975 VDDA.n889 3.4105
R1807 VDDA.n963 VDDA.n889 3.4105
R1808 VDDA.n977 VDDA.n889 3.4105
R1809 VDDA.n962 VDDA.n889 3.4105
R1810 VDDA.n979 VDDA.n889 3.4105
R1811 VDDA.n961 VDDA.n889 3.4105
R1812 VDDA.n981 VDDA.n889 3.4105
R1813 VDDA.n960 VDDA.n889 3.4105
R1814 VDDA.n983 VDDA.n889 3.4105
R1815 VDDA.n959 VDDA.n889 3.4105
R1816 VDDA.n985 VDDA.n889 3.4105
R1817 VDDA.n958 VDDA.n889 3.4105
R1818 VDDA.n987 VDDA.n889 3.4105
R1819 VDDA.n957 VDDA.n889 3.4105
R1820 VDDA.n989 VDDA.n889 3.4105
R1821 VDDA.n956 VDDA.n889 3.4105
R1822 VDDA.n991 VDDA.n889 3.4105
R1823 VDDA.n955 VDDA.n889 3.4105
R1824 VDDA.n993 VDDA.n889 3.4105
R1825 VDDA.n954 VDDA.n889 3.4105
R1826 VDDA.n995 VDDA.n889 3.4105
R1827 VDDA.n953 VDDA.n889 3.4105
R1828 VDDA.n997 VDDA.n889 3.4105
R1829 VDDA.n952 VDDA.n889 3.4105
R1830 VDDA.n889 VDDA.n18 3.4105
R1831 VDDA.n999 VDDA.n889 3.4105
R1832 VDDA.n943 VDDA.n16 3.4105
R1833 VDDA.n969 VDDA.n943 3.4105
R1834 VDDA.n966 VDDA.n943 3.4105
R1835 VDDA.n971 VDDA.n943 3.4105
R1836 VDDA.n965 VDDA.n943 3.4105
R1837 VDDA.n973 VDDA.n943 3.4105
R1838 VDDA.n964 VDDA.n943 3.4105
R1839 VDDA.n975 VDDA.n943 3.4105
R1840 VDDA.n963 VDDA.n943 3.4105
R1841 VDDA.n977 VDDA.n943 3.4105
R1842 VDDA.n962 VDDA.n943 3.4105
R1843 VDDA.n979 VDDA.n943 3.4105
R1844 VDDA.n961 VDDA.n943 3.4105
R1845 VDDA.n981 VDDA.n943 3.4105
R1846 VDDA.n960 VDDA.n943 3.4105
R1847 VDDA.n983 VDDA.n943 3.4105
R1848 VDDA.n959 VDDA.n943 3.4105
R1849 VDDA.n985 VDDA.n943 3.4105
R1850 VDDA.n958 VDDA.n943 3.4105
R1851 VDDA.n987 VDDA.n943 3.4105
R1852 VDDA.n957 VDDA.n943 3.4105
R1853 VDDA.n989 VDDA.n943 3.4105
R1854 VDDA.n956 VDDA.n943 3.4105
R1855 VDDA.n991 VDDA.n943 3.4105
R1856 VDDA.n955 VDDA.n943 3.4105
R1857 VDDA.n993 VDDA.n943 3.4105
R1858 VDDA.n954 VDDA.n943 3.4105
R1859 VDDA.n995 VDDA.n943 3.4105
R1860 VDDA.n953 VDDA.n943 3.4105
R1861 VDDA.n997 VDDA.n943 3.4105
R1862 VDDA.n952 VDDA.n943 3.4105
R1863 VDDA.n943 VDDA.n18 3.4105
R1864 VDDA.n999 VDDA.n943 3.4105
R1865 VDDA.n888 VDDA.n16 3.4105
R1866 VDDA.n969 VDDA.n888 3.4105
R1867 VDDA.n966 VDDA.n888 3.4105
R1868 VDDA.n971 VDDA.n888 3.4105
R1869 VDDA.n965 VDDA.n888 3.4105
R1870 VDDA.n973 VDDA.n888 3.4105
R1871 VDDA.n964 VDDA.n888 3.4105
R1872 VDDA.n975 VDDA.n888 3.4105
R1873 VDDA.n963 VDDA.n888 3.4105
R1874 VDDA.n977 VDDA.n888 3.4105
R1875 VDDA.n962 VDDA.n888 3.4105
R1876 VDDA.n979 VDDA.n888 3.4105
R1877 VDDA.n961 VDDA.n888 3.4105
R1878 VDDA.n981 VDDA.n888 3.4105
R1879 VDDA.n960 VDDA.n888 3.4105
R1880 VDDA.n983 VDDA.n888 3.4105
R1881 VDDA.n959 VDDA.n888 3.4105
R1882 VDDA.n985 VDDA.n888 3.4105
R1883 VDDA.n958 VDDA.n888 3.4105
R1884 VDDA.n987 VDDA.n888 3.4105
R1885 VDDA.n957 VDDA.n888 3.4105
R1886 VDDA.n989 VDDA.n888 3.4105
R1887 VDDA.n956 VDDA.n888 3.4105
R1888 VDDA.n991 VDDA.n888 3.4105
R1889 VDDA.n955 VDDA.n888 3.4105
R1890 VDDA.n993 VDDA.n888 3.4105
R1891 VDDA.n954 VDDA.n888 3.4105
R1892 VDDA.n995 VDDA.n888 3.4105
R1893 VDDA.n953 VDDA.n888 3.4105
R1894 VDDA.n997 VDDA.n888 3.4105
R1895 VDDA.n952 VDDA.n888 3.4105
R1896 VDDA.n888 VDDA.n18 3.4105
R1897 VDDA.n999 VDDA.n888 3.4105
R1898 VDDA.n946 VDDA.n16 3.4105
R1899 VDDA.n969 VDDA.n946 3.4105
R1900 VDDA.n966 VDDA.n946 3.4105
R1901 VDDA.n971 VDDA.n946 3.4105
R1902 VDDA.n965 VDDA.n946 3.4105
R1903 VDDA.n973 VDDA.n946 3.4105
R1904 VDDA.n964 VDDA.n946 3.4105
R1905 VDDA.n975 VDDA.n946 3.4105
R1906 VDDA.n963 VDDA.n946 3.4105
R1907 VDDA.n977 VDDA.n946 3.4105
R1908 VDDA.n962 VDDA.n946 3.4105
R1909 VDDA.n979 VDDA.n946 3.4105
R1910 VDDA.n961 VDDA.n946 3.4105
R1911 VDDA.n981 VDDA.n946 3.4105
R1912 VDDA.n960 VDDA.n946 3.4105
R1913 VDDA.n983 VDDA.n946 3.4105
R1914 VDDA.n959 VDDA.n946 3.4105
R1915 VDDA.n985 VDDA.n946 3.4105
R1916 VDDA.n958 VDDA.n946 3.4105
R1917 VDDA.n987 VDDA.n946 3.4105
R1918 VDDA.n957 VDDA.n946 3.4105
R1919 VDDA.n989 VDDA.n946 3.4105
R1920 VDDA.n956 VDDA.n946 3.4105
R1921 VDDA.n991 VDDA.n946 3.4105
R1922 VDDA.n955 VDDA.n946 3.4105
R1923 VDDA.n993 VDDA.n946 3.4105
R1924 VDDA.n954 VDDA.n946 3.4105
R1925 VDDA.n995 VDDA.n946 3.4105
R1926 VDDA.n953 VDDA.n946 3.4105
R1927 VDDA.n997 VDDA.n946 3.4105
R1928 VDDA.n952 VDDA.n946 3.4105
R1929 VDDA.n946 VDDA.n18 3.4105
R1930 VDDA.n999 VDDA.n946 3.4105
R1931 VDDA.n887 VDDA.n16 3.4105
R1932 VDDA.n969 VDDA.n887 3.4105
R1933 VDDA.n966 VDDA.n887 3.4105
R1934 VDDA.n971 VDDA.n887 3.4105
R1935 VDDA.n965 VDDA.n887 3.4105
R1936 VDDA.n973 VDDA.n887 3.4105
R1937 VDDA.n964 VDDA.n887 3.4105
R1938 VDDA.n975 VDDA.n887 3.4105
R1939 VDDA.n963 VDDA.n887 3.4105
R1940 VDDA.n977 VDDA.n887 3.4105
R1941 VDDA.n962 VDDA.n887 3.4105
R1942 VDDA.n979 VDDA.n887 3.4105
R1943 VDDA.n961 VDDA.n887 3.4105
R1944 VDDA.n981 VDDA.n887 3.4105
R1945 VDDA.n960 VDDA.n887 3.4105
R1946 VDDA.n983 VDDA.n887 3.4105
R1947 VDDA.n959 VDDA.n887 3.4105
R1948 VDDA.n985 VDDA.n887 3.4105
R1949 VDDA.n958 VDDA.n887 3.4105
R1950 VDDA.n987 VDDA.n887 3.4105
R1951 VDDA.n957 VDDA.n887 3.4105
R1952 VDDA.n989 VDDA.n887 3.4105
R1953 VDDA.n956 VDDA.n887 3.4105
R1954 VDDA.n991 VDDA.n887 3.4105
R1955 VDDA.n955 VDDA.n887 3.4105
R1956 VDDA.n993 VDDA.n887 3.4105
R1957 VDDA.n954 VDDA.n887 3.4105
R1958 VDDA.n995 VDDA.n887 3.4105
R1959 VDDA.n953 VDDA.n887 3.4105
R1960 VDDA.n997 VDDA.n887 3.4105
R1961 VDDA.n952 VDDA.n887 3.4105
R1962 VDDA.n887 VDDA.n18 3.4105
R1963 VDDA.n999 VDDA.n887 3.4105
R1964 VDDA.n949 VDDA.n16 3.4105
R1965 VDDA.n969 VDDA.n949 3.4105
R1966 VDDA.n966 VDDA.n949 3.4105
R1967 VDDA.n971 VDDA.n949 3.4105
R1968 VDDA.n965 VDDA.n949 3.4105
R1969 VDDA.n973 VDDA.n949 3.4105
R1970 VDDA.n964 VDDA.n949 3.4105
R1971 VDDA.n975 VDDA.n949 3.4105
R1972 VDDA.n963 VDDA.n949 3.4105
R1973 VDDA.n977 VDDA.n949 3.4105
R1974 VDDA.n962 VDDA.n949 3.4105
R1975 VDDA.n979 VDDA.n949 3.4105
R1976 VDDA.n961 VDDA.n949 3.4105
R1977 VDDA.n981 VDDA.n949 3.4105
R1978 VDDA.n960 VDDA.n949 3.4105
R1979 VDDA.n983 VDDA.n949 3.4105
R1980 VDDA.n959 VDDA.n949 3.4105
R1981 VDDA.n985 VDDA.n949 3.4105
R1982 VDDA.n958 VDDA.n949 3.4105
R1983 VDDA.n987 VDDA.n949 3.4105
R1984 VDDA.n957 VDDA.n949 3.4105
R1985 VDDA.n989 VDDA.n949 3.4105
R1986 VDDA.n956 VDDA.n949 3.4105
R1987 VDDA.n991 VDDA.n949 3.4105
R1988 VDDA.n955 VDDA.n949 3.4105
R1989 VDDA.n993 VDDA.n949 3.4105
R1990 VDDA.n954 VDDA.n949 3.4105
R1991 VDDA.n995 VDDA.n949 3.4105
R1992 VDDA.n953 VDDA.n949 3.4105
R1993 VDDA.n997 VDDA.n949 3.4105
R1994 VDDA.n952 VDDA.n949 3.4105
R1995 VDDA.n949 VDDA.n18 3.4105
R1996 VDDA.n999 VDDA.n949 3.4105
R1997 VDDA.n886 VDDA.n16 3.4105
R1998 VDDA.n969 VDDA.n886 3.4105
R1999 VDDA.n966 VDDA.n886 3.4105
R2000 VDDA.n971 VDDA.n886 3.4105
R2001 VDDA.n965 VDDA.n886 3.4105
R2002 VDDA.n973 VDDA.n886 3.4105
R2003 VDDA.n964 VDDA.n886 3.4105
R2004 VDDA.n975 VDDA.n886 3.4105
R2005 VDDA.n963 VDDA.n886 3.4105
R2006 VDDA.n977 VDDA.n886 3.4105
R2007 VDDA.n962 VDDA.n886 3.4105
R2008 VDDA.n979 VDDA.n886 3.4105
R2009 VDDA.n961 VDDA.n886 3.4105
R2010 VDDA.n981 VDDA.n886 3.4105
R2011 VDDA.n960 VDDA.n886 3.4105
R2012 VDDA.n983 VDDA.n886 3.4105
R2013 VDDA.n959 VDDA.n886 3.4105
R2014 VDDA.n985 VDDA.n886 3.4105
R2015 VDDA.n958 VDDA.n886 3.4105
R2016 VDDA.n987 VDDA.n886 3.4105
R2017 VDDA.n957 VDDA.n886 3.4105
R2018 VDDA.n989 VDDA.n886 3.4105
R2019 VDDA.n956 VDDA.n886 3.4105
R2020 VDDA.n991 VDDA.n886 3.4105
R2021 VDDA.n955 VDDA.n886 3.4105
R2022 VDDA.n993 VDDA.n886 3.4105
R2023 VDDA.n954 VDDA.n886 3.4105
R2024 VDDA.n995 VDDA.n886 3.4105
R2025 VDDA.n953 VDDA.n886 3.4105
R2026 VDDA.n997 VDDA.n886 3.4105
R2027 VDDA.n952 VDDA.n886 3.4105
R2028 VDDA.n886 VDDA.n18 3.4105
R2029 VDDA.n999 VDDA.n886 3.4105
R2030 VDDA.n998 VDDA.n969 3.4105
R2031 VDDA.n998 VDDA.n966 3.4105
R2032 VDDA.n998 VDDA.n971 3.4105
R2033 VDDA.n998 VDDA.n965 3.4105
R2034 VDDA.n998 VDDA.n973 3.4105
R2035 VDDA.n998 VDDA.n964 3.4105
R2036 VDDA.n998 VDDA.n975 3.4105
R2037 VDDA.n998 VDDA.n963 3.4105
R2038 VDDA.n998 VDDA.n977 3.4105
R2039 VDDA.n998 VDDA.n962 3.4105
R2040 VDDA.n998 VDDA.n979 3.4105
R2041 VDDA.n998 VDDA.n961 3.4105
R2042 VDDA.n998 VDDA.n981 3.4105
R2043 VDDA.n998 VDDA.n960 3.4105
R2044 VDDA.n998 VDDA.n983 3.4105
R2045 VDDA.n998 VDDA.n959 3.4105
R2046 VDDA.n998 VDDA.n985 3.4105
R2047 VDDA.n998 VDDA.n958 3.4105
R2048 VDDA.n998 VDDA.n987 3.4105
R2049 VDDA.n998 VDDA.n957 3.4105
R2050 VDDA.n998 VDDA.n989 3.4105
R2051 VDDA.n998 VDDA.n956 3.4105
R2052 VDDA.n998 VDDA.n991 3.4105
R2053 VDDA.n998 VDDA.n955 3.4105
R2054 VDDA.n998 VDDA.n993 3.4105
R2055 VDDA.n998 VDDA.n954 3.4105
R2056 VDDA.n998 VDDA.n995 3.4105
R2057 VDDA.n998 VDDA.n953 3.4105
R2058 VDDA.n998 VDDA.n997 3.4105
R2059 VDDA.n998 VDDA.n952 3.4105
R2060 VDDA.n998 VDDA.n18 3.4105
R2061 VDDA.n999 VDDA.n998 3.4105
R2062 VDDA.n445 VDDA.n444 3.11118
R2063 VDDA.n455 VDDA.n454 3.11118
R2064 VDDA.n444 VDDA.n426 3.04304
R2065 VDDA.n454 VDDA.n406 3.04304
R2066 VDDA.n882 VDDA.n881 2.97446
R2067 VDDA.n725 VDDA.n721 2.97446
R2068 VDDA.n238 VDDA.n234 2.96402
R2069 VDDA.n853 VDDA.n849 2.96402
R2070 VDDA.n779 VDDA.n778 2.8255
R2071 VDDA.n781 VDDA.n780 2.8255
R2072 VDDA.n237 VDDA.n236 2.423
R2073 VDDA.n235 VDDA.n234 2.423
R2074 VDDA.n850 VDDA.n849 2.423
R2075 VDDA.n852 VDDA.n851 2.423
R2076 VDDA.n819 VDDA.n817 2.3971
R2077 VDDA.n359 VDDA.n358 2.39683
R2078 VDDA.n750 VDDA.n206 2.39632
R2079 VDDA.n308 VDDA.n306 2.3573
R2080 VDDA.n136 VDDA.n135 2.30736
R2081 VDDA.n659 VDDA.n657 2.30736
R2082 VDDA.n99 VDDA.n98 2.30612
R2083 VDDA.n644 VDDA.n643 2.30612
R2084 VDDA.n238 VDDA.n237 2.27652
R2085 VDDA.n853 VDDA.n852 2.27652
R2086 VDDA.n400 VDDA.n392 2.26187
R2087 VDDA.n466 VDDA.n390 2.26187
R2088 VDDA.n543 VDDA.n388 2.26187
R2089 VDDA.n593 VDDA.n386 2.26187
R2090 VDDA.n770 VDDA.n761 2.26187
R2091 VDDA.n772 VDDA.n770 2.26187
R2092 VDDA.n859 VDDA.n858 2.26187
R2093 VDDA.n846 VDDA.n824 2.26187
R2094 VDDA.n830 VDDA.n827 2.26187
R2095 VDDA.n831 VDDA.n830 2.26187
R2096 VDDA.n749 VDDA.n748 2.26187
R2097 VDDA.n231 VDDA.n230 2.26187
R2098 VDDA.n724 VDDA.n723 2.26187
R2099 VDDA.n723 VDDA.n247 2.26187
R2100 VDDA.n397 VDDA.n392 2.26187
R2101 VDDA.n232 VDDA.n231 2.26187
R2102 VDDA.n243 VDDA.n242 2.26187
R2103 VDDA.n788 VDDA.n787 2.26187
R2104 VDDA.n401 VDDA.n391 2.24063
R2105 VDDA.n467 VDDA.n389 2.24063
R2106 VDDA.n544 VDDA.n387 2.24063
R2107 VDDA.n594 VDDA.n385 2.24063
R2108 VDDA.n789 VDDA.n788 2.24063
R2109 VDDA.n783 VDDA.n759 2.24063
R2110 VDDA.n785 VDDA.n784 2.24063
R2111 VDDA.n775 VDDA.n774 2.24063
R2112 VDDA.n880 VDDA.n879 2.24063
R2113 VDDA.n179 VDDA.n178 2.24063
R2114 VDDA.n857 VDDA.n182 2.24063
R2115 VDDA.n848 VDDA.n847 2.24063
R2116 VDDA.n818 VDDA.n185 2.24063
R2117 VDDA.n802 VDDA.n184 2.24063
R2118 VDDA.n792 VDDA.n791 2.24063
R2119 VDDA.n758 VDDA.n189 2.24063
R2120 VDDA.n747 VDDA.n190 2.24063
R2121 VDDA.n240 VDDA.n239 2.24063
R2122 VDDA.n242 VDDA.n241 2.24063
R2123 VDDA.n230 VDDA.n229 2.24063
R2124 VDDA.n745 VDDA.n744 2.24063
R2125 VDDA.n211 VDDA.n210 2.24063
R2126 VDDA.n397 VDDA.n396 2.24063
R2127 VDDA.n402 VDDA.n390 2.24063
R2128 VDDA.n463 VDDA.n462 2.24063
R2129 VDDA.n468 VDDA.n388 2.24063
R2130 VDDA.n540 VDDA.n539 2.24063
R2131 VDDA.n545 VDDA.n386 2.24063
R2132 VDDA.n590 VDDA.n589 2.24063
R2133 VDDA.n773 VDDA.n772 2.24063
R2134 VDDA.n881 VDDA.n176 2.24063
R2135 VDDA.n860 VDDA.n859 2.24063
R2136 VDDA.n862 VDDA.n861 2.24063
R2137 VDDA.n856 VDDA.n824 2.24063
R2138 VDDA.n855 VDDA.n854 2.24063
R2139 VDDA.n845 VDDA.n827 2.24063
R2140 VDDA.n844 VDDA.n843 2.24063
R2141 VDDA.n820 VDDA.n819 2.24063
R2142 VDDA.n750 VDDA.n749 2.24063
R2143 VDDA.n752 VDDA.n751 2.24063
R2144 VDDA.n244 VDDA.n212 2.24063
R2145 VDDA.n233 VDDA.n215 2.24063
R2146 VDDA.n746 VDDA.n208 2.24063
R2147 VDDA.n725 VDDA.n724 2.24063
R2148 VDDA.n727 VDDA.n726 2.24063
R2149 VDDA.n875 VDDA.n874 1.97758
R2150 VDDA.n873 VDDA.n872 1.97758
R2151 VDDA.n740 VDDA.n739 1.97758
R2152 VDDA.n738 VDDA.n737 1.97758
R2153 VDDA.n443 VDDA.n442 1.90331
R2154 VDDA.n768 VDDA.n767 1.888
R2155 VDDA.n766 VDDA.n765 1.888
R2156 VDDA.n814 VDDA.n813 1.888
R2157 VDDA.n816 VDDA.n815 1.888
R2158 VDDA.n205 VDDA.n204 1.888
R2159 VDDA.n203 VDDA.n202 1.888
R2160 VDDA.n876 VDDA.n875 1.88069
R2161 VDDA.n872 VDDA.n871 1.88069
R2162 VDDA.n741 VDDA.n740 1.88069
R2163 VDDA.n737 VDDA.n736 1.88069
R2164 VDDA.n451 VDDA.n450 1.77831
R2165 VDDA.n453 VDDA.n452 1.77831
R2166 VDDA.n461 VDDA.n460 1.77831
R2167 VDDA.n384 VDDA.n372 1.73971
R2168 VDDA.n646 VDDA.n372 1.70624
R2169 VDDA.n902 VDDA.n0 1.70567
R2170 VDDA.n903 VDDA.n17 1.70567
R2171 VDDA.n905 VDDA.n902 1.70567
R2172 VDDA.n906 VDDA.n17 1.70567
R2173 VDDA.n908 VDDA.n902 1.70567
R2174 VDDA.n909 VDDA.n17 1.70567
R2175 VDDA.n911 VDDA.n902 1.70567
R2176 VDDA.n912 VDDA.n17 1.70567
R2177 VDDA.n914 VDDA.n902 1.70567
R2178 VDDA.n915 VDDA.n17 1.70567
R2179 VDDA.n917 VDDA.n902 1.70567
R2180 VDDA.n918 VDDA.n17 1.70567
R2181 VDDA.n920 VDDA.n902 1.70567
R2182 VDDA.n921 VDDA.n17 1.70567
R2183 VDDA.n923 VDDA.n902 1.70567
R2184 VDDA.n924 VDDA.n17 1.70567
R2185 VDDA.n926 VDDA.n902 1.70567
R2186 VDDA.n927 VDDA.n17 1.70567
R2187 VDDA.n929 VDDA.n902 1.70567
R2188 VDDA.n930 VDDA.n17 1.70567
R2189 VDDA.n932 VDDA.n902 1.70567
R2190 VDDA.n933 VDDA.n17 1.70567
R2191 VDDA.n935 VDDA.n902 1.70567
R2192 VDDA.n936 VDDA.n17 1.70567
R2193 VDDA.n938 VDDA.n902 1.70567
R2194 VDDA.n939 VDDA.n17 1.70567
R2195 VDDA.n941 VDDA.n902 1.70567
R2196 VDDA.n942 VDDA.n17 1.70567
R2197 VDDA.n944 VDDA.n902 1.70567
R2198 VDDA.n945 VDDA.n17 1.70567
R2199 VDDA.n947 VDDA.n902 1.70567
R2200 VDDA.n948 VDDA.n17 1.70567
R2201 VDDA.n950 VDDA.n902 1.70567
R2202 VDDA.n1000 VDDA.n15 1.70566
R2203 VDDA.n1000 VDDA.n14 1.70566
R2204 VDDA.n1000 VDDA.n13 1.70566
R2205 VDDA.n1000 VDDA.n12 1.70566
R2206 VDDA.n1000 VDDA.n11 1.70566
R2207 VDDA.n1000 VDDA.n10 1.70566
R2208 VDDA.n1000 VDDA.n9 1.70566
R2209 VDDA.n1000 VDDA.n8 1.70566
R2210 VDDA.n1000 VDDA.n7 1.70566
R2211 VDDA.n1000 VDDA.n6 1.70566
R2212 VDDA.n1000 VDDA.n5 1.70566
R2213 VDDA.n1000 VDDA.n4 1.70566
R2214 VDDA.n1000 VDDA.n3 1.70566
R2215 VDDA.n1000 VDDA.n2 1.70566
R2216 VDDA.n1000 VDDA.n1 1.70566
R2217 VDDA.n968 VDDA.n904 1.70566
R2218 VDDA.n970 VDDA.n904 1.70566
R2219 VDDA.n972 VDDA.n904 1.70566
R2220 VDDA.n974 VDDA.n904 1.70566
R2221 VDDA.n976 VDDA.n904 1.70566
R2222 VDDA.n978 VDDA.n904 1.70566
R2223 VDDA.n980 VDDA.n904 1.70566
R2224 VDDA.n982 VDDA.n904 1.70566
R2225 VDDA.n984 VDDA.n904 1.70566
R2226 VDDA.n986 VDDA.n904 1.70566
R2227 VDDA.n988 VDDA.n904 1.70566
R2228 VDDA.n990 VDDA.n904 1.70566
R2229 VDDA.n992 VDDA.n904 1.70566
R2230 VDDA.n994 VDDA.n904 1.70566
R2231 VDDA.n996 VDDA.n904 1.70566
R2232 VDDA.n951 VDDA.n904 1.70566
R2233 VDDA.n998 VDDA.n967 1.70566
R2234 VDDA.n718 VDDA.n648 1.69337
R2235 VDDA.n718 VDDA.n649 1.69337
R2236 VDDA.n718 VDDA.n651 1.69337
R2237 VDDA.n718 VDDA.n652 1.69337
R2238 VDDA.n718 VDDA.n654 1.69337
R2239 VDDA.n718 VDDA.n655 1.69337
R2240 VDDA.n718 VDDA.n717 1.69337
R2241 VDDA.n646 VDDA.n363 1.69337
R2242 VDDA.n646 VDDA.n364 1.69337
R2243 VDDA.n646 VDDA.n366 1.69337
R2244 VDDA.n646 VDDA.n367 1.69337
R2245 VDDA.n646 VDDA.n369 1.69337
R2246 VDDA.n646 VDDA.n370 1.69337
R2247 VDDA.n885 VDDA.n103 1.69337
R2248 VDDA.n885 VDDA.n104 1.69337
R2249 VDDA.n885 VDDA.n106 1.69337
R2250 VDDA.n885 VDDA.n107 1.69337
R2251 VDDA.n885 VDDA.n109 1.69337
R2252 VDDA.n885 VDDA.n110 1.69337
R2253 VDDA.n885 VDDA.n112 1.69337
R2254 VDDA.n101 VDDA.n20 1.69337
R2255 VDDA.n101 VDDA.n21 1.69337
R2256 VDDA.n101 VDDA.n23 1.69337
R2257 VDDA.n101 VDDA.n24 1.69337
R2258 VDDA.n101 VDDA.n26 1.69337
R2259 VDDA.n101 VDDA.n27 1.69337
R2260 VDDA.n101 VDDA.n29 1.69337
R2261 VDDA.n361 VDDA.n253 1.69337
R2262 VDDA.n361 VDDA.n254 1.69337
R2263 VDDA.n361 VDDA.n256 1.69337
R2264 VDDA.n361 VDDA.n257 1.69337
R2265 VDDA.n361 VDDA.n259 1.69337
R2266 VDDA.n361 VDDA.n260 1.69337
R2267 VDDA.n361 VDDA.n262 1.69337
R2268 VDDA.n718 VDDA.n647 1.6924
R2269 VDDA.n718 VDDA.n650 1.6924
R2270 VDDA.n718 VDDA.n653 1.6924
R2271 VDDA.n718 VDDA.n656 1.6924
R2272 VDDA.n646 VDDA.n362 1.6924
R2273 VDDA.n646 VDDA.n365 1.6924
R2274 VDDA.n646 VDDA.n368 1.6924
R2275 VDDA.n646 VDDA.n371 1.6924
R2276 VDDA.n885 VDDA.n102 1.6924
R2277 VDDA.n885 VDDA.n105 1.6924
R2278 VDDA.n885 VDDA.n108 1.6924
R2279 VDDA.n885 VDDA.n111 1.6924
R2280 VDDA.n101 VDDA.n19 1.6924
R2281 VDDA.n101 VDDA.n22 1.6924
R2282 VDDA.n101 VDDA.n25 1.6924
R2283 VDDA.n101 VDDA.n28 1.6924
R2284 VDDA.n361 VDDA.n252 1.6924
R2285 VDDA.n361 VDDA.n255 1.6924
R2286 VDDA.n361 VDDA.n258 1.6924
R2287 VDDA.n361 VDDA.n261 1.6924
R2288 VDDA.n569 VDDA.n567 1.68456
R2289 VDDA.n285 VDDA.n276 1.68356
R2290 VDDA.n765 VDDA.n763 1.63212
R2291 VDDA.n778 VDDA.n777 1.63212
R2292 VDDA.n585 VDDA.n551 1.56997
R2293 VDDA.n580 VDDA.n554 1.56997
R2294 VDDA.n572 VDDA.n564 1.56997
R2295 VDDA.n769 VDDA.n768 1.56962
R2296 VDDA.n782 VDDA.n781 1.56962
R2297 VDDA.n306 VDDA.n276 1.50969
R2298 VDDA.n396 VDDA.n395 1.26222
R2299 VDDA.n999 VDDA.n885 1.17314
R2300 VDDA.n857 VDDA.n856 1.14633
R2301 VDDA.n743 VDDA.n244 1.14633
R2302 VDDA.n847 VDDA.n845 1.06821
R2303 VDDA.n241 VDDA.n233 1.06821
R2304 VDDA.n402 VDDA.n401 0.943208
R2305 VDDA.n755 VDDA.n752 0.932792
R2306 VDDA.n821 VDDA.n800 0.932792
R2307 VDDA.n877 VDDA.n876 0.885917
R2308 VDDA.n736 VDDA.n727 0.885917
R2309 VDDA.n539 VDDA.n538 0.880708
R2310 VDDA.n462 VDDA.n461 0.865083
R2311 VDDA.n589 VDDA.n588 0.807792
R2312 VDDA.n394 VDDA.n393 0.75233
R2313 VDDA.n468 VDDA.n467 0.672375
R2314 VDDA.n395 VDDA.n394 0.648711
R2315 VDDA.n860 VDDA.n822 0.495292
R2316 VDDA.n747 VDDA.n746 0.495292
R2317 VDDA.n595 VDDA.n594 0.448417
R2318 VDDA.n790 VDDA.n789 0.417167
R2319 VDDA.n817 VDDA.n804 0.3755
R2320 VDDA.n806 VDDA.n804 0.3755
R2321 VDDA.n808 VDDA.n806 0.3755
R2322 VDDA.n810 VDDA.n808 0.3755
R2323 VDDA.n812 VDDA.n810 0.3755
R2324 VDDA.n201 VDDA.n199 0.3755
R2325 VDDA.n199 VDDA.n197 0.3755
R2326 VDDA.n197 VDDA.n195 0.3755
R2327 VDDA.n195 VDDA.n193 0.3755
R2328 VDDA.n206 VDDA.n193 0.3755
R2329 VDDA.n452 VDDA.n451 0.333833
R2330 VDDA.n533 VDDA.n532 0.328625
R2331 VDDA.n229 VDDA.n228 0.323417
R2332 VDDA.n843 VDDA.n842 0.323417
R2333 VDDA.n586 VDDA.n585 0.292167
R2334 VDDA.n580 VDDA.n579 0.292167
R2335 VDDA.n573 VDDA.n572 0.292167
R2336 VDDA.n545 VDDA.n544 0.292167
R2337 VDDA.n239 VDDA.n238 0.266125
R2338 VDDA.n854 VDDA.n853 0.266125
R2339 VDDA.n871 VDDA.n862 0.266125
R2340 VDDA.n742 VDDA.n741 0.266125
R2341 VDDA.n450 VDDA.n449 0.2505
R2342 VDDA.n460 VDDA.n459 0.2505
R2343 VDDA.n286 VDDA.n285 0.229667
R2344 VDDA.n305 VDDA.n304 0.229667
R2345 VDDA.n538 VDDA.n533 0.229667
R2346 VDDA.n773 VDDA.n769 0.214042
R2347 VDDA.n783 VDDA.n782 0.214042
R2348 VDDA.n291 VDDA.n283 0.208833
R2349 VDDA.n287 VDDA.n283 0.208833
R2350 VDDA.n287 VDDA.n286 0.208833
R2351 VDDA.n300 VDDA.n299 0.208833
R2352 VDDA.n300 VDDA.n277 0.208833
R2353 VDDA.n304 VDDA.n277 0.208833
R2354 VDDA.n500 VDDA.n486 0.208833
R2355 VDDA.n494 VDDA.n486 0.208833
R2356 VDDA.n494 VDDA.n493 0.208833
R2357 VDDA.n509 VDDA.n507 0.208833
R2358 VDDA.n510 VDDA.n509 0.208833
R2359 VDDA.n510 VDDA.n479 0.208833
R2360 VDDA.n532 VDDA.n531 0.188
R2361 VDDA.n531 VDDA.n530 0.188
R2362 VDDA.n530 VDDA.n529 0.188
R2363 VDDA.n529 VDDA.n528 0.188
R2364 VDDA.n528 VDDA.n527 0.188
R2365 VDDA.n527 VDDA.n526 0.188
R2366 VDDA.n526 VDDA.n525 0.188
R2367 VDDA.n525 VDDA.n524 0.188
R2368 VDDA.n757 VDDA.n755 0.172375
R2369 VDDA.n792 VDDA.n757 0.172375
R2370 VDDA.n758 VDDA.n187 0.172375
R2371 VDDA.n800 VDDA.n187 0.172375
R2372 VDDA.t415 VDDA.t159 0.1603
R2373 VDDA.t387 VDDA.t128 0.1603
R2374 VDDA.t152 VDDA.t418 0.1603
R2375 VDDA.t82 VDDA.t43 0.1603
R2376 VDDA.t129 VDDA.t369 0.1603
R2377 VDDA.n43 VDDA.t15 0.159278
R2378 VDDA.n44 VDDA.t153 0.159278
R2379 VDDA.n45 VDDA.t388 0.159278
R2380 VDDA.n46 VDDA.t72 0.159278
R2381 VDDA.n310 VDDA.n309 0.146333
R2382 VDDA.n310 VDDA.n273 0.146333
R2383 VDDA.n318 VDDA.n273 0.146333
R2384 VDDA.n328 VDDA.n271 0.146333
R2385 VDDA.n329 VDDA.n328 0.146333
R2386 VDDA.n330 VDDA.n329 0.146333
R2387 VDDA.n340 VDDA.n339 0.146333
R2388 VDDA.n340 VDDA.n267 0.146333
R2389 VDDA.n348 VDDA.n267 0.146333
R2390 VDDA.n358 VDDA.n265 0.146333
R2391 VDDA.n313 VDDA.n274 0.146333
R2392 VDDA.n314 VDDA.n313 0.146333
R2393 VDDA.n317 VDDA.n314 0.146333
R2394 VDDA.n327 VDDA.n324 0.146333
R2395 VDDA.n327 VDDA.n270 0.146333
R2396 VDDA.n333 VDDA.n270 0.146333
R2397 VDDA.n343 VDDA.n268 0.146333
R2398 VDDA.n344 VDDA.n343 0.146333
R2399 VDDA.n347 VDDA.n344 0.146333
R2400 VDDA.n357 VDDA.n354 0.146333
R2401 VDDA.n357 VDDA.n264 0.146333
R2402 VDDA.n53 VDDA.n41 0.146333
R2403 VDDA.n54 VDDA.n53 0.146333
R2404 VDDA.n57 VDDA.n54 0.146333
R2405 VDDA.n67 VDDA.n64 0.146333
R2406 VDDA.n67 VDDA.n37 0.146333
R2407 VDDA.n73 VDDA.n37 0.146333
R2408 VDDA.n83 VDDA.n35 0.146333
R2409 VDDA.n84 VDDA.n83 0.146333
R2410 VDDA.n87 VDDA.n84 0.146333
R2411 VDDA.n97 VDDA.n94 0.146333
R2412 VDDA.n97 VDDA.n31 0.146333
R2413 VDDA.n598 VDDA.n384 0.146333
R2414 VDDA.n599 VDDA.n598 0.146333
R2415 VDDA.n602 VDDA.n599 0.146333
R2416 VDDA.n612 VDDA.n609 0.146333
R2417 VDDA.n612 VDDA.n380 0.146333
R2418 VDDA.n618 VDDA.n380 0.146333
R2419 VDDA.n628 VDDA.n378 0.146333
R2420 VDDA.n629 VDDA.n628 0.146333
R2421 VDDA.n632 VDDA.n629 0.146333
R2422 VDDA.n642 VDDA.n639 0.146333
R2423 VDDA.n642 VDDA.n374 0.146333
R2424 VDDA.n137 VDDA.n132 0.146333
R2425 VDDA.n138 VDDA.n137 0.146333
R2426 VDDA.n141 VDDA.n138 0.146333
R2427 VDDA.n149 VDDA.n146 0.146333
R2428 VDDA.n149 VDDA.n124 0.146333
R2429 VDDA.n153 VDDA.n124 0.146333
R2430 VDDA.n161 VDDA.n120 0.146333
R2431 VDDA.n162 VDDA.n161 0.146333
R2432 VDDA.n165 VDDA.n162 0.146333
R2433 VDDA.n173 VDDA.n170 0.146333
R2434 VDDA.n173 VDDA.n114 0.146333
R2435 VDDA.n883 VDDA.n114 0.146333
R2436 VDDA.n714 VDDA.n658 0.146333
R2437 VDDA.n714 VDDA.n713 0.146333
R2438 VDDA.n713 VDDA.n710 0.146333
R2439 VDDA.n705 VDDA.n702 0.146333
R2440 VDDA.n702 VDDA.n701 0.146333
R2441 VDDA.n701 VDDA.n698 0.146333
R2442 VDDA.n693 VDDA.n690 0.146333
R2443 VDDA.n690 VDDA.n689 0.146333
R2444 VDDA.n689 VDDA.n686 0.146333
R2445 VDDA.n681 VDDA.n678 0.146333
R2446 VDDA.n678 VDDA.n250 0.146333
R2447 VDDA.n720 VDDA.n250 0.146333
R2448 VDDA.n46 VDDA.t83 0.1368
R2449 VDDA.n46 VDDA.t415 0.1368
R2450 VDDA.n45 VDDA.t44 0.1368
R2451 VDDA.n45 VDDA.t387 0.1368
R2452 VDDA.n44 VDDA.t142 0.1368
R2453 VDDA.n44 VDDA.t152 0.1368
R2454 VDDA.n43 VDDA.t14 0.1368
R2455 VDDA.n43 VDDA.t82 0.1368
R2456 VDDA.n42 VDDA.t127 0.1368
R2457 VDDA.n42 VDDA.t129 0.1368
R2458 VDDA.n309 VDDA.n308 0.135917
R2459 VDDA.n319 VDDA.n318 0.135917
R2460 VDDA.n320 VDDA.n271 0.135917
R2461 VDDA.n330 VDDA.n269 0.135917
R2462 VDDA.n339 VDDA.n338 0.135917
R2463 VDDA.n349 VDDA.n348 0.135917
R2464 VDDA.n350 VDDA.n265 0.135917
R2465 VDDA.n307 VDDA.n274 0.135917
R2466 VDDA.n317 VDDA.n272 0.135917
R2467 VDDA.n324 VDDA.n323 0.135917
R2468 VDDA.n334 VDDA.n333 0.135917
R2469 VDDA.n337 VDDA.n268 0.135917
R2470 VDDA.n347 VDDA.n266 0.135917
R2471 VDDA.n354 VDDA.n353 0.135917
R2472 VDDA.n47 VDDA.n41 0.135917
R2473 VDDA.n57 VDDA.n39 0.135917
R2474 VDDA.n64 VDDA.n63 0.135917
R2475 VDDA.n74 VDDA.n73 0.135917
R2476 VDDA.n77 VDDA.n35 0.135917
R2477 VDDA.n87 VDDA.n33 0.135917
R2478 VDDA.n94 VDDA.n93 0.135917
R2479 VDDA.n602 VDDA.n382 0.135917
R2480 VDDA.n609 VDDA.n608 0.135917
R2481 VDDA.n619 VDDA.n618 0.135917
R2482 VDDA.n622 VDDA.n378 0.135917
R2483 VDDA.n632 VDDA.n376 0.135917
R2484 VDDA.n639 VDDA.n638 0.135917
R2485 VDDA.n141 VDDA.n128 0.135917
R2486 VDDA.n146 VDDA.n145 0.135917
R2487 VDDA.n154 VDDA.n153 0.135917
R2488 VDDA.n157 VDDA.n120 0.135917
R2489 VDDA.n165 VDDA.n116 0.135917
R2490 VDDA.n170 VDDA.n169 0.135917
R2491 VDDA.n710 VDDA.n709 0.135917
R2492 VDDA.n706 VDDA.n705 0.135917
R2493 VDDA.n698 VDDA.n697 0.135917
R2494 VDDA.n694 VDDA.n693 0.135917
R2495 VDDA.n686 VDDA.n685 0.135917
R2496 VDDA.n682 VDDA.n681 0.135917
R2497 VDDA.n320 VDDA.n319 0.1255
R2498 VDDA.n338 VDDA.n269 0.1255
R2499 VDDA.n350 VDDA.n349 0.1255
R2500 VDDA.n323 VDDA.n272 0.1255
R2501 VDDA.n337 VDDA.n334 0.1255
R2502 VDDA.n353 VDDA.n266 0.1255
R2503 VDDA.n63 VDDA.n39 0.1255
R2504 VDDA.n77 VDDA.n74 0.1255
R2505 VDDA.n93 VDDA.n33 0.1255
R2506 VDDA.n588 VDDA.n587 0.1255
R2507 VDDA.n587 VDDA.n586 0.1255
R2508 VDDA.n461 VDDA.n404 0.1255
R2509 VDDA.n408 VDDA.n404 0.1255
R2510 VDDA.n410 VDDA.n408 0.1255
R2511 VDDA.n412 VDDA.n410 0.1255
R2512 VDDA.n414 VDDA.n412 0.1255
R2513 VDDA.n416 VDDA.n414 0.1255
R2514 VDDA.n418 VDDA.n416 0.1255
R2515 VDDA.n420 VDDA.n418 0.1255
R2516 VDDA.n422 VDDA.n420 0.1255
R2517 VDDA.n452 VDDA.n422 0.1255
R2518 VDDA.n451 VDDA.n424 0.1255
R2519 VDDA.n428 VDDA.n424 0.1255
R2520 VDDA.n430 VDDA.n428 0.1255
R2521 VDDA.n432 VDDA.n430 0.1255
R2522 VDDA.n434 VDDA.n432 0.1255
R2523 VDDA.n436 VDDA.n434 0.1255
R2524 VDDA.n438 VDDA.n436 0.1255
R2525 VDDA.n440 VDDA.n438 0.1255
R2526 VDDA.n442 VDDA.n440 0.1255
R2527 VDDA.n608 VDDA.n382 0.1255
R2528 VDDA.n622 VDDA.n619 0.1255
R2529 VDDA.n638 VDDA.n376 0.1255
R2530 VDDA.n769 VDDA.n763 0.1255
R2531 VDDA.n782 VDDA.n777 0.1255
R2532 VDDA.n145 VDDA.n128 0.1255
R2533 VDDA.n157 VDDA.n154 0.1255
R2534 VDDA.n169 VDDA.n116 0.1255
R2535 VDDA.n709 VDDA.n706 0.1255
R2536 VDDA.n697 VDDA.n694 0.1255
R2537 VDDA.n685 VDDA.n682 0.1255
R2538 VDDA.n306 VDDA.n305 0.123287
R2539 VDDA.n585 VDDA.n584 0.115083
R2540 VDDA.n584 VDDA.n582 0.115083
R2541 VDDA.n582 VDDA.n580 0.115083
R2542 VDDA.n578 VDDA.n577 0.115083
R2543 VDDA.n577 VDDA.n576 0.115083
R2544 VDDA.n576 VDDA.n575 0.115083
R2545 VDDA.n575 VDDA.n574 0.115083
R2546 VDDA.n572 VDDA.n571 0.115083
R2547 VDDA.n571 VDDA.n569 0.115083
R2548 VDDA.n222 VDDA.n220 0.115083
R2549 VDDA.n224 VDDA.n222 0.115083
R2550 VDDA.n226 VDDA.n224 0.115083
R2551 VDDA.n228 VDDA.n226 0.115083
R2552 VDDA.n842 VDDA.n840 0.115083
R2553 VDDA.n840 VDDA.n838 0.115083
R2554 VDDA.n838 VDDA.n836 0.115083
R2555 VDDA.n836 VDDA.n834 0.115083
R2556 VDDA.n871 VDDA.n870 0.115083
R2557 VDDA.n870 VDDA.n868 0.115083
R2558 VDDA.n868 VDDA.n866 0.115083
R2559 VDDA.n866 VDDA.n864 0.115083
R2560 VDDA.n864 VDDA.n181 0.115083
R2561 VDDA.n876 VDDA.n181 0.115083
R2562 VDDA.n736 VDDA.n735 0.115083
R2563 VDDA.n735 VDDA.n733 0.115083
R2564 VDDA.n733 VDDA.n731 0.115083
R2565 VDDA.n731 VDDA.n729 0.115083
R2566 VDDA.n729 VDDA.n246 0.115083
R2567 VDDA.n741 VDDA.n246 0.115083
R2568 VDDA.n646 VDDA.n361 0.107733
R2569 VDDA.n785 VDDA.n775 0.09425
R2570 VDDA.n792 VDDA.n758 0.0838333
R2571 VDDA.n50 VDDA.n49 0.0734167
R2572 VDDA.n50 VDDA.n40 0.0734167
R2573 VDDA.n58 VDDA.n40 0.0734167
R2574 VDDA.n68 VDDA.n38 0.0734167
R2575 VDDA.n69 VDDA.n68 0.0734167
R2576 VDDA.n70 VDDA.n69 0.0734167
R2577 VDDA.n80 VDDA.n79 0.0734167
R2578 VDDA.n80 VDDA.n34 0.0734167
R2579 VDDA.n88 VDDA.n34 0.0734167
R2580 VDDA.n98 VDDA.n32 0.0734167
R2581 VDDA.n596 VDDA.n595 0.0734167
R2582 VDDA.n596 VDDA.n383 0.0734167
R2583 VDDA.n603 VDDA.n383 0.0734167
R2584 VDDA.n613 VDDA.n381 0.0734167
R2585 VDDA.n614 VDDA.n613 0.0734167
R2586 VDDA.n615 VDDA.n614 0.0734167
R2587 VDDA.n625 VDDA.n624 0.0734167
R2588 VDDA.n625 VDDA.n377 0.0734167
R2589 VDDA.n633 VDDA.n377 0.0734167
R2590 VDDA.n643 VDDA.n375 0.0734167
R2591 VDDA.n136 VDDA.n131 0.0734167
R2592 VDDA.n142 VDDA.n131 0.0734167
R2593 VDDA.n150 VDDA.n127 0.0734167
R2594 VDDA.n151 VDDA.n150 0.0734167
R2595 VDDA.n152 VDDA.n151 0.0734167
R2596 VDDA.n160 VDDA.n159 0.0734167
R2597 VDDA.n160 VDDA.n119 0.0734167
R2598 VDDA.n166 VDDA.n119 0.0734167
R2599 VDDA.n174 VDDA.n115 0.0734167
R2600 VDDA.n175 VDDA.n174 0.0734167
R2601 VDDA.n882 VDDA.n175 0.0734167
R2602 VDDA.n660 VDDA.n659 0.0734167
R2603 VDDA.n661 VDDA.n660 0.0734167
R2604 VDDA.n665 VDDA.n664 0.0734167
R2605 VDDA.n666 VDDA.n665 0.0734167
R2606 VDDA.n667 VDDA.n666 0.0734167
R2607 VDDA.n671 VDDA.n670 0.0734167
R2608 VDDA.n672 VDDA.n671 0.0734167
R2609 VDDA.n673 VDDA.n672 0.0734167
R2610 VDDA.n677 VDDA.n676 0.0734167
R2611 VDDA.n677 VDDA.n249 0.0734167
R2612 VDDA.n721 VDDA.n249 0.0734167
R2613 VDDA.n99 VDDA.n31 0.0721864
R2614 VDDA.n644 VDDA.n374 0.0721864
R2615 VDDA.n359 VDDA.n264 0.0716278
R2616 VDDA.n597 VDDA.n372 0.0683791
R2617 VDDA.n49 VDDA.n48 0.0682083
R2618 VDDA.n59 VDDA.n58 0.0682083
R2619 VDDA.n60 VDDA.n38 0.0682083
R2620 VDDA.n70 VDDA.n36 0.0682083
R2621 VDDA.n79 VDDA.n78 0.0682083
R2622 VDDA.n89 VDDA.n88 0.0682083
R2623 VDDA.n90 VDDA.n32 0.0682083
R2624 VDDA.n579 VDDA.n578 0.0682083
R2625 VDDA.n574 VDDA.n573 0.0682083
R2626 VDDA.n604 VDDA.n603 0.0682083
R2627 VDDA.n605 VDDA.n381 0.0682083
R2628 VDDA.n615 VDDA.n379 0.0682083
R2629 VDDA.n624 VDDA.n623 0.0682083
R2630 VDDA.n634 VDDA.n633 0.0682083
R2631 VDDA.n635 VDDA.n375 0.0682083
R2632 VDDA.n143 VDDA.n142 0.0682083
R2633 VDDA.n144 VDDA.n127 0.0682083
R2634 VDDA.n152 VDDA.n123 0.0682083
R2635 VDDA.n159 VDDA.n158 0.0682083
R2636 VDDA.n167 VDDA.n166 0.0682083
R2637 VDDA.n168 VDDA.n115 0.0682083
R2638 VDDA.n662 VDDA.n661 0.0682083
R2639 VDDA.n664 VDDA.n663 0.0682083
R2640 VDDA.n668 VDDA.n667 0.0682083
R2641 VDDA.n670 VDDA.n669 0.0682083
R2642 VDDA.n674 VDDA.n673 0.0682083
R2643 VDDA.n676 VDDA.n675 0.0682083
R2644 VDDA.n135 VDDA.n132 0.0672139
R2645 VDDA.n658 VDDA.n657 0.0672139
R2646 VDDA.n60 VDDA.n59 0.063
R2647 VDDA.n78 VDDA.n36 0.063
R2648 VDDA.n90 VDDA.n89 0.063
R2649 VDDA.n605 VDDA.n604 0.063
R2650 VDDA.n623 VDDA.n379 0.063
R2651 VDDA.n635 VDDA.n634 0.063
R2652 VDDA.n144 VDDA.n143 0.063
R2653 VDDA.n158 VDDA.n123 0.063
R2654 VDDA.n168 VDDA.n167 0.063
R2655 VDDA.n663 VDDA.n662 0.063
R2656 VDDA.n669 VDDA.n668 0.063
R2657 VDDA.n675 VDDA.n674 0.063
R2658 VDDA.n312 VDDA.n311 0.0553333
R2659 VDDA.n316 VDDA.n315 0.0553333
R2660 VDDA.n326 VDDA.n325 0.0553333
R2661 VDDA.n332 VDDA.n331 0.0553333
R2662 VDDA.n342 VDDA.n341 0.0553333
R2663 VDDA.n346 VDDA.n345 0.0553333
R2664 VDDA.n356 VDDA.n355 0.0553333
R2665 VDDA.n360 VDDA.n263 0.0553333
R2666 VDDA.n52 VDDA.n51 0.0553333
R2667 VDDA.n56 VDDA.n55 0.0553333
R2668 VDDA.n66 VDDA.n65 0.0553333
R2669 VDDA.n72 VDDA.n71 0.0553333
R2670 VDDA.n82 VDDA.n81 0.0553333
R2671 VDDA.n86 VDDA.n85 0.0553333
R2672 VDDA.n96 VDDA.n95 0.0553333
R2673 VDDA.n100 VDDA.n30 0.0553333
R2674 VDDA.n601 VDDA.n600 0.0553333
R2675 VDDA.n611 VDDA.n610 0.0553333
R2676 VDDA.n617 VDDA.n616 0.0553333
R2677 VDDA.n627 VDDA.n626 0.0553333
R2678 VDDA.n631 VDDA.n630 0.0553333
R2679 VDDA.n641 VDDA.n640 0.0553333
R2680 VDDA.n645 VDDA.n373 0.0553333
R2681 VDDA.n134 VDDA.n133 0.0553333
R2682 VDDA.n140 VDDA.n139 0.0553333
R2683 VDDA.n148 VDDA.n147 0.0553333
R2684 VDDA.n126 VDDA.n125 0.0553333
R2685 VDDA.n122 VDDA.n121 0.0553333
R2686 VDDA.n164 VDDA.n163 0.0553333
R2687 VDDA.n172 VDDA.n171 0.0553333
R2688 VDDA.n884 VDDA.n113 0.0553333
R2689 VDDA.n716 VDDA.n715 0.0553333
R2690 VDDA.n712 VDDA.n711 0.0553333
R2691 VDDA.n704 VDDA.n703 0.0553333
R2692 VDDA.n700 VDDA.n699 0.0553333
R2693 VDDA.n692 VDDA.n691 0.0553333
R2694 VDDA.n688 VDDA.n687 0.0553333
R2695 VDDA.n680 VDDA.n679 0.0553333
R2696 VDDA.n719 VDDA.n251 0.0553333
R2697 VDDA.n322 VDDA.n321 0.0475
R2698 VDDA.n336 VDDA.n335 0.0475
R2699 VDDA.n352 VDDA.n351 0.0475
R2700 VDDA.n62 VDDA.n61 0.0475
R2701 VDDA.n76 VDDA.n75 0.0475
R2702 VDDA.n92 VDDA.n91 0.0475
R2703 VDDA.n607 VDDA.n606 0.0475
R2704 VDDA.n621 VDDA.n620 0.0475
R2705 VDDA.n637 VDDA.n636 0.0475
R2706 VDDA.n130 VDDA.n129 0.0475
R2707 VDDA.n156 VDDA.n155 0.0475
R2708 VDDA.n118 VDDA.n117 0.0475
R2709 VDDA.n708 VDDA.n707 0.0475
R2710 VDDA.n696 VDDA.n695 0.0475
R2711 VDDA.n684 VDDA.n683 0.0475
R2712 VDDA.n791 VDDA.n189 0.0429747
R2713 VDDA.n879 VDDA.n178 0.0421667
R2714 VDDA.n802 VDDA.n185 0.0421667
R2715 VDDA.n744 VDDA.n210 0.0421667
R2716 VDDA.n361 VDDA.n101 0.0287913
R2717 VDDA.n885 VDDA.n101 0.0286392
R2718 VDDA.n718 VDDA.n646 0.0284871
R2719 VDDA.n315 VDDA.n261 0.028198
R2720 VDDA.n331 VDDA.n258 0.028198
R2721 VDDA.n345 VDDA.n255 0.028198
R2722 VDDA.n263 VDDA.n252 0.028198
R2723 VDDA.n55 VDDA.n28 0.028198
R2724 VDDA.n71 VDDA.n25 0.028198
R2725 VDDA.n85 VDDA.n22 0.028198
R2726 VDDA.n30 VDDA.n19 0.028198
R2727 VDDA.n600 VDDA.n371 0.028198
R2728 VDDA.n616 VDDA.n368 0.028198
R2729 VDDA.n630 VDDA.n365 0.028198
R2730 VDDA.n373 VDDA.n362 0.028198
R2731 VDDA.n139 VDDA.n111 0.028198
R2732 VDDA.n125 VDDA.n108 0.028198
R2733 VDDA.n163 VDDA.n105 0.028198
R2734 VDDA.n113 VDDA.n102 0.028198
R2735 VDDA.n712 VDDA.n656 0.028198
R2736 VDDA.n700 VDDA.n653 0.028198
R2737 VDDA.n688 VDDA.n650 0.028198
R2738 VDDA.n647 VDDA.n251 0.028198
R2739 VDDA.n679 VDDA.n647 0.028198
R2740 VDDA.n691 VDDA.n650 0.028198
R2741 VDDA.n703 VDDA.n653 0.028198
R2742 VDDA.n715 VDDA.n656 0.028198
R2743 VDDA.n641 VDDA.n362 0.028198
R2744 VDDA.n627 VDDA.n365 0.028198
R2745 VDDA.n611 VDDA.n368 0.028198
R2746 VDDA.n597 VDDA.n371 0.028198
R2747 VDDA.n172 VDDA.n102 0.028198
R2748 VDDA.n122 VDDA.n105 0.028198
R2749 VDDA.n148 VDDA.n108 0.028198
R2750 VDDA.n134 VDDA.n111 0.028198
R2751 VDDA.n96 VDDA.n19 0.028198
R2752 VDDA.n82 VDDA.n22 0.028198
R2753 VDDA.n66 VDDA.n25 0.028198
R2754 VDDA.n52 VDDA.n28 0.028198
R2755 VDDA.n356 VDDA.n252 0.028198
R2756 VDDA.n342 VDDA.n255 0.028198
R2757 VDDA.n326 VDDA.n258 0.028198
R2758 VDDA.n312 VDDA.n261 0.028198
R2759 VDDA.n311 VDDA.n262 0.0262697
R2760 VDDA.n321 VDDA.n260 0.0262697
R2761 VDDA.n325 VDDA.n259 0.0262697
R2762 VDDA.n335 VDDA.n257 0.0262697
R2763 VDDA.n341 VDDA.n256 0.0262697
R2764 VDDA.n351 VDDA.n254 0.0262697
R2765 VDDA.n355 VDDA.n253 0.0262697
R2766 VDDA.n51 VDDA.n29 0.0262697
R2767 VDDA.n61 VDDA.n27 0.0262697
R2768 VDDA.n65 VDDA.n26 0.0262697
R2769 VDDA.n75 VDDA.n24 0.0262697
R2770 VDDA.n81 VDDA.n23 0.0262697
R2771 VDDA.n91 VDDA.n21 0.0262697
R2772 VDDA.n95 VDDA.n20 0.0262697
R2773 VDDA.n606 VDDA.n370 0.0262697
R2774 VDDA.n610 VDDA.n369 0.0262697
R2775 VDDA.n620 VDDA.n367 0.0262697
R2776 VDDA.n626 VDDA.n366 0.0262697
R2777 VDDA.n636 VDDA.n364 0.0262697
R2778 VDDA.n640 VDDA.n363 0.0262697
R2779 VDDA.n133 VDDA.n112 0.0262697
R2780 VDDA.n129 VDDA.n110 0.0262697
R2781 VDDA.n147 VDDA.n109 0.0262697
R2782 VDDA.n155 VDDA.n107 0.0262697
R2783 VDDA.n121 VDDA.n106 0.0262697
R2784 VDDA.n117 VDDA.n104 0.0262697
R2785 VDDA.n171 VDDA.n103 0.0262697
R2786 VDDA.n717 VDDA.n716 0.0262697
R2787 VDDA.n708 VDDA.n655 0.0262697
R2788 VDDA.n704 VDDA.n654 0.0262697
R2789 VDDA.n696 VDDA.n652 0.0262697
R2790 VDDA.n692 VDDA.n651 0.0262697
R2791 VDDA.n684 VDDA.n649 0.0262697
R2792 VDDA.n680 VDDA.n648 0.0262697
R2793 VDDA.n683 VDDA.n648 0.0262697
R2794 VDDA.n687 VDDA.n649 0.0262697
R2795 VDDA.n695 VDDA.n651 0.0262697
R2796 VDDA.n699 VDDA.n652 0.0262697
R2797 VDDA.n707 VDDA.n654 0.0262697
R2798 VDDA.n711 VDDA.n655 0.0262697
R2799 VDDA.n637 VDDA.n363 0.0262697
R2800 VDDA.n631 VDDA.n364 0.0262697
R2801 VDDA.n621 VDDA.n366 0.0262697
R2802 VDDA.n617 VDDA.n367 0.0262697
R2803 VDDA.n607 VDDA.n369 0.0262697
R2804 VDDA.n601 VDDA.n370 0.0262697
R2805 VDDA.n118 VDDA.n103 0.0262697
R2806 VDDA.n164 VDDA.n104 0.0262697
R2807 VDDA.n156 VDDA.n106 0.0262697
R2808 VDDA.n126 VDDA.n107 0.0262697
R2809 VDDA.n130 VDDA.n109 0.0262697
R2810 VDDA.n140 VDDA.n110 0.0262697
R2811 VDDA.n92 VDDA.n20 0.0262697
R2812 VDDA.n86 VDDA.n21 0.0262697
R2813 VDDA.n76 VDDA.n23 0.0262697
R2814 VDDA.n72 VDDA.n24 0.0262697
R2815 VDDA.n62 VDDA.n26 0.0262697
R2816 VDDA.n56 VDDA.n27 0.0262697
R2817 VDDA.n352 VDDA.n253 0.0262697
R2818 VDDA.n346 VDDA.n254 0.0262697
R2819 VDDA.n336 VDDA.n256 0.0262697
R2820 VDDA.n332 VDDA.n257 0.0262697
R2821 VDDA.n322 VDDA.n259 0.0262697
R2822 VDDA.n316 VDDA.n260 0.0262697
R2823 VDDA.n589 VDDA.n385 0.0217373
R2824 VDDA.n539 VDDA.n387 0.0217373
R2825 VDDA.n462 VDDA.n389 0.0217373
R2826 VDDA.n396 VDDA.n391 0.0217373
R2827 VDDA.n400 VDDA.n399 0.0217373
R2828 VDDA.n466 VDDA.n465 0.0217373
R2829 VDDA.n543 VDDA.n542 0.0217373
R2830 VDDA.n593 VDDA.n592 0.0217373
R2831 VDDA.n398 VDDA.n391 0.0217373
R2832 VDDA.n401 VDDA.n400 0.0217373
R2833 VDDA.n464 VDDA.n389 0.0217373
R2834 VDDA.n467 VDDA.n466 0.0217373
R2835 VDDA.n541 VDDA.n387 0.0217373
R2836 VDDA.n544 VDDA.n543 0.0217373
R2837 VDDA.n591 VDDA.n385 0.0217373
R2838 VDDA.n594 VDDA.n593 0.0217373
R2839 VDDA.n774 VDDA.n773 0.0217373
R2840 VDDA.n770 VDDA.n762 0.0217373
R2841 VDDA.n784 VDDA.n760 0.0217373
R2842 VDDA.n775 VDDA.n761 0.0217373
R2843 VDDA.n789 VDDA.n759 0.0217373
R2844 VDDA.n793 VDDA.n189 0.0217373
R2845 VDDA.n788 VDDA.n760 0.0217373
R2846 VDDA.n786 VDDA.n759 0.0217373
R2847 VDDA.n784 VDDA.n783 0.0217373
R2848 VDDA.n774 VDDA.n762 0.0217373
R2849 VDDA.n771 VDDA.n761 0.0217373
R2850 VDDA.n843 VDDA.n831 0.0217373
R2851 VDDA.n854 VDDA.n848 0.0217373
R2852 VDDA.n881 VDDA.n880 0.0217373
R2853 VDDA.n878 VDDA.n179 0.0217373
R2854 VDDA.n862 VDDA.n182 0.0217373
R2855 VDDA.n880 VDDA.n177 0.0217373
R2856 VDDA.n179 VDDA.n177 0.0217373
R2857 VDDA.n819 VDDA.n818 0.0217373
R2858 VDDA.n822 VDDA.n184 0.0217373
R2859 VDDA.n858 VDDA.n183 0.0217373
R2860 VDDA.n846 VDDA.n825 0.0217373
R2861 VDDA.n830 VDDA.n828 0.0217373
R2862 VDDA.n823 VDDA.n182 0.0217373
R2863 VDDA.n858 VDDA.n857 0.0217373
R2864 VDDA.n848 VDDA.n826 0.0217373
R2865 VDDA.n847 VDDA.n846 0.0217373
R2866 VDDA.n831 VDDA.n829 0.0217373
R2867 VDDA.n752 VDDA.n190 0.0217373
R2868 VDDA.n818 VDDA.n801 0.0217373
R2869 VDDA.n801 VDDA.n184 0.0217373
R2870 VDDA.n791 VDDA.n790 0.0217373
R2871 VDDA.n748 VDDA.n191 0.0217373
R2872 VDDA.n746 VDDA.n745 0.0217373
R2873 VDDA.n743 VDDA.n211 0.0217373
R2874 VDDA.n240 VDDA.n213 0.0217373
R2875 VDDA.n230 VDDA.n216 0.0217373
R2876 VDDA.n207 VDDA.n190 0.0217373
R2877 VDDA.n748 VDDA.n747 0.0217373
R2878 VDDA.n242 VDDA.n214 0.0217373
R2879 VDDA.n241 VDDA.n240 0.0217373
R2880 VDDA.n231 VDDA.n217 0.0217373
R2881 VDDA.n727 VDDA.n247 0.0217373
R2882 VDDA.n745 VDDA.n209 0.0217373
R2883 VDDA.n211 VDDA.n209 0.0217373
R2884 VDDA.n723 VDDA.n248 0.0217373
R2885 VDDA.n722 VDDA.n247 0.0217373
R2886 VDDA.n591 VDDA.n386 0.0217373
R2887 VDDA.n541 VDDA.n388 0.0217373
R2888 VDDA.n464 VDDA.n390 0.0217373
R2889 VDDA.n398 VDDA.n392 0.0217373
R2890 VDDA.n399 VDDA.n397 0.0217373
R2891 VDDA.n465 VDDA.n463 0.0217373
R2892 VDDA.n542 VDDA.n540 0.0217373
R2893 VDDA.n592 VDDA.n590 0.0217373
R2894 VDDA.n463 VDDA.n402 0.0217373
R2895 VDDA.n540 VDDA.n468 0.0217373
R2896 VDDA.n590 VDDA.n545 0.0217373
R2897 VDDA.n217 VDDA.n215 0.0217373
R2898 VDDA.n214 VDDA.n212 0.0217373
R2899 VDDA.n787 VDDA.n785 0.0217373
R2900 VDDA.n787 VDDA.n786 0.0217373
R2901 VDDA.n772 VDDA.n771 0.0217373
R2902 VDDA.n829 VDDA.n827 0.0217373
R2903 VDDA.n826 VDDA.n824 0.0217373
R2904 VDDA.n859 VDDA.n823 0.0217373
R2905 VDDA.n877 VDDA.n176 0.0217373
R2906 VDDA.n178 VDDA.n176 0.0217373
R2907 VDDA.n861 VDDA.n183 0.0217373
R2908 VDDA.n855 VDDA.n825 0.0217373
R2909 VDDA.n844 VDDA.n828 0.0217373
R2910 VDDA.n861 VDDA.n860 0.0217373
R2911 VDDA.n856 VDDA.n855 0.0217373
R2912 VDDA.n845 VDDA.n844 0.0217373
R2913 VDDA.n749 VDDA.n207 0.0217373
R2914 VDDA.n821 VDDA.n820 0.0217373
R2915 VDDA.n820 VDDA.n802 0.0217373
R2916 VDDA.n751 VDDA.n191 0.0217373
R2917 VDDA.n243 VDDA.n213 0.0217373
R2918 VDDA.n232 VDDA.n216 0.0217373
R2919 VDDA.n751 VDDA.n750 0.0217373
R2920 VDDA.n244 VDDA.n243 0.0217373
R2921 VDDA.n239 VDDA.n212 0.0217373
R2922 VDDA.n233 VDDA.n232 0.0217373
R2923 VDDA.n229 VDDA.n215 0.0217373
R2924 VDDA.n724 VDDA.n722 0.0217373
R2925 VDDA.n742 VDDA.n208 0.0217373
R2926 VDDA.n210 VDDA.n208 0.0217373
R2927 VDDA.n726 VDDA.n248 0.0217373
R2928 VDDA.n726 VDDA.n725 0.0217373
R2929 VDDA VDDA.n1000 0.0164359
R2930 VDDA.n999 VDDA.n902 0.00186893
R2931 VDDA.n902 VDDA.n18 0.00186893
R2932 VDDA.n952 VDDA.n951 0.00168433
R2933 VDDA.n952 VDDA.n1 0.00168433
R2934 VDDA.n996 VDDA.n953 0.00168433
R2935 VDDA.n953 VDDA.n2 0.00168433
R2936 VDDA.n994 VDDA.n954 0.00168433
R2937 VDDA.n954 VDDA.n3 0.00168433
R2938 VDDA.n992 VDDA.n955 0.00168433
R2939 VDDA.n955 VDDA.n4 0.00168433
R2940 VDDA.n990 VDDA.n956 0.00168433
R2941 VDDA.n956 VDDA.n5 0.00168433
R2942 VDDA.n988 VDDA.n957 0.00168433
R2943 VDDA.n957 VDDA.n6 0.00168433
R2944 VDDA.n986 VDDA.n958 0.00168433
R2945 VDDA.n958 VDDA.n7 0.00168433
R2946 VDDA.n984 VDDA.n959 0.00168433
R2947 VDDA.n959 VDDA.n8 0.00168433
R2948 VDDA.n982 VDDA.n960 0.00168433
R2949 VDDA.n960 VDDA.n9 0.00168433
R2950 VDDA.n980 VDDA.n961 0.00168433
R2951 VDDA.n961 VDDA.n10 0.00168433
R2952 VDDA.n978 VDDA.n962 0.00168433
R2953 VDDA.n962 VDDA.n11 0.00168433
R2954 VDDA.n976 VDDA.n963 0.00168433
R2955 VDDA.n963 VDDA.n12 0.00168433
R2956 VDDA.n974 VDDA.n964 0.00168433
R2957 VDDA.n964 VDDA.n13 0.00168433
R2958 VDDA.n972 VDDA.n965 0.00168433
R2959 VDDA.n965 VDDA.n14 0.00168433
R2960 VDDA.n970 VDDA.n966 0.00168433
R2961 VDDA.n966 VDDA.n15 0.00168433
R2962 VDDA.n968 VDDA.n16 0.00168433
R2963 VDDA.n967 VDDA.n17 0.00168433
R2964 VDDA.n969 VDDA.n15 0.00168433
R2965 VDDA.n971 VDDA.n14 0.00168433
R2966 VDDA.n973 VDDA.n13 0.00168433
R2967 VDDA.n975 VDDA.n12 0.00168433
R2968 VDDA.n977 VDDA.n11 0.00168433
R2969 VDDA.n979 VDDA.n10 0.00168433
R2970 VDDA.n981 VDDA.n9 0.00168433
R2971 VDDA.n983 VDDA.n8 0.00168433
R2972 VDDA.n985 VDDA.n7 0.00168433
R2973 VDDA.n987 VDDA.n6 0.00168433
R2974 VDDA.n989 VDDA.n5 0.00168433
R2975 VDDA.n991 VDDA.n4 0.00168433
R2976 VDDA.n993 VDDA.n3 0.00168433
R2977 VDDA.n995 VDDA.n2 0.00168433
R2978 VDDA.n997 VDDA.n1 0.00168433
R2979 VDDA.n969 VDDA.n968 0.00168433
R2980 VDDA.n971 VDDA.n970 0.00168433
R2981 VDDA.n973 VDDA.n972 0.00168433
R2982 VDDA.n975 VDDA.n974 0.00168433
R2983 VDDA.n977 VDDA.n976 0.00168433
R2984 VDDA.n979 VDDA.n978 0.00168433
R2985 VDDA.n981 VDDA.n980 0.00168433
R2986 VDDA.n983 VDDA.n982 0.00168433
R2987 VDDA.n985 VDDA.n984 0.00168433
R2988 VDDA.n987 VDDA.n986 0.00168433
R2989 VDDA.n989 VDDA.n988 0.00168433
R2990 VDDA.n991 VDDA.n990 0.00168433
R2991 VDDA.n993 VDDA.n992 0.00168433
R2992 VDDA.n995 VDDA.n994 0.00168433
R2993 VDDA.n997 VDDA.n996 0.00168433
R2994 VDDA.n951 VDDA.n18 0.00168433
R2995 VDDA.n967 VDDA.n16 0.00168433
R2996 VDDA.n904 VDDA.n0 0.00166081
R2997 VDDA.n903 VDDA.n901 0.00166081
R2998 VDDA.n907 VDDA.n905 0.00166081
R2999 VDDA.n906 VDDA.n900 0.00166081
R3000 VDDA.n910 VDDA.n908 0.00166081
R3001 VDDA.n909 VDDA.n899 0.00166081
R3002 VDDA.n913 VDDA.n911 0.00166081
R3003 VDDA.n912 VDDA.n898 0.00166081
R3004 VDDA.n916 VDDA.n914 0.00166081
R3005 VDDA.n915 VDDA.n897 0.00166081
R3006 VDDA.n919 VDDA.n917 0.00166081
R3007 VDDA.n918 VDDA.n896 0.00166081
R3008 VDDA.n922 VDDA.n920 0.00166081
R3009 VDDA.n921 VDDA.n895 0.00166081
R3010 VDDA.n925 VDDA.n923 0.00166081
R3011 VDDA.n924 VDDA.n894 0.00166081
R3012 VDDA.n928 VDDA.n926 0.00166081
R3013 VDDA.n927 VDDA.n893 0.00166081
R3014 VDDA.n931 VDDA.n929 0.00166081
R3015 VDDA.n930 VDDA.n892 0.00166081
R3016 VDDA.n934 VDDA.n932 0.00166081
R3017 VDDA.n933 VDDA.n891 0.00166081
R3018 VDDA.n937 VDDA.n935 0.00166081
R3019 VDDA.n936 VDDA.n890 0.00166081
R3020 VDDA.n940 VDDA.n938 0.00166081
R3021 VDDA.n939 VDDA.n889 0.00166081
R3022 VDDA.n943 VDDA.n941 0.00166081
R3023 VDDA.n942 VDDA.n888 0.00166081
R3024 VDDA.n946 VDDA.n944 0.00166081
R3025 VDDA.n945 VDDA.n887 0.00166081
R3026 VDDA.n949 VDDA.n947 0.00166081
R3027 VDDA.n948 VDDA.n886 0.00166081
R3028 VDDA.n998 VDDA.n950 0.00166081
R3029 VDDA.n1000 VDDA.n0 0.00166081
R3030 VDDA.n904 VDDA.n903 0.00166081
R3031 VDDA.n905 VDDA.n901 0.00166081
R3032 VDDA.n907 VDDA.n906 0.00166081
R3033 VDDA.n908 VDDA.n900 0.00166081
R3034 VDDA.n910 VDDA.n909 0.00166081
R3035 VDDA.n911 VDDA.n899 0.00166081
R3036 VDDA.n913 VDDA.n912 0.00166081
R3037 VDDA.n914 VDDA.n898 0.00166081
R3038 VDDA.n916 VDDA.n915 0.00166081
R3039 VDDA.n917 VDDA.n897 0.00166081
R3040 VDDA.n919 VDDA.n918 0.00166081
R3041 VDDA.n920 VDDA.n896 0.00166081
R3042 VDDA.n922 VDDA.n921 0.00166081
R3043 VDDA.n923 VDDA.n895 0.00166081
R3044 VDDA.n925 VDDA.n924 0.00166081
R3045 VDDA.n926 VDDA.n894 0.00166081
R3046 VDDA.n928 VDDA.n927 0.00166081
R3047 VDDA.n929 VDDA.n893 0.00166081
R3048 VDDA.n931 VDDA.n930 0.00166081
R3049 VDDA.n932 VDDA.n892 0.00166081
R3050 VDDA.n934 VDDA.n933 0.00166081
R3051 VDDA.n935 VDDA.n891 0.00166081
R3052 VDDA.n937 VDDA.n936 0.00166081
R3053 VDDA.n938 VDDA.n890 0.00166081
R3054 VDDA.n940 VDDA.n939 0.00166081
R3055 VDDA.n941 VDDA.n889 0.00166081
R3056 VDDA.n943 VDDA.n942 0.00166081
R3057 VDDA.n944 VDDA.n888 0.00166081
R3058 VDDA.n946 VDDA.n945 0.00166081
R3059 VDDA.n947 VDDA.n887 0.00166081
R3060 VDDA.n949 VDDA.n948 0.00166081
R3061 VDDA.n950 VDDA.n886 0.00166081
R3062 VDDA.t15 VDDA.n42 0.00152174
R3063 VDDA.t153 VDDA.n43 0.00152174
R3064 VDDA.t388 VDDA.n44 0.00152174
R3065 VDDA.t72 VDDA.n45 0.00152174
R3066 VDDA.t141 VDDA.n46 0.00152174
R3067 two_stage_opamp_dummy_magic_29_0.Vb3.n15 two_stage_opamp_dummy_magic_29_0.Vb3.t19 793.28
R3068 two_stage_opamp_dummy_magic_29_0.Vb3.n8 two_stage_opamp_dummy_magic_29_0.Vb3.t18 752.422
R3069 two_stage_opamp_dummy_magic_29_0.Vb3.n0 two_stage_opamp_dummy_magic_29_0.Vb3.t23 752.422
R3070 two_stage_opamp_dummy_magic_29_0.Vb3.n8 two_stage_opamp_dummy_magic_29_0.Vb3.t11 752.234
R3071 two_stage_opamp_dummy_magic_29_0.Vb3.n8 two_stage_opamp_dummy_magic_29_0.Vb3.t22 752.234
R3072 two_stage_opamp_dummy_magic_29_0.Vb3.n7 two_stage_opamp_dummy_magic_29_0.Vb3.t8 752.234
R3073 two_stage_opamp_dummy_magic_29_0.Vb3.n5 two_stage_opamp_dummy_magic_29_0.Vb3.t20 752.234
R3074 two_stage_opamp_dummy_magic_29_0.Vb3.n6 two_stage_opamp_dummy_magic_29_0.Vb3.t9 752.234
R3075 two_stage_opamp_dummy_magic_29_0.Vb3.n6 two_stage_opamp_dummy_magic_29_0.Vb3.t15 752.234
R3076 two_stage_opamp_dummy_magic_29_0.Vb3.n19 two_stage_opamp_dummy_magic_29_0.Vb3.t25 752.234
R3077 two_stage_opamp_dummy_magic_29_0.Vb3.n4 two_stage_opamp_dummy_magic_29_0.Vb3.t16 752.234
R3078 two_stage_opamp_dummy_magic_29_0.Vb3.n4 two_stage_opamp_dummy_magic_29_0.Vb3.t26 752.234
R3079 two_stage_opamp_dummy_magic_29_0.Vb3.n3 two_stage_opamp_dummy_magic_29_0.Vb3.t21 752.234
R3080 two_stage_opamp_dummy_magic_29_0.Vb3.n3 two_stage_opamp_dummy_magic_29_0.Vb3.t10 752.234
R3081 two_stage_opamp_dummy_magic_29_0.Vb3.n0 two_stage_opamp_dummy_magic_29_0.Vb3.t12 752.234
R3082 two_stage_opamp_dummy_magic_29_0.Vb3.n0 two_stage_opamp_dummy_magic_29_0.Vb3.t28 752.234
R3083 two_stage_opamp_dummy_magic_29_0.Vb3.n0 two_stage_opamp_dummy_magic_29_0.Vb3.t13 752.234
R3084 two_stage_opamp_dummy_magic_29_0.Vb3.n17 two_stage_opamp_dummy_magic_29_0.Vb3.t14 747.734
R3085 two_stage_opamp_dummy_magic_29_0.Vb3.n18 two_stage_opamp_dummy_magic_29_0.Vb3.t24 747.734
R3086 two_stage_opamp_dummy_magic_29_0.Vb3.n2 two_stage_opamp_dummy_magic_29_0.Vb3.t27 747.827
R3087 two_stage_opamp_dummy_magic_29_0.Vb3.n11 two_stage_opamp_dummy_magic_29_0.Vb3.n9 139.639
R3088 two_stage_opamp_dummy_magic_29_0.Vb3.n11 two_stage_opamp_dummy_magic_29_0.Vb3.n10 139.638
R3089 two_stage_opamp_dummy_magic_29_0.Vb3.n13 two_stage_opamp_dummy_magic_29_0.Vb3.n12 134.577
R3090 two_stage_opamp_dummy_magic_29_0.Vb3.n15 two_stage_opamp_dummy_magic_29_0.Vb3.n14 72.612
R3091 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_29_0.Vb3.n13 43.0317
R3092 bgr_11_0.VB3_CUR_BIAS two_stage_opamp_dummy_magic_29_0.Vb3.n20 35.0317
R3093 two_stage_opamp_dummy_magic_29_0.Vb3.n12 two_stage_opamp_dummy_magic_29_0.Vb3.t6 24.0005
R3094 two_stage_opamp_dummy_magic_29_0.Vb3.n12 two_stage_opamp_dummy_magic_29_0.Vb3.t5 24.0005
R3095 two_stage_opamp_dummy_magic_29_0.Vb3.n10 two_stage_opamp_dummy_magic_29_0.Vb3.t3 24.0005
R3096 two_stage_opamp_dummy_magic_29_0.Vb3.n10 two_stage_opamp_dummy_magic_29_0.Vb3.t1 24.0005
R3097 two_stage_opamp_dummy_magic_29_0.Vb3.n9 two_stage_opamp_dummy_magic_29_0.Vb3.t2 24.0005
R3098 two_stage_opamp_dummy_magic_29_0.Vb3.n9 two_stage_opamp_dummy_magic_29_0.Vb3.t4 24.0005
R3099 two_stage_opamp_dummy_magic_29_0.Vb3.n14 two_stage_opamp_dummy_magic_29_0.Vb3.t7 11.2576
R3100 two_stage_opamp_dummy_magic_29_0.Vb3.n14 two_stage_opamp_dummy_magic_29_0.Vb3.t0 11.2576
R3101 two_stage_opamp_dummy_magic_29_0.Vb3.n16 two_stage_opamp_dummy_magic_29_0.Vb3.n15 11.2036
R3102 two_stage_opamp_dummy_magic_29_0.Vb3.n20 two_stage_opamp_dummy_magic_29_0.Vb3.n16 6.14112
R3103 two_stage_opamp_dummy_magic_29_0.Vb3.n13 two_stage_opamp_dummy_magic_29_0.Vb3.n11 4.5005
R3104 two_stage_opamp_dummy_magic_29_0.Vb3.n1 two_stage_opamp_dummy_magic_29_0.Vb3.n2 2.20508
R3105 two_stage_opamp_dummy_magic_29_0.Vb3.n5 two_stage_opamp_dummy_magic_29_0.Vb3.n18 4.5005
R3106 two_stage_opamp_dummy_magic_29_0.Vb3.n17 two_stage_opamp_dummy_magic_29_0.Vb3.n7 4.5005
R3107 two_stage_opamp_dummy_magic_29_0.Vb3.n16 two_stage_opamp_dummy_magic_29_0.Vb3.n4 3.21925
R3108 two_stage_opamp_dummy_magic_29_0.Vb3.n20 two_stage_opamp_dummy_magic_29_0.Vb3.n19 0.641125
R3109 two_stage_opamp_dummy_magic_29_0.Vb3.n7 two_stage_opamp_dummy_magic_29_0.Vb3.n8 0.3755
R3110 two_stage_opamp_dummy_magic_29_0.Vb3.n5 two_stage_opamp_dummy_magic_29_0.Vb3.n7 0.3755
R3111 two_stage_opamp_dummy_magic_29_0.Vb3.n6 two_stage_opamp_dummy_magic_29_0.Vb3.n5 0.3755
R3112 two_stage_opamp_dummy_magic_29_0.Vb3.n19 two_stage_opamp_dummy_magic_29_0.Vb3.n6 0.3755
R3113 two_stage_opamp_dummy_magic_29_0.Vb3.n4 two_stage_opamp_dummy_magic_29_0.Vb3.n3 0.3755
R3114 two_stage_opamp_dummy_magic_29_0.Vb3.n3 two_stage_opamp_dummy_magic_29_0.Vb3.n1 0.3755
R3115 two_stage_opamp_dummy_magic_29_0.Vb3.n18 two_stage_opamp_dummy_magic_29_0.Vb3.n17 0.188
R3116 two_stage_opamp_dummy_magic_29_0.Vb3.t17 two_stage_opamp_dummy_magic_29_0.Vb3.n2 747.827
R3117 two_stage_opamp_dummy_magic_29_0.Vb3.n1 two_stage_opamp_dummy_magic_29_0.Vb3.n0 0.7505
R3118 two_stage_opamp_dummy_magic_29_0.VD4.n20 two_stage_opamp_dummy_magic_29_0.VD4.t32 671.418
R3119 two_stage_opamp_dummy_magic_29_0.VD4.n17 two_stage_opamp_dummy_magic_29_0.VD4.t35 671.418
R3120 two_stage_opamp_dummy_magic_29_0.VD4.t36 two_stage_opamp_dummy_magic_29_0.VD4.n18 213.131
R3121 two_stage_opamp_dummy_magic_29_0.VD4.n19 two_stage_opamp_dummy_magic_29_0.VD4.t33 213.131
R3122 two_stage_opamp_dummy_magic_29_0.VD4.t2 two_stage_opamp_dummy_magic_29_0.VD4.t36 146.155
R3123 two_stage_opamp_dummy_magic_29_0.VD4.t12 two_stage_opamp_dummy_magic_29_0.VD4.t2 146.155
R3124 two_stage_opamp_dummy_magic_29_0.VD4.t8 two_stage_opamp_dummy_magic_29_0.VD4.t12 146.155
R3125 two_stage_opamp_dummy_magic_29_0.VD4.t0 two_stage_opamp_dummy_magic_29_0.VD4.t8 146.155
R3126 two_stage_opamp_dummy_magic_29_0.VD4.t4 two_stage_opamp_dummy_magic_29_0.VD4.t0 146.155
R3127 two_stage_opamp_dummy_magic_29_0.VD4.t10 two_stage_opamp_dummy_magic_29_0.VD4.t4 146.155
R3128 two_stage_opamp_dummy_magic_29_0.VD4.t14 two_stage_opamp_dummy_magic_29_0.VD4.t10 146.155
R3129 two_stage_opamp_dummy_magic_29_0.VD4.t16 two_stage_opamp_dummy_magic_29_0.VD4.t14 146.155
R3130 two_stage_opamp_dummy_magic_29_0.VD4.t6 two_stage_opamp_dummy_magic_29_0.VD4.t16 146.155
R3131 two_stage_opamp_dummy_magic_29_0.VD4.t18 two_stage_opamp_dummy_magic_29_0.VD4.t6 146.155
R3132 two_stage_opamp_dummy_magic_29_0.VD4.t33 two_stage_opamp_dummy_magic_29_0.VD4.t18 146.155
R3133 two_stage_opamp_dummy_magic_29_0.VD4.n18 two_stage_opamp_dummy_magic_29_0.VD4.t37 76.2576
R3134 two_stage_opamp_dummy_magic_29_0.VD4.n19 two_stage_opamp_dummy_magic_29_0.VD4.t34 76.2576
R3135 two_stage_opamp_dummy_magic_29_0.VD4.n0 two_stage_opamp_dummy_magic_29_0.VD4.n10 67.013
R3136 two_stage_opamp_dummy_magic_29_0.VD4.n1 two_stage_opamp_dummy_magic_29_0.VD4.n4 67.013
R3137 two_stage_opamp_dummy_magic_29_0.VD4.n0 two_stage_opamp_dummy_magic_29_0.VD4.n7 67.013
R3138 two_stage_opamp_dummy_magic_29_0.VD4.n0 two_stage_opamp_dummy_magic_29_0.VD4.n11 67.013
R3139 two_stage_opamp_dummy_magic_29_0.VD4.n3 two_stage_opamp_dummy_magic_29_0.VD4.n16 67.013
R3140 two_stage_opamp_dummy_magic_29_0.VD4.n22 two_stage_opamp_dummy_magic_29_0.VD4.n21 66.0338
R3141 two_stage_opamp_dummy_magic_29_0.VD4.n24 two_stage_opamp_dummy_magic_29_0.VD4.n23 66.0338
R3142 two_stage_opamp_dummy_magic_29_0.VD4.n9 two_stage_opamp_dummy_magic_29_0.VD4.n8 66.0338
R3143 two_stage_opamp_dummy_magic_29_0.VD4.n6 two_stage_opamp_dummy_magic_29_0.VD4.n5 66.0338
R3144 two_stage_opamp_dummy_magic_29_0.VD4.n13 two_stage_opamp_dummy_magic_29_0.VD4.n12 66.0338
R3145 two_stage_opamp_dummy_magic_29_0.VD4.n28 two_stage_opamp_dummy_magic_29_0.VD4.n27 66.0338
R3146 two_stage_opamp_dummy_magic_29_0.VD4.n10 two_stage_opamp_dummy_magic_29_0.VD4.t5 11.2576
R3147 two_stage_opamp_dummy_magic_29_0.VD4.n10 two_stage_opamp_dummy_magic_29_0.VD4.t11 11.2576
R3148 two_stage_opamp_dummy_magic_29_0.VD4.n4 two_stage_opamp_dummy_magic_29_0.VD4.t3 11.2576
R3149 two_stage_opamp_dummy_magic_29_0.VD4.n4 two_stage_opamp_dummy_magic_29_0.VD4.t13 11.2576
R3150 two_stage_opamp_dummy_magic_29_0.VD4.n7 two_stage_opamp_dummy_magic_29_0.VD4.t9 11.2576
R3151 two_stage_opamp_dummy_magic_29_0.VD4.n7 two_stage_opamp_dummy_magic_29_0.VD4.t1 11.2576
R3152 two_stage_opamp_dummy_magic_29_0.VD4.n11 two_stage_opamp_dummy_magic_29_0.VD4.t15 11.2576
R3153 two_stage_opamp_dummy_magic_29_0.VD4.n11 two_stage_opamp_dummy_magic_29_0.VD4.t17 11.2576
R3154 two_stage_opamp_dummy_magic_29_0.VD4.n21 two_stage_opamp_dummy_magic_29_0.VD4.t26 11.2576
R3155 two_stage_opamp_dummy_magic_29_0.VD4.n21 two_stage_opamp_dummy_magic_29_0.VD4.t21 11.2576
R3156 two_stage_opamp_dummy_magic_29_0.VD4.n23 two_stage_opamp_dummy_magic_29_0.VD4.t24 11.2576
R3157 two_stage_opamp_dummy_magic_29_0.VD4.n23 two_stage_opamp_dummy_magic_29_0.VD4.t29 11.2576
R3158 two_stage_opamp_dummy_magic_29_0.VD4.n8 two_stage_opamp_dummy_magic_29_0.VD4.t25 11.2576
R3159 two_stage_opamp_dummy_magic_29_0.VD4.n8 two_stage_opamp_dummy_magic_29_0.VD4.t23 11.2576
R3160 two_stage_opamp_dummy_magic_29_0.VD4.n5 two_stage_opamp_dummy_magic_29_0.VD4.t27 11.2576
R3161 two_stage_opamp_dummy_magic_29_0.VD4.n5 two_stage_opamp_dummy_magic_29_0.VD4.t30 11.2576
R3162 two_stage_opamp_dummy_magic_29_0.VD4.n12 two_stage_opamp_dummy_magic_29_0.VD4.t20 11.2576
R3163 two_stage_opamp_dummy_magic_29_0.VD4.n12 two_stage_opamp_dummy_magic_29_0.VD4.t22 11.2576
R3164 two_stage_opamp_dummy_magic_29_0.VD4.n16 two_stage_opamp_dummy_magic_29_0.VD4.t7 11.2576
R3165 two_stage_opamp_dummy_magic_29_0.VD4.n16 two_stage_opamp_dummy_magic_29_0.VD4.t19 11.2576
R3166 two_stage_opamp_dummy_magic_29_0.VD4.n27 two_stage_opamp_dummy_magic_29_0.VD4.t28 11.2576
R3167 two_stage_opamp_dummy_magic_29_0.VD4.n27 two_stage_opamp_dummy_magic_29_0.VD4.t31 11.2576
R3168 two_stage_opamp_dummy_magic_29_0.VD4.n14 two_stage_opamp_dummy_magic_29_0.VD4.n13 5.66717
R3169 two_stage_opamp_dummy_magic_29_0.VD4.n25 two_stage_opamp_dummy_magic_29_0.VD4.n22 5.66717
R3170 two_stage_opamp_dummy_magic_29_0.VD4.n25 two_stage_opamp_dummy_magic_29_0.VD4.n24 5.29217
R3171 two_stage_opamp_dummy_magic_29_0.VD4.n28 two_stage_opamp_dummy_magic_29_0.VD4.n26 5.29217
R3172 two_stage_opamp_dummy_magic_29_0.VD4.n15 two_stage_opamp_dummy_magic_29_0.VD4.n9 5.29217
R3173 two_stage_opamp_dummy_magic_29_0.VD4.n14 two_stage_opamp_dummy_magic_29_0.VD4.n6 5.29217
R3174 two_stage_opamp_dummy_magic_29_0.VD4.n18 two_stage_opamp_dummy_magic_29_0.VD4.n17 1.90883
R3175 two_stage_opamp_dummy_magic_29_0.VD4.n20 two_stage_opamp_dummy_magic_29_0.VD4.n19 1.90883
R3176 two_stage_opamp_dummy_magic_29_0.VD4.n24 two_stage_opamp_dummy_magic_29_0.VD4.n0 1.02133
R3177 two_stage_opamp_dummy_magic_29_0.VD4.n0 two_stage_opamp_dummy_magic_29_0.VD4.n9 1.02133
R3178 two_stage_opamp_dummy_magic_29_0.VD4.n1 two_stage_opamp_dummy_magic_29_0.VD4.n6 1.02133
R3179 two_stage_opamp_dummy_magic_29_0.VD4.n13 two_stage_opamp_dummy_magic_29_0.VD4.n1 1.02133
R3180 two_stage_opamp_dummy_magic_29_0.VD4.n22 two_stage_opamp_dummy_magic_29_0.VD4.n3 1.02133
R3181 two_stage_opamp_dummy_magic_29_0.VD4.n0 two_stage_opamp_dummy_magic_29_0.VD4.n28 1.02133
R3182 two_stage_opamp_dummy_magic_29_0.VD4 two_stage_opamp_dummy_magic_29_0.VD4.n1 0.325242
R3183 two_stage_opamp_dummy_magic_29_0.VD4.n0 two_stage_opamp_dummy_magic_29_0.VD4.n2 0.0450006
R3184 two_stage_opamp_dummy_magic_29_0.VD4.n15 two_stage_opamp_dummy_magic_29_0.VD4.n14 0.3755
R3185 two_stage_opamp_dummy_magic_29_0.VD4.n26 two_stage_opamp_dummy_magic_29_0.VD4.n15 0.3755
R3186 two_stage_opamp_dummy_magic_29_0.VD4.n26 two_stage_opamp_dummy_magic_29_0.VD4.n25 0.3755
R3187 two_stage_opamp_dummy_magic_29_0.VD4.n3 two_stage_opamp_dummy_magic_29_0.VD4.n20 0.132669
R3188 two_stage_opamp_dummy_magic_29_0.VD4.n3 two_stage_opamp_dummy_magic_29_0.VD4.n2 0.0716452
R3189 two_stage_opamp_dummy_magic_29_0.VD4.n1 two_stage_opamp_dummy_magic_29_0.VD4.n0 0.107643
R3190 two_stage_opamp_dummy_magic_29_0.VD4 two_stage_opamp_dummy_magic_29_0.VD4.n2 0.251159
R3191 two_stage_opamp_dummy_magic_29_0.VD4.n17 two_stage_opamp_dummy_magic_29_0.VD4.n1 0.158238
R3192 two_stage_opamp_dummy_magic_29_0.X.n70 two_stage_opamp_dummy_magic_29_0.X.t43 1172.87
R3193 two_stage_opamp_dummy_magic_29_0.X.n66 two_stage_opamp_dummy_magic_29_0.X.t36 1172.87
R3194 two_stage_opamp_dummy_magic_29_0.X.n70 two_stage_opamp_dummy_magic_29_0.X.t29 996.134
R3195 two_stage_opamp_dummy_magic_29_0.X.n71 two_stage_opamp_dummy_magic_29_0.X.t45 996.134
R3196 two_stage_opamp_dummy_magic_29_0.X.n72 two_stage_opamp_dummy_magic_29_0.X.t28 996.134
R3197 two_stage_opamp_dummy_magic_29_0.X.n73 two_stage_opamp_dummy_magic_29_0.X.t44 996.134
R3198 two_stage_opamp_dummy_magic_29_0.X.n69 two_stage_opamp_dummy_magic_29_0.X.t30 996.134
R3199 two_stage_opamp_dummy_magic_29_0.X.n68 two_stage_opamp_dummy_magic_29_0.X.t46 996.134
R3200 two_stage_opamp_dummy_magic_29_0.X.n67 two_stage_opamp_dummy_magic_29_0.X.t32 996.134
R3201 two_stage_opamp_dummy_magic_29_0.X.n66 two_stage_opamp_dummy_magic_29_0.X.t49 996.134
R3202 two_stage_opamp_dummy_magic_29_0.X.n37 two_stage_opamp_dummy_magic_29_0.X.t31 690.867
R3203 two_stage_opamp_dummy_magic_29_0.X.n36 two_stage_opamp_dummy_magic_29_0.X.t26 690.867
R3204 two_stage_opamp_dummy_magic_29_0.X.n46 two_stage_opamp_dummy_magic_29_0.X.t33 530.201
R3205 two_stage_opamp_dummy_magic_29_0.X.n45 two_stage_opamp_dummy_magic_29_0.X.t27 530.201
R3206 two_stage_opamp_dummy_magic_29_0.X.n43 two_stage_opamp_dummy_magic_29_0.X.t54 514.134
R3207 two_stage_opamp_dummy_magic_29_0.X.n42 two_stage_opamp_dummy_magic_29_0.X.t39 514.134
R3208 two_stage_opamp_dummy_magic_29_0.X.n41 two_stage_opamp_dummy_magic_29_0.X.t52 514.134
R3209 two_stage_opamp_dummy_magic_29_0.X.n40 two_stage_opamp_dummy_magic_29_0.X.t34 514.134
R3210 two_stage_opamp_dummy_magic_29_0.X.n39 two_stage_opamp_dummy_magic_29_0.X.t47 514.134
R3211 two_stage_opamp_dummy_magic_29_0.X.n38 two_stage_opamp_dummy_magic_29_0.X.t35 514.134
R3212 two_stage_opamp_dummy_magic_29_0.X.n37 two_stage_opamp_dummy_magic_29_0.X.t48 514.134
R3213 two_stage_opamp_dummy_magic_29_0.X.n36 two_stage_opamp_dummy_magic_29_0.X.t41 514.134
R3214 two_stage_opamp_dummy_magic_29_0.X.n46 two_stage_opamp_dummy_magic_29_0.X.t51 353.467
R3215 two_stage_opamp_dummy_magic_29_0.X.n47 two_stage_opamp_dummy_magic_29_0.X.t38 353.467
R3216 two_stage_opamp_dummy_magic_29_0.X.n48 two_stage_opamp_dummy_magic_29_0.X.t50 353.467
R3217 two_stage_opamp_dummy_magic_29_0.X.n49 two_stage_opamp_dummy_magic_29_0.X.t37 353.467
R3218 two_stage_opamp_dummy_magic_29_0.X.n50 two_stage_opamp_dummy_magic_29_0.X.t53 353.467
R3219 two_stage_opamp_dummy_magic_29_0.X.n51 two_stage_opamp_dummy_magic_29_0.X.t40 353.467
R3220 two_stage_opamp_dummy_magic_29_0.X.n52 two_stage_opamp_dummy_magic_29_0.X.t25 353.467
R3221 two_stage_opamp_dummy_magic_29_0.X.n45 two_stage_opamp_dummy_magic_29_0.X.t42 353.467
R3222 two_stage_opamp_dummy_magic_29_0.X.n69 two_stage_opamp_dummy_magic_29_0.X.n68 176.733
R3223 two_stage_opamp_dummy_magic_29_0.X.n68 two_stage_opamp_dummy_magic_29_0.X.n67 176.733
R3224 two_stage_opamp_dummy_magic_29_0.X.n67 two_stage_opamp_dummy_magic_29_0.X.n66 176.733
R3225 two_stage_opamp_dummy_magic_29_0.X.n71 two_stage_opamp_dummy_magic_29_0.X.n70 176.733
R3226 two_stage_opamp_dummy_magic_29_0.X.n72 two_stage_opamp_dummy_magic_29_0.X.n71 176.733
R3227 two_stage_opamp_dummy_magic_29_0.X.n73 two_stage_opamp_dummy_magic_29_0.X.n72 176.733
R3228 two_stage_opamp_dummy_magic_29_0.X.n47 two_stage_opamp_dummy_magic_29_0.X.n46 176.733
R3229 two_stage_opamp_dummy_magic_29_0.X.n48 two_stage_opamp_dummy_magic_29_0.X.n47 176.733
R3230 two_stage_opamp_dummy_magic_29_0.X.n49 two_stage_opamp_dummy_magic_29_0.X.n48 176.733
R3231 two_stage_opamp_dummy_magic_29_0.X.n50 two_stage_opamp_dummy_magic_29_0.X.n49 176.733
R3232 two_stage_opamp_dummy_magic_29_0.X.n51 two_stage_opamp_dummy_magic_29_0.X.n50 176.733
R3233 two_stage_opamp_dummy_magic_29_0.X.n52 two_stage_opamp_dummy_magic_29_0.X.n51 176.733
R3234 two_stage_opamp_dummy_magic_29_0.X.n38 two_stage_opamp_dummy_magic_29_0.X.n37 176.733
R3235 two_stage_opamp_dummy_magic_29_0.X.n39 two_stage_opamp_dummy_magic_29_0.X.n38 176.733
R3236 two_stage_opamp_dummy_magic_29_0.X.n40 two_stage_opamp_dummy_magic_29_0.X.n39 176.733
R3237 two_stage_opamp_dummy_magic_29_0.X.n41 two_stage_opamp_dummy_magic_29_0.X.n40 176.733
R3238 two_stage_opamp_dummy_magic_29_0.X.n42 two_stage_opamp_dummy_magic_29_0.X.n41 176.733
R3239 two_stage_opamp_dummy_magic_29_0.X.n43 two_stage_opamp_dummy_magic_29_0.X.n42 176.733
R3240 two_stage_opamp_dummy_magic_29_0.X.n54 two_stage_opamp_dummy_magic_29_0.X.n53 165.472
R3241 two_stage_opamp_dummy_magic_29_0.X.n54 two_stage_opamp_dummy_magic_29_0.X.n44 165.472
R3242 two_stage_opamp_dummy_magic_29_0.X.n76 two_stage_opamp_dummy_magic_29_0.X.n75 152
R3243 two_stage_opamp_dummy_magic_29_0.X.n77 two_stage_opamp_dummy_magic_29_0.X.n76 131.571
R3244 two_stage_opamp_dummy_magic_29_0.X.n76 two_stage_opamp_dummy_magic_29_0.X.n74 124.517
R3245 two_stage_opamp_dummy_magic_29_0.X.n81 two_stage_opamp_dummy_magic_29_0.X.n54 74.5362
R3246 two_stage_opamp_dummy_magic_29_0.X.n13 two_stage_opamp_dummy_magic_29_0.X.n12 66.0338
R3247 two_stage_opamp_dummy_magic_29_0.X.n29 two_stage_opamp_dummy_magic_29_0.X.n28 66.0338
R3248 two_stage_opamp_dummy_magic_29_0.X.n26 two_stage_opamp_dummy_magic_29_0.X.n25 66.0338
R3249 two_stage_opamp_dummy_magic_29_0.X.n23 two_stage_opamp_dummy_magic_29_0.X.n22 66.0338
R3250 two_stage_opamp_dummy_magic_29_0.X.n19 two_stage_opamp_dummy_magic_29_0.X.n18 66.0338
R3251 two_stage_opamp_dummy_magic_29_0.X.n16 two_stage_opamp_dummy_magic_29_0.X.n15 66.0338
R3252 two_stage_opamp_dummy_magic_29_0.X.n110 two_stage_opamp_dummy_magic_29_0.X.n108 54.7984
R3253 two_stage_opamp_dummy_magic_29_0.X.n118 two_stage_opamp_dummy_magic_29_0.X.n117 54.4547
R3254 two_stage_opamp_dummy_magic_29_0.X.n116 two_stage_opamp_dummy_magic_29_0.X.n115 54.4547
R3255 two_stage_opamp_dummy_magic_29_0.X.n114 two_stage_opamp_dummy_magic_29_0.X.n113 54.4547
R3256 two_stage_opamp_dummy_magic_29_0.X.n112 two_stage_opamp_dummy_magic_29_0.X.n111 54.4547
R3257 two_stage_opamp_dummy_magic_29_0.X.n110 two_stage_opamp_dummy_magic_29_0.X.n109 54.4547
R3258 two_stage_opamp_dummy_magic_29_0.X.n60 two_stage_opamp_dummy_magic_29_0.X.t24 41.0384
R3259 two_stage_opamp_dummy_magic_29_0.X.n74 two_stage_opamp_dummy_magic_29_0.X.n69 40.1672
R3260 two_stage_opamp_dummy_magic_29_0.X.n74 two_stage_opamp_dummy_magic_29_0.X.n73 40.1672
R3261 two_stage_opamp_dummy_magic_29_0.X.n53 two_stage_opamp_dummy_magic_29_0.X.n45 40.1672
R3262 two_stage_opamp_dummy_magic_29_0.X.n53 two_stage_opamp_dummy_magic_29_0.X.n52 40.1672
R3263 two_stage_opamp_dummy_magic_29_0.X.n44 two_stage_opamp_dummy_magic_29_0.X.n36 40.1672
R3264 two_stage_opamp_dummy_magic_29_0.X.n44 two_stage_opamp_dummy_magic_29_0.X.n43 40.1672
R3265 two_stage_opamp_dummy_magic_29_0.X.n78 two_stage_opamp_dummy_magic_29_0.X.n77 16.3217
R3266 two_stage_opamp_dummy_magic_29_0.X.n117 two_stage_opamp_dummy_magic_29_0.X.t14 16.0005
R3267 two_stage_opamp_dummy_magic_29_0.X.n117 two_stage_opamp_dummy_magic_29_0.X.t17 16.0005
R3268 two_stage_opamp_dummy_magic_29_0.X.n115 two_stage_opamp_dummy_magic_29_0.X.t5 16.0005
R3269 two_stage_opamp_dummy_magic_29_0.X.n115 two_stage_opamp_dummy_magic_29_0.X.t3 16.0005
R3270 two_stage_opamp_dummy_magic_29_0.X.n113 two_stage_opamp_dummy_magic_29_0.X.t11 16.0005
R3271 two_stage_opamp_dummy_magic_29_0.X.n113 two_stage_opamp_dummy_magic_29_0.X.t4 16.0005
R3272 two_stage_opamp_dummy_magic_29_0.X.n111 two_stage_opamp_dummy_magic_29_0.X.t15 16.0005
R3273 two_stage_opamp_dummy_magic_29_0.X.n111 two_stage_opamp_dummy_magic_29_0.X.t9 16.0005
R3274 two_stage_opamp_dummy_magic_29_0.X.n109 two_stage_opamp_dummy_magic_29_0.X.t13 16.0005
R3275 two_stage_opamp_dummy_magic_29_0.X.n109 two_stage_opamp_dummy_magic_29_0.X.t10 16.0005
R3276 two_stage_opamp_dummy_magic_29_0.X.n108 two_stage_opamp_dummy_magic_29_0.X.t12 16.0005
R3277 two_stage_opamp_dummy_magic_29_0.X.n108 two_stage_opamp_dummy_magic_29_0.X.t22 16.0005
R3278 two_stage_opamp_dummy_magic_29_0.X.n75 two_stage_opamp_dummy_magic_29_0.X.n65 12.8005
R3279 two_stage_opamp_dummy_magic_29_0.X.n12 two_stage_opamp_dummy_magic_29_0.X.t16 11.2576
R3280 two_stage_opamp_dummy_magic_29_0.X.n12 two_stage_opamp_dummy_magic_29_0.X.t20 11.2576
R3281 two_stage_opamp_dummy_magic_29_0.X.n28 two_stage_opamp_dummy_magic_29_0.X.t8 11.2576
R3282 two_stage_opamp_dummy_magic_29_0.X.n28 two_stage_opamp_dummy_magic_29_0.X.t23 11.2576
R3283 two_stage_opamp_dummy_magic_29_0.X.n25 two_stage_opamp_dummy_magic_29_0.X.t21 11.2576
R3284 two_stage_opamp_dummy_magic_29_0.X.n25 two_stage_opamp_dummy_magic_29_0.X.t0 11.2576
R3285 two_stage_opamp_dummy_magic_29_0.X.n22 two_stage_opamp_dummy_magic_29_0.X.t6 11.2576
R3286 two_stage_opamp_dummy_magic_29_0.X.n22 two_stage_opamp_dummy_magic_29_0.X.t1 11.2576
R3287 two_stage_opamp_dummy_magic_29_0.X.n18 two_stage_opamp_dummy_magic_29_0.X.t7 11.2576
R3288 two_stage_opamp_dummy_magic_29_0.X.n18 two_stage_opamp_dummy_magic_29_0.X.t19 11.2576
R3289 two_stage_opamp_dummy_magic_29_0.X.n15 two_stage_opamp_dummy_magic_29_0.X.t18 11.2576
R3290 two_stage_opamp_dummy_magic_29_0.X.n15 two_stage_opamp_dummy_magic_29_0.X.t2 11.2576
R3291 two_stage_opamp_dummy_magic_29_0.X.n119 two_stage_opamp_dummy_magic_29_0.X.n118 11.1099
R3292 two_stage_opamp_dummy_magic_29_0.X.n75 two_stage_opamp_dummy_magic_29_0.X.n63 9.36264
R3293 two_stage_opamp_dummy_magic_29_0.X.n65 two_stage_opamp_dummy_magic_29_0.X.n64 9.3005
R3294 two_stage_opamp_dummy_magic_29_0.X.n103 two_stage_opamp_dummy_magic_29_0.X.n3 5.78175
R3295 two_stage_opamp_dummy_magic_29_0.X.n29 two_stage_opamp_dummy_magic_29_0.X.n27 5.66717
R3296 two_stage_opamp_dummy_magic_29_0.X.n14 two_stage_opamp_dummy_magic_29_0.X.n13 5.66717
R3297 two_stage_opamp_dummy_magic_29_0.X.n17 two_stage_opamp_dummy_magic_29_0.X.n13 5.66717
R3298 two_stage_opamp_dummy_magic_29_0.X.n120 two_stage_opamp_dummy_magic_29_0.X.n119 5.46373
R3299 two_stage_opamp_dummy_magic_29_0.X.n103 two_stage_opamp_dummy_magic_29_0.X.n102 5.438
R3300 two_stage_opamp_dummy_magic_29_0.X.n104 two_stage_opamp_dummy_magic_29_0.X.n2 5.438
R3301 two_stage_opamp_dummy_magic_29_0.X.n123 two_stage_opamp_dummy_magic_29_0.X.n105 5.438
R3302 two_stage_opamp_dummy_magic_29_0.X.n107 two_stage_opamp_dummy_magic_29_0.X.n106 5.438
R3303 two_stage_opamp_dummy_magic_29_0.X.n77 two_stage_opamp_dummy_magic_29_0.X.n65 5.33141
R3304 two_stage_opamp_dummy_magic_29_0.X.n30 two_stage_opamp_dummy_magic_29_0.X.n29 5.29217
R3305 two_stage_opamp_dummy_magic_29_0.X.n26 two_stage_opamp_dummy_magic_29_0.X.n10 5.29217
R3306 two_stage_opamp_dummy_magic_29_0.X.n27 two_stage_opamp_dummy_magic_29_0.X.n26 5.29217
R3307 two_stage_opamp_dummy_magic_29_0.X.n23 two_stage_opamp_dummy_magic_29_0.X.n21 5.29217
R3308 two_stage_opamp_dummy_magic_29_0.X.n24 two_stage_opamp_dummy_magic_29_0.X.n23 5.29217
R3309 two_stage_opamp_dummy_magic_29_0.X.n20 two_stage_opamp_dummy_magic_29_0.X.n19 5.29217
R3310 two_stage_opamp_dummy_magic_29_0.X.n19 two_stage_opamp_dummy_magic_29_0.X.n11 5.29217
R3311 two_stage_opamp_dummy_magic_29_0.X.n17 two_stage_opamp_dummy_magic_29_0.X.n16 5.29217
R3312 two_stage_opamp_dummy_magic_29_0.X.n16 two_stage_opamp_dummy_magic_29_0.X.n14 5.29217
R3313 two_stage_opamp_dummy_magic_29_0.X.n93 two_stage_opamp_dummy_magic_29_0.X.n9 4.5005
R3314 two_stage_opamp_dummy_magic_29_0.X.n93 two_stage_opamp_dummy_magic_29_0.X.n90 4.5005
R3315 two_stage_opamp_dummy_magic_29_0.X.n93 two_stage_opamp_dummy_magic_29_0.X.n88 4.5005
R3316 two_stage_opamp_dummy_magic_29_0.X.n93 two_stage_opamp_dummy_magic_29_0.X.n92 4.5005
R3317 two_stage_opamp_dummy_magic_29_0.X.n86 two_stage_opamp_dummy_magic_29_0.X.n31 4.5005
R3318 two_stage_opamp_dummy_magic_29_0.X.n80 two_stage_opamp_dummy_magic_29_0.X.n33 4.5005
R3319 two_stage_opamp_dummy_magic_29_0.X.n82 two_stage_opamp_dummy_magic_29_0.X.n81 4.5005
R3320 two_stage_opamp_dummy_magic_29_0.X.n81 two_stage_opamp_dummy_magic_29_0.X.n80 4.5005
R3321 two_stage_opamp_dummy_magic_29_0.X.n79 two_stage_opamp_dummy_magic_29_0.X.n78 4.5005
R3322 two_stage_opamp_dummy_magic_29_0.X.n57 two_stage_opamp_dummy_magic_29_0.X.n56 4.5005
R3323 two_stage_opamp_dummy_magic_29_0.X.n95 two_stage_opamp_dummy_magic_29_0.X.n30 2.35465
R3324 two_stage_opamp_dummy_magic_29_0.X.n59 two_stage_opamp_dummy_magic_29_0.X.n58 2.26187
R3325 two_stage_opamp_dummy_magic_29_0.X.n58 two_stage_opamp_dummy_magic_29_0.X.n55 2.26187
R3326 two_stage_opamp_dummy_magic_29_0.X.n95 two_stage_opamp_dummy_magic_29_0.X.n94 2.24654
R3327 two_stage_opamp_dummy_magic_29_0.X.n85 two_stage_opamp_dummy_magic_29_0.X.n6 2.24654
R3328 two_stage_opamp_dummy_magic_29_0.X.n89 two_stage_opamp_dummy_magic_29_0.X.n31 2.24063
R3329 two_stage_opamp_dummy_magic_29_0.X.n91 two_stage_opamp_dummy_magic_29_0.X.n31 2.24063
R3330 two_stage_opamp_dummy_magic_29_0.X.n93 two_stage_opamp_dummy_magic_29_0.X.n87 2.24063
R3331 two_stage_opamp_dummy_magic_29_0.X.n83 two_stage_opamp_dummy_magic_29_0.X.n82 2.24063
R3332 two_stage_opamp_dummy_magic_29_0.X.n35 two_stage_opamp_dummy_magic_29_0.X.n34 2.24063
R3333 two_stage_opamp_dummy_magic_29_0.X.n97 two_stage_opamp_dummy_magic_29_0.X.n96 2.24063
R3334 two_stage_opamp_dummy_magic_29_0.X.n97 two_stage_opamp_dummy_magic_29_0.X.n8 2.24063
R3335 two_stage_opamp_dummy_magic_29_0.X.n97 two_stage_opamp_dummy_magic_29_0.X.n7 2.24063
R3336 two_stage_opamp_dummy_magic_29_0.X.n84 two_stage_opamp_dummy_magic_29_0.X.n32 2.24063
R3337 two_stage_opamp_dummy_magic_29_0.X.n60 two_stage_opamp_dummy_magic_29_0.X.n59 2.24063
R3338 two_stage_opamp_dummy_magic_29_0.X.n62 two_stage_opamp_dummy_magic_29_0.X.n61 2.24063
R3339 two_stage_opamp_dummy_magic_29_0.X.n79 two_stage_opamp_dummy_magic_29_0.X.n63 2.22018
R3340 two_stage_opamp_dummy_magic_29_0.X.n79 two_stage_opamp_dummy_magic_29_0.X.n62 0.682792
R3341 two_stage_opamp_dummy_magic_29_0.X.n122 two_stage_opamp_dummy_magic_29_0.X.n121 0.643357
R3342 two_stage_opamp_dummy_magic_29_0.X.n123 two_stage_opamp_dummy_magic_29_0.X.n1 0.643357
R3343 two_stage_opamp_dummy_magic_29_0.X.n125 two_stage_opamp_dummy_magic_29_0.X.n124 0.643357
R3344 two_stage_opamp_dummy_magic_29_0.X.n2 two_stage_opamp_dummy_magic_29_0.X.n0 0.643357
R3345 two_stage_opamp_dummy_magic_29_0.X.n100 two_stage_opamp_dummy_magic_29_0.X.n5 0.643357
R3346 two_stage_opamp_dummy_magic_29_0.X.n102 two_stage_opamp_dummy_magic_29_0.X.n101 0.643357
R3347 two_stage_opamp_dummy_magic_29_0.X.n99 two_stage_opamp_dummy_magic_29_0.X.n4 0.643357
R3348 two_stage_opamp_dummy_magic_29_0.X.n98 two_stage_opamp_dummy_magic_29_0.X.n3 0.643357
R3349 two_stage_opamp_dummy_magic_29_0.X.n85 two_stage_opamp_dummy_magic_29_0.X.n84 0.479667
R3350 two_stage_opamp_dummy_magic_29_0.X.n80 two_stage_opamp_dummy_magic_29_0.X.n79 0.46925
R3351 two_stage_opamp_dummy_magic_29_0.X.n14 two_stage_opamp_dummy_magic_29_0.X.n11 0.3755
R3352 two_stage_opamp_dummy_magic_29_0.X.n24 two_stage_opamp_dummy_magic_29_0.X.n11 0.3755
R3353 two_stage_opamp_dummy_magic_29_0.X.n27 two_stage_opamp_dummy_magic_29_0.X.n24 0.3755
R3354 two_stage_opamp_dummy_magic_29_0.X.n20 two_stage_opamp_dummy_magic_29_0.X.n17 0.3755
R3355 two_stage_opamp_dummy_magic_29_0.X.n21 two_stage_opamp_dummy_magic_29_0.X.n20 0.3755
R3356 two_stage_opamp_dummy_magic_29_0.X.n21 two_stage_opamp_dummy_magic_29_0.X.n10 0.3755
R3357 two_stage_opamp_dummy_magic_29_0.X.n30 two_stage_opamp_dummy_magic_29_0.X.n10 0.3755
R3358 two_stage_opamp_dummy_magic_29_0.X.n112 two_stage_opamp_dummy_magic_29_0.X.n110 0.34425
R3359 two_stage_opamp_dummy_magic_29_0.X.n114 two_stage_opamp_dummy_magic_29_0.X.n112 0.34425
R3360 two_stage_opamp_dummy_magic_29_0.X.n116 two_stage_opamp_dummy_magic_29_0.X.n114 0.34425
R3361 two_stage_opamp_dummy_magic_29_0.X.n118 two_stage_opamp_dummy_magic_29_0.X.n116 0.34425
R3362 two_stage_opamp_dummy_magic_29_0.X.n104 two_stage_opamp_dummy_magic_29_0.X.n103 0.34425
R3363 two_stage_opamp_dummy_magic_29_0.X.n105 two_stage_opamp_dummy_magic_29_0.X.n104 0.34425
R3364 two_stage_opamp_dummy_magic_29_0.X.n107 two_stage_opamp_dummy_magic_29_0.X.n105 0.34425
R3365 two_stage_opamp_dummy_magic_29_0.X.n119 two_stage_opamp_dummy_magic_29_0.X.n107 0.34425
R3366 two_stage_opamp_dummy_magic_29_0.X.n98 two_stage_opamp_dummy_magic_29_0.X.n97 0.270589
R3367 two_stage_opamp_dummy_magic_29_0.X.n121 two_stage_opamp_dummy_magic_29_0.X.n120 0.242602
R3368 two_stage_opamp_dummy_magic_29_0.X.n78 two_stage_opamp_dummy_magic_29_0.X.n64 0.1255
R3369 two_stage_opamp_dummy_magic_29_0.X.n64 two_stage_opamp_dummy_magic_29_0.X.n63 0.0626438
R3370 two_stage_opamp_dummy_magic_29_0.X.n82 two_stage_opamp_dummy_magic_29_0.X.n34 0.0421667
R3371 two_stage_opamp_dummy_magic_29_0.X.n4 two_stage_opamp_dummy_magic_29_0.X.n3 0.0250536
R3372 two_stage_opamp_dummy_magic_29_0.X.n102 two_stage_opamp_dummy_magic_29_0.X.n4 0.0250536
R3373 two_stage_opamp_dummy_magic_29_0.X.n102 two_stage_opamp_dummy_magic_29_0.X.n5 0.0250536
R3374 two_stage_opamp_dummy_magic_29_0.X.n5 two_stage_opamp_dummy_magic_29_0.X.n2 0.0250536
R3375 two_stage_opamp_dummy_magic_29_0.X.n124 two_stage_opamp_dummy_magic_29_0.X.n2 0.0250536
R3376 two_stage_opamp_dummy_magic_29_0.X.n124 two_stage_opamp_dummy_magic_29_0.X.n123 0.0250536
R3377 two_stage_opamp_dummy_magic_29_0.X.n123 two_stage_opamp_dummy_magic_29_0.X.n122 0.0250536
R3378 two_stage_opamp_dummy_magic_29_0.X.n122 two_stage_opamp_dummy_magic_29_0.X.n106 0.0250536
R3379 two_stage_opamp_dummy_magic_29_0.X.n99 two_stage_opamp_dummy_magic_29_0.X.n98 0.0250536
R3380 two_stage_opamp_dummy_magic_29_0.X.n101 two_stage_opamp_dummy_magic_29_0.X.n99 0.0250536
R3381 two_stage_opamp_dummy_magic_29_0.X.n101 two_stage_opamp_dummy_magic_29_0.X.n100 0.0250536
R3382 two_stage_opamp_dummy_magic_29_0.X.n100 two_stage_opamp_dummy_magic_29_0.X.n0 0.0250536
R3383 two_stage_opamp_dummy_magic_29_0.X.n125 two_stage_opamp_dummy_magic_29_0.X.n1 0.0250536
R3384 two_stage_opamp_dummy_magic_29_0.X.n121 two_stage_opamp_dummy_magic_29_0.X.n1 0.0250536
R3385 two_stage_opamp_dummy_magic_29_0.X.n120 two_stage_opamp_dummy_magic_29_0.X.n106 0.0241021
R3386 two_stage_opamp_dummy_magic_29_0.X.n90 two_stage_opamp_dummy_magic_29_0.X.n89 0.0217373
R3387 two_stage_opamp_dummy_magic_29_0.X.n92 two_stage_opamp_dummy_magic_29_0.X.n91 0.0217373
R3388 two_stage_opamp_dummy_magic_29_0.X.n87 two_stage_opamp_dummy_magic_29_0.X.n86 0.0217373
R3389 two_stage_opamp_dummy_magic_29_0.X.n84 two_stage_opamp_dummy_magic_29_0.X.n83 0.0217373
R3390 two_stage_opamp_dummy_magic_29_0.X.n81 two_stage_opamp_dummy_magic_29_0.X.n35 0.0217373
R3391 two_stage_opamp_dummy_magic_29_0.X.n89 two_stage_opamp_dummy_magic_29_0.X.n9 0.0217373
R3392 two_stage_opamp_dummy_magic_29_0.X.n91 two_stage_opamp_dummy_magic_29_0.X.n88 0.0217373
R3393 two_stage_opamp_dummy_magic_29_0.X.n87 two_stage_opamp_dummy_magic_29_0.X.n85 0.0217373
R3394 two_stage_opamp_dummy_magic_29_0.X.n62 two_stage_opamp_dummy_magic_29_0.X.n55 0.0217373
R3395 two_stage_opamp_dummy_magic_29_0.X.n83 two_stage_opamp_dummy_magic_29_0.X.n33 0.0217373
R3396 two_stage_opamp_dummy_magic_29_0.X.n35 two_stage_opamp_dummy_magic_29_0.X.n33 0.0217373
R3397 two_stage_opamp_dummy_magic_29_0.X.n58 two_stage_opamp_dummy_magic_29_0.X.n56 0.0217373
R3398 two_stage_opamp_dummy_magic_29_0.X.n57 two_stage_opamp_dummy_magic_29_0.X.n55 0.0217373
R3399 two_stage_opamp_dummy_magic_29_0.X.n96 two_stage_opamp_dummy_magic_29_0.X.n9 0.0217373
R3400 two_stage_opamp_dummy_magic_29_0.X.n88 two_stage_opamp_dummy_magic_29_0.X.n8 0.0217373
R3401 two_stage_opamp_dummy_magic_29_0.X.n86 two_stage_opamp_dummy_magic_29_0.X.n7 0.0217373
R3402 two_stage_opamp_dummy_magic_29_0.X.n96 two_stage_opamp_dummy_magic_29_0.X.n95 0.0217373
R3403 two_stage_opamp_dummy_magic_29_0.X.n90 two_stage_opamp_dummy_magic_29_0.X.n8 0.0217373
R3404 two_stage_opamp_dummy_magic_29_0.X.n92 two_stage_opamp_dummy_magic_29_0.X.n7 0.0217373
R3405 two_stage_opamp_dummy_magic_29_0.X.n59 two_stage_opamp_dummy_magic_29_0.X.n57 0.0217373
R3406 two_stage_opamp_dummy_magic_29_0.X.n80 two_stage_opamp_dummy_magic_29_0.X.n32 0.0217373
R3407 two_stage_opamp_dummy_magic_29_0.X.n34 two_stage_opamp_dummy_magic_29_0.X.n32 0.0217373
R3408 two_stage_opamp_dummy_magic_29_0.X.n61 two_stage_opamp_dummy_magic_29_0.X.n56 0.0217373
R3409 two_stage_opamp_dummy_magic_29_0.X.n61 two_stage_opamp_dummy_magic_29_0.X.n60 0.0217373
R3410 two_stage_opamp_dummy_magic_29_0.X two_stage_opamp_dummy_magic_29_0.X.n125 0.016125
R3411 two_stage_opamp_dummy_magic_29_0.X.n94 two_stage_opamp_dummy_magic_29_0.X.n31 0.00991089
R3412 two_stage_opamp_dummy_magic_29_0.X.n97 two_stage_opamp_dummy_magic_29_0.X.n6 0.00991089
R3413 two_stage_opamp_dummy_magic_29_0.X.n94 two_stage_opamp_dummy_magic_29_0.X.n93 0.00991089
R3414 two_stage_opamp_dummy_magic_29_0.X.n31 two_stage_opamp_dummy_magic_29_0.X.n6 0.00991089
R3415 two_stage_opamp_dummy_magic_29_0.X two_stage_opamp_dummy_magic_29_0.X.n0 0.00942857
R3416 GNDA.n4916 GNDA.n429 497659
R3417 GNDA.n1663 GNDA.n635 396244
R3418 GNDA.n4916 GNDA.n430 313500
R3419 GNDA.n4065 GNDA.n633 195549
R3420 GNDA.n4123 GNDA.n430 182270
R3421 GNDA.n4917 GNDA.n428 173869
R3422 GNDA.n4122 GNDA.n4121 158989
R3423 GNDA.n1666 GNDA.n635 148345
R3424 GNDA.n4122 GNDA.n599 145383
R3425 GNDA.n635 GNDA.n599 134933
R3426 GNDA.n3382 GNDA.n633 132035
R3427 GNDA.n4916 GNDA.n4915 132035
R3428 GNDA.n1664 GNDA.n1663 105027
R3429 GNDA.n1669 GNDA.n1663 71214.8
R3430 GNDA.n4917 GNDA.n429 62388
R3431 GNDA.t92 GNDA.n635 55812.1
R3432 GNDA.n4126 GNDA.n4122 42457
R3433 GNDA.t18 GNDA.n4916 28032.8
R3434 GNDA.t13 GNDA.n633 28031.1
R3435 GNDA.n4065 GNDA.n4064 23839.1
R3436 GNDA.n4062 GNDA.n599 21706.7
R3437 GNDA.n4126 GNDA.n4125 18170.4
R3438 GNDA.n4931 GNDA.n4930 17109.1
R3439 GNDA.n4062 GNDA.n4061 16116.7
R3440 GNDA.n4063 GNDA.n4062 13566.7
R3441 GNDA.n1667 GNDA.n1666 13527.3
R3442 GNDA.n1668 GNDA.n1667 13460.8
R3443 GNDA.n4064 GNDA.n634 13200
R3444 GNDA.n4062 GNDA.n636 13111.6
R3445 GNDA.n1666 GNDA.n428 12640.3
R3446 GNDA.n4125 GNDA.n4124 11163
R3447 GNDA.n742 GNDA.n637 11032
R3448 GNDA.n742 GNDA.n600 11032
R3449 GNDA.n728 GNDA.n637 10933.5
R3450 GNDA.n728 GNDA.n600 10933.5
R3451 GNDA.n689 GNDA.n602 10884.2
R3452 GNDA.n4120 GNDA.n602 10884.2
R3453 GNDA.n689 GNDA.n601 10441
R3454 GNDA.n4120 GNDA.n601 10441
R3455 GNDA.n4064 GNDA.n4063 10046.7
R3456 GNDA.n4059 GNDA.n746 9850
R3457 GNDA.n4045 GNDA.n746 9751.5
R3458 GNDA.n1670 GNDA.n1669 9511.11
R3459 GNDA.n1670 GNDA.n428 9423.88
R3460 GNDA.n4059 GNDA.n745 9406.75
R3461 GNDA.n4045 GNDA.n745 9308.25
R3462 GNDA.n4067 GNDA.n4066 7301.54
R3463 GNDA.n2534 GNDA.n2532 7286.54
R3464 GNDA.n4123 GNDA.n429 6794.03
R3465 GNDA.n4124 GNDA.n4123 6475.77
R3466 GNDA.n3999 GNDA.n3997 5910
R3467 GNDA.n4125 GNDA.n430 5681.89
R3468 GNDA.n3998 GNDA.n3997 5466.75
R3469 GNDA.n4004 GNDA.n3999 5319
R3470 GNDA.n4004 GNDA.n3998 4875.75
R3471 GNDA.n1665 GNDA.n1664 4738.46
R3472 GNDA.n727 GNDA.n726 4375.56
R3473 GNDA.t186 GNDA.n1670 4106.67
R3474 GNDA.n1669 GNDA.n1668 4106.67
R3475 GNDA.n676 GNDA.n672 3841.5
R3476 GNDA.n676 GNDA.n673 3841.5
R3477 GNDA.n723 GNDA.n672 3743
R3478 GNDA.n723 GNDA.n673 3743
R3479 GNDA.n1665 GNDA.n635 3156.91
R3480 GNDA.n4063 GNDA.n635 3156.91
R3481 GNDA.n1456 GNDA.n1455 1684.55
R3482 GNDA.n744 GNDA.n743 1417.78
R3483 GNDA.n676 GNDA.t63 1319.17
R3484 GNDA.t3 GNDA.n636 1161.11
R3485 GNDA.n744 GNDA.t3 1148.89
R3486 GNDA.n725 GNDA.n724 1100
R3487 GNDA.n724 GNDA.n671 1075.56
R3488 GNDA.n743 GNDA.t0 1075.56
R3489 GNDA.n760 GNDA.n759 1075.56
R3490 GNDA.n1668 GNDA.n1664 1031.25
R3491 GNDA.n727 GNDA.t0 1026.67
R3492 GNDA.n726 GNDA.t46 1002.22
R3493 GNDA.n4066 GNDA.n4065 915.982
R3494 GNDA.n4005 GNDA.t43 855.557
R3495 GNDA.n3999 GNDA.t43 854.722
R3496 GNDA.n1667 GNDA.n1665 854.477
R3497 GNDA.t46 GNDA.n725 782.222
R3498 GNDA.t47 GNDA.n760 782.222
R3499 GNDA.n3380 GNDA.t207 749.742
R3500 GNDA.n4913 GNDA.t244 749.742
R3501 GNDA.n4127 GNDA.t225 749.742
R3502 GNDA.n4069 GNDA.t214 747.734
R3503 GNDA.t186 GNDA.n102 741.376
R3504 GNDA.n2520 GNDA.n2519 686.717
R3505 GNDA.n2065 GNDA.n2064 686.717
R3506 GNDA.n2057 GNDA.n1882 686.717
R3507 GNDA.n2511 GNDA.n1560 686.717
R3508 GNDA.n730 GNDA.n729 678.4
R3509 GNDA.n729 GNDA.n670 678.4
R3510 GNDA.n688 GNDA.n687 675.201
R3511 GNDA.n687 GNDA.n604 675.201
R3512 GNDA.n2325 GNDA.t84 671.187
R3513 GNDA.n2043 GNDA.n2042 669.307
R3514 GNDA.n1928 GNDA.n1927 669.307
R3515 GNDA.n4017 GNDA.t238 659.367
R3516 GNDA.n4016 GNDA.t259 659.367
R3517 GNDA.n707 GNDA.t219 659.367
R3518 GNDA.n679 GNDA.t198 659.367
R3519 GNDA.n4972 GNDA.n357 654.447
R3520 GNDA.n686 GNDA.n603 646.4
R3521 GNDA.n691 GNDA.n686 646.4
R3522 GNDA.n4058 GNDA.n747 611.201
R3523 GNDA.n4046 GNDA.n747 604.801
R3524 GNDA.n1425 GNDA.n1424 585.003
R3525 GNDA.n1863 GNDA.n1862 585.001
R3526 GNDA.n1866 GNDA.n1865 585.001
R3527 GNDA.n1914 GNDA.n1913 585.001
R3528 GNDA.n1916 GNDA.n1915 585.001
R3529 GNDA.n1660 GNDA.n1659 585.001
R3530 GNDA.n2473 GNDA.n2472 585.001
R3531 GNDA.n2546 GNDA.n2545 585.001
R3532 GNDA.n4987 GNDA.n4986 585
R3533 GNDA.n4988 GNDA.n4987 585
R3534 GNDA.n299 GNDA.n298 585
R3535 GNDA.n4989 GNDA.n299 585
R3536 GNDA.n4992 GNDA.n4991 585
R3537 GNDA.n4991 GNDA.n4990 585
R3538 GNDA.n4993 GNDA.n297 585
R3539 GNDA.n297 GNDA.n296 585
R3540 GNDA.n4995 GNDA.n4994 585
R3541 GNDA.n4996 GNDA.n4995 585
R3542 GNDA.n295 GNDA.n294 585
R3543 GNDA.n4997 GNDA.n295 585
R3544 GNDA.n5000 GNDA.n4999 585
R3545 GNDA.n4999 GNDA.n4998 585
R3546 GNDA.n5001 GNDA.n293 585
R3547 GNDA.n293 GNDA.n292 585
R3548 GNDA.n5003 GNDA.n5002 585
R3549 GNDA.n5004 GNDA.n5003 585
R3550 GNDA.n291 GNDA.n290 585
R3551 GNDA.n5005 GNDA.n291 585
R3552 GNDA.n5008 GNDA.n5007 585
R3553 GNDA.n5007 GNDA.n5006 585
R3554 GNDA.n5009 GNDA.n289 585
R3555 GNDA.n289 GNDA.n99 585
R3556 GNDA.n4971 GNDA.n4970 585
R3557 GNDA.n4969 GNDA.n355 585
R3558 GNDA.t186 GNDA.n355 585
R3559 GNDA.n5368 GNDA.n5367 585
R3560 GNDA.n131 GNDA.n129 585
R3561 GNDA.n242 GNDA.n241 585
R3562 GNDA.n244 GNDA.n243 585
R3563 GNDA.n246 GNDA.n245 585
R3564 GNDA.n248 GNDA.n247 585
R3565 GNDA.n250 GNDA.n249 585
R3566 GNDA.n252 GNDA.n251 585
R3567 GNDA.n254 GNDA.n253 585
R3568 GNDA.n256 GNDA.n255 585
R3569 GNDA.n258 GNDA.n257 585
R3570 GNDA.n260 GNDA.n259 585
R3571 GNDA.n2174 GNDA.n2173 585
R3572 GNDA.n2171 GNDA.n2170 585
R3573 GNDA.n2169 GNDA.n2168 585
R3574 GNDA.n2167 GNDA.n2166 585
R3575 GNDA.n2165 GNDA.n2164 585
R3576 GNDA.n2163 GNDA.n2162 585
R3577 GNDA.n2161 GNDA.n2160 585
R3578 GNDA.n2159 GNDA.n2158 585
R3579 GNDA.n2157 GNDA.n2156 585
R3580 GNDA.n2155 GNDA.n2154 585
R3581 GNDA.n2153 GNDA.n2152 585
R3582 GNDA.n135 GNDA.n132 585
R3583 GNDA.n2328 GNDA.n2327 585
R3584 GNDA.n2330 GNDA.n2329 585
R3585 GNDA.n2332 GNDA.n2331 585
R3586 GNDA.n2334 GNDA.n2333 585
R3587 GNDA.n2336 GNDA.n2335 585
R3588 GNDA.n2338 GNDA.n2337 585
R3589 GNDA.n2340 GNDA.n2339 585
R3590 GNDA.n2342 GNDA.n2341 585
R3591 GNDA.n2344 GNDA.n2343 585
R3592 GNDA.n2346 GNDA.n2345 585
R3593 GNDA.n2348 GNDA.n2347 585
R3594 GNDA.n2350 GNDA.n2349 585
R3595 GNDA.n5548 GNDA.n5547 585
R3596 GNDA.n5545 GNDA.n54 585
R3597 GNDA.n59 GNDA.n58 585
R3598 GNDA.n5540 GNDA.n5539 585
R3599 GNDA.n5538 GNDA.n5537 585
R3600 GNDA.n5464 GNDA.n63 585
R3601 GNDA.n5466 GNDA.n5465 585
R3602 GNDA.n5471 GNDA.n5470 585
R3603 GNDA.n5469 GNDA.n5462 585
R3604 GNDA.n5477 GNDA.n5476 585
R3605 GNDA.n5479 GNDA.n5478 585
R3606 GNDA.n5460 GNDA.n5459 585
R3607 GNDA.n5125 GNDA.n5124 585
R3608 GNDA.n5122 GNDA.n5121 585
R3609 GNDA.n5120 GNDA.n5119 585
R3610 GNDA.n5036 GNDA.n5012 585
R3611 GNDA.n5038 GNDA.n5037 585
R3612 GNDA.n5042 GNDA.n5041 585
R3613 GNDA.n5044 GNDA.n5043 585
R3614 GNDA.n5051 GNDA.n5050 585
R3615 GNDA.n5049 GNDA.n5034 585
R3616 GNDA.n5057 GNDA.n5056 585
R3617 GNDA.n5059 GNDA.n5058 585
R3618 GNDA.n5032 GNDA.n5031 585
R3619 GNDA.n328 GNDA.n325 585
R3620 GNDA.n329 GNDA.n323 585
R3621 GNDA.n330 GNDA.n322 585
R3622 GNDA.n320 GNDA.n318 585
R3623 GNDA.n336 GNDA.n317 585
R3624 GNDA.n337 GNDA.n315 585
R3625 GNDA.n338 GNDA.n314 585
R3626 GNDA.n312 GNDA.n310 585
R3627 GNDA.n344 GNDA.n309 585
R3628 GNDA.n345 GNDA.n307 585
R3629 GNDA.n346 GNDA.n306 585
R3630 GNDA.n302 GNDA.n301 585
R3631 GNDA.n133 GNDA.n85 585
R3632 GNDA.n5457 GNDA.n85 585
R3633 GNDA.n349 GNDA.n302 585
R3634 GNDA.n347 GNDA.n346 585
R3635 GNDA.n345 GNDA.n304 585
R3636 GNDA.n344 GNDA.n343 585
R3637 GNDA.n341 GNDA.n310 585
R3638 GNDA.n339 GNDA.n338 585
R3639 GNDA.n337 GNDA.n311 585
R3640 GNDA.n336 GNDA.n335 585
R3641 GNDA.n333 GNDA.n318 585
R3642 GNDA.n331 GNDA.n330 585
R3643 GNDA.n329 GNDA.n319 585
R3644 GNDA.n328 GNDA.n327 585
R3645 GNDA.n133 GNDA.n55 585
R3646 GNDA.n5457 GNDA.n55 585
R3647 GNDA.n5343 GNDA.n159 585
R3648 GNDA.n5344 GNDA.n150 585
R3649 GNDA.n5347 GNDA.n149 585
R3650 GNDA.n5348 GNDA.n148 585
R3651 GNDA.n5351 GNDA.n147 585
R3652 GNDA.n5352 GNDA.n146 585
R3653 GNDA.n5355 GNDA.n145 585
R3654 GNDA.n5357 GNDA.n144 585
R3655 GNDA.n5358 GNDA.n143 585
R3656 GNDA.n5359 GNDA.n142 585
R3657 GNDA.n151 GNDA.n134 585
R3658 GNDA.n5365 GNDA.n130 585
R3659 GNDA.n5365 GNDA.n5364 585
R3660 GNDA.n136 GNDA.n134 585
R3661 GNDA.n5360 GNDA.n5359 585
R3662 GNDA.n5358 GNDA.n141 585
R3663 GNDA.n5357 GNDA.n5356 585
R3664 GNDA.n5355 GNDA.n5354 585
R3665 GNDA.n5353 GNDA.n5352 585
R3666 GNDA.n5351 GNDA.n5350 585
R3667 GNDA.n5349 GNDA.n5348 585
R3668 GNDA.n5347 GNDA.n5346 585
R3669 GNDA.n5345 GNDA.n5344 585
R3670 GNDA.n5343 GNDA.n5342 585
R3671 GNDA.n2089 GNDA.n1713 585
R3672 GNDA.n2090 GNDA.n1711 585
R3673 GNDA.n1710 GNDA.n1707 585
R3674 GNDA.n2096 GNDA.n1706 585
R3675 GNDA.n2097 GNDA.n1705 585
R3676 GNDA.n2098 GNDA.n1703 585
R3677 GNDA.n1702 GNDA.n1699 585
R3678 GNDA.n2103 GNDA.n1698 585
R3679 GNDA.n2104 GNDA.n1697 585
R3680 GNDA.n1695 GNDA.n1693 585
R3681 GNDA.n2108 GNDA.n1692 585
R3682 GNDA.n2109 GNDA.n1690 585
R3683 GNDA.n2110 GNDA.n2109 585
R3684 GNDA.n2108 GNDA.n2107 585
R3685 GNDA.n2106 GNDA.n1693 585
R3686 GNDA.n2106 GNDA.n1662 585
R3687 GNDA.n2105 GNDA.n2104 585
R3688 GNDA.n2103 GNDA.n2102 585
R3689 GNDA.n2101 GNDA.n1699 585
R3690 GNDA.n2099 GNDA.n2098 585
R3691 GNDA.n2097 GNDA.n1700 585
R3692 GNDA.n2096 GNDA.n2095 585
R3693 GNDA.n2093 GNDA.n1707 585
R3694 GNDA.n2091 GNDA.n2090 585
R3695 GNDA.n2089 GNDA.n1708 585
R3696 GNDA.n1708 GNDA.n1662 585
R3697 GNDA.n1812 GNDA.n1811 585
R3698 GNDA.n1813 GNDA.n1809 585
R3699 GNDA.n1815 GNDA.n1814 585
R3700 GNDA.n1817 GNDA.n1807 585
R3701 GNDA.n1819 GNDA.n1818 585
R3702 GNDA.n1820 GNDA.n1806 585
R3703 GNDA.n1822 GNDA.n1821 585
R3704 GNDA.n1824 GNDA.n1804 585
R3705 GNDA.n1826 GNDA.n1825 585
R3706 GNDA.n1827 GNDA.n1803 585
R3707 GNDA.n1829 GNDA.n1828 585
R3708 GNDA.n1831 GNDA.n1802 585
R3709 GNDA.n2135 GNDA.n2134 585
R3710 GNDA.n2131 GNDA.n1682 585
R3711 GNDA.n2130 GNDA.n2129 585
R3712 GNDA.n2128 GNDA.n2127 585
R3713 GNDA.n2126 GNDA.n1684 585
R3714 GNDA.n2124 GNDA.n2123 585
R3715 GNDA.n2122 GNDA.n1685 585
R3716 GNDA.n2121 GNDA.n2120 585
R3717 GNDA.n2118 GNDA.n1686 585
R3718 GNDA.n2116 GNDA.n2115 585
R3719 GNDA.n2114 GNDA.n1687 585
R3720 GNDA.n2113 GNDA.n2112 585
R3721 GNDA.n2422 GNDA.n2421 585
R3722 GNDA.n2423 GNDA.n2395 585
R3723 GNDA.n2425 GNDA.n2424 585
R3724 GNDA.n2427 GNDA.n2393 585
R3725 GNDA.n2429 GNDA.n2428 585
R3726 GNDA.n2430 GNDA.n2392 585
R3727 GNDA.n2432 GNDA.n2431 585
R3728 GNDA.n2434 GNDA.n2390 585
R3729 GNDA.n2436 GNDA.n2435 585
R3730 GNDA.n2437 GNDA.n2389 585
R3731 GNDA.n2439 GNDA.n2438 585
R3732 GNDA.n2441 GNDA.n2388 585
R3733 GNDA.n5179 GNDA.n162 585
R3734 GNDA.n5179 GNDA.n161 585
R3735 GNDA.n5269 GNDA.n5268 585
R3736 GNDA.n5266 GNDA.n226 585
R3737 GNDA.n5156 GNDA.n5155 585
R3738 GNDA.n5261 GNDA.n5260 585
R3739 GNDA.n5259 GNDA.n5258 585
R3740 GNDA.n5185 GNDA.n5160 585
R3741 GNDA.n5187 GNDA.n5186 585
R3742 GNDA.n5192 GNDA.n5191 585
R3743 GNDA.n5190 GNDA.n5183 585
R3744 GNDA.n5198 GNDA.n5197 585
R3745 GNDA.n5200 GNDA.n5199 585
R3746 GNDA.n5181 GNDA.n5180 585
R3747 GNDA.n5341 GNDA.n162 585
R3748 GNDA.n5341 GNDA.n161 585
R3749 GNDA.n5340 GNDA.n5339 585
R3750 GNDA.n5337 GNDA.n5336 585
R3751 GNDA.n5335 GNDA.n5334 585
R3752 GNDA.n199 GNDA.n167 585
R3753 GNDA.n219 GNDA.n218 585
R3754 GNDA.n215 GNDA.n198 585
R3755 GNDA.n202 GNDA.n201 585
R3756 GNDA.n210 GNDA.n209 585
R3757 GNDA.n208 GNDA.n207 585
R3758 GNDA.n188 GNDA.n187 585
R3759 GNDA.n5274 GNDA.n5273 585
R3760 GNDA.n2136 GNDA.n189 585
R3761 GNDA.n2263 GNDA.n2139 585
R3762 GNDA.n2287 GNDA.n2265 585
R3763 GNDA.n2289 GNDA.n2288 585
R3764 GNDA.n2285 GNDA.n2284 585
R3765 GNDA.n2283 GNDA.n2282 585
R3766 GNDA.n2278 GNDA.n2277 585
R3767 GNDA.n2276 GNDA.n2275 585
R3768 GNDA.n2271 GNDA.n2270 585
R3769 GNDA.n2269 GNDA.n2190 585
R3770 GNDA.n2297 GNDA.n2296 585
R3771 GNDA.n2299 GNDA.n2298 585
R3772 GNDA.n2302 GNDA.n2301 585
R3773 GNDA.n2531 GNDA.n2530 585
R3774 GNDA.n2532 GNDA.n2531 585
R3775 GNDA.n2528 GNDA.n1457 585
R3776 GNDA.n1457 GNDA.n1456 585
R3777 GNDA.n2535 GNDA.n1453 585
R3778 GNDA.n2538 GNDA.n2537 585
R3779 GNDA.n2537 GNDA.n2536 585
R3780 GNDA.n1452 GNDA.n1451 585
R3781 GNDA.n1454 GNDA.n1452 585
R3782 GNDA.n2405 GNDA.n2404 585
R3783 GNDA.n2407 GNDA.n2404 585
R3784 GNDA.n2409 GNDA.n2406 585
R3785 GNDA.n2409 GNDA.n2408 585
R3786 GNDA.n2410 GNDA.n2403 585
R3787 GNDA.n2410 GNDA.n1562 585
R3788 GNDA.n2412 GNDA.n2411 585
R3789 GNDA.n2411 GNDA.n1561 585
R3790 GNDA.n2413 GNDA.n2401 585
R3791 GNDA.n2401 GNDA.n2400 585
R3792 GNDA.n2415 GNDA.n2414 585
R3793 GNDA.n2416 GNDA.n2415 585
R3794 GNDA.n2402 GNDA.n2398 585
R3795 GNDA.n2417 GNDA.n2398 585
R3796 GNDA.n2419 GNDA.n2399 585
R3797 GNDA.n2419 GNDA.n2418 585
R3798 GNDA.n2420 GNDA.n2396 585
R3799 GNDA.n2420 GNDA.n102 585
R3800 GNDA.n2534 GNDA.n2533 585
R3801 GNDA.n2187 GNDA.n2186 585
R3802 GNDA.n2307 GNDA.n2306 585
R3803 GNDA.n2308 GNDA.n2307 585
R3804 GNDA.n2184 GNDA.n2183 585
R3805 GNDA.n2309 GNDA.n2184 585
R3806 GNDA.n2312 GNDA.n2311 585
R3807 GNDA.n2311 GNDA.n2310 585
R3808 GNDA.n2313 GNDA.n2182 585
R3809 GNDA.n2185 GNDA.n2182 585
R3810 GNDA.n2315 GNDA.n2314 585
R3811 GNDA.n2315 GNDA.n108 585
R3812 GNDA.n2316 GNDA.n2181 585
R3813 GNDA.n2316 GNDA.n109 585
R3814 GNDA.n2319 GNDA.n2318 585
R3815 GNDA.n2318 GNDA.n2317 585
R3816 GNDA.n2320 GNDA.n2179 585
R3817 GNDA.n2179 GNDA.n2178 585
R3818 GNDA.n2322 GNDA.n2321 585
R3819 GNDA.n2323 GNDA.n2322 585
R3820 GNDA.n2180 GNDA.n2177 585
R3821 GNDA.n2324 GNDA.n2177 585
R3822 GNDA.n2326 GNDA.n2176 585
R3823 GNDA.n2326 GNDA.n2325 585
R3824 GNDA.n2303 GNDA.n103 585
R3825 GNDA.n5382 GNDA.n5381 585
R3826 GNDA.n5384 GNDA.n88 585
R3827 GNDA.n5455 GNDA.n5454 585
R3828 GNDA.n24 GNDA.n22 585
R3829 GNDA.n5553 GNDA.n5552 585
R3830 GNDA.n32 GNDA.n25 585
R3831 GNDA.n40 GNDA.n39 585
R3832 GNDA.n35 GNDA.n31 585
R3833 GNDA.n30 GNDA.n0 585
R3834 GNDA.n5389 GNDA.n1 585
R3835 GNDA.n5391 GNDA.n5390 585
R3836 GNDA.n5395 GNDA.n5394 585
R3837 GNDA.n5397 GNDA.n5396 585
R3838 GNDA.n5386 GNDA.n5385 585
R3839 GNDA.n5376 GNDA.n89 585
R3840 GNDA.n5380 GNDA.n89 585
R3841 GNDA.n5378 GNDA.n5377 585
R3842 GNDA.n5379 GNDA.n5378 585
R3843 GNDA.n5375 GNDA.n91 585
R3844 GNDA.n91 GNDA.n90 585
R3845 GNDA.n5374 GNDA.n5373 585
R3846 GNDA.n5373 GNDA.n5372 585
R3847 GNDA.n93 GNDA.n92 585
R3848 GNDA.n5371 GNDA.n93 585
R3849 GNDA.n4919 GNDA.n4918 585
R3850 GNDA.n4918 GNDA.n110 585
R3851 GNDA.n4921 GNDA.n4920 585
R3852 GNDA.n4922 GNDA.n4921 585
R3853 GNDA.n427 GNDA.n426 585
R3854 GNDA.n4923 GNDA.n427 585
R3855 GNDA.n4926 GNDA.n4925 585
R3856 GNDA.n4925 GNDA.n4924 585
R3857 GNDA.n4927 GNDA.n425 585
R3858 GNDA.n425 GNDA.n424 585
R3859 GNDA.n4929 GNDA.n4928 585
R3860 GNDA.n4930 GNDA.n4929 585
R3861 GNDA.n423 GNDA.n422 585
R3862 GNDA.n4931 GNDA.n423 585
R3863 GNDA.n4934 GNDA.n4933 585
R3864 GNDA.n4933 GNDA.n4932 585
R3865 GNDA.n4935 GNDA.n421 585
R3866 GNDA.n421 GNDA.n420 585
R3867 GNDA.n4937 GNDA.n4936 585
R3868 GNDA.n4938 GNDA.n4937 585
R3869 GNDA.n419 GNDA.n418 585
R3870 GNDA.n4939 GNDA.n419 585
R3871 GNDA.n4942 GNDA.n4941 585
R3872 GNDA.n4941 GNDA.n4940 585
R3873 GNDA.n4943 GNDA.n417 585
R3874 GNDA.n417 GNDA.n416 585
R3875 GNDA.n4945 GNDA.n4944 585
R3876 GNDA.n4946 GNDA.n4945 585
R3877 GNDA.n415 GNDA.n414 585
R3878 GNDA.n4947 GNDA.n415 585
R3879 GNDA.n4950 GNDA.n4949 585
R3880 GNDA.n4949 GNDA.n4948 585
R3881 GNDA.n4951 GNDA.n413 585
R3882 GNDA.n413 GNDA.n367 585
R3883 GNDA.n4953 GNDA.n4952 585
R3884 GNDA.n4954 GNDA.n4953 585
R3885 GNDA.n4958 GNDA.n4957 585
R3886 GNDA.n4957 GNDA.n4956 585
R3887 GNDA.n4959 GNDA.n363 585
R3888 GNDA.n363 GNDA.n362 585
R3889 GNDA.n4961 GNDA.n4960 585
R3890 GNDA.n4962 GNDA.n4961 585
R3891 GNDA.n364 GNDA.n361 585
R3892 GNDA.n4963 GNDA.n361 585
R3893 GNDA.n4965 GNDA.n360 585
R3894 GNDA.n4965 GNDA.n4964 585
R3895 GNDA.n4967 GNDA.n4966 585
R3896 GNDA.n4966 GNDA.n356 585
R3897 GNDA.n354 GNDA.n353 585
R3898 GNDA.n4973 GNDA.n354 585
R3899 GNDA.n4976 GNDA.n4975 585
R3900 GNDA.n4975 GNDA.n4974 585
R3901 GNDA.n4977 GNDA.n352 585
R3902 GNDA.n352 GNDA.n351 585
R3903 GNDA.n4979 GNDA.n4978 585
R3904 GNDA.n4980 GNDA.n4979 585
R3905 GNDA.n350 GNDA.n303 585
R3906 GNDA.n4981 GNDA.n350 585
R3907 GNDA.n4984 GNDA.n4983 585
R3908 GNDA.n4983 GNDA.n4982 585
R3909 GNDA.n389 GNDA.n83 585
R3910 GNDA.n390 GNDA.n388 585
R3911 GNDA.n395 GNDA.n386 585
R3912 GNDA.n396 GNDA.n384 585
R3913 GNDA.n397 GNDA.n383 585
R3914 GNDA.n381 GNDA.n379 585
R3915 GNDA.n403 GNDA.n378 585
R3916 GNDA.n404 GNDA.n376 585
R3917 GNDA.n405 GNDA.n375 585
R3918 GNDA.n373 GNDA.n371 585
R3919 GNDA.n410 GNDA.n370 585
R3920 GNDA.n411 GNDA.n366 585
R3921 GNDA.n5458 GNDA.n84 585
R3922 GNDA.n5458 GNDA.n5457 585
R3923 GNDA.n412 GNDA.n411 585
R3924 GNDA.n410 GNDA.n409 585
R3925 GNDA.n408 GNDA.n371 585
R3926 GNDA.n406 GNDA.n405 585
R3927 GNDA.n404 GNDA.n372 585
R3928 GNDA.n403 GNDA.n402 585
R3929 GNDA.n400 GNDA.n379 585
R3930 GNDA.n398 GNDA.n397 585
R3931 GNDA.n396 GNDA.n380 585
R3932 GNDA.n395 GNDA.n394 585
R3933 GNDA.n392 GNDA.n390 585
R3934 GNDA.n389 GNDA.n86 585
R3935 GNDA.n5456 GNDA.n84 585
R3936 GNDA.n5457 GNDA.n5456 585
R3937 GNDA.n2383 GNDA.n2382 585
R3938 GNDA.n2380 GNDA.n2141 585
R3939 GNDA.n2379 GNDA.n2378 585
R3940 GNDA.n2370 GNDA.n2143 585
R3941 GNDA.n2372 GNDA.n2371 585
R3942 GNDA.n2368 GNDA.n2145 585
R3943 GNDA.n2367 GNDA.n2366 585
R3944 GNDA.n2358 GNDA.n2147 585
R3945 GNDA.n2360 GNDA.n2359 585
R3946 GNDA.n2356 GNDA.n2149 585
R3947 GNDA.n2355 GNDA.n2354 585
R3948 GNDA.n2172 GNDA.n2151 585
R3949 GNDA.n2386 GNDA.n2138 585
R3950 GNDA.n2138 GNDA.n161 585
R3951 GNDA.n2351 GNDA.n2151 585
R3952 GNDA.n2354 GNDA.n2353 585
R3953 GNDA.n2149 GNDA.n2148 585
R3954 GNDA.n2148 GNDA.n111 585
R3955 GNDA.n2361 GNDA.n2360 585
R3956 GNDA.n2363 GNDA.n2147 585
R3957 GNDA.n2366 GNDA.n2365 585
R3958 GNDA.n2145 GNDA.n2144 585
R3959 GNDA.n2373 GNDA.n2372 585
R3960 GNDA.n2375 GNDA.n2143 585
R3961 GNDA.n2378 GNDA.n2377 585
R3962 GNDA.n2141 GNDA.n2140 585
R3963 GNDA.n2384 GNDA.n2383 585
R3964 GNDA.n2384 GNDA.n111 585
R3965 GNDA.n2386 GNDA.n2385 585
R3966 GNDA.n2385 GNDA.n161 585
R3967 GNDA.n2477 GNDA.n2476 585
R3968 GNDA.n1676 GNDA.n1602 585
R3969 GNDA.n2469 GNDA.n2468 585
R3970 GNDA.n1677 GNDA.n1675 585
R3971 GNDA.n2462 GNDA.n2461 585
R3972 GNDA.n2460 GNDA.n2459 585
R3973 GNDA.n2458 GNDA.n2457 585
R3974 GNDA.n2449 GNDA.n1679 585
R3975 GNDA.n2451 GNDA.n2450 585
R3976 GNDA.n2448 GNDA.n2447 585
R3977 GNDA.n2446 GNDA.n2445 585
R3978 GNDA.n2133 GNDA.n1681 585
R3979 GNDA.n2442 GNDA.n1681 585
R3980 GNDA.n2445 GNDA.n2444 585
R3981 GNDA.n2448 GNDA.n1680 585
R3982 GNDA.n1680 GNDA.n1563 585
R3983 GNDA.n2452 GNDA.n2451 585
R3984 GNDA.n2454 GNDA.n1679 585
R3985 GNDA.n2457 GNDA.n2456 585
R3986 GNDA.n2460 GNDA.n1678 585
R3987 GNDA.n2463 GNDA.n2462 585
R3988 GNDA.n2465 GNDA.n1677 585
R3989 GNDA.n2468 GNDA.n2467 585
R3990 GNDA.n1602 GNDA.n1601 585
R3991 GNDA.n2478 GNDA.n2477 585
R3992 GNDA.n2478 GNDA.n1563 585
R3993 GNDA.n1926 GNDA.n1918 585
R3994 GNDA.n1920 GNDA.n1917 585
R3995 GNDA.n1929 GNDA.n1917 585
R3996 GNDA.n1897 GNDA.n1896 585
R3997 GNDA.n2046 GNDA.n2045 585
R3998 GNDA.n2045 GNDA.n2044 585
R3999 GNDA.n2055 GNDA.n1884 585
R4000 GNDA.n2062 GNDA.n1883 585
R4001 GNDA.n2066 GNDA.n1883 585
R4002 GNDA.n2060 GNDA.n2059 585
R4003 GNDA.n2514 GNDA.n1558 585
R4004 GNDA.n2517 GNDA.n2516 585
R4005 GNDA.n2518 GNDA.n2517 585
R4006 GNDA.n2509 GNDA.n2508 585
R4007 GNDA.n1718 GNDA.n1715 585
R4008 GNDA.n2084 GNDA.n1718 585
R4009 GNDA.n1856 GNDA.n1734 585
R4010 GNDA.n1734 GNDA.n1733 585
R4011 GNDA.n1860 GNDA.n1859 585
R4012 GNDA.n1861 GNDA.n1860 585
R4013 GNDA.n1731 GNDA.n1730 585
R4014 GNDA.n1864 GNDA.n1731 585
R4015 GNDA.n1870 GNDA.n1869 585
R4016 GNDA.n1869 GNDA.n1868 585
R4017 GNDA.n1732 GNDA.n1727 585
R4018 GNDA.n1867 GNDA.n1732 585
R4019 GNDA.n1878 GNDA.n1726 585
R4020 GNDA.n1726 GNDA.n106 585
R4021 GNDA.n1881 GNDA.n1880 585
R4022 GNDA.n2067 GNDA.n1881 585
R4023 GNDA.n2071 GNDA.n2070 585
R4024 GNDA.n2070 GNDA.n2069 585
R4025 GNDA.n1723 GNDA.n1719 585
R4026 GNDA.n2068 GNDA.n1719 585
R4027 GNDA.n2081 GNDA.n2080 585
R4028 GNDA.n2082 GNDA.n2081 585
R4029 GNDA.n1721 GNDA.n1717 585
R4030 GNDA.n2083 GNDA.n1717 585
R4031 GNDA.n2087 GNDA.n2086 585
R4032 GNDA.n2086 GNDA.n2085 585
R4033 GNDA.n2475 GNDA.n1600 585
R4034 GNDA.n2475 GNDA.n2474 585
R4035 GNDA.n1912 GNDA.n1715 585
R4036 GNDA.n1912 GNDA.n1661 585
R4037 GNDA.n1931 GNDA.n1714 585
R4038 GNDA.n1931 GNDA.n1930 585
R4039 GNDA.n1996 GNDA.n1932 585
R4040 GNDA.n1932 GNDA.n1911 585
R4041 GNDA.n2006 GNDA.n2005 585
R4042 GNDA.n2007 GNDA.n2006 585
R4043 GNDA.n1934 GNDA.n1910 585
R4044 GNDA.n2008 GNDA.n1910 585
R4045 GNDA.n2012 GNDA.n2011 585
R4046 GNDA.n2011 GNDA.n2010 585
R4047 GNDA.n2013 GNDA.n1905 585
R4048 GNDA.n2009 GNDA.n1905 585
R4049 GNDA.n2022 GNDA.n2021 585
R4050 GNDA.n2023 GNDA.n2022 585
R4051 GNDA.n1906 GNDA.n1904 585
R4052 GNDA.n2024 GNDA.n1904 585
R4053 GNDA.n2028 GNDA.n2027 585
R4054 GNDA.n2027 GNDA.n2026 585
R4055 GNDA.n2029 GNDA.n1898 585
R4056 GNDA.n2025 GNDA.n1898 585
R4057 GNDA.n2039 GNDA.n2038 585
R4058 GNDA.n2040 GNDA.n2039 585
R4059 GNDA.n2036 GNDA.n1658 585
R4060 GNDA.n2041 GNDA.n1658 585
R4061 GNDA.n2479 GNDA.n1600 585
R4062 GNDA.n2480 GNDA.n2479 585
R4063 GNDA.n1655 GNDA.n1599 585
R4064 GNDA.n2481 GNDA.n1599 585
R4065 GNDA.n2483 GNDA.n1597 585
R4066 GNDA.n2483 GNDA.n2482 585
R4067 GNDA.n2498 GNDA.n2497 585
R4068 GNDA.n2497 GNDA.n2496 585
R4069 GNDA.n2485 GNDA.n2484 585
R4070 GNDA.n2495 GNDA.n2484 585
R4071 GNDA.n2493 GNDA.n2492 585
R4072 GNDA.n2494 GNDA.n2493 585
R4073 GNDA.n2488 GNDA.n1564 585
R4074 GNDA.n1564 GNDA.n1559 585
R4075 GNDA.n2506 GNDA.n2505 585
R4076 GNDA.n2507 GNDA.n2506 585
R4077 GNDA.n1566 GNDA.n1565 585
R4078 GNDA.n1574 GNDA.n1565 585
R4079 GNDA.n1577 GNDA.n1576 585
R4080 GNDA.n1576 GNDA.n1575 585
R4081 GNDA.n1578 GNDA.n1446 585
R4082 GNDA.n1446 GNDA.n1444 585
R4083 GNDA.n2543 GNDA.n2542 585
R4084 GNDA.n2544 GNDA.n2543 585
R4085 GNDA.n2540 GNDA.n1447 585
R4086 GNDA.n1447 GNDA.n1445 585
R4087 GNDA.n1833 GNDA.n1832 585
R4088 GNDA.n1835 GNDA.n1834 585
R4089 GNDA.n1837 GNDA.n1836 585
R4090 GNDA.n1839 GNDA.n1838 585
R4091 GNDA.n1841 GNDA.n1840 585
R4092 GNDA.n1843 GNDA.n1842 585
R4093 GNDA.n1845 GNDA.n1844 585
R4094 GNDA.n1847 GNDA.n1846 585
R4095 GNDA.n1849 GNDA.n1848 585
R4096 GNDA.n1851 GNDA.n1850 585
R4097 GNDA.n1853 GNDA.n1852 585
R4098 GNDA.n5150 GNDA.n280 585
R4099 GNDA.n262 GNDA.n261 585
R4100 GNDA.n264 GNDA.n263 585
R4101 GNDA.n266 GNDA.n265 585
R4102 GNDA.n268 GNDA.n267 585
R4103 GNDA.n270 GNDA.n269 585
R4104 GNDA.n272 GNDA.n271 585
R4105 GNDA.n274 GNDA.n273 585
R4106 GNDA.n275 GNDA.n240 585
R4107 GNDA.n278 GNDA.n277 585
R4108 GNDA.n276 GNDA.n239 585
R4109 GNDA.n229 GNDA.n228 585
R4110 GNDA.n5150 GNDA.n229 585
R4111 GNDA.n5153 GNDA.n5152 585
R4112 GNDA.n5153 GNDA.n227 585
R4113 GNDA.n5148 GNDA.n5147 585
R4114 GNDA.n5146 GNDA.n288 585
R4115 GNDA.n5145 GNDA.n287 585
R4116 GNDA.n5150 GNDA.n287 585
R4117 GNDA.n5144 GNDA.n5143 585
R4118 GNDA.n5142 GNDA.n5141 585
R4119 GNDA.n5140 GNDA.n5139 585
R4120 GNDA.n5138 GNDA.n5137 585
R4121 GNDA.n5136 GNDA.n5135 585
R4122 GNDA.n5134 GNDA.n5133 585
R4123 GNDA.n5132 GNDA.n5131 585
R4124 GNDA.n5130 GNDA.n5129 585
R4125 GNDA.n5128 GNDA.n5127 585
R4126 GNDA.n5127 GNDA.n5126 585
R4127 GNDA.n666 GNDA.n643 582.4
R4128 GNDA.n740 GNDA.n734 582.4
R4129 GNDA.n646 GNDA.t267 548.082
R4130 GNDA.n664 GNDA.t256 546.375
R4131 GNDA.n693 GNDA.t202 546.375
R4132 GNDA.n606 GNDA.t211 546.375
R4133 GNDA.n4132 GNDA.t193 524.808
R4134 GNDA.n4281 GNDA.t179 524.808
R4135 GNDA.n3385 GNDA.t269 524.808
R4136 GNDA.n3481 GNDA.t262 524.808
R4137 GNDA.n4091 GNDA.t200 509.2
R4138 GNDA.n4089 GNDA.t196 509.2
R4139 GNDA.n4007 GNDA.t272 509.034
R4140 GNDA.n3995 GNDA.t205 509.034
R4141 GNDA.n735 GNDA.t229 492.675
R4142 GNDA.n738 GNDA.t254 492.675
R4143 GNDA.n638 GNDA.t252 492.675
R4144 GNDA.n641 GNDA.t265 492.675
R4145 GNDA.t186 GNDA.n88 486.94
R4146 GNDA.t186 GNDA.n103 486.94
R4147 GNDA.n4053 GNDA.n4052 483.2
R4148 GNDA.n4052 GNDA.n4051 476.8
R4149 GNDA.n1439 GNDA.t247 425.134
R4150 GNDA.n1429 GNDA.t231 425.134
R4151 GNDA.t47 GNDA.n4005 415.557
R4152 GNDA.n1426 GNDA.t182 409.067
R4153 GNDA.n2547 GNDA.t235 409.067
R4154 GNDA.n1440 GNDA.t190 409.067
R4155 GNDA.n1435 GNDA.t221 409.067
R4156 GNDA.n1434 GNDA.t187 409.067
R4157 GNDA.n1430 GNDA.t274 409.067
R4158 GNDA.n4930 GNDA.n424 394.817
R4159 GNDA.n4924 GNDA.n4923 394.817
R4160 GNDA.n4923 GNDA.n4922 394.817
R4161 GNDA.n4922 GNDA.n110 394.817
R4162 GNDA.n5372 GNDA.n5371 394.817
R4163 GNDA.n5372 GNDA.n90 394.817
R4164 GNDA.n5379 GNDA.n90 394.817
R4165 GNDA.n5380 GNDA.n5379 394.817
R4166 GNDA.n5381 GNDA.n5380 394.817
R4167 GNDA.n5381 GNDA.n88 394.817
R4168 GNDA.n2325 GNDA.n2324 394.817
R4169 GNDA.n2324 GNDA.n2323 394.817
R4170 GNDA.n2323 GNDA.n2178 394.817
R4171 GNDA.n2317 GNDA.n2178 394.817
R4172 GNDA.n2317 GNDA.n109 394.817
R4173 GNDA.n2185 GNDA.n108 394.817
R4174 GNDA.n2310 GNDA.n2185 394.817
R4175 GNDA.n2310 GNDA.n2309 394.817
R4176 GNDA.n2309 GNDA.n2308 394.817
R4177 GNDA.n2308 GNDA.n2186 394.817
R4178 GNDA.n2186 GNDA.n103 394.817
R4179 GNDA.n2418 GNDA.n102 394.817
R4180 GNDA.n2418 GNDA.n2417 394.817
R4181 GNDA.n2417 GNDA.n2416 394.817
R4182 GNDA.n2416 GNDA.n2400 394.817
R4183 GNDA.n2400 GNDA.n1561 394.817
R4184 GNDA.n2408 GNDA.n1562 394.817
R4185 GNDA.n2408 GNDA.n2407 394.817
R4186 GNDA.n2407 GNDA.n1454 394.817
R4187 GNDA.n2536 GNDA.n1454 394.817
R4188 GNDA.n2536 GNDA.n2535 394.817
R4189 GNDA.n2535 GNDA.n2534 394.817
R4190 GNDA.n4002 GNDA.n4001 384
R4191 GNDA.n4917 GNDA.n424 377.269
R4192 GNDA.n300 GNDA.n96 370.214
R4193 GNDA.n4955 GNDA.n98 370.214
R4194 GNDA.n300 GNDA.n95 365.957
R4195 GNDA.n4955 GNDA.n97 365.957
R4196 GNDA.n4001 GNDA.n4000 355.2
R4197 GNDA.n4003 GNDA.n4002 345.601
R4198 GNDA.t186 GNDA.n94 172.876
R4199 GNDA.t186 GNDA.n95 327.661
R4200 GNDA.t186 GNDA.n97 327.661
R4201 GNDA.n2471 GNDA.t186 172.876
R4202 GNDA.t186 GNDA.n1662 172.615
R4203 GNDA.t186 GNDA.n96 323.404
R4204 GNDA.t186 GNDA.n98 323.404
R4205 GNDA.t186 GNDA.n1563 172.615
R4206 GNDA.n4003 GNDA.n4000 316.8
R4207 GNDA.t47 GNDA.n3996 293.651
R4208 GNDA.n4006 GNDA.t47 293.651
R4209 GNDA.n4059 GNDA.n4058 292.5
R4210 GNDA.n4060 GNDA.n4059 292.5
R4211 GNDA.n644 GNDA.n600 292.5
R4212 GNDA.n4121 GNDA.n600 292.5
R4213 GNDA.n4120 GNDA.n4119 292.5
R4214 GNDA.n4121 GNDA.n4120 292.5
R4215 GNDA.n4001 GNDA.n3997 292.5
R4216 GNDA.n4005 GNDA.n3997 292.5
R4217 GNDA.n4002 GNDA.n3999 292.5
R4218 GNDA.n4004 GNDA.n4003 292.5
R4219 GNDA.n4005 GNDA.n4004 292.5
R4220 GNDA.n4000 GNDA.n3998 292.5
R4221 GNDA.n3998 GNDA.n760 292.5
R4222 GNDA.n4052 GNDA.n746 292.5
R4223 GNDA.n759 GNDA.n746 292.5
R4224 GNDA.n747 GNDA.n745 292.5
R4225 GNDA.n745 GNDA.n744 292.5
R4226 GNDA.n742 GNDA.n741 292.5
R4227 GNDA.n743 GNDA.n742 292.5
R4228 GNDA.n729 GNDA.n728 292.5
R4229 GNDA.n728 GNDA.n727 292.5
R4230 GNDA.n687 GNDA.n602 292.5
R4231 GNDA.n726 GNDA.n602 292.5
R4232 GNDA.n686 GNDA.n601 292.5
R4233 GNDA.n725 GNDA.n601 292.5
R4234 GNDA.n678 GNDA.n673 292.5
R4235 GNDA.n673 GNDA.n671 292.5
R4236 GNDA.n723 GNDA.n722 292.5
R4237 GNDA.n724 GNDA.n723 292.5
R4238 GNDA.n675 GNDA.n672 292.5
R4239 GNDA.n672 GNDA.n671 292.5
R4240 GNDA.n677 GNDA.n676 292.5
R4241 GNDA.n4046 GNDA.n4045 292.5
R4242 GNDA.n4045 GNDA.n4044 292.5
R4243 GNDA.n663 GNDA.n637 292.5
R4244 GNDA.n637 GNDA.n632 292.5
R4245 GNDA.n690 GNDA.n689 292.5
R4246 GNDA.n689 GNDA.n632 292.5
R4247 GNDA.t186 GNDA.n110 267.598
R4248 GNDA.t186 GNDA.n109 267.598
R4249 GNDA.t186 GNDA.n1561 267.598
R4250 GNDA.n2539 GNDA.n1450 264.301
R4251 GNDA.n2305 GNDA.n2304 264.301
R4252 GNDA.n5383 GNDA.n87 264.301
R4253 GNDA.n1855 GNDA.n1854 264.301
R4254 GNDA.n5151 GNDA.n5150 264.301
R4255 GNDA.n5150 GNDA.n234 264.301
R4256 GNDA.n2530 GNDA.t15 260
R4257 GNDA.n2528 GNDA.t15 260
R4258 GNDA.n2421 GNDA.n2420 259.416
R4259 GNDA.n2134 GNDA.n2133 259.416
R4260 GNDA.n1811 GNDA.n1690 259.416
R4261 GNDA.n4957 GNDA.n366 259.416
R4262 GNDA.n2327 GNDA.n2326 259.416
R4263 GNDA.n2173 GNDA.n2172 259.416
R4264 GNDA.n5368 GNDA.n130 259.416
R4265 GNDA.n4987 GNDA.n301 259.416
R4266 GNDA.n4929 GNDA.n423 259.416
R4267 GNDA.n1637 GNDA.n1636 258.334
R4268 GNDA.n1981 GNDA.n1939 258.334
R4269 GNDA.n5313 GNDA.n5312 258.334
R4270 GNDA.n5098 GNDA.n5097 258.334
R4271 GNDA.n2246 GNDA.n2245 258.334
R4272 GNDA.n5237 GNDA.n5177 258.334
R4273 GNDA.n5516 GNDA.n80 258.334
R4274 GNDA.n1784 GNDA.n1782 258.334
R4275 GNDA.n5436 GNDA.n5435 258.334
R4276 GNDA.t186 GNDA.n4972 257.779
R4277 GNDA.n759 GNDA.n636 256.668
R4278 GNDA.n5370 GNDA.n5369 254.34
R4279 GNDA.n5370 GNDA.n128 254.34
R4280 GNDA.n5370 GNDA.n127 254.34
R4281 GNDA.n5370 GNDA.n126 254.34
R4282 GNDA.n5370 GNDA.n125 254.34
R4283 GNDA.n5370 GNDA.n124 254.34
R4284 GNDA.n5370 GNDA.n123 254.34
R4285 GNDA.n5370 GNDA.n122 254.34
R4286 GNDA.n5370 GNDA.n121 254.34
R4287 GNDA.n5370 GNDA.n120 254.34
R4288 GNDA.n5370 GNDA.n119 254.34
R4289 GNDA.n5370 GNDA.n118 254.34
R4290 GNDA.n5370 GNDA.n117 254.34
R4291 GNDA.n5370 GNDA.n116 254.34
R4292 GNDA.n5370 GNDA.n115 254.34
R4293 GNDA.n5370 GNDA.n114 254.34
R4294 GNDA.n5370 GNDA.n113 254.34
R4295 GNDA.n5370 GNDA.n112 254.34
R4296 GNDA.n5550 GNDA.n5549 254.34
R4297 GNDA.n5550 GNDA.n53 254.34
R4298 GNDA.n5550 GNDA.n52 254.34
R4299 GNDA.n5550 GNDA.n51 254.34
R4300 GNDA.n5550 GNDA.n50 254.34
R4301 GNDA.n5550 GNDA.n49 254.34
R4302 GNDA.n5550 GNDA.n48 254.34
R4303 GNDA.n5550 GNDA.n47 254.34
R4304 GNDA.n5550 GNDA.n46 254.34
R4305 GNDA.n5550 GNDA.n45 254.34
R4306 GNDA.n5550 GNDA.n44 254.34
R4307 GNDA.n5550 GNDA.n43 254.34
R4308 GNDA.n324 GNDA.n95 254.34
R4309 GNDA.n321 GNDA.n95 254.34
R4310 GNDA.n316 GNDA.n95 254.34
R4311 GNDA.n313 GNDA.n95 254.34
R4312 GNDA.n308 GNDA.n95 254.34
R4313 GNDA.n305 GNDA.n95 254.34
R4314 GNDA.n348 GNDA.n96 254.34
R4315 GNDA.n342 GNDA.n96 254.34
R4316 GNDA.n340 GNDA.n96 254.34
R4317 GNDA.n334 GNDA.n96 254.34
R4318 GNDA.n332 GNDA.n96 254.34
R4319 GNDA.n326 GNDA.n96 254.34
R4320 GNDA.n158 GNDA.n157 254.34
R4321 GNDA.n157 GNDA.n156 254.34
R4322 GNDA.n157 GNDA.n155 254.34
R4323 GNDA.n157 GNDA.n154 254.34
R4324 GNDA.n157 GNDA.n153 254.34
R4325 GNDA.n157 GNDA.n152 254.34
R4326 GNDA.n5363 GNDA.n5362 254.34
R4327 GNDA.n5362 GNDA.n5361 254.34
R4328 GNDA.n5362 GNDA.n140 254.34
R4329 GNDA.n5362 GNDA.n139 254.34
R4330 GNDA.n5362 GNDA.n138 254.34
R4331 GNDA.n5362 GNDA.n137 254.34
R4332 GNDA.n1712 GNDA.n94 254.34
R4333 GNDA.n1709 GNDA.n94 254.34
R4334 GNDA.n1704 GNDA.n94 254.34
R4335 GNDA.n1701 GNDA.n94 254.34
R4336 GNDA.n1696 GNDA.n94 254.34
R4337 GNDA.n1691 GNDA.n94 254.34
R4338 GNDA.n1689 GNDA.n1662 254.34
R4339 GNDA.n1694 GNDA.n1662 254.34
R4340 GNDA.n2100 GNDA.n1662 254.34
R4341 GNDA.n2094 GNDA.n1662 254.34
R4342 GNDA.n2092 GNDA.n1662 254.34
R4343 GNDA.n1810 GNDA.n104 254.34
R4344 GNDA.n1816 GNDA.n104 254.34
R4345 GNDA.n1808 GNDA.n104 254.34
R4346 GNDA.n1823 GNDA.n104 254.34
R4347 GNDA.n1805 GNDA.n104 254.34
R4348 GNDA.n1830 GNDA.n104 254.34
R4349 GNDA.n2132 GNDA.n104 254.34
R4350 GNDA.n1683 GNDA.n104 254.34
R4351 GNDA.n2125 GNDA.n104 254.34
R4352 GNDA.n2119 GNDA.n104 254.34
R4353 GNDA.n2117 GNDA.n104 254.34
R4354 GNDA.n2111 GNDA.n104 254.34
R4355 GNDA.n2397 GNDA.n104 254.34
R4356 GNDA.n2426 GNDA.n104 254.34
R4357 GNDA.n2394 GNDA.n104 254.34
R4358 GNDA.n2433 GNDA.n104 254.34
R4359 GNDA.n2391 GNDA.n104 254.34
R4360 GNDA.n2440 GNDA.n104 254.34
R4361 GNDA.n5271 GNDA.n5270 254.34
R4362 GNDA.n5271 GNDA.n225 254.34
R4363 GNDA.n5271 GNDA.n224 254.34
R4364 GNDA.n5271 GNDA.n223 254.34
R4365 GNDA.n5271 GNDA.n222 254.34
R4366 GNDA.n5271 GNDA.n221 254.34
R4367 GNDA.n5271 GNDA.n163 254.34
R4368 GNDA.n5271 GNDA.n166 254.34
R4369 GNDA.n5271 GNDA.n220 254.34
R4370 GNDA.n5271 GNDA.n197 254.34
R4371 GNDA.n5271 GNDA.n196 254.34
R4372 GNDA.n5272 GNDA.n5271 254.34
R4373 GNDA.n5271 GNDA.n195 254.34
R4374 GNDA.n5271 GNDA.n194 254.34
R4375 GNDA.n5271 GNDA.n193 254.34
R4376 GNDA.n5271 GNDA.n192 254.34
R4377 GNDA.n5271 GNDA.n191 254.34
R4378 GNDA.n5271 GNDA.n190 254.34
R4379 GNDA.n5550 GNDA.n42 254.34
R4380 GNDA.n5551 GNDA.n5550 254.34
R4381 GNDA.n5550 GNDA.n41 254.34
R4382 GNDA.n5550 GNDA.n29 254.34
R4383 GNDA.n5550 GNDA.n28 254.34
R4384 GNDA.n5550 GNDA.n27 254.34
R4385 GNDA.n387 GNDA.n97 254.34
R4386 GNDA.n385 GNDA.n97 254.34
R4387 GNDA.n382 GNDA.n97 254.34
R4388 GNDA.n377 GNDA.n97 254.34
R4389 GNDA.n374 GNDA.n97 254.34
R4390 GNDA.n369 GNDA.n97 254.34
R4391 GNDA.n368 GNDA.n98 254.34
R4392 GNDA.n407 GNDA.n98 254.34
R4393 GNDA.n401 GNDA.n98 254.34
R4394 GNDA.n399 GNDA.n98 254.34
R4395 GNDA.n393 GNDA.n98 254.34
R4396 GNDA.n391 GNDA.n98 254.34
R4397 GNDA.n2381 GNDA.n101 254.34
R4398 GNDA.n2142 GNDA.n101 254.34
R4399 GNDA.n2369 GNDA.n101 254.34
R4400 GNDA.n2146 GNDA.n101 254.34
R4401 GNDA.n2357 GNDA.n101 254.34
R4402 GNDA.n2150 GNDA.n101 254.34
R4403 GNDA.n2352 GNDA.n111 254.34
R4404 GNDA.n2362 GNDA.n111 254.34
R4405 GNDA.n2364 GNDA.n111 254.34
R4406 GNDA.n2374 GNDA.n111 254.34
R4407 GNDA.n2376 GNDA.n111 254.34
R4408 GNDA.n2471 GNDA.n1657 254.34
R4409 GNDA.n2471 GNDA.n2470 254.34
R4410 GNDA.n2471 GNDA.n1674 254.34
R4411 GNDA.n2471 GNDA.n1673 254.34
R4412 GNDA.n2471 GNDA.n1672 254.34
R4413 GNDA.n2471 GNDA.n1671 254.34
R4414 GNDA.n2443 GNDA.n1563 254.34
R4415 GNDA.n2453 GNDA.n1563 254.34
R4416 GNDA.n2455 GNDA.n1563 254.34
R4417 GNDA.n2464 GNDA.n1563 254.34
R4418 GNDA.n2466 GNDA.n1563 254.34
R4419 GNDA.n5150 GNDA.n286 254.34
R4420 GNDA.n5150 GNDA.n285 254.34
R4421 GNDA.n5150 GNDA.n284 254.34
R4422 GNDA.n5150 GNDA.n283 254.34
R4423 GNDA.n5150 GNDA.n282 254.34
R4424 GNDA.n5150 GNDA.n281 254.34
R4425 GNDA.n5150 GNDA.n235 254.34
R4426 GNDA.n5150 GNDA.n236 254.34
R4427 GNDA.n5150 GNDA.n237 254.34
R4428 GNDA.n5150 GNDA.n238 254.34
R4429 GNDA.n5150 GNDA.n279 254.34
R4430 GNDA.n5150 GNDA.n5149 254.34
R4431 GNDA.n5150 GNDA.n230 254.34
R4432 GNDA.n5150 GNDA.n231 254.34
R4433 GNDA.n5150 GNDA.n232 254.34
R4434 GNDA.n5150 GNDA.n233 254.34
R4435 GNDA.n1929 GNDA.n1928 250.349
R4436 GNDA.n2044 GNDA.n2043 250.349
R4437 GNDA.n2442 GNDA.n2441 249.663
R4438 GNDA.n2112 GNDA.n2110 249.663
R4439 GNDA.n1832 GNDA.n1831 249.663
R4440 GNDA.n4983 GNDA.n349 249.663
R4441 GNDA.n2351 GNDA.n2350 249.663
R4442 GNDA.n5364 GNDA.n135 249.663
R4443 GNDA.n261 GNDA.n260 249.663
R4444 GNDA.n5148 GNDA.n289 249.663
R4445 GNDA.n4953 GNDA.n412 249.663
R4446 GNDA.n678 GNDA.n677 249.601
R4447 GNDA.n677 GNDA.n675 249.601
R4448 GNDA.n2517 GNDA.n1558 246.25
R4449 GNDA.n2517 GNDA.n2508 246.25
R4450 GNDA.n1884 GNDA.n1883 246.25
R4451 GNDA.n2059 GNDA.n1883 246.25
R4452 GNDA.n2531 GNDA.n1457 246.25
R4453 GNDA.n2066 GNDA.n2065 241.643
R4454 GNDA.n2066 GNDA.n1882 241.643
R4455 GNDA.n2519 GNDA.n2518 241.643
R4456 GNDA.n2518 GNDA.n1560 241.643
R4457 GNDA.t74 GNDA.t232 227.873
R4458 GNDA.n2532 GNDA.t14 219.343
R4459 GNDA.n1456 GNDA.t14 219.343
R4460 GNDA.n2045 GNDA.n1897 197
R4461 GNDA.n1918 GNDA.n1917 197
R4462 GNDA.n2533 GNDA.n1447 197
R4463 GNDA.n2475 GNDA.n1658 197
R4464 GNDA.n2086 GNDA.n1718 197
R4465 GNDA.n2303 GNDA.n2302 197
R4466 GNDA.n2138 GNDA.n189 197
R4467 GNDA.n5180 GNDA.n5179 197
R4468 GNDA.n5031 GNDA.n85 197
R4469 GNDA.n5459 GNDA.n5458 197
R4470 GNDA.n5385 GNDA.n5384 197
R4471 GNDA.n2479 GNDA.n1599 187.249
R4472 GNDA.n1931 GNDA.n1912 187.249
R4473 GNDA.n1734 GNDA.n280 187.249
R4474 GNDA.n2385 GNDA.n2139 187.249
R4475 GNDA.n5341 GNDA.n5340 187.249
R4476 GNDA.n5269 GNDA.n227 187.249
R4477 GNDA.n5126 GNDA.n5125 187.249
R4478 GNDA.n5548 GNDA.n55 187.249
R4479 GNDA.n5456 GNDA.n5455 187.249
R4480 GNDA.n1638 GNDA.n1637 185
R4481 GNDA.n1640 GNDA.n1639 185
R4482 GNDA.n1642 GNDA.n1641 185
R4483 GNDA.n1644 GNDA.n1643 185
R4484 GNDA.n1646 GNDA.n1645 185
R4485 GNDA.n1648 GNDA.n1647 185
R4486 GNDA.n1650 GNDA.n1649 185
R4487 GNDA.n1652 GNDA.n1651 185
R4488 GNDA.n1653 GNDA.n1595 185
R4489 GNDA.n1620 GNDA.n1619 185
R4490 GNDA.n1622 GNDA.n1621 185
R4491 GNDA.n1624 GNDA.n1623 185
R4492 GNDA.n1626 GNDA.n1625 185
R4493 GNDA.n1628 GNDA.n1627 185
R4494 GNDA.n1630 GNDA.n1629 185
R4495 GNDA.n1632 GNDA.n1631 185
R4496 GNDA.n1634 GNDA.n1633 185
R4497 GNDA.n1636 GNDA.n1635 185
R4498 GNDA.n1587 GNDA.n1449 185
R4499 GNDA.n1604 GNDA.n1603 185
R4500 GNDA.n1606 GNDA.n1605 185
R4501 GNDA.n1608 GNDA.n1607 185
R4502 GNDA.n1610 GNDA.n1609 185
R4503 GNDA.n1612 GNDA.n1611 185
R4504 GNDA.n1614 GNDA.n1613 185
R4505 GNDA.n1616 GNDA.n1615 185
R4506 GNDA.n1618 GNDA.n1617 185
R4507 GNDA.n1586 GNDA.n1448 185
R4508 GNDA.n1580 GNDA.n1579 185
R4509 GNDA.n1573 GNDA.n1568 185
R4510 GNDA.n2504 GNDA.n2503 185
R4511 GNDA.n2487 GNDA.n1567 185
R4512 GNDA.n2491 GNDA.n2490 185
R4513 GNDA.n2489 GNDA.n2486 185
R4514 GNDA.n1598 GNDA.n1596 185
R4515 GNDA.n2500 GNDA.n2499 185
R4516 GNDA.n1981 GNDA.n1980 185
R4517 GNDA.n1983 GNDA.n1938 185
R4518 GNDA.n1986 GNDA.n1985 185
R4519 GNDA.n1987 GNDA.n1937 185
R4520 GNDA.n1989 GNDA.n1988 185
R4521 GNDA.n1991 GNDA.n1936 185
R4522 GNDA.n1994 GNDA.n1993 185
R4523 GNDA.n1995 GNDA.n1935 185
R4524 GNDA.n1999 GNDA.n1998 185
R4525 GNDA.n1963 GNDA.n1943 185
R4526 GNDA.n1965 GNDA.n1964 185
R4527 GNDA.n1967 GNDA.n1942 185
R4528 GNDA.n1970 GNDA.n1969 185
R4529 GNDA.n1971 GNDA.n1941 185
R4530 GNDA.n1973 GNDA.n1972 185
R4531 GNDA.n1975 GNDA.n1940 185
R4532 GNDA.n1978 GNDA.n1977 185
R4533 GNDA.n1979 GNDA.n1939 185
R4534 GNDA.n2035 GNDA.n2034 185
R4535 GNDA.n1948 GNDA.n1900 185
R4536 GNDA.n1950 GNDA.n1949 185
R4537 GNDA.n1952 GNDA.n1946 185
R4538 GNDA.n1954 GNDA.n1953 185
R4539 GNDA.n1955 GNDA.n1945 185
R4540 GNDA.n1957 GNDA.n1956 185
R4541 GNDA.n1959 GNDA.n1944 185
R4542 GNDA.n1962 GNDA.n1961 185
R4543 GNDA.n2033 GNDA.n1899 185
R4544 GNDA.n2031 GNDA.n2030 185
R4545 GNDA.n1903 GNDA.n1902 185
R4546 GNDA.n2020 GNDA.n2019 185
R4547 GNDA.n2017 GNDA.n1907 185
R4548 GNDA.n2015 GNDA.n2014 185
R4549 GNDA.n1909 GNDA.n1908 185
R4550 GNDA.n2004 GNDA.n2003 185
R4551 GNDA.n2001 GNDA.n1933 185
R4552 GNDA.n5314 GNDA.n5313 185
R4553 GNDA.n5316 GNDA.n5315 185
R4554 GNDA.n5318 GNDA.n5317 185
R4555 GNDA.n5320 GNDA.n5319 185
R4556 GNDA.n5322 GNDA.n5321 185
R4557 GNDA.n5324 GNDA.n5323 185
R4558 GNDA.n5326 GNDA.n5325 185
R4559 GNDA.n5328 GNDA.n5327 185
R4560 GNDA.n5329 GNDA.n164 185
R4561 GNDA.n5296 GNDA.n5295 185
R4562 GNDA.n5298 GNDA.n5297 185
R4563 GNDA.n5300 GNDA.n5299 185
R4564 GNDA.n5302 GNDA.n5301 185
R4565 GNDA.n5304 GNDA.n5303 185
R4566 GNDA.n5306 GNDA.n5305 185
R4567 GNDA.n5308 GNDA.n5307 185
R4568 GNDA.n5310 GNDA.n5309 185
R4569 GNDA.n5312 GNDA.n5311 185
R4570 GNDA.n5278 GNDA.n5277 185
R4571 GNDA.n5280 GNDA.n5279 185
R4572 GNDA.n5282 GNDA.n5281 185
R4573 GNDA.n5284 GNDA.n5283 185
R4574 GNDA.n5286 GNDA.n5285 185
R4575 GNDA.n5288 GNDA.n5287 185
R4576 GNDA.n5290 GNDA.n5289 185
R4577 GNDA.n5292 GNDA.n5291 185
R4578 GNDA.n5294 GNDA.n5293 185
R4579 GNDA.n5276 GNDA.n5275 185
R4580 GNDA.n206 GNDA.n205 185
R4581 GNDA.n204 GNDA.n203 185
R4582 GNDA.n212 GNDA.n211 185
R4583 GNDA.n214 GNDA.n213 185
R4584 GNDA.n217 GNDA.n216 185
R4585 GNDA.n200 GNDA.n169 185
R4586 GNDA.n5333 GNDA.n5332 185
R4587 GNDA.n168 GNDA.n165 185
R4588 GNDA.n5099 GNDA.n5098 185
R4589 GNDA.n5101 GNDA.n5100 185
R4590 GNDA.n5103 GNDA.n5102 185
R4591 GNDA.n5105 GNDA.n5104 185
R4592 GNDA.n5107 GNDA.n5106 185
R4593 GNDA.n5109 GNDA.n5108 185
R4594 GNDA.n5111 GNDA.n5110 185
R4595 GNDA.n5113 GNDA.n5112 185
R4596 GNDA.n5114 GNDA.n5010 185
R4597 GNDA.n5081 GNDA.n5080 185
R4598 GNDA.n5083 GNDA.n5082 185
R4599 GNDA.n5085 GNDA.n5084 185
R4600 GNDA.n5087 GNDA.n5086 185
R4601 GNDA.n5089 GNDA.n5088 185
R4602 GNDA.n5091 GNDA.n5090 185
R4603 GNDA.n5093 GNDA.n5092 185
R4604 GNDA.n5095 GNDA.n5094 185
R4605 GNDA.n5097 GNDA.n5096 185
R4606 GNDA.n5063 GNDA.n5062 185
R4607 GNDA.n5065 GNDA.n5064 185
R4608 GNDA.n5067 GNDA.n5066 185
R4609 GNDA.n5069 GNDA.n5068 185
R4610 GNDA.n5071 GNDA.n5070 185
R4611 GNDA.n5073 GNDA.n5072 185
R4612 GNDA.n5075 GNDA.n5074 185
R4613 GNDA.n5077 GNDA.n5076 185
R4614 GNDA.n5079 GNDA.n5078 185
R4615 GNDA.n2247 GNDA.n2246 185
R4616 GNDA.n2249 GNDA.n2248 185
R4617 GNDA.n2251 GNDA.n2250 185
R4618 GNDA.n2253 GNDA.n2252 185
R4619 GNDA.n2255 GNDA.n2254 185
R4620 GNDA.n2257 GNDA.n2256 185
R4621 GNDA.n2259 GNDA.n2258 185
R4622 GNDA.n2261 GNDA.n2260 185
R4623 GNDA.n2262 GNDA.n2210 185
R4624 GNDA.n2229 GNDA.n2228 185
R4625 GNDA.n2231 GNDA.n2230 185
R4626 GNDA.n2233 GNDA.n2232 185
R4627 GNDA.n2235 GNDA.n2234 185
R4628 GNDA.n2237 GNDA.n2236 185
R4629 GNDA.n2239 GNDA.n2238 185
R4630 GNDA.n2241 GNDA.n2240 185
R4631 GNDA.n2243 GNDA.n2242 185
R4632 GNDA.n2245 GNDA.n2244 185
R4633 GNDA.n2202 GNDA.n2188 185
R4634 GNDA.n2213 GNDA.n2212 185
R4635 GNDA.n2215 GNDA.n2214 185
R4636 GNDA.n2217 GNDA.n2216 185
R4637 GNDA.n2219 GNDA.n2218 185
R4638 GNDA.n2221 GNDA.n2220 185
R4639 GNDA.n2223 GNDA.n2222 185
R4640 GNDA.n2225 GNDA.n2224 185
R4641 GNDA.n2227 GNDA.n2226 185
R4642 GNDA.n2192 GNDA.n2189 185
R4643 GNDA.n2295 GNDA.n2294 185
R4644 GNDA.n2268 GNDA.n2191 185
R4645 GNDA.n2274 GNDA.n2273 185
R4646 GNDA.n2272 GNDA.n2267 185
R4647 GNDA.n2281 GNDA.n2280 185
R4648 GNDA.n2279 GNDA.n2266 185
R4649 GNDA.n2286 GNDA.n2211 185
R4650 GNDA.n2291 GNDA.n2290 185
R4651 GNDA.n5239 GNDA.n5177 185
R4652 GNDA.n5253 GNDA.n5252 185
R4653 GNDA.n5251 GNDA.n5178 185
R4654 GNDA.n5250 GNDA.n5249 185
R4655 GNDA.n5248 GNDA.n5247 185
R4656 GNDA.n5246 GNDA.n5245 185
R4657 GNDA.n5244 GNDA.n5243 185
R4658 GNDA.n5242 GNDA.n5241 185
R4659 GNDA.n5240 GNDA.n5154 185
R4660 GNDA.n5222 GNDA.n5221 185
R4661 GNDA.n5224 GNDA.n5223 185
R4662 GNDA.n5226 GNDA.n5225 185
R4663 GNDA.n5228 GNDA.n5227 185
R4664 GNDA.n5230 GNDA.n5229 185
R4665 GNDA.n5232 GNDA.n5231 185
R4666 GNDA.n5234 GNDA.n5233 185
R4667 GNDA.n5236 GNDA.n5235 185
R4668 GNDA.n5238 GNDA.n5237 185
R4669 GNDA.n5204 GNDA.n5203 185
R4670 GNDA.n5206 GNDA.n5205 185
R4671 GNDA.n5208 GNDA.n5207 185
R4672 GNDA.n5210 GNDA.n5209 185
R4673 GNDA.n5212 GNDA.n5211 185
R4674 GNDA.n5214 GNDA.n5213 185
R4675 GNDA.n5216 GNDA.n5215 185
R4676 GNDA.n5218 GNDA.n5217 185
R4677 GNDA.n5220 GNDA.n5219 185
R4678 GNDA.n5202 GNDA.n5201 185
R4679 GNDA.n5196 GNDA.n5195 185
R4680 GNDA.n5194 GNDA.n5193 185
R4681 GNDA.n5189 GNDA.n5188 185
R4682 GNDA.n5184 GNDA.n5162 185
R4683 GNDA.n5257 GNDA.n5256 185
R4684 GNDA.n5161 GNDA.n5159 185
R4685 GNDA.n5263 GNDA.n5262 185
R4686 GNDA.n5265 GNDA.n5264 185
R4687 GNDA.n2520 GNDA.n1557 185
R4688 GNDA.n2512 GNDA.n2511 185
R4689 GNDA.n2064 GNDA.n2063 185
R4690 GNDA.n2063 GNDA.n2062 185
R4691 GNDA.n2064 GNDA.n2054 185
R4692 GNDA.n2057 GNDA.n2054 185
R4693 GNDA.n5518 GNDA.n80 185
R4694 GNDA.n5532 GNDA.n5531 185
R4695 GNDA.n5530 GNDA.n81 185
R4696 GNDA.n5529 GNDA.n5528 185
R4697 GNDA.n5527 GNDA.n5526 185
R4698 GNDA.n5525 GNDA.n5524 185
R4699 GNDA.n5523 GNDA.n5522 185
R4700 GNDA.n5521 GNDA.n5520 185
R4701 GNDA.n5519 GNDA.n57 185
R4702 GNDA.n5501 GNDA.n5500 185
R4703 GNDA.n5503 GNDA.n5502 185
R4704 GNDA.n5505 GNDA.n5504 185
R4705 GNDA.n5507 GNDA.n5506 185
R4706 GNDA.n5509 GNDA.n5508 185
R4707 GNDA.n5511 GNDA.n5510 185
R4708 GNDA.n5513 GNDA.n5512 185
R4709 GNDA.n5515 GNDA.n5514 185
R4710 GNDA.n5517 GNDA.n5516 185
R4711 GNDA.n5483 GNDA.n5482 185
R4712 GNDA.n5485 GNDA.n5484 185
R4713 GNDA.n5487 GNDA.n5486 185
R4714 GNDA.n5489 GNDA.n5488 185
R4715 GNDA.n5491 GNDA.n5490 185
R4716 GNDA.n5493 GNDA.n5492 185
R4717 GNDA.n5495 GNDA.n5494 185
R4718 GNDA.n5497 GNDA.n5496 185
R4719 GNDA.n5499 GNDA.n5498 185
R4720 GNDA.n5481 GNDA.n5480 185
R4721 GNDA.n5475 GNDA.n5474 185
R4722 GNDA.n5473 GNDA.n5472 185
R4723 GNDA.n5468 GNDA.n5467 185
R4724 GNDA.n5463 GNDA.n65 185
R4725 GNDA.n5536 GNDA.n5535 185
R4726 GNDA.n64 GNDA.n62 185
R4727 GNDA.n5542 GNDA.n5541 185
R4728 GNDA.n5544 GNDA.n5543 185
R4729 GNDA.n5061 GNDA.n5060 185
R4730 GNDA.n5055 GNDA.n5054 185
R4731 GNDA.n5053 GNDA.n5052 185
R4732 GNDA.n5048 GNDA.n5047 185
R4733 GNDA.n5046 GNDA.n5045 185
R4734 GNDA.n5040 GNDA.n5039 185
R4735 GNDA.n5035 GNDA.n5014 185
R4736 GNDA.n5118 GNDA.n5117 185
R4737 GNDA.n5013 GNDA.n5011 185
R4738 GNDA.n1785 GNDA.n1784 185
R4739 GNDA.n1786 GNDA.n1738 185
R4740 GNDA.n1788 GNDA.n1787 185
R4741 GNDA.n1790 GNDA.n1737 185
R4742 GNDA.n1793 GNDA.n1792 185
R4743 GNDA.n1794 GNDA.n1736 185
R4744 GNDA.n1796 GNDA.n1795 185
R4745 GNDA.n1798 GNDA.n1735 185
R4746 GNDA.n1801 GNDA.n1800 185
R4747 GNDA.n1766 GNDA.n1743 185
R4748 GNDA.n1769 GNDA.n1768 185
R4749 GNDA.n1770 GNDA.n1742 185
R4750 GNDA.n1772 GNDA.n1771 185
R4751 GNDA.n1774 GNDA.n1741 185
R4752 GNDA.n1777 GNDA.n1776 185
R4753 GNDA.n1778 GNDA.n1740 185
R4754 GNDA.n1780 GNDA.n1779 185
R4755 GNDA.n1782 GNDA.n1739 185
R4756 GNDA.n1748 GNDA.n1722 185
R4757 GNDA.n1752 GNDA.n1749 185
R4758 GNDA.n1754 GNDA.n1753 185
R4759 GNDA.n1755 GNDA.n1747 185
R4760 GNDA.n1757 GNDA.n1756 185
R4761 GNDA.n1759 GNDA.n1745 185
R4762 GNDA.n1761 GNDA.n1760 185
R4763 GNDA.n1762 GNDA.n1744 185
R4764 GNDA.n1764 GNDA.n1763 185
R4765 GNDA.n2079 GNDA.n2078 185
R4766 GNDA.n2076 GNDA.n1720 185
R4767 GNDA.n2075 GNDA.n1724 185
R4768 GNDA.n2073 GNDA.n2072 185
R4769 GNDA.n1879 GNDA.n1725 185
R4770 GNDA.n1877 GNDA.n1876 185
R4771 GNDA.n1874 GNDA.n1728 185
R4772 GNDA.n1872 GNDA.n1871 185
R4773 GNDA.n1858 GNDA.n1729 185
R4774 GNDA.n5437 GNDA.n5436 185
R4775 GNDA.n5439 GNDA.n5438 185
R4776 GNDA.n5441 GNDA.n5440 185
R4777 GNDA.n5443 GNDA.n5442 185
R4778 GNDA.n5445 GNDA.n5444 185
R4779 GNDA.n5447 GNDA.n5446 185
R4780 GNDA.n5449 GNDA.n5448 185
R4781 GNDA.n5451 GNDA.n5450 185
R4782 GNDA.n5452 GNDA.n20 185
R4783 GNDA.n5419 GNDA.n5418 185
R4784 GNDA.n5421 GNDA.n5420 185
R4785 GNDA.n5423 GNDA.n5422 185
R4786 GNDA.n5425 GNDA.n5424 185
R4787 GNDA.n5427 GNDA.n5426 185
R4788 GNDA.n5429 GNDA.n5428 185
R4789 GNDA.n5431 GNDA.n5430 185
R4790 GNDA.n5433 GNDA.n5432 185
R4791 GNDA.n5435 GNDA.n5434 185
R4792 GNDA.n5401 GNDA.n5400 185
R4793 GNDA.n5403 GNDA.n5402 185
R4794 GNDA.n5405 GNDA.n5404 185
R4795 GNDA.n5407 GNDA.n5406 185
R4796 GNDA.n5409 GNDA.n5408 185
R4797 GNDA.n5411 GNDA.n5410 185
R4798 GNDA.n5413 GNDA.n5412 185
R4799 GNDA.n5415 GNDA.n5414 185
R4800 GNDA.n5417 GNDA.n5416 185
R4801 GNDA.n5399 GNDA.n5398 185
R4802 GNDA.n5393 GNDA.n5392 185
R4803 GNDA.n5388 GNDA.n3 185
R4804 GNDA.n5559 GNDA.n5558 185
R4805 GNDA.n34 GNDA.n2 185
R4806 GNDA.n38 GNDA.n37 185
R4807 GNDA.n36 GNDA.n33 185
R4808 GNDA.n23 GNDA.n21 185
R4809 GNDA.n5555 GNDA.n5554 185
R4810 GNDA.n2420 GNDA.n2419 175.546
R4811 GNDA.n2419 GNDA.n2398 175.546
R4812 GNDA.n2415 GNDA.n2398 175.546
R4813 GNDA.n2415 GNDA.n2401 175.546
R4814 GNDA.n2411 GNDA.n2401 175.546
R4815 GNDA.n2411 GNDA.n2410 175.546
R4816 GNDA.n2410 GNDA.n2409 175.546
R4817 GNDA.n2409 GNDA.n2404 175.546
R4818 GNDA.n2404 GNDA.n1452 175.546
R4819 GNDA.n2537 GNDA.n1452 175.546
R4820 GNDA.n2537 GNDA.n1453 175.546
R4821 GNDA.n2483 GNDA.n1599 175.546
R4822 GNDA.n2497 GNDA.n2483 175.546
R4823 GNDA.n2497 GNDA.n2484 175.546
R4824 GNDA.n2493 GNDA.n2484 175.546
R4825 GNDA.n2493 GNDA.n1564 175.546
R4826 GNDA.n2506 GNDA.n1564 175.546
R4827 GNDA.n2506 GNDA.n1565 175.546
R4828 GNDA.n1576 GNDA.n1565 175.546
R4829 GNDA.n1576 GNDA.n1446 175.546
R4830 GNDA.n2543 GNDA.n1446 175.546
R4831 GNDA.n2543 GNDA.n1447 175.546
R4832 GNDA.n2444 GNDA.n1680 175.546
R4833 GNDA.n2452 GNDA.n1680 175.546
R4834 GNDA.n2456 GNDA.n2454 175.546
R4835 GNDA.n2463 GNDA.n1678 175.546
R4836 GNDA.n2467 GNDA.n2465 175.546
R4837 GNDA.n2478 GNDA.n1601 175.546
R4838 GNDA.n2439 GNDA.n2389 175.546
R4839 GNDA.n2435 GNDA.n2434 175.546
R4840 GNDA.n2432 GNDA.n2392 175.546
R4841 GNDA.n2428 GNDA.n2427 175.546
R4842 GNDA.n2425 GNDA.n2395 175.546
R4843 GNDA.n2447 GNDA.n2446 175.546
R4844 GNDA.n2450 GNDA.n2449 175.546
R4845 GNDA.n2459 GNDA.n2458 175.546
R4846 GNDA.n2461 GNDA.n1675 175.546
R4847 GNDA.n2469 GNDA.n1676 175.546
R4848 GNDA.n2116 GNDA.n1687 175.546
R4849 GNDA.n2120 GNDA.n2118 175.546
R4850 GNDA.n2124 GNDA.n1685 175.546
R4851 GNDA.n2127 GNDA.n2126 175.546
R4852 GNDA.n2131 GNDA.n2130 175.546
R4853 GNDA.n1932 GNDA.n1931 175.546
R4854 GNDA.n2006 GNDA.n1932 175.546
R4855 GNDA.n2006 GNDA.n1910 175.546
R4856 GNDA.n2011 GNDA.n1910 175.546
R4857 GNDA.n2011 GNDA.n1905 175.546
R4858 GNDA.n2022 GNDA.n1905 175.546
R4859 GNDA.n2022 GNDA.n1904 175.546
R4860 GNDA.n2027 GNDA.n1904 175.546
R4861 GNDA.n2027 GNDA.n1898 175.546
R4862 GNDA.n2039 GNDA.n1898 175.546
R4863 GNDA.n2039 GNDA.n1658 175.546
R4864 GNDA.n2107 GNDA.n2106 175.546
R4865 GNDA.n2106 GNDA.n2105 175.546
R4866 GNDA.n2102 GNDA.n2101 175.546
R4867 GNDA.n2099 GNDA.n1700 175.546
R4868 GNDA.n2095 GNDA.n2093 175.546
R4869 GNDA.n2091 GNDA.n1708 175.546
R4870 GNDA.n1836 GNDA.n1835 175.546
R4871 GNDA.n1840 GNDA.n1839 175.546
R4872 GNDA.n1844 GNDA.n1843 175.546
R4873 GNDA.n1848 GNDA.n1847 175.546
R4874 GNDA.n1852 GNDA.n1851 175.546
R4875 GNDA.n1829 GNDA.n1803 175.546
R4876 GNDA.n1825 GNDA.n1824 175.546
R4877 GNDA.n1822 GNDA.n1806 175.546
R4878 GNDA.n1818 GNDA.n1817 175.546
R4879 GNDA.n1815 GNDA.n1809 175.546
R4880 GNDA.n1860 GNDA.n1734 175.546
R4881 GNDA.n1860 GNDA.n1731 175.546
R4882 GNDA.n1869 GNDA.n1731 175.546
R4883 GNDA.n1869 GNDA.n1732 175.546
R4884 GNDA.n1732 GNDA.n1726 175.546
R4885 GNDA.n1881 GNDA.n1726 175.546
R4886 GNDA.n2070 GNDA.n1881 175.546
R4887 GNDA.n2070 GNDA.n1719 175.546
R4888 GNDA.n2081 GNDA.n1719 175.546
R4889 GNDA.n2081 GNDA.n1717 175.546
R4890 GNDA.n2086 GNDA.n1717 175.546
R4891 GNDA.n1695 GNDA.n1692 175.546
R4892 GNDA.n1698 GNDA.n1697 175.546
R4893 GNDA.n1703 GNDA.n1702 175.546
R4894 GNDA.n1706 GNDA.n1705 175.546
R4895 GNDA.n1711 GNDA.n1710 175.546
R4896 GNDA.n373 GNDA.n370 175.546
R4897 GNDA.n376 GNDA.n375 175.546
R4898 GNDA.n381 GNDA.n378 175.546
R4899 GNDA.n384 GNDA.n383 175.546
R4900 GNDA.n388 GNDA.n386 175.546
R4901 GNDA.n4983 GNDA.n350 175.546
R4902 GNDA.n4979 GNDA.n350 175.546
R4903 GNDA.n4979 GNDA.n352 175.546
R4904 GNDA.n4975 GNDA.n352 175.546
R4905 GNDA.n4975 GNDA.n354 175.546
R4906 GNDA.n4966 GNDA.n354 175.546
R4907 GNDA.n4966 GNDA.n4965 175.546
R4908 GNDA.n4965 GNDA.n361 175.546
R4909 GNDA.n4961 GNDA.n361 175.546
R4910 GNDA.n4961 GNDA.n363 175.546
R4911 GNDA.n4957 GNDA.n363 175.546
R4912 GNDA.n347 GNDA.n304 175.546
R4913 GNDA.n343 GNDA.n341 175.546
R4914 GNDA.n339 GNDA.n311 175.546
R4915 GNDA.n335 GNDA.n333 175.546
R4916 GNDA.n331 GNDA.n319 175.546
R4917 GNDA.n2326 GNDA.n2177 175.546
R4918 GNDA.n2322 GNDA.n2177 175.546
R4919 GNDA.n2322 GNDA.n2179 175.546
R4920 GNDA.n2318 GNDA.n2179 175.546
R4921 GNDA.n2318 GNDA.n2316 175.546
R4922 GNDA.n2316 GNDA.n2315 175.546
R4923 GNDA.n2315 GNDA.n2182 175.546
R4924 GNDA.n2311 GNDA.n2182 175.546
R4925 GNDA.n2311 GNDA.n2184 175.546
R4926 GNDA.n2307 GNDA.n2184 175.546
R4927 GNDA.n2307 GNDA.n2187 175.546
R4928 GNDA.n2288 GNDA.n2287 175.546
R4929 GNDA.n2284 GNDA.n2283 175.546
R4930 GNDA.n2277 GNDA.n2276 175.546
R4931 GNDA.n2270 GNDA.n2269 175.546
R4932 GNDA.n2298 GNDA.n2297 175.546
R4933 GNDA.n2353 GNDA.n2148 175.546
R4934 GNDA.n2361 GNDA.n2148 175.546
R4935 GNDA.n2365 GNDA.n2363 175.546
R4936 GNDA.n2373 GNDA.n2144 175.546
R4937 GNDA.n2377 GNDA.n2375 175.546
R4938 GNDA.n2384 GNDA.n2140 175.546
R4939 GNDA.n2347 GNDA.n2346 175.546
R4940 GNDA.n2343 GNDA.n2342 175.546
R4941 GNDA.n2339 GNDA.n2338 175.546
R4942 GNDA.n2335 GNDA.n2334 175.546
R4943 GNDA.n2331 GNDA.n2330 175.546
R4944 GNDA.n2356 GNDA.n2355 175.546
R4945 GNDA.n2359 GNDA.n2358 175.546
R4946 GNDA.n2368 GNDA.n2367 175.546
R4947 GNDA.n2371 GNDA.n2370 175.546
R4948 GNDA.n2380 GNDA.n2379 175.546
R4949 GNDA.n5336 GNDA.n5335 175.546
R4950 GNDA.n219 GNDA.n199 175.546
R4951 GNDA.n201 GNDA.n198 175.546
R4952 GNDA.n209 GNDA.n208 175.546
R4953 GNDA.n5273 GNDA.n188 175.546
R4954 GNDA.n5360 GNDA.n136 175.546
R4955 GNDA.n5356 GNDA.n141 175.546
R4956 GNDA.n5354 GNDA.n5353 175.546
R4957 GNDA.n5350 GNDA.n5349 175.546
R4958 GNDA.n5346 GNDA.n5345 175.546
R4959 GNDA.n2154 GNDA.n2153 175.546
R4960 GNDA.n2158 GNDA.n2157 175.546
R4961 GNDA.n2162 GNDA.n2161 175.546
R4962 GNDA.n2166 GNDA.n2165 175.546
R4963 GNDA.n2170 GNDA.n2169 175.546
R4964 GNDA.n151 GNDA.n142 175.546
R4965 GNDA.n144 GNDA.n143 175.546
R4966 GNDA.n146 GNDA.n145 175.546
R4967 GNDA.n148 GNDA.n147 175.546
R4968 GNDA.n150 GNDA.n149 175.546
R4969 GNDA.n5155 GNDA.n226 175.546
R4970 GNDA.n5260 GNDA.n5259 175.546
R4971 GNDA.n5186 GNDA.n5185 175.546
R4972 GNDA.n5191 GNDA.n5190 175.546
R4973 GNDA.n5199 GNDA.n5198 175.546
R4974 GNDA.n265 GNDA.n264 175.546
R4975 GNDA.n269 GNDA.n268 175.546
R4976 GNDA.n273 GNDA.n272 175.546
R4977 GNDA.n278 GNDA.n240 175.546
R4978 GNDA.n239 GNDA.n229 175.546
R4979 GNDA.n5152 GNDA.n229 175.546
R4980 GNDA.n257 GNDA.n256 175.546
R4981 GNDA.n253 GNDA.n252 175.546
R4982 GNDA.n249 GNDA.n248 175.546
R4983 GNDA.n245 GNDA.n244 175.546
R4984 GNDA.n241 GNDA.n129 175.546
R4985 GNDA.n307 GNDA.n306 175.546
R4986 GNDA.n312 GNDA.n309 175.546
R4987 GNDA.n315 GNDA.n314 175.546
R4988 GNDA.n320 GNDA.n317 175.546
R4989 GNDA.n323 GNDA.n322 175.546
R4990 GNDA.n5121 GNDA.n5120 175.546
R4991 GNDA.n5037 GNDA.n5036 175.546
R4992 GNDA.n5043 GNDA.n5042 175.546
R4993 GNDA.n5050 GNDA.n5049 175.546
R4994 GNDA.n5058 GNDA.n5057 175.546
R4995 GNDA.n288 GNDA.n287 175.546
R4996 GNDA.n5143 GNDA.n287 175.546
R4997 GNDA.n5141 GNDA.n5140 175.546
R4998 GNDA.n5137 GNDA.n5136 175.546
R4999 GNDA.n5133 GNDA.n5132 175.546
R5000 GNDA.n5129 GNDA.n5128 175.546
R5001 GNDA.n5007 GNDA.n289 175.546
R5002 GNDA.n5007 GNDA.n291 175.546
R5003 GNDA.n5003 GNDA.n291 175.546
R5004 GNDA.n5003 GNDA.n293 175.546
R5005 GNDA.n4999 GNDA.n293 175.546
R5006 GNDA.n4999 GNDA.n295 175.546
R5007 GNDA.n4995 GNDA.n295 175.546
R5008 GNDA.n4995 GNDA.n297 175.546
R5009 GNDA.n4991 GNDA.n297 175.546
R5010 GNDA.n4991 GNDA.n299 175.546
R5011 GNDA.n4987 GNDA.n299 175.546
R5012 GNDA.n58 GNDA.n54 175.546
R5013 GNDA.n5539 GNDA.n5538 175.546
R5014 GNDA.n5465 GNDA.n5464 175.546
R5015 GNDA.n5470 GNDA.n5469 175.546
R5016 GNDA.n5478 GNDA.n5477 175.546
R5017 GNDA.n409 GNDA.n408 175.546
R5018 GNDA.n406 GNDA.n372 175.546
R5019 GNDA.n402 GNDA.n400 175.546
R5020 GNDA.n398 GNDA.n380 175.546
R5021 GNDA.n394 GNDA.n392 175.546
R5022 GNDA.n4953 GNDA.n413 175.546
R5023 GNDA.n4949 GNDA.n413 175.546
R5024 GNDA.n4949 GNDA.n415 175.546
R5025 GNDA.n4945 GNDA.n415 175.546
R5026 GNDA.n4945 GNDA.n417 175.546
R5027 GNDA.n4941 GNDA.n417 175.546
R5028 GNDA.n4941 GNDA.n419 175.546
R5029 GNDA.n4937 GNDA.n419 175.546
R5030 GNDA.n4937 GNDA.n421 175.546
R5031 GNDA.n4933 GNDA.n421 175.546
R5032 GNDA.n4933 GNDA.n423 175.546
R5033 GNDA.n5552 GNDA.n24 175.546
R5034 GNDA.n40 GNDA.n25 175.546
R5035 GNDA.n31 GNDA.n30 175.546
R5036 GNDA.n5390 GNDA.n5389 175.546
R5037 GNDA.n5396 GNDA.n5395 175.546
R5038 GNDA.n4929 GNDA.n425 175.546
R5039 GNDA.n4925 GNDA.n425 175.546
R5040 GNDA.n4925 GNDA.n427 175.546
R5041 GNDA.n4921 GNDA.n427 175.546
R5042 GNDA.n4921 GNDA.n4918 175.546
R5043 GNDA.n4918 GNDA.n93 175.546
R5044 GNDA.n5373 GNDA.n93 175.546
R5045 GNDA.n5373 GNDA.n91 175.546
R5046 GNDA.n5378 GNDA.n91 175.546
R5047 GNDA.n5378 GNDA.n89 175.546
R5048 GNDA.n5382 GNDA.n89 175.546
R5049 GNDA.n157 GNDA.n100 173.881
R5050 GNDA.t186 GNDA.n101 172.876
R5051 GNDA.t186 GNDA.n111 172.615
R5052 GNDA.n5362 GNDA.n100 171.624
R5053 GNDA.n721 GNDA.n678 166.4
R5054 GNDA.n675 GNDA.n674 166.4
R5055 GNDA.n1587 GNDA.n1586 163.333
R5056 GNDA.n2034 GNDA.n2033 163.333
R5057 GNDA.n5277 GNDA.n5276 163.333
R5058 GNDA.n5062 GNDA.n5061 163.333
R5059 GNDA.n2202 GNDA.n2192 163.333
R5060 GNDA.n5203 GNDA.n5202 163.333
R5061 GNDA.n5482 GNDA.n5481 163.333
R5062 GNDA.n2078 GNDA.n1722 163.333
R5063 GNDA.n5400 GNDA.n5399 163.333
R5064 GNDA.n4971 GNDA.n355 157.601
R5065 GNDA.n1633 GNDA.n1632 150
R5066 GNDA.n1629 GNDA.n1628 150
R5067 GNDA.n1625 GNDA.n1624 150
R5068 GNDA.n1621 GNDA.n1620 150
R5069 GNDA.n1617 GNDA.n1616 150
R5070 GNDA.n1613 GNDA.n1612 150
R5071 GNDA.n1609 GNDA.n1608 150
R5072 GNDA.n1605 GNDA.n1604 150
R5073 GNDA.n2500 GNDA.n1596 150
R5074 GNDA.n2490 GNDA.n2489 150
R5075 GNDA.n2503 GNDA.n1567 150
R5076 GNDA.n1580 GNDA.n1568 150
R5077 GNDA.n1641 GNDA.n1640 150
R5078 GNDA.n1645 GNDA.n1644 150
R5079 GNDA.n1649 GNDA.n1648 150
R5080 GNDA.n1651 GNDA.n1595 150
R5081 GNDA.n1977 GNDA.n1975 150
R5082 GNDA.n1973 GNDA.n1941 150
R5083 GNDA.n1969 GNDA.n1967 150
R5084 GNDA.n1965 GNDA.n1943 150
R5085 GNDA.n1961 GNDA.n1959 150
R5086 GNDA.n1957 GNDA.n1945 150
R5087 GNDA.n1953 GNDA.n1952 150
R5088 GNDA.n1950 GNDA.n1948 150
R5089 GNDA.n2003 GNDA.n2001 150
R5090 GNDA.n2015 GNDA.n1908 150
R5091 GNDA.n2019 GNDA.n2017 150
R5092 GNDA.n2031 GNDA.n1902 150
R5093 GNDA.n1985 GNDA.n1983 150
R5094 GNDA.n1989 GNDA.n1937 150
R5095 GNDA.n1993 GNDA.n1991 150
R5096 GNDA.n1999 GNDA.n1935 150
R5097 GNDA.n5309 GNDA.n5308 150
R5098 GNDA.n5305 GNDA.n5304 150
R5099 GNDA.n5301 GNDA.n5300 150
R5100 GNDA.n5297 GNDA.n5296 150
R5101 GNDA.n5293 GNDA.n5292 150
R5102 GNDA.n5289 GNDA.n5288 150
R5103 GNDA.n5285 GNDA.n5284 150
R5104 GNDA.n5281 GNDA.n5280 150
R5105 GNDA.n5332 GNDA.n168 150
R5106 GNDA.n216 GNDA.n169 150
R5107 GNDA.n213 GNDA.n212 150
R5108 GNDA.n205 GNDA.n204 150
R5109 GNDA.n5317 GNDA.n5316 150
R5110 GNDA.n5321 GNDA.n5320 150
R5111 GNDA.n5325 GNDA.n5324 150
R5112 GNDA.n5329 GNDA.n5328 150
R5113 GNDA.n5094 GNDA.n5093 150
R5114 GNDA.n5090 GNDA.n5089 150
R5115 GNDA.n5086 GNDA.n5085 150
R5116 GNDA.n5082 GNDA.n5081 150
R5117 GNDA.n5078 GNDA.n5077 150
R5118 GNDA.n5074 GNDA.n5073 150
R5119 GNDA.n5070 GNDA.n5069 150
R5120 GNDA.n5066 GNDA.n5065 150
R5121 GNDA.n5117 GNDA.n5013 150
R5122 GNDA.n5039 GNDA.n5014 150
R5123 GNDA.n5047 GNDA.n5046 150
R5124 GNDA.n5054 GNDA.n5053 150
R5125 GNDA.n5102 GNDA.n5101 150
R5126 GNDA.n5106 GNDA.n5105 150
R5127 GNDA.n5110 GNDA.n5109 150
R5128 GNDA.n5114 GNDA.n5113 150
R5129 GNDA.n2242 GNDA.n2241 150
R5130 GNDA.n2238 GNDA.n2237 150
R5131 GNDA.n2234 GNDA.n2233 150
R5132 GNDA.n2230 GNDA.n2229 150
R5133 GNDA.n2226 GNDA.n2225 150
R5134 GNDA.n2222 GNDA.n2221 150
R5135 GNDA.n2218 GNDA.n2217 150
R5136 GNDA.n2214 GNDA.n2213 150
R5137 GNDA.n2291 GNDA.n2211 150
R5138 GNDA.n2280 GNDA.n2279 150
R5139 GNDA.n2273 GNDA.n2272 150
R5140 GNDA.n2294 GNDA.n2191 150
R5141 GNDA.n2250 GNDA.n2249 150
R5142 GNDA.n2254 GNDA.n2253 150
R5143 GNDA.n2258 GNDA.n2257 150
R5144 GNDA.n2260 GNDA.n2210 150
R5145 GNDA.n5235 GNDA.n5234 150
R5146 GNDA.n5231 GNDA.n5230 150
R5147 GNDA.n5227 GNDA.n5226 150
R5148 GNDA.n5223 GNDA.n5222 150
R5149 GNDA.n5219 GNDA.n5218 150
R5150 GNDA.n5215 GNDA.n5214 150
R5151 GNDA.n5211 GNDA.n5210 150
R5152 GNDA.n5207 GNDA.n5206 150
R5153 GNDA.n5264 GNDA.n5263 150
R5154 GNDA.n5256 GNDA.n5161 150
R5155 GNDA.n5188 GNDA.n5162 150
R5156 GNDA.n5195 GNDA.n5194 150
R5157 GNDA.n5253 GNDA.n5178 150
R5158 GNDA.n5249 GNDA.n5248 150
R5159 GNDA.n5245 GNDA.n5244 150
R5160 GNDA.n5241 GNDA.n5240 150
R5161 GNDA.n5514 GNDA.n5513 150
R5162 GNDA.n5510 GNDA.n5509 150
R5163 GNDA.n5506 GNDA.n5505 150
R5164 GNDA.n5502 GNDA.n5501 150
R5165 GNDA.n5498 GNDA.n5497 150
R5166 GNDA.n5494 GNDA.n5493 150
R5167 GNDA.n5490 GNDA.n5489 150
R5168 GNDA.n5486 GNDA.n5485 150
R5169 GNDA.n5543 GNDA.n5542 150
R5170 GNDA.n5535 GNDA.n64 150
R5171 GNDA.n5467 GNDA.n65 150
R5172 GNDA.n5474 GNDA.n5473 150
R5173 GNDA.n5532 GNDA.n81 150
R5174 GNDA.n5528 GNDA.n5527 150
R5175 GNDA.n5524 GNDA.n5523 150
R5176 GNDA.n5520 GNDA.n5519 150
R5177 GNDA.n1780 GNDA.n1740 150
R5178 GNDA.n1776 GNDA.n1774 150
R5179 GNDA.n1772 GNDA.n1742 150
R5180 GNDA.n1768 GNDA.n1766 150
R5181 GNDA.n1764 GNDA.n1744 150
R5182 GNDA.n1760 GNDA.n1759 150
R5183 GNDA.n1757 GNDA.n1747 150
R5184 GNDA.n1753 GNDA.n1752 150
R5185 GNDA.n1872 GNDA.n1729 150
R5186 GNDA.n1876 GNDA.n1874 150
R5187 GNDA.n2073 GNDA.n1725 150
R5188 GNDA.n2076 GNDA.n2075 150
R5189 GNDA.n1788 GNDA.n1738 150
R5190 GNDA.n1792 GNDA.n1790 150
R5191 GNDA.n1796 GNDA.n1736 150
R5192 GNDA.n1800 GNDA.n1798 150
R5193 GNDA.n5432 GNDA.n5431 150
R5194 GNDA.n5428 GNDA.n5427 150
R5195 GNDA.n5424 GNDA.n5423 150
R5196 GNDA.n5420 GNDA.n5419 150
R5197 GNDA.n5416 GNDA.n5415 150
R5198 GNDA.n5412 GNDA.n5411 150
R5199 GNDA.n5408 GNDA.n5407 150
R5200 GNDA.n5404 GNDA.n5403 150
R5201 GNDA.n5555 GNDA.n21 150
R5202 GNDA.n37 GNDA.n36 150
R5203 GNDA.n5558 GNDA.n2 150
R5204 GNDA.n5392 GNDA.n3 150
R5205 GNDA.n5440 GNDA.n5439 150
R5206 GNDA.n5444 GNDA.n5443 150
R5207 GNDA.n5448 GNDA.n5447 150
R5208 GNDA.n5450 GNDA.n20 150
R5209 GNDA.n4915 GNDA.n4914 148.017
R5210 GNDA.n4129 GNDA.n4128 148.017
R5211 GNDA.n4068 GNDA.n4067 148.017
R5212 GNDA.n3382 GNDA.n3381 148.017
R5213 GNDA.n2548 GNDA.n1443 136.145
R5214 GNDA.n2549 GNDA.n1442 136.145
R5215 GNDA.n2550 GNDA.n1441 136.145
R5216 GNDA.n2553 GNDA.n1438 136.145
R5217 GNDA.n2554 GNDA.n1437 136.145
R5218 GNDA.n2555 GNDA.n1436 136.145
R5219 GNDA.n2558 GNDA.n1433 136.145
R5220 GNDA.n2559 GNDA.n1432 136.145
R5221 GNDA.n2560 GNDA.n1431 136.145
R5222 GNDA.n2563 GNDA.n1428 136.145
R5223 GNDA.n2564 GNDA.n1427 136.145
R5224 GNDA.n2063 GNDA.n2056 134.268
R5225 GNDA.n2056 GNDA.n2054 134.268
R5226 GNDA.n1854 GNDA.n281 132.721
R5227 GNDA.n2546 GNDA.t237 130.001
R5228 GNDA.n2472 GNDA.t192 130.001
R5229 GNDA.n1659 GNDA.t250 130.001
R5230 GNDA.n1915 GNDA.t223 130.001
R5231 GNDA.n1913 GNDA.t189 130.001
R5232 GNDA.n1865 GNDA.t276 130.001
R5233 GNDA.n1862 GNDA.t234 130.001
R5234 GNDA.n1425 GNDA.t184 130
R5235 GNDA.n5371 GNDA.t186 127.219
R5236 GNDA.t186 GNDA.n108 127.219
R5237 GNDA.t186 GNDA.n1562 127.219
R5238 GNDA.n2479 GNDA.n2478 124.832
R5239 GNDA.n2476 GNDA.n2475 124.832
R5240 GNDA.n1912 GNDA.n1708 124.832
R5241 GNDA.n1718 GNDA.n1713 124.832
R5242 GNDA.n5458 GNDA.n83 124.832
R5243 GNDA.n327 GNDA.n55 124.832
R5244 GNDA.n2385 GNDA.n2384 124.832
R5245 GNDA.n2382 GNDA.n2138 124.832
R5246 GNDA.n5342 GNDA.n5341 124.832
R5247 GNDA.n5179 GNDA.n159 124.832
R5248 GNDA.n325 GNDA.n85 124.832
R5249 GNDA.n5456 GNDA.n86 124.832
R5250 GNDA.n4891 GNDA.n4889 121.251
R5251 GNDA.n1002 GNDA.n1000 121.251
R5252 GNDA.n4899 GNDA.n4898 121.136
R5253 GNDA.n4897 GNDA.n4896 121.136
R5254 GNDA.n4895 GNDA.n4894 121.136
R5255 GNDA.n4893 GNDA.n4892 121.136
R5256 GNDA.n4891 GNDA.n4890 121.136
R5257 GNDA.n1002 GNDA.n1001 121.136
R5258 GNDA.n1004 GNDA.n1003 121.136
R5259 GNDA.n1006 GNDA.n1005 121.136
R5260 GNDA.n1008 GNDA.n1007 121.136
R5261 GNDA.n1010 GNDA.n1009 121.136
R5262 GNDA.n1463 GNDA.t52 111.799
R5263 GNDA.n1462 GNDA.t108 111.331
R5264 GNDA.n2572 GNDA.t91 111.206
R5265 GNDA.n2572 GNDA.t20 111.076
R5266 GNDA.n4988 GNDA.n300 105.719
R5267 GNDA.n4956 GNDA.n4955 105.719
R5268 GNDA.n4982 GNDA.n300 103.457
R5269 GNDA.n4955 GNDA.n4954 103.457
R5270 GNDA.n2508 GNDA.n1560 101.718
R5271 GNDA.n2059 GNDA.n1882 101.718
R5272 GNDA.n2065 GNDA.n1884 101.718
R5273 GNDA.n2519 GNDA.n1558 101.718
R5274 GNDA.t186 GNDA.n104 47.6748
R5275 GNDA.t63 GNDA.n671 97.7783
R5276 GNDA.n4129 GNDA.n4126 95.3634
R5277 GNDA.n4124 GNDA.n4122 94.2862
R5278 GNDA.n4047 GNDA.n4046 92.8005
R5279 GNDA.n4058 GNDA.n4057 92.8005
R5280 GNDA.n2515 GNDA.n1557 91.069
R5281 GNDA.n2510 GNDA.n1557 91.069
R5282 GNDA.n2512 GNDA.n1556 91.069
R5283 GNDA.n2513 GNDA.n2512 91.069
R5284 GNDA.n2063 GNDA.n2058 91.069
R5285 GNDA.n2061 GNDA.n2054 91.069
R5286 GNDA.n1861 GNDA.n1733 90.1439
R5287 GNDA.n2069 GNDA.n2068 90.1439
R5288 GNDA.n2007 GNDA.n1911 90.1439
R5289 GNDA.n2495 GNDA.n2494 90.1439
R5290 GNDA.n1575 GNDA.n1444 90.1439
R5291 GNDA.n2544 GNDA.n1445 90.1439
R5292 GNDA.n741 GNDA.n643 89.6005
R5293 GNDA.n741 GNDA.n740 89.6005
R5294 GNDA.n1866 GNDA.n1864 87.1391
R5295 GNDA.t186 GNDA.n1661 87.1391
R5296 GNDA.n1928 GNDA.n1918 84.306
R5297 GNDA.n2043 GNDA.n1897 84.306
R5298 GNDA.t38 GNDA.n1867 83.1328
R5299 GNDA.t131 GNDA.n2067 82.1312
R5300 GNDA.n2010 GNDA.t277 82.1312
R5301 GNDA.n2496 GNDA.t36 82.1312
R5302 GNDA.n1455 GNDA.t146 78.5658
R5303 GNDA.n2082 GNDA.t24 78.1248
R5304 GNDA.n2024 GNDA.t129 78.1248
R5305 GNDA.t93 GNDA.n1559 78.1248
R5306 GNDA.t186 GNDA.n100 76.3879
R5307 GNDA.n2443 GNDA.n2442 76.3222
R5308 GNDA.n2453 GNDA.n2452 76.3222
R5309 GNDA.n2456 GNDA.n2455 76.3222
R5310 GNDA.n2464 GNDA.n2463 76.3222
R5311 GNDA.n2467 GNDA.n2466 76.3222
R5312 GNDA.n2440 GNDA.n2439 76.3222
R5313 GNDA.n2435 GNDA.n2391 76.3222
R5314 GNDA.n2433 GNDA.n2432 76.3222
R5315 GNDA.n2428 GNDA.n2394 76.3222
R5316 GNDA.n2426 GNDA.n2425 76.3222
R5317 GNDA.n2421 GNDA.n2397 76.3222
R5318 GNDA.n2446 GNDA.n1671 76.3222
R5319 GNDA.n2450 GNDA.n1672 76.3222
R5320 GNDA.n2458 GNDA.n1673 76.3222
R5321 GNDA.n2461 GNDA.n1674 76.3222
R5322 GNDA.n2470 GNDA.n2469 76.3222
R5323 GNDA.n2476 GNDA.n1657 76.3222
R5324 GNDA.n2111 GNDA.n1687 76.3222
R5325 GNDA.n2118 GNDA.n2117 76.3222
R5326 GNDA.n2119 GNDA.n1685 76.3222
R5327 GNDA.n2126 GNDA.n2125 76.3222
R5328 GNDA.n2130 GNDA.n1683 76.3222
R5329 GNDA.n2134 GNDA.n2132 76.3222
R5330 GNDA.n2110 GNDA.n1689 76.3222
R5331 GNDA.n2105 GNDA.n1694 76.3222
R5332 GNDA.n2101 GNDA.n2100 76.3222
R5333 GNDA.n2094 GNDA.n1700 76.3222
R5334 GNDA.n2093 GNDA.n2092 76.3222
R5335 GNDA.n1832 GNDA.n286 76.3222
R5336 GNDA.n1836 GNDA.n285 76.3222
R5337 GNDA.n1840 GNDA.n284 76.3222
R5338 GNDA.n1844 GNDA.n283 76.3222
R5339 GNDA.n1848 GNDA.n282 76.3222
R5340 GNDA.n1852 GNDA.n281 76.3222
R5341 GNDA.n1830 GNDA.n1829 76.3222
R5342 GNDA.n1825 GNDA.n1805 76.3222
R5343 GNDA.n1823 GNDA.n1822 76.3222
R5344 GNDA.n1818 GNDA.n1808 76.3222
R5345 GNDA.n1816 GNDA.n1815 76.3222
R5346 GNDA.n1811 GNDA.n1810 76.3222
R5347 GNDA.n1691 GNDA.n1690 76.3222
R5348 GNDA.n1696 GNDA.n1695 76.3222
R5349 GNDA.n1701 GNDA.n1698 76.3222
R5350 GNDA.n1704 GNDA.n1703 76.3222
R5351 GNDA.n1709 GNDA.n1706 76.3222
R5352 GNDA.n1712 GNDA.n1711 76.3222
R5353 GNDA.n370 GNDA.n369 76.3222
R5354 GNDA.n375 GNDA.n374 76.3222
R5355 GNDA.n378 GNDA.n377 76.3222
R5356 GNDA.n383 GNDA.n382 76.3222
R5357 GNDA.n386 GNDA.n385 76.3222
R5358 GNDA.n387 GNDA.n83 76.3222
R5359 GNDA.n349 GNDA.n348 76.3222
R5360 GNDA.n342 GNDA.n304 76.3222
R5361 GNDA.n341 GNDA.n340 76.3222
R5362 GNDA.n334 GNDA.n311 76.3222
R5363 GNDA.n333 GNDA.n332 76.3222
R5364 GNDA.n326 GNDA.n319 76.3222
R5365 GNDA.n2139 GNDA.n195 76.3222
R5366 GNDA.n2288 GNDA.n194 76.3222
R5367 GNDA.n2283 GNDA.n193 76.3222
R5368 GNDA.n2276 GNDA.n192 76.3222
R5369 GNDA.n2269 GNDA.n191 76.3222
R5370 GNDA.n2298 GNDA.n190 76.3222
R5371 GNDA.n2352 GNDA.n2351 76.3222
R5372 GNDA.n2362 GNDA.n2361 76.3222
R5373 GNDA.n2365 GNDA.n2364 76.3222
R5374 GNDA.n2374 GNDA.n2373 76.3222
R5375 GNDA.n2377 GNDA.n2376 76.3222
R5376 GNDA.n2347 GNDA.n112 76.3222
R5377 GNDA.n2343 GNDA.n113 76.3222
R5378 GNDA.n2339 GNDA.n114 76.3222
R5379 GNDA.n2335 GNDA.n115 76.3222
R5380 GNDA.n2331 GNDA.n116 76.3222
R5381 GNDA.n2327 GNDA.n117 76.3222
R5382 GNDA.n2355 GNDA.n2150 76.3222
R5383 GNDA.n2359 GNDA.n2357 76.3222
R5384 GNDA.n2367 GNDA.n2146 76.3222
R5385 GNDA.n2371 GNDA.n2369 76.3222
R5386 GNDA.n2379 GNDA.n2142 76.3222
R5387 GNDA.n2382 GNDA.n2381 76.3222
R5388 GNDA.n5340 GNDA.n163 76.3222
R5389 GNDA.n5335 GNDA.n166 76.3222
R5390 GNDA.n220 GNDA.n219 76.3222
R5391 GNDA.n201 GNDA.n197 76.3222
R5392 GNDA.n208 GNDA.n196 76.3222
R5393 GNDA.n5273 GNDA.n5272 76.3222
R5394 GNDA.n5364 GNDA.n5363 76.3222
R5395 GNDA.n5361 GNDA.n5360 76.3222
R5396 GNDA.n5356 GNDA.n140 76.3222
R5397 GNDA.n5353 GNDA.n139 76.3222
R5398 GNDA.n5349 GNDA.n138 76.3222
R5399 GNDA.n5345 GNDA.n137 76.3222
R5400 GNDA.n2153 GNDA.n118 76.3222
R5401 GNDA.n2157 GNDA.n119 76.3222
R5402 GNDA.n2161 GNDA.n120 76.3222
R5403 GNDA.n2165 GNDA.n121 76.3222
R5404 GNDA.n2169 GNDA.n122 76.3222
R5405 GNDA.n2173 GNDA.n123 76.3222
R5406 GNDA.n152 GNDA.n151 76.3222
R5407 GNDA.n153 GNDA.n143 76.3222
R5408 GNDA.n154 GNDA.n145 76.3222
R5409 GNDA.n155 GNDA.n147 76.3222
R5410 GNDA.n156 GNDA.n149 76.3222
R5411 GNDA.n159 GNDA.n158 76.3222
R5412 GNDA.n5270 GNDA.n5269 76.3222
R5413 GNDA.n5155 GNDA.n225 76.3222
R5414 GNDA.n5259 GNDA.n224 76.3222
R5415 GNDA.n5186 GNDA.n223 76.3222
R5416 GNDA.n5190 GNDA.n222 76.3222
R5417 GNDA.n5199 GNDA.n221 76.3222
R5418 GNDA.n261 GNDA.n235 76.3222
R5419 GNDA.n265 GNDA.n236 76.3222
R5420 GNDA.n269 GNDA.n237 76.3222
R5421 GNDA.n273 GNDA.n238 76.3222
R5422 GNDA.n279 GNDA.n278 76.3222
R5423 GNDA.n257 GNDA.n124 76.3222
R5424 GNDA.n253 GNDA.n125 76.3222
R5425 GNDA.n249 GNDA.n126 76.3222
R5426 GNDA.n245 GNDA.n127 76.3222
R5427 GNDA.n241 GNDA.n128 76.3222
R5428 GNDA.n5369 GNDA.n5368 76.3222
R5429 GNDA.n306 GNDA.n305 76.3222
R5430 GNDA.n309 GNDA.n308 76.3222
R5431 GNDA.n314 GNDA.n313 76.3222
R5432 GNDA.n317 GNDA.n316 76.3222
R5433 GNDA.n322 GNDA.n321 76.3222
R5434 GNDA.n325 GNDA.n324 76.3222
R5435 GNDA.n5121 GNDA.n48 76.3222
R5436 GNDA.n5036 GNDA.n47 76.3222
R5437 GNDA.n5042 GNDA.n46 76.3222
R5438 GNDA.n5050 GNDA.n45 76.3222
R5439 GNDA.n5057 GNDA.n44 76.3222
R5440 GNDA.n5031 GNDA.n43 76.3222
R5441 GNDA.n5149 GNDA.n5148 76.3222
R5442 GNDA.n5143 GNDA.n230 76.3222
R5443 GNDA.n5140 GNDA.n231 76.3222
R5444 GNDA.n5136 GNDA.n232 76.3222
R5445 GNDA.n5132 GNDA.n233 76.3222
R5446 GNDA.n5369 GNDA.n129 76.3222
R5447 GNDA.n244 GNDA.n128 76.3222
R5448 GNDA.n248 GNDA.n127 76.3222
R5449 GNDA.n252 GNDA.n126 76.3222
R5450 GNDA.n256 GNDA.n125 76.3222
R5451 GNDA.n260 GNDA.n124 76.3222
R5452 GNDA.n2170 GNDA.n123 76.3222
R5453 GNDA.n2166 GNDA.n122 76.3222
R5454 GNDA.n2162 GNDA.n121 76.3222
R5455 GNDA.n2158 GNDA.n120 76.3222
R5456 GNDA.n2154 GNDA.n119 76.3222
R5457 GNDA.n135 GNDA.n118 76.3222
R5458 GNDA.n2330 GNDA.n117 76.3222
R5459 GNDA.n2334 GNDA.n116 76.3222
R5460 GNDA.n2338 GNDA.n115 76.3222
R5461 GNDA.n2342 GNDA.n114 76.3222
R5462 GNDA.n2346 GNDA.n113 76.3222
R5463 GNDA.n2350 GNDA.n112 76.3222
R5464 GNDA.n5549 GNDA.n54 76.3222
R5465 GNDA.n5539 GNDA.n53 76.3222
R5466 GNDA.n5464 GNDA.n52 76.3222
R5467 GNDA.n5470 GNDA.n51 76.3222
R5468 GNDA.n5477 GNDA.n50 76.3222
R5469 GNDA.n5459 GNDA.n49 76.3222
R5470 GNDA.n5549 GNDA.n5548 76.3222
R5471 GNDA.n58 GNDA.n53 76.3222
R5472 GNDA.n5538 GNDA.n52 76.3222
R5473 GNDA.n5465 GNDA.n51 76.3222
R5474 GNDA.n5469 GNDA.n50 76.3222
R5475 GNDA.n5478 GNDA.n49 76.3222
R5476 GNDA.n5125 GNDA.n48 76.3222
R5477 GNDA.n5120 GNDA.n47 76.3222
R5478 GNDA.n5037 GNDA.n46 76.3222
R5479 GNDA.n5043 GNDA.n45 76.3222
R5480 GNDA.n5049 GNDA.n44 76.3222
R5481 GNDA.n5058 GNDA.n43 76.3222
R5482 GNDA.n324 GNDA.n323 76.3222
R5483 GNDA.n321 GNDA.n320 76.3222
R5484 GNDA.n316 GNDA.n315 76.3222
R5485 GNDA.n313 GNDA.n312 76.3222
R5486 GNDA.n308 GNDA.n307 76.3222
R5487 GNDA.n305 GNDA.n301 76.3222
R5488 GNDA.n348 GNDA.n347 76.3222
R5489 GNDA.n343 GNDA.n342 76.3222
R5490 GNDA.n340 GNDA.n339 76.3222
R5491 GNDA.n335 GNDA.n334 76.3222
R5492 GNDA.n332 GNDA.n331 76.3222
R5493 GNDA.n327 GNDA.n326 76.3222
R5494 GNDA.n158 GNDA.n150 76.3222
R5495 GNDA.n156 GNDA.n148 76.3222
R5496 GNDA.n155 GNDA.n146 76.3222
R5497 GNDA.n154 GNDA.n144 76.3222
R5498 GNDA.n153 GNDA.n142 76.3222
R5499 GNDA.n152 GNDA.n130 76.3222
R5500 GNDA.n5363 GNDA.n136 76.3222
R5501 GNDA.n5361 GNDA.n141 76.3222
R5502 GNDA.n5354 GNDA.n140 76.3222
R5503 GNDA.n5350 GNDA.n139 76.3222
R5504 GNDA.n5346 GNDA.n138 76.3222
R5505 GNDA.n5342 GNDA.n137 76.3222
R5506 GNDA.n1713 GNDA.n1712 76.3222
R5507 GNDA.n1710 GNDA.n1709 76.3222
R5508 GNDA.n1705 GNDA.n1704 76.3222
R5509 GNDA.n1702 GNDA.n1701 76.3222
R5510 GNDA.n1697 GNDA.n1696 76.3222
R5511 GNDA.n1692 GNDA.n1691 76.3222
R5512 GNDA.n2107 GNDA.n1689 76.3222
R5513 GNDA.n2102 GNDA.n1694 76.3222
R5514 GNDA.n2100 GNDA.n2099 76.3222
R5515 GNDA.n2095 GNDA.n2094 76.3222
R5516 GNDA.n2092 GNDA.n2091 76.3222
R5517 GNDA.n1810 GNDA.n1809 76.3222
R5518 GNDA.n1817 GNDA.n1816 76.3222
R5519 GNDA.n1808 GNDA.n1806 76.3222
R5520 GNDA.n1824 GNDA.n1823 76.3222
R5521 GNDA.n1805 GNDA.n1803 76.3222
R5522 GNDA.n1831 GNDA.n1830 76.3222
R5523 GNDA.n2132 GNDA.n2131 76.3222
R5524 GNDA.n2127 GNDA.n1683 76.3222
R5525 GNDA.n2125 GNDA.n2124 76.3222
R5526 GNDA.n2120 GNDA.n2119 76.3222
R5527 GNDA.n2117 GNDA.n2116 76.3222
R5528 GNDA.n2112 GNDA.n2111 76.3222
R5529 GNDA.n2397 GNDA.n2395 76.3222
R5530 GNDA.n2427 GNDA.n2426 76.3222
R5531 GNDA.n2394 GNDA.n2392 76.3222
R5532 GNDA.n2434 GNDA.n2433 76.3222
R5533 GNDA.n2391 GNDA.n2389 76.3222
R5534 GNDA.n2441 GNDA.n2440 76.3222
R5535 GNDA.n5270 GNDA.n226 76.3222
R5536 GNDA.n5260 GNDA.n225 76.3222
R5537 GNDA.n5185 GNDA.n224 76.3222
R5538 GNDA.n5191 GNDA.n223 76.3222
R5539 GNDA.n5198 GNDA.n222 76.3222
R5540 GNDA.n5180 GNDA.n221 76.3222
R5541 GNDA.n5336 GNDA.n163 76.3222
R5542 GNDA.n199 GNDA.n166 76.3222
R5543 GNDA.n220 GNDA.n198 76.3222
R5544 GNDA.n209 GNDA.n197 76.3222
R5545 GNDA.n196 GNDA.n188 76.3222
R5546 GNDA.n5272 GNDA.n189 76.3222
R5547 GNDA.n2287 GNDA.n195 76.3222
R5548 GNDA.n2284 GNDA.n194 76.3222
R5549 GNDA.n2277 GNDA.n193 76.3222
R5550 GNDA.n2270 GNDA.n192 76.3222
R5551 GNDA.n2297 GNDA.n191 76.3222
R5552 GNDA.n2302 GNDA.n190 76.3222
R5553 GNDA.n412 GNDA.n368 76.3222
R5554 GNDA.n408 GNDA.n407 76.3222
R5555 GNDA.n401 GNDA.n372 76.3222
R5556 GNDA.n400 GNDA.n399 76.3222
R5557 GNDA.n393 GNDA.n380 76.3222
R5558 GNDA.n392 GNDA.n391 76.3222
R5559 GNDA.n42 GNDA.n24 76.3222
R5560 GNDA.n5551 GNDA.n25 76.3222
R5561 GNDA.n41 GNDA.n31 76.3222
R5562 GNDA.n5389 GNDA.n29 76.3222
R5563 GNDA.n5395 GNDA.n28 76.3222
R5564 GNDA.n5385 GNDA.n27 76.3222
R5565 GNDA.n5455 GNDA.n42 76.3222
R5566 GNDA.n5552 GNDA.n5551 76.3222
R5567 GNDA.n41 GNDA.n40 76.3222
R5568 GNDA.n30 GNDA.n29 76.3222
R5569 GNDA.n5390 GNDA.n28 76.3222
R5570 GNDA.n5396 GNDA.n27 76.3222
R5571 GNDA.n388 GNDA.n387 76.3222
R5572 GNDA.n385 GNDA.n384 76.3222
R5573 GNDA.n382 GNDA.n381 76.3222
R5574 GNDA.n377 GNDA.n376 76.3222
R5575 GNDA.n374 GNDA.n373 76.3222
R5576 GNDA.n369 GNDA.n366 76.3222
R5577 GNDA.n409 GNDA.n368 76.3222
R5578 GNDA.n407 GNDA.n406 76.3222
R5579 GNDA.n402 GNDA.n401 76.3222
R5580 GNDA.n399 GNDA.n398 76.3222
R5581 GNDA.n394 GNDA.n393 76.3222
R5582 GNDA.n391 GNDA.n86 76.3222
R5583 GNDA.n2381 GNDA.n2380 76.3222
R5584 GNDA.n2370 GNDA.n2142 76.3222
R5585 GNDA.n2369 GNDA.n2368 76.3222
R5586 GNDA.n2358 GNDA.n2146 76.3222
R5587 GNDA.n2357 GNDA.n2356 76.3222
R5588 GNDA.n2172 GNDA.n2150 76.3222
R5589 GNDA.n2353 GNDA.n2352 76.3222
R5590 GNDA.n2363 GNDA.n2362 76.3222
R5591 GNDA.n2364 GNDA.n2144 76.3222
R5592 GNDA.n2375 GNDA.n2374 76.3222
R5593 GNDA.n2376 GNDA.n2140 76.3222
R5594 GNDA.n1676 GNDA.n1657 76.3222
R5595 GNDA.n2470 GNDA.n1675 76.3222
R5596 GNDA.n2459 GNDA.n1674 76.3222
R5597 GNDA.n2449 GNDA.n1673 76.3222
R5598 GNDA.n2447 GNDA.n1672 76.3222
R5599 GNDA.n2133 GNDA.n1671 76.3222
R5600 GNDA.n2444 GNDA.n2443 76.3222
R5601 GNDA.n2454 GNDA.n2453 76.3222
R5602 GNDA.n2455 GNDA.n1678 76.3222
R5603 GNDA.n2465 GNDA.n2464 76.3222
R5604 GNDA.n2466 GNDA.n1601 76.3222
R5605 GNDA.n1835 GNDA.n286 76.3222
R5606 GNDA.n1839 GNDA.n285 76.3222
R5607 GNDA.n1843 GNDA.n284 76.3222
R5608 GNDA.n1847 GNDA.n283 76.3222
R5609 GNDA.n1851 GNDA.n282 76.3222
R5610 GNDA.n264 GNDA.n235 76.3222
R5611 GNDA.n268 GNDA.n236 76.3222
R5612 GNDA.n272 GNDA.n237 76.3222
R5613 GNDA.n240 GNDA.n238 76.3222
R5614 GNDA.n279 GNDA.n239 76.3222
R5615 GNDA.n5149 GNDA.n288 76.3222
R5616 GNDA.n5141 GNDA.n230 76.3222
R5617 GNDA.n5137 GNDA.n231 76.3222
R5618 GNDA.n5133 GNDA.n232 76.3222
R5619 GNDA.n5129 GNDA.n233 76.3222
R5620 GNDA.n1620 GNDA.n1582 74.5978
R5621 GNDA.n1617 GNDA.n1582 74.5978
R5622 GNDA.n1960 GNDA.n1943 74.5978
R5623 GNDA.n1961 GNDA.n1960 74.5978
R5624 GNDA.n5296 GNDA.n175 74.5978
R5625 GNDA.n5293 GNDA.n175 74.5978
R5626 GNDA.n5081 GNDA.n5020 74.5978
R5627 GNDA.n5078 GNDA.n5020 74.5978
R5628 GNDA.n2229 GNDA.n2198 74.5978
R5629 GNDA.n2226 GNDA.n2198 74.5978
R5630 GNDA.n5222 GNDA.n5167 74.5978
R5631 GNDA.n5219 GNDA.n5167 74.5978
R5632 GNDA.n5501 GNDA.n70 74.5978
R5633 GNDA.n5498 GNDA.n70 74.5978
R5634 GNDA.n1766 GNDA.n1765 74.5978
R5635 GNDA.n1765 GNDA.n1764 74.5978
R5636 GNDA.n5419 GNDA.n9 74.5978
R5637 GNDA.n5416 GNDA.n9 74.5978
R5638 GNDA.n2474 GNDA.n1660 74.1184
R5639 GNDA.t279 GNDA.t13 72.3293
R5640 GNDA.n2085 GNDA.t110 72.1152
R5641 GNDA.n2025 GNDA.t248 72.1152
R5642 GNDA.t236 GNDA.n1574 72.1152
R5643 GNDA.t281 GNDA.t18 70.6072
R5644 GNDA.t186 GNDA.t84 70.1899
R5645 GNDA.n4972 GNDA.n4971 69.4466
R5646 GNDA.n2501 GNDA.n2500 69.3109
R5647 GNDA.n2501 GNDA.n1595 69.3109
R5648 GNDA.n2001 GNDA.n2000 69.3109
R5649 GNDA.n2000 GNDA.n1999 69.3109
R5650 GNDA.n5330 GNDA.n168 69.3109
R5651 GNDA.n5330 GNDA.n5329 69.3109
R5652 GNDA.n5115 GNDA.n5013 69.3109
R5653 GNDA.n5115 GNDA.n5114 69.3109
R5654 GNDA.n2292 GNDA.n2291 69.3109
R5655 GNDA.n2292 GNDA.n2210 69.3109
R5656 GNDA.n5264 GNDA.n5157 69.3109
R5657 GNDA.n5240 GNDA.n5157 69.3109
R5658 GNDA.n5543 GNDA.n60 69.3109
R5659 GNDA.n5519 GNDA.n60 69.3109
R5660 GNDA.n1799 GNDA.n1729 69.3109
R5661 GNDA.n1800 GNDA.n1799 69.3109
R5662 GNDA.n5556 GNDA.n5555 69.3109
R5663 GNDA.n5556 GNDA.n20 69.3109
R5664 GNDA.n2481 GNDA.t191 68.1089
R5665 GNDA.n2474 GNDA.n2473 66.1057
R5666 GNDA.t242 GNDA.n1594 65.8183
R5667 GNDA.t242 GNDA.n1593 65.8183
R5668 GNDA.t242 GNDA.n1592 65.8183
R5669 GNDA.t242 GNDA.n1591 65.8183
R5670 GNDA.t242 GNDA.n1572 65.8183
R5671 GNDA.t242 GNDA.n1589 65.8183
R5672 GNDA.t242 GNDA.n1570 65.8183
R5673 GNDA.t242 GNDA.n1590 65.8183
R5674 GNDA.t242 GNDA.n1588 65.8183
R5675 GNDA.t242 GNDA.n1585 65.8183
R5676 GNDA.t242 GNDA.n1584 65.8183
R5677 GNDA.t242 GNDA.n1583 65.8183
R5678 GNDA.t242 GNDA.n1581 65.8183
R5679 GNDA.n2502 GNDA.t242 65.8183
R5680 GNDA.t242 GNDA.n1571 65.8183
R5681 GNDA.t242 GNDA.n1569 65.8183
R5682 GNDA.n1982 GNDA.t217 65.8183
R5683 GNDA.n1984 GNDA.t217 65.8183
R5684 GNDA.n1990 GNDA.t217 65.8183
R5685 GNDA.n1992 GNDA.t217 65.8183
R5686 GNDA.n1966 GNDA.t217 65.8183
R5687 GNDA.n1968 GNDA.t217 65.8183
R5688 GNDA.n1974 GNDA.t217 65.8183
R5689 GNDA.n1976 GNDA.t217 65.8183
R5690 GNDA.t217 GNDA.n1901 65.8183
R5691 GNDA.n1951 GNDA.t217 65.8183
R5692 GNDA.n1947 GNDA.t217 65.8183
R5693 GNDA.n1958 GNDA.t217 65.8183
R5694 GNDA.n2032 GNDA.t217 65.8183
R5695 GNDA.n2018 GNDA.t217 65.8183
R5696 GNDA.n2016 GNDA.t217 65.8183
R5697 GNDA.n2002 GNDA.t217 65.8183
R5698 GNDA.t185 GNDA.n185 65.8183
R5699 GNDA.t185 GNDA.n184 65.8183
R5700 GNDA.t185 GNDA.n183 65.8183
R5701 GNDA.t185 GNDA.n182 65.8183
R5702 GNDA.t185 GNDA.n173 65.8183
R5703 GNDA.t185 GNDA.n180 65.8183
R5704 GNDA.t185 GNDA.n170 65.8183
R5705 GNDA.t185 GNDA.n181 65.8183
R5706 GNDA.t185 GNDA.n179 65.8183
R5707 GNDA.t185 GNDA.n178 65.8183
R5708 GNDA.t185 GNDA.n177 65.8183
R5709 GNDA.t185 GNDA.n176 65.8183
R5710 GNDA.t185 GNDA.n174 65.8183
R5711 GNDA.t185 GNDA.n172 65.8183
R5712 GNDA.t185 GNDA.n171 65.8183
R5713 GNDA.n5331 GNDA.t185 65.8183
R5714 GNDA.t243 GNDA.n5030 65.8183
R5715 GNDA.t243 GNDA.n5029 65.8183
R5716 GNDA.t243 GNDA.n5028 65.8183
R5717 GNDA.t243 GNDA.n5027 65.8183
R5718 GNDA.t243 GNDA.n5018 65.8183
R5719 GNDA.t243 GNDA.n5025 65.8183
R5720 GNDA.t243 GNDA.n5015 65.8183
R5721 GNDA.t243 GNDA.n5026 65.8183
R5722 GNDA.t243 GNDA.n5024 65.8183
R5723 GNDA.t243 GNDA.n5023 65.8183
R5724 GNDA.t243 GNDA.n5022 65.8183
R5725 GNDA.t243 GNDA.n5021 65.8183
R5726 GNDA.t224 GNDA.n2209 65.8183
R5727 GNDA.t224 GNDA.n2208 65.8183
R5728 GNDA.t224 GNDA.n2207 65.8183
R5729 GNDA.t224 GNDA.n2206 65.8183
R5730 GNDA.t224 GNDA.n2197 65.8183
R5731 GNDA.t224 GNDA.n2204 65.8183
R5732 GNDA.t224 GNDA.n2194 65.8183
R5733 GNDA.t224 GNDA.n2205 65.8183
R5734 GNDA.t224 GNDA.n2203 65.8183
R5735 GNDA.t224 GNDA.n2201 65.8183
R5736 GNDA.t224 GNDA.n2200 65.8183
R5737 GNDA.t224 GNDA.n2199 65.8183
R5738 GNDA.n2293 GNDA.t224 65.8183
R5739 GNDA.t224 GNDA.n2196 65.8183
R5740 GNDA.t224 GNDA.n2195 65.8183
R5741 GNDA.t224 GNDA.n2193 65.8183
R5742 GNDA.t251 GNDA.n5254 65.8183
R5743 GNDA.t251 GNDA.n5176 65.8183
R5744 GNDA.t251 GNDA.n5175 65.8183
R5745 GNDA.t251 GNDA.n5174 65.8183
R5746 GNDA.t251 GNDA.n5165 65.8183
R5747 GNDA.t251 GNDA.n5172 65.8183
R5748 GNDA.t251 GNDA.n5163 65.8183
R5749 GNDA.t251 GNDA.n5173 65.8183
R5750 GNDA.t251 GNDA.n5171 65.8183
R5751 GNDA.t251 GNDA.n5170 65.8183
R5752 GNDA.t251 GNDA.n5169 65.8183
R5753 GNDA.t251 GNDA.n5168 65.8183
R5754 GNDA.t251 GNDA.n5166 65.8183
R5755 GNDA.t251 GNDA.n5164 65.8183
R5756 GNDA.n5255 GNDA.t251 65.8183
R5757 GNDA.t251 GNDA.n5158 65.8183
R5758 GNDA.t210 GNDA.n5533 65.8183
R5759 GNDA.t210 GNDA.n79 65.8183
R5760 GNDA.t210 GNDA.n78 65.8183
R5761 GNDA.t210 GNDA.n77 65.8183
R5762 GNDA.t210 GNDA.n68 65.8183
R5763 GNDA.t210 GNDA.n75 65.8183
R5764 GNDA.t210 GNDA.n66 65.8183
R5765 GNDA.t210 GNDA.n76 65.8183
R5766 GNDA.t210 GNDA.n74 65.8183
R5767 GNDA.t210 GNDA.n73 65.8183
R5768 GNDA.t210 GNDA.n72 65.8183
R5769 GNDA.t210 GNDA.n71 65.8183
R5770 GNDA.t210 GNDA.n69 65.8183
R5771 GNDA.t210 GNDA.n67 65.8183
R5772 GNDA.n5534 GNDA.t210 65.8183
R5773 GNDA.t210 GNDA.n61 65.8183
R5774 GNDA.t243 GNDA.n5019 65.8183
R5775 GNDA.t243 GNDA.n5017 65.8183
R5776 GNDA.t243 GNDA.n5016 65.8183
R5777 GNDA.n5116 GNDA.t243 65.8183
R5778 GNDA.n1783 GNDA.t258 65.8183
R5779 GNDA.n1789 GNDA.t258 65.8183
R5780 GNDA.n1791 GNDA.t258 65.8183
R5781 GNDA.n1797 GNDA.t258 65.8183
R5782 GNDA.n1767 GNDA.t258 65.8183
R5783 GNDA.n1773 GNDA.t258 65.8183
R5784 GNDA.n1775 GNDA.t258 65.8183
R5785 GNDA.n1781 GNDA.t258 65.8183
R5786 GNDA.n1751 GNDA.t258 65.8183
R5787 GNDA.n1750 GNDA.t258 65.8183
R5788 GNDA.n1758 GNDA.t258 65.8183
R5789 GNDA.n1746 GNDA.t258 65.8183
R5790 GNDA.n2077 GNDA.t258 65.8183
R5791 GNDA.n2074 GNDA.t258 65.8183
R5792 GNDA.n1875 GNDA.t258 65.8183
R5793 GNDA.n1873 GNDA.t258 65.8183
R5794 GNDA.t228 GNDA.n19 65.8183
R5795 GNDA.t228 GNDA.n18 65.8183
R5796 GNDA.t228 GNDA.n17 65.8183
R5797 GNDA.t228 GNDA.n16 65.8183
R5798 GNDA.t228 GNDA.n7 65.8183
R5799 GNDA.t228 GNDA.n14 65.8183
R5800 GNDA.t228 GNDA.n5 65.8183
R5801 GNDA.t228 GNDA.n15 65.8183
R5802 GNDA.t228 GNDA.n13 65.8183
R5803 GNDA.t228 GNDA.n12 65.8183
R5804 GNDA.t228 GNDA.n11 65.8183
R5805 GNDA.t228 GNDA.n10 65.8183
R5806 GNDA.t228 GNDA.n8 65.8183
R5807 GNDA.n5557 GNDA.t228 65.8183
R5808 GNDA.t228 GNDA.n6 65.8183
R5809 GNDA.t228 GNDA.n4 65.8183
R5810 GNDA.n737 GNDA.t255 65.3505
R5811 GNDA.n736 GNDA.t230 65.3505
R5812 GNDA.n640 GNDA.t266 65.3505
R5813 GNDA.n639 GNDA.t253 65.3505
R5814 GNDA.n4091 GNDA.t201 65.3505
R5815 GNDA.n4089 GNDA.t197 65.3505
R5816 GNDA.n722 GNDA.n674 64.0005
R5817 GNDA.n722 GNDA.n721 64.0005
R5818 GNDA.n4006 GNDA.t273 63.4011
R5819 GNDA.n3996 GNDA.t206 63.4011
R5820 GNDA.n2545 GNDA.n2544 63.1009
R5821 GNDA.n664 GNDA.t257 62.2505
R5822 GNDA.n646 GNDA.t268 62.2505
R5823 GNDA.n693 GNDA.t204 62.2505
R5824 GNDA.n606 GNDA.t213 62.2505
R5825 GNDA.t105 GNDA.n2008 62.0993
R5826 GNDA.n2482 GNDA.t10 62.0993
R5827 GNDA.n4280 GNDA.n431 59.2425
R5828 GNDA.n3480 GNDA.n631 59.2425
R5829 GNDA.n3384 GNDA.n3383 59.2425
R5830 GNDA.n4131 GNDA.n4130 59.2425
R5831 GNDA.n2083 GNDA.t115 58.0929
R5832 GNDA.n2026 GNDA.t88 58.0929
R5833 GNDA.t242 GNDA.n2501 57.8461
R5834 GNDA.n2000 GNDA.t217 57.8461
R5835 GNDA.t185 GNDA.n5330 57.8461
R5836 GNDA.t224 GNDA.n2292 57.8461
R5837 GNDA.t251 GNDA.n5157 57.8461
R5838 GNDA.t210 GNDA.n60 57.8461
R5839 GNDA.t243 GNDA.n5115 57.8461
R5840 GNDA.n1799 GNDA.t258 57.8461
R5841 GNDA.t228 GNDA.n5556 57.8461
R5842 GNDA.n1930 GNDA.n1929 57.0913
R5843 GNDA.n1453 GNDA.n1450 56.3995
R5844 GNDA.n2304 GNDA.n2187 56.3995
R5845 GNDA.n5152 GNDA.n5151 56.3995
R5846 GNDA.n5128 GNDA.n234 56.3995
R5847 GNDA.n2533 GNDA.n1450 56.3995
R5848 GNDA.n2304 GNDA.n2303 56.3995
R5849 GNDA.n5383 GNDA.n5382 56.3995
R5850 GNDA.n5384 GNDA.n5383 56.3995
R5851 GNDA.n1854 GNDA.n280 56.3995
R5852 GNDA.n5151 GNDA.n227 56.3995
R5853 GNDA.n5126 GNDA.n234 56.3995
R5854 GNDA.t242 GNDA.n1582 55.2026
R5855 GNDA.n1960 GNDA.t217 55.2026
R5856 GNDA.t185 GNDA.n175 55.2026
R5857 GNDA.t243 GNDA.n5020 55.2026
R5858 GNDA.t224 GNDA.n2198 55.2026
R5859 GNDA.t251 GNDA.n5167 55.2026
R5860 GNDA.t210 GNDA.n70 55.2026
R5861 GNDA.n1765 GNDA.t258 55.2026
R5862 GNDA.t228 GNDA.n9 55.2026
R5863 GNDA.n1636 GNDA.n1590 53.3664
R5864 GNDA.n1632 GNDA.n1570 53.3664
R5865 GNDA.n1628 GNDA.n1589 53.3664
R5866 GNDA.n1624 GNDA.n1572 53.3664
R5867 GNDA.n1613 GNDA.n1583 53.3664
R5868 GNDA.n1609 GNDA.n1584 53.3664
R5869 GNDA.n1605 GNDA.n1585 53.3664
R5870 GNDA.n1588 GNDA.n1587 53.3664
R5871 GNDA.n1596 GNDA.n1569 53.3664
R5872 GNDA.n2490 GNDA.n1571 53.3664
R5873 GNDA.n2503 GNDA.n2502 53.3664
R5874 GNDA.n1581 GNDA.n1580 53.3664
R5875 GNDA.n1640 GNDA.n1594 53.3664
R5876 GNDA.n1641 GNDA.n1593 53.3664
R5877 GNDA.n1645 GNDA.n1592 53.3664
R5878 GNDA.n1649 GNDA.n1591 53.3664
R5879 GNDA.n1637 GNDA.n1594 53.3664
R5880 GNDA.n1644 GNDA.n1593 53.3664
R5881 GNDA.n1648 GNDA.n1592 53.3664
R5882 GNDA.n1651 GNDA.n1591 53.3664
R5883 GNDA.n1621 GNDA.n1572 53.3664
R5884 GNDA.n1625 GNDA.n1589 53.3664
R5885 GNDA.n1629 GNDA.n1570 53.3664
R5886 GNDA.n1633 GNDA.n1590 53.3664
R5887 GNDA.n1604 GNDA.n1588 53.3664
R5888 GNDA.n1608 GNDA.n1585 53.3664
R5889 GNDA.n1612 GNDA.n1584 53.3664
R5890 GNDA.n1616 GNDA.n1583 53.3664
R5891 GNDA.n1586 GNDA.n1581 53.3664
R5892 GNDA.n2502 GNDA.n1568 53.3664
R5893 GNDA.n1571 GNDA.n1567 53.3664
R5894 GNDA.n2489 GNDA.n1569 53.3664
R5895 GNDA.n1976 GNDA.n1939 53.3664
R5896 GNDA.n1975 GNDA.n1974 53.3664
R5897 GNDA.n1968 GNDA.n1941 53.3664
R5898 GNDA.n1967 GNDA.n1966 53.3664
R5899 GNDA.n1958 GNDA.n1957 53.3664
R5900 GNDA.n1953 GNDA.n1947 53.3664
R5901 GNDA.n1951 GNDA.n1950 53.3664
R5902 GNDA.n2034 GNDA.n1901 53.3664
R5903 GNDA.n2003 GNDA.n2002 53.3664
R5904 GNDA.n2016 GNDA.n2015 53.3664
R5905 GNDA.n2019 GNDA.n2018 53.3664
R5906 GNDA.n2032 GNDA.n2031 53.3664
R5907 GNDA.n1983 GNDA.n1982 53.3664
R5908 GNDA.n1985 GNDA.n1984 53.3664
R5909 GNDA.n1990 GNDA.n1989 53.3664
R5910 GNDA.n1993 GNDA.n1992 53.3664
R5911 GNDA.n1982 GNDA.n1981 53.3664
R5912 GNDA.n1984 GNDA.n1937 53.3664
R5913 GNDA.n1991 GNDA.n1990 53.3664
R5914 GNDA.n1992 GNDA.n1935 53.3664
R5915 GNDA.n1966 GNDA.n1965 53.3664
R5916 GNDA.n1969 GNDA.n1968 53.3664
R5917 GNDA.n1974 GNDA.n1973 53.3664
R5918 GNDA.n1977 GNDA.n1976 53.3664
R5919 GNDA.n1948 GNDA.n1901 53.3664
R5920 GNDA.n1952 GNDA.n1951 53.3664
R5921 GNDA.n1947 GNDA.n1945 53.3664
R5922 GNDA.n1959 GNDA.n1958 53.3664
R5923 GNDA.n2033 GNDA.n2032 53.3664
R5924 GNDA.n2018 GNDA.n1902 53.3664
R5925 GNDA.n2017 GNDA.n2016 53.3664
R5926 GNDA.n2002 GNDA.n1908 53.3664
R5927 GNDA.n5312 GNDA.n181 53.3664
R5928 GNDA.n5308 GNDA.n170 53.3664
R5929 GNDA.n5304 GNDA.n180 53.3664
R5930 GNDA.n5300 GNDA.n173 53.3664
R5931 GNDA.n5289 GNDA.n176 53.3664
R5932 GNDA.n5285 GNDA.n177 53.3664
R5933 GNDA.n5281 GNDA.n178 53.3664
R5934 GNDA.n5277 GNDA.n179 53.3664
R5935 GNDA.n5332 GNDA.n5331 53.3664
R5936 GNDA.n216 GNDA.n171 53.3664
R5937 GNDA.n212 GNDA.n172 53.3664
R5938 GNDA.n205 GNDA.n174 53.3664
R5939 GNDA.n5316 GNDA.n185 53.3664
R5940 GNDA.n5317 GNDA.n184 53.3664
R5941 GNDA.n5321 GNDA.n183 53.3664
R5942 GNDA.n5325 GNDA.n182 53.3664
R5943 GNDA.n5313 GNDA.n185 53.3664
R5944 GNDA.n5320 GNDA.n184 53.3664
R5945 GNDA.n5324 GNDA.n183 53.3664
R5946 GNDA.n5328 GNDA.n182 53.3664
R5947 GNDA.n5297 GNDA.n173 53.3664
R5948 GNDA.n5301 GNDA.n180 53.3664
R5949 GNDA.n5305 GNDA.n170 53.3664
R5950 GNDA.n5309 GNDA.n181 53.3664
R5951 GNDA.n5280 GNDA.n179 53.3664
R5952 GNDA.n5284 GNDA.n178 53.3664
R5953 GNDA.n5288 GNDA.n177 53.3664
R5954 GNDA.n5292 GNDA.n176 53.3664
R5955 GNDA.n5276 GNDA.n174 53.3664
R5956 GNDA.n204 GNDA.n172 53.3664
R5957 GNDA.n213 GNDA.n171 53.3664
R5958 GNDA.n5331 GNDA.n169 53.3664
R5959 GNDA.n5097 GNDA.n5026 53.3664
R5960 GNDA.n5093 GNDA.n5015 53.3664
R5961 GNDA.n5089 GNDA.n5025 53.3664
R5962 GNDA.n5085 GNDA.n5018 53.3664
R5963 GNDA.n5074 GNDA.n5021 53.3664
R5964 GNDA.n5070 GNDA.n5022 53.3664
R5965 GNDA.n5066 GNDA.n5023 53.3664
R5966 GNDA.n5062 GNDA.n5024 53.3664
R5967 GNDA.n5117 GNDA.n5116 53.3664
R5968 GNDA.n5039 GNDA.n5016 53.3664
R5969 GNDA.n5047 GNDA.n5017 53.3664
R5970 GNDA.n5054 GNDA.n5019 53.3664
R5971 GNDA.n5101 GNDA.n5030 53.3664
R5972 GNDA.n5102 GNDA.n5029 53.3664
R5973 GNDA.n5106 GNDA.n5028 53.3664
R5974 GNDA.n5110 GNDA.n5027 53.3664
R5975 GNDA.n5098 GNDA.n5030 53.3664
R5976 GNDA.n5105 GNDA.n5029 53.3664
R5977 GNDA.n5109 GNDA.n5028 53.3664
R5978 GNDA.n5113 GNDA.n5027 53.3664
R5979 GNDA.n5082 GNDA.n5018 53.3664
R5980 GNDA.n5086 GNDA.n5025 53.3664
R5981 GNDA.n5090 GNDA.n5015 53.3664
R5982 GNDA.n5094 GNDA.n5026 53.3664
R5983 GNDA.n5065 GNDA.n5024 53.3664
R5984 GNDA.n5069 GNDA.n5023 53.3664
R5985 GNDA.n5073 GNDA.n5022 53.3664
R5986 GNDA.n5077 GNDA.n5021 53.3664
R5987 GNDA.n2245 GNDA.n2205 53.3664
R5988 GNDA.n2241 GNDA.n2194 53.3664
R5989 GNDA.n2237 GNDA.n2204 53.3664
R5990 GNDA.n2233 GNDA.n2197 53.3664
R5991 GNDA.n2222 GNDA.n2199 53.3664
R5992 GNDA.n2218 GNDA.n2200 53.3664
R5993 GNDA.n2214 GNDA.n2201 53.3664
R5994 GNDA.n2203 GNDA.n2202 53.3664
R5995 GNDA.n2211 GNDA.n2193 53.3664
R5996 GNDA.n2280 GNDA.n2195 53.3664
R5997 GNDA.n2273 GNDA.n2196 53.3664
R5998 GNDA.n2294 GNDA.n2293 53.3664
R5999 GNDA.n2249 GNDA.n2209 53.3664
R6000 GNDA.n2250 GNDA.n2208 53.3664
R6001 GNDA.n2254 GNDA.n2207 53.3664
R6002 GNDA.n2258 GNDA.n2206 53.3664
R6003 GNDA.n2246 GNDA.n2209 53.3664
R6004 GNDA.n2253 GNDA.n2208 53.3664
R6005 GNDA.n2257 GNDA.n2207 53.3664
R6006 GNDA.n2260 GNDA.n2206 53.3664
R6007 GNDA.n2230 GNDA.n2197 53.3664
R6008 GNDA.n2234 GNDA.n2204 53.3664
R6009 GNDA.n2238 GNDA.n2194 53.3664
R6010 GNDA.n2242 GNDA.n2205 53.3664
R6011 GNDA.n2213 GNDA.n2203 53.3664
R6012 GNDA.n2217 GNDA.n2201 53.3664
R6013 GNDA.n2221 GNDA.n2200 53.3664
R6014 GNDA.n2225 GNDA.n2199 53.3664
R6015 GNDA.n2293 GNDA.n2192 53.3664
R6016 GNDA.n2196 GNDA.n2191 53.3664
R6017 GNDA.n2272 GNDA.n2195 53.3664
R6018 GNDA.n2279 GNDA.n2193 53.3664
R6019 GNDA.n5237 GNDA.n5173 53.3664
R6020 GNDA.n5234 GNDA.n5163 53.3664
R6021 GNDA.n5230 GNDA.n5172 53.3664
R6022 GNDA.n5226 GNDA.n5165 53.3664
R6023 GNDA.n5215 GNDA.n5168 53.3664
R6024 GNDA.n5211 GNDA.n5169 53.3664
R6025 GNDA.n5207 GNDA.n5170 53.3664
R6026 GNDA.n5203 GNDA.n5171 53.3664
R6027 GNDA.n5263 GNDA.n5158 53.3664
R6028 GNDA.n5256 GNDA.n5255 53.3664
R6029 GNDA.n5188 GNDA.n5164 53.3664
R6030 GNDA.n5195 GNDA.n5166 53.3664
R6031 GNDA.n5254 GNDA.n5253 53.3664
R6032 GNDA.n5178 GNDA.n5176 53.3664
R6033 GNDA.n5248 GNDA.n5175 53.3664
R6034 GNDA.n5244 GNDA.n5174 53.3664
R6035 GNDA.n5254 GNDA.n5177 53.3664
R6036 GNDA.n5249 GNDA.n5176 53.3664
R6037 GNDA.n5245 GNDA.n5175 53.3664
R6038 GNDA.n5241 GNDA.n5174 53.3664
R6039 GNDA.n5223 GNDA.n5165 53.3664
R6040 GNDA.n5227 GNDA.n5172 53.3664
R6041 GNDA.n5231 GNDA.n5163 53.3664
R6042 GNDA.n5235 GNDA.n5173 53.3664
R6043 GNDA.n5206 GNDA.n5171 53.3664
R6044 GNDA.n5210 GNDA.n5170 53.3664
R6045 GNDA.n5214 GNDA.n5169 53.3664
R6046 GNDA.n5218 GNDA.n5168 53.3664
R6047 GNDA.n5202 GNDA.n5166 53.3664
R6048 GNDA.n5194 GNDA.n5164 53.3664
R6049 GNDA.n5255 GNDA.n5162 53.3664
R6050 GNDA.n5161 GNDA.n5158 53.3664
R6051 GNDA.n5516 GNDA.n76 53.3664
R6052 GNDA.n5513 GNDA.n66 53.3664
R6053 GNDA.n5509 GNDA.n75 53.3664
R6054 GNDA.n5505 GNDA.n68 53.3664
R6055 GNDA.n5494 GNDA.n71 53.3664
R6056 GNDA.n5490 GNDA.n72 53.3664
R6057 GNDA.n5486 GNDA.n73 53.3664
R6058 GNDA.n5482 GNDA.n74 53.3664
R6059 GNDA.n5542 GNDA.n61 53.3664
R6060 GNDA.n5535 GNDA.n5534 53.3664
R6061 GNDA.n5467 GNDA.n67 53.3664
R6062 GNDA.n5474 GNDA.n69 53.3664
R6063 GNDA.n5533 GNDA.n5532 53.3664
R6064 GNDA.n81 GNDA.n79 53.3664
R6065 GNDA.n5527 GNDA.n78 53.3664
R6066 GNDA.n5523 GNDA.n77 53.3664
R6067 GNDA.n5533 GNDA.n80 53.3664
R6068 GNDA.n5528 GNDA.n79 53.3664
R6069 GNDA.n5524 GNDA.n78 53.3664
R6070 GNDA.n5520 GNDA.n77 53.3664
R6071 GNDA.n5502 GNDA.n68 53.3664
R6072 GNDA.n5506 GNDA.n75 53.3664
R6073 GNDA.n5510 GNDA.n66 53.3664
R6074 GNDA.n5514 GNDA.n76 53.3664
R6075 GNDA.n5485 GNDA.n74 53.3664
R6076 GNDA.n5489 GNDA.n73 53.3664
R6077 GNDA.n5493 GNDA.n72 53.3664
R6078 GNDA.n5497 GNDA.n71 53.3664
R6079 GNDA.n5481 GNDA.n69 53.3664
R6080 GNDA.n5473 GNDA.n67 53.3664
R6081 GNDA.n5534 GNDA.n65 53.3664
R6082 GNDA.n64 GNDA.n61 53.3664
R6083 GNDA.n5061 GNDA.n5019 53.3664
R6084 GNDA.n5053 GNDA.n5017 53.3664
R6085 GNDA.n5046 GNDA.n5016 53.3664
R6086 GNDA.n5116 GNDA.n5014 53.3664
R6087 GNDA.n1782 GNDA.n1781 53.3664
R6088 GNDA.n1775 GNDA.n1740 53.3664
R6089 GNDA.n1774 GNDA.n1773 53.3664
R6090 GNDA.n1767 GNDA.n1742 53.3664
R6091 GNDA.n1760 GNDA.n1746 53.3664
R6092 GNDA.n1758 GNDA.n1757 53.3664
R6093 GNDA.n1753 GNDA.n1750 53.3664
R6094 GNDA.n1751 GNDA.n1722 53.3664
R6095 GNDA.n1873 GNDA.n1872 53.3664
R6096 GNDA.n1876 GNDA.n1875 53.3664
R6097 GNDA.n2074 GNDA.n2073 53.3664
R6098 GNDA.n2077 GNDA.n2076 53.3664
R6099 GNDA.n1783 GNDA.n1738 53.3664
R6100 GNDA.n1789 GNDA.n1788 53.3664
R6101 GNDA.n1792 GNDA.n1791 53.3664
R6102 GNDA.n1797 GNDA.n1796 53.3664
R6103 GNDA.n1784 GNDA.n1783 53.3664
R6104 GNDA.n1790 GNDA.n1789 53.3664
R6105 GNDA.n1791 GNDA.n1736 53.3664
R6106 GNDA.n1798 GNDA.n1797 53.3664
R6107 GNDA.n1768 GNDA.n1767 53.3664
R6108 GNDA.n1773 GNDA.n1772 53.3664
R6109 GNDA.n1776 GNDA.n1775 53.3664
R6110 GNDA.n1781 GNDA.n1780 53.3664
R6111 GNDA.n1752 GNDA.n1751 53.3664
R6112 GNDA.n1750 GNDA.n1747 53.3664
R6113 GNDA.n1759 GNDA.n1758 53.3664
R6114 GNDA.n1746 GNDA.n1744 53.3664
R6115 GNDA.n2078 GNDA.n2077 53.3664
R6116 GNDA.n2075 GNDA.n2074 53.3664
R6117 GNDA.n1875 GNDA.n1725 53.3664
R6118 GNDA.n1874 GNDA.n1873 53.3664
R6119 GNDA.n5435 GNDA.n15 53.3664
R6120 GNDA.n5431 GNDA.n5 53.3664
R6121 GNDA.n5427 GNDA.n14 53.3664
R6122 GNDA.n5423 GNDA.n7 53.3664
R6123 GNDA.n5412 GNDA.n10 53.3664
R6124 GNDA.n5408 GNDA.n11 53.3664
R6125 GNDA.n5404 GNDA.n12 53.3664
R6126 GNDA.n5400 GNDA.n13 53.3664
R6127 GNDA.n21 GNDA.n4 53.3664
R6128 GNDA.n37 GNDA.n6 53.3664
R6129 GNDA.n5558 GNDA.n5557 53.3664
R6130 GNDA.n5392 GNDA.n8 53.3664
R6131 GNDA.n5439 GNDA.n19 53.3664
R6132 GNDA.n5440 GNDA.n18 53.3664
R6133 GNDA.n5444 GNDA.n17 53.3664
R6134 GNDA.n5448 GNDA.n16 53.3664
R6135 GNDA.n5436 GNDA.n19 53.3664
R6136 GNDA.n5443 GNDA.n18 53.3664
R6137 GNDA.n5447 GNDA.n17 53.3664
R6138 GNDA.n5450 GNDA.n16 53.3664
R6139 GNDA.n5420 GNDA.n7 53.3664
R6140 GNDA.n5424 GNDA.n14 53.3664
R6141 GNDA.n5428 GNDA.n5 53.3664
R6142 GNDA.n5432 GNDA.n15 53.3664
R6143 GNDA.n5403 GNDA.n13 53.3664
R6144 GNDA.n5407 GNDA.n12 53.3664
R6145 GNDA.n5411 GNDA.n11 53.3664
R6146 GNDA.n5415 GNDA.n10 53.3664
R6147 GNDA.n5399 GNDA.n8 53.3664
R6148 GNDA.n5557 GNDA.n3 53.3664
R6149 GNDA.n6 GNDA.n2 53.3664
R6150 GNDA.n36 GNDA.n4 53.3664
R6151 GNDA.n1864 GNDA.n1863 53.085
R6152 GNDA.n1930 GNDA.n1914 53.085
R6153 GNDA.n2044 GNDA.n2041 53.085
R6154 GNDA.n4121 GNDA.t212 52.2393
R6155 GNDA.t203 GNDA.n632 52.2393
R6156 GNDA.t286 GNDA.n2083 52.0834
R6157 GNDA.n2026 GNDA.t26 52.0834
R6158 GNDA.n2507 GNDA.t70 52.0834
R6159 GNDA.n5006 GNDA.n99 50.8806
R6160 GNDA.n5006 GNDA.n5005 50.8806
R6161 GNDA.n5005 GNDA.n5004 50.8806
R6162 GNDA.n5004 GNDA.n292 50.8806
R6163 GNDA.n4998 GNDA.n292 50.8806
R6164 GNDA.n4997 GNDA.n4996 50.8806
R6165 GNDA.n4996 GNDA.n296 50.8806
R6166 GNDA.n4990 GNDA.n296 50.8806
R6167 GNDA.n4990 GNDA.n4989 50.8806
R6168 GNDA.n4989 GNDA.n4988 50.8806
R6169 GNDA.n4982 GNDA.n4981 50.8806
R6170 GNDA.n4981 GNDA.n4980 50.8806
R6171 GNDA.n4980 GNDA.n351 50.8806
R6172 GNDA.n4974 GNDA.n351 50.8806
R6173 GNDA.n4974 GNDA.n4973 50.8806
R6174 GNDA.n4964 GNDA.n356 50.8806
R6175 GNDA.n4964 GNDA.n4963 50.8806
R6176 GNDA.n4963 GNDA.n4962 50.8806
R6177 GNDA.n4962 GNDA.n362 50.8806
R6178 GNDA.n4956 GNDA.n362 50.8806
R6179 GNDA.n4954 GNDA.n367 50.8806
R6180 GNDA.n4948 GNDA.n367 50.8806
R6181 GNDA.n4948 GNDA.n4947 50.8806
R6182 GNDA.n4947 GNDA.n4946 50.8806
R6183 GNDA.n4946 GNDA.n416 50.8806
R6184 GNDA.n4940 GNDA.n4939 50.8806
R6185 GNDA.n4939 GNDA.n4938 50.8806
R6186 GNDA.n4938 GNDA.n420 50.8806
R6187 GNDA.n4932 GNDA.n420 50.8806
R6188 GNDA.n4932 GNDA.n4931 50.8806
R6189 GNDA.t174 GNDA.t163 48.7908
R6190 GNDA.t171 GNDA.t164 48.7908
R6191 GNDA.t172 GNDA.t160 48.7908
R6192 GNDA.t168 GNDA.t158 48.7908
R6193 GNDA.t166 GNDA.t176 48.7908
R6194 GNDA.t121 GNDA.t86 48.7908
R6195 GNDA.t73 GNDA.t142 48.7908
R6196 GNDA.t54 GNDA.t117 48.7908
R6197 GNDA.t12 GNDA.t87 48.7908
R6198 GNDA.t285 GNDA.t85 48.7908
R6199 GNDA.t275 GNDA.n106 48.077
R6200 GNDA.n2008 GNDA.t222 48.077
R6201 GNDA.n2482 GNDA.t288 48.077
R6202 GNDA.t186 GNDA.n5370 47.6748
R6203 GNDA.t186 GNDA.n106 47.0754
R6204 GNDA.n2480 GNDA.t148 47.0754
R6205 GNDA.t208 GNDA.t270 46.5731
R6206 GNDA.t263 GNDA.t215 46.5731
R6207 GNDA.t226 GNDA.t194 46.5731
R6208 GNDA.t180 GNDA.t245 46.5731
R6209 GNDA.n2084 GNDA.t155 46.0738
R6210 GNDA.n1914 GNDA.n1661 43.069
R6211 GNDA.n2023 GNDA.t186 43.069
R6212 GNDA.t186 GNDA.n2507 43.069
R6213 GNDA.n4017 GNDA.t241 42.6297
R6214 GNDA.t261 GNDA.n4016 42.6297
R6215 GNDA.n679 GNDA.t199 42.6297
R6216 GNDA.n707 GNDA.t220 42.6297
R6217 GNDA.t222 GNDA.n2007 42.0674
R6218 GNDA.t288 GNDA.n2481 42.0674
R6219 GNDA.n2009 GNDA.t42 41.0658
R6220 GNDA.t186 GNDA.t148 40.0642
R6221 GNDA.n4066 GNDA.n632 38.8065
R6222 GNDA.n2085 GNDA.t286 38.0611
R6223 GNDA.t26 GNDA.n2025 38.0611
R6224 GNDA.t163 GNDA.t138 37.7021
R6225 GNDA.t22 GNDA.t166 37.7021
R6226 GNDA.t86 GNDA.t80 37.7021
R6227 GNDA.t136 GNDA.t285 37.7021
R6228 GNDA.n1863 GNDA.n1861 37.0595
R6229 GNDA.n1867 GNDA.t78 37.0595
R6230 GNDA.n2044 GNDA.n2040 37.0595
R6231 GNDA.t155 GNDA.t188 35.0563
R6232 GNDA.n4020 GNDA.n4019 34.5991
R6233 GNDA.n4022 GNDA.n4021 34.5991
R6234 GNDA.n4024 GNDA.n4023 34.5991
R6235 GNDA.n4026 GNDA.n4025 34.5991
R6236 GNDA.n4028 GNDA.n4027 34.5991
R6237 GNDA.n4030 GNDA.n4029 34.5991
R6238 GNDA.n4032 GNDA.n4031 34.5991
R6239 GNDA.n4034 GNDA.n4033 34.5991
R6240 GNDA.n4036 GNDA.n4035 34.5991
R6241 GNDA.n4038 GNDA.n4037 34.5991
R6242 GNDA.n4040 GNDA.n4039 34.5991
R6243 GNDA.n4042 GNDA.n4041 34.5991
R6244 GNDA.n711 GNDA.n710 34.5991
R6245 GNDA.n3383 GNDA.t208 33.2666
R6246 GNDA.t215 GNDA.n631 33.2666
R6247 GNDA.n4130 GNDA.t226 33.2666
R6248 GNDA.t245 GNDA.n431 33.2666
R6249 GNDA.t79 GNDA.t92 33.1455
R6250 GNDA.n2064 GNDA.n2053 33.0531
R6251 GNDA.n1574 GNDA.t280 33.0531
R6252 GNDA.t186 GNDA.n26 32.9056
R6253 GNDA.t186 GNDA.n107 32.9056
R6254 GNDA.t21 GNDA.t59 32.8363
R6255 GNDA.t112 GNDA.t212 32.8363
R6256 GNDA.t178 GNDA.t203 32.8363
R6257 GNDA.t97 GNDA.t41 32.8363
R6258 GNDA.n2521 GNDA.n2520 32.3969
R6259 GNDA.t88 GNDA.n2024 32.0515
R6260 GNDA.n4969 GNDA.n4968 31.3605
R6261 GNDA.n3381 GNDA.t209 31.1255
R6262 GNDA.n4914 GNDA.t246 31.1255
R6263 GNDA.n4128 GNDA.t227 31.1255
R6264 GNDA.n4068 GNDA.t216 31.1255
R6265 GNDA.t183 GNDA.t103 30.3834
R6266 GNDA.t103 GNDA.t113 30.3834
R6267 GNDA.t113 GNDA.t290 30.3834
R6268 GNDA.n1929 GNDA.n1916 30.0483
R6269 GNDA.t110 GNDA.n2084 29.0467
R6270 GNDA.t164 GNDA.t33 28.8311
R6271 GNDA.t127 GNDA.t168 28.8311
R6272 GNDA.t142 GNDA.t144 28.8311
R6273 GNDA.t7 GNDA.t12 28.8311
R6274 GNDA.n4060 GNDA.t112 28.3587
R6275 GNDA.n4044 GNDA.t178 28.3587
R6276 GNDA.n2010 GNDA.t105 28.0451
R6277 GNDA.t191 GNDA.n2480 28.0451
R6278 GNDA.n1638 GNDA.n1635 27.5561
R6279 GNDA.n1980 GNDA.n1979 27.5561
R6280 GNDA.n5314 GNDA.n5311 27.5561
R6281 GNDA.n5099 GNDA.n5096 27.5561
R6282 GNDA.n2247 GNDA.n2244 27.5561
R6283 GNDA.n5239 GNDA.n5238 27.5561
R6284 GNDA.n5518 GNDA.n5517 27.5561
R6285 GNDA.n1785 GNDA.n1739 27.5561
R6286 GNDA.n5437 GNDA.n5434 27.5561
R6287 GNDA.n4916 GNDA.t82 27.1216
R6288 GNDA.n633 GNDA.t9 27.1216
R6289 GNDA.n2041 GNDA.n1660 27.0435
R6290 GNDA.n2518 GNDA.n1559 27.0435
R6291 GNDA.n2545 GNDA.n1444 27.0435
R6292 GNDA.n1619 GNDA.n1618 26.6672
R6293 GNDA.n1963 GNDA.n1962 26.6672
R6294 GNDA.n5295 GNDA.n5294 26.6672
R6295 GNDA.n5080 GNDA.n5079 26.6672
R6296 GNDA.n2228 GNDA.n2227 26.6672
R6297 GNDA.n5221 GNDA.n5220 26.6672
R6298 GNDA.n5500 GNDA.n5499 26.6672
R6299 GNDA.n1763 GNDA.n1743 26.6672
R6300 GNDA.n5418 GNDA.n5417 26.6672
R6301 GNDA.n3383 GNDA.n3382 26.6134
R6302 GNDA.n4067 GNDA.n631 26.6134
R6303 GNDA.n4130 GNDA.n4129 26.6134
R6304 GNDA.n4915 GNDA.n431 26.6134
R6305 GNDA.n4998 GNDA.t186 26.5712
R6306 GNDA.n4973 GNDA.t186 26.5712
R6307 GNDA.t186 GNDA.n416 26.5712
R6308 GNDA.n2056 GNDA.n2055 25.3679
R6309 GNDA.t115 GNDA.t74 25.0403
R6310 GNDA.t10 GNDA.t14 25.0403
R6311 GNDA.t186 GNDA.n4997 24.3099
R6312 GNDA.t186 GNDA.n356 24.3099
R6313 GNDA.n4940 GNDA.t186 24.3099
R6314 GNDA.n1455 GNDA.n1445 24.0387
R6315 GNDA.n1443 GNDA.t62 24.0005
R6316 GNDA.n1443 GNDA.t71 24.0005
R6317 GNDA.n1442 GNDA.t37 24.0005
R6318 GNDA.n1442 GNDA.t94 24.0005
R6319 GNDA.n1441 GNDA.t289 24.0005
R6320 GNDA.n1441 GNDA.t11 24.0005
R6321 GNDA.n1438 GNDA.t27 24.0005
R6322 GNDA.n1438 GNDA.t249 24.0005
R6323 GNDA.n1437 GNDA.t130 24.0005
R6324 GNDA.n1437 GNDA.t89 24.0005
R6325 GNDA.n1436 GNDA.t106 24.0005
R6326 GNDA.n1436 GNDA.t278 24.0005
R6327 GNDA.n1433 GNDA.t287 24.0005
R6328 GNDA.n1433 GNDA.t111 24.0005
R6329 GNDA.n1432 GNDA.t25 24.0005
R6330 GNDA.n1432 GNDA.t116 24.0005
R6331 GNDA.n1431 GNDA.t96 24.0005
R6332 GNDA.n1431 GNDA.t132 24.0005
R6333 GNDA.n1428 GNDA.t291 24.0005
R6334 GNDA.n1428 GNDA.t233 24.0005
R6335 GNDA.n1427 GNDA.t104 24.0005
R6336 GNDA.n1427 GNDA.t114 24.0005
R6337 GNDA.t16 GNDA.t75 23.8245
R6338 GNDA.t282 GNDA.t283 23.8245
R6339 GNDA.n1424 GNDA.t19 23.4782
R6340 GNDA.n2067 GNDA.n2066 23.0371
R6341 GNDA.n1659 GNDA.n1439 22.53
R6342 GNDA.n4917 GNDA.t51 21.5269
R6343 GNDA.n2547 GNDA.n2546 20.8233
R6344 GNDA.n2472 GNDA.n1440 20.8233
R6345 GNDA.n1915 GNDA.n1435 20.8233
R6346 GNDA.n1913 GNDA.n1434 20.8233
R6347 GNDA.n1865 GNDA.n1430 20.8233
R6348 GNDA.n1862 GNDA.n1429 20.8233
R6349 GNDA.n1426 GNDA.n1425 20.8233
R6350 GNDA.t51 GNDA.t2 20.6659
R6351 GNDA.t2 GNDA.t281 20.6659
R6352 GNDA.t1 GNDA.t279 20.6659
R6353 GNDA.t90 GNDA.t1 20.6659
R6354 GNDA.n2473 GNDA.t186 20.0324
R6355 GNDA.t33 GNDA.t172 19.9602
R6356 GNDA.t160 GNDA.t127 19.9602
R6357 GNDA.t144 GNDA.t54 19.9602
R6358 GNDA.t117 GNDA.t7 19.9602
R6359 GNDA.n4898 GNDA.t140 19.7005
R6360 GNDA.n4898 GNDA.t151 19.7005
R6361 GNDA.n4896 GNDA.t67 19.7005
R6362 GNDA.n4896 GNDA.t72 19.7005
R6363 GNDA.n4894 GNDA.t69 19.7005
R6364 GNDA.n4894 GNDA.t50 19.7005
R6365 GNDA.n4892 GNDA.t143 19.7005
R6366 GNDA.n4892 GNDA.t55 19.7005
R6367 GNDA.n4890 GNDA.t141 19.7005
R6368 GNDA.n4890 GNDA.t60 19.7005
R6369 GNDA.n4889 GNDA.t157 19.7005
R6370 GNDA.n4889 GNDA.t68 19.7005
R6371 GNDA.n1000 GNDA.t175 19.7005
R6372 GNDA.n1000 GNDA.t154 19.7005
R6373 GNDA.n1001 GNDA.t177 19.7005
R6374 GNDA.n1001 GNDA.t165 19.7005
R6375 GNDA.n1003 GNDA.t159 19.7005
R6376 GNDA.n1003 GNDA.t167 19.7005
R6377 GNDA.n1005 GNDA.t162 19.7005
R6378 GNDA.n1005 GNDA.t170 19.7005
R6379 GNDA.n1007 GNDA.t161 19.7005
R6380 GNDA.n1007 GNDA.t169 19.7005
R6381 GNDA.n1009 GNDA.t150 19.7005
R6382 GNDA.n1009 GNDA.t173 19.7005
R6383 GNDA.n2040 GNDA.t248 18.0292
R6384 GNDA.t100 GNDA.t32 17.9109
R6385 GNDA.t56 GNDA.t239 17.9109
R6386 GNDA.t260 GNDA.t125 17.9109
R6387 GNDA.t77 GNDA.t39 17.9109
R6388 GNDA.n2422 GNDA.n2396 17.5843
R6389 GNDA.n2328 GNDA.n2176 17.5843
R6390 GNDA.n4928 GNDA.n422 17.5843
R6391 GNDA.n4924 GNDA.n4917 17.5479
R6392 GNDA.n262 GNDA.n259 16.9379
R6393 GNDA.n5147 GNDA.n5009 16.9379
R6394 GNDA.n1833 GNDA.n1802 16.9379
R6395 GNDA.n5366 GNDA.n133 16.7709
R6396 GNDA.n1688 GNDA.n162 16.7709
R6397 GNDA.n2175 GNDA.n84 16.7709
R6398 GNDA.n2387 GNDA.n2386 16.7709
R6399 GNDA.t186 GNDA.n105 16.4553
R6400 GNDA.n1639 GNDA.n1638 16.0005
R6401 GNDA.n1642 GNDA.n1639 16.0005
R6402 GNDA.n1643 GNDA.n1642 16.0005
R6403 GNDA.n1646 GNDA.n1643 16.0005
R6404 GNDA.n1647 GNDA.n1646 16.0005
R6405 GNDA.n1650 GNDA.n1647 16.0005
R6406 GNDA.n1652 GNDA.n1650 16.0005
R6407 GNDA.n1653 GNDA.n1652 16.0005
R6408 GNDA.n1635 GNDA.n1634 16.0005
R6409 GNDA.n1634 GNDA.n1631 16.0005
R6410 GNDA.n1631 GNDA.n1630 16.0005
R6411 GNDA.n1630 GNDA.n1627 16.0005
R6412 GNDA.n1627 GNDA.n1626 16.0005
R6413 GNDA.n1626 GNDA.n1623 16.0005
R6414 GNDA.n1623 GNDA.n1622 16.0005
R6415 GNDA.n1622 GNDA.n1619 16.0005
R6416 GNDA.n1618 GNDA.n1615 16.0005
R6417 GNDA.n1615 GNDA.n1614 16.0005
R6418 GNDA.n1614 GNDA.n1611 16.0005
R6419 GNDA.n1611 GNDA.n1610 16.0005
R6420 GNDA.n1610 GNDA.n1607 16.0005
R6421 GNDA.n1607 GNDA.n1606 16.0005
R6422 GNDA.n1606 GNDA.n1603 16.0005
R6423 GNDA.n1603 GNDA.n1449 16.0005
R6424 GNDA.n1980 GNDA.n1938 16.0005
R6425 GNDA.n1986 GNDA.n1938 16.0005
R6426 GNDA.n1987 GNDA.n1986 16.0005
R6427 GNDA.n1988 GNDA.n1987 16.0005
R6428 GNDA.n1988 GNDA.n1936 16.0005
R6429 GNDA.n1994 GNDA.n1936 16.0005
R6430 GNDA.n1995 GNDA.n1994 16.0005
R6431 GNDA.n1998 GNDA.n1995 16.0005
R6432 GNDA.n1979 GNDA.n1978 16.0005
R6433 GNDA.n1978 GNDA.n1940 16.0005
R6434 GNDA.n1972 GNDA.n1940 16.0005
R6435 GNDA.n1972 GNDA.n1971 16.0005
R6436 GNDA.n1971 GNDA.n1970 16.0005
R6437 GNDA.n1970 GNDA.n1942 16.0005
R6438 GNDA.n1964 GNDA.n1942 16.0005
R6439 GNDA.n1964 GNDA.n1963 16.0005
R6440 GNDA.n1962 GNDA.n1944 16.0005
R6441 GNDA.n1956 GNDA.n1944 16.0005
R6442 GNDA.n1956 GNDA.n1955 16.0005
R6443 GNDA.n1955 GNDA.n1954 16.0005
R6444 GNDA.n1954 GNDA.n1946 16.0005
R6445 GNDA.n1949 GNDA.n1946 16.0005
R6446 GNDA.n1949 GNDA.n1900 16.0005
R6447 GNDA.n2035 GNDA.n1900 16.0005
R6448 GNDA.n5315 GNDA.n5314 16.0005
R6449 GNDA.n5318 GNDA.n5315 16.0005
R6450 GNDA.n5319 GNDA.n5318 16.0005
R6451 GNDA.n5322 GNDA.n5319 16.0005
R6452 GNDA.n5323 GNDA.n5322 16.0005
R6453 GNDA.n5326 GNDA.n5323 16.0005
R6454 GNDA.n5327 GNDA.n5326 16.0005
R6455 GNDA.n5327 GNDA.n164 16.0005
R6456 GNDA.n5311 GNDA.n5310 16.0005
R6457 GNDA.n5310 GNDA.n5307 16.0005
R6458 GNDA.n5307 GNDA.n5306 16.0005
R6459 GNDA.n5306 GNDA.n5303 16.0005
R6460 GNDA.n5303 GNDA.n5302 16.0005
R6461 GNDA.n5302 GNDA.n5299 16.0005
R6462 GNDA.n5299 GNDA.n5298 16.0005
R6463 GNDA.n5298 GNDA.n5295 16.0005
R6464 GNDA.n5294 GNDA.n5291 16.0005
R6465 GNDA.n5291 GNDA.n5290 16.0005
R6466 GNDA.n5290 GNDA.n5287 16.0005
R6467 GNDA.n5287 GNDA.n5286 16.0005
R6468 GNDA.n5286 GNDA.n5283 16.0005
R6469 GNDA.n5283 GNDA.n5282 16.0005
R6470 GNDA.n5282 GNDA.n5279 16.0005
R6471 GNDA.n5279 GNDA.n5278 16.0005
R6472 GNDA.n5100 GNDA.n5099 16.0005
R6473 GNDA.n5103 GNDA.n5100 16.0005
R6474 GNDA.n5104 GNDA.n5103 16.0005
R6475 GNDA.n5107 GNDA.n5104 16.0005
R6476 GNDA.n5108 GNDA.n5107 16.0005
R6477 GNDA.n5111 GNDA.n5108 16.0005
R6478 GNDA.n5112 GNDA.n5111 16.0005
R6479 GNDA.n5112 GNDA.n5010 16.0005
R6480 GNDA.n5096 GNDA.n5095 16.0005
R6481 GNDA.n5095 GNDA.n5092 16.0005
R6482 GNDA.n5092 GNDA.n5091 16.0005
R6483 GNDA.n5091 GNDA.n5088 16.0005
R6484 GNDA.n5088 GNDA.n5087 16.0005
R6485 GNDA.n5087 GNDA.n5084 16.0005
R6486 GNDA.n5084 GNDA.n5083 16.0005
R6487 GNDA.n5083 GNDA.n5080 16.0005
R6488 GNDA.n5079 GNDA.n5076 16.0005
R6489 GNDA.n5076 GNDA.n5075 16.0005
R6490 GNDA.n5075 GNDA.n5072 16.0005
R6491 GNDA.n5072 GNDA.n5071 16.0005
R6492 GNDA.n5071 GNDA.n5068 16.0005
R6493 GNDA.n5068 GNDA.n5067 16.0005
R6494 GNDA.n5067 GNDA.n5064 16.0005
R6495 GNDA.n5064 GNDA.n5063 16.0005
R6496 GNDA.n2248 GNDA.n2247 16.0005
R6497 GNDA.n2251 GNDA.n2248 16.0005
R6498 GNDA.n2252 GNDA.n2251 16.0005
R6499 GNDA.n2255 GNDA.n2252 16.0005
R6500 GNDA.n2256 GNDA.n2255 16.0005
R6501 GNDA.n2259 GNDA.n2256 16.0005
R6502 GNDA.n2261 GNDA.n2259 16.0005
R6503 GNDA.n2262 GNDA.n2261 16.0005
R6504 GNDA.n2244 GNDA.n2243 16.0005
R6505 GNDA.n2243 GNDA.n2240 16.0005
R6506 GNDA.n2240 GNDA.n2239 16.0005
R6507 GNDA.n2239 GNDA.n2236 16.0005
R6508 GNDA.n2236 GNDA.n2235 16.0005
R6509 GNDA.n2235 GNDA.n2232 16.0005
R6510 GNDA.n2232 GNDA.n2231 16.0005
R6511 GNDA.n2231 GNDA.n2228 16.0005
R6512 GNDA.n2227 GNDA.n2224 16.0005
R6513 GNDA.n2224 GNDA.n2223 16.0005
R6514 GNDA.n2223 GNDA.n2220 16.0005
R6515 GNDA.n2220 GNDA.n2219 16.0005
R6516 GNDA.n2219 GNDA.n2216 16.0005
R6517 GNDA.n2216 GNDA.n2215 16.0005
R6518 GNDA.n2215 GNDA.n2212 16.0005
R6519 GNDA.n2212 GNDA.n2188 16.0005
R6520 GNDA.n5252 GNDA.n5239 16.0005
R6521 GNDA.n5252 GNDA.n5251 16.0005
R6522 GNDA.n5251 GNDA.n5250 16.0005
R6523 GNDA.n5250 GNDA.n5247 16.0005
R6524 GNDA.n5247 GNDA.n5246 16.0005
R6525 GNDA.n5246 GNDA.n5243 16.0005
R6526 GNDA.n5243 GNDA.n5242 16.0005
R6527 GNDA.n5242 GNDA.n5154 16.0005
R6528 GNDA.n5238 GNDA.n5236 16.0005
R6529 GNDA.n5236 GNDA.n5233 16.0005
R6530 GNDA.n5233 GNDA.n5232 16.0005
R6531 GNDA.n5232 GNDA.n5229 16.0005
R6532 GNDA.n5229 GNDA.n5228 16.0005
R6533 GNDA.n5228 GNDA.n5225 16.0005
R6534 GNDA.n5225 GNDA.n5224 16.0005
R6535 GNDA.n5224 GNDA.n5221 16.0005
R6536 GNDA.n5220 GNDA.n5217 16.0005
R6537 GNDA.n5217 GNDA.n5216 16.0005
R6538 GNDA.n5216 GNDA.n5213 16.0005
R6539 GNDA.n5213 GNDA.n5212 16.0005
R6540 GNDA.n5212 GNDA.n5209 16.0005
R6541 GNDA.n5209 GNDA.n5208 16.0005
R6542 GNDA.n5208 GNDA.n5205 16.0005
R6543 GNDA.n5205 GNDA.n5204 16.0005
R6544 GNDA.n5531 GNDA.n5518 16.0005
R6545 GNDA.n5531 GNDA.n5530 16.0005
R6546 GNDA.n5530 GNDA.n5529 16.0005
R6547 GNDA.n5529 GNDA.n5526 16.0005
R6548 GNDA.n5526 GNDA.n5525 16.0005
R6549 GNDA.n5525 GNDA.n5522 16.0005
R6550 GNDA.n5522 GNDA.n5521 16.0005
R6551 GNDA.n5521 GNDA.n57 16.0005
R6552 GNDA.n5517 GNDA.n5515 16.0005
R6553 GNDA.n5515 GNDA.n5512 16.0005
R6554 GNDA.n5512 GNDA.n5511 16.0005
R6555 GNDA.n5511 GNDA.n5508 16.0005
R6556 GNDA.n5508 GNDA.n5507 16.0005
R6557 GNDA.n5507 GNDA.n5504 16.0005
R6558 GNDA.n5504 GNDA.n5503 16.0005
R6559 GNDA.n5503 GNDA.n5500 16.0005
R6560 GNDA.n5499 GNDA.n5496 16.0005
R6561 GNDA.n5496 GNDA.n5495 16.0005
R6562 GNDA.n5495 GNDA.n5492 16.0005
R6563 GNDA.n5492 GNDA.n5491 16.0005
R6564 GNDA.n5491 GNDA.n5488 16.0005
R6565 GNDA.n5488 GNDA.n5487 16.0005
R6566 GNDA.n5487 GNDA.n5484 16.0005
R6567 GNDA.n5484 GNDA.n5483 16.0005
R6568 GNDA.n1786 GNDA.n1785 16.0005
R6569 GNDA.n1787 GNDA.n1786 16.0005
R6570 GNDA.n1787 GNDA.n1737 16.0005
R6571 GNDA.n1793 GNDA.n1737 16.0005
R6572 GNDA.n1794 GNDA.n1793 16.0005
R6573 GNDA.n1795 GNDA.n1794 16.0005
R6574 GNDA.n1795 GNDA.n1735 16.0005
R6575 GNDA.n1801 GNDA.n1735 16.0005
R6576 GNDA.n1779 GNDA.n1739 16.0005
R6577 GNDA.n1779 GNDA.n1778 16.0005
R6578 GNDA.n1778 GNDA.n1777 16.0005
R6579 GNDA.n1777 GNDA.n1741 16.0005
R6580 GNDA.n1771 GNDA.n1741 16.0005
R6581 GNDA.n1771 GNDA.n1770 16.0005
R6582 GNDA.n1770 GNDA.n1769 16.0005
R6583 GNDA.n1769 GNDA.n1743 16.0005
R6584 GNDA.n1763 GNDA.n1762 16.0005
R6585 GNDA.n1762 GNDA.n1761 16.0005
R6586 GNDA.n1761 GNDA.n1745 16.0005
R6587 GNDA.n1756 GNDA.n1745 16.0005
R6588 GNDA.n1756 GNDA.n1755 16.0005
R6589 GNDA.n1755 GNDA.n1754 16.0005
R6590 GNDA.n1754 GNDA.n1749 16.0005
R6591 GNDA.n1749 GNDA.n1748 16.0005
R6592 GNDA.n5438 GNDA.n5437 16.0005
R6593 GNDA.n5441 GNDA.n5438 16.0005
R6594 GNDA.n5442 GNDA.n5441 16.0005
R6595 GNDA.n5445 GNDA.n5442 16.0005
R6596 GNDA.n5446 GNDA.n5445 16.0005
R6597 GNDA.n5449 GNDA.n5446 16.0005
R6598 GNDA.n5451 GNDA.n5449 16.0005
R6599 GNDA.n5452 GNDA.n5451 16.0005
R6600 GNDA.n5434 GNDA.n5433 16.0005
R6601 GNDA.n5433 GNDA.n5430 16.0005
R6602 GNDA.n5430 GNDA.n5429 16.0005
R6603 GNDA.n5429 GNDA.n5426 16.0005
R6604 GNDA.n5426 GNDA.n5425 16.0005
R6605 GNDA.n5425 GNDA.n5422 16.0005
R6606 GNDA.n5422 GNDA.n5421 16.0005
R6607 GNDA.n5421 GNDA.n5418 16.0005
R6608 GNDA.n5417 GNDA.n5414 16.0005
R6609 GNDA.n5414 GNDA.n5413 16.0005
R6610 GNDA.n5413 GNDA.n5410 16.0005
R6611 GNDA.n5410 GNDA.n5409 16.0005
R6612 GNDA.n5409 GNDA.n5406 16.0005
R6613 GNDA.n5406 GNDA.n5405 16.0005
R6614 GNDA.n5405 GNDA.n5402 16.0005
R6615 GNDA.n5402 GNDA.n5401 16.0005
R6616 GNDA.t186 GNDA.t95 15.0244
R6617 GNDA.t61 GNDA.t186 15.0244
R6618 GNDA.t28 GNDA.t236 15.0244
R6619 GNDA.t32 GNDA.t5 14.9259
R6620 GNDA.t31 GNDA.t100 14.9259
R6621 GNDA.t123 GNDA.t56 14.9259
R6622 GNDA.t239 GNDA.t21 14.9259
R6623 GNDA.t41 GNDA.t260 14.9259
R6624 GNDA.t125 GNDA.t133 14.9259
R6625 GNDA.t39 GNDA.t76 14.9259
R6626 GNDA.t119 GNDA.t77 14.9259
R6627 GNDA.n5550 GNDA.n26 14.555
R6628 GNDA.n5271 GNDA.n107 14.555
R6629 GNDA.t284 GNDA.t16 14.4651
R6630 GNDA.t66 GNDA.t282 14.4651
R6631 GNDA.n740 GNDA.n739 14.238
R6632 GNDA.n643 GNDA.n642 14.238
R6633 GNDA.t19 GNDA.t183 13.8109
R6634 GNDA.n4136 GNDA.n4135 13.5941
R6635 GNDA.n3477 GNDA.n3476 13.5941
R6636 GNDA.n4278 GNDA.n479 13.5697
R6637 GNDA.n3389 GNDA.n3388 13.5697
R6638 GNDA.n4061 GNDA.t31 13.4333
R6639 GNDA.t76 GNDA.n634 13.4333
R6640 GNDA.n4057 GNDA.n748 12.8005
R6641 GNDA.n4053 GNDA.n748 12.8005
R6642 GNDA.n4047 GNDA.n750 12.8005
R6643 GNDA.n4051 GNDA.n750 12.8005
R6644 GNDA.n670 GNDA.n663 12.8005
R6645 GNDA.n666 GNDA.n663 12.8005
R6646 GNDA.n730 GNDA.n644 12.8005
R6647 GNDA.n734 GNDA.n644 12.8005
R6648 GNDA.n691 GNDA.n690 12.8005
R6649 GNDA.n690 GNDA.n688 12.8005
R6650 GNDA.n4119 GNDA.n603 12.8005
R6651 GNDA.n4119 GNDA.n604 12.8005
R6652 GNDA.n2042 GNDA.n1896 12.8005
R6653 GNDA.n2046 GNDA.n1896 12.8005
R6654 GNDA.n1927 GNDA.n1926 12.8005
R6655 GNDA.n1926 GNDA.n1920 12.8005
R6656 GNDA.n4970 GNDA.n357 12.8005
R6657 GNDA.n4970 GNDA.n4969 12.8005
R6658 GNDA.t82 GNDA.t284 12.7634
R6659 GNDA.t75 GNDA.t135 12.7634
R6660 GNDA.t135 GNDA.t109 12.7634
R6661 GNDA.t109 GNDA.t17 12.7634
R6662 GNDA.t53 GNDA.t107 12.7634
R6663 GNDA.t83 GNDA.t53 12.7634
R6664 GNDA.t283 GNDA.t83 12.7634
R6665 GNDA.t9 GNDA.t66 12.7634
R6666 GNDA.n4131 GNDA.t195 12.6791
R6667 GNDA.n4280 GNDA.t181 12.6791
R6668 GNDA.n3384 GNDA.t271 12.6791
R6669 GNDA.n3480 GNDA.t264 12.6791
R6670 GNDA.n2068 GNDA.t24 12.0196
R6671 GNDA.t129 GNDA.n2023 12.0196
R6672 GNDA.n2494 GNDA.t93 12.0196
R6673 GNDA.n2399 GNDA.n2396 11.6369
R6674 GNDA.n2402 GNDA.n2399 11.6369
R6675 GNDA.n2414 GNDA.n2402 11.6369
R6676 GNDA.n2414 GNDA.n2413 11.6369
R6677 GNDA.n2413 GNDA.n2412 11.6369
R6678 GNDA.n2412 GNDA.n2403 11.6369
R6679 GNDA.n2406 GNDA.n2403 11.6369
R6680 GNDA.n2406 GNDA.n2405 11.6369
R6681 GNDA.n2405 GNDA.n1451 11.6369
R6682 GNDA.n2538 GNDA.n1451 11.6369
R6683 GNDA.n2438 GNDA.n2388 11.6369
R6684 GNDA.n2438 GNDA.n2437 11.6369
R6685 GNDA.n2437 GNDA.n2436 11.6369
R6686 GNDA.n2436 GNDA.n2390 11.6369
R6687 GNDA.n2431 GNDA.n2390 11.6369
R6688 GNDA.n2431 GNDA.n2430 11.6369
R6689 GNDA.n2430 GNDA.n2429 11.6369
R6690 GNDA.n2429 GNDA.n2393 11.6369
R6691 GNDA.n2424 GNDA.n2393 11.6369
R6692 GNDA.n2424 GNDA.n2423 11.6369
R6693 GNDA.n2423 GNDA.n2422 11.6369
R6694 GNDA.n2114 GNDA.n2113 11.6369
R6695 GNDA.n2115 GNDA.n2114 11.6369
R6696 GNDA.n2115 GNDA.n1686 11.6369
R6697 GNDA.n2121 GNDA.n1686 11.6369
R6698 GNDA.n2122 GNDA.n2121 11.6369
R6699 GNDA.n2123 GNDA.n2122 11.6369
R6700 GNDA.n2123 GNDA.n1684 11.6369
R6701 GNDA.n2128 GNDA.n1684 11.6369
R6702 GNDA.n2129 GNDA.n2128 11.6369
R6703 GNDA.n2129 GNDA.n1682 11.6369
R6704 GNDA.n2135 GNDA.n1682 11.6369
R6705 GNDA.n2180 GNDA.n2176 11.6369
R6706 GNDA.n2321 GNDA.n2180 11.6369
R6707 GNDA.n2321 GNDA.n2320 11.6369
R6708 GNDA.n2320 GNDA.n2319 11.6369
R6709 GNDA.n2319 GNDA.n2181 11.6369
R6710 GNDA.n2314 GNDA.n2181 11.6369
R6711 GNDA.n2314 GNDA.n2313 11.6369
R6712 GNDA.n2313 GNDA.n2312 11.6369
R6713 GNDA.n2312 GNDA.n2183 11.6369
R6714 GNDA.n2306 GNDA.n2183 11.6369
R6715 GNDA.n2349 GNDA.n2348 11.6369
R6716 GNDA.n2348 GNDA.n2345 11.6369
R6717 GNDA.n2345 GNDA.n2344 11.6369
R6718 GNDA.n2344 GNDA.n2341 11.6369
R6719 GNDA.n2341 GNDA.n2340 11.6369
R6720 GNDA.n2340 GNDA.n2337 11.6369
R6721 GNDA.n2337 GNDA.n2336 11.6369
R6722 GNDA.n2336 GNDA.n2333 11.6369
R6723 GNDA.n2333 GNDA.n2332 11.6369
R6724 GNDA.n2332 GNDA.n2329 11.6369
R6725 GNDA.n2329 GNDA.n2328 11.6369
R6726 GNDA.n2152 GNDA.n132 11.6369
R6727 GNDA.n2155 GNDA.n2152 11.6369
R6728 GNDA.n2156 GNDA.n2155 11.6369
R6729 GNDA.n2159 GNDA.n2156 11.6369
R6730 GNDA.n2160 GNDA.n2159 11.6369
R6731 GNDA.n2163 GNDA.n2160 11.6369
R6732 GNDA.n2164 GNDA.n2163 11.6369
R6733 GNDA.n2167 GNDA.n2164 11.6369
R6734 GNDA.n2168 GNDA.n2167 11.6369
R6735 GNDA.n2171 GNDA.n2168 11.6369
R6736 GNDA.n2174 GNDA.n2171 11.6369
R6737 GNDA.n263 GNDA.n262 11.6369
R6738 GNDA.n266 GNDA.n263 11.6369
R6739 GNDA.n267 GNDA.n266 11.6369
R6740 GNDA.n270 GNDA.n267 11.6369
R6741 GNDA.n271 GNDA.n270 11.6369
R6742 GNDA.n274 GNDA.n271 11.6369
R6743 GNDA.n275 GNDA.n274 11.6369
R6744 GNDA.n277 GNDA.n275 11.6369
R6745 GNDA.n277 GNDA.n276 11.6369
R6746 GNDA.n276 GNDA.n228 11.6369
R6747 GNDA.n259 GNDA.n258 11.6369
R6748 GNDA.n258 GNDA.n255 11.6369
R6749 GNDA.n255 GNDA.n254 11.6369
R6750 GNDA.n254 GNDA.n251 11.6369
R6751 GNDA.n251 GNDA.n250 11.6369
R6752 GNDA.n250 GNDA.n247 11.6369
R6753 GNDA.n247 GNDA.n246 11.6369
R6754 GNDA.n246 GNDA.n243 11.6369
R6755 GNDA.n243 GNDA.n242 11.6369
R6756 GNDA.n242 GNDA.n131 11.6369
R6757 GNDA.n5367 GNDA.n131 11.6369
R6758 GNDA.n5147 GNDA.n5146 11.6369
R6759 GNDA.n5146 GNDA.n5145 11.6369
R6760 GNDA.n5145 GNDA.n5144 11.6369
R6761 GNDA.n5144 GNDA.n5142 11.6369
R6762 GNDA.n5142 GNDA.n5139 11.6369
R6763 GNDA.n5139 GNDA.n5138 11.6369
R6764 GNDA.n5138 GNDA.n5135 11.6369
R6765 GNDA.n5135 GNDA.n5134 11.6369
R6766 GNDA.n5134 GNDA.n5131 11.6369
R6767 GNDA.n5131 GNDA.n5130 11.6369
R6768 GNDA.n5009 GNDA.n5008 11.6369
R6769 GNDA.n5008 GNDA.n290 11.6369
R6770 GNDA.n5002 GNDA.n290 11.6369
R6771 GNDA.n5002 GNDA.n5001 11.6369
R6772 GNDA.n5001 GNDA.n5000 11.6369
R6773 GNDA.n5000 GNDA.n294 11.6369
R6774 GNDA.n4994 GNDA.n294 11.6369
R6775 GNDA.n4994 GNDA.n4993 11.6369
R6776 GNDA.n4993 GNDA.n4992 11.6369
R6777 GNDA.n4992 GNDA.n298 11.6369
R6778 GNDA.n4986 GNDA.n298 11.6369
R6779 GNDA.n1834 GNDA.n1833 11.6369
R6780 GNDA.n1837 GNDA.n1834 11.6369
R6781 GNDA.n1838 GNDA.n1837 11.6369
R6782 GNDA.n1841 GNDA.n1838 11.6369
R6783 GNDA.n1842 GNDA.n1841 11.6369
R6784 GNDA.n1845 GNDA.n1842 11.6369
R6785 GNDA.n1846 GNDA.n1845 11.6369
R6786 GNDA.n1849 GNDA.n1846 11.6369
R6787 GNDA.n1850 GNDA.n1849 11.6369
R6788 GNDA.n1853 GNDA.n1850 11.6369
R6789 GNDA.n1828 GNDA.n1802 11.6369
R6790 GNDA.n1828 GNDA.n1827 11.6369
R6791 GNDA.n1827 GNDA.n1826 11.6369
R6792 GNDA.n1826 GNDA.n1804 11.6369
R6793 GNDA.n1821 GNDA.n1804 11.6369
R6794 GNDA.n1821 GNDA.n1820 11.6369
R6795 GNDA.n1820 GNDA.n1819 11.6369
R6796 GNDA.n1819 GNDA.n1807 11.6369
R6797 GNDA.n1814 GNDA.n1807 11.6369
R6798 GNDA.n1814 GNDA.n1813 11.6369
R6799 GNDA.n1813 GNDA.n1812 11.6369
R6800 GNDA.n4928 GNDA.n4927 11.6369
R6801 GNDA.n4927 GNDA.n4926 11.6369
R6802 GNDA.n4926 GNDA.n426 11.6369
R6803 GNDA.n4920 GNDA.n426 11.6369
R6804 GNDA.n4920 GNDA.n4919 11.6369
R6805 GNDA.n4919 GNDA.n92 11.6369
R6806 GNDA.n5374 GNDA.n92 11.6369
R6807 GNDA.n5375 GNDA.n5374 11.6369
R6808 GNDA.n5377 GNDA.n5375 11.6369
R6809 GNDA.n5377 GNDA.n5376 11.6369
R6810 GNDA.n4952 GNDA.n4951 11.6369
R6811 GNDA.n4951 GNDA.n4950 11.6369
R6812 GNDA.n4950 GNDA.n414 11.6369
R6813 GNDA.n4944 GNDA.n414 11.6369
R6814 GNDA.n4944 GNDA.n4943 11.6369
R6815 GNDA.n4943 GNDA.n4942 11.6369
R6816 GNDA.n4942 GNDA.n418 11.6369
R6817 GNDA.n4936 GNDA.n418 11.6369
R6818 GNDA.n4936 GNDA.n4935 11.6369
R6819 GNDA.n4935 GNDA.n4934 11.6369
R6820 GNDA.n4934 GNDA.n422 11.6369
R6821 GNDA.n4984 GNDA.n303 11.6369
R6822 GNDA.n4978 GNDA.n303 11.6369
R6823 GNDA.n4978 GNDA.n4977 11.6369
R6824 GNDA.n4977 GNDA.n4976 11.6369
R6825 GNDA.n4976 GNDA.n353 11.6369
R6826 GNDA.n4967 GNDA.n360 11.6369
R6827 GNDA.n364 GNDA.n360 11.6369
R6828 GNDA.n4960 GNDA.n364 11.6369
R6829 GNDA.n4960 GNDA.n4959 11.6369
R6830 GNDA.n4959 GNDA.n4958 11.6369
R6831 GNDA.t186 GNDA.n99 11.3072
R6832 GNDA.t138 GNDA.t171 11.0892
R6833 GNDA.t158 GNDA.t22 11.0892
R6834 GNDA.t80 GNDA.t73 11.0892
R6835 GNDA.t87 GNDA.t136 11.0892
R6836 GNDA.n2548 GNDA.n2547 10.9846
R6837 GNDA.n2565 GNDA.n1426 10.87
R6838 GNDA.n2562 GNDA.n1429 10.87
R6839 GNDA.n2561 GNDA.n1430 10.87
R6840 GNDA.n2557 GNDA.n1434 10.87
R6841 GNDA.n2556 GNDA.n1435 10.87
R6842 GNDA.n2552 GNDA.n1439 10.87
R6843 GNDA.n2551 GNDA.n1440 10.87
R6844 GNDA.t5 GNDA.n636 10.4483
R6845 GNDA.n636 GNDA.t119 10.4483
R6846 GNDA.n1424 GNDA.t79 9.66779
R6847 GNDA.n4019 GNDA.t124 9.6005
R6848 GNDA.n4019 GNDA.t240 9.6005
R6849 GNDA.n4021 GNDA.t6 9.6005
R6850 GNDA.n4021 GNDA.t101 9.6005
R6851 GNDA.n4023 GNDA.t35 9.6005
R6852 GNDA.n4023 GNDA.t98 9.6005
R6853 GNDA.n4025 GNDA.t30 9.6005
R6854 GNDA.n4025 GNDA.t49 9.6005
R6855 GNDA.n4027 GNDA.t29 9.6005
R6856 GNDA.n4027 GNDA.t48 9.6005
R6857 GNDA.n4029 GNDA.t44 9.6005
R6858 GNDA.n4029 GNDA.t65 9.6005
R6859 GNDA.n4031 GNDA.t122 9.6005
R6860 GNDA.n4031 GNDA.t102 9.6005
R6861 GNDA.n4033 GNDA.t118 9.6005
R6862 GNDA.n4033 GNDA.t58 9.6005
R6863 GNDA.n4035 GNDA.t99 9.6005
R6864 GNDA.n4035 GNDA.t57 9.6005
R6865 GNDA.n4037 GNDA.t45 9.6005
R6866 GNDA.n4037 GNDA.t4 9.6005
R6867 GNDA.n4039 GNDA.t40 9.6005
R6868 GNDA.n4039 GNDA.t120 9.6005
R6869 GNDA.n4041 GNDA.t261 9.6005
R6870 GNDA.n4041 GNDA.t134 9.6005
R6871 GNDA.n710 GNDA.t126 9.6005
R6872 GNDA.n710 GNDA.t64 9.6005
R6873 GNDA.n2512 GNDA.t147 9.6005
R6874 GNDA.n1557 GNDA.t149 9.6005
R6875 GNDA.n2054 GNDA.t153 9.6005
R6876 GNDA.n2063 GNDA.t156 9.6005
R6877 GNDA.n721 GNDA.n720 9.42329
R6878 GNDA.n708 GNDA.n674 9.42293
R6879 GNDA.n4048 GNDA.n4047 9.36264
R6880 GNDA.n4057 GNDA.n4056 9.36264
R6881 GNDA.n667 GNDA.n666 9.36264
R6882 GNDA.n731 GNDA.n730 9.36264
R6883 GNDA.n688 GNDA.n684 9.36264
R6884 GNDA.n605 GNDA.n603 9.36264
R6885 GNDA.n2042 GNDA.n1894 9.36264
R6886 GNDA.n1927 GNDA.n1919 9.36264
R6887 GNDA.n1460 GNDA.n357 9.36264
R6888 GNDA.n4055 GNDA.n748 9.3005
R6889 GNDA.n4054 GNDA.n4053 9.3005
R6890 GNDA.n751 GNDA.n750 9.3005
R6891 GNDA.n4051 GNDA.n4050 9.3005
R6892 GNDA.n668 GNDA.n663 9.3005
R6893 GNDA.n670 GNDA.n669 9.3005
R6894 GNDA.n645 GNDA.n644 9.3005
R6895 GNDA.n734 GNDA.n733 9.3005
R6896 GNDA.n690 GNDA.n685 9.3005
R6897 GNDA.n692 GNDA.n691 9.3005
R6898 GNDA.n4119 GNDA.n4118 9.3005
R6899 GNDA.n4117 GNDA.n604 9.3005
R6900 GNDA.n1896 GNDA.n1895 9.3005
R6901 GNDA.n2047 GNDA.n2046 9.3005
R6902 GNDA.n1926 GNDA.n1925 9.3005
R6903 GNDA.n1924 GNDA.n1920 9.3005
R6904 GNDA.n4970 GNDA.n358 9.3005
R6905 GNDA.n4969 GNDA.n359 9.3005
R6906 GNDA.n2529 GNDA.n2527 8.62751
R6907 GNDA.n5457 GNDA.n26 8.60107
R6908 GNDA.n161 GNDA.n107 8.60107
R6909 GNDA.n1733 GNDA.t232 8.01325
R6910 GNDA.n2069 GNDA.t131 8.01325
R6911 GNDA.t277 GNDA.n2009 8.01325
R6912 GNDA.t36 GNDA.n2495 8.01325
R6913 GNDA.n1868 GNDA.t38 7.01165
R6914 GNDA.t74 GNDA.n2082 7.01165
R6915 GNDA.n2387 GNDA.n2135 6.72373
R6916 GNDA.n2175 GNDA.n2174 6.72373
R6917 GNDA.n5367 GNDA.n5366 6.72373
R6918 GNDA.n4986 GNDA.n4985 6.72373
R6919 GNDA.n1812 GNDA.n1688 6.72373
R6920 GNDA.n4958 GNDA.n365 6.72373
R6921 GNDA.n2388 GNDA.n2387 6.20656
R6922 GNDA.n2113 GNDA.n1688 6.20656
R6923 GNDA.n2349 GNDA.n2175 6.20656
R6924 GNDA.n5366 GNDA.n132 6.20656
R6925 GNDA.n4952 GNDA.n365 6.20656
R6926 GNDA.n4985 GNDA.n4984 6.20656
R6927 GNDA.n4968 GNDA.n353 6.07727
R6928 GNDA.n635 GNDA.t90 6.0279
R6929 GNDA.t42 GNDA.t186 6.01006
R6930 GNDA.n2064 GNDA.n2055 5.81868
R6931 GNDA.n2062 GNDA.n2055 5.81868
R6932 GNDA.n4968 GNDA.n4967 5.5601
R6933 GNDA.n2541 GNDA.n1449 5.51161
R6934 GNDA.n2037 GNDA.n2035 5.51161
R6935 GNDA.n5278 GNDA.n186 5.51161
R6936 GNDA.n5063 GNDA.n5033 5.51161
R6937 GNDA.n2300 GNDA.n2188 5.51161
R6938 GNDA.n5204 GNDA.n5182 5.51161
R6939 GNDA.n5483 GNDA.n5461 5.51161
R6940 GNDA.n1748 GNDA.n1716 5.51161
R6941 GNDA.n5401 GNDA.n5387 5.51161
R6942 GNDA.n2540 GNDA.n2539 5.1717
R6943 GNDA.n2305 GNDA.n2301 5.1717
R6944 GNDA.n5386 GNDA.n87 5.1717
R6945 GNDA.t78 GNDA.t275 5.00847
R6946 GNDA.n2066 GNDA.t95 5.00847
R6947 GNDA.t186 GNDA.t188 5.00847
R6948 GNDA.n2518 GNDA.t61 5.00847
R6949 GNDA.t280 GNDA.t70 5.00847
R6950 GNDA.n5268 GNDA.n5153 4.9157
R6951 GNDA.n5127 GNDA.n5124 4.9157
R6952 GNDA.n1856 GNDA.n1855 4.9157
R6953 GNDA.n665 GNDA.n664 4.663
R6954 GNDA.n732 GNDA.n646 4.663
R6955 GNDA.n694 GNDA.n693 4.663
R6956 GNDA.n4116 GNDA.n606 4.663
R6957 GNDA.n739 GNDA.n735 4.64112
R6958 GNDA.n739 GNDA.n738 4.64112
R6959 GNDA.n642 GNDA.n638 4.64112
R6960 GNDA.n642 GNDA.n641 4.64112
R6961 GNDA.n4726 GNDA.n4725 4.5005
R6962 GNDA.n4564 GNDA.n4563 4.5005
R6963 GNDA.n4671 GNDA.n4670 4.5005
R6964 GNDA.n4675 GNDA.n4672 4.5005
R6965 GNDA.n4676 GNDA.n4669 4.5005
R6966 GNDA.n4680 GNDA.n4679 4.5005
R6967 GNDA.n4681 GNDA.n4668 4.5005
R6968 GNDA.n4685 GNDA.n4682 4.5005
R6969 GNDA.n4686 GNDA.n4667 4.5005
R6970 GNDA.n4690 GNDA.n4689 4.5005
R6971 GNDA.n4691 GNDA.n4666 4.5005
R6972 GNDA.n4695 GNDA.n4692 4.5005
R6973 GNDA.n4696 GNDA.n4665 4.5005
R6974 GNDA.n4700 GNDA.n4699 4.5005
R6975 GNDA.n4701 GNDA.n4664 4.5005
R6976 GNDA.n4705 GNDA.n4702 4.5005
R6977 GNDA.n4706 GNDA.n4663 4.5005
R6978 GNDA.n4710 GNDA.n4709 4.5005
R6979 GNDA.n4711 GNDA.n4662 4.5005
R6980 GNDA.n4715 GNDA.n4712 4.5005
R6981 GNDA.n4716 GNDA.n4661 4.5005
R6982 GNDA.n4720 GNDA.n4719 4.5005
R6983 GNDA.n4591 GNDA.n4590 4.5005
R6984 GNDA.n4594 GNDA.n4593 4.5005
R6985 GNDA.n4595 GNDA.n4589 4.5005
R6986 GNDA.n4599 GNDA.n4596 4.5005
R6987 GNDA.n4600 GNDA.n4588 4.5005
R6988 GNDA.n4604 GNDA.n4603 4.5005
R6989 GNDA.n4605 GNDA.n4587 4.5005
R6990 GNDA.n4609 GNDA.n4606 4.5005
R6991 GNDA.n4610 GNDA.n4586 4.5005
R6992 GNDA.n4614 GNDA.n4613 4.5005
R6993 GNDA.n4615 GNDA.n4585 4.5005
R6994 GNDA.n4619 GNDA.n4616 4.5005
R6995 GNDA.n4620 GNDA.n4584 4.5005
R6996 GNDA.n4624 GNDA.n4623 4.5005
R6997 GNDA.n4625 GNDA.n4583 4.5005
R6998 GNDA.n4629 GNDA.n4626 4.5005
R6999 GNDA.n4630 GNDA.n4582 4.5005
R7000 GNDA.n4634 GNDA.n4633 4.5005
R7001 GNDA.n4635 GNDA.n4581 4.5005
R7002 GNDA.n4639 GNDA.n4636 4.5005
R7003 GNDA.n4640 GNDA.n4580 4.5005
R7004 GNDA.n4644 GNDA.n4643 4.5005
R7005 GNDA.n4552 GNDA.n4551 4.5005
R7006 GNDA.n4473 GNDA.n4472 4.5005
R7007 GNDA.n4495 GNDA.n4474 4.5005
R7008 GNDA.n4496 GNDA.n4475 4.5005
R7009 GNDA.n4497 GNDA.n4476 4.5005
R7010 GNDA.n4498 GNDA.n4477 4.5005
R7011 GNDA.n4499 GNDA.n4478 4.5005
R7012 GNDA.n4500 GNDA.n4479 4.5005
R7013 GNDA.n4501 GNDA.n4480 4.5005
R7014 GNDA.n4502 GNDA.n4481 4.5005
R7015 GNDA.n4503 GNDA.n4482 4.5005
R7016 GNDA.n4504 GNDA.n4483 4.5005
R7017 GNDA.n4505 GNDA.n4484 4.5005
R7018 GNDA.n4506 GNDA.n4485 4.5005
R7019 GNDA.n4507 GNDA.n4486 4.5005
R7020 GNDA.n4508 GNDA.n4487 4.5005
R7021 GNDA.n4509 GNDA.n4488 4.5005
R7022 GNDA.n4510 GNDA.n4489 4.5005
R7023 GNDA.n4511 GNDA.n4490 4.5005
R7024 GNDA.n4512 GNDA.n4491 4.5005
R7025 GNDA.n4513 GNDA.n4492 4.5005
R7026 GNDA.n4514 GNDA.n4493 4.5005
R7027 GNDA.n4751 GNDA.n4750 4.5005
R7028 GNDA.n4754 GNDA.n4753 4.5005
R7029 GNDA.n4755 GNDA.n4468 4.5005
R7030 GNDA.n4759 GNDA.n4756 4.5005
R7031 GNDA.n4760 GNDA.n4467 4.5005
R7032 GNDA.n4764 GNDA.n4763 4.5005
R7033 GNDA.n4765 GNDA.n4466 4.5005
R7034 GNDA.n4769 GNDA.n4766 4.5005
R7035 GNDA.n4770 GNDA.n4465 4.5005
R7036 GNDA.n4774 GNDA.n4773 4.5005
R7037 GNDA.n4775 GNDA.n4464 4.5005
R7038 GNDA.n4779 GNDA.n4776 4.5005
R7039 GNDA.n4780 GNDA.n4463 4.5005
R7040 GNDA.n4784 GNDA.n4783 4.5005
R7041 GNDA.n4785 GNDA.n4462 4.5005
R7042 GNDA.n4789 GNDA.n4786 4.5005
R7043 GNDA.n4790 GNDA.n4461 4.5005
R7044 GNDA.n4794 GNDA.n4793 4.5005
R7045 GNDA.n4795 GNDA.n4460 4.5005
R7046 GNDA.n4799 GNDA.n4796 4.5005
R7047 GNDA.n4800 GNDA.n4459 4.5005
R7048 GNDA.n4804 GNDA.n4803 4.5005
R7049 GNDA.n4274 GNDA.n4273 4.5005
R7050 GNDA.n484 GNDA.n483 4.5005
R7051 GNDA.n4219 GNDA.n4218 4.5005
R7052 GNDA.n4223 GNDA.n4220 4.5005
R7053 GNDA.n4224 GNDA.n4217 4.5005
R7054 GNDA.n4228 GNDA.n4227 4.5005
R7055 GNDA.n4229 GNDA.n4216 4.5005
R7056 GNDA.n4233 GNDA.n4230 4.5005
R7057 GNDA.n4234 GNDA.n4215 4.5005
R7058 GNDA.n4238 GNDA.n4237 4.5005
R7059 GNDA.n4239 GNDA.n4214 4.5005
R7060 GNDA.n4243 GNDA.n4240 4.5005
R7061 GNDA.n4244 GNDA.n4213 4.5005
R7062 GNDA.n4248 GNDA.n4247 4.5005
R7063 GNDA.n4249 GNDA.n4212 4.5005
R7064 GNDA.n4253 GNDA.n4250 4.5005
R7065 GNDA.n4254 GNDA.n4211 4.5005
R7066 GNDA.n4258 GNDA.n4257 4.5005
R7067 GNDA.n4259 GNDA.n4210 4.5005
R7068 GNDA.n4263 GNDA.n4260 4.5005
R7069 GNDA.n4264 GNDA.n4209 4.5005
R7070 GNDA.n4268 GNDA.n4267 4.5005
R7071 GNDA.n4875 GNDA.n4874 4.5005
R7072 GNDA.n444 GNDA.n443 4.5005
R7073 GNDA.n4820 GNDA.n4819 4.5005
R7074 GNDA.n4824 GNDA.n4821 4.5005
R7075 GNDA.n4825 GNDA.n4818 4.5005
R7076 GNDA.n4829 GNDA.n4828 4.5005
R7077 GNDA.n4830 GNDA.n4817 4.5005
R7078 GNDA.n4834 GNDA.n4831 4.5005
R7079 GNDA.n4835 GNDA.n4816 4.5005
R7080 GNDA.n4839 GNDA.n4838 4.5005
R7081 GNDA.n4840 GNDA.n4815 4.5005
R7082 GNDA.n4844 GNDA.n4841 4.5005
R7083 GNDA.n4845 GNDA.n4814 4.5005
R7084 GNDA.n4849 GNDA.n4848 4.5005
R7085 GNDA.n4850 GNDA.n4813 4.5005
R7086 GNDA.n4854 GNDA.n4851 4.5005
R7087 GNDA.n4855 GNDA.n4812 4.5005
R7088 GNDA.n4859 GNDA.n4858 4.5005
R7089 GNDA.n4860 GNDA.n4811 4.5005
R7090 GNDA.n4864 GNDA.n4861 4.5005
R7091 GNDA.n4865 GNDA.n4810 4.5005
R7092 GNDA.n4869 GNDA.n4868 4.5005
R7093 GNDA.n4376 GNDA.n4375 4.5005
R7094 GNDA.n4379 GNDA.n4378 4.5005
R7095 GNDA.n4380 GNDA.n470 4.5005
R7096 GNDA.n4384 GNDA.n4381 4.5005
R7097 GNDA.n4385 GNDA.n469 4.5005
R7098 GNDA.n4389 GNDA.n4388 4.5005
R7099 GNDA.n4390 GNDA.n468 4.5005
R7100 GNDA.n4394 GNDA.n4391 4.5005
R7101 GNDA.n4395 GNDA.n467 4.5005
R7102 GNDA.n4399 GNDA.n4398 4.5005
R7103 GNDA.n4400 GNDA.n466 4.5005
R7104 GNDA.n4404 GNDA.n4401 4.5005
R7105 GNDA.n4405 GNDA.n465 4.5005
R7106 GNDA.n4409 GNDA.n4408 4.5005
R7107 GNDA.n4410 GNDA.n464 4.5005
R7108 GNDA.n4414 GNDA.n4411 4.5005
R7109 GNDA.n4415 GNDA.n463 4.5005
R7110 GNDA.n4419 GNDA.n4418 4.5005
R7111 GNDA.n4420 GNDA.n462 4.5005
R7112 GNDA.n4424 GNDA.n4421 4.5005
R7113 GNDA.n4425 GNDA.n461 4.5005
R7114 GNDA.n4429 GNDA.n4428 4.5005
R7115 GNDA.n4364 GNDA.n4363 4.5005
R7116 GNDA.n4285 GNDA.n4284 4.5005
R7117 GNDA.n4307 GNDA.n4286 4.5005
R7118 GNDA.n4308 GNDA.n4287 4.5005
R7119 GNDA.n4309 GNDA.n4288 4.5005
R7120 GNDA.n4310 GNDA.n4289 4.5005
R7121 GNDA.n4311 GNDA.n4290 4.5005
R7122 GNDA.n4312 GNDA.n4291 4.5005
R7123 GNDA.n4313 GNDA.n4292 4.5005
R7124 GNDA.n4314 GNDA.n4293 4.5005
R7125 GNDA.n4315 GNDA.n4294 4.5005
R7126 GNDA.n4316 GNDA.n4295 4.5005
R7127 GNDA.n4317 GNDA.n4296 4.5005
R7128 GNDA.n4318 GNDA.n4297 4.5005
R7129 GNDA.n4319 GNDA.n4298 4.5005
R7130 GNDA.n4320 GNDA.n4299 4.5005
R7131 GNDA.n4321 GNDA.n4300 4.5005
R7132 GNDA.n4322 GNDA.n4301 4.5005
R7133 GNDA.n4323 GNDA.n4302 4.5005
R7134 GNDA.n4324 GNDA.n4303 4.5005
R7135 GNDA.n4325 GNDA.n4304 4.5005
R7136 GNDA.n4326 GNDA.n4305 4.5005
R7137 GNDA.n4139 GNDA.n4138 4.5005
R7138 GNDA.n4142 GNDA.n4141 4.5005
R7139 GNDA.n4143 GNDA.n510 4.5005
R7140 GNDA.n4147 GNDA.n4144 4.5005
R7141 GNDA.n4148 GNDA.n509 4.5005
R7142 GNDA.n4152 GNDA.n4151 4.5005
R7143 GNDA.n4153 GNDA.n508 4.5005
R7144 GNDA.n4157 GNDA.n4154 4.5005
R7145 GNDA.n4158 GNDA.n507 4.5005
R7146 GNDA.n4162 GNDA.n4161 4.5005
R7147 GNDA.n4163 GNDA.n506 4.5005
R7148 GNDA.n4167 GNDA.n4164 4.5005
R7149 GNDA.n4168 GNDA.n505 4.5005
R7150 GNDA.n4172 GNDA.n4171 4.5005
R7151 GNDA.n4173 GNDA.n504 4.5005
R7152 GNDA.n4177 GNDA.n4174 4.5005
R7153 GNDA.n4178 GNDA.n503 4.5005
R7154 GNDA.n4182 GNDA.n4181 4.5005
R7155 GNDA.n4183 GNDA.n502 4.5005
R7156 GNDA.n4187 GNDA.n4184 4.5005
R7157 GNDA.n4188 GNDA.n501 4.5005
R7158 GNDA.n4192 GNDA.n4191 4.5005
R7159 GNDA.n3987 GNDA.n3986 4.5005
R7160 GNDA.n3985 GNDA.n773 4.5005
R7161 GNDA.n3984 GNDA.n3983 4.5005
R7162 GNDA.n3982 GNDA.n777 4.5005
R7163 GNDA.n3981 GNDA.n3980 4.5005
R7164 GNDA.n3979 GNDA.n778 4.5005
R7165 GNDA.n3978 GNDA.n3977 4.5005
R7166 GNDA.n3976 GNDA.n782 4.5005
R7167 GNDA.n3975 GNDA.n3974 4.5005
R7168 GNDA.n3973 GNDA.n783 4.5005
R7169 GNDA.n3972 GNDA.n3971 4.5005
R7170 GNDA.n3970 GNDA.n787 4.5005
R7171 GNDA.n3969 GNDA.n3968 4.5005
R7172 GNDA.n3967 GNDA.n788 4.5005
R7173 GNDA.n3966 GNDA.n3965 4.5005
R7174 GNDA.n3964 GNDA.n792 4.5005
R7175 GNDA.n3963 GNDA.n3962 4.5005
R7176 GNDA.n3961 GNDA.n793 4.5005
R7177 GNDA.n3960 GNDA.n3959 4.5005
R7178 GNDA.n3958 GNDA.n797 4.5005
R7179 GNDA.n3957 GNDA.n3956 4.5005
R7180 GNDA.n3955 GNDA.n798 4.5005
R7181 GNDA.n771 GNDA.n762 4.5005
R7182 GNDA.n769 GNDA.n765 4.5005
R7183 GNDA.n770 GNDA.n764 4.5005
R7184 GNDA.n770 GNDA.n769 4.5005
R7185 GNDA.n4050 GNDA.n4049 4.5005
R7186 GNDA.n4054 GNDA.n749 4.5005
R7187 GNDA.n754 GNDA.n753 4.5005
R7188 GNDA.n757 GNDA.n756 4.5005
R7189 GNDA.n3572 GNDA.n3571 4.5005
R7190 GNDA.n3575 GNDA.n3574 4.5005
R7191 GNDA.n3576 GNDA.n3568 4.5005
R7192 GNDA.n3578 GNDA.n3577 4.5005
R7193 GNDA.n3579 GNDA.n3567 4.5005
R7194 GNDA.n3583 GNDA.n3582 4.5005
R7195 GNDA.n3584 GNDA.n3564 4.5005
R7196 GNDA.n3586 GNDA.n3585 4.5005
R7197 GNDA.n3587 GNDA.n3563 4.5005
R7198 GNDA.n3591 GNDA.n3590 4.5005
R7199 GNDA.n3592 GNDA.n3560 4.5005
R7200 GNDA.n3594 GNDA.n3593 4.5005
R7201 GNDA.n3595 GNDA.n3559 4.5005
R7202 GNDA.n3599 GNDA.n3598 4.5005
R7203 GNDA.n3600 GNDA.n3556 4.5005
R7204 GNDA.n3602 GNDA.n3601 4.5005
R7205 GNDA.n3603 GNDA.n3555 4.5005
R7206 GNDA.n3607 GNDA.n3606 4.5005
R7207 GNDA.n3608 GNDA.n3552 4.5005
R7208 GNDA.n3610 GNDA.n3609 4.5005
R7209 GNDA.n3611 GNDA.n3551 4.5005
R7210 GNDA.n3615 GNDA.n3614 4.5005
R7211 GNDA.n3888 GNDA.n3887 4.5005
R7212 GNDA.n3891 GNDA.n3890 4.5005
R7213 GNDA.n3892 GNDA.n834 4.5005
R7214 GNDA.n3894 GNDA.n3893 4.5005
R7215 GNDA.n3895 GNDA.n833 4.5005
R7216 GNDA.n3899 GNDA.n3898 4.5005
R7217 GNDA.n3900 GNDA.n830 4.5005
R7218 GNDA.n3902 GNDA.n3901 4.5005
R7219 GNDA.n3903 GNDA.n829 4.5005
R7220 GNDA.n3907 GNDA.n3906 4.5005
R7221 GNDA.n3908 GNDA.n826 4.5005
R7222 GNDA.n3910 GNDA.n3909 4.5005
R7223 GNDA.n3911 GNDA.n825 4.5005
R7224 GNDA.n3915 GNDA.n3914 4.5005
R7225 GNDA.n3916 GNDA.n822 4.5005
R7226 GNDA.n3918 GNDA.n3917 4.5005
R7227 GNDA.n3919 GNDA.n821 4.5005
R7228 GNDA.n3923 GNDA.n3922 4.5005
R7229 GNDA.n3924 GNDA.n818 4.5005
R7230 GNDA.n3926 GNDA.n3925 4.5005
R7231 GNDA.n3927 GNDA.n817 4.5005
R7232 GNDA.n3931 GNDA.n3930 4.5005
R7233 GNDA.n921 GNDA.n920 4.5005
R7234 GNDA.n919 GNDA.n841 4.5005
R7235 GNDA.n918 GNDA.n917 4.5005
R7236 GNDA.n916 GNDA.n846 4.5005
R7237 GNDA.n915 GNDA.n914 4.5005
R7238 GNDA.n913 GNDA.n847 4.5005
R7239 GNDA.n912 GNDA.n911 4.5005
R7240 GNDA.n910 GNDA.n854 4.5005
R7241 GNDA.n909 GNDA.n908 4.5005
R7242 GNDA.n907 GNDA.n855 4.5005
R7243 GNDA.n906 GNDA.n905 4.5005
R7244 GNDA.n904 GNDA.n862 4.5005
R7245 GNDA.n903 GNDA.n902 4.5005
R7246 GNDA.n901 GNDA.n863 4.5005
R7247 GNDA.n900 GNDA.n899 4.5005
R7248 GNDA.n898 GNDA.n870 4.5005
R7249 GNDA.n897 GNDA.n896 4.5005
R7250 GNDA.n895 GNDA.n871 4.5005
R7251 GNDA.n894 GNDA.n893 4.5005
R7252 GNDA.n892 GNDA.n878 4.5005
R7253 GNDA.n891 GNDA.n890 4.5005
R7254 GNDA.n889 GNDA.n879 4.5005
R7255 GNDA.n3676 GNDA.n925 4.5005
R7256 GNDA.n3679 GNDA.n3678 4.5005
R7257 GNDA.n3680 GNDA.n3673 4.5005
R7258 GNDA.n3682 GNDA.n3681 4.5005
R7259 GNDA.n3683 GNDA.n3672 4.5005
R7260 GNDA.n3687 GNDA.n3686 4.5005
R7261 GNDA.n3688 GNDA.n3669 4.5005
R7262 GNDA.n3690 GNDA.n3689 4.5005
R7263 GNDA.n3691 GNDA.n3668 4.5005
R7264 GNDA.n3695 GNDA.n3694 4.5005
R7265 GNDA.n3696 GNDA.n3665 4.5005
R7266 GNDA.n3698 GNDA.n3697 4.5005
R7267 GNDA.n3699 GNDA.n3664 4.5005
R7268 GNDA.n3703 GNDA.n3702 4.5005
R7269 GNDA.n3704 GNDA.n3661 4.5005
R7270 GNDA.n3706 GNDA.n3705 4.5005
R7271 GNDA.n3707 GNDA.n3660 4.5005
R7272 GNDA.n3711 GNDA.n3710 4.5005
R7273 GNDA.n3712 GNDA.n3657 4.5005
R7274 GNDA.n3714 GNDA.n3713 4.5005
R7275 GNDA.n3715 GNDA.n3656 4.5005
R7276 GNDA.n3719 GNDA.n3718 4.5005
R7277 GNDA.n3745 GNDA.n929 4.5005
R7278 GNDA.n3748 GNDA.n3747 4.5005
R7279 GNDA.n3749 GNDA.n3742 4.5005
R7280 GNDA.n3751 GNDA.n3750 4.5005
R7281 GNDA.n3752 GNDA.n3741 4.5005
R7282 GNDA.n3756 GNDA.n3755 4.5005
R7283 GNDA.n3757 GNDA.n3738 4.5005
R7284 GNDA.n3759 GNDA.n3758 4.5005
R7285 GNDA.n3760 GNDA.n3737 4.5005
R7286 GNDA.n3764 GNDA.n3763 4.5005
R7287 GNDA.n3765 GNDA.n3734 4.5005
R7288 GNDA.n3767 GNDA.n3766 4.5005
R7289 GNDA.n3768 GNDA.n3733 4.5005
R7290 GNDA.n3772 GNDA.n3771 4.5005
R7291 GNDA.n3773 GNDA.n3730 4.5005
R7292 GNDA.n3775 GNDA.n3774 4.5005
R7293 GNDA.n3776 GNDA.n3729 4.5005
R7294 GNDA.n3780 GNDA.n3779 4.5005
R7295 GNDA.n3781 GNDA.n3726 4.5005
R7296 GNDA.n3783 GNDA.n3782 4.5005
R7297 GNDA.n3784 GNDA.n3725 4.5005
R7298 GNDA.n3788 GNDA.n3787 4.5005
R7299 GNDA.n3868 GNDA.n3866 4.5005
R7300 GNDA.n3870 GNDA.n3869 4.5005
R7301 GNDA.n3869 GNDA.n3868 4.5005
R7302 GNDA.n3873 GNDA.n3871 4.5005
R7303 GNDA.n3875 GNDA.n3874 4.5005
R7304 GNDA.n3874 GNDA.n3873 4.5005
R7305 GNDA.n3878 GNDA.n3876 4.5005
R7306 GNDA.n3880 GNDA.n3879 4.5005
R7307 GNDA.n3879 GNDA.n3878 4.5005
R7308 GNDA.n3885 GNDA.n3881 4.5005
R7309 GNDA.n3886 GNDA.n772 4.5005
R7310 GNDA.n3886 GNDA.n3885 4.5005
R7311 GNDA.n932 GNDA.n931 4.5005
R7312 GNDA.n3859 GNDA.n3858 4.5005
R7313 GNDA.n937 GNDA.n936 4.5005
R7314 GNDA.n3804 GNDA.n3803 4.5005
R7315 GNDA.n3808 GNDA.n3805 4.5005
R7316 GNDA.n3809 GNDA.n3802 4.5005
R7317 GNDA.n3813 GNDA.n3812 4.5005
R7318 GNDA.n3814 GNDA.n3801 4.5005
R7319 GNDA.n3818 GNDA.n3815 4.5005
R7320 GNDA.n3819 GNDA.n3800 4.5005
R7321 GNDA.n3823 GNDA.n3822 4.5005
R7322 GNDA.n3824 GNDA.n3799 4.5005
R7323 GNDA.n3828 GNDA.n3825 4.5005
R7324 GNDA.n3829 GNDA.n3798 4.5005
R7325 GNDA.n3833 GNDA.n3832 4.5005
R7326 GNDA.n3834 GNDA.n3797 4.5005
R7327 GNDA.n3838 GNDA.n3835 4.5005
R7328 GNDA.n3839 GNDA.n3796 4.5005
R7329 GNDA.n3843 GNDA.n3842 4.5005
R7330 GNDA.n3844 GNDA.n3795 4.5005
R7331 GNDA.n3848 GNDA.n3845 4.5005
R7332 GNDA.n3849 GNDA.n3794 4.5005
R7333 GNDA.n3853 GNDA.n3852 4.5005
R7334 GNDA.n3475 GNDA.n3474 4.5005
R7335 GNDA.n3473 GNDA.n3395 4.5005
R7336 GNDA.n3472 GNDA.n3471 4.5005
R7337 GNDA.n3470 GNDA.n3400 4.5005
R7338 GNDA.n3469 GNDA.n3468 4.5005
R7339 GNDA.n3467 GNDA.n3401 4.5005
R7340 GNDA.n3466 GNDA.n3465 4.5005
R7341 GNDA.n3464 GNDA.n3408 4.5005
R7342 GNDA.n3463 GNDA.n3462 4.5005
R7343 GNDA.n3461 GNDA.n3409 4.5005
R7344 GNDA.n3460 GNDA.n3459 4.5005
R7345 GNDA.n3458 GNDA.n3416 4.5005
R7346 GNDA.n3457 GNDA.n3456 4.5005
R7347 GNDA.n3455 GNDA.n3417 4.5005
R7348 GNDA.n3454 GNDA.n3453 4.5005
R7349 GNDA.n3452 GNDA.n3424 4.5005
R7350 GNDA.n3451 GNDA.n3450 4.5005
R7351 GNDA.n3449 GNDA.n3425 4.5005
R7352 GNDA.n3448 GNDA.n3447 4.5005
R7353 GNDA.n3446 GNDA.n3432 4.5005
R7354 GNDA.n3445 GNDA.n3444 4.5005
R7355 GNDA.n3443 GNDA.n3433 4.5005
R7356 GNDA.n3490 GNDA.n3489 4.5005
R7357 GNDA.n3493 GNDA.n3492 4.5005
R7358 GNDA.n3494 GNDA.n971 4.5005
R7359 GNDA.n3496 GNDA.n3495 4.5005
R7360 GNDA.n3497 GNDA.n970 4.5005
R7361 GNDA.n3501 GNDA.n3500 4.5005
R7362 GNDA.n3502 GNDA.n967 4.5005
R7363 GNDA.n3504 GNDA.n3503 4.5005
R7364 GNDA.n3505 GNDA.n966 4.5005
R7365 GNDA.n3509 GNDA.n3508 4.5005
R7366 GNDA.n3510 GNDA.n963 4.5005
R7367 GNDA.n3512 GNDA.n3511 4.5005
R7368 GNDA.n3513 GNDA.n962 4.5005
R7369 GNDA.n3517 GNDA.n3516 4.5005
R7370 GNDA.n3518 GNDA.n959 4.5005
R7371 GNDA.n3520 GNDA.n3519 4.5005
R7372 GNDA.n3521 GNDA.n958 4.5005
R7373 GNDA.n3525 GNDA.n3524 4.5005
R7374 GNDA.n3526 GNDA.n955 4.5005
R7375 GNDA.n3528 GNDA.n3527 4.5005
R7376 GNDA.n3529 GNDA.n954 4.5005
R7377 GNDA.n3533 GNDA.n3532 4.5005
R7378 GNDA.n2811 GNDA.n979 4.5005
R7379 GNDA.n2814 GNDA.n2813 4.5005
R7380 GNDA.n2815 GNDA.n2808 4.5005
R7381 GNDA.n2817 GNDA.n2816 4.5005
R7382 GNDA.n2818 GNDA.n2807 4.5005
R7383 GNDA.n2822 GNDA.n2821 4.5005
R7384 GNDA.n2823 GNDA.n2804 4.5005
R7385 GNDA.n2825 GNDA.n2824 4.5005
R7386 GNDA.n2826 GNDA.n2803 4.5005
R7387 GNDA.n2830 GNDA.n2829 4.5005
R7388 GNDA.n2831 GNDA.n2800 4.5005
R7389 GNDA.n2833 GNDA.n2832 4.5005
R7390 GNDA.n2834 GNDA.n2799 4.5005
R7391 GNDA.n2838 GNDA.n2837 4.5005
R7392 GNDA.n2839 GNDA.n2796 4.5005
R7393 GNDA.n2841 GNDA.n2840 4.5005
R7394 GNDA.n2842 GNDA.n2795 4.5005
R7395 GNDA.n2846 GNDA.n2845 4.5005
R7396 GNDA.n2847 GNDA.n2792 4.5005
R7397 GNDA.n2849 GNDA.n2848 4.5005
R7398 GNDA.n2850 GNDA.n2791 4.5005
R7399 GNDA.n2854 GNDA.n2853 4.5005
R7400 GNDA.n4904 GNDA.n4903 4.5005
R7401 GNDA.n4911 GNDA.n433 4.5005
R7402 GNDA.n4910 GNDA.n4909 4.5005
R7403 GNDA.n4911 GNDA.n4910 4.5005
R7404 GNDA.n669 GNDA.n665 4.5005
R7405 GNDA.n733 GNDA.n732 4.5005
R7406 GNDA.n4096 GNDA.n4095 4.5005
R7407 GNDA.n4101 GNDA.n4087 4.5005
R7408 GNDA.n4103 GNDA.n4102 4.5005
R7409 GNDA.n4102 GNDA.n4101 4.5005
R7410 GNDA.n694 GNDA.n692 4.5005
R7411 GNDA.n4117 GNDA.n4116 4.5005
R7412 GNDA.n610 GNDA.n608 4.5005
R7413 GNDA.n613 GNDA.n612 4.5005
R7414 GNDA.n660 GNDA.n648 4.5005
R7415 GNDA.n651 GNDA.n650 4.5005
R7416 GNDA.n718 GNDA.n712 4.5005
R7417 GNDA.n715 GNDA.n609 4.5005
R7418 GNDA.n718 GNDA.n609 4.5005
R7419 GNDA.n682 GNDA.n681 4.5005
R7420 GNDA.n701 GNDA.n695 4.5005
R7421 GNDA.n701 GNDA.n700 4.5005
R7422 GNDA.n700 GNDA.n697 4.5005
R7423 GNDA.n4086 GNDA.n4085 4.5005
R7424 GNDA.n4085 GNDA.n4084 4.5005
R7425 GNDA.n4084 GNDA.n622 4.5005
R7426 GNDA.n4081 GNDA.n624 4.5005
R7427 GNDA.n4081 GNDA.n4080 4.5005
R7428 GNDA.n4080 GNDA.n625 4.5005
R7429 GNDA.n1014 GNDA.n1013 4.5005
R7430 GNDA.n1020 GNDA.n996 4.5005
R7431 GNDA.n1021 GNDA.n995 4.5005
R7432 GNDA.n1021 GNDA.n1020 4.5005
R7433 GNDA.n4071 GNDA.n627 4.5005
R7434 GNDA.n4073 GNDA.n4072 4.5005
R7435 GNDA.n4072 GNDA.n4071 4.5005
R7436 GNDA.n2880 GNDA.n983 4.5005
R7437 GNDA.n2883 GNDA.n2882 4.5005
R7438 GNDA.n2884 GNDA.n2877 4.5005
R7439 GNDA.n2886 GNDA.n2885 4.5005
R7440 GNDA.n2887 GNDA.n2876 4.5005
R7441 GNDA.n2891 GNDA.n2890 4.5005
R7442 GNDA.n2892 GNDA.n2873 4.5005
R7443 GNDA.n2894 GNDA.n2893 4.5005
R7444 GNDA.n2895 GNDA.n2872 4.5005
R7445 GNDA.n2899 GNDA.n2898 4.5005
R7446 GNDA.n2900 GNDA.n2869 4.5005
R7447 GNDA.n2902 GNDA.n2901 4.5005
R7448 GNDA.n2903 GNDA.n2868 4.5005
R7449 GNDA.n2907 GNDA.n2906 4.5005
R7450 GNDA.n2908 GNDA.n2865 4.5005
R7451 GNDA.n2910 GNDA.n2909 4.5005
R7452 GNDA.n2911 GNDA.n2864 4.5005
R7453 GNDA.n2915 GNDA.n2914 4.5005
R7454 GNDA.n2916 GNDA.n2861 4.5005
R7455 GNDA.n2918 GNDA.n2917 4.5005
R7456 GNDA.n2919 GNDA.n2860 4.5005
R7457 GNDA.n2923 GNDA.n2922 4.5005
R7458 GNDA.n2949 GNDA.n987 4.5005
R7459 GNDA.n2952 GNDA.n2951 4.5005
R7460 GNDA.n2953 GNDA.n2946 4.5005
R7461 GNDA.n2955 GNDA.n2954 4.5005
R7462 GNDA.n2956 GNDA.n2945 4.5005
R7463 GNDA.n2960 GNDA.n2959 4.5005
R7464 GNDA.n2961 GNDA.n2942 4.5005
R7465 GNDA.n2963 GNDA.n2962 4.5005
R7466 GNDA.n2964 GNDA.n2941 4.5005
R7467 GNDA.n2968 GNDA.n2967 4.5005
R7468 GNDA.n2969 GNDA.n2938 4.5005
R7469 GNDA.n2971 GNDA.n2970 4.5005
R7470 GNDA.n2972 GNDA.n2937 4.5005
R7471 GNDA.n2976 GNDA.n2975 4.5005
R7472 GNDA.n2977 GNDA.n2934 4.5005
R7473 GNDA.n2979 GNDA.n2978 4.5005
R7474 GNDA.n2980 GNDA.n2933 4.5005
R7475 GNDA.n2984 GNDA.n2983 4.5005
R7476 GNDA.n2985 GNDA.n2930 4.5005
R7477 GNDA.n2987 GNDA.n2986 4.5005
R7478 GNDA.n2988 GNDA.n2929 4.5005
R7479 GNDA.n2992 GNDA.n2991 4.5005
R7480 GNDA.n3018 GNDA.n991 4.5005
R7481 GNDA.n3021 GNDA.n3020 4.5005
R7482 GNDA.n3022 GNDA.n3015 4.5005
R7483 GNDA.n3024 GNDA.n3023 4.5005
R7484 GNDA.n3025 GNDA.n3014 4.5005
R7485 GNDA.n3029 GNDA.n3028 4.5005
R7486 GNDA.n3030 GNDA.n3011 4.5005
R7487 GNDA.n3032 GNDA.n3031 4.5005
R7488 GNDA.n3033 GNDA.n3010 4.5005
R7489 GNDA.n3037 GNDA.n3036 4.5005
R7490 GNDA.n3038 GNDA.n3007 4.5005
R7491 GNDA.n3040 GNDA.n3039 4.5005
R7492 GNDA.n3041 GNDA.n3006 4.5005
R7493 GNDA.n3045 GNDA.n3044 4.5005
R7494 GNDA.n3046 GNDA.n3003 4.5005
R7495 GNDA.n3048 GNDA.n3047 4.5005
R7496 GNDA.n3049 GNDA.n3002 4.5005
R7497 GNDA.n3053 GNDA.n3052 4.5005
R7498 GNDA.n3054 GNDA.n2999 4.5005
R7499 GNDA.n3056 GNDA.n3055 4.5005
R7500 GNDA.n3057 GNDA.n2998 4.5005
R7501 GNDA.n3061 GNDA.n3060 4.5005
R7502 GNDA.n3087 GNDA.n1026 4.5005
R7503 GNDA.n3090 GNDA.n3089 4.5005
R7504 GNDA.n3091 GNDA.n3084 4.5005
R7505 GNDA.n3093 GNDA.n3092 4.5005
R7506 GNDA.n3094 GNDA.n3083 4.5005
R7507 GNDA.n3098 GNDA.n3097 4.5005
R7508 GNDA.n3099 GNDA.n3080 4.5005
R7509 GNDA.n3101 GNDA.n3100 4.5005
R7510 GNDA.n3102 GNDA.n3079 4.5005
R7511 GNDA.n3106 GNDA.n3105 4.5005
R7512 GNDA.n3107 GNDA.n3076 4.5005
R7513 GNDA.n3109 GNDA.n3108 4.5005
R7514 GNDA.n3110 GNDA.n3075 4.5005
R7515 GNDA.n3114 GNDA.n3113 4.5005
R7516 GNDA.n3115 GNDA.n3072 4.5005
R7517 GNDA.n3117 GNDA.n3116 4.5005
R7518 GNDA.n3118 GNDA.n3071 4.5005
R7519 GNDA.n3122 GNDA.n3121 4.5005
R7520 GNDA.n3123 GNDA.n3068 4.5005
R7521 GNDA.n3125 GNDA.n3124 4.5005
R7522 GNDA.n3126 GNDA.n3067 4.5005
R7523 GNDA.n3130 GNDA.n3129 4.5005
R7524 GNDA.n3156 GNDA.n1030 4.5005
R7525 GNDA.n3159 GNDA.n3158 4.5005
R7526 GNDA.n3160 GNDA.n3153 4.5005
R7527 GNDA.n3162 GNDA.n3161 4.5005
R7528 GNDA.n3163 GNDA.n3152 4.5005
R7529 GNDA.n3167 GNDA.n3166 4.5005
R7530 GNDA.n3168 GNDA.n3149 4.5005
R7531 GNDA.n3170 GNDA.n3169 4.5005
R7532 GNDA.n3171 GNDA.n3148 4.5005
R7533 GNDA.n3175 GNDA.n3174 4.5005
R7534 GNDA.n3176 GNDA.n3145 4.5005
R7535 GNDA.n3178 GNDA.n3177 4.5005
R7536 GNDA.n3179 GNDA.n3144 4.5005
R7537 GNDA.n3183 GNDA.n3182 4.5005
R7538 GNDA.n3184 GNDA.n3141 4.5005
R7539 GNDA.n3186 GNDA.n3185 4.5005
R7540 GNDA.n3187 GNDA.n3140 4.5005
R7541 GNDA.n3191 GNDA.n3190 4.5005
R7542 GNDA.n3192 GNDA.n3137 4.5005
R7543 GNDA.n3194 GNDA.n3193 4.5005
R7544 GNDA.n3195 GNDA.n3136 4.5005
R7545 GNDA.n3199 GNDA.n3198 4.5005
R7546 GNDA.n3225 GNDA.n1034 4.5005
R7547 GNDA.n3228 GNDA.n3227 4.5005
R7548 GNDA.n3229 GNDA.n3222 4.5005
R7549 GNDA.n3231 GNDA.n3230 4.5005
R7550 GNDA.n3232 GNDA.n3221 4.5005
R7551 GNDA.n3236 GNDA.n3235 4.5005
R7552 GNDA.n3237 GNDA.n3218 4.5005
R7553 GNDA.n3239 GNDA.n3238 4.5005
R7554 GNDA.n3240 GNDA.n3217 4.5005
R7555 GNDA.n3244 GNDA.n3243 4.5005
R7556 GNDA.n3245 GNDA.n3214 4.5005
R7557 GNDA.n3247 GNDA.n3246 4.5005
R7558 GNDA.n3248 GNDA.n3213 4.5005
R7559 GNDA.n3252 GNDA.n3251 4.5005
R7560 GNDA.n3253 GNDA.n3210 4.5005
R7561 GNDA.n3255 GNDA.n3254 4.5005
R7562 GNDA.n3256 GNDA.n3209 4.5005
R7563 GNDA.n3260 GNDA.n3259 4.5005
R7564 GNDA.n3261 GNDA.n3206 4.5005
R7565 GNDA.n3263 GNDA.n3262 4.5005
R7566 GNDA.n3264 GNDA.n3205 4.5005
R7567 GNDA.n3268 GNDA.n3267 4.5005
R7568 GNDA.n3347 GNDA.n3345 4.5005
R7569 GNDA.n3349 GNDA.n3348 4.5005
R7570 GNDA.n3348 GNDA.n3347 4.5005
R7571 GNDA.n3352 GNDA.n3350 4.5005
R7572 GNDA.n3354 GNDA.n3353 4.5005
R7573 GNDA.n3353 GNDA.n3352 4.5005
R7574 GNDA.n3357 GNDA.n3355 4.5005
R7575 GNDA.n3359 GNDA.n3358 4.5005
R7576 GNDA.n3358 GNDA.n3357 4.5005
R7577 GNDA.n3367 GNDA.n3365 4.5005
R7578 GNDA.n3369 GNDA.n3368 4.5005
R7579 GNDA.n3368 GNDA.n3367 4.5005
R7580 GNDA.n3372 GNDA.n3370 4.5005
R7581 GNDA.n3374 GNDA.n3373 4.5005
R7582 GNDA.n3373 GNDA.n3372 4.5005
R7583 GNDA.n3377 GNDA.n3375 4.5005
R7584 GNDA.n3379 GNDA.n3378 4.5005
R7585 GNDA.n3378 GNDA.n3377 4.5005
R7586 GNDA.n3391 GNDA.n3387 4.5005
R7587 GNDA.n3393 GNDA.n3392 4.5005
R7588 GNDA.n3392 GNDA.n3391 4.5005
R7589 GNDA.n3487 GNDA.n3483 4.5005
R7590 GNDA.n3488 GNDA.n975 4.5005
R7591 GNDA.n3488 GNDA.n3487 4.5005
R7592 GNDA.n3364 GNDA.n3363 4.5005
R7593 GNDA.n3363 GNDA.n3362 4.5005
R7594 GNDA.n3362 GNDA.n3360 4.5005
R7595 GNDA.n1037 GNDA.n1036 4.5005
R7596 GNDA.n3339 GNDA.n3338 4.5005
R7597 GNDA.n1039 GNDA.n1038 4.5005
R7598 GNDA.n3284 GNDA.n3283 4.5005
R7599 GNDA.n3288 GNDA.n3285 4.5005
R7600 GNDA.n3289 GNDA.n3282 4.5005
R7601 GNDA.n3293 GNDA.n3292 4.5005
R7602 GNDA.n3294 GNDA.n3281 4.5005
R7603 GNDA.n3298 GNDA.n3295 4.5005
R7604 GNDA.n3299 GNDA.n3280 4.5005
R7605 GNDA.n3303 GNDA.n3302 4.5005
R7606 GNDA.n3304 GNDA.n3279 4.5005
R7607 GNDA.n3308 GNDA.n3305 4.5005
R7608 GNDA.n3309 GNDA.n3278 4.5005
R7609 GNDA.n3313 GNDA.n3312 4.5005
R7610 GNDA.n3314 GNDA.n3277 4.5005
R7611 GNDA.n3318 GNDA.n3315 4.5005
R7612 GNDA.n3319 GNDA.n3276 4.5005
R7613 GNDA.n3323 GNDA.n3322 4.5005
R7614 GNDA.n3324 GNDA.n3275 4.5005
R7615 GNDA.n3328 GNDA.n3325 4.5005
R7616 GNDA.n3329 GNDA.n3274 4.5005
R7617 GNDA.n3333 GNDA.n3332 4.5005
R7618 GNDA.n593 GNDA.n592 4.5005
R7619 GNDA.n591 GNDA.n514 4.5005
R7620 GNDA.n590 GNDA.n589 4.5005
R7621 GNDA.n588 GNDA.n518 4.5005
R7622 GNDA.n587 GNDA.n586 4.5005
R7623 GNDA.n585 GNDA.n519 4.5005
R7624 GNDA.n584 GNDA.n583 4.5005
R7625 GNDA.n582 GNDA.n526 4.5005
R7626 GNDA.n581 GNDA.n580 4.5005
R7627 GNDA.n579 GNDA.n527 4.5005
R7628 GNDA.n578 GNDA.n577 4.5005
R7629 GNDA.n576 GNDA.n534 4.5005
R7630 GNDA.n575 GNDA.n574 4.5005
R7631 GNDA.n573 GNDA.n535 4.5005
R7632 GNDA.n572 GNDA.n571 4.5005
R7633 GNDA.n570 GNDA.n542 4.5005
R7634 GNDA.n569 GNDA.n568 4.5005
R7635 GNDA.n567 GNDA.n543 4.5005
R7636 GNDA.n566 GNDA.n565 4.5005
R7637 GNDA.n564 GNDA.n550 4.5005
R7638 GNDA.n563 GNDA.n562 4.5005
R7639 GNDA.n561 GNDA.n551 4.5005
R7640 GNDA.n596 GNDA.n594 4.5005
R7641 GNDA.n598 GNDA.n597 4.5005
R7642 GNDA.n597 GNDA.n596 4.5005
R7643 GNDA.n4369 GNDA.n4368 4.5005
R7644 GNDA.n4368 GNDA.n4367 4.5005
R7645 GNDA.n4367 GNDA.n4283 4.5005
R7646 GNDA.n4370 GNDA.n441 4.5005
R7647 GNDA.n4371 GNDA.n4370 4.5005
R7648 GNDA.n4372 GNDA.n4371 4.5005
R7649 GNDA.n4880 GNDA.n4879 4.5005
R7650 GNDA.n4879 GNDA.n4878 4.5005
R7651 GNDA.n4878 GNDA.n442 4.5005
R7652 GNDA.n4279 GNDA.n4278 4.5005
R7653 GNDA.n4278 GNDA.n4277 4.5005
R7654 GNDA.n4277 GNDA.n482 4.5005
R7655 GNDA.n4745 GNDA.n4742 4.5005
R7656 GNDA.n4746 GNDA.n4745 4.5005
R7657 GNDA.n4747 GNDA.n4746 4.5005
R7658 GNDA.n4738 GNDA.n4471 4.5005
R7659 GNDA.n4741 GNDA.n4471 4.5005
R7660 GNDA.n4741 GNDA.n4470 4.5005
R7661 GNDA.n4734 GNDA.n4557 4.5005
R7662 GNDA.n4737 GNDA.n4557 4.5005
R7663 GNDA.n4737 GNDA.n4556 4.5005
R7664 GNDA.n4730 GNDA.n4562 4.5005
R7665 GNDA.n4733 GNDA.n4562 4.5005
R7666 GNDA.n4733 GNDA.n4561 4.5005
R7667 GNDA.n4886 GNDA.n437 4.5005
R7668 GNDA.n4886 GNDA.n4885 4.5005
R7669 GNDA.n4885 GNDA.n4881 4.5005
R7670 GNDA.n1924 GNDA.n1923 4.5005
R7671 GNDA.n2048 GNDA.n2047 4.5005
R7672 GNDA.n1892 GNDA.n1891 4.5005
R7673 GNDA.n2053 GNDA.n1885 4.5005
R7674 GNDA.n2052 GNDA.n1555 4.5005
R7675 GNDA.n2053 GNDA.n2052 4.5005
R7676 GNDA.n1487 GNDA.n1486 4.5005
R7677 GNDA.n1497 GNDA.n1496 4.5005
R7678 GNDA.n1498 GNDA.n1485 4.5005
R7679 GNDA.n1500 GNDA.n1499 4.5005
R7680 GNDA.n1483 GNDA.n1482 4.5005
R7681 GNDA.n1507 GNDA.n1506 4.5005
R7682 GNDA.n1508 GNDA.n1481 4.5005
R7683 GNDA.n1510 GNDA.n1509 4.5005
R7684 GNDA.n1479 GNDA.n1478 4.5005
R7685 GNDA.n1517 GNDA.n1516 4.5005
R7686 GNDA.n1518 GNDA.n1477 4.5005
R7687 GNDA.n1520 GNDA.n1519 4.5005
R7688 GNDA.n1475 GNDA.n1474 4.5005
R7689 GNDA.n1527 GNDA.n1526 4.5005
R7690 GNDA.n1528 GNDA.n1473 4.5005
R7691 GNDA.n1530 GNDA.n1529 4.5005
R7692 GNDA.n1471 GNDA.n1470 4.5005
R7693 GNDA.n1537 GNDA.n1536 4.5005
R7694 GNDA.n1538 GNDA.n1469 4.5005
R7695 GNDA.n1540 GNDA.n1539 4.5005
R7696 GNDA.n1467 GNDA.n1466 4.5005
R7697 GNDA.n1546 GNDA.n1545 4.5005
R7698 GNDA.n1554 GNDA.n1553 4.5005
R7699 GNDA.n1550 GNDA.n1464 4.5005
R7700 GNDA.n1551 GNDA.n1459 4.5005
R7701 GNDA.n1551 GNDA.n1550 4.5005
R7702 GNDA.n1461 GNDA.n359 4.5005
R7703 GNDA.n1418 GNDA.n1417 4.5005
R7704 GNDA.n1421 GNDA.n1420 4.5005
R7705 GNDA.n1365 GNDA.n1361 4.5005
R7706 GNDA.n1369 GNDA.n1366 4.5005
R7707 GNDA.n1370 GNDA.n1360 4.5005
R7708 GNDA.n1374 GNDA.n1373 4.5005
R7709 GNDA.n1375 GNDA.n1359 4.5005
R7710 GNDA.n1379 GNDA.n1376 4.5005
R7711 GNDA.n1380 GNDA.n1358 4.5005
R7712 GNDA.n1384 GNDA.n1383 4.5005
R7713 GNDA.n1385 GNDA.n1357 4.5005
R7714 GNDA.n1389 GNDA.n1386 4.5005
R7715 GNDA.n1390 GNDA.n1356 4.5005
R7716 GNDA.n1394 GNDA.n1393 4.5005
R7717 GNDA.n1395 GNDA.n1355 4.5005
R7718 GNDA.n1399 GNDA.n1396 4.5005
R7719 GNDA.n1400 GNDA.n1354 4.5005
R7720 GNDA.n1404 GNDA.n1403 4.5005
R7721 GNDA.n1405 GNDA.n1353 4.5005
R7722 GNDA.n1409 GNDA.n1406 4.5005
R7723 GNDA.n1410 GNDA.n1352 4.5005
R7724 GNDA.n1414 GNDA.n1413 4.5005
R7725 GNDA.n1415 GNDA.n1351 4.5005
R7726 GNDA.n2577 GNDA.n2576 4.5005
R7727 GNDA.n4061 GNDA.t123 4.47811
R7728 GNDA.t59 GNDA.n4060 4.47811
R7729 GNDA.n4044 GNDA.t97 4.47811
R7730 GNDA.t133 GNDA.n634 4.47811
R7731 GNDA.n346 GNDA.n302 4.26717
R7732 GNDA.n346 GNDA.n345 4.26717
R7733 GNDA.n345 GNDA.n344 4.26717
R7734 GNDA.n344 GNDA.n310 4.26717
R7735 GNDA.n338 GNDA.n310 4.26717
R7736 GNDA.n338 GNDA.n337 4.26717
R7737 GNDA.n337 GNDA.n336 4.26717
R7738 GNDA.n336 GNDA.n318 4.26717
R7739 GNDA.n330 GNDA.n318 4.26717
R7740 GNDA.n330 GNDA.n329 4.26717
R7741 GNDA.n329 GNDA.n328 4.26717
R7742 GNDA.n5365 GNDA.n134 4.26717
R7743 GNDA.n5359 GNDA.n134 4.26717
R7744 GNDA.n5359 GNDA.n5358 4.26717
R7745 GNDA.n5358 GNDA.n5357 4.26717
R7746 GNDA.n5357 GNDA.n5355 4.26717
R7747 GNDA.n5355 GNDA.n5352 4.26717
R7748 GNDA.n5352 GNDA.n5351 4.26717
R7749 GNDA.n5351 GNDA.n5348 4.26717
R7750 GNDA.n5348 GNDA.n5347 4.26717
R7751 GNDA.n5347 GNDA.n5344 4.26717
R7752 GNDA.n5344 GNDA.n5343 4.26717
R7753 GNDA.n2109 GNDA.n2108 4.26717
R7754 GNDA.n2108 GNDA.n1693 4.26717
R7755 GNDA.n2104 GNDA.n1693 4.26717
R7756 GNDA.n2104 GNDA.n2103 4.26717
R7757 GNDA.n2103 GNDA.n1699 4.26717
R7758 GNDA.n2098 GNDA.n1699 4.26717
R7759 GNDA.n2098 GNDA.n2097 4.26717
R7760 GNDA.n2097 GNDA.n2096 4.26717
R7761 GNDA.n2096 GNDA.n1707 4.26717
R7762 GNDA.n2090 GNDA.n1707 4.26717
R7763 GNDA.n2090 GNDA.n2089 4.26717
R7764 GNDA.n411 GNDA.n410 4.26717
R7765 GNDA.n410 GNDA.n371 4.26717
R7766 GNDA.n405 GNDA.n371 4.26717
R7767 GNDA.n405 GNDA.n404 4.26717
R7768 GNDA.n404 GNDA.n403 4.26717
R7769 GNDA.n403 GNDA.n379 4.26717
R7770 GNDA.n397 GNDA.n379 4.26717
R7771 GNDA.n397 GNDA.n396 4.26717
R7772 GNDA.n396 GNDA.n395 4.26717
R7773 GNDA.n395 GNDA.n390 4.26717
R7774 GNDA.n390 GNDA.n389 4.26717
R7775 GNDA.n2354 GNDA.n2151 4.26717
R7776 GNDA.n2354 GNDA.n2149 4.26717
R7777 GNDA.n2360 GNDA.n2149 4.26717
R7778 GNDA.n2360 GNDA.n2147 4.26717
R7779 GNDA.n2366 GNDA.n2147 4.26717
R7780 GNDA.n2366 GNDA.n2145 4.26717
R7781 GNDA.n2372 GNDA.n2145 4.26717
R7782 GNDA.n2372 GNDA.n2143 4.26717
R7783 GNDA.n2378 GNDA.n2143 4.26717
R7784 GNDA.n2378 GNDA.n2141 4.26717
R7785 GNDA.n2383 GNDA.n2141 4.26717
R7786 GNDA.n2445 GNDA.n1681 4.26717
R7787 GNDA.n2448 GNDA.n2445 4.26717
R7788 GNDA.n2451 GNDA.n2448 4.26717
R7789 GNDA.n2451 GNDA.n1679 4.26717
R7790 GNDA.n2457 GNDA.n1679 4.26717
R7791 GNDA.n2460 GNDA.n2457 4.26717
R7792 GNDA.n2462 GNDA.n2460 4.26717
R7793 GNDA.n2462 GNDA.n1677 4.26717
R7794 GNDA.n2468 GNDA.n1677 4.26717
R7795 GNDA.n2468 GNDA.n1602 4.26717
R7796 GNDA.n2477 GNDA.n1602 4.26717
R7797 GNDA.t290 GNDA.t152 4.14363
R7798 GNDA.n4985 GNDA.n302 3.93531
R7799 GNDA.n5366 GNDA.n5365 3.93531
R7800 GNDA.n2109 GNDA.n1688 3.93531
R7801 GNDA.n411 GNDA.n365 3.93531
R7802 GNDA.n2175 GNDA.n2151 3.93531
R7803 GNDA.n2387 GNDA.n1681 3.93531
R7804 GNDA.n4282 GNDA.n4281 3.84081
R7805 GNDA.n3482 GNDA.n3481 3.84081
R7806 GNDA.n3386 GNDA.n3385 3.84081
R7807 GNDA.n4133 GNDA.n4132 3.84045
R7808 GNDA.n2499 GNDA.n1597 3.7893
R7809 GNDA.n2498 GNDA.n1598 3.7893
R7810 GNDA.n2486 GNDA.n2485 3.7893
R7811 GNDA.n2492 GNDA.n2491 3.7893
R7812 GNDA.n2488 GNDA.n2487 3.7893
R7813 GNDA.n1573 GNDA.n1566 3.7893
R7814 GNDA.n1579 GNDA.n1577 3.7893
R7815 GNDA.n1578 GNDA.n1448 3.7893
R7816 GNDA.n1996 GNDA.n1933 3.7893
R7817 GNDA.n2005 GNDA.n2004 3.7893
R7818 GNDA.n1934 GNDA.n1909 3.7893
R7819 GNDA.n2014 GNDA.n2012 3.7893
R7820 GNDA.n2013 GNDA.n1907 3.7893
R7821 GNDA.n1906 GNDA.n1903 3.7893
R7822 GNDA.n2030 GNDA.n2028 3.7893
R7823 GNDA.n2029 GNDA.n1899 3.7893
R7824 GNDA.n5337 GNDA.n165 3.7893
R7825 GNDA.n5334 GNDA.n5333 3.7893
R7826 GNDA.n200 GNDA.n167 3.7893
R7827 GNDA.n218 GNDA.n217 3.7893
R7828 GNDA.n215 GNDA.n214 3.7893
R7829 GNDA.n210 GNDA.n203 3.7893
R7830 GNDA.n207 GNDA.n206 3.7893
R7831 GNDA.n5275 GNDA.n187 3.7893
R7832 GNDA.n2290 GNDA.n2265 3.7893
R7833 GNDA.n2289 GNDA.n2286 3.7893
R7834 GNDA.n2285 GNDA.n2266 3.7893
R7835 GNDA.n2282 GNDA.n2281 3.7893
R7836 GNDA.n2278 GNDA.n2267 3.7893
R7837 GNDA.n2271 GNDA.n2268 3.7893
R7838 GNDA.n2295 GNDA.n2190 3.7893
R7839 GNDA.n2296 GNDA.n2189 3.7893
R7840 GNDA.n5266 GNDA.n5265 3.7893
R7841 GNDA.n5262 GNDA.n5156 3.7893
R7842 GNDA.n5261 GNDA.n5159 3.7893
R7843 GNDA.n5258 GNDA.n5257 3.7893
R7844 GNDA.n5184 GNDA.n5160 3.7893
R7845 GNDA.n5193 GNDA.n5192 3.7893
R7846 GNDA.n5196 GNDA.n5183 3.7893
R7847 GNDA.n5201 GNDA.n5197 3.7893
R7848 GNDA.n5545 GNDA.n5544 3.7893
R7849 GNDA.n5541 GNDA.n59 3.7893
R7850 GNDA.n5540 GNDA.n62 3.7893
R7851 GNDA.n5537 GNDA.n5536 3.7893
R7852 GNDA.n5463 GNDA.n63 3.7893
R7853 GNDA.n5472 GNDA.n5471 3.7893
R7854 GNDA.n5475 GNDA.n5462 3.7893
R7855 GNDA.n5480 GNDA.n5476 3.7893
R7856 GNDA.n5122 GNDA.n5011 3.7893
R7857 GNDA.n5119 GNDA.n5118 3.7893
R7858 GNDA.n5035 GNDA.n5012 3.7893
R7859 GNDA.n5040 GNDA.n5038 3.7893
R7860 GNDA.n5045 GNDA.n5041 3.7893
R7861 GNDA.n5052 GNDA.n5051 3.7893
R7862 GNDA.n5055 GNDA.n5034 3.7893
R7863 GNDA.n5060 GNDA.n5056 3.7893
R7864 GNDA.n1859 GNDA.n1858 3.7893
R7865 GNDA.n1871 GNDA.n1730 3.7893
R7866 GNDA.n1870 GNDA.n1728 3.7893
R7867 GNDA.n1877 GNDA.n1727 3.7893
R7868 GNDA.n1879 GNDA.n1878 3.7893
R7869 GNDA.n2071 GNDA.n1724 3.7893
R7870 GNDA.n1723 GNDA.n1720 3.7893
R7871 GNDA.n2080 GNDA.n2079 3.7893
R7872 GNDA.n5554 GNDA.n22 3.7893
R7873 GNDA.n5553 GNDA.n23 3.7893
R7874 GNDA.n33 GNDA.n32 3.7893
R7875 GNDA.n39 GNDA.n38 3.7893
R7876 GNDA.n35 GNDA.n34 3.7893
R7877 GNDA.n5388 GNDA.n1 3.7893
R7878 GNDA.n5393 GNDA.n5391 3.7893
R7879 GNDA.n5398 GNDA.n5394 3.7893
R7880 GNDA GNDA.n2504 3.7381
R7881 GNDA GNDA.n2020 3.7381
R7882 GNDA.n211 GNDA 3.7381
R7883 GNDA GNDA.n2274 3.7381
R7884 GNDA.n5189 GNDA 3.7381
R7885 GNDA.n5468 GNDA 3.7381
R7886 GNDA.n5048 GNDA 3.7381
R7887 GNDA.n2072 GNDA 3.7381
R7888 GNDA GNDA.n5559 3.7381
R7889 GNDA.n559 GNDA.n558 3.50398
R7890 GNDA.n1364 GNDA.n1337 3.47871
R7891 GNDA.n4722 GNDA.n4721 3.47821
R7892 GNDA.n4646 GNDA.n4645 3.47821
R7893 GNDA.n4516 GNDA.n4515 3.47821
R7894 GNDA.n4806 GNDA.n4805 3.47821
R7895 GNDA.n4270 GNDA.n4269 3.47821
R7896 GNDA.n4871 GNDA.n4870 3.47821
R7897 GNDA.n4431 GNDA.n4430 3.47821
R7898 GNDA.n4328 GNDA.n4327 3.47821
R7899 GNDA.n4194 GNDA.n4193 3.47821
R7900 GNDA.n3953 GNDA.n3952 3.47821
R7901 GNDA.n3617 GNDA.n3616 3.47821
R7902 GNDA.n3933 GNDA.n3932 3.47821
R7903 GNDA.n887 GNDA.n886 3.47821
R7904 GNDA.n3721 GNDA.n3720 3.47821
R7905 GNDA.n3790 GNDA.n3789 3.47821
R7906 GNDA.n3855 GNDA.n3854 3.47821
R7907 GNDA.n3441 GNDA.n3440 3.47821
R7908 GNDA.n3535 GNDA.n3534 3.47821
R7909 GNDA.n2856 GNDA.n2855 3.47821
R7910 GNDA.n2925 GNDA.n2924 3.47821
R7911 GNDA.n2994 GNDA.n2993 3.47821
R7912 GNDA.n3063 GNDA.n3062 3.47821
R7913 GNDA.n3132 GNDA.n3131 3.47821
R7914 GNDA.n3201 GNDA.n3200 3.47821
R7915 GNDA.n3270 GNDA.n3269 3.47821
R7916 GNDA.n3335 GNDA.n3334 3.47821
R7917 GNDA.n1489 GNDA.n1488 3.47821
R7918 GNDA.n592 GNDA.n515 3.43627
R7919 GNDA.n479 GNDA.t8 3.42907
R7920 GNDA.n479 GNDA.t137 3.42907
R7921 GNDA.n4135 GNDA.t81 3.42907
R7922 GNDA.n4135 GNDA.t145 3.42907
R7923 GNDA.n3476 GNDA.t128 3.42907
R7924 GNDA.n3476 GNDA.t23 3.42907
R7925 GNDA.n3388 GNDA.t139 3.42907
R7926 GNDA.n3388 GNDA.t34 3.42907
R7927 GNDA.n4660 GNDA.n4659 3.4105
R7928 GNDA.n4719 GNDA.n4718 3.4105
R7929 GNDA.n4717 GNDA.n4716 3.4105
R7930 GNDA.n4715 GNDA.n4714 3.4105
R7931 GNDA.n4713 GNDA.n4662 3.4105
R7932 GNDA.n4709 GNDA.n4708 3.4105
R7933 GNDA.n4707 GNDA.n4706 3.4105
R7934 GNDA.n4705 GNDA.n4704 3.4105
R7935 GNDA.n4703 GNDA.n4664 3.4105
R7936 GNDA.n4699 GNDA.n4698 3.4105
R7937 GNDA.n4697 GNDA.n4696 3.4105
R7938 GNDA.n4695 GNDA.n4694 3.4105
R7939 GNDA.n4693 GNDA.n4666 3.4105
R7940 GNDA.n4689 GNDA.n4688 3.4105
R7941 GNDA.n4687 GNDA.n4686 3.4105
R7942 GNDA.n4685 GNDA.n4684 3.4105
R7943 GNDA.n4683 GNDA.n4668 3.4105
R7944 GNDA.n4679 GNDA.n4678 3.4105
R7945 GNDA.n4677 GNDA.n4676 3.4105
R7946 GNDA.n4675 GNDA.n4674 3.4105
R7947 GNDA.n4673 GNDA.n4670 3.4105
R7948 GNDA.n4565 GNDA.n4564 3.4105
R7949 GNDA.n4725 GNDA.n4724 3.4105
R7950 GNDA.n4579 GNDA.n4578 3.4105
R7951 GNDA.n4643 GNDA.n4642 3.4105
R7952 GNDA.n4641 GNDA.n4640 3.4105
R7953 GNDA.n4639 GNDA.n4638 3.4105
R7954 GNDA.n4637 GNDA.n4581 3.4105
R7955 GNDA.n4633 GNDA.n4632 3.4105
R7956 GNDA.n4631 GNDA.n4630 3.4105
R7957 GNDA.n4629 GNDA.n4628 3.4105
R7958 GNDA.n4627 GNDA.n4583 3.4105
R7959 GNDA.n4623 GNDA.n4622 3.4105
R7960 GNDA.n4621 GNDA.n4620 3.4105
R7961 GNDA.n4619 GNDA.n4618 3.4105
R7962 GNDA.n4617 GNDA.n4585 3.4105
R7963 GNDA.n4613 GNDA.n4612 3.4105
R7964 GNDA.n4611 GNDA.n4610 3.4105
R7965 GNDA.n4609 GNDA.n4608 3.4105
R7966 GNDA.n4607 GNDA.n4587 3.4105
R7967 GNDA.n4603 GNDA.n4602 3.4105
R7968 GNDA.n4601 GNDA.n4600 3.4105
R7969 GNDA.n4599 GNDA.n4598 3.4105
R7970 GNDA.n4597 GNDA.n4589 3.4105
R7971 GNDA.n4593 GNDA.n4592 3.4105
R7972 GNDA.n4591 GNDA.n4566 3.4105
R7973 GNDA.n4517 GNDA.n4494 3.4105
R7974 GNDA.n4519 GNDA.n4493 3.4105
R7975 GNDA.n4520 GNDA.n4492 3.4105
R7976 GNDA.n4522 GNDA.n4491 3.4105
R7977 GNDA.n4523 GNDA.n4490 3.4105
R7978 GNDA.n4525 GNDA.n4489 3.4105
R7979 GNDA.n4526 GNDA.n4488 3.4105
R7980 GNDA.n4528 GNDA.n4487 3.4105
R7981 GNDA.n4529 GNDA.n4486 3.4105
R7982 GNDA.n4531 GNDA.n4485 3.4105
R7983 GNDA.n4532 GNDA.n4484 3.4105
R7984 GNDA.n4534 GNDA.n4483 3.4105
R7985 GNDA.n4535 GNDA.n4482 3.4105
R7986 GNDA.n4537 GNDA.n4481 3.4105
R7987 GNDA.n4538 GNDA.n4480 3.4105
R7988 GNDA.n4540 GNDA.n4479 3.4105
R7989 GNDA.n4541 GNDA.n4478 3.4105
R7990 GNDA.n4543 GNDA.n4477 3.4105
R7991 GNDA.n4544 GNDA.n4476 3.4105
R7992 GNDA.n4546 GNDA.n4475 3.4105
R7993 GNDA.n4547 GNDA.n4474 3.4105
R7994 GNDA.n4549 GNDA.n4473 3.4105
R7995 GNDA.n4551 GNDA.n4550 3.4105
R7996 GNDA.n4458 GNDA.n4457 3.4105
R7997 GNDA.n4803 GNDA.n4802 3.4105
R7998 GNDA.n4801 GNDA.n4800 3.4105
R7999 GNDA.n4799 GNDA.n4798 3.4105
R8000 GNDA.n4797 GNDA.n4460 3.4105
R8001 GNDA.n4793 GNDA.n4792 3.4105
R8002 GNDA.n4791 GNDA.n4790 3.4105
R8003 GNDA.n4789 GNDA.n4788 3.4105
R8004 GNDA.n4787 GNDA.n4462 3.4105
R8005 GNDA.n4783 GNDA.n4782 3.4105
R8006 GNDA.n4781 GNDA.n4780 3.4105
R8007 GNDA.n4779 GNDA.n4778 3.4105
R8008 GNDA.n4777 GNDA.n4464 3.4105
R8009 GNDA.n4773 GNDA.n4772 3.4105
R8010 GNDA.n4771 GNDA.n4770 3.4105
R8011 GNDA.n4769 GNDA.n4768 3.4105
R8012 GNDA.n4767 GNDA.n4466 3.4105
R8013 GNDA.n4763 GNDA.n4762 3.4105
R8014 GNDA.n4761 GNDA.n4760 3.4105
R8015 GNDA.n4759 GNDA.n4758 3.4105
R8016 GNDA.n4757 GNDA.n4468 3.4105
R8017 GNDA.n4753 GNDA.n4752 3.4105
R8018 GNDA.n4751 GNDA.n4444 3.4105
R8019 GNDA.n4208 GNDA.n4207 3.4105
R8020 GNDA.n4267 GNDA.n4266 3.4105
R8021 GNDA.n4265 GNDA.n4264 3.4105
R8022 GNDA.n4263 GNDA.n4262 3.4105
R8023 GNDA.n4261 GNDA.n4210 3.4105
R8024 GNDA.n4257 GNDA.n4256 3.4105
R8025 GNDA.n4255 GNDA.n4254 3.4105
R8026 GNDA.n4253 GNDA.n4252 3.4105
R8027 GNDA.n4251 GNDA.n4212 3.4105
R8028 GNDA.n4247 GNDA.n4246 3.4105
R8029 GNDA.n4245 GNDA.n4244 3.4105
R8030 GNDA.n4243 GNDA.n4242 3.4105
R8031 GNDA.n4241 GNDA.n4214 3.4105
R8032 GNDA.n4237 GNDA.n4236 3.4105
R8033 GNDA.n4235 GNDA.n4234 3.4105
R8034 GNDA.n4233 GNDA.n4232 3.4105
R8035 GNDA.n4231 GNDA.n4216 3.4105
R8036 GNDA.n4227 GNDA.n4226 3.4105
R8037 GNDA.n4225 GNDA.n4224 3.4105
R8038 GNDA.n4223 GNDA.n4222 3.4105
R8039 GNDA.n4221 GNDA.n4218 3.4105
R8040 GNDA.n485 GNDA.n484 3.4105
R8041 GNDA.n4273 GNDA.n4272 3.4105
R8042 GNDA.n4809 GNDA.n4808 3.4105
R8043 GNDA.n4868 GNDA.n4867 3.4105
R8044 GNDA.n4866 GNDA.n4865 3.4105
R8045 GNDA.n4864 GNDA.n4863 3.4105
R8046 GNDA.n4862 GNDA.n4811 3.4105
R8047 GNDA.n4858 GNDA.n4857 3.4105
R8048 GNDA.n4856 GNDA.n4855 3.4105
R8049 GNDA.n4854 GNDA.n4853 3.4105
R8050 GNDA.n4852 GNDA.n4813 3.4105
R8051 GNDA.n4848 GNDA.n4847 3.4105
R8052 GNDA.n4846 GNDA.n4845 3.4105
R8053 GNDA.n4844 GNDA.n4843 3.4105
R8054 GNDA.n4842 GNDA.n4815 3.4105
R8055 GNDA.n4838 GNDA.n4837 3.4105
R8056 GNDA.n4836 GNDA.n4835 3.4105
R8057 GNDA.n4834 GNDA.n4833 3.4105
R8058 GNDA.n4832 GNDA.n4817 3.4105
R8059 GNDA.n4828 GNDA.n4827 3.4105
R8060 GNDA.n4826 GNDA.n4825 3.4105
R8061 GNDA.n4824 GNDA.n4823 3.4105
R8062 GNDA.n4822 GNDA.n4819 3.4105
R8063 GNDA.n445 GNDA.n444 3.4105
R8064 GNDA.n4874 GNDA.n4873 3.4105
R8065 GNDA.n460 GNDA.n459 3.4105
R8066 GNDA.n4428 GNDA.n4427 3.4105
R8067 GNDA.n4426 GNDA.n4425 3.4105
R8068 GNDA.n4424 GNDA.n4423 3.4105
R8069 GNDA.n4422 GNDA.n462 3.4105
R8070 GNDA.n4418 GNDA.n4417 3.4105
R8071 GNDA.n4416 GNDA.n4415 3.4105
R8072 GNDA.n4414 GNDA.n4413 3.4105
R8073 GNDA.n4412 GNDA.n464 3.4105
R8074 GNDA.n4408 GNDA.n4407 3.4105
R8075 GNDA.n4406 GNDA.n4405 3.4105
R8076 GNDA.n4404 GNDA.n4403 3.4105
R8077 GNDA.n4402 GNDA.n466 3.4105
R8078 GNDA.n4398 GNDA.n4397 3.4105
R8079 GNDA.n4396 GNDA.n4395 3.4105
R8080 GNDA.n4394 GNDA.n4393 3.4105
R8081 GNDA.n4392 GNDA.n468 3.4105
R8082 GNDA.n4388 GNDA.n4387 3.4105
R8083 GNDA.n4386 GNDA.n4385 3.4105
R8084 GNDA.n4384 GNDA.n4383 3.4105
R8085 GNDA.n4382 GNDA.n470 3.4105
R8086 GNDA.n4378 GNDA.n4377 3.4105
R8087 GNDA.n4376 GNDA.n447 3.4105
R8088 GNDA.n4329 GNDA.n4306 3.4105
R8089 GNDA.n4331 GNDA.n4305 3.4105
R8090 GNDA.n4332 GNDA.n4304 3.4105
R8091 GNDA.n4334 GNDA.n4303 3.4105
R8092 GNDA.n4335 GNDA.n4302 3.4105
R8093 GNDA.n4337 GNDA.n4301 3.4105
R8094 GNDA.n4338 GNDA.n4300 3.4105
R8095 GNDA.n4340 GNDA.n4299 3.4105
R8096 GNDA.n4341 GNDA.n4298 3.4105
R8097 GNDA.n4343 GNDA.n4297 3.4105
R8098 GNDA.n4344 GNDA.n4296 3.4105
R8099 GNDA.n4346 GNDA.n4295 3.4105
R8100 GNDA.n4347 GNDA.n4294 3.4105
R8101 GNDA.n4349 GNDA.n4293 3.4105
R8102 GNDA.n4350 GNDA.n4292 3.4105
R8103 GNDA.n4352 GNDA.n4291 3.4105
R8104 GNDA.n4353 GNDA.n4290 3.4105
R8105 GNDA.n4355 GNDA.n4289 3.4105
R8106 GNDA.n4356 GNDA.n4288 3.4105
R8107 GNDA.n4358 GNDA.n4287 3.4105
R8108 GNDA.n4359 GNDA.n4286 3.4105
R8109 GNDA.n4361 GNDA.n4285 3.4105
R8110 GNDA.n4363 GNDA.n4362 3.4105
R8111 GNDA.n500 GNDA.n499 3.4105
R8112 GNDA.n4191 GNDA.n4190 3.4105
R8113 GNDA.n4189 GNDA.n4188 3.4105
R8114 GNDA.n4187 GNDA.n4186 3.4105
R8115 GNDA.n4185 GNDA.n502 3.4105
R8116 GNDA.n4181 GNDA.n4180 3.4105
R8117 GNDA.n4179 GNDA.n4178 3.4105
R8118 GNDA.n4177 GNDA.n4176 3.4105
R8119 GNDA.n4175 GNDA.n504 3.4105
R8120 GNDA.n4171 GNDA.n4170 3.4105
R8121 GNDA.n4169 GNDA.n4168 3.4105
R8122 GNDA.n4167 GNDA.n4166 3.4105
R8123 GNDA.n4165 GNDA.n506 3.4105
R8124 GNDA.n4161 GNDA.n4160 3.4105
R8125 GNDA.n4159 GNDA.n4158 3.4105
R8126 GNDA.n4157 GNDA.n4156 3.4105
R8127 GNDA.n4155 GNDA.n508 3.4105
R8128 GNDA.n4151 GNDA.n4150 3.4105
R8129 GNDA.n4149 GNDA.n4148 3.4105
R8130 GNDA.n4147 GNDA.n4146 3.4105
R8131 GNDA.n4145 GNDA.n510 3.4105
R8132 GNDA.n4141 GNDA.n4140 3.4105
R8133 GNDA.n4139 GNDA.n487 3.4105
R8134 GNDA.n3954 GNDA.n801 3.4105
R8135 GNDA.n3955 GNDA.n800 3.4105
R8136 GNDA.n3956 GNDA.n799 3.4105
R8137 GNDA.n3948 GNDA.n797 3.4105
R8138 GNDA.n3960 GNDA.n796 3.4105
R8139 GNDA.n3961 GNDA.n795 3.4105
R8140 GNDA.n3962 GNDA.n794 3.4105
R8141 GNDA.n3945 GNDA.n792 3.4105
R8142 GNDA.n3966 GNDA.n791 3.4105
R8143 GNDA.n3967 GNDA.n790 3.4105
R8144 GNDA.n3968 GNDA.n789 3.4105
R8145 GNDA.n3942 GNDA.n787 3.4105
R8146 GNDA.n3972 GNDA.n786 3.4105
R8147 GNDA.n3973 GNDA.n785 3.4105
R8148 GNDA.n3974 GNDA.n784 3.4105
R8149 GNDA.n3939 GNDA.n782 3.4105
R8150 GNDA.n3978 GNDA.n781 3.4105
R8151 GNDA.n3979 GNDA.n780 3.4105
R8152 GNDA.n3980 GNDA.n779 3.4105
R8153 GNDA.n3936 GNDA.n777 3.4105
R8154 GNDA.n3984 GNDA.n776 3.4105
R8155 GNDA.n3985 GNDA.n775 3.4105
R8156 GNDA.n3986 GNDA.n774 3.4105
R8157 GNDA.n3550 GNDA.n3549 3.4105
R8158 GNDA.n3614 GNDA.n3613 3.4105
R8159 GNDA.n3612 GNDA.n3611 3.4105
R8160 GNDA.n3610 GNDA.n3554 3.4105
R8161 GNDA.n3553 GNDA.n3552 3.4105
R8162 GNDA.n3606 GNDA.n3605 3.4105
R8163 GNDA.n3604 GNDA.n3603 3.4105
R8164 GNDA.n3602 GNDA.n3558 3.4105
R8165 GNDA.n3557 GNDA.n3556 3.4105
R8166 GNDA.n3598 GNDA.n3597 3.4105
R8167 GNDA.n3596 GNDA.n3595 3.4105
R8168 GNDA.n3594 GNDA.n3562 3.4105
R8169 GNDA.n3561 GNDA.n3560 3.4105
R8170 GNDA.n3590 GNDA.n3589 3.4105
R8171 GNDA.n3588 GNDA.n3587 3.4105
R8172 GNDA.n3586 GNDA.n3566 3.4105
R8173 GNDA.n3565 GNDA.n3564 3.4105
R8174 GNDA.n3582 GNDA.n3581 3.4105
R8175 GNDA.n3580 GNDA.n3579 3.4105
R8176 GNDA.n3578 GNDA.n3570 3.4105
R8177 GNDA.n3569 GNDA.n3568 3.4105
R8178 GNDA.n3574 GNDA.n3573 3.4105
R8179 GNDA.n3572 GNDA.n3537 3.4105
R8180 GNDA.n816 GNDA.n815 3.4105
R8181 GNDA.n3930 GNDA.n3929 3.4105
R8182 GNDA.n3928 GNDA.n3927 3.4105
R8183 GNDA.n3926 GNDA.n820 3.4105
R8184 GNDA.n819 GNDA.n818 3.4105
R8185 GNDA.n3922 GNDA.n3921 3.4105
R8186 GNDA.n3920 GNDA.n3919 3.4105
R8187 GNDA.n3918 GNDA.n824 3.4105
R8188 GNDA.n823 GNDA.n822 3.4105
R8189 GNDA.n3914 GNDA.n3913 3.4105
R8190 GNDA.n3912 GNDA.n3911 3.4105
R8191 GNDA.n3910 GNDA.n828 3.4105
R8192 GNDA.n827 GNDA.n826 3.4105
R8193 GNDA.n3906 GNDA.n3905 3.4105
R8194 GNDA.n3904 GNDA.n3903 3.4105
R8195 GNDA.n3902 GNDA.n832 3.4105
R8196 GNDA.n831 GNDA.n830 3.4105
R8197 GNDA.n3898 GNDA.n3897 3.4105
R8198 GNDA.n3896 GNDA.n3895 3.4105
R8199 GNDA.n3894 GNDA.n836 3.4105
R8200 GNDA.n835 GNDA.n834 3.4105
R8201 GNDA.n3890 GNDA.n3889 3.4105
R8202 GNDA.n3888 GNDA.n803 3.4105
R8203 GNDA.n888 GNDA.n885 3.4105
R8204 GNDA.n889 GNDA.n883 3.4105
R8205 GNDA.n890 GNDA.n882 3.4105
R8206 GNDA.n880 GNDA.n878 3.4105
R8207 GNDA.n894 GNDA.n877 3.4105
R8208 GNDA.n895 GNDA.n875 3.4105
R8209 GNDA.n896 GNDA.n874 3.4105
R8210 GNDA.n872 GNDA.n870 3.4105
R8211 GNDA.n900 GNDA.n869 3.4105
R8212 GNDA.n901 GNDA.n867 3.4105
R8213 GNDA.n902 GNDA.n866 3.4105
R8214 GNDA.n864 GNDA.n862 3.4105
R8215 GNDA.n906 GNDA.n861 3.4105
R8216 GNDA.n907 GNDA.n859 3.4105
R8217 GNDA.n908 GNDA.n858 3.4105
R8218 GNDA.n856 GNDA.n854 3.4105
R8219 GNDA.n912 GNDA.n853 3.4105
R8220 GNDA.n913 GNDA.n851 3.4105
R8221 GNDA.n914 GNDA.n850 3.4105
R8222 GNDA.n848 GNDA.n846 3.4105
R8223 GNDA.n918 GNDA.n845 3.4105
R8224 GNDA.n919 GNDA.n843 3.4105
R8225 GNDA.n920 GNDA.n842 3.4105
R8226 GNDA.n3655 GNDA.n3654 3.4105
R8227 GNDA.n3718 GNDA.n3717 3.4105
R8228 GNDA.n3716 GNDA.n3715 3.4105
R8229 GNDA.n3714 GNDA.n3659 3.4105
R8230 GNDA.n3658 GNDA.n3657 3.4105
R8231 GNDA.n3710 GNDA.n3709 3.4105
R8232 GNDA.n3708 GNDA.n3707 3.4105
R8233 GNDA.n3706 GNDA.n3663 3.4105
R8234 GNDA.n3662 GNDA.n3661 3.4105
R8235 GNDA.n3702 GNDA.n3701 3.4105
R8236 GNDA.n3700 GNDA.n3699 3.4105
R8237 GNDA.n3698 GNDA.n3667 3.4105
R8238 GNDA.n3666 GNDA.n3665 3.4105
R8239 GNDA.n3694 GNDA.n3693 3.4105
R8240 GNDA.n3692 GNDA.n3691 3.4105
R8241 GNDA.n3690 GNDA.n3671 3.4105
R8242 GNDA.n3670 GNDA.n3669 3.4105
R8243 GNDA.n3686 GNDA.n3685 3.4105
R8244 GNDA.n3684 GNDA.n3683 3.4105
R8245 GNDA.n3682 GNDA.n3675 3.4105
R8246 GNDA.n3674 GNDA.n3673 3.4105
R8247 GNDA.n3678 GNDA.n3677 3.4105
R8248 GNDA.n3676 GNDA.n3642 3.4105
R8249 GNDA.n3724 GNDA.n3723 3.4105
R8250 GNDA.n3787 GNDA.n3786 3.4105
R8251 GNDA.n3785 GNDA.n3784 3.4105
R8252 GNDA.n3783 GNDA.n3728 3.4105
R8253 GNDA.n3727 GNDA.n3726 3.4105
R8254 GNDA.n3779 GNDA.n3778 3.4105
R8255 GNDA.n3777 GNDA.n3776 3.4105
R8256 GNDA.n3775 GNDA.n3732 3.4105
R8257 GNDA.n3731 GNDA.n3730 3.4105
R8258 GNDA.n3771 GNDA.n3770 3.4105
R8259 GNDA.n3769 GNDA.n3768 3.4105
R8260 GNDA.n3767 GNDA.n3736 3.4105
R8261 GNDA.n3735 GNDA.n3734 3.4105
R8262 GNDA.n3763 GNDA.n3762 3.4105
R8263 GNDA.n3761 GNDA.n3760 3.4105
R8264 GNDA.n3759 GNDA.n3740 3.4105
R8265 GNDA.n3739 GNDA.n3738 3.4105
R8266 GNDA.n3755 GNDA.n3754 3.4105
R8267 GNDA.n3753 GNDA.n3752 3.4105
R8268 GNDA.n3751 GNDA.n3744 3.4105
R8269 GNDA.n3743 GNDA.n3742 3.4105
R8270 GNDA.n3747 GNDA.n3746 3.4105
R8271 GNDA.n3745 GNDA.n3630 3.4105
R8272 GNDA.n3793 GNDA.n3792 3.4105
R8273 GNDA.n3852 GNDA.n3851 3.4105
R8274 GNDA.n3850 GNDA.n3849 3.4105
R8275 GNDA.n3848 GNDA.n3847 3.4105
R8276 GNDA.n3846 GNDA.n3795 3.4105
R8277 GNDA.n3842 GNDA.n3841 3.4105
R8278 GNDA.n3840 GNDA.n3839 3.4105
R8279 GNDA.n3838 GNDA.n3837 3.4105
R8280 GNDA.n3836 GNDA.n3797 3.4105
R8281 GNDA.n3832 GNDA.n3831 3.4105
R8282 GNDA.n3830 GNDA.n3829 3.4105
R8283 GNDA.n3828 GNDA.n3827 3.4105
R8284 GNDA.n3826 GNDA.n3799 3.4105
R8285 GNDA.n3822 GNDA.n3821 3.4105
R8286 GNDA.n3820 GNDA.n3819 3.4105
R8287 GNDA.n3818 GNDA.n3817 3.4105
R8288 GNDA.n3816 GNDA.n3801 3.4105
R8289 GNDA.n3812 GNDA.n3811 3.4105
R8290 GNDA.n3810 GNDA.n3809 3.4105
R8291 GNDA.n3808 GNDA.n3807 3.4105
R8292 GNDA.n3806 GNDA.n3803 3.4105
R8293 GNDA.n938 GNDA.n937 3.4105
R8294 GNDA.n3858 GNDA.n3857 3.4105
R8295 GNDA.n3442 GNDA.n3439 3.4105
R8296 GNDA.n3443 GNDA.n3437 3.4105
R8297 GNDA.n3444 GNDA.n3436 3.4105
R8298 GNDA.n3434 GNDA.n3432 3.4105
R8299 GNDA.n3448 GNDA.n3431 3.4105
R8300 GNDA.n3449 GNDA.n3429 3.4105
R8301 GNDA.n3450 GNDA.n3428 3.4105
R8302 GNDA.n3426 GNDA.n3424 3.4105
R8303 GNDA.n3454 GNDA.n3423 3.4105
R8304 GNDA.n3455 GNDA.n3421 3.4105
R8305 GNDA.n3456 GNDA.n3420 3.4105
R8306 GNDA.n3418 GNDA.n3416 3.4105
R8307 GNDA.n3460 GNDA.n3415 3.4105
R8308 GNDA.n3461 GNDA.n3413 3.4105
R8309 GNDA.n3462 GNDA.n3412 3.4105
R8310 GNDA.n3410 GNDA.n3408 3.4105
R8311 GNDA.n3466 GNDA.n3407 3.4105
R8312 GNDA.n3467 GNDA.n3405 3.4105
R8313 GNDA.n3468 GNDA.n3404 3.4105
R8314 GNDA.n3402 GNDA.n3400 3.4105
R8315 GNDA.n3472 GNDA.n3399 3.4105
R8316 GNDA.n3473 GNDA.n3397 3.4105
R8317 GNDA.n3474 GNDA.n3396 3.4105
R8318 GNDA.n953 GNDA.n952 3.4105
R8319 GNDA.n3532 GNDA.n3531 3.4105
R8320 GNDA.n3530 GNDA.n3529 3.4105
R8321 GNDA.n3528 GNDA.n957 3.4105
R8322 GNDA.n956 GNDA.n955 3.4105
R8323 GNDA.n3524 GNDA.n3523 3.4105
R8324 GNDA.n3522 GNDA.n3521 3.4105
R8325 GNDA.n3520 GNDA.n961 3.4105
R8326 GNDA.n960 GNDA.n959 3.4105
R8327 GNDA.n3516 GNDA.n3515 3.4105
R8328 GNDA.n3514 GNDA.n3513 3.4105
R8329 GNDA.n3512 GNDA.n965 3.4105
R8330 GNDA.n964 GNDA.n963 3.4105
R8331 GNDA.n3508 GNDA.n3507 3.4105
R8332 GNDA.n3506 GNDA.n3505 3.4105
R8333 GNDA.n3504 GNDA.n969 3.4105
R8334 GNDA.n968 GNDA.n967 3.4105
R8335 GNDA.n3500 GNDA.n3499 3.4105
R8336 GNDA.n3498 GNDA.n3497 3.4105
R8337 GNDA.n3496 GNDA.n973 3.4105
R8338 GNDA.n972 GNDA.n971 3.4105
R8339 GNDA.n3492 GNDA.n3491 3.4105
R8340 GNDA.n3490 GNDA.n940 3.4105
R8341 GNDA.n2790 GNDA.n2789 3.4105
R8342 GNDA.n2853 GNDA.n2852 3.4105
R8343 GNDA.n2851 GNDA.n2850 3.4105
R8344 GNDA.n2849 GNDA.n2794 3.4105
R8345 GNDA.n2793 GNDA.n2792 3.4105
R8346 GNDA.n2845 GNDA.n2844 3.4105
R8347 GNDA.n2843 GNDA.n2842 3.4105
R8348 GNDA.n2841 GNDA.n2798 3.4105
R8349 GNDA.n2797 GNDA.n2796 3.4105
R8350 GNDA.n2837 GNDA.n2836 3.4105
R8351 GNDA.n2835 GNDA.n2834 3.4105
R8352 GNDA.n2833 GNDA.n2802 3.4105
R8353 GNDA.n2801 GNDA.n2800 3.4105
R8354 GNDA.n2829 GNDA.n2828 3.4105
R8355 GNDA.n2827 GNDA.n2826 3.4105
R8356 GNDA.n2825 GNDA.n2806 3.4105
R8357 GNDA.n2805 GNDA.n2804 3.4105
R8358 GNDA.n2821 GNDA.n2820 3.4105
R8359 GNDA.n2819 GNDA.n2818 3.4105
R8360 GNDA.n2817 GNDA.n2810 3.4105
R8361 GNDA.n2809 GNDA.n2808 3.4105
R8362 GNDA.n2813 GNDA.n2812 3.4105
R8363 GNDA.n2811 GNDA.n2777 3.4105
R8364 GNDA.n2859 GNDA.n2858 3.4105
R8365 GNDA.n2922 GNDA.n2921 3.4105
R8366 GNDA.n2920 GNDA.n2919 3.4105
R8367 GNDA.n2918 GNDA.n2863 3.4105
R8368 GNDA.n2862 GNDA.n2861 3.4105
R8369 GNDA.n2914 GNDA.n2913 3.4105
R8370 GNDA.n2912 GNDA.n2911 3.4105
R8371 GNDA.n2910 GNDA.n2867 3.4105
R8372 GNDA.n2866 GNDA.n2865 3.4105
R8373 GNDA.n2906 GNDA.n2905 3.4105
R8374 GNDA.n2904 GNDA.n2903 3.4105
R8375 GNDA.n2902 GNDA.n2871 3.4105
R8376 GNDA.n2870 GNDA.n2869 3.4105
R8377 GNDA.n2898 GNDA.n2897 3.4105
R8378 GNDA.n2896 GNDA.n2895 3.4105
R8379 GNDA.n2894 GNDA.n2875 3.4105
R8380 GNDA.n2874 GNDA.n2873 3.4105
R8381 GNDA.n2890 GNDA.n2889 3.4105
R8382 GNDA.n2888 GNDA.n2887 3.4105
R8383 GNDA.n2886 GNDA.n2879 3.4105
R8384 GNDA.n2878 GNDA.n2877 3.4105
R8385 GNDA.n2882 GNDA.n2881 3.4105
R8386 GNDA.n2880 GNDA.n2765 3.4105
R8387 GNDA.n2928 GNDA.n2927 3.4105
R8388 GNDA.n2991 GNDA.n2990 3.4105
R8389 GNDA.n2989 GNDA.n2988 3.4105
R8390 GNDA.n2987 GNDA.n2932 3.4105
R8391 GNDA.n2931 GNDA.n2930 3.4105
R8392 GNDA.n2983 GNDA.n2982 3.4105
R8393 GNDA.n2981 GNDA.n2980 3.4105
R8394 GNDA.n2979 GNDA.n2936 3.4105
R8395 GNDA.n2935 GNDA.n2934 3.4105
R8396 GNDA.n2975 GNDA.n2974 3.4105
R8397 GNDA.n2973 GNDA.n2972 3.4105
R8398 GNDA.n2971 GNDA.n2940 3.4105
R8399 GNDA.n2939 GNDA.n2938 3.4105
R8400 GNDA.n2967 GNDA.n2966 3.4105
R8401 GNDA.n2965 GNDA.n2964 3.4105
R8402 GNDA.n2963 GNDA.n2944 3.4105
R8403 GNDA.n2943 GNDA.n2942 3.4105
R8404 GNDA.n2959 GNDA.n2958 3.4105
R8405 GNDA.n2957 GNDA.n2956 3.4105
R8406 GNDA.n2955 GNDA.n2948 3.4105
R8407 GNDA.n2947 GNDA.n2946 3.4105
R8408 GNDA.n2951 GNDA.n2950 3.4105
R8409 GNDA.n2949 GNDA.n2753 3.4105
R8410 GNDA.n2997 GNDA.n2996 3.4105
R8411 GNDA.n3060 GNDA.n3059 3.4105
R8412 GNDA.n3058 GNDA.n3057 3.4105
R8413 GNDA.n3056 GNDA.n3001 3.4105
R8414 GNDA.n3000 GNDA.n2999 3.4105
R8415 GNDA.n3052 GNDA.n3051 3.4105
R8416 GNDA.n3050 GNDA.n3049 3.4105
R8417 GNDA.n3048 GNDA.n3005 3.4105
R8418 GNDA.n3004 GNDA.n3003 3.4105
R8419 GNDA.n3044 GNDA.n3043 3.4105
R8420 GNDA.n3042 GNDA.n3041 3.4105
R8421 GNDA.n3040 GNDA.n3009 3.4105
R8422 GNDA.n3008 GNDA.n3007 3.4105
R8423 GNDA.n3036 GNDA.n3035 3.4105
R8424 GNDA.n3034 GNDA.n3033 3.4105
R8425 GNDA.n3032 GNDA.n3013 3.4105
R8426 GNDA.n3012 GNDA.n3011 3.4105
R8427 GNDA.n3028 GNDA.n3027 3.4105
R8428 GNDA.n3026 GNDA.n3025 3.4105
R8429 GNDA.n3024 GNDA.n3017 3.4105
R8430 GNDA.n3016 GNDA.n3015 3.4105
R8431 GNDA.n3020 GNDA.n3019 3.4105
R8432 GNDA.n3018 GNDA.n2741 3.4105
R8433 GNDA.n3066 GNDA.n3065 3.4105
R8434 GNDA.n3129 GNDA.n3128 3.4105
R8435 GNDA.n3127 GNDA.n3126 3.4105
R8436 GNDA.n3125 GNDA.n3070 3.4105
R8437 GNDA.n3069 GNDA.n3068 3.4105
R8438 GNDA.n3121 GNDA.n3120 3.4105
R8439 GNDA.n3119 GNDA.n3118 3.4105
R8440 GNDA.n3117 GNDA.n3074 3.4105
R8441 GNDA.n3073 GNDA.n3072 3.4105
R8442 GNDA.n3113 GNDA.n3112 3.4105
R8443 GNDA.n3111 GNDA.n3110 3.4105
R8444 GNDA.n3109 GNDA.n3078 3.4105
R8445 GNDA.n3077 GNDA.n3076 3.4105
R8446 GNDA.n3105 GNDA.n3104 3.4105
R8447 GNDA.n3103 GNDA.n3102 3.4105
R8448 GNDA.n3101 GNDA.n3082 3.4105
R8449 GNDA.n3081 GNDA.n3080 3.4105
R8450 GNDA.n3097 GNDA.n3096 3.4105
R8451 GNDA.n3095 GNDA.n3094 3.4105
R8452 GNDA.n3093 GNDA.n3086 3.4105
R8453 GNDA.n3085 GNDA.n3084 3.4105
R8454 GNDA.n3089 GNDA.n3088 3.4105
R8455 GNDA.n3087 GNDA.n2729 3.4105
R8456 GNDA.n3135 GNDA.n3134 3.4105
R8457 GNDA.n3198 GNDA.n3197 3.4105
R8458 GNDA.n3196 GNDA.n3195 3.4105
R8459 GNDA.n3194 GNDA.n3139 3.4105
R8460 GNDA.n3138 GNDA.n3137 3.4105
R8461 GNDA.n3190 GNDA.n3189 3.4105
R8462 GNDA.n3188 GNDA.n3187 3.4105
R8463 GNDA.n3186 GNDA.n3143 3.4105
R8464 GNDA.n3142 GNDA.n3141 3.4105
R8465 GNDA.n3182 GNDA.n3181 3.4105
R8466 GNDA.n3180 GNDA.n3179 3.4105
R8467 GNDA.n3178 GNDA.n3147 3.4105
R8468 GNDA.n3146 GNDA.n3145 3.4105
R8469 GNDA.n3174 GNDA.n3173 3.4105
R8470 GNDA.n3172 GNDA.n3171 3.4105
R8471 GNDA.n3170 GNDA.n3151 3.4105
R8472 GNDA.n3150 GNDA.n3149 3.4105
R8473 GNDA.n3166 GNDA.n3165 3.4105
R8474 GNDA.n3164 GNDA.n3163 3.4105
R8475 GNDA.n3162 GNDA.n3155 3.4105
R8476 GNDA.n3154 GNDA.n3153 3.4105
R8477 GNDA.n3158 GNDA.n3157 3.4105
R8478 GNDA.n3156 GNDA.n2717 3.4105
R8479 GNDA.n3204 GNDA.n3203 3.4105
R8480 GNDA.n3267 GNDA.n3266 3.4105
R8481 GNDA.n3265 GNDA.n3264 3.4105
R8482 GNDA.n3263 GNDA.n3208 3.4105
R8483 GNDA.n3207 GNDA.n3206 3.4105
R8484 GNDA.n3259 GNDA.n3258 3.4105
R8485 GNDA.n3257 GNDA.n3256 3.4105
R8486 GNDA.n3255 GNDA.n3212 3.4105
R8487 GNDA.n3211 GNDA.n3210 3.4105
R8488 GNDA.n3251 GNDA.n3250 3.4105
R8489 GNDA.n3249 GNDA.n3248 3.4105
R8490 GNDA.n3247 GNDA.n3216 3.4105
R8491 GNDA.n3215 GNDA.n3214 3.4105
R8492 GNDA.n3243 GNDA.n3242 3.4105
R8493 GNDA.n3241 GNDA.n3240 3.4105
R8494 GNDA.n3239 GNDA.n3220 3.4105
R8495 GNDA.n3219 GNDA.n3218 3.4105
R8496 GNDA.n3235 GNDA.n3234 3.4105
R8497 GNDA.n3233 GNDA.n3232 3.4105
R8498 GNDA.n3231 GNDA.n3224 3.4105
R8499 GNDA.n3223 GNDA.n3222 3.4105
R8500 GNDA.n3227 GNDA.n3226 3.4105
R8501 GNDA.n3225 GNDA.n2705 3.4105
R8502 GNDA.n3273 GNDA.n3272 3.4105
R8503 GNDA.n3332 GNDA.n3331 3.4105
R8504 GNDA.n3330 GNDA.n3329 3.4105
R8505 GNDA.n3328 GNDA.n3327 3.4105
R8506 GNDA.n3326 GNDA.n3275 3.4105
R8507 GNDA.n3322 GNDA.n3321 3.4105
R8508 GNDA.n3320 GNDA.n3319 3.4105
R8509 GNDA.n3318 GNDA.n3317 3.4105
R8510 GNDA.n3316 GNDA.n3277 3.4105
R8511 GNDA.n3312 GNDA.n3311 3.4105
R8512 GNDA.n3310 GNDA.n3309 3.4105
R8513 GNDA.n3308 GNDA.n3307 3.4105
R8514 GNDA.n3306 GNDA.n3279 3.4105
R8515 GNDA.n3302 GNDA.n3301 3.4105
R8516 GNDA.n3300 GNDA.n3299 3.4105
R8517 GNDA.n3298 GNDA.n3297 3.4105
R8518 GNDA.n3296 GNDA.n3281 3.4105
R8519 GNDA.n3292 GNDA.n3291 3.4105
R8520 GNDA.n3290 GNDA.n3289 3.4105
R8521 GNDA.n3288 GNDA.n3287 3.4105
R8522 GNDA.n3286 GNDA.n3283 3.4105
R8523 GNDA.n1040 GNDA.n1039 3.4105
R8524 GNDA.n3338 GNDA.n3337 3.4105
R8525 GNDA.n3337 GNDA.n3336 3.4105
R8526 GNDA.n3336 GNDA.n3335 3.4105
R8527 GNDA.n3271 GNDA.n2705 3.4105
R8528 GNDA.n3271 GNDA.n3270 3.4105
R8529 GNDA.n3202 GNDA.n2717 3.4105
R8530 GNDA.n3202 GNDA.n3201 3.4105
R8531 GNDA.n3133 GNDA.n2729 3.4105
R8532 GNDA.n3133 GNDA.n3132 3.4105
R8533 GNDA.n3064 GNDA.n2741 3.4105
R8534 GNDA.n3064 GNDA.n3063 3.4105
R8535 GNDA.n2995 GNDA.n2753 3.4105
R8536 GNDA.n2995 GNDA.n2994 3.4105
R8537 GNDA.n2926 GNDA.n2765 3.4105
R8538 GNDA.n2926 GNDA.n2925 3.4105
R8539 GNDA.n2857 GNDA.n2777 3.4105
R8540 GNDA.n2857 GNDA.n2856 3.4105
R8541 GNDA.n3536 GNDA.n940 3.4105
R8542 GNDA.n3536 GNDA.n3535 3.4105
R8543 GNDA.n3857 GNDA.n3856 3.4105
R8544 GNDA.n3856 GNDA.n3855 3.4105
R8545 GNDA.n3791 GNDA.n3630 3.4105
R8546 GNDA.n3791 GNDA.n3790 3.4105
R8547 GNDA.n3722 GNDA.n3642 3.4105
R8548 GNDA.n3722 GNDA.n3721 3.4105
R8549 GNDA.n842 GNDA.n802 3.4105
R8550 GNDA.n886 GNDA.n802 3.4105
R8551 GNDA.n3934 GNDA.n803 3.4105
R8552 GNDA.n3934 GNDA.n3933 3.4105
R8553 GNDA.n3396 GNDA.n939 3.4105
R8554 GNDA.n3440 GNDA.n939 3.4105
R8555 GNDA.n3618 GNDA.n3537 3.4105
R8556 GNDA.n3618 GNDA.n3617 3.4105
R8557 GNDA.n3951 GNDA.n774 3.4105
R8558 GNDA.n3952 GNDA.n3951 3.4105
R8559 GNDA.n4195 GNDA.n487 3.4105
R8560 GNDA.n4195 GNDA.n4194 3.4105
R8561 GNDA.n4362 GNDA.n446 3.4105
R8562 GNDA.n4328 GNDA.n446 3.4105
R8563 GNDA.n4432 GNDA.n447 3.4105
R8564 GNDA.n4432 GNDA.n4431 3.4105
R8565 GNDA.n4873 GNDA.n4872 3.4105
R8566 GNDA.n4872 GNDA.n4871 3.4105
R8567 GNDA.n4272 GNDA.n4271 3.4105
R8568 GNDA.n4271 GNDA.n4270 3.4105
R8569 GNDA.n4807 GNDA.n4444 3.4105
R8570 GNDA.n4807 GNDA.n4806 3.4105
R8571 GNDA.n4550 GNDA.n4456 3.4105
R8572 GNDA.n4516 GNDA.n4456 3.4105
R8573 GNDA.n4647 GNDA.n4566 3.4105
R8574 GNDA.n4647 GNDA.n4646 3.4105
R8575 GNDA.n4724 GNDA.n4723 3.4105
R8576 GNDA.n4723 GNDA.n4722 3.4105
R8577 GNDA.n560 GNDA.n557 3.4105
R8578 GNDA.n561 GNDA.n556 3.4105
R8579 GNDA.n562 GNDA.n554 3.4105
R8580 GNDA.n553 GNDA.n550 3.4105
R8581 GNDA.n566 GNDA.n549 3.4105
R8582 GNDA.n567 GNDA.n548 3.4105
R8583 GNDA.n568 GNDA.n546 3.4105
R8584 GNDA.n545 GNDA.n542 3.4105
R8585 GNDA.n572 GNDA.n541 3.4105
R8586 GNDA.n573 GNDA.n540 3.4105
R8587 GNDA.n574 GNDA.n538 3.4105
R8588 GNDA.n537 GNDA.n534 3.4105
R8589 GNDA.n578 GNDA.n533 3.4105
R8590 GNDA.n579 GNDA.n532 3.4105
R8591 GNDA.n580 GNDA.n530 3.4105
R8592 GNDA.n529 GNDA.n526 3.4105
R8593 GNDA.n584 GNDA.n525 3.4105
R8594 GNDA.n585 GNDA.n524 3.4105
R8595 GNDA.n586 GNDA.n522 3.4105
R8596 GNDA.n521 GNDA.n518 3.4105
R8597 GNDA.n590 GNDA.n517 3.4105
R8598 GNDA.n591 GNDA.n516 3.4105
R8599 GNDA.n1543 GNDA.n1467 3.4105
R8600 GNDA.n1541 GNDA.n1540 3.4105
R8601 GNDA.n1469 GNDA.n1468 3.4105
R8602 GNDA.n1536 GNDA.n1535 3.4105
R8603 GNDA.n1533 GNDA.n1471 3.4105
R8604 GNDA.n1531 GNDA.n1530 3.4105
R8605 GNDA.n1473 GNDA.n1472 3.4105
R8606 GNDA.n1526 GNDA.n1525 3.4105
R8607 GNDA.n1523 GNDA.n1475 3.4105
R8608 GNDA.n1521 GNDA.n1520 3.4105
R8609 GNDA.n1477 GNDA.n1476 3.4105
R8610 GNDA.n1516 GNDA.n1515 3.4105
R8611 GNDA.n1513 GNDA.n1479 3.4105
R8612 GNDA.n1511 GNDA.n1510 3.4105
R8613 GNDA.n1481 GNDA.n1480 3.4105
R8614 GNDA.n1506 GNDA.n1505 3.4105
R8615 GNDA.n1503 GNDA.n1483 3.4105
R8616 GNDA.n1501 GNDA.n1500 3.4105
R8617 GNDA.n1485 GNDA.n1484 3.4105
R8618 GNDA.n1496 GNDA.n1495 3.4105
R8619 GNDA.n1493 GNDA.n1487 3.4105
R8620 GNDA.n1491 GNDA.n1490 3.4105
R8621 GNDA.n1545 GNDA.n1544 3.4105
R8622 GNDA.n1351 GNDA.n1350 3.4105
R8623 GNDA.n1413 GNDA.n1412 3.4105
R8624 GNDA.n1411 GNDA.n1410 3.4105
R8625 GNDA.n1409 GNDA.n1408 3.4105
R8626 GNDA.n1407 GNDA.n1353 3.4105
R8627 GNDA.n1403 GNDA.n1402 3.4105
R8628 GNDA.n1401 GNDA.n1400 3.4105
R8629 GNDA.n1399 GNDA.n1398 3.4105
R8630 GNDA.n1397 GNDA.n1355 3.4105
R8631 GNDA.n1393 GNDA.n1392 3.4105
R8632 GNDA.n1391 GNDA.n1390 3.4105
R8633 GNDA.n1389 GNDA.n1388 3.4105
R8634 GNDA.n1387 GNDA.n1357 3.4105
R8635 GNDA.n1383 GNDA.n1382 3.4105
R8636 GNDA.n1381 GNDA.n1380 3.4105
R8637 GNDA.n1379 GNDA.n1378 3.4105
R8638 GNDA.n1377 GNDA.n1359 3.4105
R8639 GNDA.n1373 GNDA.n1372 3.4105
R8640 GNDA.n1371 GNDA.n1370 3.4105
R8641 GNDA.n1369 GNDA.n1368 3.4105
R8642 GNDA.n1367 GNDA.n1361 3.4105
R8643 GNDA.n1363 GNDA.n1362 3.4105
R8644 GNDA.n2578 GNDA.n2577 3.4105
R8645 GNDA.n2579 GNDA.n1337 3.4105
R8646 GNDA.n2579 GNDA.n2578 3.4105
R8647 GNDA.n1488 GNDA.n1349 3.4105
R8648 GNDA.n1544 GNDA.n1349 3.4105
R8649 GNDA.n1320 GNDA.n1287 3.4105
R8650 GNDA.n2583 GNDA.n1287 3.4105
R8651 GNDA.n2583 GNDA.n1269 3.4105
R8652 GNDA.n1320 GNDA.n1289 3.4105
R8653 GNDA.n1289 GNDA.n1222 3.4105
R8654 GNDA.n1289 GNDA.n1220 3.4105
R8655 GNDA.n1289 GNDA.n1223 3.4105
R8656 GNDA.n1289 GNDA.n1219 3.4105
R8657 GNDA.n1289 GNDA.n1224 3.4105
R8658 GNDA.n1289 GNDA.n1218 3.4105
R8659 GNDA.n1289 GNDA.n1225 3.4105
R8660 GNDA.n1289 GNDA.n1217 3.4105
R8661 GNDA.n1289 GNDA.n1226 3.4105
R8662 GNDA.n1289 GNDA.n1216 3.4105
R8663 GNDA.n1289 GNDA.n1227 3.4105
R8664 GNDA.n1289 GNDA.n1215 3.4105
R8665 GNDA.n1289 GNDA.n1228 3.4105
R8666 GNDA.n1289 GNDA.n1214 3.4105
R8667 GNDA.n1289 GNDA.n1229 3.4105
R8668 GNDA.n1289 GNDA.n1213 3.4105
R8669 GNDA.n1289 GNDA.n1230 3.4105
R8670 GNDA.n1289 GNDA.n1212 3.4105
R8671 GNDA.n1289 GNDA.n1231 3.4105
R8672 GNDA.n1289 GNDA.n1211 3.4105
R8673 GNDA.n1289 GNDA.n1232 3.4105
R8674 GNDA.n1289 GNDA.n1210 3.4105
R8675 GNDA.n1289 GNDA.n1233 3.4105
R8676 GNDA.n1289 GNDA.n1209 3.4105
R8677 GNDA.n1289 GNDA.n1234 3.4105
R8678 GNDA.n1289 GNDA.n1208 3.4105
R8679 GNDA.n1289 GNDA.n1235 3.4105
R8680 GNDA.n1289 GNDA.n1207 3.4105
R8681 GNDA.n1289 GNDA.n1236 3.4105
R8682 GNDA.n1289 GNDA.n1206 3.4105
R8683 GNDA.n1289 GNDA.n1237 3.4105
R8684 GNDA.n2583 GNDA.n1289 3.4105
R8685 GNDA.n1320 GNDA.n1253 3.4105
R8686 GNDA.n1253 GNDA.n1222 3.4105
R8687 GNDA.n1253 GNDA.n1220 3.4105
R8688 GNDA.n1253 GNDA.n1223 3.4105
R8689 GNDA.n1253 GNDA.n1219 3.4105
R8690 GNDA.n1253 GNDA.n1224 3.4105
R8691 GNDA.n1253 GNDA.n1218 3.4105
R8692 GNDA.n1253 GNDA.n1225 3.4105
R8693 GNDA.n1253 GNDA.n1217 3.4105
R8694 GNDA.n1253 GNDA.n1226 3.4105
R8695 GNDA.n1253 GNDA.n1216 3.4105
R8696 GNDA.n1253 GNDA.n1227 3.4105
R8697 GNDA.n1253 GNDA.n1215 3.4105
R8698 GNDA.n1253 GNDA.n1228 3.4105
R8699 GNDA.n1253 GNDA.n1214 3.4105
R8700 GNDA.n1253 GNDA.n1229 3.4105
R8701 GNDA.n1253 GNDA.n1213 3.4105
R8702 GNDA.n1253 GNDA.n1230 3.4105
R8703 GNDA.n1253 GNDA.n1212 3.4105
R8704 GNDA.n1253 GNDA.n1231 3.4105
R8705 GNDA.n1253 GNDA.n1211 3.4105
R8706 GNDA.n1253 GNDA.n1232 3.4105
R8707 GNDA.n1253 GNDA.n1210 3.4105
R8708 GNDA.n1253 GNDA.n1233 3.4105
R8709 GNDA.n1253 GNDA.n1209 3.4105
R8710 GNDA.n1253 GNDA.n1234 3.4105
R8711 GNDA.n1253 GNDA.n1208 3.4105
R8712 GNDA.n1253 GNDA.n1235 3.4105
R8713 GNDA.n1253 GNDA.n1207 3.4105
R8714 GNDA.n1253 GNDA.n1236 3.4105
R8715 GNDA.n1253 GNDA.n1206 3.4105
R8716 GNDA.n1253 GNDA.n1237 3.4105
R8717 GNDA.n2583 GNDA.n1253 3.4105
R8718 GNDA.n1320 GNDA.n1291 3.4105
R8719 GNDA.n1291 GNDA.n1222 3.4105
R8720 GNDA.n1291 GNDA.n1220 3.4105
R8721 GNDA.n1291 GNDA.n1223 3.4105
R8722 GNDA.n1291 GNDA.n1219 3.4105
R8723 GNDA.n1291 GNDA.n1224 3.4105
R8724 GNDA.n1291 GNDA.n1218 3.4105
R8725 GNDA.n1291 GNDA.n1225 3.4105
R8726 GNDA.n1291 GNDA.n1217 3.4105
R8727 GNDA.n1291 GNDA.n1226 3.4105
R8728 GNDA.n1291 GNDA.n1216 3.4105
R8729 GNDA.n1291 GNDA.n1227 3.4105
R8730 GNDA.n1291 GNDA.n1215 3.4105
R8731 GNDA.n1291 GNDA.n1228 3.4105
R8732 GNDA.n1291 GNDA.n1214 3.4105
R8733 GNDA.n1291 GNDA.n1229 3.4105
R8734 GNDA.n1291 GNDA.n1213 3.4105
R8735 GNDA.n1291 GNDA.n1230 3.4105
R8736 GNDA.n1291 GNDA.n1212 3.4105
R8737 GNDA.n1291 GNDA.n1231 3.4105
R8738 GNDA.n1291 GNDA.n1211 3.4105
R8739 GNDA.n1291 GNDA.n1232 3.4105
R8740 GNDA.n1291 GNDA.n1210 3.4105
R8741 GNDA.n1291 GNDA.n1233 3.4105
R8742 GNDA.n1291 GNDA.n1209 3.4105
R8743 GNDA.n1291 GNDA.n1234 3.4105
R8744 GNDA.n1291 GNDA.n1208 3.4105
R8745 GNDA.n1291 GNDA.n1235 3.4105
R8746 GNDA.n1291 GNDA.n1207 3.4105
R8747 GNDA.n1291 GNDA.n1236 3.4105
R8748 GNDA.n1291 GNDA.n1206 3.4105
R8749 GNDA.n1291 GNDA.n1237 3.4105
R8750 GNDA.n2583 GNDA.n1291 3.4105
R8751 GNDA.n1320 GNDA.n1252 3.4105
R8752 GNDA.n1252 GNDA.n1222 3.4105
R8753 GNDA.n1252 GNDA.n1220 3.4105
R8754 GNDA.n1252 GNDA.n1223 3.4105
R8755 GNDA.n1252 GNDA.n1219 3.4105
R8756 GNDA.n1252 GNDA.n1224 3.4105
R8757 GNDA.n1252 GNDA.n1218 3.4105
R8758 GNDA.n1252 GNDA.n1225 3.4105
R8759 GNDA.n1252 GNDA.n1217 3.4105
R8760 GNDA.n1252 GNDA.n1226 3.4105
R8761 GNDA.n1252 GNDA.n1216 3.4105
R8762 GNDA.n1252 GNDA.n1227 3.4105
R8763 GNDA.n1252 GNDA.n1215 3.4105
R8764 GNDA.n1252 GNDA.n1228 3.4105
R8765 GNDA.n1252 GNDA.n1214 3.4105
R8766 GNDA.n1252 GNDA.n1229 3.4105
R8767 GNDA.n1252 GNDA.n1213 3.4105
R8768 GNDA.n1252 GNDA.n1230 3.4105
R8769 GNDA.n1252 GNDA.n1212 3.4105
R8770 GNDA.n1252 GNDA.n1231 3.4105
R8771 GNDA.n1252 GNDA.n1211 3.4105
R8772 GNDA.n1252 GNDA.n1232 3.4105
R8773 GNDA.n1252 GNDA.n1210 3.4105
R8774 GNDA.n1252 GNDA.n1233 3.4105
R8775 GNDA.n1252 GNDA.n1209 3.4105
R8776 GNDA.n1252 GNDA.n1234 3.4105
R8777 GNDA.n1252 GNDA.n1208 3.4105
R8778 GNDA.n1252 GNDA.n1235 3.4105
R8779 GNDA.n1252 GNDA.n1207 3.4105
R8780 GNDA.n1252 GNDA.n1236 3.4105
R8781 GNDA.n1252 GNDA.n1206 3.4105
R8782 GNDA.n1252 GNDA.n1237 3.4105
R8783 GNDA.n2583 GNDA.n1252 3.4105
R8784 GNDA.n1320 GNDA.n1293 3.4105
R8785 GNDA.n1293 GNDA.n1222 3.4105
R8786 GNDA.n1293 GNDA.n1220 3.4105
R8787 GNDA.n1293 GNDA.n1223 3.4105
R8788 GNDA.n1293 GNDA.n1219 3.4105
R8789 GNDA.n1293 GNDA.n1224 3.4105
R8790 GNDA.n1293 GNDA.n1218 3.4105
R8791 GNDA.n1293 GNDA.n1225 3.4105
R8792 GNDA.n1293 GNDA.n1217 3.4105
R8793 GNDA.n1293 GNDA.n1226 3.4105
R8794 GNDA.n1293 GNDA.n1216 3.4105
R8795 GNDA.n1293 GNDA.n1227 3.4105
R8796 GNDA.n1293 GNDA.n1215 3.4105
R8797 GNDA.n1293 GNDA.n1228 3.4105
R8798 GNDA.n1293 GNDA.n1214 3.4105
R8799 GNDA.n1293 GNDA.n1229 3.4105
R8800 GNDA.n1293 GNDA.n1213 3.4105
R8801 GNDA.n1293 GNDA.n1230 3.4105
R8802 GNDA.n1293 GNDA.n1212 3.4105
R8803 GNDA.n1293 GNDA.n1231 3.4105
R8804 GNDA.n1293 GNDA.n1211 3.4105
R8805 GNDA.n1293 GNDA.n1232 3.4105
R8806 GNDA.n1293 GNDA.n1210 3.4105
R8807 GNDA.n1293 GNDA.n1233 3.4105
R8808 GNDA.n1293 GNDA.n1209 3.4105
R8809 GNDA.n1293 GNDA.n1234 3.4105
R8810 GNDA.n1293 GNDA.n1208 3.4105
R8811 GNDA.n1293 GNDA.n1235 3.4105
R8812 GNDA.n1293 GNDA.n1207 3.4105
R8813 GNDA.n1293 GNDA.n1236 3.4105
R8814 GNDA.n1293 GNDA.n1206 3.4105
R8815 GNDA.n1293 GNDA.n1237 3.4105
R8816 GNDA.n2583 GNDA.n1293 3.4105
R8817 GNDA.n1320 GNDA.n1251 3.4105
R8818 GNDA.n1251 GNDA.n1222 3.4105
R8819 GNDA.n1251 GNDA.n1220 3.4105
R8820 GNDA.n1251 GNDA.n1223 3.4105
R8821 GNDA.n1251 GNDA.n1219 3.4105
R8822 GNDA.n1251 GNDA.n1224 3.4105
R8823 GNDA.n1251 GNDA.n1218 3.4105
R8824 GNDA.n1251 GNDA.n1225 3.4105
R8825 GNDA.n1251 GNDA.n1217 3.4105
R8826 GNDA.n1251 GNDA.n1226 3.4105
R8827 GNDA.n1251 GNDA.n1216 3.4105
R8828 GNDA.n1251 GNDA.n1227 3.4105
R8829 GNDA.n1251 GNDA.n1215 3.4105
R8830 GNDA.n1251 GNDA.n1228 3.4105
R8831 GNDA.n1251 GNDA.n1214 3.4105
R8832 GNDA.n1251 GNDA.n1229 3.4105
R8833 GNDA.n1251 GNDA.n1213 3.4105
R8834 GNDA.n1251 GNDA.n1230 3.4105
R8835 GNDA.n1251 GNDA.n1212 3.4105
R8836 GNDA.n1251 GNDA.n1231 3.4105
R8837 GNDA.n1251 GNDA.n1211 3.4105
R8838 GNDA.n1251 GNDA.n1232 3.4105
R8839 GNDA.n1251 GNDA.n1210 3.4105
R8840 GNDA.n1251 GNDA.n1233 3.4105
R8841 GNDA.n1251 GNDA.n1209 3.4105
R8842 GNDA.n1251 GNDA.n1234 3.4105
R8843 GNDA.n1251 GNDA.n1208 3.4105
R8844 GNDA.n1251 GNDA.n1235 3.4105
R8845 GNDA.n1251 GNDA.n1207 3.4105
R8846 GNDA.n1251 GNDA.n1236 3.4105
R8847 GNDA.n1251 GNDA.n1206 3.4105
R8848 GNDA.n1251 GNDA.n1237 3.4105
R8849 GNDA.n2583 GNDA.n1251 3.4105
R8850 GNDA.n1320 GNDA.n1295 3.4105
R8851 GNDA.n1295 GNDA.n1222 3.4105
R8852 GNDA.n1295 GNDA.n1220 3.4105
R8853 GNDA.n1295 GNDA.n1223 3.4105
R8854 GNDA.n1295 GNDA.n1219 3.4105
R8855 GNDA.n1295 GNDA.n1224 3.4105
R8856 GNDA.n1295 GNDA.n1218 3.4105
R8857 GNDA.n1295 GNDA.n1225 3.4105
R8858 GNDA.n1295 GNDA.n1217 3.4105
R8859 GNDA.n1295 GNDA.n1226 3.4105
R8860 GNDA.n1295 GNDA.n1216 3.4105
R8861 GNDA.n1295 GNDA.n1227 3.4105
R8862 GNDA.n1295 GNDA.n1215 3.4105
R8863 GNDA.n1295 GNDA.n1228 3.4105
R8864 GNDA.n1295 GNDA.n1214 3.4105
R8865 GNDA.n1295 GNDA.n1229 3.4105
R8866 GNDA.n1295 GNDA.n1213 3.4105
R8867 GNDA.n1295 GNDA.n1230 3.4105
R8868 GNDA.n1295 GNDA.n1212 3.4105
R8869 GNDA.n1295 GNDA.n1231 3.4105
R8870 GNDA.n1295 GNDA.n1211 3.4105
R8871 GNDA.n1295 GNDA.n1232 3.4105
R8872 GNDA.n1295 GNDA.n1210 3.4105
R8873 GNDA.n1295 GNDA.n1233 3.4105
R8874 GNDA.n1295 GNDA.n1209 3.4105
R8875 GNDA.n1295 GNDA.n1234 3.4105
R8876 GNDA.n1295 GNDA.n1208 3.4105
R8877 GNDA.n1295 GNDA.n1235 3.4105
R8878 GNDA.n1295 GNDA.n1207 3.4105
R8879 GNDA.n1295 GNDA.n1236 3.4105
R8880 GNDA.n1295 GNDA.n1206 3.4105
R8881 GNDA.n1295 GNDA.n1237 3.4105
R8882 GNDA.n2583 GNDA.n1295 3.4105
R8883 GNDA.n1320 GNDA.n1250 3.4105
R8884 GNDA.n1250 GNDA.n1222 3.4105
R8885 GNDA.n1250 GNDA.n1220 3.4105
R8886 GNDA.n1250 GNDA.n1223 3.4105
R8887 GNDA.n1250 GNDA.n1219 3.4105
R8888 GNDA.n1250 GNDA.n1224 3.4105
R8889 GNDA.n1250 GNDA.n1218 3.4105
R8890 GNDA.n1250 GNDA.n1225 3.4105
R8891 GNDA.n1250 GNDA.n1217 3.4105
R8892 GNDA.n1250 GNDA.n1226 3.4105
R8893 GNDA.n1250 GNDA.n1216 3.4105
R8894 GNDA.n1250 GNDA.n1227 3.4105
R8895 GNDA.n1250 GNDA.n1215 3.4105
R8896 GNDA.n1250 GNDA.n1228 3.4105
R8897 GNDA.n1250 GNDA.n1214 3.4105
R8898 GNDA.n1250 GNDA.n1229 3.4105
R8899 GNDA.n1250 GNDA.n1213 3.4105
R8900 GNDA.n1250 GNDA.n1230 3.4105
R8901 GNDA.n1250 GNDA.n1212 3.4105
R8902 GNDA.n1250 GNDA.n1231 3.4105
R8903 GNDA.n1250 GNDA.n1211 3.4105
R8904 GNDA.n1250 GNDA.n1232 3.4105
R8905 GNDA.n1250 GNDA.n1210 3.4105
R8906 GNDA.n1250 GNDA.n1233 3.4105
R8907 GNDA.n1250 GNDA.n1209 3.4105
R8908 GNDA.n1250 GNDA.n1234 3.4105
R8909 GNDA.n1250 GNDA.n1208 3.4105
R8910 GNDA.n1250 GNDA.n1235 3.4105
R8911 GNDA.n1250 GNDA.n1207 3.4105
R8912 GNDA.n1250 GNDA.n1236 3.4105
R8913 GNDA.n1250 GNDA.n1206 3.4105
R8914 GNDA.n1250 GNDA.n1237 3.4105
R8915 GNDA.n2583 GNDA.n1250 3.4105
R8916 GNDA.n1320 GNDA.n1297 3.4105
R8917 GNDA.n1297 GNDA.n1222 3.4105
R8918 GNDA.n1297 GNDA.n1220 3.4105
R8919 GNDA.n1297 GNDA.n1223 3.4105
R8920 GNDA.n1297 GNDA.n1219 3.4105
R8921 GNDA.n1297 GNDA.n1224 3.4105
R8922 GNDA.n1297 GNDA.n1218 3.4105
R8923 GNDA.n1297 GNDA.n1225 3.4105
R8924 GNDA.n1297 GNDA.n1217 3.4105
R8925 GNDA.n1297 GNDA.n1226 3.4105
R8926 GNDA.n1297 GNDA.n1216 3.4105
R8927 GNDA.n1297 GNDA.n1227 3.4105
R8928 GNDA.n1297 GNDA.n1215 3.4105
R8929 GNDA.n1297 GNDA.n1228 3.4105
R8930 GNDA.n1297 GNDA.n1214 3.4105
R8931 GNDA.n1297 GNDA.n1229 3.4105
R8932 GNDA.n1297 GNDA.n1213 3.4105
R8933 GNDA.n1297 GNDA.n1230 3.4105
R8934 GNDA.n1297 GNDA.n1212 3.4105
R8935 GNDA.n1297 GNDA.n1231 3.4105
R8936 GNDA.n1297 GNDA.n1211 3.4105
R8937 GNDA.n1297 GNDA.n1232 3.4105
R8938 GNDA.n1297 GNDA.n1210 3.4105
R8939 GNDA.n1297 GNDA.n1233 3.4105
R8940 GNDA.n1297 GNDA.n1209 3.4105
R8941 GNDA.n1297 GNDA.n1234 3.4105
R8942 GNDA.n1297 GNDA.n1208 3.4105
R8943 GNDA.n1297 GNDA.n1235 3.4105
R8944 GNDA.n1297 GNDA.n1207 3.4105
R8945 GNDA.n1297 GNDA.n1236 3.4105
R8946 GNDA.n1297 GNDA.n1206 3.4105
R8947 GNDA.n1297 GNDA.n1237 3.4105
R8948 GNDA.n2583 GNDA.n1297 3.4105
R8949 GNDA.n1320 GNDA.n1249 3.4105
R8950 GNDA.n1249 GNDA.n1222 3.4105
R8951 GNDA.n1249 GNDA.n1220 3.4105
R8952 GNDA.n1249 GNDA.n1223 3.4105
R8953 GNDA.n1249 GNDA.n1219 3.4105
R8954 GNDA.n1249 GNDA.n1224 3.4105
R8955 GNDA.n1249 GNDA.n1218 3.4105
R8956 GNDA.n1249 GNDA.n1225 3.4105
R8957 GNDA.n1249 GNDA.n1217 3.4105
R8958 GNDA.n1249 GNDA.n1226 3.4105
R8959 GNDA.n1249 GNDA.n1216 3.4105
R8960 GNDA.n1249 GNDA.n1227 3.4105
R8961 GNDA.n1249 GNDA.n1215 3.4105
R8962 GNDA.n1249 GNDA.n1228 3.4105
R8963 GNDA.n1249 GNDA.n1214 3.4105
R8964 GNDA.n1249 GNDA.n1229 3.4105
R8965 GNDA.n1249 GNDA.n1213 3.4105
R8966 GNDA.n1249 GNDA.n1230 3.4105
R8967 GNDA.n1249 GNDA.n1212 3.4105
R8968 GNDA.n1249 GNDA.n1231 3.4105
R8969 GNDA.n1249 GNDA.n1211 3.4105
R8970 GNDA.n1249 GNDA.n1232 3.4105
R8971 GNDA.n1249 GNDA.n1210 3.4105
R8972 GNDA.n1249 GNDA.n1233 3.4105
R8973 GNDA.n1249 GNDA.n1209 3.4105
R8974 GNDA.n1249 GNDA.n1234 3.4105
R8975 GNDA.n1249 GNDA.n1208 3.4105
R8976 GNDA.n1249 GNDA.n1235 3.4105
R8977 GNDA.n1249 GNDA.n1207 3.4105
R8978 GNDA.n1249 GNDA.n1236 3.4105
R8979 GNDA.n1249 GNDA.n1206 3.4105
R8980 GNDA.n1249 GNDA.n1237 3.4105
R8981 GNDA.n2583 GNDA.n1249 3.4105
R8982 GNDA.n1320 GNDA.n1299 3.4105
R8983 GNDA.n1299 GNDA.n1222 3.4105
R8984 GNDA.n1299 GNDA.n1220 3.4105
R8985 GNDA.n1299 GNDA.n1223 3.4105
R8986 GNDA.n1299 GNDA.n1219 3.4105
R8987 GNDA.n1299 GNDA.n1224 3.4105
R8988 GNDA.n1299 GNDA.n1218 3.4105
R8989 GNDA.n1299 GNDA.n1225 3.4105
R8990 GNDA.n1299 GNDA.n1217 3.4105
R8991 GNDA.n1299 GNDA.n1226 3.4105
R8992 GNDA.n1299 GNDA.n1216 3.4105
R8993 GNDA.n1299 GNDA.n1227 3.4105
R8994 GNDA.n1299 GNDA.n1215 3.4105
R8995 GNDA.n1299 GNDA.n1228 3.4105
R8996 GNDA.n1299 GNDA.n1214 3.4105
R8997 GNDA.n1299 GNDA.n1229 3.4105
R8998 GNDA.n1299 GNDA.n1213 3.4105
R8999 GNDA.n1299 GNDA.n1230 3.4105
R9000 GNDA.n1299 GNDA.n1212 3.4105
R9001 GNDA.n1299 GNDA.n1231 3.4105
R9002 GNDA.n1299 GNDA.n1211 3.4105
R9003 GNDA.n1299 GNDA.n1232 3.4105
R9004 GNDA.n1299 GNDA.n1210 3.4105
R9005 GNDA.n1299 GNDA.n1233 3.4105
R9006 GNDA.n1299 GNDA.n1209 3.4105
R9007 GNDA.n1299 GNDA.n1234 3.4105
R9008 GNDA.n1299 GNDA.n1208 3.4105
R9009 GNDA.n1299 GNDA.n1235 3.4105
R9010 GNDA.n1299 GNDA.n1207 3.4105
R9011 GNDA.n1299 GNDA.n1236 3.4105
R9012 GNDA.n1299 GNDA.n1206 3.4105
R9013 GNDA.n1299 GNDA.n1237 3.4105
R9014 GNDA.n2583 GNDA.n1299 3.4105
R9015 GNDA.n1320 GNDA.n1248 3.4105
R9016 GNDA.n1248 GNDA.n1222 3.4105
R9017 GNDA.n1248 GNDA.n1220 3.4105
R9018 GNDA.n1248 GNDA.n1223 3.4105
R9019 GNDA.n1248 GNDA.n1219 3.4105
R9020 GNDA.n1248 GNDA.n1224 3.4105
R9021 GNDA.n1248 GNDA.n1218 3.4105
R9022 GNDA.n1248 GNDA.n1225 3.4105
R9023 GNDA.n1248 GNDA.n1217 3.4105
R9024 GNDA.n1248 GNDA.n1226 3.4105
R9025 GNDA.n1248 GNDA.n1216 3.4105
R9026 GNDA.n1248 GNDA.n1227 3.4105
R9027 GNDA.n1248 GNDA.n1215 3.4105
R9028 GNDA.n1248 GNDA.n1228 3.4105
R9029 GNDA.n1248 GNDA.n1214 3.4105
R9030 GNDA.n1248 GNDA.n1229 3.4105
R9031 GNDA.n1248 GNDA.n1213 3.4105
R9032 GNDA.n1248 GNDA.n1230 3.4105
R9033 GNDA.n1248 GNDA.n1212 3.4105
R9034 GNDA.n1248 GNDA.n1231 3.4105
R9035 GNDA.n1248 GNDA.n1211 3.4105
R9036 GNDA.n1248 GNDA.n1232 3.4105
R9037 GNDA.n1248 GNDA.n1210 3.4105
R9038 GNDA.n1248 GNDA.n1233 3.4105
R9039 GNDA.n1248 GNDA.n1209 3.4105
R9040 GNDA.n1248 GNDA.n1234 3.4105
R9041 GNDA.n1248 GNDA.n1208 3.4105
R9042 GNDA.n1248 GNDA.n1235 3.4105
R9043 GNDA.n1248 GNDA.n1207 3.4105
R9044 GNDA.n1248 GNDA.n1236 3.4105
R9045 GNDA.n1248 GNDA.n1206 3.4105
R9046 GNDA.n1248 GNDA.n1237 3.4105
R9047 GNDA.n2583 GNDA.n1248 3.4105
R9048 GNDA.n1320 GNDA.n1301 3.4105
R9049 GNDA.n1301 GNDA.n1222 3.4105
R9050 GNDA.n1301 GNDA.n1220 3.4105
R9051 GNDA.n1301 GNDA.n1223 3.4105
R9052 GNDA.n1301 GNDA.n1219 3.4105
R9053 GNDA.n1301 GNDA.n1224 3.4105
R9054 GNDA.n1301 GNDA.n1218 3.4105
R9055 GNDA.n1301 GNDA.n1225 3.4105
R9056 GNDA.n1301 GNDA.n1217 3.4105
R9057 GNDA.n1301 GNDA.n1226 3.4105
R9058 GNDA.n1301 GNDA.n1216 3.4105
R9059 GNDA.n1301 GNDA.n1227 3.4105
R9060 GNDA.n1301 GNDA.n1215 3.4105
R9061 GNDA.n1301 GNDA.n1228 3.4105
R9062 GNDA.n1301 GNDA.n1214 3.4105
R9063 GNDA.n1301 GNDA.n1229 3.4105
R9064 GNDA.n1301 GNDA.n1213 3.4105
R9065 GNDA.n1301 GNDA.n1230 3.4105
R9066 GNDA.n1301 GNDA.n1212 3.4105
R9067 GNDA.n1301 GNDA.n1231 3.4105
R9068 GNDA.n1301 GNDA.n1211 3.4105
R9069 GNDA.n1301 GNDA.n1232 3.4105
R9070 GNDA.n1301 GNDA.n1210 3.4105
R9071 GNDA.n1301 GNDA.n1233 3.4105
R9072 GNDA.n1301 GNDA.n1209 3.4105
R9073 GNDA.n1301 GNDA.n1234 3.4105
R9074 GNDA.n1301 GNDA.n1208 3.4105
R9075 GNDA.n1301 GNDA.n1235 3.4105
R9076 GNDA.n1301 GNDA.n1207 3.4105
R9077 GNDA.n1301 GNDA.n1236 3.4105
R9078 GNDA.n1301 GNDA.n1206 3.4105
R9079 GNDA.n1301 GNDA.n1237 3.4105
R9080 GNDA.n2583 GNDA.n1301 3.4105
R9081 GNDA.n1320 GNDA.n1247 3.4105
R9082 GNDA.n1247 GNDA.n1222 3.4105
R9083 GNDA.n1247 GNDA.n1220 3.4105
R9084 GNDA.n1247 GNDA.n1223 3.4105
R9085 GNDA.n1247 GNDA.n1219 3.4105
R9086 GNDA.n1247 GNDA.n1224 3.4105
R9087 GNDA.n1247 GNDA.n1218 3.4105
R9088 GNDA.n1247 GNDA.n1225 3.4105
R9089 GNDA.n1247 GNDA.n1217 3.4105
R9090 GNDA.n1247 GNDA.n1226 3.4105
R9091 GNDA.n1247 GNDA.n1216 3.4105
R9092 GNDA.n1247 GNDA.n1227 3.4105
R9093 GNDA.n1247 GNDA.n1215 3.4105
R9094 GNDA.n1247 GNDA.n1228 3.4105
R9095 GNDA.n1247 GNDA.n1214 3.4105
R9096 GNDA.n1247 GNDA.n1229 3.4105
R9097 GNDA.n1247 GNDA.n1213 3.4105
R9098 GNDA.n1247 GNDA.n1230 3.4105
R9099 GNDA.n1247 GNDA.n1212 3.4105
R9100 GNDA.n1247 GNDA.n1231 3.4105
R9101 GNDA.n1247 GNDA.n1211 3.4105
R9102 GNDA.n1247 GNDA.n1232 3.4105
R9103 GNDA.n1247 GNDA.n1210 3.4105
R9104 GNDA.n1247 GNDA.n1233 3.4105
R9105 GNDA.n1247 GNDA.n1209 3.4105
R9106 GNDA.n1247 GNDA.n1234 3.4105
R9107 GNDA.n1247 GNDA.n1208 3.4105
R9108 GNDA.n1247 GNDA.n1235 3.4105
R9109 GNDA.n1247 GNDA.n1207 3.4105
R9110 GNDA.n1247 GNDA.n1236 3.4105
R9111 GNDA.n1247 GNDA.n1206 3.4105
R9112 GNDA.n1247 GNDA.n1237 3.4105
R9113 GNDA.n2583 GNDA.n1247 3.4105
R9114 GNDA.n1320 GNDA.n1303 3.4105
R9115 GNDA.n1303 GNDA.n1222 3.4105
R9116 GNDA.n1303 GNDA.n1220 3.4105
R9117 GNDA.n1303 GNDA.n1223 3.4105
R9118 GNDA.n1303 GNDA.n1219 3.4105
R9119 GNDA.n1303 GNDA.n1224 3.4105
R9120 GNDA.n1303 GNDA.n1218 3.4105
R9121 GNDA.n1303 GNDA.n1225 3.4105
R9122 GNDA.n1303 GNDA.n1217 3.4105
R9123 GNDA.n1303 GNDA.n1226 3.4105
R9124 GNDA.n1303 GNDA.n1216 3.4105
R9125 GNDA.n1303 GNDA.n1227 3.4105
R9126 GNDA.n1303 GNDA.n1215 3.4105
R9127 GNDA.n1303 GNDA.n1228 3.4105
R9128 GNDA.n1303 GNDA.n1214 3.4105
R9129 GNDA.n1303 GNDA.n1229 3.4105
R9130 GNDA.n1303 GNDA.n1213 3.4105
R9131 GNDA.n1303 GNDA.n1230 3.4105
R9132 GNDA.n1303 GNDA.n1212 3.4105
R9133 GNDA.n1303 GNDA.n1231 3.4105
R9134 GNDA.n1303 GNDA.n1211 3.4105
R9135 GNDA.n1303 GNDA.n1232 3.4105
R9136 GNDA.n1303 GNDA.n1210 3.4105
R9137 GNDA.n1303 GNDA.n1233 3.4105
R9138 GNDA.n1303 GNDA.n1209 3.4105
R9139 GNDA.n1303 GNDA.n1234 3.4105
R9140 GNDA.n1303 GNDA.n1208 3.4105
R9141 GNDA.n1303 GNDA.n1235 3.4105
R9142 GNDA.n1303 GNDA.n1207 3.4105
R9143 GNDA.n1303 GNDA.n1236 3.4105
R9144 GNDA.n1303 GNDA.n1206 3.4105
R9145 GNDA.n1303 GNDA.n1237 3.4105
R9146 GNDA.n2583 GNDA.n1303 3.4105
R9147 GNDA.n1320 GNDA.n1246 3.4105
R9148 GNDA.n1246 GNDA.n1222 3.4105
R9149 GNDA.n1246 GNDA.n1220 3.4105
R9150 GNDA.n1246 GNDA.n1223 3.4105
R9151 GNDA.n1246 GNDA.n1219 3.4105
R9152 GNDA.n1246 GNDA.n1224 3.4105
R9153 GNDA.n1246 GNDA.n1218 3.4105
R9154 GNDA.n1246 GNDA.n1225 3.4105
R9155 GNDA.n1246 GNDA.n1217 3.4105
R9156 GNDA.n1246 GNDA.n1226 3.4105
R9157 GNDA.n1246 GNDA.n1216 3.4105
R9158 GNDA.n1246 GNDA.n1227 3.4105
R9159 GNDA.n1246 GNDA.n1215 3.4105
R9160 GNDA.n1246 GNDA.n1228 3.4105
R9161 GNDA.n1246 GNDA.n1214 3.4105
R9162 GNDA.n1246 GNDA.n1229 3.4105
R9163 GNDA.n1246 GNDA.n1213 3.4105
R9164 GNDA.n1246 GNDA.n1230 3.4105
R9165 GNDA.n1246 GNDA.n1212 3.4105
R9166 GNDA.n1246 GNDA.n1231 3.4105
R9167 GNDA.n1246 GNDA.n1211 3.4105
R9168 GNDA.n1246 GNDA.n1232 3.4105
R9169 GNDA.n1246 GNDA.n1210 3.4105
R9170 GNDA.n1246 GNDA.n1233 3.4105
R9171 GNDA.n1246 GNDA.n1209 3.4105
R9172 GNDA.n1246 GNDA.n1234 3.4105
R9173 GNDA.n1246 GNDA.n1208 3.4105
R9174 GNDA.n1246 GNDA.n1235 3.4105
R9175 GNDA.n1246 GNDA.n1207 3.4105
R9176 GNDA.n1246 GNDA.n1236 3.4105
R9177 GNDA.n1246 GNDA.n1206 3.4105
R9178 GNDA.n1246 GNDA.n1237 3.4105
R9179 GNDA.n2583 GNDA.n1246 3.4105
R9180 GNDA.n1320 GNDA.n1305 3.4105
R9181 GNDA.n1305 GNDA.n1222 3.4105
R9182 GNDA.n1305 GNDA.n1220 3.4105
R9183 GNDA.n1305 GNDA.n1223 3.4105
R9184 GNDA.n1305 GNDA.n1219 3.4105
R9185 GNDA.n1305 GNDA.n1224 3.4105
R9186 GNDA.n1305 GNDA.n1218 3.4105
R9187 GNDA.n1305 GNDA.n1225 3.4105
R9188 GNDA.n1305 GNDA.n1217 3.4105
R9189 GNDA.n1305 GNDA.n1226 3.4105
R9190 GNDA.n1305 GNDA.n1216 3.4105
R9191 GNDA.n1305 GNDA.n1227 3.4105
R9192 GNDA.n1305 GNDA.n1215 3.4105
R9193 GNDA.n1305 GNDA.n1228 3.4105
R9194 GNDA.n1305 GNDA.n1214 3.4105
R9195 GNDA.n1305 GNDA.n1229 3.4105
R9196 GNDA.n1305 GNDA.n1213 3.4105
R9197 GNDA.n1305 GNDA.n1230 3.4105
R9198 GNDA.n1305 GNDA.n1212 3.4105
R9199 GNDA.n1305 GNDA.n1231 3.4105
R9200 GNDA.n1305 GNDA.n1211 3.4105
R9201 GNDA.n1305 GNDA.n1232 3.4105
R9202 GNDA.n1305 GNDA.n1210 3.4105
R9203 GNDA.n1305 GNDA.n1233 3.4105
R9204 GNDA.n1305 GNDA.n1209 3.4105
R9205 GNDA.n1305 GNDA.n1234 3.4105
R9206 GNDA.n1305 GNDA.n1208 3.4105
R9207 GNDA.n1305 GNDA.n1235 3.4105
R9208 GNDA.n1305 GNDA.n1207 3.4105
R9209 GNDA.n1305 GNDA.n1236 3.4105
R9210 GNDA.n1305 GNDA.n1206 3.4105
R9211 GNDA.n1305 GNDA.n1237 3.4105
R9212 GNDA.n2583 GNDA.n1305 3.4105
R9213 GNDA.n1320 GNDA.n1245 3.4105
R9214 GNDA.n1245 GNDA.n1222 3.4105
R9215 GNDA.n1245 GNDA.n1220 3.4105
R9216 GNDA.n1245 GNDA.n1223 3.4105
R9217 GNDA.n1245 GNDA.n1219 3.4105
R9218 GNDA.n1245 GNDA.n1224 3.4105
R9219 GNDA.n1245 GNDA.n1218 3.4105
R9220 GNDA.n1245 GNDA.n1225 3.4105
R9221 GNDA.n1245 GNDA.n1217 3.4105
R9222 GNDA.n1245 GNDA.n1226 3.4105
R9223 GNDA.n1245 GNDA.n1216 3.4105
R9224 GNDA.n1245 GNDA.n1227 3.4105
R9225 GNDA.n1245 GNDA.n1215 3.4105
R9226 GNDA.n1245 GNDA.n1228 3.4105
R9227 GNDA.n1245 GNDA.n1214 3.4105
R9228 GNDA.n1245 GNDA.n1229 3.4105
R9229 GNDA.n1245 GNDA.n1213 3.4105
R9230 GNDA.n1245 GNDA.n1230 3.4105
R9231 GNDA.n1245 GNDA.n1212 3.4105
R9232 GNDA.n1245 GNDA.n1231 3.4105
R9233 GNDA.n1245 GNDA.n1211 3.4105
R9234 GNDA.n1245 GNDA.n1232 3.4105
R9235 GNDA.n1245 GNDA.n1210 3.4105
R9236 GNDA.n1245 GNDA.n1233 3.4105
R9237 GNDA.n1245 GNDA.n1209 3.4105
R9238 GNDA.n1245 GNDA.n1234 3.4105
R9239 GNDA.n1245 GNDA.n1208 3.4105
R9240 GNDA.n1245 GNDA.n1235 3.4105
R9241 GNDA.n1245 GNDA.n1207 3.4105
R9242 GNDA.n1245 GNDA.n1236 3.4105
R9243 GNDA.n1245 GNDA.n1206 3.4105
R9244 GNDA.n1245 GNDA.n1237 3.4105
R9245 GNDA.n2583 GNDA.n1245 3.4105
R9246 GNDA.n1320 GNDA.n1307 3.4105
R9247 GNDA.n1307 GNDA.n1222 3.4105
R9248 GNDA.n1307 GNDA.n1220 3.4105
R9249 GNDA.n1307 GNDA.n1223 3.4105
R9250 GNDA.n1307 GNDA.n1219 3.4105
R9251 GNDA.n1307 GNDA.n1224 3.4105
R9252 GNDA.n1307 GNDA.n1218 3.4105
R9253 GNDA.n1307 GNDA.n1225 3.4105
R9254 GNDA.n1307 GNDA.n1217 3.4105
R9255 GNDA.n1307 GNDA.n1226 3.4105
R9256 GNDA.n1307 GNDA.n1216 3.4105
R9257 GNDA.n1307 GNDA.n1227 3.4105
R9258 GNDA.n1307 GNDA.n1215 3.4105
R9259 GNDA.n1307 GNDA.n1228 3.4105
R9260 GNDA.n1307 GNDA.n1214 3.4105
R9261 GNDA.n1307 GNDA.n1229 3.4105
R9262 GNDA.n1307 GNDA.n1213 3.4105
R9263 GNDA.n1307 GNDA.n1230 3.4105
R9264 GNDA.n1307 GNDA.n1212 3.4105
R9265 GNDA.n1307 GNDA.n1231 3.4105
R9266 GNDA.n1307 GNDA.n1211 3.4105
R9267 GNDA.n1307 GNDA.n1232 3.4105
R9268 GNDA.n1307 GNDA.n1210 3.4105
R9269 GNDA.n1307 GNDA.n1233 3.4105
R9270 GNDA.n1307 GNDA.n1209 3.4105
R9271 GNDA.n1307 GNDA.n1234 3.4105
R9272 GNDA.n1307 GNDA.n1208 3.4105
R9273 GNDA.n1307 GNDA.n1235 3.4105
R9274 GNDA.n1307 GNDA.n1207 3.4105
R9275 GNDA.n1307 GNDA.n1236 3.4105
R9276 GNDA.n1307 GNDA.n1206 3.4105
R9277 GNDA.n1307 GNDA.n1237 3.4105
R9278 GNDA.n2583 GNDA.n1307 3.4105
R9279 GNDA.n1320 GNDA.n1244 3.4105
R9280 GNDA.n1244 GNDA.n1222 3.4105
R9281 GNDA.n1244 GNDA.n1220 3.4105
R9282 GNDA.n1244 GNDA.n1223 3.4105
R9283 GNDA.n1244 GNDA.n1219 3.4105
R9284 GNDA.n1244 GNDA.n1224 3.4105
R9285 GNDA.n1244 GNDA.n1218 3.4105
R9286 GNDA.n1244 GNDA.n1225 3.4105
R9287 GNDA.n1244 GNDA.n1217 3.4105
R9288 GNDA.n1244 GNDA.n1226 3.4105
R9289 GNDA.n1244 GNDA.n1216 3.4105
R9290 GNDA.n1244 GNDA.n1227 3.4105
R9291 GNDA.n1244 GNDA.n1215 3.4105
R9292 GNDA.n1244 GNDA.n1228 3.4105
R9293 GNDA.n1244 GNDA.n1214 3.4105
R9294 GNDA.n1244 GNDA.n1229 3.4105
R9295 GNDA.n1244 GNDA.n1213 3.4105
R9296 GNDA.n1244 GNDA.n1230 3.4105
R9297 GNDA.n1244 GNDA.n1212 3.4105
R9298 GNDA.n1244 GNDA.n1231 3.4105
R9299 GNDA.n1244 GNDA.n1211 3.4105
R9300 GNDA.n1244 GNDA.n1232 3.4105
R9301 GNDA.n1244 GNDA.n1210 3.4105
R9302 GNDA.n1244 GNDA.n1233 3.4105
R9303 GNDA.n1244 GNDA.n1209 3.4105
R9304 GNDA.n1244 GNDA.n1234 3.4105
R9305 GNDA.n1244 GNDA.n1208 3.4105
R9306 GNDA.n1244 GNDA.n1235 3.4105
R9307 GNDA.n1244 GNDA.n1207 3.4105
R9308 GNDA.n1244 GNDA.n1236 3.4105
R9309 GNDA.n1244 GNDA.n1206 3.4105
R9310 GNDA.n1244 GNDA.n1237 3.4105
R9311 GNDA.n2583 GNDA.n1244 3.4105
R9312 GNDA.n1320 GNDA.n1309 3.4105
R9313 GNDA.n1309 GNDA.n1222 3.4105
R9314 GNDA.n1309 GNDA.n1220 3.4105
R9315 GNDA.n1309 GNDA.n1223 3.4105
R9316 GNDA.n1309 GNDA.n1219 3.4105
R9317 GNDA.n1309 GNDA.n1224 3.4105
R9318 GNDA.n1309 GNDA.n1218 3.4105
R9319 GNDA.n1309 GNDA.n1225 3.4105
R9320 GNDA.n1309 GNDA.n1217 3.4105
R9321 GNDA.n1309 GNDA.n1226 3.4105
R9322 GNDA.n1309 GNDA.n1216 3.4105
R9323 GNDA.n1309 GNDA.n1227 3.4105
R9324 GNDA.n1309 GNDA.n1215 3.4105
R9325 GNDA.n1309 GNDA.n1228 3.4105
R9326 GNDA.n1309 GNDA.n1214 3.4105
R9327 GNDA.n1309 GNDA.n1229 3.4105
R9328 GNDA.n1309 GNDA.n1213 3.4105
R9329 GNDA.n1309 GNDA.n1230 3.4105
R9330 GNDA.n1309 GNDA.n1212 3.4105
R9331 GNDA.n1309 GNDA.n1231 3.4105
R9332 GNDA.n1309 GNDA.n1211 3.4105
R9333 GNDA.n1309 GNDA.n1232 3.4105
R9334 GNDA.n1309 GNDA.n1210 3.4105
R9335 GNDA.n1309 GNDA.n1233 3.4105
R9336 GNDA.n1309 GNDA.n1209 3.4105
R9337 GNDA.n1309 GNDA.n1234 3.4105
R9338 GNDA.n1309 GNDA.n1208 3.4105
R9339 GNDA.n1309 GNDA.n1235 3.4105
R9340 GNDA.n1309 GNDA.n1207 3.4105
R9341 GNDA.n1309 GNDA.n1236 3.4105
R9342 GNDA.n1309 GNDA.n1206 3.4105
R9343 GNDA.n1309 GNDA.n1237 3.4105
R9344 GNDA.n2583 GNDA.n1309 3.4105
R9345 GNDA.n1320 GNDA.n1243 3.4105
R9346 GNDA.n1243 GNDA.n1222 3.4105
R9347 GNDA.n1243 GNDA.n1220 3.4105
R9348 GNDA.n1243 GNDA.n1223 3.4105
R9349 GNDA.n1243 GNDA.n1219 3.4105
R9350 GNDA.n1243 GNDA.n1224 3.4105
R9351 GNDA.n1243 GNDA.n1218 3.4105
R9352 GNDA.n1243 GNDA.n1225 3.4105
R9353 GNDA.n1243 GNDA.n1217 3.4105
R9354 GNDA.n1243 GNDA.n1226 3.4105
R9355 GNDA.n1243 GNDA.n1216 3.4105
R9356 GNDA.n1243 GNDA.n1227 3.4105
R9357 GNDA.n1243 GNDA.n1215 3.4105
R9358 GNDA.n1243 GNDA.n1228 3.4105
R9359 GNDA.n1243 GNDA.n1214 3.4105
R9360 GNDA.n1243 GNDA.n1229 3.4105
R9361 GNDA.n1243 GNDA.n1213 3.4105
R9362 GNDA.n1243 GNDA.n1230 3.4105
R9363 GNDA.n1243 GNDA.n1212 3.4105
R9364 GNDA.n1243 GNDA.n1231 3.4105
R9365 GNDA.n1243 GNDA.n1211 3.4105
R9366 GNDA.n1243 GNDA.n1232 3.4105
R9367 GNDA.n1243 GNDA.n1210 3.4105
R9368 GNDA.n1243 GNDA.n1233 3.4105
R9369 GNDA.n1243 GNDA.n1209 3.4105
R9370 GNDA.n1243 GNDA.n1234 3.4105
R9371 GNDA.n1243 GNDA.n1208 3.4105
R9372 GNDA.n1243 GNDA.n1235 3.4105
R9373 GNDA.n1243 GNDA.n1207 3.4105
R9374 GNDA.n1243 GNDA.n1236 3.4105
R9375 GNDA.n1243 GNDA.n1206 3.4105
R9376 GNDA.n1243 GNDA.n1237 3.4105
R9377 GNDA.n2583 GNDA.n1243 3.4105
R9378 GNDA.n1320 GNDA.n1311 3.4105
R9379 GNDA.n1311 GNDA.n1222 3.4105
R9380 GNDA.n1311 GNDA.n1220 3.4105
R9381 GNDA.n1311 GNDA.n1223 3.4105
R9382 GNDA.n1311 GNDA.n1219 3.4105
R9383 GNDA.n1311 GNDA.n1224 3.4105
R9384 GNDA.n1311 GNDA.n1218 3.4105
R9385 GNDA.n1311 GNDA.n1225 3.4105
R9386 GNDA.n1311 GNDA.n1217 3.4105
R9387 GNDA.n1311 GNDA.n1226 3.4105
R9388 GNDA.n1311 GNDA.n1216 3.4105
R9389 GNDA.n1311 GNDA.n1227 3.4105
R9390 GNDA.n1311 GNDA.n1215 3.4105
R9391 GNDA.n1311 GNDA.n1228 3.4105
R9392 GNDA.n1311 GNDA.n1214 3.4105
R9393 GNDA.n1311 GNDA.n1229 3.4105
R9394 GNDA.n1311 GNDA.n1213 3.4105
R9395 GNDA.n1311 GNDA.n1230 3.4105
R9396 GNDA.n1311 GNDA.n1212 3.4105
R9397 GNDA.n1311 GNDA.n1231 3.4105
R9398 GNDA.n1311 GNDA.n1211 3.4105
R9399 GNDA.n1311 GNDA.n1232 3.4105
R9400 GNDA.n1311 GNDA.n1210 3.4105
R9401 GNDA.n1311 GNDA.n1233 3.4105
R9402 GNDA.n1311 GNDA.n1209 3.4105
R9403 GNDA.n1311 GNDA.n1234 3.4105
R9404 GNDA.n1311 GNDA.n1208 3.4105
R9405 GNDA.n1311 GNDA.n1235 3.4105
R9406 GNDA.n1311 GNDA.n1207 3.4105
R9407 GNDA.n1311 GNDA.n1236 3.4105
R9408 GNDA.n1311 GNDA.n1206 3.4105
R9409 GNDA.n1311 GNDA.n1237 3.4105
R9410 GNDA.n2583 GNDA.n1311 3.4105
R9411 GNDA.n1320 GNDA.n1242 3.4105
R9412 GNDA.n1242 GNDA.n1222 3.4105
R9413 GNDA.n1242 GNDA.n1220 3.4105
R9414 GNDA.n1242 GNDA.n1223 3.4105
R9415 GNDA.n1242 GNDA.n1219 3.4105
R9416 GNDA.n1242 GNDA.n1224 3.4105
R9417 GNDA.n1242 GNDA.n1218 3.4105
R9418 GNDA.n1242 GNDA.n1225 3.4105
R9419 GNDA.n1242 GNDA.n1217 3.4105
R9420 GNDA.n1242 GNDA.n1226 3.4105
R9421 GNDA.n1242 GNDA.n1216 3.4105
R9422 GNDA.n1242 GNDA.n1227 3.4105
R9423 GNDA.n1242 GNDA.n1215 3.4105
R9424 GNDA.n1242 GNDA.n1228 3.4105
R9425 GNDA.n1242 GNDA.n1214 3.4105
R9426 GNDA.n1242 GNDA.n1229 3.4105
R9427 GNDA.n1242 GNDA.n1213 3.4105
R9428 GNDA.n1242 GNDA.n1230 3.4105
R9429 GNDA.n1242 GNDA.n1212 3.4105
R9430 GNDA.n1242 GNDA.n1231 3.4105
R9431 GNDA.n1242 GNDA.n1211 3.4105
R9432 GNDA.n1242 GNDA.n1232 3.4105
R9433 GNDA.n1242 GNDA.n1210 3.4105
R9434 GNDA.n1242 GNDA.n1233 3.4105
R9435 GNDA.n1242 GNDA.n1209 3.4105
R9436 GNDA.n1242 GNDA.n1234 3.4105
R9437 GNDA.n1242 GNDA.n1208 3.4105
R9438 GNDA.n1242 GNDA.n1235 3.4105
R9439 GNDA.n1242 GNDA.n1207 3.4105
R9440 GNDA.n1242 GNDA.n1236 3.4105
R9441 GNDA.n1242 GNDA.n1206 3.4105
R9442 GNDA.n1242 GNDA.n1237 3.4105
R9443 GNDA.n2583 GNDA.n1242 3.4105
R9444 GNDA.n1320 GNDA.n1313 3.4105
R9445 GNDA.n1313 GNDA.n1222 3.4105
R9446 GNDA.n1313 GNDA.n1220 3.4105
R9447 GNDA.n1313 GNDA.n1223 3.4105
R9448 GNDA.n1313 GNDA.n1219 3.4105
R9449 GNDA.n1313 GNDA.n1224 3.4105
R9450 GNDA.n1313 GNDA.n1218 3.4105
R9451 GNDA.n1313 GNDA.n1225 3.4105
R9452 GNDA.n1313 GNDA.n1217 3.4105
R9453 GNDA.n1313 GNDA.n1226 3.4105
R9454 GNDA.n1313 GNDA.n1216 3.4105
R9455 GNDA.n1313 GNDA.n1227 3.4105
R9456 GNDA.n1313 GNDA.n1215 3.4105
R9457 GNDA.n1313 GNDA.n1228 3.4105
R9458 GNDA.n1313 GNDA.n1214 3.4105
R9459 GNDA.n1313 GNDA.n1229 3.4105
R9460 GNDA.n1313 GNDA.n1213 3.4105
R9461 GNDA.n1313 GNDA.n1230 3.4105
R9462 GNDA.n1313 GNDA.n1212 3.4105
R9463 GNDA.n1313 GNDA.n1231 3.4105
R9464 GNDA.n1313 GNDA.n1211 3.4105
R9465 GNDA.n1313 GNDA.n1232 3.4105
R9466 GNDA.n1313 GNDA.n1210 3.4105
R9467 GNDA.n1313 GNDA.n1233 3.4105
R9468 GNDA.n1313 GNDA.n1209 3.4105
R9469 GNDA.n1313 GNDA.n1234 3.4105
R9470 GNDA.n1313 GNDA.n1208 3.4105
R9471 GNDA.n1313 GNDA.n1235 3.4105
R9472 GNDA.n1313 GNDA.n1207 3.4105
R9473 GNDA.n1313 GNDA.n1236 3.4105
R9474 GNDA.n1313 GNDA.n1206 3.4105
R9475 GNDA.n1313 GNDA.n1237 3.4105
R9476 GNDA.n2583 GNDA.n1313 3.4105
R9477 GNDA.n1320 GNDA.n1241 3.4105
R9478 GNDA.n1241 GNDA.n1222 3.4105
R9479 GNDA.n1241 GNDA.n1220 3.4105
R9480 GNDA.n1241 GNDA.n1223 3.4105
R9481 GNDA.n1241 GNDA.n1219 3.4105
R9482 GNDA.n1241 GNDA.n1224 3.4105
R9483 GNDA.n1241 GNDA.n1218 3.4105
R9484 GNDA.n1241 GNDA.n1225 3.4105
R9485 GNDA.n1241 GNDA.n1217 3.4105
R9486 GNDA.n1241 GNDA.n1226 3.4105
R9487 GNDA.n1241 GNDA.n1216 3.4105
R9488 GNDA.n1241 GNDA.n1227 3.4105
R9489 GNDA.n1241 GNDA.n1215 3.4105
R9490 GNDA.n1241 GNDA.n1228 3.4105
R9491 GNDA.n1241 GNDA.n1214 3.4105
R9492 GNDA.n1241 GNDA.n1229 3.4105
R9493 GNDA.n1241 GNDA.n1213 3.4105
R9494 GNDA.n1241 GNDA.n1230 3.4105
R9495 GNDA.n1241 GNDA.n1212 3.4105
R9496 GNDA.n1241 GNDA.n1231 3.4105
R9497 GNDA.n1241 GNDA.n1211 3.4105
R9498 GNDA.n1241 GNDA.n1232 3.4105
R9499 GNDA.n1241 GNDA.n1210 3.4105
R9500 GNDA.n1241 GNDA.n1233 3.4105
R9501 GNDA.n1241 GNDA.n1209 3.4105
R9502 GNDA.n1241 GNDA.n1234 3.4105
R9503 GNDA.n1241 GNDA.n1208 3.4105
R9504 GNDA.n1241 GNDA.n1235 3.4105
R9505 GNDA.n1241 GNDA.n1207 3.4105
R9506 GNDA.n1241 GNDA.n1236 3.4105
R9507 GNDA.n1241 GNDA.n1206 3.4105
R9508 GNDA.n1241 GNDA.n1237 3.4105
R9509 GNDA.n2583 GNDA.n1241 3.4105
R9510 GNDA.n1320 GNDA.n1315 3.4105
R9511 GNDA.n1315 GNDA.n1222 3.4105
R9512 GNDA.n1315 GNDA.n1220 3.4105
R9513 GNDA.n1315 GNDA.n1223 3.4105
R9514 GNDA.n1315 GNDA.n1219 3.4105
R9515 GNDA.n1315 GNDA.n1224 3.4105
R9516 GNDA.n1315 GNDA.n1218 3.4105
R9517 GNDA.n1315 GNDA.n1225 3.4105
R9518 GNDA.n1315 GNDA.n1217 3.4105
R9519 GNDA.n1315 GNDA.n1226 3.4105
R9520 GNDA.n1315 GNDA.n1216 3.4105
R9521 GNDA.n1315 GNDA.n1227 3.4105
R9522 GNDA.n1315 GNDA.n1215 3.4105
R9523 GNDA.n1315 GNDA.n1228 3.4105
R9524 GNDA.n1315 GNDA.n1214 3.4105
R9525 GNDA.n1315 GNDA.n1229 3.4105
R9526 GNDA.n1315 GNDA.n1213 3.4105
R9527 GNDA.n1315 GNDA.n1230 3.4105
R9528 GNDA.n1315 GNDA.n1212 3.4105
R9529 GNDA.n1315 GNDA.n1231 3.4105
R9530 GNDA.n1315 GNDA.n1211 3.4105
R9531 GNDA.n1315 GNDA.n1232 3.4105
R9532 GNDA.n1315 GNDA.n1210 3.4105
R9533 GNDA.n1315 GNDA.n1233 3.4105
R9534 GNDA.n1315 GNDA.n1209 3.4105
R9535 GNDA.n1315 GNDA.n1234 3.4105
R9536 GNDA.n1315 GNDA.n1208 3.4105
R9537 GNDA.n1315 GNDA.n1235 3.4105
R9538 GNDA.n1315 GNDA.n1207 3.4105
R9539 GNDA.n1315 GNDA.n1236 3.4105
R9540 GNDA.n1315 GNDA.n1206 3.4105
R9541 GNDA.n1315 GNDA.n1237 3.4105
R9542 GNDA.n2583 GNDA.n1315 3.4105
R9543 GNDA.n1320 GNDA.n1240 3.4105
R9544 GNDA.n1240 GNDA.n1222 3.4105
R9545 GNDA.n1240 GNDA.n1220 3.4105
R9546 GNDA.n1240 GNDA.n1223 3.4105
R9547 GNDA.n1240 GNDA.n1219 3.4105
R9548 GNDA.n1240 GNDA.n1224 3.4105
R9549 GNDA.n1240 GNDA.n1218 3.4105
R9550 GNDA.n1240 GNDA.n1225 3.4105
R9551 GNDA.n1240 GNDA.n1217 3.4105
R9552 GNDA.n1240 GNDA.n1226 3.4105
R9553 GNDA.n1240 GNDA.n1216 3.4105
R9554 GNDA.n1240 GNDA.n1227 3.4105
R9555 GNDA.n1240 GNDA.n1215 3.4105
R9556 GNDA.n1240 GNDA.n1228 3.4105
R9557 GNDA.n1240 GNDA.n1214 3.4105
R9558 GNDA.n1240 GNDA.n1229 3.4105
R9559 GNDA.n1240 GNDA.n1213 3.4105
R9560 GNDA.n1240 GNDA.n1230 3.4105
R9561 GNDA.n1240 GNDA.n1212 3.4105
R9562 GNDA.n1240 GNDA.n1231 3.4105
R9563 GNDA.n1240 GNDA.n1211 3.4105
R9564 GNDA.n1240 GNDA.n1232 3.4105
R9565 GNDA.n1240 GNDA.n1210 3.4105
R9566 GNDA.n1240 GNDA.n1233 3.4105
R9567 GNDA.n1240 GNDA.n1209 3.4105
R9568 GNDA.n1240 GNDA.n1234 3.4105
R9569 GNDA.n1240 GNDA.n1208 3.4105
R9570 GNDA.n1240 GNDA.n1235 3.4105
R9571 GNDA.n1240 GNDA.n1207 3.4105
R9572 GNDA.n1240 GNDA.n1236 3.4105
R9573 GNDA.n1240 GNDA.n1206 3.4105
R9574 GNDA.n1240 GNDA.n1237 3.4105
R9575 GNDA.n2583 GNDA.n1240 3.4105
R9576 GNDA.n1320 GNDA.n1317 3.4105
R9577 GNDA.n1317 GNDA.n1222 3.4105
R9578 GNDA.n1317 GNDA.n1220 3.4105
R9579 GNDA.n1317 GNDA.n1223 3.4105
R9580 GNDA.n1317 GNDA.n1219 3.4105
R9581 GNDA.n1317 GNDA.n1224 3.4105
R9582 GNDA.n1317 GNDA.n1218 3.4105
R9583 GNDA.n1317 GNDA.n1225 3.4105
R9584 GNDA.n1317 GNDA.n1217 3.4105
R9585 GNDA.n1317 GNDA.n1226 3.4105
R9586 GNDA.n1317 GNDA.n1216 3.4105
R9587 GNDA.n1317 GNDA.n1227 3.4105
R9588 GNDA.n1317 GNDA.n1215 3.4105
R9589 GNDA.n1317 GNDA.n1228 3.4105
R9590 GNDA.n1317 GNDA.n1214 3.4105
R9591 GNDA.n1317 GNDA.n1229 3.4105
R9592 GNDA.n1317 GNDA.n1213 3.4105
R9593 GNDA.n1317 GNDA.n1230 3.4105
R9594 GNDA.n1317 GNDA.n1212 3.4105
R9595 GNDA.n1317 GNDA.n1231 3.4105
R9596 GNDA.n1317 GNDA.n1211 3.4105
R9597 GNDA.n1317 GNDA.n1232 3.4105
R9598 GNDA.n1317 GNDA.n1210 3.4105
R9599 GNDA.n1317 GNDA.n1233 3.4105
R9600 GNDA.n1317 GNDA.n1209 3.4105
R9601 GNDA.n1317 GNDA.n1234 3.4105
R9602 GNDA.n1317 GNDA.n1208 3.4105
R9603 GNDA.n1317 GNDA.n1235 3.4105
R9604 GNDA.n1317 GNDA.n1207 3.4105
R9605 GNDA.n1317 GNDA.n1236 3.4105
R9606 GNDA.n1317 GNDA.n1206 3.4105
R9607 GNDA.n1317 GNDA.n1237 3.4105
R9608 GNDA.n2583 GNDA.n1317 3.4105
R9609 GNDA.n1320 GNDA.n1239 3.4105
R9610 GNDA.n1239 GNDA.n1222 3.4105
R9611 GNDA.n1239 GNDA.n1220 3.4105
R9612 GNDA.n1239 GNDA.n1223 3.4105
R9613 GNDA.n1239 GNDA.n1219 3.4105
R9614 GNDA.n1239 GNDA.n1224 3.4105
R9615 GNDA.n1239 GNDA.n1218 3.4105
R9616 GNDA.n1239 GNDA.n1225 3.4105
R9617 GNDA.n1239 GNDA.n1217 3.4105
R9618 GNDA.n1239 GNDA.n1226 3.4105
R9619 GNDA.n1239 GNDA.n1216 3.4105
R9620 GNDA.n1239 GNDA.n1227 3.4105
R9621 GNDA.n1239 GNDA.n1215 3.4105
R9622 GNDA.n1239 GNDA.n1228 3.4105
R9623 GNDA.n1239 GNDA.n1214 3.4105
R9624 GNDA.n1239 GNDA.n1229 3.4105
R9625 GNDA.n1239 GNDA.n1213 3.4105
R9626 GNDA.n1239 GNDA.n1230 3.4105
R9627 GNDA.n1239 GNDA.n1212 3.4105
R9628 GNDA.n1239 GNDA.n1231 3.4105
R9629 GNDA.n1239 GNDA.n1211 3.4105
R9630 GNDA.n1239 GNDA.n1232 3.4105
R9631 GNDA.n1239 GNDA.n1210 3.4105
R9632 GNDA.n1239 GNDA.n1233 3.4105
R9633 GNDA.n1239 GNDA.n1209 3.4105
R9634 GNDA.n1239 GNDA.n1234 3.4105
R9635 GNDA.n1239 GNDA.n1208 3.4105
R9636 GNDA.n1239 GNDA.n1235 3.4105
R9637 GNDA.n1239 GNDA.n1207 3.4105
R9638 GNDA.n1239 GNDA.n1236 3.4105
R9639 GNDA.n1239 GNDA.n1206 3.4105
R9640 GNDA.n1239 GNDA.n1237 3.4105
R9641 GNDA.n2583 GNDA.n1239 3.4105
R9642 GNDA.n2582 GNDA.n1320 3.4105
R9643 GNDA.n2582 GNDA.n1222 3.4105
R9644 GNDA.n2582 GNDA.n1220 3.4105
R9645 GNDA.n2582 GNDA.n1223 3.4105
R9646 GNDA.n2582 GNDA.n1219 3.4105
R9647 GNDA.n2582 GNDA.n1224 3.4105
R9648 GNDA.n2582 GNDA.n1218 3.4105
R9649 GNDA.n2582 GNDA.n1225 3.4105
R9650 GNDA.n2582 GNDA.n1217 3.4105
R9651 GNDA.n2582 GNDA.n1226 3.4105
R9652 GNDA.n2582 GNDA.n1216 3.4105
R9653 GNDA.n2582 GNDA.n1227 3.4105
R9654 GNDA.n2582 GNDA.n1215 3.4105
R9655 GNDA.n2582 GNDA.n1228 3.4105
R9656 GNDA.n2582 GNDA.n1214 3.4105
R9657 GNDA.n2582 GNDA.n1229 3.4105
R9658 GNDA.n2582 GNDA.n1213 3.4105
R9659 GNDA.n2582 GNDA.n1230 3.4105
R9660 GNDA.n2582 GNDA.n1212 3.4105
R9661 GNDA.n2582 GNDA.n1231 3.4105
R9662 GNDA.n2582 GNDA.n1211 3.4105
R9663 GNDA.n2582 GNDA.n1232 3.4105
R9664 GNDA.n2582 GNDA.n1210 3.4105
R9665 GNDA.n2582 GNDA.n1233 3.4105
R9666 GNDA.n2582 GNDA.n1209 3.4105
R9667 GNDA.n2582 GNDA.n1234 3.4105
R9668 GNDA.n2582 GNDA.n1208 3.4105
R9669 GNDA.n2582 GNDA.n1235 3.4105
R9670 GNDA.n2582 GNDA.n1207 3.4105
R9671 GNDA.n2582 GNDA.n1236 3.4105
R9672 GNDA.n2582 GNDA.n1206 3.4105
R9673 GNDA.n2582 GNDA.n1237 3.4105
R9674 GNDA.n2583 GNDA.n2582 3.4105
R9675 GNDA.n1320 GNDA.n1238 3.4105
R9676 GNDA.n1238 GNDA.n1222 3.4105
R9677 GNDA.n1238 GNDA.n1220 3.4105
R9678 GNDA.n1238 GNDA.n1223 3.4105
R9679 GNDA.n1238 GNDA.n1219 3.4105
R9680 GNDA.n1238 GNDA.n1224 3.4105
R9681 GNDA.n1238 GNDA.n1218 3.4105
R9682 GNDA.n1238 GNDA.n1225 3.4105
R9683 GNDA.n1238 GNDA.n1217 3.4105
R9684 GNDA.n1238 GNDA.n1226 3.4105
R9685 GNDA.n1238 GNDA.n1216 3.4105
R9686 GNDA.n1238 GNDA.n1227 3.4105
R9687 GNDA.n1238 GNDA.n1215 3.4105
R9688 GNDA.n1238 GNDA.n1228 3.4105
R9689 GNDA.n1238 GNDA.n1214 3.4105
R9690 GNDA.n1238 GNDA.n1229 3.4105
R9691 GNDA.n1238 GNDA.n1213 3.4105
R9692 GNDA.n1238 GNDA.n1230 3.4105
R9693 GNDA.n1238 GNDA.n1212 3.4105
R9694 GNDA.n1238 GNDA.n1231 3.4105
R9695 GNDA.n1238 GNDA.n1211 3.4105
R9696 GNDA.n1238 GNDA.n1232 3.4105
R9697 GNDA.n1238 GNDA.n1210 3.4105
R9698 GNDA.n1238 GNDA.n1233 3.4105
R9699 GNDA.n1238 GNDA.n1209 3.4105
R9700 GNDA.n1238 GNDA.n1234 3.4105
R9701 GNDA.n1238 GNDA.n1208 3.4105
R9702 GNDA.n1238 GNDA.n1235 3.4105
R9703 GNDA.n1238 GNDA.n1207 3.4105
R9704 GNDA.n1238 GNDA.n1236 3.4105
R9705 GNDA.n1238 GNDA.n1206 3.4105
R9706 GNDA.n1238 GNDA.n1237 3.4105
R9707 GNDA.n2583 GNDA.n1238 3.4105
R9708 GNDA.n2584 GNDA.n1222 3.4105
R9709 GNDA.n2584 GNDA.n1220 3.4105
R9710 GNDA.n2584 GNDA.n1223 3.4105
R9711 GNDA.n2584 GNDA.n1219 3.4105
R9712 GNDA.n2584 GNDA.n1224 3.4105
R9713 GNDA.n2584 GNDA.n1218 3.4105
R9714 GNDA.n2584 GNDA.n1225 3.4105
R9715 GNDA.n2584 GNDA.n1217 3.4105
R9716 GNDA.n2584 GNDA.n1226 3.4105
R9717 GNDA.n2584 GNDA.n1216 3.4105
R9718 GNDA.n2584 GNDA.n1227 3.4105
R9719 GNDA.n2584 GNDA.n1215 3.4105
R9720 GNDA.n2584 GNDA.n1228 3.4105
R9721 GNDA.n2584 GNDA.n1214 3.4105
R9722 GNDA.n2584 GNDA.n1229 3.4105
R9723 GNDA.n2584 GNDA.n1213 3.4105
R9724 GNDA.n2584 GNDA.n1230 3.4105
R9725 GNDA.n2584 GNDA.n1212 3.4105
R9726 GNDA.n2584 GNDA.n1231 3.4105
R9727 GNDA.n2584 GNDA.n1211 3.4105
R9728 GNDA.n2584 GNDA.n1232 3.4105
R9729 GNDA.n2584 GNDA.n1210 3.4105
R9730 GNDA.n2584 GNDA.n1233 3.4105
R9731 GNDA.n2584 GNDA.n1209 3.4105
R9732 GNDA.n2584 GNDA.n1234 3.4105
R9733 GNDA.n2584 GNDA.n1208 3.4105
R9734 GNDA.n2584 GNDA.n1235 3.4105
R9735 GNDA.n2584 GNDA.n1207 3.4105
R9736 GNDA.n2584 GNDA.n1236 3.4105
R9737 GNDA.n2584 GNDA.n1206 3.4105
R9738 GNDA.n2584 GNDA.n1237 3.4105
R9739 GNDA.n2584 GNDA.n2583 3.4105
R9740 GNDA.n2690 GNDA.n2689 3.4105
R9741 GNDA.n2691 GNDA.n2690 3.4105
R9742 GNDA.n2693 GNDA.n1057 3.4105
R9743 GNDA.n2689 GNDA.n1057 3.4105
R9744 GNDA.n2691 GNDA.n1057 3.4105
R9745 GNDA.n2693 GNDA.n1059 3.4105
R9746 GNDA.n1090 GNDA.n1059 3.4105
R9747 GNDA.n1092 GNDA.n1059 3.4105
R9748 GNDA.n1089 GNDA.n1059 3.4105
R9749 GNDA.n1094 GNDA.n1059 3.4105
R9750 GNDA.n1088 GNDA.n1059 3.4105
R9751 GNDA.n1096 GNDA.n1059 3.4105
R9752 GNDA.n1087 GNDA.n1059 3.4105
R9753 GNDA.n1098 GNDA.n1059 3.4105
R9754 GNDA.n1086 GNDA.n1059 3.4105
R9755 GNDA.n1100 GNDA.n1059 3.4105
R9756 GNDA.n1085 GNDA.n1059 3.4105
R9757 GNDA.n1102 GNDA.n1059 3.4105
R9758 GNDA.n1084 GNDA.n1059 3.4105
R9759 GNDA.n1104 GNDA.n1059 3.4105
R9760 GNDA.n1083 GNDA.n1059 3.4105
R9761 GNDA.n1106 GNDA.n1059 3.4105
R9762 GNDA.n1082 GNDA.n1059 3.4105
R9763 GNDA.n1108 GNDA.n1059 3.4105
R9764 GNDA.n1081 GNDA.n1059 3.4105
R9765 GNDA.n1110 GNDA.n1059 3.4105
R9766 GNDA.n1080 GNDA.n1059 3.4105
R9767 GNDA.n1112 GNDA.n1059 3.4105
R9768 GNDA.n1079 GNDA.n1059 3.4105
R9769 GNDA.n1114 GNDA.n1059 3.4105
R9770 GNDA.n1078 GNDA.n1059 3.4105
R9771 GNDA.n1116 GNDA.n1059 3.4105
R9772 GNDA.n1077 GNDA.n1059 3.4105
R9773 GNDA.n1118 GNDA.n1059 3.4105
R9774 GNDA.n1076 GNDA.n1059 3.4105
R9775 GNDA.n1120 GNDA.n1059 3.4105
R9776 GNDA.n2689 GNDA.n1059 3.4105
R9777 GNDA.n2691 GNDA.n1059 3.4105
R9778 GNDA.n2693 GNDA.n1056 3.4105
R9779 GNDA.n1090 GNDA.n1056 3.4105
R9780 GNDA.n1092 GNDA.n1056 3.4105
R9781 GNDA.n1089 GNDA.n1056 3.4105
R9782 GNDA.n1094 GNDA.n1056 3.4105
R9783 GNDA.n1088 GNDA.n1056 3.4105
R9784 GNDA.n1096 GNDA.n1056 3.4105
R9785 GNDA.n1087 GNDA.n1056 3.4105
R9786 GNDA.n1098 GNDA.n1056 3.4105
R9787 GNDA.n1086 GNDA.n1056 3.4105
R9788 GNDA.n1100 GNDA.n1056 3.4105
R9789 GNDA.n1085 GNDA.n1056 3.4105
R9790 GNDA.n1102 GNDA.n1056 3.4105
R9791 GNDA.n1084 GNDA.n1056 3.4105
R9792 GNDA.n1104 GNDA.n1056 3.4105
R9793 GNDA.n1083 GNDA.n1056 3.4105
R9794 GNDA.n1106 GNDA.n1056 3.4105
R9795 GNDA.n1082 GNDA.n1056 3.4105
R9796 GNDA.n1108 GNDA.n1056 3.4105
R9797 GNDA.n1081 GNDA.n1056 3.4105
R9798 GNDA.n1110 GNDA.n1056 3.4105
R9799 GNDA.n1080 GNDA.n1056 3.4105
R9800 GNDA.n1112 GNDA.n1056 3.4105
R9801 GNDA.n1079 GNDA.n1056 3.4105
R9802 GNDA.n1114 GNDA.n1056 3.4105
R9803 GNDA.n1078 GNDA.n1056 3.4105
R9804 GNDA.n1116 GNDA.n1056 3.4105
R9805 GNDA.n1077 GNDA.n1056 3.4105
R9806 GNDA.n1118 GNDA.n1056 3.4105
R9807 GNDA.n1076 GNDA.n1056 3.4105
R9808 GNDA.n1120 GNDA.n1056 3.4105
R9809 GNDA.n2689 GNDA.n1056 3.4105
R9810 GNDA.n2691 GNDA.n1056 3.4105
R9811 GNDA.n2693 GNDA.n1060 3.4105
R9812 GNDA.n1090 GNDA.n1060 3.4105
R9813 GNDA.n1092 GNDA.n1060 3.4105
R9814 GNDA.n1089 GNDA.n1060 3.4105
R9815 GNDA.n1094 GNDA.n1060 3.4105
R9816 GNDA.n1088 GNDA.n1060 3.4105
R9817 GNDA.n1096 GNDA.n1060 3.4105
R9818 GNDA.n1087 GNDA.n1060 3.4105
R9819 GNDA.n1098 GNDA.n1060 3.4105
R9820 GNDA.n1086 GNDA.n1060 3.4105
R9821 GNDA.n1100 GNDA.n1060 3.4105
R9822 GNDA.n1085 GNDA.n1060 3.4105
R9823 GNDA.n1102 GNDA.n1060 3.4105
R9824 GNDA.n1084 GNDA.n1060 3.4105
R9825 GNDA.n1104 GNDA.n1060 3.4105
R9826 GNDA.n1083 GNDA.n1060 3.4105
R9827 GNDA.n1106 GNDA.n1060 3.4105
R9828 GNDA.n1082 GNDA.n1060 3.4105
R9829 GNDA.n1108 GNDA.n1060 3.4105
R9830 GNDA.n1081 GNDA.n1060 3.4105
R9831 GNDA.n1110 GNDA.n1060 3.4105
R9832 GNDA.n1080 GNDA.n1060 3.4105
R9833 GNDA.n1112 GNDA.n1060 3.4105
R9834 GNDA.n1079 GNDA.n1060 3.4105
R9835 GNDA.n1114 GNDA.n1060 3.4105
R9836 GNDA.n1078 GNDA.n1060 3.4105
R9837 GNDA.n1116 GNDA.n1060 3.4105
R9838 GNDA.n1077 GNDA.n1060 3.4105
R9839 GNDA.n1118 GNDA.n1060 3.4105
R9840 GNDA.n1076 GNDA.n1060 3.4105
R9841 GNDA.n1120 GNDA.n1060 3.4105
R9842 GNDA.n2689 GNDA.n1060 3.4105
R9843 GNDA.n2691 GNDA.n1060 3.4105
R9844 GNDA.n2693 GNDA.n1055 3.4105
R9845 GNDA.n1090 GNDA.n1055 3.4105
R9846 GNDA.n1092 GNDA.n1055 3.4105
R9847 GNDA.n1089 GNDA.n1055 3.4105
R9848 GNDA.n1094 GNDA.n1055 3.4105
R9849 GNDA.n1088 GNDA.n1055 3.4105
R9850 GNDA.n1096 GNDA.n1055 3.4105
R9851 GNDA.n1087 GNDA.n1055 3.4105
R9852 GNDA.n1098 GNDA.n1055 3.4105
R9853 GNDA.n1086 GNDA.n1055 3.4105
R9854 GNDA.n1100 GNDA.n1055 3.4105
R9855 GNDA.n1085 GNDA.n1055 3.4105
R9856 GNDA.n1102 GNDA.n1055 3.4105
R9857 GNDA.n1084 GNDA.n1055 3.4105
R9858 GNDA.n1104 GNDA.n1055 3.4105
R9859 GNDA.n1083 GNDA.n1055 3.4105
R9860 GNDA.n1106 GNDA.n1055 3.4105
R9861 GNDA.n1082 GNDA.n1055 3.4105
R9862 GNDA.n1108 GNDA.n1055 3.4105
R9863 GNDA.n1081 GNDA.n1055 3.4105
R9864 GNDA.n1110 GNDA.n1055 3.4105
R9865 GNDA.n1080 GNDA.n1055 3.4105
R9866 GNDA.n1112 GNDA.n1055 3.4105
R9867 GNDA.n1079 GNDA.n1055 3.4105
R9868 GNDA.n1114 GNDA.n1055 3.4105
R9869 GNDA.n1078 GNDA.n1055 3.4105
R9870 GNDA.n1116 GNDA.n1055 3.4105
R9871 GNDA.n1077 GNDA.n1055 3.4105
R9872 GNDA.n1118 GNDA.n1055 3.4105
R9873 GNDA.n1076 GNDA.n1055 3.4105
R9874 GNDA.n1120 GNDA.n1055 3.4105
R9875 GNDA.n2689 GNDA.n1055 3.4105
R9876 GNDA.n2691 GNDA.n1055 3.4105
R9877 GNDA.n2693 GNDA.n1061 3.4105
R9878 GNDA.n1090 GNDA.n1061 3.4105
R9879 GNDA.n1092 GNDA.n1061 3.4105
R9880 GNDA.n1089 GNDA.n1061 3.4105
R9881 GNDA.n1094 GNDA.n1061 3.4105
R9882 GNDA.n1088 GNDA.n1061 3.4105
R9883 GNDA.n1096 GNDA.n1061 3.4105
R9884 GNDA.n1087 GNDA.n1061 3.4105
R9885 GNDA.n1098 GNDA.n1061 3.4105
R9886 GNDA.n1086 GNDA.n1061 3.4105
R9887 GNDA.n1100 GNDA.n1061 3.4105
R9888 GNDA.n1085 GNDA.n1061 3.4105
R9889 GNDA.n1102 GNDA.n1061 3.4105
R9890 GNDA.n1084 GNDA.n1061 3.4105
R9891 GNDA.n1104 GNDA.n1061 3.4105
R9892 GNDA.n1083 GNDA.n1061 3.4105
R9893 GNDA.n1106 GNDA.n1061 3.4105
R9894 GNDA.n1082 GNDA.n1061 3.4105
R9895 GNDA.n1108 GNDA.n1061 3.4105
R9896 GNDA.n1081 GNDA.n1061 3.4105
R9897 GNDA.n1110 GNDA.n1061 3.4105
R9898 GNDA.n1080 GNDA.n1061 3.4105
R9899 GNDA.n1112 GNDA.n1061 3.4105
R9900 GNDA.n1079 GNDA.n1061 3.4105
R9901 GNDA.n1114 GNDA.n1061 3.4105
R9902 GNDA.n1078 GNDA.n1061 3.4105
R9903 GNDA.n1116 GNDA.n1061 3.4105
R9904 GNDA.n1077 GNDA.n1061 3.4105
R9905 GNDA.n1118 GNDA.n1061 3.4105
R9906 GNDA.n1076 GNDA.n1061 3.4105
R9907 GNDA.n1120 GNDA.n1061 3.4105
R9908 GNDA.n2689 GNDA.n1061 3.4105
R9909 GNDA.n2691 GNDA.n1061 3.4105
R9910 GNDA.n2693 GNDA.n1054 3.4105
R9911 GNDA.n1090 GNDA.n1054 3.4105
R9912 GNDA.n1092 GNDA.n1054 3.4105
R9913 GNDA.n1089 GNDA.n1054 3.4105
R9914 GNDA.n1094 GNDA.n1054 3.4105
R9915 GNDA.n1088 GNDA.n1054 3.4105
R9916 GNDA.n1096 GNDA.n1054 3.4105
R9917 GNDA.n1087 GNDA.n1054 3.4105
R9918 GNDA.n1098 GNDA.n1054 3.4105
R9919 GNDA.n1086 GNDA.n1054 3.4105
R9920 GNDA.n1100 GNDA.n1054 3.4105
R9921 GNDA.n1085 GNDA.n1054 3.4105
R9922 GNDA.n1102 GNDA.n1054 3.4105
R9923 GNDA.n1084 GNDA.n1054 3.4105
R9924 GNDA.n1104 GNDA.n1054 3.4105
R9925 GNDA.n1083 GNDA.n1054 3.4105
R9926 GNDA.n1106 GNDA.n1054 3.4105
R9927 GNDA.n1082 GNDA.n1054 3.4105
R9928 GNDA.n1108 GNDA.n1054 3.4105
R9929 GNDA.n1081 GNDA.n1054 3.4105
R9930 GNDA.n1110 GNDA.n1054 3.4105
R9931 GNDA.n1080 GNDA.n1054 3.4105
R9932 GNDA.n1112 GNDA.n1054 3.4105
R9933 GNDA.n1079 GNDA.n1054 3.4105
R9934 GNDA.n1114 GNDA.n1054 3.4105
R9935 GNDA.n1078 GNDA.n1054 3.4105
R9936 GNDA.n1116 GNDA.n1054 3.4105
R9937 GNDA.n1077 GNDA.n1054 3.4105
R9938 GNDA.n1118 GNDA.n1054 3.4105
R9939 GNDA.n1076 GNDA.n1054 3.4105
R9940 GNDA.n1120 GNDA.n1054 3.4105
R9941 GNDA.n2689 GNDA.n1054 3.4105
R9942 GNDA.n2691 GNDA.n1054 3.4105
R9943 GNDA.n2693 GNDA.n1062 3.4105
R9944 GNDA.n1090 GNDA.n1062 3.4105
R9945 GNDA.n1092 GNDA.n1062 3.4105
R9946 GNDA.n1089 GNDA.n1062 3.4105
R9947 GNDA.n1094 GNDA.n1062 3.4105
R9948 GNDA.n1088 GNDA.n1062 3.4105
R9949 GNDA.n1096 GNDA.n1062 3.4105
R9950 GNDA.n1087 GNDA.n1062 3.4105
R9951 GNDA.n1098 GNDA.n1062 3.4105
R9952 GNDA.n1086 GNDA.n1062 3.4105
R9953 GNDA.n1100 GNDA.n1062 3.4105
R9954 GNDA.n1085 GNDA.n1062 3.4105
R9955 GNDA.n1102 GNDA.n1062 3.4105
R9956 GNDA.n1084 GNDA.n1062 3.4105
R9957 GNDA.n1104 GNDA.n1062 3.4105
R9958 GNDA.n1083 GNDA.n1062 3.4105
R9959 GNDA.n1106 GNDA.n1062 3.4105
R9960 GNDA.n1082 GNDA.n1062 3.4105
R9961 GNDA.n1108 GNDA.n1062 3.4105
R9962 GNDA.n1081 GNDA.n1062 3.4105
R9963 GNDA.n1110 GNDA.n1062 3.4105
R9964 GNDA.n1080 GNDA.n1062 3.4105
R9965 GNDA.n1112 GNDA.n1062 3.4105
R9966 GNDA.n1079 GNDA.n1062 3.4105
R9967 GNDA.n1114 GNDA.n1062 3.4105
R9968 GNDA.n1078 GNDA.n1062 3.4105
R9969 GNDA.n1116 GNDA.n1062 3.4105
R9970 GNDA.n1077 GNDA.n1062 3.4105
R9971 GNDA.n1118 GNDA.n1062 3.4105
R9972 GNDA.n1076 GNDA.n1062 3.4105
R9973 GNDA.n1120 GNDA.n1062 3.4105
R9974 GNDA.n2689 GNDA.n1062 3.4105
R9975 GNDA.n2691 GNDA.n1062 3.4105
R9976 GNDA.n2693 GNDA.n1053 3.4105
R9977 GNDA.n1090 GNDA.n1053 3.4105
R9978 GNDA.n1092 GNDA.n1053 3.4105
R9979 GNDA.n1089 GNDA.n1053 3.4105
R9980 GNDA.n1094 GNDA.n1053 3.4105
R9981 GNDA.n1088 GNDA.n1053 3.4105
R9982 GNDA.n1096 GNDA.n1053 3.4105
R9983 GNDA.n1087 GNDA.n1053 3.4105
R9984 GNDA.n1098 GNDA.n1053 3.4105
R9985 GNDA.n1086 GNDA.n1053 3.4105
R9986 GNDA.n1100 GNDA.n1053 3.4105
R9987 GNDA.n1085 GNDA.n1053 3.4105
R9988 GNDA.n1102 GNDA.n1053 3.4105
R9989 GNDA.n1084 GNDA.n1053 3.4105
R9990 GNDA.n1104 GNDA.n1053 3.4105
R9991 GNDA.n1083 GNDA.n1053 3.4105
R9992 GNDA.n1106 GNDA.n1053 3.4105
R9993 GNDA.n1082 GNDA.n1053 3.4105
R9994 GNDA.n1108 GNDA.n1053 3.4105
R9995 GNDA.n1081 GNDA.n1053 3.4105
R9996 GNDA.n1110 GNDA.n1053 3.4105
R9997 GNDA.n1080 GNDA.n1053 3.4105
R9998 GNDA.n1112 GNDA.n1053 3.4105
R9999 GNDA.n1079 GNDA.n1053 3.4105
R10000 GNDA.n1114 GNDA.n1053 3.4105
R10001 GNDA.n1078 GNDA.n1053 3.4105
R10002 GNDA.n1116 GNDA.n1053 3.4105
R10003 GNDA.n1077 GNDA.n1053 3.4105
R10004 GNDA.n1118 GNDA.n1053 3.4105
R10005 GNDA.n1076 GNDA.n1053 3.4105
R10006 GNDA.n1120 GNDA.n1053 3.4105
R10007 GNDA.n2689 GNDA.n1053 3.4105
R10008 GNDA.n2691 GNDA.n1053 3.4105
R10009 GNDA.n2693 GNDA.n1063 3.4105
R10010 GNDA.n1090 GNDA.n1063 3.4105
R10011 GNDA.n1092 GNDA.n1063 3.4105
R10012 GNDA.n1089 GNDA.n1063 3.4105
R10013 GNDA.n1094 GNDA.n1063 3.4105
R10014 GNDA.n1088 GNDA.n1063 3.4105
R10015 GNDA.n1096 GNDA.n1063 3.4105
R10016 GNDA.n1087 GNDA.n1063 3.4105
R10017 GNDA.n1098 GNDA.n1063 3.4105
R10018 GNDA.n1086 GNDA.n1063 3.4105
R10019 GNDA.n1100 GNDA.n1063 3.4105
R10020 GNDA.n1085 GNDA.n1063 3.4105
R10021 GNDA.n1102 GNDA.n1063 3.4105
R10022 GNDA.n1084 GNDA.n1063 3.4105
R10023 GNDA.n1104 GNDA.n1063 3.4105
R10024 GNDA.n1083 GNDA.n1063 3.4105
R10025 GNDA.n1106 GNDA.n1063 3.4105
R10026 GNDA.n1082 GNDA.n1063 3.4105
R10027 GNDA.n1108 GNDA.n1063 3.4105
R10028 GNDA.n1081 GNDA.n1063 3.4105
R10029 GNDA.n1110 GNDA.n1063 3.4105
R10030 GNDA.n1080 GNDA.n1063 3.4105
R10031 GNDA.n1112 GNDA.n1063 3.4105
R10032 GNDA.n1079 GNDA.n1063 3.4105
R10033 GNDA.n1114 GNDA.n1063 3.4105
R10034 GNDA.n1078 GNDA.n1063 3.4105
R10035 GNDA.n1116 GNDA.n1063 3.4105
R10036 GNDA.n1077 GNDA.n1063 3.4105
R10037 GNDA.n1118 GNDA.n1063 3.4105
R10038 GNDA.n1076 GNDA.n1063 3.4105
R10039 GNDA.n1120 GNDA.n1063 3.4105
R10040 GNDA.n2689 GNDA.n1063 3.4105
R10041 GNDA.n2691 GNDA.n1063 3.4105
R10042 GNDA.n2693 GNDA.n1052 3.4105
R10043 GNDA.n1090 GNDA.n1052 3.4105
R10044 GNDA.n1092 GNDA.n1052 3.4105
R10045 GNDA.n1089 GNDA.n1052 3.4105
R10046 GNDA.n1094 GNDA.n1052 3.4105
R10047 GNDA.n1088 GNDA.n1052 3.4105
R10048 GNDA.n1096 GNDA.n1052 3.4105
R10049 GNDA.n1087 GNDA.n1052 3.4105
R10050 GNDA.n1098 GNDA.n1052 3.4105
R10051 GNDA.n1086 GNDA.n1052 3.4105
R10052 GNDA.n1100 GNDA.n1052 3.4105
R10053 GNDA.n1085 GNDA.n1052 3.4105
R10054 GNDA.n1102 GNDA.n1052 3.4105
R10055 GNDA.n1084 GNDA.n1052 3.4105
R10056 GNDA.n1104 GNDA.n1052 3.4105
R10057 GNDA.n1083 GNDA.n1052 3.4105
R10058 GNDA.n1106 GNDA.n1052 3.4105
R10059 GNDA.n1082 GNDA.n1052 3.4105
R10060 GNDA.n1108 GNDA.n1052 3.4105
R10061 GNDA.n1081 GNDA.n1052 3.4105
R10062 GNDA.n1110 GNDA.n1052 3.4105
R10063 GNDA.n1080 GNDA.n1052 3.4105
R10064 GNDA.n1112 GNDA.n1052 3.4105
R10065 GNDA.n1079 GNDA.n1052 3.4105
R10066 GNDA.n1114 GNDA.n1052 3.4105
R10067 GNDA.n1078 GNDA.n1052 3.4105
R10068 GNDA.n1116 GNDA.n1052 3.4105
R10069 GNDA.n1077 GNDA.n1052 3.4105
R10070 GNDA.n1118 GNDA.n1052 3.4105
R10071 GNDA.n1076 GNDA.n1052 3.4105
R10072 GNDA.n1120 GNDA.n1052 3.4105
R10073 GNDA.n2689 GNDA.n1052 3.4105
R10074 GNDA.n2691 GNDA.n1052 3.4105
R10075 GNDA.n2693 GNDA.n1064 3.4105
R10076 GNDA.n1090 GNDA.n1064 3.4105
R10077 GNDA.n1092 GNDA.n1064 3.4105
R10078 GNDA.n1089 GNDA.n1064 3.4105
R10079 GNDA.n1094 GNDA.n1064 3.4105
R10080 GNDA.n1088 GNDA.n1064 3.4105
R10081 GNDA.n1096 GNDA.n1064 3.4105
R10082 GNDA.n1087 GNDA.n1064 3.4105
R10083 GNDA.n1098 GNDA.n1064 3.4105
R10084 GNDA.n1086 GNDA.n1064 3.4105
R10085 GNDA.n1100 GNDA.n1064 3.4105
R10086 GNDA.n1085 GNDA.n1064 3.4105
R10087 GNDA.n1102 GNDA.n1064 3.4105
R10088 GNDA.n1084 GNDA.n1064 3.4105
R10089 GNDA.n1104 GNDA.n1064 3.4105
R10090 GNDA.n1083 GNDA.n1064 3.4105
R10091 GNDA.n1106 GNDA.n1064 3.4105
R10092 GNDA.n1082 GNDA.n1064 3.4105
R10093 GNDA.n1108 GNDA.n1064 3.4105
R10094 GNDA.n1081 GNDA.n1064 3.4105
R10095 GNDA.n1110 GNDA.n1064 3.4105
R10096 GNDA.n1080 GNDA.n1064 3.4105
R10097 GNDA.n1112 GNDA.n1064 3.4105
R10098 GNDA.n1079 GNDA.n1064 3.4105
R10099 GNDA.n1114 GNDA.n1064 3.4105
R10100 GNDA.n1078 GNDA.n1064 3.4105
R10101 GNDA.n1116 GNDA.n1064 3.4105
R10102 GNDA.n1077 GNDA.n1064 3.4105
R10103 GNDA.n1118 GNDA.n1064 3.4105
R10104 GNDA.n1076 GNDA.n1064 3.4105
R10105 GNDA.n1120 GNDA.n1064 3.4105
R10106 GNDA.n2689 GNDA.n1064 3.4105
R10107 GNDA.n2691 GNDA.n1064 3.4105
R10108 GNDA.n2693 GNDA.n1051 3.4105
R10109 GNDA.n1090 GNDA.n1051 3.4105
R10110 GNDA.n1092 GNDA.n1051 3.4105
R10111 GNDA.n1089 GNDA.n1051 3.4105
R10112 GNDA.n1094 GNDA.n1051 3.4105
R10113 GNDA.n1088 GNDA.n1051 3.4105
R10114 GNDA.n1096 GNDA.n1051 3.4105
R10115 GNDA.n1087 GNDA.n1051 3.4105
R10116 GNDA.n1098 GNDA.n1051 3.4105
R10117 GNDA.n1086 GNDA.n1051 3.4105
R10118 GNDA.n1100 GNDA.n1051 3.4105
R10119 GNDA.n1085 GNDA.n1051 3.4105
R10120 GNDA.n1102 GNDA.n1051 3.4105
R10121 GNDA.n1084 GNDA.n1051 3.4105
R10122 GNDA.n1104 GNDA.n1051 3.4105
R10123 GNDA.n1083 GNDA.n1051 3.4105
R10124 GNDA.n1106 GNDA.n1051 3.4105
R10125 GNDA.n1082 GNDA.n1051 3.4105
R10126 GNDA.n1108 GNDA.n1051 3.4105
R10127 GNDA.n1081 GNDA.n1051 3.4105
R10128 GNDA.n1110 GNDA.n1051 3.4105
R10129 GNDA.n1080 GNDA.n1051 3.4105
R10130 GNDA.n1112 GNDA.n1051 3.4105
R10131 GNDA.n1079 GNDA.n1051 3.4105
R10132 GNDA.n1114 GNDA.n1051 3.4105
R10133 GNDA.n1078 GNDA.n1051 3.4105
R10134 GNDA.n1116 GNDA.n1051 3.4105
R10135 GNDA.n1077 GNDA.n1051 3.4105
R10136 GNDA.n1118 GNDA.n1051 3.4105
R10137 GNDA.n1076 GNDA.n1051 3.4105
R10138 GNDA.n1120 GNDA.n1051 3.4105
R10139 GNDA.n2689 GNDA.n1051 3.4105
R10140 GNDA.n2691 GNDA.n1051 3.4105
R10141 GNDA.n2693 GNDA.n1065 3.4105
R10142 GNDA.n1090 GNDA.n1065 3.4105
R10143 GNDA.n1092 GNDA.n1065 3.4105
R10144 GNDA.n1089 GNDA.n1065 3.4105
R10145 GNDA.n1094 GNDA.n1065 3.4105
R10146 GNDA.n1088 GNDA.n1065 3.4105
R10147 GNDA.n1096 GNDA.n1065 3.4105
R10148 GNDA.n1087 GNDA.n1065 3.4105
R10149 GNDA.n1098 GNDA.n1065 3.4105
R10150 GNDA.n1086 GNDA.n1065 3.4105
R10151 GNDA.n1100 GNDA.n1065 3.4105
R10152 GNDA.n1085 GNDA.n1065 3.4105
R10153 GNDA.n1102 GNDA.n1065 3.4105
R10154 GNDA.n1084 GNDA.n1065 3.4105
R10155 GNDA.n1104 GNDA.n1065 3.4105
R10156 GNDA.n1083 GNDA.n1065 3.4105
R10157 GNDA.n1106 GNDA.n1065 3.4105
R10158 GNDA.n1082 GNDA.n1065 3.4105
R10159 GNDA.n1108 GNDA.n1065 3.4105
R10160 GNDA.n1081 GNDA.n1065 3.4105
R10161 GNDA.n1110 GNDA.n1065 3.4105
R10162 GNDA.n1080 GNDA.n1065 3.4105
R10163 GNDA.n1112 GNDA.n1065 3.4105
R10164 GNDA.n1079 GNDA.n1065 3.4105
R10165 GNDA.n1114 GNDA.n1065 3.4105
R10166 GNDA.n1078 GNDA.n1065 3.4105
R10167 GNDA.n1116 GNDA.n1065 3.4105
R10168 GNDA.n1077 GNDA.n1065 3.4105
R10169 GNDA.n1118 GNDA.n1065 3.4105
R10170 GNDA.n1076 GNDA.n1065 3.4105
R10171 GNDA.n1120 GNDA.n1065 3.4105
R10172 GNDA.n2689 GNDA.n1065 3.4105
R10173 GNDA.n2691 GNDA.n1065 3.4105
R10174 GNDA.n2693 GNDA.n1050 3.4105
R10175 GNDA.n1090 GNDA.n1050 3.4105
R10176 GNDA.n1092 GNDA.n1050 3.4105
R10177 GNDA.n1089 GNDA.n1050 3.4105
R10178 GNDA.n1094 GNDA.n1050 3.4105
R10179 GNDA.n1088 GNDA.n1050 3.4105
R10180 GNDA.n1096 GNDA.n1050 3.4105
R10181 GNDA.n1087 GNDA.n1050 3.4105
R10182 GNDA.n1098 GNDA.n1050 3.4105
R10183 GNDA.n1086 GNDA.n1050 3.4105
R10184 GNDA.n1100 GNDA.n1050 3.4105
R10185 GNDA.n1085 GNDA.n1050 3.4105
R10186 GNDA.n1102 GNDA.n1050 3.4105
R10187 GNDA.n1084 GNDA.n1050 3.4105
R10188 GNDA.n1104 GNDA.n1050 3.4105
R10189 GNDA.n1083 GNDA.n1050 3.4105
R10190 GNDA.n1106 GNDA.n1050 3.4105
R10191 GNDA.n1082 GNDA.n1050 3.4105
R10192 GNDA.n1108 GNDA.n1050 3.4105
R10193 GNDA.n1081 GNDA.n1050 3.4105
R10194 GNDA.n1110 GNDA.n1050 3.4105
R10195 GNDA.n1080 GNDA.n1050 3.4105
R10196 GNDA.n1112 GNDA.n1050 3.4105
R10197 GNDA.n1079 GNDA.n1050 3.4105
R10198 GNDA.n1114 GNDA.n1050 3.4105
R10199 GNDA.n1078 GNDA.n1050 3.4105
R10200 GNDA.n1116 GNDA.n1050 3.4105
R10201 GNDA.n1077 GNDA.n1050 3.4105
R10202 GNDA.n1118 GNDA.n1050 3.4105
R10203 GNDA.n1076 GNDA.n1050 3.4105
R10204 GNDA.n1120 GNDA.n1050 3.4105
R10205 GNDA.n2689 GNDA.n1050 3.4105
R10206 GNDA.n2691 GNDA.n1050 3.4105
R10207 GNDA.n2693 GNDA.n1066 3.4105
R10208 GNDA.n1090 GNDA.n1066 3.4105
R10209 GNDA.n1092 GNDA.n1066 3.4105
R10210 GNDA.n1089 GNDA.n1066 3.4105
R10211 GNDA.n1094 GNDA.n1066 3.4105
R10212 GNDA.n1088 GNDA.n1066 3.4105
R10213 GNDA.n1096 GNDA.n1066 3.4105
R10214 GNDA.n1087 GNDA.n1066 3.4105
R10215 GNDA.n1098 GNDA.n1066 3.4105
R10216 GNDA.n1086 GNDA.n1066 3.4105
R10217 GNDA.n1100 GNDA.n1066 3.4105
R10218 GNDA.n1085 GNDA.n1066 3.4105
R10219 GNDA.n1102 GNDA.n1066 3.4105
R10220 GNDA.n1084 GNDA.n1066 3.4105
R10221 GNDA.n1104 GNDA.n1066 3.4105
R10222 GNDA.n1083 GNDA.n1066 3.4105
R10223 GNDA.n1106 GNDA.n1066 3.4105
R10224 GNDA.n1082 GNDA.n1066 3.4105
R10225 GNDA.n1108 GNDA.n1066 3.4105
R10226 GNDA.n1081 GNDA.n1066 3.4105
R10227 GNDA.n1110 GNDA.n1066 3.4105
R10228 GNDA.n1080 GNDA.n1066 3.4105
R10229 GNDA.n1112 GNDA.n1066 3.4105
R10230 GNDA.n1079 GNDA.n1066 3.4105
R10231 GNDA.n1114 GNDA.n1066 3.4105
R10232 GNDA.n1078 GNDA.n1066 3.4105
R10233 GNDA.n1116 GNDA.n1066 3.4105
R10234 GNDA.n1077 GNDA.n1066 3.4105
R10235 GNDA.n1118 GNDA.n1066 3.4105
R10236 GNDA.n1076 GNDA.n1066 3.4105
R10237 GNDA.n1120 GNDA.n1066 3.4105
R10238 GNDA.n2689 GNDA.n1066 3.4105
R10239 GNDA.n2691 GNDA.n1066 3.4105
R10240 GNDA.n2693 GNDA.n1049 3.4105
R10241 GNDA.n1090 GNDA.n1049 3.4105
R10242 GNDA.n1092 GNDA.n1049 3.4105
R10243 GNDA.n1089 GNDA.n1049 3.4105
R10244 GNDA.n1094 GNDA.n1049 3.4105
R10245 GNDA.n1088 GNDA.n1049 3.4105
R10246 GNDA.n1096 GNDA.n1049 3.4105
R10247 GNDA.n1087 GNDA.n1049 3.4105
R10248 GNDA.n1098 GNDA.n1049 3.4105
R10249 GNDA.n1086 GNDA.n1049 3.4105
R10250 GNDA.n1100 GNDA.n1049 3.4105
R10251 GNDA.n1085 GNDA.n1049 3.4105
R10252 GNDA.n1102 GNDA.n1049 3.4105
R10253 GNDA.n1084 GNDA.n1049 3.4105
R10254 GNDA.n1104 GNDA.n1049 3.4105
R10255 GNDA.n1083 GNDA.n1049 3.4105
R10256 GNDA.n1106 GNDA.n1049 3.4105
R10257 GNDA.n1082 GNDA.n1049 3.4105
R10258 GNDA.n1108 GNDA.n1049 3.4105
R10259 GNDA.n1081 GNDA.n1049 3.4105
R10260 GNDA.n1110 GNDA.n1049 3.4105
R10261 GNDA.n1080 GNDA.n1049 3.4105
R10262 GNDA.n1112 GNDA.n1049 3.4105
R10263 GNDA.n1079 GNDA.n1049 3.4105
R10264 GNDA.n1114 GNDA.n1049 3.4105
R10265 GNDA.n1078 GNDA.n1049 3.4105
R10266 GNDA.n1116 GNDA.n1049 3.4105
R10267 GNDA.n1077 GNDA.n1049 3.4105
R10268 GNDA.n1118 GNDA.n1049 3.4105
R10269 GNDA.n1076 GNDA.n1049 3.4105
R10270 GNDA.n1120 GNDA.n1049 3.4105
R10271 GNDA.n2689 GNDA.n1049 3.4105
R10272 GNDA.n2691 GNDA.n1049 3.4105
R10273 GNDA.n2693 GNDA.n1067 3.4105
R10274 GNDA.n1090 GNDA.n1067 3.4105
R10275 GNDA.n1092 GNDA.n1067 3.4105
R10276 GNDA.n1089 GNDA.n1067 3.4105
R10277 GNDA.n1094 GNDA.n1067 3.4105
R10278 GNDA.n1088 GNDA.n1067 3.4105
R10279 GNDA.n1096 GNDA.n1067 3.4105
R10280 GNDA.n1087 GNDA.n1067 3.4105
R10281 GNDA.n1098 GNDA.n1067 3.4105
R10282 GNDA.n1086 GNDA.n1067 3.4105
R10283 GNDA.n1100 GNDA.n1067 3.4105
R10284 GNDA.n1085 GNDA.n1067 3.4105
R10285 GNDA.n1102 GNDA.n1067 3.4105
R10286 GNDA.n1084 GNDA.n1067 3.4105
R10287 GNDA.n1104 GNDA.n1067 3.4105
R10288 GNDA.n1083 GNDA.n1067 3.4105
R10289 GNDA.n1106 GNDA.n1067 3.4105
R10290 GNDA.n1082 GNDA.n1067 3.4105
R10291 GNDA.n1108 GNDA.n1067 3.4105
R10292 GNDA.n1081 GNDA.n1067 3.4105
R10293 GNDA.n1110 GNDA.n1067 3.4105
R10294 GNDA.n1080 GNDA.n1067 3.4105
R10295 GNDA.n1112 GNDA.n1067 3.4105
R10296 GNDA.n1079 GNDA.n1067 3.4105
R10297 GNDA.n1114 GNDA.n1067 3.4105
R10298 GNDA.n1078 GNDA.n1067 3.4105
R10299 GNDA.n1116 GNDA.n1067 3.4105
R10300 GNDA.n1077 GNDA.n1067 3.4105
R10301 GNDA.n1118 GNDA.n1067 3.4105
R10302 GNDA.n1076 GNDA.n1067 3.4105
R10303 GNDA.n1120 GNDA.n1067 3.4105
R10304 GNDA.n2689 GNDA.n1067 3.4105
R10305 GNDA.n2691 GNDA.n1067 3.4105
R10306 GNDA.n2693 GNDA.n1048 3.4105
R10307 GNDA.n1090 GNDA.n1048 3.4105
R10308 GNDA.n1092 GNDA.n1048 3.4105
R10309 GNDA.n1089 GNDA.n1048 3.4105
R10310 GNDA.n1094 GNDA.n1048 3.4105
R10311 GNDA.n1088 GNDA.n1048 3.4105
R10312 GNDA.n1096 GNDA.n1048 3.4105
R10313 GNDA.n1087 GNDA.n1048 3.4105
R10314 GNDA.n1098 GNDA.n1048 3.4105
R10315 GNDA.n1086 GNDA.n1048 3.4105
R10316 GNDA.n1100 GNDA.n1048 3.4105
R10317 GNDA.n1085 GNDA.n1048 3.4105
R10318 GNDA.n1102 GNDA.n1048 3.4105
R10319 GNDA.n1084 GNDA.n1048 3.4105
R10320 GNDA.n1104 GNDA.n1048 3.4105
R10321 GNDA.n1083 GNDA.n1048 3.4105
R10322 GNDA.n1106 GNDA.n1048 3.4105
R10323 GNDA.n1082 GNDA.n1048 3.4105
R10324 GNDA.n1108 GNDA.n1048 3.4105
R10325 GNDA.n1081 GNDA.n1048 3.4105
R10326 GNDA.n1110 GNDA.n1048 3.4105
R10327 GNDA.n1080 GNDA.n1048 3.4105
R10328 GNDA.n1112 GNDA.n1048 3.4105
R10329 GNDA.n1079 GNDA.n1048 3.4105
R10330 GNDA.n1114 GNDA.n1048 3.4105
R10331 GNDA.n1078 GNDA.n1048 3.4105
R10332 GNDA.n1116 GNDA.n1048 3.4105
R10333 GNDA.n1077 GNDA.n1048 3.4105
R10334 GNDA.n1118 GNDA.n1048 3.4105
R10335 GNDA.n1076 GNDA.n1048 3.4105
R10336 GNDA.n1120 GNDA.n1048 3.4105
R10337 GNDA.n2689 GNDA.n1048 3.4105
R10338 GNDA.n2691 GNDA.n1048 3.4105
R10339 GNDA.n2693 GNDA.n1068 3.4105
R10340 GNDA.n1090 GNDA.n1068 3.4105
R10341 GNDA.n1092 GNDA.n1068 3.4105
R10342 GNDA.n1089 GNDA.n1068 3.4105
R10343 GNDA.n1094 GNDA.n1068 3.4105
R10344 GNDA.n1088 GNDA.n1068 3.4105
R10345 GNDA.n1096 GNDA.n1068 3.4105
R10346 GNDA.n1087 GNDA.n1068 3.4105
R10347 GNDA.n1098 GNDA.n1068 3.4105
R10348 GNDA.n1086 GNDA.n1068 3.4105
R10349 GNDA.n1100 GNDA.n1068 3.4105
R10350 GNDA.n1085 GNDA.n1068 3.4105
R10351 GNDA.n1102 GNDA.n1068 3.4105
R10352 GNDA.n1084 GNDA.n1068 3.4105
R10353 GNDA.n1104 GNDA.n1068 3.4105
R10354 GNDA.n1083 GNDA.n1068 3.4105
R10355 GNDA.n1106 GNDA.n1068 3.4105
R10356 GNDA.n1082 GNDA.n1068 3.4105
R10357 GNDA.n1108 GNDA.n1068 3.4105
R10358 GNDA.n1081 GNDA.n1068 3.4105
R10359 GNDA.n1110 GNDA.n1068 3.4105
R10360 GNDA.n1080 GNDA.n1068 3.4105
R10361 GNDA.n1112 GNDA.n1068 3.4105
R10362 GNDA.n1079 GNDA.n1068 3.4105
R10363 GNDA.n1114 GNDA.n1068 3.4105
R10364 GNDA.n1078 GNDA.n1068 3.4105
R10365 GNDA.n1116 GNDA.n1068 3.4105
R10366 GNDA.n1077 GNDA.n1068 3.4105
R10367 GNDA.n1118 GNDA.n1068 3.4105
R10368 GNDA.n1076 GNDA.n1068 3.4105
R10369 GNDA.n1120 GNDA.n1068 3.4105
R10370 GNDA.n2689 GNDA.n1068 3.4105
R10371 GNDA.n2691 GNDA.n1068 3.4105
R10372 GNDA.n2693 GNDA.n1047 3.4105
R10373 GNDA.n1090 GNDA.n1047 3.4105
R10374 GNDA.n1092 GNDA.n1047 3.4105
R10375 GNDA.n1089 GNDA.n1047 3.4105
R10376 GNDA.n1094 GNDA.n1047 3.4105
R10377 GNDA.n1088 GNDA.n1047 3.4105
R10378 GNDA.n1096 GNDA.n1047 3.4105
R10379 GNDA.n1087 GNDA.n1047 3.4105
R10380 GNDA.n1098 GNDA.n1047 3.4105
R10381 GNDA.n1086 GNDA.n1047 3.4105
R10382 GNDA.n1100 GNDA.n1047 3.4105
R10383 GNDA.n1085 GNDA.n1047 3.4105
R10384 GNDA.n1102 GNDA.n1047 3.4105
R10385 GNDA.n1084 GNDA.n1047 3.4105
R10386 GNDA.n1104 GNDA.n1047 3.4105
R10387 GNDA.n1083 GNDA.n1047 3.4105
R10388 GNDA.n1106 GNDA.n1047 3.4105
R10389 GNDA.n1082 GNDA.n1047 3.4105
R10390 GNDA.n1108 GNDA.n1047 3.4105
R10391 GNDA.n1081 GNDA.n1047 3.4105
R10392 GNDA.n1110 GNDA.n1047 3.4105
R10393 GNDA.n1080 GNDA.n1047 3.4105
R10394 GNDA.n1112 GNDA.n1047 3.4105
R10395 GNDA.n1079 GNDA.n1047 3.4105
R10396 GNDA.n1114 GNDA.n1047 3.4105
R10397 GNDA.n1078 GNDA.n1047 3.4105
R10398 GNDA.n1116 GNDA.n1047 3.4105
R10399 GNDA.n1077 GNDA.n1047 3.4105
R10400 GNDA.n1118 GNDA.n1047 3.4105
R10401 GNDA.n1076 GNDA.n1047 3.4105
R10402 GNDA.n1120 GNDA.n1047 3.4105
R10403 GNDA.n2689 GNDA.n1047 3.4105
R10404 GNDA.n2691 GNDA.n1047 3.4105
R10405 GNDA.n2693 GNDA.n1069 3.4105
R10406 GNDA.n1090 GNDA.n1069 3.4105
R10407 GNDA.n1092 GNDA.n1069 3.4105
R10408 GNDA.n1089 GNDA.n1069 3.4105
R10409 GNDA.n1094 GNDA.n1069 3.4105
R10410 GNDA.n1088 GNDA.n1069 3.4105
R10411 GNDA.n1096 GNDA.n1069 3.4105
R10412 GNDA.n1087 GNDA.n1069 3.4105
R10413 GNDA.n1098 GNDA.n1069 3.4105
R10414 GNDA.n1086 GNDA.n1069 3.4105
R10415 GNDA.n1100 GNDA.n1069 3.4105
R10416 GNDA.n1085 GNDA.n1069 3.4105
R10417 GNDA.n1102 GNDA.n1069 3.4105
R10418 GNDA.n1084 GNDA.n1069 3.4105
R10419 GNDA.n1104 GNDA.n1069 3.4105
R10420 GNDA.n1083 GNDA.n1069 3.4105
R10421 GNDA.n1106 GNDA.n1069 3.4105
R10422 GNDA.n1082 GNDA.n1069 3.4105
R10423 GNDA.n1108 GNDA.n1069 3.4105
R10424 GNDA.n1081 GNDA.n1069 3.4105
R10425 GNDA.n1110 GNDA.n1069 3.4105
R10426 GNDA.n1080 GNDA.n1069 3.4105
R10427 GNDA.n1112 GNDA.n1069 3.4105
R10428 GNDA.n1079 GNDA.n1069 3.4105
R10429 GNDA.n1114 GNDA.n1069 3.4105
R10430 GNDA.n1078 GNDA.n1069 3.4105
R10431 GNDA.n1116 GNDA.n1069 3.4105
R10432 GNDA.n1077 GNDA.n1069 3.4105
R10433 GNDA.n1118 GNDA.n1069 3.4105
R10434 GNDA.n1076 GNDA.n1069 3.4105
R10435 GNDA.n1120 GNDA.n1069 3.4105
R10436 GNDA.n2689 GNDA.n1069 3.4105
R10437 GNDA.n2691 GNDA.n1069 3.4105
R10438 GNDA.n2693 GNDA.n1046 3.4105
R10439 GNDA.n1090 GNDA.n1046 3.4105
R10440 GNDA.n1092 GNDA.n1046 3.4105
R10441 GNDA.n1089 GNDA.n1046 3.4105
R10442 GNDA.n1094 GNDA.n1046 3.4105
R10443 GNDA.n1088 GNDA.n1046 3.4105
R10444 GNDA.n1096 GNDA.n1046 3.4105
R10445 GNDA.n1087 GNDA.n1046 3.4105
R10446 GNDA.n1098 GNDA.n1046 3.4105
R10447 GNDA.n1086 GNDA.n1046 3.4105
R10448 GNDA.n1100 GNDA.n1046 3.4105
R10449 GNDA.n1085 GNDA.n1046 3.4105
R10450 GNDA.n1102 GNDA.n1046 3.4105
R10451 GNDA.n1084 GNDA.n1046 3.4105
R10452 GNDA.n1104 GNDA.n1046 3.4105
R10453 GNDA.n1083 GNDA.n1046 3.4105
R10454 GNDA.n1106 GNDA.n1046 3.4105
R10455 GNDA.n1082 GNDA.n1046 3.4105
R10456 GNDA.n1108 GNDA.n1046 3.4105
R10457 GNDA.n1081 GNDA.n1046 3.4105
R10458 GNDA.n1110 GNDA.n1046 3.4105
R10459 GNDA.n1080 GNDA.n1046 3.4105
R10460 GNDA.n1112 GNDA.n1046 3.4105
R10461 GNDA.n1079 GNDA.n1046 3.4105
R10462 GNDA.n1114 GNDA.n1046 3.4105
R10463 GNDA.n1078 GNDA.n1046 3.4105
R10464 GNDA.n1116 GNDA.n1046 3.4105
R10465 GNDA.n1077 GNDA.n1046 3.4105
R10466 GNDA.n1118 GNDA.n1046 3.4105
R10467 GNDA.n1076 GNDA.n1046 3.4105
R10468 GNDA.n1120 GNDA.n1046 3.4105
R10469 GNDA.n2689 GNDA.n1046 3.4105
R10470 GNDA.n2691 GNDA.n1046 3.4105
R10471 GNDA.n2693 GNDA.n1070 3.4105
R10472 GNDA.n1090 GNDA.n1070 3.4105
R10473 GNDA.n1092 GNDA.n1070 3.4105
R10474 GNDA.n1089 GNDA.n1070 3.4105
R10475 GNDA.n1094 GNDA.n1070 3.4105
R10476 GNDA.n1088 GNDA.n1070 3.4105
R10477 GNDA.n1096 GNDA.n1070 3.4105
R10478 GNDA.n1087 GNDA.n1070 3.4105
R10479 GNDA.n1098 GNDA.n1070 3.4105
R10480 GNDA.n1086 GNDA.n1070 3.4105
R10481 GNDA.n1100 GNDA.n1070 3.4105
R10482 GNDA.n1085 GNDA.n1070 3.4105
R10483 GNDA.n1102 GNDA.n1070 3.4105
R10484 GNDA.n1084 GNDA.n1070 3.4105
R10485 GNDA.n1104 GNDA.n1070 3.4105
R10486 GNDA.n1083 GNDA.n1070 3.4105
R10487 GNDA.n1106 GNDA.n1070 3.4105
R10488 GNDA.n1082 GNDA.n1070 3.4105
R10489 GNDA.n1108 GNDA.n1070 3.4105
R10490 GNDA.n1081 GNDA.n1070 3.4105
R10491 GNDA.n1110 GNDA.n1070 3.4105
R10492 GNDA.n1080 GNDA.n1070 3.4105
R10493 GNDA.n1112 GNDA.n1070 3.4105
R10494 GNDA.n1079 GNDA.n1070 3.4105
R10495 GNDA.n1114 GNDA.n1070 3.4105
R10496 GNDA.n1078 GNDA.n1070 3.4105
R10497 GNDA.n1116 GNDA.n1070 3.4105
R10498 GNDA.n1077 GNDA.n1070 3.4105
R10499 GNDA.n1118 GNDA.n1070 3.4105
R10500 GNDA.n1076 GNDA.n1070 3.4105
R10501 GNDA.n1120 GNDA.n1070 3.4105
R10502 GNDA.n2689 GNDA.n1070 3.4105
R10503 GNDA.n2691 GNDA.n1070 3.4105
R10504 GNDA.n2693 GNDA.n1045 3.4105
R10505 GNDA.n1090 GNDA.n1045 3.4105
R10506 GNDA.n1092 GNDA.n1045 3.4105
R10507 GNDA.n1089 GNDA.n1045 3.4105
R10508 GNDA.n1094 GNDA.n1045 3.4105
R10509 GNDA.n1088 GNDA.n1045 3.4105
R10510 GNDA.n1096 GNDA.n1045 3.4105
R10511 GNDA.n1087 GNDA.n1045 3.4105
R10512 GNDA.n1098 GNDA.n1045 3.4105
R10513 GNDA.n1086 GNDA.n1045 3.4105
R10514 GNDA.n1100 GNDA.n1045 3.4105
R10515 GNDA.n1085 GNDA.n1045 3.4105
R10516 GNDA.n1102 GNDA.n1045 3.4105
R10517 GNDA.n1084 GNDA.n1045 3.4105
R10518 GNDA.n1104 GNDA.n1045 3.4105
R10519 GNDA.n1083 GNDA.n1045 3.4105
R10520 GNDA.n1106 GNDA.n1045 3.4105
R10521 GNDA.n1082 GNDA.n1045 3.4105
R10522 GNDA.n1108 GNDA.n1045 3.4105
R10523 GNDA.n1081 GNDA.n1045 3.4105
R10524 GNDA.n1110 GNDA.n1045 3.4105
R10525 GNDA.n1080 GNDA.n1045 3.4105
R10526 GNDA.n1112 GNDA.n1045 3.4105
R10527 GNDA.n1079 GNDA.n1045 3.4105
R10528 GNDA.n1114 GNDA.n1045 3.4105
R10529 GNDA.n1078 GNDA.n1045 3.4105
R10530 GNDA.n1116 GNDA.n1045 3.4105
R10531 GNDA.n1077 GNDA.n1045 3.4105
R10532 GNDA.n1118 GNDA.n1045 3.4105
R10533 GNDA.n1076 GNDA.n1045 3.4105
R10534 GNDA.n1120 GNDA.n1045 3.4105
R10535 GNDA.n2689 GNDA.n1045 3.4105
R10536 GNDA.n2691 GNDA.n1045 3.4105
R10537 GNDA.n2693 GNDA.n1071 3.4105
R10538 GNDA.n1090 GNDA.n1071 3.4105
R10539 GNDA.n1092 GNDA.n1071 3.4105
R10540 GNDA.n1089 GNDA.n1071 3.4105
R10541 GNDA.n1094 GNDA.n1071 3.4105
R10542 GNDA.n1088 GNDA.n1071 3.4105
R10543 GNDA.n1096 GNDA.n1071 3.4105
R10544 GNDA.n1087 GNDA.n1071 3.4105
R10545 GNDA.n1098 GNDA.n1071 3.4105
R10546 GNDA.n1086 GNDA.n1071 3.4105
R10547 GNDA.n1100 GNDA.n1071 3.4105
R10548 GNDA.n1085 GNDA.n1071 3.4105
R10549 GNDA.n1102 GNDA.n1071 3.4105
R10550 GNDA.n1084 GNDA.n1071 3.4105
R10551 GNDA.n1104 GNDA.n1071 3.4105
R10552 GNDA.n1083 GNDA.n1071 3.4105
R10553 GNDA.n1106 GNDA.n1071 3.4105
R10554 GNDA.n1082 GNDA.n1071 3.4105
R10555 GNDA.n1108 GNDA.n1071 3.4105
R10556 GNDA.n1081 GNDA.n1071 3.4105
R10557 GNDA.n1110 GNDA.n1071 3.4105
R10558 GNDA.n1080 GNDA.n1071 3.4105
R10559 GNDA.n1112 GNDA.n1071 3.4105
R10560 GNDA.n1079 GNDA.n1071 3.4105
R10561 GNDA.n1114 GNDA.n1071 3.4105
R10562 GNDA.n1078 GNDA.n1071 3.4105
R10563 GNDA.n1116 GNDA.n1071 3.4105
R10564 GNDA.n1077 GNDA.n1071 3.4105
R10565 GNDA.n1118 GNDA.n1071 3.4105
R10566 GNDA.n1076 GNDA.n1071 3.4105
R10567 GNDA.n1120 GNDA.n1071 3.4105
R10568 GNDA.n2689 GNDA.n1071 3.4105
R10569 GNDA.n2691 GNDA.n1071 3.4105
R10570 GNDA.n2693 GNDA.n1044 3.4105
R10571 GNDA.n1090 GNDA.n1044 3.4105
R10572 GNDA.n1092 GNDA.n1044 3.4105
R10573 GNDA.n1089 GNDA.n1044 3.4105
R10574 GNDA.n1094 GNDA.n1044 3.4105
R10575 GNDA.n1088 GNDA.n1044 3.4105
R10576 GNDA.n1096 GNDA.n1044 3.4105
R10577 GNDA.n1087 GNDA.n1044 3.4105
R10578 GNDA.n1098 GNDA.n1044 3.4105
R10579 GNDA.n1086 GNDA.n1044 3.4105
R10580 GNDA.n1100 GNDA.n1044 3.4105
R10581 GNDA.n1085 GNDA.n1044 3.4105
R10582 GNDA.n1102 GNDA.n1044 3.4105
R10583 GNDA.n1084 GNDA.n1044 3.4105
R10584 GNDA.n1104 GNDA.n1044 3.4105
R10585 GNDA.n1083 GNDA.n1044 3.4105
R10586 GNDA.n1106 GNDA.n1044 3.4105
R10587 GNDA.n1082 GNDA.n1044 3.4105
R10588 GNDA.n1108 GNDA.n1044 3.4105
R10589 GNDA.n1081 GNDA.n1044 3.4105
R10590 GNDA.n1110 GNDA.n1044 3.4105
R10591 GNDA.n1080 GNDA.n1044 3.4105
R10592 GNDA.n1112 GNDA.n1044 3.4105
R10593 GNDA.n1079 GNDA.n1044 3.4105
R10594 GNDA.n1114 GNDA.n1044 3.4105
R10595 GNDA.n1078 GNDA.n1044 3.4105
R10596 GNDA.n1116 GNDA.n1044 3.4105
R10597 GNDA.n1077 GNDA.n1044 3.4105
R10598 GNDA.n1118 GNDA.n1044 3.4105
R10599 GNDA.n1076 GNDA.n1044 3.4105
R10600 GNDA.n1120 GNDA.n1044 3.4105
R10601 GNDA.n2689 GNDA.n1044 3.4105
R10602 GNDA.n2691 GNDA.n1044 3.4105
R10603 GNDA.n2693 GNDA.n1072 3.4105
R10604 GNDA.n1090 GNDA.n1072 3.4105
R10605 GNDA.n1092 GNDA.n1072 3.4105
R10606 GNDA.n1089 GNDA.n1072 3.4105
R10607 GNDA.n1094 GNDA.n1072 3.4105
R10608 GNDA.n1088 GNDA.n1072 3.4105
R10609 GNDA.n1096 GNDA.n1072 3.4105
R10610 GNDA.n1087 GNDA.n1072 3.4105
R10611 GNDA.n1098 GNDA.n1072 3.4105
R10612 GNDA.n1086 GNDA.n1072 3.4105
R10613 GNDA.n1100 GNDA.n1072 3.4105
R10614 GNDA.n1085 GNDA.n1072 3.4105
R10615 GNDA.n1102 GNDA.n1072 3.4105
R10616 GNDA.n1084 GNDA.n1072 3.4105
R10617 GNDA.n1104 GNDA.n1072 3.4105
R10618 GNDA.n1083 GNDA.n1072 3.4105
R10619 GNDA.n1106 GNDA.n1072 3.4105
R10620 GNDA.n1082 GNDA.n1072 3.4105
R10621 GNDA.n1108 GNDA.n1072 3.4105
R10622 GNDA.n1081 GNDA.n1072 3.4105
R10623 GNDA.n1110 GNDA.n1072 3.4105
R10624 GNDA.n1080 GNDA.n1072 3.4105
R10625 GNDA.n1112 GNDA.n1072 3.4105
R10626 GNDA.n1079 GNDA.n1072 3.4105
R10627 GNDA.n1114 GNDA.n1072 3.4105
R10628 GNDA.n1078 GNDA.n1072 3.4105
R10629 GNDA.n1116 GNDA.n1072 3.4105
R10630 GNDA.n1077 GNDA.n1072 3.4105
R10631 GNDA.n1118 GNDA.n1072 3.4105
R10632 GNDA.n1076 GNDA.n1072 3.4105
R10633 GNDA.n1120 GNDA.n1072 3.4105
R10634 GNDA.n2689 GNDA.n1072 3.4105
R10635 GNDA.n2691 GNDA.n1072 3.4105
R10636 GNDA.n2693 GNDA.n1043 3.4105
R10637 GNDA.n1090 GNDA.n1043 3.4105
R10638 GNDA.n1092 GNDA.n1043 3.4105
R10639 GNDA.n1089 GNDA.n1043 3.4105
R10640 GNDA.n1094 GNDA.n1043 3.4105
R10641 GNDA.n1088 GNDA.n1043 3.4105
R10642 GNDA.n1096 GNDA.n1043 3.4105
R10643 GNDA.n1087 GNDA.n1043 3.4105
R10644 GNDA.n1098 GNDA.n1043 3.4105
R10645 GNDA.n1086 GNDA.n1043 3.4105
R10646 GNDA.n1100 GNDA.n1043 3.4105
R10647 GNDA.n1085 GNDA.n1043 3.4105
R10648 GNDA.n1102 GNDA.n1043 3.4105
R10649 GNDA.n1084 GNDA.n1043 3.4105
R10650 GNDA.n1104 GNDA.n1043 3.4105
R10651 GNDA.n1083 GNDA.n1043 3.4105
R10652 GNDA.n1106 GNDA.n1043 3.4105
R10653 GNDA.n1082 GNDA.n1043 3.4105
R10654 GNDA.n1108 GNDA.n1043 3.4105
R10655 GNDA.n1081 GNDA.n1043 3.4105
R10656 GNDA.n1110 GNDA.n1043 3.4105
R10657 GNDA.n1080 GNDA.n1043 3.4105
R10658 GNDA.n1112 GNDA.n1043 3.4105
R10659 GNDA.n1079 GNDA.n1043 3.4105
R10660 GNDA.n1114 GNDA.n1043 3.4105
R10661 GNDA.n1078 GNDA.n1043 3.4105
R10662 GNDA.n1116 GNDA.n1043 3.4105
R10663 GNDA.n1077 GNDA.n1043 3.4105
R10664 GNDA.n1118 GNDA.n1043 3.4105
R10665 GNDA.n1076 GNDA.n1043 3.4105
R10666 GNDA.n1120 GNDA.n1043 3.4105
R10667 GNDA.n2689 GNDA.n1043 3.4105
R10668 GNDA.n2691 GNDA.n1043 3.4105
R10669 GNDA.n2693 GNDA.n1073 3.4105
R10670 GNDA.n1090 GNDA.n1073 3.4105
R10671 GNDA.n1092 GNDA.n1073 3.4105
R10672 GNDA.n1089 GNDA.n1073 3.4105
R10673 GNDA.n1094 GNDA.n1073 3.4105
R10674 GNDA.n1088 GNDA.n1073 3.4105
R10675 GNDA.n1096 GNDA.n1073 3.4105
R10676 GNDA.n1087 GNDA.n1073 3.4105
R10677 GNDA.n1098 GNDA.n1073 3.4105
R10678 GNDA.n1086 GNDA.n1073 3.4105
R10679 GNDA.n1100 GNDA.n1073 3.4105
R10680 GNDA.n1085 GNDA.n1073 3.4105
R10681 GNDA.n1102 GNDA.n1073 3.4105
R10682 GNDA.n1084 GNDA.n1073 3.4105
R10683 GNDA.n1104 GNDA.n1073 3.4105
R10684 GNDA.n1083 GNDA.n1073 3.4105
R10685 GNDA.n1106 GNDA.n1073 3.4105
R10686 GNDA.n1082 GNDA.n1073 3.4105
R10687 GNDA.n1108 GNDA.n1073 3.4105
R10688 GNDA.n1081 GNDA.n1073 3.4105
R10689 GNDA.n1110 GNDA.n1073 3.4105
R10690 GNDA.n1080 GNDA.n1073 3.4105
R10691 GNDA.n1112 GNDA.n1073 3.4105
R10692 GNDA.n1079 GNDA.n1073 3.4105
R10693 GNDA.n1114 GNDA.n1073 3.4105
R10694 GNDA.n1078 GNDA.n1073 3.4105
R10695 GNDA.n1116 GNDA.n1073 3.4105
R10696 GNDA.n1077 GNDA.n1073 3.4105
R10697 GNDA.n1118 GNDA.n1073 3.4105
R10698 GNDA.n1076 GNDA.n1073 3.4105
R10699 GNDA.n1120 GNDA.n1073 3.4105
R10700 GNDA.n2689 GNDA.n1073 3.4105
R10701 GNDA.n2691 GNDA.n1073 3.4105
R10702 GNDA.n2693 GNDA.n1042 3.4105
R10703 GNDA.n1090 GNDA.n1042 3.4105
R10704 GNDA.n1092 GNDA.n1042 3.4105
R10705 GNDA.n1089 GNDA.n1042 3.4105
R10706 GNDA.n1094 GNDA.n1042 3.4105
R10707 GNDA.n1088 GNDA.n1042 3.4105
R10708 GNDA.n1096 GNDA.n1042 3.4105
R10709 GNDA.n1087 GNDA.n1042 3.4105
R10710 GNDA.n1098 GNDA.n1042 3.4105
R10711 GNDA.n1086 GNDA.n1042 3.4105
R10712 GNDA.n1100 GNDA.n1042 3.4105
R10713 GNDA.n1085 GNDA.n1042 3.4105
R10714 GNDA.n1102 GNDA.n1042 3.4105
R10715 GNDA.n1084 GNDA.n1042 3.4105
R10716 GNDA.n1104 GNDA.n1042 3.4105
R10717 GNDA.n1083 GNDA.n1042 3.4105
R10718 GNDA.n1106 GNDA.n1042 3.4105
R10719 GNDA.n1082 GNDA.n1042 3.4105
R10720 GNDA.n1108 GNDA.n1042 3.4105
R10721 GNDA.n1081 GNDA.n1042 3.4105
R10722 GNDA.n1110 GNDA.n1042 3.4105
R10723 GNDA.n1080 GNDA.n1042 3.4105
R10724 GNDA.n1112 GNDA.n1042 3.4105
R10725 GNDA.n1079 GNDA.n1042 3.4105
R10726 GNDA.n1114 GNDA.n1042 3.4105
R10727 GNDA.n1078 GNDA.n1042 3.4105
R10728 GNDA.n1116 GNDA.n1042 3.4105
R10729 GNDA.n1077 GNDA.n1042 3.4105
R10730 GNDA.n1118 GNDA.n1042 3.4105
R10731 GNDA.n1076 GNDA.n1042 3.4105
R10732 GNDA.n1120 GNDA.n1042 3.4105
R10733 GNDA.n2689 GNDA.n1042 3.4105
R10734 GNDA.n2691 GNDA.n1042 3.4105
R10735 GNDA.n2693 GNDA.n1074 3.4105
R10736 GNDA.n1090 GNDA.n1074 3.4105
R10737 GNDA.n1092 GNDA.n1074 3.4105
R10738 GNDA.n1089 GNDA.n1074 3.4105
R10739 GNDA.n1094 GNDA.n1074 3.4105
R10740 GNDA.n1088 GNDA.n1074 3.4105
R10741 GNDA.n1096 GNDA.n1074 3.4105
R10742 GNDA.n1087 GNDA.n1074 3.4105
R10743 GNDA.n1098 GNDA.n1074 3.4105
R10744 GNDA.n1086 GNDA.n1074 3.4105
R10745 GNDA.n1100 GNDA.n1074 3.4105
R10746 GNDA.n1085 GNDA.n1074 3.4105
R10747 GNDA.n1102 GNDA.n1074 3.4105
R10748 GNDA.n1084 GNDA.n1074 3.4105
R10749 GNDA.n1104 GNDA.n1074 3.4105
R10750 GNDA.n1083 GNDA.n1074 3.4105
R10751 GNDA.n1106 GNDA.n1074 3.4105
R10752 GNDA.n1082 GNDA.n1074 3.4105
R10753 GNDA.n1108 GNDA.n1074 3.4105
R10754 GNDA.n1081 GNDA.n1074 3.4105
R10755 GNDA.n1110 GNDA.n1074 3.4105
R10756 GNDA.n1080 GNDA.n1074 3.4105
R10757 GNDA.n1112 GNDA.n1074 3.4105
R10758 GNDA.n1079 GNDA.n1074 3.4105
R10759 GNDA.n1114 GNDA.n1074 3.4105
R10760 GNDA.n1078 GNDA.n1074 3.4105
R10761 GNDA.n1116 GNDA.n1074 3.4105
R10762 GNDA.n1077 GNDA.n1074 3.4105
R10763 GNDA.n1118 GNDA.n1074 3.4105
R10764 GNDA.n1076 GNDA.n1074 3.4105
R10765 GNDA.n1120 GNDA.n1074 3.4105
R10766 GNDA.n2689 GNDA.n1074 3.4105
R10767 GNDA.n2691 GNDA.n1074 3.4105
R10768 GNDA.n2693 GNDA.n1041 3.4105
R10769 GNDA.n1090 GNDA.n1041 3.4105
R10770 GNDA.n1092 GNDA.n1041 3.4105
R10771 GNDA.n1089 GNDA.n1041 3.4105
R10772 GNDA.n1094 GNDA.n1041 3.4105
R10773 GNDA.n1088 GNDA.n1041 3.4105
R10774 GNDA.n1096 GNDA.n1041 3.4105
R10775 GNDA.n1087 GNDA.n1041 3.4105
R10776 GNDA.n1098 GNDA.n1041 3.4105
R10777 GNDA.n1086 GNDA.n1041 3.4105
R10778 GNDA.n1100 GNDA.n1041 3.4105
R10779 GNDA.n1085 GNDA.n1041 3.4105
R10780 GNDA.n1102 GNDA.n1041 3.4105
R10781 GNDA.n1084 GNDA.n1041 3.4105
R10782 GNDA.n1104 GNDA.n1041 3.4105
R10783 GNDA.n1083 GNDA.n1041 3.4105
R10784 GNDA.n1106 GNDA.n1041 3.4105
R10785 GNDA.n1082 GNDA.n1041 3.4105
R10786 GNDA.n1108 GNDA.n1041 3.4105
R10787 GNDA.n1081 GNDA.n1041 3.4105
R10788 GNDA.n1110 GNDA.n1041 3.4105
R10789 GNDA.n1080 GNDA.n1041 3.4105
R10790 GNDA.n1112 GNDA.n1041 3.4105
R10791 GNDA.n1079 GNDA.n1041 3.4105
R10792 GNDA.n1114 GNDA.n1041 3.4105
R10793 GNDA.n1078 GNDA.n1041 3.4105
R10794 GNDA.n1116 GNDA.n1041 3.4105
R10795 GNDA.n1077 GNDA.n1041 3.4105
R10796 GNDA.n1118 GNDA.n1041 3.4105
R10797 GNDA.n1076 GNDA.n1041 3.4105
R10798 GNDA.n1120 GNDA.n1041 3.4105
R10799 GNDA.n2689 GNDA.n1041 3.4105
R10800 GNDA.n2691 GNDA.n1041 3.4105
R10801 GNDA.n2693 GNDA.n2692 3.4105
R10802 GNDA.n2692 GNDA.n1090 3.4105
R10803 GNDA.n2692 GNDA.n1092 3.4105
R10804 GNDA.n2692 GNDA.n1089 3.4105
R10805 GNDA.n2692 GNDA.n1094 3.4105
R10806 GNDA.n2692 GNDA.n1088 3.4105
R10807 GNDA.n2692 GNDA.n1096 3.4105
R10808 GNDA.n2692 GNDA.n1087 3.4105
R10809 GNDA.n2692 GNDA.n1098 3.4105
R10810 GNDA.n2692 GNDA.n1086 3.4105
R10811 GNDA.n2692 GNDA.n1100 3.4105
R10812 GNDA.n2692 GNDA.n1085 3.4105
R10813 GNDA.n2692 GNDA.n1102 3.4105
R10814 GNDA.n2692 GNDA.n1084 3.4105
R10815 GNDA.n2692 GNDA.n1104 3.4105
R10816 GNDA.n2692 GNDA.n1083 3.4105
R10817 GNDA.n2692 GNDA.n1106 3.4105
R10818 GNDA.n2692 GNDA.n1082 3.4105
R10819 GNDA.n2692 GNDA.n1108 3.4105
R10820 GNDA.n2692 GNDA.n1081 3.4105
R10821 GNDA.n2692 GNDA.n1110 3.4105
R10822 GNDA.n2692 GNDA.n1080 3.4105
R10823 GNDA.n2692 GNDA.n1112 3.4105
R10824 GNDA.n2692 GNDA.n1079 3.4105
R10825 GNDA.n2692 GNDA.n1114 3.4105
R10826 GNDA.n2692 GNDA.n1078 3.4105
R10827 GNDA.n2692 GNDA.n1116 3.4105
R10828 GNDA.n2692 GNDA.n1077 3.4105
R10829 GNDA.n2692 GNDA.n1118 3.4105
R10830 GNDA.n2692 GNDA.n1076 3.4105
R10831 GNDA.n2692 GNDA.n1120 3.4105
R10832 GNDA.n2692 GNDA.n2691 3.4105
R10833 GNDA.n1204 GNDA.n1155 3.4105
R10834 GNDA.n1204 GNDA.n1172 3.4105
R10835 GNDA.n2654 GNDA.n1204 3.4105
R10836 GNDA.n2606 GNDA.n1157 3.4105
R10837 GNDA.n2606 GNDA.n1154 3.4105
R10838 GNDA.n2606 GNDA.n1158 3.4105
R10839 GNDA.n2606 GNDA.n1153 3.4105
R10840 GNDA.n2606 GNDA.n1159 3.4105
R10841 GNDA.n2606 GNDA.n1152 3.4105
R10842 GNDA.n2606 GNDA.n1160 3.4105
R10843 GNDA.n2606 GNDA.n1151 3.4105
R10844 GNDA.n2606 GNDA.n1161 3.4105
R10845 GNDA.n2606 GNDA.n1150 3.4105
R10846 GNDA.n2606 GNDA.n1162 3.4105
R10847 GNDA.n2606 GNDA.n1149 3.4105
R10848 GNDA.n2606 GNDA.n1163 3.4105
R10849 GNDA.n2606 GNDA.n1148 3.4105
R10850 GNDA.n2606 GNDA.n1164 3.4105
R10851 GNDA.n2606 GNDA.n1147 3.4105
R10852 GNDA.n2606 GNDA.n1165 3.4105
R10853 GNDA.n2606 GNDA.n1146 3.4105
R10854 GNDA.n2606 GNDA.n1166 3.4105
R10855 GNDA.n2606 GNDA.n1145 3.4105
R10856 GNDA.n2606 GNDA.n1167 3.4105
R10857 GNDA.n2606 GNDA.n1144 3.4105
R10858 GNDA.n2606 GNDA.n1168 3.4105
R10859 GNDA.n2606 GNDA.n1143 3.4105
R10860 GNDA.n2606 GNDA.n1169 3.4105
R10861 GNDA.n2606 GNDA.n1142 3.4105
R10862 GNDA.n2606 GNDA.n1170 3.4105
R10863 GNDA.n2606 GNDA.n1141 3.4105
R10864 GNDA.n2606 GNDA.n1171 3.4105
R10865 GNDA.n2606 GNDA.n1172 3.4105
R10866 GNDA.n2654 GNDA.n2606 3.4105
R10867 GNDA.n1188 GNDA.n1156 3.4105
R10868 GNDA.n1188 GNDA.n1155 3.4105
R10869 GNDA.n1188 GNDA.n1157 3.4105
R10870 GNDA.n1188 GNDA.n1154 3.4105
R10871 GNDA.n1188 GNDA.n1158 3.4105
R10872 GNDA.n1188 GNDA.n1153 3.4105
R10873 GNDA.n1188 GNDA.n1159 3.4105
R10874 GNDA.n1188 GNDA.n1152 3.4105
R10875 GNDA.n1188 GNDA.n1160 3.4105
R10876 GNDA.n1188 GNDA.n1151 3.4105
R10877 GNDA.n1188 GNDA.n1161 3.4105
R10878 GNDA.n1188 GNDA.n1150 3.4105
R10879 GNDA.n1188 GNDA.n1162 3.4105
R10880 GNDA.n1188 GNDA.n1149 3.4105
R10881 GNDA.n1188 GNDA.n1163 3.4105
R10882 GNDA.n1188 GNDA.n1148 3.4105
R10883 GNDA.n1188 GNDA.n1164 3.4105
R10884 GNDA.n1188 GNDA.n1147 3.4105
R10885 GNDA.n1188 GNDA.n1165 3.4105
R10886 GNDA.n1188 GNDA.n1146 3.4105
R10887 GNDA.n1188 GNDA.n1166 3.4105
R10888 GNDA.n1188 GNDA.n1145 3.4105
R10889 GNDA.n1188 GNDA.n1167 3.4105
R10890 GNDA.n1188 GNDA.n1144 3.4105
R10891 GNDA.n1188 GNDA.n1168 3.4105
R10892 GNDA.n1188 GNDA.n1143 3.4105
R10893 GNDA.n1188 GNDA.n1169 3.4105
R10894 GNDA.n1188 GNDA.n1142 3.4105
R10895 GNDA.n1188 GNDA.n1170 3.4105
R10896 GNDA.n1188 GNDA.n1141 3.4105
R10897 GNDA.n1188 GNDA.n1171 3.4105
R10898 GNDA.n1188 GNDA.n1172 3.4105
R10899 GNDA.n2654 GNDA.n1188 3.4105
R10900 GNDA.n2608 GNDA.n1156 3.4105
R10901 GNDA.n2608 GNDA.n1155 3.4105
R10902 GNDA.n2608 GNDA.n1157 3.4105
R10903 GNDA.n2608 GNDA.n1154 3.4105
R10904 GNDA.n2608 GNDA.n1158 3.4105
R10905 GNDA.n2608 GNDA.n1153 3.4105
R10906 GNDA.n2608 GNDA.n1159 3.4105
R10907 GNDA.n2608 GNDA.n1152 3.4105
R10908 GNDA.n2608 GNDA.n1160 3.4105
R10909 GNDA.n2608 GNDA.n1151 3.4105
R10910 GNDA.n2608 GNDA.n1161 3.4105
R10911 GNDA.n2608 GNDA.n1150 3.4105
R10912 GNDA.n2608 GNDA.n1162 3.4105
R10913 GNDA.n2608 GNDA.n1149 3.4105
R10914 GNDA.n2608 GNDA.n1163 3.4105
R10915 GNDA.n2608 GNDA.n1148 3.4105
R10916 GNDA.n2608 GNDA.n1164 3.4105
R10917 GNDA.n2608 GNDA.n1147 3.4105
R10918 GNDA.n2608 GNDA.n1165 3.4105
R10919 GNDA.n2608 GNDA.n1146 3.4105
R10920 GNDA.n2608 GNDA.n1166 3.4105
R10921 GNDA.n2608 GNDA.n1145 3.4105
R10922 GNDA.n2608 GNDA.n1167 3.4105
R10923 GNDA.n2608 GNDA.n1144 3.4105
R10924 GNDA.n2608 GNDA.n1168 3.4105
R10925 GNDA.n2608 GNDA.n1143 3.4105
R10926 GNDA.n2608 GNDA.n1169 3.4105
R10927 GNDA.n2608 GNDA.n1142 3.4105
R10928 GNDA.n2608 GNDA.n1170 3.4105
R10929 GNDA.n2608 GNDA.n1141 3.4105
R10930 GNDA.n2608 GNDA.n1171 3.4105
R10931 GNDA.n2608 GNDA.n1172 3.4105
R10932 GNDA.n2654 GNDA.n2608 3.4105
R10933 GNDA.n1187 GNDA.n1156 3.4105
R10934 GNDA.n1187 GNDA.n1155 3.4105
R10935 GNDA.n1187 GNDA.n1157 3.4105
R10936 GNDA.n1187 GNDA.n1154 3.4105
R10937 GNDA.n1187 GNDA.n1158 3.4105
R10938 GNDA.n1187 GNDA.n1153 3.4105
R10939 GNDA.n1187 GNDA.n1159 3.4105
R10940 GNDA.n1187 GNDA.n1152 3.4105
R10941 GNDA.n1187 GNDA.n1160 3.4105
R10942 GNDA.n1187 GNDA.n1151 3.4105
R10943 GNDA.n1187 GNDA.n1161 3.4105
R10944 GNDA.n1187 GNDA.n1150 3.4105
R10945 GNDA.n1187 GNDA.n1162 3.4105
R10946 GNDA.n1187 GNDA.n1149 3.4105
R10947 GNDA.n1187 GNDA.n1163 3.4105
R10948 GNDA.n1187 GNDA.n1148 3.4105
R10949 GNDA.n1187 GNDA.n1164 3.4105
R10950 GNDA.n1187 GNDA.n1147 3.4105
R10951 GNDA.n1187 GNDA.n1165 3.4105
R10952 GNDA.n1187 GNDA.n1146 3.4105
R10953 GNDA.n1187 GNDA.n1166 3.4105
R10954 GNDA.n1187 GNDA.n1145 3.4105
R10955 GNDA.n1187 GNDA.n1167 3.4105
R10956 GNDA.n1187 GNDA.n1144 3.4105
R10957 GNDA.n1187 GNDA.n1168 3.4105
R10958 GNDA.n1187 GNDA.n1143 3.4105
R10959 GNDA.n1187 GNDA.n1169 3.4105
R10960 GNDA.n1187 GNDA.n1142 3.4105
R10961 GNDA.n1187 GNDA.n1170 3.4105
R10962 GNDA.n1187 GNDA.n1141 3.4105
R10963 GNDA.n1187 GNDA.n1171 3.4105
R10964 GNDA.n1187 GNDA.n1172 3.4105
R10965 GNDA.n2654 GNDA.n1187 3.4105
R10966 GNDA.n2610 GNDA.n1156 3.4105
R10967 GNDA.n2610 GNDA.n1155 3.4105
R10968 GNDA.n2610 GNDA.n1157 3.4105
R10969 GNDA.n2610 GNDA.n1154 3.4105
R10970 GNDA.n2610 GNDA.n1158 3.4105
R10971 GNDA.n2610 GNDA.n1153 3.4105
R10972 GNDA.n2610 GNDA.n1159 3.4105
R10973 GNDA.n2610 GNDA.n1152 3.4105
R10974 GNDA.n2610 GNDA.n1160 3.4105
R10975 GNDA.n2610 GNDA.n1151 3.4105
R10976 GNDA.n2610 GNDA.n1161 3.4105
R10977 GNDA.n2610 GNDA.n1150 3.4105
R10978 GNDA.n2610 GNDA.n1162 3.4105
R10979 GNDA.n2610 GNDA.n1149 3.4105
R10980 GNDA.n2610 GNDA.n1163 3.4105
R10981 GNDA.n2610 GNDA.n1148 3.4105
R10982 GNDA.n2610 GNDA.n1164 3.4105
R10983 GNDA.n2610 GNDA.n1147 3.4105
R10984 GNDA.n2610 GNDA.n1165 3.4105
R10985 GNDA.n2610 GNDA.n1146 3.4105
R10986 GNDA.n2610 GNDA.n1166 3.4105
R10987 GNDA.n2610 GNDA.n1145 3.4105
R10988 GNDA.n2610 GNDA.n1167 3.4105
R10989 GNDA.n2610 GNDA.n1144 3.4105
R10990 GNDA.n2610 GNDA.n1168 3.4105
R10991 GNDA.n2610 GNDA.n1143 3.4105
R10992 GNDA.n2610 GNDA.n1169 3.4105
R10993 GNDA.n2610 GNDA.n1142 3.4105
R10994 GNDA.n2610 GNDA.n1170 3.4105
R10995 GNDA.n2610 GNDA.n1141 3.4105
R10996 GNDA.n2610 GNDA.n1171 3.4105
R10997 GNDA.n2610 GNDA.n1172 3.4105
R10998 GNDA.n2654 GNDA.n2610 3.4105
R10999 GNDA.n1186 GNDA.n1156 3.4105
R11000 GNDA.n1186 GNDA.n1155 3.4105
R11001 GNDA.n1186 GNDA.n1157 3.4105
R11002 GNDA.n1186 GNDA.n1154 3.4105
R11003 GNDA.n1186 GNDA.n1158 3.4105
R11004 GNDA.n1186 GNDA.n1153 3.4105
R11005 GNDA.n1186 GNDA.n1159 3.4105
R11006 GNDA.n1186 GNDA.n1152 3.4105
R11007 GNDA.n1186 GNDA.n1160 3.4105
R11008 GNDA.n1186 GNDA.n1151 3.4105
R11009 GNDA.n1186 GNDA.n1161 3.4105
R11010 GNDA.n1186 GNDA.n1150 3.4105
R11011 GNDA.n1186 GNDA.n1162 3.4105
R11012 GNDA.n1186 GNDA.n1149 3.4105
R11013 GNDA.n1186 GNDA.n1163 3.4105
R11014 GNDA.n1186 GNDA.n1148 3.4105
R11015 GNDA.n1186 GNDA.n1164 3.4105
R11016 GNDA.n1186 GNDA.n1147 3.4105
R11017 GNDA.n1186 GNDA.n1165 3.4105
R11018 GNDA.n1186 GNDA.n1146 3.4105
R11019 GNDA.n1186 GNDA.n1166 3.4105
R11020 GNDA.n1186 GNDA.n1145 3.4105
R11021 GNDA.n1186 GNDA.n1167 3.4105
R11022 GNDA.n1186 GNDA.n1144 3.4105
R11023 GNDA.n1186 GNDA.n1168 3.4105
R11024 GNDA.n1186 GNDA.n1143 3.4105
R11025 GNDA.n1186 GNDA.n1169 3.4105
R11026 GNDA.n1186 GNDA.n1142 3.4105
R11027 GNDA.n1186 GNDA.n1170 3.4105
R11028 GNDA.n1186 GNDA.n1141 3.4105
R11029 GNDA.n1186 GNDA.n1171 3.4105
R11030 GNDA.n1186 GNDA.n1172 3.4105
R11031 GNDA.n2654 GNDA.n1186 3.4105
R11032 GNDA.n2612 GNDA.n1156 3.4105
R11033 GNDA.n2612 GNDA.n1155 3.4105
R11034 GNDA.n2612 GNDA.n1157 3.4105
R11035 GNDA.n2612 GNDA.n1154 3.4105
R11036 GNDA.n2612 GNDA.n1158 3.4105
R11037 GNDA.n2612 GNDA.n1153 3.4105
R11038 GNDA.n2612 GNDA.n1159 3.4105
R11039 GNDA.n2612 GNDA.n1152 3.4105
R11040 GNDA.n2612 GNDA.n1160 3.4105
R11041 GNDA.n2612 GNDA.n1151 3.4105
R11042 GNDA.n2612 GNDA.n1161 3.4105
R11043 GNDA.n2612 GNDA.n1150 3.4105
R11044 GNDA.n2612 GNDA.n1162 3.4105
R11045 GNDA.n2612 GNDA.n1149 3.4105
R11046 GNDA.n2612 GNDA.n1163 3.4105
R11047 GNDA.n2612 GNDA.n1148 3.4105
R11048 GNDA.n2612 GNDA.n1164 3.4105
R11049 GNDA.n2612 GNDA.n1147 3.4105
R11050 GNDA.n2612 GNDA.n1165 3.4105
R11051 GNDA.n2612 GNDA.n1146 3.4105
R11052 GNDA.n2612 GNDA.n1166 3.4105
R11053 GNDA.n2612 GNDA.n1145 3.4105
R11054 GNDA.n2612 GNDA.n1167 3.4105
R11055 GNDA.n2612 GNDA.n1144 3.4105
R11056 GNDA.n2612 GNDA.n1168 3.4105
R11057 GNDA.n2612 GNDA.n1143 3.4105
R11058 GNDA.n2612 GNDA.n1169 3.4105
R11059 GNDA.n2612 GNDA.n1142 3.4105
R11060 GNDA.n2612 GNDA.n1170 3.4105
R11061 GNDA.n2612 GNDA.n1141 3.4105
R11062 GNDA.n2612 GNDA.n1171 3.4105
R11063 GNDA.n2612 GNDA.n1172 3.4105
R11064 GNDA.n2654 GNDA.n2612 3.4105
R11065 GNDA.n1185 GNDA.n1156 3.4105
R11066 GNDA.n1185 GNDA.n1155 3.4105
R11067 GNDA.n1185 GNDA.n1157 3.4105
R11068 GNDA.n1185 GNDA.n1154 3.4105
R11069 GNDA.n1185 GNDA.n1158 3.4105
R11070 GNDA.n1185 GNDA.n1153 3.4105
R11071 GNDA.n1185 GNDA.n1159 3.4105
R11072 GNDA.n1185 GNDA.n1152 3.4105
R11073 GNDA.n1185 GNDA.n1160 3.4105
R11074 GNDA.n1185 GNDA.n1151 3.4105
R11075 GNDA.n1185 GNDA.n1161 3.4105
R11076 GNDA.n1185 GNDA.n1150 3.4105
R11077 GNDA.n1185 GNDA.n1162 3.4105
R11078 GNDA.n1185 GNDA.n1149 3.4105
R11079 GNDA.n1185 GNDA.n1163 3.4105
R11080 GNDA.n1185 GNDA.n1148 3.4105
R11081 GNDA.n1185 GNDA.n1164 3.4105
R11082 GNDA.n1185 GNDA.n1147 3.4105
R11083 GNDA.n1185 GNDA.n1165 3.4105
R11084 GNDA.n1185 GNDA.n1146 3.4105
R11085 GNDA.n1185 GNDA.n1166 3.4105
R11086 GNDA.n1185 GNDA.n1145 3.4105
R11087 GNDA.n1185 GNDA.n1167 3.4105
R11088 GNDA.n1185 GNDA.n1144 3.4105
R11089 GNDA.n1185 GNDA.n1168 3.4105
R11090 GNDA.n1185 GNDA.n1143 3.4105
R11091 GNDA.n1185 GNDA.n1169 3.4105
R11092 GNDA.n1185 GNDA.n1142 3.4105
R11093 GNDA.n1185 GNDA.n1170 3.4105
R11094 GNDA.n1185 GNDA.n1141 3.4105
R11095 GNDA.n1185 GNDA.n1171 3.4105
R11096 GNDA.n1185 GNDA.n1172 3.4105
R11097 GNDA.n2654 GNDA.n1185 3.4105
R11098 GNDA.n2614 GNDA.n1156 3.4105
R11099 GNDA.n2614 GNDA.n1155 3.4105
R11100 GNDA.n2614 GNDA.n1157 3.4105
R11101 GNDA.n2614 GNDA.n1154 3.4105
R11102 GNDA.n2614 GNDA.n1158 3.4105
R11103 GNDA.n2614 GNDA.n1153 3.4105
R11104 GNDA.n2614 GNDA.n1159 3.4105
R11105 GNDA.n2614 GNDA.n1152 3.4105
R11106 GNDA.n2614 GNDA.n1160 3.4105
R11107 GNDA.n2614 GNDA.n1151 3.4105
R11108 GNDA.n2614 GNDA.n1161 3.4105
R11109 GNDA.n2614 GNDA.n1150 3.4105
R11110 GNDA.n2614 GNDA.n1162 3.4105
R11111 GNDA.n2614 GNDA.n1149 3.4105
R11112 GNDA.n2614 GNDA.n1163 3.4105
R11113 GNDA.n2614 GNDA.n1148 3.4105
R11114 GNDA.n2614 GNDA.n1164 3.4105
R11115 GNDA.n2614 GNDA.n1147 3.4105
R11116 GNDA.n2614 GNDA.n1165 3.4105
R11117 GNDA.n2614 GNDA.n1146 3.4105
R11118 GNDA.n2614 GNDA.n1166 3.4105
R11119 GNDA.n2614 GNDA.n1145 3.4105
R11120 GNDA.n2614 GNDA.n1167 3.4105
R11121 GNDA.n2614 GNDA.n1144 3.4105
R11122 GNDA.n2614 GNDA.n1168 3.4105
R11123 GNDA.n2614 GNDA.n1143 3.4105
R11124 GNDA.n2614 GNDA.n1169 3.4105
R11125 GNDA.n2614 GNDA.n1142 3.4105
R11126 GNDA.n2614 GNDA.n1170 3.4105
R11127 GNDA.n2614 GNDA.n1141 3.4105
R11128 GNDA.n2614 GNDA.n1171 3.4105
R11129 GNDA.n2614 GNDA.n1172 3.4105
R11130 GNDA.n2654 GNDA.n2614 3.4105
R11131 GNDA.n1184 GNDA.n1156 3.4105
R11132 GNDA.n1184 GNDA.n1155 3.4105
R11133 GNDA.n1184 GNDA.n1157 3.4105
R11134 GNDA.n1184 GNDA.n1154 3.4105
R11135 GNDA.n1184 GNDA.n1158 3.4105
R11136 GNDA.n1184 GNDA.n1153 3.4105
R11137 GNDA.n1184 GNDA.n1159 3.4105
R11138 GNDA.n1184 GNDA.n1152 3.4105
R11139 GNDA.n1184 GNDA.n1160 3.4105
R11140 GNDA.n1184 GNDA.n1151 3.4105
R11141 GNDA.n1184 GNDA.n1161 3.4105
R11142 GNDA.n1184 GNDA.n1150 3.4105
R11143 GNDA.n1184 GNDA.n1162 3.4105
R11144 GNDA.n1184 GNDA.n1149 3.4105
R11145 GNDA.n1184 GNDA.n1163 3.4105
R11146 GNDA.n1184 GNDA.n1148 3.4105
R11147 GNDA.n1184 GNDA.n1164 3.4105
R11148 GNDA.n1184 GNDA.n1147 3.4105
R11149 GNDA.n1184 GNDA.n1165 3.4105
R11150 GNDA.n1184 GNDA.n1146 3.4105
R11151 GNDA.n1184 GNDA.n1166 3.4105
R11152 GNDA.n1184 GNDA.n1145 3.4105
R11153 GNDA.n1184 GNDA.n1167 3.4105
R11154 GNDA.n1184 GNDA.n1144 3.4105
R11155 GNDA.n1184 GNDA.n1168 3.4105
R11156 GNDA.n1184 GNDA.n1143 3.4105
R11157 GNDA.n1184 GNDA.n1169 3.4105
R11158 GNDA.n1184 GNDA.n1142 3.4105
R11159 GNDA.n1184 GNDA.n1170 3.4105
R11160 GNDA.n1184 GNDA.n1141 3.4105
R11161 GNDA.n1184 GNDA.n1171 3.4105
R11162 GNDA.n1184 GNDA.n1172 3.4105
R11163 GNDA.n2654 GNDA.n1184 3.4105
R11164 GNDA.n2616 GNDA.n1156 3.4105
R11165 GNDA.n2616 GNDA.n1155 3.4105
R11166 GNDA.n2616 GNDA.n1157 3.4105
R11167 GNDA.n2616 GNDA.n1154 3.4105
R11168 GNDA.n2616 GNDA.n1158 3.4105
R11169 GNDA.n2616 GNDA.n1153 3.4105
R11170 GNDA.n2616 GNDA.n1159 3.4105
R11171 GNDA.n2616 GNDA.n1152 3.4105
R11172 GNDA.n2616 GNDA.n1160 3.4105
R11173 GNDA.n2616 GNDA.n1151 3.4105
R11174 GNDA.n2616 GNDA.n1161 3.4105
R11175 GNDA.n2616 GNDA.n1150 3.4105
R11176 GNDA.n2616 GNDA.n1162 3.4105
R11177 GNDA.n2616 GNDA.n1149 3.4105
R11178 GNDA.n2616 GNDA.n1163 3.4105
R11179 GNDA.n2616 GNDA.n1148 3.4105
R11180 GNDA.n2616 GNDA.n1164 3.4105
R11181 GNDA.n2616 GNDA.n1147 3.4105
R11182 GNDA.n2616 GNDA.n1165 3.4105
R11183 GNDA.n2616 GNDA.n1146 3.4105
R11184 GNDA.n2616 GNDA.n1166 3.4105
R11185 GNDA.n2616 GNDA.n1145 3.4105
R11186 GNDA.n2616 GNDA.n1167 3.4105
R11187 GNDA.n2616 GNDA.n1144 3.4105
R11188 GNDA.n2616 GNDA.n1168 3.4105
R11189 GNDA.n2616 GNDA.n1143 3.4105
R11190 GNDA.n2616 GNDA.n1169 3.4105
R11191 GNDA.n2616 GNDA.n1142 3.4105
R11192 GNDA.n2616 GNDA.n1170 3.4105
R11193 GNDA.n2616 GNDA.n1141 3.4105
R11194 GNDA.n2616 GNDA.n1171 3.4105
R11195 GNDA.n2616 GNDA.n1172 3.4105
R11196 GNDA.n2654 GNDA.n2616 3.4105
R11197 GNDA.n1183 GNDA.n1156 3.4105
R11198 GNDA.n1183 GNDA.n1155 3.4105
R11199 GNDA.n1183 GNDA.n1157 3.4105
R11200 GNDA.n1183 GNDA.n1154 3.4105
R11201 GNDA.n1183 GNDA.n1158 3.4105
R11202 GNDA.n1183 GNDA.n1153 3.4105
R11203 GNDA.n1183 GNDA.n1159 3.4105
R11204 GNDA.n1183 GNDA.n1152 3.4105
R11205 GNDA.n1183 GNDA.n1160 3.4105
R11206 GNDA.n1183 GNDA.n1151 3.4105
R11207 GNDA.n1183 GNDA.n1161 3.4105
R11208 GNDA.n1183 GNDA.n1150 3.4105
R11209 GNDA.n1183 GNDA.n1162 3.4105
R11210 GNDA.n1183 GNDA.n1149 3.4105
R11211 GNDA.n1183 GNDA.n1163 3.4105
R11212 GNDA.n1183 GNDA.n1148 3.4105
R11213 GNDA.n1183 GNDA.n1164 3.4105
R11214 GNDA.n1183 GNDA.n1147 3.4105
R11215 GNDA.n1183 GNDA.n1165 3.4105
R11216 GNDA.n1183 GNDA.n1146 3.4105
R11217 GNDA.n1183 GNDA.n1166 3.4105
R11218 GNDA.n1183 GNDA.n1145 3.4105
R11219 GNDA.n1183 GNDA.n1167 3.4105
R11220 GNDA.n1183 GNDA.n1144 3.4105
R11221 GNDA.n1183 GNDA.n1168 3.4105
R11222 GNDA.n1183 GNDA.n1143 3.4105
R11223 GNDA.n1183 GNDA.n1169 3.4105
R11224 GNDA.n1183 GNDA.n1142 3.4105
R11225 GNDA.n1183 GNDA.n1170 3.4105
R11226 GNDA.n1183 GNDA.n1141 3.4105
R11227 GNDA.n1183 GNDA.n1171 3.4105
R11228 GNDA.n1183 GNDA.n1172 3.4105
R11229 GNDA.n2654 GNDA.n1183 3.4105
R11230 GNDA.n2618 GNDA.n1156 3.4105
R11231 GNDA.n2618 GNDA.n1155 3.4105
R11232 GNDA.n2618 GNDA.n1157 3.4105
R11233 GNDA.n2618 GNDA.n1154 3.4105
R11234 GNDA.n2618 GNDA.n1158 3.4105
R11235 GNDA.n2618 GNDA.n1153 3.4105
R11236 GNDA.n2618 GNDA.n1159 3.4105
R11237 GNDA.n2618 GNDA.n1152 3.4105
R11238 GNDA.n2618 GNDA.n1160 3.4105
R11239 GNDA.n2618 GNDA.n1151 3.4105
R11240 GNDA.n2618 GNDA.n1161 3.4105
R11241 GNDA.n2618 GNDA.n1150 3.4105
R11242 GNDA.n2618 GNDA.n1162 3.4105
R11243 GNDA.n2618 GNDA.n1149 3.4105
R11244 GNDA.n2618 GNDA.n1163 3.4105
R11245 GNDA.n2618 GNDA.n1148 3.4105
R11246 GNDA.n2618 GNDA.n1164 3.4105
R11247 GNDA.n2618 GNDA.n1147 3.4105
R11248 GNDA.n2618 GNDA.n1165 3.4105
R11249 GNDA.n2618 GNDA.n1146 3.4105
R11250 GNDA.n2618 GNDA.n1166 3.4105
R11251 GNDA.n2618 GNDA.n1145 3.4105
R11252 GNDA.n2618 GNDA.n1167 3.4105
R11253 GNDA.n2618 GNDA.n1144 3.4105
R11254 GNDA.n2618 GNDA.n1168 3.4105
R11255 GNDA.n2618 GNDA.n1143 3.4105
R11256 GNDA.n2618 GNDA.n1169 3.4105
R11257 GNDA.n2618 GNDA.n1142 3.4105
R11258 GNDA.n2618 GNDA.n1170 3.4105
R11259 GNDA.n2618 GNDA.n1141 3.4105
R11260 GNDA.n2618 GNDA.n1171 3.4105
R11261 GNDA.n2618 GNDA.n1172 3.4105
R11262 GNDA.n2654 GNDA.n2618 3.4105
R11263 GNDA.n1182 GNDA.n1156 3.4105
R11264 GNDA.n1182 GNDA.n1155 3.4105
R11265 GNDA.n1182 GNDA.n1157 3.4105
R11266 GNDA.n1182 GNDA.n1154 3.4105
R11267 GNDA.n1182 GNDA.n1158 3.4105
R11268 GNDA.n1182 GNDA.n1153 3.4105
R11269 GNDA.n1182 GNDA.n1159 3.4105
R11270 GNDA.n1182 GNDA.n1152 3.4105
R11271 GNDA.n1182 GNDA.n1160 3.4105
R11272 GNDA.n1182 GNDA.n1151 3.4105
R11273 GNDA.n1182 GNDA.n1161 3.4105
R11274 GNDA.n1182 GNDA.n1150 3.4105
R11275 GNDA.n1182 GNDA.n1162 3.4105
R11276 GNDA.n1182 GNDA.n1149 3.4105
R11277 GNDA.n1182 GNDA.n1163 3.4105
R11278 GNDA.n1182 GNDA.n1148 3.4105
R11279 GNDA.n1182 GNDA.n1164 3.4105
R11280 GNDA.n1182 GNDA.n1147 3.4105
R11281 GNDA.n1182 GNDA.n1165 3.4105
R11282 GNDA.n1182 GNDA.n1146 3.4105
R11283 GNDA.n1182 GNDA.n1166 3.4105
R11284 GNDA.n1182 GNDA.n1145 3.4105
R11285 GNDA.n1182 GNDA.n1167 3.4105
R11286 GNDA.n1182 GNDA.n1144 3.4105
R11287 GNDA.n1182 GNDA.n1168 3.4105
R11288 GNDA.n1182 GNDA.n1143 3.4105
R11289 GNDA.n1182 GNDA.n1169 3.4105
R11290 GNDA.n1182 GNDA.n1142 3.4105
R11291 GNDA.n1182 GNDA.n1170 3.4105
R11292 GNDA.n1182 GNDA.n1141 3.4105
R11293 GNDA.n1182 GNDA.n1171 3.4105
R11294 GNDA.n1182 GNDA.n1172 3.4105
R11295 GNDA.n2654 GNDA.n1182 3.4105
R11296 GNDA.n2620 GNDA.n1156 3.4105
R11297 GNDA.n2620 GNDA.n1155 3.4105
R11298 GNDA.n2620 GNDA.n1157 3.4105
R11299 GNDA.n2620 GNDA.n1154 3.4105
R11300 GNDA.n2620 GNDA.n1158 3.4105
R11301 GNDA.n2620 GNDA.n1153 3.4105
R11302 GNDA.n2620 GNDA.n1159 3.4105
R11303 GNDA.n2620 GNDA.n1152 3.4105
R11304 GNDA.n2620 GNDA.n1160 3.4105
R11305 GNDA.n2620 GNDA.n1151 3.4105
R11306 GNDA.n2620 GNDA.n1161 3.4105
R11307 GNDA.n2620 GNDA.n1150 3.4105
R11308 GNDA.n2620 GNDA.n1162 3.4105
R11309 GNDA.n2620 GNDA.n1149 3.4105
R11310 GNDA.n2620 GNDA.n1163 3.4105
R11311 GNDA.n2620 GNDA.n1148 3.4105
R11312 GNDA.n2620 GNDA.n1164 3.4105
R11313 GNDA.n2620 GNDA.n1147 3.4105
R11314 GNDA.n2620 GNDA.n1165 3.4105
R11315 GNDA.n2620 GNDA.n1146 3.4105
R11316 GNDA.n2620 GNDA.n1166 3.4105
R11317 GNDA.n2620 GNDA.n1145 3.4105
R11318 GNDA.n2620 GNDA.n1167 3.4105
R11319 GNDA.n2620 GNDA.n1144 3.4105
R11320 GNDA.n2620 GNDA.n1168 3.4105
R11321 GNDA.n2620 GNDA.n1143 3.4105
R11322 GNDA.n2620 GNDA.n1169 3.4105
R11323 GNDA.n2620 GNDA.n1142 3.4105
R11324 GNDA.n2620 GNDA.n1170 3.4105
R11325 GNDA.n2620 GNDA.n1141 3.4105
R11326 GNDA.n2620 GNDA.n1171 3.4105
R11327 GNDA.n2620 GNDA.n1172 3.4105
R11328 GNDA.n2654 GNDA.n2620 3.4105
R11329 GNDA.n1181 GNDA.n1156 3.4105
R11330 GNDA.n1181 GNDA.n1155 3.4105
R11331 GNDA.n1181 GNDA.n1157 3.4105
R11332 GNDA.n1181 GNDA.n1154 3.4105
R11333 GNDA.n1181 GNDA.n1158 3.4105
R11334 GNDA.n1181 GNDA.n1153 3.4105
R11335 GNDA.n1181 GNDA.n1159 3.4105
R11336 GNDA.n1181 GNDA.n1152 3.4105
R11337 GNDA.n1181 GNDA.n1160 3.4105
R11338 GNDA.n1181 GNDA.n1151 3.4105
R11339 GNDA.n1181 GNDA.n1161 3.4105
R11340 GNDA.n1181 GNDA.n1150 3.4105
R11341 GNDA.n1181 GNDA.n1162 3.4105
R11342 GNDA.n1181 GNDA.n1149 3.4105
R11343 GNDA.n1181 GNDA.n1163 3.4105
R11344 GNDA.n1181 GNDA.n1148 3.4105
R11345 GNDA.n1181 GNDA.n1164 3.4105
R11346 GNDA.n1181 GNDA.n1147 3.4105
R11347 GNDA.n1181 GNDA.n1165 3.4105
R11348 GNDA.n1181 GNDA.n1146 3.4105
R11349 GNDA.n1181 GNDA.n1166 3.4105
R11350 GNDA.n1181 GNDA.n1145 3.4105
R11351 GNDA.n1181 GNDA.n1167 3.4105
R11352 GNDA.n1181 GNDA.n1144 3.4105
R11353 GNDA.n1181 GNDA.n1168 3.4105
R11354 GNDA.n1181 GNDA.n1143 3.4105
R11355 GNDA.n1181 GNDA.n1169 3.4105
R11356 GNDA.n1181 GNDA.n1142 3.4105
R11357 GNDA.n1181 GNDA.n1170 3.4105
R11358 GNDA.n1181 GNDA.n1141 3.4105
R11359 GNDA.n1181 GNDA.n1171 3.4105
R11360 GNDA.n1181 GNDA.n1172 3.4105
R11361 GNDA.n2654 GNDA.n1181 3.4105
R11362 GNDA.n2622 GNDA.n1156 3.4105
R11363 GNDA.n2622 GNDA.n1155 3.4105
R11364 GNDA.n2622 GNDA.n1157 3.4105
R11365 GNDA.n2622 GNDA.n1154 3.4105
R11366 GNDA.n2622 GNDA.n1158 3.4105
R11367 GNDA.n2622 GNDA.n1153 3.4105
R11368 GNDA.n2622 GNDA.n1159 3.4105
R11369 GNDA.n2622 GNDA.n1152 3.4105
R11370 GNDA.n2622 GNDA.n1160 3.4105
R11371 GNDA.n2622 GNDA.n1151 3.4105
R11372 GNDA.n2622 GNDA.n1161 3.4105
R11373 GNDA.n2622 GNDA.n1150 3.4105
R11374 GNDA.n2622 GNDA.n1162 3.4105
R11375 GNDA.n2622 GNDA.n1149 3.4105
R11376 GNDA.n2622 GNDA.n1163 3.4105
R11377 GNDA.n2622 GNDA.n1148 3.4105
R11378 GNDA.n2622 GNDA.n1164 3.4105
R11379 GNDA.n2622 GNDA.n1147 3.4105
R11380 GNDA.n2622 GNDA.n1165 3.4105
R11381 GNDA.n2622 GNDA.n1146 3.4105
R11382 GNDA.n2622 GNDA.n1166 3.4105
R11383 GNDA.n2622 GNDA.n1145 3.4105
R11384 GNDA.n2622 GNDA.n1167 3.4105
R11385 GNDA.n2622 GNDA.n1144 3.4105
R11386 GNDA.n2622 GNDA.n1168 3.4105
R11387 GNDA.n2622 GNDA.n1143 3.4105
R11388 GNDA.n2622 GNDA.n1169 3.4105
R11389 GNDA.n2622 GNDA.n1142 3.4105
R11390 GNDA.n2622 GNDA.n1170 3.4105
R11391 GNDA.n2622 GNDA.n1141 3.4105
R11392 GNDA.n2622 GNDA.n1171 3.4105
R11393 GNDA.n2622 GNDA.n1172 3.4105
R11394 GNDA.n2654 GNDA.n2622 3.4105
R11395 GNDA.n1180 GNDA.n1156 3.4105
R11396 GNDA.n1180 GNDA.n1155 3.4105
R11397 GNDA.n1180 GNDA.n1157 3.4105
R11398 GNDA.n1180 GNDA.n1154 3.4105
R11399 GNDA.n1180 GNDA.n1158 3.4105
R11400 GNDA.n1180 GNDA.n1153 3.4105
R11401 GNDA.n1180 GNDA.n1159 3.4105
R11402 GNDA.n1180 GNDA.n1152 3.4105
R11403 GNDA.n1180 GNDA.n1160 3.4105
R11404 GNDA.n1180 GNDA.n1151 3.4105
R11405 GNDA.n1180 GNDA.n1161 3.4105
R11406 GNDA.n1180 GNDA.n1150 3.4105
R11407 GNDA.n1180 GNDA.n1162 3.4105
R11408 GNDA.n1180 GNDA.n1149 3.4105
R11409 GNDA.n1180 GNDA.n1163 3.4105
R11410 GNDA.n1180 GNDA.n1148 3.4105
R11411 GNDA.n1180 GNDA.n1164 3.4105
R11412 GNDA.n1180 GNDA.n1147 3.4105
R11413 GNDA.n1180 GNDA.n1165 3.4105
R11414 GNDA.n1180 GNDA.n1146 3.4105
R11415 GNDA.n1180 GNDA.n1166 3.4105
R11416 GNDA.n1180 GNDA.n1145 3.4105
R11417 GNDA.n1180 GNDA.n1167 3.4105
R11418 GNDA.n1180 GNDA.n1144 3.4105
R11419 GNDA.n1180 GNDA.n1168 3.4105
R11420 GNDA.n1180 GNDA.n1143 3.4105
R11421 GNDA.n1180 GNDA.n1169 3.4105
R11422 GNDA.n1180 GNDA.n1142 3.4105
R11423 GNDA.n1180 GNDA.n1170 3.4105
R11424 GNDA.n1180 GNDA.n1141 3.4105
R11425 GNDA.n1180 GNDA.n1171 3.4105
R11426 GNDA.n1180 GNDA.n1172 3.4105
R11427 GNDA.n2654 GNDA.n1180 3.4105
R11428 GNDA.n2624 GNDA.n1156 3.4105
R11429 GNDA.n2624 GNDA.n1155 3.4105
R11430 GNDA.n2624 GNDA.n1157 3.4105
R11431 GNDA.n2624 GNDA.n1154 3.4105
R11432 GNDA.n2624 GNDA.n1158 3.4105
R11433 GNDA.n2624 GNDA.n1153 3.4105
R11434 GNDA.n2624 GNDA.n1159 3.4105
R11435 GNDA.n2624 GNDA.n1152 3.4105
R11436 GNDA.n2624 GNDA.n1160 3.4105
R11437 GNDA.n2624 GNDA.n1151 3.4105
R11438 GNDA.n2624 GNDA.n1161 3.4105
R11439 GNDA.n2624 GNDA.n1150 3.4105
R11440 GNDA.n2624 GNDA.n1162 3.4105
R11441 GNDA.n2624 GNDA.n1149 3.4105
R11442 GNDA.n2624 GNDA.n1163 3.4105
R11443 GNDA.n2624 GNDA.n1148 3.4105
R11444 GNDA.n2624 GNDA.n1164 3.4105
R11445 GNDA.n2624 GNDA.n1147 3.4105
R11446 GNDA.n2624 GNDA.n1165 3.4105
R11447 GNDA.n2624 GNDA.n1146 3.4105
R11448 GNDA.n2624 GNDA.n1166 3.4105
R11449 GNDA.n2624 GNDA.n1145 3.4105
R11450 GNDA.n2624 GNDA.n1167 3.4105
R11451 GNDA.n2624 GNDA.n1144 3.4105
R11452 GNDA.n2624 GNDA.n1168 3.4105
R11453 GNDA.n2624 GNDA.n1143 3.4105
R11454 GNDA.n2624 GNDA.n1169 3.4105
R11455 GNDA.n2624 GNDA.n1142 3.4105
R11456 GNDA.n2624 GNDA.n1170 3.4105
R11457 GNDA.n2624 GNDA.n1141 3.4105
R11458 GNDA.n2624 GNDA.n1171 3.4105
R11459 GNDA.n2624 GNDA.n1172 3.4105
R11460 GNDA.n2654 GNDA.n2624 3.4105
R11461 GNDA.n1179 GNDA.n1156 3.4105
R11462 GNDA.n1179 GNDA.n1155 3.4105
R11463 GNDA.n1179 GNDA.n1157 3.4105
R11464 GNDA.n1179 GNDA.n1154 3.4105
R11465 GNDA.n1179 GNDA.n1158 3.4105
R11466 GNDA.n1179 GNDA.n1153 3.4105
R11467 GNDA.n1179 GNDA.n1159 3.4105
R11468 GNDA.n1179 GNDA.n1152 3.4105
R11469 GNDA.n1179 GNDA.n1160 3.4105
R11470 GNDA.n1179 GNDA.n1151 3.4105
R11471 GNDA.n1179 GNDA.n1161 3.4105
R11472 GNDA.n1179 GNDA.n1150 3.4105
R11473 GNDA.n1179 GNDA.n1162 3.4105
R11474 GNDA.n1179 GNDA.n1149 3.4105
R11475 GNDA.n1179 GNDA.n1163 3.4105
R11476 GNDA.n1179 GNDA.n1148 3.4105
R11477 GNDA.n1179 GNDA.n1164 3.4105
R11478 GNDA.n1179 GNDA.n1147 3.4105
R11479 GNDA.n1179 GNDA.n1165 3.4105
R11480 GNDA.n1179 GNDA.n1146 3.4105
R11481 GNDA.n1179 GNDA.n1166 3.4105
R11482 GNDA.n1179 GNDA.n1145 3.4105
R11483 GNDA.n1179 GNDA.n1167 3.4105
R11484 GNDA.n1179 GNDA.n1144 3.4105
R11485 GNDA.n1179 GNDA.n1168 3.4105
R11486 GNDA.n1179 GNDA.n1143 3.4105
R11487 GNDA.n1179 GNDA.n1169 3.4105
R11488 GNDA.n1179 GNDA.n1142 3.4105
R11489 GNDA.n1179 GNDA.n1170 3.4105
R11490 GNDA.n1179 GNDA.n1141 3.4105
R11491 GNDA.n1179 GNDA.n1171 3.4105
R11492 GNDA.n1179 GNDA.n1172 3.4105
R11493 GNDA.n2654 GNDA.n1179 3.4105
R11494 GNDA.n2626 GNDA.n1156 3.4105
R11495 GNDA.n2626 GNDA.n1155 3.4105
R11496 GNDA.n2626 GNDA.n1157 3.4105
R11497 GNDA.n2626 GNDA.n1154 3.4105
R11498 GNDA.n2626 GNDA.n1158 3.4105
R11499 GNDA.n2626 GNDA.n1153 3.4105
R11500 GNDA.n2626 GNDA.n1159 3.4105
R11501 GNDA.n2626 GNDA.n1152 3.4105
R11502 GNDA.n2626 GNDA.n1160 3.4105
R11503 GNDA.n2626 GNDA.n1151 3.4105
R11504 GNDA.n2626 GNDA.n1161 3.4105
R11505 GNDA.n2626 GNDA.n1150 3.4105
R11506 GNDA.n2626 GNDA.n1162 3.4105
R11507 GNDA.n2626 GNDA.n1149 3.4105
R11508 GNDA.n2626 GNDA.n1163 3.4105
R11509 GNDA.n2626 GNDA.n1148 3.4105
R11510 GNDA.n2626 GNDA.n1164 3.4105
R11511 GNDA.n2626 GNDA.n1147 3.4105
R11512 GNDA.n2626 GNDA.n1165 3.4105
R11513 GNDA.n2626 GNDA.n1146 3.4105
R11514 GNDA.n2626 GNDA.n1166 3.4105
R11515 GNDA.n2626 GNDA.n1145 3.4105
R11516 GNDA.n2626 GNDA.n1167 3.4105
R11517 GNDA.n2626 GNDA.n1144 3.4105
R11518 GNDA.n2626 GNDA.n1168 3.4105
R11519 GNDA.n2626 GNDA.n1143 3.4105
R11520 GNDA.n2626 GNDA.n1169 3.4105
R11521 GNDA.n2626 GNDA.n1142 3.4105
R11522 GNDA.n2626 GNDA.n1170 3.4105
R11523 GNDA.n2626 GNDA.n1141 3.4105
R11524 GNDA.n2626 GNDA.n1171 3.4105
R11525 GNDA.n2626 GNDA.n1172 3.4105
R11526 GNDA.n2654 GNDA.n2626 3.4105
R11527 GNDA.n1178 GNDA.n1156 3.4105
R11528 GNDA.n1178 GNDA.n1155 3.4105
R11529 GNDA.n1178 GNDA.n1157 3.4105
R11530 GNDA.n1178 GNDA.n1154 3.4105
R11531 GNDA.n1178 GNDA.n1158 3.4105
R11532 GNDA.n1178 GNDA.n1153 3.4105
R11533 GNDA.n1178 GNDA.n1159 3.4105
R11534 GNDA.n1178 GNDA.n1152 3.4105
R11535 GNDA.n1178 GNDA.n1160 3.4105
R11536 GNDA.n1178 GNDA.n1151 3.4105
R11537 GNDA.n1178 GNDA.n1161 3.4105
R11538 GNDA.n1178 GNDA.n1150 3.4105
R11539 GNDA.n1178 GNDA.n1162 3.4105
R11540 GNDA.n1178 GNDA.n1149 3.4105
R11541 GNDA.n1178 GNDA.n1163 3.4105
R11542 GNDA.n1178 GNDA.n1148 3.4105
R11543 GNDA.n1178 GNDA.n1164 3.4105
R11544 GNDA.n1178 GNDA.n1147 3.4105
R11545 GNDA.n1178 GNDA.n1165 3.4105
R11546 GNDA.n1178 GNDA.n1146 3.4105
R11547 GNDA.n1178 GNDA.n1166 3.4105
R11548 GNDA.n1178 GNDA.n1145 3.4105
R11549 GNDA.n1178 GNDA.n1167 3.4105
R11550 GNDA.n1178 GNDA.n1144 3.4105
R11551 GNDA.n1178 GNDA.n1168 3.4105
R11552 GNDA.n1178 GNDA.n1143 3.4105
R11553 GNDA.n1178 GNDA.n1169 3.4105
R11554 GNDA.n1178 GNDA.n1142 3.4105
R11555 GNDA.n1178 GNDA.n1170 3.4105
R11556 GNDA.n1178 GNDA.n1141 3.4105
R11557 GNDA.n1178 GNDA.n1171 3.4105
R11558 GNDA.n1178 GNDA.n1172 3.4105
R11559 GNDA.n2654 GNDA.n1178 3.4105
R11560 GNDA.n2628 GNDA.n1156 3.4105
R11561 GNDA.n2628 GNDA.n1155 3.4105
R11562 GNDA.n2628 GNDA.n1157 3.4105
R11563 GNDA.n2628 GNDA.n1154 3.4105
R11564 GNDA.n2628 GNDA.n1158 3.4105
R11565 GNDA.n2628 GNDA.n1153 3.4105
R11566 GNDA.n2628 GNDA.n1159 3.4105
R11567 GNDA.n2628 GNDA.n1152 3.4105
R11568 GNDA.n2628 GNDA.n1160 3.4105
R11569 GNDA.n2628 GNDA.n1151 3.4105
R11570 GNDA.n2628 GNDA.n1161 3.4105
R11571 GNDA.n2628 GNDA.n1150 3.4105
R11572 GNDA.n2628 GNDA.n1162 3.4105
R11573 GNDA.n2628 GNDA.n1149 3.4105
R11574 GNDA.n2628 GNDA.n1163 3.4105
R11575 GNDA.n2628 GNDA.n1148 3.4105
R11576 GNDA.n2628 GNDA.n1164 3.4105
R11577 GNDA.n2628 GNDA.n1147 3.4105
R11578 GNDA.n2628 GNDA.n1165 3.4105
R11579 GNDA.n2628 GNDA.n1146 3.4105
R11580 GNDA.n2628 GNDA.n1166 3.4105
R11581 GNDA.n2628 GNDA.n1145 3.4105
R11582 GNDA.n2628 GNDA.n1167 3.4105
R11583 GNDA.n2628 GNDA.n1144 3.4105
R11584 GNDA.n2628 GNDA.n1168 3.4105
R11585 GNDA.n2628 GNDA.n1143 3.4105
R11586 GNDA.n2628 GNDA.n1169 3.4105
R11587 GNDA.n2628 GNDA.n1142 3.4105
R11588 GNDA.n2628 GNDA.n1170 3.4105
R11589 GNDA.n2628 GNDA.n1141 3.4105
R11590 GNDA.n2628 GNDA.n1171 3.4105
R11591 GNDA.n2628 GNDA.n1172 3.4105
R11592 GNDA.n2654 GNDA.n2628 3.4105
R11593 GNDA.n1177 GNDA.n1156 3.4105
R11594 GNDA.n1177 GNDA.n1155 3.4105
R11595 GNDA.n1177 GNDA.n1157 3.4105
R11596 GNDA.n1177 GNDA.n1154 3.4105
R11597 GNDA.n1177 GNDA.n1158 3.4105
R11598 GNDA.n1177 GNDA.n1153 3.4105
R11599 GNDA.n1177 GNDA.n1159 3.4105
R11600 GNDA.n1177 GNDA.n1152 3.4105
R11601 GNDA.n1177 GNDA.n1160 3.4105
R11602 GNDA.n1177 GNDA.n1151 3.4105
R11603 GNDA.n1177 GNDA.n1161 3.4105
R11604 GNDA.n1177 GNDA.n1150 3.4105
R11605 GNDA.n1177 GNDA.n1162 3.4105
R11606 GNDA.n1177 GNDA.n1149 3.4105
R11607 GNDA.n1177 GNDA.n1163 3.4105
R11608 GNDA.n1177 GNDA.n1148 3.4105
R11609 GNDA.n1177 GNDA.n1164 3.4105
R11610 GNDA.n1177 GNDA.n1147 3.4105
R11611 GNDA.n1177 GNDA.n1165 3.4105
R11612 GNDA.n1177 GNDA.n1146 3.4105
R11613 GNDA.n1177 GNDA.n1166 3.4105
R11614 GNDA.n1177 GNDA.n1145 3.4105
R11615 GNDA.n1177 GNDA.n1167 3.4105
R11616 GNDA.n1177 GNDA.n1144 3.4105
R11617 GNDA.n1177 GNDA.n1168 3.4105
R11618 GNDA.n1177 GNDA.n1143 3.4105
R11619 GNDA.n1177 GNDA.n1169 3.4105
R11620 GNDA.n1177 GNDA.n1142 3.4105
R11621 GNDA.n1177 GNDA.n1170 3.4105
R11622 GNDA.n1177 GNDA.n1141 3.4105
R11623 GNDA.n1177 GNDA.n1171 3.4105
R11624 GNDA.n1177 GNDA.n1172 3.4105
R11625 GNDA.n2654 GNDA.n1177 3.4105
R11626 GNDA.n2630 GNDA.n1156 3.4105
R11627 GNDA.n2630 GNDA.n1155 3.4105
R11628 GNDA.n2630 GNDA.n1157 3.4105
R11629 GNDA.n2630 GNDA.n1154 3.4105
R11630 GNDA.n2630 GNDA.n1158 3.4105
R11631 GNDA.n2630 GNDA.n1153 3.4105
R11632 GNDA.n2630 GNDA.n1159 3.4105
R11633 GNDA.n2630 GNDA.n1152 3.4105
R11634 GNDA.n2630 GNDA.n1160 3.4105
R11635 GNDA.n2630 GNDA.n1151 3.4105
R11636 GNDA.n2630 GNDA.n1161 3.4105
R11637 GNDA.n2630 GNDA.n1150 3.4105
R11638 GNDA.n2630 GNDA.n1162 3.4105
R11639 GNDA.n2630 GNDA.n1149 3.4105
R11640 GNDA.n2630 GNDA.n1163 3.4105
R11641 GNDA.n2630 GNDA.n1148 3.4105
R11642 GNDA.n2630 GNDA.n1164 3.4105
R11643 GNDA.n2630 GNDA.n1147 3.4105
R11644 GNDA.n2630 GNDA.n1165 3.4105
R11645 GNDA.n2630 GNDA.n1146 3.4105
R11646 GNDA.n2630 GNDA.n1166 3.4105
R11647 GNDA.n2630 GNDA.n1145 3.4105
R11648 GNDA.n2630 GNDA.n1167 3.4105
R11649 GNDA.n2630 GNDA.n1144 3.4105
R11650 GNDA.n2630 GNDA.n1168 3.4105
R11651 GNDA.n2630 GNDA.n1143 3.4105
R11652 GNDA.n2630 GNDA.n1169 3.4105
R11653 GNDA.n2630 GNDA.n1142 3.4105
R11654 GNDA.n2630 GNDA.n1170 3.4105
R11655 GNDA.n2630 GNDA.n1141 3.4105
R11656 GNDA.n2630 GNDA.n1171 3.4105
R11657 GNDA.n2630 GNDA.n1172 3.4105
R11658 GNDA.n2654 GNDA.n2630 3.4105
R11659 GNDA.n1176 GNDA.n1156 3.4105
R11660 GNDA.n1176 GNDA.n1155 3.4105
R11661 GNDA.n1176 GNDA.n1157 3.4105
R11662 GNDA.n1176 GNDA.n1154 3.4105
R11663 GNDA.n1176 GNDA.n1158 3.4105
R11664 GNDA.n1176 GNDA.n1153 3.4105
R11665 GNDA.n1176 GNDA.n1159 3.4105
R11666 GNDA.n1176 GNDA.n1152 3.4105
R11667 GNDA.n1176 GNDA.n1160 3.4105
R11668 GNDA.n1176 GNDA.n1151 3.4105
R11669 GNDA.n1176 GNDA.n1161 3.4105
R11670 GNDA.n1176 GNDA.n1150 3.4105
R11671 GNDA.n1176 GNDA.n1162 3.4105
R11672 GNDA.n1176 GNDA.n1149 3.4105
R11673 GNDA.n1176 GNDA.n1163 3.4105
R11674 GNDA.n1176 GNDA.n1148 3.4105
R11675 GNDA.n1176 GNDA.n1164 3.4105
R11676 GNDA.n1176 GNDA.n1147 3.4105
R11677 GNDA.n1176 GNDA.n1165 3.4105
R11678 GNDA.n1176 GNDA.n1146 3.4105
R11679 GNDA.n1176 GNDA.n1166 3.4105
R11680 GNDA.n1176 GNDA.n1145 3.4105
R11681 GNDA.n1176 GNDA.n1167 3.4105
R11682 GNDA.n1176 GNDA.n1144 3.4105
R11683 GNDA.n1176 GNDA.n1168 3.4105
R11684 GNDA.n1176 GNDA.n1143 3.4105
R11685 GNDA.n1176 GNDA.n1169 3.4105
R11686 GNDA.n1176 GNDA.n1142 3.4105
R11687 GNDA.n1176 GNDA.n1170 3.4105
R11688 GNDA.n1176 GNDA.n1141 3.4105
R11689 GNDA.n1176 GNDA.n1171 3.4105
R11690 GNDA.n1176 GNDA.n1172 3.4105
R11691 GNDA.n2654 GNDA.n1176 3.4105
R11692 GNDA.n2632 GNDA.n1156 3.4105
R11693 GNDA.n2632 GNDA.n1155 3.4105
R11694 GNDA.n2632 GNDA.n1157 3.4105
R11695 GNDA.n2632 GNDA.n1154 3.4105
R11696 GNDA.n2632 GNDA.n1158 3.4105
R11697 GNDA.n2632 GNDA.n1153 3.4105
R11698 GNDA.n2632 GNDA.n1159 3.4105
R11699 GNDA.n2632 GNDA.n1152 3.4105
R11700 GNDA.n2632 GNDA.n1160 3.4105
R11701 GNDA.n2632 GNDA.n1151 3.4105
R11702 GNDA.n2632 GNDA.n1161 3.4105
R11703 GNDA.n2632 GNDA.n1150 3.4105
R11704 GNDA.n2632 GNDA.n1162 3.4105
R11705 GNDA.n2632 GNDA.n1149 3.4105
R11706 GNDA.n2632 GNDA.n1163 3.4105
R11707 GNDA.n2632 GNDA.n1148 3.4105
R11708 GNDA.n2632 GNDA.n1164 3.4105
R11709 GNDA.n2632 GNDA.n1147 3.4105
R11710 GNDA.n2632 GNDA.n1165 3.4105
R11711 GNDA.n2632 GNDA.n1146 3.4105
R11712 GNDA.n2632 GNDA.n1166 3.4105
R11713 GNDA.n2632 GNDA.n1145 3.4105
R11714 GNDA.n2632 GNDA.n1167 3.4105
R11715 GNDA.n2632 GNDA.n1144 3.4105
R11716 GNDA.n2632 GNDA.n1168 3.4105
R11717 GNDA.n2632 GNDA.n1143 3.4105
R11718 GNDA.n2632 GNDA.n1169 3.4105
R11719 GNDA.n2632 GNDA.n1142 3.4105
R11720 GNDA.n2632 GNDA.n1170 3.4105
R11721 GNDA.n2632 GNDA.n1141 3.4105
R11722 GNDA.n2632 GNDA.n1171 3.4105
R11723 GNDA.n2632 GNDA.n1172 3.4105
R11724 GNDA.n2654 GNDA.n2632 3.4105
R11725 GNDA.n1175 GNDA.n1156 3.4105
R11726 GNDA.n1175 GNDA.n1155 3.4105
R11727 GNDA.n1175 GNDA.n1157 3.4105
R11728 GNDA.n1175 GNDA.n1154 3.4105
R11729 GNDA.n1175 GNDA.n1158 3.4105
R11730 GNDA.n1175 GNDA.n1153 3.4105
R11731 GNDA.n1175 GNDA.n1159 3.4105
R11732 GNDA.n1175 GNDA.n1152 3.4105
R11733 GNDA.n1175 GNDA.n1160 3.4105
R11734 GNDA.n1175 GNDA.n1151 3.4105
R11735 GNDA.n1175 GNDA.n1161 3.4105
R11736 GNDA.n1175 GNDA.n1150 3.4105
R11737 GNDA.n1175 GNDA.n1162 3.4105
R11738 GNDA.n1175 GNDA.n1149 3.4105
R11739 GNDA.n1175 GNDA.n1163 3.4105
R11740 GNDA.n1175 GNDA.n1148 3.4105
R11741 GNDA.n1175 GNDA.n1164 3.4105
R11742 GNDA.n1175 GNDA.n1147 3.4105
R11743 GNDA.n1175 GNDA.n1165 3.4105
R11744 GNDA.n1175 GNDA.n1146 3.4105
R11745 GNDA.n1175 GNDA.n1166 3.4105
R11746 GNDA.n1175 GNDA.n1145 3.4105
R11747 GNDA.n1175 GNDA.n1167 3.4105
R11748 GNDA.n1175 GNDA.n1144 3.4105
R11749 GNDA.n1175 GNDA.n1168 3.4105
R11750 GNDA.n1175 GNDA.n1143 3.4105
R11751 GNDA.n1175 GNDA.n1169 3.4105
R11752 GNDA.n1175 GNDA.n1142 3.4105
R11753 GNDA.n1175 GNDA.n1170 3.4105
R11754 GNDA.n1175 GNDA.n1141 3.4105
R11755 GNDA.n1175 GNDA.n1171 3.4105
R11756 GNDA.n1175 GNDA.n1172 3.4105
R11757 GNDA.n2654 GNDA.n1175 3.4105
R11758 GNDA.n2634 GNDA.n1156 3.4105
R11759 GNDA.n2634 GNDA.n1155 3.4105
R11760 GNDA.n2634 GNDA.n1157 3.4105
R11761 GNDA.n2634 GNDA.n1154 3.4105
R11762 GNDA.n2634 GNDA.n1158 3.4105
R11763 GNDA.n2634 GNDA.n1153 3.4105
R11764 GNDA.n2634 GNDA.n1159 3.4105
R11765 GNDA.n2634 GNDA.n1152 3.4105
R11766 GNDA.n2634 GNDA.n1160 3.4105
R11767 GNDA.n2634 GNDA.n1151 3.4105
R11768 GNDA.n2634 GNDA.n1161 3.4105
R11769 GNDA.n2634 GNDA.n1150 3.4105
R11770 GNDA.n2634 GNDA.n1162 3.4105
R11771 GNDA.n2634 GNDA.n1149 3.4105
R11772 GNDA.n2634 GNDA.n1163 3.4105
R11773 GNDA.n2634 GNDA.n1148 3.4105
R11774 GNDA.n2634 GNDA.n1164 3.4105
R11775 GNDA.n2634 GNDA.n1147 3.4105
R11776 GNDA.n2634 GNDA.n1165 3.4105
R11777 GNDA.n2634 GNDA.n1146 3.4105
R11778 GNDA.n2634 GNDA.n1166 3.4105
R11779 GNDA.n2634 GNDA.n1145 3.4105
R11780 GNDA.n2634 GNDA.n1167 3.4105
R11781 GNDA.n2634 GNDA.n1144 3.4105
R11782 GNDA.n2634 GNDA.n1168 3.4105
R11783 GNDA.n2634 GNDA.n1143 3.4105
R11784 GNDA.n2634 GNDA.n1169 3.4105
R11785 GNDA.n2634 GNDA.n1142 3.4105
R11786 GNDA.n2634 GNDA.n1170 3.4105
R11787 GNDA.n2634 GNDA.n1141 3.4105
R11788 GNDA.n2634 GNDA.n1171 3.4105
R11789 GNDA.n2634 GNDA.n1172 3.4105
R11790 GNDA.n2654 GNDA.n2634 3.4105
R11791 GNDA.n1174 GNDA.n1156 3.4105
R11792 GNDA.n1174 GNDA.n1155 3.4105
R11793 GNDA.n1174 GNDA.n1157 3.4105
R11794 GNDA.n1174 GNDA.n1154 3.4105
R11795 GNDA.n1174 GNDA.n1158 3.4105
R11796 GNDA.n1174 GNDA.n1153 3.4105
R11797 GNDA.n1174 GNDA.n1159 3.4105
R11798 GNDA.n1174 GNDA.n1152 3.4105
R11799 GNDA.n1174 GNDA.n1160 3.4105
R11800 GNDA.n1174 GNDA.n1151 3.4105
R11801 GNDA.n1174 GNDA.n1161 3.4105
R11802 GNDA.n1174 GNDA.n1150 3.4105
R11803 GNDA.n1174 GNDA.n1162 3.4105
R11804 GNDA.n1174 GNDA.n1149 3.4105
R11805 GNDA.n1174 GNDA.n1163 3.4105
R11806 GNDA.n1174 GNDA.n1148 3.4105
R11807 GNDA.n1174 GNDA.n1164 3.4105
R11808 GNDA.n1174 GNDA.n1147 3.4105
R11809 GNDA.n1174 GNDA.n1165 3.4105
R11810 GNDA.n1174 GNDA.n1146 3.4105
R11811 GNDA.n1174 GNDA.n1166 3.4105
R11812 GNDA.n1174 GNDA.n1145 3.4105
R11813 GNDA.n1174 GNDA.n1167 3.4105
R11814 GNDA.n1174 GNDA.n1144 3.4105
R11815 GNDA.n1174 GNDA.n1168 3.4105
R11816 GNDA.n1174 GNDA.n1143 3.4105
R11817 GNDA.n1174 GNDA.n1169 3.4105
R11818 GNDA.n1174 GNDA.n1142 3.4105
R11819 GNDA.n1174 GNDA.n1170 3.4105
R11820 GNDA.n1174 GNDA.n1141 3.4105
R11821 GNDA.n1174 GNDA.n1171 3.4105
R11822 GNDA.n1174 GNDA.n1172 3.4105
R11823 GNDA.n2654 GNDA.n1174 3.4105
R11824 GNDA.n2653 GNDA.n1156 3.4105
R11825 GNDA.n2653 GNDA.n1155 3.4105
R11826 GNDA.n2653 GNDA.n1157 3.4105
R11827 GNDA.n2653 GNDA.n1154 3.4105
R11828 GNDA.n2653 GNDA.n1158 3.4105
R11829 GNDA.n2653 GNDA.n1153 3.4105
R11830 GNDA.n2653 GNDA.n1159 3.4105
R11831 GNDA.n2653 GNDA.n1152 3.4105
R11832 GNDA.n2653 GNDA.n1160 3.4105
R11833 GNDA.n2653 GNDA.n1151 3.4105
R11834 GNDA.n2653 GNDA.n1161 3.4105
R11835 GNDA.n2653 GNDA.n1150 3.4105
R11836 GNDA.n2653 GNDA.n1162 3.4105
R11837 GNDA.n2653 GNDA.n1149 3.4105
R11838 GNDA.n2653 GNDA.n1163 3.4105
R11839 GNDA.n2653 GNDA.n1148 3.4105
R11840 GNDA.n2653 GNDA.n1164 3.4105
R11841 GNDA.n2653 GNDA.n1147 3.4105
R11842 GNDA.n2653 GNDA.n1165 3.4105
R11843 GNDA.n2653 GNDA.n1146 3.4105
R11844 GNDA.n2653 GNDA.n1166 3.4105
R11845 GNDA.n2653 GNDA.n1145 3.4105
R11846 GNDA.n2653 GNDA.n1167 3.4105
R11847 GNDA.n2653 GNDA.n1144 3.4105
R11848 GNDA.n2653 GNDA.n1168 3.4105
R11849 GNDA.n2653 GNDA.n1143 3.4105
R11850 GNDA.n2653 GNDA.n1169 3.4105
R11851 GNDA.n2653 GNDA.n1142 3.4105
R11852 GNDA.n2653 GNDA.n1170 3.4105
R11853 GNDA.n2653 GNDA.n1141 3.4105
R11854 GNDA.n2653 GNDA.n1171 3.4105
R11855 GNDA.n2653 GNDA.n1172 3.4105
R11856 GNDA.n2654 GNDA.n2653 3.4105
R11857 GNDA.n1173 GNDA.n1156 3.4105
R11858 GNDA.n1173 GNDA.n1155 3.4105
R11859 GNDA.n1173 GNDA.n1157 3.4105
R11860 GNDA.n1173 GNDA.n1154 3.4105
R11861 GNDA.n1173 GNDA.n1158 3.4105
R11862 GNDA.n1173 GNDA.n1153 3.4105
R11863 GNDA.n1173 GNDA.n1159 3.4105
R11864 GNDA.n1173 GNDA.n1152 3.4105
R11865 GNDA.n1173 GNDA.n1160 3.4105
R11866 GNDA.n1173 GNDA.n1151 3.4105
R11867 GNDA.n1173 GNDA.n1161 3.4105
R11868 GNDA.n1173 GNDA.n1150 3.4105
R11869 GNDA.n1173 GNDA.n1162 3.4105
R11870 GNDA.n1173 GNDA.n1149 3.4105
R11871 GNDA.n1173 GNDA.n1163 3.4105
R11872 GNDA.n1173 GNDA.n1148 3.4105
R11873 GNDA.n1173 GNDA.n1164 3.4105
R11874 GNDA.n1173 GNDA.n1147 3.4105
R11875 GNDA.n1173 GNDA.n1165 3.4105
R11876 GNDA.n1173 GNDA.n1146 3.4105
R11877 GNDA.n1173 GNDA.n1166 3.4105
R11878 GNDA.n1173 GNDA.n1145 3.4105
R11879 GNDA.n1173 GNDA.n1167 3.4105
R11880 GNDA.n1173 GNDA.n1144 3.4105
R11881 GNDA.n1173 GNDA.n1168 3.4105
R11882 GNDA.n1173 GNDA.n1143 3.4105
R11883 GNDA.n1173 GNDA.n1169 3.4105
R11884 GNDA.n1173 GNDA.n1142 3.4105
R11885 GNDA.n1173 GNDA.n1170 3.4105
R11886 GNDA.n1173 GNDA.n1141 3.4105
R11887 GNDA.n1173 GNDA.n1171 3.4105
R11888 GNDA.n1173 GNDA.n1172 3.4105
R11889 GNDA.n2654 GNDA.n1173 3.4105
R11890 GNDA.n2655 GNDA.n1156 3.4105
R11891 GNDA.n2655 GNDA.n1155 3.4105
R11892 GNDA.n2655 GNDA.n1157 3.4105
R11893 GNDA.n2655 GNDA.n1154 3.4105
R11894 GNDA.n2655 GNDA.n1158 3.4105
R11895 GNDA.n2655 GNDA.n1153 3.4105
R11896 GNDA.n2655 GNDA.n1159 3.4105
R11897 GNDA.n2655 GNDA.n1152 3.4105
R11898 GNDA.n2655 GNDA.n1160 3.4105
R11899 GNDA.n2655 GNDA.n1151 3.4105
R11900 GNDA.n2655 GNDA.n1161 3.4105
R11901 GNDA.n2655 GNDA.n1150 3.4105
R11902 GNDA.n2655 GNDA.n1162 3.4105
R11903 GNDA.n2655 GNDA.n1149 3.4105
R11904 GNDA.n2655 GNDA.n1163 3.4105
R11905 GNDA.n2655 GNDA.n1148 3.4105
R11906 GNDA.n2655 GNDA.n1164 3.4105
R11907 GNDA.n2655 GNDA.n1147 3.4105
R11908 GNDA.n2655 GNDA.n1165 3.4105
R11909 GNDA.n2655 GNDA.n1146 3.4105
R11910 GNDA.n2655 GNDA.n1166 3.4105
R11911 GNDA.n2655 GNDA.n1145 3.4105
R11912 GNDA.n2655 GNDA.n1167 3.4105
R11913 GNDA.n2655 GNDA.n1144 3.4105
R11914 GNDA.n2655 GNDA.n1168 3.4105
R11915 GNDA.n2655 GNDA.n1143 3.4105
R11916 GNDA.n2655 GNDA.n1169 3.4105
R11917 GNDA.n2655 GNDA.n1142 3.4105
R11918 GNDA.n2655 GNDA.n1170 3.4105
R11919 GNDA.n2655 GNDA.n1141 3.4105
R11920 GNDA.n2655 GNDA.n1171 3.4105
R11921 GNDA.n2655 GNDA.n1140 3.4105
R11922 GNDA.n2655 GNDA.n1172 3.4105
R11923 GNDA.n2655 GNDA.n2654 3.4105
R11924 GNDA.n737 GNDA.n736 3.08383
R11925 GNDA.n640 GNDA.n639 3.08383
R11926 GNDA.n2527 GNDA.n1551 3.04346
R11927 GNDA.n1868 GNDA.n1866 3.00528
R11928 GNDA.n1916 GNDA.n1911 3.00528
R11929 GNDA.n2496 GNDA.t14 3.00528
R11930 GNDA.n1575 GNDA.t28 3.00528
R11931 GNDA.n2514 GNDA.n1556 2.86505
R11932 GNDA.n2515 GNDA.n2514 2.86505
R11933 GNDA.n2513 GNDA.n2509 2.86505
R11934 GNDA.n2510 GNDA.n2509 2.86505
R11935 GNDA.n2516 GNDA.n2515 2.86505
R11936 GNDA.n2511 GNDA.n2510 2.86505
R11937 GNDA.n2520 GNDA.n1556 2.86505
R11938 GNDA.n2516 GNDA.n2513 2.86505
R11939 GNDA.n2061 GNDA.n2060 2.86505
R11940 GNDA.n2060 GNDA.n2058 2.86505
R11941 GNDA.n2058 GNDA.n2057 2.86505
R11942 GNDA.n2062 GNDA.n2061 2.86505
R11943 GNDA.n2570 GNDA.n2568 2.69842
R11944 GNDA.n1655 GNDA.n1654 2.6629
R11945 GNDA.n1997 GNDA.n1714 2.6629
R11946 GNDA.n2036 GNDA.n1656 2.6629
R11947 GNDA.n5339 GNDA.n5338 2.6629
R11948 GNDA.n2137 GNDA.n2136 2.6629
R11949 GNDA.n2264 GNDA.n2263 2.6629
R11950 GNDA.n5268 GNDA.n5267 2.6629
R11951 GNDA.n5181 GNDA.n160 2.6629
R11952 GNDA.n5547 GNDA.n5546 2.6629
R11953 GNDA.n5460 GNDA.n82 2.6629
R11954 GNDA.n5124 GNDA.n5123 2.6629
R11955 GNDA.n5032 GNDA.n56 2.6629
R11956 GNDA.n1857 GNDA.n1856 2.6629
R11957 GNDA.n2088 GNDA.n2087 2.6629
R11958 GNDA.n5454 GNDA.n5453 2.6629
R11959 GNDA.t186 GNDA.t232 2.59854
R11960 GNDA.n4008 GNDA.n4007 2.46404
R11961 GNDA.n3995 GNDA.n3994 2.46404
R11962 GNDA.n1656 GNDA.n1655 2.4581
R11963 GNDA.n2541 GNDA.n2540 2.4581
R11964 GNDA.n2088 GNDA.n1714 2.4581
R11965 GNDA.n2037 GNDA.n2036 2.4581
R11966 GNDA.n5339 GNDA.n160 2.4581
R11967 GNDA.n2136 GNDA.n186 2.4581
R11968 GNDA.n2263 GNDA.n2137 2.4581
R11969 GNDA.n2301 GNDA.n2300 2.4581
R11970 GNDA.n5182 GNDA.n5181 2.4581
R11971 GNDA.n5547 GNDA.n56 2.4581
R11972 GNDA.n5461 GNDA.n5460 2.4581
R11973 GNDA.n5033 GNDA.n5032 2.4581
R11974 GNDA.n2087 GNDA.n1716 2.4581
R11975 GNDA.n5454 GNDA.n82 2.4581
R11976 GNDA.n5387 GNDA.n5386 2.4581
R11977 GNDA.n2530 GNDA.n2529 2.44675
R11978 GNDA.n2529 GNDA.n2528 2.44675
R11979 GNDA.n1365 GNDA.n1364 2.39683
R11980 GNDA.n1489 GNDA.n1486 2.30736
R11981 GNDA.n4721 GNDA.n4720 2.30736
R11982 GNDA.n4645 GNDA.n4644 2.30736
R11983 GNDA.n4515 GNDA.n4514 2.30736
R11984 GNDA.n4805 GNDA.n4804 2.30736
R11985 GNDA.n4269 GNDA.n4268 2.30736
R11986 GNDA.n4870 GNDA.n4869 2.30736
R11987 GNDA.n4430 GNDA.n4429 2.30736
R11988 GNDA.n4327 GNDA.n4326 2.30736
R11989 GNDA.n4193 GNDA.n4192 2.30736
R11990 GNDA.n3953 GNDA.n798 2.30736
R11991 GNDA.n3616 GNDA.n3615 2.30736
R11992 GNDA.n3932 GNDA.n3931 2.30736
R11993 GNDA.n887 GNDA.n879 2.30736
R11994 GNDA.n3720 GNDA.n3719 2.30736
R11995 GNDA.n3789 GNDA.n3788 2.30736
R11996 GNDA.n3854 GNDA.n3853 2.30736
R11997 GNDA.n3441 GNDA.n3433 2.30736
R11998 GNDA.n3534 GNDA.n3533 2.30736
R11999 GNDA.n2855 GNDA.n2854 2.30736
R12000 GNDA.n2924 GNDA.n2923 2.30736
R12001 GNDA.n2993 GNDA.n2992 2.30736
R12002 GNDA.n3062 GNDA.n3061 2.30736
R12003 GNDA.n3131 GNDA.n3130 2.30736
R12004 GNDA.n3200 GNDA.n3199 2.30736
R12005 GNDA.n3269 GNDA.n3268 2.30736
R12006 GNDA.n3334 GNDA.n3333 2.30736
R12007 GNDA.n559 GNDA.n551 2.30736
R12008 GNDA.n4913 GNDA.n4912 2.29914
R12009 GNDA.n4127 GNDA.n432 2.29914
R12010 GNDA.n4070 GNDA.n4069 2.29914
R12011 GNDA.n3380 GNDA.n630 2.29878
R12012 GNDA.n2576 GNDA.n2575 2.29738
R12013 GNDA.n4013 GNDA.n4012 2.26187
R12014 GNDA.n933 GNDA.n755 2.26187
R12015 GNDA.n652 GNDA.n649 2.26187
R12016 GNDA.n653 GNDA.n652 2.26187
R12017 GNDA.n704 GNDA.n703 2.26187
R12018 GNDA.n1015 GNDA.n999 2.26187
R12019 GNDA.n3361 GNDA.n993 2.26187
R12020 GNDA.n3342 GNDA.n3341 2.26187
R12021 GNDA.n4884 GNDA.n4882 2.26187
R12022 GNDA.n1921 GNDA.n1893 2.26187
R12023 GNDA.n2524 GNDA.n2523 2.26187
R12024 GNDA.n2569 GNDA.n1416 2.26187
R12025 GNDA.n1422 GNDA.n1419 2.26187
R12026 GNDA.n1423 GNDA.n1422 2.26187
R12027 GNDA.n3991 GNDA.n3990 2.26187
R12028 GNDA.n768 GNDA.n767 2.26187
R12029 GNDA.n4014 GNDA.n4013 2.26187
R12030 GNDA.n3867 GNDA.n927 2.26187
R12031 GNDA.n3872 GNDA.n923 2.26187
R12032 GNDA.n3877 GNDA.n839 2.26187
R12033 GNDA.n3884 GNDA.n3883 2.26187
R12034 GNDA.n3864 GNDA.n3863 2.26187
R12035 GNDA.n4901 GNDA.n4888 2.26187
R12036 GNDA.n4902 GNDA.n4901 2.26187
R12037 GNDA.n659 GNDA.n658 2.26187
R12038 GNDA.n4094 GNDA.n4093 2.26187
R12039 GNDA.n4108 GNDA.n4107 2.26187
R12040 GNDA.n4112 GNDA.n4111 2.26187
R12041 GNDA.n717 GNDA.n716 2.26187
R12042 GNDA.n705 GNDA.n704 2.26187
R12043 GNDA.n1012 GNDA.n999 2.26187
R12044 GNDA.n3346 GNDA.n1032 2.26187
R12045 GNDA.n3351 GNDA.n1028 2.26187
R12046 GNDA.n3356 GNDA.n1024 2.26187
R12047 GNDA.n3366 GNDA.n989 2.26187
R12048 GNDA.n3371 GNDA.n985 2.26187
R12049 GNDA.n3376 GNDA.n981 2.26187
R12050 GNDA.n3486 GNDA.n3485 2.26187
R12051 GNDA.n3343 GNDA.n3342 2.26187
R12052 GNDA.n595 GNDA.n512 2.26187
R12053 GNDA.n2525 GNDA.n2524 2.26187
R12054 GNDA.n1887 GNDA.n1886 2.26187
R12055 GNDA.n3393 GNDA.n977 2.24241
R12056 GNDA.n978 GNDA.n976 2.24241
R12057 GNDA.n4279 GNDA.n478 2.24241
R12058 GNDA.n480 GNDA.n477 2.24241
R12059 GNDA.n3994 GNDA.n761 2.24063
R12060 GNDA.n3990 GNDA.n3989 2.24063
R12061 GNDA.n767 GNDA.n764 2.24063
R12062 GNDA.n766 GNDA.n763 2.24063
R12063 GNDA.n4011 GNDA.n752 2.24063
R12064 GNDA.n934 GNDA.n758 2.24063
R12065 GNDA.n3870 GNDA.n927 2.24063
R12066 GNDA.n928 GNDA.n926 2.24063
R12067 GNDA.n3875 GNDA.n923 2.24063
R12068 GNDA.n924 GNDA.n922 2.24063
R12069 GNDA.n3880 GNDA.n839 2.24063
R12070 GNDA.n840 GNDA.n838 2.24063
R12071 GNDA.n3883 GNDA.n772 2.24063
R12072 GNDA.n3882 GNDA.n837 2.24063
R12073 GNDA.n3862 GNDA.n3861 2.24063
R12074 GNDA.n3860 GNDA.n930 2.24063
R12075 GNDA.n4905 GNDA.n4900 2.24063
R12076 GNDA.n4906 GNDA.n4888 2.24063
R12077 GNDA.n4909 GNDA.n4908 2.24063
R12078 GNDA.n4887 GNDA.n435 2.24063
R12079 GNDA.n4097 GNDA.n4090 2.24063
R12080 GNDA.n4098 GNDA.n4088 2.24063
R12081 GNDA.n4103 GNDA.n616 2.24063
R12082 GNDA.n617 GNDA.n615 2.24063
R12083 GNDA.n4115 GNDA.n607 2.24063
R12084 GNDA.n4111 GNDA.n4110 2.24063
R12085 GNDA.n4105 GNDA.n4104 2.24063
R12086 GNDA.n4107 GNDA.n4106 2.24063
R12087 GNDA.n662 GNDA.n647 2.24063
R12088 GNDA.n659 GNDA.n657 2.24063
R12089 GNDA.n716 GNDA.n715 2.24063
R12090 GNDA.n714 GNDA.n713 2.24063
R12091 GNDA.n702 GNDA.n680 2.24063
R12092 GNDA.n696 GNDA.n695 2.24063
R12093 GNDA.n698 GNDA.n683 2.24063
R12094 GNDA.n699 GNDA.n620 2.24063
R12095 GNDA.n4086 GNDA.n619 2.24063
R12096 GNDA.n621 GNDA.n618 2.24063
R12097 GNDA.n4083 GNDA.n4082 2.24063
R12098 GNDA.n4076 GNDA.n624 2.24063
R12099 GNDA.n4078 GNDA.n623 2.24063
R12100 GNDA.n4079 GNDA.n4077 2.24063
R12101 GNDA.n1016 GNDA.n998 2.24063
R12102 GNDA.n1017 GNDA.n995 2.24063
R12103 GNDA.n997 GNDA.n994 2.24063
R12104 GNDA.n4074 GNDA.n4073 2.24063
R12105 GNDA.n629 GNDA.n628 2.24063
R12106 GNDA.n3349 GNDA.n1032 2.24063
R12107 GNDA.n1033 GNDA.n1031 2.24063
R12108 GNDA.n3354 GNDA.n1028 2.24063
R12109 GNDA.n1029 GNDA.n1027 2.24063
R12110 GNDA.n3359 GNDA.n1024 2.24063
R12111 GNDA.n1025 GNDA.n1023 2.24063
R12112 GNDA.n3369 GNDA.n989 2.24063
R12113 GNDA.n990 GNDA.n988 2.24063
R12114 GNDA.n3374 GNDA.n985 2.24063
R12115 GNDA.n986 GNDA.n984 2.24063
R12116 GNDA.n3379 GNDA.n981 2.24063
R12117 GNDA.n982 GNDA.n980 2.24063
R12118 GNDA.n3485 GNDA.n975 2.24063
R12119 GNDA.n3484 GNDA.n974 2.24063
R12120 GNDA.n3364 GNDA.n993 2.24063
R12121 GNDA.n1022 GNDA.n992 2.24063
R12122 GNDA.n3340 GNDA.n1035 2.24063
R12123 GNDA.n598 GNDA.n512 2.24063
R12124 GNDA.n513 GNDA.n511 2.24063
R12125 GNDA.n4369 GNDA.n475 2.24063
R12126 GNDA.n476 GNDA.n474 2.24063
R12127 GNDA.n4366 GNDA.n4365 2.24063
R12128 GNDA.n4373 GNDA.n441 2.24063
R12129 GNDA.n473 GNDA.n472 2.24063
R12130 GNDA.n4374 GNDA.n471 2.24063
R12131 GNDA.n4880 GNDA.n439 2.24063
R12132 GNDA.n440 GNDA.n438 2.24063
R12133 GNDA.n4877 GNDA.n4876 2.24063
R12134 GNDA.n4276 GNDA.n4275 2.24063
R12135 GNDA.n4748 GNDA.n4742 2.24063
R12136 GNDA.n4744 GNDA.n4743 2.24063
R12137 GNDA.n4749 GNDA.n4469 2.24063
R12138 GNDA.n4738 GNDA.n4555 2.24063
R12139 GNDA.n4739 GNDA.n4554 2.24063
R12140 GNDA.n4740 GNDA.n4553 2.24063
R12141 GNDA.n4734 GNDA.n4560 2.24063
R12142 GNDA.n4735 GNDA.n4559 2.24063
R12143 GNDA.n4736 GNDA.n4558 2.24063
R12144 GNDA.n4730 GNDA.n4729 2.24063
R12145 GNDA.n4731 GNDA.n4728 2.24063
R12146 GNDA.n4732 GNDA.n4727 2.24063
R12147 GNDA.n4882 GNDA.n437 2.24063
R12148 GNDA.n4883 GNDA.n436 2.24063
R12149 GNDA.n1922 GNDA.n1921 2.24063
R12150 GNDA.n1886 GNDA.n1555 2.24063
R12151 GNDA.n1889 GNDA.n1888 2.24063
R12152 GNDA.n2523 GNDA.n2522 2.24063
R12153 GNDA.n1547 GNDA.n1459 2.24063
R12154 GNDA.n1465 GNDA.n1458 2.24063
R12155 GNDA.n2571 GNDA.n2570 2.24063
R12156 GNDA.n3993 GNDA.n3992 2.24063
R12157 GNDA.n4015 GNDA.n4014 2.24063
R12158 GNDA.n4010 GNDA.n755 2.24063
R12159 GNDA.n4009 GNDA.n4008 2.24063
R12160 GNDA.n3865 GNDA.n3864 2.24063
R12161 GNDA.n4907 GNDA.n434 2.24063
R12162 GNDA.n4093 GNDA.n4092 2.24063
R12163 GNDA.n4100 GNDA.n4099 2.24063
R12164 GNDA.n4114 GNDA.n4113 2.24063
R12165 GNDA.n4109 GNDA.n611 2.24063
R12166 GNDA.n661 GNDA.n614 2.24063
R12167 GNDA.n656 GNDA.n649 2.24063
R12168 GNDA.n655 GNDA.n654 2.24063
R12169 GNDA.n706 GNDA.n705 2.24063
R12170 GNDA.n1012 GNDA.n1011 2.24063
R12171 GNDA.n1019 GNDA.n1018 2.24063
R12172 GNDA.n4075 GNDA.n626 2.24063
R12173 GNDA.n3390 GNDA.n3389 2.24063
R12174 GNDA.n3344 GNDA.n3343 2.24063
R12175 GNDA.n2051 GNDA.n1890 2.24063
R12176 GNDA.n2050 GNDA.n2049 2.24063
R12177 GNDA.n2526 GNDA.n1552 2.24063
R12178 GNDA.n1549 GNDA.n1548 2.24063
R12179 GNDA.n2575 GNDA.n1416 2.24063
R12180 GNDA.n2574 GNDA.n2573 2.24063
R12181 GNDA.n2568 GNDA.n1419 2.24063
R12182 GNDA.n2567 GNDA.n2566 2.24063
R12183 GNDA.n4049 GNDA.n4048 2.22018
R12184 GNDA.n4056 GNDA.n749 2.22018
R12185 GNDA.n667 GNDA.n665 2.22018
R12186 GNDA.n732 GNDA.n731 2.22018
R12187 GNDA.n694 GNDA.n684 2.22018
R12188 GNDA.n4116 GNDA.n605 2.22018
R12189 GNDA.n1923 GNDA.n1919 2.22018
R12190 GNDA.n2048 GNDA.n1894 2.22018
R12191 GNDA.n1461 GNDA.n1460 2.22018
R12192 GNDA.t270 GNDA.t174 2.21824
R12193 GNDA.t176 GNDA.t263 2.21824
R12194 GNDA.t194 GNDA.t121 2.21824
R12195 GNDA.t85 GNDA.t180 2.21824
R12196 GNDA.n328 GNDA.n56 2.18124
R12197 GNDA.n5343 GNDA.n160 2.18124
R12198 GNDA.n2089 GNDA.n2088 2.18124
R12199 GNDA.n389 GNDA.n82 2.18124
R12200 GNDA.n2383 GNDA.n2137 2.18124
R12201 GNDA.n2477 GNDA.n1656 2.18124
R12202 GNDA.n1548 GNDA.n1546 2.16717
R12203 GNDA.n2542 GNDA.n2541 2.1509
R12204 GNDA.n2038 GNDA.n2037 2.1509
R12205 GNDA.n5274 GNDA.n186 2.1509
R12206 GNDA.n2300 GNDA.n2299 2.1509
R12207 GNDA.n5200 GNDA.n5182 2.1509
R12208 GNDA.n5479 GNDA.n5461 2.1509
R12209 GNDA.n5059 GNDA.n5033 2.1509
R12210 GNDA.n1721 GNDA.n1716 2.1509
R12211 GNDA.n5397 GNDA.n5387 2.1509
R12212 GNDA.n1654 GNDA.n1653 2.13383
R12213 GNDA.n1998 GNDA.n1997 2.13383
R12214 GNDA.n5338 GNDA.n164 2.13383
R12215 GNDA.n5123 GNDA.n5010 2.13383
R12216 GNDA.n2264 GNDA.n2262 2.13383
R12217 GNDA.n5267 GNDA.n5154 2.13383
R12218 GNDA.n5546 GNDA.n57 2.13383
R12219 GNDA.n1857 GNDA.n1801 2.13383
R12220 GNDA.n5453 GNDA.n5452 2.13383
R12221 GNDA.n4281 GNDA.n4280 2.09414
R12222 GNDA.n3481 GNDA.n3480 2.09414
R12223 GNDA.n3385 GNDA.n3384 2.09414
R12224 GNDA.n4132 GNDA.n4131 2.09414
R12225 GNDA.n133 GNDA.n56 2.08643
R12226 GNDA.n162 GNDA.n160 2.08643
R12227 GNDA.n2088 GNDA.n1715 2.08643
R12228 GNDA.n84 GNDA.n82 2.08643
R12229 GNDA.n2386 GNDA.n2137 2.08643
R12230 GNDA.n1656 GNDA.n1600 2.08643
R12231 GNDA.n1654 GNDA.n1597 1.9461
R12232 GNDA.n1997 GNDA.n1996 1.9461
R12233 GNDA.n5338 GNDA.n5337 1.9461
R12234 GNDA.n2265 GNDA.n2264 1.9461
R12235 GNDA.n5267 GNDA.n5266 1.9461
R12236 GNDA.n5546 GNDA.n5545 1.9461
R12237 GNDA.n5123 GNDA.n5122 1.9461
R12238 GNDA.n1859 GNDA.n1857 1.9461
R12239 GNDA.n5453 GNDA.n22 1.9461
R12240 GNDA.n4914 GNDA.n4913 1.93383
R12241 GNDA.n4128 GNDA.n4127 1.93383
R12242 GNDA.n4069 GNDA.n4068 1.93383
R12243 GNDA.n3381 GNDA.n3380 1.93383
R12244 GNDA.n4910 GNDA.n4886 1.82342
R12245 GNDA.n3363 GNDA.n1021 1.82342
R12246 GNDA.n2522 GNDA.n2521 1.71925
R12247 GNDA.n1287 GNDA.n1286 1.70567
R12248 GNDA.n1287 GNDA.n1285 1.70567
R12249 GNDA.n1287 GNDA.n1284 1.70567
R12250 GNDA.n1287 GNDA.n1283 1.70567
R12251 GNDA.n1287 GNDA.n1282 1.70567
R12252 GNDA.n1287 GNDA.n1281 1.70567
R12253 GNDA.n1287 GNDA.n1280 1.70567
R12254 GNDA.n1287 GNDA.n1279 1.70567
R12255 GNDA.n1287 GNDA.n1278 1.70567
R12256 GNDA.n1287 GNDA.n1277 1.70567
R12257 GNDA.n1287 GNDA.n1276 1.70567
R12258 GNDA.n1287 GNDA.n1275 1.70567
R12259 GNDA.n1287 GNDA.n1274 1.70567
R12260 GNDA.n1287 GNDA.n1273 1.70567
R12261 GNDA.n1287 GNDA.n1272 1.70567
R12262 GNDA.n1287 GNDA.n1271 1.70567
R12263 GNDA.n2580 GNDA.n1336 1.70567
R12264 GNDA.n1319 GNDA.n1269 1.70567
R12265 GNDA.n1269 GNDA.n1268 1.70567
R12266 GNDA.n1269 GNDA.n1267 1.70567
R12267 GNDA.n1269 GNDA.n1266 1.70567
R12268 GNDA.n1269 GNDA.n1265 1.70567
R12269 GNDA.n1269 GNDA.n1264 1.70567
R12270 GNDA.n1269 GNDA.n1263 1.70567
R12271 GNDA.n1269 GNDA.n1262 1.70567
R12272 GNDA.n1269 GNDA.n1261 1.70567
R12273 GNDA.n1269 GNDA.n1260 1.70567
R12274 GNDA.n1269 GNDA.n1259 1.70567
R12275 GNDA.n1269 GNDA.n1258 1.70567
R12276 GNDA.n1269 GNDA.n1257 1.70567
R12277 GNDA.n1269 GNDA.n1256 1.70567
R12278 GNDA.n1269 GNDA.n1255 1.70567
R12279 GNDA.n1269 GNDA.n1254 1.70567
R12280 GNDA.n1288 GNDA.n1270 1.70567
R12281 GNDA.n2580 GNDA.n1335 1.70567
R12282 GNDA.n1290 GNDA.n1270 1.70567
R12283 GNDA.n2580 GNDA.n1334 1.70567
R12284 GNDA.n1292 GNDA.n1270 1.70567
R12285 GNDA.n2580 GNDA.n1333 1.70567
R12286 GNDA.n1294 GNDA.n1270 1.70567
R12287 GNDA.n2580 GNDA.n1332 1.70567
R12288 GNDA.n1296 GNDA.n1270 1.70567
R12289 GNDA.n2580 GNDA.n1331 1.70567
R12290 GNDA.n1298 GNDA.n1270 1.70567
R12291 GNDA.n2580 GNDA.n1330 1.70567
R12292 GNDA.n1300 GNDA.n1270 1.70567
R12293 GNDA.n2580 GNDA.n1329 1.70567
R12294 GNDA.n1302 GNDA.n1270 1.70567
R12295 GNDA.n2580 GNDA.n1328 1.70567
R12296 GNDA.n1304 GNDA.n1270 1.70567
R12297 GNDA.n2580 GNDA.n1327 1.70567
R12298 GNDA.n1306 GNDA.n1270 1.70567
R12299 GNDA.n2580 GNDA.n1326 1.70567
R12300 GNDA.n1308 GNDA.n1270 1.70567
R12301 GNDA.n2580 GNDA.n1325 1.70567
R12302 GNDA.n1310 GNDA.n1270 1.70567
R12303 GNDA.n2580 GNDA.n1324 1.70567
R12304 GNDA.n1312 GNDA.n1270 1.70567
R12305 GNDA.n2580 GNDA.n1323 1.70567
R12306 GNDA.n1314 GNDA.n1270 1.70567
R12307 GNDA.n2580 GNDA.n1322 1.70567
R12308 GNDA.n1316 GNDA.n1270 1.70567
R12309 GNDA.n2580 GNDA.n1321 1.70567
R12310 GNDA.n1318 GNDA.n1270 1.70567
R12311 GNDA.n2581 GNDA.n2580 1.70567
R12312 GNDA.n2584 GNDA.n1221 1.70567
R12313 GNDA.n1270 GNDA.n1205 1.70567
R12314 GNDA.n2690 GNDA.n1058 1.70567
R12315 GNDA.n2690 GNDA.n2671 1.70567
R12316 GNDA.n2690 GNDA.n2670 1.70567
R12317 GNDA.n2690 GNDA.n2669 1.70567
R12318 GNDA.n2690 GNDA.n2668 1.70567
R12319 GNDA.n2690 GNDA.n2667 1.70567
R12320 GNDA.n2690 GNDA.n2666 1.70567
R12321 GNDA.n2690 GNDA.n2665 1.70567
R12322 GNDA.n2690 GNDA.n2664 1.70567
R12323 GNDA.n2690 GNDA.n2663 1.70567
R12324 GNDA.n2690 GNDA.n2662 1.70567
R12325 GNDA.n2690 GNDA.n2661 1.70567
R12326 GNDA.n2690 GNDA.n2660 1.70567
R12327 GNDA.n2690 GNDA.n2659 1.70567
R12328 GNDA.n2690 GNDA.n2658 1.70567
R12329 GNDA.n2690 GNDA.n2657 1.70567
R12330 GNDA.n1091 GNDA.n1057 1.70567
R12331 GNDA.n1093 GNDA.n1057 1.70567
R12332 GNDA.n1095 GNDA.n1057 1.70567
R12333 GNDA.n1097 GNDA.n1057 1.70567
R12334 GNDA.n1099 GNDA.n1057 1.70567
R12335 GNDA.n1101 GNDA.n1057 1.70567
R12336 GNDA.n1103 GNDA.n1057 1.70567
R12337 GNDA.n1105 GNDA.n1057 1.70567
R12338 GNDA.n1107 GNDA.n1057 1.70567
R12339 GNDA.n1109 GNDA.n1057 1.70567
R12340 GNDA.n1111 GNDA.n1057 1.70567
R12341 GNDA.n1113 GNDA.n1057 1.70567
R12342 GNDA.n1115 GNDA.n1057 1.70567
R12343 GNDA.n1117 GNDA.n1057 1.70567
R12344 GNDA.n1119 GNDA.n1057 1.70567
R12345 GNDA.n2656 GNDA.n1138 1.70567
R12346 GNDA.n2688 GNDA.n2672 1.70567
R12347 GNDA.n1138 GNDA.n1137 1.70567
R12348 GNDA.n2688 GNDA.n2673 1.70567
R12349 GNDA.n1138 GNDA.n1136 1.70567
R12350 GNDA.n2688 GNDA.n2674 1.70567
R12351 GNDA.n1138 GNDA.n1135 1.70567
R12352 GNDA.n2688 GNDA.n2675 1.70567
R12353 GNDA.n1138 GNDA.n1134 1.70567
R12354 GNDA.n2688 GNDA.n2676 1.70567
R12355 GNDA.n1138 GNDA.n1133 1.70567
R12356 GNDA.n2688 GNDA.n2677 1.70567
R12357 GNDA.n1138 GNDA.n1132 1.70567
R12358 GNDA.n2688 GNDA.n2678 1.70567
R12359 GNDA.n1138 GNDA.n1131 1.70567
R12360 GNDA.n2688 GNDA.n2679 1.70567
R12361 GNDA.n1138 GNDA.n1130 1.70567
R12362 GNDA.n2688 GNDA.n2680 1.70567
R12363 GNDA.n1138 GNDA.n1129 1.70567
R12364 GNDA.n2688 GNDA.n2681 1.70567
R12365 GNDA.n1138 GNDA.n1128 1.70567
R12366 GNDA.n2688 GNDA.n2682 1.70567
R12367 GNDA.n1138 GNDA.n1127 1.70567
R12368 GNDA.n2688 GNDA.n2683 1.70567
R12369 GNDA.n1138 GNDA.n1126 1.70567
R12370 GNDA.n2688 GNDA.n2684 1.70567
R12371 GNDA.n1138 GNDA.n1125 1.70567
R12372 GNDA.n2688 GNDA.n2685 1.70567
R12373 GNDA.n1138 GNDA.n1124 1.70567
R12374 GNDA.n2688 GNDA.n2686 1.70567
R12375 GNDA.n1138 GNDA.n1123 1.70567
R12376 GNDA.n2688 GNDA.n2687 1.70567
R12377 GNDA.n1138 GNDA.n1122 1.70567
R12378 GNDA.n2688 GNDA.n1075 1.70567
R12379 GNDA.n2692 GNDA.n1121 1.70567
R12380 GNDA.n2601 GNDA.n1156 1.70567
R12381 GNDA.n2602 GNDA.n2600 1.70567
R12382 GNDA.n2602 GNDA.n2599 1.70567
R12383 GNDA.n2602 GNDA.n2598 1.70567
R12384 GNDA.n2602 GNDA.n2597 1.70567
R12385 GNDA.n2602 GNDA.n2596 1.70567
R12386 GNDA.n2602 GNDA.n2595 1.70567
R12387 GNDA.n2602 GNDA.n2594 1.70567
R12388 GNDA.n2602 GNDA.n2593 1.70567
R12389 GNDA.n2602 GNDA.n2592 1.70567
R12390 GNDA.n2602 GNDA.n2591 1.70567
R12391 GNDA.n2602 GNDA.n2590 1.70567
R12392 GNDA.n2602 GNDA.n2589 1.70567
R12393 GNDA.n2602 GNDA.n2588 1.70567
R12394 GNDA.n2602 GNDA.n2587 1.70567
R12395 GNDA.n2602 GNDA.n2586 1.70567
R12396 GNDA.n2602 GNDA.n2585 1.70567
R12397 GNDA.n2603 GNDA.n2602 1.70567
R12398 GNDA.n1204 GNDA.n1203 1.70567
R12399 GNDA.n1204 GNDA.n1202 1.70567
R12400 GNDA.n1204 GNDA.n1201 1.70567
R12401 GNDA.n1204 GNDA.n1200 1.70567
R12402 GNDA.n1204 GNDA.n1199 1.70567
R12403 GNDA.n1204 GNDA.n1198 1.70567
R12404 GNDA.n1204 GNDA.n1197 1.70567
R12405 GNDA.n1204 GNDA.n1196 1.70567
R12406 GNDA.n1204 GNDA.n1195 1.70567
R12407 GNDA.n1204 GNDA.n1194 1.70567
R12408 GNDA.n1204 GNDA.n1193 1.70567
R12409 GNDA.n1204 GNDA.n1192 1.70567
R12410 GNDA.n1204 GNDA.n1191 1.70567
R12411 GNDA.n1204 GNDA.n1190 1.70567
R12412 GNDA.n1204 GNDA.n1189 1.70567
R12413 GNDA.n2606 GNDA.n2605 1.70567
R12414 GNDA.n2650 GNDA.n2635 1.70567
R12415 GNDA.n2604 GNDA.n1140 1.70567
R12416 GNDA.n2650 GNDA.n2636 1.70567
R12417 GNDA.n2607 GNDA.n1140 1.70567
R12418 GNDA.n2650 GNDA.n2637 1.70567
R12419 GNDA.n2609 GNDA.n1140 1.70567
R12420 GNDA.n2650 GNDA.n2638 1.70567
R12421 GNDA.n2611 GNDA.n1140 1.70567
R12422 GNDA.n2650 GNDA.n2639 1.70567
R12423 GNDA.n2613 GNDA.n1140 1.70567
R12424 GNDA.n2650 GNDA.n2640 1.70567
R12425 GNDA.n2615 GNDA.n1140 1.70567
R12426 GNDA.n2650 GNDA.n2641 1.70567
R12427 GNDA.n2617 GNDA.n1140 1.70567
R12428 GNDA.n2650 GNDA.n2642 1.70567
R12429 GNDA.n2619 GNDA.n1140 1.70567
R12430 GNDA.n2650 GNDA.n2643 1.70567
R12431 GNDA.n2621 GNDA.n1140 1.70567
R12432 GNDA.n2650 GNDA.n2644 1.70567
R12433 GNDA.n2623 GNDA.n1140 1.70567
R12434 GNDA.n2650 GNDA.n2645 1.70567
R12435 GNDA.n2625 GNDA.n1140 1.70567
R12436 GNDA.n2650 GNDA.n2646 1.70567
R12437 GNDA.n2627 GNDA.n1140 1.70567
R12438 GNDA.n2650 GNDA.n2647 1.70567
R12439 GNDA.n2629 GNDA.n1140 1.70567
R12440 GNDA.n2650 GNDA.n2648 1.70567
R12441 GNDA.n2631 GNDA.n1140 1.70567
R12442 GNDA.n2650 GNDA.n2649 1.70567
R12443 GNDA.n2633 GNDA.n1140 1.70567
R12444 GNDA.n2651 GNDA.n2650 1.70567
R12445 GNDA.n2652 GNDA.n1140 1.70567
R12446 GNDA.n2650 GNDA.n1139 1.70567
R12447 GNDA.n3336 GNDA.n2702 1.69433
R12448 GNDA.n3336 GNDA.n2699 1.69433
R12449 GNDA.n3336 GNDA.n2696 1.69433
R12450 GNDA.n3271 GNDA.n2714 1.69433
R12451 GNDA.n3271 GNDA.n2711 1.69433
R12452 GNDA.n3271 GNDA.n2708 1.69433
R12453 GNDA.n3202 GNDA.n2726 1.69433
R12454 GNDA.n3202 GNDA.n2723 1.69433
R12455 GNDA.n3202 GNDA.n2720 1.69433
R12456 GNDA.n3133 GNDA.n2738 1.69433
R12457 GNDA.n3133 GNDA.n2735 1.69433
R12458 GNDA.n3133 GNDA.n2732 1.69433
R12459 GNDA.n3064 GNDA.n2750 1.69433
R12460 GNDA.n3064 GNDA.n2747 1.69433
R12461 GNDA.n3064 GNDA.n2744 1.69433
R12462 GNDA.n2995 GNDA.n2762 1.69433
R12463 GNDA.n2995 GNDA.n2759 1.69433
R12464 GNDA.n2995 GNDA.n2756 1.69433
R12465 GNDA.n2926 GNDA.n2774 1.69433
R12466 GNDA.n2926 GNDA.n2771 1.69433
R12467 GNDA.n2926 GNDA.n2768 1.69433
R12468 GNDA.n2857 GNDA.n2786 1.69433
R12469 GNDA.n2857 GNDA.n2783 1.69433
R12470 GNDA.n2857 GNDA.n2780 1.69433
R12471 GNDA.n3536 GNDA.n949 1.69433
R12472 GNDA.n3536 GNDA.n946 1.69433
R12473 GNDA.n3536 GNDA.n943 1.69433
R12474 GNDA.n3856 GNDA.n3627 1.69433
R12475 GNDA.n3856 GNDA.n3624 1.69433
R12476 GNDA.n3856 GNDA.n3621 1.69433
R12477 GNDA.n3791 GNDA.n3639 1.69433
R12478 GNDA.n3791 GNDA.n3636 1.69433
R12479 GNDA.n3791 GNDA.n3633 1.69433
R12480 GNDA.n3722 GNDA.n3651 1.69433
R12481 GNDA.n3722 GNDA.n3648 1.69433
R12482 GNDA.n3722 GNDA.n3645 1.69433
R12483 GNDA.n876 GNDA.n802 1.69433
R12484 GNDA.n865 GNDA.n802 1.69433
R12485 GNDA.n852 GNDA.n802 1.69433
R12486 GNDA.n3934 GNDA.n812 1.69433
R12487 GNDA.n3934 GNDA.n809 1.69433
R12488 GNDA.n3934 GNDA.n806 1.69433
R12489 GNDA.n3430 GNDA.n939 1.69433
R12490 GNDA.n3419 GNDA.n939 1.69433
R12491 GNDA.n3406 GNDA.n939 1.69433
R12492 GNDA.n3618 GNDA.n3546 1.69433
R12493 GNDA.n3618 GNDA.n3543 1.69433
R12494 GNDA.n3618 GNDA.n3540 1.69433
R12495 GNDA.n3951 GNDA.n3947 1.69433
R12496 GNDA.n3951 GNDA.n3943 1.69433
R12497 GNDA.n3951 GNDA.n3938 1.69433
R12498 GNDA.n4195 GNDA.n496 1.69433
R12499 GNDA.n4195 GNDA.n493 1.69433
R12500 GNDA.n4195 GNDA.n490 1.69433
R12501 GNDA.n4336 GNDA.n446 1.69433
R12502 GNDA.n4345 GNDA.n446 1.69433
R12503 GNDA.n4354 GNDA.n446 1.69433
R12504 GNDA.n4432 GNDA.n456 1.69433
R12505 GNDA.n4432 GNDA.n453 1.69433
R12506 GNDA.n4432 GNDA.n450 1.69433
R12507 GNDA.n4872 GNDA.n4441 1.69433
R12508 GNDA.n4872 GNDA.n4438 1.69433
R12509 GNDA.n4872 GNDA.n4435 1.69433
R12510 GNDA.n4271 GNDA.n4204 1.69433
R12511 GNDA.n4271 GNDA.n4201 1.69433
R12512 GNDA.n4271 GNDA.n4198 1.69433
R12513 GNDA.n4807 GNDA.n4453 1.69433
R12514 GNDA.n4807 GNDA.n4450 1.69433
R12515 GNDA.n4807 GNDA.n4447 1.69433
R12516 GNDA.n4524 GNDA.n4456 1.69433
R12517 GNDA.n4533 GNDA.n4456 1.69433
R12518 GNDA.n4542 GNDA.n4456 1.69433
R12519 GNDA.n4647 GNDA.n4575 1.69433
R12520 GNDA.n4647 GNDA.n4572 1.69433
R12521 GNDA.n4647 GNDA.n4569 1.69433
R12522 GNDA.n4723 GNDA.n4656 1.69433
R12523 GNDA.n4723 GNDA.n4653 1.69433
R12524 GNDA.n4723 GNDA.n4650 1.69433
R12525 GNDA.n2579 GNDA.n1346 1.69433
R12526 GNDA.n2579 GNDA.n1343 1.69433
R12527 GNDA.n2579 GNDA.n1340 1.69433
R12528 GNDA.n1532 GNDA.n1349 1.69433
R12529 GNDA.n1514 GNDA.n1349 1.69433
R12530 GNDA.n1502 GNDA.n1349 1.69433
R12531 GNDA.n552 GNDA.n486 1.69337
R12532 GNDA.n547 GNDA.n486 1.69337
R12533 GNDA.n539 GNDA.n486 1.69337
R12534 GNDA.n536 GNDA.n486 1.69337
R12535 GNDA.n528 GNDA.n486 1.69337
R12536 GNDA.n523 GNDA.n486 1.69337
R12537 GNDA.n515 GNDA.n486 1.69337
R12538 GNDA.n558 GNDA.n486 1.69337
R12539 GNDA.n3336 GNDA.n2704 1.6924
R12540 GNDA.n3336 GNDA.n2703 1.6924
R12541 GNDA.n3336 GNDA.n2701 1.6924
R12542 GNDA.n3336 GNDA.n2700 1.6924
R12543 GNDA.n3336 GNDA.n2698 1.6924
R12544 GNDA.n3336 GNDA.n2697 1.6924
R12545 GNDA.n3336 GNDA.n2695 1.6924
R12546 GNDA.n3336 GNDA.n2694 1.6924
R12547 GNDA.n3271 GNDA.n2716 1.6924
R12548 GNDA.n3271 GNDA.n2715 1.6924
R12549 GNDA.n3271 GNDA.n2713 1.6924
R12550 GNDA.n3271 GNDA.n2712 1.6924
R12551 GNDA.n3271 GNDA.n2710 1.6924
R12552 GNDA.n3271 GNDA.n2709 1.6924
R12553 GNDA.n3271 GNDA.n2707 1.6924
R12554 GNDA.n3271 GNDA.n2706 1.6924
R12555 GNDA.n3202 GNDA.n2728 1.6924
R12556 GNDA.n3202 GNDA.n2727 1.6924
R12557 GNDA.n3202 GNDA.n2725 1.6924
R12558 GNDA.n3202 GNDA.n2724 1.6924
R12559 GNDA.n3202 GNDA.n2722 1.6924
R12560 GNDA.n3202 GNDA.n2721 1.6924
R12561 GNDA.n3202 GNDA.n2719 1.6924
R12562 GNDA.n3202 GNDA.n2718 1.6924
R12563 GNDA.n3133 GNDA.n2740 1.6924
R12564 GNDA.n3133 GNDA.n2739 1.6924
R12565 GNDA.n3133 GNDA.n2737 1.6924
R12566 GNDA.n3133 GNDA.n2736 1.6924
R12567 GNDA.n3133 GNDA.n2734 1.6924
R12568 GNDA.n3133 GNDA.n2733 1.6924
R12569 GNDA.n3133 GNDA.n2731 1.6924
R12570 GNDA.n3133 GNDA.n2730 1.6924
R12571 GNDA.n3064 GNDA.n2752 1.6924
R12572 GNDA.n3064 GNDA.n2751 1.6924
R12573 GNDA.n3064 GNDA.n2749 1.6924
R12574 GNDA.n3064 GNDA.n2748 1.6924
R12575 GNDA.n3064 GNDA.n2746 1.6924
R12576 GNDA.n3064 GNDA.n2745 1.6924
R12577 GNDA.n3064 GNDA.n2743 1.6924
R12578 GNDA.n3064 GNDA.n2742 1.6924
R12579 GNDA.n2995 GNDA.n2764 1.6924
R12580 GNDA.n2995 GNDA.n2763 1.6924
R12581 GNDA.n2995 GNDA.n2761 1.6924
R12582 GNDA.n2995 GNDA.n2760 1.6924
R12583 GNDA.n2995 GNDA.n2758 1.6924
R12584 GNDA.n2995 GNDA.n2757 1.6924
R12585 GNDA.n2995 GNDA.n2755 1.6924
R12586 GNDA.n2995 GNDA.n2754 1.6924
R12587 GNDA.n2926 GNDA.n2776 1.6924
R12588 GNDA.n2926 GNDA.n2775 1.6924
R12589 GNDA.n2926 GNDA.n2773 1.6924
R12590 GNDA.n2926 GNDA.n2772 1.6924
R12591 GNDA.n2926 GNDA.n2770 1.6924
R12592 GNDA.n2926 GNDA.n2769 1.6924
R12593 GNDA.n2926 GNDA.n2767 1.6924
R12594 GNDA.n2926 GNDA.n2766 1.6924
R12595 GNDA.n2857 GNDA.n2788 1.6924
R12596 GNDA.n2857 GNDA.n2787 1.6924
R12597 GNDA.n2857 GNDA.n2785 1.6924
R12598 GNDA.n2857 GNDA.n2784 1.6924
R12599 GNDA.n2857 GNDA.n2782 1.6924
R12600 GNDA.n2857 GNDA.n2781 1.6924
R12601 GNDA.n2857 GNDA.n2779 1.6924
R12602 GNDA.n2857 GNDA.n2778 1.6924
R12603 GNDA.n3536 GNDA.n951 1.6924
R12604 GNDA.n3536 GNDA.n950 1.6924
R12605 GNDA.n3536 GNDA.n948 1.6924
R12606 GNDA.n3536 GNDA.n947 1.6924
R12607 GNDA.n3536 GNDA.n945 1.6924
R12608 GNDA.n3536 GNDA.n944 1.6924
R12609 GNDA.n3536 GNDA.n942 1.6924
R12610 GNDA.n3536 GNDA.n941 1.6924
R12611 GNDA.n3856 GNDA.n3629 1.6924
R12612 GNDA.n3856 GNDA.n3628 1.6924
R12613 GNDA.n3856 GNDA.n3626 1.6924
R12614 GNDA.n3856 GNDA.n3625 1.6924
R12615 GNDA.n3856 GNDA.n3623 1.6924
R12616 GNDA.n3856 GNDA.n3622 1.6924
R12617 GNDA.n3856 GNDA.n3620 1.6924
R12618 GNDA.n3856 GNDA.n3619 1.6924
R12619 GNDA.n3791 GNDA.n3641 1.6924
R12620 GNDA.n3791 GNDA.n3640 1.6924
R12621 GNDA.n3791 GNDA.n3638 1.6924
R12622 GNDA.n3791 GNDA.n3637 1.6924
R12623 GNDA.n3791 GNDA.n3635 1.6924
R12624 GNDA.n3791 GNDA.n3634 1.6924
R12625 GNDA.n3791 GNDA.n3632 1.6924
R12626 GNDA.n3791 GNDA.n3631 1.6924
R12627 GNDA.n3722 GNDA.n3653 1.6924
R12628 GNDA.n3722 GNDA.n3652 1.6924
R12629 GNDA.n3722 GNDA.n3650 1.6924
R12630 GNDA.n3722 GNDA.n3649 1.6924
R12631 GNDA.n3722 GNDA.n3647 1.6924
R12632 GNDA.n3722 GNDA.n3646 1.6924
R12633 GNDA.n3722 GNDA.n3644 1.6924
R12634 GNDA.n3722 GNDA.n3643 1.6924
R12635 GNDA.n884 GNDA.n802 1.6924
R12636 GNDA.n881 GNDA.n802 1.6924
R12637 GNDA.n873 GNDA.n802 1.6924
R12638 GNDA.n868 GNDA.n802 1.6924
R12639 GNDA.n860 GNDA.n802 1.6924
R12640 GNDA.n857 GNDA.n802 1.6924
R12641 GNDA.n849 GNDA.n802 1.6924
R12642 GNDA.n844 GNDA.n802 1.6924
R12643 GNDA.n3934 GNDA.n814 1.6924
R12644 GNDA.n3934 GNDA.n813 1.6924
R12645 GNDA.n3934 GNDA.n811 1.6924
R12646 GNDA.n3934 GNDA.n810 1.6924
R12647 GNDA.n3934 GNDA.n808 1.6924
R12648 GNDA.n3934 GNDA.n807 1.6924
R12649 GNDA.n3934 GNDA.n805 1.6924
R12650 GNDA.n3934 GNDA.n804 1.6924
R12651 GNDA.n3438 GNDA.n939 1.6924
R12652 GNDA.n3435 GNDA.n939 1.6924
R12653 GNDA.n3427 GNDA.n939 1.6924
R12654 GNDA.n3422 GNDA.n939 1.6924
R12655 GNDA.n3414 GNDA.n939 1.6924
R12656 GNDA.n3411 GNDA.n939 1.6924
R12657 GNDA.n3403 GNDA.n939 1.6924
R12658 GNDA.n3398 GNDA.n939 1.6924
R12659 GNDA.n3618 GNDA.n3548 1.6924
R12660 GNDA.n3618 GNDA.n3547 1.6924
R12661 GNDA.n3618 GNDA.n3545 1.6924
R12662 GNDA.n3618 GNDA.n3544 1.6924
R12663 GNDA.n3618 GNDA.n3542 1.6924
R12664 GNDA.n3618 GNDA.n3541 1.6924
R12665 GNDA.n3618 GNDA.n3539 1.6924
R12666 GNDA.n3618 GNDA.n3538 1.6924
R12667 GNDA.n3951 GNDA.n3950 1.6924
R12668 GNDA.n3951 GNDA.n3949 1.6924
R12669 GNDA.n3951 GNDA.n3946 1.6924
R12670 GNDA.n3951 GNDA.n3944 1.6924
R12671 GNDA.n3951 GNDA.n3941 1.6924
R12672 GNDA.n3951 GNDA.n3940 1.6924
R12673 GNDA.n3951 GNDA.n3937 1.6924
R12674 GNDA.n3951 GNDA.n3935 1.6924
R12675 GNDA.n4195 GNDA.n498 1.6924
R12676 GNDA.n4195 GNDA.n497 1.6924
R12677 GNDA.n4195 GNDA.n495 1.6924
R12678 GNDA.n4195 GNDA.n494 1.6924
R12679 GNDA.n4195 GNDA.n492 1.6924
R12680 GNDA.n4195 GNDA.n491 1.6924
R12681 GNDA.n4195 GNDA.n489 1.6924
R12682 GNDA.n4195 GNDA.n488 1.6924
R12683 GNDA.n4330 GNDA.n446 1.6924
R12684 GNDA.n4333 GNDA.n446 1.6924
R12685 GNDA.n4339 GNDA.n446 1.6924
R12686 GNDA.n4342 GNDA.n446 1.6924
R12687 GNDA.n4348 GNDA.n446 1.6924
R12688 GNDA.n4351 GNDA.n446 1.6924
R12689 GNDA.n4357 GNDA.n446 1.6924
R12690 GNDA.n4360 GNDA.n446 1.6924
R12691 GNDA.n4432 GNDA.n458 1.6924
R12692 GNDA.n4432 GNDA.n457 1.6924
R12693 GNDA.n4432 GNDA.n455 1.6924
R12694 GNDA.n4432 GNDA.n454 1.6924
R12695 GNDA.n4432 GNDA.n452 1.6924
R12696 GNDA.n4432 GNDA.n451 1.6924
R12697 GNDA.n4432 GNDA.n449 1.6924
R12698 GNDA.n4432 GNDA.n448 1.6924
R12699 GNDA.n4872 GNDA.n4443 1.6924
R12700 GNDA.n4872 GNDA.n4442 1.6924
R12701 GNDA.n4872 GNDA.n4440 1.6924
R12702 GNDA.n4872 GNDA.n4439 1.6924
R12703 GNDA.n4872 GNDA.n4437 1.6924
R12704 GNDA.n4872 GNDA.n4436 1.6924
R12705 GNDA.n4872 GNDA.n4434 1.6924
R12706 GNDA.n4872 GNDA.n4433 1.6924
R12707 GNDA.n4271 GNDA.n4206 1.6924
R12708 GNDA.n4271 GNDA.n4205 1.6924
R12709 GNDA.n4271 GNDA.n4203 1.6924
R12710 GNDA.n4271 GNDA.n4202 1.6924
R12711 GNDA.n4271 GNDA.n4200 1.6924
R12712 GNDA.n4271 GNDA.n4199 1.6924
R12713 GNDA.n4271 GNDA.n4197 1.6924
R12714 GNDA.n4271 GNDA.n4196 1.6924
R12715 GNDA.n4807 GNDA.n4455 1.6924
R12716 GNDA.n4807 GNDA.n4454 1.6924
R12717 GNDA.n4807 GNDA.n4452 1.6924
R12718 GNDA.n4807 GNDA.n4451 1.6924
R12719 GNDA.n4807 GNDA.n4449 1.6924
R12720 GNDA.n4807 GNDA.n4448 1.6924
R12721 GNDA.n4807 GNDA.n4446 1.6924
R12722 GNDA.n4807 GNDA.n4445 1.6924
R12723 GNDA.n4518 GNDA.n4456 1.6924
R12724 GNDA.n4521 GNDA.n4456 1.6924
R12725 GNDA.n4527 GNDA.n4456 1.6924
R12726 GNDA.n4530 GNDA.n4456 1.6924
R12727 GNDA.n4536 GNDA.n4456 1.6924
R12728 GNDA.n4539 GNDA.n4456 1.6924
R12729 GNDA.n4545 GNDA.n4456 1.6924
R12730 GNDA.n4548 GNDA.n4456 1.6924
R12731 GNDA.n4647 GNDA.n4577 1.6924
R12732 GNDA.n4647 GNDA.n4576 1.6924
R12733 GNDA.n4647 GNDA.n4574 1.6924
R12734 GNDA.n4647 GNDA.n4573 1.6924
R12735 GNDA.n4647 GNDA.n4571 1.6924
R12736 GNDA.n4647 GNDA.n4570 1.6924
R12737 GNDA.n4647 GNDA.n4568 1.6924
R12738 GNDA.n4647 GNDA.n4567 1.6924
R12739 GNDA.n4723 GNDA.n4658 1.6924
R12740 GNDA.n4723 GNDA.n4657 1.6924
R12741 GNDA.n4723 GNDA.n4655 1.6924
R12742 GNDA.n4723 GNDA.n4654 1.6924
R12743 GNDA.n4723 GNDA.n4652 1.6924
R12744 GNDA.n4723 GNDA.n4651 1.6924
R12745 GNDA.n4723 GNDA.n4649 1.6924
R12746 GNDA.n4723 GNDA.n4648 1.6924
R12747 GNDA.n2579 GNDA.n1348 1.6924
R12748 GNDA.n2579 GNDA.n1347 1.6924
R12749 GNDA.n2579 GNDA.n1345 1.6924
R12750 GNDA.n2579 GNDA.n1344 1.6924
R12751 GNDA.n2579 GNDA.n1342 1.6924
R12752 GNDA.n2579 GNDA.n1341 1.6924
R12753 GNDA.n2579 GNDA.n1339 1.6924
R12754 GNDA.n2579 GNDA.n1338 1.6924
R12755 GNDA.n1542 GNDA.n1349 1.6924
R12756 GNDA.n1534 GNDA.n1349 1.6924
R12757 GNDA.n1524 GNDA.n1349 1.6924
R12758 GNDA.n1522 GNDA.n1349 1.6924
R12759 GNDA.n1512 GNDA.n1349 1.6924
R12760 GNDA.n1504 GNDA.n1349 1.6924
R12761 GNDA.n1494 GNDA.n1349 1.6924
R12762 GNDA.n1492 GNDA.n1349 1.6924
R12763 GNDA.n555 GNDA.n486 1.6924
R12764 GNDA.n544 GNDA.n486 1.6924
R12765 GNDA.n531 GNDA.n486 1.6924
R12766 GNDA.n520 GNDA.n486 1.6924
R12767 GNDA.n4090 GNDA.n4089 1.65675
R12768 GNDA.n4092 GNDA.n4091 1.65675
R12769 GNDA.n4043 GNDA.n4016 1.56997
R12770 GNDA.n4018 GNDA.n4017 1.56997
R12771 GNDA.t152 GNDA.n105 1.51652
R12772 GNDA.n3477 GNDA.n3394 1.5005
R12773 GNDA.n4136 GNDA.n481 1.5005
R12774 GNDA.n2539 GNDA.n2538 1.47392
R12775 GNDA.n2306 GNDA.n2305 1.47392
R12776 GNDA.n5153 GNDA.n228 1.47392
R12777 GNDA.n5130 GNDA.n5127 1.47392
R12778 GNDA.n1855 GNDA.n1853 1.47392
R12779 GNDA.n5376 GNDA.n87 1.47392
R12780 GNDA.n709 GNDA.n708 1.44719
R12781 GNDA.n720 GNDA.n719 1.44719
R12782 GNDA.n1462 GNDA.n1461 1.22446
R12783 GNDA.n4900 GNDA.n4899 1.15154
R12784 GNDA.n1011 GNDA.n1010 1.15154
R12785 GNDA.n4101 GNDA.n4086 1.13592
R12786 GNDA.n4104 GNDA.n4103 1.13592
R12787 GNDA.n4912 GNDA.n4911 1.09425
R12788 GNDA.n995 GNDA.n630 1.09425
R12789 GNDA.n4907 GNDA.n4906 1.07342
R12790 GNDA.n1018 GNDA.n1016 1.06821
R12791 GNDA.n709 GNDA.n706 1.063
R12792 GNDA.n719 GNDA.n718 1.063
R12793 GNDA.n2566 GNDA.n2565 1.05258
R12794 GNDA.n4106 GNDA.n614 0.984875
R12795 GNDA.n4082 GNDA.n4081 0.984875
R12796 GNDA.n4007 GNDA.n4006 0.975928
R12797 GNDA.n3996 GNDA.n3995 0.975928
R12798 GNDA.n1550 GNDA.n1463 0.854667
R12799 GNDA.n2499 GNDA.n2498 0.8197
R12800 GNDA.n2485 GNDA.n1598 0.8197
R12801 GNDA.n2492 GNDA.n2486 0.8197
R12802 GNDA.n2491 GNDA.n2488 0.8197
R12803 GNDA.n2504 GNDA.n1566 0.8197
R12804 GNDA.n1577 GNDA.n1573 0.8197
R12805 GNDA.n1579 GNDA.n1578 0.8197
R12806 GNDA.n2542 GNDA.n1448 0.8197
R12807 GNDA.n2005 GNDA.n1933 0.8197
R12808 GNDA.n2004 GNDA.n1934 0.8197
R12809 GNDA.n2012 GNDA.n1909 0.8197
R12810 GNDA.n2014 GNDA.n2013 0.8197
R12811 GNDA.n2020 GNDA.n1906 0.8197
R12812 GNDA.n2028 GNDA.n1903 0.8197
R12813 GNDA.n2030 GNDA.n2029 0.8197
R12814 GNDA.n2038 GNDA.n1899 0.8197
R12815 GNDA.n5334 GNDA.n165 0.8197
R12816 GNDA.n5333 GNDA.n167 0.8197
R12817 GNDA.n218 GNDA.n200 0.8197
R12818 GNDA.n217 GNDA.n215 0.8197
R12819 GNDA.n211 GNDA.n210 0.8197
R12820 GNDA.n207 GNDA.n203 0.8197
R12821 GNDA.n206 GNDA.n187 0.8197
R12822 GNDA.n5275 GNDA.n5274 0.8197
R12823 GNDA.n2290 GNDA.n2289 0.8197
R12824 GNDA.n2286 GNDA.n2285 0.8197
R12825 GNDA.n2282 GNDA.n2266 0.8197
R12826 GNDA.n2281 GNDA.n2278 0.8197
R12827 GNDA.n2274 GNDA.n2271 0.8197
R12828 GNDA.n2268 GNDA.n2190 0.8197
R12829 GNDA.n2296 GNDA.n2295 0.8197
R12830 GNDA.n2299 GNDA.n2189 0.8197
R12831 GNDA.n5265 GNDA.n5156 0.8197
R12832 GNDA.n5262 GNDA.n5261 0.8197
R12833 GNDA.n5258 GNDA.n5159 0.8197
R12834 GNDA.n5257 GNDA.n5160 0.8197
R12835 GNDA.n5192 GNDA.n5189 0.8197
R12836 GNDA.n5193 GNDA.n5183 0.8197
R12837 GNDA.n5197 GNDA.n5196 0.8197
R12838 GNDA.n5201 GNDA.n5200 0.8197
R12839 GNDA.n5544 GNDA.n59 0.8197
R12840 GNDA.n5541 GNDA.n5540 0.8197
R12841 GNDA.n5537 GNDA.n62 0.8197
R12842 GNDA.n5536 GNDA.n63 0.8197
R12843 GNDA.n5471 GNDA.n5468 0.8197
R12844 GNDA.n5472 GNDA.n5462 0.8197
R12845 GNDA.n5476 GNDA.n5475 0.8197
R12846 GNDA.n5480 GNDA.n5479 0.8197
R12847 GNDA.n5119 GNDA.n5011 0.8197
R12848 GNDA.n5118 GNDA.n5012 0.8197
R12849 GNDA.n5038 GNDA.n5035 0.8197
R12850 GNDA.n5041 GNDA.n5040 0.8197
R12851 GNDA.n5051 GNDA.n5048 0.8197
R12852 GNDA.n5052 GNDA.n5034 0.8197
R12853 GNDA.n5056 GNDA.n5055 0.8197
R12854 GNDA.n5060 GNDA.n5059 0.8197
R12855 GNDA.n1858 GNDA.n1730 0.8197
R12856 GNDA.n1871 GNDA.n1870 0.8197
R12857 GNDA.n1728 GNDA.n1727 0.8197
R12858 GNDA.n1878 GNDA.n1877 0.8197
R12859 GNDA.n2072 GNDA.n2071 0.8197
R12860 GNDA.n1724 GNDA.n1723 0.8197
R12861 GNDA.n2080 GNDA.n1720 0.8197
R12862 GNDA.n2079 GNDA.n1721 0.8197
R12863 GNDA.n5554 GNDA.n5553 0.8197
R12864 GNDA.n32 GNDA.n23 0.8197
R12865 GNDA.n39 GNDA.n33 0.8197
R12866 GNDA.n38 GNDA.n35 0.8197
R12867 GNDA.n5559 GNDA.n1 0.8197
R12868 GNDA.n5391 GNDA.n5388 0.8197
R12869 GNDA.n5394 GNDA.n5393 0.8197
R12870 GNDA.n5398 GNDA.n5397 0.8197
R12871 GNDA.n3988 GNDA.n3987 0.808944
R12872 GNDA.n3571 GNDA.n935 0.808539
R12873 GNDA.n4727 GNDA.n4726 0.776542
R12874 GNDA.n4590 GNDA.n4558 0.776542
R12875 GNDA.n4553 GNDA.n4552 0.776542
R12876 GNDA.n4750 GNDA.n4749 0.776542
R12877 GNDA.n4876 GNDA.n4875 0.776542
R12878 GNDA.n4375 GNDA.n4374 0.776542
R12879 GNDA.n4365 GNDA.n4364 0.776542
R12880 GNDA.n3887 GNDA.n3886 0.776542
R12881 GNDA.n3879 GNDA.n921 0.776542
R12882 GNDA.n3874 GNDA.n925 0.776542
R12883 GNDA.n3869 GNDA.n929 0.776542
R12884 GNDA.n3860 GNDA.n3859 0.776542
R12885 GNDA.n3489 GNDA.n3488 0.776542
R12886 GNDA.n3373 GNDA.n987 0.776542
R12887 GNDA.n3368 GNDA.n991 0.776542
R12888 GNDA.n3358 GNDA.n1026 0.776542
R12889 GNDA.n3353 GNDA.n1030 0.776542
R12890 GNDA.n3348 GNDA.n1034 0.776542
R12891 GNDA.n3340 GNDA.n3339 0.776542
R12892 GNDA.n597 GNDA.n593 0.776542
R12893 GNDA.n2052 GNDA.n2051 0.776542
R12894 GNDA.n3378 GNDA.n983 0.776542
R12895 GNDA.n4275 GNDA.n4274 0.77295
R12896 GNDA.n3392 GNDA.n979 0.77295
R12897 GNDA.n4138 GNDA.n4137 0.755708
R12898 GNDA.n3478 GNDA.n3475 0.755708
R12899 GNDA.n3479 GNDA.n3478 0.751386
R12900 GNDA.n4137 GNDA.n4134 0.751
R12901 GNDA.n2580 GNDA.n2579 0.723198
R12902 GNDA.n2573 GNDA.n2572 0.71925
R12903 GNDA.n4912 GNDA.n432 0.688
R12904 GNDA.n4070 GNDA.n630 0.688
R12905 GNDA.n2521 GNDA.n1555 0.65675
R12906 GNDA.n3336 GNDA.n2693 0.655048
R12907 GNDA.n3989 GNDA.n3988 0.577365
R12908 GNDA.n935 GNDA.n934 0.576819
R12909 GNDA.n3862 GNDA.n935 0.5696
R12910 GNDA.n3988 GNDA.n772 0.567414
R12911 GNDA.n2487 GNDA 0.5637
R12912 GNDA.n1907 GNDA 0.5637
R12913 GNDA.n214 GNDA 0.5637
R12914 GNDA GNDA.n2267 0.5637
R12915 GNDA GNDA.n5184 0.5637
R12916 GNDA GNDA.n5463 0.5637
R12917 GNDA.n5045 GNDA 0.5637
R12918 GNDA GNDA.n1879 0.5637
R12919 GNDA.n34 GNDA 0.5637
R12920 GNDA.n738 GNDA.n737 0.5005
R12921 GNDA.n736 GNDA.n735 0.5005
R12922 GNDA.n641 GNDA.n640 0.5005
R12923 GNDA.n639 GNDA.n638 0.5005
R12924 GNDA.n4049 GNDA.n4015 0.427583
R12925 GNDA.n769 GNDA.n749 0.427583
R12926 GNDA.n3992 GNDA.n770 0.40675
R12927 GNDA.n4011 GNDA.n4010 0.40675
R12928 GNDA.n654 GNDA.n432 0.40675
R12929 GNDA.n4071 GNDA.n4070 0.40675
R12930 GNDA.n5150 GNDA.n105 0.383687
R12931 GNDA.n4113 GNDA.n609 0.359875
R12932 GNDA.n702 GNDA.n701 0.359875
R12933 GNDA.n1463 GNDA.n1462 0.339042
R12934 GNDA.n3868 GNDA.n3865 0.28175
R12935 GNDA.n3873 GNDA.n3870 0.28175
R12936 GNDA.n3878 GNDA.n3875 0.28175
R12937 GNDA.n3885 GNDA.n3880 0.28175
R12938 GNDA.n3347 GNDA.n3344 0.28175
R12939 GNDA.n3352 GNDA.n3349 0.28175
R12940 GNDA.n3357 GNDA.n3354 0.28175
R12941 GNDA.n3372 GNDA.n3369 0.28175
R12942 GNDA.n3394 GNDA.n3393 0.28175
R12943 GNDA.n4277 GNDA.n481 0.28175
R12944 GNDA.n4371 GNDA.n4369 0.28175
R12945 GNDA.n4878 GNDA.n441 0.28175
R12946 GNDA.n4742 GNDA.n4741 0.28175
R12947 GNDA.n4738 GNDA.n4737 0.28175
R12948 GNDA.n4734 GNDA.n4733 0.28175
R12949 GNDA.n3386 GNDA.n3379 0.271333
R12950 GNDA.n2690 GNDA.n2655 0.258413
R12951 GNDA.n2505 GNDA 0.2565
R12952 GNDA.n2021 GNDA 0.2565
R12953 GNDA.n202 GNDA 0.2565
R12954 GNDA.n2275 GNDA 0.2565
R12955 GNDA.n5187 GNDA 0.2565
R12956 GNDA.n5466 GNDA 0.2565
R12957 GNDA GNDA.n5044 0.2565
R12958 GNDA.n1880 GNDA 0.2565
R12959 GNDA GNDA.n0 0.2565
R12960 GNDA.n665 GNDA.n624 0.229667
R12961 GNDA.n732 GNDA.n662 0.229667
R12962 GNDA.n695 GNDA.n694 0.229667
R12963 GNDA.n4116 GNDA.n4115 0.229667
R12964 GNDA.n4099 GNDA.n4098 0.214042
R12965 GNDA.n4110 GNDA.n4109 0.214042
R12966 GNDA.n4085 GNDA.n620 0.214042
R12967 GNDA.n2602 GNDA.n2584 0.213322
R12968 GNDA.n3377 GNDA.n3374 0.198417
R12969 GNDA.n3487 GNDA.n3482 0.198417
R12970 GNDA.n4133 GNDA.n598 0.198417
R12971 GNDA.n4367 GNDA.n4282 0.188
R12972 GNDA.n1923 GNDA.n1922 0.188
R12973 GNDA.n2049 GNDA.n2048 0.188
R12974 GNDA.n2557 GNDA.n2556 0.15675
R12975 GNDA.n2562 GNDA.n2561 0.151542
R12976 GNDA.n2552 GNDA.n2551 0.151542
R12977 GNDA.n2527 GNDA.n2526 0.147453
R12978 GNDA.n4670 GNDA.n4564 0.146333
R12979 GNDA.n4675 GNDA.n4670 0.146333
R12980 GNDA.n4676 GNDA.n4675 0.146333
R12981 GNDA.n4686 GNDA.n4685 0.146333
R12982 GNDA.n4689 GNDA.n4686 0.146333
R12983 GNDA.n4689 GNDA.n4666 0.146333
R12984 GNDA.n4699 GNDA.n4664 0.146333
R12985 GNDA.n4705 GNDA.n4664 0.146333
R12986 GNDA.n4706 GNDA.n4705 0.146333
R12987 GNDA.n4716 GNDA.n4715 0.146333
R12988 GNDA.n4719 GNDA.n4716 0.146333
R12989 GNDA.n4719 GNDA.n4660 0.146333
R12990 GNDA.n4593 GNDA.n4589 0.146333
R12991 GNDA.n4599 GNDA.n4589 0.146333
R12992 GNDA.n4600 GNDA.n4599 0.146333
R12993 GNDA.n4610 GNDA.n4609 0.146333
R12994 GNDA.n4613 GNDA.n4610 0.146333
R12995 GNDA.n4613 GNDA.n4585 0.146333
R12996 GNDA.n4623 GNDA.n4583 0.146333
R12997 GNDA.n4629 GNDA.n4583 0.146333
R12998 GNDA.n4630 GNDA.n4629 0.146333
R12999 GNDA.n4640 GNDA.n4639 0.146333
R13000 GNDA.n4643 GNDA.n4640 0.146333
R13001 GNDA.n4643 GNDA.n4579 0.146333
R13002 GNDA.n4474 GNDA.n4473 0.146333
R13003 GNDA.n4475 GNDA.n4474 0.146333
R13004 GNDA.n4476 GNDA.n4475 0.146333
R13005 GNDA.n4480 GNDA.n4479 0.146333
R13006 GNDA.n4481 GNDA.n4480 0.146333
R13007 GNDA.n4482 GNDA.n4481 0.146333
R13008 GNDA.n4486 GNDA.n4485 0.146333
R13009 GNDA.n4487 GNDA.n4486 0.146333
R13010 GNDA.n4488 GNDA.n4487 0.146333
R13011 GNDA.n4492 GNDA.n4491 0.146333
R13012 GNDA.n4493 GNDA.n4492 0.146333
R13013 GNDA.n4494 GNDA.n4493 0.146333
R13014 GNDA.n4753 GNDA.n4468 0.146333
R13015 GNDA.n4759 GNDA.n4468 0.146333
R13016 GNDA.n4760 GNDA.n4759 0.146333
R13017 GNDA.n4770 GNDA.n4769 0.146333
R13018 GNDA.n4773 GNDA.n4770 0.146333
R13019 GNDA.n4773 GNDA.n4464 0.146333
R13020 GNDA.n4783 GNDA.n4462 0.146333
R13021 GNDA.n4789 GNDA.n4462 0.146333
R13022 GNDA.n4790 GNDA.n4789 0.146333
R13023 GNDA.n4800 GNDA.n4799 0.146333
R13024 GNDA.n4803 GNDA.n4800 0.146333
R13025 GNDA.n4803 GNDA.n4458 0.146333
R13026 GNDA.n4218 GNDA.n484 0.146333
R13027 GNDA.n4223 GNDA.n4218 0.146333
R13028 GNDA.n4224 GNDA.n4223 0.146333
R13029 GNDA.n4234 GNDA.n4233 0.146333
R13030 GNDA.n4237 GNDA.n4234 0.146333
R13031 GNDA.n4237 GNDA.n4214 0.146333
R13032 GNDA.n4247 GNDA.n4212 0.146333
R13033 GNDA.n4253 GNDA.n4212 0.146333
R13034 GNDA.n4254 GNDA.n4253 0.146333
R13035 GNDA.n4264 GNDA.n4263 0.146333
R13036 GNDA.n4267 GNDA.n4264 0.146333
R13037 GNDA.n4267 GNDA.n4208 0.146333
R13038 GNDA.n4819 GNDA.n444 0.146333
R13039 GNDA.n4824 GNDA.n4819 0.146333
R13040 GNDA.n4825 GNDA.n4824 0.146333
R13041 GNDA.n4835 GNDA.n4834 0.146333
R13042 GNDA.n4838 GNDA.n4835 0.146333
R13043 GNDA.n4838 GNDA.n4815 0.146333
R13044 GNDA.n4848 GNDA.n4813 0.146333
R13045 GNDA.n4854 GNDA.n4813 0.146333
R13046 GNDA.n4855 GNDA.n4854 0.146333
R13047 GNDA.n4865 GNDA.n4864 0.146333
R13048 GNDA.n4868 GNDA.n4865 0.146333
R13049 GNDA.n4868 GNDA.n4809 0.146333
R13050 GNDA.n4378 GNDA.n470 0.146333
R13051 GNDA.n4384 GNDA.n470 0.146333
R13052 GNDA.n4385 GNDA.n4384 0.146333
R13053 GNDA.n4395 GNDA.n4394 0.146333
R13054 GNDA.n4398 GNDA.n4395 0.146333
R13055 GNDA.n4398 GNDA.n466 0.146333
R13056 GNDA.n4408 GNDA.n464 0.146333
R13057 GNDA.n4414 GNDA.n464 0.146333
R13058 GNDA.n4415 GNDA.n4414 0.146333
R13059 GNDA.n4425 GNDA.n4424 0.146333
R13060 GNDA.n4428 GNDA.n4425 0.146333
R13061 GNDA.n4428 GNDA.n460 0.146333
R13062 GNDA.n4286 GNDA.n4285 0.146333
R13063 GNDA.n4287 GNDA.n4286 0.146333
R13064 GNDA.n4288 GNDA.n4287 0.146333
R13065 GNDA.n4292 GNDA.n4291 0.146333
R13066 GNDA.n4293 GNDA.n4292 0.146333
R13067 GNDA.n4294 GNDA.n4293 0.146333
R13068 GNDA.n4298 GNDA.n4297 0.146333
R13069 GNDA.n4299 GNDA.n4298 0.146333
R13070 GNDA.n4300 GNDA.n4299 0.146333
R13071 GNDA.n4304 GNDA.n4303 0.146333
R13072 GNDA.n4305 GNDA.n4304 0.146333
R13073 GNDA.n4306 GNDA.n4305 0.146333
R13074 GNDA.n4141 GNDA.n510 0.146333
R13075 GNDA.n4147 GNDA.n510 0.146333
R13076 GNDA.n4148 GNDA.n4147 0.146333
R13077 GNDA.n4158 GNDA.n4157 0.146333
R13078 GNDA.n4161 GNDA.n4158 0.146333
R13079 GNDA.n4161 GNDA.n506 0.146333
R13080 GNDA.n4171 GNDA.n504 0.146333
R13081 GNDA.n4177 GNDA.n504 0.146333
R13082 GNDA.n4178 GNDA.n4177 0.146333
R13083 GNDA.n4188 GNDA.n4187 0.146333
R13084 GNDA.n4191 GNDA.n4188 0.146333
R13085 GNDA.n4191 GNDA.n500 0.146333
R13086 GNDA.n3985 GNDA.n3984 0.146333
R13087 GNDA.n3984 GNDA.n777 0.146333
R13088 GNDA.n3980 GNDA.n777 0.146333
R13089 GNDA.n3974 GNDA.n782 0.146333
R13090 GNDA.n3974 GNDA.n3973 0.146333
R13091 GNDA.n3973 GNDA.n3972 0.146333
R13092 GNDA.n3967 GNDA.n3966 0.146333
R13093 GNDA.n3966 GNDA.n792 0.146333
R13094 GNDA.n3962 GNDA.n792 0.146333
R13095 GNDA.n3956 GNDA.n797 0.146333
R13096 GNDA.n3956 GNDA.n3955 0.146333
R13097 GNDA.n3955 GNDA.n3954 0.146333
R13098 GNDA.n3574 GNDA.n3568 0.146333
R13099 GNDA.n3578 GNDA.n3568 0.146333
R13100 GNDA.n3579 GNDA.n3578 0.146333
R13101 GNDA.n3587 GNDA.n3586 0.146333
R13102 GNDA.n3590 GNDA.n3587 0.146333
R13103 GNDA.n3590 GNDA.n3560 0.146333
R13104 GNDA.n3598 GNDA.n3556 0.146333
R13105 GNDA.n3602 GNDA.n3556 0.146333
R13106 GNDA.n3603 GNDA.n3602 0.146333
R13107 GNDA.n3611 GNDA.n3610 0.146333
R13108 GNDA.n3614 GNDA.n3611 0.146333
R13109 GNDA.n3614 GNDA.n3550 0.146333
R13110 GNDA.n3890 GNDA.n834 0.146333
R13111 GNDA.n3894 GNDA.n834 0.146333
R13112 GNDA.n3895 GNDA.n3894 0.146333
R13113 GNDA.n3903 GNDA.n3902 0.146333
R13114 GNDA.n3906 GNDA.n3903 0.146333
R13115 GNDA.n3906 GNDA.n826 0.146333
R13116 GNDA.n3914 GNDA.n822 0.146333
R13117 GNDA.n3918 GNDA.n822 0.146333
R13118 GNDA.n3919 GNDA.n3918 0.146333
R13119 GNDA.n3927 GNDA.n3926 0.146333
R13120 GNDA.n3930 GNDA.n3927 0.146333
R13121 GNDA.n3930 GNDA.n816 0.146333
R13122 GNDA.n919 GNDA.n918 0.146333
R13123 GNDA.n918 GNDA.n846 0.146333
R13124 GNDA.n914 GNDA.n846 0.146333
R13125 GNDA.n908 GNDA.n854 0.146333
R13126 GNDA.n908 GNDA.n907 0.146333
R13127 GNDA.n907 GNDA.n906 0.146333
R13128 GNDA.n901 GNDA.n900 0.146333
R13129 GNDA.n900 GNDA.n870 0.146333
R13130 GNDA.n896 GNDA.n870 0.146333
R13131 GNDA.n890 GNDA.n878 0.146333
R13132 GNDA.n890 GNDA.n889 0.146333
R13133 GNDA.n889 GNDA.n888 0.146333
R13134 GNDA.n3678 GNDA.n3673 0.146333
R13135 GNDA.n3682 GNDA.n3673 0.146333
R13136 GNDA.n3683 GNDA.n3682 0.146333
R13137 GNDA.n3691 GNDA.n3690 0.146333
R13138 GNDA.n3694 GNDA.n3691 0.146333
R13139 GNDA.n3694 GNDA.n3665 0.146333
R13140 GNDA.n3702 GNDA.n3661 0.146333
R13141 GNDA.n3706 GNDA.n3661 0.146333
R13142 GNDA.n3707 GNDA.n3706 0.146333
R13143 GNDA.n3715 GNDA.n3714 0.146333
R13144 GNDA.n3718 GNDA.n3715 0.146333
R13145 GNDA.n3718 GNDA.n3655 0.146333
R13146 GNDA.n3747 GNDA.n3742 0.146333
R13147 GNDA.n3751 GNDA.n3742 0.146333
R13148 GNDA.n3752 GNDA.n3751 0.146333
R13149 GNDA.n3760 GNDA.n3759 0.146333
R13150 GNDA.n3763 GNDA.n3760 0.146333
R13151 GNDA.n3763 GNDA.n3734 0.146333
R13152 GNDA.n3771 GNDA.n3730 0.146333
R13153 GNDA.n3775 GNDA.n3730 0.146333
R13154 GNDA.n3776 GNDA.n3775 0.146333
R13155 GNDA.n3784 GNDA.n3783 0.146333
R13156 GNDA.n3787 GNDA.n3784 0.146333
R13157 GNDA.n3787 GNDA.n3724 0.146333
R13158 GNDA.n3803 GNDA.n937 0.146333
R13159 GNDA.n3808 GNDA.n3803 0.146333
R13160 GNDA.n3809 GNDA.n3808 0.146333
R13161 GNDA.n3819 GNDA.n3818 0.146333
R13162 GNDA.n3822 GNDA.n3819 0.146333
R13163 GNDA.n3822 GNDA.n3799 0.146333
R13164 GNDA.n3832 GNDA.n3797 0.146333
R13165 GNDA.n3838 GNDA.n3797 0.146333
R13166 GNDA.n3839 GNDA.n3838 0.146333
R13167 GNDA.n3849 GNDA.n3848 0.146333
R13168 GNDA.n3852 GNDA.n3849 0.146333
R13169 GNDA.n3852 GNDA.n3793 0.146333
R13170 GNDA.n3473 GNDA.n3472 0.146333
R13171 GNDA.n3472 GNDA.n3400 0.146333
R13172 GNDA.n3468 GNDA.n3400 0.146333
R13173 GNDA.n3462 GNDA.n3408 0.146333
R13174 GNDA.n3462 GNDA.n3461 0.146333
R13175 GNDA.n3461 GNDA.n3460 0.146333
R13176 GNDA.n3455 GNDA.n3454 0.146333
R13177 GNDA.n3454 GNDA.n3424 0.146333
R13178 GNDA.n3450 GNDA.n3424 0.146333
R13179 GNDA.n3444 GNDA.n3432 0.146333
R13180 GNDA.n3444 GNDA.n3443 0.146333
R13181 GNDA.n3443 GNDA.n3442 0.146333
R13182 GNDA.n3492 GNDA.n971 0.146333
R13183 GNDA.n3496 GNDA.n971 0.146333
R13184 GNDA.n3497 GNDA.n3496 0.146333
R13185 GNDA.n3505 GNDA.n3504 0.146333
R13186 GNDA.n3508 GNDA.n3505 0.146333
R13187 GNDA.n3508 GNDA.n963 0.146333
R13188 GNDA.n3516 GNDA.n959 0.146333
R13189 GNDA.n3520 GNDA.n959 0.146333
R13190 GNDA.n3521 GNDA.n3520 0.146333
R13191 GNDA.n3529 GNDA.n3528 0.146333
R13192 GNDA.n3532 GNDA.n3529 0.146333
R13193 GNDA.n3532 GNDA.n953 0.146333
R13194 GNDA.n2813 GNDA.n2808 0.146333
R13195 GNDA.n2817 GNDA.n2808 0.146333
R13196 GNDA.n2818 GNDA.n2817 0.146333
R13197 GNDA.n2826 GNDA.n2825 0.146333
R13198 GNDA.n2829 GNDA.n2826 0.146333
R13199 GNDA.n2829 GNDA.n2800 0.146333
R13200 GNDA.n2837 GNDA.n2796 0.146333
R13201 GNDA.n2841 GNDA.n2796 0.146333
R13202 GNDA.n2842 GNDA.n2841 0.146333
R13203 GNDA.n2850 GNDA.n2849 0.146333
R13204 GNDA.n2853 GNDA.n2850 0.146333
R13205 GNDA.n2853 GNDA.n2790 0.146333
R13206 GNDA.n2882 GNDA.n2877 0.146333
R13207 GNDA.n2886 GNDA.n2877 0.146333
R13208 GNDA.n2887 GNDA.n2886 0.146333
R13209 GNDA.n2895 GNDA.n2894 0.146333
R13210 GNDA.n2898 GNDA.n2895 0.146333
R13211 GNDA.n2898 GNDA.n2869 0.146333
R13212 GNDA.n2906 GNDA.n2865 0.146333
R13213 GNDA.n2910 GNDA.n2865 0.146333
R13214 GNDA.n2911 GNDA.n2910 0.146333
R13215 GNDA.n2919 GNDA.n2918 0.146333
R13216 GNDA.n2922 GNDA.n2919 0.146333
R13217 GNDA.n2922 GNDA.n2859 0.146333
R13218 GNDA.n2951 GNDA.n2946 0.146333
R13219 GNDA.n2955 GNDA.n2946 0.146333
R13220 GNDA.n2956 GNDA.n2955 0.146333
R13221 GNDA.n2964 GNDA.n2963 0.146333
R13222 GNDA.n2967 GNDA.n2964 0.146333
R13223 GNDA.n2967 GNDA.n2938 0.146333
R13224 GNDA.n2975 GNDA.n2934 0.146333
R13225 GNDA.n2979 GNDA.n2934 0.146333
R13226 GNDA.n2980 GNDA.n2979 0.146333
R13227 GNDA.n2988 GNDA.n2987 0.146333
R13228 GNDA.n2991 GNDA.n2988 0.146333
R13229 GNDA.n2991 GNDA.n2928 0.146333
R13230 GNDA.n3020 GNDA.n3015 0.146333
R13231 GNDA.n3024 GNDA.n3015 0.146333
R13232 GNDA.n3025 GNDA.n3024 0.146333
R13233 GNDA.n3033 GNDA.n3032 0.146333
R13234 GNDA.n3036 GNDA.n3033 0.146333
R13235 GNDA.n3036 GNDA.n3007 0.146333
R13236 GNDA.n3044 GNDA.n3003 0.146333
R13237 GNDA.n3048 GNDA.n3003 0.146333
R13238 GNDA.n3049 GNDA.n3048 0.146333
R13239 GNDA.n3057 GNDA.n3056 0.146333
R13240 GNDA.n3060 GNDA.n3057 0.146333
R13241 GNDA.n3060 GNDA.n2997 0.146333
R13242 GNDA.n3089 GNDA.n3084 0.146333
R13243 GNDA.n3093 GNDA.n3084 0.146333
R13244 GNDA.n3094 GNDA.n3093 0.146333
R13245 GNDA.n3102 GNDA.n3101 0.146333
R13246 GNDA.n3105 GNDA.n3102 0.146333
R13247 GNDA.n3105 GNDA.n3076 0.146333
R13248 GNDA.n3113 GNDA.n3072 0.146333
R13249 GNDA.n3117 GNDA.n3072 0.146333
R13250 GNDA.n3118 GNDA.n3117 0.146333
R13251 GNDA.n3126 GNDA.n3125 0.146333
R13252 GNDA.n3129 GNDA.n3126 0.146333
R13253 GNDA.n3129 GNDA.n3066 0.146333
R13254 GNDA.n3158 GNDA.n3153 0.146333
R13255 GNDA.n3162 GNDA.n3153 0.146333
R13256 GNDA.n3163 GNDA.n3162 0.146333
R13257 GNDA.n3171 GNDA.n3170 0.146333
R13258 GNDA.n3174 GNDA.n3171 0.146333
R13259 GNDA.n3174 GNDA.n3145 0.146333
R13260 GNDA.n3182 GNDA.n3141 0.146333
R13261 GNDA.n3186 GNDA.n3141 0.146333
R13262 GNDA.n3187 GNDA.n3186 0.146333
R13263 GNDA.n3195 GNDA.n3194 0.146333
R13264 GNDA.n3198 GNDA.n3195 0.146333
R13265 GNDA.n3198 GNDA.n3135 0.146333
R13266 GNDA.n3227 GNDA.n3222 0.146333
R13267 GNDA.n3231 GNDA.n3222 0.146333
R13268 GNDA.n3232 GNDA.n3231 0.146333
R13269 GNDA.n3240 GNDA.n3239 0.146333
R13270 GNDA.n3243 GNDA.n3240 0.146333
R13271 GNDA.n3243 GNDA.n3214 0.146333
R13272 GNDA.n3251 GNDA.n3210 0.146333
R13273 GNDA.n3255 GNDA.n3210 0.146333
R13274 GNDA.n3256 GNDA.n3255 0.146333
R13275 GNDA.n3264 GNDA.n3263 0.146333
R13276 GNDA.n3267 GNDA.n3264 0.146333
R13277 GNDA.n3267 GNDA.n3204 0.146333
R13278 GNDA.n3283 GNDA.n1039 0.146333
R13279 GNDA.n3288 GNDA.n3283 0.146333
R13280 GNDA.n3289 GNDA.n3288 0.146333
R13281 GNDA.n3299 GNDA.n3298 0.146333
R13282 GNDA.n3302 GNDA.n3299 0.146333
R13283 GNDA.n3302 GNDA.n3279 0.146333
R13284 GNDA.n3312 GNDA.n3277 0.146333
R13285 GNDA.n3318 GNDA.n3277 0.146333
R13286 GNDA.n3319 GNDA.n3318 0.146333
R13287 GNDA.n3329 GNDA.n3328 0.146333
R13288 GNDA.n3332 GNDA.n3329 0.146333
R13289 GNDA.n3332 GNDA.n3273 0.146333
R13290 GNDA.n591 GNDA.n590 0.146333
R13291 GNDA.n590 GNDA.n518 0.146333
R13292 GNDA.n586 GNDA.n518 0.146333
R13293 GNDA.n580 GNDA.n526 0.146333
R13294 GNDA.n580 GNDA.n579 0.146333
R13295 GNDA.n579 GNDA.n578 0.146333
R13296 GNDA.n573 GNDA.n572 0.146333
R13297 GNDA.n572 GNDA.n542 0.146333
R13298 GNDA.n568 GNDA.n542 0.146333
R13299 GNDA.n562 GNDA.n550 0.146333
R13300 GNDA.n562 GNDA.n561 0.146333
R13301 GNDA.n561 GNDA.n560 0.146333
R13302 GNDA.n1490 GNDA.n1487 0.146333
R13303 GNDA.n1496 GNDA.n1487 0.146333
R13304 GNDA.n1496 GNDA.n1485 0.146333
R13305 GNDA.n1506 GNDA.n1481 0.146333
R13306 GNDA.n1510 GNDA.n1481 0.146333
R13307 GNDA.n1510 GNDA.n1479 0.146333
R13308 GNDA.n1520 GNDA.n1475 0.146333
R13309 GNDA.n1526 GNDA.n1475 0.146333
R13310 GNDA.n1526 GNDA.n1473 0.146333
R13311 GNDA.n1536 GNDA.n1469 0.146333
R13312 GNDA.n1540 GNDA.n1469 0.146333
R13313 GNDA.n1540 GNDA.n1467 0.146333
R13314 GNDA.n1366 GNDA.n1365 0.146333
R13315 GNDA.n1366 GNDA.n1360 0.146333
R13316 GNDA.n1376 GNDA.n1358 0.146333
R13317 GNDA.n1384 GNDA.n1358 0.146333
R13318 GNDA.n1385 GNDA.n1384 0.146333
R13319 GNDA.n1395 GNDA.n1394 0.146333
R13320 GNDA.n1396 GNDA.n1395 0.146333
R13321 GNDA.n1396 GNDA.n1354 0.146333
R13322 GNDA.n1406 GNDA.n1352 0.146333
R13323 GNDA.n1414 GNDA.n1352 0.146333
R13324 GNDA.n1415 GNDA.n1414 0.146333
R13325 GNDA.n1363 GNDA.n1361 0.146333
R13326 GNDA.n1369 GNDA.n1361 0.146333
R13327 GNDA.n1370 GNDA.n1369 0.146333
R13328 GNDA.n1380 GNDA.n1379 0.146333
R13329 GNDA.n1383 GNDA.n1380 0.146333
R13330 GNDA.n1383 GNDA.n1357 0.146333
R13331 GNDA.n1393 GNDA.n1355 0.146333
R13332 GNDA.n1399 GNDA.n1355 0.146333
R13333 GNDA.n1400 GNDA.n1399 0.146333
R13334 GNDA.n1410 GNDA.n1409 0.146333
R13335 GNDA.n1413 GNDA.n1410 0.146333
R13336 GNDA.n1413 GNDA.n1351 0.146333
R13337 GNDA.n4725 GNDA.n4564 0.135917
R13338 GNDA.n4679 GNDA.n4676 0.135917
R13339 GNDA.n4685 GNDA.n4668 0.135917
R13340 GNDA.n4695 GNDA.n4666 0.135917
R13341 GNDA.n4699 GNDA.n4696 0.135917
R13342 GNDA.n4709 GNDA.n4706 0.135917
R13343 GNDA.n4715 GNDA.n4662 0.135917
R13344 GNDA.n4593 GNDA.n4591 0.135917
R13345 GNDA.n4603 GNDA.n4600 0.135917
R13346 GNDA.n4609 GNDA.n4587 0.135917
R13347 GNDA.n4619 GNDA.n4585 0.135917
R13348 GNDA.n4623 GNDA.n4620 0.135917
R13349 GNDA.n4633 GNDA.n4630 0.135917
R13350 GNDA.n4639 GNDA.n4581 0.135917
R13351 GNDA.n4551 GNDA.n4473 0.135917
R13352 GNDA.n4477 GNDA.n4476 0.135917
R13353 GNDA.n4479 GNDA.n4478 0.135917
R13354 GNDA.n4483 GNDA.n4482 0.135917
R13355 GNDA.n4485 GNDA.n4484 0.135917
R13356 GNDA.n4489 GNDA.n4488 0.135917
R13357 GNDA.n4491 GNDA.n4490 0.135917
R13358 GNDA.n4753 GNDA.n4751 0.135917
R13359 GNDA.n4763 GNDA.n4760 0.135917
R13360 GNDA.n4769 GNDA.n4466 0.135917
R13361 GNDA.n4779 GNDA.n4464 0.135917
R13362 GNDA.n4783 GNDA.n4780 0.135917
R13363 GNDA.n4793 GNDA.n4790 0.135917
R13364 GNDA.n4799 GNDA.n4460 0.135917
R13365 GNDA.n4273 GNDA.n484 0.135917
R13366 GNDA.n4227 GNDA.n4224 0.135917
R13367 GNDA.n4233 GNDA.n4216 0.135917
R13368 GNDA.n4243 GNDA.n4214 0.135917
R13369 GNDA.n4247 GNDA.n4244 0.135917
R13370 GNDA.n4257 GNDA.n4254 0.135917
R13371 GNDA.n4263 GNDA.n4210 0.135917
R13372 GNDA.n4874 GNDA.n444 0.135917
R13373 GNDA.n4828 GNDA.n4825 0.135917
R13374 GNDA.n4834 GNDA.n4817 0.135917
R13375 GNDA.n4844 GNDA.n4815 0.135917
R13376 GNDA.n4848 GNDA.n4845 0.135917
R13377 GNDA.n4858 GNDA.n4855 0.135917
R13378 GNDA.n4864 GNDA.n4811 0.135917
R13379 GNDA.n4378 GNDA.n4376 0.135917
R13380 GNDA.n4388 GNDA.n4385 0.135917
R13381 GNDA.n4394 GNDA.n468 0.135917
R13382 GNDA.n4404 GNDA.n466 0.135917
R13383 GNDA.n4408 GNDA.n4405 0.135917
R13384 GNDA.n4418 GNDA.n4415 0.135917
R13385 GNDA.n4424 GNDA.n462 0.135917
R13386 GNDA.n4363 GNDA.n4285 0.135917
R13387 GNDA.n4289 GNDA.n4288 0.135917
R13388 GNDA.n4291 GNDA.n4290 0.135917
R13389 GNDA.n4295 GNDA.n4294 0.135917
R13390 GNDA.n4297 GNDA.n4296 0.135917
R13391 GNDA.n4301 GNDA.n4300 0.135917
R13392 GNDA.n4303 GNDA.n4302 0.135917
R13393 GNDA.n4141 GNDA.n4139 0.135917
R13394 GNDA.n4151 GNDA.n4148 0.135917
R13395 GNDA.n4157 GNDA.n508 0.135917
R13396 GNDA.n4167 GNDA.n506 0.135917
R13397 GNDA.n4171 GNDA.n4168 0.135917
R13398 GNDA.n4181 GNDA.n4178 0.135917
R13399 GNDA.n4187 GNDA.n502 0.135917
R13400 GNDA.n3986 GNDA.n3985 0.135917
R13401 GNDA.n3980 GNDA.n3979 0.135917
R13402 GNDA.n3978 GNDA.n782 0.135917
R13403 GNDA.n3972 GNDA.n787 0.135917
R13404 GNDA.n3968 GNDA.n3967 0.135917
R13405 GNDA.n3962 GNDA.n3961 0.135917
R13406 GNDA.n3960 GNDA.n797 0.135917
R13407 GNDA.n3574 GNDA.n3572 0.135917
R13408 GNDA.n3582 GNDA.n3579 0.135917
R13409 GNDA.n3586 GNDA.n3564 0.135917
R13410 GNDA.n3594 GNDA.n3560 0.135917
R13411 GNDA.n3598 GNDA.n3595 0.135917
R13412 GNDA.n3606 GNDA.n3603 0.135917
R13413 GNDA.n3610 GNDA.n3552 0.135917
R13414 GNDA.n3890 GNDA.n3888 0.135917
R13415 GNDA.n3898 GNDA.n3895 0.135917
R13416 GNDA.n3902 GNDA.n830 0.135917
R13417 GNDA.n3910 GNDA.n826 0.135917
R13418 GNDA.n3914 GNDA.n3911 0.135917
R13419 GNDA.n3922 GNDA.n3919 0.135917
R13420 GNDA.n3926 GNDA.n818 0.135917
R13421 GNDA.n920 GNDA.n919 0.135917
R13422 GNDA.n914 GNDA.n913 0.135917
R13423 GNDA.n912 GNDA.n854 0.135917
R13424 GNDA.n906 GNDA.n862 0.135917
R13425 GNDA.n902 GNDA.n901 0.135917
R13426 GNDA.n896 GNDA.n895 0.135917
R13427 GNDA.n894 GNDA.n878 0.135917
R13428 GNDA.n3678 GNDA.n3676 0.135917
R13429 GNDA.n3686 GNDA.n3683 0.135917
R13430 GNDA.n3690 GNDA.n3669 0.135917
R13431 GNDA.n3698 GNDA.n3665 0.135917
R13432 GNDA.n3702 GNDA.n3699 0.135917
R13433 GNDA.n3710 GNDA.n3707 0.135917
R13434 GNDA.n3714 GNDA.n3657 0.135917
R13435 GNDA.n3747 GNDA.n3745 0.135917
R13436 GNDA.n3755 GNDA.n3752 0.135917
R13437 GNDA.n3759 GNDA.n3738 0.135917
R13438 GNDA.n3767 GNDA.n3734 0.135917
R13439 GNDA.n3771 GNDA.n3768 0.135917
R13440 GNDA.n3779 GNDA.n3776 0.135917
R13441 GNDA.n3783 GNDA.n3726 0.135917
R13442 GNDA.n3858 GNDA.n937 0.135917
R13443 GNDA.n3812 GNDA.n3809 0.135917
R13444 GNDA.n3818 GNDA.n3801 0.135917
R13445 GNDA.n3828 GNDA.n3799 0.135917
R13446 GNDA.n3832 GNDA.n3829 0.135917
R13447 GNDA.n3842 GNDA.n3839 0.135917
R13448 GNDA.n3848 GNDA.n3795 0.135917
R13449 GNDA.n3474 GNDA.n3473 0.135917
R13450 GNDA.n3468 GNDA.n3467 0.135917
R13451 GNDA.n3466 GNDA.n3408 0.135917
R13452 GNDA.n3460 GNDA.n3416 0.135917
R13453 GNDA.n3456 GNDA.n3455 0.135917
R13454 GNDA.n3450 GNDA.n3449 0.135917
R13455 GNDA.n3448 GNDA.n3432 0.135917
R13456 GNDA.n3492 GNDA.n3490 0.135917
R13457 GNDA.n3500 GNDA.n3497 0.135917
R13458 GNDA.n3504 GNDA.n967 0.135917
R13459 GNDA.n3512 GNDA.n963 0.135917
R13460 GNDA.n3516 GNDA.n3513 0.135917
R13461 GNDA.n3524 GNDA.n3521 0.135917
R13462 GNDA.n3528 GNDA.n955 0.135917
R13463 GNDA.n2813 GNDA.n2811 0.135917
R13464 GNDA.n2821 GNDA.n2818 0.135917
R13465 GNDA.n2825 GNDA.n2804 0.135917
R13466 GNDA.n2833 GNDA.n2800 0.135917
R13467 GNDA.n2837 GNDA.n2834 0.135917
R13468 GNDA.n2845 GNDA.n2842 0.135917
R13469 GNDA.n2849 GNDA.n2792 0.135917
R13470 GNDA.n2882 GNDA.n2880 0.135917
R13471 GNDA.n2890 GNDA.n2887 0.135917
R13472 GNDA.n2894 GNDA.n2873 0.135917
R13473 GNDA.n2902 GNDA.n2869 0.135917
R13474 GNDA.n2906 GNDA.n2903 0.135917
R13475 GNDA.n2914 GNDA.n2911 0.135917
R13476 GNDA.n2918 GNDA.n2861 0.135917
R13477 GNDA.n2951 GNDA.n2949 0.135917
R13478 GNDA.n2959 GNDA.n2956 0.135917
R13479 GNDA.n2963 GNDA.n2942 0.135917
R13480 GNDA.n2971 GNDA.n2938 0.135917
R13481 GNDA.n2975 GNDA.n2972 0.135917
R13482 GNDA.n2983 GNDA.n2980 0.135917
R13483 GNDA.n2987 GNDA.n2930 0.135917
R13484 GNDA.n3020 GNDA.n3018 0.135917
R13485 GNDA.n3028 GNDA.n3025 0.135917
R13486 GNDA.n3032 GNDA.n3011 0.135917
R13487 GNDA.n3040 GNDA.n3007 0.135917
R13488 GNDA.n3044 GNDA.n3041 0.135917
R13489 GNDA.n3052 GNDA.n3049 0.135917
R13490 GNDA.n3056 GNDA.n2999 0.135917
R13491 GNDA.n3089 GNDA.n3087 0.135917
R13492 GNDA.n3097 GNDA.n3094 0.135917
R13493 GNDA.n3101 GNDA.n3080 0.135917
R13494 GNDA.n3109 GNDA.n3076 0.135917
R13495 GNDA.n3113 GNDA.n3110 0.135917
R13496 GNDA.n3121 GNDA.n3118 0.135917
R13497 GNDA.n3125 GNDA.n3068 0.135917
R13498 GNDA.n3158 GNDA.n3156 0.135917
R13499 GNDA.n3166 GNDA.n3163 0.135917
R13500 GNDA.n3170 GNDA.n3149 0.135917
R13501 GNDA.n3178 GNDA.n3145 0.135917
R13502 GNDA.n3182 GNDA.n3179 0.135917
R13503 GNDA.n3190 GNDA.n3187 0.135917
R13504 GNDA.n3194 GNDA.n3137 0.135917
R13505 GNDA.n3227 GNDA.n3225 0.135917
R13506 GNDA.n3235 GNDA.n3232 0.135917
R13507 GNDA.n3239 GNDA.n3218 0.135917
R13508 GNDA.n3247 GNDA.n3214 0.135917
R13509 GNDA.n3251 GNDA.n3248 0.135917
R13510 GNDA.n3259 GNDA.n3256 0.135917
R13511 GNDA.n3263 GNDA.n3206 0.135917
R13512 GNDA.n3338 GNDA.n1039 0.135917
R13513 GNDA.n3292 GNDA.n3289 0.135917
R13514 GNDA.n3298 GNDA.n3281 0.135917
R13515 GNDA.n3308 GNDA.n3279 0.135917
R13516 GNDA.n3312 GNDA.n3309 0.135917
R13517 GNDA.n3322 GNDA.n3319 0.135917
R13518 GNDA.n3328 GNDA.n3275 0.135917
R13519 GNDA.n592 GNDA.n591 0.135917
R13520 GNDA.n586 GNDA.n585 0.135917
R13521 GNDA.n584 GNDA.n526 0.135917
R13522 GNDA.n578 GNDA.n534 0.135917
R13523 GNDA.n574 GNDA.n573 0.135917
R13524 GNDA.n568 GNDA.n567 0.135917
R13525 GNDA.n566 GNDA.n550 0.135917
R13526 GNDA.n1500 GNDA.n1485 0.135917
R13527 GNDA.n1506 GNDA.n1483 0.135917
R13528 GNDA.n1516 GNDA.n1479 0.135917
R13529 GNDA.n1520 GNDA.n1477 0.135917
R13530 GNDA.n1530 GNDA.n1473 0.135917
R13531 GNDA.n1536 GNDA.n1471 0.135917
R13532 GNDA.n1545 GNDA.n1467 0.135917
R13533 GNDA.n1374 GNDA.n1360 0.135917
R13534 GNDA.n1376 GNDA.n1375 0.135917
R13535 GNDA.n1386 GNDA.n1385 0.135917
R13536 GNDA.n1394 GNDA.n1356 0.135917
R13537 GNDA.n1404 GNDA.n1354 0.135917
R13538 GNDA.n1406 GNDA.n1405 0.135917
R13539 GNDA.n2576 GNDA.n1415 0.135917
R13540 GNDA.n1373 GNDA.n1370 0.135917
R13541 GNDA.n1379 GNDA.n1359 0.135917
R13542 GNDA.n1389 GNDA.n1357 0.135917
R13543 GNDA.n1393 GNDA.n1390 0.135917
R13544 GNDA.n1403 GNDA.n1400 0.135917
R13545 GNDA.n1409 GNDA.n1353 0.135917
R13546 GNDA.n2577 GNDA.n1351 0.135917
R13547 GNDA.n2579 GNDA.n1349 0.135331
R13548 GNDA.n4679 GNDA.n4668 0.1255
R13549 GNDA.n4696 GNDA.n4695 0.1255
R13550 GNDA.n4709 GNDA.n4662 0.1255
R13551 GNDA.n4603 GNDA.n4587 0.1255
R13552 GNDA.n4620 GNDA.n4619 0.1255
R13553 GNDA.n4633 GNDA.n4581 0.1255
R13554 GNDA.n4478 GNDA.n4477 0.1255
R13555 GNDA.n4484 GNDA.n4483 0.1255
R13556 GNDA.n4490 GNDA.n4489 0.1255
R13557 GNDA.n4763 GNDA.n4466 0.1255
R13558 GNDA.n4780 GNDA.n4779 0.1255
R13559 GNDA.n4793 GNDA.n4460 0.1255
R13560 GNDA.n4227 GNDA.n4216 0.1255
R13561 GNDA.n4244 GNDA.n4243 0.1255
R13562 GNDA.n4257 GNDA.n4210 0.1255
R13563 GNDA.n4828 GNDA.n4817 0.1255
R13564 GNDA.n4845 GNDA.n4844 0.1255
R13565 GNDA.n4858 GNDA.n4811 0.1255
R13566 GNDA.n4388 GNDA.n468 0.1255
R13567 GNDA.n4405 GNDA.n4404 0.1255
R13568 GNDA.n4418 GNDA.n462 0.1255
R13569 GNDA.n4290 GNDA.n4289 0.1255
R13570 GNDA.n4296 GNDA.n4295 0.1255
R13571 GNDA.n4302 GNDA.n4301 0.1255
R13572 GNDA.n4151 GNDA.n508 0.1255
R13573 GNDA.n4168 GNDA.n4167 0.1255
R13574 GNDA.n4181 GNDA.n502 0.1255
R13575 GNDA.n3979 GNDA.n3978 0.1255
R13576 GNDA.n3968 GNDA.n787 0.1255
R13577 GNDA.n3961 GNDA.n3960 0.1255
R13578 GNDA.n4055 GNDA.n4054 0.1255
R13579 GNDA.n4050 GNDA.n751 0.1255
R13580 GNDA.n3582 GNDA.n3564 0.1255
R13581 GNDA.n3595 GNDA.n3594 0.1255
R13582 GNDA.n3606 GNDA.n3552 0.1255
R13583 GNDA.n3898 GNDA.n830 0.1255
R13584 GNDA.n3911 GNDA.n3910 0.1255
R13585 GNDA.n3922 GNDA.n818 0.1255
R13586 GNDA.n913 GNDA.n912 0.1255
R13587 GNDA.n902 GNDA.n862 0.1255
R13588 GNDA.n895 GNDA.n894 0.1255
R13589 GNDA.n3686 GNDA.n3669 0.1255
R13590 GNDA.n3699 GNDA.n3698 0.1255
R13591 GNDA.n3710 GNDA.n3657 0.1255
R13592 GNDA.n3755 GNDA.n3738 0.1255
R13593 GNDA.n3768 GNDA.n3767 0.1255
R13594 GNDA.n3779 GNDA.n3726 0.1255
R13595 GNDA.n3812 GNDA.n3801 0.1255
R13596 GNDA.n3829 GNDA.n3828 0.1255
R13597 GNDA.n3842 GNDA.n3795 0.1255
R13598 GNDA.n3467 GNDA.n3466 0.1255
R13599 GNDA.n3456 GNDA.n3416 0.1255
R13600 GNDA.n3449 GNDA.n3448 0.1255
R13601 GNDA.n3500 GNDA.n967 0.1255
R13602 GNDA.n3513 GNDA.n3512 0.1255
R13603 GNDA.n3524 GNDA.n955 0.1255
R13604 GNDA.n2821 GNDA.n2804 0.1255
R13605 GNDA.n2834 GNDA.n2833 0.1255
R13606 GNDA.n2845 GNDA.n2792 0.1255
R13607 GNDA.n669 GNDA.n668 0.1255
R13608 GNDA.n733 GNDA.n645 0.1255
R13609 GNDA.n692 GNDA.n685 0.1255
R13610 GNDA.n4118 GNDA.n4117 0.1255
R13611 GNDA.n2890 GNDA.n2873 0.1255
R13612 GNDA.n2903 GNDA.n2902 0.1255
R13613 GNDA.n2914 GNDA.n2861 0.1255
R13614 GNDA.n2959 GNDA.n2942 0.1255
R13615 GNDA.n2972 GNDA.n2971 0.1255
R13616 GNDA.n2983 GNDA.n2930 0.1255
R13617 GNDA.n3028 GNDA.n3011 0.1255
R13618 GNDA.n3041 GNDA.n3040 0.1255
R13619 GNDA.n3052 GNDA.n2999 0.1255
R13620 GNDA.n3097 GNDA.n3080 0.1255
R13621 GNDA.n3110 GNDA.n3109 0.1255
R13622 GNDA.n3121 GNDA.n3068 0.1255
R13623 GNDA.n3166 GNDA.n3149 0.1255
R13624 GNDA.n3179 GNDA.n3178 0.1255
R13625 GNDA.n3190 GNDA.n3137 0.1255
R13626 GNDA.n3235 GNDA.n3218 0.1255
R13627 GNDA.n3248 GNDA.n3247 0.1255
R13628 GNDA.n3259 GNDA.n3206 0.1255
R13629 GNDA.n3367 GNDA.n3364 0.1255
R13630 GNDA.n3292 GNDA.n3281 0.1255
R13631 GNDA.n3309 GNDA.n3308 0.1255
R13632 GNDA.n3322 GNDA.n3275 0.1255
R13633 GNDA.n585 GNDA.n584 0.1255
R13634 GNDA.n574 GNDA.n534 0.1255
R13635 GNDA.n567 GNDA.n566 0.1255
R13636 GNDA.n4885 GNDA.n4880 0.1255
R13637 GNDA.n2047 GNDA.n1895 0.1255
R13638 GNDA.n1925 GNDA.n1924 0.1255
R13639 GNDA.n1500 GNDA.n1483 0.1255
R13640 GNDA.n1516 GNDA.n1477 0.1255
R13641 GNDA.n1530 GNDA.n1471 0.1255
R13642 GNDA.n359 GNDA.n358 0.1255
R13643 GNDA.n1375 GNDA.n1374 0.1255
R13644 GNDA.n1386 GNDA.n1356 0.1255
R13645 GNDA.n1405 GNDA.n1404 0.1255
R13646 GNDA.n1373 GNDA.n1359 0.1255
R13647 GNDA.n1390 GNDA.n1389 0.1255
R13648 GNDA.n1403 GNDA.n1353 0.1255
R13649 GNDA.n708 GNDA.n707 0.123287
R13650 GNDA.n720 GNDA.n679 0.12293
R13651 GNDA.n4042 GNDA.n4040 0.115083
R13652 GNDA.n4040 GNDA.n4038 0.115083
R13653 GNDA.n4038 GNDA.n4036 0.115083
R13654 GNDA.n4036 GNDA.n4034 0.115083
R13655 GNDA.n4034 GNDA.n4032 0.115083
R13656 GNDA.n4032 GNDA.n4030 0.115083
R13657 GNDA.n4030 GNDA.n4028 0.115083
R13658 GNDA.n4028 GNDA.n4026 0.115083
R13659 GNDA.n4026 GNDA.n4024 0.115083
R13660 GNDA.n4024 GNDA.n4022 0.115083
R13661 GNDA.n4022 GNDA.n4020 0.115083
R13662 GNDA.n4893 GNDA.n4891 0.115083
R13663 GNDA.n4895 GNDA.n4893 0.115083
R13664 GNDA.n4897 GNDA.n4895 0.115083
R13665 GNDA.n4899 GNDA.n4897 0.115083
R13666 GNDA.n711 GNDA.n709 0.115083
R13667 GNDA.n719 GNDA.n711 0.115083
R13668 GNDA.n1010 GNDA.n1008 0.115083
R13669 GNDA.n1008 GNDA.n1006 0.115083
R13670 GNDA.n1006 GNDA.n1004 0.115083
R13671 GNDA.n1004 GNDA.n1002 0.115083
R13672 GNDA.n2565 GNDA.n2564 0.115083
R13673 GNDA.n2564 GNDA.n2563 0.115083
R13674 GNDA.n2561 GNDA.n2560 0.115083
R13675 GNDA.n2560 GNDA.n2559 0.115083
R13676 GNDA.n2559 GNDA.n2558 0.115083
R13677 GNDA.n2558 GNDA.n2557 0.115083
R13678 GNDA.n2556 GNDA.n2555 0.115083
R13679 GNDA.n2555 GNDA.n2554 0.115083
R13680 GNDA.n2554 GNDA.n2553 0.115083
R13681 GNDA.n2551 GNDA.n2550 0.115083
R13682 GNDA.n2550 GNDA.n2549 0.115083
R13683 GNDA.n2549 GNDA.n2548 0.115083
R13684 GNDA.n3482 GNDA.n3479 0.10642
R13685 GNDA.n4134 GNDA.n4133 0.105167
R13686 GNDA.n657 GNDA.n656 0.0994583
R13687 GNDA.n4077 GNDA.n4075 0.0994583
R13688 GNDA.n3391 GNDA.n3386 0.09425
R13689 GNDA.n4282 GNDA.n4279 0.09425
R13690 GNDA.n2654 GNDA 0.0817953
R13691 GNDA.n4671 GNDA.n4563 0.0734167
R13692 GNDA.n4672 GNDA.n4671 0.0734167
R13693 GNDA.n4672 GNDA.n4669 0.0734167
R13694 GNDA.n4682 GNDA.n4667 0.0734167
R13695 GNDA.n4690 GNDA.n4667 0.0734167
R13696 GNDA.n4691 GNDA.n4690 0.0734167
R13697 GNDA.n4701 GNDA.n4700 0.0734167
R13698 GNDA.n4702 GNDA.n4701 0.0734167
R13699 GNDA.n4702 GNDA.n4663 0.0734167
R13700 GNDA.n4712 GNDA.n4661 0.0734167
R13701 GNDA.n4720 GNDA.n4661 0.0734167
R13702 GNDA.n4595 GNDA.n4594 0.0734167
R13703 GNDA.n4596 GNDA.n4595 0.0734167
R13704 GNDA.n4596 GNDA.n4588 0.0734167
R13705 GNDA.n4606 GNDA.n4586 0.0734167
R13706 GNDA.n4614 GNDA.n4586 0.0734167
R13707 GNDA.n4615 GNDA.n4614 0.0734167
R13708 GNDA.n4625 GNDA.n4624 0.0734167
R13709 GNDA.n4626 GNDA.n4625 0.0734167
R13710 GNDA.n4626 GNDA.n4582 0.0734167
R13711 GNDA.n4636 GNDA.n4580 0.0734167
R13712 GNDA.n4644 GNDA.n4580 0.0734167
R13713 GNDA.n4495 GNDA.n4472 0.0734167
R13714 GNDA.n4496 GNDA.n4495 0.0734167
R13715 GNDA.n4497 GNDA.n4496 0.0734167
R13716 GNDA.n4501 GNDA.n4500 0.0734167
R13717 GNDA.n4502 GNDA.n4501 0.0734167
R13718 GNDA.n4503 GNDA.n4502 0.0734167
R13719 GNDA.n4507 GNDA.n4506 0.0734167
R13720 GNDA.n4508 GNDA.n4507 0.0734167
R13721 GNDA.n4509 GNDA.n4508 0.0734167
R13722 GNDA.n4513 GNDA.n4512 0.0734167
R13723 GNDA.n4514 GNDA.n4513 0.0734167
R13724 GNDA.n4755 GNDA.n4754 0.0734167
R13725 GNDA.n4756 GNDA.n4755 0.0734167
R13726 GNDA.n4756 GNDA.n4467 0.0734167
R13727 GNDA.n4766 GNDA.n4465 0.0734167
R13728 GNDA.n4774 GNDA.n4465 0.0734167
R13729 GNDA.n4775 GNDA.n4774 0.0734167
R13730 GNDA.n4785 GNDA.n4784 0.0734167
R13731 GNDA.n4786 GNDA.n4785 0.0734167
R13732 GNDA.n4786 GNDA.n4461 0.0734167
R13733 GNDA.n4796 GNDA.n4459 0.0734167
R13734 GNDA.n4804 GNDA.n4459 0.0734167
R13735 GNDA.n4219 GNDA.n483 0.0734167
R13736 GNDA.n4220 GNDA.n4219 0.0734167
R13737 GNDA.n4220 GNDA.n4217 0.0734167
R13738 GNDA.n4230 GNDA.n4215 0.0734167
R13739 GNDA.n4238 GNDA.n4215 0.0734167
R13740 GNDA.n4239 GNDA.n4238 0.0734167
R13741 GNDA.n4249 GNDA.n4248 0.0734167
R13742 GNDA.n4250 GNDA.n4249 0.0734167
R13743 GNDA.n4250 GNDA.n4211 0.0734167
R13744 GNDA.n4260 GNDA.n4209 0.0734167
R13745 GNDA.n4268 GNDA.n4209 0.0734167
R13746 GNDA.n4820 GNDA.n443 0.0734167
R13747 GNDA.n4821 GNDA.n4820 0.0734167
R13748 GNDA.n4821 GNDA.n4818 0.0734167
R13749 GNDA.n4831 GNDA.n4816 0.0734167
R13750 GNDA.n4839 GNDA.n4816 0.0734167
R13751 GNDA.n4840 GNDA.n4839 0.0734167
R13752 GNDA.n4850 GNDA.n4849 0.0734167
R13753 GNDA.n4851 GNDA.n4850 0.0734167
R13754 GNDA.n4851 GNDA.n4812 0.0734167
R13755 GNDA.n4861 GNDA.n4810 0.0734167
R13756 GNDA.n4869 GNDA.n4810 0.0734167
R13757 GNDA.n4380 GNDA.n4379 0.0734167
R13758 GNDA.n4381 GNDA.n4380 0.0734167
R13759 GNDA.n4381 GNDA.n469 0.0734167
R13760 GNDA.n4391 GNDA.n467 0.0734167
R13761 GNDA.n4399 GNDA.n467 0.0734167
R13762 GNDA.n4400 GNDA.n4399 0.0734167
R13763 GNDA.n4410 GNDA.n4409 0.0734167
R13764 GNDA.n4411 GNDA.n4410 0.0734167
R13765 GNDA.n4411 GNDA.n463 0.0734167
R13766 GNDA.n4421 GNDA.n461 0.0734167
R13767 GNDA.n4429 GNDA.n461 0.0734167
R13768 GNDA.n4307 GNDA.n4284 0.0734167
R13769 GNDA.n4308 GNDA.n4307 0.0734167
R13770 GNDA.n4309 GNDA.n4308 0.0734167
R13771 GNDA.n4313 GNDA.n4312 0.0734167
R13772 GNDA.n4314 GNDA.n4313 0.0734167
R13773 GNDA.n4315 GNDA.n4314 0.0734167
R13774 GNDA.n4319 GNDA.n4318 0.0734167
R13775 GNDA.n4320 GNDA.n4319 0.0734167
R13776 GNDA.n4321 GNDA.n4320 0.0734167
R13777 GNDA.n4325 GNDA.n4324 0.0734167
R13778 GNDA.n4326 GNDA.n4325 0.0734167
R13779 GNDA.n4143 GNDA.n4142 0.0734167
R13780 GNDA.n4144 GNDA.n4143 0.0734167
R13781 GNDA.n4144 GNDA.n509 0.0734167
R13782 GNDA.n4154 GNDA.n507 0.0734167
R13783 GNDA.n4162 GNDA.n507 0.0734167
R13784 GNDA.n4163 GNDA.n4162 0.0734167
R13785 GNDA.n4173 GNDA.n4172 0.0734167
R13786 GNDA.n4174 GNDA.n4173 0.0734167
R13787 GNDA.n4174 GNDA.n503 0.0734167
R13788 GNDA.n4184 GNDA.n501 0.0734167
R13789 GNDA.n4192 GNDA.n501 0.0734167
R13790 GNDA.n3983 GNDA.n773 0.0734167
R13791 GNDA.n3983 GNDA.n3982 0.0734167
R13792 GNDA.n3982 GNDA.n3981 0.0734167
R13793 GNDA.n3976 GNDA.n3975 0.0734167
R13794 GNDA.n3975 GNDA.n783 0.0734167
R13795 GNDA.n3971 GNDA.n783 0.0734167
R13796 GNDA.n3965 GNDA.n788 0.0734167
R13797 GNDA.n3965 GNDA.n3964 0.0734167
R13798 GNDA.n3964 GNDA.n3963 0.0734167
R13799 GNDA.n3958 GNDA.n3957 0.0734167
R13800 GNDA.n3957 GNDA.n798 0.0734167
R13801 GNDA.n3576 GNDA.n3575 0.0734167
R13802 GNDA.n3577 GNDA.n3576 0.0734167
R13803 GNDA.n3577 GNDA.n3567 0.0734167
R13804 GNDA.n3585 GNDA.n3563 0.0734167
R13805 GNDA.n3591 GNDA.n3563 0.0734167
R13806 GNDA.n3592 GNDA.n3591 0.0734167
R13807 GNDA.n3600 GNDA.n3599 0.0734167
R13808 GNDA.n3601 GNDA.n3600 0.0734167
R13809 GNDA.n3601 GNDA.n3555 0.0734167
R13810 GNDA.n3609 GNDA.n3551 0.0734167
R13811 GNDA.n3615 GNDA.n3551 0.0734167
R13812 GNDA.n3892 GNDA.n3891 0.0734167
R13813 GNDA.n3893 GNDA.n3892 0.0734167
R13814 GNDA.n3893 GNDA.n833 0.0734167
R13815 GNDA.n3901 GNDA.n829 0.0734167
R13816 GNDA.n3907 GNDA.n829 0.0734167
R13817 GNDA.n3908 GNDA.n3907 0.0734167
R13818 GNDA.n3916 GNDA.n3915 0.0734167
R13819 GNDA.n3917 GNDA.n3916 0.0734167
R13820 GNDA.n3917 GNDA.n821 0.0734167
R13821 GNDA.n3925 GNDA.n817 0.0734167
R13822 GNDA.n3931 GNDA.n817 0.0734167
R13823 GNDA.n917 GNDA.n841 0.0734167
R13824 GNDA.n917 GNDA.n916 0.0734167
R13825 GNDA.n916 GNDA.n915 0.0734167
R13826 GNDA.n910 GNDA.n909 0.0734167
R13827 GNDA.n909 GNDA.n855 0.0734167
R13828 GNDA.n905 GNDA.n855 0.0734167
R13829 GNDA.n899 GNDA.n863 0.0734167
R13830 GNDA.n899 GNDA.n898 0.0734167
R13831 GNDA.n898 GNDA.n897 0.0734167
R13832 GNDA.n892 GNDA.n891 0.0734167
R13833 GNDA.n891 GNDA.n879 0.0734167
R13834 GNDA.n3680 GNDA.n3679 0.0734167
R13835 GNDA.n3681 GNDA.n3680 0.0734167
R13836 GNDA.n3681 GNDA.n3672 0.0734167
R13837 GNDA.n3689 GNDA.n3668 0.0734167
R13838 GNDA.n3695 GNDA.n3668 0.0734167
R13839 GNDA.n3696 GNDA.n3695 0.0734167
R13840 GNDA.n3704 GNDA.n3703 0.0734167
R13841 GNDA.n3705 GNDA.n3704 0.0734167
R13842 GNDA.n3705 GNDA.n3660 0.0734167
R13843 GNDA.n3713 GNDA.n3656 0.0734167
R13844 GNDA.n3719 GNDA.n3656 0.0734167
R13845 GNDA.n3749 GNDA.n3748 0.0734167
R13846 GNDA.n3750 GNDA.n3749 0.0734167
R13847 GNDA.n3750 GNDA.n3741 0.0734167
R13848 GNDA.n3758 GNDA.n3737 0.0734167
R13849 GNDA.n3764 GNDA.n3737 0.0734167
R13850 GNDA.n3765 GNDA.n3764 0.0734167
R13851 GNDA.n3773 GNDA.n3772 0.0734167
R13852 GNDA.n3774 GNDA.n3773 0.0734167
R13853 GNDA.n3774 GNDA.n3729 0.0734167
R13854 GNDA.n3782 GNDA.n3725 0.0734167
R13855 GNDA.n3788 GNDA.n3725 0.0734167
R13856 GNDA.n3804 GNDA.n936 0.0734167
R13857 GNDA.n3805 GNDA.n3804 0.0734167
R13858 GNDA.n3805 GNDA.n3802 0.0734167
R13859 GNDA.n3815 GNDA.n3800 0.0734167
R13860 GNDA.n3823 GNDA.n3800 0.0734167
R13861 GNDA.n3824 GNDA.n3823 0.0734167
R13862 GNDA.n3834 GNDA.n3833 0.0734167
R13863 GNDA.n3835 GNDA.n3834 0.0734167
R13864 GNDA.n3835 GNDA.n3796 0.0734167
R13865 GNDA.n3845 GNDA.n3794 0.0734167
R13866 GNDA.n3853 GNDA.n3794 0.0734167
R13867 GNDA.n3471 GNDA.n3395 0.0734167
R13868 GNDA.n3471 GNDA.n3470 0.0734167
R13869 GNDA.n3470 GNDA.n3469 0.0734167
R13870 GNDA.n3464 GNDA.n3463 0.0734167
R13871 GNDA.n3463 GNDA.n3409 0.0734167
R13872 GNDA.n3459 GNDA.n3409 0.0734167
R13873 GNDA.n3453 GNDA.n3417 0.0734167
R13874 GNDA.n3453 GNDA.n3452 0.0734167
R13875 GNDA.n3452 GNDA.n3451 0.0734167
R13876 GNDA.n3446 GNDA.n3445 0.0734167
R13877 GNDA.n3445 GNDA.n3433 0.0734167
R13878 GNDA.n3494 GNDA.n3493 0.0734167
R13879 GNDA.n3495 GNDA.n3494 0.0734167
R13880 GNDA.n3495 GNDA.n970 0.0734167
R13881 GNDA.n3503 GNDA.n966 0.0734167
R13882 GNDA.n3509 GNDA.n966 0.0734167
R13883 GNDA.n3510 GNDA.n3509 0.0734167
R13884 GNDA.n3518 GNDA.n3517 0.0734167
R13885 GNDA.n3519 GNDA.n3518 0.0734167
R13886 GNDA.n3519 GNDA.n958 0.0734167
R13887 GNDA.n3527 GNDA.n954 0.0734167
R13888 GNDA.n3533 GNDA.n954 0.0734167
R13889 GNDA.n2815 GNDA.n2814 0.0734167
R13890 GNDA.n2816 GNDA.n2815 0.0734167
R13891 GNDA.n2816 GNDA.n2807 0.0734167
R13892 GNDA.n2824 GNDA.n2803 0.0734167
R13893 GNDA.n2830 GNDA.n2803 0.0734167
R13894 GNDA.n2831 GNDA.n2830 0.0734167
R13895 GNDA.n2839 GNDA.n2838 0.0734167
R13896 GNDA.n2840 GNDA.n2839 0.0734167
R13897 GNDA.n2840 GNDA.n2795 0.0734167
R13898 GNDA.n2848 GNDA.n2791 0.0734167
R13899 GNDA.n2854 GNDA.n2791 0.0734167
R13900 GNDA.n2884 GNDA.n2883 0.0734167
R13901 GNDA.n2885 GNDA.n2884 0.0734167
R13902 GNDA.n2885 GNDA.n2876 0.0734167
R13903 GNDA.n2893 GNDA.n2872 0.0734167
R13904 GNDA.n2899 GNDA.n2872 0.0734167
R13905 GNDA.n2900 GNDA.n2899 0.0734167
R13906 GNDA.n2908 GNDA.n2907 0.0734167
R13907 GNDA.n2909 GNDA.n2908 0.0734167
R13908 GNDA.n2909 GNDA.n2864 0.0734167
R13909 GNDA.n2917 GNDA.n2860 0.0734167
R13910 GNDA.n2923 GNDA.n2860 0.0734167
R13911 GNDA.n2953 GNDA.n2952 0.0734167
R13912 GNDA.n2954 GNDA.n2953 0.0734167
R13913 GNDA.n2954 GNDA.n2945 0.0734167
R13914 GNDA.n2962 GNDA.n2941 0.0734167
R13915 GNDA.n2968 GNDA.n2941 0.0734167
R13916 GNDA.n2969 GNDA.n2968 0.0734167
R13917 GNDA.n2977 GNDA.n2976 0.0734167
R13918 GNDA.n2978 GNDA.n2977 0.0734167
R13919 GNDA.n2978 GNDA.n2933 0.0734167
R13920 GNDA.n2986 GNDA.n2929 0.0734167
R13921 GNDA.n2992 GNDA.n2929 0.0734167
R13922 GNDA.n3022 GNDA.n3021 0.0734167
R13923 GNDA.n3023 GNDA.n3022 0.0734167
R13924 GNDA.n3023 GNDA.n3014 0.0734167
R13925 GNDA.n3031 GNDA.n3010 0.0734167
R13926 GNDA.n3037 GNDA.n3010 0.0734167
R13927 GNDA.n3038 GNDA.n3037 0.0734167
R13928 GNDA.n3046 GNDA.n3045 0.0734167
R13929 GNDA.n3047 GNDA.n3046 0.0734167
R13930 GNDA.n3047 GNDA.n3002 0.0734167
R13931 GNDA.n3055 GNDA.n2998 0.0734167
R13932 GNDA.n3061 GNDA.n2998 0.0734167
R13933 GNDA.n3091 GNDA.n3090 0.0734167
R13934 GNDA.n3092 GNDA.n3091 0.0734167
R13935 GNDA.n3092 GNDA.n3083 0.0734167
R13936 GNDA.n3100 GNDA.n3079 0.0734167
R13937 GNDA.n3106 GNDA.n3079 0.0734167
R13938 GNDA.n3107 GNDA.n3106 0.0734167
R13939 GNDA.n3115 GNDA.n3114 0.0734167
R13940 GNDA.n3116 GNDA.n3115 0.0734167
R13941 GNDA.n3116 GNDA.n3071 0.0734167
R13942 GNDA.n3124 GNDA.n3067 0.0734167
R13943 GNDA.n3130 GNDA.n3067 0.0734167
R13944 GNDA.n3160 GNDA.n3159 0.0734167
R13945 GNDA.n3161 GNDA.n3160 0.0734167
R13946 GNDA.n3161 GNDA.n3152 0.0734167
R13947 GNDA.n3169 GNDA.n3148 0.0734167
R13948 GNDA.n3175 GNDA.n3148 0.0734167
R13949 GNDA.n3176 GNDA.n3175 0.0734167
R13950 GNDA.n3184 GNDA.n3183 0.0734167
R13951 GNDA.n3185 GNDA.n3184 0.0734167
R13952 GNDA.n3185 GNDA.n3140 0.0734167
R13953 GNDA.n3193 GNDA.n3136 0.0734167
R13954 GNDA.n3199 GNDA.n3136 0.0734167
R13955 GNDA.n3229 GNDA.n3228 0.0734167
R13956 GNDA.n3230 GNDA.n3229 0.0734167
R13957 GNDA.n3230 GNDA.n3221 0.0734167
R13958 GNDA.n3238 GNDA.n3217 0.0734167
R13959 GNDA.n3244 GNDA.n3217 0.0734167
R13960 GNDA.n3245 GNDA.n3244 0.0734167
R13961 GNDA.n3253 GNDA.n3252 0.0734167
R13962 GNDA.n3254 GNDA.n3253 0.0734167
R13963 GNDA.n3254 GNDA.n3209 0.0734167
R13964 GNDA.n3262 GNDA.n3205 0.0734167
R13965 GNDA.n3268 GNDA.n3205 0.0734167
R13966 GNDA.n3362 GNDA.n3359 0.0734167
R13967 GNDA.n3284 GNDA.n1038 0.0734167
R13968 GNDA.n3285 GNDA.n3284 0.0734167
R13969 GNDA.n3285 GNDA.n3282 0.0734167
R13970 GNDA.n3295 GNDA.n3280 0.0734167
R13971 GNDA.n3303 GNDA.n3280 0.0734167
R13972 GNDA.n3304 GNDA.n3303 0.0734167
R13973 GNDA.n3314 GNDA.n3313 0.0734167
R13974 GNDA.n3315 GNDA.n3314 0.0734167
R13975 GNDA.n3315 GNDA.n3276 0.0734167
R13976 GNDA.n3325 GNDA.n3274 0.0734167
R13977 GNDA.n3333 GNDA.n3274 0.0734167
R13978 GNDA.n589 GNDA.n514 0.0734167
R13979 GNDA.n589 GNDA.n588 0.0734167
R13980 GNDA.n588 GNDA.n587 0.0734167
R13981 GNDA.n582 GNDA.n581 0.0734167
R13982 GNDA.n581 GNDA.n527 0.0734167
R13983 GNDA.n577 GNDA.n527 0.0734167
R13984 GNDA.n571 GNDA.n535 0.0734167
R13985 GNDA.n571 GNDA.n570 0.0734167
R13986 GNDA.n570 GNDA.n569 0.0734167
R13987 GNDA.n564 GNDA.n563 0.0734167
R13988 GNDA.n563 GNDA.n551 0.0734167
R13989 GNDA.n4746 GNDA.n437 0.0734167
R13990 GNDA.n1497 GNDA.n1486 0.0734167
R13991 GNDA.n1498 GNDA.n1497 0.0734167
R13992 GNDA.n1508 GNDA.n1507 0.0734167
R13993 GNDA.n1509 GNDA.n1508 0.0734167
R13994 GNDA.n1509 GNDA.n1478 0.0734167
R13995 GNDA.n1519 GNDA.n1474 0.0734167
R13996 GNDA.n1527 GNDA.n1474 0.0734167
R13997 GNDA.n1528 GNDA.n1527 0.0734167
R13998 GNDA.n1538 GNDA.n1537 0.0734167
R13999 GNDA.n1539 GNDA.n1538 0.0734167
R14000 GNDA.n1539 GNDA.n1466 0.0734167
R14001 GNDA.n4726 GNDA.n4563 0.0682083
R14002 GNDA.n4680 GNDA.n4669 0.0682083
R14003 GNDA.n4682 GNDA.n4681 0.0682083
R14004 GNDA.n4692 GNDA.n4691 0.0682083
R14005 GNDA.n4700 GNDA.n4665 0.0682083
R14006 GNDA.n4710 GNDA.n4663 0.0682083
R14007 GNDA.n4712 GNDA.n4711 0.0682083
R14008 GNDA.n4594 GNDA.n4590 0.0682083
R14009 GNDA.n4604 GNDA.n4588 0.0682083
R14010 GNDA.n4606 GNDA.n4605 0.0682083
R14011 GNDA.n4616 GNDA.n4615 0.0682083
R14012 GNDA.n4624 GNDA.n4584 0.0682083
R14013 GNDA.n4634 GNDA.n4582 0.0682083
R14014 GNDA.n4636 GNDA.n4635 0.0682083
R14015 GNDA.n4552 GNDA.n4472 0.0682083
R14016 GNDA.n4498 GNDA.n4497 0.0682083
R14017 GNDA.n4500 GNDA.n4499 0.0682083
R14018 GNDA.n4504 GNDA.n4503 0.0682083
R14019 GNDA.n4506 GNDA.n4505 0.0682083
R14020 GNDA.n4510 GNDA.n4509 0.0682083
R14021 GNDA.n4512 GNDA.n4511 0.0682083
R14022 GNDA.n4754 GNDA.n4750 0.0682083
R14023 GNDA.n4764 GNDA.n4467 0.0682083
R14024 GNDA.n4766 GNDA.n4765 0.0682083
R14025 GNDA.n4776 GNDA.n4775 0.0682083
R14026 GNDA.n4784 GNDA.n4463 0.0682083
R14027 GNDA.n4794 GNDA.n4461 0.0682083
R14028 GNDA.n4796 GNDA.n4795 0.0682083
R14029 GNDA.n4274 GNDA.n483 0.0682083
R14030 GNDA.n4228 GNDA.n4217 0.0682083
R14031 GNDA.n4230 GNDA.n4229 0.0682083
R14032 GNDA.n4240 GNDA.n4239 0.0682083
R14033 GNDA.n4248 GNDA.n4213 0.0682083
R14034 GNDA.n4258 GNDA.n4211 0.0682083
R14035 GNDA.n4260 GNDA.n4259 0.0682083
R14036 GNDA.n4875 GNDA.n443 0.0682083
R14037 GNDA.n4829 GNDA.n4818 0.0682083
R14038 GNDA.n4831 GNDA.n4830 0.0682083
R14039 GNDA.n4841 GNDA.n4840 0.0682083
R14040 GNDA.n4849 GNDA.n4814 0.0682083
R14041 GNDA.n4859 GNDA.n4812 0.0682083
R14042 GNDA.n4861 GNDA.n4860 0.0682083
R14043 GNDA.n4379 GNDA.n4375 0.0682083
R14044 GNDA.n4389 GNDA.n469 0.0682083
R14045 GNDA.n4391 GNDA.n4390 0.0682083
R14046 GNDA.n4401 GNDA.n4400 0.0682083
R14047 GNDA.n4409 GNDA.n465 0.0682083
R14048 GNDA.n4419 GNDA.n463 0.0682083
R14049 GNDA.n4421 GNDA.n4420 0.0682083
R14050 GNDA.n4364 GNDA.n4284 0.0682083
R14051 GNDA.n4310 GNDA.n4309 0.0682083
R14052 GNDA.n4312 GNDA.n4311 0.0682083
R14053 GNDA.n4316 GNDA.n4315 0.0682083
R14054 GNDA.n4318 GNDA.n4317 0.0682083
R14055 GNDA.n4322 GNDA.n4321 0.0682083
R14056 GNDA.n4324 GNDA.n4323 0.0682083
R14057 GNDA.n4142 GNDA.n4138 0.0682083
R14058 GNDA.n4152 GNDA.n509 0.0682083
R14059 GNDA.n4154 GNDA.n4153 0.0682083
R14060 GNDA.n4164 GNDA.n4163 0.0682083
R14061 GNDA.n4172 GNDA.n505 0.0682083
R14062 GNDA.n4182 GNDA.n503 0.0682083
R14063 GNDA.n4184 GNDA.n4183 0.0682083
R14064 GNDA.n3987 GNDA.n773 0.0682083
R14065 GNDA.n3981 GNDA.n778 0.0682083
R14066 GNDA.n3977 GNDA.n3976 0.0682083
R14067 GNDA.n3971 GNDA.n3970 0.0682083
R14068 GNDA.n3969 GNDA.n788 0.0682083
R14069 GNDA.n3963 GNDA.n793 0.0682083
R14070 GNDA.n3959 GNDA.n3958 0.0682083
R14071 GNDA.n3575 GNDA.n3571 0.0682083
R14072 GNDA.n3583 GNDA.n3567 0.0682083
R14073 GNDA.n3585 GNDA.n3584 0.0682083
R14074 GNDA.n3593 GNDA.n3592 0.0682083
R14075 GNDA.n3599 GNDA.n3559 0.0682083
R14076 GNDA.n3607 GNDA.n3555 0.0682083
R14077 GNDA.n3609 GNDA.n3608 0.0682083
R14078 GNDA.n3891 GNDA.n3887 0.0682083
R14079 GNDA.n3899 GNDA.n833 0.0682083
R14080 GNDA.n3901 GNDA.n3900 0.0682083
R14081 GNDA.n3909 GNDA.n3908 0.0682083
R14082 GNDA.n3915 GNDA.n825 0.0682083
R14083 GNDA.n3923 GNDA.n821 0.0682083
R14084 GNDA.n3925 GNDA.n3924 0.0682083
R14085 GNDA.n921 GNDA.n841 0.0682083
R14086 GNDA.n915 GNDA.n847 0.0682083
R14087 GNDA.n911 GNDA.n910 0.0682083
R14088 GNDA.n905 GNDA.n904 0.0682083
R14089 GNDA.n903 GNDA.n863 0.0682083
R14090 GNDA.n897 GNDA.n871 0.0682083
R14091 GNDA.n893 GNDA.n892 0.0682083
R14092 GNDA.n3679 GNDA.n925 0.0682083
R14093 GNDA.n3687 GNDA.n3672 0.0682083
R14094 GNDA.n3689 GNDA.n3688 0.0682083
R14095 GNDA.n3697 GNDA.n3696 0.0682083
R14096 GNDA.n3703 GNDA.n3664 0.0682083
R14097 GNDA.n3711 GNDA.n3660 0.0682083
R14098 GNDA.n3713 GNDA.n3712 0.0682083
R14099 GNDA.n3748 GNDA.n929 0.0682083
R14100 GNDA.n3756 GNDA.n3741 0.0682083
R14101 GNDA.n3758 GNDA.n3757 0.0682083
R14102 GNDA.n3766 GNDA.n3765 0.0682083
R14103 GNDA.n3772 GNDA.n3733 0.0682083
R14104 GNDA.n3780 GNDA.n3729 0.0682083
R14105 GNDA.n3782 GNDA.n3781 0.0682083
R14106 GNDA.n3859 GNDA.n936 0.0682083
R14107 GNDA.n3813 GNDA.n3802 0.0682083
R14108 GNDA.n3815 GNDA.n3814 0.0682083
R14109 GNDA.n3825 GNDA.n3824 0.0682083
R14110 GNDA.n3833 GNDA.n3798 0.0682083
R14111 GNDA.n3843 GNDA.n3796 0.0682083
R14112 GNDA.n3845 GNDA.n3844 0.0682083
R14113 GNDA.n3475 GNDA.n3395 0.0682083
R14114 GNDA.n3469 GNDA.n3401 0.0682083
R14115 GNDA.n3465 GNDA.n3464 0.0682083
R14116 GNDA.n3459 GNDA.n3458 0.0682083
R14117 GNDA.n3457 GNDA.n3417 0.0682083
R14118 GNDA.n3451 GNDA.n3425 0.0682083
R14119 GNDA.n3447 GNDA.n3446 0.0682083
R14120 GNDA.n3493 GNDA.n3489 0.0682083
R14121 GNDA.n3501 GNDA.n970 0.0682083
R14122 GNDA.n3503 GNDA.n3502 0.0682083
R14123 GNDA.n3511 GNDA.n3510 0.0682083
R14124 GNDA.n3517 GNDA.n962 0.0682083
R14125 GNDA.n3525 GNDA.n958 0.0682083
R14126 GNDA.n3527 GNDA.n3526 0.0682083
R14127 GNDA.n2814 GNDA.n979 0.0682083
R14128 GNDA.n2822 GNDA.n2807 0.0682083
R14129 GNDA.n2824 GNDA.n2823 0.0682083
R14130 GNDA.n2832 GNDA.n2831 0.0682083
R14131 GNDA.n2838 GNDA.n2799 0.0682083
R14132 GNDA.n2846 GNDA.n2795 0.0682083
R14133 GNDA.n2848 GNDA.n2847 0.0682083
R14134 GNDA.n2883 GNDA.n983 0.0682083
R14135 GNDA.n2891 GNDA.n2876 0.0682083
R14136 GNDA.n2893 GNDA.n2892 0.0682083
R14137 GNDA.n2901 GNDA.n2900 0.0682083
R14138 GNDA.n2907 GNDA.n2868 0.0682083
R14139 GNDA.n2915 GNDA.n2864 0.0682083
R14140 GNDA.n2917 GNDA.n2916 0.0682083
R14141 GNDA.n2952 GNDA.n987 0.0682083
R14142 GNDA.n2960 GNDA.n2945 0.0682083
R14143 GNDA.n2962 GNDA.n2961 0.0682083
R14144 GNDA.n2970 GNDA.n2969 0.0682083
R14145 GNDA.n2976 GNDA.n2937 0.0682083
R14146 GNDA.n2984 GNDA.n2933 0.0682083
R14147 GNDA.n2986 GNDA.n2985 0.0682083
R14148 GNDA.n3021 GNDA.n991 0.0682083
R14149 GNDA.n3029 GNDA.n3014 0.0682083
R14150 GNDA.n3031 GNDA.n3030 0.0682083
R14151 GNDA.n3039 GNDA.n3038 0.0682083
R14152 GNDA.n3045 GNDA.n3006 0.0682083
R14153 GNDA.n3053 GNDA.n3002 0.0682083
R14154 GNDA.n3055 GNDA.n3054 0.0682083
R14155 GNDA.n3090 GNDA.n1026 0.0682083
R14156 GNDA.n3098 GNDA.n3083 0.0682083
R14157 GNDA.n3100 GNDA.n3099 0.0682083
R14158 GNDA.n3108 GNDA.n3107 0.0682083
R14159 GNDA.n3114 GNDA.n3075 0.0682083
R14160 GNDA.n3122 GNDA.n3071 0.0682083
R14161 GNDA.n3124 GNDA.n3123 0.0682083
R14162 GNDA.n3159 GNDA.n1030 0.0682083
R14163 GNDA.n3167 GNDA.n3152 0.0682083
R14164 GNDA.n3169 GNDA.n3168 0.0682083
R14165 GNDA.n3177 GNDA.n3176 0.0682083
R14166 GNDA.n3183 GNDA.n3144 0.0682083
R14167 GNDA.n3191 GNDA.n3140 0.0682083
R14168 GNDA.n3193 GNDA.n3192 0.0682083
R14169 GNDA.n3228 GNDA.n1034 0.0682083
R14170 GNDA.n3236 GNDA.n3221 0.0682083
R14171 GNDA.n3238 GNDA.n3237 0.0682083
R14172 GNDA.n3246 GNDA.n3245 0.0682083
R14173 GNDA.n3252 GNDA.n3213 0.0682083
R14174 GNDA.n3260 GNDA.n3209 0.0682083
R14175 GNDA.n3262 GNDA.n3261 0.0682083
R14176 GNDA.n3339 GNDA.n1038 0.0682083
R14177 GNDA.n3293 GNDA.n3282 0.0682083
R14178 GNDA.n3295 GNDA.n3294 0.0682083
R14179 GNDA.n3305 GNDA.n3304 0.0682083
R14180 GNDA.n3313 GNDA.n3278 0.0682083
R14181 GNDA.n3323 GNDA.n3276 0.0682083
R14182 GNDA.n3325 GNDA.n3324 0.0682083
R14183 GNDA.n593 GNDA.n514 0.0682083
R14184 GNDA.n587 GNDA.n519 0.0682083
R14185 GNDA.n583 GNDA.n582 0.0682083
R14186 GNDA.n577 GNDA.n576 0.0682083
R14187 GNDA.n575 GNDA.n535 0.0682083
R14188 GNDA.n569 GNDA.n543 0.0682083
R14189 GNDA.n565 GNDA.n564 0.0682083
R14190 GNDA.n1499 GNDA.n1498 0.0682083
R14191 GNDA.n1507 GNDA.n1482 0.0682083
R14192 GNDA.n1517 GNDA.n1478 0.0682083
R14193 GNDA.n1519 GNDA.n1518 0.0682083
R14194 GNDA.n1529 GNDA.n1528 0.0682083
R14195 GNDA.n1537 GNDA.n1470 0.0682083
R14196 GNDA.n1546 GNDA.n1466 0.0682083
R14197 GNDA.n1490 GNDA.n1489 0.0672139
R14198 GNDA.n4721 GNDA.n4660 0.0672139
R14199 GNDA.n4645 GNDA.n4579 0.0672139
R14200 GNDA.n4515 GNDA.n4494 0.0672139
R14201 GNDA.n4805 GNDA.n4458 0.0672139
R14202 GNDA.n4269 GNDA.n4208 0.0672139
R14203 GNDA.n4870 GNDA.n4809 0.0672139
R14204 GNDA.n4430 GNDA.n460 0.0672139
R14205 GNDA.n4327 GNDA.n4306 0.0672139
R14206 GNDA.n4193 GNDA.n500 0.0672139
R14207 GNDA.n3954 GNDA.n3953 0.0672139
R14208 GNDA.n3616 GNDA.n3550 0.0672139
R14209 GNDA.n3932 GNDA.n816 0.0672139
R14210 GNDA.n888 GNDA.n887 0.0672139
R14211 GNDA.n3720 GNDA.n3655 0.0672139
R14212 GNDA.n3789 GNDA.n3724 0.0672139
R14213 GNDA.n3854 GNDA.n3793 0.0672139
R14214 GNDA.n3442 GNDA.n3441 0.0672139
R14215 GNDA.n3534 GNDA.n953 0.0672139
R14216 GNDA.n2855 GNDA.n2790 0.0672139
R14217 GNDA.n2924 GNDA.n2859 0.0672139
R14218 GNDA.n2993 GNDA.n2928 0.0672139
R14219 GNDA.n3062 GNDA.n2997 0.0672139
R14220 GNDA.n3131 GNDA.n3066 0.0672139
R14221 GNDA.n3200 GNDA.n3135 0.0672139
R14222 GNDA.n3269 GNDA.n3204 0.0672139
R14223 GNDA.n3334 GNDA.n3273 0.0672139
R14224 GNDA.n560 GNDA.n559 0.0672139
R14225 GNDA.n1364 GNDA.n1363 0.0667303
R14226 GNDA.n3479 GNDA.n3394 0.0636702
R14227 GNDA.n4681 GNDA.n4680 0.063
R14228 GNDA.n4692 GNDA.n4665 0.063
R14229 GNDA.n4711 GNDA.n4710 0.063
R14230 GNDA.n4605 GNDA.n4604 0.063
R14231 GNDA.n4616 GNDA.n4584 0.063
R14232 GNDA.n4635 GNDA.n4634 0.063
R14233 GNDA.n4499 GNDA.n4498 0.063
R14234 GNDA.n4505 GNDA.n4504 0.063
R14235 GNDA.n4511 GNDA.n4510 0.063
R14236 GNDA.n4765 GNDA.n4764 0.063
R14237 GNDA.n4776 GNDA.n4463 0.063
R14238 GNDA.n4795 GNDA.n4794 0.063
R14239 GNDA.n4229 GNDA.n4228 0.063
R14240 GNDA.n4240 GNDA.n4213 0.063
R14241 GNDA.n4259 GNDA.n4258 0.063
R14242 GNDA.n4830 GNDA.n4829 0.063
R14243 GNDA.n4841 GNDA.n4814 0.063
R14244 GNDA.n4860 GNDA.n4859 0.063
R14245 GNDA.n4390 GNDA.n4389 0.063
R14246 GNDA.n4401 GNDA.n465 0.063
R14247 GNDA.n4420 GNDA.n4419 0.063
R14248 GNDA.n4311 GNDA.n4310 0.063
R14249 GNDA.n4317 GNDA.n4316 0.063
R14250 GNDA.n4323 GNDA.n4322 0.063
R14251 GNDA.n4153 GNDA.n4152 0.063
R14252 GNDA.n4164 GNDA.n505 0.063
R14253 GNDA.n4183 GNDA.n4182 0.063
R14254 GNDA.n3977 GNDA.n778 0.063
R14255 GNDA.n3970 GNDA.n3969 0.063
R14256 GNDA.n3959 GNDA.n793 0.063
R14257 GNDA.n4049 GNDA.n4043 0.063
R14258 GNDA.n4018 GNDA.n749 0.063
R14259 GNDA.n3584 GNDA.n3583 0.063
R14260 GNDA.n3593 GNDA.n3559 0.063
R14261 GNDA.n3608 GNDA.n3607 0.063
R14262 GNDA.n3900 GNDA.n3899 0.063
R14263 GNDA.n3909 GNDA.n825 0.063
R14264 GNDA.n3924 GNDA.n3923 0.063
R14265 GNDA.n911 GNDA.n847 0.063
R14266 GNDA.n904 GNDA.n903 0.063
R14267 GNDA.n893 GNDA.n871 0.063
R14268 GNDA.n3688 GNDA.n3687 0.063
R14269 GNDA.n3697 GNDA.n3664 0.063
R14270 GNDA.n3712 GNDA.n3711 0.063
R14271 GNDA.n3757 GNDA.n3756 0.063
R14272 GNDA.n3766 GNDA.n3733 0.063
R14273 GNDA.n3781 GNDA.n3780 0.063
R14274 GNDA.n3814 GNDA.n3813 0.063
R14275 GNDA.n3825 GNDA.n3798 0.063
R14276 GNDA.n3844 GNDA.n3843 0.063
R14277 GNDA.n3465 GNDA.n3401 0.063
R14278 GNDA.n3458 GNDA.n3457 0.063
R14279 GNDA.n3447 GNDA.n3425 0.063
R14280 GNDA.n3502 GNDA.n3501 0.063
R14281 GNDA.n3511 GNDA.n962 0.063
R14282 GNDA.n3526 GNDA.n3525 0.063
R14283 GNDA.n2823 GNDA.n2822 0.063
R14284 GNDA.n2832 GNDA.n2799 0.063
R14285 GNDA.n2847 GNDA.n2846 0.063
R14286 GNDA.n2892 GNDA.n2891 0.063
R14287 GNDA.n2901 GNDA.n2868 0.063
R14288 GNDA.n2916 GNDA.n2915 0.063
R14289 GNDA.n2961 GNDA.n2960 0.063
R14290 GNDA.n2970 GNDA.n2937 0.063
R14291 GNDA.n2985 GNDA.n2984 0.063
R14292 GNDA.n3030 GNDA.n3029 0.063
R14293 GNDA.n3039 GNDA.n3006 0.063
R14294 GNDA.n3054 GNDA.n3053 0.063
R14295 GNDA.n3099 GNDA.n3098 0.063
R14296 GNDA.n3108 GNDA.n3075 0.063
R14297 GNDA.n3123 GNDA.n3122 0.063
R14298 GNDA.n3168 GNDA.n3167 0.063
R14299 GNDA.n3177 GNDA.n3144 0.063
R14300 GNDA.n3192 GNDA.n3191 0.063
R14301 GNDA.n3237 GNDA.n3236 0.063
R14302 GNDA.n3246 GNDA.n3213 0.063
R14303 GNDA.n3261 GNDA.n3260 0.063
R14304 GNDA.n3294 GNDA.n3293 0.063
R14305 GNDA.n3305 GNDA.n3278 0.063
R14306 GNDA.n3324 GNDA.n3323 0.063
R14307 GNDA.n583 GNDA.n519 0.063
R14308 GNDA.n576 GNDA.n575 0.063
R14309 GNDA.n565 GNDA.n543 0.063
R14310 GNDA.n1499 GNDA.n1482 0.063
R14311 GNDA.n1518 GNDA.n1517 0.063
R14312 GNDA.n1529 GNDA.n1470 0.063
R14313 GNDA.n2563 GNDA.n2562 0.063
R14314 GNDA.n2553 GNDA.n2552 0.063
R14315 GNDA.n4134 GNDA.n481 0.0629369
R14316 GNDA.n4056 GNDA.n4055 0.0626438
R14317 GNDA.n4048 GNDA.n751 0.0626438
R14318 GNDA.n668 GNDA.n667 0.0626438
R14319 GNDA.n731 GNDA.n645 0.0626438
R14320 GNDA.n685 GNDA.n684 0.0626438
R14321 GNDA.n4118 GNDA.n605 0.0626438
R14322 GNDA.n1895 GNDA.n1894 0.0626438
R14323 GNDA.n1925 GNDA.n1919 0.0626438
R14324 GNDA.n1460 GNDA.n358 0.0626438
R14325 GNDA.n4043 GNDA.n4042 0.0577917
R14326 GNDA.n4020 GNDA.n4018 0.0577917
R14327 GNDA.n4674 GNDA.n4673 0.0553333
R14328 GNDA.n4688 GNDA.n4687 0.0553333
R14329 GNDA.n4704 GNDA.n4703 0.0553333
R14330 GNDA.n4718 GNDA.n4717 0.0553333
R14331 GNDA.n4598 GNDA.n4597 0.0553333
R14332 GNDA.n4612 GNDA.n4611 0.0553333
R14333 GNDA.n4628 GNDA.n4627 0.0553333
R14334 GNDA.n4642 GNDA.n4641 0.0553333
R14335 GNDA.n4547 GNDA.n4546 0.0553333
R14336 GNDA.n4538 GNDA.n4537 0.0553333
R14337 GNDA.n4529 GNDA.n4528 0.0553333
R14338 GNDA.n4520 GNDA.n4519 0.0553333
R14339 GNDA.n4758 GNDA.n4757 0.0553333
R14340 GNDA.n4772 GNDA.n4771 0.0553333
R14341 GNDA.n4788 GNDA.n4787 0.0553333
R14342 GNDA.n4802 GNDA.n4801 0.0553333
R14343 GNDA.n4222 GNDA.n4221 0.0553333
R14344 GNDA.n4236 GNDA.n4235 0.0553333
R14345 GNDA.n4252 GNDA.n4251 0.0553333
R14346 GNDA.n4266 GNDA.n4265 0.0553333
R14347 GNDA.n4823 GNDA.n4822 0.0553333
R14348 GNDA.n4837 GNDA.n4836 0.0553333
R14349 GNDA.n4853 GNDA.n4852 0.0553333
R14350 GNDA.n4867 GNDA.n4866 0.0553333
R14351 GNDA.n4383 GNDA.n4382 0.0553333
R14352 GNDA.n4397 GNDA.n4396 0.0553333
R14353 GNDA.n4413 GNDA.n4412 0.0553333
R14354 GNDA.n4427 GNDA.n4426 0.0553333
R14355 GNDA.n4359 GNDA.n4358 0.0553333
R14356 GNDA.n4350 GNDA.n4349 0.0553333
R14357 GNDA.n4341 GNDA.n4340 0.0553333
R14358 GNDA.n4332 GNDA.n4331 0.0553333
R14359 GNDA.n4146 GNDA.n4145 0.0553333
R14360 GNDA.n4160 GNDA.n4159 0.0553333
R14361 GNDA.n4176 GNDA.n4175 0.0553333
R14362 GNDA.n4190 GNDA.n4189 0.0553333
R14363 GNDA.n3936 GNDA.n776 0.0553333
R14364 GNDA.n785 GNDA.n784 0.0553333
R14365 GNDA.n3945 GNDA.n791 0.0553333
R14366 GNDA.n800 GNDA.n799 0.0553333
R14367 GNDA.n3570 GNDA.n3569 0.0553333
R14368 GNDA.n3589 GNDA.n3588 0.0553333
R14369 GNDA.n3558 GNDA.n3557 0.0553333
R14370 GNDA.n3613 GNDA.n3612 0.0553333
R14371 GNDA.n836 GNDA.n835 0.0553333
R14372 GNDA.n3905 GNDA.n3904 0.0553333
R14373 GNDA.n824 GNDA.n823 0.0553333
R14374 GNDA.n3929 GNDA.n3928 0.0553333
R14375 GNDA.n848 GNDA.n845 0.0553333
R14376 GNDA.n859 GNDA.n858 0.0553333
R14377 GNDA.n872 GNDA.n869 0.0553333
R14378 GNDA.n883 GNDA.n882 0.0553333
R14379 GNDA.n3675 GNDA.n3674 0.0553333
R14380 GNDA.n3693 GNDA.n3692 0.0553333
R14381 GNDA.n3663 GNDA.n3662 0.0553333
R14382 GNDA.n3717 GNDA.n3716 0.0553333
R14383 GNDA.n3744 GNDA.n3743 0.0553333
R14384 GNDA.n3762 GNDA.n3761 0.0553333
R14385 GNDA.n3732 GNDA.n3731 0.0553333
R14386 GNDA.n3786 GNDA.n3785 0.0553333
R14387 GNDA.n3807 GNDA.n3806 0.0553333
R14388 GNDA.n3821 GNDA.n3820 0.0553333
R14389 GNDA.n3837 GNDA.n3836 0.0553333
R14390 GNDA.n3851 GNDA.n3850 0.0553333
R14391 GNDA.n3402 GNDA.n3399 0.0553333
R14392 GNDA.n3413 GNDA.n3412 0.0553333
R14393 GNDA.n3426 GNDA.n3423 0.0553333
R14394 GNDA.n3437 GNDA.n3436 0.0553333
R14395 GNDA.n973 GNDA.n972 0.0553333
R14396 GNDA.n3507 GNDA.n3506 0.0553333
R14397 GNDA.n961 GNDA.n960 0.0553333
R14398 GNDA.n3531 GNDA.n3530 0.0553333
R14399 GNDA.n2810 GNDA.n2809 0.0553333
R14400 GNDA.n2828 GNDA.n2827 0.0553333
R14401 GNDA.n2798 GNDA.n2797 0.0553333
R14402 GNDA.n2852 GNDA.n2851 0.0553333
R14403 GNDA.n2879 GNDA.n2878 0.0553333
R14404 GNDA.n2897 GNDA.n2896 0.0553333
R14405 GNDA.n2867 GNDA.n2866 0.0553333
R14406 GNDA.n2921 GNDA.n2920 0.0553333
R14407 GNDA.n2948 GNDA.n2947 0.0553333
R14408 GNDA.n2966 GNDA.n2965 0.0553333
R14409 GNDA.n2936 GNDA.n2935 0.0553333
R14410 GNDA.n2990 GNDA.n2989 0.0553333
R14411 GNDA.n3017 GNDA.n3016 0.0553333
R14412 GNDA.n3035 GNDA.n3034 0.0553333
R14413 GNDA.n3005 GNDA.n3004 0.0553333
R14414 GNDA.n3059 GNDA.n3058 0.0553333
R14415 GNDA.n3086 GNDA.n3085 0.0553333
R14416 GNDA.n3104 GNDA.n3103 0.0553333
R14417 GNDA.n3074 GNDA.n3073 0.0553333
R14418 GNDA.n3128 GNDA.n3127 0.0553333
R14419 GNDA.n3155 GNDA.n3154 0.0553333
R14420 GNDA.n3173 GNDA.n3172 0.0553333
R14421 GNDA.n3143 GNDA.n3142 0.0553333
R14422 GNDA.n3197 GNDA.n3196 0.0553333
R14423 GNDA.n3224 GNDA.n3223 0.0553333
R14424 GNDA.n3242 GNDA.n3241 0.0553333
R14425 GNDA.n3212 GNDA.n3211 0.0553333
R14426 GNDA.n3266 GNDA.n3265 0.0553333
R14427 GNDA.n3287 GNDA.n3286 0.0553333
R14428 GNDA.n3301 GNDA.n3300 0.0553333
R14429 GNDA.n3317 GNDA.n3316 0.0553333
R14430 GNDA.n3331 GNDA.n3330 0.0553333
R14431 GNDA.n517 GNDA.n516 0.0553333
R14432 GNDA.n522 GNDA.n521 0.0553333
R14433 GNDA.n530 GNDA.n529 0.0553333
R14434 GNDA.n533 GNDA.n532 0.0553333
R14435 GNDA.n541 GNDA.n540 0.0553333
R14436 GNDA.n546 GNDA.n545 0.0553333
R14437 GNDA.n554 GNDA.n553 0.0553333
R14438 GNDA.n557 GNDA.n556 0.0553333
R14439 GNDA.n1495 GNDA.n1493 0.0553333
R14440 GNDA.n1511 GNDA.n1480 0.0553333
R14441 GNDA.n1525 GNDA.n1523 0.0553333
R14442 GNDA.n1541 GNDA.n1468 0.0553333
R14443 GNDA.n1368 GNDA.n1367 0.0553333
R14444 GNDA.n1382 GNDA.n1381 0.0553333
R14445 GNDA.n1398 GNDA.n1397 0.0553333
R14446 GNDA.n1412 GNDA.n1411 0.0553333
R14447 GNDA.n2505 GNDA 0.0517
R14448 GNDA.n2021 GNDA 0.0517
R14449 GNDA GNDA.n202 0.0517
R14450 GNDA.n2275 GNDA 0.0517
R14451 GNDA GNDA.n5187 0.0517
R14452 GNDA GNDA.n5466 0.0517
R14453 GNDA.n5044 GNDA 0.0517
R14454 GNDA.n1880 GNDA 0.0517
R14455 GNDA GNDA.n0 0.0517
R14456 GNDA.n4724 GNDA.n4565 0.0514167
R14457 GNDA.n4678 GNDA.n4677 0.0514167
R14458 GNDA.n4684 GNDA.n4683 0.0514167
R14459 GNDA.n4694 GNDA.n4693 0.0514167
R14460 GNDA.n4698 GNDA.n4697 0.0514167
R14461 GNDA.n4708 GNDA.n4707 0.0514167
R14462 GNDA.n4714 GNDA.n4713 0.0514167
R14463 GNDA.n4722 GNDA.n4659 0.0514167
R14464 GNDA.n4592 GNDA.n4566 0.0514167
R14465 GNDA.n4602 GNDA.n4601 0.0514167
R14466 GNDA.n4608 GNDA.n4607 0.0514167
R14467 GNDA.n4618 GNDA.n4617 0.0514167
R14468 GNDA.n4622 GNDA.n4621 0.0514167
R14469 GNDA.n4632 GNDA.n4631 0.0514167
R14470 GNDA.n4638 GNDA.n4637 0.0514167
R14471 GNDA.n4646 GNDA.n4578 0.0514167
R14472 GNDA.n4550 GNDA.n4549 0.0514167
R14473 GNDA.n4544 GNDA.n4543 0.0514167
R14474 GNDA.n4541 GNDA.n4540 0.0514167
R14475 GNDA.n4535 GNDA.n4534 0.0514167
R14476 GNDA.n4532 GNDA.n4531 0.0514167
R14477 GNDA.n4526 GNDA.n4525 0.0514167
R14478 GNDA.n4523 GNDA.n4522 0.0514167
R14479 GNDA.n4517 GNDA.n4516 0.0514167
R14480 GNDA.n4752 GNDA.n4444 0.0514167
R14481 GNDA.n4762 GNDA.n4761 0.0514167
R14482 GNDA.n4768 GNDA.n4767 0.0514167
R14483 GNDA.n4778 GNDA.n4777 0.0514167
R14484 GNDA.n4782 GNDA.n4781 0.0514167
R14485 GNDA.n4792 GNDA.n4791 0.0514167
R14486 GNDA.n4798 GNDA.n4797 0.0514167
R14487 GNDA.n4806 GNDA.n4457 0.0514167
R14488 GNDA.n4272 GNDA.n485 0.0514167
R14489 GNDA.n4226 GNDA.n4225 0.0514167
R14490 GNDA.n4232 GNDA.n4231 0.0514167
R14491 GNDA.n4242 GNDA.n4241 0.0514167
R14492 GNDA.n4246 GNDA.n4245 0.0514167
R14493 GNDA.n4256 GNDA.n4255 0.0514167
R14494 GNDA.n4262 GNDA.n4261 0.0514167
R14495 GNDA.n4270 GNDA.n4207 0.0514167
R14496 GNDA.n4873 GNDA.n445 0.0514167
R14497 GNDA.n4827 GNDA.n4826 0.0514167
R14498 GNDA.n4833 GNDA.n4832 0.0514167
R14499 GNDA.n4843 GNDA.n4842 0.0514167
R14500 GNDA.n4847 GNDA.n4846 0.0514167
R14501 GNDA.n4857 GNDA.n4856 0.0514167
R14502 GNDA.n4863 GNDA.n4862 0.0514167
R14503 GNDA.n4871 GNDA.n4808 0.0514167
R14504 GNDA.n4377 GNDA.n447 0.0514167
R14505 GNDA.n4387 GNDA.n4386 0.0514167
R14506 GNDA.n4393 GNDA.n4392 0.0514167
R14507 GNDA.n4403 GNDA.n4402 0.0514167
R14508 GNDA.n4407 GNDA.n4406 0.0514167
R14509 GNDA.n4417 GNDA.n4416 0.0514167
R14510 GNDA.n4423 GNDA.n4422 0.0514167
R14511 GNDA.n4431 GNDA.n459 0.0514167
R14512 GNDA.n4362 GNDA.n4361 0.0514167
R14513 GNDA.n4356 GNDA.n4355 0.0514167
R14514 GNDA.n4353 GNDA.n4352 0.0514167
R14515 GNDA.n4347 GNDA.n4346 0.0514167
R14516 GNDA.n4344 GNDA.n4343 0.0514167
R14517 GNDA.n4338 GNDA.n4337 0.0514167
R14518 GNDA.n4335 GNDA.n4334 0.0514167
R14519 GNDA.n4329 GNDA.n4328 0.0514167
R14520 GNDA.n4140 GNDA.n487 0.0514167
R14521 GNDA.n4150 GNDA.n4149 0.0514167
R14522 GNDA.n4156 GNDA.n4155 0.0514167
R14523 GNDA.n4166 GNDA.n4165 0.0514167
R14524 GNDA.n4170 GNDA.n4169 0.0514167
R14525 GNDA.n4180 GNDA.n4179 0.0514167
R14526 GNDA.n4186 GNDA.n4185 0.0514167
R14527 GNDA.n4194 GNDA.n499 0.0514167
R14528 GNDA.n775 GNDA.n774 0.0514167
R14529 GNDA.n780 GNDA.n779 0.0514167
R14530 GNDA.n3939 GNDA.n781 0.0514167
R14531 GNDA.n3942 GNDA.n786 0.0514167
R14532 GNDA.n790 GNDA.n789 0.0514167
R14533 GNDA.n795 GNDA.n794 0.0514167
R14534 GNDA.n3948 GNDA.n796 0.0514167
R14535 GNDA.n3952 GNDA.n801 0.0514167
R14536 GNDA.n3573 GNDA.n3537 0.0514167
R14537 GNDA.n3581 GNDA.n3580 0.0514167
R14538 GNDA.n3566 GNDA.n3565 0.0514167
R14539 GNDA.n3562 GNDA.n3561 0.0514167
R14540 GNDA.n3597 GNDA.n3596 0.0514167
R14541 GNDA.n3605 GNDA.n3604 0.0514167
R14542 GNDA.n3554 GNDA.n3553 0.0514167
R14543 GNDA.n3617 GNDA.n3549 0.0514167
R14544 GNDA.n3889 GNDA.n803 0.0514167
R14545 GNDA.n3897 GNDA.n3896 0.0514167
R14546 GNDA.n832 GNDA.n831 0.0514167
R14547 GNDA.n828 GNDA.n827 0.0514167
R14548 GNDA.n3913 GNDA.n3912 0.0514167
R14549 GNDA.n3921 GNDA.n3920 0.0514167
R14550 GNDA.n820 GNDA.n819 0.0514167
R14551 GNDA.n3933 GNDA.n815 0.0514167
R14552 GNDA.n843 GNDA.n842 0.0514167
R14553 GNDA.n851 GNDA.n850 0.0514167
R14554 GNDA.n856 GNDA.n853 0.0514167
R14555 GNDA.n864 GNDA.n861 0.0514167
R14556 GNDA.n867 GNDA.n866 0.0514167
R14557 GNDA.n875 GNDA.n874 0.0514167
R14558 GNDA.n880 GNDA.n877 0.0514167
R14559 GNDA.n886 GNDA.n885 0.0514167
R14560 GNDA.n3677 GNDA.n3642 0.0514167
R14561 GNDA.n3685 GNDA.n3684 0.0514167
R14562 GNDA.n3671 GNDA.n3670 0.0514167
R14563 GNDA.n3667 GNDA.n3666 0.0514167
R14564 GNDA.n3701 GNDA.n3700 0.0514167
R14565 GNDA.n3709 GNDA.n3708 0.0514167
R14566 GNDA.n3659 GNDA.n3658 0.0514167
R14567 GNDA.n3721 GNDA.n3654 0.0514167
R14568 GNDA.n3746 GNDA.n3630 0.0514167
R14569 GNDA.n3754 GNDA.n3753 0.0514167
R14570 GNDA.n3740 GNDA.n3739 0.0514167
R14571 GNDA.n3736 GNDA.n3735 0.0514167
R14572 GNDA.n3770 GNDA.n3769 0.0514167
R14573 GNDA.n3778 GNDA.n3777 0.0514167
R14574 GNDA.n3728 GNDA.n3727 0.0514167
R14575 GNDA.n3790 GNDA.n3723 0.0514167
R14576 GNDA.n3857 GNDA.n938 0.0514167
R14577 GNDA.n3811 GNDA.n3810 0.0514167
R14578 GNDA.n3817 GNDA.n3816 0.0514167
R14579 GNDA.n3827 GNDA.n3826 0.0514167
R14580 GNDA.n3831 GNDA.n3830 0.0514167
R14581 GNDA.n3841 GNDA.n3840 0.0514167
R14582 GNDA.n3847 GNDA.n3846 0.0514167
R14583 GNDA.n3855 GNDA.n3792 0.0514167
R14584 GNDA.n3397 GNDA.n3396 0.0514167
R14585 GNDA.n3405 GNDA.n3404 0.0514167
R14586 GNDA.n3410 GNDA.n3407 0.0514167
R14587 GNDA.n3418 GNDA.n3415 0.0514167
R14588 GNDA.n3421 GNDA.n3420 0.0514167
R14589 GNDA.n3429 GNDA.n3428 0.0514167
R14590 GNDA.n3434 GNDA.n3431 0.0514167
R14591 GNDA.n3440 GNDA.n3439 0.0514167
R14592 GNDA.n3491 GNDA.n940 0.0514167
R14593 GNDA.n3499 GNDA.n3498 0.0514167
R14594 GNDA.n969 GNDA.n968 0.0514167
R14595 GNDA.n965 GNDA.n964 0.0514167
R14596 GNDA.n3515 GNDA.n3514 0.0514167
R14597 GNDA.n3523 GNDA.n3522 0.0514167
R14598 GNDA.n957 GNDA.n956 0.0514167
R14599 GNDA.n3535 GNDA.n952 0.0514167
R14600 GNDA.n2812 GNDA.n2777 0.0514167
R14601 GNDA.n2820 GNDA.n2819 0.0514167
R14602 GNDA.n2806 GNDA.n2805 0.0514167
R14603 GNDA.n2802 GNDA.n2801 0.0514167
R14604 GNDA.n2836 GNDA.n2835 0.0514167
R14605 GNDA.n2844 GNDA.n2843 0.0514167
R14606 GNDA.n2794 GNDA.n2793 0.0514167
R14607 GNDA.n2856 GNDA.n2789 0.0514167
R14608 GNDA.n2881 GNDA.n2765 0.0514167
R14609 GNDA.n2889 GNDA.n2888 0.0514167
R14610 GNDA.n2875 GNDA.n2874 0.0514167
R14611 GNDA.n2871 GNDA.n2870 0.0514167
R14612 GNDA.n2905 GNDA.n2904 0.0514167
R14613 GNDA.n2913 GNDA.n2912 0.0514167
R14614 GNDA.n2863 GNDA.n2862 0.0514167
R14615 GNDA.n2925 GNDA.n2858 0.0514167
R14616 GNDA.n2950 GNDA.n2753 0.0514167
R14617 GNDA.n2958 GNDA.n2957 0.0514167
R14618 GNDA.n2944 GNDA.n2943 0.0514167
R14619 GNDA.n2940 GNDA.n2939 0.0514167
R14620 GNDA.n2974 GNDA.n2973 0.0514167
R14621 GNDA.n2982 GNDA.n2981 0.0514167
R14622 GNDA.n2932 GNDA.n2931 0.0514167
R14623 GNDA.n2994 GNDA.n2927 0.0514167
R14624 GNDA.n3019 GNDA.n2741 0.0514167
R14625 GNDA.n3027 GNDA.n3026 0.0514167
R14626 GNDA.n3013 GNDA.n3012 0.0514167
R14627 GNDA.n3009 GNDA.n3008 0.0514167
R14628 GNDA.n3043 GNDA.n3042 0.0514167
R14629 GNDA.n3051 GNDA.n3050 0.0514167
R14630 GNDA.n3001 GNDA.n3000 0.0514167
R14631 GNDA.n3063 GNDA.n2996 0.0514167
R14632 GNDA.n3088 GNDA.n2729 0.0514167
R14633 GNDA.n3096 GNDA.n3095 0.0514167
R14634 GNDA.n3082 GNDA.n3081 0.0514167
R14635 GNDA.n3078 GNDA.n3077 0.0514167
R14636 GNDA.n3112 GNDA.n3111 0.0514167
R14637 GNDA.n3120 GNDA.n3119 0.0514167
R14638 GNDA.n3070 GNDA.n3069 0.0514167
R14639 GNDA.n3132 GNDA.n3065 0.0514167
R14640 GNDA.n3157 GNDA.n2717 0.0514167
R14641 GNDA.n3165 GNDA.n3164 0.0514167
R14642 GNDA.n3151 GNDA.n3150 0.0514167
R14643 GNDA.n3147 GNDA.n3146 0.0514167
R14644 GNDA.n3181 GNDA.n3180 0.0514167
R14645 GNDA.n3189 GNDA.n3188 0.0514167
R14646 GNDA.n3139 GNDA.n3138 0.0514167
R14647 GNDA.n3201 GNDA.n3134 0.0514167
R14648 GNDA.n3226 GNDA.n2705 0.0514167
R14649 GNDA.n3234 GNDA.n3233 0.0514167
R14650 GNDA.n3220 GNDA.n3219 0.0514167
R14651 GNDA.n3216 GNDA.n3215 0.0514167
R14652 GNDA.n3250 GNDA.n3249 0.0514167
R14653 GNDA.n3258 GNDA.n3257 0.0514167
R14654 GNDA.n3208 GNDA.n3207 0.0514167
R14655 GNDA.n3270 GNDA.n3203 0.0514167
R14656 GNDA.n3337 GNDA.n1040 0.0514167
R14657 GNDA.n3291 GNDA.n3290 0.0514167
R14658 GNDA.n3297 GNDA.n3296 0.0514167
R14659 GNDA.n3307 GNDA.n3306 0.0514167
R14660 GNDA.n3311 GNDA.n3310 0.0514167
R14661 GNDA.n3321 GNDA.n3320 0.0514167
R14662 GNDA.n3327 GNDA.n3326 0.0514167
R14663 GNDA.n3335 GNDA.n3272 0.0514167
R14664 GNDA.n1491 GNDA.n1488 0.0514167
R14665 GNDA.n1501 GNDA.n1484 0.0514167
R14666 GNDA.n1505 GNDA.n1503 0.0514167
R14667 GNDA.n1515 GNDA.n1513 0.0514167
R14668 GNDA.n1521 GNDA.n1476 0.0514167
R14669 GNDA.n1531 GNDA.n1472 0.0514167
R14670 GNDA.n1535 GNDA.n1533 0.0514167
R14671 GNDA.n1544 GNDA.n1543 0.0514167
R14672 GNDA.n1362 GNDA.n1337 0.0514167
R14673 GNDA.n1372 GNDA.n1371 0.0514167
R14674 GNDA.n1378 GNDA.n1377 0.0514167
R14675 GNDA.n1388 GNDA.n1387 0.0514167
R14676 GNDA.n1392 GNDA.n1391 0.0514167
R14677 GNDA.n1402 GNDA.n1401 0.0514167
R14678 GNDA.n1408 GNDA.n1407 0.0514167
R14679 GNDA.n2578 GNDA.n1350 0.0514167
R14680 GNDA.n525 GNDA.n524 0.0475
R14681 GNDA.n538 GNDA.n537 0.0475
R14682 GNDA.n549 GNDA.n548 0.0475
R14683 GNDA.n4137 GNDA.n4136 0.0421667
R14684 GNDA.n766 GNDA.n764 0.0421667
R14685 GNDA.n3870 GNDA.n926 0.0421667
R14686 GNDA.n3875 GNDA.n922 0.0421667
R14687 GNDA.n3880 GNDA.n838 0.0421667
R14688 GNDA.n3882 GNDA.n772 0.0421667
R14689 GNDA.n3478 GNDA.n3477 0.0421667
R14690 GNDA.n4909 GNDA.n4887 0.0421667
R14691 GNDA.n4078 GNDA.n624 0.0421667
R14692 GNDA.n4086 GNDA.n618 0.0421667
R14693 GNDA.n4103 GNDA.n615 0.0421667
R14694 GNDA.n698 GNDA.n695 0.0421667
R14695 GNDA.n715 GNDA.n714 0.0421667
R14696 GNDA.n997 GNDA.n995 0.0421667
R14697 GNDA.n4073 GNDA.n628 0.0421667
R14698 GNDA.n3349 GNDA.n1031 0.0421667
R14699 GNDA.n3354 GNDA.n1027 0.0421667
R14700 GNDA.n3359 GNDA.n1023 0.0421667
R14701 GNDA.n3364 GNDA.n992 0.0421667
R14702 GNDA.n3369 GNDA.n988 0.0421667
R14703 GNDA.n3374 GNDA.n984 0.0421667
R14704 GNDA.n3379 GNDA.n980 0.0421667
R14705 GNDA.n3393 GNDA.n976 0.0421667
R14706 GNDA.n3484 GNDA.n975 0.0421667
R14707 GNDA.n598 GNDA.n511 0.0421667
R14708 GNDA.n4279 GNDA.n477 0.0421667
R14709 GNDA.n4369 GNDA.n474 0.0421667
R14710 GNDA.n472 GNDA.n441 0.0421667
R14711 GNDA.n4880 GNDA.n438 0.0421667
R14712 GNDA.n4883 GNDA.n437 0.0421667
R14713 GNDA.n4743 GNDA.n4742 0.0421667
R14714 GNDA.n4739 GNDA.n4738 0.0421667
R14715 GNDA.n4735 GNDA.n4734 0.0421667
R14716 GNDA.n4731 GNDA.n4730 0.0421667
R14717 GNDA.n1888 GNDA.n1555 0.0421667
R14718 GNDA.n1465 GNDA.n1459 0.0421667
R14719 GNDA.n4673 GNDA.n4648 0.028198
R14720 GNDA.n4677 GNDA.n4649 0.028198
R14721 GNDA.n4687 GNDA.n4651 0.028198
R14722 GNDA.n4693 GNDA.n4652 0.028198
R14723 GNDA.n4703 GNDA.n4654 0.028198
R14724 GNDA.n4707 GNDA.n4655 0.028198
R14725 GNDA.n4717 GNDA.n4657 0.028198
R14726 GNDA.n4659 GNDA.n4658 0.028198
R14727 GNDA.n4597 GNDA.n4567 0.028198
R14728 GNDA.n4601 GNDA.n4568 0.028198
R14729 GNDA.n4611 GNDA.n4570 0.028198
R14730 GNDA.n4617 GNDA.n4571 0.028198
R14731 GNDA.n4627 GNDA.n4573 0.028198
R14732 GNDA.n4631 GNDA.n4574 0.028198
R14733 GNDA.n4641 GNDA.n4576 0.028198
R14734 GNDA.n4578 GNDA.n4577 0.028198
R14735 GNDA.n4548 GNDA.n4547 0.028198
R14736 GNDA.n4545 GNDA.n4544 0.028198
R14737 GNDA.n4539 GNDA.n4538 0.028198
R14738 GNDA.n4536 GNDA.n4535 0.028198
R14739 GNDA.n4530 GNDA.n4529 0.028198
R14740 GNDA.n4527 GNDA.n4526 0.028198
R14741 GNDA.n4521 GNDA.n4520 0.028198
R14742 GNDA.n4518 GNDA.n4517 0.028198
R14743 GNDA.n4757 GNDA.n4445 0.028198
R14744 GNDA.n4761 GNDA.n4446 0.028198
R14745 GNDA.n4771 GNDA.n4448 0.028198
R14746 GNDA.n4777 GNDA.n4449 0.028198
R14747 GNDA.n4787 GNDA.n4451 0.028198
R14748 GNDA.n4791 GNDA.n4452 0.028198
R14749 GNDA.n4801 GNDA.n4454 0.028198
R14750 GNDA.n4457 GNDA.n4455 0.028198
R14751 GNDA.n4221 GNDA.n4196 0.028198
R14752 GNDA.n4225 GNDA.n4197 0.028198
R14753 GNDA.n4235 GNDA.n4199 0.028198
R14754 GNDA.n4241 GNDA.n4200 0.028198
R14755 GNDA.n4251 GNDA.n4202 0.028198
R14756 GNDA.n4255 GNDA.n4203 0.028198
R14757 GNDA.n4265 GNDA.n4205 0.028198
R14758 GNDA.n4207 GNDA.n4206 0.028198
R14759 GNDA.n4822 GNDA.n4433 0.028198
R14760 GNDA.n4826 GNDA.n4434 0.028198
R14761 GNDA.n4836 GNDA.n4436 0.028198
R14762 GNDA.n4842 GNDA.n4437 0.028198
R14763 GNDA.n4852 GNDA.n4439 0.028198
R14764 GNDA.n4856 GNDA.n4440 0.028198
R14765 GNDA.n4866 GNDA.n4442 0.028198
R14766 GNDA.n4808 GNDA.n4443 0.028198
R14767 GNDA.n4382 GNDA.n448 0.028198
R14768 GNDA.n4386 GNDA.n449 0.028198
R14769 GNDA.n4396 GNDA.n451 0.028198
R14770 GNDA.n4402 GNDA.n452 0.028198
R14771 GNDA.n4412 GNDA.n454 0.028198
R14772 GNDA.n4416 GNDA.n455 0.028198
R14773 GNDA.n4426 GNDA.n457 0.028198
R14774 GNDA.n459 GNDA.n458 0.028198
R14775 GNDA.n4360 GNDA.n4359 0.028198
R14776 GNDA.n4357 GNDA.n4356 0.028198
R14777 GNDA.n4351 GNDA.n4350 0.028198
R14778 GNDA.n4348 GNDA.n4347 0.028198
R14779 GNDA.n4342 GNDA.n4341 0.028198
R14780 GNDA.n4339 GNDA.n4338 0.028198
R14781 GNDA.n4333 GNDA.n4332 0.028198
R14782 GNDA.n4330 GNDA.n4329 0.028198
R14783 GNDA.n4145 GNDA.n488 0.028198
R14784 GNDA.n4149 GNDA.n489 0.028198
R14785 GNDA.n4159 GNDA.n491 0.028198
R14786 GNDA.n4165 GNDA.n492 0.028198
R14787 GNDA.n4175 GNDA.n494 0.028198
R14788 GNDA.n4179 GNDA.n495 0.028198
R14789 GNDA.n4189 GNDA.n497 0.028198
R14790 GNDA.n499 GNDA.n498 0.028198
R14791 GNDA.n3935 GNDA.n776 0.028198
R14792 GNDA.n3937 GNDA.n779 0.028198
R14793 GNDA.n3940 GNDA.n784 0.028198
R14794 GNDA.n3941 GNDA.n786 0.028198
R14795 GNDA.n3944 GNDA.n791 0.028198
R14796 GNDA.n3946 GNDA.n794 0.028198
R14797 GNDA.n3949 GNDA.n799 0.028198
R14798 GNDA.n3950 GNDA.n801 0.028198
R14799 GNDA.n3569 GNDA.n3538 0.028198
R14800 GNDA.n3580 GNDA.n3539 0.028198
R14801 GNDA.n3588 GNDA.n3541 0.028198
R14802 GNDA.n3561 GNDA.n3542 0.028198
R14803 GNDA.n3557 GNDA.n3544 0.028198
R14804 GNDA.n3604 GNDA.n3545 0.028198
R14805 GNDA.n3612 GNDA.n3547 0.028198
R14806 GNDA.n3549 GNDA.n3548 0.028198
R14807 GNDA.n835 GNDA.n804 0.028198
R14808 GNDA.n3896 GNDA.n805 0.028198
R14809 GNDA.n3904 GNDA.n807 0.028198
R14810 GNDA.n827 GNDA.n808 0.028198
R14811 GNDA.n823 GNDA.n810 0.028198
R14812 GNDA.n3920 GNDA.n811 0.028198
R14813 GNDA.n3928 GNDA.n813 0.028198
R14814 GNDA.n815 GNDA.n814 0.028198
R14815 GNDA.n845 GNDA.n844 0.028198
R14816 GNDA.n850 GNDA.n849 0.028198
R14817 GNDA.n858 GNDA.n857 0.028198
R14818 GNDA.n861 GNDA.n860 0.028198
R14819 GNDA.n869 GNDA.n868 0.028198
R14820 GNDA.n874 GNDA.n873 0.028198
R14821 GNDA.n882 GNDA.n881 0.028198
R14822 GNDA.n885 GNDA.n884 0.028198
R14823 GNDA.n3674 GNDA.n3643 0.028198
R14824 GNDA.n3684 GNDA.n3644 0.028198
R14825 GNDA.n3692 GNDA.n3646 0.028198
R14826 GNDA.n3666 GNDA.n3647 0.028198
R14827 GNDA.n3662 GNDA.n3649 0.028198
R14828 GNDA.n3708 GNDA.n3650 0.028198
R14829 GNDA.n3716 GNDA.n3652 0.028198
R14830 GNDA.n3654 GNDA.n3653 0.028198
R14831 GNDA.n3743 GNDA.n3631 0.028198
R14832 GNDA.n3753 GNDA.n3632 0.028198
R14833 GNDA.n3761 GNDA.n3634 0.028198
R14834 GNDA.n3735 GNDA.n3635 0.028198
R14835 GNDA.n3731 GNDA.n3637 0.028198
R14836 GNDA.n3777 GNDA.n3638 0.028198
R14837 GNDA.n3785 GNDA.n3640 0.028198
R14838 GNDA.n3723 GNDA.n3641 0.028198
R14839 GNDA.n3806 GNDA.n3619 0.028198
R14840 GNDA.n3810 GNDA.n3620 0.028198
R14841 GNDA.n3820 GNDA.n3622 0.028198
R14842 GNDA.n3826 GNDA.n3623 0.028198
R14843 GNDA.n3836 GNDA.n3625 0.028198
R14844 GNDA.n3840 GNDA.n3626 0.028198
R14845 GNDA.n3850 GNDA.n3628 0.028198
R14846 GNDA.n3792 GNDA.n3629 0.028198
R14847 GNDA.n3399 GNDA.n3398 0.028198
R14848 GNDA.n3404 GNDA.n3403 0.028198
R14849 GNDA.n3412 GNDA.n3411 0.028198
R14850 GNDA.n3415 GNDA.n3414 0.028198
R14851 GNDA.n3423 GNDA.n3422 0.028198
R14852 GNDA.n3428 GNDA.n3427 0.028198
R14853 GNDA.n3436 GNDA.n3435 0.028198
R14854 GNDA.n3439 GNDA.n3438 0.028198
R14855 GNDA.n972 GNDA.n941 0.028198
R14856 GNDA.n3498 GNDA.n942 0.028198
R14857 GNDA.n3506 GNDA.n944 0.028198
R14858 GNDA.n964 GNDA.n945 0.028198
R14859 GNDA.n960 GNDA.n947 0.028198
R14860 GNDA.n3522 GNDA.n948 0.028198
R14861 GNDA.n3530 GNDA.n950 0.028198
R14862 GNDA.n952 GNDA.n951 0.028198
R14863 GNDA.n2809 GNDA.n2778 0.028198
R14864 GNDA.n2819 GNDA.n2779 0.028198
R14865 GNDA.n2827 GNDA.n2781 0.028198
R14866 GNDA.n2801 GNDA.n2782 0.028198
R14867 GNDA.n2797 GNDA.n2784 0.028198
R14868 GNDA.n2843 GNDA.n2785 0.028198
R14869 GNDA.n2851 GNDA.n2787 0.028198
R14870 GNDA.n2789 GNDA.n2788 0.028198
R14871 GNDA.n2878 GNDA.n2766 0.028198
R14872 GNDA.n2888 GNDA.n2767 0.028198
R14873 GNDA.n2896 GNDA.n2769 0.028198
R14874 GNDA.n2870 GNDA.n2770 0.028198
R14875 GNDA.n2866 GNDA.n2772 0.028198
R14876 GNDA.n2912 GNDA.n2773 0.028198
R14877 GNDA.n2920 GNDA.n2775 0.028198
R14878 GNDA.n2858 GNDA.n2776 0.028198
R14879 GNDA.n2947 GNDA.n2754 0.028198
R14880 GNDA.n2957 GNDA.n2755 0.028198
R14881 GNDA.n2965 GNDA.n2757 0.028198
R14882 GNDA.n2939 GNDA.n2758 0.028198
R14883 GNDA.n2935 GNDA.n2760 0.028198
R14884 GNDA.n2981 GNDA.n2761 0.028198
R14885 GNDA.n2989 GNDA.n2763 0.028198
R14886 GNDA.n2927 GNDA.n2764 0.028198
R14887 GNDA.n3016 GNDA.n2742 0.028198
R14888 GNDA.n3026 GNDA.n2743 0.028198
R14889 GNDA.n3034 GNDA.n2745 0.028198
R14890 GNDA.n3008 GNDA.n2746 0.028198
R14891 GNDA.n3004 GNDA.n2748 0.028198
R14892 GNDA.n3050 GNDA.n2749 0.028198
R14893 GNDA.n3058 GNDA.n2751 0.028198
R14894 GNDA.n2996 GNDA.n2752 0.028198
R14895 GNDA.n3085 GNDA.n2730 0.028198
R14896 GNDA.n3095 GNDA.n2731 0.028198
R14897 GNDA.n3103 GNDA.n2733 0.028198
R14898 GNDA.n3077 GNDA.n2734 0.028198
R14899 GNDA.n3073 GNDA.n2736 0.028198
R14900 GNDA.n3119 GNDA.n2737 0.028198
R14901 GNDA.n3127 GNDA.n2739 0.028198
R14902 GNDA.n3065 GNDA.n2740 0.028198
R14903 GNDA.n3154 GNDA.n2718 0.028198
R14904 GNDA.n3164 GNDA.n2719 0.028198
R14905 GNDA.n3172 GNDA.n2721 0.028198
R14906 GNDA.n3146 GNDA.n2722 0.028198
R14907 GNDA.n3142 GNDA.n2724 0.028198
R14908 GNDA.n3188 GNDA.n2725 0.028198
R14909 GNDA.n3196 GNDA.n2727 0.028198
R14910 GNDA.n3134 GNDA.n2728 0.028198
R14911 GNDA.n3223 GNDA.n2706 0.028198
R14912 GNDA.n3233 GNDA.n2707 0.028198
R14913 GNDA.n3241 GNDA.n2709 0.028198
R14914 GNDA.n3215 GNDA.n2710 0.028198
R14915 GNDA.n3211 GNDA.n2712 0.028198
R14916 GNDA.n3257 GNDA.n2713 0.028198
R14917 GNDA.n3265 GNDA.n2715 0.028198
R14918 GNDA.n3203 GNDA.n2716 0.028198
R14919 GNDA.n3286 GNDA.n2694 0.028198
R14920 GNDA.n3290 GNDA.n2695 0.028198
R14921 GNDA.n3300 GNDA.n2697 0.028198
R14922 GNDA.n3306 GNDA.n2698 0.028198
R14923 GNDA.n3316 GNDA.n2700 0.028198
R14924 GNDA.n3320 GNDA.n2701 0.028198
R14925 GNDA.n3330 GNDA.n2703 0.028198
R14926 GNDA.n3272 GNDA.n2704 0.028198
R14927 GNDA.n3331 GNDA.n2704 0.028198
R14928 GNDA.n3327 GNDA.n2703 0.028198
R14929 GNDA.n3317 GNDA.n2701 0.028198
R14930 GNDA.n3311 GNDA.n2700 0.028198
R14931 GNDA.n3301 GNDA.n2698 0.028198
R14932 GNDA.n3297 GNDA.n2697 0.028198
R14933 GNDA.n3287 GNDA.n2695 0.028198
R14934 GNDA.n2694 GNDA.n1040 0.028198
R14935 GNDA.n3266 GNDA.n2716 0.028198
R14936 GNDA.n3208 GNDA.n2715 0.028198
R14937 GNDA.n3212 GNDA.n2713 0.028198
R14938 GNDA.n3250 GNDA.n2712 0.028198
R14939 GNDA.n3242 GNDA.n2710 0.028198
R14940 GNDA.n3220 GNDA.n2709 0.028198
R14941 GNDA.n3224 GNDA.n2707 0.028198
R14942 GNDA.n3226 GNDA.n2706 0.028198
R14943 GNDA.n3197 GNDA.n2728 0.028198
R14944 GNDA.n3139 GNDA.n2727 0.028198
R14945 GNDA.n3143 GNDA.n2725 0.028198
R14946 GNDA.n3181 GNDA.n2724 0.028198
R14947 GNDA.n3173 GNDA.n2722 0.028198
R14948 GNDA.n3151 GNDA.n2721 0.028198
R14949 GNDA.n3155 GNDA.n2719 0.028198
R14950 GNDA.n3157 GNDA.n2718 0.028198
R14951 GNDA.n3128 GNDA.n2740 0.028198
R14952 GNDA.n3070 GNDA.n2739 0.028198
R14953 GNDA.n3074 GNDA.n2737 0.028198
R14954 GNDA.n3112 GNDA.n2736 0.028198
R14955 GNDA.n3104 GNDA.n2734 0.028198
R14956 GNDA.n3082 GNDA.n2733 0.028198
R14957 GNDA.n3086 GNDA.n2731 0.028198
R14958 GNDA.n3088 GNDA.n2730 0.028198
R14959 GNDA.n3059 GNDA.n2752 0.028198
R14960 GNDA.n3001 GNDA.n2751 0.028198
R14961 GNDA.n3005 GNDA.n2749 0.028198
R14962 GNDA.n3043 GNDA.n2748 0.028198
R14963 GNDA.n3035 GNDA.n2746 0.028198
R14964 GNDA.n3013 GNDA.n2745 0.028198
R14965 GNDA.n3017 GNDA.n2743 0.028198
R14966 GNDA.n3019 GNDA.n2742 0.028198
R14967 GNDA.n2990 GNDA.n2764 0.028198
R14968 GNDA.n2932 GNDA.n2763 0.028198
R14969 GNDA.n2936 GNDA.n2761 0.028198
R14970 GNDA.n2974 GNDA.n2760 0.028198
R14971 GNDA.n2966 GNDA.n2758 0.028198
R14972 GNDA.n2944 GNDA.n2757 0.028198
R14973 GNDA.n2948 GNDA.n2755 0.028198
R14974 GNDA.n2950 GNDA.n2754 0.028198
R14975 GNDA.n2921 GNDA.n2776 0.028198
R14976 GNDA.n2863 GNDA.n2775 0.028198
R14977 GNDA.n2867 GNDA.n2773 0.028198
R14978 GNDA.n2905 GNDA.n2772 0.028198
R14979 GNDA.n2897 GNDA.n2770 0.028198
R14980 GNDA.n2875 GNDA.n2769 0.028198
R14981 GNDA.n2879 GNDA.n2767 0.028198
R14982 GNDA.n2881 GNDA.n2766 0.028198
R14983 GNDA.n2852 GNDA.n2788 0.028198
R14984 GNDA.n2794 GNDA.n2787 0.028198
R14985 GNDA.n2798 GNDA.n2785 0.028198
R14986 GNDA.n2836 GNDA.n2784 0.028198
R14987 GNDA.n2828 GNDA.n2782 0.028198
R14988 GNDA.n2806 GNDA.n2781 0.028198
R14989 GNDA.n2810 GNDA.n2779 0.028198
R14990 GNDA.n2812 GNDA.n2778 0.028198
R14991 GNDA.n3531 GNDA.n951 0.028198
R14992 GNDA.n957 GNDA.n950 0.028198
R14993 GNDA.n961 GNDA.n948 0.028198
R14994 GNDA.n3515 GNDA.n947 0.028198
R14995 GNDA.n3507 GNDA.n945 0.028198
R14996 GNDA.n969 GNDA.n944 0.028198
R14997 GNDA.n973 GNDA.n942 0.028198
R14998 GNDA.n3491 GNDA.n941 0.028198
R14999 GNDA.n3851 GNDA.n3629 0.028198
R15000 GNDA.n3847 GNDA.n3628 0.028198
R15001 GNDA.n3837 GNDA.n3626 0.028198
R15002 GNDA.n3831 GNDA.n3625 0.028198
R15003 GNDA.n3821 GNDA.n3623 0.028198
R15004 GNDA.n3817 GNDA.n3622 0.028198
R15005 GNDA.n3807 GNDA.n3620 0.028198
R15006 GNDA.n3619 GNDA.n938 0.028198
R15007 GNDA.n3786 GNDA.n3641 0.028198
R15008 GNDA.n3728 GNDA.n3640 0.028198
R15009 GNDA.n3732 GNDA.n3638 0.028198
R15010 GNDA.n3770 GNDA.n3637 0.028198
R15011 GNDA.n3762 GNDA.n3635 0.028198
R15012 GNDA.n3740 GNDA.n3634 0.028198
R15013 GNDA.n3744 GNDA.n3632 0.028198
R15014 GNDA.n3746 GNDA.n3631 0.028198
R15015 GNDA.n3717 GNDA.n3653 0.028198
R15016 GNDA.n3659 GNDA.n3652 0.028198
R15017 GNDA.n3663 GNDA.n3650 0.028198
R15018 GNDA.n3701 GNDA.n3649 0.028198
R15019 GNDA.n3693 GNDA.n3647 0.028198
R15020 GNDA.n3671 GNDA.n3646 0.028198
R15021 GNDA.n3675 GNDA.n3644 0.028198
R15022 GNDA.n3677 GNDA.n3643 0.028198
R15023 GNDA.n884 GNDA.n883 0.028198
R15024 GNDA.n881 GNDA.n880 0.028198
R15025 GNDA.n873 GNDA.n872 0.028198
R15026 GNDA.n868 GNDA.n867 0.028198
R15027 GNDA.n860 GNDA.n859 0.028198
R15028 GNDA.n857 GNDA.n856 0.028198
R15029 GNDA.n849 GNDA.n848 0.028198
R15030 GNDA.n844 GNDA.n843 0.028198
R15031 GNDA.n3929 GNDA.n814 0.028198
R15032 GNDA.n820 GNDA.n813 0.028198
R15033 GNDA.n824 GNDA.n811 0.028198
R15034 GNDA.n3913 GNDA.n810 0.028198
R15035 GNDA.n3905 GNDA.n808 0.028198
R15036 GNDA.n832 GNDA.n807 0.028198
R15037 GNDA.n836 GNDA.n805 0.028198
R15038 GNDA.n3889 GNDA.n804 0.028198
R15039 GNDA.n3438 GNDA.n3437 0.028198
R15040 GNDA.n3435 GNDA.n3434 0.028198
R15041 GNDA.n3427 GNDA.n3426 0.028198
R15042 GNDA.n3422 GNDA.n3421 0.028198
R15043 GNDA.n3414 GNDA.n3413 0.028198
R15044 GNDA.n3411 GNDA.n3410 0.028198
R15045 GNDA.n3403 GNDA.n3402 0.028198
R15046 GNDA.n3398 GNDA.n3397 0.028198
R15047 GNDA.n3613 GNDA.n3548 0.028198
R15048 GNDA.n3554 GNDA.n3547 0.028198
R15049 GNDA.n3558 GNDA.n3545 0.028198
R15050 GNDA.n3597 GNDA.n3544 0.028198
R15051 GNDA.n3589 GNDA.n3542 0.028198
R15052 GNDA.n3566 GNDA.n3541 0.028198
R15053 GNDA.n3570 GNDA.n3539 0.028198
R15054 GNDA.n3573 GNDA.n3538 0.028198
R15055 GNDA.n3950 GNDA.n800 0.028198
R15056 GNDA.n3949 GNDA.n3948 0.028198
R15057 GNDA.n3946 GNDA.n3945 0.028198
R15058 GNDA.n3944 GNDA.n790 0.028198
R15059 GNDA.n3941 GNDA.n785 0.028198
R15060 GNDA.n3940 GNDA.n3939 0.028198
R15061 GNDA.n3937 GNDA.n3936 0.028198
R15062 GNDA.n3935 GNDA.n775 0.028198
R15063 GNDA.n4190 GNDA.n498 0.028198
R15064 GNDA.n4186 GNDA.n497 0.028198
R15065 GNDA.n4176 GNDA.n495 0.028198
R15066 GNDA.n4170 GNDA.n494 0.028198
R15067 GNDA.n4160 GNDA.n492 0.028198
R15068 GNDA.n4156 GNDA.n491 0.028198
R15069 GNDA.n4146 GNDA.n489 0.028198
R15070 GNDA.n4140 GNDA.n488 0.028198
R15071 GNDA.n4331 GNDA.n4330 0.028198
R15072 GNDA.n4334 GNDA.n4333 0.028198
R15073 GNDA.n4340 GNDA.n4339 0.028198
R15074 GNDA.n4343 GNDA.n4342 0.028198
R15075 GNDA.n4349 GNDA.n4348 0.028198
R15076 GNDA.n4352 GNDA.n4351 0.028198
R15077 GNDA.n4358 GNDA.n4357 0.028198
R15078 GNDA.n4361 GNDA.n4360 0.028198
R15079 GNDA.n4427 GNDA.n458 0.028198
R15080 GNDA.n4423 GNDA.n457 0.028198
R15081 GNDA.n4413 GNDA.n455 0.028198
R15082 GNDA.n4407 GNDA.n454 0.028198
R15083 GNDA.n4397 GNDA.n452 0.028198
R15084 GNDA.n4393 GNDA.n451 0.028198
R15085 GNDA.n4383 GNDA.n449 0.028198
R15086 GNDA.n4377 GNDA.n448 0.028198
R15087 GNDA.n4867 GNDA.n4443 0.028198
R15088 GNDA.n4863 GNDA.n4442 0.028198
R15089 GNDA.n4853 GNDA.n4440 0.028198
R15090 GNDA.n4847 GNDA.n4439 0.028198
R15091 GNDA.n4837 GNDA.n4437 0.028198
R15092 GNDA.n4833 GNDA.n4436 0.028198
R15093 GNDA.n4823 GNDA.n4434 0.028198
R15094 GNDA.n4433 GNDA.n445 0.028198
R15095 GNDA.n4266 GNDA.n4206 0.028198
R15096 GNDA.n4262 GNDA.n4205 0.028198
R15097 GNDA.n4252 GNDA.n4203 0.028198
R15098 GNDA.n4246 GNDA.n4202 0.028198
R15099 GNDA.n4236 GNDA.n4200 0.028198
R15100 GNDA.n4232 GNDA.n4199 0.028198
R15101 GNDA.n4222 GNDA.n4197 0.028198
R15102 GNDA.n4196 GNDA.n485 0.028198
R15103 GNDA.n4802 GNDA.n4455 0.028198
R15104 GNDA.n4798 GNDA.n4454 0.028198
R15105 GNDA.n4788 GNDA.n4452 0.028198
R15106 GNDA.n4782 GNDA.n4451 0.028198
R15107 GNDA.n4772 GNDA.n4449 0.028198
R15108 GNDA.n4768 GNDA.n4448 0.028198
R15109 GNDA.n4758 GNDA.n4446 0.028198
R15110 GNDA.n4752 GNDA.n4445 0.028198
R15111 GNDA.n4519 GNDA.n4518 0.028198
R15112 GNDA.n4522 GNDA.n4521 0.028198
R15113 GNDA.n4528 GNDA.n4527 0.028198
R15114 GNDA.n4531 GNDA.n4530 0.028198
R15115 GNDA.n4537 GNDA.n4536 0.028198
R15116 GNDA.n4540 GNDA.n4539 0.028198
R15117 GNDA.n4546 GNDA.n4545 0.028198
R15118 GNDA.n4549 GNDA.n4548 0.028198
R15119 GNDA.n4642 GNDA.n4577 0.028198
R15120 GNDA.n4638 GNDA.n4576 0.028198
R15121 GNDA.n4628 GNDA.n4574 0.028198
R15122 GNDA.n4622 GNDA.n4573 0.028198
R15123 GNDA.n4612 GNDA.n4571 0.028198
R15124 GNDA.n4608 GNDA.n4570 0.028198
R15125 GNDA.n4598 GNDA.n4568 0.028198
R15126 GNDA.n4592 GNDA.n4567 0.028198
R15127 GNDA.n4718 GNDA.n4658 0.028198
R15128 GNDA.n4714 GNDA.n4657 0.028198
R15129 GNDA.n4704 GNDA.n4655 0.028198
R15130 GNDA.n4698 GNDA.n4654 0.028198
R15131 GNDA.n4688 GNDA.n4652 0.028198
R15132 GNDA.n4684 GNDA.n4651 0.028198
R15133 GNDA.n4674 GNDA.n4649 0.028198
R15134 GNDA.n4648 GNDA.n4565 0.028198
R15135 GNDA.n1493 GNDA.n1492 0.028198
R15136 GNDA.n1494 GNDA.n1484 0.028198
R15137 GNDA.n1504 GNDA.n1480 0.028198
R15138 GNDA.n1513 GNDA.n1512 0.028198
R15139 GNDA.n1523 GNDA.n1522 0.028198
R15140 GNDA.n1524 GNDA.n1472 0.028198
R15141 GNDA.n1534 GNDA.n1468 0.028198
R15142 GNDA.n1543 GNDA.n1542 0.028198
R15143 GNDA.n1367 GNDA.n1338 0.028198
R15144 GNDA.n1371 GNDA.n1339 0.028198
R15145 GNDA.n1381 GNDA.n1341 0.028198
R15146 GNDA.n1387 GNDA.n1342 0.028198
R15147 GNDA.n1397 GNDA.n1344 0.028198
R15148 GNDA.n1401 GNDA.n1345 0.028198
R15149 GNDA.n1411 GNDA.n1347 0.028198
R15150 GNDA.n1350 GNDA.n1348 0.028198
R15151 GNDA.n1412 GNDA.n1348 0.028198
R15152 GNDA.n1408 GNDA.n1347 0.028198
R15153 GNDA.n1398 GNDA.n1345 0.028198
R15154 GNDA.n1392 GNDA.n1344 0.028198
R15155 GNDA.n1382 GNDA.n1342 0.028198
R15156 GNDA.n1378 GNDA.n1341 0.028198
R15157 GNDA.n1368 GNDA.n1339 0.028198
R15158 GNDA.n1362 GNDA.n1338 0.028198
R15159 GNDA.n1542 GNDA.n1541 0.028198
R15160 GNDA.n1535 GNDA.n1534 0.028198
R15161 GNDA.n1525 GNDA.n1524 0.028198
R15162 GNDA.n1522 GNDA.n1521 0.028198
R15163 GNDA.n1512 GNDA.n1511 0.028198
R15164 GNDA.n1505 GNDA.n1504 0.028198
R15165 GNDA.n1495 GNDA.n1494 0.028198
R15166 GNDA.n1492 GNDA.n1491 0.028198
R15167 GNDA.n520 GNDA.n517 0.028198
R15168 GNDA.n531 GNDA.n530 0.028198
R15169 GNDA.n544 GNDA.n541 0.028198
R15170 GNDA.n555 GNDA.n554 0.028198
R15171 GNDA.n556 GNDA.n555 0.028198
R15172 GNDA.n545 GNDA.n544 0.028198
R15173 GNDA.n532 GNDA.n531 0.028198
R15174 GNDA.n521 GNDA.n520 0.028198
R15175 GNDA.n523 GNDA.n522 0.0262697
R15176 GNDA.n528 GNDA.n525 0.0262697
R15177 GNDA.n536 GNDA.n533 0.0262697
R15178 GNDA.n539 GNDA.n538 0.0262697
R15179 GNDA.n547 GNDA.n546 0.0262697
R15180 GNDA.n552 GNDA.n549 0.0262697
R15181 GNDA.n558 GNDA.n557 0.0262697
R15182 GNDA.n553 GNDA.n552 0.0262697
R15183 GNDA.n548 GNDA.n547 0.0262697
R15184 GNDA.n540 GNDA.n539 0.0262697
R15185 GNDA.n537 GNDA.n536 0.0262697
R15186 GNDA.n529 GNDA.n528 0.0262697
R15187 GNDA.n524 GNDA.n523 0.0262697
R15188 GNDA.n516 GNDA.n515 0.0262697
R15189 GNDA.n4683 GNDA.n4650 0.0243392
R15190 GNDA.n4697 GNDA.n4653 0.0243392
R15191 GNDA.n4713 GNDA.n4656 0.0243392
R15192 GNDA.n4607 GNDA.n4569 0.0243392
R15193 GNDA.n4621 GNDA.n4572 0.0243392
R15194 GNDA.n4637 GNDA.n4575 0.0243392
R15195 GNDA.n4542 GNDA.n4541 0.0243392
R15196 GNDA.n4533 GNDA.n4532 0.0243392
R15197 GNDA.n4524 GNDA.n4523 0.0243392
R15198 GNDA.n4767 GNDA.n4447 0.0243392
R15199 GNDA.n4781 GNDA.n4450 0.0243392
R15200 GNDA.n4797 GNDA.n4453 0.0243392
R15201 GNDA.n4231 GNDA.n4198 0.0243392
R15202 GNDA.n4245 GNDA.n4201 0.0243392
R15203 GNDA.n4261 GNDA.n4204 0.0243392
R15204 GNDA.n4832 GNDA.n4435 0.0243392
R15205 GNDA.n4846 GNDA.n4438 0.0243392
R15206 GNDA.n4862 GNDA.n4441 0.0243392
R15207 GNDA.n4392 GNDA.n450 0.0243392
R15208 GNDA.n4406 GNDA.n453 0.0243392
R15209 GNDA.n4422 GNDA.n456 0.0243392
R15210 GNDA.n4354 GNDA.n4353 0.0243392
R15211 GNDA.n4345 GNDA.n4344 0.0243392
R15212 GNDA.n4336 GNDA.n4335 0.0243392
R15213 GNDA.n4155 GNDA.n490 0.0243392
R15214 GNDA.n4169 GNDA.n493 0.0243392
R15215 GNDA.n4185 GNDA.n496 0.0243392
R15216 GNDA.n3938 GNDA.n781 0.0243392
R15217 GNDA.n3943 GNDA.n789 0.0243392
R15218 GNDA.n3947 GNDA.n796 0.0243392
R15219 GNDA.n3565 GNDA.n3540 0.0243392
R15220 GNDA.n3596 GNDA.n3543 0.0243392
R15221 GNDA.n3553 GNDA.n3546 0.0243392
R15222 GNDA.n831 GNDA.n806 0.0243392
R15223 GNDA.n3912 GNDA.n809 0.0243392
R15224 GNDA.n819 GNDA.n812 0.0243392
R15225 GNDA.n853 GNDA.n852 0.0243392
R15226 GNDA.n866 GNDA.n865 0.0243392
R15227 GNDA.n877 GNDA.n876 0.0243392
R15228 GNDA.n3670 GNDA.n3645 0.0243392
R15229 GNDA.n3700 GNDA.n3648 0.0243392
R15230 GNDA.n3658 GNDA.n3651 0.0243392
R15231 GNDA.n3739 GNDA.n3633 0.0243392
R15232 GNDA.n3769 GNDA.n3636 0.0243392
R15233 GNDA.n3727 GNDA.n3639 0.0243392
R15234 GNDA.n3816 GNDA.n3621 0.0243392
R15235 GNDA.n3830 GNDA.n3624 0.0243392
R15236 GNDA.n3846 GNDA.n3627 0.0243392
R15237 GNDA.n3407 GNDA.n3406 0.0243392
R15238 GNDA.n3420 GNDA.n3419 0.0243392
R15239 GNDA.n3431 GNDA.n3430 0.0243392
R15240 GNDA.n968 GNDA.n943 0.0243392
R15241 GNDA.n3514 GNDA.n946 0.0243392
R15242 GNDA.n956 GNDA.n949 0.0243392
R15243 GNDA.n2805 GNDA.n2780 0.0243392
R15244 GNDA.n2835 GNDA.n2783 0.0243392
R15245 GNDA.n2793 GNDA.n2786 0.0243392
R15246 GNDA.n2874 GNDA.n2768 0.0243392
R15247 GNDA.n2904 GNDA.n2771 0.0243392
R15248 GNDA.n2862 GNDA.n2774 0.0243392
R15249 GNDA.n2943 GNDA.n2756 0.0243392
R15250 GNDA.n2973 GNDA.n2759 0.0243392
R15251 GNDA.n2931 GNDA.n2762 0.0243392
R15252 GNDA.n3012 GNDA.n2744 0.0243392
R15253 GNDA.n3042 GNDA.n2747 0.0243392
R15254 GNDA.n3000 GNDA.n2750 0.0243392
R15255 GNDA.n3081 GNDA.n2732 0.0243392
R15256 GNDA.n3111 GNDA.n2735 0.0243392
R15257 GNDA.n3069 GNDA.n2738 0.0243392
R15258 GNDA.n3150 GNDA.n2720 0.0243392
R15259 GNDA.n3180 GNDA.n2723 0.0243392
R15260 GNDA.n3138 GNDA.n2726 0.0243392
R15261 GNDA.n3219 GNDA.n2708 0.0243392
R15262 GNDA.n3249 GNDA.n2711 0.0243392
R15263 GNDA.n3207 GNDA.n2714 0.0243392
R15264 GNDA.n3296 GNDA.n2696 0.0243392
R15265 GNDA.n3310 GNDA.n2699 0.0243392
R15266 GNDA.n3326 GNDA.n2702 0.0243392
R15267 GNDA.n3321 GNDA.n2702 0.0243392
R15268 GNDA.n3307 GNDA.n2699 0.0243392
R15269 GNDA.n3291 GNDA.n2696 0.0243392
R15270 GNDA.n3258 GNDA.n2714 0.0243392
R15271 GNDA.n3216 GNDA.n2711 0.0243392
R15272 GNDA.n3234 GNDA.n2708 0.0243392
R15273 GNDA.n3189 GNDA.n2726 0.0243392
R15274 GNDA.n3147 GNDA.n2723 0.0243392
R15275 GNDA.n3165 GNDA.n2720 0.0243392
R15276 GNDA.n3120 GNDA.n2738 0.0243392
R15277 GNDA.n3078 GNDA.n2735 0.0243392
R15278 GNDA.n3096 GNDA.n2732 0.0243392
R15279 GNDA.n3051 GNDA.n2750 0.0243392
R15280 GNDA.n3009 GNDA.n2747 0.0243392
R15281 GNDA.n3027 GNDA.n2744 0.0243392
R15282 GNDA.n2982 GNDA.n2762 0.0243392
R15283 GNDA.n2940 GNDA.n2759 0.0243392
R15284 GNDA.n2958 GNDA.n2756 0.0243392
R15285 GNDA.n2913 GNDA.n2774 0.0243392
R15286 GNDA.n2871 GNDA.n2771 0.0243392
R15287 GNDA.n2889 GNDA.n2768 0.0243392
R15288 GNDA.n2844 GNDA.n2786 0.0243392
R15289 GNDA.n2802 GNDA.n2783 0.0243392
R15290 GNDA.n2820 GNDA.n2780 0.0243392
R15291 GNDA.n3523 GNDA.n949 0.0243392
R15292 GNDA.n965 GNDA.n946 0.0243392
R15293 GNDA.n3499 GNDA.n943 0.0243392
R15294 GNDA.n3841 GNDA.n3627 0.0243392
R15295 GNDA.n3827 GNDA.n3624 0.0243392
R15296 GNDA.n3811 GNDA.n3621 0.0243392
R15297 GNDA.n3778 GNDA.n3639 0.0243392
R15298 GNDA.n3736 GNDA.n3636 0.0243392
R15299 GNDA.n3754 GNDA.n3633 0.0243392
R15300 GNDA.n3709 GNDA.n3651 0.0243392
R15301 GNDA.n3667 GNDA.n3648 0.0243392
R15302 GNDA.n3685 GNDA.n3645 0.0243392
R15303 GNDA.n876 GNDA.n875 0.0243392
R15304 GNDA.n865 GNDA.n864 0.0243392
R15305 GNDA.n852 GNDA.n851 0.0243392
R15306 GNDA.n3921 GNDA.n812 0.0243392
R15307 GNDA.n828 GNDA.n809 0.0243392
R15308 GNDA.n3897 GNDA.n806 0.0243392
R15309 GNDA.n3430 GNDA.n3429 0.0243392
R15310 GNDA.n3419 GNDA.n3418 0.0243392
R15311 GNDA.n3406 GNDA.n3405 0.0243392
R15312 GNDA.n3605 GNDA.n3546 0.0243392
R15313 GNDA.n3562 GNDA.n3543 0.0243392
R15314 GNDA.n3581 GNDA.n3540 0.0243392
R15315 GNDA.n3947 GNDA.n795 0.0243392
R15316 GNDA.n3943 GNDA.n3942 0.0243392
R15317 GNDA.n3938 GNDA.n780 0.0243392
R15318 GNDA.n4180 GNDA.n496 0.0243392
R15319 GNDA.n4166 GNDA.n493 0.0243392
R15320 GNDA.n4150 GNDA.n490 0.0243392
R15321 GNDA.n4337 GNDA.n4336 0.0243392
R15322 GNDA.n4346 GNDA.n4345 0.0243392
R15323 GNDA.n4355 GNDA.n4354 0.0243392
R15324 GNDA.n4417 GNDA.n456 0.0243392
R15325 GNDA.n4403 GNDA.n453 0.0243392
R15326 GNDA.n4387 GNDA.n450 0.0243392
R15327 GNDA.n4857 GNDA.n4441 0.0243392
R15328 GNDA.n4843 GNDA.n4438 0.0243392
R15329 GNDA.n4827 GNDA.n4435 0.0243392
R15330 GNDA.n4256 GNDA.n4204 0.0243392
R15331 GNDA.n4242 GNDA.n4201 0.0243392
R15332 GNDA.n4226 GNDA.n4198 0.0243392
R15333 GNDA.n4792 GNDA.n4453 0.0243392
R15334 GNDA.n4778 GNDA.n4450 0.0243392
R15335 GNDA.n4762 GNDA.n4447 0.0243392
R15336 GNDA.n4525 GNDA.n4524 0.0243392
R15337 GNDA.n4534 GNDA.n4533 0.0243392
R15338 GNDA.n4543 GNDA.n4542 0.0243392
R15339 GNDA.n4632 GNDA.n4575 0.0243392
R15340 GNDA.n4618 GNDA.n4572 0.0243392
R15341 GNDA.n4602 GNDA.n4569 0.0243392
R15342 GNDA.n4708 GNDA.n4656 0.0243392
R15343 GNDA.n4694 GNDA.n4653 0.0243392
R15344 GNDA.n4678 GNDA.n4650 0.0243392
R15345 GNDA.n1503 GNDA.n1502 0.0243392
R15346 GNDA.n1514 GNDA.n1476 0.0243392
R15347 GNDA.n1533 GNDA.n1532 0.0243392
R15348 GNDA.n1377 GNDA.n1340 0.0243392
R15349 GNDA.n1391 GNDA.n1343 0.0243392
R15350 GNDA.n1407 GNDA.n1346 0.0243392
R15351 GNDA.n1402 GNDA.n1346 0.0243392
R15352 GNDA.n1388 GNDA.n1343 0.0243392
R15353 GNDA.n1372 GNDA.n1340 0.0243392
R15354 GNDA.n1532 GNDA.n1531 0.0243392
R15355 GNDA.n1515 GNDA.n1514 0.0243392
R15356 GNDA.n1502 GNDA.n1501 0.0243392
R15357 GNDA.n4728 GNDA.n4561 0.0217373
R15358 GNDA.n4729 GNDA.n4561 0.0217373
R15359 GNDA.n4559 GNDA.n4556 0.0217373
R15360 GNDA.n4560 GNDA.n4556 0.0217373
R15361 GNDA.n4554 GNDA.n4470 0.0217373
R15362 GNDA.n4555 GNDA.n4470 0.0217373
R15363 GNDA.n4747 GNDA.n4744 0.0217373
R15364 GNDA.n4748 GNDA.n4747 0.0217373
R15365 GNDA.n442 GNDA.n440 0.0217373
R15366 GNDA.n442 GNDA.n439 0.0217373
R15367 GNDA.n4372 GNDA.n473 0.0217373
R15368 GNDA.n4373 GNDA.n4372 0.0217373
R15369 GNDA.n4283 GNDA.n476 0.0217373
R15370 GNDA.n4283 GNDA.n475 0.0217373
R15371 GNDA.n4008 GNDA.n758 0.0217373
R15372 GNDA.n770 GNDA.n763 0.0217373
R15373 GNDA.n771 GNDA.n761 0.0217373
R15374 GNDA.n3990 GNDA.n762 0.0217373
R15375 GNDA.n3989 GNDA.n761 0.0217373
R15376 GNDA.n4015 GNDA.n752 0.0217373
R15377 GNDA.n767 GNDA.n765 0.0217373
R15378 GNDA.n765 GNDA.n763 0.0217373
R15379 GNDA.n4012 GNDA.n753 0.0217373
R15380 GNDA.n933 GNDA.n756 0.0217373
R15381 GNDA.n754 GNDA.n752 0.0217373
R15382 GNDA.n4012 GNDA.n4011 0.0217373
R15383 GNDA.n758 GNDA.n757 0.0217373
R15384 GNDA.n934 GNDA.n933 0.0217373
R15385 GNDA.n3886 GNDA.n837 0.0217373
R15386 GNDA.n3879 GNDA.n840 0.0217373
R15387 GNDA.n3874 GNDA.n924 0.0217373
R15388 GNDA.n3869 GNDA.n928 0.0217373
R15389 GNDA.n3865 GNDA.n930 0.0217373
R15390 GNDA.n3866 GNDA.n927 0.0217373
R15391 GNDA.n3866 GNDA.n928 0.0217373
R15392 GNDA.n3871 GNDA.n923 0.0217373
R15393 GNDA.n3871 GNDA.n924 0.0217373
R15394 GNDA.n3876 GNDA.n839 0.0217373
R15395 GNDA.n3876 GNDA.n840 0.0217373
R15396 GNDA.n3883 GNDA.n3881 0.0217373
R15397 GNDA.n3881 GNDA.n837 0.0217373
R15398 GNDA.n3861 GNDA.n931 0.0217373
R15399 GNDA.n932 GNDA.n930 0.0217373
R15400 GNDA.n3861 GNDA.n3860 0.0217373
R15401 GNDA.n3488 GNDA.n974 0.0217373
R15402 GNDA.n4905 GNDA.n4904 0.0217373
R15403 GNDA.n4908 GNDA.n4907 0.0217373
R15404 GNDA.n4910 GNDA.n435 0.0217373
R15405 GNDA.n4881 GNDA.n436 0.0217373
R15406 GNDA.n4882 GNDA.n4881 0.0217373
R15407 GNDA.n4903 GNDA.n4888 0.0217373
R15408 GNDA.n4906 GNDA.n4905 0.0217373
R15409 GNDA.n654 GNDA.n653 0.0217373
R15410 GNDA.n4908 GNDA.n433 0.0217373
R15411 GNDA.n435 GNDA.n433 0.0217373
R15412 GNDA.n4079 GNDA.n4078 0.0217373
R15413 GNDA.n4092 GNDA.n4088 0.0217373
R15414 GNDA.n4097 GNDA.n4096 0.0217373
R15415 GNDA.n4099 GNDA.n616 0.0217373
R15416 GNDA.n4102 GNDA.n617 0.0217373
R15417 GNDA.n4095 GNDA.n4088 0.0217373
R15418 GNDA.n4098 GNDA.n4097 0.0217373
R15419 GNDA.n4083 GNDA.n618 0.0217373
R15420 GNDA.n4087 GNDA.n616 0.0217373
R15421 GNDA.n4087 GNDA.n617 0.0217373
R15422 GNDA.n699 GNDA.n698 0.0217373
R15423 GNDA.n713 GNDA.n609 0.0217373
R15424 GNDA.n610 GNDA.n607 0.0217373
R15425 GNDA.n4105 GNDA.n612 0.0217373
R15426 GNDA.n648 GNDA.n647 0.0217373
R15427 GNDA.n652 GNDA.n650 0.0217373
R15428 GNDA.n4111 GNDA.n608 0.0217373
R15429 GNDA.n4110 GNDA.n607 0.0217373
R15430 GNDA.n4107 GNDA.n613 0.0217373
R15431 GNDA.n4106 GNDA.n4105 0.0217373
R15432 GNDA.n660 GNDA.n659 0.0217373
R15433 GNDA.n657 GNDA.n647 0.0217373
R15434 GNDA.n653 GNDA.n651 0.0217373
R15435 GNDA.n706 GNDA.n680 0.0217373
R15436 GNDA.n716 GNDA.n712 0.0217373
R15437 GNDA.n713 GNDA.n712 0.0217373
R15438 GNDA.n703 GNDA.n681 0.0217373
R15439 GNDA.n697 GNDA.n683 0.0217373
R15440 GNDA.n697 GNDA.n696 0.0217373
R15441 GNDA.n622 GNDA.n621 0.0217373
R15442 GNDA.n622 GNDA.n619 0.0217373
R15443 GNDA.n625 GNDA.n623 0.0217373
R15444 GNDA.n4076 GNDA.n625 0.0217373
R15445 GNDA.n4075 GNDA.n4074 0.0217373
R15446 GNDA.n4072 GNDA.n629 0.0217373
R15447 GNDA.n682 GNDA.n680 0.0217373
R15448 GNDA.n703 GNDA.n702 0.0217373
R15449 GNDA.n701 GNDA.n683 0.0217373
R15450 GNDA.n696 GNDA.n620 0.0217373
R15451 GNDA.n700 GNDA.n699 0.0217373
R15452 GNDA.n4085 GNDA.n621 0.0217373
R15453 GNDA.n4082 GNDA.n619 0.0217373
R15454 GNDA.n4084 GNDA.n4083 0.0217373
R15455 GNDA.n4081 GNDA.n623 0.0217373
R15456 GNDA.n4077 GNDA.n4076 0.0217373
R15457 GNDA.n4080 GNDA.n4079 0.0217373
R15458 GNDA.n1011 GNDA.n998 0.0217373
R15459 GNDA.n1015 GNDA.n1014 0.0217373
R15460 GNDA.n1018 GNDA.n1017 0.0217373
R15461 GNDA.n1021 GNDA.n994 0.0217373
R15462 GNDA.n3360 GNDA.n1022 0.0217373
R15463 GNDA.n3360 GNDA.n993 0.0217373
R15464 GNDA.n1013 GNDA.n998 0.0217373
R15465 GNDA.n1016 GNDA.n1015 0.0217373
R15466 GNDA.n1017 GNDA.n996 0.0217373
R15467 GNDA.n996 GNDA.n994 0.0217373
R15468 GNDA.n4074 GNDA.n627 0.0217373
R15469 GNDA.n629 GNDA.n627 0.0217373
R15470 GNDA.n3378 GNDA.n982 0.0217373
R15471 GNDA.n3373 GNDA.n986 0.0217373
R15472 GNDA.n3368 GNDA.n990 0.0217373
R15473 GNDA.n3358 GNDA.n1025 0.0217373
R15474 GNDA.n3353 GNDA.n1029 0.0217373
R15475 GNDA.n3348 GNDA.n1033 0.0217373
R15476 GNDA.n3344 GNDA.n1035 0.0217373
R15477 GNDA.n3361 GNDA.n992 0.0217373
R15478 GNDA.n3345 GNDA.n1032 0.0217373
R15479 GNDA.n3345 GNDA.n1033 0.0217373
R15480 GNDA.n3350 GNDA.n1028 0.0217373
R15481 GNDA.n3350 GNDA.n1029 0.0217373
R15482 GNDA.n3355 GNDA.n1024 0.0217373
R15483 GNDA.n3355 GNDA.n1025 0.0217373
R15484 GNDA.n3365 GNDA.n989 0.0217373
R15485 GNDA.n3365 GNDA.n990 0.0217373
R15486 GNDA.n3370 GNDA.n985 0.0217373
R15487 GNDA.n3370 GNDA.n986 0.0217373
R15488 GNDA.n3375 GNDA.n981 0.0217373
R15489 GNDA.n3375 GNDA.n982 0.0217373
R15490 GNDA.n3485 GNDA.n3483 0.0217373
R15491 GNDA.n3483 GNDA.n974 0.0217373
R15492 GNDA.n3363 GNDA.n1022 0.0217373
R15493 GNDA.n3362 GNDA.n3361 0.0217373
R15494 GNDA.n3341 GNDA.n1036 0.0217373
R15495 GNDA.n1037 GNDA.n1035 0.0217373
R15496 GNDA.n3341 GNDA.n3340 0.0217373
R15497 GNDA.n597 GNDA.n513 0.0217373
R15498 GNDA.n4276 GNDA.n477 0.0217373
R15499 GNDA.n4366 GNDA.n474 0.0217373
R15500 GNDA.n472 GNDA.n471 0.0217373
R15501 GNDA.n4877 GNDA.n438 0.0217373
R15502 GNDA.n4884 GNDA.n4883 0.0217373
R15503 GNDA.n4743 GNDA.n4469 0.0217373
R15504 GNDA.n4740 GNDA.n4739 0.0217373
R15505 GNDA.n4736 GNDA.n4735 0.0217373
R15506 GNDA.n4732 GNDA.n4731 0.0217373
R15507 GNDA.n594 GNDA.n512 0.0217373
R15508 GNDA.n594 GNDA.n513 0.0217373
R15509 GNDA.n4368 GNDA.n476 0.0217373
R15510 GNDA.n4365 GNDA.n475 0.0217373
R15511 GNDA.n4367 GNDA.n4366 0.0217373
R15512 GNDA.n4370 GNDA.n473 0.0217373
R15513 GNDA.n4374 GNDA.n4373 0.0217373
R15514 GNDA.n4371 GNDA.n471 0.0217373
R15515 GNDA.n4879 GNDA.n440 0.0217373
R15516 GNDA.n4876 GNDA.n439 0.0217373
R15517 GNDA.n4878 GNDA.n4877 0.0217373
R15518 GNDA.n4277 GNDA.n4276 0.0217373
R15519 GNDA.n4745 GNDA.n4744 0.0217373
R15520 GNDA.n4749 GNDA.n4748 0.0217373
R15521 GNDA.n4746 GNDA.n4469 0.0217373
R15522 GNDA.n4554 GNDA.n4471 0.0217373
R15523 GNDA.n4555 GNDA.n4553 0.0217373
R15524 GNDA.n4741 GNDA.n4740 0.0217373
R15525 GNDA.n4559 GNDA.n4557 0.0217373
R15526 GNDA.n4560 GNDA.n4558 0.0217373
R15527 GNDA.n4737 GNDA.n4736 0.0217373
R15528 GNDA.n4728 GNDA.n4562 0.0217373
R15529 GNDA.n4729 GNDA.n4727 0.0217373
R15530 GNDA.n4733 GNDA.n4732 0.0217373
R15531 GNDA.n4886 GNDA.n436 0.0217373
R15532 GNDA.n4885 GNDA.n4884 0.0217373
R15533 GNDA.n2049 GNDA.n1893 0.0217373
R15534 GNDA.n2052 GNDA.n1889 0.0217373
R15535 GNDA.n1921 GNDA.n1891 0.0217373
R15536 GNDA.n1893 GNDA.n1892 0.0217373
R15537 GNDA.n1886 GNDA.n1885 0.0217373
R15538 GNDA.n1889 GNDA.n1885 0.0217373
R15539 GNDA.n1548 GNDA.n1547 0.0217373
R15540 GNDA.n1551 GNDA.n1458 0.0217373
R15541 GNDA.n2523 GNDA.n1553 0.0217373
R15542 GNDA.n2524 GNDA.n1554 0.0217373
R15543 GNDA.n1547 GNDA.n1464 0.0217373
R15544 GNDA.n1464 GNDA.n1458 0.0217373
R15545 GNDA.n2566 GNDA.n1423 0.0217373
R15546 GNDA.n2573 GNDA.n2571 0.0217373
R15547 GNDA.n2569 GNDA.n1417 0.0217373
R15548 GNDA.n1422 GNDA.n1420 0.0217373
R15549 GNDA.n2571 GNDA.n1418 0.0217373
R15550 GNDA.n2570 GNDA.n2569 0.0217373
R15551 GNDA.n1423 GNDA.n1421 0.0217373
R15552 GNDA.n757 GNDA.n755 0.0217373
R15553 GNDA.n3993 GNDA.n762 0.0217373
R15554 GNDA.n3991 GNDA.n771 0.0217373
R15555 GNDA.n3992 GNDA.n3991 0.0217373
R15556 GNDA.n3994 GNDA.n3993 0.0217373
R15557 GNDA.n4013 GNDA.n754 0.0217373
R15558 GNDA.n769 GNDA.n768 0.0217373
R15559 GNDA.n768 GNDA.n766 0.0217373
R15560 GNDA.n4014 GNDA.n753 0.0217373
R15561 GNDA.n4009 GNDA.n756 0.0217373
R15562 GNDA.n4010 GNDA.n4009 0.0217373
R15563 GNDA.n3863 GNDA.n932 0.0217373
R15564 GNDA.n3868 GNDA.n3867 0.0217373
R15565 GNDA.n3873 GNDA.n3872 0.0217373
R15566 GNDA.n3878 GNDA.n3877 0.0217373
R15567 GNDA.n3885 GNDA.n3884 0.0217373
R15568 GNDA.n3867 GNDA.n926 0.0217373
R15569 GNDA.n3872 GNDA.n922 0.0217373
R15570 GNDA.n3877 GNDA.n838 0.0217373
R15571 GNDA.n3884 GNDA.n3882 0.0217373
R15572 GNDA.n3864 GNDA.n931 0.0217373
R15573 GNDA.n3863 GNDA.n3862 0.0217373
R15574 GNDA.n4903 GNDA.n4902 0.0217373
R15575 GNDA.n4904 GNDA.n4901 0.0217373
R15576 GNDA.n4902 GNDA.n4900 0.0217373
R15577 GNDA.n651 GNDA.n649 0.0217373
R15578 GNDA.n4911 GNDA.n434 0.0217373
R15579 GNDA.n4887 GNDA.n434 0.0217373
R15580 GNDA.n661 GNDA.n660 0.0217373
R15581 GNDA.n4095 GNDA.n4094 0.0217373
R15582 GNDA.n4096 GNDA.n4093 0.0217373
R15583 GNDA.n4094 GNDA.n4090 0.0217373
R15584 GNDA.n4101 GNDA.n4100 0.0217373
R15585 GNDA.n613 GNDA.n611 0.0217373
R15586 GNDA.n4100 GNDA.n615 0.0217373
R15587 GNDA.n4114 GNDA.n608 0.0217373
R15588 GNDA.n4112 GNDA.n610 0.0217373
R15589 GNDA.n4108 GNDA.n612 0.0217373
R15590 GNDA.n658 GNDA.n648 0.0217373
R15591 GNDA.n655 GNDA.n650 0.0217373
R15592 GNDA.n4113 GNDA.n4112 0.0217373
R15593 GNDA.n4115 GNDA.n4114 0.0217373
R15594 GNDA.n4109 GNDA.n4108 0.0217373
R15595 GNDA.n4104 GNDA.n611 0.0217373
R15596 GNDA.n658 GNDA.n614 0.0217373
R15597 GNDA.n662 GNDA.n661 0.0217373
R15598 GNDA.n656 GNDA.n655 0.0217373
R15599 GNDA.n704 GNDA.n682 0.0217373
R15600 GNDA.n718 GNDA.n717 0.0217373
R15601 GNDA.n717 GNDA.n714 0.0217373
R15602 GNDA.n705 GNDA.n681 0.0217373
R15603 GNDA.n1013 GNDA.n999 0.0217373
R15604 GNDA.n1014 GNDA.n1012 0.0217373
R15605 GNDA.n1020 GNDA.n1019 0.0217373
R15606 GNDA.n4071 GNDA.n626 0.0217373
R15607 GNDA.n1019 GNDA.n997 0.0217373
R15608 GNDA.n628 GNDA.n626 0.0217373
R15609 GNDA.n3342 GNDA.n1037 0.0217373
R15610 GNDA.n3347 GNDA.n3346 0.0217373
R15611 GNDA.n3352 GNDA.n3351 0.0217373
R15612 GNDA.n3357 GNDA.n3356 0.0217373
R15613 GNDA.n3367 GNDA.n3366 0.0217373
R15614 GNDA.n3372 GNDA.n3371 0.0217373
R15615 GNDA.n3377 GNDA.n3376 0.0217373
R15616 GNDA.n3391 GNDA.n3390 0.0217373
R15617 GNDA.n3487 GNDA.n3486 0.0217373
R15618 GNDA.n3346 GNDA.n1031 0.0217373
R15619 GNDA.n3351 GNDA.n1027 0.0217373
R15620 GNDA.n3356 GNDA.n1023 0.0217373
R15621 GNDA.n3366 GNDA.n988 0.0217373
R15622 GNDA.n3371 GNDA.n984 0.0217373
R15623 GNDA.n3376 GNDA.n980 0.0217373
R15624 GNDA.n3390 GNDA.n976 0.0217373
R15625 GNDA.n3486 GNDA.n3484 0.0217373
R15626 GNDA.n3343 GNDA.n1036 0.0217373
R15627 GNDA.n596 GNDA.n595 0.0217373
R15628 GNDA.n595 GNDA.n511 0.0217373
R15629 GNDA.n1892 GNDA.n1890 0.0217373
R15630 GNDA.n2050 GNDA.n1891 0.0217373
R15631 GNDA.n2051 GNDA.n2050 0.0217373
R15632 GNDA.n1922 GNDA.n1890 0.0217373
R15633 GNDA.n2053 GNDA.n1887 0.0217373
R15634 GNDA.n1554 GNDA.n1552 0.0217373
R15635 GNDA.n1888 GNDA.n1887 0.0217373
R15636 GNDA.n2525 GNDA.n1553 0.0217373
R15637 GNDA.n2526 GNDA.n2525 0.0217373
R15638 GNDA.n2522 GNDA.n1552 0.0217373
R15639 GNDA.n1550 GNDA.n1549 0.0217373
R15640 GNDA.n1549 GNDA.n1465 0.0217373
R15641 GNDA.n1421 GNDA.n1419 0.0217373
R15642 GNDA.n1418 GNDA.n1416 0.0217373
R15643 GNDA.n2574 GNDA.n1417 0.0217373
R15644 GNDA.n2567 GNDA.n1420 0.0217373
R15645 GNDA.n2575 GNDA.n2574 0.0217373
R15646 GNDA.n2568 GNDA.n2567 0.0217373
R15647 GNDA.n482 GNDA.n480 0.0181756
R15648 GNDA.n482 GNDA.n478 0.0181756
R15649 GNDA.n3389 GNDA.n977 0.0181756
R15650 GNDA.n3392 GNDA.n978 0.0181756
R15651 GNDA.n3387 GNDA.n977 0.0181756
R15652 GNDA.n3387 GNDA.n978 0.0181756
R15653 GNDA.n4278 GNDA.n480 0.0181756
R15654 GNDA.n4275 GNDA.n478 0.0181756
R15655 GNDA.n3336 GNDA.n3271 0.0107812
R15656 GNDA.n3271 GNDA.n3202 0.0107812
R15657 GNDA.n3202 GNDA.n3133 0.0107812
R15658 GNDA.n3133 GNDA.n3064 0.0107812
R15659 GNDA.n3064 GNDA.n2995 0.0107812
R15660 GNDA.n2995 GNDA.n2926 0.0107812
R15661 GNDA.n2926 GNDA.n2857 0.0107812
R15662 GNDA.n2857 GNDA.n939 0.0107812
R15663 GNDA.n3536 GNDA.n939 0.0107812
R15664 GNDA.n3618 GNDA.n3536 0.0107812
R15665 GNDA.n3856 GNDA.n3618 0.0107812
R15666 GNDA.n3856 GNDA.n3791 0.0107812
R15667 GNDA.n3791 GNDA.n3722 0.0107812
R15668 GNDA.n3722 GNDA.n802 0.0107812
R15669 GNDA.n3934 GNDA.n802 0.0107812
R15670 GNDA.n3951 GNDA.n3934 0.0107812
R15671 GNDA.n3951 GNDA.n486 0.0107812
R15672 GNDA.n4195 GNDA.n486 0.0107812
R15673 GNDA.n4271 GNDA.n4195 0.0107812
R15674 GNDA.n4271 GNDA.n446 0.0107812
R15675 GNDA.n4432 GNDA.n446 0.0107812
R15676 GNDA.n4872 GNDA.n4432 0.0107812
R15677 GNDA.n4872 GNDA.n4807 0.0107812
R15678 GNDA.n4807 GNDA.n4456 0.0107812
R15679 GNDA.n4647 GNDA.n4456 0.0107812
R15680 GNDA.n4723 GNDA.n4647 0.0107812
R15681 GNDA.n2691 GNDA.n1138 0.00182188
R15682 GNDA.n2689 GNDA.n2688 0.00182188
R15683 GNDA.n2583 GNDA.n1270 0.00182188
R15684 GNDA.n2650 GNDA.n1172 0.00182188
R15685 GNDA.n2689 GNDA.n1121 0.00166081
R15686 GNDA.n2688 GNDA.n2657 0.00166081
R15687 GNDA.n1119 GNDA.n1076 0.00166081
R15688 GNDA.n2658 GNDA.n1076 0.00166081
R15689 GNDA.n1117 GNDA.n1077 0.00166081
R15690 GNDA.n2659 GNDA.n1077 0.00166081
R15691 GNDA.n1115 GNDA.n1078 0.00166081
R15692 GNDA.n2660 GNDA.n1078 0.00166081
R15693 GNDA.n1113 GNDA.n1079 0.00166081
R15694 GNDA.n2661 GNDA.n1079 0.00166081
R15695 GNDA.n1111 GNDA.n1080 0.00166081
R15696 GNDA.n2662 GNDA.n1080 0.00166081
R15697 GNDA.n1109 GNDA.n1081 0.00166081
R15698 GNDA.n2663 GNDA.n1081 0.00166081
R15699 GNDA.n1107 GNDA.n1082 0.00166081
R15700 GNDA.n2664 GNDA.n1082 0.00166081
R15701 GNDA.n1105 GNDA.n1083 0.00166081
R15702 GNDA.n2665 GNDA.n1083 0.00166081
R15703 GNDA.n1103 GNDA.n1084 0.00166081
R15704 GNDA.n2666 GNDA.n1084 0.00166081
R15705 GNDA.n1101 GNDA.n1085 0.00166081
R15706 GNDA.n2667 GNDA.n1085 0.00166081
R15707 GNDA.n1099 GNDA.n1086 0.00166081
R15708 GNDA.n2668 GNDA.n1086 0.00166081
R15709 GNDA.n1097 GNDA.n1087 0.00166081
R15710 GNDA.n2669 GNDA.n1087 0.00166081
R15711 GNDA.n1095 GNDA.n1088 0.00166081
R15712 GNDA.n2670 GNDA.n1088 0.00166081
R15713 GNDA.n1093 GNDA.n1089 0.00166081
R15714 GNDA.n2671 GNDA.n1089 0.00166081
R15715 GNDA.n1091 GNDA.n1090 0.00166081
R15716 GNDA.n1090 GNDA.n1058 0.00166081
R15717 GNDA.n1271 GNDA.n1270 0.00166081
R15718 GNDA.n1254 GNDA.n1206 0.00166081
R15719 GNDA.n1272 GNDA.n1206 0.00166081
R15720 GNDA.n1255 GNDA.n1207 0.00166081
R15721 GNDA.n1273 GNDA.n1207 0.00166081
R15722 GNDA.n1256 GNDA.n1208 0.00166081
R15723 GNDA.n1274 GNDA.n1208 0.00166081
R15724 GNDA.n1257 GNDA.n1209 0.00166081
R15725 GNDA.n1275 GNDA.n1209 0.00166081
R15726 GNDA.n1258 GNDA.n1210 0.00166081
R15727 GNDA.n1276 GNDA.n1210 0.00166081
R15728 GNDA.n1259 GNDA.n1211 0.00166081
R15729 GNDA.n1277 GNDA.n1211 0.00166081
R15730 GNDA.n1260 GNDA.n1212 0.00166081
R15731 GNDA.n1278 GNDA.n1212 0.00166081
R15732 GNDA.n1261 GNDA.n1213 0.00166081
R15733 GNDA.n1279 GNDA.n1213 0.00166081
R15734 GNDA.n1262 GNDA.n1214 0.00166081
R15735 GNDA.n1280 GNDA.n1214 0.00166081
R15736 GNDA.n1263 GNDA.n1215 0.00166081
R15737 GNDA.n1281 GNDA.n1215 0.00166081
R15738 GNDA.n1264 GNDA.n1216 0.00166081
R15739 GNDA.n1282 GNDA.n1216 0.00166081
R15740 GNDA.n1265 GNDA.n1217 0.00166081
R15741 GNDA.n1283 GNDA.n1217 0.00166081
R15742 GNDA.n1266 GNDA.n1218 0.00166081
R15743 GNDA.n1284 GNDA.n1218 0.00166081
R15744 GNDA.n1267 GNDA.n1219 0.00166081
R15745 GNDA.n1285 GNDA.n1219 0.00166081
R15746 GNDA.n1268 GNDA.n1220 0.00166081
R15747 GNDA.n1286 GNDA.n1220 0.00166081
R15748 GNDA.n1320 GNDA.n1319 0.00166081
R15749 GNDA.n2580 GNDA.n1221 0.00166081
R15750 GNDA.n1336 GNDA.n1269 0.00166081
R15751 GNDA.n1289 GNDA.n1288 0.00166081
R15752 GNDA.n1335 GNDA.n1253 0.00166081
R15753 GNDA.n1291 GNDA.n1290 0.00166081
R15754 GNDA.n1334 GNDA.n1252 0.00166081
R15755 GNDA.n1293 GNDA.n1292 0.00166081
R15756 GNDA.n1333 GNDA.n1251 0.00166081
R15757 GNDA.n1295 GNDA.n1294 0.00166081
R15758 GNDA.n1332 GNDA.n1250 0.00166081
R15759 GNDA.n1297 GNDA.n1296 0.00166081
R15760 GNDA.n1331 GNDA.n1249 0.00166081
R15761 GNDA.n1299 GNDA.n1298 0.00166081
R15762 GNDA.n1330 GNDA.n1248 0.00166081
R15763 GNDA.n1301 GNDA.n1300 0.00166081
R15764 GNDA.n1329 GNDA.n1247 0.00166081
R15765 GNDA.n1303 GNDA.n1302 0.00166081
R15766 GNDA.n1328 GNDA.n1246 0.00166081
R15767 GNDA.n1305 GNDA.n1304 0.00166081
R15768 GNDA.n1327 GNDA.n1245 0.00166081
R15769 GNDA.n1307 GNDA.n1306 0.00166081
R15770 GNDA.n1326 GNDA.n1244 0.00166081
R15771 GNDA.n1309 GNDA.n1308 0.00166081
R15772 GNDA.n1325 GNDA.n1243 0.00166081
R15773 GNDA.n1311 GNDA.n1310 0.00166081
R15774 GNDA.n1324 GNDA.n1242 0.00166081
R15775 GNDA.n1313 GNDA.n1312 0.00166081
R15776 GNDA.n1323 GNDA.n1241 0.00166081
R15777 GNDA.n1315 GNDA.n1314 0.00166081
R15778 GNDA.n1322 GNDA.n1240 0.00166081
R15779 GNDA.n1317 GNDA.n1316 0.00166081
R15780 GNDA.n1321 GNDA.n1239 0.00166081
R15781 GNDA.n2582 GNDA.n1318 0.00166081
R15782 GNDA.n2581 GNDA.n1238 0.00166081
R15783 GNDA.n2584 GNDA.n1205 0.00166081
R15784 GNDA.n2602 GNDA.n2601 0.00166081
R15785 GNDA.n2635 GNDA.n2606 0.00166081
R15786 GNDA.n2604 GNDA.n1188 0.00166081
R15787 GNDA.n2636 GNDA.n2608 0.00166081
R15788 GNDA.n2607 GNDA.n1187 0.00166081
R15789 GNDA.n2637 GNDA.n2610 0.00166081
R15790 GNDA.n2609 GNDA.n1186 0.00166081
R15791 GNDA.n2638 GNDA.n2612 0.00166081
R15792 GNDA.n2611 GNDA.n1185 0.00166081
R15793 GNDA.n2639 GNDA.n2614 0.00166081
R15794 GNDA.n2613 GNDA.n1184 0.00166081
R15795 GNDA.n2640 GNDA.n2616 0.00166081
R15796 GNDA.n2615 GNDA.n1183 0.00166081
R15797 GNDA.n2641 GNDA.n2618 0.00166081
R15798 GNDA.n2617 GNDA.n1182 0.00166081
R15799 GNDA.n2642 GNDA.n2620 0.00166081
R15800 GNDA.n2619 GNDA.n1181 0.00166081
R15801 GNDA.n2643 GNDA.n2622 0.00166081
R15802 GNDA.n2621 GNDA.n1180 0.00166081
R15803 GNDA.n2644 GNDA.n2624 0.00166081
R15804 GNDA.n2623 GNDA.n1179 0.00166081
R15805 GNDA.n2645 GNDA.n2626 0.00166081
R15806 GNDA.n2625 GNDA.n1178 0.00166081
R15807 GNDA.n2646 GNDA.n2628 0.00166081
R15808 GNDA.n2627 GNDA.n1177 0.00166081
R15809 GNDA.n2647 GNDA.n2630 0.00166081
R15810 GNDA.n2629 GNDA.n1176 0.00166081
R15811 GNDA.n2648 GNDA.n2632 0.00166081
R15812 GNDA.n2631 GNDA.n1175 0.00166081
R15813 GNDA.n2649 GNDA.n2634 0.00166081
R15814 GNDA.n2633 GNDA.n1174 0.00166081
R15815 GNDA.n2653 GNDA.n2651 0.00166081
R15816 GNDA.n2652 GNDA.n1173 0.00166081
R15817 GNDA.n2655 GNDA.n1139 0.00166081
R15818 GNDA.n2656 GNDA.n1057 0.00166081
R15819 GNDA.n2672 GNDA.n1059 0.00166081
R15820 GNDA.n1137 GNDA.n1056 0.00166081
R15821 GNDA.n2673 GNDA.n1060 0.00166081
R15822 GNDA.n1136 GNDA.n1055 0.00166081
R15823 GNDA.n2674 GNDA.n1061 0.00166081
R15824 GNDA.n1135 GNDA.n1054 0.00166081
R15825 GNDA.n2675 GNDA.n1062 0.00166081
R15826 GNDA.n1134 GNDA.n1053 0.00166081
R15827 GNDA.n2676 GNDA.n1063 0.00166081
R15828 GNDA.n1133 GNDA.n1052 0.00166081
R15829 GNDA.n2677 GNDA.n1064 0.00166081
R15830 GNDA.n1132 GNDA.n1051 0.00166081
R15831 GNDA.n2678 GNDA.n1065 0.00166081
R15832 GNDA.n1131 GNDA.n1050 0.00166081
R15833 GNDA.n2679 GNDA.n1066 0.00166081
R15834 GNDA.n1130 GNDA.n1049 0.00166081
R15835 GNDA.n2680 GNDA.n1067 0.00166081
R15836 GNDA.n1129 GNDA.n1048 0.00166081
R15837 GNDA.n2681 GNDA.n1068 0.00166081
R15838 GNDA.n1128 GNDA.n1047 0.00166081
R15839 GNDA.n2682 GNDA.n1069 0.00166081
R15840 GNDA.n1127 GNDA.n1046 0.00166081
R15841 GNDA.n2683 GNDA.n1070 0.00166081
R15842 GNDA.n1126 GNDA.n1045 0.00166081
R15843 GNDA.n2684 GNDA.n1071 0.00166081
R15844 GNDA.n1125 GNDA.n1044 0.00166081
R15845 GNDA.n2685 GNDA.n1072 0.00166081
R15846 GNDA.n1124 GNDA.n1043 0.00166081
R15847 GNDA.n2686 GNDA.n1073 0.00166081
R15848 GNDA.n1123 GNDA.n1042 0.00166081
R15849 GNDA.n2687 GNDA.n1074 0.00166081
R15850 GNDA.n1122 GNDA.n1041 0.00166081
R15851 GNDA.n2692 GNDA.n1075 0.00166081
R15852 GNDA.n1336 GNDA.n1287 0.00166081
R15853 GNDA.n1286 GNDA.n1222 0.00166081
R15854 GNDA.n1285 GNDA.n1223 0.00166081
R15855 GNDA.n1284 GNDA.n1224 0.00166081
R15856 GNDA.n1283 GNDA.n1225 0.00166081
R15857 GNDA.n1282 GNDA.n1226 0.00166081
R15858 GNDA.n1281 GNDA.n1227 0.00166081
R15859 GNDA.n1280 GNDA.n1228 0.00166081
R15860 GNDA.n1279 GNDA.n1229 0.00166081
R15861 GNDA.n1278 GNDA.n1230 0.00166081
R15862 GNDA.n1277 GNDA.n1231 0.00166081
R15863 GNDA.n1276 GNDA.n1232 0.00166081
R15864 GNDA.n1275 GNDA.n1233 0.00166081
R15865 GNDA.n1274 GNDA.n1234 0.00166081
R15866 GNDA.n1273 GNDA.n1235 0.00166081
R15867 GNDA.n1272 GNDA.n1236 0.00166081
R15868 GNDA.n1271 GNDA.n1237 0.00166081
R15869 GNDA.n1319 GNDA.n1222 0.00166081
R15870 GNDA.n1268 GNDA.n1223 0.00166081
R15871 GNDA.n1267 GNDA.n1224 0.00166081
R15872 GNDA.n1266 GNDA.n1225 0.00166081
R15873 GNDA.n1265 GNDA.n1226 0.00166081
R15874 GNDA.n1264 GNDA.n1227 0.00166081
R15875 GNDA.n1263 GNDA.n1228 0.00166081
R15876 GNDA.n1262 GNDA.n1229 0.00166081
R15877 GNDA.n1261 GNDA.n1230 0.00166081
R15878 GNDA.n1260 GNDA.n1231 0.00166081
R15879 GNDA.n1259 GNDA.n1232 0.00166081
R15880 GNDA.n1258 GNDA.n1233 0.00166081
R15881 GNDA.n1257 GNDA.n1234 0.00166081
R15882 GNDA.n1256 GNDA.n1235 0.00166081
R15883 GNDA.n1255 GNDA.n1236 0.00166081
R15884 GNDA.n1254 GNDA.n1237 0.00166081
R15885 GNDA.n1288 GNDA.n1269 0.00166081
R15886 GNDA.n1335 GNDA.n1289 0.00166081
R15887 GNDA.n1290 GNDA.n1253 0.00166081
R15888 GNDA.n1334 GNDA.n1291 0.00166081
R15889 GNDA.n1292 GNDA.n1252 0.00166081
R15890 GNDA.n1333 GNDA.n1293 0.00166081
R15891 GNDA.n1294 GNDA.n1251 0.00166081
R15892 GNDA.n1332 GNDA.n1295 0.00166081
R15893 GNDA.n1296 GNDA.n1250 0.00166081
R15894 GNDA.n1331 GNDA.n1297 0.00166081
R15895 GNDA.n1298 GNDA.n1249 0.00166081
R15896 GNDA.n1330 GNDA.n1299 0.00166081
R15897 GNDA.n1300 GNDA.n1248 0.00166081
R15898 GNDA.n1329 GNDA.n1301 0.00166081
R15899 GNDA.n1302 GNDA.n1247 0.00166081
R15900 GNDA.n1328 GNDA.n1303 0.00166081
R15901 GNDA.n1304 GNDA.n1246 0.00166081
R15902 GNDA.n1327 GNDA.n1305 0.00166081
R15903 GNDA.n1306 GNDA.n1245 0.00166081
R15904 GNDA.n1326 GNDA.n1307 0.00166081
R15905 GNDA.n1308 GNDA.n1244 0.00166081
R15906 GNDA.n1325 GNDA.n1309 0.00166081
R15907 GNDA.n1310 GNDA.n1243 0.00166081
R15908 GNDA.n1324 GNDA.n1311 0.00166081
R15909 GNDA.n1312 GNDA.n1242 0.00166081
R15910 GNDA.n1323 GNDA.n1313 0.00166081
R15911 GNDA.n1314 GNDA.n1241 0.00166081
R15912 GNDA.n1322 GNDA.n1315 0.00166081
R15913 GNDA.n1316 GNDA.n1240 0.00166081
R15914 GNDA.n1321 GNDA.n1317 0.00166081
R15915 GNDA.n1318 GNDA.n1239 0.00166081
R15916 GNDA.n2582 GNDA.n2581 0.00166081
R15917 GNDA.n1238 GNDA.n1205 0.00166081
R15918 GNDA.n1320 GNDA.n1221 0.00166081
R15919 GNDA.n2693 GNDA.n1058 0.00166081
R15920 GNDA.n2671 GNDA.n1092 0.00166081
R15921 GNDA.n2670 GNDA.n1094 0.00166081
R15922 GNDA.n2669 GNDA.n1096 0.00166081
R15923 GNDA.n2668 GNDA.n1098 0.00166081
R15924 GNDA.n2667 GNDA.n1100 0.00166081
R15925 GNDA.n2666 GNDA.n1102 0.00166081
R15926 GNDA.n2665 GNDA.n1104 0.00166081
R15927 GNDA.n2664 GNDA.n1106 0.00166081
R15928 GNDA.n2663 GNDA.n1108 0.00166081
R15929 GNDA.n2662 GNDA.n1110 0.00166081
R15930 GNDA.n2661 GNDA.n1112 0.00166081
R15931 GNDA.n2660 GNDA.n1114 0.00166081
R15932 GNDA.n2659 GNDA.n1116 0.00166081
R15933 GNDA.n2658 GNDA.n1118 0.00166081
R15934 GNDA.n2657 GNDA.n1120 0.00166081
R15935 GNDA.n2690 GNDA.n2656 0.00166081
R15936 GNDA.n1092 GNDA.n1091 0.00166081
R15937 GNDA.n1094 GNDA.n1093 0.00166081
R15938 GNDA.n1096 GNDA.n1095 0.00166081
R15939 GNDA.n1098 GNDA.n1097 0.00166081
R15940 GNDA.n1100 GNDA.n1099 0.00166081
R15941 GNDA.n1102 GNDA.n1101 0.00166081
R15942 GNDA.n1104 GNDA.n1103 0.00166081
R15943 GNDA.n1106 GNDA.n1105 0.00166081
R15944 GNDA.n1108 GNDA.n1107 0.00166081
R15945 GNDA.n1110 GNDA.n1109 0.00166081
R15946 GNDA.n1112 GNDA.n1111 0.00166081
R15947 GNDA.n1114 GNDA.n1113 0.00166081
R15948 GNDA.n1116 GNDA.n1115 0.00166081
R15949 GNDA.n1118 GNDA.n1117 0.00166081
R15950 GNDA.n1120 GNDA.n1119 0.00166081
R15951 GNDA.n2672 GNDA.n1057 0.00166081
R15952 GNDA.n1137 GNDA.n1059 0.00166081
R15953 GNDA.n2673 GNDA.n1056 0.00166081
R15954 GNDA.n1136 GNDA.n1060 0.00166081
R15955 GNDA.n2674 GNDA.n1055 0.00166081
R15956 GNDA.n1135 GNDA.n1061 0.00166081
R15957 GNDA.n2675 GNDA.n1054 0.00166081
R15958 GNDA.n1134 GNDA.n1062 0.00166081
R15959 GNDA.n2676 GNDA.n1053 0.00166081
R15960 GNDA.n1133 GNDA.n1063 0.00166081
R15961 GNDA.n2677 GNDA.n1052 0.00166081
R15962 GNDA.n1132 GNDA.n1064 0.00166081
R15963 GNDA.n2678 GNDA.n1051 0.00166081
R15964 GNDA.n1131 GNDA.n1065 0.00166081
R15965 GNDA.n2679 GNDA.n1050 0.00166081
R15966 GNDA.n1130 GNDA.n1066 0.00166081
R15967 GNDA.n2680 GNDA.n1049 0.00166081
R15968 GNDA.n1129 GNDA.n1067 0.00166081
R15969 GNDA.n2681 GNDA.n1048 0.00166081
R15970 GNDA.n1128 GNDA.n1068 0.00166081
R15971 GNDA.n2682 GNDA.n1047 0.00166081
R15972 GNDA.n1127 GNDA.n1069 0.00166081
R15973 GNDA.n2683 GNDA.n1046 0.00166081
R15974 GNDA.n1126 GNDA.n1070 0.00166081
R15975 GNDA.n2684 GNDA.n1045 0.00166081
R15976 GNDA.n1125 GNDA.n1071 0.00166081
R15977 GNDA.n2685 GNDA.n1044 0.00166081
R15978 GNDA.n1124 GNDA.n1072 0.00166081
R15979 GNDA.n2686 GNDA.n1043 0.00166081
R15980 GNDA.n1123 GNDA.n1073 0.00166081
R15981 GNDA.n2687 GNDA.n1042 0.00166081
R15982 GNDA.n1122 GNDA.n1074 0.00166081
R15983 GNDA.n1075 GNDA.n1041 0.00166081
R15984 GNDA.n1138 GNDA.n1121 0.00166081
R15985 GNDA.n2654 GNDA.n2603 0.00166081
R15986 GNDA.n2585 GNDA.n1172 0.00166081
R15987 GNDA.n1189 GNDA.n1140 0.00166081
R15988 GNDA.n2586 GNDA.n1171 0.00166081
R15989 GNDA.n1190 GNDA.n1141 0.00166081
R15990 GNDA.n2587 GNDA.n1170 0.00166081
R15991 GNDA.n1191 GNDA.n1142 0.00166081
R15992 GNDA.n2588 GNDA.n1169 0.00166081
R15993 GNDA.n1192 GNDA.n1143 0.00166081
R15994 GNDA.n2589 GNDA.n1168 0.00166081
R15995 GNDA.n1193 GNDA.n1144 0.00166081
R15996 GNDA.n2590 GNDA.n1167 0.00166081
R15997 GNDA.n1194 GNDA.n1145 0.00166081
R15998 GNDA.n2591 GNDA.n1166 0.00166081
R15999 GNDA.n1195 GNDA.n1146 0.00166081
R16000 GNDA.n2592 GNDA.n1165 0.00166081
R16001 GNDA.n1196 GNDA.n1147 0.00166081
R16002 GNDA.n2593 GNDA.n1164 0.00166081
R16003 GNDA.n1197 GNDA.n1148 0.00166081
R16004 GNDA.n2594 GNDA.n1163 0.00166081
R16005 GNDA.n1198 GNDA.n1149 0.00166081
R16006 GNDA.n2595 GNDA.n1162 0.00166081
R16007 GNDA.n1199 GNDA.n1150 0.00166081
R16008 GNDA.n2596 GNDA.n1161 0.00166081
R16009 GNDA.n1200 GNDA.n1151 0.00166081
R16010 GNDA.n2597 GNDA.n1160 0.00166081
R16011 GNDA.n1201 GNDA.n1152 0.00166081
R16012 GNDA.n2598 GNDA.n1159 0.00166081
R16013 GNDA.n1202 GNDA.n1153 0.00166081
R16014 GNDA.n2599 GNDA.n1158 0.00166081
R16015 GNDA.n1203 GNDA.n1154 0.00166081
R16016 GNDA.n2600 GNDA.n1157 0.00166081
R16017 GNDA.n2605 GNDA.n1155 0.00166081
R16018 GNDA.n2600 GNDA.n1155 0.00166081
R16019 GNDA.n2599 GNDA.n1154 0.00166081
R16020 GNDA.n2598 GNDA.n1153 0.00166081
R16021 GNDA.n2597 GNDA.n1152 0.00166081
R16022 GNDA.n2596 GNDA.n1151 0.00166081
R16023 GNDA.n2595 GNDA.n1150 0.00166081
R16024 GNDA.n2594 GNDA.n1149 0.00166081
R16025 GNDA.n2593 GNDA.n1148 0.00166081
R16026 GNDA.n2592 GNDA.n1147 0.00166081
R16027 GNDA.n2591 GNDA.n1146 0.00166081
R16028 GNDA.n2590 GNDA.n1145 0.00166081
R16029 GNDA.n2589 GNDA.n1144 0.00166081
R16030 GNDA.n2588 GNDA.n1143 0.00166081
R16031 GNDA.n2587 GNDA.n1142 0.00166081
R16032 GNDA.n2586 GNDA.n1141 0.00166081
R16033 GNDA.n2585 GNDA.n1140 0.00166081
R16034 GNDA.n2650 GNDA.n2603 0.00166081
R16035 GNDA.n2601 GNDA.n1204 0.00166081
R16036 GNDA.n1203 GNDA.n1157 0.00166081
R16037 GNDA.n1202 GNDA.n1158 0.00166081
R16038 GNDA.n1201 GNDA.n1159 0.00166081
R16039 GNDA.n1200 GNDA.n1160 0.00166081
R16040 GNDA.n1199 GNDA.n1161 0.00166081
R16041 GNDA.n1198 GNDA.n1162 0.00166081
R16042 GNDA.n1197 GNDA.n1163 0.00166081
R16043 GNDA.n1196 GNDA.n1164 0.00166081
R16044 GNDA.n1195 GNDA.n1165 0.00166081
R16045 GNDA.n1194 GNDA.n1166 0.00166081
R16046 GNDA.n1193 GNDA.n1167 0.00166081
R16047 GNDA.n1192 GNDA.n1168 0.00166081
R16048 GNDA.n1191 GNDA.n1169 0.00166081
R16049 GNDA.n1190 GNDA.n1170 0.00166081
R16050 GNDA.n1189 GNDA.n1171 0.00166081
R16051 GNDA.n2635 GNDA.n1204 0.00166081
R16052 GNDA.n2605 GNDA.n1156 0.00166081
R16053 GNDA.n2606 GNDA.n2604 0.00166081
R16054 GNDA.n2636 GNDA.n1188 0.00166081
R16055 GNDA.n2608 GNDA.n2607 0.00166081
R16056 GNDA.n2637 GNDA.n1187 0.00166081
R16057 GNDA.n2610 GNDA.n2609 0.00166081
R16058 GNDA.n2638 GNDA.n1186 0.00166081
R16059 GNDA.n2612 GNDA.n2611 0.00166081
R16060 GNDA.n2639 GNDA.n1185 0.00166081
R16061 GNDA.n2614 GNDA.n2613 0.00166081
R16062 GNDA.n2640 GNDA.n1184 0.00166081
R16063 GNDA.n2616 GNDA.n2615 0.00166081
R16064 GNDA.n2641 GNDA.n1183 0.00166081
R16065 GNDA.n2618 GNDA.n2617 0.00166081
R16066 GNDA.n2642 GNDA.n1182 0.00166081
R16067 GNDA.n2620 GNDA.n2619 0.00166081
R16068 GNDA.n2643 GNDA.n1181 0.00166081
R16069 GNDA.n2622 GNDA.n2621 0.00166081
R16070 GNDA.n2644 GNDA.n1180 0.00166081
R16071 GNDA.n2624 GNDA.n2623 0.00166081
R16072 GNDA.n2645 GNDA.n1179 0.00166081
R16073 GNDA.n2626 GNDA.n2625 0.00166081
R16074 GNDA.n2646 GNDA.n1178 0.00166081
R16075 GNDA.n2628 GNDA.n2627 0.00166081
R16076 GNDA.n2647 GNDA.n1177 0.00166081
R16077 GNDA.n2630 GNDA.n2629 0.00166081
R16078 GNDA.n2648 GNDA.n1176 0.00166081
R16079 GNDA.n2632 GNDA.n2631 0.00166081
R16080 GNDA.n2649 GNDA.n1175 0.00166081
R16081 GNDA.n2634 GNDA.n2633 0.00166081
R16082 GNDA.n2651 GNDA.n1174 0.00166081
R16083 GNDA.n2653 GNDA.n2652 0.00166081
R16084 GNDA.n1173 GNDA.n1139 0.00166081
R16085 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n7 301.983
R16086 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n9 297.151
R16087 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n6 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n5 297.151
R16088 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n27 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n26 118.861
R16089 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n29 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n28 118.861
R16090 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n33 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n32 118.861
R16091 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n35 118.861
R16092 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n39 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n38 118.861
R16093 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n41 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t0 115.672
R16094 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t5 39.4005
R16095 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t2 39.4005
R16096 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t4 39.4005
R16097 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t3 39.4005
R16098 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t1 39.4005
R16099 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t6 39.4005
R16100 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n26 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t10 19.7005
R16101 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n26 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t15 19.7005
R16102 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n28 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t11 19.7005
R16103 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n28 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t16 19.7005
R16104 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n32 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t13 19.7005
R16105 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n32 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t7 19.7005
R16106 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n35 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t12 19.7005
R16107 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n35 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t9 19.7005
R16108 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n38 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t14 19.7005
R16109 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n38 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t8 19.7005
R16110 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n6 11.9588
R16111 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n11 11.6211
R16112 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 9.92238
R16113 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n30 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n27 5.60467
R16114 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n39 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n37 5.54217
R16115 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n27 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n25 5.54217
R16116 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n6 5.39633
R16117 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n10 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n8 5.39633
R16118 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n30 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n29 5.04217
R16119 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n33 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n31 5.04217
R16120 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n24 5.04217
R16121 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n40 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n39 5.04217
R16122 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n29 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n25 4.97967
R16123 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n34 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n33 4.97967
R16124 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n37 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n36 4.97967
R16125 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n4 4.5005
R16126 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n15 4.5005
R16127 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n14 4.5005
R16128 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n20 4.5005
R16129 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n41 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n40 2.99085
R16130 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n0 2.26187
R16131 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n18 2.26187
R16132 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n2 2.24063
R16133 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n1 2.24063
R16134 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n17 2.24063
R16135 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n23 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n0 2.24063
R16136 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n12 2.24063
R16137 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n10 1.34946
R16138 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n37 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n34 0.563
R16139 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n34 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n25 0.563
R16140 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n23 0.443208
R16141 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n40 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n24 0.34425
R16142 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n31 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n24 0.34425
R16143 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n31 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n30 0.34425
R16144 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n16 0.078625
R16145 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n1 0.0421667
R16146 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n2 0.0217373
R16147 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n3 0.0217373
R16148 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n2 0.0217373
R16149 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n4 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n3 0.0217373
R16150 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n22 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n21 0.0217373
R16151 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n0 0.0217373
R16152 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n23 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n22 0.0217373
R16153 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n14 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n13 0.0217373
R16154 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n19 0.0217373
R16155 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n1 0.0217373
R16156 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n21 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n18 0.0217373
R16157 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n17 0.0217373
R16158 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n41 0.0213333
R16159 two_stage_opamp_dummy_magic_29_0.Y.n53 two_stage_opamp_dummy_magic_29_0.Y.t38 1172.87
R16160 two_stage_opamp_dummy_magic_29_0.Y.n49 two_stage_opamp_dummy_magic_29_0.Y.t29 1172.87
R16161 two_stage_opamp_dummy_magic_29_0.Y.n53 two_stage_opamp_dummy_magic_29_0.Y.t30 996.134
R16162 two_stage_opamp_dummy_magic_29_0.Y.n54 two_stage_opamp_dummy_magic_29_0.Y.t44 996.134
R16163 two_stage_opamp_dummy_magic_29_0.Y.n55 two_stage_opamp_dummy_magic_29_0.Y.t32 996.134
R16164 two_stage_opamp_dummy_magic_29_0.Y.n56 two_stage_opamp_dummy_magic_29_0.Y.t46 996.134
R16165 two_stage_opamp_dummy_magic_29_0.Y.n52 two_stage_opamp_dummy_magic_29_0.Y.t35 996.134
R16166 two_stage_opamp_dummy_magic_29_0.Y.n51 two_stage_opamp_dummy_magic_29_0.Y.t42 996.134
R16167 two_stage_opamp_dummy_magic_29_0.Y.n50 two_stage_opamp_dummy_magic_29_0.Y.t27 996.134
R16168 two_stage_opamp_dummy_magic_29_0.Y.n49 two_stage_opamp_dummy_magic_29_0.Y.t43 996.134
R16169 two_stage_opamp_dummy_magic_29_0.Y.n71 two_stage_opamp_dummy_magic_29_0.Y.t25 690.867
R16170 two_stage_opamp_dummy_magic_29_0.Y.n64 two_stage_opamp_dummy_magic_29_0.Y.t48 690.867
R16171 two_stage_opamp_dummy_magic_29_0.Y.n80 two_stage_opamp_dummy_magic_29_0.Y.t28 530.201
R16172 two_stage_opamp_dummy_magic_29_0.Y.n73 two_stage_opamp_dummy_magic_29_0.Y.t50 530.201
R16173 two_stage_opamp_dummy_magic_29_0.Y.n71 two_stage_opamp_dummy_magic_29_0.Y.t49 514.134
R16174 two_stage_opamp_dummy_magic_29_0.Y.n64 two_stage_opamp_dummy_magic_29_0.Y.t34 514.134
R16175 two_stage_opamp_dummy_magic_29_0.Y.n65 two_stage_opamp_dummy_magic_29_0.Y.t45 514.134
R16176 two_stage_opamp_dummy_magic_29_0.Y.n66 two_stage_opamp_dummy_magic_29_0.Y.t31 514.134
R16177 two_stage_opamp_dummy_magic_29_0.Y.n67 two_stage_opamp_dummy_magic_29_0.Y.t54 514.134
R16178 two_stage_opamp_dummy_magic_29_0.Y.n68 two_stage_opamp_dummy_magic_29_0.Y.t40 514.134
R16179 two_stage_opamp_dummy_magic_29_0.Y.n69 two_stage_opamp_dummy_magic_29_0.Y.t52 514.134
R16180 two_stage_opamp_dummy_magic_29_0.Y.n70 two_stage_opamp_dummy_magic_29_0.Y.t37 514.134
R16181 two_stage_opamp_dummy_magic_29_0.Y.n80 two_stage_opamp_dummy_magic_29_0.Y.t51 353.467
R16182 two_stage_opamp_dummy_magic_29_0.Y.n79 two_stage_opamp_dummy_magic_29_0.Y.t39 353.467
R16183 two_stage_opamp_dummy_magic_29_0.Y.n78 two_stage_opamp_dummy_magic_29_0.Y.t53 353.467
R16184 two_stage_opamp_dummy_magic_29_0.Y.n77 two_stage_opamp_dummy_magic_29_0.Y.t41 353.467
R16185 two_stage_opamp_dummy_magic_29_0.Y.n76 two_stage_opamp_dummy_magic_29_0.Y.t26 353.467
R16186 two_stage_opamp_dummy_magic_29_0.Y.n75 two_stage_opamp_dummy_magic_29_0.Y.t33 353.467
R16187 two_stage_opamp_dummy_magic_29_0.Y.n74 two_stage_opamp_dummy_magic_29_0.Y.t47 353.467
R16188 two_stage_opamp_dummy_magic_29_0.Y.n73 two_stage_opamp_dummy_magic_29_0.Y.t36 353.467
R16189 two_stage_opamp_dummy_magic_29_0.Y.n52 two_stage_opamp_dummy_magic_29_0.Y.n51 176.733
R16190 two_stage_opamp_dummy_magic_29_0.Y.n51 two_stage_opamp_dummy_magic_29_0.Y.n50 176.733
R16191 two_stage_opamp_dummy_magic_29_0.Y.n50 two_stage_opamp_dummy_magic_29_0.Y.n49 176.733
R16192 two_stage_opamp_dummy_magic_29_0.Y.n54 two_stage_opamp_dummy_magic_29_0.Y.n53 176.733
R16193 two_stage_opamp_dummy_magic_29_0.Y.n55 two_stage_opamp_dummy_magic_29_0.Y.n54 176.733
R16194 two_stage_opamp_dummy_magic_29_0.Y.n56 two_stage_opamp_dummy_magic_29_0.Y.n55 176.733
R16195 two_stage_opamp_dummy_magic_29_0.Y.n79 two_stage_opamp_dummy_magic_29_0.Y.n78 176.733
R16196 two_stage_opamp_dummy_magic_29_0.Y.n78 two_stage_opamp_dummy_magic_29_0.Y.n77 176.733
R16197 two_stage_opamp_dummy_magic_29_0.Y.n77 two_stage_opamp_dummy_magic_29_0.Y.n76 176.733
R16198 two_stage_opamp_dummy_magic_29_0.Y.n76 two_stage_opamp_dummy_magic_29_0.Y.n75 176.733
R16199 two_stage_opamp_dummy_magic_29_0.Y.n75 two_stage_opamp_dummy_magic_29_0.Y.n74 176.733
R16200 two_stage_opamp_dummy_magic_29_0.Y.n74 two_stage_opamp_dummy_magic_29_0.Y.n73 176.733
R16201 two_stage_opamp_dummy_magic_29_0.Y.n70 two_stage_opamp_dummy_magic_29_0.Y.n69 176.733
R16202 two_stage_opamp_dummy_magic_29_0.Y.n69 two_stage_opamp_dummy_magic_29_0.Y.n68 176.733
R16203 two_stage_opamp_dummy_magic_29_0.Y.n68 two_stage_opamp_dummy_magic_29_0.Y.n67 176.733
R16204 two_stage_opamp_dummy_magic_29_0.Y.n67 two_stage_opamp_dummy_magic_29_0.Y.n66 176.733
R16205 two_stage_opamp_dummy_magic_29_0.Y.n66 two_stage_opamp_dummy_magic_29_0.Y.n65 176.733
R16206 two_stage_opamp_dummy_magic_29_0.Y.n65 two_stage_opamp_dummy_magic_29_0.Y.n64 176.733
R16207 two_stage_opamp_dummy_magic_29_0.Y.n82 two_stage_opamp_dummy_magic_29_0.Y.n81 165.472
R16208 two_stage_opamp_dummy_magic_29_0.Y.n82 two_stage_opamp_dummy_magic_29_0.Y.n72 165.472
R16209 two_stage_opamp_dummy_magic_29_0.Y.n59 two_stage_opamp_dummy_magic_29_0.Y.n58 152
R16210 two_stage_opamp_dummy_magic_29_0.Y.n60 two_stage_opamp_dummy_magic_29_0.Y.n59 131.571
R16211 two_stage_opamp_dummy_magic_29_0.Y.n59 two_stage_opamp_dummy_magic_29_0.Y.n57 124.517
R16212 two_stage_opamp_dummy_magic_29_0.Y.n84 two_stage_opamp_dummy_magic_29_0.Y.n82 74.5372
R16213 two_stage_opamp_dummy_magic_29_0.Y.n110 two_stage_opamp_dummy_magic_29_0.Y.n109 66.0338
R16214 two_stage_opamp_dummy_magic_29_0.Y.n94 two_stage_opamp_dummy_magic_29_0.Y.n93 66.0338
R16215 two_stage_opamp_dummy_magic_29_0.Y.n97 two_stage_opamp_dummy_magic_29_0.Y.n96 66.0338
R16216 two_stage_opamp_dummy_magic_29_0.Y.n100 two_stage_opamp_dummy_magic_29_0.Y.n99 66.0338
R16217 two_stage_opamp_dummy_magic_29_0.Y.n104 two_stage_opamp_dummy_magic_29_0.Y.n103 66.0338
R16218 two_stage_opamp_dummy_magic_29_0.Y.n107 two_stage_opamp_dummy_magic_29_0.Y.n106 66.0338
R16219 two_stage_opamp_dummy_magic_29_0.Y.n8 two_stage_opamp_dummy_magic_29_0.Y.n6 54.7984
R16220 two_stage_opamp_dummy_magic_29_0.Y.n8 two_stage_opamp_dummy_magic_29_0.Y.n7 54.4547
R16221 two_stage_opamp_dummy_magic_29_0.Y.n10 two_stage_opamp_dummy_magic_29_0.Y.n9 54.4547
R16222 two_stage_opamp_dummy_magic_29_0.Y.n12 two_stage_opamp_dummy_magic_29_0.Y.n11 54.4547
R16223 two_stage_opamp_dummy_magic_29_0.Y.n14 two_stage_opamp_dummy_magic_29_0.Y.n13 54.4547
R16224 two_stage_opamp_dummy_magic_29_0.Y.n16 two_stage_opamp_dummy_magic_29_0.Y.n15 54.4547
R16225 two_stage_opamp_dummy_magic_29_0.Y.n43 two_stage_opamp_dummy_magic_29_0.Y.t0 41.0384
R16226 two_stage_opamp_dummy_magic_29_0.Y.n57 two_stage_opamp_dummy_magic_29_0.Y.n52 40.1672
R16227 two_stage_opamp_dummy_magic_29_0.Y.n57 two_stage_opamp_dummy_magic_29_0.Y.n56 40.1672
R16228 two_stage_opamp_dummy_magic_29_0.Y.n81 two_stage_opamp_dummy_magic_29_0.Y.n79 40.1672
R16229 two_stage_opamp_dummy_magic_29_0.Y.n81 two_stage_opamp_dummy_magic_29_0.Y.n80 40.1672
R16230 two_stage_opamp_dummy_magic_29_0.Y.n72 two_stage_opamp_dummy_magic_29_0.Y.n70 40.1672
R16231 two_stage_opamp_dummy_magic_29_0.Y.n72 two_stage_opamp_dummy_magic_29_0.Y.n71 40.1672
R16232 two_stage_opamp_dummy_magic_29_0.Y.n61 two_stage_opamp_dummy_magic_29_0.Y.n60 16.3217
R16233 two_stage_opamp_dummy_magic_29_0.Y.n6 two_stage_opamp_dummy_magic_29_0.Y.t15 16.0005
R16234 two_stage_opamp_dummy_magic_29_0.Y.n6 two_stage_opamp_dummy_magic_29_0.Y.t23 16.0005
R16235 two_stage_opamp_dummy_magic_29_0.Y.n7 two_stage_opamp_dummy_magic_29_0.Y.t16 16.0005
R16236 two_stage_opamp_dummy_magic_29_0.Y.n7 two_stage_opamp_dummy_magic_29_0.Y.t13 16.0005
R16237 two_stage_opamp_dummy_magic_29_0.Y.n9 two_stage_opamp_dummy_magic_29_0.Y.t4 16.0005
R16238 two_stage_opamp_dummy_magic_29_0.Y.n9 two_stage_opamp_dummy_magic_29_0.Y.t14 16.0005
R16239 two_stage_opamp_dummy_magic_29_0.Y.n11 two_stage_opamp_dummy_magic_29_0.Y.t11 16.0005
R16240 two_stage_opamp_dummy_magic_29_0.Y.n11 two_stage_opamp_dummy_magic_29_0.Y.t5 16.0005
R16241 two_stage_opamp_dummy_magic_29_0.Y.n13 two_stage_opamp_dummy_magic_29_0.Y.t12 16.0005
R16242 two_stage_opamp_dummy_magic_29_0.Y.n13 two_stage_opamp_dummy_magic_29_0.Y.t8 16.0005
R16243 two_stage_opamp_dummy_magic_29_0.Y.n15 two_stage_opamp_dummy_magic_29_0.Y.t22 16.0005
R16244 two_stage_opamp_dummy_magic_29_0.Y.n15 two_stage_opamp_dummy_magic_29_0.Y.t24 16.0005
R16245 two_stage_opamp_dummy_magic_29_0.Y.n58 two_stage_opamp_dummy_magic_29_0.Y.n48 12.8005
R16246 two_stage_opamp_dummy_magic_29_0.Y.n109 two_stage_opamp_dummy_magic_29_0.Y.t21 11.2576
R16247 two_stage_opamp_dummy_magic_29_0.Y.n109 two_stage_opamp_dummy_magic_29_0.Y.t2 11.2576
R16248 two_stage_opamp_dummy_magic_29_0.Y.n93 two_stage_opamp_dummy_magic_29_0.Y.t19 11.2576
R16249 two_stage_opamp_dummy_magic_29_0.Y.n93 two_stage_opamp_dummy_magic_29_0.Y.t20 11.2576
R16250 two_stage_opamp_dummy_magic_29_0.Y.n96 two_stage_opamp_dummy_magic_29_0.Y.t18 11.2576
R16251 two_stage_opamp_dummy_magic_29_0.Y.n96 two_stage_opamp_dummy_magic_29_0.Y.t6 11.2576
R16252 two_stage_opamp_dummy_magic_29_0.Y.n99 two_stage_opamp_dummy_magic_29_0.Y.t9 11.2576
R16253 two_stage_opamp_dummy_magic_29_0.Y.n99 two_stage_opamp_dummy_magic_29_0.Y.t17 11.2576
R16254 two_stage_opamp_dummy_magic_29_0.Y.n103 two_stage_opamp_dummy_magic_29_0.Y.t1 11.2576
R16255 two_stage_opamp_dummy_magic_29_0.Y.n103 two_stage_opamp_dummy_magic_29_0.Y.t3 11.2576
R16256 two_stage_opamp_dummy_magic_29_0.Y.n106 two_stage_opamp_dummy_magic_29_0.Y.t10 11.2576
R16257 two_stage_opamp_dummy_magic_29_0.Y.n106 two_stage_opamp_dummy_magic_29_0.Y.t7 11.2576
R16258 two_stage_opamp_dummy_magic_29_0.Y.n17 two_stage_opamp_dummy_magic_29_0.Y.n16 11.1099
R16259 two_stage_opamp_dummy_magic_29_0.Y.n58 two_stage_opamp_dummy_magic_29_0.Y.n46 9.36264
R16260 two_stage_opamp_dummy_magic_29_0.Y.n48 two_stage_opamp_dummy_magic_29_0.Y.n47 9.3005
R16261 two_stage_opamp_dummy_magic_29_0.Y.n119 two_stage_opamp_dummy_magic_29_0.Y.n25 5.78175
R16262 two_stage_opamp_dummy_magic_29_0.Y.n98 two_stage_opamp_dummy_magic_29_0.Y.n94 5.66717
R16263 two_stage_opamp_dummy_magic_29_0.Y.n95 two_stage_opamp_dummy_magic_29_0.Y.n94 5.66717
R16264 two_stage_opamp_dummy_magic_29_0.Y.n110 two_stage_opamp_dummy_magic_29_0.Y.n108 5.66717
R16265 two_stage_opamp_dummy_magic_29_0.Y.n18 two_stage_opamp_dummy_magic_29_0.Y.n17 5.46373
R16266 two_stage_opamp_dummy_magic_29_0.Y.n19 two_stage_opamp_dummy_magic_29_0.Y.n5 5.438
R16267 two_stage_opamp_dummy_magic_29_0.Y.n21 two_stage_opamp_dummy_magic_29_0.Y.n4 5.438
R16268 two_stage_opamp_dummy_magic_29_0.Y.n125 two_stage_opamp_dummy_magic_29_0.Y.n1 5.438
R16269 two_stage_opamp_dummy_magic_29_0.Y.n121 two_stage_opamp_dummy_magic_29_0.Y.n25 5.438
R16270 two_stage_opamp_dummy_magic_29_0.Y.n60 two_stage_opamp_dummy_magic_29_0.Y.n48 5.33141
R16271 two_stage_opamp_dummy_magic_29_0.Y.n98 two_stage_opamp_dummy_magic_29_0.Y.n97 5.29217
R16272 two_stage_opamp_dummy_magic_29_0.Y.n97 two_stage_opamp_dummy_magic_29_0.Y.n95 5.29217
R16273 two_stage_opamp_dummy_magic_29_0.Y.n101 two_stage_opamp_dummy_magic_29_0.Y.n100 5.29217
R16274 two_stage_opamp_dummy_magic_29_0.Y.n100 two_stage_opamp_dummy_magic_29_0.Y.n92 5.29217
R16275 two_stage_opamp_dummy_magic_29_0.Y.n104 two_stage_opamp_dummy_magic_29_0.Y.n102 5.29217
R16276 two_stage_opamp_dummy_magic_29_0.Y.n105 two_stage_opamp_dummy_magic_29_0.Y.n104 5.29217
R16277 two_stage_opamp_dummy_magic_29_0.Y.n107 two_stage_opamp_dummy_magic_29_0.Y.n91 5.29217
R16278 two_stage_opamp_dummy_magic_29_0.Y.n108 two_stage_opamp_dummy_magic_29_0.Y.n107 5.29217
R16279 two_stage_opamp_dummy_magic_29_0.Y.n111 two_stage_opamp_dummy_magic_29_0.Y.n110 5.29217
R16280 two_stage_opamp_dummy_magic_29_0.Y.n117 two_stage_opamp_dummy_magic_29_0.Y.n28 4.5005
R16281 two_stage_opamp_dummy_magic_29_0.Y.n117 two_stage_opamp_dummy_magic_29_0.Y.n30 4.5005
R16282 two_stage_opamp_dummy_magic_29_0.Y.n117 two_stage_opamp_dummy_magic_29_0.Y.n27 4.5005
R16283 two_stage_opamp_dummy_magic_29_0.Y.n117 two_stage_opamp_dummy_magic_29_0.Y.n116 4.5005
R16284 two_stage_opamp_dummy_magic_29_0.Y.n34 two_stage_opamp_dummy_magic_29_0.Y.n32 4.5005
R16285 two_stage_opamp_dummy_magic_29_0.Y.n83 two_stage_opamp_dummy_magic_29_0.Y.n36 4.5005
R16286 two_stage_opamp_dummy_magic_29_0.Y.n85 two_stage_opamp_dummy_magic_29_0.Y.n84 4.5005
R16287 two_stage_opamp_dummy_magic_29_0.Y.n84 two_stage_opamp_dummy_magic_29_0.Y.n83 4.5005
R16288 two_stage_opamp_dummy_magic_29_0.Y.n62 two_stage_opamp_dummy_magic_29_0.Y.n61 4.5005
R16289 two_stage_opamp_dummy_magic_29_0.Y.n40 two_stage_opamp_dummy_magic_29_0.Y.n39 4.5005
R16290 two_stage_opamp_dummy_magic_29_0.Y.n112 two_stage_opamp_dummy_magic_29_0.Y.n111 2.35543
R16291 two_stage_opamp_dummy_magic_29_0.Y.n41 two_stage_opamp_dummy_magic_29_0.Y.n38 2.26187
R16292 two_stage_opamp_dummy_magic_29_0.Y.n42 two_stage_opamp_dummy_magic_29_0.Y.n41 2.26187
R16293 two_stage_opamp_dummy_magic_29_0.Y.n112 two_stage_opamp_dummy_magic_29_0.Y.n29 2.24654
R16294 two_stage_opamp_dummy_magic_29_0.Y.n89 two_stage_opamp_dummy_magic_29_0.Y.n88 2.24654
R16295 two_stage_opamp_dummy_magic_29_0.Y.n34 two_stage_opamp_dummy_magic_29_0.Y.n33 2.24063
R16296 two_stage_opamp_dummy_magic_29_0.Y.n34 two_stage_opamp_dummy_magic_29_0.Y.n31 2.24063
R16297 two_stage_opamp_dummy_magic_29_0.Y.n117 two_stage_opamp_dummy_magic_29_0.Y.n26 2.24063
R16298 two_stage_opamp_dummy_magic_29_0.Y.n86 two_stage_opamp_dummy_magic_29_0.Y.n85 2.24063
R16299 two_stage_opamp_dummy_magic_29_0.Y.n63 two_stage_opamp_dummy_magic_29_0.Y.n37 2.24063
R16300 two_stage_opamp_dummy_magic_29_0.Y.n45 two_stage_opamp_dummy_magic_29_0.Y.n38 2.24063
R16301 two_stage_opamp_dummy_magic_29_0.Y.n114 two_stage_opamp_dummy_magic_29_0.Y.n113 2.24063
R16302 two_stage_opamp_dummy_magic_29_0.Y.n114 two_stage_opamp_dummy_magic_29_0.Y.n90 2.24063
R16303 two_stage_opamp_dummy_magic_29_0.Y.n115 two_stage_opamp_dummy_magic_29_0.Y.n114 2.24063
R16304 two_stage_opamp_dummy_magic_29_0.Y.n87 two_stage_opamp_dummy_magic_29_0.Y.n35 2.24063
R16305 two_stage_opamp_dummy_magic_29_0.Y.n44 two_stage_opamp_dummy_magic_29_0.Y.n43 2.24063
R16306 two_stage_opamp_dummy_magic_29_0.Y.n62 two_stage_opamp_dummy_magic_29_0.Y.n46 2.22018
R16307 two_stage_opamp_dummy_magic_29_0.Y.n62 two_stage_opamp_dummy_magic_29_0.Y.n45 0.682792
R16308 two_stage_opamp_dummy_magic_29_0.Y.n119 two_stage_opamp_dummy_magic_29_0.Y.n118 0.643357
R16309 two_stage_opamp_dummy_magic_29_0.Y.n120 two_stage_opamp_dummy_magic_29_0.Y.n24 0.643357
R16310 two_stage_opamp_dummy_magic_29_0.Y.n122 two_stage_opamp_dummy_magic_29_0.Y.n121 0.643357
R16311 two_stage_opamp_dummy_magic_29_0.Y.n123 two_stage_opamp_dummy_magic_29_0.Y.n2 0.643357
R16312 two_stage_opamp_dummy_magic_29_0.Y.n125 two_stage_opamp_dummy_magic_29_0.Y.n124 0.643357
R16313 two_stage_opamp_dummy_magic_29_0.Y.n23 two_stage_opamp_dummy_magic_29_0.Y.n0 0.643357
R16314 two_stage_opamp_dummy_magic_29_0.Y.n22 two_stage_opamp_dummy_magic_29_0.Y.n21 0.643357
R16315 two_stage_opamp_dummy_magic_29_0.Y.n20 two_stage_opamp_dummy_magic_29_0.Y.n3 0.643357
R16316 two_stage_opamp_dummy_magic_29_0.Y.n88 two_stage_opamp_dummy_magic_29_0.Y.n87 0.479667
R16317 two_stage_opamp_dummy_magic_29_0.Y.n85 two_stage_opamp_dummy_magic_29_0.Y.n62 0.46925
R16318 two_stage_opamp_dummy_magic_29_0.Y.n108 two_stage_opamp_dummy_magic_29_0.Y.n105 0.3755
R16319 two_stage_opamp_dummy_magic_29_0.Y.n105 two_stage_opamp_dummy_magic_29_0.Y.n92 0.3755
R16320 two_stage_opamp_dummy_magic_29_0.Y.n95 two_stage_opamp_dummy_magic_29_0.Y.n92 0.3755
R16321 two_stage_opamp_dummy_magic_29_0.Y.n111 two_stage_opamp_dummy_magic_29_0.Y.n91 0.3755
R16322 two_stage_opamp_dummy_magic_29_0.Y.n102 two_stage_opamp_dummy_magic_29_0.Y.n91 0.3755
R16323 two_stage_opamp_dummy_magic_29_0.Y.n102 two_stage_opamp_dummy_magic_29_0.Y.n101 0.3755
R16324 two_stage_opamp_dummy_magic_29_0.Y.n101 two_stage_opamp_dummy_magic_29_0.Y.n98 0.3755
R16325 two_stage_opamp_dummy_magic_29_0.Y.n16 two_stage_opamp_dummy_magic_29_0.Y.n14 0.34425
R16326 two_stage_opamp_dummy_magic_29_0.Y.n14 two_stage_opamp_dummy_magic_29_0.Y.n12 0.34425
R16327 two_stage_opamp_dummy_magic_29_0.Y.n12 two_stage_opamp_dummy_magic_29_0.Y.n10 0.34425
R16328 two_stage_opamp_dummy_magic_29_0.Y.n10 two_stage_opamp_dummy_magic_29_0.Y.n8 0.34425
R16329 two_stage_opamp_dummy_magic_29_0.Y.n17 two_stage_opamp_dummy_magic_29_0.Y.n5 0.34425
R16330 two_stage_opamp_dummy_magic_29_0.Y.n5 two_stage_opamp_dummy_magic_29_0.Y.n4 0.34425
R16331 two_stage_opamp_dummy_magic_29_0.Y.n4 two_stage_opamp_dummy_magic_29_0.Y.n1 0.34425
R16332 two_stage_opamp_dummy_magic_29_0.Y.n25 two_stage_opamp_dummy_magic_29_0.Y.n1 0.34425
R16333 two_stage_opamp_dummy_magic_29_0.Y.n118 two_stage_opamp_dummy_magic_29_0.Y.n117 0.270589
R16334 two_stage_opamp_dummy_magic_29_0.Y.n18 two_stage_opamp_dummy_magic_29_0.Y.n3 0.242602
R16335 two_stage_opamp_dummy_magic_29_0.Y.n61 two_stage_opamp_dummy_magic_29_0.Y.n47 0.1255
R16336 two_stage_opamp_dummy_magic_29_0.Y.n47 two_stage_opamp_dummy_magic_29_0.Y.n46 0.0626438
R16337 two_stage_opamp_dummy_magic_29_0.Y.n85 two_stage_opamp_dummy_magic_29_0.Y.n37 0.0421667
R16338 two_stage_opamp_dummy_magic_29_0.Y.n20 two_stage_opamp_dummy_magic_29_0.Y.n19 0.0250536
R16339 two_stage_opamp_dummy_magic_29_0.Y.n21 two_stage_opamp_dummy_magic_29_0.Y.n20 0.0250536
R16340 two_stage_opamp_dummy_magic_29_0.Y.n21 two_stage_opamp_dummy_magic_29_0.Y.n0 0.0250536
R16341 two_stage_opamp_dummy_magic_29_0.Y.n125 two_stage_opamp_dummy_magic_29_0.Y.n2 0.0250536
R16342 two_stage_opamp_dummy_magic_29_0.Y.n121 two_stage_opamp_dummy_magic_29_0.Y.n2 0.0250536
R16343 two_stage_opamp_dummy_magic_29_0.Y.n121 two_stage_opamp_dummy_magic_29_0.Y.n120 0.0250536
R16344 two_stage_opamp_dummy_magic_29_0.Y.n120 two_stage_opamp_dummy_magic_29_0.Y.n119 0.0250536
R16345 two_stage_opamp_dummy_magic_29_0.Y.n22 two_stage_opamp_dummy_magic_29_0.Y.n3 0.0250536
R16346 two_stage_opamp_dummy_magic_29_0.Y.n23 two_stage_opamp_dummy_magic_29_0.Y.n22 0.0250536
R16347 two_stage_opamp_dummy_magic_29_0.Y.n124 two_stage_opamp_dummy_magic_29_0.Y.n23 0.0250536
R16348 two_stage_opamp_dummy_magic_29_0.Y.n124 two_stage_opamp_dummy_magic_29_0.Y.n123 0.0250536
R16349 two_stage_opamp_dummy_magic_29_0.Y.n123 two_stage_opamp_dummy_magic_29_0.Y.n122 0.0250536
R16350 two_stage_opamp_dummy_magic_29_0.Y.n122 two_stage_opamp_dummy_magic_29_0.Y.n24 0.0250536
R16351 two_stage_opamp_dummy_magic_29_0.Y.n118 two_stage_opamp_dummy_magic_29_0.Y.n24 0.0250536
R16352 two_stage_opamp_dummy_magic_29_0.Y.n19 two_stage_opamp_dummy_magic_29_0.Y.n18 0.024102
R16353 two_stage_opamp_dummy_magic_29_0.Y.n33 two_stage_opamp_dummy_magic_29_0.Y.n30 0.0217373
R16354 two_stage_opamp_dummy_magic_29_0.Y.n116 two_stage_opamp_dummy_magic_29_0.Y.n31 0.0217373
R16355 two_stage_opamp_dummy_magic_29_0.Y.n32 two_stage_opamp_dummy_magic_29_0.Y.n26 0.0217373
R16356 two_stage_opamp_dummy_magic_29_0.Y.n87 two_stage_opamp_dummy_magic_29_0.Y.n86 0.0217373
R16357 two_stage_opamp_dummy_magic_29_0.Y.n84 two_stage_opamp_dummy_magic_29_0.Y.n63 0.0217373
R16358 two_stage_opamp_dummy_magic_29_0.Y.n33 two_stage_opamp_dummy_magic_29_0.Y.n28 0.0217373
R16359 two_stage_opamp_dummy_magic_29_0.Y.n31 two_stage_opamp_dummy_magic_29_0.Y.n27 0.0217373
R16360 two_stage_opamp_dummy_magic_29_0.Y.n88 two_stage_opamp_dummy_magic_29_0.Y.n26 0.0217373
R16361 two_stage_opamp_dummy_magic_29_0.Y.n86 two_stage_opamp_dummy_magic_29_0.Y.n36 0.0217373
R16362 two_stage_opamp_dummy_magic_29_0.Y.n63 two_stage_opamp_dummy_magic_29_0.Y.n36 0.0217373
R16363 two_stage_opamp_dummy_magic_29_0.Y.n40 two_stage_opamp_dummy_magic_29_0.Y.n38 0.0217373
R16364 two_stage_opamp_dummy_magic_29_0.Y.n41 two_stage_opamp_dummy_magic_29_0.Y.n39 0.0217373
R16365 two_stage_opamp_dummy_magic_29_0.Y.n113 two_stage_opamp_dummy_magic_29_0.Y.n28 0.0217373
R16366 two_stage_opamp_dummy_magic_29_0.Y.n90 two_stage_opamp_dummy_magic_29_0.Y.n27 0.0217373
R16367 two_stage_opamp_dummy_magic_29_0.Y.n115 two_stage_opamp_dummy_magic_29_0.Y.n32 0.0217373
R16368 two_stage_opamp_dummy_magic_29_0.Y.n113 two_stage_opamp_dummy_magic_29_0.Y.n112 0.0217373
R16369 two_stage_opamp_dummy_magic_29_0.Y.n90 two_stage_opamp_dummy_magic_29_0.Y.n30 0.0217373
R16370 two_stage_opamp_dummy_magic_29_0.Y.n116 two_stage_opamp_dummy_magic_29_0.Y.n115 0.0217373
R16371 two_stage_opamp_dummy_magic_29_0.Y.n83 two_stage_opamp_dummy_magic_29_0.Y.n35 0.0217373
R16372 two_stage_opamp_dummy_magic_29_0.Y.n44 two_stage_opamp_dummy_magic_29_0.Y.n39 0.0217373
R16373 two_stage_opamp_dummy_magic_29_0.Y.n37 two_stage_opamp_dummy_magic_29_0.Y.n35 0.0217373
R16374 two_stage_opamp_dummy_magic_29_0.Y.n42 two_stage_opamp_dummy_magic_29_0.Y.n40 0.0217373
R16375 two_stage_opamp_dummy_magic_29_0.Y.n43 two_stage_opamp_dummy_magic_29_0.Y.n42 0.0217373
R16376 two_stage_opamp_dummy_magic_29_0.Y.n45 two_stage_opamp_dummy_magic_29_0.Y.n44 0.0217373
R16377 two_stage_opamp_dummy_magic_29_0.Y two_stage_opamp_dummy_magic_29_0.Y.n0 0.016125
R16378 two_stage_opamp_dummy_magic_29_0.Y.n34 two_stage_opamp_dummy_magic_29_0.Y.n29 0.00991089
R16379 two_stage_opamp_dummy_magic_29_0.Y.n114 two_stage_opamp_dummy_magic_29_0.Y.n89 0.00991089
R16380 two_stage_opamp_dummy_magic_29_0.Y.n117 two_stage_opamp_dummy_magic_29_0.Y.n29 0.00991089
R16381 two_stage_opamp_dummy_magic_29_0.Y.n89 two_stage_opamp_dummy_magic_29_0.Y.n34 0.00991089
R16382 two_stage_opamp_dummy_magic_29_0.Y two_stage_opamp_dummy_magic_29_0.Y.n125 0.00942857
R16383 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t11 115.6
R16384 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n0 107.121
R16385 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n1 97.4332
R16386 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n2 28.6724
R16387 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n5 24.288
R16388 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n7 24.288
R16389 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n11 24.288
R16390 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n14 24.288
R16391 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n17 24.288
R16392 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t13 24.0005
R16393 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t14 24.0005
R16394 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t12 24.0005
R16395 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t0 24.0005
R16396 bgr_11_0.V_CMFB_S4 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n20 17.464
R16397 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t10 8.0005
R16398 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t3 8.0005
R16399 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t7 8.0005
R16400 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t2 8.0005
R16401 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t6 8.0005
R16402 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t1 8.0005
R16403 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t9 8.0005
R16404 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n14 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t5 8.0005
R16405 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t8 8.0005
R16406 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t4 8.0005
R16407 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n16 5.7505
R16408 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n6 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n4 5.7505
R16409 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n6 5.53175
R16410 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n8 5.188
R16411 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n4 5.188
R16412 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n10 5.188
R16413 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n12 5.188
R16414 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n3 5.188
R16415 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n15 5.188
R16416 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n18 5.188
R16417 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n19 2.38069
R16418 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n13 0.563
R16419 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n4 0.563
R16420 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n9 0.34425
R16421 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n10 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n3 0.34425
R16422 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n3 0.34425
R16423 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t28 610.534
R16424 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t26 610.534
R16425 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n27 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t17 433.8
R16426 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t14 433.8
R16427 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t23 433.8
R16428 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t31 433.8
R16429 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t20 433.8
R16430 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t30 433.8
R16431 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t19 433.8
R16432 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n34 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t29 433.8
R16433 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n35 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t12 433.8
R16434 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t27 433.8
R16435 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t16 433.8
R16436 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t25 433.8
R16437 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t15 433.8
R16438 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t24 433.8
R16439 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t13 433.8
R16440 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n6 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t22 433.8
R16441 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t21 433.8
R16442 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t18 433.8
R16443 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n2 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n14 287.264
R16444 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n18 287.264
R16445 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n15 287.264
R16446 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n21 287.264
R16447 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n35 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n34 176.733
R16448 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n34 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n33 176.733
R16449 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n33 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n32 176.733
R16450 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n32 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n31 176.733
R16451 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n31 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n30 176.733
R16452 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n30 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n29 176.733
R16453 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n29 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n28 176.733
R16454 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n28 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n27 176.733
R16455 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n7 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n6 176.733
R16456 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n8 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n7 176.733
R16457 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n9 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n8 176.733
R16458 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n10 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n9 176.733
R16459 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n11 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n10 176.733
R16460 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n12 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n11 176.733
R16461 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n26 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n25 176.733
R16462 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n37 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n36 161.986
R16463 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_tail_gate.n13 161.986
R16464 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n0 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n22 56.7378
R16465 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n19 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n0 56.737
R16466 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n2 56.737
R16467 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n2 52.5725
R16468 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n22 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n20 52.5725
R16469 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n19 52.01
R16470 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n17 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n16 52.01
R16471 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n23 49.7255
R16472 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n5 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n4 49.7255
R16473 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n16 two_stage_opamp_dummy_magic_29_0.V_tail_gate 46.7517
R16474 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n36 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n35 45.5227
R16475 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n13 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n12 45.5227
R16476 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n25 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n13 45.5227
R16477 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n36 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n26 45.5227
R16478 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t6 39.4005
R16479 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n21 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t2 39.4005
R16480 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t8 39.4005
R16481 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n18 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t5 39.4005
R16482 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t7 39.4005
R16483 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n15 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t3 39.4005
R16484 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t4 39.4005
R16485 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n14 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t9 39.4005
R16486 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t0 16.0005
R16487 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n23 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t10 16.0005
R16488 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t11 16.0005
R16489 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n4 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t1 16.0005
R16490 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_tail_gate.n3 9.98584
R16491 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n24 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n5 9.563
R16492 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n0 6.53418
R16493 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_tail_gate.n1 1.56177
R16494 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n1 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n37 1.44719
R16495 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n37 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n24 0.842037
R16496 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_tail_gate.n5 0.842037
R16497 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n20 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n17 0.563
R16498 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n3 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n0 0.340844
R16499 two_stage_opamp_dummy_magic_29_0.V_source.n59 two_stage_opamp_dummy_magic_29_0.V_source.t5 67.545
R16500 two_stage_opamp_dummy_magic_29_0.V_source.n28 two_stage_opamp_dummy_magic_29_0.V_source.n27 49.3505
R16501 two_stage_opamp_dummy_magic_29_0.V_source.n26 two_stage_opamp_dummy_magic_29_0.V_source.n25 49.3505
R16502 two_stage_opamp_dummy_magic_29_0.V_source.n16 two_stage_opamp_dummy_magic_29_0.V_source.n15 49.3505
R16503 two_stage_opamp_dummy_magic_29_0.V_source.n34 two_stage_opamp_dummy_magic_29_0.V_source.n33 49.3505
R16504 two_stage_opamp_dummy_magic_29_0.V_source.n31 two_stage_opamp_dummy_magic_29_0.V_source.n30 49.3505
R16505 two_stage_opamp_dummy_magic_29_0.V_source.n43 two_stage_opamp_dummy_magic_29_0.V_source.n42 49.3505
R16506 two_stage_opamp_dummy_magic_29_0.V_source.n39 two_stage_opamp_dummy_magic_29_0.V_source.n38 49.3505
R16507 two_stage_opamp_dummy_magic_29_0.V_source.n37 two_stage_opamp_dummy_magic_29_0.V_source.n36 49.3505
R16508 two_stage_opamp_dummy_magic_29_0.V_source.n22 two_stage_opamp_dummy_magic_29_0.V_source.n21 49.3505
R16509 two_stage_opamp_dummy_magic_29_0.V_source.n18 two_stage_opamp_dummy_magic_29_0.V_source.n17 49.3505
R16510 two_stage_opamp_dummy_magic_29_0.V_source.n6 two_stage_opamp_dummy_magic_29_0.V_source.n5 32.3838
R16511 two_stage_opamp_dummy_magic_29_0.V_source.n68 two_stage_opamp_dummy_magic_29_0.V_source.n67 32.3838
R16512 two_stage_opamp_dummy_magic_29_0.V_source.n49 two_stage_opamp_dummy_magic_29_0.V_source.n48 32.3838
R16513 two_stage_opamp_dummy_magic_29_0.V_source.n47 two_stage_opamp_dummy_magic_29_0.V_source.n46 32.3838
R16514 two_stage_opamp_dummy_magic_29_0.V_source.n53 two_stage_opamp_dummy_magic_29_0.V_source.n52 32.3838
R16515 two_stage_opamp_dummy_magic_29_0.V_source.n56 two_stage_opamp_dummy_magic_29_0.V_source.n55 32.3838
R16516 two_stage_opamp_dummy_magic_29_0.V_source.n9 two_stage_opamp_dummy_magic_29_0.V_source.n8 32.3838
R16517 two_stage_opamp_dummy_magic_29_0.V_source.n74 two_stage_opamp_dummy_magic_29_0.V_source.n73 32.3838
R16518 two_stage_opamp_dummy_magic_29_0.V_source.n78 two_stage_opamp_dummy_magic_29_0.V_source.n77 32.3838
R16519 two_stage_opamp_dummy_magic_29_0.V_source.n71 two_stage_opamp_dummy_magic_29_0.V_source.n70 32.3838
R16520 two_stage_opamp_dummy_magic_29_0.V_source.n27 two_stage_opamp_dummy_magic_29_0.V_source.t18 16.0005
R16521 two_stage_opamp_dummy_magic_29_0.V_source.n27 two_stage_opamp_dummy_magic_29_0.V_source.t17 16.0005
R16522 two_stage_opamp_dummy_magic_29_0.V_source.n25 two_stage_opamp_dummy_magic_29_0.V_source.t0 16.0005
R16523 two_stage_opamp_dummy_magic_29_0.V_source.n25 two_stage_opamp_dummy_magic_29_0.V_source.t21 16.0005
R16524 two_stage_opamp_dummy_magic_29_0.V_source.n15 two_stage_opamp_dummy_magic_29_0.V_source.t14 16.0005
R16525 two_stage_opamp_dummy_magic_29_0.V_source.n15 two_stage_opamp_dummy_magic_29_0.V_source.t19 16.0005
R16526 two_stage_opamp_dummy_magic_29_0.V_source.n33 two_stage_opamp_dummy_magic_29_0.V_source.t1 16.0005
R16527 two_stage_opamp_dummy_magic_29_0.V_source.n33 two_stage_opamp_dummy_magic_29_0.V_source.t10 16.0005
R16528 two_stage_opamp_dummy_magic_29_0.V_source.n30 two_stage_opamp_dummy_magic_29_0.V_source.t12 16.0005
R16529 two_stage_opamp_dummy_magic_29_0.V_source.n30 two_stage_opamp_dummy_magic_29_0.V_source.t40 16.0005
R16530 two_stage_opamp_dummy_magic_29_0.V_source.n42 two_stage_opamp_dummy_magic_29_0.V_source.t8 16.0005
R16531 two_stage_opamp_dummy_magic_29_0.V_source.n42 two_stage_opamp_dummy_magic_29_0.V_source.t9 16.0005
R16532 two_stage_opamp_dummy_magic_29_0.V_source.n38 two_stage_opamp_dummy_magic_29_0.V_source.t6 16.0005
R16533 two_stage_opamp_dummy_magic_29_0.V_source.n38 two_stage_opamp_dummy_magic_29_0.V_source.t2 16.0005
R16534 two_stage_opamp_dummy_magic_29_0.V_source.n36 two_stage_opamp_dummy_magic_29_0.V_source.t7 16.0005
R16535 two_stage_opamp_dummy_magic_29_0.V_source.n36 two_stage_opamp_dummy_magic_29_0.V_source.t11 16.0005
R16536 two_stage_opamp_dummy_magic_29_0.V_source.n21 two_stage_opamp_dummy_magic_29_0.V_source.t20 16.0005
R16537 two_stage_opamp_dummy_magic_29_0.V_source.n21 two_stage_opamp_dummy_magic_29_0.V_source.t16 16.0005
R16538 two_stage_opamp_dummy_magic_29_0.V_source.n17 two_stage_opamp_dummy_magic_29_0.V_source.t4 16.0005
R16539 two_stage_opamp_dummy_magic_29_0.V_source.n17 two_stage_opamp_dummy_magic_29_0.V_source.t15 16.0005
R16540 two_stage_opamp_dummy_magic_29_0.V_source.n5 two_stage_opamp_dummy_magic_29_0.V_source.t13 9.6005
R16541 two_stage_opamp_dummy_magic_29_0.V_source.n5 two_stage_opamp_dummy_magic_29_0.V_source.t3 9.6005
R16542 two_stage_opamp_dummy_magic_29_0.V_source.n67 two_stage_opamp_dummy_magic_29_0.V_source.t32 9.6005
R16543 two_stage_opamp_dummy_magic_29_0.V_source.n67 two_stage_opamp_dummy_magic_29_0.V_source.t22 9.6005
R16544 two_stage_opamp_dummy_magic_29_0.V_source.n48 two_stage_opamp_dummy_magic_29_0.V_source.t33 9.6005
R16545 two_stage_opamp_dummy_magic_29_0.V_source.n48 two_stage_opamp_dummy_magic_29_0.V_source.t23 9.6005
R16546 two_stage_opamp_dummy_magic_29_0.V_source.n46 two_stage_opamp_dummy_magic_29_0.V_source.t29 9.6005
R16547 two_stage_opamp_dummy_magic_29_0.V_source.n46 two_stage_opamp_dummy_magic_29_0.V_source.t37 9.6005
R16548 two_stage_opamp_dummy_magic_29_0.V_source.n52 two_stage_opamp_dummy_magic_29_0.V_source.t38 9.6005
R16549 two_stage_opamp_dummy_magic_29_0.V_source.n52 two_stage_opamp_dummy_magic_29_0.V_source.t28 9.6005
R16550 two_stage_opamp_dummy_magic_29_0.V_source.n55 two_stage_opamp_dummy_magic_29_0.V_source.t26 9.6005
R16551 two_stage_opamp_dummy_magic_29_0.V_source.n55 two_stage_opamp_dummy_magic_29_0.V_source.t30 9.6005
R16552 two_stage_opamp_dummy_magic_29_0.V_source.n8 two_stage_opamp_dummy_magic_29_0.V_source.t36 9.6005
R16553 two_stage_opamp_dummy_magic_29_0.V_source.n8 two_stage_opamp_dummy_magic_29_0.V_source.t27 9.6005
R16554 two_stage_opamp_dummy_magic_29_0.V_source.n73 two_stage_opamp_dummy_magic_29_0.V_source.t34 9.6005
R16555 two_stage_opamp_dummy_magic_29_0.V_source.n73 two_stage_opamp_dummy_magic_29_0.V_source.t31 9.6005
R16556 two_stage_opamp_dummy_magic_29_0.V_source.n77 two_stage_opamp_dummy_magic_29_0.V_source.t35 9.6005
R16557 two_stage_opamp_dummy_magic_29_0.V_source.n77 two_stage_opamp_dummy_magic_29_0.V_source.t25 9.6005
R16558 two_stage_opamp_dummy_magic_29_0.V_source.n70 two_stage_opamp_dummy_magic_29_0.V_source.t39 9.6005
R16559 two_stage_opamp_dummy_magic_29_0.V_source.n70 two_stage_opamp_dummy_magic_29_0.V_source.t24 9.6005
R16560 two_stage_opamp_dummy_magic_29_0.V_source.n80 two_stage_opamp_dummy_magic_29_0.V_source.n6 5.85227
R16561 two_stage_opamp_dummy_magic_29_0.V_source.n37 two_stage_opamp_dummy_magic_29_0.V_source.n13 5.51092
R16562 two_stage_opamp_dummy_magic_29_0.V_source.n19 two_stage_opamp_dummy_magic_29_0.V_source.n16 5.51092
R16563 two_stage_opamp_dummy_magic_29_0.V_source.n40 two_stage_opamp_dummy_magic_29_0.V_source.n37 5.45883
R16564 two_stage_opamp_dummy_magic_29_0.V_source.n16 two_stage_opamp_dummy_magic_29_0.V_source.n14 5.45883
R16565 two_stage_opamp_dummy_magic_29_0.V_source.n71 two_stage_opamp_dummy_magic_29_0.V_source.n69 5.188
R16566 two_stage_opamp_dummy_magic_29_0.V_source.n74 two_stage_opamp_dummy_magic_29_0.V_source.n7 5.188
R16567 two_stage_opamp_dummy_magic_29_0.V_source.n79 two_stage_opamp_dummy_magic_29_0.V_source.n78 5.188
R16568 two_stage_opamp_dummy_magic_29_0.V_source.n44 two_stage_opamp_dummy_magic_29_0.V_source.n43 5.16717
R16569 two_stage_opamp_dummy_magic_29_0.V_source.n39 two_stage_opamp_dummy_magic_29_0.V_source.n13 5.16717
R16570 two_stage_opamp_dummy_magic_29_0.V_source.n22 two_stage_opamp_dummy_magic_29_0.V_source.n20 5.16717
R16571 two_stage_opamp_dummy_magic_29_0.V_source.n19 two_stage_opamp_dummy_magic_29_0.V_source.n18 5.16717
R16572 two_stage_opamp_dummy_magic_29_0.V_source.n35 two_stage_opamp_dummy_magic_29_0.V_source.n34 4.89633
R16573 two_stage_opamp_dummy_magic_29_0.V_source.n43 two_stage_opamp_dummy_magic_29_0.V_source.n41 4.89633
R16574 two_stage_opamp_dummy_magic_29_0.V_source.n40 two_stage_opamp_dummy_magic_29_0.V_source.n39 4.89633
R16575 two_stage_opamp_dummy_magic_29_0.V_source.n29 two_stage_opamp_dummy_magic_29_0.V_source.n28 4.89633
R16576 two_stage_opamp_dummy_magic_29_0.V_source.n32 two_stage_opamp_dummy_magic_29_0.V_source.n31 4.89633
R16577 two_stage_opamp_dummy_magic_29_0.V_source.n23 two_stage_opamp_dummy_magic_29_0.V_source.n22 4.89633
R16578 two_stage_opamp_dummy_magic_29_0.V_source.n18 two_stage_opamp_dummy_magic_29_0.V_source.n14 4.89633
R16579 two_stage_opamp_dummy_magic_29_0.V_source.n26 two_stage_opamp_dummy_magic_29_0.V_source.n24 4.89633
R16580 two_stage_opamp_dummy_magic_29_0.V_source.n60 two_stage_opamp_dummy_magic_29_0.V_source.n50 4.5005
R16581 two_stage_opamp_dummy_magic_29_0.V_source.n62 two_stage_opamp_dummy_magic_29_0.V_source.n61 4.5005
R16582 two_stage_opamp_dummy_magic_29_0.V_source.n61 two_stage_opamp_dummy_magic_29_0.V_source.n60 4.5005
R16583 two_stage_opamp_dummy_magic_29_0.V_source.n32 two_stage_opamp_dummy_magic_29_0.V_source.n29 3.6255
R16584 two_stage_opamp_dummy_magic_29_0.V_source.n68 two_stage_opamp_dummy_magic_29_0.V_source.n66 2.98664
R16585 two_stage_opamp_dummy_magic_29_0.V_source.n49 two_stage_opamp_dummy_magic_29_0.V_source.n11 2.98664
R16586 two_stage_opamp_dummy_magic_29_0.V_source.n65 two_stage_opamp_dummy_magic_29_0.V_source.n47 2.98664
R16587 two_stage_opamp_dummy_magic_29_0.V_source.n54 two_stage_opamp_dummy_magic_29_0.V_source.n53 2.98664
R16588 two_stage_opamp_dummy_magic_29_0.V_source.n57 two_stage_opamp_dummy_magic_29_0.V_source.n56 2.98664
R16589 two_stage_opamp_dummy_magic_29_0.V_source.n10 two_stage_opamp_dummy_magic_29_0.V_source.n9 2.98664
R16590 two_stage_opamp_dummy_magic_29_0.V_source.n75 two_stage_opamp_dummy_magic_29_0.V_source.n74 2.98664
R16591 two_stage_opamp_dummy_magic_29_0.V_source.n78 two_stage_opamp_dummy_magic_29_0.V_source.n76 2.98664
R16592 two_stage_opamp_dummy_magic_29_0.V_source.n58 two_stage_opamp_dummy_magic_29_0.V_source.n6 2.98664
R16593 two_stage_opamp_dummy_magic_29_0.V_source.n72 two_stage_opamp_dummy_magic_29_0.V_source.n71 2.98628
R16594 two_stage_opamp_dummy_magic_29_0.V_source.n63 two_stage_opamp_dummy_magic_29_0.V_source.n62 2.24063
R16595 two_stage_opamp_dummy_magic_29_0.V_source.n51 two_stage_opamp_dummy_magic_29_0.V_source.n0 2.24063
R16596 two_stage_opamp_dummy_magic_29_0.V_source.n64 two_stage_opamp_dummy_magic_29_0.V_source.n0 2.24063
R16597 two_stage_opamp_dummy_magic_29_0.V_source.n45 two_stage_opamp_dummy_magic_29_0.V_source.n12 2.2076
R16598 two_stage_opamp_dummy_magic_29_0.V_source.n1 two_stage_opamp_dummy_magic_29_0.V_source.n45 2.16822
R16599 two_stage_opamp_dummy_magic_29_0.V_source.n12 two_stage_opamp_dummy_magic_29_0.V_source.n3 2.16822
R16600 two_stage_opamp_dummy_magic_29_0.V_source.n69 two_stage_opamp_dummy_magic_29_0.V_source.n2 2.02255
R16601 two_stage_opamp_dummy_magic_29_0.V_source.n4 two_stage_opamp_dummy_magic_29_0.V_source.n80 1.36007
R16602 two_stage_opamp_dummy_magic_29_0.V_source.n60 two_stage_opamp_dummy_magic_29_0.V_source.n59 0.922375
R16603 two_stage_opamp_dummy_magic_29_0.V_source.n59 two_stage_opamp_dummy_magic_29_0.V_source.n58 2.52416
R16604 two_stage_opamp_dummy_magic_29_0.V_source.n80 two_stage_opamp_dummy_magic_29_0.V_source.n79 0.664374
R16605 two_stage_opamp_dummy_magic_29_0.V_source.n2 two_stage_opamp_dummy_magic_29_0.V_source.n47 0.6255
R16606 two_stage_opamp_dummy_magic_29_0.V_source.n2 two_stage_opamp_dummy_magic_29_0.V_source.n49 0.6255
R16607 two_stage_opamp_dummy_magic_29_0.V_source.n2 two_stage_opamp_dummy_magic_29_0.V_source.n68 0.6255
R16608 two_stage_opamp_dummy_magic_29_0.V_source.n9 two_stage_opamp_dummy_magic_29_0.V_source.n4 0.6255
R16609 two_stage_opamp_dummy_magic_29_0.V_source.n56 two_stage_opamp_dummy_magic_29_0.V_source.n4 0.6255
R16610 two_stage_opamp_dummy_magic_29_0.V_source.n53 two_stage_opamp_dummy_magic_29_0.V_source.n4 0.6255
R16611 two_stage_opamp_dummy_magic_29_0.V_source.n31 two_stage_opamp_dummy_magic_29_0.V_source.n1 0.604667
R16612 two_stage_opamp_dummy_magic_29_0.V_source.n34 two_stage_opamp_dummy_magic_29_0.V_source.n1 0.604667
R16613 two_stage_opamp_dummy_magic_29_0.V_source.n3 two_stage_opamp_dummy_magic_29_0.V_source.n26 0.604667
R16614 two_stage_opamp_dummy_magic_29_0.V_source.n28 two_stage_opamp_dummy_magic_29_0.V_source.n3 0.604667
R16615 two_stage_opamp_dummy_magic_29_0.V_source.n41 two_stage_opamp_dummy_magic_29_0.V_source.n40 0.563
R16616 two_stage_opamp_dummy_magic_29_0.V_source.n41 two_stage_opamp_dummy_magic_29_0.V_source.n35 0.563
R16617 two_stage_opamp_dummy_magic_29_0.V_source.n35 two_stage_opamp_dummy_magic_29_0.V_source.n32 0.563
R16618 two_stage_opamp_dummy_magic_29_0.V_source.n29 two_stage_opamp_dummy_magic_29_0.V_source.n24 0.563
R16619 two_stage_opamp_dummy_magic_29_0.V_source.n23 two_stage_opamp_dummy_magic_29_0.V_source.n14 0.563
R16620 two_stage_opamp_dummy_magic_29_0.V_source.n24 two_stage_opamp_dummy_magic_29_0.V_source.n23 0.563
R16621 two_stage_opamp_dummy_magic_29_0.V_source.n20 two_stage_opamp_dummy_magic_29_0.V_source.n12 0.510302
R16622 two_stage_opamp_dummy_magic_29_0.V_source.n45 two_stage_opamp_dummy_magic_29_0.V_source.n44 0.510302
R16623 two_stage_opamp_dummy_magic_29_0.V_source.n20 two_stage_opamp_dummy_magic_29_0.V_source.n19 0.34425
R16624 two_stage_opamp_dummy_magic_29_0.V_source.n44 two_stage_opamp_dummy_magic_29_0.V_source.n13 0.34425
R16625 two_stage_opamp_dummy_magic_29_0.V_source.n79 two_stage_opamp_dummy_magic_29_0.V_source.n7 0.34425
R16626 two_stage_opamp_dummy_magic_29_0.V_source.n69 two_stage_opamp_dummy_magic_29_0.V_source.n7 0.34425
R16627 two_stage_opamp_dummy_magic_29_0.V_source.n65 two_stage_opamp_dummy_magic_29_0.V_source.n64 1.51368
R16628 two_stage_opamp_dummy_magic_29_0.V_source.n2 two_stage_opamp_dummy_magic_29_0.V_source.n1 0.216846
R16629 two_stage_opamp_dummy_magic_29_0.V_source two_stage_opamp_dummy_magic_29_0.V_source.n3 0.120692
R16630 two_stage_opamp_dummy_magic_29_0.V_source.n58 two_stage_opamp_dummy_magic_29_0.V_source.n57 0.115083
R16631 two_stage_opamp_dummy_magic_29_0.V_source.n57 two_stage_opamp_dummy_magic_29_0.V_source.n54 0.115083
R16632 two_stage_opamp_dummy_magic_29_0.V_source.n54 two_stage_opamp_dummy_magic_29_0.V_source.n10 0.115083
R16633 two_stage_opamp_dummy_magic_29_0.V_source.n76 two_stage_opamp_dummy_magic_29_0.V_source.n10 0.115083
R16634 two_stage_opamp_dummy_magic_29_0.V_source.n76 two_stage_opamp_dummy_magic_29_0.V_source.n75 0.115083
R16635 two_stage_opamp_dummy_magic_29_0.V_source.n75 two_stage_opamp_dummy_magic_29_0.V_source.n72 0.115083
R16636 two_stage_opamp_dummy_magic_29_0.V_source.n72 two_stage_opamp_dummy_magic_29_0.V_source.n11 0.115083
R16637 two_stage_opamp_dummy_magic_29_0.V_source.n66 two_stage_opamp_dummy_magic_29_0.V_source.n11 0.115083
R16638 two_stage_opamp_dummy_magic_29_0.V_source.n66 two_stage_opamp_dummy_magic_29_0.V_source.n65 0.115083
R16639 two_stage_opamp_dummy_magic_29_0.V_source two_stage_opamp_dummy_magic_29_0.V_source.n4 0.0966538
R16640 two_stage_opamp_dummy_magic_29_0.V_source.n62 two_stage_opamp_dummy_magic_29_0.V_source.n0 0.0421667
R16641 two_stage_opamp_dummy_magic_29_0.V_source.n64 two_stage_opamp_dummy_magic_29_0.V_source.n63 0.0217373
R16642 two_stage_opamp_dummy_magic_29_0.V_source.n61 two_stage_opamp_dummy_magic_29_0.V_source.n51 0.0217373
R16643 two_stage_opamp_dummy_magic_29_0.V_source.n63 two_stage_opamp_dummy_magic_29_0.V_source.n50 0.0217373
R16644 two_stage_opamp_dummy_magic_29_0.V_source.n51 two_stage_opamp_dummy_magic_29_0.V_source.n50 0.0217373
R16645 two_stage_opamp_dummy_magic_29_0.V_source.n60 two_stage_opamp_dummy_magic_29_0.V_source.n0 0.0429746
R16646 two_stage_opamp_dummy_magic_29_0.Vb2.n2 two_stage_opamp_dummy_magic_29_0.Vb2.t17 752.422
R16647 two_stage_opamp_dummy_magic_29_0.Vb2.n0 two_stage_opamp_dummy_magic_29_0.Vb2.t18 752.422
R16648 two_stage_opamp_dummy_magic_29_0.Vb2.n2 two_stage_opamp_dummy_magic_29_0.Vb2.t26 752.234
R16649 two_stage_opamp_dummy_magic_29_0.Vb2.n2 two_stage_opamp_dummy_magic_29_0.Vb2.t19 752.234
R16650 two_stage_opamp_dummy_magic_29_0.Vb2.n3 two_stage_opamp_dummy_magic_29_0.Vb2.t30 752.234
R16651 two_stage_opamp_dummy_magic_29_0.Vb2.n3 two_stage_opamp_dummy_magic_29_0.Vb2.t14 752.234
R16652 two_stage_opamp_dummy_magic_29_0.Vb2.n3 two_stage_opamp_dummy_magic_29_0.Vb2.t23 752.234
R16653 two_stage_opamp_dummy_magic_29_0.Vb2.n3 two_stage_opamp_dummy_magic_29_0.Vb2.t32 752.234
R16654 two_stage_opamp_dummy_magic_29_0.Vb2.n4 two_stage_opamp_dummy_magic_29_0.Vb2.t27 752.234
R16655 two_stage_opamp_dummy_magic_29_0.Vb2.n4 two_stage_opamp_dummy_magic_29_0.Vb2.t15 752.234
R16656 two_stage_opamp_dummy_magic_29_0.Vb2.n4 two_stage_opamp_dummy_magic_29_0.Vb2.t24 752.234
R16657 two_stage_opamp_dummy_magic_29_0.Vb2.n5 two_stage_opamp_dummy_magic_29_0.Vb2.t11 752.234
R16658 two_stage_opamp_dummy_magic_29_0.Vb2.n5 two_stage_opamp_dummy_magic_29_0.Vb2.t28 752.234
R16659 two_stage_opamp_dummy_magic_29_0.Vb2.n1 two_stage_opamp_dummy_magic_29_0.Vb2.t16 752.234
R16660 two_stage_opamp_dummy_magic_29_0.Vb2.n1 two_stage_opamp_dummy_magic_29_0.Vb2.t25 752.234
R16661 two_stage_opamp_dummy_magic_29_0.Vb2.n1 two_stage_opamp_dummy_magic_29_0.Vb2.t12 752.234
R16662 two_stage_opamp_dummy_magic_29_0.Vb2.n1 two_stage_opamp_dummy_magic_29_0.Vb2.t21 752.234
R16663 two_stage_opamp_dummy_magic_29_0.Vb2.n0 two_stage_opamp_dummy_magic_29_0.Vb2.t13 752.234
R16664 two_stage_opamp_dummy_magic_29_0.Vb2.n0 two_stage_opamp_dummy_magic_29_0.Vb2.t22 752.234
R16665 two_stage_opamp_dummy_magic_29_0.Vb2.n0 two_stage_opamp_dummy_magic_29_0.Vb2.t31 752.234
R16666 two_stage_opamp_dummy_magic_29_0.Vb2.n17 two_stage_opamp_dummy_magic_29_0.Vb2.t29 746.673
R16667 two_stage_opamp_dummy_magic_29_0.Vb2.n14 two_stage_opamp_dummy_magic_29_0.Vb2.t4 745.726
R16668 two_stage_opamp_dummy_magic_29_0.Vb2.n16 two_stage_opamp_dummy_magic_29_0.Vb2.t20 587.551
R16669 two_stage_opamp_dummy_magic_29_0.Vb2.n8 two_stage_opamp_dummy_magic_29_0.Vb2.n6 140.546
R16670 two_stage_opamp_dummy_magic_29_0.Vb2.n12 two_stage_opamp_dummy_magic_29_0.Vb2.n11 139.297
R16671 two_stage_opamp_dummy_magic_29_0.Vb2.n10 two_stage_opamp_dummy_magic_29_0.Vb2.n9 139.297
R16672 two_stage_opamp_dummy_magic_29_0.Vb2.n8 two_stage_opamp_dummy_magic_29_0.Vb2.n7 139.297
R16673 two_stage_opamp_dummy_magic_29_0.Vb2.n14 two_stage_opamp_dummy_magic_29_0.Vb2.n13 67.0547
R16674 bgr_11_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_29_0.Vb2.n18 36.2193
R16675 two_stage_opamp_dummy_magic_29_0.Vb2.n11 two_stage_opamp_dummy_magic_29_0.Vb2.t9 24.0005
R16676 two_stage_opamp_dummy_magic_29_0.Vb2.n11 two_stage_opamp_dummy_magic_29_0.Vb2.t6 24.0005
R16677 two_stage_opamp_dummy_magic_29_0.Vb2.n9 two_stage_opamp_dummy_magic_29_0.Vb2.t7 24.0005
R16678 two_stage_opamp_dummy_magic_29_0.Vb2.n9 two_stage_opamp_dummy_magic_29_0.Vb2.t10 24.0005
R16679 two_stage_opamp_dummy_magic_29_0.Vb2.n7 two_stage_opamp_dummy_magic_29_0.Vb2.t0 24.0005
R16680 two_stage_opamp_dummy_magic_29_0.Vb2.n7 two_stage_opamp_dummy_magic_29_0.Vb2.t1 24.0005
R16681 two_stage_opamp_dummy_magic_29_0.Vb2.n6 two_stage_opamp_dummy_magic_29_0.Vb2.t2 24.0005
R16682 two_stage_opamp_dummy_magic_29_0.Vb2.n6 two_stage_opamp_dummy_magic_29_0.Vb2.t8 24.0005
R16683 bgr_11_0.VB2_CUR_BIAS two_stage_opamp_dummy_magic_29_0.Vb2.n12 21.5317
R16684 two_stage_opamp_dummy_magic_29_0.Vb2.n15 two_stage_opamp_dummy_magic_29_0.Vb2.n4 13.5005
R16685 two_stage_opamp_dummy_magic_29_0.Vb2.n18 two_stage_opamp_dummy_magic_29_0.Vb2.n5 12.5005
R16686 two_stage_opamp_dummy_magic_29_0.Vb2.n13 two_stage_opamp_dummy_magic_29_0.Vb2.t5 11.2576
R16687 two_stage_opamp_dummy_magic_29_0.Vb2.n13 two_stage_opamp_dummy_magic_29_0.Vb2.t3 11.2576
R16688 two_stage_opamp_dummy_magic_29_0.Vb2.n10 two_stage_opamp_dummy_magic_29_0.Vb2.n8 6.21925
R16689 two_stage_opamp_dummy_magic_29_0.Vb2.n15 two_stage_opamp_dummy_magic_29_0.Vb2.n14 4.5005
R16690 two_stage_opamp_dummy_magic_29_0.Vb2.n17 two_stage_opamp_dummy_magic_29_0.Vb2.n16 3.58175
R16691 two_stage_opamp_dummy_magic_29_0.Vb2.n16 two_stage_opamp_dummy_magic_29_0.Vb2.n15 1.48488
R16692 two_stage_opamp_dummy_magic_29_0.Vb2.n12 two_stage_opamp_dummy_magic_29_0.Vb2.n10 1.2505
R16693 two_stage_opamp_dummy_magic_29_0.Vb2.n18 two_stage_opamp_dummy_magic_29_0.Vb2.n17 1.12238
R16694 two_stage_opamp_dummy_magic_29_0.Vb2.n4 two_stage_opamp_dummy_magic_29_0.Vb2.n3 0.7505
R16695 two_stage_opamp_dummy_magic_29_0.Vb2.n3 two_stage_opamp_dummy_magic_29_0.Vb2.n2 0.7505
R16696 two_stage_opamp_dummy_magic_29_0.Vb2.n1 two_stage_opamp_dummy_magic_29_0.Vb2.n0 0.7505
R16697 two_stage_opamp_dummy_magic_29_0.Vb2.n5 two_stage_opamp_dummy_magic_29_0.Vb2.n1 0.7505
R16698 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t14 115.6
R16699 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n0 107.121
R16700 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n1 97.4332
R16701 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n2 24.5317
R16702 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n17 24.288
R16703 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n14 24.288
R16704 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n11 24.288
R16705 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n7 24.288
R16706 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n5 24.288
R16707 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t1 24.0005
R16708 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t13 24.0005
R16709 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t2 24.0005
R16710 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t0 24.0005
R16711 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t11 8.0005
R16712 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t5 8.0005
R16713 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t9 8.0005
R16714 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n14 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t6 8.0005
R16715 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t10 8.0005
R16716 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n11 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t4 8.0005
R16717 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t8 8.0005
R16718 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t3 8.0005
R16719 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t7 8.0005
R16720 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t12 8.0005
R16721 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n6 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n4 5.7505
R16722 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n16 5.7505
R16723 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n6 5.53175
R16724 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n3 5.188
R16725 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n15 5.188
R16726 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n10 5.188
R16727 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n12 5.188
R16728 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n8 5.188
R16729 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n4 5.188
R16730 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n18 5.188
R16731 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n19 2.38147
R16732 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n13 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n4 0.563
R16733 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n13 0.563
R16734 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n3 0.34425
R16735 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n3 0.34425
R16736 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n10 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n9 0.34425
R16737 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n20 0.0213333
R16738 VOUT-.n179 VOUT-.t0 110.386
R16739 VOUT-.n39 VOUT-.n38 34.9935
R16740 VOUT-.n28 VOUT-.n27 34.9935
R16741 VOUT-.n30 VOUT-.n29 34.9935
R16742 VOUT-.n33 VOUT-.n32 34.9935
R16743 VOUT-.n36 VOUT-.n35 34.9935
R16744 VOUT-.n42 VOUT-.n41 34.9935
R16745 VOUT-.n186 VOUT-.n185 9.73997
R16746 VOUT-.n182 VOUT-.n181 9.73997
R16747 VOUT-.n189 VOUT-.n188 9.73997
R16748 VOUT-.n187 VOUT-.n182 6.64633
R16749 VOUT-.n187 VOUT-.n186 6.64633
R16750 VOUT-.n38 VOUT-.t12 6.56717
R16751 VOUT-.n38 VOUT-.t5 6.56717
R16752 VOUT-.n27 VOUT-.t6 6.56717
R16753 VOUT-.n27 VOUT-.t11 6.56717
R16754 VOUT-.n29 VOUT-.t15 6.56717
R16755 VOUT-.n29 VOUT-.t9 6.56717
R16756 VOUT-.n32 VOUT-.t16 6.56717
R16757 VOUT-.n32 VOUT-.t10 6.56717
R16758 VOUT-.n35 VOUT-.t14 6.56717
R16759 VOUT-.n35 VOUT-.t8 6.56717
R16760 VOUT-.n41 VOUT-.t13 6.56717
R16761 VOUT-.n41 VOUT-.t7 6.56717
R16762 VOUT-.n31 VOUT-.n28 6.3755
R16763 VOUT-.n40 VOUT-.n39 6.3755
R16764 VOUT-.n189 VOUT-.n187 6.02133
R16765 VOUT-.n31 VOUT-.n30 5.813
R16766 VOUT-.n34 VOUT-.n33 5.813
R16767 VOUT-.n37 VOUT-.n36 5.813
R16768 VOUT-.n42 VOUT-.n40 5.813
R16769 VOUT-.n46 VOUT-.n26 5.063
R16770 VOUT-.n43 VOUT-.n19 5.063
R16771 VOUT-.n111 VOUT-.t86 4.8295
R16772 VOUT-.n110 VOUT-.t63 4.8295
R16773 VOUT-.n109 VOUT-.t103 4.8295
R16774 VOUT-.n108 VOUT-.t110 4.8295
R16775 VOUT-.n125 VOUT-.t68 4.8295
R16776 VOUT-.n126 VOUT-.t41 4.8295
R16777 VOUT-.n128 VOUT-.t31 4.8295
R16778 VOUT-.n129 VOUT-.t143 4.8295
R16779 VOUT-.n131 VOUT-.t132 4.8295
R16780 VOUT-.n132 VOUT-.t101 4.8295
R16781 VOUT-.n134 VOUT-.t26 4.8295
R16782 VOUT-.n135 VOUT-.t138 4.8295
R16783 VOUT-.n137 VOUT-.t126 4.8295
R16784 VOUT-.n138 VOUT-.t97 4.8295
R16785 VOUT-.n140 VOUT-.t30 4.8295
R16786 VOUT-.n141 VOUT-.t140 4.8295
R16787 VOUT-.n143 VOUT-.t64 4.8295
R16788 VOUT-.n144 VOUT-.t32 4.8295
R16789 VOUT-.n146 VOUT-.t24 4.8295
R16790 VOUT-.n147 VOUT-.t133 4.8295
R16791 VOUT-.n149 VOUT-.t123 4.8295
R16792 VOUT-.n150 VOUT-.t92 4.8295
R16793 VOUT-.n71 VOUT-.t113 4.8295
R16794 VOUT-.n73 VOUT-.t131 4.8295
R16795 VOUT-.n87 VOUT-.t29 4.8295
R16796 VOUT-.n88 VOUT-.t141 4.8295
R16797 VOUT-.n90 VOUT-.t137 4.8295
R16798 VOUT-.n91 VOUT-.t104 4.8295
R16799 VOUT-.n93 VOUT-.t35 4.8295
R16800 VOUT-.n94 VOUT-.t146 4.8295
R16801 VOUT-.n96 VOUT-.t75 4.8295
R16802 VOUT-.n97 VOUT-.t44 4.8295
R16803 VOUT-.n99 VOUT-.t40 4.8295
R16804 VOUT-.n100 VOUT-.t150 4.8295
R16805 VOUT-.n102 VOUT-.t79 4.8295
R16806 VOUT-.n103 VOUT-.t49 4.8295
R16807 VOUT-.n105 VOUT-.t121 4.8295
R16808 VOUT-.n106 VOUT-.t87 4.8295
R16809 VOUT-.n152 VOUT-.t21 4.8295
R16810 VOUT-.n112 VOUT-.t144 4.8154
R16811 VOUT-.n115 VOUT-.t34 4.8154
R16812 VOUT-.n113 VOUT-.t117 4.81305
R16813 VOUT-.n116 VOUT-.t156 4.81305
R16814 VOUT-.n114 VOUT-.t139 4.806
R16815 VOUT-.n117 VOUT-.t54 4.806
R16816 VOUT-.n118 VOUT-.t88 4.806
R16817 VOUT-.n74 VOUT-.t108 4.806
R16818 VOUT-.n75 VOUT-.t154 4.806
R16819 VOUT-.n76 VOUT-.t72 4.806
R16820 VOUT-.n77 VOUT-.t22 4.806
R16821 VOUT-.n78 VOUT-.t65 4.806
R16822 VOUT-.n79 VOUT-.t160 4.806
R16823 VOUT-.n80 VOUT-.t105 4.806
R16824 VOUT-.n81 VOUT-.t56 4.806
R16825 VOUT-.n82 VOUT-.t96 4.806
R16826 VOUT-.n83 VOUT-.t47 4.806
R16827 VOUT-.n84 VOUT-.t134 4.806
R16828 VOUT-.n85 VOUT-.t36 4.806
R16829 VOUT-.n111 VOUT-.t125 4.5005
R16830 VOUT-.n110 VOUT-.t106 4.5005
R16831 VOUT-.n109 VOUT-.t145 4.5005
R16832 VOUT-.n108 VOUT-.t135 4.5005
R16833 VOUT-.n124 VOUT-.t98 4.5005
R16834 VOUT-.n123 VOUT-.t60 4.5005
R16835 VOUT-.n122 VOUT-.t80 4.5005
R16836 VOUT-.n121 VOUT-.t43 4.5005
R16837 VOUT-.n120 VOUT-.t149 4.5005
R16838 VOUT-.n119 VOUT-.t25 4.5005
R16839 VOUT-.n118 VOUT-.t128 4.5005
R16840 VOUT-.n117 VOUT-.t90 4.5005
R16841 VOUT-.n116 VOUT-.t55 4.5005
R16842 VOUT-.n115 VOUT-.t74 4.5005
R16843 VOUT-.n114 VOUT-.t37 4.5005
R16844 VOUT-.n113 VOUT-.t20 4.5005
R16845 VOUT-.n112 VOUT-.t42 4.5005
R16846 VOUT-.n125 VOUT-.t94 4.5005
R16847 VOUT-.n127 VOUT-.t59 4.5005
R16848 VOUT-.n126 VOUT-.t19 4.5005
R16849 VOUT-.n128 VOUT-.t58 4.5005
R16850 VOUT-.n130 VOUT-.t161 4.5005
R16851 VOUT-.n129 VOUT-.t116 4.5005
R16852 VOUT-.n131 VOUT-.t159 4.5005
R16853 VOUT-.n133 VOUT-.t114 4.5005
R16854 VOUT-.n132 VOUT-.t76 4.5005
R16855 VOUT-.n134 VOUT-.t53 4.5005
R16856 VOUT-.n136 VOUT-.t153 4.5005
R16857 VOUT-.n135 VOUT-.t111 4.5005
R16858 VOUT-.n137 VOUT-.t152 4.5005
R16859 VOUT-.n139 VOUT-.t109 4.5005
R16860 VOUT-.n138 VOUT-.t69 4.5005
R16861 VOUT-.n140 VOUT-.t120 4.5005
R16862 VOUT-.n142 VOUT-.t85 4.5005
R16863 VOUT-.n141 VOUT-.t50 4.5005
R16864 VOUT-.n143 VOUT-.t157 4.5005
R16865 VOUT-.n145 VOUT-.t118 4.5005
R16866 VOUT-.n144 VOUT-.t82 4.5005
R16867 VOUT-.n146 VOUT-.t112 4.5005
R16868 VOUT-.n148 VOUT-.t77 4.5005
R16869 VOUT-.n147 VOUT-.t45 4.5005
R16870 VOUT-.n149 VOUT-.t71 4.5005
R16871 VOUT-.n151 VOUT-.t39 4.5005
R16872 VOUT-.n150 VOUT-.t148 4.5005
R16873 VOUT-.n71 VOUT-.t73 4.5005
R16874 VOUT-.n72 VOUT-.t124 4.5005
R16875 VOUT-.n73 VOUT-.t78 4.5005
R16876 VOUT-.n86 VOUT-.t46 4.5005
R16877 VOUT-.n85 VOUT-.t151 4.5005
R16878 VOUT-.n84 VOUT-.t99 4.5005
R16879 VOUT-.n83 VOUT-.t62 4.5005
R16880 VOUT-.n82 VOUT-.t27 4.5005
R16881 VOUT-.n81 VOUT-.t115 4.5005
R16882 VOUT-.n80 VOUT-.t81 4.5005
R16883 VOUT-.n79 VOUT-.t48 4.5005
R16884 VOUT-.n78 VOUT-.t155 4.5005
R16885 VOUT-.n77 VOUT-.t102 4.5005
R16886 VOUT-.n76 VOUT-.t66 4.5005
R16887 VOUT-.n75 VOUT-.t147 4.5005
R16888 VOUT-.n74 VOUT-.t91 4.5005
R16889 VOUT-.n87 VOUT-.t119 4.5005
R16890 VOUT-.n89 VOUT-.t84 4.5005
R16891 VOUT-.n88 VOUT-.t52 4.5005
R16892 VOUT-.n90 VOUT-.t83 4.5005
R16893 VOUT-.n92 VOUT-.t51 4.5005
R16894 VOUT-.n91 VOUT-.t158 4.5005
R16895 VOUT-.n93 VOUT-.t122 4.5005
R16896 VOUT-.n95 VOUT-.t89 4.5005
R16897 VOUT-.n94 VOUT-.t57 4.5005
R16898 VOUT-.n96 VOUT-.t23 4.5005
R16899 VOUT-.n98 VOUT-.t129 4.5005
R16900 VOUT-.n97 VOUT-.t93 4.5005
R16901 VOUT-.n99 VOUT-.t130 4.5005
R16902 VOUT-.n101 VOUT-.t95 4.5005
R16903 VOUT-.n100 VOUT-.t61 4.5005
R16904 VOUT-.n102 VOUT-.t28 4.5005
R16905 VOUT-.n104 VOUT-.t136 4.5005
R16906 VOUT-.n103 VOUT-.t100 4.5005
R16907 VOUT-.n105 VOUT-.t67 4.5005
R16908 VOUT-.n107 VOUT-.t33 4.5005
R16909 VOUT-.n106 VOUT-.t142 4.5005
R16910 VOUT-.n152 VOUT-.t107 4.5005
R16911 VOUT-.n153 VOUT-.t70 4.5005
R16912 VOUT-.n154 VOUT-.t38 4.5005
R16913 VOUT-.n155 VOUT-.t127 4.5005
R16914 VOUT-.n47 VOUT-.n46 4.5005
R16915 VOUT-.n45 VOUT-.n24 4.5005
R16916 VOUT-.n44 VOUT-.n23 4.5005
R16917 VOUT-.n43 VOUT-.n20 4.5005
R16918 VOUT-.n65 VOUT-.n64 4.5005
R16919 VOUT-.n16 VOUT-.n13 4.5005
R16920 VOUT-.n65 VOUT-.n13 4.5005
R16921 VOUT-.n66 VOUT-.n9 4.5005
R16922 VOUT-.n66 VOUT-.n11 4.5005
R16923 VOUT-.n66 VOUT-.n65 4.5005
R16924 VOUT-.n164 VOUT-.n69 4.5005
R16925 VOUT-.n165 VOUT-.n164 4.5005
R16926 VOUT-.n165 VOUT-.n5 4.5005
R16927 VOUT-.n166 VOUT-.n4 4.5005
R16928 VOUT-.n166 VOUT-.n165 4.5005
R16929 VOUT-.n178 VOUT-.n177 4.5005
R16930 VOUT-.n178 VOUT-.n1 4.5005
R16931 VOUT-.n174 VOUT-.n1 4.5005
R16932 VOUT-.n171 VOUT-.n1 4.5005
R16933 VOUT-.n172 VOUT-.n1 4.5005
R16934 VOUT-.n174 VOUT-.n173 4.5005
R16935 VOUT-.n173 VOUT-.n171 4.5005
R16936 VOUT-.n173 VOUT-.n172 4.5005
R16937 VOUT-.n185 VOUT-.t1 3.42907
R16938 VOUT-.n185 VOUT-.t17 3.42907
R16939 VOUT-.n181 VOUT-.t18 3.42907
R16940 VOUT-.n181 VOUT-.t4 3.42907
R16941 VOUT-.n188 VOUT-.t2 3.42907
R16942 VOUT-.n188 VOUT-.t3 3.42907
R16943 VOUT-.n63 VOUT-.n62 2.24601
R16944 VOUT-.n14 VOUT-.n8 2.24601
R16945 VOUT-.n176 VOUT-.n175 2.24601
R16946 VOUT-.n170 VOUT-.n169 2.24601
R16947 VOUT-.n163 VOUT-.n162 2.24477
R16948 VOUT-.n7 VOUT-.n2 2.24477
R16949 VOUT-.n66 VOUT-.n10 2.24063
R16950 VOUT-.n166 VOUT-.n3 2.24063
R16951 VOUT-.n173 VOUT-.n0 2.24063
R16952 VOUT-.n13 VOUT-.n12 2.24063
R16953 VOUT-.n164 VOUT-.n67 2.24063
R16954 VOUT-.n68 VOUT-.n5 2.24063
R16955 VOUT-.n177 VOUT-.n168 2.24063
R16956 VOUT-.n177 VOUT-.n167 2.24063
R16957 VOUT-.n64 VOUT-.n17 2.23934
R16958 VOUT-.n64 VOUT-.n15 2.23934
R16959 VOUT-.n186 VOUT-.n184 1.83719
R16960 VOUT-.n197 VOUT-.n182 1.72967
R16961 VOUT-.n190 VOUT-.n189 1.72967
R16962 VOUT-.n50 VOUT-.n25 1.5005
R16963 VOUT-.n52 VOUT-.n51 1.5005
R16964 VOUT-.n53 VOUT-.n22 1.5005
R16965 VOUT-.n55 VOUT-.n54 1.5005
R16966 VOUT-.n56 VOUT-.n21 1.5005
R16967 VOUT-.n58 VOUT-.n57 1.5005
R16968 VOUT-.n59 VOUT-.n18 1.5005
R16969 VOUT-.n61 VOUT-.n60 1.5005
R16970 VOUT-.n192 VOUT-.n191 1.5005
R16971 VOUT-.n193 VOUT-.n183 1.5005
R16972 VOUT-.n195 VOUT-.n194 1.5005
R16973 VOUT-.n196 VOUT-.n180 1.5005
R16974 VOUT-.n198 VOUT-.n197 1.5005
R16975 VOUT-.n30 VOUT-.n20 1.313
R16976 VOUT-.n33 VOUT-.n23 1.313
R16977 VOUT-.n36 VOUT-.n24 1.313
R16978 VOUT-.n47 VOUT-.n42 1.313
R16979 VOUT-.n28 VOUT-.n19 1.313
R16980 VOUT-.n39 VOUT-.n26 1.313
R16981 VOUT-.n162 VOUT-.n161 1.1455
R16982 VOUT-.n156 VOUT-.n6 1.13717
R16983 VOUT-.n158 VOUT-.n157 1.13717
R16984 VOUT-.n160 VOUT-.n159 1.13717
R16985 VOUT-.n165 VOUT-.n6 1.13717
R16986 VOUT-.n158 VOUT-.n7 1.13717
R16987 VOUT-.n159 VOUT-.n4 1.13717
R16988 VOUT-.n70 VOUT-.n69 1.13717
R16989 VOUT-.n62 VOUT-.n61 0.859875
R16990 VOUT-.n49 VOUT-.n26 0.715216
R16991 VOUT-.n58 VOUT-.n20 0.65675
R16992 VOUT-.n54 VOUT-.n23 0.65675
R16993 VOUT-.n52 VOUT-.n24 0.65675
R16994 VOUT-.n48 VOUT-.n47 0.65675
R16995 VOUT-.n60 VOUT-.n19 0.65675
R16996 VOUT-.n161 VOUT-.n160 0.585
R16997 VOUT-.n50 VOUT-.n49 0.564601
R16998 VOUT-.n46 VOUT-.n45 0.563
R16999 VOUT-.n45 VOUT-.n44 0.563
R17000 VOUT-.n44 VOUT-.n43 0.563
R17001 VOUT-.n34 VOUT-.n31 0.563
R17002 VOUT-.n37 VOUT-.n34 0.563
R17003 VOUT-.n40 VOUT-.n37 0.563
R17004 VOUT-.n179 VOUT-.n178 0.557792
R17005 VOUT-.n177 VOUT-.n166 0.5455
R17006 VOUT-.n124 VOUT-.n108 0.3295
R17007 VOUT-.n124 VOUT-.n123 0.3295
R17008 VOUT-.n123 VOUT-.n122 0.3295
R17009 VOUT-.n122 VOUT-.n121 0.3295
R17010 VOUT-.n121 VOUT-.n120 0.3295
R17011 VOUT-.n120 VOUT-.n119 0.3295
R17012 VOUT-.n119 VOUT-.n118 0.3295
R17013 VOUT-.n118 VOUT-.n117 0.3295
R17014 VOUT-.n117 VOUT-.n116 0.3295
R17015 VOUT-.n116 VOUT-.n115 0.3295
R17016 VOUT-.n115 VOUT-.n114 0.3295
R17017 VOUT-.n114 VOUT-.n113 0.3295
R17018 VOUT-.n113 VOUT-.n112 0.3295
R17019 VOUT-.n127 VOUT-.n125 0.3295
R17020 VOUT-.n127 VOUT-.n126 0.3295
R17021 VOUT-.n130 VOUT-.n128 0.3295
R17022 VOUT-.n130 VOUT-.n129 0.3295
R17023 VOUT-.n133 VOUT-.n131 0.3295
R17024 VOUT-.n133 VOUT-.n132 0.3295
R17025 VOUT-.n136 VOUT-.n134 0.3295
R17026 VOUT-.n136 VOUT-.n135 0.3295
R17027 VOUT-.n139 VOUT-.n137 0.3295
R17028 VOUT-.n139 VOUT-.n138 0.3295
R17029 VOUT-.n142 VOUT-.n140 0.3295
R17030 VOUT-.n142 VOUT-.n141 0.3295
R17031 VOUT-.n145 VOUT-.n143 0.3295
R17032 VOUT-.n145 VOUT-.n144 0.3295
R17033 VOUT-.n148 VOUT-.n146 0.3295
R17034 VOUT-.n148 VOUT-.n147 0.3295
R17035 VOUT-.n151 VOUT-.n149 0.3295
R17036 VOUT-.n151 VOUT-.n150 0.3295
R17037 VOUT-.n72 VOUT-.n71 0.3295
R17038 VOUT-.n86 VOUT-.n73 0.3295
R17039 VOUT-.n86 VOUT-.n85 0.3295
R17040 VOUT-.n85 VOUT-.n84 0.3295
R17041 VOUT-.n84 VOUT-.n83 0.3295
R17042 VOUT-.n83 VOUT-.n82 0.3295
R17043 VOUT-.n82 VOUT-.n81 0.3295
R17044 VOUT-.n81 VOUT-.n80 0.3295
R17045 VOUT-.n80 VOUT-.n79 0.3295
R17046 VOUT-.n79 VOUT-.n78 0.3295
R17047 VOUT-.n78 VOUT-.n77 0.3295
R17048 VOUT-.n77 VOUT-.n76 0.3295
R17049 VOUT-.n76 VOUT-.n75 0.3295
R17050 VOUT-.n75 VOUT-.n74 0.3295
R17051 VOUT-.n89 VOUT-.n87 0.3295
R17052 VOUT-.n89 VOUT-.n88 0.3295
R17053 VOUT-.n92 VOUT-.n90 0.3295
R17054 VOUT-.n92 VOUT-.n91 0.3295
R17055 VOUT-.n95 VOUT-.n93 0.3295
R17056 VOUT-.n95 VOUT-.n94 0.3295
R17057 VOUT-.n98 VOUT-.n96 0.3295
R17058 VOUT-.n98 VOUT-.n97 0.3295
R17059 VOUT-.n101 VOUT-.n99 0.3295
R17060 VOUT-.n101 VOUT-.n100 0.3295
R17061 VOUT-.n104 VOUT-.n102 0.3295
R17062 VOUT-.n104 VOUT-.n103 0.3295
R17063 VOUT-.n107 VOUT-.n105 0.3295
R17064 VOUT-.n107 VOUT-.n106 0.3295
R17065 VOUT-.n153 VOUT-.n152 0.3295
R17066 VOUT-.n154 VOUT-.n153 0.3295
R17067 VOUT-.n192 VOUT-.n184 0.314966
R17068 VOUT-.n155 VOUT-.n154 0.3107
R17069 VOUT-.n119 VOUT-.n111 0.306
R17070 VOUT-.n120 VOUT-.n110 0.306
R17071 VOUT-.n121 VOUT-.n109 0.306
R17072 VOUT-.n127 VOUT-.n124 0.2825
R17073 VOUT-.n130 VOUT-.n127 0.2825
R17074 VOUT-.n133 VOUT-.n130 0.2825
R17075 VOUT-.n136 VOUT-.n133 0.2825
R17076 VOUT-.n139 VOUT-.n136 0.2825
R17077 VOUT-.n142 VOUT-.n139 0.2825
R17078 VOUT-.n145 VOUT-.n142 0.2825
R17079 VOUT-.n148 VOUT-.n145 0.2825
R17080 VOUT-.n151 VOUT-.n148 0.2825
R17081 VOUT-.n86 VOUT-.n72 0.2825
R17082 VOUT-.n89 VOUT-.n86 0.2825
R17083 VOUT-.n92 VOUT-.n89 0.2825
R17084 VOUT-.n95 VOUT-.n92 0.2825
R17085 VOUT-.n98 VOUT-.n95 0.2825
R17086 VOUT-.n101 VOUT-.n98 0.2825
R17087 VOUT-.n104 VOUT-.n101 0.2825
R17088 VOUT-.n107 VOUT-.n104 0.2825
R17089 VOUT-.n153 VOUT-.n107 0.2825
R17090 VOUT-.n153 VOUT-.n151 0.2825
R17091 VOUT-.n164 VOUT-.n66 0.2455
R17092 VOUT- VOUT-.n179 0.198417
R17093 VOUT- VOUT-.n198 0.182792
R17094 VOUT-.n156 VOUT-.n155 0.138367
R17095 VOUT-.n190 VOUT-.n184 0.0891864
R17096 VOUT-.n60 VOUT-.n59 0.0577917
R17097 VOUT-.n59 VOUT-.n58 0.0577917
R17098 VOUT-.n58 VOUT-.n21 0.0577917
R17099 VOUT-.n54 VOUT-.n21 0.0577917
R17100 VOUT-.n54 VOUT-.n53 0.0577917
R17101 VOUT-.n53 VOUT-.n52 0.0577917
R17102 VOUT-.n52 VOUT-.n25 0.0577917
R17103 VOUT-.n48 VOUT-.n25 0.0577917
R17104 VOUT-.n61 VOUT-.n18 0.0577917
R17105 VOUT-.n57 VOUT-.n18 0.0577917
R17106 VOUT-.n57 VOUT-.n56 0.0577917
R17107 VOUT-.n56 VOUT-.n55 0.0577917
R17108 VOUT-.n55 VOUT-.n22 0.0577917
R17109 VOUT-.n51 VOUT-.n22 0.0577917
R17110 VOUT-.n51 VOUT-.n50 0.0577917
R17111 VOUT-.n49 VOUT-.n48 0.054517
R17112 VOUT-.n171 VOUT-.n170 0.047375
R17113 VOUT-.n175 VOUT-.n174 0.047375
R17114 VOUT-.n165 VOUT-.n7 0.0421667
R17115 VOUT-.n65 VOUT-.n14 0.0421667
R17116 VOUT-.n197 VOUT-.n196 0.0421667
R17117 VOUT-.n196 VOUT-.n195 0.0421667
R17118 VOUT-.n195 VOUT-.n183 0.0421667
R17119 VOUT-.n191 VOUT-.n183 0.0421667
R17120 VOUT-.n191 VOUT-.n190 0.0421667
R17121 VOUT-.n198 VOUT-.n180 0.0421667
R17122 VOUT-.n194 VOUT-.n180 0.0421667
R17123 VOUT-.n194 VOUT-.n193 0.0421667
R17124 VOUT-.n193 VOUT-.n192 0.0421667
R17125 VOUT-.n15 VOUT-.n14 0.0243161
R17126 VOUT-.n17 VOUT-.n9 0.0243161
R17127 VOUT-.n17 VOUT-.n16 0.0243161
R17128 VOUT-.n15 VOUT-.n11 0.0243161
R17129 VOUT-.n162 VOUT-.n3 0.0217373
R17130 VOUT-.n62 VOUT-.n10 0.0217373
R17131 VOUT-.n16 VOUT-.n10 0.0217373
R17132 VOUT-.n69 VOUT-.n3 0.0217373
R17133 VOUT-.n178 VOUT-.n0 0.0217373
R17134 VOUT-.n175 VOUT-.n0 0.0217373
R17135 VOUT-.n67 VOUT-.n7 0.0217373
R17136 VOUT-.n69 VOUT-.n68 0.0217373
R17137 VOUT-.n12 VOUT-.n9 0.0217373
R17138 VOUT-.n12 VOUT-.n11 0.0217373
R17139 VOUT-.n67 VOUT-.n4 0.0217373
R17140 VOUT-.n68 VOUT-.n4 0.0217373
R17141 VOUT-.n172 VOUT-.n167 0.0217373
R17142 VOUT-.n171 VOUT-.n168 0.0217373
R17143 VOUT-.n174 VOUT-.n168 0.0217373
R17144 VOUT-.n170 VOUT-.n167 0.0217373
R17145 VOUT-.n157 VOUT-.n156 0.0161667
R17146 VOUT-.n160 VOUT-.n157 0.0161667
R17147 VOUT-.n158 VOUT-.n6 0.0161667
R17148 VOUT-.n159 VOUT-.n158 0.0161667
R17149 VOUT-.n159 VOUT-.n70 0.0161667
R17150 VOUT-.n163 VOUT-.n5 0.0134654
R17151 VOUT-.n166 VOUT-.n2 0.0134654
R17152 VOUT-.n164 VOUT-.n163 0.0134654
R17153 VOUT-.n5 VOUT-.n2 0.0134654
R17154 VOUT-.n63 VOUT-.n13 0.0109778
R17155 VOUT-.n66 VOUT-.n8 0.0109778
R17156 VOUT-.n176 VOUT-.n1 0.0109778
R17157 VOUT-.n173 VOUT-.n169 0.0109778
R17158 VOUT-.n64 VOUT-.n63 0.0109778
R17159 VOUT-.n13 VOUT-.n8 0.0109778
R17160 VOUT-.n177 VOUT-.n176 0.0109778
R17161 VOUT-.n169 VOUT-.n1 0.0109778
R17162 VOUT-.n161 VOUT-.n70 0.00872683
R17163 two_stage_opamp_dummy_magic_29_0.cap_res_X two_stage_opamp_dummy_magic_29_0.cap_res_X.t143 49.8942
R17164 two_stage_opamp_dummy_magic_29_0.cap_res_X two_stage_opamp_dummy_magic_29_0.cap_res_X.t75 0.9405
R17165 two_stage_opamp_dummy_magic_29_0.cap_res_X.t119 two_stage_opamp_dummy_magic_29_0.cap_res_X.t17 0.1603
R17166 two_stage_opamp_dummy_magic_29_0.cap_res_X.t141 two_stage_opamp_dummy_magic_29_0.cap_res_X.t44 0.1603
R17167 two_stage_opamp_dummy_magic_29_0.cap_res_X.t124 two_stage_opamp_dummy_magic_29_0.cap_res_X.t22 0.1603
R17168 two_stage_opamp_dummy_magic_29_0.cap_res_X.t87 two_stage_opamp_dummy_magic_29_0.cap_res_X.t127 0.1603
R17169 two_stage_opamp_dummy_magic_29_0.cap_res_X.t106 two_stage_opamp_dummy_magic_29_0.cap_res_X.t5 0.1603
R17170 two_stage_opamp_dummy_magic_29_0.cap_res_X.t71 two_stage_opamp_dummy_magic_29_0.cap_res_X.t107 0.1603
R17171 two_stage_opamp_dummy_magic_29_0.cap_res_X.t33 two_stage_opamp_dummy_magic_29_0.cap_res_X.t73 0.1603
R17172 two_stage_opamp_dummy_magic_29_0.cap_res_X.t26 two_stage_opamp_dummy_magic_29_0.cap_res_X.t51 0.1603
R17173 two_stage_opamp_dummy_magic_29_0.cap_res_X.t142 two_stage_opamp_dummy_magic_29_0.cap_res_X.t120 0.1603
R17174 two_stage_opamp_dummy_magic_29_0.cap_res_X.t67 two_stage_opamp_dummy_magic_29_0.cap_res_X.t93 0.1603
R17175 two_stage_opamp_dummy_magic_29_0.cap_res_X.t45 two_stage_opamp_dummy_magic_29_0.cap_res_X.t18 0.1603
R17176 two_stage_opamp_dummy_magic_29_0.cap_res_X.t103 two_stage_opamp_dummy_magic_29_0.cap_res_X.t130 0.1603
R17177 two_stage_opamp_dummy_magic_29_0.cap_res_X.t85 two_stage_opamp_dummy_magic_29_0.cap_res_X.t60 0.1603
R17178 two_stage_opamp_dummy_magic_29_0.cap_res_X.t2 two_stage_opamp_dummy_magic_29_0.cap_res_X.t29 0.1603
R17179 two_stage_opamp_dummy_magic_29_0.cap_res_X.t50 two_stage_opamp_dummy_magic_29_0.cap_res_X.t23 0.1603
R17180 two_stage_opamp_dummy_magic_29_0.cap_res_X.t108 two_stage_opamp_dummy_magic_29_0.cap_res_X.t135 0.1603
R17181 two_stage_opamp_dummy_magic_29_0.cap_res_X.t92 two_stage_opamp_dummy_magic_29_0.cap_res_X.t64 0.1603
R17182 two_stage_opamp_dummy_magic_29_0.cap_res_X.t9 two_stage_opamp_dummy_magic_29_0.cap_res_X.t35 0.1603
R17183 two_stage_opamp_dummy_magic_29_0.cap_res_X.t111 two_stage_opamp_dummy_magic_29_0.cap_res_X.t21 0.1603
R17184 two_stage_opamp_dummy_magic_29_0.cap_res_X.t41 two_stage_opamp_dummy_magic_29_0.cap_res_X.t131 0.1603
R17185 two_stage_opamp_dummy_magic_29_0.cap_res_X.t79 two_stage_opamp_dummy_magic_29_0.cap_res_X.t129 0.1603
R17186 two_stage_opamp_dummy_magic_29_0.cap_res_X.t4 two_stage_opamp_dummy_magic_29_0.cap_res_X.t97 0.1603
R17187 two_stage_opamp_dummy_magic_29_0.cap_res_X.t116 two_stage_opamp_dummy_magic_29_0.cap_res_X.t28 0.1603
R17188 two_stage_opamp_dummy_magic_29_0.cap_res_X.t49 two_stage_opamp_dummy_magic_29_0.cap_res_X.t137 0.1603
R17189 two_stage_opamp_dummy_magic_29_0.cap_res_X.t13 two_stage_opamp_dummy_magic_29_0.cap_res_X.t69 0.1603
R17190 two_stage_opamp_dummy_magic_29_0.cap_res_X.t90 two_stage_opamp_dummy_magic_29_0.cap_res_X.t38 0.1603
R17191 two_stage_opamp_dummy_magic_29_0.cap_res_X.t123 two_stage_opamp_dummy_magic_29_0.cap_res_X.t34 0.1603
R17192 two_stage_opamp_dummy_magic_29_0.cap_res_X.t54 two_stage_opamp_dummy_magic_29_0.cap_res_X.t140 0.1603
R17193 two_stage_opamp_dummy_magic_29_0.cap_res_X.t19 two_stage_opamp_dummy_magic_29_0.cap_res_X.t74 0.1603
R17194 two_stage_opamp_dummy_magic_29_0.cap_res_X.t94 two_stage_opamp_dummy_magic_29_0.cap_res_X.t40 0.1603
R17195 two_stage_opamp_dummy_magic_29_0.cap_res_X.t61 two_stage_opamp_dummy_magic_29_0.cap_res_X.t112 0.1603
R17196 two_stage_opamp_dummy_magic_29_0.cap_res_X.t133 two_stage_opamp_dummy_magic_29_0.cap_res_X.t82 0.1603
R17197 two_stage_opamp_dummy_magic_29_0.cap_res_X.t100 two_stage_opamp_dummy_magic_29_0.cap_res_X.t11 0.1603
R17198 two_stage_opamp_dummy_magic_29_0.cap_res_X.t31 two_stage_opamp_dummy_magic_29_0.cap_res_X.t121 0.1603
R17199 two_stage_opamp_dummy_magic_29_0.cap_res_X.t68 two_stage_opamp_dummy_magic_29_0.cap_res_X.t117 0.1603
R17200 two_stage_opamp_dummy_magic_29_0.cap_res_X.t138 two_stage_opamp_dummy_magic_29_0.cap_res_X.t86 0.1603
R17201 two_stage_opamp_dummy_magic_29_0.cap_res_X.t104 two_stage_opamp_dummy_magic_29_0.cap_res_X.t15 0.1603
R17202 two_stage_opamp_dummy_magic_29_0.cap_res_X.t39 two_stage_opamp_dummy_magic_29_0.cap_res_X.t126 0.1603
R17203 two_stage_opamp_dummy_magic_29_0.cap_res_X.t3 two_stage_opamp_dummy_magic_29_0.cap_res_X.t57 0.1603
R17204 two_stage_opamp_dummy_magic_29_0.cap_res_X.t78 two_stage_opamp_dummy_magic_29_0.cap_res_X.t24 0.1603
R17205 two_stage_opamp_dummy_magic_29_0.cap_res_X.t109 two_stage_opamp_dummy_magic_29_0.cap_res_X.t20 0.1603
R17206 two_stage_opamp_dummy_magic_29_0.cap_res_X.t42 two_stage_opamp_dummy_magic_29_0.cap_res_X.t132 0.1603
R17207 two_stage_opamp_dummy_magic_29_0.cap_res_X.t70 two_stage_opamp_dummy_magic_29_0.cap_res_X.t53 0.1603
R17208 two_stage_opamp_dummy_magic_29_0.cap_res_X.t14 two_stage_opamp_dummy_magic_29_0.cap_res_X.t7 0.1603
R17209 two_stage_opamp_dummy_magic_29_0.cap_res_X.t95 two_stage_opamp_dummy_magic_29_0.cap_res_X.t89 0.1603
R17210 two_stage_opamp_dummy_magic_29_0.cap_res_X.t59 two_stage_opamp_dummy_magic_29_0.cap_res_X.t139 0.1603
R17211 two_stage_opamp_dummy_magic_29_0.cap_res_X.t6 two_stage_opamp_dummy_magic_29_0.cap_res_X.t96 0.1603
R17212 two_stage_opamp_dummy_magic_29_0.cap_res_X.t113 two_stage_opamp_dummy_magic_29_0.cap_res_X.t1 0.1603
R17213 two_stage_opamp_dummy_magic_29_0.cap_res_X.t80 two_stage_opamp_dummy_magic_29_0.cap_res_X.t56 0.1603
R17214 two_stage_opamp_dummy_magic_29_0.cap_res_X.t46 two_stage_opamp_dummy_magic_29_0.cap_res_X.t105 0.1603
R17215 two_stage_opamp_dummy_magic_29_0.cap_res_X.t134 two_stage_opamp_dummy_magic_29_0.cap_res_X.t65 0.1603
R17216 two_stage_opamp_dummy_magic_29_0.cap_res_X.t99 two_stage_opamp_dummy_magic_29_0.cap_res_X.t114 0.1603
R17217 two_stage_opamp_dummy_magic_29_0.cap_res_X.t62 two_stage_opamp_dummy_magic_29_0.cap_res_X.t27 0.1603
R17218 two_stage_opamp_dummy_magic_29_0.cap_res_X.t10 two_stage_opamp_dummy_magic_29_0.cap_res_X.t125 0.1603
R17219 two_stage_opamp_dummy_magic_29_0.cap_res_X.t83 two_stage_opamp_dummy_magic_29_0.cap_res_X.t30 0.1603
R17220 two_stage_opamp_dummy_magic_29_0.cap_res_X.t88 two_stage_opamp_dummy_magic_29_0.cap_res_X.t48 0.1603
R17221 two_stage_opamp_dummy_magic_29_0.cap_res_X.t81 two_stage_opamp_dummy_magic_29_0.cap_res_X.t101 0.1603
R17222 two_stage_opamp_dummy_magic_29_0.cap_res_X.t16 two_stage_opamp_dummy_magic_29_0.cap_res_X.t58 0.1603
R17223 two_stage_opamp_dummy_magic_29_0.cap_res_X.t118 two_stage_opamp_dummy_magic_29_0.cap_res_X.t16 0.1603
R17224 two_stage_opamp_dummy_magic_29_0.cap_res_X.t55 two_stage_opamp_dummy_magic_29_0.cap_res_X.t98 0.1603
R17225 two_stage_opamp_dummy_magic_29_0.cap_res_X.t12 two_stage_opamp_dummy_magic_29_0.cap_res_X.t55 0.1603
R17226 two_stage_opamp_dummy_magic_29_0.cap_res_X.t36 two_stage_opamp_dummy_magic_29_0.cap_res_X.t136 0.1603
R17227 two_stage_opamp_dummy_magic_29_0.cap_res_X.t75 two_stage_opamp_dummy_magic_29_0.cap_res_X.t36 0.1603
R17228 two_stage_opamp_dummy_magic_29_0.cap_res_X.t115 two_stage_opamp_dummy_magic_29_0.cap_res_X.n11 0.159278
R17229 two_stage_opamp_dummy_magic_29_0.cap_res_X.t77 two_stage_opamp_dummy_magic_29_0.cap_res_X.n12 0.159278
R17230 two_stage_opamp_dummy_magic_29_0.cap_res_X.t110 two_stage_opamp_dummy_magic_29_0.cap_res_X.n13 0.159278
R17231 two_stage_opamp_dummy_magic_29_0.cap_res_X.t72 two_stage_opamp_dummy_magic_29_0.cap_res_X.n14 0.159278
R17232 two_stage_opamp_dummy_magic_29_0.cap_res_X.t32 two_stage_opamp_dummy_magic_29_0.cap_res_X.n15 0.159278
R17233 two_stage_opamp_dummy_magic_29_0.cap_res_X.t66 two_stage_opamp_dummy_magic_29_0.cap_res_X.n16 0.159278
R17234 two_stage_opamp_dummy_magic_29_0.cap_res_X.t25 two_stage_opamp_dummy_magic_29_0.cap_res_X.n17 0.159278
R17235 two_stage_opamp_dummy_magic_29_0.cap_res_X.t128 two_stage_opamp_dummy_magic_29_0.cap_res_X.n18 0.159278
R17236 two_stage_opamp_dummy_magic_29_0.cap_res_X.t91 two_stage_opamp_dummy_magic_29_0.cap_res_X.n19 0.159278
R17237 two_stage_opamp_dummy_magic_29_0.cap_res_X.t122 two_stage_opamp_dummy_magic_29_0.cap_res_X.n20 0.159278
R17238 two_stage_opamp_dummy_magic_29_0.cap_res_X.t84 two_stage_opamp_dummy_magic_29_0.cap_res_X.n21 0.159278
R17239 two_stage_opamp_dummy_magic_29_0.cap_res_X.t43 two_stage_opamp_dummy_magic_29_0.cap_res_X.n22 0.159278
R17240 two_stage_opamp_dummy_magic_29_0.cap_res_X.t76 two_stage_opamp_dummy_magic_29_0.cap_res_X.n23 0.159278
R17241 two_stage_opamp_dummy_magic_29_0.cap_res_X.t52 two_stage_opamp_dummy_magic_29_0.cap_res_X.n24 0.159278
R17242 two_stage_opamp_dummy_magic_29_0.cap_res_X.t8 two_stage_opamp_dummy_magic_29_0.cap_res_X.n25 0.159278
R17243 two_stage_opamp_dummy_magic_29_0.cap_res_X.t47 two_stage_opamp_dummy_magic_29_0.cap_res_X.n26 0.159278
R17244 two_stage_opamp_dummy_magic_29_0.cap_res_X.t0 two_stage_opamp_dummy_magic_29_0.cap_res_X.n27 0.159278
R17245 two_stage_opamp_dummy_magic_29_0.cap_res_X.t102 two_stage_opamp_dummy_magic_29_0.cap_res_X.n28 0.159278
R17246 two_stage_opamp_dummy_magic_29_0.cap_res_X.t63 two_stage_opamp_dummy_magic_29_0.cap_res_X.n29 0.159278
R17247 two_stage_opamp_dummy_magic_29_0.cap_res_X.n30 two_stage_opamp_dummy_magic_29_0.cap_res_X.t26 0.1368
R17248 two_stage_opamp_dummy_magic_29_0.cap_res_X.n29 two_stage_opamp_dummy_magic_29_0.cap_res_X.t142 0.1368
R17249 two_stage_opamp_dummy_magic_29_0.cap_res_X.n29 two_stage_opamp_dummy_magic_29_0.cap_res_X.t67 0.1368
R17250 two_stage_opamp_dummy_magic_29_0.cap_res_X.n28 two_stage_opamp_dummy_magic_29_0.cap_res_X.t45 0.1368
R17251 two_stage_opamp_dummy_magic_29_0.cap_res_X.n28 two_stage_opamp_dummy_magic_29_0.cap_res_X.t103 0.1368
R17252 two_stage_opamp_dummy_magic_29_0.cap_res_X.n27 two_stage_opamp_dummy_magic_29_0.cap_res_X.t85 0.1368
R17253 two_stage_opamp_dummy_magic_29_0.cap_res_X.n27 two_stage_opamp_dummy_magic_29_0.cap_res_X.t2 0.1368
R17254 two_stage_opamp_dummy_magic_29_0.cap_res_X.n26 two_stage_opamp_dummy_magic_29_0.cap_res_X.t50 0.1368
R17255 two_stage_opamp_dummy_magic_29_0.cap_res_X.n26 two_stage_opamp_dummy_magic_29_0.cap_res_X.t108 0.1368
R17256 two_stage_opamp_dummy_magic_29_0.cap_res_X.n25 two_stage_opamp_dummy_magic_29_0.cap_res_X.t92 0.1368
R17257 two_stage_opamp_dummy_magic_29_0.cap_res_X.n25 two_stage_opamp_dummy_magic_29_0.cap_res_X.t9 0.1368
R17258 two_stage_opamp_dummy_magic_29_0.cap_res_X.n24 two_stage_opamp_dummy_magic_29_0.cap_res_X.t111 0.1368
R17259 two_stage_opamp_dummy_magic_29_0.cap_res_X.n24 two_stage_opamp_dummy_magic_29_0.cap_res_X.t41 0.1368
R17260 two_stage_opamp_dummy_magic_29_0.cap_res_X.n23 two_stage_opamp_dummy_magic_29_0.cap_res_X.t79 0.1368
R17261 two_stage_opamp_dummy_magic_29_0.cap_res_X.n23 two_stage_opamp_dummy_magic_29_0.cap_res_X.t4 0.1368
R17262 two_stage_opamp_dummy_magic_29_0.cap_res_X.n22 two_stage_opamp_dummy_magic_29_0.cap_res_X.t116 0.1368
R17263 two_stage_opamp_dummy_magic_29_0.cap_res_X.n22 two_stage_opamp_dummy_magic_29_0.cap_res_X.t49 0.1368
R17264 two_stage_opamp_dummy_magic_29_0.cap_res_X.n21 two_stage_opamp_dummy_magic_29_0.cap_res_X.t13 0.1368
R17265 two_stage_opamp_dummy_magic_29_0.cap_res_X.n21 two_stage_opamp_dummy_magic_29_0.cap_res_X.t90 0.1368
R17266 two_stage_opamp_dummy_magic_29_0.cap_res_X.n20 two_stage_opamp_dummy_magic_29_0.cap_res_X.t123 0.1368
R17267 two_stage_opamp_dummy_magic_29_0.cap_res_X.n20 two_stage_opamp_dummy_magic_29_0.cap_res_X.t54 0.1368
R17268 two_stage_opamp_dummy_magic_29_0.cap_res_X.n19 two_stage_opamp_dummy_magic_29_0.cap_res_X.t19 0.1368
R17269 two_stage_opamp_dummy_magic_29_0.cap_res_X.n19 two_stage_opamp_dummy_magic_29_0.cap_res_X.t94 0.1368
R17270 two_stage_opamp_dummy_magic_29_0.cap_res_X.n18 two_stage_opamp_dummy_magic_29_0.cap_res_X.t61 0.1368
R17271 two_stage_opamp_dummy_magic_29_0.cap_res_X.n18 two_stage_opamp_dummy_magic_29_0.cap_res_X.t133 0.1368
R17272 two_stage_opamp_dummy_magic_29_0.cap_res_X.n17 two_stage_opamp_dummy_magic_29_0.cap_res_X.t100 0.1368
R17273 two_stage_opamp_dummy_magic_29_0.cap_res_X.n17 two_stage_opamp_dummy_magic_29_0.cap_res_X.t31 0.1368
R17274 two_stage_opamp_dummy_magic_29_0.cap_res_X.n16 two_stage_opamp_dummy_magic_29_0.cap_res_X.t68 0.1368
R17275 two_stage_opamp_dummy_magic_29_0.cap_res_X.n16 two_stage_opamp_dummy_magic_29_0.cap_res_X.t138 0.1368
R17276 two_stage_opamp_dummy_magic_29_0.cap_res_X.n15 two_stage_opamp_dummy_magic_29_0.cap_res_X.t104 0.1368
R17277 two_stage_opamp_dummy_magic_29_0.cap_res_X.n15 two_stage_opamp_dummy_magic_29_0.cap_res_X.t39 0.1368
R17278 two_stage_opamp_dummy_magic_29_0.cap_res_X.n14 two_stage_opamp_dummy_magic_29_0.cap_res_X.t3 0.1368
R17279 two_stage_opamp_dummy_magic_29_0.cap_res_X.n14 two_stage_opamp_dummy_magic_29_0.cap_res_X.t78 0.1368
R17280 two_stage_opamp_dummy_magic_29_0.cap_res_X.n13 two_stage_opamp_dummy_magic_29_0.cap_res_X.t109 0.1368
R17281 two_stage_opamp_dummy_magic_29_0.cap_res_X.n13 two_stage_opamp_dummy_magic_29_0.cap_res_X.t42 0.1368
R17282 two_stage_opamp_dummy_magic_29_0.cap_res_X.n12 two_stage_opamp_dummy_magic_29_0.cap_res_X.t83 0.1368
R17283 two_stage_opamp_dummy_magic_29_0.cap_res_X.n11 two_stage_opamp_dummy_magic_29_0.cap_res_X.t88 0.1368
R17284 two_stage_opamp_dummy_magic_29_0.cap_res_X.t101 two_stage_opamp_dummy_magic_29_0.cap_res_X.n30 0.1368
R17285 two_stage_opamp_dummy_magic_29_0.cap_res_X.n31 two_stage_opamp_dummy_magic_29_0.cap_res_X.t81 0.1368
R17286 two_stage_opamp_dummy_magic_29_0.cap_res_X.n33 two_stage_opamp_dummy_magic_29_0.cap_res_X.t119 0.114322
R17287 two_stage_opamp_dummy_magic_29_0.cap_res_X.n0 two_stage_opamp_dummy_magic_29_0.cap_res_X.t70 0.114322
R17288 two_stage_opamp_dummy_magic_29_0.cap_res_X.n34 two_stage_opamp_dummy_magic_29_0.cap_res_X.n33 0.1133
R17289 two_stage_opamp_dummy_magic_29_0.cap_res_X.n35 two_stage_opamp_dummy_magic_29_0.cap_res_X.n34 0.1133
R17290 two_stage_opamp_dummy_magic_29_0.cap_res_X.n36 two_stage_opamp_dummy_magic_29_0.cap_res_X.n35 0.1133
R17291 two_stage_opamp_dummy_magic_29_0.cap_res_X.n37 two_stage_opamp_dummy_magic_29_0.cap_res_X.n36 0.1133
R17292 two_stage_opamp_dummy_magic_29_0.cap_res_X.n38 two_stage_opamp_dummy_magic_29_0.cap_res_X.n37 0.1133
R17293 two_stage_opamp_dummy_magic_29_0.cap_res_X.n1 two_stage_opamp_dummy_magic_29_0.cap_res_X.n0 0.1133
R17294 two_stage_opamp_dummy_magic_29_0.cap_res_X.n2 two_stage_opamp_dummy_magic_29_0.cap_res_X.n1 0.1133
R17295 two_stage_opamp_dummy_magic_29_0.cap_res_X.n3 two_stage_opamp_dummy_magic_29_0.cap_res_X.n2 0.1133
R17296 two_stage_opamp_dummy_magic_29_0.cap_res_X.n4 two_stage_opamp_dummy_magic_29_0.cap_res_X.n3 0.1133
R17297 two_stage_opamp_dummy_magic_29_0.cap_res_X.n5 two_stage_opamp_dummy_magic_29_0.cap_res_X.n4 0.1133
R17298 two_stage_opamp_dummy_magic_29_0.cap_res_X.n6 two_stage_opamp_dummy_magic_29_0.cap_res_X.n5 0.1133
R17299 two_stage_opamp_dummy_magic_29_0.cap_res_X.n7 two_stage_opamp_dummy_magic_29_0.cap_res_X.n6 0.1133
R17300 two_stage_opamp_dummy_magic_29_0.cap_res_X.n8 two_stage_opamp_dummy_magic_29_0.cap_res_X.n7 0.1133
R17301 two_stage_opamp_dummy_magic_29_0.cap_res_X.n9 two_stage_opamp_dummy_magic_29_0.cap_res_X.n8 0.1133
R17302 two_stage_opamp_dummy_magic_29_0.cap_res_X.n10 two_stage_opamp_dummy_magic_29_0.cap_res_X.n9 0.1133
R17303 two_stage_opamp_dummy_magic_29_0.cap_res_X.n12 two_stage_opamp_dummy_magic_29_0.cap_res_X.n10 0.1133
R17304 two_stage_opamp_dummy_magic_29_0.cap_res_X.n32 two_stage_opamp_dummy_magic_29_0.cap_res_X.n31 0.1133
R17305 two_stage_opamp_dummy_magic_29_0.cap_res_X.n39 two_stage_opamp_dummy_magic_29_0.cap_res_X.n32 0.1133
R17306 two_stage_opamp_dummy_magic_29_0.cap_res_X.n39 two_stage_opamp_dummy_magic_29_0.cap_res_X.n38 0.1133
R17307 two_stage_opamp_dummy_magic_29_0.cap_res_X.n33 two_stage_opamp_dummy_magic_29_0.cap_res_X.t141 0.00152174
R17308 two_stage_opamp_dummy_magic_29_0.cap_res_X.n34 two_stage_opamp_dummy_magic_29_0.cap_res_X.t124 0.00152174
R17309 two_stage_opamp_dummy_magic_29_0.cap_res_X.n35 two_stage_opamp_dummy_magic_29_0.cap_res_X.t87 0.00152174
R17310 two_stage_opamp_dummy_magic_29_0.cap_res_X.n36 two_stage_opamp_dummy_magic_29_0.cap_res_X.t106 0.00152174
R17311 two_stage_opamp_dummy_magic_29_0.cap_res_X.n37 two_stage_opamp_dummy_magic_29_0.cap_res_X.t71 0.00152174
R17312 two_stage_opamp_dummy_magic_29_0.cap_res_X.n38 two_stage_opamp_dummy_magic_29_0.cap_res_X.t33 0.00152174
R17313 two_stage_opamp_dummy_magic_29_0.cap_res_X.n0 two_stage_opamp_dummy_magic_29_0.cap_res_X.t14 0.00152174
R17314 two_stage_opamp_dummy_magic_29_0.cap_res_X.n1 two_stage_opamp_dummy_magic_29_0.cap_res_X.t95 0.00152174
R17315 two_stage_opamp_dummy_magic_29_0.cap_res_X.n2 two_stage_opamp_dummy_magic_29_0.cap_res_X.t59 0.00152174
R17316 two_stage_opamp_dummy_magic_29_0.cap_res_X.n3 two_stage_opamp_dummy_magic_29_0.cap_res_X.t6 0.00152174
R17317 two_stage_opamp_dummy_magic_29_0.cap_res_X.n4 two_stage_opamp_dummy_magic_29_0.cap_res_X.t113 0.00152174
R17318 two_stage_opamp_dummy_magic_29_0.cap_res_X.n5 two_stage_opamp_dummy_magic_29_0.cap_res_X.t80 0.00152174
R17319 two_stage_opamp_dummy_magic_29_0.cap_res_X.n6 two_stage_opamp_dummy_magic_29_0.cap_res_X.t46 0.00152174
R17320 two_stage_opamp_dummy_magic_29_0.cap_res_X.n7 two_stage_opamp_dummy_magic_29_0.cap_res_X.t134 0.00152174
R17321 two_stage_opamp_dummy_magic_29_0.cap_res_X.n8 two_stage_opamp_dummy_magic_29_0.cap_res_X.t99 0.00152174
R17322 two_stage_opamp_dummy_magic_29_0.cap_res_X.n9 two_stage_opamp_dummy_magic_29_0.cap_res_X.t62 0.00152174
R17323 two_stage_opamp_dummy_magic_29_0.cap_res_X.n10 two_stage_opamp_dummy_magic_29_0.cap_res_X.t10 0.00152174
R17324 two_stage_opamp_dummy_magic_29_0.cap_res_X.n11 two_stage_opamp_dummy_magic_29_0.cap_res_X.t37 0.00152174
R17325 two_stage_opamp_dummy_magic_29_0.cap_res_X.n12 two_stage_opamp_dummy_magic_29_0.cap_res_X.t115 0.00152174
R17326 two_stage_opamp_dummy_magic_29_0.cap_res_X.n13 two_stage_opamp_dummy_magic_29_0.cap_res_X.t77 0.00152174
R17327 two_stage_opamp_dummy_magic_29_0.cap_res_X.n14 two_stage_opamp_dummy_magic_29_0.cap_res_X.t110 0.00152174
R17328 two_stage_opamp_dummy_magic_29_0.cap_res_X.n15 two_stage_opamp_dummy_magic_29_0.cap_res_X.t72 0.00152174
R17329 two_stage_opamp_dummy_magic_29_0.cap_res_X.n16 two_stage_opamp_dummy_magic_29_0.cap_res_X.t32 0.00152174
R17330 two_stage_opamp_dummy_magic_29_0.cap_res_X.n17 two_stage_opamp_dummy_magic_29_0.cap_res_X.t66 0.00152174
R17331 two_stage_opamp_dummy_magic_29_0.cap_res_X.n18 two_stage_opamp_dummy_magic_29_0.cap_res_X.t25 0.00152174
R17332 two_stage_opamp_dummy_magic_29_0.cap_res_X.n19 two_stage_opamp_dummy_magic_29_0.cap_res_X.t128 0.00152174
R17333 two_stage_opamp_dummy_magic_29_0.cap_res_X.n20 two_stage_opamp_dummy_magic_29_0.cap_res_X.t91 0.00152174
R17334 two_stage_opamp_dummy_magic_29_0.cap_res_X.n21 two_stage_opamp_dummy_magic_29_0.cap_res_X.t122 0.00152174
R17335 two_stage_opamp_dummy_magic_29_0.cap_res_X.n22 two_stage_opamp_dummy_magic_29_0.cap_res_X.t84 0.00152174
R17336 two_stage_opamp_dummy_magic_29_0.cap_res_X.n23 two_stage_opamp_dummy_magic_29_0.cap_res_X.t43 0.00152174
R17337 two_stage_opamp_dummy_magic_29_0.cap_res_X.n24 two_stage_opamp_dummy_magic_29_0.cap_res_X.t76 0.00152174
R17338 two_stage_opamp_dummy_magic_29_0.cap_res_X.n25 two_stage_opamp_dummy_magic_29_0.cap_res_X.t52 0.00152174
R17339 two_stage_opamp_dummy_magic_29_0.cap_res_X.n26 two_stage_opamp_dummy_magic_29_0.cap_res_X.t8 0.00152174
R17340 two_stage_opamp_dummy_magic_29_0.cap_res_X.n27 two_stage_opamp_dummy_magic_29_0.cap_res_X.t47 0.00152174
R17341 two_stage_opamp_dummy_magic_29_0.cap_res_X.n28 two_stage_opamp_dummy_magic_29_0.cap_res_X.t0 0.00152174
R17342 two_stage_opamp_dummy_magic_29_0.cap_res_X.n29 two_stage_opamp_dummy_magic_29_0.cap_res_X.t102 0.00152174
R17343 two_stage_opamp_dummy_magic_29_0.cap_res_X.n30 two_stage_opamp_dummy_magic_29_0.cap_res_X.t63 0.00152174
R17344 two_stage_opamp_dummy_magic_29_0.cap_res_X.n31 two_stage_opamp_dummy_magic_29_0.cap_res_X.t118 0.00152174
R17345 two_stage_opamp_dummy_magic_29_0.cap_res_X.n32 two_stage_opamp_dummy_magic_29_0.cap_res_X.t12 0.00152174
R17346 two_stage_opamp_dummy_magic_29_0.cap_res_X.t136 two_stage_opamp_dummy_magic_29_0.cap_res_X.n39 0.00152174
R17347 two_stage_opamp_dummy_magic_29_0.cap_res_Y two_stage_opamp_dummy_magic_29_0.cap_res_Y.t3 49.895
R17348 two_stage_opamp_dummy_magic_29_0.cap_res_Y two_stage_opamp_dummy_magic_29_0.cap_res_Y.t26 0.9405
R17349 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t46 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t60 0.1603
R17350 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t1 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t138 0.1603
R17351 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t65 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t15 0.1603
R17352 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t108 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t79 0.1603
R17353 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t77 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t68 0.1603
R17354 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t84 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t28 0.1603
R17355 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t88 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t81 0.1603
R17356 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t57 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t21 0.1603
R17357 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t78 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t0 0.1603
R17358 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t40 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t83 0.1603
R17359 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t56 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t89 0.1603
R17360 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t17 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t110 0.1603
R17361 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t29 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t43 0.1603
R17362 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t115 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t48 0.1603
R17363 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t71 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t129 0.1603
R17364 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t14 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t113 0.1603
R17365 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t112 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t38 0.1603
R17366 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t18 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t126 0.1603
R17367 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t87 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t61 0.1603
R17368 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t64 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t59 0.1603
R17369 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t58 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t51 0.1603
R17370 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t76 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t63 0.1603
R17371 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t62 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t116 0.1603
R17372 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t55 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t142 0.1603
R17373 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t69 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t120 0.1603
R17374 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t24 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t130 0.1603
R17375 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t107 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t70 0.1603
R17376 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t135 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t99 0.1603
R17377 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t75 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t140 0.1603
R17378 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t33 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t133 0.1603
R17379 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t132 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t6 0.1603
R17380 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t103 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t23 0.1603
R17381 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t22 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t11 0.1603
R17382 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t12 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t34 0.1603
R17383 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t35 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t42 0.1603
R17384 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t93 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t44 0.1603
R17385 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t27 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t122 0.1603
R17386 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t123 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t136 0.1603
R17387 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t105 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t67 0.1603
R17388 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t30 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t36 0.1603
R17389 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t119 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t49 0.1603
R17390 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t92 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t47 0.1603
R17391 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t8 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t74 0.1603
R17392 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t73 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t86 0.1603
R17393 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t66 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t53 0.1603
R17394 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t39 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t25 0.1603
R17395 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t37 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t50 0.1603
R17396 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t41 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t137 0.1603
R17397 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t96 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t125 0.1603
R17398 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t10 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t31 0.1603
R17399 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t114 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t118 0.1603
R17400 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t100 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t114 0.1603
R17401 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t85 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t2 0.1603
R17402 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t109 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t85 0.1603
R17403 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t19 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t80 0.1603
R17404 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t106 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t97 0.1603
R17405 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t20 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t91 0.1603
R17406 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t82 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t13 0.1603
R17407 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t32 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t102 0.1603
R17408 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t128 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t124 0.1603
R17409 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t139 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t4 0.1603
R17410 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t54 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t5 0.1603
R17411 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t26 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t54 0.1603
R17412 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t45 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n17 0.159278
R17413 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t111 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n18 0.159278
R17414 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t72 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n19 0.159278
R17415 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t52 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n20 0.159278
R17416 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t98 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n21 0.159278
R17417 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t131 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n22 0.159278
R17418 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t143 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n23 0.159278
R17419 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t16 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n24 0.159278
R17420 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t90 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n25 0.159278
R17421 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t127 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n26 0.159278
R17422 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t134 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n27 0.159278
R17423 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t94 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n28 0.159278
R17424 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t9 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n29 0.159278
R17425 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t7 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n30 0.159278
R17426 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t141 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n31 0.159278
R17427 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t95 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n32 0.159278
R17428 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t121 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n33 0.159278
R17429 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t117 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n34 0.159278
R17430 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t104 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n35 0.159278
R17431 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n36 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t46 0.1368
R17432 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t1 0.1368
R17433 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t65 0.1368
R17434 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t108 0.1368
R17435 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t77 0.1368
R17436 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t84 0.1368
R17437 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t88 0.1368
R17438 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t57 0.1368
R17439 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t78 0.1368
R17440 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t40 0.1368
R17441 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t56 0.1368
R17442 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t17 0.1368
R17443 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t29 0.1368
R17444 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t115 0.1368
R17445 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t71 0.1368
R17446 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t14 0.1368
R17447 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t112 0.1368
R17448 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t18 0.1368
R17449 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t87 0.1368
R17450 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t64 0.1368
R17451 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t58 0.1368
R17452 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t76 0.1368
R17453 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t62 0.1368
R17454 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t55 0.1368
R17455 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t69 0.1368
R17456 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t24 0.1368
R17457 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t107 0.1368
R17458 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t135 0.1368
R17459 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t75 0.1368
R17460 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t33 0.1368
R17461 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t132 0.1368
R17462 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t103 0.1368
R17463 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t22 0.1368
R17464 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t12 0.1368
R17465 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t35 0.1368
R17466 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t93 0.1368
R17467 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t96 0.1368
R17468 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t31 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n36 0.1368
R17469 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n37 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t10 0.1368
R17470 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t27 0.114322
R17471 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t19 0.114322
R17472 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n6 0.1133
R17473 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n7 0.1133
R17474 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n8 0.1133
R17475 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n9 0.1133
R17476 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n10 0.1133
R17477 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n11 0.1133
R17478 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n12 0.1133
R17479 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n13 0.1133
R17480 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n14 0.1133
R17481 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n15 0.1133
R17482 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n16 0.1133
R17483 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n38 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n37 0.1133
R17484 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n0 0.1133
R17485 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n1 0.1133
R17486 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n2 0.1133
R17487 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n3 0.1133
R17488 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n4 0.1133
R17489 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n39 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n5 0.1133
R17490 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n39 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n38 0.1133
R17491 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n6 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t123 0.00152174
R17492 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n7 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t105 0.00152174
R17493 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n8 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t30 0.00152174
R17494 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n9 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t119 0.00152174
R17495 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n10 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t92 0.00152174
R17496 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n11 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t8 0.00152174
R17497 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n12 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t73 0.00152174
R17498 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n13 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t66 0.00152174
R17499 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n14 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t39 0.00152174
R17500 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n15 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t37 0.00152174
R17501 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n16 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t41 0.00152174
R17502 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n17 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t101 0.00152174
R17503 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n18 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t45 0.00152174
R17504 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n19 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t111 0.00152174
R17505 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n20 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t72 0.00152174
R17506 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n21 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t52 0.00152174
R17507 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n22 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t98 0.00152174
R17508 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n23 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t131 0.00152174
R17509 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n24 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t143 0.00152174
R17510 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n25 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t16 0.00152174
R17511 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n26 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t90 0.00152174
R17512 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n27 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t127 0.00152174
R17513 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n28 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t134 0.00152174
R17514 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n29 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t94 0.00152174
R17515 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n30 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t9 0.00152174
R17516 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n31 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t7 0.00152174
R17517 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n32 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t141 0.00152174
R17518 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n33 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t95 0.00152174
R17519 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n34 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t121 0.00152174
R17520 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n35 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t117 0.00152174
R17521 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n36 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t104 0.00152174
R17522 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n37 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t100 0.00152174
R17523 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n38 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t109 0.00152174
R17524 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n0 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t106 0.00152174
R17525 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n1 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t20 0.00152174
R17526 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n2 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t82 0.00152174
R17527 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n3 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t32 0.00152174
R17528 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n4 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t128 0.00152174
R17529 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n5 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t139 0.00152174
R17530 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t5 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n39 0.00152174
R17531 VOUT+.n197 VOUT+.t12 110.386
R17532 VOUT+.n47 VOUT+.n46 34.9935
R17533 VOUT+.n45 VOUT+.n44 34.9935
R17534 VOUT+.n59 VOUT+.n58 34.9935
R17535 VOUT+.n55 VOUT+.n54 34.9935
R17536 VOUT+.n52 VOUT+.n51 34.9935
R17537 VOUT+.n49 VOUT+.n48 34.9935
R17538 VOUT+.n2 VOUT+.n1 9.73997
R17539 VOUT+.n6 VOUT+.n5 9.73997
R17540 VOUT+.n9 VOUT+.n8 9.73997
R17541 VOUT+.n7 VOUT+.n6 6.64633
R17542 VOUT+.n7 VOUT+.n2 6.64633
R17543 VOUT+.n46 VOUT+.t9 6.56717
R17544 VOUT+.n46 VOUT+.t16 6.56717
R17545 VOUT+.n44 VOUT+.t15 6.56717
R17546 VOUT+.n44 VOUT+.t5 6.56717
R17547 VOUT+.n58 VOUT+.t8 6.56717
R17548 VOUT+.n58 VOUT+.t2 6.56717
R17549 VOUT+.n54 VOUT+.t7 6.56717
R17550 VOUT+.n54 VOUT+.t1 6.56717
R17551 VOUT+.n51 VOUT+.t6 6.56717
R17552 VOUT+.n51 VOUT+.t4 6.56717
R17553 VOUT+.n48 VOUT+.t10 6.56717
R17554 VOUT+.n48 VOUT+.t3 6.56717
R17555 VOUT+.n57 VOUT+.n45 6.3755
R17556 VOUT+.n50 VOUT+.n47 6.3755
R17557 VOUT+.n9 VOUT+.n7 6.02133
R17558 VOUT+.n59 VOUT+.n57 5.813
R17559 VOUT+.n56 VOUT+.n55 5.813
R17560 VOUT+.n53 VOUT+.n52 5.813
R17561 VOUT+.n50 VOUT+.n49 5.813
R17562 VOUT+.n60 VOUT+.n36 5.063
R17563 VOUT+.n63 VOUT+.n43 5.063
R17564 VOUT+.n134 VOUT+.t34 4.8295
R17565 VOUT+.n135 VOUT+.t19 4.8295
R17566 VOUT+.n136 VOUT+.t54 4.8295
R17567 VOUT+.n149 VOUT+.t70 4.8295
R17568 VOUT+.n151 VOUT+.t37 4.8295
R17569 VOUT+.n152 VOUT+.t28 4.8295
R17570 VOUT+.n154 VOUT+.t152 4.8295
R17571 VOUT+.n155 VOUT+.t139 4.8295
R17572 VOUT+.n157 VOUT+.t111 4.8295
R17573 VOUT+.n158 VOUT+.t92 4.8295
R17574 VOUT+.n160 VOUT+.t144 4.8295
R17575 VOUT+.n161 VOUT+.t131 4.8295
R17576 VOUT+.n163 VOUT+.t103 4.8295
R17577 VOUT+.n164 VOUT+.t85 4.8295
R17578 VOUT+.n166 VOUT+.t125 4.8295
R17579 VOUT+.n167 VOUT+.t96 4.8295
R17580 VOUT+.n169 VOUT+.t161 4.8295
R17581 VOUT+.n170 VOUT+.t134 4.8295
R17582 VOUT+.n172 VOUT+.t122 4.8295
R17583 VOUT+.n173 VOUT+.t87 4.8295
R17584 VOUT+.n175 VOUT+.t71 4.8295
R17585 VOUT+.n176 VOUT+.t46 4.8295
R17586 VOUT+.n97 VOUT+.t121 4.8295
R17587 VOUT+.n111 VOUT+.t52 4.8295
R17588 VOUT+.n113 VOUT+.t124 4.8295
R17589 VOUT+.n114 VOUT+.t94 4.8295
R17590 VOUT+.n116 VOUT+.t79 4.8295
R17591 VOUT+.n117 VOUT+.t61 4.8295
R17592 VOUT+.n119 VOUT+.t128 4.8295
R17593 VOUT+.n120 VOUT+.t107 4.8295
R17594 VOUT+.n122 VOUT+.t22 4.8295
R17595 VOUT+.n123 VOUT+.t149 4.8295
R17596 VOUT+.n125 VOUT+.t132 4.8295
R17597 VOUT+.n126 VOUT+.t114 4.8295
R17598 VOUT+.n128 VOUT+.t26 4.8295
R17599 VOUT+.n129 VOUT+.t154 4.8295
R17600 VOUT+.n131 VOUT+.t66 4.8295
R17601 VOUT+.n132 VOUT+.t39 4.8295
R17602 VOUT+.n178 VOUT+.t81 4.8295
R17603 VOUT+.n141 VOUT+.t158 4.8154
R17604 VOUT+.n140 VOUT+.t43 4.8154
R17605 VOUT+.n138 VOUT+.t65 4.8154
R17606 VOUT+.n137 VOUT+.t110 4.8154
R17607 VOUT+.n143 VOUT+.t140 4.806
R17608 VOUT+.n142 VOUT+.t120 4.806
R17609 VOUT+.n139 VOUT+.t83 4.806
R17610 VOUT+.n110 VOUT+.t69 4.806
R17611 VOUT+.n109 VOUT+.t116 4.806
R17612 VOUT+.n108 VOUT+.t57 4.806
R17613 VOUT+.n107 VOUT+.t109 4.806
R17614 VOUT+.n106 VOUT+.t44 4.806
R17615 VOUT+.n105 VOUT+.t146 4.806
R17616 VOUT+.n104 VOUT+.t33 4.806
R17617 VOUT+.n103 VOUT+.t135 4.806
R17618 VOUT+.n102 VOUT+.t74 4.806
R17619 VOUT+.n101 VOUT+.t25 4.806
R17620 VOUT+.n100 VOUT+.t68 4.806
R17621 VOUT+.n99 VOUT+.t20 4.806
R17622 VOUT+.n134 VOUT+.t76 4.5005
R17623 VOUT+.n135 VOUT+.t59 4.5005
R17624 VOUT+.n136 VOUT+.t100 4.5005
R17625 VOUT+.n137 VOUT+.t151 4.5005
R17626 VOUT+.n138 VOUT+.t112 4.5005
R17627 VOUT+.n139 VOUT+.t130 4.5005
R17628 VOUT+.n140 VOUT+.t84 4.5005
R17629 VOUT+.n141 VOUT+.t48 4.5005
R17630 VOUT+.n142 VOUT+.t160 4.5005
R17631 VOUT+.n143 VOUT+.t29 4.5005
R17632 VOUT+.n144 VOUT+.t141 4.5005
R17633 VOUT+.n145 VOUT+.t105 4.5005
R17634 VOUT+.n146 VOUT+.t126 4.5005
R17635 VOUT+.n147 VOUT+.t78 4.5005
R17636 VOUT+.n148 VOUT+.t73 4.5005
R17637 VOUT+.n150 VOUT+.t118 4.5005
R17638 VOUT+.n149 VOUT+.t32 4.5005
R17639 VOUT+.n151 VOUT+.t31 4.5005
R17640 VOUT+.n153 VOUT+.t67 4.5005
R17641 VOUT+.n152 VOUT+.t145 4.5005
R17642 VOUT+.n154 VOUT+.t143 4.5005
R17643 VOUT+.n156 VOUT+.t27 4.5005
R17644 VOUT+.n155 VOUT+.t104 4.5005
R17645 VOUT+.n157 VOUT+.t102 4.5005
R17646 VOUT+.n159 VOUT+.t137 4.5005
R17647 VOUT+.n158 VOUT+.t58 4.5005
R17648 VOUT+.n160 VOUT+.t138 4.5005
R17649 VOUT+.n162 VOUT+.t23 4.5005
R17650 VOUT+.n161 VOUT+.t91 4.5005
R17651 VOUT+.n163 VOUT+.t90 4.5005
R17652 VOUT+.n165 VOUT+.t129 4.5005
R17653 VOUT+.n164 VOUT+.t50 4.5005
R17654 VOUT+.n166 VOUT+.t93 4.5005
R17655 VOUT+.n168 VOUT+.t99 4.5005
R17656 VOUT+.n167 VOUT+.t41 4.5005
R17657 VOUT+.n169 VOUT+.t133 4.5005
R17658 VOUT+.n171 VOUT+.t136 4.5005
R17659 VOUT+.n170 VOUT+.t77 4.5005
R17660 VOUT+.n172 VOUT+.t86 4.5005
R17661 VOUT+.n174 VOUT+.t88 4.5005
R17662 VOUT+.n173 VOUT+.t36 4.5005
R17663 VOUT+.n175 VOUT+.t45 4.5005
R17664 VOUT+.n177 VOUT+.t47 4.5005
R17665 VOUT+.n176 VOUT+.t150 4.5005
R17666 VOUT+.n98 VOUT+.t127 4.5005
R17667 VOUT+.n97 VOUT+.t64 4.5005
R17668 VOUT+.n99 VOUT+.t55 4.5005
R17669 VOUT+.n100 VOUT+.t21 4.5005
R17670 VOUT+.n101 VOUT+.t119 4.5005
R17671 VOUT+.n102 VOUT+.t72 4.5005
R17672 VOUT+.n103 VOUT+.t35 4.5005
R17673 VOUT+.n104 VOUT+.t156 4.5005
R17674 VOUT+.n105 VOUT+.t98 4.5005
R17675 VOUT+.n106 VOUT+.t63 4.5005
R17676 VOUT+.n107 VOUT+.t24 4.5005
R17677 VOUT+.n108 VOUT+.t123 4.5005
R17678 VOUT+.n109 VOUT+.t75 4.5005
R17679 VOUT+.n110 VOUT+.t51 4.5005
R17680 VOUT+.n112 VOUT+.t53 4.5005
R17681 VOUT+.n111 VOUT+.t157 4.5005
R17682 VOUT+.n113 VOUT+.t95 4.5005
R17683 VOUT+.n115 VOUT+.t97 4.5005
R17684 VOUT+.n114 VOUT+.t42 4.5005
R17685 VOUT+.n116 VOUT+.t60 4.5005
R17686 VOUT+.n118 VOUT+.t62 4.5005
R17687 VOUT+.n117 VOUT+.t159 4.5005
R17688 VOUT+.n119 VOUT+.t106 4.5005
R17689 VOUT+.n121 VOUT+.t108 4.5005
R17690 VOUT+.n120 VOUT+.t49 4.5005
R17691 VOUT+.n122 VOUT+.t147 4.5005
R17692 VOUT+.n124 VOUT+.t148 4.5005
R17693 VOUT+.n123 VOUT+.t89 4.5005
R17694 VOUT+.n125 VOUT+.t113 4.5005
R17695 VOUT+.n127 VOUT+.t115 4.5005
R17696 VOUT+.n126 VOUT+.t56 4.5005
R17697 VOUT+.n128 VOUT+.t153 4.5005
R17698 VOUT+.n130 VOUT+.t155 4.5005
R17699 VOUT+.n129 VOUT+.t101 4.5005
R17700 VOUT+.n131 VOUT+.t38 4.5005
R17701 VOUT+.n133 VOUT+.t40 4.5005
R17702 VOUT+.n132 VOUT+.t142 4.5005
R17703 VOUT+.n180 VOUT+.t80 4.5005
R17704 VOUT+.n179 VOUT+.t82 4.5005
R17705 VOUT+.n178 VOUT+.t30 4.5005
R17706 VOUT+.n181 VOUT+.t117 4.5005
R17707 VOUT+.n60 VOUT+.n37 4.5005
R17708 VOUT+.n61 VOUT+.n40 4.5005
R17709 VOUT+.n62 VOUT+.n41 4.5005
R17710 VOUT+.n64 VOUT+.n63 4.5005
R17711 VOUT+.n87 VOUT+.n86 4.5005
R17712 VOUT+.n83 VOUT+.n80 4.5005
R17713 VOUT+.n87 VOUT+.n80 4.5005
R17714 VOUT+.n88 VOUT+.n32 4.5005
R17715 VOUT+.n88 VOUT+.n34 4.5005
R17716 VOUT+.n88 VOUT+.n87 4.5005
R17717 VOUT+.n186 VOUT+.n91 4.5005
R17718 VOUT+.n187 VOUT+.n186 4.5005
R17719 VOUT+.n187 VOUT+.n28 4.5005
R17720 VOUT+.n188 VOUT+.n27 4.5005
R17721 VOUT+.n188 VOUT+.n187 4.5005
R17722 VOUT+.n192 VOUT+.n191 4.5005
R17723 VOUT+.n191 VOUT+.n19 4.5005
R17724 VOUT+.n22 VOUT+.n19 4.5005
R17725 VOUT+.n194 VOUT+.n19 4.5005
R17726 VOUT+.n196 VOUT+.n19 4.5005
R17727 VOUT+.n195 VOUT+.n22 4.5005
R17728 VOUT+.n195 VOUT+.n194 4.5005
R17729 VOUT+.n196 VOUT+.n195 4.5005
R17730 VOUT+.n1 VOUT+.t13 3.42907
R17731 VOUT+.n1 VOUT+.t17 3.42907
R17732 VOUT+.n5 VOUT+.t18 3.42907
R17733 VOUT+.n5 VOUT+.t11 3.42907
R17734 VOUT+.n8 VOUT+.t14 3.42907
R17735 VOUT+.n8 VOUT+.t0 3.42907
R17736 VOUT+.n85 VOUT+.n33 2.26725
R17737 VOUT+.n81 VOUT+.n31 2.24601
R17738 VOUT+.n190 VOUT+.n189 2.24601
R17739 VOUT+.n24 VOUT+.n21 2.24601
R17740 VOUT+.n185 VOUT+.n184 2.24477
R17741 VOUT+.n30 VOUT+.n25 2.24477
R17742 VOUT+.n88 VOUT+.n33 2.24063
R17743 VOUT+.n188 VOUT+.n26 2.24063
R17744 VOUT+.n195 VOUT+.n23 2.24063
R17745 VOUT+.n80 VOUT+.n79 2.24063
R17746 VOUT+.n186 VOUT+.n89 2.24063
R17747 VOUT+.n90 VOUT+.n28 2.24063
R17748 VOUT+.n193 VOUT+.n192 2.24063
R17749 VOUT+.n192 VOUT+.n20 2.24063
R17750 VOUT+.n86 VOUT+.n84 2.23934
R17751 VOUT+.n86 VOUT+.n82 2.23934
R17752 VOUT+.n6 VOUT+.n4 1.83719
R17753 VOUT+.n10 VOUT+.n9 1.72967
R17754 VOUT+.n17 VOUT+.n2 1.72967
R17755 VOUT+.n78 VOUT+.n77 1.5005
R17756 VOUT+.n76 VOUT+.n35 1.5005
R17757 VOUT+.n75 VOUT+.n74 1.5005
R17758 VOUT+.n73 VOUT+.n38 1.5005
R17759 VOUT+.n72 VOUT+.n71 1.5005
R17760 VOUT+.n70 VOUT+.n39 1.5005
R17761 VOUT+.n69 VOUT+.n68 1.5005
R17762 VOUT+.n67 VOUT+.n42 1.5005
R17763 VOUT+.n18 VOUT+.n17 1.5005
R17764 VOUT+.n16 VOUT+.n0 1.5005
R17765 VOUT+.n15 VOUT+.n14 1.5005
R17766 VOUT+.n13 VOUT+.n3 1.5005
R17767 VOUT+.n12 VOUT+.n11 1.5005
R17768 VOUT+.n64 VOUT+.n59 1.313
R17769 VOUT+.n55 VOUT+.n41 1.313
R17770 VOUT+.n52 VOUT+.n40 1.313
R17771 VOUT+.n49 VOUT+.n37 1.313
R17772 VOUT+.n45 VOUT+.n43 1.313
R17773 VOUT+.n47 VOUT+.n36 1.313
R17774 VOUT+.n187 VOUT+.n29 1.1455
R17775 VOUT+.n95 VOUT+.n94 1.13717
R17776 VOUT+.n96 VOUT+.n92 1.13717
R17777 VOUT+.n183 VOUT+.n182 1.13717
R17778 VOUT+.n93 VOUT+.n30 1.13717
R17779 VOUT+.n94 VOUT+.n27 1.13717
R17780 VOUT+.n92 VOUT+.n91 1.13717
R17781 VOUT+.n184 VOUT+.n183 1.13717
R17782 VOUT+.n87 VOUT+.n78 0.859875
R17783 VOUT+.n66 VOUT+.n43 0.715216
R17784 VOUT+.n65 VOUT+.n64 0.65675
R17785 VOUT+.n69 VOUT+.n41 0.65675
R17786 VOUT+.n71 VOUT+.n40 0.65675
R17787 VOUT+.n75 VOUT+.n37 0.65675
R17788 VOUT+.n77 VOUT+.n36 0.65675
R17789 VOUT+.n95 VOUT+.n29 0.585
R17790 VOUT+.n67 VOUT+.n66 0.564601
R17791 VOUT+.n61 VOUT+.n60 0.563
R17792 VOUT+.n62 VOUT+.n61 0.563
R17793 VOUT+.n63 VOUT+.n62 0.563
R17794 VOUT+.n57 VOUT+.n56 0.563
R17795 VOUT+.n56 VOUT+.n53 0.563
R17796 VOUT+.n53 VOUT+.n50 0.563
R17797 VOUT+.n197 VOUT+.n196 0.557792
R17798 VOUT+.n192 VOUT+.n188 0.5455
R17799 VOUT+.n138 VOUT+.n137 0.3295
R17800 VOUT+.n139 VOUT+.n138 0.3295
R17801 VOUT+.n140 VOUT+.n139 0.3295
R17802 VOUT+.n141 VOUT+.n140 0.3295
R17803 VOUT+.n142 VOUT+.n141 0.3295
R17804 VOUT+.n143 VOUT+.n142 0.3295
R17805 VOUT+.n144 VOUT+.n143 0.3295
R17806 VOUT+.n145 VOUT+.n144 0.3295
R17807 VOUT+.n146 VOUT+.n145 0.3295
R17808 VOUT+.n147 VOUT+.n146 0.3295
R17809 VOUT+.n148 VOUT+.n147 0.3295
R17810 VOUT+.n150 VOUT+.n148 0.3295
R17811 VOUT+.n150 VOUT+.n149 0.3295
R17812 VOUT+.n153 VOUT+.n151 0.3295
R17813 VOUT+.n153 VOUT+.n152 0.3295
R17814 VOUT+.n156 VOUT+.n154 0.3295
R17815 VOUT+.n156 VOUT+.n155 0.3295
R17816 VOUT+.n159 VOUT+.n157 0.3295
R17817 VOUT+.n159 VOUT+.n158 0.3295
R17818 VOUT+.n162 VOUT+.n160 0.3295
R17819 VOUT+.n162 VOUT+.n161 0.3295
R17820 VOUT+.n165 VOUT+.n163 0.3295
R17821 VOUT+.n165 VOUT+.n164 0.3295
R17822 VOUT+.n168 VOUT+.n166 0.3295
R17823 VOUT+.n168 VOUT+.n167 0.3295
R17824 VOUT+.n171 VOUT+.n169 0.3295
R17825 VOUT+.n171 VOUT+.n170 0.3295
R17826 VOUT+.n174 VOUT+.n172 0.3295
R17827 VOUT+.n174 VOUT+.n173 0.3295
R17828 VOUT+.n177 VOUT+.n175 0.3295
R17829 VOUT+.n177 VOUT+.n176 0.3295
R17830 VOUT+.n98 VOUT+.n97 0.3295
R17831 VOUT+.n100 VOUT+.n99 0.3295
R17832 VOUT+.n101 VOUT+.n100 0.3295
R17833 VOUT+.n102 VOUT+.n101 0.3295
R17834 VOUT+.n103 VOUT+.n102 0.3295
R17835 VOUT+.n104 VOUT+.n103 0.3295
R17836 VOUT+.n105 VOUT+.n104 0.3295
R17837 VOUT+.n106 VOUT+.n105 0.3295
R17838 VOUT+.n107 VOUT+.n106 0.3295
R17839 VOUT+.n108 VOUT+.n107 0.3295
R17840 VOUT+.n109 VOUT+.n108 0.3295
R17841 VOUT+.n110 VOUT+.n109 0.3295
R17842 VOUT+.n112 VOUT+.n110 0.3295
R17843 VOUT+.n112 VOUT+.n111 0.3295
R17844 VOUT+.n115 VOUT+.n113 0.3295
R17845 VOUT+.n115 VOUT+.n114 0.3295
R17846 VOUT+.n118 VOUT+.n116 0.3295
R17847 VOUT+.n118 VOUT+.n117 0.3295
R17848 VOUT+.n121 VOUT+.n119 0.3295
R17849 VOUT+.n121 VOUT+.n120 0.3295
R17850 VOUT+.n124 VOUT+.n122 0.3295
R17851 VOUT+.n124 VOUT+.n123 0.3295
R17852 VOUT+.n127 VOUT+.n125 0.3295
R17853 VOUT+.n127 VOUT+.n126 0.3295
R17854 VOUT+.n130 VOUT+.n128 0.3295
R17855 VOUT+.n130 VOUT+.n129 0.3295
R17856 VOUT+.n133 VOUT+.n131 0.3295
R17857 VOUT+.n133 VOUT+.n132 0.3295
R17858 VOUT+.n180 VOUT+.n179 0.3295
R17859 VOUT+.n179 VOUT+.n178 0.3295
R17860 VOUT+.n12 VOUT+.n4 0.314966
R17861 VOUT+.n181 VOUT+.n180 0.313833
R17862 VOUT+.n146 VOUT+.n134 0.306
R17863 VOUT+.n145 VOUT+.n135 0.306
R17864 VOUT+.n144 VOUT+.n136 0.306
R17865 VOUT+.n153 VOUT+.n150 0.2825
R17866 VOUT+.n156 VOUT+.n153 0.2825
R17867 VOUT+.n159 VOUT+.n156 0.2825
R17868 VOUT+.n162 VOUT+.n159 0.2825
R17869 VOUT+.n165 VOUT+.n162 0.2825
R17870 VOUT+.n168 VOUT+.n165 0.2825
R17871 VOUT+.n171 VOUT+.n168 0.2825
R17872 VOUT+.n174 VOUT+.n171 0.2825
R17873 VOUT+.n177 VOUT+.n174 0.2825
R17874 VOUT+.n112 VOUT+.n98 0.2825
R17875 VOUT+.n115 VOUT+.n112 0.2825
R17876 VOUT+.n118 VOUT+.n115 0.2825
R17877 VOUT+.n121 VOUT+.n118 0.2825
R17878 VOUT+.n124 VOUT+.n121 0.2825
R17879 VOUT+.n127 VOUT+.n124 0.2825
R17880 VOUT+.n130 VOUT+.n127 0.2825
R17881 VOUT+.n133 VOUT+.n130 0.2825
R17882 VOUT+.n179 VOUT+.n133 0.2825
R17883 VOUT+.n179 VOUT+.n177 0.2825
R17884 VOUT+.n186 VOUT+.n88 0.2455
R17885 VOUT+ VOUT+.n197 0.198417
R17886 VOUT+ VOUT+.n18 0.182792
R17887 VOUT+.n182 VOUT+.n181 0.138367
R17888 VOUT+.n10 VOUT+.n4 0.0891864
R17889 VOUT+.n65 VOUT+.n42 0.0577917
R17890 VOUT+.n69 VOUT+.n42 0.0577917
R17891 VOUT+.n70 VOUT+.n69 0.0577917
R17892 VOUT+.n71 VOUT+.n70 0.0577917
R17893 VOUT+.n71 VOUT+.n38 0.0577917
R17894 VOUT+.n75 VOUT+.n38 0.0577917
R17895 VOUT+.n76 VOUT+.n75 0.0577917
R17896 VOUT+.n77 VOUT+.n76 0.0577917
R17897 VOUT+.n68 VOUT+.n67 0.0577917
R17898 VOUT+.n68 VOUT+.n39 0.0577917
R17899 VOUT+.n72 VOUT+.n39 0.0577917
R17900 VOUT+.n73 VOUT+.n72 0.0577917
R17901 VOUT+.n74 VOUT+.n73 0.0577917
R17902 VOUT+.n74 VOUT+.n35 0.0577917
R17903 VOUT+.n78 VOUT+.n35 0.0577917
R17904 VOUT+.n66 VOUT+.n65 0.054517
R17905 VOUT+.n194 VOUT+.n24 0.047375
R17906 VOUT+.n189 VOUT+.n22 0.047375
R17907 VOUT+.n187 VOUT+.n30 0.0421667
R17908 VOUT+.n87 VOUT+.n81 0.0421667
R17909 VOUT+.n11 VOUT+.n10 0.0421667
R17910 VOUT+.n11 VOUT+.n3 0.0421667
R17911 VOUT+.n15 VOUT+.n3 0.0421667
R17912 VOUT+.n16 VOUT+.n15 0.0421667
R17913 VOUT+.n17 VOUT+.n16 0.0421667
R17914 VOUT+.n13 VOUT+.n12 0.0421667
R17915 VOUT+.n14 VOUT+.n13 0.0421667
R17916 VOUT+.n14 VOUT+.n0 0.0421667
R17917 VOUT+.n18 VOUT+.n0 0.0421667
R17918 VOUT+.n82 VOUT+.n81 0.0243161
R17919 VOUT+.n84 VOUT+.n32 0.0243161
R17920 VOUT+.n84 VOUT+.n83 0.0243161
R17921 VOUT+.n82 VOUT+.n34 0.0243161
R17922 VOUT+.n184 VOUT+.n26 0.0217373
R17923 VOUT+.n83 VOUT+.n33 0.0217373
R17924 VOUT+.n91 VOUT+.n26 0.0217373
R17925 VOUT+.n191 VOUT+.n23 0.0217373
R17926 VOUT+.n189 VOUT+.n23 0.0217373
R17927 VOUT+.n89 VOUT+.n30 0.0217373
R17928 VOUT+.n91 VOUT+.n90 0.0217373
R17929 VOUT+.n79 VOUT+.n32 0.0217373
R17930 VOUT+.n79 VOUT+.n34 0.0217373
R17931 VOUT+.n89 VOUT+.n27 0.0217373
R17932 VOUT+.n90 VOUT+.n27 0.0217373
R17933 VOUT+.n196 VOUT+.n20 0.0217373
R17934 VOUT+.n194 VOUT+.n193 0.0217373
R17935 VOUT+.n193 VOUT+.n22 0.0217373
R17936 VOUT+.n24 VOUT+.n20 0.0217373
R17937 VOUT+.n96 VOUT+.n95 0.0161667
R17938 VOUT+.n182 VOUT+.n96 0.0161667
R17939 VOUT+.n94 VOUT+.n93 0.0161667
R17940 VOUT+.n94 VOUT+.n92 0.0161667
R17941 VOUT+.n183 VOUT+.n92 0.0161667
R17942 VOUT+.n185 VOUT+.n28 0.0134654
R17943 VOUT+.n188 VOUT+.n25 0.0134654
R17944 VOUT+.n186 VOUT+.n185 0.0134654
R17945 VOUT+.n28 VOUT+.n25 0.0134654
R17946 VOUT+.n85 VOUT+.n80 0.0109778
R17947 VOUT+.n88 VOUT+.n31 0.0109778
R17948 VOUT+.n190 VOUT+.n19 0.0109778
R17949 VOUT+.n195 VOUT+.n21 0.0109778
R17950 VOUT+.n86 VOUT+.n85 0.0109778
R17951 VOUT+.n80 VOUT+.n31 0.0109778
R17952 VOUT+.n192 VOUT+.n190 0.0109778
R17953 VOUT+.n21 VOUT+.n19 0.0109778
R17954 VOUT+.n93 VOUT+.n29 0.00872683
R17955 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n21 344.178
R17956 bgr_11_0.V_TOP.n23 bgr_11_0.V_TOP.n22 334.772
R17957 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.t37 312.798
R17958 bgr_11_0.V_TOP bgr_11_0.V_TOP.t21 312.639
R17959 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.t45 312.5
R17960 bgr_11_0.V_TOP.n42 bgr_11_0.V_TOP.t33 310.401
R17961 bgr_11_0.V_TOP.n41 bgr_11_0.V_TOP.t42 310.401
R17962 bgr_11_0.V_TOP.n40 bgr_11_0.V_TOP.t49 310.401
R17963 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.t26 310.401
R17964 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.t25 310.401
R17965 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.t36 310.401
R17966 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.t27 310.401
R17967 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.t39 310.401
R17968 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.t48 310.401
R17969 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.t23 310.401
R17970 bgr_11_0.V_TOP.n1 bgr_11_0.V_TOP.t38 310.401
R17971 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.t14 308
R17972 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.t29 305.901
R17973 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n30 301.933
R17974 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n28 301.933
R17975 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n26 301.933
R17976 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n20 297.433
R17977 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.t0 108.424
R17978 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.t13 99.5675
R17979 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t10 39.4005
R17980 bgr_11_0.V_TOP.n22 bgr_11_0.V_TOP.t6 39.4005
R17981 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t5 39.4005
R17982 bgr_11_0.V_TOP.n21 bgr_11_0.V_TOP.t12 39.4005
R17983 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t11 39.4005
R17984 bgr_11_0.V_TOP.n20 bgr_11_0.V_TOP.t4 39.4005
R17985 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.t7 39.4005
R17986 bgr_11_0.V_TOP.n30 bgr_11_0.V_TOP.t9 39.4005
R17987 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t3 39.4005
R17988 bgr_11_0.V_TOP.n28 bgr_11_0.V_TOP.t8 39.4005
R17989 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t1 39.4005
R17990 bgr_11_0.V_TOP.n26 bgr_11_0.V_TOP.t2 39.4005
R17991 bgr_11_0.V_TOP.n19 bgr_11_0.V_TOP.n18 29.1779
R17992 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n19 16.5063
R17993 bgr_11_0.V_TOP.n32 bgr_11_0.V_TOP.n31 4.90675
R17994 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t24 4.8295
R17995 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t46 4.8295
R17996 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t34 4.8295
R17997 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t18 4.8295
R17998 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t22 4.8295
R17999 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t44 4.8295
R18000 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t47 4.8295
R18001 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.t35 4.8295
R18002 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.t41 4.8295
R18003 bgr_11_0.V_TOP.n8 bgr_11_0.V_TOP.t32 4.5005
R18004 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.t19 4.5005
R18005 bgr_11_0.V_TOP.n10 bgr_11_0.V_TOP.t40 4.5005
R18006 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.t31 4.5005
R18007 bgr_11_0.V_TOP.n12 bgr_11_0.V_TOP.t30 4.5005
R18008 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.t17 4.5005
R18009 bgr_11_0.V_TOP.n14 bgr_11_0.V_TOP.t16 4.5005
R18010 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.t43 4.5005
R18011 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.t20 4.5005
R18012 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.t28 4.5005
R18013 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.t15 4.5005
R18014 bgr_11_0.V_TOP.n7 bgr_11_0.V_TOP.n6 4.5005
R18015 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n0 4.5005
R18016 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.n34 4.5005
R18017 bgr_11_0.V_TOP.n25 bgr_11_0.V_TOP.n24 4.5005
R18018 bgr_11_0.V_TOP.n24 bgr_11_0.V_TOP.n23 1.59425
R18019 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n32 1.21925
R18020 bgr_11_0.V_TOP.n27 bgr_11_0.V_TOP.n25 1.1255
R18021 bgr_11_0.V_TOP.n29 bgr_11_0.V_TOP.n27 1.1255
R18022 bgr_11_0.V_TOP.n31 bgr_11_0.V_TOP.n29 1.1255
R18023 bgr_11_0.V_TOP.n9 bgr_11_0.V_TOP.n8 0.3295
R18024 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n10 0.3295
R18025 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n12 0.3295
R18026 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.n14 0.3295
R18027 bgr_11_0.V_TOP.n18 bgr_11_0.V_TOP.n17 0.3295
R18028 bgr_11_0.V_TOP.n17 bgr_11_0.V_TOP.n16 0.3295
R18029 bgr_11_0.V_TOP.n11 bgr_11_0.V_TOP.n9 0.2825
R18030 bgr_11_0.V_TOP.n13 bgr_11_0.V_TOP.n11 0.2825
R18031 bgr_11_0.V_TOP.n15 bgr_11_0.V_TOP.n13 0.2825
R18032 bgr_11_0.V_TOP.n16 bgr_11_0.V_TOP.n15 0.2825
R18033 bgr_11_0.V_TOP.n2 bgr_11_0.V_TOP.n1 0.28175
R18034 bgr_11_0.V_TOP.n3 bgr_11_0.V_TOP.n2 0.28175
R18035 bgr_11_0.V_TOP.n4 bgr_11_0.V_TOP.n3 0.28175
R18036 bgr_11_0.V_TOP.n5 bgr_11_0.V_TOP.n4 0.28175
R18037 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.n5 0.28175
R18038 bgr_11_0.V_TOP.n36 bgr_11_0.V_TOP.n35 0.28175
R18039 bgr_11_0.V_TOP.n37 bgr_11_0.V_TOP.n36 0.28175
R18040 bgr_11_0.V_TOP.n38 bgr_11_0.V_TOP.n37 0.28175
R18041 bgr_11_0.V_TOP.n39 bgr_11_0.V_TOP.n38 0.28175
R18042 bgr_11_0.V_TOP.n40 bgr_11_0.V_TOP.n39 0.28175
R18043 bgr_11_0.V_TOP.n41 bgr_11_0.V_TOP.n40 0.28175
R18044 bgr_11_0.V_TOP.n42 bgr_11_0.V_TOP.n41 0.28175
R18045 bgr_11_0.V_TOP.n6 bgr_11_0.V_TOP.n0 0.141125
R18046 bgr_11_0.V_TOP.n35 bgr_11_0.V_TOP.n0 0.141125
R18047 bgr_11_0.V_TOP bgr_11_0.V_TOP.n42 0.141125
R18048 bgr_11_0.V_TOP.n33 bgr_11_0.V_TOP.n7 0.141125
R18049 bgr_11_0.V_TOP.n34 bgr_11_0.V_TOP.n33 0.141125
R18050 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t9 651.343
R18051 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n7 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t8 647.968
R18052 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t7 537.922
R18053 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n0 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t6 117.243
R18054 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n1 107.266
R18055 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n4 105.016
R18056 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n3 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n2 105.016
R18057 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t2 13.1338
R18058 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n4 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t5 13.1338
R18059 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t3 13.1338
R18060 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n2 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t0 13.1338
R18061 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t4 13.1338
R18062 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n1 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t1 13.1338
R18063 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n5 7.32862
R18064 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n6 3.98488
R18065 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n5 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n3 2.2505
R18066 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n6 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n0 1.73488
R18067 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n7 1.53175
R18068 two_stage_opamp_dummy_magic_29_0.Vb1.n2 two_stage_opamp_dummy_magic_29_0.Vb1.t15 484.212
R18069 two_stage_opamp_dummy_magic_29_0.Vb1.n2 two_stage_opamp_dummy_magic_29_0.Vb1.t26 484.212
R18070 two_stage_opamp_dummy_magic_29_0.Vb1.n2 two_stage_opamp_dummy_magic_29_0.Vb1.t12 484.212
R18071 two_stage_opamp_dummy_magic_29_0.Vb1.n2 two_stage_opamp_dummy_magic_29_0.Vb1.t25 484.212
R18072 two_stage_opamp_dummy_magic_29_0.Vb1.n3 two_stage_opamp_dummy_magic_29_0.Vb1.t32 484.212
R18073 two_stage_opamp_dummy_magic_29_0.Vb1.n3 two_stage_opamp_dummy_magic_29_0.Vb1.t23 484.212
R18074 two_stage_opamp_dummy_magic_29_0.Vb1.n3 two_stage_opamp_dummy_magic_29_0.Vb1.t18 484.212
R18075 two_stage_opamp_dummy_magic_29_0.Vb1.n3 two_stage_opamp_dummy_magic_29_0.Vb1.t24 484.212
R18076 two_stage_opamp_dummy_magic_29_0.Vb1.n7 two_stage_opamp_dummy_magic_29_0.Vb1.t31 484.212
R18077 two_stage_opamp_dummy_magic_29_0.Vb1.n7 two_stage_opamp_dummy_magic_29_0.Vb1.t22 484.212
R18078 two_stage_opamp_dummy_magic_29_0.Vb1.n4 two_stage_opamp_dummy_magic_29_0.Vb1.t20 484.212
R18079 two_stage_opamp_dummy_magic_29_0.Vb1.n4 two_stage_opamp_dummy_magic_29_0.Vb1.t30 484.212
R18080 two_stage_opamp_dummy_magic_29_0.Vb1.n4 two_stage_opamp_dummy_magic_29_0.Vb1.t19 484.212
R18081 two_stage_opamp_dummy_magic_29_0.Vb1.n4 two_stage_opamp_dummy_magic_29_0.Vb1.t28 484.212
R18082 two_stage_opamp_dummy_magic_29_0.Vb1.n5 two_stage_opamp_dummy_magic_29_0.Vb1.t16 484.212
R18083 two_stage_opamp_dummy_magic_29_0.Vb1.n5 two_stage_opamp_dummy_magic_29_0.Vb1.t29 484.212
R18084 two_stage_opamp_dummy_magic_29_0.Vb1.n5 two_stage_opamp_dummy_magic_29_0.Vb1.t17 484.212
R18085 two_stage_opamp_dummy_magic_29_0.Vb1.n5 two_stage_opamp_dummy_magic_29_0.Vb1.t27 484.212
R18086 two_stage_opamp_dummy_magic_29_0.Vb1.n6 two_stage_opamp_dummy_magic_29_0.Vb1.t14 484.212
R18087 two_stage_opamp_dummy_magic_29_0.Vb1.n6 two_stage_opamp_dummy_magic_29_0.Vb1.t21 484.212
R18088 two_stage_opamp_dummy_magic_29_0.Vb1.n9 two_stage_opamp_dummy_magic_29_0.Vb1.t6 449.868
R18089 two_stage_opamp_dummy_magic_29_0.Vb1.n8 two_stage_opamp_dummy_magic_29_0.Vb1.t0 449.868
R18090 two_stage_opamp_dummy_magic_29_0.Vb1.n9 two_stage_opamp_dummy_magic_29_0.Vb1.t2 273.134
R18091 two_stage_opamp_dummy_magic_29_0.Vb1.n8 two_stage_opamp_dummy_magic_29_0.Vb1.t4 273.134
R18092 two_stage_opamp_dummy_magic_29_0.Vb1.n12 two_stage_opamp_dummy_magic_29_0.Vb1.t13 161.363
R18093 two_stage_opamp_dummy_magic_29_0.Vb1.n1 two_stage_opamp_dummy_magic_29_0.Vb1.n10 161.3
R18094 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.Vb1.n19 151.042
R18095 two_stage_opamp_dummy_magic_29_0.Vb1.n18 two_stage_opamp_dummy_magic_29_0.Vb1.n17 49.3505
R18096 two_stage_opamp_dummy_magic_29_0.Vb1.n1 two_stage_opamp_dummy_magic_29_0.Vb1.n11 49.3505
R18097 two_stage_opamp_dummy_magic_29_0.Vb1.n15 two_stage_opamp_dummy_magic_29_0.Vb1.n14 49.3505
R18098 two_stage_opamp_dummy_magic_29_0.Vb1.n10 two_stage_opamp_dummy_magic_29_0.Vb1.n9 45.5227
R18099 two_stage_opamp_dummy_magic_29_0.Vb1.n10 two_stage_opamp_dummy_magic_29_0.Vb1.n8 45.5227
R18100 two_stage_opamp_dummy_magic_29_0.Vb1.n2 two_stage_opamp_dummy_magic_29_0.Vb1.n0 21.4927
R18101 two_stage_opamp_dummy_magic_29_0.Vb1.n13 two_stage_opamp_dummy_magic_29_0.Vb1.n6 21.4927
R18102 two_stage_opamp_dummy_magic_29_0.Vb1.n19 two_stage_opamp_dummy_magic_29_0.Vb1.t9 19.7005
R18103 two_stage_opamp_dummy_magic_29_0.Vb1.n19 two_stage_opamp_dummy_magic_29_0.Vb1.t8 19.7005
R18104 two_stage_opamp_dummy_magic_29_0.Vb1.n17 two_stage_opamp_dummy_magic_29_0.Vb1.t7 16.0005
R18105 two_stage_opamp_dummy_magic_29_0.Vb1.n17 two_stage_opamp_dummy_magic_29_0.Vb1.t10 16.0005
R18106 two_stage_opamp_dummy_magic_29_0.Vb1.n11 two_stage_opamp_dummy_magic_29_0.Vb1.t5 16.0005
R18107 two_stage_opamp_dummy_magic_29_0.Vb1.n11 two_stage_opamp_dummy_magic_29_0.Vb1.t3 16.0005
R18108 two_stage_opamp_dummy_magic_29_0.Vb1.n14 two_stage_opamp_dummy_magic_29_0.Vb1.t11 16.0005
R18109 two_stage_opamp_dummy_magic_29_0.Vb1.n14 two_stage_opamp_dummy_magic_29_0.Vb1.t1 16.0005
R18110 two_stage_opamp_dummy_magic_29_0.Vb1.n18 two_stage_opamp_dummy_magic_29_0.Vb1.n16 5.28175
R18111 two_stage_opamp_dummy_magic_29_0.Vb1.n16 two_stage_opamp_dummy_magic_29_0.Vb1.n15 5.28175
R18112 two_stage_opamp_dummy_magic_29_0.Vb1.n15 two_stage_opamp_dummy_magic_29_0.Vb1.n13 4.938
R18113 two_stage_opamp_dummy_magic_29_0.Vb1.n0 two_stage_opamp_dummy_magic_29_0.Vb1.n18 4.938
R18114 two_stage_opamp_dummy_magic_29_0.Vb1.n1 two_stage_opamp_dummy_magic_29_0.Vb1.n0 4.5005
R18115 two_stage_opamp_dummy_magic_29_0.Vb1.n16 two_stage_opamp_dummy_magic_29_0.Vb1.n12 2.23569
R18116 two_stage_opamp_dummy_magic_29_0.Vb1.n5 two_stage_opamp_dummy_magic_29_0.Vb1.n4 1.03175
R18117 two_stage_opamp_dummy_magic_29_0.Vb1.n3 two_stage_opamp_dummy_magic_29_0.Vb1.n2 1.03175
R18118 two_stage_opamp_dummy_magic_29_0.Vb1.n12 two_stage_opamp_dummy_magic_29_0.Vb1.n1 0.937224
R18119 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.Vb1.n4 0.852062
R18120 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.Vb1.n7 0.852062
R18121 two_stage_opamp_dummy_magic_29_0.Vb1.n13 two_stage_opamp_dummy_magic_29_0.Vb1.n0 0.688
R18122 two_stage_opamp_dummy_magic_29_0.Vb1.n7 two_stage_opamp_dummy_magic_29_0.Vb1.n3 0.516125
R18123 two_stage_opamp_dummy_magic_29_0.Vb1.n6 two_stage_opamp_dummy_magic_29_0.Vb1.n5 0.516125
R18124 two_stage_opamp_dummy_magic_29_0.VD2.n1 two_stage_opamp_dummy_magic_29_0.VD2.n0 49.7255
R18125 two_stage_opamp_dummy_magic_29_0.VD2.n21 two_stage_opamp_dummy_magic_29_0.VD2.n12 49.7255
R18126 two_stage_opamp_dummy_magic_29_0.VD2.n11 two_stage_opamp_dummy_magic_29_0.VD2.n10 49.7255
R18127 two_stage_opamp_dummy_magic_29_0.VD2.n27 two_stage_opamp_dummy_magic_29_0.VD2.n9 49.7255
R18128 two_stage_opamp_dummy_magic_29_0.VD2.n25 two_stage_opamp_dummy_magic_29_0.VD2.n24 49.7255
R18129 two_stage_opamp_dummy_magic_29_0.VD2.n15 two_stage_opamp_dummy_magic_29_0.VD2.n14 49.3505
R18130 two_stage_opamp_dummy_magic_29_0.VD2.n18 two_stage_opamp_dummy_magic_29_0.VD2.n17 49.3505
R18131 two_stage_opamp_dummy_magic_29_0.VD2.n5 two_stage_opamp_dummy_magic_29_0.VD2.n4 49.3505
R18132 two_stage_opamp_dummy_magic_29_0.VD2.n35 two_stage_opamp_dummy_magic_29_0.VD2.n34 49.3505
R18133 two_stage_opamp_dummy_magic_29_0.VD2.n8 two_stage_opamp_dummy_magic_29_0.VD2.n7 49.3505
R18134 two_stage_opamp_dummy_magic_29_0.VD2.n31 two_stage_opamp_dummy_magic_29_0.VD2.n30 49.3505
R18135 two_stage_opamp_dummy_magic_29_0.VD2.n14 two_stage_opamp_dummy_magic_29_0.VD2.t19 16.0005
R18136 two_stage_opamp_dummy_magic_29_0.VD2.n14 two_stage_opamp_dummy_magic_29_0.VD2.t18 16.0005
R18137 two_stage_opamp_dummy_magic_29_0.VD2.n17 two_stage_opamp_dummy_magic_29_0.VD2.t21 16.0005
R18138 two_stage_opamp_dummy_magic_29_0.VD2.n17 two_stage_opamp_dummy_magic_29_0.VD2.t0 16.0005
R18139 two_stage_opamp_dummy_magic_29_0.VD2.n4 two_stage_opamp_dummy_magic_29_0.VD2.t6 16.0005
R18140 two_stage_opamp_dummy_magic_29_0.VD2.n4 two_stage_opamp_dummy_magic_29_0.VD2.t4 16.0005
R18141 two_stage_opamp_dummy_magic_29_0.VD2.n34 two_stage_opamp_dummy_magic_29_0.VD2.t5 16.0005
R18142 two_stage_opamp_dummy_magic_29_0.VD2.n34 two_stage_opamp_dummy_magic_29_0.VD2.t2 16.0005
R18143 two_stage_opamp_dummy_magic_29_0.VD2.n7 two_stage_opamp_dummy_magic_29_0.VD2.t7 16.0005
R18144 two_stage_opamp_dummy_magic_29_0.VD2.n7 two_stage_opamp_dummy_magic_29_0.VD2.t20 16.0005
R18145 two_stage_opamp_dummy_magic_29_0.VD2.n0 two_stage_opamp_dummy_magic_29_0.VD2.t13 16.0005
R18146 two_stage_opamp_dummy_magic_29_0.VD2.n0 two_stage_opamp_dummy_magic_29_0.VD2.t8 16.0005
R18147 two_stage_opamp_dummy_magic_29_0.VD2.n12 two_stage_opamp_dummy_magic_29_0.VD2.t12 16.0005
R18148 two_stage_opamp_dummy_magic_29_0.VD2.n12 two_stage_opamp_dummy_magic_29_0.VD2.t15 16.0005
R18149 two_stage_opamp_dummy_magic_29_0.VD2.n10 two_stage_opamp_dummy_magic_29_0.VD2.t14 16.0005
R18150 two_stage_opamp_dummy_magic_29_0.VD2.n10 two_stage_opamp_dummy_magic_29_0.VD2.t9 16.0005
R18151 two_stage_opamp_dummy_magic_29_0.VD2.n9 two_stage_opamp_dummy_magic_29_0.VD2.t10 16.0005
R18152 two_stage_opamp_dummy_magic_29_0.VD2.n9 two_stage_opamp_dummy_magic_29_0.VD2.t16 16.0005
R18153 two_stage_opamp_dummy_magic_29_0.VD2.n30 two_stage_opamp_dummy_magic_29_0.VD2.t1 16.0005
R18154 two_stage_opamp_dummy_magic_29_0.VD2.n30 two_stage_opamp_dummy_magic_29_0.VD2.t3 16.0005
R18155 two_stage_opamp_dummy_magic_29_0.VD2.n24 two_stage_opamp_dummy_magic_29_0.VD2.t11 16.0005
R18156 two_stage_opamp_dummy_magic_29_0.VD2.n24 two_stage_opamp_dummy_magic_29_0.VD2.t17 16.0005
R18157 two_stage_opamp_dummy_magic_29_0.VD2.n21 two_stage_opamp_dummy_magic_29_0.VD2.n20 8.89633
R18158 two_stage_opamp_dummy_magic_29_0.VD2.n13 two_stage_opamp_dummy_magic_29_0.VD2.n11 8.89633
R18159 two_stage_opamp_dummy_magic_29_0.VD2.n28 two_stage_opamp_dummy_magic_29_0.VD2.n27 8.89633
R18160 two_stage_opamp_dummy_magic_29_0.VD2.n25 two_stage_opamp_dummy_magic_29_0.VD2.n3 8.89633
R18161 two_stage_opamp_dummy_magic_29_0.VD2.n32 two_stage_opamp_dummy_magic_29_0.VD2.n8 5.438
R18162 two_stage_opamp_dummy_magic_29_0.VD2.n16 two_stage_opamp_dummy_magic_29_0.VD2.n15 5.438
R18163 two_stage_opamp_dummy_magic_29_0.VD2.n28 two_stage_opamp_dummy_magic_29_0.VD2.n8 5.31821
R18164 two_stage_opamp_dummy_magic_29_0.VD2.n15 two_stage_opamp_dummy_magic_29_0.VD2.n13 5.31821
R18165 two_stage_opamp_dummy_magic_29_0.VD2.n19 two_stage_opamp_dummy_magic_29_0.VD2.n18 5.08383
R18166 two_stage_opamp_dummy_magic_29_0.VD2.n5 two_stage_opamp_dummy_magic_29_0.VD2.n2 5.08383
R18167 two_stage_opamp_dummy_magic_29_0.VD2.n36 two_stage_opamp_dummy_magic_29_0.VD2.n35 5.08383
R18168 two_stage_opamp_dummy_magic_29_0.VD2.n31 two_stage_opamp_dummy_magic_29_0.VD2.n29 5.08383
R18169 two_stage_opamp_dummy_magic_29_0.VD2.n22 two_stage_opamp_dummy_magic_29_0.VD2.n11 5.063
R18170 two_stage_opamp_dummy_magic_29_0.VD2.n27 two_stage_opamp_dummy_magic_29_0.VD2.n26 5.063
R18171 two_stage_opamp_dummy_magic_29_0.VD2.n18 two_stage_opamp_dummy_magic_29_0.VD2.n16 4.8755
R18172 two_stage_opamp_dummy_magic_29_0.VD2.n6 two_stage_opamp_dummy_magic_29_0.VD2.n5 4.8755
R18173 two_stage_opamp_dummy_magic_29_0.VD2.n35 two_stage_opamp_dummy_magic_29_0.VD2.n33 4.8755
R18174 two_stage_opamp_dummy_magic_29_0.VD2.n32 two_stage_opamp_dummy_magic_29_0.VD2.n31 4.8755
R18175 two_stage_opamp_dummy_magic_29_0.VD2 two_stage_opamp_dummy_magic_29_0.VD2.n37 4.60467
R18176 two_stage_opamp_dummy_magic_29_0.VD2.n22 two_stage_opamp_dummy_magic_29_0.VD2.n21 4.5005
R18177 two_stage_opamp_dummy_magic_29_0.VD2.n23 two_stage_opamp_dummy_magic_29_0.VD2.n1 4.5005
R18178 two_stage_opamp_dummy_magic_29_0.VD2.n26 two_stage_opamp_dummy_magic_29_0.VD2.n25 4.5005
R18179 two_stage_opamp_dummy_magic_29_0.VD2 two_stage_opamp_dummy_magic_29_0.VD2.n1 4.29217
R18180 two_stage_opamp_dummy_magic_29_0.VD2.n23 two_stage_opamp_dummy_magic_29_0.VD2.n22 0.563
R18181 two_stage_opamp_dummy_magic_29_0.VD2.n26 two_stage_opamp_dummy_magic_29_0.VD2.n23 0.563
R18182 two_stage_opamp_dummy_magic_29_0.VD2.n33 two_stage_opamp_dummy_magic_29_0.VD2.n32 0.563
R18183 two_stage_opamp_dummy_magic_29_0.VD2.n33 two_stage_opamp_dummy_magic_29_0.VD2.n6 0.563
R18184 two_stage_opamp_dummy_magic_29_0.VD2.n16 two_stage_opamp_dummy_magic_29_0.VD2.n6 0.563
R18185 two_stage_opamp_dummy_magic_29_0.VD2.n29 two_stage_opamp_dummy_magic_29_0.VD2.n3 0.234875
R18186 two_stage_opamp_dummy_magic_29_0.VD2.n29 two_stage_opamp_dummy_magic_29_0.VD2.n28 0.234875
R18187 two_stage_opamp_dummy_magic_29_0.VD2.n19 two_stage_opamp_dummy_magic_29_0.VD2.n13 0.234875
R18188 two_stage_opamp_dummy_magic_29_0.VD2.n20 two_stage_opamp_dummy_magic_29_0.VD2.n19 0.234875
R18189 two_stage_opamp_dummy_magic_29_0.VD2.n20 two_stage_opamp_dummy_magic_29_0.VD2.n2 0.234875
R18190 two_stage_opamp_dummy_magic_29_0.VD2.n37 two_stage_opamp_dummy_magic_29_0.VD2.n2 0.234875
R18191 two_stage_opamp_dummy_magic_29_0.VD2.n37 two_stage_opamp_dummy_magic_29_0.VD2.n36 0.234875
R18192 two_stage_opamp_dummy_magic_29_0.VD2.n36 two_stage_opamp_dummy_magic_29_0.VD2.n3 0.234875
R18193 bgr_11_0.1st_Vout_1.n12 bgr_11_0.1st_Vout_1.t29 363.909
R18194 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.t13 351.88
R18195 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n22 299.25
R18196 bgr_11_0.1st_Vout_1.n14 bgr_11_0.1st_Vout_1.n13 299.25
R18197 bgr_11_0.1st_Vout_1.n18 bgr_11_0.1st_Vout_1.n17 297.807
R18198 bgr_11_0.1st_Vout_1.n20 bgr_11_0.1st_Vout_1.t30 194.809
R18199 bgr_11_0.1st_Vout_1.n20 bgr_11_0.1st_Vout_1.t10 194.809
R18200 bgr_11_0.1st_Vout_1.n15 bgr_11_0.1st_Vout_1.t28 194.809
R18201 bgr_11_0.1st_Vout_1.n15 bgr_11_0.1st_Vout_1.t19 194.809
R18202 bgr_11_0.1st_Vout_1.n21 bgr_11_0.1st_Vout_1.n20 163.097
R18203 bgr_11_0.1st_Vout_1.n16 bgr_11_0.1st_Vout_1.n15 163.097
R18204 bgr_11_0.1st_Vout_1.n18 bgr_11_0.1st_Vout_1.t3 49.4474
R18205 bgr_11_0.1st_Vout_1.n22 bgr_11_0.1st_Vout_1.t0 39.4005
R18206 bgr_11_0.1st_Vout_1.n22 bgr_11_0.1st_Vout_1.t1 39.4005
R18207 bgr_11_0.1st_Vout_1.n13 bgr_11_0.1st_Vout_1.t5 39.4005
R18208 bgr_11_0.1st_Vout_1.n13 bgr_11_0.1st_Vout_1.t4 39.4005
R18209 bgr_11_0.1st_Vout_1.n17 bgr_11_0.1st_Vout_1.t2 39.4005
R18210 bgr_11_0.1st_Vout_1.n17 bgr_11_0.1st_Vout_1.t6 39.4005
R18211 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t27 4.8295
R18212 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t14 4.8295
R18213 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.t32 4.8295
R18214 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t22 4.8295
R18215 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t25 4.8295
R18216 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t12 4.8295
R18217 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t16 4.8295
R18218 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t7 4.8295
R18219 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.t24 4.8295
R18220 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.t18 4.5005
R18221 bgr_11_0.1st_Vout_1.n1 bgr_11_0.1st_Vout_1.t23 4.5005
R18222 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.t26 4.5005
R18223 bgr_11_0.1st_Vout_1.n3 bgr_11_0.1st_Vout_1.t31 4.5005
R18224 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.t17 4.5005
R18225 bgr_11_0.1st_Vout_1.n5 bgr_11_0.1st_Vout_1.t21 4.5005
R18226 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.t8 4.5005
R18227 bgr_11_0.1st_Vout_1.n7 bgr_11_0.1st_Vout_1.t11 4.5005
R18228 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.t15 4.5005
R18229 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.t20 4.5005
R18230 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.t9 4.5005
R18231 bgr_11_0.1st_Vout_1.n19 bgr_11_0.1st_Vout_1.n18 1.44719
R18232 bgr_11_0.1st_Vout_1.n2 bgr_11_0.1st_Vout_1.n1 0.3295
R18233 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n3 0.3295
R18234 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.n5 0.3295
R18235 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.n7 0.3295
R18236 bgr_11_0.1st_Vout_1.n10 bgr_11_0.1st_Vout_1.n9 0.3295
R18237 bgr_11_0.1st_Vout_1.n11 bgr_11_0.1st_Vout_1.n10 0.3295
R18238 bgr_11_0.1st_Vout_1.n4 bgr_11_0.1st_Vout_1.n2 0.2825
R18239 bgr_11_0.1st_Vout_1.n6 bgr_11_0.1st_Vout_1.n4 0.2825
R18240 bgr_11_0.1st_Vout_1.n8 bgr_11_0.1st_Vout_1.n6 0.2825
R18241 bgr_11_0.1st_Vout_1.n9 bgr_11_0.1st_Vout_1.n8 0.2825
R18242 bgr_11_0.1st_Vout_1.n19 bgr_11_0.1st_Vout_1.n16 0.2505
R18243 bgr_11_0.1st_Vout_1.n0 bgr_11_0.1st_Vout_1.n21 0.2505
R18244 bgr_11_0.1st_Vout_1.n14 bgr_11_0.1st_Vout_1.n12 0.21925
R18245 bgr_11_0.1st_Vout_1.n16 bgr_11_0.1st_Vout_1.n14 0.1255
R18246 bgr_11_0.1st_Vout_1.n21 bgr_11_0.1st_Vout_1.n19 0.1255
R18247 bgr_11_0.1st_Vout_1 bgr_11_0.1st_Vout_1.n0 0.09425
R18248 bgr_11_0.1st_Vout_1.n12 bgr_11_0.1st_Vout_1.n11 10.102
R18249 bgr_11_0.cap_res1.t0 bgr_11_0.cap_res1.t14 121.983
R18250 bgr_11_0.cap_res1.t10 bgr_11_0.cap_res1.t18 0.1603
R18251 bgr_11_0.cap_res1.t17 bgr_11_0.cap_res1.t20 0.1603
R18252 bgr_11_0.cap_res1.t9 bgr_11_0.cap_res1.t16 0.1603
R18253 bgr_11_0.cap_res1.t2 bgr_11_0.cap_res1.t8 0.1603
R18254 bgr_11_0.cap_res1.t7 bgr_11_0.cap_res1.t15 0.1603
R18255 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t11 0.159278
R18256 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t4 0.159278
R18257 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t12 0.159278
R18258 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t19 0.159278
R18259 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t10 0.1368
R18260 bgr_11_0.cap_res1.n4 bgr_11_0.cap_res1.t6 0.1368
R18261 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t17 0.1368
R18262 bgr_11_0.cap_res1.n3 bgr_11_0.cap_res1.t13 0.1368
R18263 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t9 0.1368
R18264 bgr_11_0.cap_res1.n2 bgr_11_0.cap_res1.t5 0.1368
R18265 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t2 0.1368
R18266 bgr_11_0.cap_res1.n1 bgr_11_0.cap_res1.t1 0.1368
R18267 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t7 0.1368
R18268 bgr_11_0.cap_res1.n0 bgr_11_0.cap_res1.t3 0.1368
R18269 bgr_11_0.cap_res1.t11 bgr_11_0.cap_res1.n0 0.00152174
R18270 bgr_11_0.cap_res1.t4 bgr_11_0.cap_res1.n1 0.00152174
R18271 bgr_11_0.cap_res1.t12 bgr_11_0.cap_res1.n2 0.00152174
R18272 bgr_11_0.cap_res1.t19 bgr_11_0.cap_res1.n3 0.00152174
R18273 bgr_11_0.cap_res1.t14 bgr_11_0.cap_res1.n4 0.00152174
R18274 two_stage_opamp_dummy_magic_29_0.VD3.n3 two_stage_opamp_dummy_magic_29_0.VD3.t35 671.418
R18275 two_stage_opamp_dummy_magic_29_0.VD3.n15 two_stage_opamp_dummy_magic_29_0.VD3.t32 671.418
R18276 two_stage_opamp_dummy_magic_29_0.VD3.n14 two_stage_opamp_dummy_magic_29_0.VD3.t33 213.131
R18277 two_stage_opamp_dummy_magic_29_0.VD3.t36 two_stage_opamp_dummy_magic_29_0.VD3.n13 213.131
R18278 two_stage_opamp_dummy_magic_29_0.VD3.t33 two_stage_opamp_dummy_magic_29_0.VD3.t10 146.155
R18279 two_stage_opamp_dummy_magic_29_0.VD3.t10 two_stage_opamp_dummy_magic_29_0.VD3.t0 146.155
R18280 two_stage_opamp_dummy_magic_29_0.VD3.t0 two_stage_opamp_dummy_magic_29_0.VD3.t6 146.155
R18281 two_stage_opamp_dummy_magic_29_0.VD3.t6 two_stage_opamp_dummy_magic_29_0.VD3.t14 146.155
R18282 two_stage_opamp_dummy_magic_29_0.VD3.t14 two_stage_opamp_dummy_magic_29_0.VD3.t8 146.155
R18283 two_stage_opamp_dummy_magic_29_0.VD3.t8 two_stage_opamp_dummy_magic_29_0.VD3.t16 146.155
R18284 two_stage_opamp_dummy_magic_29_0.VD3.t16 two_stage_opamp_dummy_magic_29_0.VD3.t4 146.155
R18285 two_stage_opamp_dummy_magic_29_0.VD3.t4 two_stage_opamp_dummy_magic_29_0.VD3.t12 146.155
R18286 two_stage_opamp_dummy_magic_29_0.VD3.t12 two_stage_opamp_dummy_magic_29_0.VD3.t2 146.155
R18287 two_stage_opamp_dummy_magic_29_0.VD3.t2 two_stage_opamp_dummy_magic_29_0.VD3.t18 146.155
R18288 two_stage_opamp_dummy_magic_29_0.VD3.t18 two_stage_opamp_dummy_magic_29_0.VD3.t36 146.155
R18289 two_stage_opamp_dummy_magic_29_0.VD3.n14 two_stage_opamp_dummy_magic_29_0.VD3.t34 76.2576
R18290 two_stage_opamp_dummy_magic_29_0.VD3.n13 two_stage_opamp_dummy_magic_29_0.VD3.t37 76.2576
R18291 two_stage_opamp_dummy_magic_29_0.VD3.n0 two_stage_opamp_dummy_magic_29_0.VD3.n19 67.013
R18292 two_stage_opamp_dummy_magic_29_0.VD3.n28 two_stage_opamp_dummy_magic_29_0.VD3.n16 67.013
R18293 two_stage_opamp_dummy_magic_29_0.VD3.n12 two_stage_opamp_dummy_magic_29_0.VD3.n11 67.013
R18294 two_stage_opamp_dummy_magic_29_0.VD3.n31 two_stage_opamp_dummy_magic_29_0.VD3.n8 67.013
R18295 two_stage_opamp_dummy_magic_29_0.VD3.n33 two_stage_opamp_dummy_magic_29_0.VD3.n32 67.013
R18296 two_stage_opamp_dummy_magic_29_0.VD3.n5 two_stage_opamp_dummy_magic_29_0.VD3.n4 66.0338
R18297 two_stage_opamp_dummy_magic_29_0.VD3.n7 two_stage_opamp_dummy_magic_29_0.VD3.n6 66.0338
R18298 two_stage_opamp_dummy_magic_29_0.VD3.n10 two_stage_opamp_dummy_magic_29_0.VD3.n9 66.0338
R18299 two_stage_opamp_dummy_magic_29_0.VD3.n23 two_stage_opamp_dummy_magic_29_0.VD3.n22 66.0338
R18300 two_stage_opamp_dummy_magic_29_0.VD3.n18 two_stage_opamp_dummy_magic_29_0.VD3.n17 66.0338
R18301 two_stage_opamp_dummy_magic_29_0.VD3.n27 two_stage_opamp_dummy_magic_29_0.VD3.n26 66.0338
R18302 two_stage_opamp_dummy_magic_29_0.VD3.n19 two_stage_opamp_dummy_magic_29_0.VD3.t11 11.2576
R18303 two_stage_opamp_dummy_magic_29_0.VD3.n19 two_stage_opamp_dummy_magic_29_0.VD3.t1 11.2576
R18304 two_stage_opamp_dummy_magic_29_0.VD3.n16 two_stage_opamp_dummy_magic_29_0.VD3.t7 11.2576
R18305 two_stage_opamp_dummy_magic_29_0.VD3.n16 two_stage_opamp_dummy_magic_29_0.VD3.t15 11.2576
R18306 two_stage_opamp_dummy_magic_29_0.VD3.n11 two_stage_opamp_dummy_magic_29_0.VD3.t9 11.2576
R18307 two_stage_opamp_dummy_magic_29_0.VD3.n11 two_stage_opamp_dummy_magic_29_0.VD3.t17 11.2576
R18308 two_stage_opamp_dummy_magic_29_0.VD3.n8 two_stage_opamp_dummy_magic_29_0.VD3.t5 11.2576
R18309 two_stage_opamp_dummy_magic_29_0.VD3.n8 two_stage_opamp_dummy_magic_29_0.VD3.t13 11.2576
R18310 two_stage_opamp_dummy_magic_29_0.VD3.n4 two_stage_opamp_dummy_magic_29_0.VD3.t28 11.2576
R18311 two_stage_opamp_dummy_magic_29_0.VD3.n4 two_stage_opamp_dummy_magic_29_0.VD3.t21 11.2576
R18312 two_stage_opamp_dummy_magic_29_0.VD3.n6 two_stage_opamp_dummy_magic_29_0.VD3.t26 11.2576
R18313 two_stage_opamp_dummy_magic_29_0.VD3.n6 two_stage_opamp_dummy_magic_29_0.VD3.t24 11.2576
R18314 two_stage_opamp_dummy_magic_29_0.VD3.n9 two_stage_opamp_dummy_magic_29_0.VD3.t27 11.2576
R18315 two_stage_opamp_dummy_magic_29_0.VD3.n9 two_stage_opamp_dummy_magic_29_0.VD3.t31 11.2576
R18316 two_stage_opamp_dummy_magic_29_0.VD3.n22 two_stage_opamp_dummy_magic_29_0.VD3.t30 11.2576
R18317 two_stage_opamp_dummy_magic_29_0.VD3.n22 two_stage_opamp_dummy_magic_29_0.VD3.t23 11.2576
R18318 two_stage_opamp_dummy_magic_29_0.VD3.n17 two_stage_opamp_dummy_magic_29_0.VD3.t29 11.2576
R18319 two_stage_opamp_dummy_magic_29_0.VD3.n17 two_stage_opamp_dummy_magic_29_0.VD3.t22 11.2576
R18320 two_stage_opamp_dummy_magic_29_0.VD3.n26 two_stage_opamp_dummy_magic_29_0.VD3.t20 11.2576
R18321 two_stage_opamp_dummy_magic_29_0.VD3.n26 two_stage_opamp_dummy_magic_29_0.VD3.t25 11.2576
R18322 two_stage_opamp_dummy_magic_29_0.VD3.n32 two_stage_opamp_dummy_magic_29_0.VD3.t3 11.2576
R18323 two_stage_opamp_dummy_magic_29_0.VD3.n32 two_stage_opamp_dummy_magic_29_0.VD3.t19 11.2576
R18324 two_stage_opamp_dummy_magic_29_0.VD3.n27 two_stage_opamp_dummy_magic_29_0.VD3.n25 5.66717
R18325 two_stage_opamp_dummy_magic_29_0.VD3.n20 two_stage_opamp_dummy_magic_29_0.VD3.n5 5.66717
R18326 two_stage_opamp_dummy_magic_29_0.VD3.n20 two_stage_opamp_dummy_magic_29_0.VD3.n7 5.29217
R18327 two_stage_opamp_dummy_magic_29_0.VD3.n21 two_stage_opamp_dummy_magic_29_0.VD3.n10 5.29217
R18328 two_stage_opamp_dummy_magic_29_0.VD3.n24 two_stage_opamp_dummy_magic_29_0.VD3.n23 5.29217
R18329 two_stage_opamp_dummy_magic_29_0.VD3.n25 two_stage_opamp_dummy_magic_29_0.VD3.n18 5.29217
R18330 two_stage_opamp_dummy_magic_29_0.VD3.n15 two_stage_opamp_dummy_magic_29_0.VD3.n14 1.90883
R18331 two_stage_opamp_dummy_magic_29_0.VD3.n13 two_stage_opamp_dummy_magic_29_0.VD3.n3 1.90883
R18332 two_stage_opamp_dummy_magic_29_0.VD3.n33 two_stage_opamp_dummy_magic_29_0.VD3.n7 1.02133
R18333 two_stage_opamp_dummy_magic_29_0.VD3.n31 two_stage_opamp_dummy_magic_29_0.VD3.n10 1.02133
R18334 two_stage_opamp_dummy_magic_29_0.VD3.n23 two_stage_opamp_dummy_magic_29_0.VD3.n12 1.02133
R18335 two_stage_opamp_dummy_magic_29_0.VD3.n28 two_stage_opamp_dummy_magic_29_0.VD3.n18 1.02133
R18336 two_stage_opamp_dummy_magic_29_0.VD3.n0 two_stage_opamp_dummy_magic_29_0.VD3.n27 1.02133
R18337 two_stage_opamp_dummy_magic_29_0.VD3.n34 two_stage_opamp_dummy_magic_29_0.VD3.n5 1.02133
R18338 two_stage_opamp_dummy_magic_29_0.VD3 two_stage_opamp_dummy_magic_29_0.VD3.n34 0.65675
R18339 two_stage_opamp_dummy_magic_29_0.VD3.n33 two_stage_opamp_dummy_magic_29_0.VD3.n2 0.643357
R18340 two_stage_opamp_dummy_magic_29_0.VD3.n31 two_stage_opamp_dummy_magic_29_0.VD3.n30 0.643357
R18341 two_stage_opamp_dummy_magic_29_0.VD3.n29 two_stage_opamp_dummy_magic_29_0.VD3.n12 0.643357
R18342 two_stage_opamp_dummy_magic_29_0.VD3.n1 two_stage_opamp_dummy_magic_29_0.VD3.n0 0.0279681
R18343 two_stage_opamp_dummy_magic_29_0.VD3.n25 two_stage_opamp_dummy_magic_29_0.VD3.n24 0.3755
R18344 two_stage_opamp_dummy_magic_29_0.VD3.n24 two_stage_opamp_dummy_magic_29_0.VD3.n21 0.3755
R18345 two_stage_opamp_dummy_magic_29_0.VD3.n21 two_stage_opamp_dummy_magic_29_0.VD3.n20 0.3755
R18346 two_stage_opamp_dummy_magic_29_0.VD3.n0 two_stage_opamp_dummy_magic_29_0.VD3.n15 0.131952
R18347 two_stage_opamp_dummy_magic_29_0.VD3.n34 two_stage_opamp_dummy_magic_29_0.VD3.n3 0.104667
R18348 two_stage_opamp_dummy_magic_29_0.VD3.n28 two_stage_opamp_dummy_magic_29_0.VD3.n1 0.0471695
R18349 two_stage_opamp_dummy_magic_29_0.VD3.n29 two_stage_opamp_dummy_magic_29_0.VD3.n1 0.274589
R18350 two_stage_opamp_dummy_magic_29_0.VD3.n30 two_stage_opamp_dummy_magic_29_0.VD3.n29 0.0540714
R18351 two_stage_opamp_dummy_magic_29_0.VD3.n30 two_stage_opamp_dummy_magic_29_0.VD3.n2 0.0540714
R18352 two_stage_opamp_dummy_magic_29_0.VD3.n28 two_stage_opamp_dummy_magic_29_0.VD3.n12 0.0540714
R18353 two_stage_opamp_dummy_magic_29_0.VD3.n31 two_stage_opamp_dummy_magic_29_0.VD3.n12 0.0540714
R18354 two_stage_opamp_dummy_magic_29_0.VD3.n33 two_stage_opamp_dummy_magic_29_0.VD3.n31 0.0540714
R18355 two_stage_opamp_dummy_magic_29_0.VD3.n34 two_stage_opamp_dummy_magic_29_0.VD3.n33 0.0540714
R18356 two_stage_opamp_dummy_magic_29_0.VD3 two_stage_opamp_dummy_magic_29_0.VD3.n2 0.0406786
R18357 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t6 369.534
R18358 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t9 369.534
R18359 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.t22 369.534
R18360 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t20 369.534
R18361 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.t13 369.534
R18362 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.t11 369.534
R18363 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.t0 369.534
R18364 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n1 360.288
R18365 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.t7 249.034
R18366 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.t5 192.8
R18367 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.t12 192.8
R18368 bgr_11_0.NFET_GATE_10uA.n3 bgr_11_0.NFET_GATE_10uA.t19 192.8
R18369 bgr_11_0.NFET_GATE_10uA.n2 bgr_11_0.NFET_GATE_10uA.t18 192.8
R18370 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.t15 192.8
R18371 bgr_11_0.NFET_GATE_10uA.n8 bgr_11_0.NFET_GATE_10uA.t23 192.8
R18372 bgr_11_0.NFET_GATE_10uA.n7 bgr_11_0.NFET_GATE_10uA.t8 192.8
R18373 bgr_11_0.NFET_GATE_10uA.n15 bgr_11_0.NFET_GATE_10uA.t10 192.8
R18374 bgr_11_0.NFET_GATE_10uA.n12 bgr_11_0.NFET_GATE_10uA.t17 192.8
R18375 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.t16 192.8
R18376 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.t21 192.8
R18377 bgr_11_0.NFET_GATE_10uA.n18 bgr_11_0.NFET_GATE_10uA.t14 192.8
R18378 bgr_11_0.NFET_GATE_10uA.n5 bgr_11_0.NFET_GATE_10uA.n4 176.733
R18379 bgr_11_0.NFET_GATE_10uA.n4 bgr_11_0.NFET_GATE_10uA.n3 176.733
R18380 bgr_11_0.NFET_GATE_10uA.n9 bgr_11_0.NFET_GATE_10uA.n8 176.733
R18381 bgr_11_0.NFET_GATE_10uA.n13 bgr_11_0.NFET_GATE_10uA.n12 176.733
R18382 bgr_11_0.NFET_GATE_10uA.n14 bgr_11_0.NFET_GATE_10uA.n13 176.733
R18383 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.n6 168.014
R18384 bgr_11_0.NFET_GATE_10uA.n11 bgr_11_0.NFET_GATE_10uA.n10 166.343
R18385 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.n16 166.343
R18386 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n19 166.343
R18387 bgr_11_0.NFET_GATE_10uA.n20 bgr_11_0.NFET_GATE_10uA.n0 141.752
R18388 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n5 56.2338
R18389 bgr_11_0.NFET_GATE_10uA.n6 bgr_11_0.NFET_GATE_10uA.n2 56.2338
R18390 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.n9 56.2338
R18391 bgr_11_0.NFET_GATE_10uA.n10 bgr_11_0.NFET_GATE_10uA.n7 56.2338
R18392 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n15 56.2338
R18393 bgr_11_0.NFET_GATE_10uA.n16 bgr_11_0.NFET_GATE_10uA.n14 56.2338
R18394 bgr_11_0.NFET_GATE_10uA.n19 bgr_11_0.NFET_GATE_10uA.n18 56.2338
R18395 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t3 39.4005
R18396 bgr_11_0.NFET_GATE_10uA.n1 bgr_11_0.NFET_GATE_10uA.t2 39.4005
R18397 bgr_11_0.NFET_GATE_10uA.n20 bgr_11_0.NFET_GATE_10uA.t4 24.0005
R18398 bgr_11_0.NFET_GATE_10uA.t1 bgr_11_0.NFET_GATE_10uA.n20 24.0005
R18399 bgr_11_0.NFET_GATE_10uA.n0 bgr_11_0.NFET_GATE_10uA.n17 2.01612
R18400 bgr_11_0.NFET_GATE_10uA.n17 bgr_11_0.NFET_GATE_10uA.n11 1.5005
R18401 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP_NFET1.t0 141.653
R18402 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.t18 310.488
R18403 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t13 310.488
R18404 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t17 310.488
R18405 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n8 297.433
R18406 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n3 297.433
R18407 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.n14 297.433
R18408 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.t10 184.097
R18409 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.t8 184.097
R18410 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.t6 184.097
R18411 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.n11 167.094
R18412 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.n5 167.094
R18413 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.n0 167.094
R18414 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.n13 161.3
R18415 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.n7 161.3
R18416 bgr_11_0.V_mir1.n4 bgr_11_0.V_mir1.n2 161.3
R18417 bgr_11_0.V_mir1.n11 bgr_11_0.V_mir1.t14 120.501
R18418 bgr_11_0.V_mir1.n12 bgr_11_0.V_mir1.t4 120.501
R18419 bgr_11_0.V_mir1.n5 bgr_11_0.V_mir1.t15 120.501
R18420 bgr_11_0.V_mir1.n6 bgr_11_0.V_mir1.t2 120.501
R18421 bgr_11_0.V_mir1.n0 bgr_11_0.V_mir1.t16 120.501
R18422 bgr_11_0.V_mir1.n1 bgr_11_0.V_mir1.t0 120.501
R18423 bgr_11_0.V_mir1.n9 bgr_11_0.V_mir1.t12 50.2004
R18424 bgr_11_0.V_mir1.n13 bgr_11_0.V_mir1.n12 40.7027
R18425 bgr_11_0.V_mir1.n7 bgr_11_0.V_mir1.n6 40.7027
R18426 bgr_11_0.V_mir1.n2 bgr_11_0.V_mir1.n1 40.7027
R18427 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t9 39.4005
R18428 bgr_11_0.V_mir1.n8 bgr_11_0.V_mir1.t3 39.4005
R18429 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t7 39.4005
R18430 bgr_11_0.V_mir1.n3 bgr_11_0.V_mir1.t1 39.4005
R18431 bgr_11_0.V_mir1.t11 bgr_11_0.V_mir1.n15 39.4005
R18432 bgr_11_0.V_mir1.n15 bgr_11_0.V_mir1.t5 39.4005
R18433 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n4 6.6255
R18434 bgr_11_0.V_mir1.n14 bgr_11_0.V_mir1.n10 6.6255
R18435 bgr_11_0.V_mir1.n10 bgr_11_0.V_mir1.n9 4.5005
R18436 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n2 301.983
R18437 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n4 297.151
R18438 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n0 297.151
R18439 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n15 118.861
R18440 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n17 118.861
R18441 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n21 118.861
R18442 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n25 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n24 118.861
R18443 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n28 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n27 118.861
R18444 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n30 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t10 115.672
R18445 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t15 39.4005
R18446 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n4 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t14 39.4005
R18447 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t12 39.4005
R18448 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t11 39.4005
R18449 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t13 39.4005
R18450 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n0 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t16 39.4005
R18451 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t8 19.7005
R18452 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n15 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t1 19.7005
R18453 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t5 19.7005
R18454 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n17 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t0 19.7005
R18455 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t4 19.7005
R18456 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n21 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t9 19.7005
R18457 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n24 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t7 19.7005
R18458 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n24 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t3 19.7005
R18459 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n27 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t6 19.7005
R18460 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n27 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t2 19.7005
R18461 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n41 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n5 11.9588
R18462 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n41 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n40 11.6203
R18463 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n41 9.92238
R18464 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n28 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n26 5.54217
R18465 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n16 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n14 5.54217
R18466 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n1 5.39633
R18467 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n5 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n3 5.39633
R18468 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n16 5.38592
R18469 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n18 5.04217
R18470 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n22 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n20 5.04217
R18471 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n25 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n13 5.04217
R18472 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n29 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n28 5.04217
R18473 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n18 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n14 4.97967
R18474 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n23 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n22 4.97967
R18475 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n26 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n25 4.97967
R18476 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n7 4.5005
R18477 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n38 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n37 4.5005
R18478 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n37 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n36 4.5005
R18479 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n11 4.5005
R18480 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n30 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n29 2.99007
R18481 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n33 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n32 2.26187
R18482 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n34 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n33 2.26187
R18483 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n39 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n38 2.24063
R18484 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n8 2.24063
R18485 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n31 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n10 2.24063
R18486 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n40 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n6 2.24063
R18487 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n35 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n34 2.24063
R18488 bgr_11_0.V_CMFB_S3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n1 1.34946
R18489 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n26 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n23 0.563
R18490 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n23 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n14 0.563
R18491 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n31 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n30 0.464042
R18492 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n19 0.34425
R18493 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n20 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n13 0.34425
R18494 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n29 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n13 0.34425
R18495 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n35 0.078625
R18496 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n38 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n8 0.0421667
R18497 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n40 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n39 0.0217373
R18498 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n37 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n9 0.0217373
R18499 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n35 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n10 0.0217373
R18500 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n39 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n7 0.0217373
R18501 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n9 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n7 0.0217373
R18502 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n32 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n11 0.0217373
R18503 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n12 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n10 0.0217373
R18504 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n32 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n31 0.0217373
R18505 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n33 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n12 0.0217373
R18506 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n36 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n6 0.0217373
R18507 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n8 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n6 0.0217373
R18508 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n34 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n11 0.0217373
R18509 a_3230_6968.t0 a_3230_6968.t1 169.905
R18510 VIN+.n0 VIN+.t9 1097.62
R18511 VIN+ VIN+.n9 433.019
R18512 VIN+.n9 VIN+.t4 273.134
R18513 VIN+.n0 VIN+.t6 273.134
R18514 VIN+.n8 VIN+.t0 273.134
R18515 VIN+.n7 VIN+.t3 273.134
R18516 VIN+.n6 VIN+.t10 273.134
R18517 VIN+.n5 VIN+.t2 273.134
R18518 VIN+.n4 VIN+.t7 273.134
R18519 VIN+.n3 VIN+.t5 273.134
R18520 VIN+.n2 VIN+.t8 273.134
R18521 VIN+.n1 VIN+.t1 273.134
R18522 VIN+.n1 VIN+.n0 176.733
R18523 VIN+.n2 VIN+.n1 176.733
R18524 VIN+.n3 VIN+.n2 176.733
R18525 VIN+.n4 VIN+.n3 176.733
R18526 VIN+.n5 VIN+.n4 176.733
R18527 VIN+.n6 VIN+.n5 176.733
R18528 VIN+.n7 VIN+.n6 176.733
R18529 VIN+.n8 VIN+.n7 176.733
R18530 VIN+.n9 VIN+.n8 176.733
R18531 a_6350_30238.t0 a_6350_30238.t1 178.133
R18532 bgr_11_0.Vin+ bgr_11_0.Vin+.t6 529.879
R18533 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t0 148.653
R18534 bgr_11_0.Vin+.n0 bgr_11_0.Vin+.t5 125.418
R18535 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n1 106.609
R18536 bgr_11_0.Vin+.n3 bgr_11_0.Vin+.n2 104.484
R18537 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n0 25.0809
R18538 bgr_11_0.Vin+.n4 bgr_11_0.Vin+.n3 18.7817
R18539 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t3 13.1338
R18540 bgr_11_0.Vin+.n2 bgr_11_0.Vin+.t2 13.1338
R18541 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t1 13.1338
R18542 bgr_11_0.Vin+.n1 bgr_11_0.Vin+.t4 13.1338
R18543 bgr_11_0.Vin+ bgr_11_0.Vin+.n4 6.53175
R18544 two_stage_opamp_dummy_magic_29_0.V_err_gate.n2 two_stage_opamp_dummy_magic_29_0.V_err_gate.t9 479.322
R18545 two_stage_opamp_dummy_magic_29_0.V_err_gate.n2 two_stage_opamp_dummy_magic_29_0.V_err_gate.t7 479.322
R18546 two_stage_opamp_dummy_magic_29_0.V_err_gate.n6 two_stage_opamp_dummy_magic_29_0.V_err_gate.t8 479.322
R18547 two_stage_opamp_dummy_magic_29_0.V_err_gate.n6 two_stage_opamp_dummy_magic_29_0.V_err_gate.t6 479.322
R18548 two_stage_opamp_dummy_magic_29_0.V_err_gate.n3 two_stage_opamp_dummy_magic_29_0.V_err_gate.n1 178.075
R18549 two_stage_opamp_dummy_magic_29_0.V_err_gate.n5 two_stage_opamp_dummy_magic_29_0.V_err_gate.n4 177.434
R18550 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_err_gate.n0 170.357
R18551 two_stage_opamp_dummy_magic_29_0.V_err_gate.n3 two_stage_opamp_dummy_magic_29_0.V_err_gate.n2 165.8
R18552 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_err_gate.n6 165.8
R18553 two_stage_opamp_dummy_magic_29_0.V_err_gate.n0 two_stage_opamp_dummy_magic_29_0.V_err_gate.t1 24.0005
R18554 two_stage_opamp_dummy_magic_29_0.V_err_gate.n0 two_stage_opamp_dummy_magic_29_0.V_err_gate.t2 24.0005
R18555 two_stage_opamp_dummy_magic_29_0.V_err_gate.n4 two_stage_opamp_dummy_magic_29_0.V_err_gate.t3 15.7605
R18556 two_stage_opamp_dummy_magic_29_0.V_err_gate.n4 two_stage_opamp_dummy_magic_29_0.V_err_gate.t5 15.7605
R18557 two_stage_opamp_dummy_magic_29_0.V_err_gate.n1 two_stage_opamp_dummy_magic_29_0.V_err_gate.t0 15.7605
R18558 two_stage_opamp_dummy_magic_29_0.V_err_gate.n1 two_stage_opamp_dummy_magic_29_0.V_err_gate.t4 15.7605
R18559 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_err_gate.n5 1.76612
R18560 two_stage_opamp_dummy_magic_29_0.V_err_gate.n5 two_stage_opamp_dummy_magic_29_0.V_err_gate.n3 0.641125
R18561 a_6540_22450.n11 a_6540_22450.t18 310.488
R18562 a_6540_22450.n5 a_6540_22450.t13 310.488
R18563 a_6540_22450.n0 a_6540_22450.t14 310.488
R18564 a_6540_22450.n9 a_6540_22450.n8 297.433
R18565 a_6540_22450.n4 a_6540_22450.n3 297.433
R18566 a_6540_22450.n15 a_6540_22450.n14 297.433
R18567 a_6540_22450.n13 a_6540_22450.t7 184.097
R18568 a_6540_22450.n7 a_6540_22450.t5 184.097
R18569 a_6540_22450.n2 a_6540_22450.t3 184.097
R18570 a_6540_22450.n12 a_6540_22450.n11 167.094
R18571 a_6540_22450.n6 a_6540_22450.n5 167.094
R18572 a_6540_22450.n1 a_6540_22450.n0 167.094
R18573 a_6540_22450.n14 a_6540_22450.n13 161.3
R18574 a_6540_22450.n9 a_6540_22450.n7 161.3
R18575 a_6540_22450.n4 a_6540_22450.n2 161.3
R18576 a_6540_22450.n11 a_6540_22450.t15 120.501
R18577 a_6540_22450.n12 a_6540_22450.t11 120.501
R18578 a_6540_22450.n5 a_6540_22450.t17 120.501
R18579 a_6540_22450.n6 a_6540_22450.t1 120.501
R18580 a_6540_22450.n0 a_6540_22450.t16 120.501
R18581 a_6540_22450.n1 a_6540_22450.t9 120.501
R18582 a_6540_22450.n9 a_6540_22450.t0 50.2004
R18583 a_6540_22450.n13 a_6540_22450.n12 40.7027
R18584 a_6540_22450.n7 a_6540_22450.n6 40.7027
R18585 a_6540_22450.n2 a_6540_22450.n1 40.7027
R18586 a_6540_22450.n8 a_6540_22450.t2 39.4005
R18587 a_6540_22450.n8 a_6540_22450.t6 39.4005
R18588 a_6540_22450.n3 a_6540_22450.t10 39.4005
R18589 a_6540_22450.n3 a_6540_22450.t4 39.4005
R18590 a_6540_22450.t12 a_6540_22450.n15 39.4005
R18591 a_6540_22450.n15 a_6540_22450.t8 39.4005
R18592 a_6540_22450.n10 a_6540_22450.n4 6.6255
R18593 a_6540_22450.n14 a_6540_22450.n10 6.6255
R18594 a_6540_22450.n10 a_6540_22450.n9 4.5005
R18595 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t5 573.044
R18596 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n1 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t0 433.8
R18597 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n0 184.09
R18598 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n2 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n1 163.978
R18599 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n2 33.0088
R18600 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t2 15.7605
R18601 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n0 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t3 15.7605
R18602 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t1 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n3 9.6005
R18603 two_stage_opamp_dummy_magic_29_0.err_amp_mir.n3 two_stage_opamp_dummy_magic_29_0.err_amp_mir.t4 9.6005
R18604 two_stage_opamp_dummy_magic_29_0.err_amp_out.n0 two_stage_opamp_dummy_magic_29_0.err_amp_out.t4 610.534
R18605 two_stage_opamp_dummy_magic_29_0.err_amp_out.n0 two_stage_opamp_dummy_magic_29_0.err_amp_out.t5 433.8
R18606 two_stage_opamp_dummy_magic_29_0.err_amp_out two_stage_opamp_dummy_magic_29_0.err_amp_out.n0 267.139
R18607 two_stage_opamp_dummy_magic_29_0.err_amp_out.n3 two_stage_opamp_dummy_magic_29_0.err_amp_out.n2 178.829
R18608 two_stage_opamp_dummy_magic_29_0.err_amp_out.n3 two_stage_opamp_dummy_magic_29_0.err_amp_out.n1 38.5609
R18609 two_stage_opamp_dummy_magic_29_0.err_amp_out.n2 two_stage_opamp_dummy_magic_29_0.err_amp_out.t2 15.7605
R18610 two_stage_opamp_dummy_magic_29_0.err_amp_out.n2 two_stage_opamp_dummy_magic_29_0.err_amp_out.t0 15.7605
R18611 two_stage_opamp_dummy_magic_29_0.err_amp_out.n1 two_stage_opamp_dummy_magic_29_0.err_amp_out.t3 9.6005
R18612 two_stage_opamp_dummy_magic_29_0.err_amp_out.n1 two_stage_opamp_dummy_magic_29_0.err_amp_out.t1 9.6005
R18613 two_stage_opamp_dummy_magic_29_0.err_amp_out two_stage_opamp_dummy_magic_29_0.err_amp_out.n3 0.922375
R18614 two_stage_opamp_dummy_magic_29_0.Vb1_2 two_stage_opamp_dummy_magic_29_0.Vb1_2.t0 74.8571
R18615 two_stage_opamp_dummy_magic_29_0.Vb1_2 two_stage_opamp_dummy_magic_29_0.Vb1_2.n1 54.689
R18616 two_stage_opamp_dummy_magic_29_0.Vb1_2 two_stage_opamp_dummy_magic_29_0.Vb1_2.n0 54.689
R18617 two_stage_opamp_dummy_magic_29_0.Vb1_2.n0 two_stage_opamp_dummy_magic_29_0.Vb1_2.t2 16.0005
R18618 two_stage_opamp_dummy_magic_29_0.Vb1_2.n0 two_stage_opamp_dummy_magic_29_0.Vb1_2.t4 16.0005
R18619 two_stage_opamp_dummy_magic_29_0.Vb1_2.n1 two_stage_opamp_dummy_magic_29_0.Vb1_2.t3 16.0005
R18620 two_stage_opamp_dummy_magic_29_0.Vb1_2.n1 two_stage_opamp_dummy_magic_29_0.Vb1_2.t1 16.0005
R18621 two_stage_opamp_dummy_magic_29_0.VD1.n1 two_stage_opamp_dummy_magic_29_0.VD1.n0 49.7255
R18622 two_stage_opamp_dummy_magic_29_0.VD1.n25 two_stage_opamp_dummy_magic_29_0.VD1.n24 49.7255
R18623 two_stage_opamp_dummy_magic_29_0.VD1.n27 two_stage_opamp_dummy_magic_29_0.VD1.n9 49.7255
R18624 two_stage_opamp_dummy_magic_29_0.VD1.n21 two_stage_opamp_dummy_magic_29_0.VD1.n12 49.7255
R18625 two_stage_opamp_dummy_magic_29_0.VD1.n11 two_stage_opamp_dummy_magic_29_0.VD1.n10 49.7255
R18626 two_stage_opamp_dummy_magic_29_0.VD1.n15 two_stage_opamp_dummy_magic_29_0.VD1.n14 49.3505
R18627 two_stage_opamp_dummy_magic_29_0.VD1.n8 two_stage_opamp_dummy_magic_29_0.VD1.n7 49.3505
R18628 two_stage_opamp_dummy_magic_29_0.VD1.n31 two_stage_opamp_dummy_magic_29_0.VD1.n30 49.3505
R18629 two_stage_opamp_dummy_magic_29_0.VD1.n35 two_stage_opamp_dummy_magic_29_0.VD1.n34 49.3505
R18630 two_stage_opamp_dummy_magic_29_0.VD1.n5 two_stage_opamp_dummy_magic_29_0.VD1.n4 49.3505
R18631 two_stage_opamp_dummy_magic_29_0.VD1.n18 two_stage_opamp_dummy_magic_29_0.VD1.n17 49.3505
R18632 two_stage_opamp_dummy_magic_29_0.VD1.n14 two_stage_opamp_dummy_magic_29_0.VD1.t15 16.0005
R18633 two_stage_opamp_dummy_magic_29_0.VD1.n14 two_stage_opamp_dummy_magic_29_0.VD1.t12 16.0005
R18634 two_stage_opamp_dummy_magic_29_0.VD1.n7 two_stage_opamp_dummy_magic_29_0.VD1.t17 16.0005
R18635 two_stage_opamp_dummy_magic_29_0.VD1.n7 two_stage_opamp_dummy_magic_29_0.VD1.t14 16.0005
R18636 two_stage_opamp_dummy_magic_29_0.VD1.n30 two_stage_opamp_dummy_magic_29_0.VD1.t21 16.0005
R18637 two_stage_opamp_dummy_magic_29_0.VD1.n30 two_stage_opamp_dummy_magic_29_0.VD1.t18 16.0005
R18638 two_stage_opamp_dummy_magic_29_0.VD1.n34 two_stage_opamp_dummy_magic_29_0.VD1.t16 16.0005
R18639 two_stage_opamp_dummy_magic_29_0.VD1.n34 two_stage_opamp_dummy_magic_29_0.VD1.t0 16.0005
R18640 two_stage_opamp_dummy_magic_29_0.VD1.n4 two_stage_opamp_dummy_magic_29_0.VD1.t13 16.0005
R18641 two_stage_opamp_dummy_magic_29_0.VD1.n4 two_stage_opamp_dummy_magic_29_0.VD1.t20 16.0005
R18642 two_stage_opamp_dummy_magic_29_0.VD1.n0 two_stage_opamp_dummy_magic_29_0.VD1.t3 16.0005
R18643 two_stage_opamp_dummy_magic_29_0.VD1.n0 two_stage_opamp_dummy_magic_29_0.VD1.t10 16.0005
R18644 two_stage_opamp_dummy_magic_29_0.VD1.n24 two_stage_opamp_dummy_magic_29_0.VD1.t4 16.0005
R18645 two_stage_opamp_dummy_magic_29_0.VD1.n24 two_stage_opamp_dummy_magic_29_0.VD1.t8 16.0005
R18646 two_stage_opamp_dummy_magic_29_0.VD1.n9 two_stage_opamp_dummy_magic_29_0.VD1.t2 16.0005
R18647 two_stage_opamp_dummy_magic_29_0.VD1.n9 two_stage_opamp_dummy_magic_29_0.VD1.t7 16.0005
R18648 two_stage_opamp_dummy_magic_29_0.VD1.n12 two_stage_opamp_dummy_magic_29_0.VD1.t5 16.0005
R18649 two_stage_opamp_dummy_magic_29_0.VD1.n12 two_stage_opamp_dummy_magic_29_0.VD1.t9 16.0005
R18650 two_stage_opamp_dummy_magic_29_0.VD1.n17 two_stage_opamp_dummy_magic_29_0.VD1.t19 16.0005
R18651 two_stage_opamp_dummy_magic_29_0.VD1.n17 two_stage_opamp_dummy_magic_29_0.VD1.t1 16.0005
R18652 two_stage_opamp_dummy_magic_29_0.VD1.n10 two_stage_opamp_dummy_magic_29_0.VD1.t6 16.0005
R18653 two_stage_opamp_dummy_magic_29_0.VD1.n10 two_stage_opamp_dummy_magic_29_0.VD1.t11 16.0005
R18654 two_stage_opamp_dummy_magic_29_0.VD1.n25 two_stage_opamp_dummy_magic_29_0.VD1.n3 8.89633
R18655 two_stage_opamp_dummy_magic_29_0.VD1.n28 two_stage_opamp_dummy_magic_29_0.VD1.n27 8.89633
R18656 two_stage_opamp_dummy_magic_29_0.VD1.n21 two_stage_opamp_dummy_magic_29_0.VD1.n20 8.89633
R18657 two_stage_opamp_dummy_magic_29_0.VD1.n13 two_stage_opamp_dummy_magic_29_0.VD1.n11 8.89633
R18658 two_stage_opamp_dummy_magic_29_0.VD1.n32 two_stage_opamp_dummy_magic_29_0.VD1.n8 5.438
R18659 two_stage_opamp_dummy_magic_29_0.VD1.n16 two_stage_opamp_dummy_magic_29_0.VD1.n15 5.438
R18660 two_stage_opamp_dummy_magic_29_0.VD1.n28 two_stage_opamp_dummy_magic_29_0.VD1.n8 5.31821
R18661 two_stage_opamp_dummy_magic_29_0.VD1.n15 two_stage_opamp_dummy_magic_29_0.VD1.n13 5.31821
R18662 two_stage_opamp_dummy_magic_29_0.VD1.n31 two_stage_opamp_dummy_magic_29_0.VD1.n29 5.08383
R18663 two_stage_opamp_dummy_magic_29_0.VD1.n36 two_stage_opamp_dummy_magic_29_0.VD1.n35 5.08383
R18664 two_stage_opamp_dummy_magic_29_0.VD1.n5 two_stage_opamp_dummy_magic_29_0.VD1.n2 5.08383
R18665 two_stage_opamp_dummy_magic_29_0.VD1.n19 two_stage_opamp_dummy_magic_29_0.VD1.n18 5.08383
R18666 two_stage_opamp_dummy_magic_29_0.VD1.n27 two_stage_opamp_dummy_magic_29_0.VD1.n26 5.063
R18667 two_stage_opamp_dummy_magic_29_0.VD1.n22 two_stage_opamp_dummy_magic_29_0.VD1.n11 5.063
R18668 two_stage_opamp_dummy_magic_29_0.VD1.n32 two_stage_opamp_dummy_magic_29_0.VD1.n31 4.8755
R18669 two_stage_opamp_dummy_magic_29_0.VD1.n35 two_stage_opamp_dummy_magic_29_0.VD1.n33 4.8755
R18670 two_stage_opamp_dummy_magic_29_0.VD1.n6 two_stage_opamp_dummy_magic_29_0.VD1.n5 4.8755
R18671 two_stage_opamp_dummy_magic_29_0.VD1.n18 two_stage_opamp_dummy_magic_29_0.VD1.n16 4.8755
R18672 two_stage_opamp_dummy_magic_29_0.VD1 two_stage_opamp_dummy_magic_29_0.VD1.n37 4.60467
R18673 two_stage_opamp_dummy_magic_29_0.VD1.n26 two_stage_opamp_dummy_magic_29_0.VD1.n25 4.5005
R18674 two_stage_opamp_dummy_magic_29_0.VD1.n23 two_stage_opamp_dummy_magic_29_0.VD1.n1 4.5005
R18675 two_stage_opamp_dummy_magic_29_0.VD1.n22 two_stage_opamp_dummy_magic_29_0.VD1.n21 4.5005
R18676 two_stage_opamp_dummy_magic_29_0.VD1 two_stage_opamp_dummy_magic_29_0.VD1.n1 4.29217
R18677 two_stage_opamp_dummy_magic_29_0.VD1.n26 two_stage_opamp_dummy_magic_29_0.VD1.n23 0.563
R18678 two_stage_opamp_dummy_magic_29_0.VD1.n23 two_stage_opamp_dummy_magic_29_0.VD1.n22 0.563
R18679 two_stage_opamp_dummy_magic_29_0.VD1.n33 two_stage_opamp_dummy_magic_29_0.VD1.n32 0.563
R18680 two_stage_opamp_dummy_magic_29_0.VD1.n33 two_stage_opamp_dummy_magic_29_0.VD1.n6 0.563
R18681 two_stage_opamp_dummy_magic_29_0.VD1.n16 two_stage_opamp_dummy_magic_29_0.VD1.n6 0.563
R18682 two_stage_opamp_dummy_magic_29_0.VD1.n19 two_stage_opamp_dummy_magic_29_0.VD1.n13 0.234875
R18683 two_stage_opamp_dummy_magic_29_0.VD1.n20 two_stage_opamp_dummy_magic_29_0.VD1.n19 0.234875
R18684 two_stage_opamp_dummy_magic_29_0.VD1.n20 two_stage_opamp_dummy_magic_29_0.VD1.n2 0.234875
R18685 two_stage_opamp_dummy_magic_29_0.VD1.n37 two_stage_opamp_dummy_magic_29_0.VD1.n2 0.234875
R18686 two_stage_opamp_dummy_magic_29_0.VD1.n37 two_stage_opamp_dummy_magic_29_0.VD1.n36 0.234875
R18687 two_stage_opamp_dummy_magic_29_0.VD1.n36 two_stage_opamp_dummy_magic_29_0.VD1.n3 0.234875
R18688 two_stage_opamp_dummy_magic_29_0.VD1.n29 two_stage_opamp_dummy_magic_29_0.VD1.n3 0.234875
R18689 two_stage_opamp_dummy_magic_29_0.VD1.n29 two_stage_opamp_dummy_magic_29_0.VD1.n28 0.234875
R18690 bgr_11_0.cap_res2.t0 bgr_11_0.cap_res2.t15 121.931
R18691 bgr_11_0.cap_res2.t10 bgr_11_0.cap_res2.t4 0.1603
R18692 bgr_11_0.cap_res2.t14 bgr_11_0.cap_res2.t9 0.1603
R18693 bgr_11_0.cap_res2.t8 bgr_11_0.cap_res2.t3 0.1603
R18694 bgr_11_0.cap_res2.t2 bgr_11_0.cap_res2.t16 0.1603
R18695 bgr_11_0.cap_res2.t6 bgr_11_0.cap_res2.t1 0.1603
R18696 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t11 0.159278
R18697 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t7 0.159278
R18698 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t13 0.159278
R18699 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t19 0.159278
R18700 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t20 0.1368
R18701 bgr_11_0.cap_res2.n4 bgr_11_0.cap_res2.t10 0.1368
R18702 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t5 0.1368
R18703 bgr_11_0.cap_res2.n3 bgr_11_0.cap_res2.t14 0.1368
R18704 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t18 0.1368
R18705 bgr_11_0.cap_res2.n2 bgr_11_0.cap_res2.t8 0.1368
R18706 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t12 0.1368
R18707 bgr_11_0.cap_res2.n1 bgr_11_0.cap_res2.t2 0.1368
R18708 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t17 0.1368
R18709 bgr_11_0.cap_res2.n0 bgr_11_0.cap_res2.t6 0.1368
R18710 bgr_11_0.cap_res2.t11 bgr_11_0.cap_res2.n0 0.00152174
R18711 bgr_11_0.cap_res2.t7 bgr_11_0.cap_res2.n1 0.00152174
R18712 bgr_11_0.cap_res2.t13 bgr_11_0.cap_res2.n2 0.00152174
R18713 bgr_11_0.cap_res2.t19 bgr_11_0.cap_res2.n3 0.00152174
R18714 bgr_11_0.cap_res2.t15 bgr_11_0.cap_res2.n4 0.00152174
R18715 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t6 447.279
R18716 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n0 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t2 446.967
R18717 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t7 446.967
R18718 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t5 446.967
R18719 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t3 344.772
R18720 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n8 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t4 281.168
R18721 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t9 281.168
R18722 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t8 281.168
R18723 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n8 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n7 205.946
R18724 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n6 205.946
R18725 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n7 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n4 165.8
R18726 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n9 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n8 165.8
R18727 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n10 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t1 108.615
R18728 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t0 108.615
R18729 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n6 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n5 63.4857
R18730 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n5 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n4 51.5193
R18731 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n10 15.6567
R18732 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n3 10.5317
R18733 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n10 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n9 6.0005
R18734 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n3 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n2 6.0005
R18735 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n9 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n4 0.313
R18736 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n2 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n1 0.313
R18737 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n1 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n0 0.313
R18738 a_3830_3166.t0 a_3830_3166.t1 169.905
R18739 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 172.969
R18740 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R18741 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 83.5719
R18742 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R18743 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R18744 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R18745 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 83.5719
R18746 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 83.5719
R18747 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 83.5719
R18748 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 83.5719
R18749 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 83.5719
R18750 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 83.5719
R18751 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 83.5719
R18752 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 83.5719
R18753 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 83.5719
R18754 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 83.5719
R18755 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 83.5719
R18756 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 83.5719
R18757 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 83.5719
R18758 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R18759 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R18760 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R18761 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 83.5719
R18762 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 73.8495
R18763 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.8495
R18764 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 73.3165
R18765 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 73.3165
R18766 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 73.3165
R18767 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 73.3165
R18768 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 73.3165
R18769 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.3165
R18770 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.19
R18771 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 73.19
R18772 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 73.19
R18773 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 73.19
R18774 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 73.19
R18775 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.19
R18776 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 65.0299
R18777 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 65.0299
R18778 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 26.074
R18779 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 26.074
R18780 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 26.074
R18781 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 26.074
R18782 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 26.074
R18783 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 26.074
R18784 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 26.074
R18785 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 26.074
R18786 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 25.7843
R18787 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 25.7843
R18788 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 25.7843
R18789 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 25.7843
R18790 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R18791 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 25.7843
R18792 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R18793 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R18794 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R18795 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 9.3005
R18796 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R18797 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R18798 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R18799 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 9.3005
R18800 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R18801 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R18802 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R18803 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R18804 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 9.3005
R18805 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 9.3005
R18806 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R18807 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R18808 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R18809 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R18810 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 9.3005
R18811 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R18812 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R18813 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 9.3005
R18814 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 9.3005
R18815 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R18816 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R18817 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 9.3005
R18818 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R18819 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 9.3005
R18820 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R18821 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R18822 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R18823 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 9.3005
R18824 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R18825 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R18826 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R18827 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 9.3005
R18828 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R18829 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R18830 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R18831 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R18832 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R18833 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R18834 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R18835 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R18836 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R18837 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R18838 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R18839 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R18840 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R18841 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 9.3005
R18842 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R18843 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 9.3005
R18844 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 9.3005
R18845 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 9.3005
R18846 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 4.64654
R18847 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 4.64654
R18848 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 4.64654
R18849 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 4.64654
R18850 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 4.64654
R18851 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 4.64654
R18852 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 4.64654
R18853 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 4.64654
R18854 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R18855 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 2.36206
R18856 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 2.36206
R18857 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 2.36206
R18858 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 2.36206
R18859 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 2.19742
R18860 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 2.19742
R18861 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 2.19742
R18862 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.19742
R18863 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 1.56363
R18864 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.56363
R18865 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 1.5505
R18866 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R18867 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R18868 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 1.5505
R18869 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 1.5505
R18870 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R18871 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 1.5505
R18872 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.5505
R18873 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 1.5505
R18874 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 1.5505
R18875 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 1.5505
R18876 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 1.5505
R18877 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 1.5505
R18878 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 1.5505
R18879 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.5505
R18880 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 1.5505
R18881 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.5505
R18882 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 1.5505
R18883 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.25468
R18884 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 1.25468
R18885 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.25468
R18886 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.25468
R18887 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 1.25468
R18888 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 1.25468
R18889 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 1.19225
R18890 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.19225
R18891 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 1.19225
R18892 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 1.19225
R18893 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.19225
R18894 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.19225
R18895 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 1.07024
R18896 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 1.07024
R18897 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R18898 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 1.07024
R18899 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R18900 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R18901 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 1.0237
R18902 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.0237
R18903 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 1.0237
R18904 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 1.0237
R18905 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.0237
R18906 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.0237
R18907 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.885803
R18908 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 0.885803
R18909 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 0.885803
R18910 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 0.885803
R18911 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.885803
R18912 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.885803
R18913 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R18914 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.885803
R18915 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 0.812055
R18916 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 0.812055
R18917 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.77514
R18918 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 0.77514
R18919 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.77514
R18920 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.77514
R18921 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 0.77514
R18922 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.77514
R18923 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R18924 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 0.77514
R18925 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.756696
R18926 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R18927 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.756696
R18928 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.756696
R18929 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R18930 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.756696
R18931 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R18932 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.756696
R18933 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 0.711459
R18934 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.711459
R18935 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.647417
R18936 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.647417
R18937 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R18938 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.590702
R18939 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.590702
R18940 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 0.590702
R18941 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.590702
R18942 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.590702
R18943 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.576566
R18944 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.576566
R18945 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 0.530034
R18946 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.530034
R18947 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 0.290206
R18948 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 0.290206
R18949 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 0.290206
R18950 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 0.290206
R18951 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 0.290206
R18952 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 0.290206
R18953 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 0.290206
R18954 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 0.290206
R18955 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R18956 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R18957 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R18958 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.203382
R18959 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.203382
R18960 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n141 0.203382
R18961 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 0.154071
R18962 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 0.154071
R18963 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 0.154071
R18964 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.154071
R18965 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 0.137464
R18966 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 0.137464
R18967 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 0.134964
R18968 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.134964
R18969 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R18970 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n140 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n139 0.0183571
R18971 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n138 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R18972 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R18973 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 0.0183571
R18974 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R18975 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R18976 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 0.0183571
R18977 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0183571
R18978 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R18979 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.0183571
R18980 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R18981 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.0183571
R18982 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 0.0183571
R18983 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R18984 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.0183571
R18985 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.0183571
R18986 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0183571
R18987 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 0.0106786
R18988 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.0106786
R18989 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.0106786
R18990 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 0.00992001
R18991 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 0.00992001
R18992 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R18993 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 0.00992001
R18994 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R18995 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 0.00992001
R18996 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R18997 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R18998 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.00992001
R18999 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.00992001
R19000 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R19001 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R19002 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R19003 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R19004 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00992001
R19005 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.00992001
R19006 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.00992001
R19007 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 0.00992001
R19008 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.00817857
R19009 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R19010 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 0.00817857
R19011 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.00817857
R19012 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.00817857
R19013 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t0 661.375
R19014 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n0 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t4 661.375
R19015 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t5 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n1 213.131
R19016 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t1 213.131
R19017 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t7 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t5 146.155
R19018 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t1 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t7 146.155
R19019 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t6 76.2576
R19020 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n2 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t3 76.2576
R19021 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n6 66.0338
R19022 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n8 66.0338
R19023 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n9 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n7 13.3963
R19024 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t8 11.2576
R19025 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n6 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t2 11.2576
R19026 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t10 11.2576
R19027 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n8 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t9 11.2576
R19028 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n9 6.72967
R19029 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n5 5.57862
R19030 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n0 5.1255
R19031 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n4 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n3 4.7505
R19032 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n5 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n4 4.5005
R19033 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n1 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n0 1.888
R19034 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n3 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n2 1.888
R19035 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n7 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n5 0.854667
R19036 VIN-.n0 VIN-.t7 1097.62
R19037 VIN- VIN-.n9 433.019
R19038 VIN-.n9 VIN-.t10 273.134
R19039 VIN-.n0 VIN-.t9 273.134
R19040 VIN-.n1 VIN-.t3 273.134
R19041 VIN-.n2 VIN-.t8 273.134
R19042 VIN-.n3 VIN-.t1 273.134
R19043 VIN-.n4 VIN-.t5 273.134
R19044 VIN-.n5 VIN-.t2 273.134
R19045 VIN-.n6 VIN-.t6 273.134
R19046 VIN-.n7 VIN-.t0 273.134
R19047 VIN-.n8 VIN-.t4 273.134
R19048 VIN-.n9 VIN-.n8 176.733
R19049 VIN-.n8 VIN-.n7 176.733
R19050 VIN-.n7 VIN-.n6 176.733
R19051 VIN-.n6 VIN-.n5 176.733
R19052 VIN-.n5 VIN-.n4 176.733
R19053 VIN-.n4 VIN-.n3 176.733
R19054 VIN-.n3 VIN-.n2 176.733
R19055 VIN-.n2 VIN-.n1 176.733
R19056 VIN-.n1 VIN-.n0 176.733
R19057 a_3110_6968.t0 a_3110_6968.t1 294.339
R19058 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t7 238.322
R19059 bgr_11_0.START_UP.n4 bgr_11_0.START_UP.t6 238.322
R19060 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n4 167.332
R19061 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t5 130.001
R19062 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n1 111.796
R19063 bgr_11_0.START_UP.n3 bgr_11_0.START_UP.n2 105.171
R19064 bgr_11_0.START_UP.n0 bgr_11_0.START_UP.t4 81.7074
R19065 bgr_11_0.START_UP bgr_11_0.START_UP.n0 36.8552
R19066 bgr_11_0.START_UP bgr_11_0.START_UP.n5 15.3755
R19067 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t0 13.1338
R19068 bgr_11_0.START_UP.n1 bgr_11_0.START_UP.t2 13.1338
R19069 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t1 13.1338
R19070 bgr_11_0.START_UP.n2 bgr_11_0.START_UP.t3 13.1338
R19071 bgr_11_0.START_UP.n5 bgr_11_0.START_UP.n3 4.21925
R19072 a_11420_30238.t0 a_11420_30238.t1 178.133
R19073 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.t8 539.797
R19074 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.n5 351.865
R19075 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.t6 117.817
R19076 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.n2 109.204
R19077 bgr_11_0.Vin-.n4 bgr_11_0.Vin-.n3 104.829
R19078 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n11 83.5719
R19079 bgr_11_0.Vin-.n1 bgr_11_0.Vin-.n0 83.5719
R19080 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n1 73.8495
R19081 bgr_11_0.Vin-.t7 bgr_11_0.Vin-.n10 65.0341
R19082 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.t5 39.4005
R19083 bgr_11_0.Vin-.n5 bgr_11_0.Vin-.t4 39.4005
R19084 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.n1 26.074
R19085 bgr_11_0.Vin-.n9 bgr_11_0.Vin-.n8 24.3755
R19086 bgr_11_0.Vin-.n8 bgr_11_0.Vin-.n7 17.6255
R19087 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t1 13.1338
R19088 bgr_11_0.Vin-.n3 bgr_11_0.Vin-.t2 13.1338
R19089 bgr_11_0.Vin-.n2 bgr_11_0.Vin-.t3 13.1338
R19090 bgr_11_0.Vin-.n2 bgr_11_0.Vin-.t0 13.1338
R19091 bgr_11_0.Vin-.n7 bgr_11_0.Vin-.n6 11.6567
R19092 bgr_11_0.Vin-.n6 bgr_11_0.Vin-.n4 3.8755
R19093 bgr_11_0.Vin-.n12 bgr_11_0.Vin-.n10 1.56483
R19094 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.n13 1.5505
R19095 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n0 0.885803
R19096 bgr_11_0.Vin-.n13 bgr_11_0.Vin-.n12 0.77514
R19097 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n0 0.756696
R19098 bgr_11_0.Vin-.n15 bgr_11_0.Vin-.n14 0.711459
R19099 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter bgr_11_0.Vin-.n15 0.576566
R19100 bgr_11_0.Vin-.n10 bgr_11_0.Vin-.n9 0.531499
R19101 bgr_11_0.Vin-.n11 bgr_11_0.Vin-.t7 0.290206
R19102 bgr_11_0.Vin-.n14 bgr_11_0.Vin-.n9 0.00817857
R19103 a_11950_28880.t0 a_11950_28880.t1 178.133
R19104 two_stage_opamp_dummy_magic_29_0.Vb2_2.n2 two_stage_opamp_dummy_magic_29_0.Vb2_2.t7 661.375
R19105 two_stage_opamp_dummy_magic_29_0.Vb2_2.n4 two_stage_opamp_dummy_magic_29_0.Vb2_2.t4 661.375
R19106 two_stage_opamp_dummy_magic_29_0.Vb2_2.t8 two_stage_opamp_dummy_magic_29_0.Vb2_2.n0 213.131
R19107 two_stage_opamp_dummy_magic_29_0.Vb2_2.n3 two_stage_opamp_dummy_magic_29_0.Vb2_2.t5 213.131
R19108 two_stage_opamp_dummy_magic_29_0.Vb2_2.n6 two_stage_opamp_dummy_magic_29_0.Vb2_2.n1 154.851
R19109 two_stage_opamp_dummy_magic_29_0.Vb2_2.t1 two_stage_opamp_dummy_magic_29_0.Vb2_2.t8 146.155
R19110 two_stage_opamp_dummy_magic_29_0.Vb2_2.t5 two_stage_opamp_dummy_magic_29_0.Vb2_2.t1 146.155
R19111 two_stage_opamp_dummy_magic_29_0.Vb2_2.t9 two_stage_opamp_dummy_magic_29_0.Vb2_2.n0 76.2576
R19112 two_stage_opamp_dummy_magic_29_0.Vb2_2.n3 two_stage_opamp_dummy_magic_29_0.Vb2_2.t6 76.2576
R19113 two_stage_opamp_dummy_magic_29_0.Vb2_2.n7 two_stage_opamp_dummy_magic_29_0.Vb2_2.n6 66.4503
R19114 two_stage_opamp_dummy_magic_29_0.Vb2_2.n1 two_stage_opamp_dummy_magic_29_0.Vb2_2.t3 21.8894
R19115 two_stage_opamp_dummy_magic_29_0.Vb2_2.n1 two_stage_opamp_dummy_magic_29_0.Vb2_2.t0 21.8894
R19116 two_stage_opamp_dummy_magic_29_0.Vb2_2.t9 two_stage_opamp_dummy_magic_29_0.Vb2_2.n7 11.2576
R19117 two_stage_opamp_dummy_magic_29_0.Vb2_2.n7 two_stage_opamp_dummy_magic_29_0.Vb2_2.t2 11.2576
R19118 two_stage_opamp_dummy_magic_29_0.Vb2_2.n5 two_stage_opamp_dummy_magic_29_0.Vb2_2.n4 5.1255
R19119 two_stage_opamp_dummy_magic_29_0.Vb2_2.n6 two_stage_opamp_dummy_magic_29_0.Vb2_2.n5 4.91195
R19120 two_stage_opamp_dummy_magic_29_0.Vb2_2.n5 two_stage_opamp_dummy_magic_29_0.Vb2_2.n2 4.7505
R19121 two_stage_opamp_dummy_magic_29_0.Vb2_2.n4 two_stage_opamp_dummy_magic_29_0.Vb2_2.n3 1.888
R19122 two_stage_opamp_dummy_magic_29_0.Vb2_2.n2 two_stage_opamp_dummy_magic_29_0.Vb2_2.n0 1.888
R19123 two_stage_opamp_dummy_magic_29_0.V_tot.n2 two_stage_opamp_dummy_magic_29_0.V_tot.t4 648.343
R19124 two_stage_opamp_dummy_magic_29_0.V_tot.n3 two_stage_opamp_dummy_magic_29_0.V_tot.t5 648.343
R19125 two_stage_opamp_dummy_magic_29_0.V_tot.n1 two_stage_opamp_dummy_magic_29_0.V_tot.t3 117.591
R19126 two_stage_opamp_dummy_magic_29_0.V_tot.n0 two_stage_opamp_dummy_magic_29_0.V_tot.t1 117.591
R19127 two_stage_opamp_dummy_magic_29_0.V_tot.n0 two_stage_opamp_dummy_magic_29_0.V_tot.t2 108.424
R19128 two_stage_opamp_dummy_magic_29_0.V_tot.n1 two_stage_opamp_dummy_magic_29_0.V_tot.t0 108.424
R19129 two_stage_opamp_dummy_magic_29_0.V_tot.n2 two_stage_opamp_dummy_magic_29_0.V_tot.n1 31.2036
R19130 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.V_tot.n0 29.5027
R19131 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.V_tot.n3 1.70362
R19132 two_stage_opamp_dummy_magic_29_0.V_tot.n3 two_stage_opamp_dummy_magic_29_0.V_tot.n2 0.84425
R19133 two_stage_opamp_dummy_magic_29_0.V_err_mir_p two_stage_opamp_dummy_magic_29_0.V_err_mir_p.n0 186.762
R19134 two_stage_opamp_dummy_magic_29_0.V_err_mir_p two_stage_opamp_dummy_magic_29_0.V_err_mir_p.n1 177.201
R19135 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t1 15.7605
R19136 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.n0 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t3 15.7605
R19137 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t2 15.7605
R19138 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.n1 two_stage_opamp_dummy_magic_29_0.V_err_mir_p.t0 15.7605
R19139 two_stage_opamp_dummy_magic_29_0.V_err_p.n1 two_stage_opamp_dummy_magic_29_0.V_err_p.n0 363.962
R19140 two_stage_opamp_dummy_magic_29_0.V_err_p.n0 two_stage_opamp_dummy_magic_29_0.V_err_p.t0 15.7605
R19141 two_stage_opamp_dummy_magic_29_0.V_err_p.n0 two_stage_opamp_dummy_magic_29_0.V_err_p.t3 15.7605
R19142 two_stage_opamp_dummy_magic_29_0.V_err_p.t2 two_stage_opamp_dummy_magic_29_0.V_err_p.n1 15.7605
R19143 two_stage_opamp_dummy_magic_29_0.V_err_p.n1 two_stage_opamp_dummy_magic_29_0.V_err_p.t1 15.7605
R19144 two_stage_opamp_dummy_magic_29_0.V_p_mir.n1 two_stage_opamp_dummy_magic_29_0.V_p_mir.n0 95.5151
R19145 two_stage_opamp_dummy_magic_29_0.V_p_mir.n0 two_stage_opamp_dummy_magic_29_0.V_p_mir.t0 16.0005
R19146 two_stage_opamp_dummy_magic_29_0.V_p_mir.n0 two_stage_opamp_dummy_magic_29_0.V_p_mir.t3 16.0005
R19147 two_stage_opamp_dummy_magic_29_0.V_p_mir.t2 two_stage_opamp_dummy_magic_29_0.V_p_mir.n1 9.6005
R19148 two_stage_opamp_dummy_magic_29_0.V_p_mir.n1 two_stage_opamp_dummy_magic_29_0.V_p_mir.t1 9.6005
R19149 a_11300_28630.t0 a_11300_28630.t1 178.133
R19150 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t1 99.8322
R19151 bgr_11_0.V_p_1.t0 bgr_11_0.V_p_1.n0 9.6005
R19152 bgr_11_0.V_p_1.n0 bgr_11_0.V_p_1.t2 9.6005
R19153 a_5700_30088.t0 a_5700_30088.t1 178.133
R19154 a_5820_28824.t0 a_5820_28824.t1 178.133
R19155 a_13940_3166.t0 a_13940_3166.t1 169.905
R19156 a_6470_28630.t0 a_6470_28630.t1 178.133
R19157 a_14420_6968.t0 a_14420_6968.t1 294.339
R19158 a_12070_30088.t0 a_12070_30088.t1 178.133
R19159 bgr_11_0.V_CUR_REF_REG bgr_11_0.V_CUR_REF_REG.t3 701.501
R19160 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.n0 357.647
R19161 bgr_11_0.V_CUR_REF_REG.n1 bgr_11_0.V_CUR_REF_REG.t2 135.239
R19162 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t0 39.4005
R19163 bgr_11_0.V_CUR_REF_REG.n0 bgr_11_0.V_CUR_REF_REG.t1 39.4005
R19164 bgr_11_0.V_CUR_REF_REG bgr_11_0.V_CUR_REF_REG.n1 5.79738
R19165 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t2 142.558
R19166 bgr_11_0.V_p_2.n0 bgr_11_0.V_p_2.t1 9.6005
R19167 bgr_11_0.V_p_2.t0 bgr_11_0.V_p_2.n0 9.6005
R19168 a_14540_6968.t0 a_14540_6968.t1 169.905
C0 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage VOUT+ 4.69775f
C1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 VOUT- 1.16944f
C2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 VDDA 9.28062f
C3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.V_err_gate 0.774203f
C4 m2_4090_7620# m2_4000_7510# 0.065657f
C5 two_stage_opamp_dummy_magic_29_0.V_tail_gate VOUT- 1.55445f
C6 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.163671f
C7 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.X 1.27179f
C8 bgr_11_0.PFET_GATE_10uA bgr_11_0.V_TOP 0.198366f
C9 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref bgr_11_0.V_CUR_REF_REG 2.48263f
C10 two_stage_opamp_dummy_magic_29_0.cap_res_X VDDA 1.32028f
C11 two_stage_opamp_dummy_magic_29_0.cap_res_Y two_stage_opamp_dummy_magic_29_0.cap_res_X 0.477735f
C12 two_stage_opamp_dummy_magic_29_0.VD3 VDDA 8.70244f
C13 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.cap_res_X 0.162723f
C14 bgr_11_0.START_UP_NFET1 VDDA 0.18791f
C15 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.V_source 0.040248f
C16 two_stage_opamp_dummy_magic_29_0.X two_stage_opamp_dummy_magic_29_0.cap_res_X 0.058941f
C17 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage VOUT- 4.67194f
C18 two_stage_opamp_dummy_magic_29_0.VD4 VDDA 8.70244f
C19 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 bgr_11_0.START_UP 0.011661f
C20 two_stage_opamp_dummy_magic_29_0.VD3 two_stage_opamp_dummy_magic_29_0.X 7.95637f
C21 two_stage_opamp_dummy_magic_29_0.VD4 two_stage_opamp_dummy_magic_29_0.cap_res_Y 0.168036f
C22 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.V_source 1.30282f
C23 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 VDDA 1.83425f
C24 bgr_11_0.Vin+ bgr_11_0.1st_Vout_1 0.275724f
C25 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 two_stage_opamp_dummy_magic_29_0.V_err_gate 0.274513f
C26 bgr_11_0.PFET_GATE_10uA VDDA 10.236f
C27 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.V_err_mir_p 0.047221f
C28 two_stage_opamp_dummy_magic_29_0.V_tail_gate VIN+ 0.060774f
C29 bgr_11_0.START_UP_NFET1 bgr_11_0.START_UP 0.145663f
C30 two_stage_opamp_dummy_magic_29_0.err_amp_out VDDA 0.228909f
C31 VIN+ VIN- 0.096614f
C32 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.err_amp_out 0.068782f
C33 two_stage_opamp_dummy_magic_29_0.cap_res_X VOUT+ 0.02055f
C34 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.V_tot 1.87985f
C35 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 0.939925f
C36 two_stage_opamp_dummy_magic_29_0.Y two_stage_opamp_dummy_magic_29_0.V_tot 0.803388f
C37 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 0.295226f
C38 two_stage_opamp_dummy_magic_29_0.err_amp_out two_stage_opamp_dummy_magic_29_0.X 1.31029f
C39 two_stage_opamp_dummy_magic_29_0.VD4 VOUT+ 0.034338f
C40 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.Y 2.31404f
C41 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.403953f
C42 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 VOUT- 0.666476f
C43 two_stage_opamp_dummy_magic_29_0.V_tail_gate VIN- 0.058275f
C44 bgr_11_0.V_TOP bgr_11_0.1st_Vout_1 2.62306f
C45 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage 5.93798f
C46 two_stage_opamp_dummy_magic_29_0.cap_res_X VOUT- 52.7123f
C47 two_stage_opamp_dummy_magic_29_0.VD3 VOUT- 0.027349f
C48 two_stage_opamp_dummy_magic_29_0.cap_res_Y two_stage_opamp_dummy_magic_29_0.V_source 0.066068f
C49 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 VOUT- 0.014192f
C50 bgr_11_0.1st_Vout_1 VDDA 2.66764f
C51 two_stage_opamp_dummy_magic_29_0.VD1 two_stage_opamp_dummy_magic_29_0.V_source 5.0157f
C52 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_29_0.V_err_amp_ref 0.792332f
C53 two_stage_opamp_dummy_magic_29_0.V_err_gate bgr_11_0.1st_Vout_1 0.131319f
C54 bgr_11_0.Vin+ bgr_11_0.V_TOP 1.8967f
C55 two_stage_opamp_dummy_magic_29_0.VD2 two_stage_opamp_dummy_magic_29_0.V_source 5.01421f
C56 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 3.24484f
C57 two_stage_opamp_dummy_magic_29_0.V_err_mir_p VDDA 0.661231f
C58 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.err_amp_out 0.158625f
C59 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_err_mir_p 0.429395f
C60 bgr_11_0.Vin+ bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 1.06291f
C61 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.456148f
C62 two_stage_opamp_dummy_magic_29_0.V_tot VDDA 0.140302f
C63 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_tot 0.611029f
C64 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 0.160792f
C65 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 two_stage_opamp_dummy_magic_29_0.cap_res_X 1.12766f
C66 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.VD1 0.222452f
C67 bgr_11_0.START_UP bgr_11_0.1st_Vout_1 0.13011f
C68 two_stage_opamp_dummy_magic_29_0.Vb1 VDDA 3.64542f
C69 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.cap_res_Y 0.238456f
C70 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.Vb1 1.79025f
C71 two_stage_opamp_dummy_magic_29_0.Y VDDA 7.31689f
C72 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.X 0.518118f
C73 two_stage_opamp_dummy_magic_29_0.Y two_stage_opamp_dummy_magic_29_0.cap_res_Y 0.058941f
C74 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.VD1 0.556757f
C75 bgr_11_0.Vin+ VDDA 1.72765f
C76 two_stage_opamp_dummy_magic_29_0.V_source VOUT+ 0.052538f
C77 bgr_11_0.Vin+ two_stage_opamp_dummy_magic_29_0.V_err_gate 0.066808f
C78 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.VD2 0.222452f
C79 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.X 2.28638f
C80 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.cap_res_X 2.021f
C81 two_stage_opamp_dummy_magic_29_0.Y two_stage_opamp_dummy_magic_29_0.X 0.056155f
C82 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.VD2 0.556757f
C83 two_stage_opamp_dummy_magic_29_0.Y two_stage_opamp_dummy_magic_29_0.VD2 4.15353f
C84 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 0.358499f
C85 two_stage_opamp_dummy_magic_29_0.V_tot VOUT+ 0.210263f
C86 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.573655f
C87 bgr_11_0.Vin+ bgr_11_0.START_UP 0.170134f
C88 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.V_TOP 0.04106f
C89 bgr_11_0.PFET_GATE_10uA bgr_11_0.V_CUR_REF_REG 0.344339f
C90 two_stage_opamp_dummy_magic_29_0.Vb1 VOUT+ 0.074784f
C91 two_stage_opamp_dummy_magic_29_0.V_source VOUT- 0.054787f
C92 two_stage_opamp_dummy_magic_29_0.Y VOUT+ 3.91972f
C93 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.err_amp_out 0.168894f
C94 bgr_11_0.V_TOP VDDA 16.3441f
C95 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_29_0.V_err_gate 0.103375f
C96 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.V_err_mir_p 0.047283f
C97 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter VDDA 0.023423f
C98 two_stage_opamp_dummy_magic_29_0.err_amp_out two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage 0.328005f
C99 two_stage_opamp_dummy_magic_29_0.V_tot VOUT- 0.210256f
C100 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.V_tot 1.21201f
C101 m2_4090_7620# VDDA 0.012155f
C102 two_stage_opamp_dummy_magic_29_0.Vb1 VOUT- 0.072458f
C103 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.Vb1 2.71797f
C104 two_stage_opamp_dummy_magic_29_0.V_source VIN+ 0.523933f
C105 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 two_stage_opamp_dummy_magic_29_0.cap_res_X 1.00943f
C106 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.Y 0.043425f
C107 two_stage_opamp_dummy_magic_29_0.VD3 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 0.421441f
C108 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref bgr_11_0.Vin+ 0.25235f
C109 two_stage_opamp_dummy_magic_29_0.cap_res_Y VDDA 1.28042f
C110 bgr_11_0.V_TOP bgr_11_0.START_UP 1.37378f
C111 two_stage_opamp_dummy_magic_29_0.V_err_gate VDDA 2.07498f
C112 two_stage_opamp_dummy_magic_29_0.X VDDA 7.32388f
C113 two_stage_opamp_dummy_magic_29_0.X two_stage_opamp_dummy_magic_29_0.VD1 4.15353f
C114 two_stage_opamp_dummy_magic_29_0.VD3 two_stage_opamp_dummy_magic_29_0.cap_res_X 0.167711f
C115 two_stage_opamp_dummy_magic_29_0.VD2 two_stage_opamp_dummy_magic_29_0.VD1 0.068381f
C116 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_source 3.43886f
C117 two_stage_opamp_dummy_magic_29_0.V_tot VIN+ 0.020171f
C118 bgr_11_0.START_UP VDDA 2.29043f
C119 two_stage_opamp_dummy_magic_29_0.V_err_gate bgr_11_0.START_UP 0.743841f
C120 two_stage_opamp_dummy_magic_29_0.V_source VIN- 0.524384f
C121 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 two_stage_opamp_dummy_magic_29_0.cap_res_X 0.063357f
C122 VDDA VOUT+ 13.9096f
C123 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 two_stage_opamp_dummy_magic_29_0.V_tot 0.438905f
C124 two_stage_opamp_dummy_magic_29_0.cap_res_Y VOUT+ 52.8086f
C125 two_stage_opamp_dummy_magic_29_0.V_source two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage 1.17205f
C126 bgr_11_0.PFET_GATE_10uA bgr_11_0.START_UP_NFET1 0.010791f
C127 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 0.146367f
C128 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref bgr_11_0.V_TOP 0.939477f
C129 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.V_tot 4.4704f
C130 two_stage_opamp_dummy_magic_29_0.V_source two_stage_opamp_dummy_magic_29_0.Vb1_2 0.443345f
C131 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.V_tail_gate 3.91616f
C132 two_stage_opamp_dummy_magic_29_0.V_tot VIN- 0.020171f
C133 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_29_0.Vb1 0.085081f
C134 bgr_11_0.Vin+ two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.014649f
C135 bgr_11_0.Vin+ bgr_11_0.V_CUR_REF_REG 1.57077f
C136 VDDA VOUT- 13.919099f
C137 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref VDDA 5.52057f
C138 two_stage_opamp_dummy_magic_29_0.cap_res_Y VOUT- 0.02055f
C139 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.cap_res_Y 0.143029f
C140 two_stage_opamp_dummy_magic_29_0.V_err_gate VOUT- 0.022304f
C141 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage 0.167852f
C142 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.V_err_gate 0.804531f
C143 two_stage_opamp_dummy_magic_29_0.X VOUT- 3.91972f
C144 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref two_stage_opamp_dummy_magic_29_0.X 0.010624f
C145 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.Vb1_2 2.00615f
C146 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 bgr_11_0.1st_Vout_1 1.93991f
C147 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref bgr_11_0.START_UP 1.39993f
C148 two_stage_opamp_dummy_magic_29_0.cap_res_X two_stage_opamp_dummy_magic_29_0.V_source 0.073057f
C149 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.028061f
C150 bgr_11_0.V_CUR_REF_REG bgr_11_0.V_TOP 0.308375f
C151 VOUT+ VOUT- 0.213277f
C152 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref VOUT+ 0.022237f
C153 two_stage_opamp_dummy_magic_29_0.VD2 VIN+ 0.532103f
C154 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 VDDA 4.0986f
C155 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter bgr_11_0.V_CUR_REF_REG 0.779503f
C156 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 0.733522f
C157 bgr_11_0.Vin+ two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 0.055084f
C158 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 two_stage_opamp_dummy_magic_29_0.X 0.90004f
C159 two_stage_opamp_dummy_magic_29_0.V_tail_gate VDDA 5.3725f
C160 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.cap_res_Y 2.02156f
C161 two_stage_opamp_dummy_magic_29_0.V_err_gate two_stage_opamp_dummy_magic_29_0.V_tail_gate 0.271999f
C162 bgr_11_0.V_CUR_REF_REG VDDA 3.71392f
C163 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.VD1 0.021061f
C164 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.cap_res_X 0.233991f
C165 bgr_11_0.V_CUR_REF_REG two_stage_opamp_dummy_magic_29_0.V_err_gate 0.375039f
C166 two_stage_opamp_dummy_magic_29_0.err_amp_out two_stage_opamp_dummy_magic_29_0.V_source 0.184635f
C167 two_stage_opamp_dummy_magic_29_0.V_tail_gate two_stage_opamp_dummy_magic_29_0.VD2 0.02134f
C168 two_stage_opamp_dummy_magic_29_0.VD1 VIN- 0.532103f
C169 two_stage_opamp_dummy_magic_29_0.VD4 two_stage_opamp_dummy_magic_29_0.Y 7.95637f
C170 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage VDDA 0.015355f
C171 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 two_stage_opamp_dummy_magic_29_0.Vb1 0.010591f
C172 bgr_11_0.PFET_GATE_10uA two_stage_opamp_dummy_magic_29_0.Vb1 0.129493f
C173 two_stage_opamp_dummy_magic_29_0.V_tot two_stage_opamp_dummy_magic_29_0.err_amp_out 3.37378f
C174 bgr_11_0.V_TOP two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 0.230311f
C175 two_stage_opamp_dummy_magic_29_0.V_tail_gate VOUT+ 1.55338f
C176 two_stage_opamp_dummy_magic_29_0.Vb1 two_stage_opamp_dummy_magic_29_0.err_amp_out 2.98002f
C177 VIN- GNDA 2.03908f
C178 VIN+ GNDA 2.04027f
C179 VOUT- GNDA 27.274624f
C180 VOUT+ GNDA 27.268608f
C181 VDDA GNDA 0.235252p
C182 m2_4000_7510# GNDA 0.039661f $ **FLOATING
C183 m2_4090_7620# GNDA 0.122312f $ **FLOATING
C184 two_stage_opamp_dummy_magic_29_0.Vb1_2 GNDA 2.88117f
C185 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage GNDA 10.256769f
C186 two_stage_opamp_dummy_magic_29_0.V_source GNDA 25.211973f
C187 two_stage_opamp_dummy_magic_29_0.VD1 GNDA 4.927533f
C188 two_stage_opamp_dummy_magic_29_0.VD2 GNDA 4.928203f
C189 two_stage_opamp_dummy_magic_29_0.cap_res_X GNDA 44.14486f
C190 two_stage_opamp_dummy_magic_29_0.cap_res_Y GNDA 44.14584f
C191 two_stage_opamp_dummy_magic_29_0.X GNDA 12.037578f
C192 two_stage_opamp_dummy_magic_29_0.err_amp_out GNDA 7.38754f
C193 two_stage_opamp_dummy_magic_29_0.V_err_mir_p GNDA 0.117954f
C194 two_stage_opamp_dummy_magic_29_0.V_tot GNDA 12.801761f
C195 two_stage_opamp_dummy_magic_29_0.Y GNDA 12.153778f
C196 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1 GNDA 13.922949f
C197 two_stage_opamp_dummy_magic_29_0.V_tail_gate GNDA 28.692923f
C198 two_stage_opamp_dummy_magic_29_0.Vb1 GNDA 36.095592f
C199 bgr_11_0.1st_Vout_1 GNDA 12.002972f
C200 bgr_11_0.START_UP GNDA 6.619071f
C201 bgr_11_0.START_UP_NFET1 GNDA 5.23862f
C202 two_stage_opamp_dummy_magic_29_0.V_err_gate GNDA 8.62121f
C203 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2 GNDA 18.00985f
C204 bgr_11_0.V_TOP GNDA 11.556623f
C205 bgr_11_0.V_CUR_REF_REG GNDA 4.852433f
C206 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 16.8453f
C207 bgr_11_0.Vin+ GNDA 4.646547f
C208 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref GNDA 9.27974f
C209 bgr_11_0.PFET_GATE_10uA GNDA 8.622524f
C210 two_stage_opamp_dummy_magic_29_0.VD3 GNDA 5.799711f
C211 two_stage_opamp_dummy_magic_29_0.VD4 GNDA 7.07405f
C212 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3 GNDA 2.394186f
C213 bgr_11_0.V_CUR_REF_REG.t3 GNDA 0.065688f
C214 bgr_11_0.V_CUR_REF_REG.t2 GNDA 0.445118f
C215 bgr_11_0.V_CUR_REF_REG.t0 GNDA 0.012849f
C216 bgr_11_0.V_CUR_REF_REG.t1 GNDA 0.012849f
C217 bgr_11_0.V_CUR_REF_REG.n0 GNDA 0.098435f
C218 bgr_11_0.V_CUR_REF_REG.n1 GNDA 5.0575f
C219 two_stage_opamp_dummy_magic_29_0.V_tot.t1 GNDA 0.164539f
C220 two_stage_opamp_dummy_magic_29_0.V_tot.t2 GNDA 0.154461f
C221 two_stage_opamp_dummy_magic_29_0.V_tot.n0 GNDA 1.65862f
C222 two_stage_opamp_dummy_magic_29_0.V_tot.t3 GNDA 0.164539f
C223 two_stage_opamp_dummy_magic_29_0.V_tot.t0 GNDA 0.154461f
C224 two_stage_opamp_dummy_magic_29_0.V_tot.n1 GNDA 1.74658f
C225 two_stage_opamp_dummy_magic_29_0.V_tot.t4 GNDA 0.046802f
C226 two_stage_opamp_dummy_magic_29_0.V_tot.n2 GNDA 1.83779f
C227 two_stage_opamp_dummy_magic_29_0.V_tot.t5 GNDA 0.046802f
C228 two_stage_opamp_dummy_magic_29_0.V_tot.n3 GNDA 0.322038f
C229 bgr_11_0.Vin-.n0 GNDA 0.07858f
C230 bgr_11_0.Vin-.n1 GNDA 0.356191f
C231 bgr_11_0.Vin-.t3 GNDA 0.030534f
C232 bgr_11_0.Vin-.t0 GNDA 0.030534f
C233 bgr_11_0.Vin-.n2 GNDA 0.085799f
C234 bgr_11_0.Vin-.t1 GNDA 0.030534f
C235 bgr_11_0.Vin-.t2 GNDA 0.030534f
C236 bgr_11_0.Vin-.n3 GNDA 0.074088f
C237 bgr_11_0.Vin-.n4 GNDA 0.633984f
C238 bgr_11_0.Vin-.t5 GNDA 0.010178f
C239 bgr_11_0.Vin-.t4 GNDA 0.010178f
C240 bgr_11_0.Vin-.n5 GNDA 0.031534f
C241 bgr_11_0.Vin-.n6 GNDA 0.428495f
C242 bgr_11_0.Vin-.t8 GNDA 0.049457f
C243 bgr_11_0.Vin-.n7 GNDA 0.623119f
C244 bgr_11_0.Vin-.t6 GNDA 0.128901f
C245 bgr_11_0.Vin-.n8 GNDA 0.734405f
C246 bgr_11_0.Vin-.n9 GNDA 1.36078f
C247 bgr_11_0.Vin-.n10 GNDA 0.531021f
C248 bgr_11_0.Vin-.t7 GNDA 0.294769f
C249 bgr_11_0.Vin-.n11 GNDA 0.078726f
C250 bgr_11_0.Vin-.n12 GNDA 0.134741f
C251 bgr_11_0.Vin-.n13 GNDA 0.079464f
C252 bgr_11_0.Vin-.n14 GNDA 0.652368f
C253 bgr_11_0.Vin-.n15 GNDA 0.403588f
C254 bgr_11_0.sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.097499f
C255 bgr_11_0.START_UP.t4 GNDA 1.72724f
C256 bgr_11_0.START_UP.t5 GNDA 0.045404f
C257 bgr_11_0.START_UP.n0 GNDA 1.15615f
C258 bgr_11_0.START_UP.t0 GNDA 0.04333f
C259 bgr_11_0.START_UP.t2 GNDA 0.04333f
C260 bgr_11_0.START_UP.n1 GNDA 0.135247f
C261 bgr_11_0.START_UP.t1 GNDA 0.04333f
C262 bgr_11_0.START_UP.t3 GNDA 0.04333f
C263 bgr_11_0.START_UP.n2 GNDA 0.106737f
C264 bgr_11_0.START_UP.n3 GNDA 1.0283f
C265 bgr_11_0.START_UP.t6 GNDA 0.016282f
C266 bgr_11_0.START_UP.t7 GNDA 0.016282f
C267 bgr_11_0.START_UP.n4 GNDA 0.046713f
C268 bgr_11_0.START_UP.n5 GNDA 0.477587f
C269 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t4 GNDA 0.038831f
C270 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n0 GNDA 0.08326f
C271 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t6 GNDA 0.078001f
C272 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n1 GNDA 0.249488f
C273 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t5 GNDA 0.186912f
C274 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t7 GNDA 0.146604f
C275 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t1 GNDA 0.186912f
C276 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t3 GNDA 0.078001f
C277 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n2 GNDA 0.249488f
C278 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t0 GNDA 0.038831f
C279 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n3 GNDA 0.08202f
C280 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n4 GNDA 0.040176f
C281 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n5 GNDA 0.062249f
C282 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t8 GNDA 0.021928f
C283 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t2 GNDA 0.021928f
C284 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n6 GNDA 0.044856f
C285 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n7 GNDA 0.16213f
C286 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t10 GNDA 0.021928f
C287 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.t9 GNDA 0.021928f
C288 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n8 GNDA 0.044856f
C289 two_stage_opamp_dummy_magic_29_0.Vb2_Vb3.n9 GNDA 0.210199f
C290 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t0 GNDA 0.245842f
C291 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t6 GNDA 0.773204f
C292 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t2 GNDA 0.772991f
C293 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n0 GNDA 0.636556f
C294 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t7 GNDA 0.772991f
C295 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n1 GNDA 0.331481f
C296 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t5 GNDA 0.772991f
C297 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n2 GNDA 0.667625f
C298 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n3 GNDA 0.790893f
C299 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t1 GNDA 0.245842f
C300 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n4 GNDA 0.431779f
C301 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t4 GNDA 0.667922f
C302 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t9 GNDA 0.667922f
C303 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t8 GNDA 0.667922f
C304 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.t3 GNDA 0.722234f
C305 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n5 GNDA 0.241787f
C306 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n6 GNDA 0.300709f
C307 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n7 GNDA 0.300709f
C308 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n8 GNDA 0.294161f
C309 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n9 GNDA 0.489447f
C310 two_stage_opamp_dummy_magic_29_0.V_b_2nd_stage.n10 GNDA 1.39879f
C311 bgr_11_0.cap_res2.t4 GNDA 0.334798f
C312 bgr_11_0.cap_res2.t10 GNDA 0.336011f
C313 bgr_11_0.cap_res2.t20 GNDA 0.318043f
C314 bgr_11_0.cap_res2.t9 GNDA 0.334798f
C315 bgr_11_0.cap_res2.t14 GNDA 0.336011f
C316 bgr_11_0.cap_res2.t5 GNDA 0.318043f
C317 bgr_11_0.cap_res2.t3 GNDA 0.334798f
C318 bgr_11_0.cap_res2.t8 GNDA 0.336011f
C319 bgr_11_0.cap_res2.t18 GNDA 0.318043f
C320 bgr_11_0.cap_res2.t16 GNDA 0.334798f
C321 bgr_11_0.cap_res2.t2 GNDA 0.336011f
C322 bgr_11_0.cap_res2.t12 GNDA 0.318043f
C323 bgr_11_0.cap_res2.t1 GNDA 0.334798f
C324 bgr_11_0.cap_res2.t6 GNDA 0.336011f
C325 bgr_11_0.cap_res2.t17 GNDA 0.318043f
C326 bgr_11_0.cap_res2.n0 GNDA 0.224415f
C327 bgr_11_0.cap_res2.t11 GNDA 0.178714f
C328 bgr_11_0.cap_res2.n1 GNDA 0.243496f
C329 bgr_11_0.cap_res2.t7 GNDA 0.178714f
C330 bgr_11_0.cap_res2.n2 GNDA 0.243496f
C331 bgr_11_0.cap_res2.t13 GNDA 0.178714f
C332 bgr_11_0.cap_res2.n3 GNDA 0.243496f
C333 bgr_11_0.cap_res2.t19 GNDA 0.178714f
C334 bgr_11_0.cap_res2.n4 GNDA 0.243496f
C335 bgr_11_0.cap_res2.t15 GNDA 0.360089f
C336 bgr_11_0.cap_res2.t0 GNDA 0.082395f
C337 two_stage_opamp_dummy_magic_29_0.VD1.t3 GNDA 0.033932f
C338 two_stage_opamp_dummy_magic_29_0.VD1.t10 GNDA 0.033932f
C339 two_stage_opamp_dummy_magic_29_0.VD1.n0 GNDA 0.075122f
C340 two_stage_opamp_dummy_magic_29_0.VD1.n1 GNDA 0.564997f
C341 two_stage_opamp_dummy_magic_29_0.VD1.n2 GNDA 0.050916f
C342 two_stage_opamp_dummy_magic_29_0.VD1.n3 GNDA 0.222536f
C343 two_stage_opamp_dummy_magic_29_0.VD1.t13 GNDA 0.033932f
C344 two_stage_opamp_dummy_magic_29_0.VD1.t20 GNDA 0.033932f
C345 two_stage_opamp_dummy_magic_29_0.VD1.n4 GNDA 0.073831f
C346 two_stage_opamp_dummy_magic_29_0.VD1.n5 GNDA 0.284467f
C347 two_stage_opamp_dummy_magic_29_0.VD1.n6 GNDA 0.072163f
C348 two_stage_opamp_dummy_magic_29_0.VD1.t17 GNDA 0.033932f
C349 two_stage_opamp_dummy_magic_29_0.VD1.t14 GNDA 0.033932f
C350 two_stage_opamp_dummy_magic_29_0.VD1.n7 GNDA 0.073831f
C351 two_stage_opamp_dummy_magic_29_0.VD1.n8 GNDA 0.292399f
C352 two_stage_opamp_dummy_magic_29_0.VD1.t2 GNDA 0.033932f
C353 two_stage_opamp_dummy_magic_29_0.VD1.t7 GNDA 0.033932f
C354 two_stage_opamp_dummy_magic_29_0.VD1.n9 GNDA 0.075122f
C355 two_stage_opamp_dummy_magic_29_0.VD1.t6 GNDA 0.033932f
C356 two_stage_opamp_dummy_magic_29_0.VD1.t11 GNDA 0.033932f
C357 two_stage_opamp_dummy_magic_29_0.VD1.n10 GNDA 0.075122f
C358 two_stage_opamp_dummy_magic_29_0.VD1.n11 GNDA 0.767242f
C359 two_stage_opamp_dummy_magic_29_0.VD1.t5 GNDA 0.033932f
C360 two_stage_opamp_dummy_magic_29_0.VD1.t9 GNDA 0.033932f
C361 two_stage_opamp_dummy_magic_29_0.VD1.n12 GNDA 0.075122f
C362 two_stage_opamp_dummy_magic_29_0.VD1.n13 GNDA 0.268181f
C363 two_stage_opamp_dummy_magic_29_0.VD1.t15 GNDA 0.033932f
C364 two_stage_opamp_dummy_magic_29_0.VD1.t12 GNDA 0.033932f
C365 two_stage_opamp_dummy_magic_29_0.VD1.n14 GNDA 0.073831f
C366 two_stage_opamp_dummy_magic_29_0.VD1.n15 GNDA 0.292399f
C367 two_stage_opamp_dummy_magic_29_0.VD1.n16 GNDA 0.122664f
C368 two_stage_opamp_dummy_magic_29_0.VD1.t19 GNDA 0.033932f
C369 two_stage_opamp_dummy_magic_29_0.VD1.t1 GNDA 0.033932f
C370 two_stage_opamp_dummy_magic_29_0.VD1.n17 GNDA 0.073831f
C371 two_stage_opamp_dummy_magic_29_0.VD1.n18 GNDA 0.284467f
C372 two_stage_opamp_dummy_magic_29_0.VD1.n19 GNDA 0.050916f
C373 two_stage_opamp_dummy_magic_29_0.VD1.n20 GNDA 0.222536f
C374 two_stage_opamp_dummy_magic_29_0.VD1.n21 GNDA 0.761461f
C375 two_stage_opamp_dummy_magic_29_0.VD1.n22 GNDA 0.114111f
C376 two_stage_opamp_dummy_magic_29_0.VD1.n23 GNDA 0.067863f
C377 two_stage_opamp_dummy_magic_29_0.VD1.t4 GNDA 0.033932f
C378 two_stage_opamp_dummy_magic_29_0.VD1.t8 GNDA 0.033932f
C379 two_stage_opamp_dummy_magic_29_0.VD1.n24 GNDA 0.075122f
C380 two_stage_opamp_dummy_magic_29_0.VD1.n25 GNDA 0.761461f
C381 two_stage_opamp_dummy_magic_29_0.VD1.n26 GNDA 0.114111f
C382 two_stage_opamp_dummy_magic_29_0.VD1.n27 GNDA 0.767242f
C383 two_stage_opamp_dummy_magic_29_0.VD1.n28 GNDA 0.268181f
C384 two_stage_opamp_dummy_magic_29_0.VD1.n29 GNDA 0.050916f
C385 two_stage_opamp_dummy_magic_29_0.VD1.t21 GNDA 0.033932f
C386 two_stage_opamp_dummy_magic_29_0.VD1.t18 GNDA 0.033932f
C387 two_stage_opamp_dummy_magic_29_0.VD1.n30 GNDA 0.073831f
C388 two_stage_opamp_dummy_magic_29_0.VD1.n31 GNDA 0.284467f
C389 two_stage_opamp_dummy_magic_29_0.VD1.n32 GNDA 0.122664f
C390 two_stage_opamp_dummy_magic_29_0.VD1.n33 GNDA 0.072163f
C391 two_stage_opamp_dummy_magic_29_0.VD1.t16 GNDA 0.033932f
C392 two_stage_opamp_dummy_magic_29_0.VD1.t0 GNDA 0.033932f
C393 two_stage_opamp_dummy_magic_29_0.VD1.n34 GNDA 0.073831f
C394 two_stage_opamp_dummy_magic_29_0.VD1.n35 GNDA 0.284467f
C395 two_stage_opamp_dummy_magic_29_0.VD1.n36 GNDA 0.050916f
C396 two_stage_opamp_dummy_magic_29_0.VD1.n37 GNDA 0.039407f
C397 two_stage_opamp_dummy_magic_29_0.Vb1_2.t2 GNDA 0.029732f
C398 two_stage_opamp_dummy_magic_29_0.Vb1_2.t4 GNDA 0.029732f
C399 two_stage_opamp_dummy_magic_29_0.Vb1_2.n0 GNDA 0.087151f
C400 two_stage_opamp_dummy_magic_29_0.Vb1_2.t0 GNDA 0.189479f
C401 two_stage_opamp_dummy_magic_29_0.Vb1_2.t3 GNDA 0.029732f
C402 two_stage_opamp_dummy_magic_29_0.Vb1_2.t1 GNDA 0.029732f
C403 two_stage_opamp_dummy_magic_29_0.Vb1_2.n1 GNDA 0.086354f
C404 two_stage_opamp_dummy_magic_29_0.err_amp_out.t5 GNDA 0.072503f
C405 two_stage_opamp_dummy_magic_29_0.err_amp_out.t4 GNDA 0.084623f
C406 two_stage_opamp_dummy_magic_29_0.err_amp_out.n0 GNDA 0.280015f
C407 two_stage_opamp_dummy_magic_29_0.err_amp_out.t3 GNDA 0.068078f
C408 two_stage_opamp_dummy_magic_29_0.err_amp_out.t1 GNDA 0.068078f
C409 two_stage_opamp_dummy_magic_29_0.err_amp_out.n1 GNDA 0.220809f
C410 two_stage_opamp_dummy_magic_29_0.err_amp_out.t2 GNDA 0.068078f
C411 two_stage_opamp_dummy_magic_29_0.err_amp_out.t0 GNDA 0.068078f
C412 two_stage_opamp_dummy_magic_29_0.err_amp_out.n2 GNDA 0.22061f
C413 two_stage_opamp_dummy_magic_29_0.err_amp_out.n3 GNDA 1.20062f
C414 two_stage_opamp_dummy_magic_29_0.V_err_gate.t1 GNDA 0.018464f
C415 two_stage_opamp_dummy_magic_29_0.V_err_gate.t2 GNDA 0.018464f
C416 two_stage_opamp_dummy_magic_29_0.V_err_gate.n0 GNDA 0.226134f
C417 two_stage_opamp_dummy_magic_29_0.V_err_gate.t0 GNDA 0.046159f
C418 two_stage_opamp_dummy_magic_29_0.V_err_gate.t4 GNDA 0.046159f
C419 two_stage_opamp_dummy_magic_29_0.V_err_gate.n1 GNDA 0.146296f
C420 two_stage_opamp_dummy_magic_29_0.V_err_gate.t7 GNDA 0.051544f
C421 two_stage_opamp_dummy_magic_29_0.V_err_gate.t9 GNDA 0.051544f
C422 two_stage_opamp_dummy_magic_29_0.V_err_gate.n2 GNDA 0.077423f
C423 two_stage_opamp_dummy_magic_29_0.V_err_gate.n3 GNDA 0.280869f
C424 two_stage_opamp_dummy_magic_29_0.V_err_gate.t3 GNDA 0.046159f
C425 two_stage_opamp_dummy_magic_29_0.V_err_gate.t5 GNDA 0.046159f
C426 two_stage_opamp_dummy_magic_29_0.V_err_gate.n4 GNDA 0.145699f
C427 two_stage_opamp_dummy_magic_29_0.V_err_gate.n5 GNDA 0.213743f
C428 two_stage_opamp_dummy_magic_29_0.V_err_gate.t6 GNDA 0.051544f
C429 two_stage_opamp_dummy_magic_29_0.V_err_gate.t8 GNDA 0.051544f
C430 two_stage_opamp_dummy_magic_29_0.V_err_gate.n6 GNDA 0.077423f
C431 bgr_11_0.Vin+.t5 GNDA 0.221779f
C432 bgr_11_0.Vin+.t0 GNDA 0.096124f
C433 bgr_11_0.Vin+.n0 GNDA 1.46352f
C434 bgr_11_0.Vin+.t1 GNDA 0.033039f
C435 bgr_11_0.Vin+.t4 GNDA 0.033039f
C436 bgr_11_0.Vin+.n1 GNDA 0.084276f
C437 bgr_11_0.Vin+.t3 GNDA 0.033039f
C438 bgr_11_0.Vin+.t2 GNDA 0.033039f
C439 bgr_11_0.Vin+.n2 GNDA 0.078979f
C440 bgr_11_0.Vin+.n3 GNDA 0.79622f
C441 bgr_11_0.Vin+.n4 GNDA 0.652102f
C442 bgr_11_0.Vin+.t6 GNDA 0.052809f
C443 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n0 GNDA 0.013013f
C444 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n1 GNDA 0.088324f
C445 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n2 GNDA 0.013768f
C446 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n3 GNDA 0.0946f
C447 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n4 GNDA 0.013013f
C448 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n5 GNDA 0.432823f
C449 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n7 GNDA 0.030586f
C450 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n8 GNDA 0.030586f
C451 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n11 GNDA 0.030586f
C452 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n12 GNDA 0.030586f
C453 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t10 GNDA 0.07743f
C454 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n13 GNDA 0.02905f
C455 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n14 GNDA 0.035605f
C456 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t8 GNDA 0.012744f
C457 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t1 GNDA 0.012744f
C458 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n15 GNDA 0.026057f
C459 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n16 GNDA 0.087236f
C460 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t5 GNDA 0.012744f
C461 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t0 GNDA 0.012744f
C462 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n17 GNDA 0.026057f
C463 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n18 GNDA 0.084286f
C464 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n19 GNDA 0.047895f
C465 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n20 GNDA 0.02905f
C466 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t4 GNDA 0.012744f
C467 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t9 GNDA 0.012744f
C468 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n21 GNDA 0.026057f
C469 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n22 GNDA 0.084286f
C470 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n23 GNDA 0.020865f
C471 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t7 GNDA 0.012744f
C472 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t3 GNDA 0.012744f
C473 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n24 GNDA 0.026057f
C474 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n25 GNDA 0.084286f
C475 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n26 GNDA 0.035605f
C476 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t6 GNDA 0.012744f
C477 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.t2 GNDA 0.012744f
C478 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n27 GNDA 0.026057f
C479 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n28 GNDA 0.085951f
C480 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n29 GNDA 0.116098f
C481 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n30 GNDA 0.772694f
C482 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n31 GNDA 0.185427f
C483 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n33 GNDA 0.030586f
C484 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n34 GNDA 0.030299f
C485 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n35 GNDA 0.043967f
C486 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n36 GNDA 0.043967f
C487 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n37 GNDA 0.030586f
C488 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n38 GNDA 0.030586f
C489 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n40 GNDA 2.62079f
C490 two_stage_opamp_dummy_magic_29_0.V_CMFB_S3.n41 GNDA 1.24119f
C491 bgr_11_0.V_CMFB_S3 GNDA 0.378144f
C492 two_stage_opamp_dummy_magic_29_0.VD3.n0 GNDA 1.11096f
C493 two_stage_opamp_dummy_magic_29_0.VD3.n1 GNDA 0.20151f
C494 two_stage_opamp_dummy_magic_29_0.VD3.n2 GNDA 0.378259f
C495 two_stage_opamp_dummy_magic_29_0.VD3.t35 GNDA 0.078836f
C496 two_stage_opamp_dummy_magic_29_0.VD3.n3 GNDA 0.149757f
C497 two_stage_opamp_dummy_magic_29_0.VD3.t28 GNDA 0.045031f
C498 two_stage_opamp_dummy_magic_29_0.VD3.t21 GNDA 0.045031f
C499 two_stage_opamp_dummy_magic_29_0.VD3.n4 GNDA 0.092115f
C500 two_stage_opamp_dummy_magic_29_0.VD3.n5 GNDA 0.260153f
C501 two_stage_opamp_dummy_magic_29_0.VD3.t26 GNDA 0.045031f
C502 two_stage_opamp_dummy_magic_29_0.VD3.t24 GNDA 0.045031f
C503 two_stage_opamp_dummy_magic_29_0.VD3.n6 GNDA 0.092115f
C504 two_stage_opamp_dummy_magic_29_0.VD3.n7 GNDA 0.25692f
C505 two_stage_opamp_dummy_magic_29_0.VD3.t5 GNDA 0.045031f
C506 two_stage_opamp_dummy_magic_29_0.VD3.t13 GNDA 0.045031f
C507 two_stage_opamp_dummy_magic_29_0.VD3.n8 GNDA 0.095624f
C508 two_stage_opamp_dummy_magic_29_0.VD3.t27 GNDA 0.045031f
C509 two_stage_opamp_dummy_magic_29_0.VD3.t31 GNDA 0.045031f
C510 two_stage_opamp_dummy_magic_29_0.VD3.n9 GNDA 0.092115f
C511 two_stage_opamp_dummy_magic_29_0.VD3.n10 GNDA 0.25692f
C512 two_stage_opamp_dummy_magic_29_0.VD3.t9 GNDA 0.045031f
C513 two_stage_opamp_dummy_magic_29_0.VD3.t17 GNDA 0.045031f
C514 two_stage_opamp_dummy_magic_29_0.VD3.n11 GNDA 0.095624f
C515 two_stage_opamp_dummy_magic_29_0.VD3.n12 GNDA 0.76157f
C516 two_stage_opamp_dummy_magic_29_0.VD3.t37 GNDA 0.160181f
C517 two_stage_opamp_dummy_magic_29_0.VD3.n13 GNDA 0.51334f
C518 two_stage_opamp_dummy_magic_29_0.VD3.t36 GNDA 0.383839f
C519 two_stage_opamp_dummy_magic_29_0.VD3.t18 GNDA 0.301063f
C520 two_stage_opamp_dummy_magic_29_0.VD3.t2 GNDA 0.301063f
C521 two_stage_opamp_dummy_magic_29_0.VD3.t12 GNDA 0.301063f
C522 two_stage_opamp_dummy_magic_29_0.VD3.t4 GNDA 0.301063f
C523 two_stage_opamp_dummy_magic_29_0.VD3.t16 GNDA 0.301063f
C524 two_stage_opamp_dummy_magic_29_0.VD3.t8 GNDA 0.301063f
C525 two_stage_opamp_dummy_magic_29_0.VD3.t14 GNDA 0.301063f
C526 two_stage_opamp_dummy_magic_29_0.VD3.t6 GNDA 0.301063f
C527 two_stage_opamp_dummy_magic_29_0.VD3.t0 GNDA 0.301063f
C528 two_stage_opamp_dummy_magic_29_0.VD3.t10 GNDA 0.301063f
C529 two_stage_opamp_dummy_magic_29_0.VD3.t33 GNDA 0.383839f
C530 two_stage_opamp_dummy_magic_29_0.VD3.t34 GNDA 0.160181f
C531 two_stage_opamp_dummy_magic_29_0.VD3.n14 GNDA 0.51334f
C532 two_stage_opamp_dummy_magic_29_0.VD3.t32 GNDA 0.078836f
C533 two_stage_opamp_dummy_magic_29_0.VD3.n15 GNDA 0.215181f
C534 two_stage_opamp_dummy_magic_29_0.VD3.t7 GNDA 0.045031f
C535 two_stage_opamp_dummy_magic_29_0.VD3.t15 GNDA 0.045031f
C536 two_stage_opamp_dummy_magic_29_0.VD3.n16 GNDA 0.095624f
C537 two_stage_opamp_dummy_magic_29_0.VD3.t29 GNDA 0.045031f
C538 two_stage_opamp_dummy_magic_29_0.VD3.t22 GNDA 0.045031f
C539 two_stage_opamp_dummy_magic_29_0.VD3.n17 GNDA 0.092115f
C540 two_stage_opamp_dummy_magic_29_0.VD3.n18 GNDA 0.25692f
C541 two_stage_opamp_dummy_magic_29_0.VD3.t11 GNDA 0.045031f
C542 two_stage_opamp_dummy_magic_29_0.VD3.t1 GNDA 0.045031f
C543 two_stage_opamp_dummy_magic_29_0.VD3.n19 GNDA 0.095624f
C544 two_stage_opamp_dummy_magic_29_0.VD3.n20 GNDA 0.115041f
C545 two_stage_opamp_dummy_magic_29_0.VD3.n21 GNDA 0.069429f
C546 two_stage_opamp_dummy_magic_29_0.VD3.t30 GNDA 0.045031f
C547 two_stage_opamp_dummy_magic_29_0.VD3.t23 GNDA 0.045031f
C548 two_stage_opamp_dummy_magic_29_0.VD3.n22 GNDA 0.092115f
C549 two_stage_opamp_dummy_magic_29_0.VD3.n23 GNDA 0.25692f
C550 two_stage_opamp_dummy_magic_29_0.VD3.n24 GNDA 0.069429f
C551 two_stage_opamp_dummy_magic_29_0.VD3.n25 GNDA 0.115041f
C552 two_stage_opamp_dummy_magic_29_0.VD3.t20 GNDA 0.045031f
C553 two_stage_opamp_dummy_magic_29_0.VD3.t25 GNDA 0.045031f
C554 two_stage_opamp_dummy_magic_29_0.VD3.n26 GNDA 0.092115f
C555 two_stage_opamp_dummy_magic_29_0.VD3.n27 GNDA 0.260153f
C556 two_stage_opamp_dummy_magic_29_0.VD3.n28 GNDA 0.76157f
C557 two_stage_opamp_dummy_magic_29_0.VD3.n29 GNDA 1.26178f
C558 two_stage_opamp_dummy_magic_29_0.VD3.n30 GNDA 0.432296f
C559 two_stage_opamp_dummy_magic_29_0.VD3.n31 GNDA 0.76157f
C560 two_stage_opamp_dummy_magic_29_0.VD3.t3 GNDA 0.045031f
C561 two_stage_opamp_dummy_magic_29_0.VD3.t19 GNDA 0.045031f
C562 two_stage_opamp_dummy_magic_29_0.VD3.n32 GNDA 0.095624f
C563 two_stage_opamp_dummy_magic_29_0.VD3.n33 GNDA 0.76157f
C564 two_stage_opamp_dummy_magic_29_0.VD3.n34 GNDA 0.342878f
C565 bgr_11_0.cap_res1.t6 GNDA 0.339883f
C566 bgr_11_0.cap_res1.t18 GNDA 0.357788f
C567 bgr_11_0.cap_res1.t10 GNDA 0.359085f
C568 bgr_11_0.cap_res1.t13 GNDA 0.339883f
C569 bgr_11_0.cap_res1.t20 GNDA 0.357788f
C570 bgr_11_0.cap_res1.t17 GNDA 0.359085f
C571 bgr_11_0.cap_res1.t5 GNDA 0.339883f
C572 bgr_11_0.cap_res1.t16 GNDA 0.357788f
C573 bgr_11_0.cap_res1.t9 GNDA 0.359085f
C574 bgr_11_0.cap_res1.t1 GNDA 0.339883f
C575 bgr_11_0.cap_res1.t8 GNDA 0.357788f
C576 bgr_11_0.cap_res1.t2 GNDA 0.359085f
C577 bgr_11_0.cap_res1.t3 GNDA 0.339883f
C578 bgr_11_0.cap_res1.t15 GNDA 0.357788f
C579 bgr_11_0.cap_res1.t7 GNDA 0.359085f
C580 bgr_11_0.cap_res1.n0 GNDA 0.239826f
C581 bgr_11_0.cap_res1.t11 GNDA 0.190986f
C582 bgr_11_0.cap_res1.n1 GNDA 0.260216f
C583 bgr_11_0.cap_res1.t4 GNDA 0.190986f
C584 bgr_11_0.cap_res1.n2 GNDA 0.260216f
C585 bgr_11_0.cap_res1.t12 GNDA 0.190986f
C586 bgr_11_0.cap_res1.n3 GNDA 0.260216f
C587 bgr_11_0.cap_res1.t19 GNDA 0.190986f
C588 bgr_11_0.cap_res1.n4 GNDA 0.260216f
C589 bgr_11_0.cap_res1.t14 GNDA 0.383393f
C590 bgr_11_0.cap_res1.t0 GNDA 0.088196f
C591 bgr_11_0.1st_Vout_1.n0 GNDA 0.191219f
C592 bgr_11_0.1st_Vout_1.t27 GNDA 0.240973f
C593 bgr_11_0.1st_Vout_1.t18 GNDA 0.236938f
C594 bgr_11_0.1st_Vout_1.t14 GNDA 0.240973f
C595 bgr_11_0.1st_Vout_1.t23 GNDA 0.236938f
C596 bgr_11_0.1st_Vout_1.n1 GNDA 0.158859f
C597 bgr_11_0.1st_Vout_1.n2 GNDA 0.203285f
C598 bgr_11_0.1st_Vout_1.t32 GNDA 0.240973f
C599 bgr_11_0.1st_Vout_1.t26 GNDA 0.236938f
C600 bgr_11_0.1st_Vout_1.t22 GNDA 0.240973f
C601 bgr_11_0.1st_Vout_1.t31 GNDA 0.236938f
C602 bgr_11_0.1st_Vout_1.n3 GNDA 0.158859f
C603 bgr_11_0.1st_Vout_1.n4 GNDA 0.247711f
C604 bgr_11_0.1st_Vout_1.t25 GNDA 0.240973f
C605 bgr_11_0.1st_Vout_1.t17 GNDA 0.236938f
C606 bgr_11_0.1st_Vout_1.t12 GNDA 0.240973f
C607 bgr_11_0.1st_Vout_1.t21 GNDA 0.236938f
C608 bgr_11_0.1st_Vout_1.n5 GNDA 0.158859f
C609 bgr_11_0.1st_Vout_1.n6 GNDA 0.247711f
C610 bgr_11_0.1st_Vout_1.t16 GNDA 0.240973f
C611 bgr_11_0.1st_Vout_1.t8 GNDA 0.236938f
C612 bgr_11_0.1st_Vout_1.t7 GNDA 0.240973f
C613 bgr_11_0.1st_Vout_1.t11 GNDA 0.236938f
C614 bgr_11_0.1st_Vout_1.n7 GNDA 0.158859f
C615 bgr_11_0.1st_Vout_1.n8 GNDA 0.247711f
C616 bgr_11_0.1st_Vout_1.t24 GNDA 0.240973f
C617 bgr_11_0.1st_Vout_1.t15 GNDA 0.236938f
C618 bgr_11_0.1st_Vout_1.n9 GNDA 0.203285f
C619 bgr_11_0.1st_Vout_1.t20 GNDA 0.236938f
C620 bgr_11_0.1st_Vout_1.n10 GNDA 0.10366f
C621 bgr_11_0.1st_Vout_1.t9 GNDA 0.236938f
C622 bgr_11_0.1st_Vout_1.n11 GNDA 2.00975f
C623 bgr_11_0.1st_Vout_1.t29 GNDA 0.01424f
C624 bgr_11_0.1st_Vout_1.n12 GNDA 3.07165f
C625 bgr_11_0.1st_Vout_1.n13 GNDA 0.012548f
C626 bgr_11_0.1st_Vout_1.n14 GNDA 0.191219f
C627 bgr_11_0.1st_Vout_1.n15 GNDA 0.017467f
C628 bgr_11_0.1st_Vout_1.n16 GNDA 0.173289f
C629 bgr_11_0.1st_Vout_1.n17 GNDA 0.012189f
C630 bgr_11_0.1st_Vout_1.t3 GNDA 0.054022f
C631 bgr_11_0.1st_Vout_1.n18 GNDA 0.173688f
C632 bgr_11_0.1st_Vout_1.n19 GNDA 0.127946f
C633 bgr_11_0.1st_Vout_1.n20 GNDA 0.017467f
C634 bgr_11_0.1st_Vout_1.n21 GNDA 0.173289f
C635 bgr_11_0.1st_Vout_1.n22 GNDA 0.012548f
C636 bgr_11_0.1st_Vout_1.t13 GNDA 0.013988f
C637 two_stage_opamp_dummy_magic_29_0.VD2.t13 GNDA 0.033932f
C638 two_stage_opamp_dummy_magic_29_0.VD2.t8 GNDA 0.033932f
C639 two_stage_opamp_dummy_magic_29_0.VD2.n0 GNDA 0.075122f
C640 two_stage_opamp_dummy_magic_29_0.VD2.n1 GNDA 0.564997f
C641 two_stage_opamp_dummy_magic_29_0.VD2.n2 GNDA 0.050916f
C642 two_stage_opamp_dummy_magic_29_0.VD2.n3 GNDA 0.222536f
C643 two_stage_opamp_dummy_magic_29_0.VD2.t6 GNDA 0.033932f
C644 two_stage_opamp_dummy_magic_29_0.VD2.t4 GNDA 0.033932f
C645 two_stage_opamp_dummy_magic_29_0.VD2.n4 GNDA 0.073831f
C646 two_stage_opamp_dummy_magic_29_0.VD2.n5 GNDA 0.284467f
C647 two_stage_opamp_dummy_magic_29_0.VD2.n6 GNDA 0.072163f
C648 two_stage_opamp_dummy_magic_29_0.VD2.t7 GNDA 0.033932f
C649 two_stage_opamp_dummy_magic_29_0.VD2.t20 GNDA 0.033932f
C650 two_stage_opamp_dummy_magic_29_0.VD2.n7 GNDA 0.073831f
C651 two_stage_opamp_dummy_magic_29_0.VD2.n8 GNDA 0.292399f
C652 two_stage_opamp_dummy_magic_29_0.VD2.t10 GNDA 0.033932f
C653 two_stage_opamp_dummy_magic_29_0.VD2.t16 GNDA 0.033932f
C654 two_stage_opamp_dummy_magic_29_0.VD2.n9 GNDA 0.075122f
C655 two_stage_opamp_dummy_magic_29_0.VD2.t14 GNDA 0.033932f
C656 two_stage_opamp_dummy_magic_29_0.VD2.t9 GNDA 0.033932f
C657 two_stage_opamp_dummy_magic_29_0.VD2.n10 GNDA 0.075122f
C658 two_stage_opamp_dummy_magic_29_0.VD2.n11 GNDA 0.767242f
C659 two_stage_opamp_dummy_magic_29_0.VD2.t12 GNDA 0.033932f
C660 two_stage_opamp_dummy_magic_29_0.VD2.t15 GNDA 0.033932f
C661 two_stage_opamp_dummy_magic_29_0.VD2.n12 GNDA 0.075122f
C662 two_stage_opamp_dummy_magic_29_0.VD2.n13 GNDA 0.268181f
C663 two_stage_opamp_dummy_magic_29_0.VD2.t19 GNDA 0.033932f
C664 two_stage_opamp_dummy_magic_29_0.VD2.t18 GNDA 0.033932f
C665 two_stage_opamp_dummy_magic_29_0.VD2.n14 GNDA 0.073831f
C666 two_stage_opamp_dummy_magic_29_0.VD2.n15 GNDA 0.292399f
C667 two_stage_opamp_dummy_magic_29_0.VD2.n16 GNDA 0.122664f
C668 two_stage_opamp_dummy_magic_29_0.VD2.t21 GNDA 0.033932f
C669 two_stage_opamp_dummy_magic_29_0.VD2.t0 GNDA 0.033932f
C670 two_stage_opamp_dummy_magic_29_0.VD2.n17 GNDA 0.073831f
C671 two_stage_opamp_dummy_magic_29_0.VD2.n18 GNDA 0.284467f
C672 two_stage_opamp_dummy_magic_29_0.VD2.n19 GNDA 0.050916f
C673 two_stage_opamp_dummy_magic_29_0.VD2.n20 GNDA 0.222536f
C674 two_stage_opamp_dummy_magic_29_0.VD2.n21 GNDA 0.761461f
C675 two_stage_opamp_dummy_magic_29_0.VD2.n22 GNDA 0.114111f
C676 two_stage_opamp_dummy_magic_29_0.VD2.n23 GNDA 0.067863f
C677 two_stage_opamp_dummy_magic_29_0.VD2.t11 GNDA 0.033932f
C678 two_stage_opamp_dummy_magic_29_0.VD2.t17 GNDA 0.033932f
C679 two_stage_opamp_dummy_magic_29_0.VD2.n24 GNDA 0.075122f
C680 two_stage_opamp_dummy_magic_29_0.VD2.n25 GNDA 0.761461f
C681 two_stage_opamp_dummy_magic_29_0.VD2.n26 GNDA 0.114111f
C682 two_stage_opamp_dummy_magic_29_0.VD2.n27 GNDA 0.767242f
C683 two_stage_opamp_dummy_magic_29_0.VD2.n28 GNDA 0.268181f
C684 two_stage_opamp_dummy_magic_29_0.VD2.n29 GNDA 0.050916f
C685 two_stage_opamp_dummy_magic_29_0.VD2.t1 GNDA 0.033932f
C686 two_stage_opamp_dummy_magic_29_0.VD2.t3 GNDA 0.033932f
C687 two_stage_opamp_dummy_magic_29_0.VD2.n30 GNDA 0.073831f
C688 two_stage_opamp_dummy_magic_29_0.VD2.n31 GNDA 0.284467f
C689 two_stage_opamp_dummy_magic_29_0.VD2.n32 GNDA 0.122664f
C690 two_stage_opamp_dummy_magic_29_0.VD2.n33 GNDA 0.072163f
C691 two_stage_opamp_dummy_magic_29_0.VD2.t5 GNDA 0.033932f
C692 two_stage_opamp_dummy_magic_29_0.VD2.t2 GNDA 0.033932f
C693 two_stage_opamp_dummy_magic_29_0.VD2.n34 GNDA 0.073831f
C694 two_stage_opamp_dummy_magic_29_0.VD2.n35 GNDA 0.284467f
C695 two_stage_opamp_dummy_magic_29_0.VD2.n36 GNDA 0.050916f
C696 two_stage_opamp_dummy_magic_29_0.VD2.n37 GNDA 0.039407f
C697 two_stage_opamp_dummy_magic_29_0.Vb1.n0 GNDA 1.31165f
C698 two_stage_opamp_dummy_magic_29_0.Vb1.n1 GNDA 0.163394f
C699 two_stage_opamp_dummy_magic_29_0.Vb1.n2 GNDA 1.38887f
C700 two_stage_opamp_dummy_magic_29_0.Vb1.n3 GNDA 0.338122f
C701 two_stage_opamp_dummy_magic_29_0.Vb1.n4 GNDA 0.398987f
C702 two_stage_opamp_dummy_magic_29_0.Vb1.n5 GNDA 0.338122f
C703 two_stage_opamp_dummy_magic_29_0.Vb1.n6 GNDA 1.2198f
C704 two_stage_opamp_dummy_magic_29_0.Vb1.n7 GNDA 0.229926f
C705 two_stage_opamp_dummy_magic_29_0.Vb1.t20 GNDA 0.033142f
C706 two_stage_opamp_dummy_magic_29_0.Vb1.t4 GNDA 0.021513f
C707 two_stage_opamp_dummy_magic_29_0.Vb1.t0 GNDA 0.027903f
C708 two_stage_opamp_dummy_magic_29_0.Vb1.n8 GNDA 0.028688f
C709 two_stage_opamp_dummy_magic_29_0.Vb1.t2 GNDA 0.021513f
C710 two_stage_opamp_dummy_magic_29_0.Vb1.t6 GNDA 0.027903f
C711 two_stage_opamp_dummy_magic_29_0.Vb1.n9 GNDA 0.028688f
C712 two_stage_opamp_dummy_magic_29_0.Vb1.n10 GNDA 0.021384f
C713 two_stage_opamp_dummy_magic_29_0.Vb1.t5 GNDA 0.020988f
C714 two_stage_opamp_dummy_magic_29_0.Vb1.t3 GNDA 0.020988f
C715 two_stage_opamp_dummy_magic_29_0.Vb1.n11 GNDA 0.045667f
C716 two_stage_opamp_dummy_magic_29_0.Vb1.t13 GNDA 0.653332f
C717 two_stage_opamp_dummy_magic_29_0.Vb1.n12 GNDA 0.076804f
C718 two_stage_opamp_dummy_magic_29_0.Vb1.t30 GNDA 0.033142f
C719 two_stage_opamp_dummy_magic_29_0.Vb1.t19 GNDA 0.033142f
C720 two_stage_opamp_dummy_magic_29_0.Vb1.t28 GNDA 0.033142f
C721 two_stage_opamp_dummy_magic_29_0.Vb1.t16 GNDA 0.033142f
C722 two_stage_opamp_dummy_magic_29_0.Vb1.t29 GNDA 0.033142f
C723 two_stage_opamp_dummy_magic_29_0.Vb1.t17 GNDA 0.033142f
C724 two_stage_opamp_dummy_magic_29_0.Vb1.t27 GNDA 0.033142f
C725 two_stage_opamp_dummy_magic_29_0.Vb1.t14 GNDA 0.033142f
C726 two_stage_opamp_dummy_magic_29_0.Vb1.t21 GNDA 0.033142f
C727 two_stage_opamp_dummy_magic_29_0.Vb1.n13 GNDA 1.25008f
C728 two_stage_opamp_dummy_magic_29_0.Vb1.t11 GNDA 0.020988f
C729 two_stage_opamp_dummy_magic_29_0.Vb1.t1 GNDA 0.020988f
C730 two_stage_opamp_dummy_magic_29_0.Vb1.n14 GNDA 0.045667f
C731 two_stage_opamp_dummy_magic_29_0.Vb1.n15 GNDA 0.171661f
C732 two_stage_opamp_dummy_magic_29_0.Vb1.n16 GNDA 0.168468f
C733 two_stage_opamp_dummy_magic_29_0.Vb1.t7 GNDA 0.020988f
C734 two_stage_opamp_dummy_magic_29_0.Vb1.t10 GNDA 0.020988f
C735 two_stage_opamp_dummy_magic_29_0.Vb1.n17 GNDA 0.045667f
C736 two_stage_opamp_dummy_magic_29_0.Vb1.n18 GNDA 0.171661f
C737 two_stage_opamp_dummy_magic_29_0.Vb1.t15 GNDA 0.033142f
C738 two_stage_opamp_dummy_magic_29_0.Vb1.t26 GNDA 0.033142f
C739 two_stage_opamp_dummy_magic_29_0.Vb1.t12 GNDA 0.033142f
C740 two_stage_opamp_dummy_magic_29_0.Vb1.t25 GNDA 0.033142f
C741 two_stage_opamp_dummy_magic_29_0.Vb1.t32 GNDA 0.033142f
C742 two_stage_opamp_dummy_magic_29_0.Vb1.t23 GNDA 0.033142f
C743 two_stage_opamp_dummy_magic_29_0.Vb1.t18 GNDA 0.033142f
C744 two_stage_opamp_dummy_magic_29_0.Vb1.t24 GNDA 0.033142f
C745 two_stage_opamp_dummy_magic_29_0.Vb1.t31 GNDA 0.033142f
C746 two_stage_opamp_dummy_magic_29_0.Vb1.t22 GNDA 0.033142f
C747 two_stage_opamp_dummy_magic_29_0.Vb1.t9 GNDA 0.027984f
C748 two_stage_opamp_dummy_magic_29_0.Vb1.t8 GNDA 0.027984f
C749 two_stage_opamp_dummy_magic_29_0.Vb1.n19 GNDA 0.063321f
C750 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t6 GNDA 0.339505f
C751 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t7 GNDA 0.107388f
C752 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n0 GNDA 3.49192f
C753 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t4 GNDA 0.064242f
C754 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t1 GNDA 0.064242f
C755 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n1 GNDA 0.179204f
C756 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t3 GNDA 0.064242f
C757 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t0 GNDA 0.064242f
C758 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n2 GNDA 0.161296f
C759 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n3 GNDA 1.98079f
C760 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t2 GNDA 0.064242f
C761 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t5 GNDA 0.064242f
C762 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n4 GNDA 0.161296f
C763 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n5 GNDA 1.47273f
C764 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n6 GNDA 0.939954f
C765 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t9 GNDA 0.073772f
C766 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.t8 GNDA 0.072531f
C767 two_stage_opamp_dummy_magic_29_0.V_err_amp_ref.n7 GNDA 0.525625f
C768 bgr_11_0.V_TOP.n0 GNDA 0.016831f
C769 bgr_11_0.V_TOP.t29 GNDA 0.128711f
C770 bgr_11_0.V_TOP.t37 GNDA 0.128973f
C771 bgr_11_0.V_TOP.t38 GNDA 0.129529f
C772 bgr_11_0.V_TOP.n1 GNDA 0.162971f
C773 bgr_11_0.V_TOP.t23 GNDA 0.129529f
C774 bgr_11_0.V_TOP.n2 GNDA 0.089272f
C775 bgr_11_0.V_TOP.t48 GNDA 0.129529f
C776 bgr_11_0.V_TOP.n3 GNDA 0.089272f
C777 bgr_11_0.V_TOP.t39 GNDA 0.129529f
C778 bgr_11_0.V_TOP.n4 GNDA 0.089272f
C779 bgr_11_0.V_TOP.t27 GNDA 0.129529f
C780 bgr_11_0.V_TOP.n5 GNDA 0.089272f
C781 bgr_11_0.V_TOP.n6 GNDA 0.025246f
C782 bgr_11_0.V_TOP.n7 GNDA 0.057364f
C783 bgr_11_0.V_TOP.t13 GNDA 0.129887f
C784 bgr_11_0.V_TOP.t20 GNDA 0.374019f
C785 bgr_11_0.V_TOP.t24 GNDA 0.38039f
C786 bgr_11_0.V_TOP.t32 GNDA 0.374019f
C787 bgr_11_0.V_TOP.n8 GNDA 0.250768f
C788 bgr_11_0.V_TOP.t19 GNDA 0.374019f
C789 bgr_11_0.V_TOP.t46 GNDA 0.38039f
C790 bgr_11_0.V_TOP.n9 GNDA 0.320897f
C791 bgr_11_0.V_TOP.t34 GNDA 0.38039f
C792 bgr_11_0.V_TOP.t40 GNDA 0.374019f
C793 bgr_11_0.V_TOP.n10 GNDA 0.250768f
C794 bgr_11_0.V_TOP.t31 GNDA 0.374019f
C795 bgr_11_0.V_TOP.t18 GNDA 0.38039f
C796 bgr_11_0.V_TOP.n11 GNDA 0.391025f
C797 bgr_11_0.V_TOP.t22 GNDA 0.38039f
C798 bgr_11_0.V_TOP.t30 GNDA 0.374019f
C799 bgr_11_0.V_TOP.n12 GNDA 0.250768f
C800 bgr_11_0.V_TOP.t17 GNDA 0.374019f
C801 bgr_11_0.V_TOP.t44 GNDA 0.38039f
C802 bgr_11_0.V_TOP.n13 GNDA 0.391025f
C803 bgr_11_0.V_TOP.t47 GNDA 0.38039f
C804 bgr_11_0.V_TOP.t16 GNDA 0.374019f
C805 bgr_11_0.V_TOP.n14 GNDA 0.250768f
C806 bgr_11_0.V_TOP.t43 GNDA 0.374019f
C807 bgr_11_0.V_TOP.t35 GNDA 0.38039f
C808 bgr_11_0.V_TOP.n15 GNDA 0.391025f
C809 bgr_11_0.V_TOP.t41 GNDA 0.38039f
C810 bgr_11_0.V_TOP.t15 GNDA 0.374019f
C811 bgr_11_0.V_TOP.n16 GNDA 0.320897f
C812 bgr_11_0.V_TOP.t28 GNDA 0.374019f
C813 bgr_11_0.V_TOP.n17 GNDA 0.163634f
C814 bgr_11_0.V_TOP.n18 GNDA 0.875119f
C815 bgr_11_0.V_TOP.t0 GNDA 0.105245f
C816 bgr_11_0.V_TOP.n19 GNDA 1.42428f
C817 bgr_11_0.V_TOP.n20 GNDA 0.019145f
C818 bgr_11_0.V_TOP.n21 GNDA 0.024925f
C819 bgr_11_0.V_TOP.n22 GNDA 0.022551f
C820 bgr_11_0.V_TOP.n23 GNDA 0.25922f
C821 bgr_11_0.V_TOP.n24 GNDA 0.158514f
C822 bgr_11_0.V_TOP.n25 GNDA 0.655866f
C823 bgr_11_0.V_TOP.n26 GNDA 0.020198f
C824 bgr_11_0.V_TOP.n27 GNDA 0.198604f
C825 bgr_11_0.V_TOP.n28 GNDA 0.020198f
C826 bgr_11_0.V_TOP.n29 GNDA 0.204214f
C827 bgr_11_0.V_TOP.n30 GNDA 0.020198f
C828 bgr_11_0.V_TOP.n31 GNDA 0.190361f
C829 bgr_11_0.V_TOP.n32 GNDA 0.391697f
C830 bgr_11_0.V_TOP.n33 GNDA 0.089765f
C831 bgr_11_0.V_TOP.t14 GNDA 0.127788f
C832 bgr_11_0.V_TOP.n34 GNDA 0.052677f
C833 bgr_11_0.V_TOP.n35 GNDA 0.025246f
C834 bgr_11_0.V_TOP.t45 GNDA 0.128533f
C835 bgr_11_0.V_TOP.n36 GNDA 0.084658f
C836 bgr_11_0.V_TOP.t36 GNDA 0.129529f
C837 bgr_11_0.V_TOP.n37 GNDA 0.089272f
C838 bgr_11_0.V_TOP.t25 GNDA 0.129529f
C839 bgr_11_0.V_TOP.n38 GNDA 0.089272f
C840 bgr_11_0.V_TOP.t26 GNDA 0.129529f
C841 bgr_11_0.V_TOP.n39 GNDA 0.089272f
C842 bgr_11_0.V_TOP.t49 GNDA 0.129529f
C843 bgr_11_0.V_TOP.n40 GNDA 0.089272f
C844 bgr_11_0.V_TOP.t42 GNDA 0.129529f
C845 bgr_11_0.V_TOP.n41 GNDA 0.089272f
C846 bgr_11_0.V_TOP.t33 GNDA 0.129529f
C847 bgr_11_0.V_TOP.n42 GNDA 0.080857f
C848 bgr_11_0.V_TOP.t21 GNDA 0.128562f
C849 VOUT+.n0 GNDA 0.035859f
C850 VOUT+.t13 GNDA 0.052295f
C851 VOUT+.t17 GNDA 0.052295f
C852 VOUT+.n1 GNDA 0.112362f
C853 VOUT+.n2 GNDA 0.275831f
C854 VOUT+.n3 GNDA 0.035859f
C855 VOUT+.n4 GNDA 0.237916f
C856 VOUT+.t18 GNDA 0.052295f
C857 VOUT+.t11 GNDA 0.052295f
C858 VOUT+.n5 GNDA 0.112362f
C859 VOUT+.n6 GNDA 0.284527f
C860 VOUT+.n7 GNDA 0.159855f
C861 VOUT+.t14 GNDA 0.052295f
C862 VOUT+.t0 GNDA 0.052295f
C863 VOUT+.n8 GNDA 0.112362f
C864 VOUT+.n9 GNDA 0.271284f
C865 VOUT+.n10 GNDA 0.127531f
C866 VOUT+.n11 GNDA 0.035859f
C867 VOUT+.n12 GNDA 0.185038f
C868 VOUT+.n13 GNDA 0.035859f
C869 VOUT+.n14 GNDA 0.035859f
C870 VOUT+.n15 GNDA 0.035859f
C871 VOUT+.n16 GNDA 0.035859f
C872 VOUT+.n17 GNDA 0.082365f
C873 VOUT+.n18 GNDA 0.096372f
C874 VOUT+.n19 GNDA 0.074707f
C875 VOUT+.n22 GNDA 0.038101f
C876 VOUT+.n24 GNDA 0.038101f
C877 VOUT+.n27 GNDA 0.05603f
C878 VOUT+.n28 GNDA 0.093384f
C879 VOUT+.n29 GNDA 0.059362f
C880 VOUT+.n30 GNDA 0.05603f
C881 VOUT+.n32 GNDA 0.038101f
C882 VOUT+.n33 GNDA 0.035523f
C883 VOUT+.n34 GNDA 0.038101f
C884 VOUT+.n35 GNDA 0.049307f
C885 VOUT+.n36 GNDA 0.071138f
C886 VOUT+.n37 GNDA 0.069229f
C887 VOUT+.n38 GNDA 0.049307f
C888 VOUT+.n39 GNDA 0.049307f
C889 VOUT+.n40 GNDA 0.069229f
C890 VOUT+.n41 GNDA 0.069229f
C891 VOUT+.n42 GNDA 0.049307f
C892 VOUT+.n43 GNDA 0.078936f
C893 VOUT+.t15 GNDA 0.044824f
C894 VOUT+.t5 GNDA 0.044824f
C895 VOUT+.n44 GNDA 0.091845f
C896 VOUT+.n45 GNDA 0.237078f
C897 VOUT+.t9 GNDA 0.044824f
C898 VOUT+.t16 GNDA 0.044824f
C899 VOUT+.n46 GNDA 0.091845f
C900 VOUT+.n47 GNDA 0.237078f
C901 VOUT+.t10 GNDA 0.044824f
C902 VOUT+.t3 GNDA 0.044824f
C903 VOUT+.n48 GNDA 0.091845f
C904 VOUT+.n49 GNDA 0.234689f
C905 VOUT+.n50 GNDA 0.056999f
C906 VOUT+.t6 GNDA 0.044824f
C907 VOUT+.t4 GNDA 0.044824f
C908 VOUT+.n51 GNDA 0.091845f
C909 VOUT+.n52 GNDA 0.234689f
C910 VOUT+.n53 GNDA 0.032309f
C911 VOUT+.t7 GNDA 0.044824f
C912 VOUT+.t1 GNDA 0.044824f
C913 VOUT+.n54 GNDA 0.091845f
C914 VOUT+.n55 GNDA 0.234689f
C915 VOUT+.n56 GNDA 0.032309f
C916 VOUT+.n57 GNDA 0.056999f
C917 VOUT+.t8 GNDA 0.044824f
C918 VOUT+.t2 GNDA 0.044824f
C919 VOUT+.n58 GNDA 0.091845f
C920 VOUT+.n59 GNDA 0.234689f
C921 VOUT+.n60 GNDA 0.037686f
C922 VOUT+.n61 GNDA 0.022412f
C923 VOUT+.n62 GNDA 0.022412f
C924 VOUT+.n63 GNDA 0.037686f
C925 VOUT+.n64 GNDA 0.069229f
C926 VOUT+.n65 GNDA 0.096906f
C927 VOUT+.n66 GNDA 0.120749f
C928 VOUT+.n67 GNDA 0.169f
C929 VOUT+.n68 GNDA 0.049307f
C930 VOUT+.n69 GNDA 0.080684f
C931 VOUT+.n70 GNDA 0.049307f
C932 VOUT+.n71 GNDA 0.080684f
C933 VOUT+.n72 GNDA 0.049307f
C934 VOUT+.n73 GNDA 0.049307f
C935 VOUT+.n74 GNDA 0.049307f
C936 VOUT+.n75 GNDA 0.080684f
C937 VOUT+.n76 GNDA 0.049307f
C938 VOUT+.n77 GNDA 0.07396f
C939 VOUT+.n78 GNDA 0.394453f
C940 VOUT+.n80 GNDA 0.074707f
C941 VOUT+.n81 GNDA 0.038101f
C942 VOUT+.n83 GNDA 0.038101f
C943 VOUT+.n86 GNDA 0.074707f
C944 VOUT+.n87 GNDA 0.387729f
C945 VOUT+.n88 GNDA 0.494934f
C946 VOUT+.n91 GNDA 0.05603f
C947 VOUT+.n92 GNDA 0.05603f
C948 VOUT+.n93 GNDA 0.05603f
C949 VOUT+.n94 GNDA 0.05603f
C950 VOUT+.n95 GNDA 0.164346f
C951 VOUT+.n96 GNDA 0.05603f
C952 VOUT+.t127 GNDA 0.298828f
C953 VOUT+.t121 GNDA 0.303918f
C954 VOUT+.t64 GNDA 0.298828f
C955 VOUT+.n97 GNDA 0.200354f
C956 VOUT+.n98 GNDA 0.130737f
C957 VOUT+.t69 GNDA 0.303281f
C958 VOUT+.t116 GNDA 0.303281f
C959 VOUT+.t57 GNDA 0.303281f
C960 VOUT+.t109 GNDA 0.303281f
C961 VOUT+.t44 GNDA 0.303281f
C962 VOUT+.t146 GNDA 0.303281f
C963 VOUT+.t33 GNDA 0.303281f
C964 VOUT+.t135 GNDA 0.303281f
C965 VOUT+.t74 GNDA 0.303281f
C966 VOUT+.t25 GNDA 0.303281f
C967 VOUT+.t68 GNDA 0.303281f
C968 VOUT+.t20 GNDA 0.303281f
C969 VOUT+.t55 GNDA 0.298828f
C970 VOUT+.n99 GNDA 0.200992f
C971 VOUT+.t21 GNDA 0.298828f
C972 VOUT+.n100 GNDA 0.257022f
C973 VOUT+.t119 GNDA 0.298828f
C974 VOUT+.n101 GNDA 0.257022f
C975 VOUT+.t72 GNDA 0.298828f
C976 VOUT+.n102 GNDA 0.257022f
C977 VOUT+.t35 GNDA 0.298828f
C978 VOUT+.n103 GNDA 0.257022f
C979 VOUT+.t156 GNDA 0.298828f
C980 VOUT+.n104 GNDA 0.257022f
C981 VOUT+.t98 GNDA 0.298828f
C982 VOUT+.n105 GNDA 0.257022f
C983 VOUT+.t63 GNDA 0.298828f
C984 VOUT+.n106 GNDA 0.257022f
C985 VOUT+.t24 GNDA 0.298828f
C986 VOUT+.n107 GNDA 0.257022f
C987 VOUT+.t123 GNDA 0.298828f
C988 VOUT+.n108 GNDA 0.257022f
C989 VOUT+.t75 GNDA 0.298828f
C990 VOUT+.n109 GNDA 0.257022f
C991 VOUT+.t51 GNDA 0.298828f
C992 VOUT+.n110 GNDA 0.257022f
C993 VOUT+.t53 GNDA 0.298828f
C994 VOUT+.t52 GNDA 0.303918f
C995 VOUT+.t157 GNDA 0.298828f
C996 VOUT+.n111 GNDA 0.200354f
C997 VOUT+.n112 GNDA 0.242798f
C998 VOUT+.t124 GNDA 0.303918f
C999 VOUT+.t95 GNDA 0.298828f
C1000 VOUT+.n113 GNDA 0.200354f
C1001 VOUT+.t97 GNDA 0.298828f
C1002 VOUT+.t94 GNDA 0.303918f
C1003 VOUT+.t42 GNDA 0.298828f
C1004 VOUT+.n114 GNDA 0.200354f
C1005 VOUT+.n115 GNDA 0.242798f
C1006 VOUT+.t79 GNDA 0.303918f
C1007 VOUT+.t60 GNDA 0.298828f
C1008 VOUT+.n116 GNDA 0.200354f
C1009 VOUT+.t62 GNDA 0.298828f
C1010 VOUT+.t61 GNDA 0.303918f
C1011 VOUT+.t159 GNDA 0.298828f
C1012 VOUT+.n117 GNDA 0.200354f
C1013 VOUT+.n118 GNDA 0.242798f
C1014 VOUT+.t128 GNDA 0.303918f
C1015 VOUT+.t106 GNDA 0.298828f
C1016 VOUT+.n119 GNDA 0.200354f
C1017 VOUT+.t108 GNDA 0.298828f
C1018 VOUT+.t107 GNDA 0.303918f
C1019 VOUT+.t49 GNDA 0.298828f
C1020 VOUT+.n120 GNDA 0.200354f
C1021 VOUT+.n121 GNDA 0.242798f
C1022 VOUT+.t22 GNDA 0.303918f
C1023 VOUT+.t147 GNDA 0.298828f
C1024 VOUT+.n122 GNDA 0.200354f
C1025 VOUT+.t148 GNDA 0.298828f
C1026 VOUT+.t149 GNDA 0.303918f
C1027 VOUT+.t89 GNDA 0.298828f
C1028 VOUT+.n123 GNDA 0.200354f
C1029 VOUT+.n124 GNDA 0.242798f
C1030 VOUT+.t132 GNDA 0.303918f
C1031 VOUT+.t113 GNDA 0.298828f
C1032 VOUT+.n125 GNDA 0.200354f
C1033 VOUT+.t115 GNDA 0.298828f
C1034 VOUT+.t114 GNDA 0.303918f
C1035 VOUT+.t56 GNDA 0.298828f
C1036 VOUT+.n126 GNDA 0.200354f
C1037 VOUT+.n127 GNDA 0.242798f
C1038 VOUT+.t26 GNDA 0.303918f
C1039 VOUT+.t153 GNDA 0.298828f
C1040 VOUT+.n128 GNDA 0.200354f
C1041 VOUT+.t155 GNDA 0.298828f
C1042 VOUT+.t154 GNDA 0.303918f
C1043 VOUT+.t101 GNDA 0.298828f
C1044 VOUT+.n129 GNDA 0.200354f
C1045 VOUT+.n130 GNDA 0.242798f
C1046 VOUT+.t66 GNDA 0.303918f
C1047 VOUT+.t38 GNDA 0.298828f
C1048 VOUT+.n131 GNDA 0.200354f
C1049 VOUT+.t40 GNDA 0.298828f
C1050 VOUT+.t39 GNDA 0.303918f
C1051 VOUT+.t142 GNDA 0.298828f
C1052 VOUT+.n132 GNDA 0.200354f
C1053 VOUT+.n133 GNDA 0.242798f
C1054 VOUT+.t34 GNDA 0.303918f
C1055 VOUT+.t76 GNDA 0.298828f
C1056 VOUT+.n134 GNDA 0.195685f
C1057 VOUT+.t19 GNDA 0.303918f
C1058 VOUT+.t59 GNDA 0.298828f
C1059 VOUT+.n135 GNDA 0.195685f
C1060 VOUT+.t54 GNDA 0.303918f
C1061 VOUT+.t100 GNDA 0.298828f
C1062 VOUT+.n136 GNDA 0.195685f
C1063 VOUT+.t140 GNDA 0.303518f
C1064 VOUT+.t120 GNDA 0.303518f
C1065 VOUT+.t158 GNDA 0.303531f
C1066 VOUT+.t43 GNDA 0.303531f
C1067 VOUT+.t83 GNDA 0.303518f
C1068 VOUT+.t65 GNDA 0.303531f
C1069 VOUT+.t110 GNDA 0.303531f
C1070 VOUT+.t151 GNDA 0.298828f
C1071 VOUT+.n137 GNDA 0.204477f
C1072 VOUT+.t112 GNDA 0.298828f
C1073 VOUT+.n138 GNDA 0.260507f
C1074 VOUT+.t130 GNDA 0.298828f
C1075 VOUT+.n139 GNDA 0.26052f
C1076 VOUT+.t84 GNDA 0.298828f
C1077 VOUT+.n140 GNDA 0.260507f
C1078 VOUT+.t48 GNDA 0.298828f
C1079 VOUT+.n141 GNDA 0.260507f
C1080 VOUT+.t160 GNDA 0.298828f
C1081 VOUT+.n142 GNDA 0.26052f
C1082 VOUT+.t29 GNDA 0.298828f
C1083 VOUT+.n143 GNDA 0.26052f
C1084 VOUT+.t141 GNDA 0.298828f
C1085 VOUT+.n144 GNDA 0.191437f
C1086 VOUT+.t105 GNDA 0.298828f
C1087 VOUT+.n145 GNDA 0.191437f
C1088 VOUT+.t126 GNDA 0.298828f
C1089 VOUT+.n146 GNDA 0.191437f
C1090 VOUT+.t78 GNDA 0.298828f
C1091 VOUT+.n147 GNDA 0.130737f
C1092 VOUT+.t73 GNDA 0.298828f
C1093 VOUT+.n148 GNDA 0.130737f
C1094 VOUT+.t118 GNDA 0.298828f
C1095 VOUT+.t70 GNDA 0.303918f
C1096 VOUT+.t32 GNDA 0.298828f
C1097 VOUT+.n149 GNDA 0.200354f
C1098 VOUT+.n150 GNDA 0.186768f
C1099 VOUT+.t37 GNDA 0.303918f
C1100 VOUT+.t31 GNDA 0.298828f
C1101 VOUT+.n151 GNDA 0.200354f
C1102 VOUT+.t67 GNDA 0.298828f
C1103 VOUT+.t28 GNDA 0.303918f
C1104 VOUT+.t145 GNDA 0.298828f
C1105 VOUT+.n152 GNDA 0.200354f
C1106 VOUT+.n153 GNDA 0.242798f
C1107 VOUT+.t152 GNDA 0.303918f
C1108 VOUT+.t143 GNDA 0.298828f
C1109 VOUT+.n154 GNDA 0.200354f
C1110 VOUT+.t27 GNDA 0.298828f
C1111 VOUT+.t139 GNDA 0.303918f
C1112 VOUT+.t104 GNDA 0.298828f
C1113 VOUT+.n155 GNDA 0.200354f
C1114 VOUT+.n156 GNDA 0.242798f
C1115 VOUT+.t111 GNDA 0.303918f
C1116 VOUT+.t102 GNDA 0.298828f
C1117 VOUT+.n157 GNDA 0.200354f
C1118 VOUT+.t137 GNDA 0.298828f
C1119 VOUT+.t92 GNDA 0.303918f
C1120 VOUT+.t58 GNDA 0.298828f
C1121 VOUT+.n158 GNDA 0.200354f
C1122 VOUT+.n159 GNDA 0.242798f
C1123 VOUT+.t144 GNDA 0.303918f
C1124 VOUT+.t138 GNDA 0.298828f
C1125 VOUT+.n160 GNDA 0.200354f
C1126 VOUT+.t23 GNDA 0.298828f
C1127 VOUT+.t131 GNDA 0.303918f
C1128 VOUT+.t91 GNDA 0.298828f
C1129 VOUT+.n161 GNDA 0.200354f
C1130 VOUT+.n162 GNDA 0.242798f
C1131 VOUT+.t103 GNDA 0.303918f
C1132 VOUT+.t90 GNDA 0.298828f
C1133 VOUT+.n163 GNDA 0.200354f
C1134 VOUT+.t129 GNDA 0.298828f
C1135 VOUT+.t85 GNDA 0.303918f
C1136 VOUT+.t50 GNDA 0.298828f
C1137 VOUT+.n164 GNDA 0.200354f
C1138 VOUT+.n165 GNDA 0.242798f
C1139 VOUT+.t125 GNDA 0.303918f
C1140 VOUT+.t93 GNDA 0.298828f
C1141 VOUT+.n166 GNDA 0.200354f
C1142 VOUT+.t99 GNDA 0.298828f
C1143 VOUT+.t96 GNDA 0.303918f
C1144 VOUT+.t41 GNDA 0.298828f
C1145 VOUT+.n167 GNDA 0.200354f
C1146 VOUT+.n168 GNDA 0.242798f
C1147 VOUT+.t161 GNDA 0.303918f
C1148 VOUT+.t133 GNDA 0.298828f
C1149 VOUT+.n169 GNDA 0.200354f
C1150 VOUT+.t136 GNDA 0.298828f
C1151 VOUT+.t134 GNDA 0.303918f
C1152 VOUT+.t77 GNDA 0.298828f
C1153 VOUT+.n170 GNDA 0.200354f
C1154 VOUT+.n171 GNDA 0.242798f
C1155 VOUT+.t122 GNDA 0.303918f
C1156 VOUT+.t86 GNDA 0.298828f
C1157 VOUT+.n172 GNDA 0.200354f
C1158 VOUT+.t88 GNDA 0.298828f
C1159 VOUT+.t87 GNDA 0.303918f
C1160 VOUT+.t36 GNDA 0.298828f
C1161 VOUT+.n173 GNDA 0.200354f
C1162 VOUT+.n174 GNDA 0.242798f
C1163 VOUT+.t71 GNDA 0.303918f
C1164 VOUT+.t45 GNDA 0.298828f
C1165 VOUT+.n175 GNDA 0.200354f
C1166 VOUT+.t47 GNDA 0.298828f
C1167 VOUT+.t46 GNDA 0.303918f
C1168 VOUT+.t150 GNDA 0.298828f
C1169 VOUT+.n176 GNDA 0.200354f
C1170 VOUT+.n177 GNDA 0.242798f
C1171 VOUT+.t81 GNDA 0.303918f
C1172 VOUT+.t30 GNDA 0.298828f
C1173 VOUT+.n178 GNDA 0.200354f
C1174 VOUT+.t82 GNDA 0.298828f
C1175 VOUT+.n179 GNDA 0.242798f
C1176 VOUT+.t80 GNDA 0.298828f
C1177 VOUT+.n180 GNDA 0.127936f
C1178 VOUT+.t117 GNDA 0.298828f
C1179 VOUT+.n181 GNDA 0.33338f
C1180 VOUT+.n182 GNDA 0.274548f
C1181 VOUT+.n183 GNDA 0.05603f
C1182 VOUT+.n184 GNDA 0.05603f
C1183 VOUT+.n186 GNDA 0.504272f
C1184 VOUT+.n187 GNDA 0.056444f
C1185 VOUT+.n188 GNDA 1.06457f
C1186 VOUT+.n189 GNDA 0.038101f
C1187 VOUT+.n191 GNDA 0.035859f
C1188 VOUT+.n192 GNDA 1.05524f
C1189 VOUT+.n194 GNDA 0.038101f
C1190 VOUT+.n195 GNDA 0.074707f
C1191 VOUT+.n196 GNDA 0.257739f
C1192 VOUT+.t12 GNDA 0.085603f
C1193 VOUT+.n197 GNDA 0.42035f
C1194 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t80 GNDA 0.35871f
C1195 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t19 GNDA 0.376298f
C1196 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t97 GNDA 0.35871f
C1197 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t106 GNDA 0.19267f
C1198 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n0 GNDA 0.206205f
C1199 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t91 GNDA 0.35871f
C1200 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t20 GNDA 0.19267f
C1201 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n1 GNDA 0.204542f
C1202 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t13 GNDA 0.35871f
C1203 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t82 GNDA 0.19267f
C1204 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n2 GNDA 0.204542f
C1205 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t102 GNDA 0.35871f
C1206 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t32 GNDA 0.19267f
C1207 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n3 GNDA 0.204542f
C1208 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t124 GNDA 0.35871f
C1209 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t128 GNDA 0.19267f
C1210 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n4 GNDA 0.204542f
C1211 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t4 GNDA 0.35871f
C1212 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t139 GNDA 0.19267f
C1213 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n5 GNDA 0.204542f
C1214 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t60 GNDA 0.35871f
C1215 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t46 GNDA 0.36001f
C1216 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t15 GNDA 0.35871f
C1217 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t65 GNDA 0.36001f
C1218 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t138 GNDA 0.35871f
C1219 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t1 GNDA 0.36001f
C1220 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t68 GNDA 0.35871f
C1221 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t77 GNDA 0.36001f
C1222 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t79 GNDA 0.35871f
C1223 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t108 GNDA 0.36001f
C1224 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t81 GNDA 0.35871f
C1225 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t88 GNDA 0.36001f
C1226 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t28 GNDA 0.35871f
C1227 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t84 GNDA 0.36001f
C1228 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t0 GNDA 0.35871f
C1229 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t78 GNDA 0.36001f
C1230 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t21 GNDA 0.35871f
C1231 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t57 GNDA 0.36001f
C1232 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t89 GNDA 0.35871f
C1233 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t56 GNDA 0.36001f
C1234 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t83 GNDA 0.35871f
C1235 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t40 GNDA 0.36001f
C1236 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t43 GNDA 0.35871f
C1237 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t29 GNDA 0.36001f
C1238 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t110 GNDA 0.35871f
C1239 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t17 GNDA 0.36001f
C1240 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t129 GNDA 0.35871f
C1241 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t71 GNDA 0.36001f
C1242 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t48 GNDA 0.35871f
C1243 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t115 GNDA 0.36001f
C1244 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t38 GNDA 0.35871f
C1245 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t112 GNDA 0.36001f
C1246 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t113 GNDA 0.35871f
C1247 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t14 GNDA 0.36001f
C1248 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t61 GNDA 0.35871f
C1249 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t87 GNDA 0.36001f
C1250 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t126 GNDA 0.35871f
C1251 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t18 GNDA 0.36001f
C1252 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t51 GNDA 0.35871f
C1253 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t58 GNDA 0.36001f
C1254 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t59 GNDA 0.35871f
C1255 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t64 GNDA 0.36001f
C1256 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t116 GNDA 0.35871f
C1257 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t62 GNDA 0.36001f
C1258 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t63 GNDA 0.35871f
C1259 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t76 GNDA 0.36001f
C1260 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t120 GNDA 0.35871f
C1261 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t69 GNDA 0.36001f
C1262 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t142 GNDA 0.35871f
C1263 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t55 GNDA 0.36001f
C1264 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t70 GNDA 0.35871f
C1265 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t107 GNDA 0.36001f
C1266 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t130 GNDA 0.35871f
C1267 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t24 GNDA 0.36001f
C1268 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t140 GNDA 0.35871f
C1269 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t75 GNDA 0.36001f
C1270 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t99 GNDA 0.35871f
C1271 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t135 GNDA 0.36001f
C1272 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t6 GNDA 0.35871f
C1273 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t132 GNDA 0.36001f
C1274 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t133 GNDA 0.35871f
C1275 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t33 GNDA 0.36001f
C1276 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t11 GNDA 0.35871f
C1277 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t22 GNDA 0.36001f
C1278 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t23 GNDA 0.35871f
C1279 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t103 GNDA 0.36001f
C1280 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t42 GNDA 0.35871f
C1281 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t35 GNDA 0.36001f
C1282 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t34 GNDA 0.35871f
C1283 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t12 GNDA 0.36001f
C1284 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t122 GNDA 0.35871f
C1285 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t27 GNDA 0.376298f
C1286 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t136 GNDA 0.35871f
C1287 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t123 GNDA 0.19267f
C1288 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n6 GNDA 0.206205f
C1289 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t67 GNDA 0.35871f
C1290 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t105 GNDA 0.19267f
C1291 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n7 GNDA 0.204542f
C1292 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t36 GNDA 0.35871f
C1293 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t30 GNDA 0.19267f
C1294 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n8 GNDA 0.204542f
C1295 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t49 GNDA 0.35871f
C1296 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t119 GNDA 0.19267f
C1297 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n9 GNDA 0.204542f
C1298 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t47 GNDA 0.35871f
C1299 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t92 GNDA 0.19267f
C1300 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n10 GNDA 0.204542f
C1301 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t74 GNDA 0.35871f
C1302 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t8 GNDA 0.19267f
C1303 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n11 GNDA 0.204542f
C1304 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t86 GNDA 0.35871f
C1305 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t73 GNDA 0.19267f
C1306 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n12 GNDA 0.204542f
C1307 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t53 GNDA 0.35871f
C1308 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t66 GNDA 0.19267f
C1309 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n13 GNDA 0.204542f
C1310 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t25 GNDA 0.35871f
C1311 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t39 GNDA 0.19267f
C1312 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n14 GNDA 0.204542f
C1313 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t50 GNDA 0.35871f
C1314 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t37 GNDA 0.19267f
C1315 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n15 GNDA 0.204542f
C1316 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t137 GNDA 0.35871f
C1317 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t41 GNDA 0.19267f
C1318 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n16 GNDA 0.204542f
C1319 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t44 GNDA 0.35871f
C1320 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t93 GNDA 0.36001f
C1321 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t125 GNDA 0.35871f
C1322 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t96 GNDA 0.36001f
C1323 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t101 GNDA 0.173419f
C1324 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n17 GNDA 0.223685f
C1325 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t45 GNDA 0.191478f
C1326 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n18 GNDA 0.242936f
C1327 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t111 GNDA 0.191478f
C1328 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n19 GNDA 0.260887f
C1329 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t72 GNDA 0.191478f
C1330 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n20 GNDA 0.260887f
C1331 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t52 GNDA 0.191478f
C1332 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n21 GNDA 0.260887f
C1333 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t98 GNDA 0.191478f
C1334 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n22 GNDA 0.260887f
C1335 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t131 GNDA 0.191478f
C1336 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n23 GNDA 0.260887f
C1337 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t143 GNDA 0.191478f
C1338 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n24 GNDA 0.260887f
C1339 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t16 GNDA 0.191478f
C1340 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n25 GNDA 0.260887f
C1341 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t90 GNDA 0.191478f
C1342 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n26 GNDA 0.260887f
C1343 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t127 GNDA 0.191478f
C1344 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n27 GNDA 0.260887f
C1345 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t134 GNDA 0.191478f
C1346 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n28 GNDA 0.260887f
C1347 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t94 GNDA 0.191478f
C1348 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n29 GNDA 0.260887f
C1349 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t9 GNDA 0.191478f
C1350 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n30 GNDA 0.260887f
C1351 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t7 GNDA 0.191478f
C1352 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n31 GNDA 0.260887f
C1353 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t141 GNDA 0.191478f
C1354 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n32 GNDA 0.260887f
C1355 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t95 GNDA 0.191478f
C1356 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n33 GNDA 0.260887f
C1357 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t121 GNDA 0.191478f
C1358 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n34 GNDA 0.260887f
C1359 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t117 GNDA 0.191478f
C1360 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n35 GNDA 0.260887f
C1361 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t104 GNDA 0.191478f
C1362 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n36 GNDA 0.240444f
C1363 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t31 GNDA 0.36001f
C1364 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t10 GNDA 0.36001f
C1365 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t118 GNDA 0.35871f
C1366 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t114 GNDA 0.377961f
C1367 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t100 GNDA 0.19267f
C1368 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n37 GNDA 0.222493f
C1369 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t2 GNDA 0.35871f
C1370 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t85 GNDA 0.377961f
C1371 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t109 GNDA 0.19267f
C1372 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n38 GNDA 0.204542f
C1373 two_stage_opamp_dummy_magic_29_0.cap_res_Y.n39 GNDA 0.204542f
C1374 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t5 GNDA 0.19267f
C1375 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t54 GNDA 0.377961f
C1376 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t26 GNDA 0.454191f
C1377 two_stage_opamp_dummy_magic_29_0.cap_res_Y.t3 GNDA 0.317638f
C1378 two_stage_opamp_dummy_magic_29_0.cap_res_X.t51 GNDA 0.358056f
C1379 two_stage_opamp_dummy_magic_29_0.cap_res_X.t26 GNDA 0.359353f
C1380 two_stage_opamp_dummy_magic_29_0.cap_res_X.t93 GNDA 0.358056f
C1381 two_stage_opamp_dummy_magic_29_0.cap_res_X.t67 GNDA 0.359353f
C1382 two_stage_opamp_dummy_magic_29_0.cap_res_X.t120 GNDA 0.358056f
C1383 two_stage_opamp_dummy_magic_29_0.cap_res_X.t142 GNDA 0.359353f
C1384 two_stage_opamp_dummy_magic_29_0.cap_res_X.t130 GNDA 0.358056f
C1385 two_stage_opamp_dummy_magic_29_0.cap_res_X.t103 GNDA 0.359353f
C1386 two_stage_opamp_dummy_magic_29_0.cap_res_X.t18 GNDA 0.358056f
C1387 two_stage_opamp_dummy_magic_29_0.cap_res_X.t45 GNDA 0.359353f
C1388 two_stage_opamp_dummy_magic_29_0.cap_res_X.t29 GNDA 0.358056f
C1389 two_stage_opamp_dummy_magic_29_0.cap_res_X.t2 GNDA 0.359353f
C1390 two_stage_opamp_dummy_magic_29_0.cap_res_X.t60 GNDA 0.358056f
C1391 two_stage_opamp_dummy_magic_29_0.cap_res_X.t85 GNDA 0.359353f
C1392 two_stage_opamp_dummy_magic_29_0.cap_res_X.t135 GNDA 0.358056f
C1393 two_stage_opamp_dummy_magic_29_0.cap_res_X.t108 GNDA 0.359353f
C1394 two_stage_opamp_dummy_magic_29_0.cap_res_X.t23 GNDA 0.358056f
C1395 two_stage_opamp_dummy_magic_29_0.cap_res_X.t50 GNDA 0.359353f
C1396 two_stage_opamp_dummy_magic_29_0.cap_res_X.t35 GNDA 0.358056f
C1397 two_stage_opamp_dummy_magic_29_0.cap_res_X.t9 GNDA 0.359353f
C1398 two_stage_opamp_dummy_magic_29_0.cap_res_X.t64 GNDA 0.358056f
C1399 two_stage_opamp_dummy_magic_29_0.cap_res_X.t92 GNDA 0.359353f
C1400 two_stage_opamp_dummy_magic_29_0.cap_res_X.t131 GNDA 0.358056f
C1401 two_stage_opamp_dummy_magic_29_0.cap_res_X.t41 GNDA 0.359353f
C1402 two_stage_opamp_dummy_magic_29_0.cap_res_X.t21 GNDA 0.358056f
C1403 two_stage_opamp_dummy_magic_29_0.cap_res_X.t111 GNDA 0.359353f
C1404 two_stage_opamp_dummy_magic_29_0.cap_res_X.t97 GNDA 0.358056f
C1405 two_stage_opamp_dummy_magic_29_0.cap_res_X.t4 GNDA 0.359353f
C1406 two_stage_opamp_dummy_magic_29_0.cap_res_X.t129 GNDA 0.358056f
C1407 two_stage_opamp_dummy_magic_29_0.cap_res_X.t79 GNDA 0.359353f
C1408 two_stage_opamp_dummy_magic_29_0.cap_res_X.t137 GNDA 0.358056f
C1409 two_stage_opamp_dummy_magic_29_0.cap_res_X.t49 GNDA 0.359353f
C1410 two_stage_opamp_dummy_magic_29_0.cap_res_X.t28 GNDA 0.358056f
C1411 two_stage_opamp_dummy_magic_29_0.cap_res_X.t116 GNDA 0.359353f
C1412 two_stage_opamp_dummy_magic_29_0.cap_res_X.t38 GNDA 0.358056f
C1413 two_stage_opamp_dummy_magic_29_0.cap_res_X.t90 GNDA 0.359353f
C1414 two_stage_opamp_dummy_magic_29_0.cap_res_X.t69 GNDA 0.358056f
C1415 two_stage_opamp_dummy_magic_29_0.cap_res_X.t13 GNDA 0.359353f
C1416 two_stage_opamp_dummy_magic_29_0.cap_res_X.t140 GNDA 0.358056f
C1417 two_stage_opamp_dummy_magic_29_0.cap_res_X.t54 GNDA 0.359353f
C1418 two_stage_opamp_dummy_magic_29_0.cap_res_X.t34 GNDA 0.358056f
C1419 two_stage_opamp_dummy_magic_29_0.cap_res_X.t123 GNDA 0.359353f
C1420 two_stage_opamp_dummy_magic_29_0.cap_res_X.t40 GNDA 0.358056f
C1421 two_stage_opamp_dummy_magic_29_0.cap_res_X.t94 GNDA 0.359353f
C1422 two_stage_opamp_dummy_magic_29_0.cap_res_X.t74 GNDA 0.358056f
C1423 two_stage_opamp_dummy_magic_29_0.cap_res_X.t19 GNDA 0.359353f
C1424 two_stage_opamp_dummy_magic_29_0.cap_res_X.t82 GNDA 0.358056f
C1425 two_stage_opamp_dummy_magic_29_0.cap_res_X.t133 GNDA 0.359353f
C1426 two_stage_opamp_dummy_magic_29_0.cap_res_X.t112 GNDA 0.358056f
C1427 two_stage_opamp_dummy_magic_29_0.cap_res_X.t61 GNDA 0.359353f
C1428 two_stage_opamp_dummy_magic_29_0.cap_res_X.t121 GNDA 0.358056f
C1429 two_stage_opamp_dummy_magic_29_0.cap_res_X.t31 GNDA 0.359353f
C1430 two_stage_opamp_dummy_magic_29_0.cap_res_X.t11 GNDA 0.358056f
C1431 two_stage_opamp_dummy_magic_29_0.cap_res_X.t100 GNDA 0.359353f
C1432 two_stage_opamp_dummy_magic_29_0.cap_res_X.t86 GNDA 0.358056f
C1433 two_stage_opamp_dummy_magic_29_0.cap_res_X.t138 GNDA 0.359353f
C1434 two_stage_opamp_dummy_magic_29_0.cap_res_X.t117 GNDA 0.358056f
C1435 two_stage_opamp_dummy_magic_29_0.cap_res_X.t68 GNDA 0.359353f
C1436 two_stage_opamp_dummy_magic_29_0.cap_res_X.t126 GNDA 0.358056f
C1437 two_stage_opamp_dummy_magic_29_0.cap_res_X.t39 GNDA 0.359353f
C1438 two_stage_opamp_dummy_magic_29_0.cap_res_X.t15 GNDA 0.358056f
C1439 two_stage_opamp_dummy_magic_29_0.cap_res_X.t104 GNDA 0.359353f
C1440 two_stage_opamp_dummy_magic_29_0.cap_res_X.t24 GNDA 0.358056f
C1441 two_stage_opamp_dummy_magic_29_0.cap_res_X.t78 GNDA 0.359353f
C1442 two_stage_opamp_dummy_magic_29_0.cap_res_X.t57 GNDA 0.358056f
C1443 two_stage_opamp_dummy_magic_29_0.cap_res_X.t3 GNDA 0.359353f
C1444 two_stage_opamp_dummy_magic_29_0.cap_res_X.t132 GNDA 0.358056f
C1445 two_stage_opamp_dummy_magic_29_0.cap_res_X.t42 GNDA 0.359353f
C1446 two_stage_opamp_dummy_magic_29_0.cap_res_X.t20 GNDA 0.358056f
C1447 two_stage_opamp_dummy_magic_29_0.cap_res_X.t109 GNDA 0.359353f
C1448 two_stage_opamp_dummy_magic_29_0.cap_res_X.t30 GNDA 0.358056f
C1449 two_stage_opamp_dummy_magic_29_0.cap_res_X.t83 GNDA 0.359353f
C1450 two_stage_opamp_dummy_magic_29_0.cap_res_X.t53 GNDA 0.358056f
C1451 two_stage_opamp_dummy_magic_29_0.cap_res_X.t70 GNDA 0.375611f
C1452 two_stage_opamp_dummy_magic_29_0.cap_res_X.t7 GNDA 0.358056f
C1453 two_stage_opamp_dummy_magic_29_0.cap_res_X.t14 GNDA 0.192319f
C1454 two_stage_opamp_dummy_magic_29_0.cap_res_X.n0 GNDA 0.205829f
C1455 two_stage_opamp_dummy_magic_29_0.cap_res_X.t89 GNDA 0.358056f
C1456 two_stage_opamp_dummy_magic_29_0.cap_res_X.t95 GNDA 0.192319f
C1457 two_stage_opamp_dummy_magic_29_0.cap_res_X.n1 GNDA 0.204169f
C1458 two_stage_opamp_dummy_magic_29_0.cap_res_X.t139 GNDA 0.358056f
C1459 two_stage_opamp_dummy_magic_29_0.cap_res_X.t59 GNDA 0.192319f
C1460 two_stage_opamp_dummy_magic_29_0.cap_res_X.n2 GNDA 0.204169f
C1461 two_stage_opamp_dummy_magic_29_0.cap_res_X.t96 GNDA 0.358056f
C1462 two_stage_opamp_dummy_magic_29_0.cap_res_X.t6 GNDA 0.192319f
C1463 two_stage_opamp_dummy_magic_29_0.cap_res_X.n3 GNDA 0.204169f
C1464 two_stage_opamp_dummy_magic_29_0.cap_res_X.t1 GNDA 0.358056f
C1465 two_stage_opamp_dummy_magic_29_0.cap_res_X.t113 GNDA 0.192319f
C1466 two_stage_opamp_dummy_magic_29_0.cap_res_X.n4 GNDA 0.204169f
C1467 two_stage_opamp_dummy_magic_29_0.cap_res_X.t56 GNDA 0.358056f
C1468 two_stage_opamp_dummy_magic_29_0.cap_res_X.t80 GNDA 0.192319f
C1469 two_stage_opamp_dummy_magic_29_0.cap_res_X.n5 GNDA 0.204169f
C1470 two_stage_opamp_dummy_magic_29_0.cap_res_X.t105 GNDA 0.358056f
C1471 two_stage_opamp_dummy_magic_29_0.cap_res_X.t46 GNDA 0.192319f
C1472 two_stage_opamp_dummy_magic_29_0.cap_res_X.n6 GNDA 0.204169f
C1473 two_stage_opamp_dummy_magic_29_0.cap_res_X.t65 GNDA 0.358056f
C1474 two_stage_opamp_dummy_magic_29_0.cap_res_X.t134 GNDA 0.192319f
C1475 two_stage_opamp_dummy_magic_29_0.cap_res_X.n7 GNDA 0.204169f
C1476 two_stage_opamp_dummy_magic_29_0.cap_res_X.t114 GNDA 0.358056f
C1477 two_stage_opamp_dummy_magic_29_0.cap_res_X.t99 GNDA 0.192319f
C1478 two_stage_opamp_dummy_magic_29_0.cap_res_X.n8 GNDA 0.204169f
C1479 two_stage_opamp_dummy_magic_29_0.cap_res_X.t27 GNDA 0.358056f
C1480 two_stage_opamp_dummy_magic_29_0.cap_res_X.t62 GNDA 0.192319f
C1481 two_stage_opamp_dummy_magic_29_0.cap_res_X.n9 GNDA 0.204169f
C1482 two_stage_opamp_dummy_magic_29_0.cap_res_X.t125 GNDA 0.358056f
C1483 two_stage_opamp_dummy_magic_29_0.cap_res_X.t10 GNDA 0.192319f
C1484 two_stage_opamp_dummy_magic_29_0.cap_res_X.n10 GNDA 0.204169f
C1485 two_stage_opamp_dummy_magic_29_0.cap_res_X.t48 GNDA 0.358056f
C1486 two_stage_opamp_dummy_magic_29_0.cap_res_X.t88 GNDA 0.359353f
C1487 two_stage_opamp_dummy_magic_29_0.cap_res_X.t37 GNDA 0.173103f
C1488 two_stage_opamp_dummy_magic_29_0.cap_res_X.n11 GNDA 0.223277f
C1489 two_stage_opamp_dummy_magic_29_0.cap_res_X.t115 GNDA 0.191129f
C1490 two_stage_opamp_dummy_magic_29_0.cap_res_X.n12 GNDA 0.242493f
C1491 two_stage_opamp_dummy_magic_29_0.cap_res_X.t77 GNDA 0.191129f
C1492 two_stage_opamp_dummy_magic_29_0.cap_res_X.n13 GNDA 0.260411f
C1493 two_stage_opamp_dummy_magic_29_0.cap_res_X.t110 GNDA 0.191129f
C1494 two_stage_opamp_dummy_magic_29_0.cap_res_X.n14 GNDA 0.260411f
C1495 two_stage_opamp_dummy_magic_29_0.cap_res_X.t72 GNDA 0.191129f
C1496 two_stage_opamp_dummy_magic_29_0.cap_res_X.n15 GNDA 0.260411f
C1497 two_stage_opamp_dummy_magic_29_0.cap_res_X.t32 GNDA 0.191129f
C1498 two_stage_opamp_dummy_magic_29_0.cap_res_X.n16 GNDA 0.260411f
C1499 two_stage_opamp_dummy_magic_29_0.cap_res_X.t66 GNDA 0.191129f
C1500 two_stage_opamp_dummy_magic_29_0.cap_res_X.n17 GNDA 0.260411f
C1501 two_stage_opamp_dummy_magic_29_0.cap_res_X.t25 GNDA 0.191129f
C1502 two_stage_opamp_dummy_magic_29_0.cap_res_X.n18 GNDA 0.260411f
C1503 two_stage_opamp_dummy_magic_29_0.cap_res_X.t128 GNDA 0.191129f
C1504 two_stage_opamp_dummy_magic_29_0.cap_res_X.n19 GNDA 0.260411f
C1505 two_stage_opamp_dummy_magic_29_0.cap_res_X.t91 GNDA 0.191129f
C1506 two_stage_opamp_dummy_magic_29_0.cap_res_X.n20 GNDA 0.260411f
C1507 two_stage_opamp_dummy_magic_29_0.cap_res_X.t122 GNDA 0.191129f
C1508 two_stage_opamp_dummy_magic_29_0.cap_res_X.n21 GNDA 0.260411f
C1509 two_stage_opamp_dummy_magic_29_0.cap_res_X.t84 GNDA 0.191129f
C1510 two_stage_opamp_dummy_magic_29_0.cap_res_X.n22 GNDA 0.260411f
C1511 two_stage_opamp_dummy_magic_29_0.cap_res_X.t43 GNDA 0.191129f
C1512 two_stage_opamp_dummy_magic_29_0.cap_res_X.n23 GNDA 0.260411f
C1513 two_stage_opamp_dummy_magic_29_0.cap_res_X.t76 GNDA 0.191129f
C1514 two_stage_opamp_dummy_magic_29_0.cap_res_X.n24 GNDA 0.260411f
C1515 two_stage_opamp_dummy_magic_29_0.cap_res_X.t52 GNDA 0.191129f
C1516 two_stage_opamp_dummy_magic_29_0.cap_res_X.n25 GNDA 0.260411f
C1517 two_stage_opamp_dummy_magic_29_0.cap_res_X.t8 GNDA 0.191129f
C1518 two_stage_opamp_dummy_magic_29_0.cap_res_X.n26 GNDA 0.260411f
C1519 two_stage_opamp_dummy_magic_29_0.cap_res_X.t47 GNDA 0.191129f
C1520 two_stage_opamp_dummy_magic_29_0.cap_res_X.n27 GNDA 0.260411f
C1521 two_stage_opamp_dummy_magic_29_0.cap_res_X.t0 GNDA 0.191129f
C1522 two_stage_opamp_dummy_magic_29_0.cap_res_X.n28 GNDA 0.260411f
C1523 two_stage_opamp_dummy_magic_29_0.cap_res_X.t102 GNDA 0.191129f
C1524 two_stage_opamp_dummy_magic_29_0.cap_res_X.n29 GNDA 0.260411f
C1525 two_stage_opamp_dummy_magic_29_0.cap_res_X.t63 GNDA 0.191129f
C1526 two_stage_opamp_dummy_magic_29_0.cap_res_X.n30 GNDA 0.240005f
C1527 two_stage_opamp_dummy_magic_29_0.cap_res_X.t101 GNDA 0.359353f
C1528 two_stage_opamp_dummy_magic_29_0.cap_res_X.t81 GNDA 0.359353f
C1529 two_stage_opamp_dummy_magic_29_0.cap_res_X.t58 GNDA 0.358056f
C1530 two_stage_opamp_dummy_magic_29_0.cap_res_X.t16 GNDA 0.377272f
C1531 two_stage_opamp_dummy_magic_29_0.cap_res_X.t118 GNDA 0.192319f
C1532 two_stage_opamp_dummy_magic_29_0.cap_res_X.n31 GNDA 0.222087f
C1533 two_stage_opamp_dummy_magic_29_0.cap_res_X.t98 GNDA 0.358056f
C1534 two_stage_opamp_dummy_magic_29_0.cap_res_X.t55 GNDA 0.377272f
C1535 two_stage_opamp_dummy_magic_29_0.cap_res_X.t12 GNDA 0.192319f
C1536 two_stage_opamp_dummy_magic_29_0.cap_res_X.n32 GNDA 0.204169f
C1537 two_stage_opamp_dummy_magic_29_0.cap_res_X.t17 GNDA 0.358056f
C1538 two_stage_opamp_dummy_magic_29_0.cap_res_X.t119 GNDA 0.375611f
C1539 two_stage_opamp_dummy_magic_29_0.cap_res_X.t44 GNDA 0.358056f
C1540 two_stage_opamp_dummy_magic_29_0.cap_res_X.t141 GNDA 0.192319f
C1541 two_stage_opamp_dummy_magic_29_0.cap_res_X.n33 GNDA 0.205829f
C1542 two_stage_opamp_dummy_magic_29_0.cap_res_X.t22 GNDA 0.358056f
C1543 two_stage_opamp_dummy_magic_29_0.cap_res_X.t124 GNDA 0.192319f
C1544 two_stage_opamp_dummy_magic_29_0.cap_res_X.n34 GNDA 0.204169f
C1545 two_stage_opamp_dummy_magic_29_0.cap_res_X.t127 GNDA 0.358056f
C1546 two_stage_opamp_dummy_magic_29_0.cap_res_X.t87 GNDA 0.192319f
C1547 two_stage_opamp_dummy_magic_29_0.cap_res_X.n35 GNDA 0.204169f
C1548 two_stage_opamp_dummy_magic_29_0.cap_res_X.t5 GNDA 0.358056f
C1549 two_stage_opamp_dummy_magic_29_0.cap_res_X.t106 GNDA 0.192319f
C1550 two_stage_opamp_dummy_magic_29_0.cap_res_X.n36 GNDA 0.204169f
C1551 two_stage_opamp_dummy_magic_29_0.cap_res_X.t107 GNDA 0.358056f
C1552 two_stage_opamp_dummy_magic_29_0.cap_res_X.t71 GNDA 0.192319f
C1553 two_stage_opamp_dummy_magic_29_0.cap_res_X.n37 GNDA 0.204169f
C1554 two_stage_opamp_dummy_magic_29_0.cap_res_X.t73 GNDA 0.358056f
C1555 two_stage_opamp_dummy_magic_29_0.cap_res_X.t33 GNDA 0.192319f
C1556 two_stage_opamp_dummy_magic_29_0.cap_res_X.n38 GNDA 0.204169f
C1557 two_stage_opamp_dummy_magic_29_0.cap_res_X.n39 GNDA 0.204169f
C1558 two_stage_opamp_dummy_magic_29_0.cap_res_X.t136 GNDA 0.192319f
C1559 two_stage_opamp_dummy_magic_29_0.cap_res_X.t36 GNDA 0.377272f
C1560 two_stage_opamp_dummy_magic_29_0.cap_res_X.t75 GNDA 0.453363f
C1561 two_stage_opamp_dummy_magic_29_0.cap_res_X.t143 GNDA 0.317057f
C1562 VOUT-.n1 GNDA 0.074623f
C1563 VOUT-.n4 GNDA 0.055967f
C1564 VOUT-.n5 GNDA 0.093278f
C1565 VOUT-.n6 GNDA 0.055967f
C1566 VOUT-.n7 GNDA 0.055967f
C1567 VOUT-.n9 GNDA 0.038057f
C1568 VOUT-.n11 GNDA 0.038057f
C1569 VOUT-.n13 GNDA 0.074623f
C1570 VOUT-.n14 GNDA 0.038057f
C1571 VOUT-.n16 GNDA 0.038057f
C1572 VOUT-.n18 GNDA 0.049251f
C1573 VOUT-.n19 GNDA 0.071057f
C1574 VOUT-.n20 GNDA 0.06915f
C1575 VOUT-.n21 GNDA 0.049251f
C1576 VOUT-.n22 GNDA 0.049251f
C1577 VOUT-.n23 GNDA 0.06915f
C1578 VOUT-.n24 GNDA 0.06915f
C1579 VOUT-.n25 GNDA 0.049251f
C1580 VOUT-.n26 GNDA 0.078847f
C1581 VOUT-.t6 GNDA 0.044774f
C1582 VOUT-.t11 GNDA 0.044774f
C1583 VOUT-.n27 GNDA 0.091741f
C1584 VOUT-.n28 GNDA 0.236811f
C1585 VOUT-.t15 GNDA 0.044774f
C1586 VOUT-.t9 GNDA 0.044774f
C1587 VOUT-.n29 GNDA 0.091741f
C1588 VOUT-.n30 GNDA 0.234424f
C1589 VOUT-.n31 GNDA 0.056934f
C1590 VOUT-.t16 GNDA 0.044774f
C1591 VOUT-.t10 GNDA 0.044774f
C1592 VOUT-.n32 GNDA 0.091741f
C1593 VOUT-.n33 GNDA 0.234424f
C1594 VOUT-.n34 GNDA 0.032272f
C1595 VOUT-.t14 GNDA 0.044774f
C1596 VOUT-.t8 GNDA 0.044774f
C1597 VOUT-.n35 GNDA 0.091741f
C1598 VOUT-.n36 GNDA 0.234424f
C1599 VOUT-.n37 GNDA 0.032272f
C1600 VOUT-.t12 GNDA 0.044774f
C1601 VOUT-.t5 GNDA 0.044774f
C1602 VOUT-.n38 GNDA 0.091741f
C1603 VOUT-.n39 GNDA 0.236811f
C1604 VOUT-.n40 GNDA 0.056934f
C1605 VOUT-.t13 GNDA 0.044774f
C1606 VOUT-.t7 GNDA 0.044774f
C1607 VOUT-.n41 GNDA 0.091741f
C1608 VOUT-.n42 GNDA 0.234424f
C1609 VOUT-.n43 GNDA 0.037643f
C1610 VOUT-.n44 GNDA 0.022387f
C1611 VOUT-.n45 GNDA 0.022387f
C1612 VOUT-.n46 GNDA 0.037643f
C1613 VOUT-.n47 GNDA 0.06915f
C1614 VOUT-.n48 GNDA 0.096796f
C1615 VOUT-.n49 GNDA 0.120613f
C1616 VOUT-.n50 GNDA 0.168809f
C1617 VOUT-.n51 GNDA 0.049251f
C1618 VOUT-.n52 GNDA 0.080592f
C1619 VOUT-.n53 GNDA 0.049251f
C1620 VOUT-.n54 GNDA 0.080592f
C1621 VOUT-.n55 GNDA 0.049251f
C1622 VOUT-.n56 GNDA 0.049251f
C1623 VOUT-.n57 GNDA 0.049251f
C1624 VOUT-.n58 GNDA 0.080592f
C1625 VOUT-.n59 GNDA 0.049251f
C1626 VOUT-.n60 GNDA 0.073876f
C1627 VOUT-.n61 GNDA 0.394007f
C1628 VOUT-.n62 GNDA 0.387291f
C1629 VOUT-.n64 GNDA 0.074623f
C1630 VOUT-.n65 GNDA 0.035819f
C1631 VOUT-.n66 GNDA 0.494375f
C1632 VOUT-.n69 GNDA 0.055967f
C1633 VOUT-.n70 GNDA 0.055967f
C1634 VOUT-.t113 GNDA 0.303574f
C1635 VOUT-.t73 GNDA 0.29849f
C1636 VOUT-.n71 GNDA 0.200128f
C1637 VOUT-.t124 GNDA 0.29849f
C1638 VOUT-.n72 GNDA 0.13059f
C1639 VOUT-.t131 GNDA 0.303574f
C1640 VOUT-.t78 GNDA 0.29849f
C1641 VOUT-.n73 GNDA 0.200128f
C1642 VOUT-.t46 GNDA 0.29849f
C1643 VOUT-.t36 GNDA 0.302938f
C1644 VOUT-.t134 GNDA 0.302938f
C1645 VOUT-.t47 GNDA 0.302938f
C1646 VOUT-.t96 GNDA 0.302938f
C1647 VOUT-.t56 GNDA 0.302938f
C1648 VOUT-.t105 GNDA 0.302938f
C1649 VOUT-.t160 GNDA 0.302938f
C1650 VOUT-.t65 GNDA 0.302938f
C1651 VOUT-.t22 GNDA 0.302938f
C1652 VOUT-.t72 GNDA 0.302938f
C1653 VOUT-.t154 GNDA 0.302938f
C1654 VOUT-.t108 GNDA 0.302938f
C1655 VOUT-.t91 GNDA 0.29849f
C1656 VOUT-.n74 GNDA 0.200765f
C1657 VOUT-.t147 GNDA 0.29849f
C1658 VOUT-.n75 GNDA 0.256732f
C1659 VOUT-.t66 GNDA 0.29849f
C1660 VOUT-.n76 GNDA 0.256732f
C1661 VOUT-.t102 GNDA 0.29849f
C1662 VOUT-.n77 GNDA 0.256732f
C1663 VOUT-.t155 GNDA 0.29849f
C1664 VOUT-.n78 GNDA 0.256732f
C1665 VOUT-.t48 GNDA 0.29849f
C1666 VOUT-.n79 GNDA 0.256732f
C1667 VOUT-.t81 GNDA 0.29849f
C1668 VOUT-.n80 GNDA 0.256732f
C1669 VOUT-.t115 GNDA 0.29849f
C1670 VOUT-.n81 GNDA 0.256732f
C1671 VOUT-.t27 GNDA 0.29849f
C1672 VOUT-.n82 GNDA 0.256732f
C1673 VOUT-.t62 GNDA 0.29849f
C1674 VOUT-.n83 GNDA 0.256732f
C1675 VOUT-.t99 GNDA 0.29849f
C1676 VOUT-.n84 GNDA 0.256732f
C1677 VOUT-.t151 GNDA 0.29849f
C1678 VOUT-.n85 GNDA 0.256732f
C1679 VOUT-.n86 GNDA 0.242523f
C1680 VOUT-.t29 GNDA 0.303574f
C1681 VOUT-.t119 GNDA 0.29849f
C1682 VOUT-.n87 GNDA 0.200128f
C1683 VOUT-.t84 GNDA 0.29849f
C1684 VOUT-.t141 GNDA 0.303574f
C1685 VOUT-.t52 GNDA 0.29849f
C1686 VOUT-.n88 GNDA 0.200128f
C1687 VOUT-.n89 GNDA 0.242523f
C1688 VOUT-.t137 GNDA 0.303574f
C1689 VOUT-.t83 GNDA 0.29849f
C1690 VOUT-.n90 GNDA 0.200128f
C1691 VOUT-.t51 GNDA 0.29849f
C1692 VOUT-.t104 GNDA 0.303574f
C1693 VOUT-.t158 GNDA 0.29849f
C1694 VOUT-.n91 GNDA 0.200128f
C1695 VOUT-.n92 GNDA 0.242523f
C1696 VOUT-.t35 GNDA 0.303574f
C1697 VOUT-.t122 GNDA 0.29849f
C1698 VOUT-.n93 GNDA 0.200128f
C1699 VOUT-.t89 GNDA 0.29849f
C1700 VOUT-.t146 GNDA 0.303574f
C1701 VOUT-.t57 GNDA 0.29849f
C1702 VOUT-.n94 GNDA 0.200128f
C1703 VOUT-.n95 GNDA 0.242523f
C1704 VOUT-.t75 GNDA 0.303574f
C1705 VOUT-.t23 GNDA 0.29849f
C1706 VOUT-.n96 GNDA 0.200128f
C1707 VOUT-.t129 GNDA 0.29849f
C1708 VOUT-.t44 GNDA 0.303574f
C1709 VOUT-.t93 GNDA 0.29849f
C1710 VOUT-.n97 GNDA 0.200128f
C1711 VOUT-.n98 GNDA 0.242523f
C1712 VOUT-.t40 GNDA 0.303574f
C1713 VOUT-.t130 GNDA 0.29849f
C1714 VOUT-.n99 GNDA 0.200128f
C1715 VOUT-.t95 GNDA 0.29849f
C1716 VOUT-.t150 GNDA 0.303574f
C1717 VOUT-.t61 GNDA 0.29849f
C1718 VOUT-.n100 GNDA 0.200128f
C1719 VOUT-.n101 GNDA 0.242523f
C1720 VOUT-.t79 GNDA 0.303574f
C1721 VOUT-.t28 GNDA 0.29849f
C1722 VOUT-.n102 GNDA 0.200128f
C1723 VOUT-.t136 GNDA 0.29849f
C1724 VOUT-.t49 GNDA 0.303574f
C1725 VOUT-.t100 GNDA 0.29849f
C1726 VOUT-.n103 GNDA 0.200128f
C1727 VOUT-.n104 GNDA 0.242523f
C1728 VOUT-.t121 GNDA 0.303574f
C1729 VOUT-.t67 GNDA 0.29849f
C1730 VOUT-.n105 GNDA 0.200128f
C1731 VOUT-.t33 GNDA 0.29849f
C1732 VOUT-.t87 GNDA 0.303574f
C1733 VOUT-.t142 GNDA 0.29849f
C1734 VOUT-.n106 GNDA 0.200128f
C1735 VOUT-.n107 GNDA 0.242523f
C1736 VOUT-.t110 GNDA 0.303574f
C1737 VOUT-.t135 GNDA 0.29849f
C1738 VOUT-.n108 GNDA 0.200128f
C1739 VOUT-.t98 GNDA 0.29849f
C1740 VOUT-.t103 GNDA 0.303574f
C1741 VOUT-.t145 GNDA 0.29849f
C1742 VOUT-.n109 GNDA 0.195464f
C1743 VOUT-.t63 GNDA 0.303574f
C1744 VOUT-.t106 GNDA 0.29849f
C1745 VOUT-.n110 GNDA 0.195464f
C1746 VOUT-.t86 GNDA 0.303574f
C1747 VOUT-.t125 GNDA 0.29849f
C1748 VOUT-.n111 GNDA 0.195464f
C1749 VOUT-.t88 GNDA 0.302938f
C1750 VOUT-.t54 GNDA 0.302938f
C1751 VOUT-.t156 GNDA 0.302943f
C1752 VOUT-.t34 GNDA 0.303188f
C1753 VOUT-.t139 GNDA 0.302938f
C1754 VOUT-.t117 GNDA 0.302943f
C1755 VOUT-.t144 GNDA 0.303188f
C1756 VOUT-.t42 GNDA 0.29849f
C1757 VOUT-.n112 GNDA 0.204246f
C1758 VOUT-.t20 GNDA 0.29849f
C1759 VOUT-.n113 GNDA 0.256727f
C1760 VOUT-.t37 GNDA 0.29849f
C1761 VOUT-.n114 GNDA 0.256732f
C1762 VOUT-.t74 GNDA 0.29849f
C1763 VOUT-.n115 GNDA 0.260213f
C1764 VOUT-.t55 GNDA 0.29849f
C1765 VOUT-.n116 GNDA 0.256727f
C1766 VOUT-.t90 GNDA 0.29849f
C1767 VOUT-.n117 GNDA 0.256732f
C1768 VOUT-.t128 GNDA 0.29849f
C1769 VOUT-.n118 GNDA 0.256732f
C1770 VOUT-.t25 GNDA 0.29849f
C1771 VOUT-.n119 GNDA 0.19122f
C1772 VOUT-.t149 GNDA 0.29849f
C1773 VOUT-.n120 GNDA 0.19122f
C1774 VOUT-.t43 GNDA 0.29849f
C1775 VOUT-.n121 GNDA 0.19122f
C1776 VOUT-.t80 GNDA 0.29849f
C1777 VOUT-.n122 GNDA 0.13059f
C1778 VOUT-.t60 GNDA 0.29849f
C1779 VOUT-.n123 GNDA 0.13059f
C1780 VOUT-.n124 GNDA 0.186556f
C1781 VOUT-.t68 GNDA 0.303574f
C1782 VOUT-.t94 GNDA 0.29849f
C1783 VOUT-.n125 GNDA 0.200128f
C1784 VOUT-.t59 GNDA 0.29849f
C1785 VOUT-.t41 GNDA 0.303574f
C1786 VOUT-.t19 GNDA 0.29849f
C1787 VOUT-.n126 GNDA 0.200128f
C1788 VOUT-.n127 GNDA 0.242523f
C1789 VOUT-.t31 GNDA 0.303574f
C1790 VOUT-.t58 GNDA 0.29849f
C1791 VOUT-.n128 GNDA 0.200128f
C1792 VOUT-.t161 GNDA 0.29849f
C1793 VOUT-.t143 GNDA 0.303574f
C1794 VOUT-.t116 GNDA 0.29849f
C1795 VOUT-.n129 GNDA 0.200128f
C1796 VOUT-.n130 GNDA 0.242523f
C1797 VOUT-.t132 GNDA 0.303574f
C1798 VOUT-.t159 GNDA 0.29849f
C1799 VOUT-.n131 GNDA 0.200128f
C1800 VOUT-.t114 GNDA 0.29849f
C1801 VOUT-.t101 GNDA 0.303574f
C1802 VOUT-.t76 GNDA 0.29849f
C1803 VOUT-.n132 GNDA 0.200128f
C1804 VOUT-.n133 GNDA 0.242523f
C1805 VOUT-.t26 GNDA 0.303574f
C1806 VOUT-.t53 GNDA 0.29849f
C1807 VOUT-.n134 GNDA 0.200128f
C1808 VOUT-.t153 GNDA 0.29849f
C1809 VOUT-.t138 GNDA 0.303574f
C1810 VOUT-.t111 GNDA 0.29849f
C1811 VOUT-.n135 GNDA 0.200128f
C1812 VOUT-.n136 GNDA 0.242523f
C1813 VOUT-.t126 GNDA 0.303574f
C1814 VOUT-.t152 GNDA 0.29849f
C1815 VOUT-.n137 GNDA 0.200128f
C1816 VOUT-.t109 GNDA 0.29849f
C1817 VOUT-.t97 GNDA 0.303574f
C1818 VOUT-.t69 GNDA 0.29849f
C1819 VOUT-.n138 GNDA 0.200128f
C1820 VOUT-.n139 GNDA 0.242523f
C1821 VOUT-.t30 GNDA 0.303574f
C1822 VOUT-.t120 GNDA 0.29849f
C1823 VOUT-.n140 GNDA 0.200128f
C1824 VOUT-.t85 GNDA 0.29849f
C1825 VOUT-.t140 GNDA 0.303574f
C1826 VOUT-.t50 GNDA 0.29849f
C1827 VOUT-.n141 GNDA 0.200128f
C1828 VOUT-.n142 GNDA 0.242523f
C1829 VOUT-.t64 GNDA 0.303574f
C1830 VOUT-.t157 GNDA 0.29849f
C1831 VOUT-.n143 GNDA 0.200128f
C1832 VOUT-.t118 GNDA 0.29849f
C1833 VOUT-.t32 GNDA 0.303574f
C1834 VOUT-.t82 GNDA 0.29849f
C1835 VOUT-.n144 GNDA 0.200128f
C1836 VOUT-.n145 GNDA 0.242523f
C1837 VOUT-.t24 GNDA 0.303574f
C1838 VOUT-.t112 GNDA 0.29849f
C1839 VOUT-.n146 GNDA 0.200128f
C1840 VOUT-.t77 GNDA 0.29849f
C1841 VOUT-.t133 GNDA 0.303574f
C1842 VOUT-.t45 GNDA 0.29849f
C1843 VOUT-.n147 GNDA 0.200128f
C1844 VOUT-.n148 GNDA 0.242523f
C1845 VOUT-.t123 GNDA 0.303574f
C1846 VOUT-.t71 GNDA 0.29849f
C1847 VOUT-.n149 GNDA 0.200128f
C1848 VOUT-.t39 GNDA 0.29849f
C1849 VOUT-.t92 GNDA 0.303574f
C1850 VOUT-.t148 GNDA 0.29849f
C1851 VOUT-.n150 GNDA 0.200128f
C1852 VOUT-.n151 GNDA 0.242523f
C1853 VOUT-.t21 GNDA 0.303574f
C1854 VOUT-.t107 GNDA 0.29849f
C1855 VOUT-.n152 GNDA 0.200128f
C1856 VOUT-.t70 GNDA 0.29849f
C1857 VOUT-.n153 GNDA 0.242523f
C1858 VOUT-.t38 GNDA 0.29849f
C1859 VOUT-.n154 GNDA 0.127311f
C1860 VOUT-.t127 GNDA 0.29849f
C1861 VOUT-.n155 GNDA 0.337215f
C1862 VOUT-.n156 GNDA 0.274238f
C1863 VOUT-.n157 GNDA 0.055967f
C1864 VOUT-.n158 GNDA 0.055967f
C1865 VOUT-.n159 GNDA 0.055967f
C1866 VOUT-.n160 GNDA 0.16416f
C1867 VOUT-.n161 GNDA 0.059295f
C1868 VOUT-.n162 GNDA 0.05638f
C1869 VOUT-.n164 GNDA 0.503703f
C1870 VOUT-.n165 GNDA 0.055967f
C1871 VOUT-.n166 GNDA 1.06337f
C1872 VOUT-.n170 GNDA 0.038057f
C1873 VOUT-.n171 GNDA 0.038057f
C1874 VOUT-.n172 GNDA 0.035819f
C1875 VOUT-.n173 GNDA 0.074623f
C1876 VOUT-.n174 GNDA 0.038057f
C1877 VOUT-.n175 GNDA 0.038057f
C1878 VOUT-.n177 GNDA 1.05404f
C1879 VOUT-.n178 GNDA 0.257448f
C1880 VOUT-.t0 GNDA 0.085506f
C1881 VOUT-.n179 GNDA 0.419876f
C1882 VOUT-.n180 GNDA 0.035819f
C1883 VOUT-.t18 GNDA 0.052236f
C1884 VOUT-.t4 GNDA 0.052236f
C1885 VOUT-.n181 GNDA 0.112235f
C1886 VOUT-.n182 GNDA 0.275519f
C1887 VOUT-.n183 GNDA 0.035819f
C1888 VOUT-.n184 GNDA 0.237647f
C1889 VOUT-.t1 GNDA 0.052236f
C1890 VOUT-.t17 GNDA 0.052236f
C1891 VOUT-.n185 GNDA 0.112235f
C1892 VOUT-.n186 GNDA 0.284206f
C1893 VOUT-.n187 GNDA 0.159675f
C1894 VOUT-.t2 GNDA 0.052236f
C1895 VOUT-.t3 GNDA 0.052236f
C1896 VOUT-.n188 GNDA 0.112235f
C1897 VOUT-.n189 GNDA 0.270977f
C1898 VOUT-.n190 GNDA 0.127387f
C1899 VOUT-.n191 GNDA 0.035819f
C1900 VOUT-.n192 GNDA 0.184829f
C1901 VOUT-.n193 GNDA 0.035819f
C1902 VOUT-.n194 GNDA 0.035819f
C1903 VOUT-.n195 GNDA 0.035819f
C1904 VOUT-.n196 GNDA 0.035819f
C1905 VOUT-.n197 GNDA 0.082271f
C1906 VOUT-.n198 GNDA 0.096263f
C1907 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t1 GNDA 0.0126f
C1908 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t13 GNDA 0.0126f
C1909 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n0 GNDA 0.039625f
C1910 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t2 GNDA 0.0126f
C1911 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t0 GNDA 0.0126f
C1912 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n1 GNDA 0.027028f
C1913 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n2 GNDA 1.22783f
C1914 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t14 GNDA 0.151689f
C1915 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n3 GNDA 0.061466f
C1916 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n4 GNDA 0.075408f
C1917 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t7 GNDA 0.0378f
C1918 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t12 GNDA 0.0378f
C1919 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n5 GNDA 0.080846f
C1920 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n6 GNDA 0.252186f
C1921 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t8 GNDA 0.0378f
C1922 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t3 GNDA 0.0378f
C1923 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n7 GNDA 0.080846f
C1924 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n8 GNDA 0.246038f
C1925 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n9 GNDA 0.102569f
C1926 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n10 GNDA 0.061466f
C1927 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t10 GNDA 0.0378f
C1928 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t4 GNDA 0.0378f
C1929 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n11 GNDA 0.080846f
C1930 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n12 GNDA 0.246038f
C1931 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n13 GNDA 0.043826f
C1932 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t9 GNDA 0.0378f
C1933 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t6 GNDA 0.0378f
C1934 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n14 GNDA 0.080846f
C1935 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n15 GNDA 0.246038f
C1936 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n16 GNDA 0.075408f
C1937 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t11 GNDA 0.0378f
C1938 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.t5 GNDA 0.0378f
C1939 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n17 GNDA 0.080846f
C1940 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n18 GNDA 0.249462f
C1941 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n19 GNDA 0.173897f
C1942 two_stage_opamp_dummy_magic_29_0.V_CMFB_S2.n20 GNDA 0.834277f
C1943 two_stage_opamp_dummy_magic_29_0.Vb2.n0 GNDA 0.53194f
C1944 two_stage_opamp_dummy_magic_29_0.Vb2.n1 GNDA 0.542995f
C1945 two_stage_opamp_dummy_magic_29_0.Vb2.n2 GNDA 0.396191f
C1946 two_stage_opamp_dummy_magic_29_0.Vb2.n3 GNDA 0.542995f
C1947 two_stage_opamp_dummy_magic_29_0.Vb2.n4 GNDA 0.960424f
C1948 two_stage_opamp_dummy_magic_29_0.Vb2.n5 GNDA 0.790732f
C1949 two_stage_opamp_dummy_magic_29_0.Vb2.t2 GNDA 0.018374f
C1950 two_stage_opamp_dummy_magic_29_0.Vb2.t8 GNDA 0.018374f
C1951 two_stage_opamp_dummy_magic_29_0.Vb2.n6 GNDA 0.061604f
C1952 two_stage_opamp_dummy_magic_29_0.Vb2.t0 GNDA 0.018374f
C1953 two_stage_opamp_dummy_magic_29_0.Vb2.t1 GNDA 0.018374f
C1954 two_stage_opamp_dummy_magic_29_0.Vb2.n7 GNDA 0.059914f
C1955 two_stage_opamp_dummy_magic_29_0.Vb2.n8 GNDA 0.557382f
C1956 two_stage_opamp_dummy_magic_29_0.Vb2.t7 GNDA 0.018374f
C1957 two_stage_opamp_dummy_magic_29_0.Vb2.t10 GNDA 0.018374f
C1958 two_stage_opamp_dummy_magic_29_0.Vb2.n9 GNDA 0.059914f
C1959 two_stage_opamp_dummy_magic_29_0.Vb2.n10 GNDA 0.369107f
C1960 two_stage_opamp_dummy_magic_29_0.Vb2.t9 GNDA 0.018374f
C1961 two_stage_opamp_dummy_magic_29_0.Vb2.t6 GNDA 0.018374f
C1962 two_stage_opamp_dummy_magic_29_0.Vb2.n11 GNDA 0.059914f
C1963 two_stage_opamp_dummy_magic_29_0.Vb2.n12 GNDA 1.14638f
C1964 two_stage_opamp_dummy_magic_29_0.Vb2.t18 GNDA 0.117836f
C1965 two_stage_opamp_dummy_magic_29_0.Vb2.t31 GNDA 0.117805f
C1966 two_stage_opamp_dummy_magic_29_0.Vb2.t22 GNDA 0.117805f
C1967 two_stage_opamp_dummy_magic_29_0.Vb2.t13 GNDA 0.117805f
C1968 two_stage_opamp_dummy_magic_29_0.Vb2.t21 GNDA 0.117805f
C1969 two_stage_opamp_dummy_magic_29_0.Vb2.t12 GNDA 0.117805f
C1970 two_stage_opamp_dummy_magic_29_0.Vb2.t25 GNDA 0.117805f
C1971 two_stage_opamp_dummy_magic_29_0.Vb2.t16 GNDA 0.117805f
C1972 two_stage_opamp_dummy_magic_29_0.Vb2.t28 GNDA 0.117805f
C1973 two_stage_opamp_dummy_magic_29_0.Vb2.t11 GNDA 0.117805f
C1974 two_stage_opamp_dummy_magic_29_0.Vb2.t17 GNDA 0.117836f
C1975 two_stage_opamp_dummy_magic_29_0.Vb2.t26 GNDA 0.117805f
C1976 two_stage_opamp_dummy_magic_29_0.Vb2.t19 GNDA 0.117805f
C1977 two_stage_opamp_dummy_magic_29_0.Vb2.t30 GNDA 0.117805f
C1978 two_stage_opamp_dummy_magic_29_0.Vb2.t14 GNDA 0.117805f
C1979 two_stage_opamp_dummy_magic_29_0.Vb2.t23 GNDA 0.117805f
C1980 two_stage_opamp_dummy_magic_29_0.Vb2.t32 GNDA 0.117805f
C1981 two_stage_opamp_dummy_magic_29_0.Vb2.t27 GNDA 0.117805f
C1982 two_stage_opamp_dummy_magic_29_0.Vb2.t15 GNDA 0.117805f
C1983 two_stage_opamp_dummy_magic_29_0.Vb2.t24 GNDA 0.117805f
C1984 two_stage_opamp_dummy_magic_29_0.Vb2.t5 GNDA 0.064307f
C1985 two_stage_opamp_dummy_magic_29_0.Vb2.t3 GNDA 0.064307f
C1986 two_stage_opamp_dummy_magic_29_0.Vb2.n13 GNDA 0.136813f
C1987 two_stage_opamp_dummy_magic_29_0.Vb2.t4 GNDA 0.12168f
C1988 two_stage_opamp_dummy_magic_29_0.Vb2.n14 GNDA 0.520543f
C1989 two_stage_opamp_dummy_magic_29_0.Vb2.n15 GNDA 0.716429f
C1990 two_stage_opamp_dummy_magic_29_0.Vb2.t20 GNDA 0.073864f
C1991 two_stage_opamp_dummy_magic_29_0.Vb2.n16 GNDA 0.672925f
C1992 two_stage_opamp_dummy_magic_29_0.Vb2.t29 GNDA 0.118193f
C1993 two_stage_opamp_dummy_magic_29_0.Vb2.n17 GNDA 0.646787f
C1994 two_stage_opamp_dummy_magic_29_0.Vb2.n18 GNDA 1.5502f
C1995 bgr_11_0.VB2_CUR_BIAS GNDA 4.23131f
C1996 two_stage_opamp_dummy_magic_29_0.V_source.n0 GNDA 0.041306f
C1997 two_stage_opamp_dummy_magic_29_0.V_source.n1 GNDA 0.540854f
C1998 two_stage_opamp_dummy_magic_29_0.V_source.n2 GNDA 0.586883f
C1999 two_stage_opamp_dummy_magic_29_0.V_source.n3 GNDA 0.339486f
C2000 two_stage_opamp_dummy_magic_29_0.V_source.n4 GNDA 0.304203f
C2001 two_stage_opamp_dummy_magic_29_0.V_source.t13 GNDA 0.021514f
C2002 two_stage_opamp_dummy_magic_29_0.V_source.t3 GNDA 0.021514f
C2003 two_stage_opamp_dummy_magic_29_0.V_source.n5 GNDA 0.045993f
C2004 two_stage_opamp_dummy_magic_29_0.V_source.n6 GNDA 0.199232f
C2005 two_stage_opamp_dummy_magic_29_0.V_source.n7 GNDA 0.04198f
C2006 two_stage_opamp_dummy_magic_29_0.V_source.t36 GNDA 0.021514f
C2007 two_stage_opamp_dummy_magic_29_0.V_source.t27 GNDA 0.021514f
C2008 two_stage_opamp_dummy_magic_29_0.V_source.n8 GNDA 0.045993f
C2009 two_stage_opamp_dummy_magic_29_0.V_source.n9 GNDA 0.164071f
C2010 two_stage_opamp_dummy_magic_29_0.V_source.n10 GNDA 0.153086f
C2011 two_stage_opamp_dummy_magic_29_0.V_source.n11 GNDA 0.153086f
C2012 two_stage_opamp_dummy_magic_29_0.V_source.n12 GNDA 0.147729f
C2013 two_stage_opamp_dummy_magic_29_0.V_source.n13 GNDA 0.069673f
C2014 two_stage_opamp_dummy_magic_29_0.V_source.n14 GNDA 0.046931f
C2015 two_stage_opamp_dummy_magic_29_0.V_source.t14 GNDA 0.012908f
C2016 two_stage_opamp_dummy_magic_29_0.V_source.t19 GNDA 0.012908f
C2017 two_stage_opamp_dummy_magic_29_0.V_source.n15 GNDA 0.028087f
C2018 two_stage_opamp_dummy_magic_29_0.V_source.n16 GNDA 0.117879f
C2019 two_stage_opamp_dummy_magic_29_0.V_source.t4 GNDA 0.012908f
C2020 two_stage_opamp_dummy_magic_29_0.V_source.t15 GNDA 0.012908f
C2021 two_stage_opamp_dummy_magic_29_0.V_source.n17 GNDA 0.028087f
C2022 two_stage_opamp_dummy_magic_29_0.V_source.n18 GNDA 0.113801f
C2023 two_stage_opamp_dummy_magic_29_0.V_source.n19 GNDA 0.069673f
C2024 two_stage_opamp_dummy_magic_29_0.V_source.n20 GNDA 0.054121f
C2025 two_stage_opamp_dummy_magic_29_0.V_source.t20 GNDA 0.012908f
C2026 two_stage_opamp_dummy_magic_29_0.V_source.t16 GNDA 0.012908f
C2027 two_stage_opamp_dummy_magic_29_0.V_source.n21 GNDA 0.028087f
C2028 two_stage_opamp_dummy_magic_29_0.V_source.n22 GNDA 0.113801f
C2029 two_stage_opamp_dummy_magic_29_0.V_source.n23 GNDA 0.027589f
C2030 two_stage_opamp_dummy_magic_29_0.V_source.n24 GNDA 0.027589f
C2031 two_stage_opamp_dummy_magic_29_0.V_source.t0 GNDA 0.012908f
C2032 two_stage_opamp_dummy_magic_29_0.V_source.t21 GNDA 0.012908f
C2033 two_stage_opamp_dummy_magic_29_0.V_source.n25 GNDA 0.028087f
C2034 two_stage_opamp_dummy_magic_29_0.V_source.n26 GNDA 0.085239f
C2035 two_stage_opamp_dummy_magic_29_0.V_source.t18 GNDA 0.012908f
C2036 two_stage_opamp_dummy_magic_29_0.V_source.t17 GNDA 0.012908f
C2037 two_stage_opamp_dummy_magic_29_0.V_source.n27 GNDA 0.028087f
C2038 two_stage_opamp_dummy_magic_29_0.V_source.n28 GNDA 0.085239f
C2039 two_stage_opamp_dummy_magic_29_0.V_source.n29 GNDA 0.069756f
C2040 two_stage_opamp_dummy_magic_29_0.V_source.t12 GNDA 0.012908f
C2041 two_stage_opamp_dummy_magic_29_0.V_source.t40 GNDA 0.012908f
C2042 two_stage_opamp_dummy_magic_29_0.V_source.n30 GNDA 0.028087f
C2043 two_stage_opamp_dummy_magic_29_0.V_source.n31 GNDA 0.085239f
C2044 two_stage_opamp_dummy_magic_29_0.V_source.n32 GNDA 0.069756f
C2045 two_stage_opamp_dummy_magic_29_0.V_source.t1 GNDA 0.012908f
C2046 two_stage_opamp_dummy_magic_29_0.V_source.t10 GNDA 0.012908f
C2047 two_stage_opamp_dummy_magic_29_0.V_source.n33 GNDA 0.028087f
C2048 two_stage_opamp_dummy_magic_29_0.V_source.n34 GNDA 0.085239f
C2049 two_stage_opamp_dummy_magic_29_0.V_source.n35 GNDA 0.027589f
C2050 two_stage_opamp_dummy_magic_29_0.V_source.t7 GNDA 0.012908f
C2051 two_stage_opamp_dummy_magic_29_0.V_source.t11 GNDA 0.012908f
C2052 two_stage_opamp_dummy_magic_29_0.V_source.n36 GNDA 0.028087f
C2053 two_stage_opamp_dummy_magic_29_0.V_source.n37 GNDA 0.117879f
C2054 two_stage_opamp_dummy_magic_29_0.V_source.t6 GNDA 0.012908f
C2055 two_stage_opamp_dummy_magic_29_0.V_source.t2 GNDA 0.012908f
C2056 two_stage_opamp_dummy_magic_29_0.V_source.n38 GNDA 0.028087f
C2057 two_stage_opamp_dummy_magic_29_0.V_source.n39 GNDA 0.113801f
C2058 two_stage_opamp_dummy_magic_29_0.V_source.n40 GNDA 0.046931f
C2059 two_stage_opamp_dummy_magic_29_0.V_source.n41 GNDA 0.027589f
C2060 two_stage_opamp_dummy_magic_29_0.V_source.t8 GNDA 0.012908f
C2061 two_stage_opamp_dummy_magic_29_0.V_source.t9 GNDA 0.012908f
C2062 two_stage_opamp_dummy_magic_29_0.V_source.n42 GNDA 0.028087f
C2063 two_stage_opamp_dummy_magic_29_0.V_source.n43 GNDA 0.113801f
C2064 two_stage_opamp_dummy_magic_29_0.V_source.n44 GNDA 0.054121f
C2065 two_stage_opamp_dummy_magic_29_0.V_source.n45 GNDA 0.147729f
C2066 two_stage_opamp_dummy_magic_29_0.V_source.t29 GNDA 0.021514f
C2067 two_stage_opamp_dummy_magic_29_0.V_source.t37 GNDA 0.021514f
C2068 two_stage_opamp_dummy_magic_29_0.V_source.n46 GNDA 0.045993f
C2069 two_stage_opamp_dummy_magic_29_0.V_source.n47 GNDA 0.164071f
C2070 two_stage_opamp_dummy_magic_29_0.V_source.t33 GNDA 0.021514f
C2071 two_stage_opamp_dummy_magic_29_0.V_source.t23 GNDA 0.021514f
C2072 two_stage_opamp_dummy_magic_29_0.V_source.n48 GNDA 0.045993f
C2073 two_stage_opamp_dummy_magic_29_0.V_source.n49 GNDA 0.164071f
C2074 two_stage_opamp_dummy_magic_29_0.V_source.n50 GNDA 0.041306f
C2075 two_stage_opamp_dummy_magic_29_0.V_source.t38 GNDA 0.021514f
C2076 two_stage_opamp_dummy_magic_29_0.V_source.t28 GNDA 0.021514f
C2077 two_stage_opamp_dummy_magic_29_0.V_source.n52 GNDA 0.045993f
C2078 two_stage_opamp_dummy_magic_29_0.V_source.n53 GNDA 0.164071f
C2079 two_stage_opamp_dummy_magic_29_0.V_source.n54 GNDA 0.153086f
C2080 two_stage_opamp_dummy_magic_29_0.V_source.t26 GNDA 0.021514f
C2081 two_stage_opamp_dummy_magic_29_0.V_source.t30 GNDA 0.021514f
C2082 two_stage_opamp_dummy_magic_29_0.V_source.n55 GNDA 0.045993f
C2083 two_stage_opamp_dummy_magic_29_0.V_source.n56 GNDA 0.164071f
C2084 two_stage_opamp_dummy_magic_29_0.V_source.n57 GNDA 0.153086f
C2085 two_stage_opamp_dummy_magic_29_0.V_source.n58 GNDA 0.95652f
C2086 two_stage_opamp_dummy_magic_29_0.V_source.t5 GNDA 0.047788f
C2087 two_stage_opamp_dummy_magic_29_0.V_source.n59 GNDA 1.55874f
C2088 two_stage_opamp_dummy_magic_29_0.V_source.n60 GNDA 0.477603f
C2089 two_stage_opamp_dummy_magic_29_0.V_source.n61 GNDA 0.041306f
C2090 two_stage_opamp_dummy_magic_29_0.V_source.n62 GNDA 0.041306f
C2091 two_stage_opamp_dummy_magic_29_0.V_source.n64 GNDA 0.649838f
C2092 two_stage_opamp_dummy_magic_29_0.V_source.n65 GNDA 0.63917f
C2093 two_stage_opamp_dummy_magic_29_0.V_source.n66 GNDA 0.153086f
C2094 two_stage_opamp_dummy_magic_29_0.V_source.t32 GNDA 0.021514f
C2095 two_stage_opamp_dummy_magic_29_0.V_source.t22 GNDA 0.021514f
C2096 two_stage_opamp_dummy_magic_29_0.V_source.n67 GNDA 0.045993f
C2097 two_stage_opamp_dummy_magic_29_0.V_source.n68 GNDA 0.164071f
C2098 two_stage_opamp_dummy_magic_29_0.V_source.n69 GNDA 0.118148f
C2099 two_stage_opamp_dummy_magic_29_0.V_source.t39 GNDA 0.021514f
C2100 two_stage_opamp_dummy_magic_29_0.V_source.t24 GNDA 0.021514f
C2101 two_stage_opamp_dummy_magic_29_0.V_source.n70 GNDA 0.045993f
C2102 two_stage_opamp_dummy_magic_29_0.V_source.n71 GNDA 0.193086f
C2103 two_stage_opamp_dummy_magic_29_0.V_source.n72 GNDA 0.153087f
C2104 two_stage_opamp_dummy_magic_29_0.V_source.t34 GNDA 0.021514f
C2105 two_stage_opamp_dummy_magic_29_0.V_source.t31 GNDA 0.021514f
C2106 two_stage_opamp_dummy_magic_29_0.V_source.n73 GNDA 0.045993f
C2107 two_stage_opamp_dummy_magic_29_0.V_source.n74 GNDA 0.193086f
C2108 two_stage_opamp_dummy_magic_29_0.V_source.n75 GNDA 0.153086f
C2109 two_stage_opamp_dummy_magic_29_0.V_source.n76 GNDA 0.153086f
C2110 two_stage_opamp_dummy_magic_29_0.V_source.t35 GNDA 0.021514f
C2111 two_stage_opamp_dummy_magic_29_0.V_source.t25 GNDA 0.021514f
C2112 two_stage_opamp_dummy_magic_29_0.V_source.n77 GNDA 0.045993f
C2113 two_stage_opamp_dummy_magic_29_0.V_source.n78 GNDA 0.193086f
C2114 two_stage_opamp_dummy_magic_29_0.V_source.n79 GNDA 0.066185f
C2115 two_stage_opamp_dummy_magic_29_0.V_source.n80 GNDA 0.113174f
C2116 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n0 GNDA 6.84231f
C2117 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n1 GNDA 11.403501f
C2118 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n2 GNDA 0.093773f
C2119 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n3 GNDA 6.53761f
C2120 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t11 GNDA 0.0117f
C2121 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t1 GNDA 0.0117f
C2122 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n4 GNDA 0.025895f
C2123 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n5 GNDA 0.121918f
C2124 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t27 GNDA 0.020768f
C2125 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t16 GNDA 0.020768f
C2126 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t25 GNDA 0.020768f
C2127 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t15 GNDA 0.020768f
C2128 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t24 GNDA 0.020768f
C2129 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t13 GNDA 0.020768f
C2130 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t22 GNDA 0.020768f
C2131 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t26 GNDA 0.024239f
C2132 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n6 GNDA 0.022854f
C2133 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n7 GNDA 0.014333f
C2134 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n8 GNDA 0.014333f
C2135 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n9 GNDA 0.014333f
C2136 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n10 GNDA 0.014333f
C2137 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n11 GNDA 0.014333f
C2138 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n12 GNDA 0.013412f
C2139 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n13 GNDA 0.012145f
C2140 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n14 GNDA 0.0156f
C2141 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n15 GNDA 0.0156f
C2142 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n16 GNDA 0.028327f
C2143 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n17 GNDA 0.089319f
C2144 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n18 GNDA 0.0156f
C2145 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n19 GNDA 0.093322f
C2146 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n20 GNDA 0.089319f
C2147 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n21 GNDA 0.0156f
C2148 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n22 GNDA 0.093781f
C2149 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t0 GNDA 0.0117f
C2150 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t10 GNDA 0.0117f
C2151 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n23 GNDA 0.025895f
C2152 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n24 GNDA 0.131005f
C2153 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t21 GNDA 0.020768f
C2154 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t18 GNDA 0.020768f
C2155 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n25 GNDA 0.013412f
C2156 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n26 GNDA 0.013412f
C2157 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t12 GNDA 0.020768f
C2158 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t29 GNDA 0.020768f
C2159 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t19 GNDA 0.020768f
C2160 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t30 GNDA 0.020768f
C2161 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t20 GNDA 0.020768f
C2162 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t31 GNDA 0.020768f
C2163 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t23 GNDA 0.020768f
C2164 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t14 GNDA 0.020768f
C2165 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t17 GNDA 0.020768f
C2166 two_stage_opamp_dummy_magic_29_0.V_tail_gate.t28 GNDA 0.024239f
C2167 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n27 GNDA 0.022854f
C2168 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n28 GNDA 0.014333f
C2169 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n29 GNDA 0.014333f
C2170 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n30 GNDA 0.014333f
C2171 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n31 GNDA 0.014333f
C2172 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n32 GNDA 0.014333f
C2173 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n33 GNDA 0.014333f
C2174 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n34 GNDA 0.014333f
C2175 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n35 GNDA 0.013412f
C2176 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n36 GNDA 0.012145f
C2177 two_stage_opamp_dummy_magic_29_0.V_tail_gate.n37 GNDA 0.128032f
C2178 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t13 GNDA 0.010731f
C2179 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t14 GNDA 0.010731f
C2180 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n0 GNDA 0.033748f
C2181 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t12 GNDA 0.010731f
C2182 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t0 GNDA 0.010731f
C2183 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n1 GNDA 0.023019f
C2184 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n2 GNDA 0.754767f
C2185 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t11 GNDA 0.129193f
C2186 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n3 GNDA 0.05235f
C2187 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n4 GNDA 0.064224f
C2188 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t10 GNDA 0.032194f
C2189 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t3 GNDA 0.032194f
C2190 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n5 GNDA 0.068856f
C2191 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n6 GNDA 0.214783f
C2192 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t7 GNDA 0.032194f
C2193 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t2 GNDA 0.032194f
C2194 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n7 GNDA 0.068856f
C2195 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n8 GNDA 0.209547f
C2196 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n9 GNDA 0.087357f
C2197 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n10 GNDA 0.05235f
C2198 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t6 GNDA 0.032194f
C2199 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t1 GNDA 0.032194f
C2200 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n11 GNDA 0.068856f
C2201 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n12 GNDA 0.209547f
C2202 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n13 GNDA 0.037326f
C2203 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t9 GNDA 0.032194f
C2204 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t5 GNDA 0.032194f
C2205 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n14 GNDA 0.068856f
C2206 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n15 GNDA 0.209547f
C2207 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n16 GNDA 0.064224f
C2208 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t8 GNDA 0.032194f
C2209 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.t4 GNDA 0.032194f
C2210 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n17 GNDA 0.068856f
C2211 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n18 GNDA 0.212464f
C2212 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n19 GNDA 0.148104f
C2213 two_stage_opamp_dummy_magic_29_0.V_CMFB_S4.n20 GNDA 6.12768f
C2214 bgr_11_0.V_CMFB_S4 GNDA 2.86063f
C2215 two_stage_opamp_dummy_magic_29_0.Y.n0 GNDA 0.194525f
C2216 two_stage_opamp_dummy_magic_29_0.Y.n1 GNDA 0.08603f
C2217 two_stage_opamp_dummy_magic_29_0.Y.n2 GNDA 0.237753f
C2218 two_stage_opamp_dummy_magic_29_0.Y.n3 GNDA 0.815021f
C2219 two_stage_opamp_dummy_magic_29_0.Y.n4 GNDA 0.08603f
C2220 two_stage_opamp_dummy_magic_29_0.Y.n5 GNDA 0.08603f
C2221 two_stage_opamp_dummy_magic_29_0.Y.t15 GNDA 0.023158f
C2222 two_stage_opamp_dummy_magic_29_0.Y.t23 GNDA 0.023158f
C2223 two_stage_opamp_dummy_magic_29_0.Y.n6 GNDA 0.068053f
C2224 two_stage_opamp_dummy_magic_29_0.Y.t16 GNDA 0.023158f
C2225 two_stage_opamp_dummy_magic_29_0.Y.t13 GNDA 0.023158f
C2226 two_stage_opamp_dummy_magic_29_0.Y.n7 GNDA 0.066733f
C2227 two_stage_opamp_dummy_magic_29_0.Y.n8 GNDA 0.441071f
C2228 two_stage_opamp_dummy_magic_29_0.Y.t4 GNDA 0.023158f
C2229 two_stage_opamp_dummy_magic_29_0.Y.t14 GNDA 0.023158f
C2230 two_stage_opamp_dummy_magic_29_0.Y.n9 GNDA 0.066733f
C2231 two_stage_opamp_dummy_magic_29_0.Y.n10 GNDA 0.232002f
C2232 two_stage_opamp_dummy_magic_29_0.Y.t11 GNDA 0.023158f
C2233 two_stage_opamp_dummy_magic_29_0.Y.t5 GNDA 0.023158f
C2234 two_stage_opamp_dummy_magic_29_0.Y.n11 GNDA 0.066733f
C2235 two_stage_opamp_dummy_magic_29_0.Y.n12 GNDA 0.232002f
C2236 two_stage_opamp_dummy_magic_29_0.Y.t12 GNDA 0.023158f
C2237 two_stage_opamp_dummy_magic_29_0.Y.t8 GNDA 0.023158f
C2238 two_stage_opamp_dummy_magic_29_0.Y.n13 GNDA 0.066733f
C2239 two_stage_opamp_dummy_magic_29_0.Y.n14 GNDA 0.232002f
C2240 two_stage_opamp_dummy_magic_29_0.Y.t22 GNDA 0.023158f
C2241 two_stage_opamp_dummy_magic_29_0.Y.t24 GNDA 0.023158f
C2242 two_stage_opamp_dummy_magic_29_0.Y.n15 GNDA 0.066733f
C2243 two_stage_opamp_dummy_magic_29_0.Y.n16 GNDA 0.431159f
C2244 two_stage_opamp_dummy_magic_29_0.Y.n17 GNDA 0.287483f
C2245 two_stage_opamp_dummy_magic_29_0.Y.n18 GNDA 0.644415f
C2246 two_stage_opamp_dummy_magic_29_0.Y.n19 GNDA 0.496725f
C2247 two_stage_opamp_dummy_magic_29_0.Y.n20 GNDA 0.237753f
C2248 two_stage_opamp_dummy_magic_29_0.Y.n21 GNDA 0.417266f
C2249 two_stage_opamp_dummy_magic_29_0.Y.n22 GNDA 0.237753f
C2250 two_stage_opamp_dummy_magic_29_0.Y.n23 GNDA 0.237753f
C2251 two_stage_opamp_dummy_magic_29_0.Y.n24 GNDA 0.237753f
C2252 two_stage_opamp_dummy_magic_29_0.Y.n25 GNDA 0.146616f
C2253 two_stage_opamp_dummy_magic_29_0.Y.n27 GNDA 0.074105f
C2254 two_stage_opamp_dummy_magic_29_0.Y.n28 GNDA 0.074105f
C2255 two_stage_opamp_dummy_magic_29_0.Y.n30 GNDA 0.074105f
C2256 two_stage_opamp_dummy_magic_29_0.Y.n32 GNDA 0.074105f
C2257 two_stage_opamp_dummy_magic_29_0.Y.n34 GNDA 0.172912f
C2258 two_stage_opamp_dummy_magic_29_0.Y.n36 GNDA 0.074105f
C2259 two_stage_opamp_dummy_magic_29_0.Y.n37 GNDA 0.074105f
C2260 two_stage_opamp_dummy_magic_29_0.Y.n38 GNDA 0.073409f
C2261 two_stage_opamp_dummy_magic_29_0.Y.n39 GNDA 0.074105f
C2262 two_stage_opamp_dummy_magic_29_0.Y.t0 GNDA 0.640789f
C2263 two_stage_opamp_dummy_magic_29_0.Y.n40 GNDA 0.074105f
C2264 two_stage_opamp_dummy_magic_29_0.Y.n41 GNDA 0.074105f
C2265 two_stage_opamp_dummy_magic_29_0.Y.n43 GNDA 0.687542f
C2266 two_stage_opamp_dummy_magic_29_0.Y.n45 GNDA 0.643787f
C2267 two_stage_opamp_dummy_magic_29_0.Y.n46 GNDA 0.024538f
C2268 two_stage_opamp_dummy_magic_29_0.Y.n47 GNDA 0.024702f
C2269 two_stage_opamp_dummy_magic_29_0.Y.n48 GNDA 0.024702f
C2270 two_stage_opamp_dummy_magic_29_0.Y.t35 GNDA 0.101894f
C2271 two_stage_opamp_dummy_magic_29_0.Y.t42 GNDA 0.101894f
C2272 two_stage_opamp_dummy_magic_29_0.Y.t27 GNDA 0.101894f
C2273 two_stage_opamp_dummy_magic_29_0.Y.t43 GNDA 0.101894f
C2274 two_stage_opamp_dummy_magic_29_0.Y.t29 GNDA 0.108524f
C2275 two_stage_opamp_dummy_magic_29_0.Y.n49 GNDA 0.086001f
C2276 two_stage_opamp_dummy_magic_29_0.Y.n50 GNDA 0.048631f
C2277 two_stage_opamp_dummy_magic_29_0.Y.n51 GNDA 0.048631f
C2278 two_stage_opamp_dummy_magic_29_0.Y.n52 GNDA 0.04371f
C2279 two_stage_opamp_dummy_magic_29_0.Y.t46 GNDA 0.101894f
C2280 two_stage_opamp_dummy_magic_29_0.Y.t32 GNDA 0.101894f
C2281 two_stage_opamp_dummy_magic_29_0.Y.t44 GNDA 0.101894f
C2282 two_stage_opamp_dummy_magic_29_0.Y.t30 GNDA 0.101894f
C2283 two_stage_opamp_dummy_magic_29_0.Y.t38 GNDA 0.108524f
C2284 two_stage_opamp_dummy_magic_29_0.Y.n53 GNDA 0.086001f
C2285 two_stage_opamp_dummy_magic_29_0.Y.n54 GNDA 0.048631f
C2286 two_stage_opamp_dummy_magic_29_0.Y.n55 GNDA 0.048631f
C2287 two_stage_opamp_dummy_magic_29_0.Y.n56 GNDA 0.04371f
C2288 two_stage_opamp_dummy_magic_29_0.Y.n57 GNDA 0.010496f
C2289 two_stage_opamp_dummy_magic_29_0.Y.n58 GNDA 0.024866f
C2290 two_stage_opamp_dummy_magic_29_0.Y.n59 GNDA 0.058532f
C2291 two_stage_opamp_dummy_magic_29_0.Y.n60 GNDA 0.033384f
C2292 two_stage_opamp_dummy_magic_29_0.Y.n61 GNDA 0.037886f
C2293 two_stage_opamp_dummy_magic_29_0.Y.n62 GNDA 1.02357f
C2294 two_stage_opamp_dummy_magic_29_0.Y.t37 GNDA 0.049789f
C2295 two_stage_opamp_dummy_magic_29_0.Y.t52 GNDA 0.049789f
C2296 two_stage_opamp_dummy_magic_29_0.Y.t40 GNDA 0.049789f
C2297 two_stage_opamp_dummy_magic_29_0.Y.t54 GNDA 0.049789f
C2298 two_stage_opamp_dummy_magic_29_0.Y.t31 GNDA 0.049789f
C2299 two_stage_opamp_dummy_magic_29_0.Y.t45 GNDA 0.049789f
C2300 two_stage_opamp_dummy_magic_29_0.Y.t34 GNDA 0.049789f
C2301 two_stage_opamp_dummy_magic_29_0.Y.t48 GNDA 0.056602f
C2302 two_stage_opamp_dummy_magic_29_0.Y.n64 GNDA 0.051082f
C2303 two_stage_opamp_dummy_magic_29_0.Y.n65 GNDA 0.031263f
C2304 two_stage_opamp_dummy_magic_29_0.Y.n66 GNDA 0.031263f
C2305 two_stage_opamp_dummy_magic_29_0.Y.n67 GNDA 0.031263f
C2306 two_stage_opamp_dummy_magic_29_0.Y.n68 GNDA 0.031263f
C2307 two_stage_opamp_dummy_magic_29_0.Y.n69 GNDA 0.031263f
C2308 two_stage_opamp_dummy_magic_29_0.Y.n70 GNDA 0.026342f
C2309 two_stage_opamp_dummy_magic_29_0.Y.t49 GNDA 0.049789f
C2310 two_stage_opamp_dummy_magic_29_0.Y.t25 GNDA 0.056602f
C2311 two_stage_opamp_dummy_magic_29_0.Y.n71 GNDA 0.046161f
C2312 two_stage_opamp_dummy_magic_29_0.Y.n72 GNDA 0.012791f
C2313 two_stage_opamp_dummy_magic_29_0.Y.t39 GNDA 0.032421f
C2314 two_stage_opamp_dummy_magic_29_0.Y.t53 GNDA 0.032421f
C2315 two_stage_opamp_dummy_magic_29_0.Y.t41 GNDA 0.032421f
C2316 two_stage_opamp_dummy_magic_29_0.Y.t26 GNDA 0.032421f
C2317 two_stage_opamp_dummy_magic_29_0.Y.t33 GNDA 0.032421f
C2318 two_stage_opamp_dummy_magic_29_0.Y.t47 GNDA 0.032421f
C2319 two_stage_opamp_dummy_magic_29_0.Y.t36 GNDA 0.032421f
C2320 two_stage_opamp_dummy_magic_29_0.Y.t50 GNDA 0.039368f
C2321 two_stage_opamp_dummy_magic_29_0.Y.n73 GNDA 0.039368f
C2322 two_stage_opamp_dummy_magic_29_0.Y.n74 GNDA 0.025474f
C2323 two_stage_opamp_dummy_magic_29_0.Y.n75 GNDA 0.025474f
C2324 two_stage_opamp_dummy_magic_29_0.Y.n76 GNDA 0.025474f
C2325 two_stage_opamp_dummy_magic_29_0.Y.n77 GNDA 0.025474f
C2326 two_stage_opamp_dummy_magic_29_0.Y.n78 GNDA 0.025474f
C2327 two_stage_opamp_dummy_magic_29_0.Y.n79 GNDA 0.020552f
C2328 two_stage_opamp_dummy_magic_29_0.Y.t51 GNDA 0.032421f
C2329 two_stage_opamp_dummy_magic_29_0.Y.t28 GNDA 0.039368f
C2330 two_stage_opamp_dummy_magic_29_0.Y.n80 GNDA 0.034447f
C2331 two_stage_opamp_dummy_magic_29_0.Y.n81 GNDA 0.012791f
C2332 two_stage_opamp_dummy_magic_29_0.Y.n82 GNDA 0.079795f
C2333 two_stage_opamp_dummy_magic_29_0.Y.n83 GNDA 0.074105f
C2334 two_stage_opamp_dummy_magic_29_0.Y.n84 GNDA 2.18995f
C2335 two_stage_opamp_dummy_magic_29_0.Y.n85 GNDA 0.453893f
C2336 two_stage_opamp_dummy_magic_29_0.Y.n87 GNDA 0.463156f
C2337 two_stage_opamp_dummy_magic_29_0.Y.n88 GNDA 0.463156f
C2338 two_stage_opamp_dummy_magic_29_0.Y.n91 GNDA 0.083312f
C2339 two_stage_opamp_dummy_magic_29_0.Y.n92 GNDA 0.083312f
C2340 two_stage_opamp_dummy_magic_29_0.Y.t19 GNDA 0.054035f
C2341 two_stage_opamp_dummy_magic_29_0.Y.t20 GNDA 0.054035f
C2342 two_stage_opamp_dummy_magic_29_0.Y.n93 GNDA 0.110534f
C2343 two_stage_opamp_dummy_magic_29_0.Y.n94 GNDA 0.35586f
C2344 two_stage_opamp_dummy_magic_29_0.Y.n95 GNDA 0.138043f
C2345 two_stage_opamp_dummy_magic_29_0.Y.t18 GNDA 0.054035f
C2346 two_stage_opamp_dummy_magic_29_0.Y.t6 GNDA 0.054035f
C2347 two_stage_opamp_dummy_magic_29_0.Y.n96 GNDA 0.110534f
C2348 two_stage_opamp_dummy_magic_29_0.Y.n97 GNDA 0.348103f
C2349 two_stage_opamp_dummy_magic_29_0.Y.n98 GNDA 0.138043f
C2350 two_stage_opamp_dummy_magic_29_0.Y.t9 GNDA 0.054035f
C2351 two_stage_opamp_dummy_magic_29_0.Y.t17 GNDA 0.054035f
C2352 two_stage_opamp_dummy_magic_29_0.Y.n99 GNDA 0.110534f
C2353 two_stage_opamp_dummy_magic_29_0.Y.n100 GNDA 0.348103f
C2354 two_stage_opamp_dummy_magic_29_0.Y.n101 GNDA 0.083312f
C2355 two_stage_opamp_dummy_magic_29_0.Y.n102 GNDA 0.083312f
C2356 two_stage_opamp_dummy_magic_29_0.Y.t1 GNDA 0.054035f
C2357 two_stage_opamp_dummy_magic_29_0.Y.t3 GNDA 0.054035f
C2358 two_stage_opamp_dummy_magic_29_0.Y.n103 GNDA 0.110534f
C2359 two_stage_opamp_dummy_magic_29_0.Y.n104 GNDA 0.348103f
C2360 two_stage_opamp_dummy_magic_29_0.Y.n105 GNDA 0.083312f
C2361 two_stage_opamp_dummy_magic_29_0.Y.t10 GNDA 0.054035f
C2362 two_stage_opamp_dummy_magic_29_0.Y.t7 GNDA 0.054035f
C2363 two_stage_opamp_dummy_magic_29_0.Y.n106 GNDA 0.110534f
C2364 two_stage_opamp_dummy_magic_29_0.Y.n107 GNDA 0.348103f
C2365 two_stage_opamp_dummy_magic_29_0.Y.n108 GNDA 0.138043f
C2366 two_stage_opamp_dummy_magic_29_0.Y.t21 GNDA 0.054035f
C2367 two_stage_opamp_dummy_magic_29_0.Y.t2 GNDA 0.054035f
C2368 two_stage_opamp_dummy_magic_29_0.Y.n109 GNDA 0.110534f
C2369 two_stage_opamp_dummy_magic_29_0.Y.n110 GNDA 0.351981f
C2370 two_stage_opamp_dummy_magic_29_0.Y.n111 GNDA 0.220104f
C2371 two_stage_opamp_dummy_magic_29_0.Y.n112 GNDA 0.619696f
C2372 two_stage_opamp_dummy_magic_29_0.Y.n114 GNDA 0.172912f
C2373 two_stage_opamp_dummy_magic_29_0.Y.n116 GNDA 0.074105f
C2374 two_stage_opamp_dummy_magic_29_0.Y.n117 GNDA 1.3941f
C2375 two_stage_opamp_dummy_magic_29_0.Y.n118 GNDA 1.42652f
C2376 two_stage_opamp_dummy_magic_29_0.Y.n119 GNDA 0.388675f
C2377 two_stage_opamp_dummy_magic_29_0.Y.n120 GNDA 0.237753f
C2378 two_stage_opamp_dummy_magic_29_0.Y.n121 GNDA 0.417266f
C2379 two_stage_opamp_dummy_magic_29_0.Y.n122 GNDA 0.237753f
C2380 two_stage_opamp_dummy_magic_29_0.Y.n123 GNDA 0.237753f
C2381 two_stage_opamp_dummy_magic_29_0.Y.n124 GNDA 0.237753f
C2382 two_stage_opamp_dummy_magic_29_0.Y.n125 GNDA 0.341617f
C2383 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n0 GNDA 0.030336f
C2384 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n1 GNDA 0.030623f
C2385 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n4 GNDA 0.030623f
C2386 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n5 GNDA 0.013029f
C2387 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n6 GNDA 0.433353f
C2388 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n7 GNDA 0.013785f
C2389 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n8 GNDA 0.094716f
C2390 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n9 GNDA 0.013029f
C2391 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n10 GNDA 0.088432f
C2392 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n11 GNDA 1.24268f
C2393 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n12 GNDA 2.62402f
C2394 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n14 GNDA 0.030623f
C2395 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n15 GNDA 0.030623f
C2396 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n16 GNDA 0.044021f
C2397 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n17 GNDA 0.044021f
C2398 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n18 GNDA 0.030623f
C2399 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n20 GNDA 0.030623f
C2400 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n21 GNDA 0.030623f
C2401 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n23 GNDA 0.177998f
C2402 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t0 GNDA 0.077525f
C2403 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n24 GNDA 0.029086f
C2404 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n25 GNDA 0.035648f
C2405 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t10 GNDA 0.01276f
C2406 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t15 GNDA 0.01276f
C2407 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n26 GNDA 0.026088f
C2408 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n27 GNDA 0.08763f
C2409 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t11 GNDA 0.01276f
C2410 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t16 GNDA 0.01276f
C2411 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n28 GNDA 0.026088f
C2412 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n29 GNDA 0.084389f
C2413 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n30 GNDA 0.038733f
C2414 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n31 GNDA 0.029086f
C2415 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t13 GNDA 0.01276f
C2416 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t7 GNDA 0.01276f
C2417 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n32 GNDA 0.026088f
C2418 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n33 GNDA 0.084389f
C2419 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n34 GNDA 0.020891f
C2420 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t12 GNDA 0.01276f
C2421 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t9 GNDA 0.01276f
C2422 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n35 GNDA 0.026088f
C2423 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n36 GNDA 0.084389f
C2424 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n37 GNDA 0.035648f
C2425 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t14 GNDA 0.01276f
C2426 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.t8 GNDA 0.01276f
C2427 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n38 GNDA 0.026088f
C2428 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n39 GNDA 0.086056f
C2429 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n40 GNDA 0.116246f
C2430 two_stage_opamp_dummy_magic_29_0.V_CMFB_S1.n41 GNDA 0.610947f
C2431 two_stage_opamp_dummy_magic_29_0.X.n0 GNDA 0.162105f
C2432 two_stage_opamp_dummy_magic_29_0.X.n1 GNDA 0.237753f
C2433 two_stage_opamp_dummy_magic_29_0.X.n2 GNDA 0.417266f
C2434 two_stage_opamp_dummy_magic_29_0.X.n3 GNDA 0.388675f
C2435 two_stage_opamp_dummy_magic_29_0.X.n4 GNDA 0.237753f
C2436 two_stage_opamp_dummy_magic_29_0.X.n5 GNDA 0.237753f
C2437 two_stage_opamp_dummy_magic_29_0.X.n9 GNDA 0.074105f
C2438 two_stage_opamp_dummy_magic_29_0.X.n10 GNDA 0.083312f
C2439 two_stage_opamp_dummy_magic_29_0.X.n11 GNDA 0.083312f
C2440 two_stage_opamp_dummy_magic_29_0.X.t16 GNDA 0.054035f
C2441 two_stage_opamp_dummy_magic_29_0.X.t20 GNDA 0.054035f
C2442 two_stage_opamp_dummy_magic_29_0.X.n12 GNDA 0.110534f
C2443 two_stage_opamp_dummy_magic_29_0.X.n13 GNDA 0.35586f
C2444 two_stage_opamp_dummy_magic_29_0.X.n14 GNDA 0.138043f
C2445 two_stage_opamp_dummy_magic_29_0.X.t18 GNDA 0.054035f
C2446 two_stage_opamp_dummy_magic_29_0.X.t2 GNDA 0.054035f
C2447 two_stage_opamp_dummy_magic_29_0.X.n15 GNDA 0.110534f
C2448 two_stage_opamp_dummy_magic_29_0.X.n16 GNDA 0.348103f
C2449 two_stage_opamp_dummy_magic_29_0.X.n17 GNDA 0.138043f
C2450 two_stage_opamp_dummy_magic_29_0.X.t7 GNDA 0.054035f
C2451 two_stage_opamp_dummy_magic_29_0.X.t19 GNDA 0.054035f
C2452 two_stage_opamp_dummy_magic_29_0.X.n18 GNDA 0.110534f
C2453 two_stage_opamp_dummy_magic_29_0.X.n19 GNDA 0.348103f
C2454 two_stage_opamp_dummy_magic_29_0.X.n20 GNDA 0.083312f
C2455 two_stage_opamp_dummy_magic_29_0.X.n21 GNDA 0.083312f
C2456 two_stage_opamp_dummy_magic_29_0.X.t6 GNDA 0.054035f
C2457 two_stage_opamp_dummy_magic_29_0.X.t1 GNDA 0.054035f
C2458 two_stage_opamp_dummy_magic_29_0.X.n22 GNDA 0.110534f
C2459 two_stage_opamp_dummy_magic_29_0.X.n23 GNDA 0.348103f
C2460 two_stage_opamp_dummy_magic_29_0.X.n24 GNDA 0.083312f
C2461 two_stage_opamp_dummy_magic_29_0.X.t21 GNDA 0.054035f
C2462 two_stage_opamp_dummy_magic_29_0.X.t0 GNDA 0.054035f
C2463 two_stage_opamp_dummy_magic_29_0.X.n25 GNDA 0.110534f
C2464 two_stage_opamp_dummy_magic_29_0.X.n26 GNDA 0.348103f
C2465 two_stage_opamp_dummy_magic_29_0.X.n27 GNDA 0.138043f
C2466 two_stage_opamp_dummy_magic_29_0.X.t8 GNDA 0.054035f
C2467 two_stage_opamp_dummy_magic_29_0.X.t23 GNDA 0.054035f
C2468 two_stage_opamp_dummy_magic_29_0.X.n28 GNDA 0.110534f
C2469 two_stage_opamp_dummy_magic_29_0.X.n29 GNDA 0.351981f
C2470 two_stage_opamp_dummy_magic_29_0.X.n30 GNDA 0.220124f
C2471 two_stage_opamp_dummy_magic_29_0.X.n31 GNDA 0.172911f
C2472 two_stage_opamp_dummy_magic_29_0.X.n33 GNDA 0.074105f
C2473 two_stage_opamp_dummy_magic_29_0.X.n34 GNDA 0.074105f
C2474 two_stage_opamp_dummy_magic_29_0.X.t41 GNDA 0.049789f
C2475 two_stage_opamp_dummy_magic_29_0.X.t26 GNDA 0.056602f
C2476 two_stage_opamp_dummy_magic_29_0.X.n36 GNDA 0.046161f
C2477 two_stage_opamp_dummy_magic_29_0.X.t54 GNDA 0.049789f
C2478 two_stage_opamp_dummy_magic_29_0.X.t39 GNDA 0.049789f
C2479 two_stage_opamp_dummy_magic_29_0.X.t52 GNDA 0.049789f
C2480 two_stage_opamp_dummy_magic_29_0.X.t34 GNDA 0.049789f
C2481 two_stage_opamp_dummy_magic_29_0.X.t47 GNDA 0.049789f
C2482 two_stage_opamp_dummy_magic_29_0.X.t35 GNDA 0.049789f
C2483 two_stage_opamp_dummy_magic_29_0.X.t48 GNDA 0.049789f
C2484 two_stage_opamp_dummy_magic_29_0.X.t31 GNDA 0.056602f
C2485 two_stage_opamp_dummy_magic_29_0.X.n37 GNDA 0.051082f
C2486 two_stage_opamp_dummy_magic_29_0.X.n38 GNDA 0.031263f
C2487 two_stage_opamp_dummy_magic_29_0.X.n39 GNDA 0.031263f
C2488 two_stage_opamp_dummy_magic_29_0.X.n40 GNDA 0.031263f
C2489 two_stage_opamp_dummy_magic_29_0.X.n41 GNDA 0.031263f
C2490 two_stage_opamp_dummy_magic_29_0.X.n42 GNDA 0.031263f
C2491 two_stage_opamp_dummy_magic_29_0.X.n43 GNDA 0.026342f
C2492 two_stage_opamp_dummy_magic_29_0.X.n44 GNDA 0.012791f
C2493 two_stage_opamp_dummy_magic_29_0.X.t42 GNDA 0.032421f
C2494 two_stage_opamp_dummy_magic_29_0.X.t27 GNDA 0.039368f
C2495 two_stage_opamp_dummy_magic_29_0.X.n45 GNDA 0.034447f
C2496 two_stage_opamp_dummy_magic_29_0.X.t25 GNDA 0.032421f
C2497 two_stage_opamp_dummy_magic_29_0.X.t40 GNDA 0.032421f
C2498 two_stage_opamp_dummy_magic_29_0.X.t53 GNDA 0.032421f
C2499 two_stage_opamp_dummy_magic_29_0.X.t37 GNDA 0.032421f
C2500 two_stage_opamp_dummy_magic_29_0.X.t50 GNDA 0.032421f
C2501 two_stage_opamp_dummy_magic_29_0.X.t38 GNDA 0.032421f
C2502 two_stage_opamp_dummy_magic_29_0.X.t51 GNDA 0.032421f
C2503 two_stage_opamp_dummy_magic_29_0.X.t33 GNDA 0.039368f
C2504 two_stage_opamp_dummy_magic_29_0.X.n46 GNDA 0.039368f
C2505 two_stage_opamp_dummy_magic_29_0.X.n47 GNDA 0.025474f
C2506 two_stage_opamp_dummy_magic_29_0.X.n48 GNDA 0.025474f
C2507 two_stage_opamp_dummy_magic_29_0.X.n49 GNDA 0.025474f
C2508 two_stage_opamp_dummy_magic_29_0.X.n50 GNDA 0.025474f
C2509 two_stage_opamp_dummy_magic_29_0.X.n51 GNDA 0.025474f
C2510 two_stage_opamp_dummy_magic_29_0.X.n52 GNDA 0.020552f
C2511 two_stage_opamp_dummy_magic_29_0.X.n53 GNDA 0.012791f
C2512 two_stage_opamp_dummy_magic_29_0.X.n54 GNDA 0.079789f
C2513 two_stage_opamp_dummy_magic_29_0.X.n56 GNDA 0.074105f
C2514 two_stage_opamp_dummy_magic_29_0.X.t24 GNDA 0.640789f
C2515 two_stage_opamp_dummy_magic_29_0.X.n57 GNDA 0.074105f
C2516 two_stage_opamp_dummy_magic_29_0.X.n58 GNDA 0.074105f
C2517 two_stage_opamp_dummy_magic_29_0.X.n59 GNDA 0.073409f
C2518 two_stage_opamp_dummy_magic_29_0.X.n60 GNDA 0.687542f
C2519 two_stage_opamp_dummy_magic_29_0.X.n62 GNDA 0.643787f
C2520 two_stage_opamp_dummy_magic_29_0.X.n63 GNDA 0.024538f
C2521 two_stage_opamp_dummy_magic_29_0.X.n64 GNDA 0.024702f
C2522 two_stage_opamp_dummy_magic_29_0.X.n65 GNDA 0.024702f
C2523 two_stage_opamp_dummy_magic_29_0.X.t30 GNDA 0.101894f
C2524 two_stage_opamp_dummy_magic_29_0.X.t46 GNDA 0.101894f
C2525 two_stage_opamp_dummy_magic_29_0.X.t32 GNDA 0.101894f
C2526 two_stage_opamp_dummy_magic_29_0.X.t49 GNDA 0.101894f
C2527 two_stage_opamp_dummy_magic_29_0.X.t36 GNDA 0.108524f
C2528 two_stage_opamp_dummy_magic_29_0.X.n66 GNDA 0.086001f
C2529 two_stage_opamp_dummy_magic_29_0.X.n67 GNDA 0.048631f
C2530 two_stage_opamp_dummy_magic_29_0.X.n68 GNDA 0.048631f
C2531 two_stage_opamp_dummy_magic_29_0.X.n69 GNDA 0.04371f
C2532 two_stage_opamp_dummy_magic_29_0.X.t44 GNDA 0.101894f
C2533 two_stage_opamp_dummy_magic_29_0.X.t28 GNDA 0.101894f
C2534 two_stage_opamp_dummy_magic_29_0.X.t45 GNDA 0.101894f
C2535 two_stage_opamp_dummy_magic_29_0.X.t29 GNDA 0.101894f
C2536 two_stage_opamp_dummy_magic_29_0.X.t43 GNDA 0.108524f
C2537 two_stage_opamp_dummy_magic_29_0.X.n70 GNDA 0.086001f
C2538 two_stage_opamp_dummy_magic_29_0.X.n71 GNDA 0.048631f
C2539 two_stage_opamp_dummy_magic_29_0.X.n72 GNDA 0.048631f
C2540 two_stage_opamp_dummy_magic_29_0.X.n73 GNDA 0.04371f
C2541 two_stage_opamp_dummy_magic_29_0.X.n74 GNDA 0.010496f
C2542 two_stage_opamp_dummy_magic_29_0.X.n75 GNDA 0.024866f
C2543 two_stage_opamp_dummy_magic_29_0.X.n76 GNDA 0.058532f
C2544 two_stage_opamp_dummy_magic_29_0.X.n77 GNDA 0.033384f
C2545 two_stage_opamp_dummy_magic_29_0.X.n78 GNDA 0.037886f
C2546 two_stage_opamp_dummy_magic_29_0.X.n79 GNDA 1.02357f
C2547 two_stage_opamp_dummy_magic_29_0.X.n80 GNDA 0.453893f
C2548 two_stage_opamp_dummy_magic_29_0.X.n81 GNDA 2.18995f
C2549 two_stage_opamp_dummy_magic_29_0.X.n82 GNDA 0.074105f
C2550 two_stage_opamp_dummy_magic_29_0.X.n84 GNDA 0.463156f
C2551 two_stage_opamp_dummy_magic_29_0.X.n85 GNDA 0.463156f
C2552 two_stage_opamp_dummy_magic_29_0.X.n86 GNDA 0.074105f
C2553 two_stage_opamp_dummy_magic_29_0.X.n88 GNDA 0.074105f
C2554 two_stage_opamp_dummy_magic_29_0.X.n90 GNDA 0.074105f
C2555 two_stage_opamp_dummy_magic_29_0.X.n92 GNDA 0.074105f
C2556 two_stage_opamp_dummy_magic_29_0.X.n93 GNDA 0.172911f
C2557 two_stage_opamp_dummy_magic_29_0.X.n95 GNDA 0.619675f
C2558 two_stage_opamp_dummy_magic_29_0.X.n97 GNDA 1.3941f
C2559 two_stage_opamp_dummy_magic_29_0.X.n98 GNDA 1.42652f
C2560 two_stage_opamp_dummy_magic_29_0.X.n99 GNDA 0.237753f
C2561 two_stage_opamp_dummy_magic_29_0.X.n100 GNDA 0.237753f
C2562 two_stage_opamp_dummy_magic_29_0.X.n101 GNDA 0.237753f
C2563 two_stage_opamp_dummy_magic_29_0.X.n102 GNDA 0.417266f
C2564 two_stage_opamp_dummy_magic_29_0.X.n103 GNDA 0.146616f
C2565 two_stage_opamp_dummy_magic_29_0.X.n104 GNDA 0.08603f
C2566 two_stage_opamp_dummy_magic_29_0.X.n105 GNDA 0.08603f
C2567 two_stage_opamp_dummy_magic_29_0.X.n106 GNDA 0.496725f
C2568 two_stage_opamp_dummy_magic_29_0.X.n107 GNDA 0.08603f
C2569 two_stage_opamp_dummy_magic_29_0.X.t12 GNDA 0.023158f
C2570 two_stage_opamp_dummy_magic_29_0.X.t22 GNDA 0.023158f
C2571 two_stage_opamp_dummy_magic_29_0.X.n108 GNDA 0.068053f
C2572 two_stage_opamp_dummy_magic_29_0.X.t13 GNDA 0.023158f
C2573 two_stage_opamp_dummy_magic_29_0.X.t10 GNDA 0.023158f
C2574 two_stage_opamp_dummy_magic_29_0.X.n109 GNDA 0.066733f
C2575 two_stage_opamp_dummy_magic_29_0.X.n110 GNDA 0.44107f
C2576 two_stage_opamp_dummy_magic_29_0.X.t15 GNDA 0.023158f
C2577 two_stage_opamp_dummy_magic_29_0.X.t9 GNDA 0.023158f
C2578 two_stage_opamp_dummy_magic_29_0.X.n111 GNDA 0.066733f
C2579 two_stage_opamp_dummy_magic_29_0.X.n112 GNDA 0.232002f
C2580 two_stage_opamp_dummy_magic_29_0.X.t11 GNDA 0.023158f
C2581 two_stage_opamp_dummy_magic_29_0.X.t4 GNDA 0.023158f
C2582 two_stage_opamp_dummy_magic_29_0.X.n113 GNDA 0.066733f
C2583 two_stage_opamp_dummy_magic_29_0.X.n114 GNDA 0.232002f
C2584 two_stage_opamp_dummy_magic_29_0.X.t5 GNDA 0.023158f
C2585 two_stage_opamp_dummy_magic_29_0.X.t3 GNDA 0.023158f
C2586 two_stage_opamp_dummy_magic_29_0.X.n115 GNDA 0.066733f
C2587 two_stage_opamp_dummy_magic_29_0.X.n116 GNDA 0.232002f
C2588 two_stage_opamp_dummy_magic_29_0.X.t14 GNDA 0.023158f
C2589 two_stage_opamp_dummy_magic_29_0.X.t17 GNDA 0.023158f
C2590 two_stage_opamp_dummy_magic_29_0.X.n117 GNDA 0.066733f
C2591 two_stage_opamp_dummy_magic_29_0.X.n118 GNDA 0.431159f
C2592 two_stage_opamp_dummy_magic_29_0.X.n119 GNDA 0.287483f
C2593 two_stage_opamp_dummy_magic_29_0.X.n120 GNDA 0.644415f
C2594 two_stage_opamp_dummy_magic_29_0.X.n121 GNDA 0.815021f
C2595 two_stage_opamp_dummy_magic_29_0.X.n122 GNDA 0.237753f
C2596 two_stage_opamp_dummy_magic_29_0.X.n123 GNDA 0.417266f
C2597 two_stage_opamp_dummy_magic_29_0.X.n124 GNDA 0.237753f
C2598 two_stage_opamp_dummy_magic_29_0.X.n125 GNDA 0.194525f
C2599 two_stage_opamp_dummy_magic_29_0.VD4.n0 GNDA 2.28471f
C2600 two_stage_opamp_dummy_magic_29_0.VD4.n1 GNDA 1.10445f
C2601 two_stage_opamp_dummy_magic_29_0.VD4.n2 GNDA 0.830716f
C2602 two_stage_opamp_dummy_magic_29_0.VD4.n3 GNDA 1.30021f
C2603 two_stage_opamp_dummy_magic_29_0.VD4.t3 GNDA 0.045031f
C2604 two_stage_opamp_dummy_magic_29_0.VD4.t13 GNDA 0.045031f
C2605 two_stage_opamp_dummy_magic_29_0.VD4.n4 GNDA 0.095624f
C2606 two_stage_opamp_dummy_magic_29_0.VD4.t27 GNDA 0.045031f
C2607 two_stage_opamp_dummy_magic_29_0.VD4.t30 GNDA 0.045031f
C2608 two_stage_opamp_dummy_magic_29_0.VD4.n5 GNDA 0.092115f
C2609 two_stage_opamp_dummy_magic_29_0.VD4.n6 GNDA 0.25692f
C2610 two_stage_opamp_dummy_magic_29_0.VD4.t9 GNDA 0.045031f
C2611 two_stage_opamp_dummy_magic_29_0.VD4.t1 GNDA 0.045031f
C2612 two_stage_opamp_dummy_magic_29_0.VD4.n7 GNDA 0.095624f
C2613 two_stage_opamp_dummy_magic_29_0.VD4.t25 GNDA 0.045031f
C2614 two_stage_opamp_dummy_magic_29_0.VD4.t23 GNDA 0.045031f
C2615 two_stage_opamp_dummy_magic_29_0.VD4.n8 GNDA 0.092115f
C2616 two_stage_opamp_dummy_magic_29_0.VD4.n9 GNDA 0.25692f
C2617 two_stage_opamp_dummy_magic_29_0.VD4.t5 GNDA 0.045031f
C2618 two_stage_opamp_dummy_magic_29_0.VD4.t11 GNDA 0.045031f
C2619 two_stage_opamp_dummy_magic_29_0.VD4.n10 GNDA 0.095624f
C2620 two_stage_opamp_dummy_magic_29_0.VD4.t15 GNDA 0.045031f
C2621 two_stage_opamp_dummy_magic_29_0.VD4.t17 GNDA 0.045031f
C2622 two_stage_opamp_dummy_magic_29_0.VD4.n11 GNDA 0.095624f
C2623 two_stage_opamp_dummy_magic_29_0.VD4.t20 GNDA 0.045031f
C2624 two_stage_opamp_dummy_magic_29_0.VD4.t22 GNDA 0.045031f
C2625 two_stage_opamp_dummy_magic_29_0.VD4.n12 GNDA 0.092115f
C2626 two_stage_opamp_dummy_magic_29_0.VD4.n13 GNDA 0.260153f
C2627 two_stage_opamp_dummy_magic_29_0.VD4.n14 GNDA 0.115041f
C2628 two_stage_opamp_dummy_magic_29_0.VD4.n15 GNDA 0.069429f
C2629 two_stage_opamp_dummy_magic_29_0.VD4.t7 GNDA 0.045031f
C2630 two_stage_opamp_dummy_magic_29_0.VD4.t19 GNDA 0.045031f
C2631 two_stage_opamp_dummy_magic_29_0.VD4.n16 GNDA 0.095624f
C2632 two_stage_opamp_dummy_magic_29_0.VD4.t34 GNDA 0.160181f
C2633 two_stage_opamp_dummy_magic_29_0.VD4.t35 GNDA 0.078836f
C2634 two_stage_opamp_dummy_magic_29_0.VD4.n17 GNDA 0.149757f
C2635 two_stage_opamp_dummy_magic_29_0.VD4.t37 GNDA 0.160181f
C2636 two_stage_opamp_dummy_magic_29_0.VD4.n18 GNDA 0.51334f
C2637 two_stage_opamp_dummy_magic_29_0.VD4.t36 GNDA 0.383839f
C2638 two_stage_opamp_dummy_magic_29_0.VD4.t2 GNDA 0.301063f
C2639 two_stage_opamp_dummy_magic_29_0.VD4.t12 GNDA 0.301063f
C2640 two_stage_opamp_dummy_magic_29_0.VD4.t8 GNDA 0.301063f
C2641 two_stage_opamp_dummy_magic_29_0.VD4.t0 GNDA 0.301063f
C2642 two_stage_opamp_dummy_magic_29_0.VD4.t4 GNDA 0.301063f
C2643 two_stage_opamp_dummy_magic_29_0.VD4.t10 GNDA 0.301063f
C2644 two_stage_opamp_dummy_magic_29_0.VD4.t14 GNDA 0.301063f
C2645 two_stage_opamp_dummy_magic_29_0.VD4.t16 GNDA 0.301063f
C2646 two_stage_opamp_dummy_magic_29_0.VD4.t6 GNDA 0.301063f
C2647 two_stage_opamp_dummy_magic_29_0.VD4.t18 GNDA 0.301063f
C2648 two_stage_opamp_dummy_magic_29_0.VD4.t33 GNDA 0.383839f
C2649 two_stage_opamp_dummy_magic_29_0.VD4.n19 GNDA 0.51334f
C2650 two_stage_opamp_dummy_magic_29_0.VD4.t32 GNDA 0.078836f
C2651 two_stage_opamp_dummy_magic_29_0.VD4.n20 GNDA 0.216535f
C2652 two_stage_opamp_dummy_magic_29_0.VD4.t26 GNDA 0.045031f
C2653 two_stage_opamp_dummy_magic_29_0.VD4.t21 GNDA 0.045031f
C2654 two_stage_opamp_dummy_magic_29_0.VD4.n21 GNDA 0.092115f
C2655 two_stage_opamp_dummy_magic_29_0.VD4.n22 GNDA 0.260153f
C2656 two_stage_opamp_dummy_magic_29_0.VD4.t24 GNDA 0.045031f
C2657 two_stage_opamp_dummy_magic_29_0.VD4.t29 GNDA 0.045031f
C2658 two_stage_opamp_dummy_magic_29_0.VD4.n23 GNDA 0.092115f
C2659 two_stage_opamp_dummy_magic_29_0.VD4.n24 GNDA 0.25692f
C2660 two_stage_opamp_dummy_magic_29_0.VD4.n25 GNDA 0.115041f
C2661 two_stage_opamp_dummy_magic_29_0.VD4.n26 GNDA 0.069429f
C2662 two_stage_opamp_dummy_magic_29_0.VD4.t28 GNDA 0.045031f
C2663 two_stage_opamp_dummy_magic_29_0.VD4.t31 GNDA 0.045031f
C2664 two_stage_opamp_dummy_magic_29_0.VD4.n27 GNDA 0.092115f
C2665 two_stage_opamp_dummy_magic_29_0.VD4.n28 GNDA 0.25692f
C2666 two_stage_opamp_dummy_magic_29_0.Vb3.n0 GNDA 0.409529f
C2667 two_stage_opamp_dummy_magic_29_0.Vb3.n1 GNDA 0.067898f
C2668 two_stage_opamp_dummy_magic_29_0.Vb3.n2 GNDA 0.158927f
C2669 two_stage_opamp_dummy_magic_29_0.Vb3.n3 GNDA 0.20902f
C2670 two_stage_opamp_dummy_magic_29_0.Vb3.n4 GNDA 0.483439f
C2671 two_stage_opamp_dummy_magic_29_0.Vb3.n5 GNDA 0.138459f
C2672 two_stage_opamp_dummy_magic_29_0.Vb3.n6 GNDA 0.20902f
C2673 two_stage_opamp_dummy_magic_29_0.Vb3.n7 GNDA 0.138459f
C2674 two_stage_opamp_dummy_magic_29_0.Vb3.n8 GNDA 0.305019f
C2675 two_stage_opamp_dummy_magic_29_0.Vb3.t2 GNDA 0.014145f
C2676 two_stage_opamp_dummy_magic_29_0.Vb3.t4 GNDA 0.014145f
C2677 two_stage_opamp_dummy_magic_29_0.Vb3.n9 GNDA 0.045564f
C2678 two_stage_opamp_dummy_magic_29_0.Vb3.t3 GNDA 0.014145f
C2679 two_stage_opamp_dummy_magic_29_0.Vb3.t1 GNDA 0.014145f
C2680 two_stage_opamp_dummy_magic_29_0.Vb3.n10 GNDA 0.045564f
C2681 two_stage_opamp_dummy_magic_29_0.Vb3.n11 GNDA 0.25119f
C2682 two_stage_opamp_dummy_magic_29_0.Vb3.t6 GNDA 0.014145f
C2683 two_stage_opamp_dummy_magic_29_0.Vb3.t5 GNDA 0.014145f
C2684 two_stage_opamp_dummy_magic_29_0.Vb3.n12 GNDA 0.042725f
C2685 two_stage_opamp_dummy_magic_29_0.Vb3.n13 GNDA 0.801828f
C2686 two_stage_opamp_dummy_magic_29_0.Vb3.t23 GNDA 0.090719f
C2687 two_stage_opamp_dummy_magic_29_0.Vb3.t13 GNDA 0.090696f
C2688 two_stage_opamp_dummy_magic_29_0.Vb3.t28 GNDA 0.090696f
C2689 two_stage_opamp_dummy_magic_29_0.Vb3.t12 GNDA 0.090696f
C2690 two_stage_opamp_dummy_magic_29_0.Vb3.t27 GNDA 0.090281f
C2691 two_stage_opamp_dummy_magic_29_0.Vb3.t17 GNDA 0.090281f
C2692 two_stage_opamp_dummy_magic_29_0.Vb3.t10 GNDA 0.090696f
C2693 two_stage_opamp_dummy_magic_29_0.Vb3.t21 GNDA 0.090696f
C2694 two_stage_opamp_dummy_magic_29_0.Vb3.t26 GNDA 0.090696f
C2695 two_stage_opamp_dummy_magic_29_0.Vb3.t16 GNDA 0.090696f
C2696 two_stage_opamp_dummy_magic_29_0.Vb3.t7 GNDA 0.049509f
C2697 two_stage_opamp_dummy_magic_29_0.Vb3.t0 GNDA 0.049509f
C2698 two_stage_opamp_dummy_magic_29_0.Vb3.n14 GNDA 0.133295f
C2699 two_stage_opamp_dummy_magic_29_0.Vb3.t19 GNDA 0.092967f
C2700 two_stage_opamp_dummy_magic_29_0.Vb3.n15 GNDA 0.93118f
C2701 two_stage_opamp_dummy_magic_29_0.Vb3.n16 GNDA 1.05807f
C2702 two_stage_opamp_dummy_magic_29_0.Vb3.t18 GNDA 0.090719f
C2703 two_stage_opamp_dummy_magic_29_0.Vb3.t11 GNDA 0.090696f
C2704 two_stage_opamp_dummy_magic_29_0.Vb3.t22 GNDA 0.090696f
C2705 two_stage_opamp_dummy_magic_29_0.Vb3.t8 GNDA 0.090696f
C2706 two_stage_opamp_dummy_magic_29_0.Vb3.t24 GNDA 0.090271f
C2707 two_stage_opamp_dummy_magic_29_0.Vb3.t14 GNDA 0.090271f
C2708 two_stage_opamp_dummy_magic_29_0.Vb3.n17 GNDA 0.079473f
C2709 two_stage_opamp_dummy_magic_29_0.Vb3.n18 GNDA 0.079473f
C2710 two_stage_opamp_dummy_magic_29_0.Vb3.t20 GNDA 0.090696f
C2711 two_stage_opamp_dummy_magic_29_0.Vb3.t9 GNDA 0.090696f
C2712 two_stage_opamp_dummy_magic_29_0.Vb3.t15 GNDA 0.090696f
C2713 two_stage_opamp_dummy_magic_29_0.Vb3.t25 GNDA 0.090696f
C2714 two_stage_opamp_dummy_magic_29_0.Vb3.n19 GNDA 0.145531f
C2715 two_stage_opamp_dummy_magic_29_0.Vb3.n20 GNDA 1.07033f
C2716 bgr_11_0.VB3_CUR_BIAS GNDA 1.50687f
C2717 VDDA.n16 GNDA 0.112326f
C2718 VDDA.n17 GNDA 0.137288f
C2719 VDDA.n18 GNDA 0.112326f
C2720 VDDA.n32 GNDA 0.013087f
C2721 VDDA.n34 GNDA 0.013571f
C2722 VDDA.n36 GNDA 0.012117f
C2723 VDDA.n38 GNDA 0.013087f
C2724 VDDA.n40 GNDA 0.013571f
C2725 VDDA.t159 GNDA 0.090313f
C2726 VDDA.t415 GNDA 0.090641f
C2727 VDDA.t83 GNDA 0.085794f
C2728 VDDA.t128 GNDA 0.090313f
C2729 VDDA.t387 GNDA 0.090641f
C2730 VDDA.t44 GNDA 0.085794f
C2731 VDDA.t418 GNDA 0.090313f
C2732 VDDA.t152 GNDA 0.090641f
C2733 VDDA.t142 GNDA 0.085794f
C2734 VDDA.t43 GNDA 0.090313f
C2735 VDDA.t82 GNDA 0.090641f
C2736 VDDA.t14 GNDA 0.085794f
C2737 VDDA.t369 GNDA 0.090313f
C2738 VDDA.t129 GNDA 0.090641f
C2739 VDDA.t127 GNDA 0.085794f
C2740 VDDA.n42 GNDA 0.060537f
C2741 VDDA.t15 GNDA 0.048209f
C2742 VDDA.n43 GNDA 0.065684f
C2743 VDDA.t153 GNDA 0.048209f
C2744 VDDA.n44 GNDA 0.065684f
C2745 VDDA.t388 GNDA 0.048209f
C2746 VDDA.n45 GNDA 0.065684f
C2747 VDDA.t72 GNDA 0.048209f
C2748 VDDA.n46 GNDA 0.065684f
C2749 VDDA.t141 GNDA 0.258312f
C2750 VDDA.n48 GNDA 1.09384f
C2751 VDDA.n49 GNDA 0.013087f
C2752 VDDA.n50 GNDA 0.013571f
C2753 VDDA.n58 GNDA 0.013087f
C2754 VDDA.n59 GNDA 0.012117f
C2755 VDDA.n60 GNDA 0.012117f
C2756 VDDA.n68 GNDA 0.013571f
C2757 VDDA.n69 GNDA 0.013571f
C2758 VDDA.n70 GNDA 0.013087f
C2759 VDDA.n78 GNDA 0.012117f
C2760 VDDA.n79 GNDA 0.013087f
C2761 VDDA.n80 GNDA 0.013571f
C2762 VDDA.n88 GNDA 0.013087f
C2763 VDDA.n89 GNDA 0.012117f
C2764 VDDA.n90 GNDA 0.012117f
C2765 VDDA.n98 GNDA 0.040569f
C2766 VDDA.n101 GNDA 2.31517f
C2767 VDDA.n115 GNDA 0.013087f
C2768 VDDA.n119 GNDA 0.013571f
C2769 VDDA.n123 GNDA 0.012117f
C2770 VDDA.n127 GNDA 0.013087f
C2771 VDDA.n131 GNDA 0.013571f
C2772 VDDA.n136 GNDA 0.037804f
C2773 VDDA.n142 GNDA 0.013087f
C2774 VDDA.n143 GNDA 0.012117f
C2775 VDDA.n144 GNDA 0.012117f
C2776 VDDA.n150 GNDA 0.013571f
C2777 VDDA.n151 GNDA 0.013571f
C2778 VDDA.n152 GNDA 0.013087f
C2779 VDDA.n158 GNDA 0.012117f
C2780 VDDA.n159 GNDA 0.013087f
C2781 VDDA.n160 GNDA 0.013571f
C2782 VDDA.n166 GNDA 0.013087f
C2783 VDDA.n167 GNDA 0.012117f
C2784 VDDA.n168 GNDA 0.012117f
C2785 VDDA.n174 GNDA 0.013571f
C2786 VDDA.n175 GNDA 0.013571f
C2787 VDDA.n180 GNDA 0.025026f
C2788 VDDA.n181 GNDA 0.085483f
C2789 VDDA.t276 GNDA 0.034115f
C2790 VDDA.n186 GNDA 0.014673f
C2791 VDDA.n187 GNDA 0.047529f
C2792 VDDA.t338 GNDA 0.01447f
C2793 VDDA.t326 GNDA 0.028698f
C2794 VDDA.n192 GNDA 0.014205f
C2795 VDDA.n193 GNDA 0.041373f
C2796 VDDA.t321 GNDA 0.020115f
C2797 VDDA.t319 GNDA 0.010014f
C2798 VDDA.n194 GNDA 0.014205f
C2799 VDDA.n195 GNDA 0.041373f
C2800 VDDA.n196 GNDA 0.014205f
C2801 VDDA.n197 GNDA 0.041373f
C2802 VDDA.n198 GNDA 0.014205f
C2803 VDDA.n199 GNDA 0.041373f
C2804 VDDA.n200 GNDA 0.014205f
C2805 VDDA.n201 GNDA 0.046145f
C2806 VDDA.n202 GNDA 0.021395f
C2807 VDDA.n203 GNDA 0.064337f
C2808 VDDA.t320 GNDA 0.0482f
C2809 VDDA.t378 GNDA 0.037806f
C2810 VDDA.t60 GNDA 0.037806f
C2811 VDDA.t29 GNDA 0.037806f
C2812 VDDA.t1 GNDA 0.037806f
C2813 VDDA.t196 GNDA 0.037806f
C2814 VDDA.t374 GNDA 0.037806f
C2815 VDDA.t89 GNDA 0.037806f
C2816 VDDA.t25 GNDA 0.037806f
C2817 VDDA.t376 GNDA 0.037806f
C2818 VDDA.t93 GNDA 0.037806f
C2819 VDDA.t358 GNDA 0.0482f
C2820 VDDA.t359 GNDA 0.020115f
C2821 VDDA.n204 GNDA 0.064337f
C2822 VDDA.t357 GNDA 0.010014f
C2823 VDDA.n205 GNDA 0.020998f
C2824 VDDA.n206 GNDA 0.022545f
C2825 VDDA.n218 GNDA 0.013673f
C2826 VDDA.n219 GNDA 0.013462f
C2827 VDDA.n220 GNDA 0.105669f
C2828 VDDA.n221 GNDA 0.013462f
C2829 VDDA.n222 GNDA 0.056333f
C2830 VDDA.n223 GNDA 0.013462f
C2831 VDDA.n224 GNDA 0.056333f
C2832 VDDA.n225 GNDA 0.013462f
C2833 VDDA.n226 GNDA 0.056333f
C2834 VDDA.n227 GNDA 0.013462f
C2835 VDDA.n228 GNDA 0.07572f
C2836 VDDA.n229 GNDA 0.033928f
C2837 VDDA.n233 GNDA 0.103238f
C2838 VDDA.n234 GNDA 0.041982f
C2839 VDDA.t285 GNDA 0.011528f
C2840 VDDA.n235 GNDA 0.035415f
C2841 VDDA.t284 GNDA 0.02872f
C2842 VDDA.t156 GNDA 0.021326f
C2843 VDDA.t187 GNDA 0.021326f
C2844 VDDA.t45 GNDA 0.021326f
C2845 VDDA.t123 GNDA 0.021326f
C2846 VDDA.t37 GNDA 0.021326f
C2847 VDDA.t134 GNDA 0.021326f
C2848 VDDA.t186 GNDA 0.021326f
C2849 VDDA.t106 GNDA 0.021326f
C2850 VDDA.t76 GNDA 0.021326f
C2851 VDDA.t103 GNDA 0.021326f
C2852 VDDA.t290 GNDA 0.02872f
C2853 VDDA.t291 GNDA 0.011528f
C2854 VDDA.n236 GNDA 0.035415f
C2855 VDDA.n237 GNDA 0.025384f
C2856 VDDA.n238 GNDA 0.14734f
C2857 VDDA.n239 GNDA 0.028596f
C2858 VDDA.n241 GNDA 0.103238f
C2859 VDDA.n244 GNDA 0.110509f
C2860 VDDA.n245 GNDA 0.025026f
C2861 VDDA.n246 GNDA 0.085483f
C2862 VDDA.t366 GNDA 0.034115f
C2863 VDDA.n249 GNDA 0.013571f
C2864 VDDA.n276 GNDA 0.063748f
C2865 VDDA.n280 GNDA 0.010116f
C2866 VDDA.n281 GNDA 0.01161f
C2867 VDDA.n282 GNDA 0.010116f
C2868 VDDA.n285 GNDA 0.014085f
C2869 VDDA.n291 GNDA 0.010434f
C2870 VDDA.n294 GNDA 0.046165f
C2871 VDDA.t296 GNDA 0.067887f
C2872 VDDA.n295 GNDA 0.019771f
C2873 VDDA.t216 GNDA 0.02067f
C2874 VDDA.t333 GNDA 0.069976f
C2875 VDDA.n296 GNDA 0.048736f
C2876 VDDA.n299 GNDA 0.010434f
C2877 VDDA.n306 GNDA 0.025239f
C2878 VDDA.n308 GNDA 0.02916f
C2879 VDDA.n358 GNDA 0.019772f
C2880 VDDA.n361 GNDA 5.56015f
C2881 VDDA.n372 GNDA 0.01148f
C2882 VDDA.n375 GNDA 0.013087f
C2883 VDDA.n377 GNDA 0.013571f
C2884 VDDA.n379 GNDA 0.012117f
C2885 VDDA.n381 GNDA 0.013087f
C2886 VDDA.n383 GNDA 0.013571f
C2887 VDDA.n384 GNDA 0.012418f
C2888 VDDA.t421 GNDA 0.190858f
C2889 VDDA.t423 GNDA 0.190858f
C2890 VDDA.t424 GNDA 0.181324f
C2891 VDDA.n393 GNDA 0.350946f
C2892 VDDA.n394 GNDA 0.185299f
C2893 VDDA.t422 GNDA 0.179114f
C2894 VDDA.n395 GNDA 0.240449f
C2895 VDDA.n396 GNDA 0.127152f
C2896 VDDA.n401 GNDA 0.091606f
C2897 VDDA.n402 GNDA 0.091606f
C2898 VDDA.n404 GNDA 0.04319f
C2899 VDDA.n408 GNDA 0.04319f
C2900 VDDA.n410 GNDA 0.04319f
C2901 VDDA.n412 GNDA 0.04319f
C2902 VDDA.n414 GNDA 0.04319f
C2903 VDDA.n416 GNDA 0.04319f
C2904 VDDA.n418 GNDA 0.04319f
C2905 VDDA.n420 GNDA 0.04319f
C2906 VDDA.n422 GNDA 0.04319f
C2907 VDDA.n424 GNDA 0.04319f
C2908 VDDA.n428 GNDA 0.04319f
C2909 VDDA.n430 GNDA 0.04319f
C2910 VDDA.n432 GNDA 0.04319f
C2911 VDDA.n434 GNDA 0.04319f
C2912 VDDA.n436 GNDA 0.04319f
C2913 VDDA.n438 GNDA 0.04319f
C2914 VDDA.n440 GNDA 0.04319f
C2915 VDDA.n442 GNDA 0.058853f
C2916 VDDA.n443 GNDA 0.018888f
C2917 VDDA.n446 GNDA 0.019915f
C2918 VDDA.t257 GNDA 0.016767f
C2919 VDDA.t204 GNDA 0.013571f
C2920 VDDA.t157 GNDA 0.013571f
C2921 VDDA.t389 GNDA 0.013571f
C2922 VDDA.t405 GNDA 0.013571f
C2923 VDDA.t382 GNDA 0.013571f
C2924 VDDA.t200 GNDA 0.013571f
C2925 VDDA.t208 GNDA 0.013571f
C2926 VDDA.t77 GNDA 0.013571f
C2927 VDDA.t178 GNDA 0.013571f
C2928 VDDA.t56 GNDA 0.013571f
C2929 VDDA.t192 GNDA 0.013571f
C2930 VDDA.t202 GNDA 0.013571f
C2931 VDDA.t210 GNDA 0.013571f
C2932 VDDA.t12 GNDA 0.013571f
C2933 VDDA.t170 GNDA 0.013571f
C2934 VDDA.t20 GNDA 0.013571f
C2935 VDDA.t99 GNDA 0.013571f
C2936 VDDA.t206 GNDA 0.013571f
C2937 VDDA.t278 GNDA 0.020622f
C2938 VDDA.n447 GNDA 0.017191f
C2939 VDDA.n450 GNDA 0.013339f
C2940 VDDA.n451 GNDA 0.043906f
C2941 VDDA.n452 GNDA 0.043906f
C2942 VDDA.n453 GNDA 0.017787f
C2943 VDDA.n456 GNDA 0.020909f
C2944 VDDA.t266 GNDA 0.016904f
C2945 VDDA.t176 GNDA 0.013571f
C2946 VDDA.t67 GNDA 0.013571f
C2947 VDDA.t49 GNDA 0.013571f
C2948 VDDA.t10 GNDA 0.013571f
C2949 VDDA.t395 GNDA 0.013571f
C2950 VDDA.t190 GNDA 0.013571f
C2951 VDDA.t136 GNDA 0.013571f
C2952 VDDA.t413 GNDA 0.013571f
C2953 VDDA.t79 GNDA 0.013571f
C2954 VDDA.t18 GNDA 0.013571f
C2955 VDDA.t180 GNDA 0.013571f
C2956 VDDA.t47 GNDA 0.013571f
C2957 VDDA.t40 GNDA 0.013571f
C2958 VDDA.t163 GNDA 0.013571f
C2959 VDDA.t172 GNDA 0.013571f
C2960 VDDA.t165 GNDA 0.013571f
C2961 VDDA.t384 GNDA 0.013571f
C2962 VDDA.t150 GNDA 0.013571f
C2963 VDDA.t323 GNDA 0.020307f
C2964 VDDA.n457 GNDA 0.016375f
C2965 VDDA.n460 GNDA 0.013339f
C2966 VDDA.n461 GNDA 0.093344f
C2967 VDDA.n462 GNDA 0.084336f
C2968 VDDA.n467 GNDA 0.066402f
C2969 VDDA.n468 GNDA 0.066402f
C2970 VDDA.t268 GNDA 0.023112f
C2971 VDDA.n470 GNDA 0.018859f
C2972 VDDA.n471 GNDA 0.018859f
C2973 VDDA.n472 GNDA 0.018859f
C2974 VDDA.n473 GNDA 0.018859f
C2975 VDDA.n474 GNDA 0.018859f
C2976 VDDA.n475 GNDA 0.018859f
C2977 VDDA.n476 GNDA 0.018859f
C2978 VDDA.n477 GNDA 0.018859f
C2979 VDDA.n503 GNDA 0.045318f
C2980 VDDA.t269 GNDA 0.048065f
C2981 VDDA.t33 GNDA 0.049438f
C2982 VDDA.t119 GNDA 0.049438f
C2983 VDDA.t419 GNDA 0.049438f
C2984 VDDA.t397 GNDA 0.049438f
C2985 VDDA.t121 GNDA 0.049438f
C2986 VDDA.t403 GNDA 0.049438f
C2987 VDDA.t416 GNDA 0.049438f
C2988 VDDA.t139 GNDA 0.049438f
C2989 VDDA.t143 GNDA 0.049438f
C2990 VDDA.t31 GNDA 0.049438f
C2991 VDDA.t370 GNDA 0.049438f
C2992 VDDA.t401 GNDA 0.049438f
C2993 VDDA.t399 GNDA 0.049438f
C2994 VDDA.t70 GNDA 0.049438f
C2995 VDDA.t130 GNDA 0.049438f
C2996 VDDA.t160 GNDA 0.049438f
C2997 VDDA.t346 GNDA 0.048065f
C2998 VDDA.n520 GNDA 0.045318f
C2999 VDDA.t345 GNDA 0.023112f
C3000 VDDA.n524 GNDA 0.092366f
C3001 VDDA.n525 GNDA 0.06483f
C3002 VDDA.n526 GNDA 0.06483f
C3003 VDDA.n527 GNDA 0.06483f
C3004 VDDA.n528 GNDA 0.06483f
C3005 VDDA.n529 GNDA 0.06483f
C3006 VDDA.n530 GNDA 0.06483f
C3007 VDDA.n531 GNDA 0.06483f
C3008 VDDA.n532 GNDA 0.054668f
C3009 VDDA.n533 GNDA 0.062336f
C3010 VDDA.n535 GNDA 0.02965f
C3011 VDDA.t343 GNDA 0.020036f
C3012 VDDA.t162 GNDA 0.01244f
C3013 VDDA.t169 GNDA 0.01244f
C3014 VDDA.t299 GNDA 0.019604f
C3015 VDDA.n536 GNDA 0.02831f
C3016 VDDA.n538 GNDA 0.113712f
C3017 VDDA.n539 GNDA 0.08579f
C3018 VDDA.n544 GNDA 0.03102f
C3019 VDDA.n545 GNDA 0.03102f
C3020 VDDA.n548 GNDA 0.028154f
C3021 VDDA.t314 GNDA 0.019603f
C3022 VDDA.t228 GNDA 0.01244f
C3023 VDDA.t212 GNDA 0.01244f
C3024 VDDA.t251 GNDA 0.019603f
C3025 VDDA.n549 GNDA 0.028154f
C3026 VDDA.n551 GNDA 0.017139f
C3027 VDDA.n552 GNDA 0.017282f
C3028 VDDA.t272 GNDA 0.017824f
C3029 VDDA.t220 GNDA 0.01244f
C3030 VDDA.t242 GNDA 0.01244f
C3031 VDDA.t234 GNDA 0.01244f
C3032 VDDA.t218 GNDA 0.01244f
C3033 VDDA.t349 GNDA 0.017824f
C3034 VDDA.n553 GNDA 0.017282f
C3035 VDDA.n554 GNDA 0.017139f
C3036 VDDA.n561 GNDA 0.028154f
C3037 VDDA.t305 GNDA 0.019603f
C3038 VDDA.t224 GNDA 0.01244f
C3039 VDDA.t244 GNDA 0.01244f
C3040 VDDA.t236 GNDA 0.01244f
C3041 VDDA.t222 GNDA 0.01244f
C3042 VDDA.t240 GNDA 0.01244f
C3043 VDDA.t230 GNDA 0.01244f
C3044 VDDA.t232 GNDA 0.01244f
C3045 VDDA.t214 GNDA 0.01244f
C3046 VDDA.t329 GNDA 0.019603f
C3047 VDDA.n562 GNDA 0.028154f
C3048 VDDA.n564 GNDA 0.017139f
C3049 VDDA.n565 GNDA 0.017282f
C3050 VDDA.t281 GNDA 0.017824f
C3051 VDDA.t248 GNDA 0.01244f
C3052 VDDA.t238 GNDA 0.01244f
C3053 VDDA.t226 GNDA 0.01244f
C3054 VDDA.t246 GNDA 0.01244f
C3055 VDDA.t308 GNDA 0.017824f
C3056 VDDA.n566 GNDA 0.017282f
C3057 VDDA.n567 GNDA 0.018151f
C3058 VDDA.n569 GNDA 0.052474f
C3059 VDDA.n571 GNDA 0.038608f
C3060 VDDA.n572 GNDA 0.038143f
C3061 VDDA.n573 GNDA 0.040127f
C3062 VDDA.n574 GNDA 0.03158f
C3063 VDDA.n575 GNDA 0.035942f
C3064 VDDA.n576 GNDA 0.035942f
C3065 VDDA.n577 GNDA 0.035942f
C3066 VDDA.n578 GNDA 0.03158f
C3067 VDDA.n579 GNDA 0.040127f
C3068 VDDA.n580 GNDA 0.038143f
C3069 VDDA.n582 GNDA 0.038608f
C3070 VDDA.n584 GNDA 0.038608f
C3071 VDDA.n585 GNDA 0.038143f
C3072 VDDA.n586 GNDA 0.045459f
C3073 VDDA.n587 GNDA 0.037881f
C3074 VDDA.n588 GNDA 0.093443f
C3075 VDDA.n589 GNDA 0.079004f
C3076 VDDA.n594 GNDA 0.045561f
C3077 VDDA.n595 GNDA 0.048469f
C3078 VDDA.n596 GNDA 0.013571f
C3079 VDDA.n603 GNDA 0.013087f
C3080 VDDA.n604 GNDA 0.012117f
C3081 VDDA.n605 GNDA 0.012117f
C3082 VDDA.n613 GNDA 0.013571f
C3083 VDDA.n614 GNDA 0.013571f
C3084 VDDA.n615 GNDA 0.013087f
C3085 VDDA.n623 GNDA 0.012117f
C3086 VDDA.n624 GNDA 0.013087f
C3087 VDDA.n625 GNDA 0.013571f
C3088 VDDA.n633 GNDA 0.013087f
C3089 VDDA.n634 GNDA 0.012117f
C3090 VDDA.n635 GNDA 0.012117f
C3091 VDDA.n643 GNDA 0.040569f
C3092 VDDA.n646 GNDA 5.54772f
C3093 VDDA.n659 GNDA 0.037804f
C3094 VDDA.n660 GNDA 0.013571f
C3095 VDDA.n661 GNDA 0.013087f
C3096 VDDA.n662 GNDA 0.012117f
C3097 VDDA.n663 GNDA 0.012117f
C3098 VDDA.n664 GNDA 0.013087f
C3099 VDDA.n665 GNDA 0.013571f
C3100 VDDA.n666 GNDA 0.013571f
C3101 VDDA.n667 GNDA 0.013087f
C3102 VDDA.n668 GNDA 0.012117f
C3103 VDDA.n669 GNDA 0.012117f
C3104 VDDA.n670 GNDA 0.013087f
C3105 VDDA.n671 GNDA 0.013571f
C3106 VDDA.n672 GNDA 0.013571f
C3107 VDDA.n673 GNDA 0.013087f
C3108 VDDA.n674 GNDA 0.012117f
C3109 VDDA.n675 GNDA 0.012117f
C3110 VDDA.n676 GNDA 0.013087f
C3111 VDDA.n677 GNDA 0.013571f
C3112 VDDA.n718 GNDA 1.29799f
C3113 VDDA.n721 GNDA 0.283542f
C3114 VDDA.n725 GNDA 0.280634f
C3115 VDDA.n727 GNDA 0.086274f
C3116 VDDA.n728 GNDA 0.025026f
C3117 VDDA.n729 GNDA 0.085483f
C3118 VDDA.n730 GNDA 0.025026f
C3119 VDDA.n731 GNDA 0.085483f
C3120 VDDA.n732 GNDA 0.025026f
C3121 VDDA.n733 GNDA 0.085483f
C3122 VDDA.n734 GNDA 0.025026f
C3123 VDDA.n735 GNDA 0.085483f
C3124 VDDA.n736 GNDA 0.0948f
C3125 VDDA.t364 GNDA 0.011761f
C3126 VDDA.n737 GNDA 0.030774f
C3127 VDDA.n738 GNDA 0.114117f
C3128 VDDA.t365 GNDA 0.07391f
C3129 VDDA.t35 GNDA 0.05687f
C3130 VDDA.t372 GNDA 0.05651f
C3131 VDDA.t391 GNDA 0.056099f
C3132 VDDA.t84 GNDA 0.05687f
C3133 VDDA.t111 GNDA 0.05687f
C3134 VDDA.t154 GNDA 0.05687f
C3135 VDDA.t23 GNDA 0.05687f
C3136 VDDA.t104 GNDA 0.05687f
C3137 VDDA.t408 GNDA 0.05687f
C3138 VDDA.t101 GNDA 0.05687f
C3139 VDDA.t260 GNDA 0.07391f
C3140 VDDA.t261 GNDA 0.034115f
C3141 VDDA.n739 GNDA 0.114117f
C3142 VDDA.t259 GNDA 0.011761f
C3143 VDDA.n740 GNDA 0.030774f
C3144 VDDA.n741 GNDA 0.037122f
C3145 VDDA.n742 GNDA 0.028596f
C3146 VDDA.n743 GNDA 0.110509f
C3147 VDDA.n746 GNDA 0.049923f
C3148 VDDA.n747 GNDA 0.049923f
C3149 VDDA.n750 GNDA 0.064376f
C3150 VDDA.n752 GNDA 0.090636f
C3151 VDDA.t138 GNDA 0.025769f
C3152 VDDA.t174 GNDA 0.025769f
C3153 VDDA.t188 GNDA 0.025769f
C3154 VDDA.t42 GNDA 0.025769f
C3155 VDDA.t293 GNDA 0.034471f
C3156 VDDA.t294 GNDA 0.01447f
C3157 VDDA.n753 GNDA 0.040819f
C3158 VDDA.n754 GNDA 0.011338f
C3159 VDDA.n755 GNDA 0.109438f
C3160 VDDA.n756 GNDA 0.014673f
C3161 VDDA.n757 GNDA 0.047529f
C3162 VDDA.n758 GNDA 0.02375f
C3163 VDDA.n763 GNDA 0.067211f
C3164 VDDA.t351 GNDA 0.010014f
C3165 VDDA.n764 GNDA 0.012876f
C3166 VDDA.t255 GNDA 0.025769f
C3167 VDDA.t253 GNDA 0.010014f
C3168 VDDA.n765 GNDA 0.026216f
C3169 VDDA.n766 GNDA 0.064337f
C3170 VDDA.t254 GNDA 0.0482f
C3171 VDDA.t38 GNDA 0.037806f
C3172 VDDA.t352 GNDA 0.0482f
C3173 VDDA.t353 GNDA 0.020115f
C3174 VDDA.n767 GNDA 0.064337f
C3175 VDDA.n768 GNDA 0.025831f
C3176 VDDA.n769 GNDA 0.031841f
C3177 VDDA.n773 GNDA 0.02375f
C3178 VDDA.n775 GNDA 0.012602f
C3179 VDDA.n777 GNDA 0.051862f
C3180 VDDA.n778 GNDA 0.021155f
C3181 VDDA.t363 GNDA 0.010497f
C3182 VDDA.n779 GNDA 0.031604f
C3183 VDDA.t361 GNDA 0.028136f
C3184 VDDA.t194 GNDA 0.021326f
C3185 VDDA.t340 GNDA 0.028136f
C3186 VDDA.t341 GNDA 0.010497f
C3187 VDDA.n780 GNDA 0.031604f
C3188 VDDA.n781 GNDA 0.020771f
C3189 VDDA.n782 GNDA 0.031841f
C3190 VDDA.n783 GNDA 0.02375f
C3191 VDDA.n785 GNDA 0.012602f
C3192 VDDA.n789 GNDA 0.042652f
C3193 VDDA.n790 GNDA 0.042652f
C3194 VDDA.n792 GNDA 0.02375f
C3195 VDDA.n795 GNDA 0.013835f
C3196 VDDA.t264 GNDA 0.01447f
C3197 VDDA.t327 GNDA 0.01447f
C3198 VDDA.n796 GNDA 0.027283f
C3199 VDDA.n797 GNDA 0.023548f
C3200 VDDA.t263 GNDA 0.028698f
C3201 VDDA.t407 GNDA 0.025769f
C3202 VDDA.t16 GNDA 0.025769f
C3203 VDDA.t132 GNDA 0.025769f
C3204 VDDA.t22 GNDA 0.025769f
C3205 VDDA.t337 GNDA 0.034471f
C3206 VDDA.n798 GNDA 0.040819f
C3207 VDDA.n799 GNDA 0.011337f
C3208 VDDA.n800 GNDA 0.109438f
C3209 VDDA.n803 GNDA 0.014205f
C3210 VDDA.n804 GNDA 0.041373f
C3211 VDDA.t354 GNDA 0.010014f
C3212 VDDA.n805 GNDA 0.014205f
C3213 VDDA.n806 GNDA 0.041373f
C3214 VDDA.n807 GNDA 0.014205f
C3215 VDDA.n808 GNDA 0.041373f
C3216 VDDA.n809 GNDA 0.014205f
C3217 VDDA.n810 GNDA 0.041373f
C3218 VDDA.n811 GNDA 0.014205f
C3219 VDDA.n812 GNDA 0.046145f
C3220 VDDA.n813 GNDA 0.021395f
C3221 VDDA.t356 GNDA 0.020115f
C3222 VDDA.n814 GNDA 0.064337f
C3223 VDDA.t355 GNDA 0.0482f
C3224 VDDA.t95 GNDA 0.037806f
C3225 VDDA.t27 GNDA 0.037806f
C3226 VDDA.t97 GNDA 0.037806f
C3227 VDDA.t52 GNDA 0.037806f
C3228 VDDA.t380 GNDA 0.037806f
C3229 VDDA.t198 GNDA 0.037806f
C3230 VDDA.t58 GNDA 0.037806f
C3231 VDDA.t54 GNDA 0.037806f
C3232 VDDA.t91 GNDA 0.037806f
C3233 VDDA.t62 GNDA 0.037806f
C3234 VDDA.t317 GNDA 0.0482f
C3235 VDDA.t318 GNDA 0.020115f
C3236 VDDA.n815 GNDA 0.064337f
C3237 VDDA.t316 GNDA 0.010014f
C3238 VDDA.n816 GNDA 0.020998f
C3239 VDDA.n817 GNDA 0.022543f
C3240 VDDA.n819 GNDA 0.064378f
C3241 VDDA.n821 GNDA 0.090636f
C3242 VDDA.n822 GNDA 0.049923f
C3243 VDDA.n832 GNDA 0.013673f
C3244 VDDA.n833 GNDA 0.013462f
C3245 VDDA.n834 GNDA 0.105669f
C3246 VDDA.n835 GNDA 0.013462f
C3247 VDDA.n836 GNDA 0.056333f
C3248 VDDA.n837 GNDA 0.013462f
C3249 VDDA.n838 GNDA 0.056333f
C3250 VDDA.n839 GNDA 0.013462f
C3251 VDDA.n840 GNDA 0.056333f
C3252 VDDA.n841 GNDA 0.013462f
C3253 VDDA.n842 GNDA 0.07572f
C3254 VDDA.n843 GNDA 0.033928f
C3255 VDDA.n845 GNDA 0.103238f
C3256 VDDA.n847 GNDA 0.103238f
C3257 VDDA.n849 GNDA 0.041982f
C3258 VDDA.t312 GNDA 0.011528f
C3259 VDDA.n850 GNDA 0.035415f
C3260 VDDA.t311 GNDA 0.02872f
C3261 VDDA.t182 GNDA 0.021326f
C3262 VDDA.t125 GNDA 0.021326f
C3263 VDDA.t110 GNDA 0.021326f
C3264 VDDA.t66 GNDA 0.021326f
C3265 VDDA.t116 GNDA 0.021326f
C3266 VDDA.t75 GNDA 0.021326f
C3267 VDDA.t185 GNDA 0.021326f
C3268 VDDA.t88 GNDA 0.021326f
C3269 VDDA.t183 GNDA 0.021326f
C3270 VDDA.t113 GNDA 0.021326f
C3271 VDDA.t302 GNDA 0.02872f
C3272 VDDA.t303 GNDA 0.011528f
C3273 VDDA.n851 GNDA 0.035415f
C3274 VDDA.n852 GNDA 0.025384f
C3275 VDDA.n853 GNDA 0.14734f
C3276 VDDA.n854 GNDA 0.028596f
C3277 VDDA.n856 GNDA 0.110509f
C3278 VDDA.n857 GNDA 0.110509f
C3279 VDDA.n860 GNDA 0.049923f
C3280 VDDA.n862 GNDA 0.028596f
C3281 VDDA.n863 GNDA 0.025026f
C3282 VDDA.n864 GNDA 0.085483f
C3283 VDDA.n865 GNDA 0.025026f
C3284 VDDA.n866 GNDA 0.085483f
C3285 VDDA.n867 GNDA 0.025026f
C3286 VDDA.n868 GNDA 0.085483f
C3287 VDDA.n869 GNDA 0.025026f
C3288 VDDA.n870 GNDA 0.085483f
C3289 VDDA.n871 GNDA 0.037122f
C3290 VDDA.t274 GNDA 0.011761f
C3291 VDDA.n872 GNDA 0.030774f
C3292 VDDA.n873 GNDA 0.114117f
C3293 VDDA.t275 GNDA 0.07391f
C3294 VDDA.t86 GNDA 0.05687f
C3295 VDDA.t7 GNDA 0.05687f
C3296 VDDA.t147 GNDA 0.05687f
C3297 VDDA.t64 GNDA 0.05687f
C3298 VDDA.t108 GNDA 0.05687f
C3299 VDDA.t411 GNDA 0.05687f
C3300 VDDA.t3 GNDA 0.05687f
C3301 VDDA.t117 GNDA 0.05687f
C3302 VDDA.t5 GNDA 0.05687f
C3303 VDDA.t114 GNDA 0.05687f
C3304 VDDA.t287 GNDA 0.07391f
C3305 VDDA.t288 GNDA 0.034115f
C3306 VDDA.n874 GNDA 0.114117f
C3307 VDDA.t286 GNDA 0.011761f
C3308 VDDA.n875 GNDA 0.030774f
C3309 VDDA.n876 GNDA 0.0948f
C3310 VDDA.n877 GNDA 0.086274f
C3311 VDDA.n881 GNDA 0.280634f
C3312 VDDA.n882 GNDA 0.283542f
C3313 VDDA.n885 GNDA 49.264397f
C3314 VDDA.n886 GNDA 0.116325f
C3315 VDDA.n887 GNDA 0.116325f
C3316 VDDA.n888 GNDA 0.116325f
C3317 VDDA.n889 GNDA 0.116325f
C3318 VDDA.n890 GNDA 0.116325f
C3319 VDDA.n891 GNDA 0.116325f
C3320 VDDA.n892 GNDA 0.116325f
C3321 VDDA.n893 GNDA 0.116325f
C3322 VDDA.n894 GNDA 0.116325f
C3323 VDDA.n895 GNDA 0.116325f
C3324 VDDA.n896 GNDA 0.116325f
C3325 VDDA.n897 GNDA 0.116325f
C3326 VDDA.n898 GNDA 0.116325f
C3327 VDDA.n899 GNDA 0.116325f
C3328 VDDA.n900 GNDA 0.116325f
C3329 VDDA.n901 GNDA 0.116325f
C3330 VDDA.n902 GNDA 0.112326f
C3331 VDDA.n904 GNDA 0.116325f
C3332 VDDA.n907 GNDA 0.116325f
C3333 VDDA.n910 GNDA 0.116325f
C3334 VDDA.n913 GNDA 0.116325f
C3335 VDDA.n916 GNDA 0.116325f
C3336 VDDA.n919 GNDA 0.116325f
C3337 VDDA.n922 GNDA 0.116325f
C3338 VDDA.n925 GNDA 0.116325f
C3339 VDDA.n928 GNDA 0.116325f
C3340 VDDA.n931 GNDA 0.116325f
C3341 VDDA.n934 GNDA 0.116325f
C3342 VDDA.n937 GNDA 0.116325f
C3343 VDDA.n940 GNDA 0.116325f
C3344 VDDA.n943 GNDA 0.116325f
C3345 VDDA.n946 GNDA 0.116325f
C3346 VDDA.n949 GNDA 0.116325f
C3347 VDDA.n952 GNDA 0.112326f
C3348 VDDA.n953 GNDA 0.112326f
C3349 VDDA.n954 GNDA 0.112326f
C3350 VDDA.n955 GNDA 0.112326f
C3351 VDDA.n956 GNDA 0.112326f
C3352 VDDA.n957 GNDA 0.112326f
C3353 VDDA.n958 GNDA 0.112326f
C3354 VDDA.n959 GNDA 0.112326f
C3355 VDDA.n960 GNDA 0.112326f
C3356 VDDA.n961 GNDA 0.112326f
C3357 VDDA.n962 GNDA 0.112326f
C3358 VDDA.n963 GNDA 0.112326f
C3359 VDDA.n964 GNDA 0.112326f
C3360 VDDA.n965 GNDA 0.112326f
C3361 VDDA.n966 GNDA 0.112326f
C3362 VDDA.n969 GNDA 0.112326f
C3363 VDDA.n971 GNDA 0.112326f
C3364 VDDA.n973 GNDA 0.112326f
C3365 VDDA.n975 GNDA 0.112326f
C3366 VDDA.n977 GNDA 0.112326f
C3367 VDDA.n979 GNDA 0.112326f
C3368 VDDA.n981 GNDA 0.112326f
C3369 VDDA.n983 GNDA 0.112326f
C3370 VDDA.n985 GNDA 0.112326f
C3371 VDDA.n987 GNDA 0.112326f
C3372 VDDA.n989 GNDA 0.112326f
C3373 VDDA.n991 GNDA 0.112326f
C3374 VDDA.n993 GNDA 0.112326f
C3375 VDDA.n995 GNDA 0.112326f
C3376 VDDA.n997 GNDA 0.112326f
C3377 VDDA.n998 GNDA 0.116325f
C3378 VDDA.n999 GNDA 48.166103f
C3379 VDDA.n1000 GNDA 0.759343f
C3380 bgr_11_0.PFET_GATE_10uA.t28 GNDA 0.023794f
C3381 bgr_11_0.PFET_GATE_10uA.t20 GNDA 0.023794f
C3382 bgr_11_0.PFET_GATE_10uA.n0 GNDA 0.083312f
C3383 bgr_11_0.PFET_GATE_10uA.t13 GNDA 0.0205f
C3384 bgr_11_0.PFET_GATE_10uA.t24 GNDA 0.030304f
C3385 bgr_11_0.PFET_GATE_10uA.n1 GNDA 0.033392f
C3386 bgr_11_0.PFET_GATE_10uA.t17 GNDA 0.0205f
C3387 bgr_11_0.PFET_GATE_10uA.t25 GNDA 0.030304f
C3388 bgr_11_0.PFET_GATE_10uA.n2 GNDA 0.033392f
C3389 bgr_11_0.PFET_GATE_10uA.n3 GNDA 0.032711f
C3390 bgr_11_0.PFET_GATE_10uA.n4 GNDA 1.04203f
C3391 bgr_11_0.PFET_GATE_10uA.t0 GNDA 0.366192f
C3392 bgr_11_0.PFET_GATE_10uA.t1 GNDA 0.326518f
C3393 bgr_11_0.PFET_GATE_10uA.t3 GNDA 0.021026f
C3394 bgr_11_0.PFET_GATE_10uA.t6 GNDA 0.021026f
C3395 bgr_11_0.PFET_GATE_10uA.n5 GNDA 0.045417f
C3396 bgr_11_0.PFET_GATE_10uA.n6 GNDA 1.1272f
C3397 bgr_11_0.PFET_GATE_10uA.t8 GNDA 0.021026f
C3398 bgr_11_0.PFET_GATE_10uA.t4 GNDA 0.021026f
C3399 bgr_11_0.PFET_GATE_10uA.n7 GNDA 0.045417f
C3400 bgr_11_0.PFET_GATE_10uA.n8 GNDA 0.4592f
C3401 bgr_11_0.PFET_GATE_10uA.t7 GNDA 0.021026f
C3402 bgr_11_0.PFET_GATE_10uA.t9 GNDA 0.021026f
C3403 bgr_11_0.PFET_GATE_10uA.n9 GNDA 0.045417f
C3404 bgr_11_0.PFET_GATE_10uA.n10 GNDA 0.449738f
C3405 bgr_11_0.PFET_GATE_10uA.t5 GNDA 0.021026f
C3406 bgr_11_0.PFET_GATE_10uA.t2 GNDA 0.021026f
C3407 bgr_11_0.PFET_GATE_10uA.n11 GNDA 0.045417f
C3408 bgr_11_0.PFET_GATE_10uA.n12 GNDA 0.705894f
C3409 bgr_11_0.PFET_GATE_10uA.n13 GNDA 3.0232f
C3410 bgr_11_0.PFET_GATE_10uA.t26 GNDA 0.070186f
C3411 bgr_11_0.PFET_GATE_10uA.n14 GNDA 1.60401f
C3412 bgr_11_0.PFET_GATE_10uA.t15 GNDA 0.0205f
C3413 bgr_11_0.PFET_GATE_10uA.t10 GNDA 0.030304f
C3414 bgr_11_0.PFET_GATE_10uA.n15 GNDA 0.033392f
C3415 bgr_11_0.PFET_GATE_10uA.t21 GNDA 0.0205f
C3416 bgr_11_0.PFET_GATE_10uA.t11 GNDA 0.030304f
C3417 bgr_11_0.PFET_GATE_10uA.n16 GNDA 0.033392f
C3418 bgr_11_0.PFET_GATE_10uA.n17 GNDA 0.032711f
C3419 bgr_11_0.PFET_GATE_10uA.n18 GNDA 1.30957f
C3420 bgr_11_0.PFET_GATE_10uA.t14 GNDA 0.0205f
C3421 bgr_11_0.PFET_GATE_10uA.t19 GNDA 0.0205f
C3422 bgr_11_0.PFET_GATE_10uA.t18 GNDA 0.0205f
C3423 bgr_11_0.PFET_GATE_10uA.t27 GNDA 0.030304f
C3424 bgr_11_0.PFET_GATE_10uA.n19 GNDA 0.037504f
C3425 bgr_11_0.PFET_GATE_10uA.n20 GNDA 0.026808f
C3426 bgr_11_0.PFET_GATE_10uA.n21 GNDA 0.020894f
C3427 bgr_11_0.PFET_GATE_10uA.t23 GNDA 0.0205f
C3428 bgr_11_0.PFET_GATE_10uA.t16 GNDA 0.0205f
C3429 bgr_11_0.PFET_GATE_10uA.t12 GNDA 0.0205f
C3430 bgr_11_0.PFET_GATE_10uA.t22 GNDA 0.030304f
C3431 bgr_11_0.PFET_GATE_10uA.n22 GNDA 0.037504f
C3432 bgr_11_0.PFET_GATE_10uA.n23 GNDA 0.026808f
C3433 bgr_11_0.PFET_GATE_10uA.n24 GNDA 0.020894f
C3434 bgr_11_0.PFET_GATE_10uA.n25 GNDA 0.059482f
C3435 bgr_11_0.1st_Vout_2.n0 GNDA 1.07305f
C3436 bgr_11_0.1st_Vout_2.n1 GNDA 0.297625f
C3437 bgr_11_0.1st_Vout_2.n2 GNDA 0.668271f
C3438 bgr_11_0.1st_Vout_2.n3 GNDA 0.091542f
C3439 bgr_11_0.1st_Vout_2.n4 GNDA 0.158156f
C3440 bgr_11_0.1st_Vout_2.t14 GNDA 0.011681f
C3441 bgr_11_0.1st_Vout_2.n6 GNDA 0.010675f
C3442 bgr_11_0.1st_Vout_2.n7 GNDA 0.115898f
C3443 bgr_11_0.1st_Vout_2.n8 GNDA 0.0146f
C3444 bgr_11_0.1st_Vout_2.t15 GNDA 0.011528f
C3445 bgr_11_0.1st_Vout_2.t29 GNDA 0.194725f
C3446 bgr_11_0.1st_Vout_2.t32 GNDA 0.198042f
C3447 bgr_11_0.1st_Vout_2.t27 GNDA 0.194725f
C3448 bgr_11_0.1st_Vout_2.t20 GNDA 0.194725f
C3449 bgr_11_0.1st_Vout_2.t12 GNDA 0.198042f
C3450 bgr_11_0.1st_Vout_2.t13 GNDA 0.198042f
C3451 bgr_11_0.1st_Vout_2.t31 GNDA 0.194725f
C3452 bgr_11_0.1st_Vout_2.t25 GNDA 0.194725f
C3453 bgr_11_0.1st_Vout_2.t19 GNDA 0.198042f
C3454 bgr_11_0.1st_Vout_2.t30 GNDA 0.198042f
C3455 bgr_11_0.1st_Vout_2.t24 GNDA 0.194725f
C3456 bgr_11_0.1st_Vout_2.t18 GNDA 0.194725f
C3457 bgr_11_0.1st_Vout_2.t11 GNDA 0.198042f
C3458 bgr_11_0.1st_Vout_2.t23 GNDA 0.198042f
C3459 bgr_11_0.1st_Vout_2.t17 GNDA 0.194725f
C3460 bgr_11_0.1st_Vout_2.t10 GNDA 0.194725f
C3461 bgr_11_0.1st_Vout_2.t28 GNDA 0.198042f
C3462 bgr_11_0.1st_Vout_2.t8 GNDA 0.198042f
C3463 bgr_11_0.1st_Vout_2.t16 GNDA 0.194725f
C3464 bgr_11_0.1st_Vout_2.t22 GNDA 0.194725f
C3465 bgr_11_0.1st_Vout_2.n9 GNDA 0.641071f
C3466 bgr_11_0.1st_Vout_2.n10 GNDA 0.010675f
C3467 bgr_11_0.1st_Vout_2.n11 GNDA 0.0146f
C3468 bgr_11_0.1st_Vout_2.n12 GNDA 0.14235f
C3469 bgr_11_0.1st_Vout_2.t5 GNDA 0.044569f
.ends

