magic
tech sky130A
timestamp 1748793413
<< metal3 >>
rect -15 130 215 215
rect 335 130 565 215
rect 685 130 915 215
rect 1035 130 1265 215
rect 1385 130 1615 215
rect -15 80 1615 130
rect -15 -15 215 80
rect 335 -15 565 80
rect 685 -15 915 80
rect 1035 -15 1265 80
rect 1385 -15 1615 80
rect 75 -135 125 -15
rect -15 -220 215 -135
rect 335 -220 565 -135
rect 685 -220 915 -135
rect 1035 -220 1265 -135
rect 1385 -220 1615 -135
rect -15 -270 1615 -220
rect -15 -365 215 -270
rect 335 -365 565 -270
rect 685 -365 915 -270
rect 1035 -365 1265 -270
rect 1385 -365 1615 -270
rect 75 -485 125 -365
rect -15 -570 215 -485
rect 335 -570 565 -485
rect 685 -570 915 -485
rect 1035 -570 1265 -485
rect 1385 -570 1615 -485
rect -15 -620 1615 -570
rect -15 -715 215 -620
rect 335 -715 565 -620
rect 685 -715 915 -620
rect 1035 -715 1265 -620
rect 1385 -715 1615 -620
rect 75 -835 125 -715
rect -15 -920 215 -835
rect 335 -920 565 -835
rect 685 -920 915 -835
rect 1035 -920 1265 -835
rect 1385 -920 1615 -835
rect -15 -970 1615 -920
rect -15 -1065 215 -970
rect 335 -1065 565 -970
rect 685 -1065 915 -970
rect 1035 -1065 1265 -970
rect 1385 -1065 1615 -970
rect 75 -1185 125 -1065
rect -15 -1270 215 -1185
rect 335 -1270 565 -1185
rect 685 -1270 915 -1185
rect 1035 -1270 1265 -1185
rect 1385 -1270 1615 -1185
rect -15 -1320 1615 -1270
rect -15 -1415 215 -1320
rect 335 -1415 565 -1320
rect 685 -1415 915 -1320
rect 1035 -1415 1265 -1320
rect 1385 -1415 1615 -1320
<< mimcap >>
rect 0 125 200 200
rect 0 85 80 125
rect 120 85 200 125
rect 0 0 200 85
rect 350 125 550 200
rect 350 85 430 125
rect 470 85 550 125
rect 350 0 550 85
rect 700 125 900 200
rect 700 85 780 125
rect 820 85 900 125
rect 700 0 900 85
rect 1050 125 1250 200
rect 1050 85 1130 125
rect 1170 85 1250 125
rect 1050 0 1250 85
rect 1400 125 1600 200
rect 1400 85 1480 125
rect 1520 85 1600 125
rect 1400 0 1600 85
rect 0 -225 200 -150
rect 0 -265 80 -225
rect 120 -265 200 -225
rect 0 -350 200 -265
rect 350 -225 550 -150
rect 350 -265 430 -225
rect 470 -265 550 -225
rect 350 -350 550 -265
rect 700 -225 900 -150
rect 700 -265 780 -225
rect 820 -265 900 -225
rect 700 -350 900 -265
rect 1050 -225 1250 -150
rect 1050 -265 1130 -225
rect 1170 -265 1250 -225
rect 1050 -350 1250 -265
rect 1400 -225 1600 -150
rect 1400 -265 1480 -225
rect 1520 -265 1600 -225
rect 1400 -350 1600 -265
rect 0 -575 200 -500
rect 0 -615 80 -575
rect 120 -615 200 -575
rect 0 -700 200 -615
rect 350 -575 550 -500
rect 350 -615 430 -575
rect 470 -615 550 -575
rect 350 -700 550 -615
rect 700 -575 900 -500
rect 700 -615 780 -575
rect 820 -615 900 -575
rect 700 -700 900 -615
rect 1050 -575 1250 -500
rect 1050 -615 1130 -575
rect 1170 -615 1250 -575
rect 1050 -700 1250 -615
rect 1400 -575 1600 -500
rect 1400 -615 1480 -575
rect 1520 -615 1600 -575
rect 1400 -700 1600 -615
rect 0 -925 200 -850
rect 0 -965 80 -925
rect 120 -965 200 -925
rect 0 -1050 200 -965
rect 350 -925 550 -850
rect 350 -965 430 -925
rect 470 -965 550 -925
rect 350 -1050 550 -965
rect 700 -925 900 -850
rect 700 -965 780 -925
rect 820 -965 900 -925
rect 700 -1050 900 -965
rect 1050 -925 1250 -850
rect 1050 -965 1130 -925
rect 1170 -965 1250 -925
rect 1050 -1050 1250 -965
rect 1400 -925 1600 -850
rect 1400 -965 1480 -925
rect 1520 -965 1600 -925
rect 1400 -1050 1600 -965
rect 0 -1275 200 -1200
rect 0 -1315 80 -1275
rect 120 -1315 200 -1275
rect 0 -1400 200 -1315
rect 350 -1275 550 -1200
rect 350 -1315 430 -1275
rect 470 -1315 550 -1275
rect 350 -1400 550 -1315
rect 700 -1275 900 -1200
rect 700 -1315 780 -1275
rect 820 -1315 900 -1275
rect 700 -1400 900 -1315
rect 1050 -1275 1250 -1200
rect 1050 -1315 1130 -1275
rect 1170 -1315 1250 -1275
rect 1050 -1400 1250 -1315
rect 1400 -1275 1600 -1200
rect 1400 -1315 1480 -1275
rect 1520 -1315 1600 -1275
rect 1400 -1400 1600 -1315
<< mimcapcontact >>
rect 80 85 120 125
rect 430 85 470 125
rect 780 85 820 125
rect 1130 85 1170 125
rect 1480 85 1520 125
rect 80 -265 120 -225
rect 430 -265 470 -225
rect 780 -265 820 -225
rect 1130 -265 1170 -225
rect 1480 -265 1520 -225
rect 80 -615 120 -575
rect 430 -615 470 -575
rect 780 -615 820 -575
rect 1130 -615 1170 -575
rect 1480 -615 1520 -575
rect 80 -965 120 -925
rect 430 -965 470 -925
rect 780 -965 820 -925
rect 1130 -965 1170 -925
rect 1480 -965 1520 -925
rect 80 -1315 120 -1275
rect 430 -1315 470 -1275
rect 780 -1315 820 -1275
rect 1130 -1315 1170 -1275
rect 1480 -1315 1520 -1275
<< metal4 >>
rect 75 125 1525 130
rect 75 85 80 125
rect 120 85 430 125
rect 470 85 780 125
rect 820 85 1130 125
rect 1170 85 1480 125
rect 1520 85 1525 125
rect 75 80 1525 85
rect 75 -220 125 80
rect 75 -225 1525 -220
rect 75 -265 80 -225
rect 120 -265 430 -225
rect 470 -265 780 -225
rect 820 -265 1130 -225
rect 1170 -265 1480 -225
rect 1520 -265 1525 -225
rect 75 -270 1525 -265
rect 75 -570 125 -270
rect 75 -575 1525 -570
rect 75 -615 80 -575
rect 120 -615 430 -575
rect 470 -615 780 -575
rect 820 -615 1130 -575
rect 1170 -615 1480 -575
rect 1520 -615 1525 -575
rect 75 -620 1525 -615
rect 75 -920 125 -620
rect 75 -925 1525 -920
rect 75 -965 80 -925
rect 120 -965 430 -925
rect 470 -965 780 -925
rect 820 -965 1130 -925
rect 1170 -965 1480 -925
rect 1520 -965 1525 -925
rect 75 -970 1525 -965
rect 75 -1270 125 -970
rect 75 -1275 1525 -1270
rect 75 -1315 80 -1275
rect 120 -1315 430 -1275
rect 470 -1315 780 -1275
rect 820 -1315 1130 -1275
rect 1170 -1315 1480 -1275
rect 1520 -1315 1525 -1275
rect 75 -1320 1525 -1315
<< end >>
