magic
tech sky130A
timestamp 1754058664
<< nwell >>
rect 16315 1270 16695 1410
rect 16825 1270 17315 1410
rect 17445 1270 18155 1410
rect 18285 1270 18775 1410
rect 16375 705 16760 845
rect 16910 605 18690 945
rect 18845 705 19170 945
rect 16360 -35 17725 105
rect 17880 -35 19240 105
<< pwell >>
rect 17780 -4300 17820 -4120
<< nmos >>
rect 17000 -450 17020 -200
rect 17060 -450 17080 -200
rect 18520 -450 18540 -200
rect 18580 -450 18600 -200
rect 16570 -985 17070 -735
rect 17190 -985 17690 -735
rect 17910 -985 18410 -735
rect 18530 -985 19030 -735
rect 16780 -1290 17780 -1190
rect 17820 -1290 18820 -1190
rect 16580 -1640 16595 -1540
rect 16635 -1640 16650 -1540
rect 16690 -1640 16705 -1540
rect 16745 -1640 16760 -1540
rect 16800 -1640 16815 -1540
rect 17065 -1640 17080 -1540
rect 17120 -1640 17135 -1540
rect 17175 -1640 17190 -1540
rect 17230 -1640 17245 -1540
rect 17285 -1640 17300 -1540
rect 17340 -1640 17355 -1540
rect 17395 -1640 17410 -1540
rect 17450 -1640 17465 -1540
rect 17655 -1640 17670 -1540
rect 17710 -1640 17725 -1540
rect 17765 -1640 17780 -1540
rect 17820 -1640 17835 -1540
rect 17875 -1640 17890 -1540
rect 17930 -1640 17945 -1540
rect 18135 -1640 18150 -1540
rect 18190 -1640 18205 -1540
rect 18245 -1640 18260 -1540
rect 18300 -1640 18315 -1540
rect 18355 -1640 18370 -1540
rect 18410 -1640 18425 -1540
rect 18465 -1640 18480 -1540
rect 18520 -1640 18535 -1540
<< pmos >>
rect 16415 1290 16430 1390
rect 16470 1290 16485 1390
rect 16525 1290 16540 1390
rect 16580 1290 16595 1390
rect 16925 1290 16940 1390
rect 16980 1290 16995 1390
rect 17035 1290 17050 1390
rect 17090 1290 17105 1390
rect 17145 1290 17160 1390
rect 17200 1290 17215 1390
rect 17545 1290 17560 1390
rect 17600 1290 17615 1390
rect 17655 1290 17670 1390
rect 17710 1290 17725 1390
rect 17765 1290 17780 1390
rect 17820 1290 17835 1390
rect 17875 1290 17890 1390
rect 17930 1290 17945 1390
rect 17985 1290 18000 1390
rect 18040 1290 18055 1390
rect 18385 1290 18400 1390
rect 18440 1290 18455 1390
rect 18495 1290 18510 1390
rect 18550 1290 18565 1390
rect 18605 1290 18620 1390
rect 18660 1290 18675 1390
rect 16475 725 16490 825
rect 16530 725 16545 825
rect 16585 725 16600 825
rect 16640 725 16655 825
rect 17010 625 17060 925
rect 17100 625 17150 925
rect 17190 625 17240 925
rect 17280 625 17330 925
rect 17370 625 17420 925
rect 17460 625 17510 925
rect 17550 625 17600 925
rect 17640 625 17690 925
rect 17730 625 17780 925
rect 17820 625 17870 925
rect 17910 625 17960 925
rect 18000 625 18050 925
rect 18090 625 18140 925
rect 18180 625 18230 925
rect 18270 625 18320 925
rect 18360 625 18410 925
rect 18450 625 18500 925
rect 18540 625 18590 925
rect 18945 725 18960 925
rect 19000 725 19015 925
rect 19055 725 19070 925
rect 16460 -15 16480 85
rect 16520 -15 16540 85
rect 16580 -15 16600 85
rect 16640 -15 16660 85
rect 16700 -15 16720 85
rect 16760 -15 16780 85
rect 16820 -15 16840 85
rect 16880 -15 16900 85
rect 16940 -15 16960 85
rect 17000 -15 17020 85
rect 17060 -15 17080 85
rect 17120 -15 17140 85
rect 17180 -15 17200 85
rect 17240 -15 17260 85
rect 17300 -15 17320 85
rect 17360 -15 17380 85
rect 17420 -15 17440 85
rect 17480 -15 17500 85
rect 17540 -15 17560 85
rect 17600 -15 17620 85
rect 17980 -15 18000 85
rect 18040 -15 18060 85
rect 18100 -15 18120 85
rect 18160 -15 18180 85
rect 18220 -15 18240 85
rect 18280 -15 18300 85
rect 18340 -15 18360 85
rect 18400 -15 18420 85
rect 18460 -15 18480 85
rect 18520 -15 18540 85
rect 18580 -15 18600 85
rect 18640 -15 18660 85
rect 18700 -15 18720 85
rect 18760 -15 18780 85
rect 18820 -15 18840 85
rect 18880 -15 18900 85
rect 18940 -15 18960 85
rect 19000 -15 19020 85
rect 19060 -15 19080 85
rect 19120 -15 19140 85
<< ndiff >>
rect 16960 -215 17000 -200
rect 16960 -235 16970 -215
rect 16990 -235 17000 -215
rect 16960 -265 17000 -235
rect 16960 -285 16970 -265
rect 16990 -285 17000 -265
rect 16960 -315 17000 -285
rect 16960 -335 16970 -315
rect 16990 -335 17000 -315
rect 16960 -365 17000 -335
rect 16960 -385 16970 -365
rect 16990 -385 17000 -365
rect 16960 -415 17000 -385
rect 16960 -435 16970 -415
rect 16990 -435 17000 -415
rect 16960 -450 17000 -435
rect 17020 -215 17060 -200
rect 17020 -235 17030 -215
rect 17050 -235 17060 -215
rect 17020 -265 17060 -235
rect 17020 -285 17030 -265
rect 17050 -285 17060 -265
rect 17020 -315 17060 -285
rect 17020 -335 17030 -315
rect 17050 -335 17060 -315
rect 17020 -365 17060 -335
rect 17020 -385 17030 -365
rect 17050 -385 17060 -365
rect 17020 -415 17060 -385
rect 17020 -435 17030 -415
rect 17050 -435 17060 -415
rect 17020 -450 17060 -435
rect 17080 -215 17120 -200
rect 17080 -235 17090 -215
rect 17110 -235 17120 -215
rect 17080 -265 17120 -235
rect 17080 -285 17090 -265
rect 17110 -285 17120 -265
rect 17080 -315 17120 -285
rect 17080 -335 17090 -315
rect 17110 -335 17120 -315
rect 18480 -215 18520 -200
rect 18480 -235 18490 -215
rect 18510 -235 18520 -215
rect 18480 -265 18520 -235
rect 18480 -285 18490 -265
rect 18510 -285 18520 -265
rect 18480 -315 18520 -285
rect 17080 -365 17120 -335
rect 17080 -385 17090 -365
rect 17110 -385 17120 -365
rect 17080 -415 17120 -385
rect 17080 -435 17090 -415
rect 17110 -435 17120 -415
rect 17080 -450 17120 -435
rect 18480 -335 18490 -315
rect 18510 -335 18520 -315
rect 18480 -365 18520 -335
rect 18480 -385 18490 -365
rect 18510 -385 18520 -365
rect 18480 -415 18520 -385
rect 18480 -435 18490 -415
rect 18510 -435 18520 -415
rect 18480 -450 18520 -435
rect 18540 -215 18580 -200
rect 18540 -235 18550 -215
rect 18570 -235 18580 -215
rect 18540 -265 18580 -235
rect 18540 -285 18550 -265
rect 18570 -285 18580 -265
rect 18540 -315 18580 -285
rect 18540 -335 18550 -315
rect 18570 -335 18580 -315
rect 18540 -365 18580 -335
rect 18540 -385 18550 -365
rect 18570 -385 18580 -365
rect 18540 -415 18580 -385
rect 18540 -435 18550 -415
rect 18570 -435 18580 -415
rect 18540 -450 18580 -435
rect 18600 -215 18640 -200
rect 18600 -235 18610 -215
rect 18630 -235 18640 -215
rect 18600 -265 18640 -235
rect 18600 -285 18610 -265
rect 18630 -285 18640 -265
rect 18600 -315 18640 -285
rect 18600 -335 18610 -315
rect 18630 -335 18640 -315
rect 18600 -365 18640 -335
rect 18600 -385 18610 -365
rect 18630 -385 18640 -365
rect 18600 -415 18640 -385
rect 18600 -435 18610 -415
rect 18630 -435 18640 -415
rect 18600 -450 18640 -435
rect 16530 -750 16570 -735
rect 16530 -770 16540 -750
rect 16560 -770 16570 -750
rect 16530 -800 16570 -770
rect 16530 -820 16540 -800
rect 16560 -820 16570 -800
rect 16530 -850 16570 -820
rect 16530 -870 16540 -850
rect 16560 -870 16570 -850
rect 16530 -900 16570 -870
rect 16530 -920 16540 -900
rect 16560 -920 16570 -900
rect 16530 -950 16570 -920
rect 16530 -970 16540 -950
rect 16560 -970 16570 -950
rect 16530 -985 16570 -970
rect 17070 -750 17110 -735
rect 17150 -750 17190 -735
rect 17070 -770 17080 -750
rect 17100 -770 17110 -750
rect 17150 -770 17160 -750
rect 17180 -770 17190 -750
rect 17070 -800 17110 -770
rect 17150 -800 17190 -770
rect 17070 -820 17080 -800
rect 17100 -820 17110 -800
rect 17150 -820 17160 -800
rect 17180 -820 17190 -800
rect 17070 -850 17110 -820
rect 17150 -850 17190 -820
rect 17070 -870 17080 -850
rect 17100 -870 17110 -850
rect 17150 -870 17160 -850
rect 17180 -870 17190 -850
rect 17070 -900 17110 -870
rect 17150 -900 17190 -870
rect 17070 -920 17080 -900
rect 17100 -920 17110 -900
rect 17150 -920 17160 -900
rect 17180 -920 17190 -900
rect 17070 -950 17110 -920
rect 17150 -950 17190 -920
rect 17070 -970 17080 -950
rect 17100 -970 17110 -950
rect 17150 -970 17160 -950
rect 17180 -970 17190 -950
rect 17070 -980 17110 -970
rect 17150 -980 17190 -970
rect 17070 -985 17190 -980
rect 17690 -750 17730 -735
rect 17690 -770 17700 -750
rect 17720 -770 17730 -750
rect 17690 -800 17730 -770
rect 17690 -820 17700 -800
rect 17720 -820 17730 -800
rect 17690 -850 17730 -820
rect 17690 -870 17700 -850
rect 17720 -870 17730 -850
rect 17690 -900 17730 -870
rect 17690 -920 17700 -900
rect 17720 -920 17730 -900
rect 17690 -950 17730 -920
rect 17690 -970 17700 -950
rect 17720 -970 17730 -950
rect 17690 -985 17730 -970
rect 17870 -750 17910 -735
rect 17870 -770 17880 -750
rect 17900 -770 17910 -750
rect 17870 -800 17910 -770
rect 17870 -820 17880 -800
rect 17900 -820 17910 -800
rect 17870 -850 17910 -820
rect 17870 -870 17880 -850
rect 17900 -870 17910 -850
rect 17870 -900 17910 -870
rect 17870 -920 17880 -900
rect 17900 -920 17910 -900
rect 17870 -950 17910 -920
rect 17870 -970 17880 -950
rect 17900 -970 17910 -950
rect 17870 -985 17910 -970
rect 18410 -750 18450 -735
rect 18490 -750 18530 -735
rect 18410 -770 18420 -750
rect 18440 -770 18450 -750
rect 18490 -770 18500 -750
rect 18520 -770 18530 -750
rect 18410 -800 18450 -770
rect 18490 -800 18530 -770
rect 18410 -820 18420 -800
rect 18440 -820 18450 -800
rect 18490 -820 18500 -800
rect 18520 -820 18530 -800
rect 18410 -850 18450 -820
rect 18490 -850 18530 -820
rect 18410 -870 18420 -850
rect 18440 -870 18450 -850
rect 18490 -870 18500 -850
rect 18520 -870 18530 -850
rect 18410 -900 18450 -870
rect 18490 -900 18530 -870
rect 18410 -920 18420 -900
rect 18440 -920 18450 -900
rect 18490 -920 18500 -900
rect 18520 -920 18530 -900
rect 18410 -950 18450 -920
rect 18490 -950 18530 -920
rect 18410 -970 18420 -950
rect 18440 -970 18450 -950
rect 18490 -970 18500 -950
rect 18520 -970 18530 -950
rect 18410 -985 18450 -970
rect 18490 -985 18530 -970
rect 19030 -750 19070 -735
rect 19030 -770 19040 -750
rect 19060 -770 19070 -750
rect 19030 -800 19070 -770
rect 19030 -820 19040 -800
rect 19060 -820 19070 -800
rect 19030 -850 19070 -820
rect 19030 -870 19040 -850
rect 19060 -870 19070 -850
rect 19030 -900 19070 -870
rect 19030 -920 19040 -900
rect 19060 -920 19070 -900
rect 19030 -950 19070 -920
rect 19030 -970 19040 -950
rect 19060 -970 19070 -950
rect 19030 -985 19070 -970
rect 16740 -1205 16780 -1190
rect 16740 -1225 16750 -1205
rect 16770 -1225 16780 -1205
rect 16740 -1255 16780 -1225
rect 16740 -1275 16750 -1255
rect 16770 -1275 16780 -1255
rect 16740 -1290 16780 -1275
rect 17780 -1205 17820 -1190
rect 17780 -1225 17790 -1205
rect 17810 -1225 17820 -1205
rect 17780 -1255 17820 -1225
rect 17780 -1275 17790 -1255
rect 17810 -1275 17820 -1255
rect 17780 -1290 17820 -1275
rect 18820 -1205 18860 -1190
rect 18820 -1225 18830 -1205
rect 18850 -1225 18860 -1205
rect 18820 -1255 18860 -1225
rect 18820 -1275 18830 -1255
rect 18850 -1275 18860 -1255
rect 18820 -1290 18860 -1275
rect 16540 -1555 16580 -1540
rect 16540 -1575 16550 -1555
rect 16570 -1575 16580 -1555
rect 16540 -1605 16580 -1575
rect 16540 -1625 16550 -1605
rect 16570 -1625 16580 -1605
rect 16540 -1640 16580 -1625
rect 16595 -1555 16635 -1540
rect 16595 -1575 16605 -1555
rect 16625 -1575 16635 -1555
rect 16595 -1605 16635 -1575
rect 16595 -1625 16605 -1605
rect 16625 -1625 16635 -1605
rect 16595 -1640 16635 -1625
rect 16650 -1555 16690 -1540
rect 16650 -1575 16660 -1555
rect 16680 -1575 16690 -1555
rect 16650 -1605 16690 -1575
rect 16650 -1625 16660 -1605
rect 16680 -1625 16690 -1605
rect 16650 -1640 16690 -1625
rect 16705 -1555 16745 -1540
rect 16705 -1575 16715 -1555
rect 16735 -1575 16745 -1555
rect 16705 -1605 16745 -1575
rect 16705 -1625 16715 -1605
rect 16735 -1625 16745 -1605
rect 16705 -1640 16745 -1625
rect 16760 -1555 16800 -1540
rect 16760 -1575 16770 -1555
rect 16790 -1575 16800 -1555
rect 16760 -1605 16800 -1575
rect 16760 -1625 16770 -1605
rect 16790 -1625 16800 -1605
rect 16760 -1640 16800 -1625
rect 16815 -1555 16855 -1540
rect 16815 -1575 16825 -1555
rect 16845 -1575 16855 -1555
rect 16815 -1605 16855 -1575
rect 16815 -1625 16825 -1605
rect 16845 -1625 16855 -1605
rect 16815 -1640 16855 -1625
rect 17025 -1555 17065 -1540
rect 17025 -1575 17035 -1555
rect 17055 -1575 17065 -1555
rect 17025 -1605 17065 -1575
rect 17025 -1625 17035 -1605
rect 17055 -1625 17065 -1605
rect 17025 -1640 17065 -1625
rect 17080 -1555 17120 -1540
rect 17080 -1575 17090 -1555
rect 17110 -1575 17120 -1555
rect 17080 -1605 17120 -1575
rect 17080 -1625 17090 -1605
rect 17110 -1625 17120 -1605
rect 17080 -1640 17120 -1625
rect 17135 -1555 17175 -1540
rect 17135 -1575 17145 -1555
rect 17165 -1575 17175 -1555
rect 17135 -1605 17175 -1575
rect 17135 -1625 17145 -1605
rect 17165 -1625 17175 -1605
rect 17135 -1640 17175 -1625
rect 17190 -1555 17230 -1540
rect 17190 -1575 17200 -1555
rect 17220 -1575 17230 -1555
rect 17190 -1605 17230 -1575
rect 17190 -1625 17200 -1605
rect 17220 -1625 17230 -1605
rect 17190 -1640 17230 -1625
rect 17245 -1555 17285 -1540
rect 17245 -1575 17255 -1555
rect 17275 -1575 17285 -1555
rect 17245 -1605 17285 -1575
rect 17245 -1625 17255 -1605
rect 17275 -1625 17285 -1605
rect 17245 -1640 17285 -1625
rect 17300 -1555 17340 -1540
rect 17300 -1575 17310 -1555
rect 17330 -1575 17340 -1555
rect 17300 -1605 17340 -1575
rect 17300 -1625 17310 -1605
rect 17330 -1625 17340 -1605
rect 17300 -1640 17340 -1625
rect 17355 -1555 17395 -1540
rect 17355 -1575 17365 -1555
rect 17385 -1575 17395 -1555
rect 17355 -1605 17395 -1575
rect 17355 -1625 17365 -1605
rect 17385 -1625 17395 -1605
rect 17355 -1640 17395 -1625
rect 17410 -1555 17450 -1540
rect 17410 -1575 17420 -1555
rect 17440 -1575 17450 -1555
rect 17410 -1605 17450 -1575
rect 17410 -1625 17420 -1605
rect 17440 -1625 17450 -1605
rect 17410 -1640 17450 -1625
rect 17465 -1555 17505 -1540
rect 17465 -1575 17475 -1555
rect 17495 -1575 17505 -1555
rect 17465 -1605 17505 -1575
rect 17465 -1625 17475 -1605
rect 17495 -1625 17505 -1605
rect 17465 -1640 17505 -1625
rect 17615 -1555 17655 -1540
rect 17615 -1575 17625 -1555
rect 17645 -1575 17655 -1555
rect 17615 -1605 17655 -1575
rect 17615 -1625 17625 -1605
rect 17645 -1625 17655 -1605
rect 17615 -1640 17655 -1625
rect 17670 -1555 17710 -1540
rect 17670 -1575 17680 -1555
rect 17700 -1575 17710 -1555
rect 17670 -1605 17710 -1575
rect 17670 -1625 17680 -1605
rect 17700 -1625 17710 -1605
rect 17670 -1640 17710 -1625
rect 17725 -1555 17765 -1540
rect 17725 -1575 17735 -1555
rect 17755 -1575 17765 -1555
rect 17725 -1605 17765 -1575
rect 17725 -1625 17735 -1605
rect 17755 -1625 17765 -1605
rect 17725 -1640 17765 -1625
rect 17780 -1555 17820 -1540
rect 17780 -1575 17790 -1555
rect 17810 -1575 17820 -1555
rect 17780 -1605 17820 -1575
rect 17780 -1625 17790 -1605
rect 17810 -1625 17820 -1605
rect 17780 -1640 17820 -1625
rect 17835 -1555 17875 -1540
rect 17835 -1575 17845 -1555
rect 17865 -1575 17875 -1555
rect 17835 -1605 17875 -1575
rect 17835 -1625 17845 -1605
rect 17865 -1625 17875 -1605
rect 17835 -1640 17875 -1625
rect 17890 -1555 17930 -1540
rect 17890 -1575 17900 -1555
rect 17920 -1575 17930 -1555
rect 17890 -1605 17930 -1575
rect 17890 -1625 17900 -1605
rect 17920 -1625 17930 -1605
rect 17890 -1640 17930 -1625
rect 17945 -1555 17985 -1540
rect 17945 -1575 17955 -1555
rect 17975 -1575 17985 -1555
rect 17945 -1605 17985 -1575
rect 17945 -1625 17955 -1605
rect 17975 -1625 17985 -1605
rect 17945 -1640 17985 -1625
rect 18095 -1555 18135 -1540
rect 18095 -1575 18105 -1555
rect 18125 -1575 18135 -1555
rect 18095 -1605 18135 -1575
rect 18095 -1625 18105 -1605
rect 18125 -1625 18135 -1605
rect 18095 -1640 18135 -1625
rect 18150 -1555 18190 -1540
rect 18150 -1575 18160 -1555
rect 18180 -1575 18190 -1555
rect 18150 -1605 18190 -1575
rect 18150 -1625 18160 -1605
rect 18180 -1625 18190 -1605
rect 18150 -1640 18190 -1625
rect 18205 -1555 18245 -1540
rect 18205 -1575 18215 -1555
rect 18235 -1575 18245 -1555
rect 18205 -1605 18245 -1575
rect 18205 -1625 18215 -1605
rect 18235 -1625 18245 -1605
rect 18205 -1640 18245 -1625
rect 18260 -1555 18300 -1540
rect 18260 -1575 18270 -1555
rect 18290 -1575 18300 -1555
rect 18260 -1605 18300 -1575
rect 18260 -1625 18270 -1605
rect 18290 -1625 18300 -1605
rect 18260 -1640 18300 -1625
rect 18315 -1555 18355 -1540
rect 18315 -1575 18325 -1555
rect 18345 -1575 18355 -1555
rect 18315 -1605 18355 -1575
rect 18315 -1625 18325 -1605
rect 18345 -1625 18355 -1605
rect 18315 -1640 18355 -1625
rect 18370 -1555 18410 -1540
rect 18370 -1575 18380 -1555
rect 18400 -1575 18410 -1555
rect 18370 -1605 18410 -1575
rect 18370 -1625 18380 -1605
rect 18400 -1625 18410 -1605
rect 18370 -1640 18410 -1625
rect 18425 -1555 18465 -1540
rect 18425 -1575 18435 -1555
rect 18455 -1575 18465 -1555
rect 18425 -1605 18465 -1575
rect 18425 -1625 18435 -1605
rect 18455 -1625 18465 -1605
rect 18425 -1640 18465 -1625
rect 18480 -1555 18520 -1540
rect 18480 -1575 18490 -1555
rect 18510 -1575 18520 -1555
rect 18480 -1605 18520 -1575
rect 18480 -1625 18490 -1605
rect 18510 -1625 18520 -1605
rect 18480 -1640 18520 -1625
rect 18535 -1555 18575 -1540
rect 18535 -1575 18545 -1555
rect 18565 -1575 18575 -1555
rect 18535 -1605 18575 -1575
rect 18535 -1625 18545 -1605
rect 18565 -1625 18575 -1605
rect 18535 -1640 18575 -1625
<< pdiff >>
rect 16375 1375 16415 1390
rect 16375 1355 16385 1375
rect 16405 1355 16415 1375
rect 16375 1325 16415 1355
rect 16375 1305 16385 1325
rect 16405 1305 16415 1325
rect 16375 1290 16415 1305
rect 16430 1375 16470 1390
rect 16430 1355 16440 1375
rect 16460 1355 16470 1375
rect 16430 1325 16470 1355
rect 16430 1305 16440 1325
rect 16460 1305 16470 1325
rect 16430 1290 16470 1305
rect 16485 1375 16525 1390
rect 16485 1355 16495 1375
rect 16515 1355 16525 1375
rect 16485 1325 16525 1355
rect 16485 1305 16495 1325
rect 16515 1305 16525 1325
rect 16485 1290 16525 1305
rect 16540 1375 16580 1390
rect 16540 1355 16550 1375
rect 16570 1355 16580 1375
rect 16540 1325 16580 1355
rect 16540 1305 16550 1325
rect 16570 1305 16580 1325
rect 16540 1290 16580 1305
rect 16595 1375 16635 1390
rect 16595 1355 16605 1375
rect 16625 1355 16635 1375
rect 16595 1325 16635 1355
rect 16595 1305 16605 1325
rect 16625 1305 16635 1325
rect 16595 1290 16635 1305
rect 16885 1375 16925 1390
rect 16885 1303 16895 1375
rect 16915 1303 16925 1375
rect 16885 1290 16925 1303
rect 16940 1375 16980 1390
rect 16940 1303 16950 1375
rect 16970 1303 16980 1375
rect 16940 1290 16980 1303
rect 16995 1375 17035 1390
rect 16995 1303 17005 1375
rect 17025 1303 17035 1375
rect 16995 1290 17035 1303
rect 17050 1375 17090 1390
rect 17050 1303 17060 1375
rect 17080 1303 17090 1375
rect 17050 1290 17090 1303
rect 17105 1375 17145 1390
rect 17105 1303 17115 1375
rect 17135 1303 17145 1375
rect 17105 1290 17145 1303
rect 17160 1375 17200 1390
rect 17160 1303 17170 1375
rect 17190 1303 17200 1375
rect 17160 1290 17200 1303
rect 17215 1375 17255 1390
rect 17215 1303 17225 1375
rect 17245 1303 17255 1375
rect 17215 1290 17255 1303
rect 17505 1375 17545 1390
rect 17505 1355 17515 1375
rect 17535 1355 17545 1375
rect 17505 1325 17545 1355
rect 17505 1305 17515 1325
rect 17535 1305 17545 1325
rect 17505 1290 17545 1305
rect 17560 1375 17600 1390
rect 17560 1355 17570 1375
rect 17590 1355 17600 1375
rect 17560 1325 17600 1355
rect 17560 1305 17570 1325
rect 17590 1305 17600 1325
rect 17560 1290 17600 1305
rect 17615 1375 17655 1390
rect 17615 1355 17625 1375
rect 17645 1355 17655 1375
rect 17615 1325 17655 1355
rect 17615 1305 17625 1325
rect 17645 1305 17655 1325
rect 17615 1290 17655 1305
rect 17670 1375 17710 1390
rect 17670 1355 17680 1375
rect 17700 1355 17710 1375
rect 17670 1325 17710 1355
rect 17670 1305 17680 1325
rect 17700 1305 17710 1325
rect 17670 1290 17710 1305
rect 17725 1375 17765 1390
rect 17725 1355 17735 1375
rect 17755 1355 17765 1375
rect 17725 1325 17765 1355
rect 17725 1305 17735 1325
rect 17755 1305 17765 1325
rect 17725 1290 17765 1305
rect 17780 1375 17820 1390
rect 17780 1355 17790 1375
rect 17810 1355 17820 1375
rect 17780 1325 17820 1355
rect 17780 1305 17790 1325
rect 17810 1305 17820 1325
rect 17780 1290 17820 1305
rect 17835 1375 17875 1390
rect 17835 1355 17845 1375
rect 17865 1355 17875 1375
rect 17835 1325 17875 1355
rect 17835 1305 17845 1325
rect 17865 1305 17875 1325
rect 17835 1290 17875 1305
rect 17890 1375 17930 1390
rect 17890 1355 17900 1375
rect 17920 1355 17930 1375
rect 17890 1325 17930 1355
rect 17890 1305 17900 1325
rect 17920 1305 17930 1325
rect 17890 1290 17930 1305
rect 17945 1375 17985 1390
rect 17945 1355 17955 1375
rect 17975 1355 17985 1375
rect 17945 1325 17985 1355
rect 17945 1305 17955 1325
rect 17975 1305 17985 1325
rect 17945 1290 17985 1305
rect 18000 1375 18040 1390
rect 18000 1355 18010 1375
rect 18030 1355 18040 1375
rect 18000 1325 18040 1355
rect 18000 1305 18010 1325
rect 18030 1305 18040 1325
rect 18000 1290 18040 1305
rect 18055 1375 18095 1390
rect 18055 1355 18065 1375
rect 18085 1355 18095 1375
rect 18055 1325 18095 1355
rect 18055 1305 18065 1325
rect 18085 1305 18095 1325
rect 18055 1290 18095 1305
rect 18345 1375 18385 1390
rect 18345 1305 18355 1375
rect 18375 1305 18385 1375
rect 18345 1290 18385 1305
rect 18400 1375 18440 1390
rect 18400 1305 18410 1375
rect 18430 1305 18440 1375
rect 18400 1290 18440 1305
rect 18455 1375 18495 1390
rect 18455 1305 18465 1375
rect 18485 1305 18495 1375
rect 18455 1290 18495 1305
rect 18510 1375 18550 1390
rect 18510 1305 18520 1375
rect 18540 1305 18550 1375
rect 18510 1290 18550 1305
rect 18565 1375 18605 1390
rect 18565 1305 18575 1375
rect 18595 1305 18605 1375
rect 18565 1290 18605 1305
rect 18620 1375 18660 1390
rect 18620 1305 18630 1375
rect 18650 1305 18660 1375
rect 18620 1290 18660 1305
rect 18675 1375 18715 1390
rect 18675 1305 18685 1375
rect 18705 1305 18715 1375
rect 18675 1290 18715 1305
rect 16970 910 17010 925
rect 16970 890 16980 910
rect 17000 890 17010 910
rect 16970 860 17010 890
rect 16970 840 16980 860
rect 17000 840 17010 860
rect 16435 810 16475 825
rect 16435 790 16445 810
rect 16465 790 16475 810
rect 16435 760 16475 790
rect 16435 740 16445 760
rect 16465 740 16475 760
rect 16435 725 16475 740
rect 16490 810 16530 825
rect 16490 790 16500 810
rect 16520 790 16530 810
rect 16490 760 16530 790
rect 16490 740 16500 760
rect 16520 740 16530 760
rect 16490 725 16530 740
rect 16545 810 16585 825
rect 16545 790 16555 810
rect 16575 790 16585 810
rect 16545 760 16585 790
rect 16545 740 16555 760
rect 16575 740 16585 760
rect 16545 725 16585 740
rect 16600 810 16640 825
rect 16600 790 16610 810
rect 16630 790 16640 810
rect 16600 760 16640 790
rect 16600 740 16610 760
rect 16630 740 16640 760
rect 16600 725 16640 740
rect 16655 810 16700 825
rect 16655 790 16665 810
rect 16685 790 16700 810
rect 16655 760 16700 790
rect 16655 740 16665 760
rect 16685 740 16700 760
rect 16655 725 16700 740
rect 16970 810 17010 840
rect 16970 790 16980 810
rect 17000 790 17010 810
rect 16970 760 17010 790
rect 16970 740 16980 760
rect 17000 740 17010 760
rect 16970 710 17010 740
rect 16970 690 16980 710
rect 17000 690 17010 710
rect 16970 660 17010 690
rect 16970 640 16980 660
rect 17000 640 17010 660
rect 16970 625 17010 640
rect 17060 910 17100 925
rect 17060 890 17070 910
rect 17090 890 17100 910
rect 17060 860 17100 890
rect 17060 840 17070 860
rect 17090 840 17100 860
rect 17060 810 17100 840
rect 17060 790 17070 810
rect 17090 790 17100 810
rect 17060 760 17100 790
rect 17060 740 17070 760
rect 17090 740 17100 760
rect 17060 710 17100 740
rect 17060 690 17070 710
rect 17090 690 17100 710
rect 17060 660 17100 690
rect 17060 640 17070 660
rect 17090 640 17100 660
rect 17060 625 17100 640
rect 17150 910 17190 925
rect 17150 890 17160 910
rect 17180 890 17190 910
rect 17150 860 17190 890
rect 17150 840 17160 860
rect 17180 840 17190 860
rect 17150 810 17190 840
rect 17150 790 17160 810
rect 17180 790 17190 810
rect 17150 760 17190 790
rect 17150 740 17160 760
rect 17180 740 17190 760
rect 17150 710 17190 740
rect 17150 690 17160 710
rect 17180 690 17190 710
rect 17150 660 17190 690
rect 17150 640 17160 660
rect 17180 640 17190 660
rect 17150 625 17190 640
rect 17240 910 17280 925
rect 17240 890 17250 910
rect 17270 890 17280 910
rect 17240 860 17280 890
rect 17240 840 17250 860
rect 17270 840 17280 860
rect 17240 810 17280 840
rect 17240 790 17250 810
rect 17270 790 17280 810
rect 17240 760 17280 790
rect 17240 740 17250 760
rect 17270 740 17280 760
rect 17240 710 17280 740
rect 17240 690 17250 710
rect 17270 690 17280 710
rect 17240 660 17280 690
rect 17240 640 17250 660
rect 17270 640 17280 660
rect 17240 625 17280 640
rect 17330 910 17370 925
rect 17330 890 17340 910
rect 17360 890 17370 910
rect 17330 860 17370 890
rect 17330 840 17340 860
rect 17360 840 17370 860
rect 17330 810 17370 840
rect 17330 790 17340 810
rect 17360 790 17370 810
rect 17330 760 17370 790
rect 17330 740 17340 760
rect 17360 740 17370 760
rect 17330 710 17370 740
rect 17330 690 17340 710
rect 17360 690 17370 710
rect 17330 660 17370 690
rect 17330 640 17340 660
rect 17360 640 17370 660
rect 17330 625 17370 640
rect 17420 910 17460 925
rect 17420 890 17430 910
rect 17450 890 17460 910
rect 17420 860 17460 890
rect 17420 840 17430 860
rect 17450 840 17460 860
rect 17420 810 17460 840
rect 17420 790 17430 810
rect 17450 790 17460 810
rect 17420 760 17460 790
rect 17420 740 17430 760
rect 17450 740 17460 760
rect 17420 710 17460 740
rect 17420 690 17430 710
rect 17450 690 17460 710
rect 17420 660 17460 690
rect 17420 640 17430 660
rect 17450 640 17460 660
rect 17420 625 17460 640
rect 17510 910 17550 925
rect 17510 890 17520 910
rect 17540 890 17550 910
rect 17510 860 17550 890
rect 17510 840 17520 860
rect 17540 840 17550 860
rect 17510 810 17550 840
rect 17510 790 17520 810
rect 17540 790 17550 810
rect 17510 760 17550 790
rect 17510 740 17520 760
rect 17540 740 17550 760
rect 17510 710 17550 740
rect 17510 690 17520 710
rect 17540 690 17550 710
rect 17510 660 17550 690
rect 17510 640 17520 660
rect 17540 640 17550 660
rect 17510 625 17550 640
rect 17600 910 17640 925
rect 17600 890 17610 910
rect 17630 890 17640 910
rect 17600 860 17640 890
rect 17600 840 17610 860
rect 17630 840 17640 860
rect 17600 810 17640 840
rect 17600 790 17610 810
rect 17630 790 17640 810
rect 17600 760 17640 790
rect 17600 740 17610 760
rect 17630 740 17640 760
rect 17600 710 17640 740
rect 17600 690 17610 710
rect 17630 690 17640 710
rect 17600 660 17640 690
rect 17600 640 17610 660
rect 17630 640 17640 660
rect 17600 625 17640 640
rect 17690 910 17730 925
rect 17690 890 17700 910
rect 17720 890 17730 910
rect 17690 860 17730 890
rect 17690 840 17700 860
rect 17720 840 17730 860
rect 17690 810 17730 840
rect 17690 790 17700 810
rect 17720 790 17730 810
rect 17690 760 17730 790
rect 17690 740 17700 760
rect 17720 740 17730 760
rect 17690 710 17730 740
rect 17690 690 17700 710
rect 17720 690 17730 710
rect 17690 660 17730 690
rect 17690 640 17700 660
rect 17720 640 17730 660
rect 17690 625 17730 640
rect 17780 910 17820 925
rect 17780 890 17790 910
rect 17810 890 17820 910
rect 17780 860 17820 890
rect 17780 840 17790 860
rect 17810 840 17820 860
rect 17780 810 17820 840
rect 17780 790 17790 810
rect 17810 790 17820 810
rect 17780 760 17820 790
rect 17780 740 17790 760
rect 17810 740 17820 760
rect 17780 710 17820 740
rect 17780 690 17790 710
rect 17810 690 17820 710
rect 17780 660 17820 690
rect 17780 640 17790 660
rect 17810 640 17820 660
rect 17780 625 17820 640
rect 17870 910 17910 925
rect 17870 890 17880 910
rect 17900 890 17910 910
rect 17870 860 17910 890
rect 17870 840 17880 860
rect 17900 840 17910 860
rect 17870 810 17910 840
rect 17870 790 17880 810
rect 17900 790 17910 810
rect 17870 760 17910 790
rect 17870 740 17880 760
rect 17900 740 17910 760
rect 17870 710 17910 740
rect 17870 690 17880 710
rect 17900 690 17910 710
rect 17870 660 17910 690
rect 17870 640 17880 660
rect 17900 640 17910 660
rect 17870 625 17910 640
rect 17960 910 18000 925
rect 17960 890 17970 910
rect 17990 890 18000 910
rect 17960 860 18000 890
rect 17960 840 17970 860
rect 17990 840 18000 860
rect 17960 810 18000 840
rect 17960 790 17970 810
rect 17990 790 18000 810
rect 17960 760 18000 790
rect 17960 740 17970 760
rect 17990 740 18000 760
rect 17960 710 18000 740
rect 17960 690 17970 710
rect 17990 690 18000 710
rect 17960 660 18000 690
rect 17960 640 17970 660
rect 17990 640 18000 660
rect 17960 625 18000 640
rect 18050 910 18090 925
rect 18050 890 18060 910
rect 18080 890 18090 910
rect 18050 860 18090 890
rect 18050 840 18060 860
rect 18080 840 18090 860
rect 18050 810 18090 840
rect 18050 790 18060 810
rect 18080 790 18090 810
rect 18050 760 18090 790
rect 18050 740 18060 760
rect 18080 740 18090 760
rect 18050 710 18090 740
rect 18050 690 18060 710
rect 18080 690 18090 710
rect 18050 660 18090 690
rect 18050 640 18060 660
rect 18080 640 18090 660
rect 18050 625 18090 640
rect 18140 910 18180 925
rect 18140 890 18150 910
rect 18170 890 18180 910
rect 18140 860 18180 890
rect 18140 840 18150 860
rect 18170 840 18180 860
rect 18140 810 18180 840
rect 18140 790 18150 810
rect 18170 790 18180 810
rect 18140 760 18180 790
rect 18140 740 18150 760
rect 18170 740 18180 760
rect 18140 710 18180 740
rect 18140 690 18150 710
rect 18170 690 18180 710
rect 18140 660 18180 690
rect 18140 640 18150 660
rect 18170 640 18180 660
rect 18140 625 18180 640
rect 18230 910 18270 925
rect 18230 890 18240 910
rect 18260 890 18270 910
rect 18230 860 18270 890
rect 18230 840 18240 860
rect 18260 840 18270 860
rect 18230 810 18270 840
rect 18230 790 18240 810
rect 18260 790 18270 810
rect 18230 760 18270 790
rect 18230 740 18240 760
rect 18260 740 18270 760
rect 18230 710 18270 740
rect 18230 690 18240 710
rect 18260 690 18270 710
rect 18230 660 18270 690
rect 18230 640 18240 660
rect 18260 640 18270 660
rect 18230 625 18270 640
rect 18320 910 18360 925
rect 18320 890 18330 910
rect 18350 890 18360 910
rect 18320 860 18360 890
rect 18320 840 18330 860
rect 18350 840 18360 860
rect 18320 810 18360 840
rect 18320 790 18330 810
rect 18350 790 18360 810
rect 18320 760 18360 790
rect 18320 740 18330 760
rect 18350 740 18360 760
rect 18320 710 18360 740
rect 18320 690 18330 710
rect 18350 690 18360 710
rect 18320 660 18360 690
rect 18320 640 18330 660
rect 18350 640 18360 660
rect 18320 625 18360 640
rect 18410 910 18450 925
rect 18410 890 18420 910
rect 18440 890 18450 910
rect 18410 860 18450 890
rect 18410 840 18420 860
rect 18440 840 18450 860
rect 18410 810 18450 840
rect 18410 790 18420 810
rect 18440 790 18450 810
rect 18410 760 18450 790
rect 18410 740 18420 760
rect 18440 740 18450 760
rect 18410 710 18450 740
rect 18410 690 18420 710
rect 18440 690 18450 710
rect 18410 660 18450 690
rect 18410 640 18420 660
rect 18440 640 18450 660
rect 18410 625 18450 640
rect 18500 910 18540 925
rect 18500 890 18510 910
rect 18530 890 18540 910
rect 18500 860 18540 890
rect 18500 840 18510 860
rect 18530 840 18540 860
rect 18500 810 18540 840
rect 18500 790 18510 810
rect 18530 790 18540 810
rect 18500 760 18540 790
rect 18500 740 18510 760
rect 18530 740 18540 760
rect 18500 710 18540 740
rect 18500 690 18510 710
rect 18530 690 18540 710
rect 18500 660 18540 690
rect 18500 640 18510 660
rect 18530 640 18540 660
rect 18500 625 18540 640
rect 18590 910 18630 925
rect 18590 890 18600 910
rect 18620 890 18630 910
rect 18590 860 18630 890
rect 18590 840 18600 860
rect 18620 840 18630 860
rect 18590 810 18630 840
rect 18590 790 18600 810
rect 18620 790 18630 810
rect 18590 760 18630 790
rect 18590 740 18600 760
rect 18620 740 18630 760
rect 18590 710 18630 740
rect 18905 910 18945 925
rect 18905 890 18915 910
rect 18935 890 18945 910
rect 18905 860 18945 890
rect 18905 840 18915 860
rect 18935 840 18945 860
rect 18905 810 18945 840
rect 18905 790 18915 810
rect 18935 790 18945 810
rect 18905 760 18945 790
rect 18905 740 18915 760
rect 18935 740 18945 760
rect 18905 725 18945 740
rect 18960 910 19000 925
rect 18960 890 18970 910
rect 18990 890 19000 910
rect 18960 860 19000 890
rect 18960 840 18970 860
rect 18990 840 19000 860
rect 18960 810 19000 840
rect 18960 790 18970 810
rect 18990 790 19000 810
rect 18960 760 19000 790
rect 18960 740 18970 760
rect 18990 740 19000 760
rect 18960 725 19000 740
rect 19015 910 19055 925
rect 19015 890 19025 910
rect 19045 890 19055 910
rect 19015 860 19055 890
rect 19015 840 19025 860
rect 19045 840 19055 860
rect 19015 810 19055 840
rect 19015 790 19025 810
rect 19045 790 19055 810
rect 19015 760 19055 790
rect 19015 740 19025 760
rect 19045 740 19055 760
rect 19015 725 19055 740
rect 19070 910 19110 925
rect 19070 890 19080 910
rect 19100 890 19110 910
rect 19070 860 19110 890
rect 19070 840 19080 860
rect 19100 840 19110 860
rect 19070 810 19110 840
rect 19070 790 19080 810
rect 19100 790 19110 810
rect 19070 760 19110 790
rect 19070 740 19080 760
rect 19100 740 19110 760
rect 19070 725 19110 740
rect 18590 690 18600 710
rect 18620 690 18630 710
rect 18590 660 18630 690
rect 18590 640 18600 660
rect 18620 640 18630 660
rect 18590 625 18630 640
rect 16420 70 16460 85
rect 16420 50 16430 70
rect 16450 50 16460 70
rect 16420 20 16460 50
rect 16420 0 16430 20
rect 16450 0 16460 20
rect 16420 -15 16460 0
rect 16480 70 16520 85
rect 16480 50 16490 70
rect 16510 50 16520 70
rect 16480 20 16520 50
rect 16480 0 16490 20
rect 16510 0 16520 20
rect 16480 -15 16520 0
rect 16540 70 16580 85
rect 16540 50 16550 70
rect 16570 50 16580 70
rect 16540 20 16580 50
rect 16540 0 16550 20
rect 16570 0 16580 20
rect 16540 -15 16580 0
rect 16600 70 16640 85
rect 16600 50 16610 70
rect 16630 50 16640 70
rect 16600 20 16640 50
rect 16600 0 16610 20
rect 16630 0 16640 20
rect 16600 -15 16640 0
rect 16660 70 16700 85
rect 16660 50 16670 70
rect 16690 50 16700 70
rect 16660 20 16700 50
rect 16660 0 16670 20
rect 16690 0 16700 20
rect 16660 -15 16700 0
rect 16720 70 16760 85
rect 16720 50 16730 70
rect 16750 50 16760 70
rect 16720 20 16760 50
rect 16720 0 16730 20
rect 16750 0 16760 20
rect 16720 -15 16760 0
rect 16780 70 16820 85
rect 16780 50 16790 70
rect 16810 50 16820 70
rect 16780 20 16820 50
rect 16780 0 16790 20
rect 16810 0 16820 20
rect 16780 -15 16820 0
rect 16840 70 16880 85
rect 16840 50 16850 70
rect 16870 50 16880 70
rect 16840 20 16880 50
rect 16840 0 16850 20
rect 16870 0 16880 20
rect 16840 -15 16880 0
rect 16900 70 16940 85
rect 16900 50 16910 70
rect 16930 50 16940 70
rect 16900 20 16940 50
rect 16900 0 16910 20
rect 16930 0 16940 20
rect 16900 -15 16940 0
rect 16960 70 17000 85
rect 16960 50 16970 70
rect 16990 50 17000 70
rect 16960 20 17000 50
rect 16960 0 16970 20
rect 16990 0 17000 20
rect 16960 -15 17000 0
rect 17020 70 17060 85
rect 17020 50 17030 70
rect 17050 50 17060 70
rect 17020 20 17060 50
rect 17020 0 17030 20
rect 17050 0 17060 20
rect 17020 -15 17060 0
rect 17080 70 17120 85
rect 17080 50 17090 70
rect 17110 50 17120 70
rect 17080 20 17120 50
rect 17080 0 17090 20
rect 17110 0 17120 20
rect 17080 -15 17120 0
rect 17140 70 17180 85
rect 17140 50 17150 70
rect 17170 50 17180 70
rect 17140 20 17180 50
rect 17140 0 17150 20
rect 17170 0 17180 20
rect 17140 -15 17180 0
rect 17200 70 17240 85
rect 17200 50 17210 70
rect 17230 50 17240 70
rect 17200 20 17240 50
rect 17200 0 17210 20
rect 17230 0 17240 20
rect 17200 -15 17240 0
rect 17260 70 17300 85
rect 17260 50 17270 70
rect 17290 50 17300 70
rect 17260 20 17300 50
rect 17260 0 17270 20
rect 17290 0 17300 20
rect 17260 -15 17300 0
rect 17320 70 17360 85
rect 17320 50 17330 70
rect 17350 50 17360 70
rect 17320 20 17360 50
rect 17320 0 17330 20
rect 17350 0 17360 20
rect 17320 -15 17360 0
rect 17380 70 17420 85
rect 17380 50 17390 70
rect 17410 50 17420 70
rect 17380 20 17420 50
rect 17380 0 17390 20
rect 17410 0 17420 20
rect 17380 -15 17420 0
rect 17440 70 17480 85
rect 17440 50 17450 70
rect 17470 50 17480 70
rect 17440 20 17480 50
rect 17440 0 17450 20
rect 17470 0 17480 20
rect 17440 -15 17480 0
rect 17500 70 17540 85
rect 17500 50 17510 70
rect 17530 50 17540 70
rect 17500 20 17540 50
rect 17500 0 17510 20
rect 17530 0 17540 20
rect 17500 -15 17540 0
rect 17560 70 17600 85
rect 17560 50 17570 70
rect 17590 50 17600 70
rect 17560 20 17600 50
rect 17560 0 17570 20
rect 17590 0 17600 20
rect 17560 -15 17600 0
rect 17620 70 17660 85
rect 17620 50 17630 70
rect 17650 50 17660 70
rect 17620 20 17660 50
rect 17620 0 17630 20
rect 17650 0 17660 20
rect 17620 -15 17660 0
rect 17940 70 17980 85
rect 17940 50 17950 70
rect 17970 50 17980 70
rect 17940 20 17980 50
rect 17940 0 17950 20
rect 17970 0 17980 20
rect 17940 -15 17980 0
rect 18000 70 18040 85
rect 18000 50 18010 70
rect 18030 50 18040 70
rect 18000 20 18040 50
rect 18000 0 18010 20
rect 18030 0 18040 20
rect 18000 -15 18040 0
rect 18060 70 18100 85
rect 18060 50 18070 70
rect 18090 50 18100 70
rect 18060 20 18100 50
rect 18060 0 18070 20
rect 18090 0 18100 20
rect 18060 -15 18100 0
rect 18120 70 18160 85
rect 18120 50 18130 70
rect 18150 50 18160 70
rect 18120 20 18160 50
rect 18120 0 18130 20
rect 18150 0 18160 20
rect 18120 -15 18160 0
rect 18180 70 18220 85
rect 18180 50 18190 70
rect 18210 50 18220 70
rect 18180 20 18220 50
rect 18180 0 18190 20
rect 18210 0 18220 20
rect 18180 -15 18220 0
rect 18240 70 18280 85
rect 18240 50 18250 70
rect 18270 50 18280 70
rect 18240 20 18280 50
rect 18240 0 18250 20
rect 18270 0 18280 20
rect 18240 -15 18280 0
rect 18300 70 18340 85
rect 18300 50 18310 70
rect 18330 50 18340 70
rect 18300 20 18340 50
rect 18300 0 18310 20
rect 18330 0 18340 20
rect 18300 -15 18340 0
rect 18360 70 18400 85
rect 18360 50 18370 70
rect 18390 50 18400 70
rect 18360 20 18400 50
rect 18360 0 18370 20
rect 18390 0 18400 20
rect 18360 -15 18400 0
rect 18420 70 18460 85
rect 18420 50 18430 70
rect 18450 50 18460 70
rect 18420 20 18460 50
rect 18420 0 18430 20
rect 18450 0 18460 20
rect 18420 -15 18460 0
rect 18480 70 18520 85
rect 18480 50 18490 70
rect 18510 50 18520 70
rect 18480 20 18520 50
rect 18480 0 18490 20
rect 18510 0 18520 20
rect 18480 -15 18520 0
rect 18540 70 18580 85
rect 18540 50 18550 70
rect 18570 50 18580 70
rect 18540 20 18580 50
rect 18540 0 18550 20
rect 18570 0 18580 20
rect 18540 -15 18580 0
rect 18600 70 18640 85
rect 18600 50 18610 70
rect 18630 50 18640 70
rect 18600 20 18640 50
rect 18600 0 18610 20
rect 18630 0 18640 20
rect 18600 -15 18640 0
rect 18660 70 18700 85
rect 18660 50 18670 70
rect 18690 50 18700 70
rect 18660 20 18700 50
rect 18660 0 18670 20
rect 18690 0 18700 20
rect 18660 -15 18700 0
rect 18720 70 18760 85
rect 18720 50 18730 70
rect 18750 50 18760 70
rect 18720 20 18760 50
rect 18720 0 18730 20
rect 18750 0 18760 20
rect 18720 -15 18760 0
rect 18780 70 18820 85
rect 18780 50 18790 70
rect 18810 50 18820 70
rect 18780 20 18820 50
rect 18780 0 18790 20
rect 18810 0 18820 20
rect 18780 -15 18820 0
rect 18840 70 18880 85
rect 18840 50 18850 70
rect 18870 50 18880 70
rect 18840 20 18880 50
rect 18840 0 18850 20
rect 18870 0 18880 20
rect 18840 -15 18880 0
rect 18900 70 18940 85
rect 18900 50 18910 70
rect 18930 50 18940 70
rect 18900 20 18940 50
rect 18900 0 18910 20
rect 18930 0 18940 20
rect 18900 -15 18940 0
rect 18960 70 19000 85
rect 18960 50 18970 70
rect 18990 50 19000 70
rect 18960 20 19000 50
rect 18960 0 18970 20
rect 18990 0 19000 20
rect 18960 -15 19000 0
rect 19020 70 19060 85
rect 19020 50 19030 70
rect 19050 50 19060 70
rect 19020 20 19060 50
rect 19020 0 19030 20
rect 19050 0 19060 20
rect 19020 -15 19060 0
rect 19080 70 19120 85
rect 19080 50 19090 70
rect 19110 50 19120 70
rect 19080 20 19120 50
rect 19080 0 19090 20
rect 19110 0 19120 20
rect 19080 -15 19120 0
rect 19140 70 19180 85
rect 19140 50 19150 70
rect 19170 50 19180 70
rect 19140 20 19180 50
rect 19140 0 19150 20
rect 19170 0 19180 20
rect 19140 -15 19180 0
<< ndiffc >>
rect 16970 -235 16990 -215
rect 16970 -285 16990 -265
rect 16970 -335 16990 -315
rect 16970 -385 16990 -365
rect 16970 -435 16990 -415
rect 17030 -235 17050 -215
rect 17030 -285 17050 -265
rect 17030 -335 17050 -315
rect 17030 -385 17050 -365
rect 17030 -435 17050 -415
rect 17090 -235 17110 -215
rect 17090 -285 17110 -265
rect 17090 -335 17110 -315
rect 18490 -235 18510 -215
rect 18490 -285 18510 -265
rect 17090 -385 17110 -365
rect 17090 -435 17110 -415
rect 18490 -335 18510 -315
rect 18490 -385 18510 -365
rect 18490 -435 18510 -415
rect 18550 -235 18570 -215
rect 18550 -285 18570 -265
rect 18550 -335 18570 -315
rect 18550 -385 18570 -365
rect 18550 -435 18570 -415
rect 18610 -235 18630 -215
rect 18610 -285 18630 -265
rect 18610 -335 18630 -315
rect 18610 -385 18630 -365
rect 18610 -435 18630 -415
rect 16540 -770 16560 -750
rect 16540 -820 16560 -800
rect 16540 -870 16560 -850
rect 16540 -920 16560 -900
rect 16540 -970 16560 -950
rect 17080 -770 17100 -750
rect 17160 -770 17180 -750
rect 17080 -820 17100 -800
rect 17160 -820 17180 -800
rect 17080 -870 17100 -850
rect 17160 -870 17180 -850
rect 17080 -920 17100 -900
rect 17160 -920 17180 -900
rect 17080 -970 17100 -950
rect 17160 -970 17180 -950
rect 17700 -770 17720 -750
rect 17700 -820 17720 -800
rect 17700 -870 17720 -850
rect 17700 -920 17720 -900
rect 17700 -970 17720 -950
rect 17880 -770 17900 -750
rect 17880 -820 17900 -800
rect 17880 -870 17900 -850
rect 17880 -920 17900 -900
rect 17880 -970 17900 -950
rect 18420 -770 18440 -750
rect 18500 -770 18520 -750
rect 18420 -820 18440 -800
rect 18500 -820 18520 -800
rect 18420 -870 18440 -850
rect 18500 -870 18520 -850
rect 18420 -920 18440 -900
rect 18500 -920 18520 -900
rect 18420 -970 18440 -950
rect 18500 -970 18520 -950
rect 19040 -770 19060 -750
rect 19040 -820 19060 -800
rect 19040 -870 19060 -850
rect 19040 -920 19060 -900
rect 19040 -970 19060 -950
rect 16750 -1225 16770 -1205
rect 16750 -1275 16770 -1255
rect 17790 -1225 17810 -1205
rect 17790 -1275 17810 -1255
rect 18830 -1225 18850 -1205
rect 18830 -1275 18850 -1255
rect 16550 -1575 16570 -1555
rect 16550 -1625 16570 -1605
rect 16605 -1575 16625 -1555
rect 16605 -1625 16625 -1605
rect 16660 -1575 16680 -1555
rect 16660 -1625 16680 -1605
rect 16715 -1575 16735 -1555
rect 16715 -1625 16735 -1605
rect 16770 -1575 16790 -1555
rect 16770 -1625 16790 -1605
rect 16825 -1575 16845 -1555
rect 16825 -1625 16845 -1605
rect 17035 -1575 17055 -1555
rect 17035 -1625 17055 -1605
rect 17090 -1575 17110 -1555
rect 17090 -1625 17110 -1605
rect 17145 -1575 17165 -1555
rect 17145 -1625 17165 -1605
rect 17200 -1575 17220 -1555
rect 17200 -1625 17220 -1605
rect 17255 -1575 17275 -1555
rect 17255 -1625 17275 -1605
rect 17310 -1575 17330 -1555
rect 17310 -1625 17330 -1605
rect 17365 -1575 17385 -1555
rect 17365 -1625 17385 -1605
rect 17420 -1575 17440 -1555
rect 17420 -1625 17440 -1605
rect 17475 -1575 17495 -1555
rect 17475 -1625 17495 -1605
rect 17625 -1575 17645 -1555
rect 17625 -1625 17645 -1605
rect 17680 -1575 17700 -1555
rect 17680 -1625 17700 -1605
rect 17735 -1575 17755 -1555
rect 17735 -1625 17755 -1605
rect 17790 -1575 17810 -1555
rect 17790 -1625 17810 -1605
rect 17845 -1575 17865 -1555
rect 17845 -1625 17865 -1605
rect 17900 -1575 17920 -1555
rect 17900 -1625 17920 -1605
rect 17955 -1575 17975 -1555
rect 17955 -1625 17975 -1605
rect 18105 -1575 18125 -1555
rect 18105 -1625 18125 -1605
rect 18160 -1575 18180 -1555
rect 18160 -1625 18180 -1605
rect 18215 -1575 18235 -1555
rect 18215 -1625 18235 -1605
rect 18270 -1575 18290 -1555
rect 18270 -1625 18290 -1605
rect 18325 -1575 18345 -1555
rect 18325 -1625 18345 -1605
rect 18380 -1575 18400 -1555
rect 18380 -1625 18400 -1605
rect 18435 -1575 18455 -1555
rect 18435 -1625 18455 -1605
rect 18490 -1575 18510 -1555
rect 18490 -1625 18510 -1605
rect 18545 -1575 18565 -1555
rect 18545 -1625 18565 -1605
<< pdiffc >>
rect 16385 1355 16405 1375
rect 16385 1305 16405 1325
rect 16440 1355 16460 1375
rect 16440 1305 16460 1325
rect 16495 1355 16515 1375
rect 16495 1305 16515 1325
rect 16550 1355 16570 1375
rect 16550 1305 16570 1325
rect 16605 1355 16625 1375
rect 16605 1305 16625 1325
rect 16895 1303 16915 1375
rect 16950 1303 16970 1375
rect 17005 1303 17025 1375
rect 17060 1303 17080 1375
rect 17115 1303 17135 1375
rect 17170 1303 17190 1375
rect 17225 1303 17245 1375
rect 17515 1355 17535 1375
rect 17515 1305 17535 1325
rect 17570 1355 17590 1375
rect 17570 1305 17590 1325
rect 17625 1355 17645 1375
rect 17625 1305 17645 1325
rect 17680 1355 17700 1375
rect 17680 1305 17700 1325
rect 17735 1355 17755 1375
rect 17735 1305 17755 1325
rect 17790 1355 17810 1375
rect 17790 1305 17810 1325
rect 17845 1355 17865 1375
rect 17845 1305 17865 1325
rect 17900 1355 17920 1375
rect 17900 1305 17920 1325
rect 17955 1355 17975 1375
rect 17955 1305 17975 1325
rect 18010 1355 18030 1375
rect 18010 1305 18030 1325
rect 18065 1355 18085 1375
rect 18065 1305 18085 1325
rect 18355 1305 18375 1375
rect 18410 1305 18430 1375
rect 18465 1305 18485 1375
rect 18520 1305 18540 1375
rect 18575 1305 18595 1375
rect 18630 1305 18650 1375
rect 18685 1305 18705 1375
rect 16980 890 17000 910
rect 16980 840 17000 860
rect 16445 790 16465 810
rect 16445 740 16465 760
rect 16500 790 16520 810
rect 16500 740 16520 760
rect 16555 790 16575 810
rect 16555 740 16575 760
rect 16610 790 16630 810
rect 16610 740 16630 760
rect 16665 790 16685 810
rect 16665 740 16685 760
rect 16980 790 17000 810
rect 16980 740 17000 760
rect 16980 690 17000 710
rect 16980 640 17000 660
rect 17070 890 17090 910
rect 17070 840 17090 860
rect 17070 790 17090 810
rect 17070 740 17090 760
rect 17070 690 17090 710
rect 17070 640 17090 660
rect 17160 890 17180 910
rect 17160 840 17180 860
rect 17160 790 17180 810
rect 17160 740 17180 760
rect 17160 690 17180 710
rect 17160 640 17180 660
rect 17250 890 17270 910
rect 17250 840 17270 860
rect 17250 790 17270 810
rect 17250 740 17270 760
rect 17250 690 17270 710
rect 17250 640 17270 660
rect 17340 890 17360 910
rect 17340 840 17360 860
rect 17340 790 17360 810
rect 17340 740 17360 760
rect 17340 690 17360 710
rect 17340 640 17360 660
rect 17430 890 17450 910
rect 17430 840 17450 860
rect 17430 790 17450 810
rect 17430 740 17450 760
rect 17430 690 17450 710
rect 17430 640 17450 660
rect 17520 890 17540 910
rect 17520 840 17540 860
rect 17520 790 17540 810
rect 17520 740 17540 760
rect 17520 690 17540 710
rect 17520 640 17540 660
rect 17610 890 17630 910
rect 17610 840 17630 860
rect 17610 790 17630 810
rect 17610 740 17630 760
rect 17610 690 17630 710
rect 17610 640 17630 660
rect 17700 890 17720 910
rect 17700 840 17720 860
rect 17700 790 17720 810
rect 17700 740 17720 760
rect 17700 690 17720 710
rect 17700 640 17720 660
rect 17790 890 17810 910
rect 17790 840 17810 860
rect 17790 790 17810 810
rect 17790 740 17810 760
rect 17790 690 17810 710
rect 17790 640 17810 660
rect 17880 890 17900 910
rect 17880 840 17900 860
rect 17880 790 17900 810
rect 17880 740 17900 760
rect 17880 690 17900 710
rect 17880 640 17900 660
rect 17970 890 17990 910
rect 17970 840 17990 860
rect 17970 790 17990 810
rect 17970 740 17990 760
rect 17970 690 17990 710
rect 17970 640 17990 660
rect 18060 890 18080 910
rect 18060 840 18080 860
rect 18060 790 18080 810
rect 18060 740 18080 760
rect 18060 690 18080 710
rect 18060 640 18080 660
rect 18150 890 18170 910
rect 18150 840 18170 860
rect 18150 790 18170 810
rect 18150 740 18170 760
rect 18150 690 18170 710
rect 18150 640 18170 660
rect 18240 890 18260 910
rect 18240 840 18260 860
rect 18240 790 18260 810
rect 18240 740 18260 760
rect 18240 690 18260 710
rect 18240 640 18260 660
rect 18330 890 18350 910
rect 18330 840 18350 860
rect 18330 790 18350 810
rect 18330 740 18350 760
rect 18330 690 18350 710
rect 18330 640 18350 660
rect 18420 890 18440 910
rect 18420 840 18440 860
rect 18420 790 18440 810
rect 18420 740 18440 760
rect 18420 690 18440 710
rect 18420 640 18440 660
rect 18510 890 18530 910
rect 18510 840 18530 860
rect 18510 790 18530 810
rect 18510 740 18530 760
rect 18510 690 18530 710
rect 18510 640 18530 660
rect 18600 890 18620 910
rect 18600 840 18620 860
rect 18600 790 18620 810
rect 18600 740 18620 760
rect 18915 890 18935 910
rect 18915 840 18935 860
rect 18915 790 18935 810
rect 18915 740 18935 760
rect 18970 890 18990 910
rect 18970 840 18990 860
rect 18970 790 18990 810
rect 18970 740 18990 760
rect 19025 890 19045 910
rect 19025 840 19045 860
rect 19025 790 19045 810
rect 19025 740 19045 760
rect 19080 890 19100 910
rect 19080 840 19100 860
rect 19080 790 19100 810
rect 19080 740 19100 760
rect 18600 690 18620 710
rect 18600 640 18620 660
rect 16430 50 16450 70
rect 16430 0 16450 20
rect 16490 50 16510 70
rect 16490 0 16510 20
rect 16550 50 16570 70
rect 16550 0 16570 20
rect 16610 50 16630 70
rect 16610 0 16630 20
rect 16670 50 16690 70
rect 16670 0 16690 20
rect 16730 50 16750 70
rect 16730 0 16750 20
rect 16790 50 16810 70
rect 16790 0 16810 20
rect 16850 50 16870 70
rect 16850 0 16870 20
rect 16910 50 16930 70
rect 16910 0 16930 20
rect 16970 50 16990 70
rect 16970 0 16990 20
rect 17030 50 17050 70
rect 17030 0 17050 20
rect 17090 50 17110 70
rect 17090 0 17110 20
rect 17150 50 17170 70
rect 17150 0 17170 20
rect 17210 50 17230 70
rect 17210 0 17230 20
rect 17270 50 17290 70
rect 17270 0 17290 20
rect 17330 50 17350 70
rect 17330 0 17350 20
rect 17390 50 17410 70
rect 17390 0 17410 20
rect 17450 50 17470 70
rect 17450 0 17470 20
rect 17510 50 17530 70
rect 17510 0 17530 20
rect 17570 50 17590 70
rect 17570 0 17590 20
rect 17630 50 17650 70
rect 17630 0 17650 20
rect 17950 50 17970 70
rect 17950 0 17970 20
rect 18010 50 18030 70
rect 18010 0 18030 20
rect 18070 50 18090 70
rect 18070 0 18090 20
rect 18130 50 18150 70
rect 18130 0 18150 20
rect 18190 50 18210 70
rect 18190 0 18210 20
rect 18250 50 18270 70
rect 18250 0 18270 20
rect 18310 50 18330 70
rect 18310 0 18330 20
rect 18370 50 18390 70
rect 18370 0 18390 20
rect 18430 50 18450 70
rect 18430 0 18450 20
rect 18490 50 18510 70
rect 18490 0 18510 20
rect 18550 50 18570 70
rect 18550 0 18570 20
rect 18610 50 18630 70
rect 18610 0 18630 20
rect 18670 50 18690 70
rect 18670 0 18690 20
rect 18730 50 18750 70
rect 18730 0 18750 20
rect 18790 50 18810 70
rect 18790 0 18810 20
rect 18850 50 18870 70
rect 18850 0 18870 20
rect 18910 50 18930 70
rect 18910 0 18930 20
rect 18970 50 18990 70
rect 18970 0 18990 20
rect 19030 50 19050 70
rect 19030 0 19050 20
rect 19090 50 19110 70
rect 19090 0 19110 20
rect 19150 50 19170 70
rect 19150 0 19170 20
<< psubdiff >>
rect 17560 -215 17600 -200
rect 17560 -235 17570 -215
rect 17590 -235 17600 -215
rect 17560 -255 17600 -235
rect 17560 -275 17570 -255
rect 17590 -275 17600 -255
rect 17560 -295 17600 -275
rect 17560 -315 17570 -295
rect 17590 -315 17600 -295
rect 17560 -330 17600 -315
rect 18000 -215 18040 -200
rect 18000 -235 18010 -215
rect 18030 -235 18040 -215
rect 18000 -255 18040 -235
rect 18000 -275 18010 -255
rect 18030 -275 18040 -255
rect 18000 -295 18040 -275
rect 18000 -315 18010 -295
rect 18030 -315 18040 -295
rect 18000 -330 18040 -315
rect 17110 -750 17150 -735
rect 17110 -770 17120 -750
rect 17140 -770 17150 -750
rect 17110 -800 17150 -770
rect 17110 -820 17120 -800
rect 17140 -820 17150 -800
rect 17110 -850 17150 -820
rect 17110 -870 17120 -850
rect 17140 -870 17150 -850
rect 17110 -900 17150 -870
rect 17110 -920 17120 -900
rect 17140 -920 17150 -900
rect 17110 -950 17150 -920
rect 17110 -970 17120 -950
rect 17140 -970 17150 -950
rect 17110 -980 17150 -970
rect 18450 -750 18490 -735
rect 18450 -770 18460 -750
rect 18480 -770 18490 -750
rect 18450 -800 18490 -770
rect 18450 -820 18460 -800
rect 18480 -820 18490 -800
rect 18450 -850 18490 -820
rect 18450 -870 18460 -850
rect 18480 -870 18490 -850
rect 18450 -900 18490 -870
rect 18450 -920 18460 -900
rect 18480 -920 18490 -900
rect 18450 -950 18490 -920
rect 18450 -970 18460 -950
rect 18480 -970 18490 -950
rect 18450 -985 18490 -970
rect 18860 -1205 18900 -1190
rect 18860 -1225 18870 -1205
rect 18890 -1225 18900 -1205
rect 18860 -1255 18900 -1225
rect 18860 -1275 18870 -1255
rect 18890 -1275 18900 -1255
rect 18860 -1290 18900 -1275
rect 16500 -1555 16540 -1540
rect 16500 -1575 16510 -1555
rect 16530 -1575 16540 -1555
rect 16500 -1605 16540 -1575
rect 16500 -1625 16510 -1605
rect 16530 -1625 16540 -1605
rect 16500 -1640 16540 -1625
rect 16855 -1555 16895 -1540
rect 16855 -1575 16865 -1555
rect 16885 -1575 16895 -1555
rect 16855 -1605 16895 -1575
rect 16855 -1625 16865 -1605
rect 16885 -1625 16895 -1605
rect 16855 -1640 16895 -1625
rect 16985 -1555 17025 -1540
rect 16985 -1575 16995 -1555
rect 17015 -1575 17025 -1555
rect 16985 -1605 17025 -1575
rect 16985 -1625 16995 -1605
rect 17015 -1625 17025 -1605
rect 16985 -1640 17025 -1625
rect 17505 -1555 17545 -1540
rect 17505 -1575 17515 -1555
rect 17535 -1575 17545 -1555
rect 17505 -1605 17545 -1575
rect 17505 -1625 17515 -1605
rect 17535 -1625 17545 -1605
rect 17505 -1640 17545 -1625
rect 17575 -1555 17615 -1540
rect 17575 -1575 17585 -1555
rect 17605 -1575 17615 -1555
rect 17575 -1605 17615 -1575
rect 17575 -1625 17585 -1605
rect 17605 -1625 17615 -1605
rect 17575 -1640 17615 -1625
rect 17985 -1555 18025 -1540
rect 17985 -1575 17995 -1555
rect 18015 -1575 18025 -1555
rect 17985 -1605 18025 -1575
rect 17985 -1625 17995 -1605
rect 18015 -1625 18025 -1605
rect 17985 -1640 18025 -1625
rect 18055 -1555 18095 -1540
rect 18055 -1575 18065 -1555
rect 18085 -1575 18095 -1555
rect 18055 -1605 18095 -1575
rect 18055 -1625 18065 -1605
rect 18085 -1625 18095 -1605
rect 18055 -1640 18095 -1625
rect 18575 -1555 18615 -1540
rect 18575 -1575 18585 -1555
rect 18605 -1575 18615 -1555
rect 18575 -1605 18615 -1575
rect 18575 -1625 18585 -1605
rect 18605 -1625 18615 -1605
rect 18575 -1640 18615 -1625
rect 17775 -4170 17825 -4155
rect 17775 -4190 17790 -4170
rect 17810 -4190 17825 -4170
rect 17775 -4220 17825 -4190
rect 17775 -4240 17790 -4220
rect 17810 -4240 17825 -4220
rect 17775 -4270 17825 -4240
rect 17775 -4290 17790 -4270
rect 17810 -4290 17825 -4270
rect 17775 -4305 17825 -4290
<< nsubdiff >>
rect 16335 1377 16375 1390
rect 16335 1355 16345 1377
rect 16365 1355 16375 1377
rect 16335 1325 16375 1355
rect 16335 1305 16345 1325
rect 16365 1305 16375 1325
rect 16335 1290 16375 1305
rect 16635 1377 16675 1390
rect 16635 1355 16645 1377
rect 16665 1355 16675 1377
rect 16635 1325 16675 1355
rect 16635 1305 16645 1325
rect 16665 1305 16675 1325
rect 16635 1290 16675 1305
rect 16845 1377 16885 1390
rect 16845 1305 16855 1377
rect 16875 1305 16885 1377
rect 16845 1290 16885 1305
rect 17255 1377 17295 1390
rect 17255 1305 17265 1377
rect 17285 1305 17295 1377
rect 17255 1290 17295 1305
rect 17465 1377 17505 1390
rect 17465 1355 17475 1377
rect 17495 1355 17505 1377
rect 17465 1325 17505 1355
rect 17465 1305 17475 1325
rect 17495 1305 17505 1325
rect 17465 1290 17505 1305
rect 18095 1377 18135 1390
rect 18095 1355 18105 1377
rect 18125 1355 18135 1377
rect 18095 1325 18135 1355
rect 18095 1305 18105 1325
rect 18125 1305 18135 1325
rect 18095 1290 18135 1305
rect 18305 1377 18345 1390
rect 18305 1305 18315 1377
rect 18335 1305 18345 1377
rect 18305 1290 18345 1305
rect 18715 1377 18755 1390
rect 18715 1305 18725 1377
rect 18745 1305 18755 1377
rect 18715 1290 18755 1305
rect 16930 910 16970 925
rect 16930 890 16940 910
rect 16960 890 16970 910
rect 16930 860 16970 890
rect 16930 840 16940 860
rect 16960 840 16970 860
rect 16395 810 16435 825
rect 16395 790 16405 810
rect 16425 790 16435 810
rect 16395 760 16435 790
rect 16395 740 16405 760
rect 16425 740 16435 760
rect 16395 725 16435 740
rect 16700 810 16740 825
rect 16700 790 16710 810
rect 16730 790 16740 810
rect 16700 760 16740 790
rect 16700 740 16710 760
rect 16730 740 16740 760
rect 16700 725 16740 740
rect 16930 810 16970 840
rect 16930 790 16940 810
rect 16960 790 16970 810
rect 16930 760 16970 790
rect 16930 740 16940 760
rect 16960 740 16970 760
rect 16930 710 16970 740
rect 16930 690 16940 710
rect 16960 690 16970 710
rect 16930 660 16970 690
rect 16930 640 16940 660
rect 16960 640 16970 660
rect 16930 625 16970 640
rect 18630 910 18670 925
rect 18630 890 18640 910
rect 18660 890 18670 910
rect 18630 860 18670 890
rect 18630 840 18640 860
rect 18660 840 18670 860
rect 18630 810 18670 840
rect 18630 790 18640 810
rect 18660 790 18670 810
rect 18630 760 18670 790
rect 18630 740 18640 760
rect 18660 740 18670 760
rect 18630 710 18670 740
rect 18865 910 18905 925
rect 18865 890 18875 910
rect 18895 890 18905 910
rect 18865 860 18905 890
rect 18865 840 18875 860
rect 18895 840 18905 860
rect 18865 810 18905 840
rect 18865 790 18875 810
rect 18895 790 18905 810
rect 18865 760 18905 790
rect 18865 740 18875 760
rect 18895 740 18905 760
rect 18865 725 18905 740
rect 19110 910 19150 925
rect 19110 890 19120 910
rect 19140 890 19150 910
rect 19110 860 19150 890
rect 19110 840 19120 860
rect 19140 840 19150 860
rect 19110 810 19150 840
rect 19110 790 19120 810
rect 19140 790 19150 810
rect 19110 760 19150 790
rect 19110 740 19120 760
rect 19140 740 19150 760
rect 19110 725 19150 740
rect 18630 690 18640 710
rect 18660 690 18670 710
rect 18630 660 18670 690
rect 18630 640 18640 660
rect 18660 640 18670 660
rect 18630 625 18670 640
rect 16380 70 16420 85
rect 16380 50 16390 70
rect 16410 50 16420 70
rect 16380 20 16420 50
rect 16380 0 16390 20
rect 16410 0 16420 20
rect 16380 -15 16420 0
rect 17660 70 17700 85
rect 17660 50 17670 70
rect 17690 50 17700 70
rect 17660 20 17700 50
rect 17660 0 17670 20
rect 17690 0 17700 20
rect 17660 -15 17700 0
rect 17900 70 17940 85
rect 17900 50 17910 70
rect 17930 50 17940 70
rect 17900 20 17940 50
rect 17900 0 17910 20
rect 17930 0 17940 20
rect 17900 -15 17940 0
rect 19180 70 19220 85
rect 19180 50 19190 70
rect 19210 50 19220 70
rect 19180 20 19220 50
rect 19180 0 19190 20
rect 19210 0 19220 20
rect 19180 -15 19220 0
<< psubdiffcont >>
rect 17570 -235 17590 -215
rect 17570 -275 17590 -255
rect 17570 -315 17590 -295
rect 18010 -235 18030 -215
rect 18010 -275 18030 -255
rect 18010 -315 18030 -295
rect 17120 -770 17140 -750
rect 17120 -820 17140 -800
rect 17120 -870 17140 -850
rect 17120 -920 17140 -900
rect 17120 -970 17140 -950
rect 18460 -770 18480 -750
rect 18460 -820 18480 -800
rect 18460 -870 18480 -850
rect 18460 -920 18480 -900
rect 18460 -970 18480 -950
rect 18870 -1225 18890 -1205
rect 18870 -1275 18890 -1255
rect 16510 -1575 16530 -1555
rect 16510 -1625 16530 -1605
rect 16865 -1575 16885 -1555
rect 16865 -1625 16885 -1605
rect 16995 -1575 17015 -1555
rect 16995 -1625 17015 -1605
rect 17515 -1575 17535 -1555
rect 17515 -1625 17535 -1605
rect 17585 -1575 17605 -1555
rect 17585 -1625 17605 -1605
rect 17995 -1575 18015 -1555
rect 17995 -1625 18015 -1605
rect 18065 -1575 18085 -1555
rect 18065 -1625 18085 -1605
rect 18585 -1575 18605 -1555
rect 18585 -1625 18605 -1605
rect 17790 -4190 17810 -4170
rect 17790 -4240 17810 -4220
rect 17790 -4290 17810 -4270
<< nsubdiffcont >>
rect 16345 1355 16365 1377
rect 16345 1305 16365 1325
rect 16645 1355 16665 1377
rect 16645 1305 16665 1325
rect 16855 1305 16875 1377
rect 17265 1305 17285 1377
rect 17475 1355 17495 1377
rect 17475 1305 17495 1325
rect 18105 1355 18125 1377
rect 18105 1305 18125 1325
rect 18315 1305 18335 1377
rect 18725 1305 18745 1377
rect 16940 890 16960 910
rect 16940 840 16960 860
rect 16405 790 16425 810
rect 16405 740 16425 760
rect 16710 790 16730 810
rect 16710 740 16730 760
rect 16940 790 16960 810
rect 16940 740 16960 760
rect 16940 690 16960 710
rect 16940 640 16960 660
rect 18640 890 18660 910
rect 18640 840 18660 860
rect 18640 790 18660 810
rect 18640 740 18660 760
rect 18875 890 18895 910
rect 18875 840 18895 860
rect 18875 790 18895 810
rect 18875 740 18895 760
rect 19120 890 19140 910
rect 19120 840 19140 860
rect 19120 790 19140 810
rect 19120 740 19140 760
rect 18640 690 18660 710
rect 18640 640 18660 660
rect 16390 50 16410 70
rect 16390 0 16410 20
rect 17670 50 17690 70
rect 17670 0 17690 20
rect 17910 50 17930 70
rect 17910 0 17930 20
rect 19190 50 19210 70
rect 19190 0 19210 20
<< poly >>
rect 16485 1615 16525 1625
rect 16485 1595 16495 1615
rect 16515 1595 16525 1615
rect 16485 1585 16525 1595
rect 17780 1615 17820 1625
rect 17780 1595 17790 1615
rect 17810 1595 17820 1615
rect 17780 1585 17820 1595
rect 16365 1435 16405 1445
rect 16365 1415 16375 1435
rect 16395 1420 16405 1435
rect 16395 1415 16430 1420
rect 16495 1415 16515 1585
rect 16605 1435 16645 1445
rect 16605 1420 16615 1435
rect 16580 1415 16615 1420
rect 16635 1415 16645 1435
rect 16365 1405 16430 1415
rect 16415 1390 16430 1405
rect 16470 1400 16540 1415
rect 16470 1390 16485 1400
rect 16525 1390 16540 1400
rect 16580 1405 16645 1415
rect 16885 1435 16925 1445
rect 16885 1415 16895 1435
rect 16915 1415 16925 1435
rect 17055 1435 17085 1445
rect 17055 1415 17060 1435
rect 17080 1415 17085 1435
rect 17215 1435 17255 1445
rect 17215 1415 17225 1435
rect 17245 1415 17255 1435
rect 16580 1390 16595 1405
rect 16885 1400 16940 1415
rect 16925 1390 16940 1400
rect 16980 1400 17160 1415
rect 16980 1390 16995 1400
rect 17035 1390 17050 1400
rect 17090 1390 17105 1400
rect 17145 1390 17160 1400
rect 17200 1400 17255 1415
rect 17495 1435 17535 1445
rect 17495 1415 17505 1435
rect 17525 1420 17535 1435
rect 17525 1415 17560 1420
rect 17790 1415 17810 1585
rect 18065 1435 18105 1445
rect 18065 1420 18075 1435
rect 18040 1415 18075 1420
rect 18095 1415 18105 1435
rect 17495 1405 17560 1415
rect 17200 1390 17215 1400
rect 17545 1390 17560 1405
rect 17600 1400 18000 1415
rect 17600 1390 17615 1400
rect 17655 1390 17670 1400
rect 17710 1390 17725 1400
rect 17765 1390 17780 1400
rect 17820 1390 17835 1400
rect 17875 1390 17890 1400
rect 17930 1390 17945 1400
rect 17985 1390 18000 1400
rect 18040 1405 18105 1415
rect 18345 1435 18385 1445
rect 18345 1415 18355 1435
rect 18375 1420 18385 1435
rect 18515 1435 18545 1445
rect 18375 1415 18400 1420
rect 18515 1415 18520 1435
rect 18540 1415 18545 1435
rect 18675 1435 18715 1445
rect 18675 1420 18685 1435
rect 18660 1415 18685 1420
rect 18705 1415 18715 1435
rect 18345 1405 18400 1415
rect 18040 1390 18055 1405
rect 18385 1390 18400 1405
rect 18440 1400 18620 1415
rect 18440 1390 18455 1400
rect 18495 1390 18510 1400
rect 18550 1390 18565 1400
rect 18605 1390 18620 1400
rect 18660 1405 18715 1415
rect 18660 1390 18675 1405
rect 16415 1275 16430 1290
rect 16470 1275 16485 1290
rect 16525 1275 16540 1290
rect 16580 1275 16595 1290
rect 16925 1275 16940 1290
rect 16980 1275 16995 1290
rect 17035 1275 17050 1290
rect 17090 1275 17105 1290
rect 17145 1275 17160 1290
rect 17200 1275 17215 1290
rect 17545 1275 17560 1290
rect 17600 1275 17615 1290
rect 17655 1275 17670 1290
rect 17710 1275 17725 1290
rect 17765 1275 17780 1290
rect 17820 1275 17835 1290
rect 17875 1275 17890 1290
rect 17930 1275 17945 1290
rect 17985 1275 18000 1290
rect 18040 1275 18055 1290
rect 18385 1275 18400 1290
rect 18440 1275 18455 1290
rect 18495 1275 18510 1290
rect 18550 1275 18565 1290
rect 18605 1275 18620 1290
rect 18660 1275 18675 1290
rect 16970 970 17010 980
rect 16970 950 16980 970
rect 17000 955 17010 970
rect 18590 970 18630 980
rect 18590 955 18600 970
rect 17000 950 17060 955
rect 16970 940 17060 950
rect 18540 950 18600 955
rect 18620 950 18630 970
rect 18540 940 18630 950
rect 18910 970 18940 980
rect 18910 950 18915 970
rect 18935 955 18940 970
rect 19080 970 19110 980
rect 19080 955 19085 970
rect 18935 950 18960 955
rect 18910 940 18960 950
rect 19055 950 19085 955
rect 19105 950 19110 970
rect 19055 940 19110 950
rect 17010 925 17060 940
rect 17100 925 17150 940
rect 17190 925 17240 940
rect 17280 925 17330 940
rect 17370 925 17420 940
rect 17460 925 17510 940
rect 17550 925 17600 940
rect 17640 925 17690 940
rect 17730 925 17780 940
rect 17820 925 17870 940
rect 17910 925 17960 940
rect 18000 925 18050 940
rect 18090 925 18140 940
rect 18180 925 18230 940
rect 18270 925 18320 940
rect 18360 925 18410 940
rect 18450 925 18500 940
rect 18540 925 18590 940
rect 18945 925 18960 940
rect 19000 925 19015 940
rect 19055 925 19070 940
rect 16440 870 16470 880
rect 16440 850 16445 870
rect 16465 850 16470 870
rect 16660 870 16690 880
rect 16660 850 16665 870
rect 16685 850 16690 870
rect 16440 835 16490 850
rect 16475 825 16490 835
rect 16530 825 16545 840
rect 16585 825 16600 840
rect 16640 835 16690 850
rect 16640 825 16655 835
rect 16475 710 16490 725
rect 16530 715 16545 725
rect 16585 715 16600 725
rect 16530 700 16600 715
rect 16640 710 16655 725
rect 16545 680 16555 700
rect 16575 680 16585 700
rect 16545 670 16585 680
rect 18945 710 18960 725
rect 19000 655 19015 725
rect 19055 710 19070 725
rect 19000 650 19040 655
rect 19000 630 19010 650
rect 19030 630 19040 650
rect 19000 625 19040 630
rect 17010 610 17060 625
rect 17100 615 17150 625
rect 17190 615 17240 625
rect 17280 615 17330 625
rect 17370 615 17420 625
rect 17460 615 17510 625
rect 17550 615 17600 625
rect 17640 615 17690 625
rect 17730 615 17780 625
rect 17820 615 17870 625
rect 17910 615 17960 625
rect 18000 615 18050 625
rect 18090 615 18140 625
rect 18180 615 18230 625
rect 18270 615 18320 625
rect 18360 615 18410 625
rect 18450 615 18500 625
rect 17100 600 18500 615
rect 18540 610 18590 625
rect 17690 580 17700 600
rect 17720 580 17730 600
rect 17690 570 17730 580
rect 18410 580 18420 600
rect 18440 580 18450 600
rect 18410 570 18450 580
rect 16425 130 16455 140
rect 16425 110 16430 130
rect 16450 110 16455 130
rect 17625 130 17655 140
rect 17625 110 17630 130
rect 17650 110 17655 130
rect 16425 95 16480 110
rect 16460 85 16480 95
rect 16520 85 16540 100
rect 16580 85 16600 100
rect 16640 85 16660 100
rect 16700 85 16720 100
rect 16760 85 16780 100
rect 16820 85 16840 100
rect 16880 85 16900 100
rect 16940 85 16960 100
rect 17000 85 17020 100
rect 17060 85 17080 100
rect 17120 85 17140 100
rect 17180 85 17200 100
rect 17240 85 17260 100
rect 17300 85 17320 100
rect 17360 85 17380 100
rect 17420 85 17440 100
rect 17480 85 17500 100
rect 17540 85 17560 100
rect 17600 95 17655 110
rect 17945 130 17975 140
rect 17945 110 17950 130
rect 17970 110 17975 130
rect 19145 130 19175 140
rect 19145 110 19150 130
rect 19170 110 19175 130
rect 17945 95 18000 110
rect 17600 85 17620 95
rect 17980 85 18000 95
rect 18040 85 18060 100
rect 18100 85 18120 100
rect 18160 85 18180 100
rect 18220 85 18240 100
rect 18280 85 18300 100
rect 18340 85 18360 100
rect 18400 85 18420 100
rect 18460 85 18480 100
rect 18520 85 18540 100
rect 18580 85 18600 100
rect 18640 85 18660 100
rect 18700 85 18720 100
rect 18760 85 18780 100
rect 18820 85 18840 100
rect 18880 85 18900 100
rect 18940 85 18960 100
rect 19000 85 19020 100
rect 19060 85 19080 100
rect 19120 95 19175 110
rect 19120 85 19140 95
rect 16460 -25 16480 -15
rect 16425 -40 16480 -25
rect 16520 -30 16540 -15
rect 16580 -25 16600 -15
rect 16640 -25 16660 -15
rect 16700 -25 16720 -15
rect 16760 -25 16780 -15
rect 16510 -40 16550 -30
rect 16580 -40 16780 -25
rect 16820 -25 16840 -15
rect 16880 -25 16900 -15
rect 16820 -40 16900 -25
rect 16940 -25 16960 -15
rect 17000 -25 17020 -15
rect 17060 -25 17080 -15
rect 17120 -25 17140 -15
rect 16940 -40 17140 -25
rect 17180 -25 17200 -15
rect 17240 -25 17260 -15
rect 17180 -40 17260 -25
rect 17300 -25 17320 -15
rect 17360 -25 17380 -15
rect 17420 -25 17440 -15
rect 17480 -25 17500 -15
rect 17300 -40 17500 -25
rect 17540 -30 17560 -15
rect 17600 -30 17620 -15
rect 17980 -25 18000 -15
rect 17535 -40 17565 -30
rect 16425 -60 16430 -40
rect 16450 -60 16455 -40
rect 16425 -70 16455 -60
rect 16510 -60 16520 -40
rect 16540 -60 16550 -40
rect 16510 -70 16550 -60
rect 16600 -60 16610 -40
rect 16630 -60 16640 -40
rect 16600 -70 16640 -60
rect 16840 -60 16850 -40
rect 16870 -60 16880 -40
rect 16840 -70 16880 -60
rect 16960 -60 16970 -40
rect 16990 -60 17000 -40
rect 16960 -70 17000 -60
rect 17200 -60 17210 -40
rect 17230 -60 17240 -40
rect 17200 -70 17240 -60
rect 17320 -60 17330 -40
rect 17350 -60 17360 -40
rect 17320 -70 17360 -60
rect 17535 -60 17540 -40
rect 17560 -60 17565 -40
rect 17535 -70 17565 -60
rect 17945 -40 18000 -25
rect 18040 -30 18060 -15
rect 18100 -25 18120 -15
rect 18160 -25 18180 -15
rect 18220 -25 18240 -15
rect 18280 -25 18300 -15
rect 18035 -40 18065 -30
rect 18100 -40 18300 -25
rect 18340 -25 18360 -15
rect 18400 -25 18420 -15
rect 18340 -40 18420 -25
rect 18460 -25 18480 -15
rect 18520 -25 18540 -15
rect 18580 -25 18600 -15
rect 18640 -25 18660 -15
rect 18460 -40 18660 -25
rect 18700 -25 18720 -15
rect 18760 -25 18780 -15
rect 18700 -40 18780 -25
rect 18820 -25 18840 -15
rect 18880 -25 18900 -15
rect 18940 -25 18960 -15
rect 19000 -25 19020 -15
rect 18820 -40 19020 -25
rect 19060 -30 19080 -15
rect 19120 -25 19140 -15
rect 19050 -40 19090 -30
rect 19120 -40 19175 -25
rect 17945 -60 17950 -40
rect 17970 -60 17975 -40
rect 17945 -70 17975 -60
rect 18035 -60 18040 -40
rect 18060 -60 18065 -40
rect 18035 -70 18065 -60
rect 18240 -60 18250 -40
rect 18270 -60 18280 -40
rect 18240 -70 18280 -60
rect 18360 -60 18370 -40
rect 18390 -60 18400 -40
rect 18360 -70 18400 -60
rect 18600 -60 18610 -40
rect 18630 -60 18640 -40
rect 18600 -70 18640 -60
rect 18720 -60 18730 -40
rect 18750 -60 18760 -40
rect 18720 -70 18760 -60
rect 18960 -60 18970 -40
rect 18990 -60 19000 -40
rect 18960 -70 19000 -60
rect 19050 -60 19060 -40
rect 19080 -60 19090 -40
rect 19050 -70 19090 -60
rect 19145 -60 19150 -40
rect 19170 -60 19175 -40
rect 19145 -70 19175 -60
rect 17007 -155 17037 -145
rect 17007 -170 17012 -155
rect 17000 -175 17012 -170
rect 17032 -175 17037 -155
rect 17000 -185 17037 -175
rect 18563 -155 18593 -145
rect 18563 -175 18568 -155
rect 18588 -170 18593 -155
rect 18588 -175 18600 -170
rect 18563 -185 18600 -175
rect 17000 -200 17020 -185
rect 17060 -200 17080 -185
rect 18520 -200 18540 -185
rect 18580 -200 18600 -185
rect 17000 -465 17020 -450
rect 17060 -465 17080 -450
rect 18520 -465 18540 -450
rect 18580 -465 18600 -450
rect 17060 -475 17105 -465
rect 17060 -495 17080 -475
rect 17100 -495 17105 -475
rect 17060 -505 17105 -495
rect 18495 -475 18540 -465
rect 18495 -495 18500 -475
rect 18520 -495 18540 -475
rect 18495 -505 18540 -495
rect 16620 -690 16660 -680
rect 16620 -710 16630 -690
rect 16650 -710 16660 -690
rect 16620 -720 16660 -710
rect 16740 -690 16780 -680
rect 16740 -710 16750 -690
rect 16770 -710 16780 -690
rect 16740 -720 16780 -710
rect 16860 -690 16900 -680
rect 16860 -710 16870 -690
rect 16890 -710 16900 -690
rect 16860 -720 16900 -710
rect 16980 -690 17020 -680
rect 16980 -710 16990 -690
rect 17010 -710 17020 -690
rect 16980 -720 17020 -710
rect 17300 -690 17340 -680
rect 17300 -710 17310 -690
rect 17330 -710 17340 -690
rect 17300 -720 17340 -710
rect 17420 -690 17460 -680
rect 17420 -710 17430 -690
rect 17450 -710 17460 -690
rect 17420 -720 17460 -710
rect 17540 -690 17580 -680
rect 17540 -710 17550 -690
rect 17570 -710 17580 -690
rect 17540 -720 17580 -710
rect 18020 -690 18060 -680
rect 18020 -710 18030 -690
rect 18050 -710 18060 -690
rect 18020 -720 18060 -710
rect 18140 -690 18180 -680
rect 18140 -710 18150 -690
rect 18170 -710 18180 -690
rect 18140 -720 18180 -710
rect 18260 -690 18300 -680
rect 18260 -710 18270 -690
rect 18290 -710 18300 -690
rect 18260 -720 18300 -710
rect 18580 -690 18620 -680
rect 18580 -710 18590 -690
rect 18610 -710 18620 -690
rect 18580 -720 18620 -710
rect 18700 -690 18740 -680
rect 18700 -710 18710 -690
rect 18730 -710 18740 -690
rect 18700 -720 18740 -710
rect 18820 -690 18860 -680
rect 18820 -710 18830 -690
rect 18850 -710 18860 -690
rect 18820 -720 18860 -710
rect 18940 -690 18980 -680
rect 18940 -710 18950 -690
rect 18970 -710 18980 -690
rect 18940 -720 18980 -710
rect 16570 -735 17070 -720
rect 17190 -735 17690 -720
rect 17910 -735 18410 -720
rect 18530 -735 19030 -720
rect 16570 -1000 17070 -985
rect 17190 -1000 17690 -985
rect 17910 -1000 18410 -985
rect 18530 -1000 19030 -985
rect 16820 -1145 16860 -1135
rect 16820 -1165 16830 -1145
rect 16850 -1165 16860 -1145
rect 16820 -1175 16860 -1165
rect 16900 -1145 16940 -1135
rect 16900 -1165 16910 -1145
rect 16930 -1165 16940 -1145
rect 16900 -1175 16940 -1165
rect 16980 -1145 17020 -1135
rect 16980 -1165 16990 -1145
rect 17010 -1165 17020 -1145
rect 16980 -1175 17020 -1165
rect 17060 -1145 17100 -1135
rect 17060 -1165 17070 -1145
rect 17090 -1165 17100 -1145
rect 17060 -1175 17100 -1165
rect 17140 -1145 17180 -1135
rect 17140 -1165 17150 -1145
rect 17170 -1165 17180 -1145
rect 17140 -1175 17180 -1165
rect 17220 -1145 17260 -1135
rect 17220 -1165 17230 -1145
rect 17250 -1165 17260 -1145
rect 17220 -1175 17260 -1165
rect 17300 -1145 17340 -1135
rect 17300 -1165 17310 -1145
rect 17330 -1165 17340 -1145
rect 17300 -1175 17340 -1165
rect 17380 -1145 17420 -1135
rect 17380 -1165 17390 -1145
rect 17410 -1165 17420 -1145
rect 17380 -1175 17420 -1165
rect 17460 -1145 17500 -1135
rect 17460 -1165 17470 -1145
rect 17490 -1165 17500 -1145
rect 17460 -1175 17500 -1165
rect 17540 -1145 17580 -1135
rect 17540 -1165 17550 -1145
rect 17570 -1165 17580 -1145
rect 17540 -1175 17580 -1165
rect 17620 -1145 17660 -1135
rect 17620 -1165 17630 -1145
rect 17650 -1165 17660 -1145
rect 17620 -1175 17660 -1165
rect 17700 -1145 17740 -1135
rect 17700 -1165 17710 -1145
rect 17730 -1165 17740 -1145
rect 17700 -1175 17740 -1165
rect 17860 -1145 17900 -1135
rect 17860 -1165 17870 -1145
rect 17890 -1165 17900 -1145
rect 17860 -1175 17900 -1165
rect 17940 -1145 17980 -1135
rect 17940 -1165 17950 -1145
rect 17970 -1165 17980 -1145
rect 17940 -1175 17980 -1165
rect 18020 -1145 18060 -1135
rect 18020 -1165 18030 -1145
rect 18050 -1165 18060 -1145
rect 18020 -1175 18060 -1165
rect 18100 -1145 18140 -1135
rect 18100 -1165 18110 -1145
rect 18130 -1165 18140 -1145
rect 18100 -1175 18140 -1165
rect 18180 -1145 18220 -1135
rect 18180 -1165 18190 -1145
rect 18210 -1165 18220 -1145
rect 18180 -1175 18220 -1165
rect 18260 -1145 18300 -1135
rect 18260 -1165 18270 -1145
rect 18290 -1165 18300 -1145
rect 18260 -1175 18300 -1165
rect 18340 -1145 18380 -1135
rect 18340 -1165 18350 -1145
rect 18370 -1165 18380 -1145
rect 18340 -1175 18380 -1165
rect 18420 -1145 18460 -1135
rect 18420 -1165 18430 -1145
rect 18450 -1165 18460 -1145
rect 18420 -1175 18460 -1165
rect 18500 -1145 18540 -1135
rect 18500 -1165 18510 -1145
rect 18530 -1165 18540 -1145
rect 18500 -1175 18540 -1165
rect 18580 -1145 18620 -1135
rect 18580 -1165 18590 -1145
rect 18610 -1165 18620 -1145
rect 18580 -1175 18620 -1165
rect 18660 -1145 18700 -1135
rect 18660 -1165 18670 -1145
rect 18690 -1165 18700 -1145
rect 18660 -1175 18700 -1165
rect 18740 -1145 18780 -1135
rect 18740 -1165 18750 -1145
rect 18770 -1165 18780 -1145
rect 18740 -1175 18780 -1165
rect 16780 -1190 17780 -1175
rect 17820 -1190 18820 -1175
rect 16780 -1305 17780 -1290
rect 17820 -1305 18820 -1290
rect 16540 -1495 16580 -1485
rect 16540 -1515 16550 -1495
rect 16570 -1510 16580 -1495
rect 16710 -1495 16740 -1485
rect 16570 -1515 16595 -1510
rect 16710 -1515 16715 -1495
rect 16735 -1515 16740 -1495
rect 16820 -1495 16860 -1485
rect 16820 -1510 16830 -1495
rect 16800 -1515 16830 -1510
rect 16850 -1515 16860 -1495
rect 16540 -1525 16595 -1515
rect 16580 -1540 16595 -1525
rect 16635 -1530 16760 -1515
rect 16635 -1540 16650 -1530
rect 16690 -1540 16705 -1530
rect 16745 -1540 16760 -1530
rect 16800 -1525 16860 -1515
rect 17025 -1495 17065 -1485
rect 17025 -1515 17035 -1495
rect 17055 -1510 17065 -1495
rect 17305 -1495 17335 -1485
rect 17055 -1515 17080 -1510
rect 17305 -1515 17310 -1495
rect 17330 -1515 17335 -1495
rect 17465 -1495 17505 -1485
rect 17465 -1510 17475 -1495
rect 17450 -1515 17475 -1510
rect 17495 -1515 17505 -1495
rect 17025 -1525 17080 -1515
rect 16800 -1540 16815 -1525
rect 17065 -1540 17080 -1525
rect 17120 -1530 17410 -1515
rect 17120 -1540 17135 -1530
rect 17175 -1540 17190 -1530
rect 17230 -1540 17245 -1530
rect 17285 -1540 17300 -1530
rect 17340 -1540 17355 -1530
rect 17395 -1540 17410 -1530
rect 17450 -1525 17505 -1515
rect 17615 -1495 17655 -1485
rect 17615 -1515 17625 -1495
rect 17645 -1510 17655 -1495
rect 17785 -1495 17815 -1485
rect 17645 -1515 17670 -1510
rect 17785 -1515 17790 -1495
rect 17810 -1515 17815 -1495
rect 17945 -1495 17985 -1485
rect 17945 -1510 17955 -1495
rect 17930 -1515 17955 -1510
rect 17975 -1515 17985 -1495
rect 17615 -1525 17670 -1515
rect 17450 -1540 17465 -1525
rect 17655 -1540 17670 -1525
rect 17710 -1530 17890 -1515
rect 17710 -1540 17725 -1530
rect 17765 -1540 17780 -1530
rect 17820 -1540 17835 -1530
rect 17875 -1540 17890 -1530
rect 17930 -1525 17985 -1515
rect 18095 -1495 18135 -1485
rect 18095 -1515 18105 -1495
rect 18125 -1510 18135 -1495
rect 18265 -1495 18295 -1485
rect 18125 -1515 18150 -1510
rect 18265 -1515 18270 -1495
rect 18290 -1515 18295 -1495
rect 18535 -1495 18575 -1485
rect 18535 -1510 18545 -1495
rect 18520 -1515 18545 -1510
rect 18565 -1515 18575 -1495
rect 18095 -1525 18150 -1515
rect 17930 -1540 17945 -1525
rect 18135 -1540 18150 -1525
rect 18190 -1530 18480 -1515
rect 18190 -1540 18205 -1530
rect 18245 -1540 18260 -1530
rect 18300 -1540 18315 -1530
rect 18355 -1540 18370 -1530
rect 18410 -1540 18425 -1530
rect 18465 -1540 18480 -1530
rect 18520 -1525 18575 -1515
rect 18520 -1540 18535 -1525
rect 16580 -1655 16595 -1640
rect 16635 -1655 16650 -1640
rect 16690 -1655 16705 -1640
rect 16745 -1655 16760 -1640
rect 16800 -1655 16815 -1640
rect 17065 -1655 17080 -1640
rect 17120 -1655 17135 -1640
rect 17175 -1655 17190 -1640
rect 17230 -1655 17245 -1640
rect 17285 -1655 17300 -1640
rect 17340 -1655 17355 -1640
rect 17395 -1655 17410 -1640
rect 17450 -1655 17465 -1640
rect 17655 -1655 17670 -1640
rect 17710 -1655 17725 -1640
rect 17765 -1655 17780 -1640
rect 17820 -1655 17835 -1640
rect 17875 -1655 17890 -1640
rect 17930 -1655 17945 -1640
rect 18135 -1655 18150 -1640
rect 18190 -1655 18205 -1640
rect 18245 -1655 18260 -1640
rect 18300 -1655 18315 -1640
rect 18355 -1655 18370 -1640
rect 18410 -1655 18425 -1640
rect 18465 -1655 18480 -1640
rect 18520 -1655 18535 -1640
<< polycont >>
rect 16495 1595 16515 1615
rect 17790 1595 17810 1615
rect 16375 1415 16395 1435
rect 16615 1415 16635 1435
rect 16895 1415 16915 1435
rect 17060 1415 17080 1435
rect 17225 1415 17245 1435
rect 17505 1415 17525 1435
rect 18075 1415 18095 1435
rect 18355 1415 18375 1435
rect 18520 1415 18540 1435
rect 18685 1415 18705 1435
rect 16980 950 17000 970
rect 18600 950 18620 970
rect 18915 950 18935 970
rect 19085 950 19105 970
rect 16445 850 16465 870
rect 16665 850 16685 870
rect 16555 680 16575 700
rect 19010 630 19030 650
rect 17700 580 17720 600
rect 18420 580 18440 600
rect 16430 110 16450 130
rect 17630 110 17650 130
rect 17950 110 17970 130
rect 19150 110 19170 130
rect 16430 -60 16450 -40
rect 16520 -60 16540 -40
rect 16610 -60 16630 -40
rect 16850 -60 16870 -40
rect 16970 -60 16990 -40
rect 17210 -60 17230 -40
rect 17330 -60 17350 -40
rect 17540 -60 17560 -40
rect 17950 -60 17970 -40
rect 18040 -60 18060 -40
rect 18250 -60 18270 -40
rect 18370 -60 18390 -40
rect 18610 -60 18630 -40
rect 18730 -60 18750 -40
rect 18970 -60 18990 -40
rect 19060 -60 19080 -40
rect 19150 -60 19170 -40
rect 17012 -175 17032 -155
rect 18568 -175 18588 -155
rect 17080 -495 17100 -475
rect 18500 -495 18520 -475
rect 16630 -710 16650 -690
rect 16750 -710 16770 -690
rect 16870 -710 16890 -690
rect 16990 -710 17010 -690
rect 17310 -710 17330 -690
rect 17430 -710 17450 -690
rect 17550 -710 17570 -690
rect 18030 -710 18050 -690
rect 18150 -710 18170 -690
rect 18270 -710 18290 -690
rect 18590 -710 18610 -690
rect 18710 -710 18730 -690
rect 18830 -710 18850 -690
rect 18950 -710 18970 -690
rect 16830 -1165 16850 -1145
rect 16910 -1165 16930 -1145
rect 16990 -1165 17010 -1145
rect 17070 -1165 17090 -1145
rect 17150 -1165 17170 -1145
rect 17230 -1165 17250 -1145
rect 17310 -1165 17330 -1145
rect 17390 -1165 17410 -1145
rect 17470 -1165 17490 -1145
rect 17550 -1165 17570 -1145
rect 17630 -1165 17650 -1145
rect 17710 -1165 17730 -1145
rect 17870 -1165 17890 -1145
rect 17950 -1165 17970 -1145
rect 18030 -1165 18050 -1145
rect 18110 -1165 18130 -1145
rect 18190 -1165 18210 -1145
rect 18270 -1165 18290 -1145
rect 18350 -1165 18370 -1145
rect 18430 -1165 18450 -1145
rect 18510 -1165 18530 -1145
rect 18590 -1165 18610 -1145
rect 18670 -1165 18690 -1145
rect 18750 -1165 18770 -1145
rect 16550 -1515 16570 -1495
rect 16715 -1515 16735 -1495
rect 16830 -1515 16850 -1495
rect 17035 -1515 17055 -1495
rect 17310 -1515 17330 -1495
rect 17475 -1515 17495 -1495
rect 17625 -1515 17645 -1495
rect 17790 -1515 17810 -1495
rect 17955 -1515 17975 -1495
rect 18105 -1515 18125 -1495
rect 18270 -1515 18290 -1495
rect 18545 -1515 18565 -1495
<< xpolycontact >>
rect 17470 -2035 17690 -2000
rect 17904 -2035 18124 -2000
rect 15950 -3376 15985 -3156
rect 15950 -3784 15985 -3565
rect 16160 -3285 16195 -3065
rect 16160 -3889 16195 -3669
rect 16220 -3285 16255 -3065
rect 16220 -3889 16255 -3669
rect 16280 -3285 16315 -3065
rect 16280 -3889 16315 -3669
rect 16485 -3160 16520 -2940
rect 16485 -3964 16520 -3744
rect 16545 -3160 16580 -2940
rect 16545 -3964 16580 -3744
rect 16605 -3160 16640 -2940
rect 16605 -3964 16640 -3744
rect 18960 -3160 18995 -2940
rect 18960 -3964 18995 -3744
rect 19020 -3160 19055 -2940
rect 19020 -3964 19055 -3744
rect 19080 -3160 19115 -2940
rect 19080 -3964 19115 -3744
rect 19285 -3257 19320 -3037
rect 19285 -3889 19320 -3669
rect 19345 -3257 19380 -3037
rect 19345 -3889 19380 -3669
rect 19405 -3257 19440 -3037
rect 19405 -3889 19440 -3669
rect 19610 -3376 19645 -3156
rect 19610 -3784 19645 -3565
<< ppolyres >>
rect 15950 -3565 15985 -3376
rect 19610 -3565 19645 -3376
<< xpolyres >>
rect 17690 -2035 17904 -2000
rect 16160 -3669 16195 -3285
rect 16220 -3669 16255 -3285
rect 16280 -3669 16315 -3285
rect 16485 -3744 16520 -3160
rect 16545 -3744 16580 -3160
rect 16605 -3744 16640 -3160
rect 18960 -3744 18995 -3160
rect 19020 -3744 19055 -3160
rect 19080 -3744 19115 -3160
rect 19285 -3669 19320 -3257
rect 19345 -3669 19380 -3257
rect 19405 -3669 19440 -3257
<< locali >>
rect 16485 1615 16525 1625
rect 16485 1595 16495 1615
rect 16515 1595 16525 1615
rect 16485 1585 16525 1595
rect 17780 1615 17820 1625
rect 17780 1595 17790 1615
rect 17810 1595 17820 1615
rect 17780 1585 17820 1595
rect 16365 1435 16405 1445
rect 16365 1415 16375 1435
rect 16395 1415 16405 1435
rect 16365 1405 16405 1415
rect 16485 1435 16525 1445
rect 16485 1415 16495 1435
rect 16515 1415 16525 1435
rect 16485 1405 16525 1415
rect 16605 1435 16645 1445
rect 16605 1415 16615 1435
rect 16635 1415 16645 1435
rect 16605 1405 16645 1415
rect 16885 1435 16925 1445
rect 16885 1415 16895 1435
rect 16915 1415 16925 1435
rect 16885 1405 16925 1415
rect 16945 1435 16975 1445
rect 16945 1415 16950 1435
rect 16970 1415 16975 1435
rect 16945 1405 16975 1415
rect 16995 1435 17035 1445
rect 16995 1415 17005 1435
rect 17025 1415 17035 1435
rect 16995 1405 17035 1415
rect 17055 1435 17085 1445
rect 17055 1415 17060 1435
rect 17080 1415 17085 1435
rect 17055 1405 17085 1415
rect 17105 1435 17145 1445
rect 17105 1415 17115 1435
rect 17135 1415 17145 1435
rect 17105 1405 17145 1415
rect 17215 1435 17255 1445
rect 17215 1415 17225 1435
rect 17245 1415 17255 1435
rect 17215 1405 17255 1415
rect 17495 1435 17535 1445
rect 17495 1415 17505 1435
rect 17525 1415 17535 1435
rect 17495 1405 17535 1415
rect 17560 1435 17600 1445
rect 17560 1415 17570 1435
rect 17590 1415 17600 1435
rect 17560 1405 17600 1415
rect 17620 1435 17650 1445
rect 17620 1415 17625 1435
rect 17645 1415 17650 1435
rect 16385 1385 16405 1405
rect 16495 1385 16515 1405
rect 16605 1385 16625 1405
rect 16895 1385 16915 1405
rect 16950 1385 16970 1405
rect 17005 1385 17025 1405
rect 17115 1385 17135 1405
rect 17225 1385 17245 1405
rect 17515 1385 17535 1405
rect 17570 1385 17590 1405
rect 16340 1377 16410 1385
rect 16340 1355 16345 1377
rect 16365 1375 16410 1377
rect 16365 1355 16385 1375
rect 16405 1355 16410 1375
rect 16340 1325 16410 1355
rect 16340 1305 16345 1325
rect 16365 1305 16385 1325
rect 16405 1305 16410 1325
rect 16340 1295 16410 1305
rect 16435 1375 16465 1385
rect 16435 1355 16440 1375
rect 16460 1355 16465 1375
rect 16435 1325 16465 1355
rect 16435 1305 16440 1325
rect 16460 1305 16465 1325
rect 16435 1295 16465 1305
rect 16490 1375 16520 1385
rect 16490 1355 16495 1375
rect 16515 1355 16520 1375
rect 16490 1325 16520 1355
rect 16490 1305 16495 1325
rect 16515 1305 16520 1325
rect 16490 1295 16520 1305
rect 16545 1375 16575 1385
rect 16545 1355 16550 1375
rect 16570 1355 16575 1375
rect 16545 1325 16575 1355
rect 16545 1305 16550 1325
rect 16570 1305 16575 1325
rect 16545 1295 16575 1305
rect 16600 1377 16670 1385
rect 16600 1375 16645 1377
rect 16600 1355 16605 1375
rect 16625 1355 16645 1375
rect 16665 1355 16670 1377
rect 16600 1325 16670 1355
rect 16600 1305 16605 1325
rect 16625 1305 16645 1325
rect 16665 1305 16670 1325
rect 16600 1295 16670 1305
rect 16850 1377 16920 1385
rect 16850 1305 16855 1377
rect 16875 1375 16920 1377
rect 16875 1305 16895 1375
rect 16850 1303 16895 1305
rect 16915 1303 16920 1375
rect 16850 1295 16920 1303
rect 16945 1375 16975 1385
rect 16945 1303 16950 1375
rect 16970 1303 16975 1375
rect 16945 1295 16975 1303
rect 17000 1375 17030 1385
rect 17000 1303 17005 1375
rect 17025 1303 17030 1375
rect 17000 1295 17030 1303
rect 17055 1375 17085 1385
rect 17055 1303 17060 1375
rect 17080 1303 17085 1375
rect 17055 1295 17085 1303
rect 17110 1375 17140 1385
rect 17110 1303 17115 1375
rect 17135 1303 17140 1375
rect 17110 1295 17140 1303
rect 17165 1375 17195 1385
rect 17165 1303 17170 1375
rect 17190 1303 17195 1375
rect 17165 1295 17195 1303
rect 17220 1377 17290 1385
rect 17220 1375 17265 1377
rect 17220 1303 17225 1375
rect 17245 1305 17265 1375
rect 17285 1305 17290 1377
rect 17245 1303 17290 1305
rect 17220 1295 17290 1303
rect 17470 1377 17540 1385
rect 17470 1355 17475 1377
rect 17495 1375 17540 1377
rect 17495 1355 17515 1375
rect 17535 1355 17540 1375
rect 17470 1325 17540 1355
rect 17470 1305 17475 1325
rect 17495 1305 17515 1325
rect 17535 1305 17540 1325
rect 17470 1295 17540 1305
rect 17565 1375 17595 1385
rect 17565 1355 17570 1375
rect 17590 1355 17595 1375
rect 17565 1325 17595 1355
rect 17565 1305 17570 1325
rect 17590 1305 17595 1325
rect 17565 1295 17595 1305
rect 17620 1375 17650 1415
rect 17670 1435 17710 1445
rect 17670 1415 17680 1435
rect 17700 1415 17710 1435
rect 17670 1405 17710 1415
rect 17730 1435 17760 1445
rect 17730 1415 17735 1435
rect 17755 1415 17760 1435
rect 17680 1385 17700 1405
rect 17620 1355 17625 1375
rect 17645 1355 17650 1375
rect 17620 1325 17650 1355
rect 17620 1305 17625 1325
rect 17645 1305 17650 1325
rect 17620 1295 17650 1305
rect 17675 1375 17705 1385
rect 17675 1355 17680 1375
rect 17700 1355 17705 1375
rect 17675 1325 17705 1355
rect 17675 1305 17680 1325
rect 17700 1305 17705 1325
rect 17675 1295 17705 1305
rect 17730 1375 17760 1415
rect 17780 1435 17820 1445
rect 17780 1415 17790 1435
rect 17810 1415 17820 1435
rect 17780 1405 17820 1415
rect 17840 1435 17870 1445
rect 17840 1415 17845 1435
rect 17865 1415 17870 1435
rect 17790 1385 17810 1405
rect 17730 1355 17735 1375
rect 17755 1355 17760 1375
rect 17730 1325 17760 1355
rect 17730 1305 17735 1325
rect 17755 1305 17760 1325
rect 17730 1295 17760 1305
rect 17785 1375 17815 1385
rect 17785 1355 17790 1375
rect 17810 1355 17815 1375
rect 17785 1325 17815 1355
rect 17785 1305 17790 1325
rect 17810 1305 17815 1325
rect 17785 1295 17815 1305
rect 17840 1375 17870 1415
rect 17890 1435 17930 1445
rect 17890 1415 17900 1435
rect 17920 1415 17930 1435
rect 17890 1405 17930 1415
rect 17950 1435 17980 1445
rect 17950 1415 17955 1435
rect 17975 1415 17980 1435
rect 17900 1385 17920 1405
rect 17840 1355 17845 1375
rect 17865 1355 17870 1375
rect 17840 1325 17870 1355
rect 17840 1305 17845 1325
rect 17865 1305 17870 1325
rect 17840 1295 17870 1305
rect 17895 1375 17925 1385
rect 17895 1355 17900 1375
rect 17920 1355 17925 1375
rect 17895 1325 17925 1355
rect 17895 1305 17900 1325
rect 17920 1305 17925 1325
rect 17895 1295 17925 1305
rect 17950 1375 17980 1415
rect 18000 1435 18040 1445
rect 18000 1415 18010 1435
rect 18030 1415 18040 1435
rect 18000 1405 18040 1415
rect 18065 1435 18105 1445
rect 18065 1415 18075 1435
rect 18095 1415 18105 1435
rect 18065 1405 18105 1415
rect 18345 1435 18385 1445
rect 18345 1415 18355 1435
rect 18375 1415 18385 1435
rect 18345 1405 18385 1415
rect 18455 1435 18495 1445
rect 18455 1415 18465 1435
rect 18485 1415 18495 1435
rect 18455 1405 18495 1415
rect 18515 1435 18545 1445
rect 18515 1415 18520 1435
rect 18540 1415 18545 1435
rect 18515 1405 18545 1415
rect 18565 1435 18605 1445
rect 18565 1415 18575 1435
rect 18595 1415 18605 1435
rect 18565 1405 18605 1415
rect 18625 1435 18655 1445
rect 18625 1415 18630 1435
rect 18650 1415 18655 1435
rect 18625 1405 18655 1415
rect 18675 1435 18715 1445
rect 18675 1415 18685 1435
rect 18705 1415 18715 1435
rect 18675 1405 18715 1415
rect 18010 1385 18030 1405
rect 18065 1385 18085 1405
rect 18355 1385 18375 1405
rect 18465 1385 18485 1405
rect 18575 1385 18595 1405
rect 18630 1385 18650 1405
rect 18685 1385 18705 1405
rect 17950 1355 17955 1375
rect 17975 1355 17980 1375
rect 17950 1325 17980 1355
rect 17950 1305 17955 1325
rect 17975 1305 17980 1325
rect 17950 1295 17980 1305
rect 18005 1375 18035 1385
rect 18005 1355 18010 1375
rect 18030 1355 18035 1375
rect 18005 1325 18035 1355
rect 18005 1305 18010 1325
rect 18030 1305 18035 1325
rect 18005 1295 18035 1305
rect 18060 1377 18130 1385
rect 18060 1375 18105 1377
rect 18060 1355 18065 1375
rect 18085 1355 18105 1375
rect 18125 1355 18130 1377
rect 18060 1325 18130 1355
rect 18060 1305 18065 1325
rect 18085 1305 18105 1325
rect 18125 1305 18130 1325
rect 18060 1295 18130 1305
rect 18310 1377 18380 1385
rect 18310 1305 18315 1377
rect 18335 1375 18380 1377
rect 18335 1305 18355 1375
rect 18375 1305 18380 1375
rect 18310 1295 18380 1305
rect 18405 1375 18435 1385
rect 18405 1305 18410 1375
rect 18430 1305 18435 1375
rect 18405 1295 18435 1305
rect 18460 1375 18490 1385
rect 18460 1305 18465 1375
rect 18485 1305 18490 1375
rect 18460 1295 18490 1305
rect 18515 1375 18545 1385
rect 18515 1305 18520 1375
rect 18540 1305 18545 1375
rect 18515 1295 18545 1305
rect 18570 1375 18600 1385
rect 18570 1305 18575 1375
rect 18595 1305 18600 1375
rect 18570 1295 18600 1305
rect 18625 1375 18655 1385
rect 18625 1305 18630 1375
rect 18650 1305 18655 1375
rect 18625 1295 18655 1305
rect 18680 1377 18750 1385
rect 18680 1375 18725 1377
rect 18680 1305 18685 1375
rect 18705 1305 18725 1375
rect 18745 1305 18750 1377
rect 18680 1295 18750 1305
rect 16440 1275 16460 1295
rect 16550 1275 16570 1295
rect 16950 1275 16970 1295
rect 17060 1275 17080 1295
rect 17170 1275 17190 1295
rect 17625 1275 17645 1295
rect 17735 1275 17755 1295
rect 17845 1275 17865 1295
rect 17955 1275 17975 1295
rect 18410 1275 18430 1295
rect 18520 1275 18540 1295
rect 18630 1275 18650 1295
rect 16430 1265 16470 1275
rect 16430 1245 16440 1265
rect 16460 1245 16470 1265
rect 16430 1235 16470 1245
rect 16540 1265 16580 1275
rect 16540 1245 16550 1265
rect 16570 1245 16580 1265
rect 16540 1235 16580 1245
rect 16940 1265 16980 1275
rect 16940 1245 16950 1265
rect 16970 1245 16980 1265
rect 16940 1235 16980 1245
rect 17050 1265 17090 1275
rect 17050 1245 17060 1265
rect 17080 1245 17090 1265
rect 17050 1235 17090 1245
rect 17160 1265 17200 1275
rect 17160 1245 17170 1265
rect 17190 1245 17200 1265
rect 17160 1235 17200 1245
rect 17615 1265 17655 1275
rect 17615 1245 17625 1265
rect 17645 1245 17655 1265
rect 17615 1235 17655 1245
rect 17725 1265 17765 1275
rect 17725 1245 17735 1265
rect 17755 1245 17765 1265
rect 17725 1235 17765 1245
rect 17835 1265 17875 1275
rect 17835 1245 17845 1265
rect 17865 1245 17875 1265
rect 17835 1235 17875 1245
rect 17945 1265 17985 1275
rect 17945 1245 17955 1265
rect 17975 1245 17985 1265
rect 17945 1235 17985 1245
rect 18400 1265 18440 1275
rect 18400 1245 18410 1265
rect 18430 1245 18440 1265
rect 18400 1235 18440 1245
rect 18510 1265 18550 1275
rect 18510 1245 18520 1265
rect 18540 1245 18550 1265
rect 18510 1235 18550 1245
rect 18620 1265 18660 1275
rect 18620 1245 18630 1265
rect 18650 1245 18660 1265
rect 18620 1235 18660 1245
rect 16970 970 17010 980
rect 16970 950 16980 970
rect 17000 950 17010 970
rect 16970 940 17010 950
rect 17150 970 17190 980
rect 17150 950 17160 970
rect 17180 950 17190 970
rect 17150 940 17190 950
rect 17330 970 17370 980
rect 17330 950 17340 970
rect 17360 950 17370 970
rect 17330 940 17370 950
rect 17510 970 17550 980
rect 17510 950 17520 970
rect 17540 950 17550 970
rect 17510 940 17550 950
rect 17690 970 17730 980
rect 17690 950 17700 970
rect 17720 950 17730 970
rect 17690 940 17730 950
rect 17870 970 17910 980
rect 17870 950 17880 970
rect 17900 950 17910 970
rect 17870 940 17910 950
rect 18050 970 18090 980
rect 18050 950 18060 970
rect 18080 950 18090 970
rect 18050 940 18090 950
rect 18230 970 18270 980
rect 18230 950 18240 970
rect 18260 950 18270 970
rect 18230 940 18270 950
rect 18410 970 18450 980
rect 18410 950 18420 970
rect 18440 950 18450 970
rect 18410 940 18450 950
rect 18590 970 18630 980
rect 18590 950 18600 970
rect 18620 950 18630 970
rect 18590 940 18630 950
rect 18905 970 18945 980
rect 18905 950 18915 970
rect 18935 950 18945 970
rect 18905 940 18945 950
rect 19015 970 19055 980
rect 19015 950 19025 970
rect 19045 950 19055 970
rect 19015 940 19055 950
rect 19075 970 19115 980
rect 19075 950 19085 970
rect 19105 950 19115 970
rect 19075 940 19115 950
rect 16980 920 17000 940
rect 17160 920 17180 940
rect 17340 920 17360 940
rect 17520 920 17540 940
rect 17700 920 17720 940
rect 17880 920 17900 940
rect 18060 920 18080 940
rect 18240 920 18260 940
rect 18420 920 18440 940
rect 18600 920 18620 940
rect 18915 920 18935 940
rect 19025 920 19045 940
rect 19080 920 19100 940
rect 16935 910 17005 920
rect 16935 890 16940 910
rect 16960 890 16980 910
rect 17000 890 17005 910
rect 16440 870 16470 880
rect 16440 850 16445 870
rect 16465 850 16470 870
rect 16440 820 16470 850
rect 16545 870 16585 880
rect 16545 850 16555 870
rect 16575 850 16585 870
rect 16545 840 16585 850
rect 16655 870 16695 880
rect 16655 850 16665 870
rect 16685 850 16695 870
rect 16655 840 16695 850
rect 16935 860 17005 890
rect 16935 840 16940 860
rect 16960 840 16980 860
rect 17000 840 17005 860
rect 16555 820 16575 840
rect 16660 820 16690 840
rect 16400 810 16470 820
rect 16400 790 16405 810
rect 16425 790 16445 810
rect 16465 790 16470 810
rect 16400 760 16470 790
rect 16400 740 16405 760
rect 16425 740 16445 760
rect 16465 740 16470 760
rect 16400 730 16470 740
rect 16495 810 16525 820
rect 16495 790 16500 810
rect 16520 790 16525 810
rect 16495 760 16525 790
rect 16495 740 16500 760
rect 16520 740 16525 760
rect 16495 730 16525 740
rect 16550 810 16580 820
rect 16550 790 16555 810
rect 16575 790 16580 810
rect 16550 760 16580 790
rect 16550 740 16555 760
rect 16575 740 16580 760
rect 16550 730 16580 740
rect 16605 810 16635 820
rect 16605 790 16610 810
rect 16630 790 16635 810
rect 16605 760 16635 790
rect 16605 740 16610 760
rect 16630 740 16635 760
rect 16605 730 16635 740
rect 16660 810 16735 820
rect 16660 790 16665 810
rect 16685 790 16710 810
rect 16730 790 16735 810
rect 16660 760 16735 790
rect 16660 740 16665 760
rect 16685 740 16710 760
rect 16730 740 16735 760
rect 16660 730 16735 740
rect 16935 810 17005 840
rect 16935 790 16940 810
rect 16960 790 16980 810
rect 17000 790 17005 810
rect 16935 760 17005 790
rect 16935 740 16940 760
rect 16960 740 16980 760
rect 17000 740 17005 760
rect 16500 710 16520 730
rect 16610 710 16630 730
rect 16935 710 17005 740
rect 16480 700 16520 710
rect 16480 680 16490 700
rect 16510 680 16520 700
rect 16480 670 16520 680
rect 16545 700 16585 710
rect 16545 680 16555 700
rect 16575 680 16585 700
rect 16545 670 16585 680
rect 16610 700 16650 710
rect 16610 680 16620 700
rect 16640 680 16650 700
rect 16610 670 16650 680
rect 16935 690 16940 710
rect 16960 690 16980 710
rect 17000 690 17005 710
rect 16935 660 17005 690
rect 16935 640 16940 660
rect 16960 640 16980 660
rect 17000 640 17005 660
rect 16935 630 17005 640
rect 17065 910 17095 920
rect 17065 890 17070 910
rect 17090 890 17095 910
rect 17065 860 17095 890
rect 17065 840 17070 860
rect 17090 840 17095 860
rect 17065 810 17095 840
rect 17065 790 17070 810
rect 17090 790 17095 810
rect 17065 760 17095 790
rect 17065 740 17070 760
rect 17090 740 17095 760
rect 17065 710 17095 740
rect 17065 690 17070 710
rect 17090 690 17095 710
rect 17065 660 17095 690
rect 17065 640 17070 660
rect 17090 640 17095 660
rect 17065 630 17095 640
rect 17155 910 17185 920
rect 17155 890 17160 910
rect 17180 890 17185 910
rect 17155 860 17185 890
rect 17155 840 17160 860
rect 17180 840 17185 860
rect 17155 810 17185 840
rect 17155 790 17160 810
rect 17180 790 17185 810
rect 17155 760 17185 790
rect 17155 740 17160 760
rect 17180 740 17185 760
rect 17155 710 17185 740
rect 17155 690 17160 710
rect 17180 690 17185 710
rect 17155 660 17185 690
rect 17155 640 17160 660
rect 17180 640 17185 660
rect 17155 630 17185 640
rect 17245 910 17275 920
rect 17245 890 17250 910
rect 17270 890 17275 910
rect 17245 860 17275 890
rect 17245 840 17250 860
rect 17270 840 17275 860
rect 17245 810 17275 840
rect 17245 790 17250 810
rect 17270 790 17275 810
rect 17245 760 17275 790
rect 17245 740 17250 760
rect 17270 740 17275 760
rect 17245 710 17275 740
rect 17245 690 17250 710
rect 17270 690 17275 710
rect 17245 660 17275 690
rect 17245 640 17250 660
rect 17270 640 17275 660
rect 17245 630 17275 640
rect 17335 910 17365 920
rect 17335 890 17340 910
rect 17360 890 17365 910
rect 17335 860 17365 890
rect 17335 840 17340 860
rect 17360 840 17365 860
rect 17335 810 17365 840
rect 17335 790 17340 810
rect 17360 790 17365 810
rect 17335 760 17365 790
rect 17335 740 17340 760
rect 17360 740 17365 760
rect 17335 710 17365 740
rect 17335 690 17340 710
rect 17360 690 17365 710
rect 17335 660 17365 690
rect 17335 640 17340 660
rect 17360 640 17365 660
rect 17335 630 17365 640
rect 17425 910 17455 920
rect 17425 890 17430 910
rect 17450 890 17455 910
rect 17425 860 17455 890
rect 17425 840 17430 860
rect 17450 840 17455 860
rect 17425 810 17455 840
rect 17425 790 17430 810
rect 17450 790 17455 810
rect 17425 760 17455 790
rect 17425 740 17430 760
rect 17450 740 17455 760
rect 17425 710 17455 740
rect 17425 690 17430 710
rect 17450 690 17455 710
rect 17425 660 17455 690
rect 17425 640 17430 660
rect 17450 640 17455 660
rect 17425 630 17455 640
rect 17515 910 17545 920
rect 17515 890 17520 910
rect 17540 890 17545 910
rect 17515 860 17545 890
rect 17515 840 17520 860
rect 17540 840 17545 860
rect 17515 810 17545 840
rect 17515 790 17520 810
rect 17540 790 17545 810
rect 17515 760 17545 790
rect 17515 740 17520 760
rect 17540 740 17545 760
rect 17515 710 17545 740
rect 17515 690 17520 710
rect 17540 690 17545 710
rect 17515 660 17545 690
rect 17515 640 17520 660
rect 17540 640 17545 660
rect 17515 630 17545 640
rect 17605 910 17635 920
rect 17605 890 17610 910
rect 17630 890 17635 910
rect 17605 860 17635 890
rect 17605 840 17610 860
rect 17630 840 17635 860
rect 17605 810 17635 840
rect 17605 790 17610 810
rect 17630 790 17635 810
rect 17605 760 17635 790
rect 17605 740 17610 760
rect 17630 740 17635 760
rect 17605 710 17635 740
rect 17605 690 17610 710
rect 17630 690 17635 710
rect 17605 660 17635 690
rect 17605 640 17610 660
rect 17630 640 17635 660
rect 17605 630 17635 640
rect 17695 910 17725 920
rect 17695 890 17700 910
rect 17720 890 17725 910
rect 17695 860 17725 890
rect 17695 840 17700 860
rect 17720 840 17725 860
rect 17695 810 17725 840
rect 17695 790 17700 810
rect 17720 790 17725 810
rect 17695 760 17725 790
rect 17695 740 17700 760
rect 17720 740 17725 760
rect 17695 710 17725 740
rect 17695 690 17700 710
rect 17720 690 17725 710
rect 17695 660 17725 690
rect 17695 640 17700 660
rect 17720 640 17725 660
rect 17695 630 17725 640
rect 17785 910 17815 920
rect 17785 890 17790 910
rect 17810 890 17815 910
rect 17785 860 17815 890
rect 17785 840 17790 860
rect 17810 840 17815 860
rect 17785 810 17815 840
rect 17785 790 17790 810
rect 17810 790 17815 810
rect 17785 760 17815 790
rect 17785 740 17790 760
rect 17810 740 17815 760
rect 17785 710 17815 740
rect 17785 690 17790 710
rect 17810 690 17815 710
rect 17785 660 17815 690
rect 17785 640 17790 660
rect 17810 640 17815 660
rect 17785 630 17815 640
rect 17875 910 17905 920
rect 17875 890 17880 910
rect 17900 890 17905 910
rect 17875 860 17905 890
rect 17875 840 17880 860
rect 17900 840 17905 860
rect 17875 810 17905 840
rect 17875 790 17880 810
rect 17900 790 17905 810
rect 17875 760 17905 790
rect 17875 740 17880 760
rect 17900 740 17905 760
rect 17875 710 17905 740
rect 17875 690 17880 710
rect 17900 690 17905 710
rect 17875 660 17905 690
rect 17875 640 17880 660
rect 17900 640 17905 660
rect 17875 630 17905 640
rect 17965 910 17995 920
rect 17965 890 17970 910
rect 17990 890 17995 910
rect 17965 860 17995 890
rect 17965 840 17970 860
rect 17990 840 17995 860
rect 17965 810 17995 840
rect 17965 790 17970 810
rect 17990 790 17995 810
rect 17965 760 17995 790
rect 17965 740 17970 760
rect 17990 740 17995 760
rect 17965 710 17995 740
rect 17965 690 17970 710
rect 17990 690 17995 710
rect 17965 660 17995 690
rect 17965 640 17970 660
rect 17990 640 17995 660
rect 17965 630 17995 640
rect 18055 910 18085 920
rect 18055 890 18060 910
rect 18080 890 18085 910
rect 18055 860 18085 890
rect 18055 840 18060 860
rect 18080 840 18085 860
rect 18055 810 18085 840
rect 18055 790 18060 810
rect 18080 790 18085 810
rect 18055 760 18085 790
rect 18055 740 18060 760
rect 18080 740 18085 760
rect 18055 710 18085 740
rect 18055 690 18060 710
rect 18080 690 18085 710
rect 18055 660 18085 690
rect 18055 640 18060 660
rect 18080 640 18085 660
rect 18055 630 18085 640
rect 18145 910 18175 920
rect 18145 890 18150 910
rect 18170 890 18175 910
rect 18145 860 18175 890
rect 18145 840 18150 860
rect 18170 840 18175 860
rect 18145 810 18175 840
rect 18145 790 18150 810
rect 18170 790 18175 810
rect 18145 760 18175 790
rect 18145 740 18150 760
rect 18170 740 18175 760
rect 18145 710 18175 740
rect 18145 690 18150 710
rect 18170 690 18175 710
rect 18145 660 18175 690
rect 18145 640 18150 660
rect 18170 640 18175 660
rect 18145 630 18175 640
rect 18235 910 18265 920
rect 18235 890 18240 910
rect 18260 890 18265 910
rect 18235 860 18265 890
rect 18235 840 18240 860
rect 18260 840 18265 860
rect 18235 810 18265 840
rect 18235 790 18240 810
rect 18260 790 18265 810
rect 18235 760 18265 790
rect 18235 740 18240 760
rect 18260 740 18265 760
rect 18235 710 18265 740
rect 18235 690 18240 710
rect 18260 690 18265 710
rect 18235 660 18265 690
rect 18235 640 18240 660
rect 18260 640 18265 660
rect 18235 630 18265 640
rect 18325 910 18355 920
rect 18325 890 18330 910
rect 18350 890 18355 910
rect 18325 860 18355 890
rect 18325 840 18330 860
rect 18350 840 18355 860
rect 18325 810 18355 840
rect 18325 790 18330 810
rect 18350 790 18355 810
rect 18325 760 18355 790
rect 18325 740 18330 760
rect 18350 740 18355 760
rect 18325 710 18355 740
rect 18325 690 18330 710
rect 18350 690 18355 710
rect 18325 660 18355 690
rect 18325 640 18330 660
rect 18350 640 18355 660
rect 18325 630 18355 640
rect 18415 910 18445 920
rect 18415 890 18420 910
rect 18440 890 18445 910
rect 18415 860 18445 890
rect 18415 840 18420 860
rect 18440 840 18445 860
rect 18415 810 18445 840
rect 18415 790 18420 810
rect 18440 790 18445 810
rect 18415 760 18445 790
rect 18415 740 18420 760
rect 18440 740 18445 760
rect 18415 710 18445 740
rect 18415 690 18420 710
rect 18440 690 18445 710
rect 18415 660 18445 690
rect 18415 640 18420 660
rect 18440 640 18445 660
rect 18415 630 18445 640
rect 18505 910 18535 920
rect 18505 890 18510 910
rect 18530 890 18535 910
rect 18505 860 18535 890
rect 18505 840 18510 860
rect 18530 840 18535 860
rect 18505 810 18535 840
rect 18505 790 18510 810
rect 18530 790 18535 810
rect 18505 760 18535 790
rect 18505 740 18510 760
rect 18530 740 18535 760
rect 18505 710 18535 740
rect 18505 690 18510 710
rect 18530 690 18535 710
rect 18505 660 18535 690
rect 18505 640 18510 660
rect 18530 640 18535 660
rect 18505 630 18535 640
rect 18595 910 18665 920
rect 18595 890 18600 910
rect 18620 890 18640 910
rect 18660 890 18665 910
rect 18595 860 18665 890
rect 18595 840 18600 860
rect 18620 840 18640 860
rect 18660 840 18665 860
rect 18595 810 18665 840
rect 18595 790 18600 810
rect 18620 790 18640 810
rect 18660 790 18665 810
rect 18595 760 18665 790
rect 18595 740 18600 760
rect 18620 740 18640 760
rect 18660 740 18665 760
rect 18595 710 18665 740
rect 18870 910 18940 920
rect 18870 890 18875 910
rect 18895 890 18915 910
rect 18935 890 18940 910
rect 18870 860 18940 890
rect 18870 840 18875 860
rect 18895 840 18915 860
rect 18935 840 18940 860
rect 18870 810 18940 840
rect 18870 790 18875 810
rect 18895 790 18915 810
rect 18935 790 18940 810
rect 18870 760 18940 790
rect 18870 740 18875 760
rect 18895 740 18915 760
rect 18935 740 18940 760
rect 18870 730 18940 740
rect 18965 910 18995 920
rect 18965 890 18970 910
rect 18990 890 18995 910
rect 18965 860 18995 890
rect 18965 840 18970 860
rect 18990 840 18995 860
rect 18965 810 18995 840
rect 18965 790 18970 810
rect 18990 790 18995 810
rect 18965 760 18995 790
rect 18965 740 18970 760
rect 18990 740 18995 760
rect 18965 730 18995 740
rect 19020 910 19050 920
rect 19020 890 19025 910
rect 19045 890 19050 910
rect 19020 860 19050 890
rect 19020 840 19025 860
rect 19045 840 19050 860
rect 19020 810 19050 840
rect 19020 790 19025 810
rect 19045 790 19050 810
rect 19020 760 19050 790
rect 19020 740 19025 760
rect 19045 740 19050 760
rect 19020 730 19050 740
rect 19075 910 19145 920
rect 19075 890 19080 910
rect 19100 890 19120 910
rect 19140 890 19145 910
rect 19075 860 19145 890
rect 19075 840 19080 860
rect 19100 840 19120 860
rect 19140 840 19145 860
rect 19075 810 19145 840
rect 19075 790 19080 810
rect 19100 790 19120 810
rect 19140 790 19145 810
rect 19075 760 19145 790
rect 19075 740 19080 760
rect 19100 740 19120 760
rect 19140 740 19145 760
rect 19075 730 19145 740
rect 18970 710 18990 730
rect 18595 690 18600 710
rect 18620 690 18640 710
rect 18660 690 18665 710
rect 18595 660 18665 690
rect 18950 700 18990 710
rect 18950 680 18960 700
rect 18980 680 18990 700
rect 18950 670 18990 680
rect 18595 640 18600 660
rect 18620 640 18640 660
rect 18660 640 18665 660
rect 18595 630 18665 640
rect 19000 650 19040 655
rect 19000 630 19010 650
rect 19030 630 19040 650
rect 17070 610 17090 630
rect 17250 610 17270 630
rect 17430 610 17450 630
rect 17610 610 17630 630
rect 17790 610 17810 630
rect 17970 610 17990 630
rect 18150 610 18170 630
rect 18330 610 18350 630
rect 18510 610 18530 630
rect 19000 625 19040 630
rect 17060 600 17100 610
rect 17060 580 17070 600
rect 17090 580 17100 600
rect 17060 570 17100 580
rect 17240 600 17280 610
rect 17240 580 17250 600
rect 17270 580 17280 600
rect 17240 570 17280 580
rect 17420 600 17460 610
rect 17420 580 17430 600
rect 17450 580 17460 600
rect 17420 570 17460 580
rect 17600 600 17640 610
rect 17600 580 17610 600
rect 17630 580 17640 600
rect 17600 570 17640 580
rect 17690 600 17730 610
rect 17690 580 17700 600
rect 17720 580 17730 600
rect 17690 570 17730 580
rect 17780 600 17820 610
rect 17780 580 17790 600
rect 17810 580 17820 600
rect 17780 570 17820 580
rect 17960 600 18000 610
rect 17960 580 17970 600
rect 17990 580 18000 600
rect 17960 570 18000 580
rect 18140 600 18180 610
rect 18140 580 18150 600
rect 18170 580 18180 600
rect 18140 570 18180 580
rect 18320 600 18360 610
rect 18320 580 18330 600
rect 18350 580 18360 600
rect 18320 570 18360 580
rect 18410 600 18450 610
rect 18410 580 18420 600
rect 18440 580 18450 600
rect 18410 570 18450 580
rect 18500 600 18540 610
rect 18500 580 18510 600
rect 18530 580 18540 600
rect 18500 570 18540 580
rect 16425 130 16455 140
rect 16425 110 16430 130
rect 16450 110 16455 130
rect 16425 80 16455 110
rect 16480 130 16520 140
rect 16480 110 16490 130
rect 16510 110 16520 130
rect 16480 100 16520 110
rect 16545 130 16575 140
rect 16545 110 16550 130
rect 16570 110 16575 130
rect 16545 100 16575 110
rect 16665 130 16695 140
rect 16665 110 16670 130
rect 16690 110 16695 130
rect 16665 100 16695 110
rect 16785 130 16815 140
rect 16785 110 16790 130
rect 16810 110 16815 130
rect 16785 100 16815 110
rect 16840 130 16880 140
rect 16840 110 16850 130
rect 16870 110 16880 130
rect 16840 100 16880 110
rect 16905 130 16935 140
rect 16905 110 16910 130
rect 16930 110 16935 130
rect 16905 100 16935 110
rect 17025 130 17055 140
rect 17025 110 17030 130
rect 17050 110 17055 130
rect 17025 100 17055 110
rect 17145 130 17175 140
rect 17145 110 17150 130
rect 17170 110 17175 130
rect 17145 100 17175 110
rect 17200 130 17240 140
rect 17200 110 17210 130
rect 17230 110 17240 130
rect 17200 100 17240 110
rect 17265 130 17295 140
rect 17265 110 17270 130
rect 17290 110 17295 130
rect 17265 100 17295 110
rect 17385 130 17415 140
rect 17385 110 17390 130
rect 17410 110 17415 130
rect 17385 100 17415 110
rect 17505 130 17535 140
rect 17505 110 17510 130
rect 17530 110 17535 130
rect 17505 100 17535 110
rect 17560 130 17600 140
rect 17560 110 17570 130
rect 17590 110 17600 130
rect 17560 100 17600 110
rect 17625 130 17655 140
rect 17625 110 17630 130
rect 17650 110 17655 130
rect 16490 80 16510 100
rect 16550 80 16570 100
rect 16670 80 16690 100
rect 16790 80 16810 100
rect 16850 80 16870 100
rect 16910 80 16930 100
rect 17030 80 17050 100
rect 17150 80 17170 100
rect 17210 80 17230 100
rect 17270 80 17290 100
rect 17390 80 17410 100
rect 17510 80 17530 100
rect 17570 80 17590 100
rect 17625 80 17655 110
rect 17945 130 17975 140
rect 17945 110 17950 130
rect 17970 110 17975 130
rect 17945 80 17975 110
rect 18000 130 18040 140
rect 18000 110 18010 130
rect 18030 110 18040 130
rect 18000 100 18040 110
rect 18065 130 18095 140
rect 18065 110 18070 130
rect 18090 110 18095 130
rect 18065 100 18095 110
rect 18185 130 18215 140
rect 18185 110 18190 130
rect 18210 110 18215 130
rect 18185 100 18215 110
rect 18305 130 18335 140
rect 18305 110 18310 130
rect 18330 110 18335 130
rect 18305 100 18335 110
rect 18360 130 18400 140
rect 18360 110 18370 130
rect 18390 110 18400 130
rect 18360 100 18400 110
rect 18425 130 18455 140
rect 18425 110 18430 130
rect 18450 110 18455 130
rect 18425 100 18455 110
rect 18545 130 18575 140
rect 18545 110 18550 130
rect 18570 110 18575 130
rect 18545 100 18575 110
rect 18665 130 18695 140
rect 18665 110 18670 130
rect 18690 110 18695 130
rect 18665 100 18695 110
rect 18720 130 18760 140
rect 18720 110 18730 130
rect 18750 110 18760 130
rect 18720 100 18760 110
rect 18785 130 18815 140
rect 18785 110 18790 130
rect 18810 110 18815 130
rect 18785 100 18815 110
rect 18905 130 18935 140
rect 18905 110 18910 130
rect 18930 110 18935 130
rect 18905 100 18935 110
rect 19025 130 19055 140
rect 19025 110 19030 130
rect 19050 110 19055 130
rect 19025 100 19055 110
rect 19080 130 19120 140
rect 19080 110 19090 130
rect 19110 110 19120 130
rect 19080 100 19120 110
rect 19145 130 19175 140
rect 19145 110 19150 130
rect 19170 110 19175 130
rect 18010 80 18030 100
rect 18070 80 18090 100
rect 18190 80 18210 100
rect 18310 80 18330 100
rect 18370 80 18390 100
rect 18430 80 18450 100
rect 18550 80 18570 100
rect 18670 80 18690 100
rect 18730 80 18750 100
rect 18790 80 18810 100
rect 18910 80 18930 100
rect 19030 80 19050 100
rect 19090 80 19110 100
rect 19145 80 19175 110
rect 16385 70 16455 80
rect 16385 50 16390 70
rect 16410 50 16430 70
rect 16450 50 16455 70
rect 16385 20 16455 50
rect 16385 0 16390 20
rect 16410 0 16430 20
rect 16450 0 16455 20
rect 16385 -10 16455 0
rect 16485 70 16515 80
rect 16485 50 16490 70
rect 16510 50 16515 70
rect 16485 20 16515 50
rect 16485 0 16490 20
rect 16510 0 16515 20
rect 16485 -10 16515 0
rect 16545 70 16575 80
rect 16545 50 16550 70
rect 16570 50 16575 70
rect 16545 20 16575 50
rect 16545 0 16550 20
rect 16570 0 16575 20
rect 16545 -10 16575 0
rect 16605 70 16635 80
rect 16605 50 16610 70
rect 16630 50 16635 70
rect 16605 20 16635 50
rect 16605 0 16610 20
rect 16630 0 16635 20
rect 16605 -10 16635 0
rect 16665 70 16695 80
rect 16665 50 16670 70
rect 16690 50 16695 70
rect 16665 20 16695 50
rect 16665 0 16670 20
rect 16690 0 16695 20
rect 16665 -10 16695 0
rect 16725 70 16755 80
rect 16725 50 16730 70
rect 16750 50 16755 70
rect 16725 20 16755 50
rect 16725 0 16730 20
rect 16750 0 16755 20
rect 16725 -10 16755 0
rect 16785 70 16815 80
rect 16785 50 16790 70
rect 16810 50 16815 70
rect 16785 20 16815 50
rect 16785 0 16790 20
rect 16810 0 16815 20
rect 16785 -10 16815 0
rect 16845 70 16875 80
rect 16845 50 16850 70
rect 16870 50 16875 70
rect 16845 20 16875 50
rect 16845 0 16850 20
rect 16870 0 16875 20
rect 16845 -10 16875 0
rect 16905 70 16935 80
rect 16905 50 16910 70
rect 16930 50 16935 70
rect 16905 20 16935 50
rect 16905 0 16910 20
rect 16930 0 16935 20
rect 16905 -10 16935 0
rect 16965 70 16995 80
rect 16965 50 16970 70
rect 16990 50 16995 70
rect 16965 20 16995 50
rect 16965 0 16970 20
rect 16990 0 16995 20
rect 16965 -10 16995 0
rect 17025 70 17055 80
rect 17025 50 17030 70
rect 17050 50 17055 70
rect 17025 20 17055 50
rect 17025 0 17030 20
rect 17050 0 17055 20
rect 17025 -10 17055 0
rect 17085 70 17115 80
rect 17085 50 17090 70
rect 17110 50 17115 70
rect 17085 20 17115 50
rect 17085 0 17090 20
rect 17110 0 17115 20
rect 17085 -10 17115 0
rect 17145 70 17175 80
rect 17145 50 17150 70
rect 17170 50 17175 70
rect 17145 20 17175 50
rect 17145 0 17150 20
rect 17170 0 17175 20
rect 17145 -10 17175 0
rect 17205 70 17235 80
rect 17205 50 17210 70
rect 17230 50 17235 70
rect 17205 20 17235 50
rect 17205 0 17210 20
rect 17230 0 17235 20
rect 17205 -10 17235 0
rect 17265 70 17295 80
rect 17265 50 17270 70
rect 17290 50 17295 70
rect 17265 20 17295 50
rect 17265 0 17270 20
rect 17290 0 17295 20
rect 17265 -10 17295 0
rect 17325 70 17355 80
rect 17325 50 17330 70
rect 17350 50 17355 70
rect 17325 20 17355 50
rect 17325 0 17330 20
rect 17350 0 17355 20
rect 17325 -10 17355 0
rect 17385 70 17415 80
rect 17385 50 17390 70
rect 17410 50 17415 70
rect 17385 20 17415 50
rect 17385 0 17390 20
rect 17410 0 17415 20
rect 17385 -10 17415 0
rect 17445 70 17475 80
rect 17445 50 17450 70
rect 17470 50 17475 70
rect 17445 20 17475 50
rect 17445 0 17450 20
rect 17470 0 17475 20
rect 17445 -10 17475 0
rect 17505 70 17535 80
rect 17505 50 17510 70
rect 17530 50 17535 70
rect 17505 20 17535 50
rect 17505 0 17510 20
rect 17530 0 17535 20
rect 17505 -10 17535 0
rect 17565 70 17595 80
rect 17565 50 17570 70
rect 17590 50 17595 70
rect 17565 20 17595 50
rect 17565 0 17570 20
rect 17590 0 17595 20
rect 17565 -10 17595 0
rect 17625 70 17695 80
rect 17625 50 17630 70
rect 17650 50 17670 70
rect 17690 50 17695 70
rect 17625 20 17695 50
rect 17625 0 17630 20
rect 17650 0 17670 20
rect 17690 0 17695 20
rect 17625 -10 17695 0
rect 17905 70 17975 80
rect 17905 50 17910 70
rect 17930 50 17950 70
rect 17970 50 17975 70
rect 17905 20 17975 50
rect 17905 0 17910 20
rect 17930 0 17950 20
rect 17970 0 17975 20
rect 17905 -10 17975 0
rect 18005 70 18035 80
rect 18005 50 18010 70
rect 18030 50 18035 70
rect 18005 20 18035 50
rect 18005 0 18010 20
rect 18030 0 18035 20
rect 18005 -10 18035 0
rect 18065 70 18095 80
rect 18065 50 18070 70
rect 18090 50 18095 70
rect 18065 20 18095 50
rect 18065 0 18070 20
rect 18090 0 18095 20
rect 18065 -10 18095 0
rect 18125 70 18155 80
rect 18125 50 18130 70
rect 18150 50 18155 70
rect 18125 20 18155 50
rect 18125 0 18130 20
rect 18150 0 18155 20
rect 18125 -10 18155 0
rect 18185 70 18215 80
rect 18185 50 18190 70
rect 18210 50 18215 70
rect 18185 20 18215 50
rect 18185 0 18190 20
rect 18210 0 18215 20
rect 18185 -10 18215 0
rect 18245 70 18275 80
rect 18245 50 18250 70
rect 18270 50 18275 70
rect 18245 20 18275 50
rect 18245 0 18250 20
rect 18270 0 18275 20
rect 18245 -10 18275 0
rect 18305 70 18335 80
rect 18305 50 18310 70
rect 18330 50 18335 70
rect 18305 20 18335 50
rect 18305 0 18310 20
rect 18330 0 18335 20
rect 18305 -10 18335 0
rect 18365 70 18395 80
rect 18365 50 18370 70
rect 18390 50 18395 70
rect 18365 20 18395 50
rect 18365 0 18370 20
rect 18390 0 18395 20
rect 18365 -10 18395 0
rect 18425 70 18455 80
rect 18425 50 18430 70
rect 18450 50 18455 70
rect 18425 20 18455 50
rect 18425 0 18430 20
rect 18450 0 18455 20
rect 18425 -10 18455 0
rect 18485 70 18515 80
rect 18485 50 18490 70
rect 18510 50 18515 70
rect 18485 20 18515 50
rect 18485 0 18490 20
rect 18510 0 18515 20
rect 18485 -10 18515 0
rect 18545 70 18575 80
rect 18545 50 18550 70
rect 18570 50 18575 70
rect 18545 20 18575 50
rect 18545 0 18550 20
rect 18570 0 18575 20
rect 18545 -10 18575 0
rect 18605 70 18635 80
rect 18605 50 18610 70
rect 18630 50 18635 70
rect 18605 20 18635 50
rect 18605 0 18610 20
rect 18630 0 18635 20
rect 18605 -10 18635 0
rect 18665 70 18695 80
rect 18665 50 18670 70
rect 18690 50 18695 70
rect 18665 20 18695 50
rect 18665 0 18670 20
rect 18690 0 18695 20
rect 18665 -10 18695 0
rect 18725 70 18755 80
rect 18725 50 18730 70
rect 18750 50 18755 70
rect 18725 20 18755 50
rect 18725 0 18730 20
rect 18750 0 18755 20
rect 18725 -10 18755 0
rect 18785 70 18815 80
rect 18785 50 18790 70
rect 18810 50 18815 70
rect 18785 20 18815 50
rect 18785 0 18790 20
rect 18810 0 18815 20
rect 18785 -10 18815 0
rect 18845 70 18875 80
rect 18845 50 18850 70
rect 18870 50 18875 70
rect 18845 20 18875 50
rect 18845 0 18850 20
rect 18870 0 18875 20
rect 18845 -10 18875 0
rect 18905 70 18935 80
rect 18905 50 18910 70
rect 18930 50 18935 70
rect 18905 20 18935 50
rect 18905 0 18910 20
rect 18930 0 18935 20
rect 18905 -10 18935 0
rect 18965 70 18995 80
rect 18965 50 18970 70
rect 18990 50 18995 70
rect 18965 20 18995 50
rect 18965 0 18970 20
rect 18990 0 18995 20
rect 18965 -10 18995 0
rect 19025 70 19055 80
rect 19025 50 19030 70
rect 19050 50 19055 70
rect 19025 20 19055 50
rect 19025 0 19030 20
rect 19050 0 19055 20
rect 19025 -10 19055 0
rect 19085 70 19115 80
rect 19085 50 19090 70
rect 19110 50 19115 70
rect 19085 20 19115 50
rect 19085 0 19090 20
rect 19110 0 19115 20
rect 19085 -10 19115 0
rect 19145 70 19215 80
rect 19145 50 19150 70
rect 19170 50 19190 70
rect 19210 50 19215 70
rect 19145 20 19215 50
rect 19145 0 19150 20
rect 19170 0 19190 20
rect 19210 0 19215 20
rect 19145 -10 19215 0
rect 16425 -40 16455 -10
rect 16610 -30 16630 -10
rect 16730 -30 16750 -10
rect 16970 -30 16990 -10
rect 17090 -30 17110 -10
rect 17330 -30 17350 -10
rect 17450 -30 17470 -10
rect 16425 -60 16430 -40
rect 16450 -60 16455 -40
rect 16425 -70 16455 -60
rect 16510 -40 16550 -30
rect 16510 -60 16520 -40
rect 16540 -60 16550 -40
rect 16510 -70 16550 -60
rect 16600 -40 16640 -30
rect 16600 -60 16610 -40
rect 16630 -60 16640 -40
rect 16600 -70 16640 -60
rect 16720 -40 16760 -30
rect 16720 -60 16730 -40
rect 16750 -60 16760 -40
rect 16720 -70 16760 -60
rect 16840 -40 16880 -30
rect 16840 -60 16850 -40
rect 16870 -60 16880 -40
rect 16840 -70 16880 -60
rect 16960 -40 17000 -30
rect 16960 -60 16970 -40
rect 16990 -60 17000 -40
rect 16960 -70 17000 -60
rect 17080 -40 17120 -30
rect 17080 -60 17090 -40
rect 17110 -60 17120 -40
rect 17080 -70 17120 -60
rect 17200 -40 17240 -30
rect 17200 -60 17210 -40
rect 17230 -60 17240 -40
rect 17200 -70 17240 -60
rect 17320 -40 17360 -30
rect 17320 -60 17330 -40
rect 17350 -60 17360 -40
rect 17320 -70 17360 -60
rect 17440 -40 17480 -30
rect 17440 -60 17450 -40
rect 17470 -60 17480 -40
rect 17440 -70 17480 -60
rect 17535 -40 17565 -30
rect 17535 -60 17540 -40
rect 17560 -60 17565 -40
rect 17535 -70 17565 -60
rect 17945 -40 17975 -10
rect 18130 -30 18150 -10
rect 18250 -30 18270 -10
rect 18490 -30 18510 -10
rect 18610 -30 18630 -10
rect 18850 -30 18870 -10
rect 18970 -30 18990 -10
rect 19145 -15 19180 -10
rect 17945 -60 17950 -40
rect 17970 -60 17975 -40
rect 17945 -70 17975 -60
rect 18035 -40 18065 -30
rect 18035 -60 18040 -40
rect 18060 -60 18065 -40
rect 18035 -70 18065 -60
rect 18120 -40 18160 -30
rect 18120 -60 18130 -40
rect 18150 -60 18160 -40
rect 18120 -70 18160 -60
rect 18240 -40 18280 -30
rect 18240 -60 18250 -40
rect 18270 -60 18280 -40
rect 18240 -70 18280 -60
rect 18360 -40 18400 -30
rect 18360 -60 18370 -40
rect 18390 -60 18400 -40
rect 18360 -70 18400 -60
rect 18480 -40 18520 -30
rect 18480 -60 18490 -40
rect 18510 -60 18520 -40
rect 18480 -70 18520 -60
rect 18600 -40 18640 -30
rect 18600 -60 18610 -40
rect 18630 -60 18640 -40
rect 18600 -70 18640 -60
rect 18720 -40 18760 -30
rect 18720 -60 18730 -40
rect 18750 -60 18760 -40
rect 18720 -70 18760 -60
rect 18840 -40 18880 -30
rect 18840 -60 18850 -40
rect 18870 -60 18880 -40
rect 18840 -70 18880 -60
rect 18960 -40 19000 -30
rect 18960 -60 18970 -40
rect 18990 -60 19000 -40
rect 18960 -70 19000 -60
rect 19050 -40 19090 -30
rect 19050 -60 19060 -40
rect 19080 -60 19090 -40
rect 19050 -70 19090 -60
rect 19145 -40 19175 -15
rect 19145 -60 19150 -40
rect 19170 -60 19175 -40
rect 19145 -70 19175 -60
rect 16960 -155 16990 -145
rect 16960 -175 16965 -155
rect 16985 -175 16990 -155
rect 16960 -185 16990 -175
rect 17007 -155 17037 -145
rect 17007 -175 17012 -155
rect 17032 -175 17037 -155
rect 17007 -185 17037 -175
rect 17090 -155 17120 -145
rect 17090 -175 17095 -155
rect 17115 -175 17120 -155
rect 17090 -185 17120 -175
rect 18480 -155 18510 -145
rect 18480 -175 18485 -155
rect 18505 -175 18510 -155
rect 18480 -185 18510 -175
rect 18563 -155 18593 -145
rect 18563 -175 18568 -155
rect 18588 -175 18593 -155
rect 18563 -185 18593 -175
rect 18610 -155 18640 -145
rect 18610 -175 18615 -155
rect 18635 -175 18640 -155
rect 18610 -185 18640 -175
rect 16970 -205 16990 -185
rect 17090 -205 17110 -185
rect 18490 -205 18510 -185
rect 18610 -205 18630 -185
rect 16965 -215 16995 -205
rect 16965 -235 16970 -215
rect 16990 -235 16995 -215
rect 16965 -265 16995 -235
rect 16965 -285 16970 -265
rect 16990 -285 16995 -265
rect 16965 -315 16995 -285
rect 16965 -335 16970 -315
rect 16990 -335 16995 -315
rect 16965 -365 16995 -335
rect 16965 -385 16970 -365
rect 16990 -385 16995 -365
rect 16965 -415 16995 -385
rect 16965 -435 16970 -415
rect 16990 -435 16995 -415
rect 16965 -445 16995 -435
rect 17025 -215 17055 -205
rect 17025 -235 17030 -215
rect 17050 -235 17055 -215
rect 17025 -265 17055 -235
rect 17025 -285 17030 -265
rect 17050 -285 17055 -265
rect 17025 -315 17055 -285
rect 17025 -335 17030 -315
rect 17050 -335 17055 -315
rect 17025 -365 17055 -335
rect 17025 -385 17030 -365
rect 17050 -385 17055 -365
rect 17025 -415 17055 -385
rect 17025 -435 17030 -415
rect 17050 -435 17055 -415
rect 17025 -445 17055 -435
rect 17085 -215 17115 -205
rect 17085 -235 17090 -215
rect 17110 -235 17115 -215
rect 17085 -265 17115 -235
rect 17085 -285 17090 -265
rect 17110 -285 17115 -265
rect 17085 -315 17115 -285
rect 17085 -335 17090 -315
rect 17110 -335 17115 -315
rect 17560 -215 17600 -205
rect 17560 -235 17570 -215
rect 17590 -235 17600 -215
rect 17560 -255 17600 -235
rect 17560 -275 17570 -255
rect 17590 -275 17600 -255
rect 17560 -295 17600 -275
rect 17560 -315 17570 -295
rect 17590 -315 17600 -295
rect 17560 -325 17600 -315
rect 18000 -215 18040 -205
rect 18000 -235 18010 -215
rect 18030 -235 18040 -215
rect 18000 -255 18040 -235
rect 18000 -275 18010 -255
rect 18030 -275 18040 -255
rect 18000 -295 18040 -275
rect 18000 -315 18010 -295
rect 18030 -315 18040 -295
rect 18000 -325 18040 -315
rect 18485 -215 18515 -205
rect 18485 -235 18490 -215
rect 18510 -235 18515 -215
rect 18485 -265 18515 -235
rect 18485 -285 18490 -265
rect 18510 -285 18515 -265
rect 18485 -315 18515 -285
rect 17085 -365 17115 -335
rect 17085 -385 17090 -365
rect 17110 -385 17115 -365
rect 17085 -415 17115 -385
rect 17085 -435 17090 -415
rect 17110 -435 17115 -415
rect 17085 -445 17115 -435
rect 18485 -335 18490 -315
rect 18510 -335 18515 -315
rect 18485 -365 18515 -335
rect 18485 -385 18490 -365
rect 18510 -385 18515 -365
rect 18485 -415 18515 -385
rect 18485 -435 18490 -415
rect 18510 -435 18515 -415
rect 18485 -445 18515 -435
rect 18545 -215 18575 -205
rect 18545 -235 18550 -215
rect 18570 -235 18575 -215
rect 18545 -265 18575 -235
rect 18545 -285 18550 -265
rect 18570 -285 18575 -265
rect 18545 -315 18575 -285
rect 18545 -335 18550 -315
rect 18570 -335 18575 -315
rect 18545 -365 18575 -335
rect 18545 -385 18550 -365
rect 18570 -385 18575 -365
rect 18545 -415 18575 -385
rect 18545 -435 18550 -415
rect 18570 -435 18575 -415
rect 18545 -445 18575 -435
rect 18605 -215 18635 -205
rect 18605 -235 18610 -215
rect 18630 -235 18635 -215
rect 18605 -265 18635 -235
rect 18605 -285 18610 -265
rect 18630 -285 18635 -265
rect 18605 -315 18635 -285
rect 18605 -335 18610 -315
rect 18630 -335 18635 -315
rect 18605 -365 18635 -335
rect 18605 -385 18610 -365
rect 18630 -385 18635 -365
rect 18605 -415 18635 -385
rect 18605 -435 18610 -415
rect 18630 -435 18635 -415
rect 18605 -445 18635 -435
rect 18550 -465 18570 -445
rect 17075 -475 17105 -465
rect 17075 -495 17080 -475
rect 17100 -495 17105 -475
rect 17075 -505 17105 -495
rect 18495 -475 18525 -465
rect 18495 -495 18500 -475
rect 18520 -495 18525 -475
rect 18495 -505 18525 -495
rect 18545 -475 18575 -465
rect 18545 -495 18550 -475
rect 18570 -495 18575 -475
rect 18545 -505 18575 -495
rect 16620 -690 16660 -680
rect 16620 -710 16630 -690
rect 16650 -710 16660 -690
rect 16620 -720 16660 -710
rect 16740 -690 16780 -680
rect 16740 -710 16750 -690
rect 16770 -710 16780 -690
rect 16740 -720 16780 -710
rect 16860 -690 16900 -680
rect 16860 -710 16870 -690
rect 16890 -710 16900 -690
rect 16860 -720 16900 -710
rect 16980 -690 17020 -680
rect 16980 -710 16990 -690
rect 17010 -710 17020 -690
rect 16980 -720 17020 -710
rect 17300 -690 17340 -680
rect 17300 -710 17310 -690
rect 17330 -710 17340 -690
rect 17300 -720 17340 -710
rect 17420 -690 17460 -680
rect 17420 -710 17430 -690
rect 17450 -710 17460 -690
rect 17420 -720 17460 -710
rect 17540 -690 17580 -680
rect 17540 -710 17550 -690
rect 17570 -710 17580 -690
rect 18020 -690 18060 -680
rect 17540 -720 17580 -710
rect 17695 -705 17725 -695
rect 17695 -725 17700 -705
rect 17720 -725 17725 -705
rect 16535 -750 16565 -740
rect 16535 -770 16540 -750
rect 16560 -770 16565 -750
rect 16535 -800 16565 -770
rect 16535 -820 16540 -800
rect 16560 -820 16565 -800
rect 16535 -850 16565 -820
rect 16535 -870 16540 -850
rect 16560 -870 16565 -850
rect 16535 -900 16565 -870
rect 16535 -920 16540 -900
rect 16560 -920 16565 -900
rect 16535 -950 16565 -920
rect 16535 -970 16540 -950
rect 16560 -970 16565 -950
rect 16535 -980 16565 -970
rect 17075 -750 17185 -740
rect 17075 -770 17080 -750
rect 17100 -770 17120 -750
rect 17140 -770 17160 -750
rect 17180 -770 17185 -750
rect 17075 -800 17185 -770
rect 17075 -820 17080 -800
rect 17100 -820 17120 -800
rect 17140 -820 17160 -800
rect 17180 -820 17185 -800
rect 17075 -850 17185 -820
rect 17075 -870 17080 -850
rect 17100 -870 17120 -850
rect 17140 -870 17160 -850
rect 17180 -870 17185 -850
rect 17075 -900 17185 -870
rect 17075 -920 17080 -900
rect 17100 -920 17120 -900
rect 17140 -920 17160 -900
rect 17180 -920 17185 -900
rect 17075 -950 17185 -920
rect 17075 -970 17080 -950
rect 17100 -970 17120 -950
rect 17140 -970 17160 -950
rect 17180 -970 17185 -950
rect 17075 -980 17185 -970
rect 17695 -750 17725 -725
rect 17695 -770 17700 -750
rect 17720 -770 17725 -750
rect 17695 -800 17725 -770
rect 17695 -820 17700 -800
rect 17720 -820 17725 -800
rect 17695 -850 17725 -820
rect 17695 -870 17700 -850
rect 17720 -870 17725 -850
rect 17695 -900 17725 -870
rect 17695 -920 17700 -900
rect 17720 -920 17725 -900
rect 17695 -950 17725 -920
rect 17695 -970 17700 -950
rect 17720 -970 17725 -950
rect 17695 -980 17725 -970
rect 17875 -705 17905 -695
rect 17875 -725 17880 -705
rect 17900 -725 17905 -705
rect 18020 -710 18030 -690
rect 18050 -710 18060 -690
rect 18020 -720 18060 -710
rect 18140 -690 18180 -680
rect 18140 -710 18150 -690
rect 18170 -710 18180 -690
rect 18140 -720 18180 -710
rect 18260 -690 18300 -680
rect 18260 -710 18270 -690
rect 18290 -710 18300 -690
rect 18260 -720 18300 -710
rect 18580 -690 18620 -680
rect 18580 -710 18590 -690
rect 18610 -710 18620 -690
rect 18580 -720 18620 -710
rect 18700 -690 18740 -680
rect 18700 -710 18710 -690
rect 18730 -710 18740 -690
rect 18700 -720 18740 -710
rect 18820 -690 18860 -680
rect 18820 -710 18830 -690
rect 18850 -710 18860 -690
rect 18820 -720 18860 -710
rect 18940 -690 18980 -680
rect 18940 -710 18950 -690
rect 18970 -710 18980 -690
rect 18940 -720 18980 -710
rect 19030 -710 19070 -700
rect 17875 -750 17905 -725
rect 19030 -730 19040 -710
rect 19060 -730 19070 -710
rect 19030 -740 19070 -730
rect 17875 -770 17880 -750
rect 17900 -770 17905 -750
rect 17875 -800 17905 -770
rect 17875 -820 17880 -800
rect 17900 -820 17905 -800
rect 17875 -850 17905 -820
rect 17875 -870 17880 -850
rect 17900 -870 17905 -850
rect 17875 -900 17905 -870
rect 17875 -920 17880 -900
rect 17900 -920 17905 -900
rect 17875 -950 17905 -920
rect 17875 -970 17880 -950
rect 17900 -970 17905 -950
rect 17875 -980 17905 -970
rect 18415 -750 18525 -740
rect 18415 -770 18420 -750
rect 18440 -770 18460 -750
rect 18480 -770 18500 -750
rect 18520 -770 18525 -750
rect 18415 -800 18525 -770
rect 18415 -820 18420 -800
rect 18440 -820 18460 -800
rect 18480 -820 18500 -800
rect 18520 -820 18525 -800
rect 18415 -850 18525 -820
rect 18415 -870 18420 -850
rect 18440 -870 18460 -850
rect 18480 -870 18500 -850
rect 18520 -870 18525 -850
rect 18415 -900 18525 -870
rect 18415 -920 18420 -900
rect 18440 -920 18460 -900
rect 18480 -920 18500 -900
rect 18520 -920 18525 -900
rect 18415 -950 18525 -920
rect 18415 -970 18420 -950
rect 18440 -970 18460 -950
rect 18480 -970 18500 -950
rect 18520 -970 18525 -950
rect 18415 -980 18525 -970
rect 19035 -750 19065 -740
rect 19035 -770 19040 -750
rect 19060 -770 19065 -750
rect 19035 -800 19065 -770
rect 19035 -820 19040 -800
rect 19060 -820 19065 -800
rect 19035 -850 19065 -820
rect 19035 -870 19040 -850
rect 19060 -870 19065 -850
rect 19035 -900 19065 -870
rect 19035 -920 19040 -900
rect 19060 -920 19065 -900
rect 19035 -950 19065 -920
rect 19035 -970 19040 -950
rect 19060 -970 19065 -950
rect 19035 -980 19065 -970
rect 17120 -1000 17140 -980
rect 18460 -1000 18480 -980
rect 17110 -1010 17150 -1000
rect 17110 -1030 17120 -1010
rect 17140 -1030 17150 -1010
rect 17110 -1040 17150 -1030
rect 18450 -1010 18490 -1000
rect 18450 -1030 18460 -1010
rect 18480 -1030 18490 -1010
rect 18450 -1040 18490 -1030
rect 16740 -1145 16780 -1135
rect 16740 -1165 16750 -1145
rect 16770 -1165 16780 -1145
rect 16740 -1175 16780 -1165
rect 16820 -1145 16860 -1135
rect 16820 -1165 16830 -1145
rect 16850 -1165 16860 -1145
rect 16820 -1175 16860 -1165
rect 16900 -1145 16940 -1135
rect 16900 -1165 16910 -1145
rect 16930 -1165 16940 -1145
rect 16900 -1175 16940 -1165
rect 16980 -1145 17020 -1135
rect 16980 -1165 16990 -1145
rect 17010 -1165 17020 -1145
rect 16980 -1175 17020 -1165
rect 17060 -1145 17100 -1135
rect 17060 -1165 17070 -1145
rect 17090 -1165 17100 -1145
rect 17060 -1175 17100 -1165
rect 17140 -1145 17180 -1135
rect 17140 -1165 17150 -1145
rect 17170 -1165 17180 -1145
rect 17140 -1175 17180 -1165
rect 17220 -1145 17260 -1135
rect 17220 -1165 17230 -1145
rect 17250 -1165 17260 -1145
rect 17220 -1175 17260 -1165
rect 17300 -1145 17340 -1135
rect 17300 -1165 17310 -1145
rect 17330 -1165 17340 -1145
rect 17300 -1175 17340 -1165
rect 17380 -1145 17420 -1135
rect 17380 -1165 17390 -1145
rect 17410 -1165 17420 -1145
rect 17380 -1175 17420 -1165
rect 17460 -1145 17500 -1135
rect 17460 -1165 17470 -1145
rect 17490 -1165 17500 -1145
rect 17460 -1175 17500 -1165
rect 17540 -1145 17580 -1135
rect 17540 -1165 17550 -1145
rect 17570 -1165 17580 -1145
rect 17540 -1175 17580 -1165
rect 17620 -1145 17660 -1135
rect 17620 -1165 17630 -1145
rect 17650 -1165 17660 -1145
rect 17620 -1175 17660 -1165
rect 17700 -1145 17740 -1135
rect 17700 -1165 17710 -1145
rect 17730 -1165 17740 -1145
rect 17700 -1175 17740 -1165
rect 17780 -1145 17820 -1135
rect 17780 -1165 17790 -1145
rect 17810 -1165 17820 -1145
rect 17780 -1175 17820 -1165
rect 17860 -1145 17900 -1135
rect 17860 -1165 17870 -1145
rect 17890 -1165 17900 -1145
rect 17860 -1175 17900 -1165
rect 17940 -1145 17980 -1135
rect 17940 -1165 17950 -1145
rect 17970 -1165 17980 -1145
rect 17940 -1175 17980 -1165
rect 18020 -1145 18060 -1135
rect 18020 -1165 18030 -1145
rect 18050 -1165 18060 -1145
rect 18020 -1175 18060 -1165
rect 18100 -1145 18140 -1135
rect 18100 -1165 18110 -1145
rect 18130 -1165 18140 -1145
rect 18100 -1175 18140 -1165
rect 18180 -1145 18220 -1135
rect 18180 -1165 18190 -1145
rect 18210 -1165 18220 -1145
rect 18180 -1175 18220 -1165
rect 18260 -1145 18300 -1135
rect 18260 -1165 18270 -1145
rect 18290 -1165 18300 -1145
rect 18260 -1175 18300 -1165
rect 18340 -1145 18380 -1135
rect 18340 -1165 18350 -1145
rect 18370 -1165 18380 -1145
rect 18340 -1175 18380 -1165
rect 18420 -1145 18460 -1135
rect 18420 -1165 18430 -1145
rect 18450 -1165 18460 -1145
rect 18420 -1175 18460 -1165
rect 18500 -1145 18540 -1135
rect 18500 -1165 18510 -1145
rect 18530 -1165 18540 -1145
rect 18500 -1175 18540 -1165
rect 18580 -1145 18620 -1135
rect 18580 -1165 18590 -1145
rect 18610 -1165 18620 -1145
rect 18580 -1175 18620 -1165
rect 18660 -1145 18700 -1135
rect 18660 -1165 18670 -1145
rect 18690 -1165 18700 -1145
rect 18660 -1175 18700 -1165
rect 18740 -1145 18780 -1135
rect 18740 -1165 18750 -1145
rect 18770 -1165 18780 -1145
rect 18740 -1175 18780 -1165
rect 16750 -1195 16770 -1175
rect 17790 -1195 17810 -1175
rect 16745 -1205 16775 -1195
rect 16745 -1220 16750 -1205
rect 16700 -1225 16750 -1220
rect 16770 -1225 16775 -1205
rect 16700 -1230 16775 -1225
rect 16700 -1250 16710 -1230
rect 16730 -1250 16775 -1230
rect 16700 -1255 16775 -1250
rect 16700 -1260 16750 -1255
rect 16745 -1275 16750 -1260
rect 16770 -1275 16775 -1255
rect 16745 -1285 16775 -1275
rect 17785 -1205 17815 -1195
rect 17785 -1225 17790 -1205
rect 17810 -1225 17815 -1205
rect 17785 -1255 17815 -1225
rect 17785 -1275 17790 -1255
rect 17810 -1275 17815 -1255
rect 17785 -1285 17815 -1275
rect 18825 -1200 18895 -1195
rect 18825 -1205 18935 -1200
rect 18825 -1225 18830 -1205
rect 18850 -1225 18870 -1205
rect 18890 -1210 18935 -1205
rect 18890 -1225 18905 -1210
rect 18825 -1230 18905 -1225
rect 18925 -1230 18935 -1210
rect 18825 -1250 18935 -1230
rect 18825 -1255 18905 -1250
rect 18825 -1275 18830 -1255
rect 18850 -1275 18870 -1255
rect 18890 -1270 18905 -1255
rect 18925 -1270 18935 -1250
rect 18890 -1275 18935 -1270
rect 18825 -1280 18935 -1275
rect 18825 -1285 18895 -1280
rect 16540 -1495 16580 -1485
rect 16540 -1515 16550 -1495
rect 16570 -1515 16580 -1495
rect 16540 -1525 16580 -1515
rect 16600 -1495 16630 -1485
rect 16600 -1515 16605 -1495
rect 16625 -1515 16630 -1495
rect 16600 -1525 16630 -1515
rect 16650 -1495 16690 -1485
rect 16650 -1515 16660 -1495
rect 16680 -1515 16690 -1495
rect 16650 -1525 16690 -1515
rect 16710 -1495 16740 -1485
rect 16710 -1515 16715 -1495
rect 16735 -1515 16740 -1495
rect 16710 -1525 16740 -1515
rect 16760 -1495 16800 -1485
rect 16760 -1515 16770 -1495
rect 16790 -1515 16800 -1495
rect 16760 -1525 16800 -1515
rect 16820 -1495 16860 -1485
rect 16820 -1515 16830 -1495
rect 16850 -1515 16860 -1495
rect 16820 -1525 16860 -1515
rect 17025 -1495 17065 -1485
rect 17025 -1515 17035 -1495
rect 17055 -1515 17065 -1495
rect 17025 -1525 17065 -1515
rect 17135 -1495 17175 -1485
rect 17135 -1515 17145 -1495
rect 17165 -1515 17175 -1495
rect 17135 -1525 17175 -1515
rect 17245 -1495 17285 -1485
rect 17245 -1515 17255 -1495
rect 17275 -1515 17285 -1495
rect 17245 -1525 17285 -1515
rect 17305 -1495 17335 -1485
rect 17305 -1515 17310 -1495
rect 17330 -1515 17335 -1495
rect 17305 -1525 17335 -1515
rect 17355 -1495 17395 -1485
rect 17355 -1515 17365 -1495
rect 17385 -1515 17395 -1495
rect 17355 -1525 17395 -1515
rect 17465 -1495 17505 -1485
rect 17465 -1515 17475 -1495
rect 17495 -1515 17505 -1495
rect 17465 -1525 17505 -1515
rect 17615 -1495 17655 -1485
rect 17615 -1515 17625 -1495
rect 17645 -1515 17655 -1495
rect 17615 -1525 17655 -1515
rect 17725 -1495 17765 -1485
rect 17725 -1515 17735 -1495
rect 17755 -1515 17765 -1495
rect 17725 -1525 17765 -1515
rect 17785 -1495 17815 -1485
rect 17785 -1515 17790 -1495
rect 17810 -1515 17815 -1495
rect 17785 -1525 17815 -1515
rect 17835 -1495 17875 -1485
rect 17835 -1515 17845 -1495
rect 17865 -1515 17875 -1495
rect 17835 -1525 17875 -1515
rect 17945 -1495 17985 -1485
rect 17945 -1515 17955 -1495
rect 17975 -1515 17985 -1495
rect 17945 -1525 17985 -1515
rect 18095 -1495 18135 -1485
rect 18095 -1515 18105 -1495
rect 18125 -1515 18135 -1495
rect 18095 -1525 18135 -1515
rect 18205 -1495 18245 -1485
rect 18205 -1515 18215 -1495
rect 18235 -1515 18245 -1495
rect 18205 -1525 18245 -1515
rect 18265 -1495 18295 -1485
rect 18265 -1515 18270 -1495
rect 18290 -1515 18295 -1495
rect 18265 -1525 18295 -1515
rect 18315 -1495 18355 -1485
rect 18315 -1515 18325 -1495
rect 18345 -1515 18355 -1495
rect 18315 -1525 18355 -1515
rect 18425 -1495 18465 -1485
rect 18425 -1515 18435 -1495
rect 18455 -1515 18465 -1495
rect 18425 -1525 18465 -1515
rect 18535 -1495 18575 -1485
rect 18535 -1515 18545 -1495
rect 18565 -1515 18575 -1495
rect 18535 -1525 18575 -1515
rect 16545 -1545 16575 -1525
rect 16605 -1545 16625 -1525
rect 16660 -1545 16680 -1525
rect 16770 -1545 16790 -1525
rect 16820 -1545 16850 -1525
rect 17030 -1545 17060 -1525
rect 17145 -1545 17165 -1525
rect 17255 -1545 17275 -1525
rect 17365 -1545 17385 -1525
rect 17470 -1545 17500 -1525
rect 17620 -1545 17650 -1525
rect 17735 -1545 17755 -1525
rect 17845 -1545 17865 -1525
rect 17950 -1545 17980 -1525
rect 18100 -1545 18130 -1525
rect 18215 -1545 18235 -1525
rect 18325 -1545 18345 -1525
rect 18435 -1545 18455 -1525
rect 18540 -1545 18570 -1525
rect 16505 -1555 16575 -1545
rect 16505 -1575 16510 -1555
rect 16530 -1575 16550 -1555
rect 16570 -1575 16575 -1555
rect 16505 -1605 16575 -1575
rect 16505 -1625 16510 -1605
rect 16530 -1625 16550 -1605
rect 16570 -1625 16575 -1605
rect 16505 -1635 16575 -1625
rect 16600 -1555 16630 -1545
rect 16600 -1575 16605 -1555
rect 16625 -1575 16630 -1555
rect 16600 -1605 16630 -1575
rect 16600 -1625 16605 -1605
rect 16625 -1625 16630 -1605
rect 16600 -1635 16630 -1625
rect 16655 -1555 16685 -1545
rect 16655 -1575 16660 -1555
rect 16680 -1575 16685 -1555
rect 16655 -1605 16685 -1575
rect 16655 -1625 16660 -1605
rect 16680 -1625 16685 -1605
rect 16655 -1635 16685 -1625
rect 16710 -1555 16740 -1545
rect 16710 -1575 16715 -1555
rect 16735 -1575 16740 -1555
rect 16710 -1605 16740 -1575
rect 16710 -1625 16715 -1605
rect 16735 -1625 16740 -1605
rect 16710 -1635 16740 -1625
rect 16765 -1555 16795 -1545
rect 16765 -1575 16770 -1555
rect 16790 -1575 16795 -1555
rect 16765 -1605 16795 -1575
rect 16765 -1625 16770 -1605
rect 16790 -1625 16795 -1605
rect 16765 -1635 16795 -1625
rect 16820 -1555 16890 -1545
rect 16820 -1575 16825 -1555
rect 16845 -1575 16865 -1555
rect 16885 -1575 16890 -1555
rect 16820 -1605 16890 -1575
rect 16820 -1625 16825 -1605
rect 16845 -1625 16865 -1605
rect 16885 -1625 16890 -1605
rect 16820 -1635 16890 -1625
rect 16990 -1555 17060 -1545
rect 16990 -1575 16995 -1555
rect 17015 -1575 17035 -1555
rect 17055 -1575 17060 -1555
rect 16990 -1605 17060 -1575
rect 16990 -1625 16995 -1605
rect 17015 -1625 17035 -1605
rect 17055 -1625 17060 -1605
rect 16990 -1635 17060 -1625
rect 17085 -1555 17115 -1545
rect 17085 -1575 17090 -1555
rect 17110 -1575 17115 -1555
rect 17085 -1605 17115 -1575
rect 17085 -1625 17090 -1605
rect 17110 -1625 17115 -1605
rect 17085 -1635 17115 -1625
rect 17140 -1555 17170 -1545
rect 17140 -1575 17145 -1555
rect 17165 -1575 17170 -1555
rect 17140 -1605 17170 -1575
rect 17140 -1625 17145 -1605
rect 17165 -1625 17170 -1605
rect 17140 -1635 17170 -1625
rect 17195 -1555 17225 -1545
rect 17195 -1575 17200 -1555
rect 17220 -1575 17225 -1555
rect 17195 -1605 17225 -1575
rect 17195 -1625 17200 -1605
rect 17220 -1625 17225 -1605
rect 17195 -1635 17225 -1625
rect 17250 -1555 17280 -1545
rect 17250 -1575 17255 -1555
rect 17275 -1575 17280 -1555
rect 17250 -1605 17280 -1575
rect 17250 -1625 17255 -1605
rect 17275 -1625 17280 -1605
rect 17250 -1635 17280 -1625
rect 17305 -1555 17335 -1545
rect 17305 -1575 17310 -1555
rect 17330 -1575 17335 -1555
rect 17305 -1605 17335 -1575
rect 17305 -1625 17310 -1605
rect 17330 -1625 17335 -1605
rect 17305 -1635 17335 -1625
rect 17360 -1555 17390 -1545
rect 17360 -1575 17365 -1555
rect 17385 -1575 17390 -1555
rect 17360 -1605 17390 -1575
rect 17360 -1625 17365 -1605
rect 17385 -1625 17390 -1605
rect 17360 -1635 17390 -1625
rect 17415 -1555 17445 -1545
rect 17415 -1575 17420 -1555
rect 17440 -1575 17445 -1555
rect 17415 -1605 17445 -1575
rect 17415 -1625 17420 -1605
rect 17440 -1625 17445 -1605
rect 17415 -1635 17445 -1625
rect 17470 -1555 17540 -1545
rect 17470 -1575 17475 -1555
rect 17495 -1575 17515 -1555
rect 17535 -1575 17540 -1555
rect 17470 -1605 17540 -1575
rect 17470 -1625 17475 -1605
rect 17495 -1625 17515 -1605
rect 17535 -1625 17540 -1605
rect 17470 -1635 17540 -1625
rect 17580 -1555 17650 -1545
rect 17580 -1575 17585 -1555
rect 17605 -1575 17625 -1555
rect 17645 -1575 17650 -1555
rect 17580 -1605 17650 -1575
rect 17580 -1625 17585 -1605
rect 17605 -1625 17625 -1605
rect 17645 -1625 17650 -1605
rect 17580 -1635 17650 -1625
rect 17675 -1555 17705 -1545
rect 17675 -1575 17680 -1555
rect 17700 -1575 17705 -1555
rect 17675 -1605 17705 -1575
rect 17675 -1625 17680 -1605
rect 17700 -1625 17705 -1605
rect 17675 -1635 17705 -1625
rect 17730 -1555 17760 -1545
rect 17730 -1575 17735 -1555
rect 17755 -1575 17760 -1555
rect 17730 -1605 17760 -1575
rect 17730 -1625 17735 -1605
rect 17755 -1625 17760 -1605
rect 17730 -1635 17760 -1625
rect 17785 -1555 17815 -1545
rect 17785 -1575 17790 -1555
rect 17810 -1575 17815 -1555
rect 17785 -1605 17815 -1575
rect 17785 -1625 17790 -1605
rect 17810 -1625 17815 -1605
rect 17785 -1635 17815 -1625
rect 17840 -1555 17870 -1545
rect 17840 -1575 17845 -1555
rect 17865 -1575 17870 -1555
rect 17840 -1605 17870 -1575
rect 17840 -1625 17845 -1605
rect 17865 -1625 17870 -1605
rect 17840 -1635 17870 -1625
rect 17895 -1555 17925 -1545
rect 17895 -1575 17900 -1555
rect 17920 -1575 17925 -1555
rect 17895 -1605 17925 -1575
rect 17895 -1625 17900 -1605
rect 17920 -1625 17925 -1605
rect 17895 -1635 17925 -1625
rect 17950 -1555 18020 -1545
rect 17950 -1575 17955 -1555
rect 17975 -1575 17995 -1555
rect 18015 -1575 18020 -1555
rect 17950 -1605 18020 -1575
rect 17950 -1625 17955 -1605
rect 17975 -1625 17995 -1605
rect 18015 -1625 18020 -1605
rect 17950 -1635 18020 -1625
rect 18060 -1555 18130 -1545
rect 18060 -1575 18065 -1555
rect 18085 -1575 18105 -1555
rect 18125 -1575 18130 -1555
rect 18060 -1605 18130 -1575
rect 18060 -1625 18065 -1605
rect 18085 -1625 18105 -1605
rect 18125 -1625 18130 -1605
rect 18060 -1635 18130 -1625
rect 18155 -1555 18185 -1545
rect 18155 -1575 18160 -1555
rect 18180 -1575 18185 -1555
rect 18155 -1605 18185 -1575
rect 18155 -1625 18160 -1605
rect 18180 -1625 18185 -1605
rect 18155 -1635 18185 -1625
rect 18210 -1555 18240 -1545
rect 18210 -1575 18215 -1555
rect 18235 -1575 18240 -1555
rect 18210 -1605 18240 -1575
rect 18210 -1625 18215 -1605
rect 18235 -1625 18240 -1605
rect 18210 -1635 18240 -1625
rect 18265 -1555 18295 -1545
rect 18265 -1575 18270 -1555
rect 18290 -1575 18295 -1555
rect 18265 -1605 18295 -1575
rect 18265 -1625 18270 -1605
rect 18290 -1625 18295 -1605
rect 18265 -1635 18295 -1625
rect 18320 -1555 18350 -1545
rect 18320 -1575 18325 -1555
rect 18345 -1575 18350 -1555
rect 18320 -1605 18350 -1575
rect 18320 -1625 18325 -1605
rect 18345 -1625 18350 -1605
rect 18320 -1635 18350 -1625
rect 18375 -1555 18405 -1545
rect 18375 -1575 18380 -1555
rect 18400 -1575 18405 -1555
rect 18375 -1605 18405 -1575
rect 18375 -1625 18380 -1605
rect 18400 -1625 18405 -1605
rect 18375 -1635 18405 -1625
rect 18430 -1555 18460 -1545
rect 18430 -1575 18435 -1555
rect 18455 -1575 18460 -1555
rect 18430 -1605 18460 -1575
rect 18430 -1625 18435 -1605
rect 18455 -1625 18460 -1605
rect 18430 -1635 18460 -1625
rect 18485 -1555 18515 -1545
rect 18485 -1575 18490 -1555
rect 18510 -1575 18515 -1555
rect 18485 -1605 18515 -1575
rect 18485 -1625 18490 -1605
rect 18510 -1625 18515 -1605
rect 18485 -1635 18515 -1625
rect 18540 -1555 18610 -1545
rect 18540 -1575 18545 -1555
rect 18565 -1575 18585 -1555
rect 18605 -1575 18610 -1555
rect 18540 -1605 18610 -1575
rect 18540 -1625 18545 -1605
rect 18565 -1625 18585 -1605
rect 18605 -1625 18610 -1605
rect 18540 -1635 18610 -1625
rect 16715 -1655 16735 -1635
rect 17090 -1655 17110 -1635
rect 17310 -1655 17330 -1635
rect 17680 -1655 17700 -1635
rect 17790 -1655 17810 -1635
rect 17900 -1655 17920 -1635
rect 18270 -1655 18290 -1635
rect 18490 -1655 18510 -1635
rect 16705 -1665 16745 -1655
rect 16705 -1685 16715 -1665
rect 16735 -1685 16745 -1665
rect 16705 -1695 16745 -1685
rect 17080 -1665 17120 -1655
rect 17080 -1685 17090 -1665
rect 17110 -1685 17120 -1665
rect 17080 -1695 17120 -1685
rect 17190 -1665 17230 -1655
rect 17190 -1685 17200 -1665
rect 17220 -1685 17230 -1665
rect 17190 -1695 17230 -1685
rect 17300 -1665 17340 -1655
rect 17300 -1685 17310 -1665
rect 17330 -1685 17340 -1665
rect 17300 -1695 17340 -1685
rect 17410 -1665 17450 -1655
rect 17410 -1685 17420 -1665
rect 17440 -1685 17450 -1665
rect 17410 -1695 17450 -1685
rect 17670 -1665 17710 -1655
rect 17670 -1685 17680 -1665
rect 17700 -1685 17710 -1665
rect 17670 -1695 17710 -1685
rect 17780 -1665 17820 -1655
rect 17780 -1685 17790 -1665
rect 17810 -1685 17820 -1665
rect 17780 -1695 17820 -1685
rect 17890 -1665 17930 -1655
rect 17890 -1685 17900 -1665
rect 17920 -1685 17930 -1665
rect 17890 -1695 17930 -1685
rect 18150 -1665 18190 -1655
rect 18150 -1685 18160 -1665
rect 18180 -1685 18190 -1665
rect 18150 -1695 18190 -1685
rect 18260 -1665 18300 -1655
rect 18260 -1685 18270 -1665
rect 18290 -1685 18300 -1665
rect 18260 -1695 18300 -1685
rect 18370 -1665 18410 -1655
rect 18370 -1685 18380 -1665
rect 18400 -1685 18410 -1665
rect 18370 -1695 18410 -1685
rect 18480 -1665 18520 -1655
rect 18480 -1685 18490 -1665
rect 18510 -1685 18520 -1665
rect 18480 -1695 18520 -1685
rect 17425 -2005 17470 -2000
rect 17425 -2030 17435 -2005
rect 17460 -2030 17470 -2005
rect 17425 -2035 17470 -2030
rect 18124 -2005 18169 -2000
rect 18124 -2030 18134 -2005
rect 18159 -2030 18169 -2005
rect 18124 -2035 18169 -2030
rect 16795 -2240 18805 -2115
rect 17440 -2795 17480 -2240
rect 18120 -2795 18160 -2240
rect 16485 -2905 16520 -2895
rect 16485 -2930 16490 -2905
rect 16515 -2930 16520 -2905
rect 16795 -2920 18805 -2795
rect 19080 -2905 19115 -2895
rect 16485 -2940 16520 -2930
rect 16160 -3030 16195 -3020
rect 16160 -3055 16165 -3030
rect 16190 -3055 16195 -3030
rect 16160 -3065 16195 -3055
rect 15950 -3121 15985 -3111
rect 15950 -3146 15955 -3121
rect 15980 -3146 15985 -3121
rect 15950 -3156 15985 -3146
rect 16255 -3100 16280 -3065
rect 16580 -2975 16605 -2940
rect 17440 -3475 17480 -2920
rect 18120 -3475 18160 -2920
rect 19080 -2930 19085 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2940 19115 -2930
rect 18995 -2975 19020 -2940
rect 19405 -3002 19440 -2992
rect 19405 -3027 19410 -3002
rect 19435 -3027 19440 -3002
rect 19405 -3037 19440 -3027
rect 19320 -3072 19345 -3037
rect 19610 -3121 19645 -3111
rect 19610 -3146 19615 -3121
rect 19640 -3146 19645 -3121
rect 19610 -3156 19645 -3146
rect 16795 -3600 18805 -3475
rect 15950 -3794 15985 -3784
rect 15950 -3819 15955 -3794
rect 15980 -3819 15985 -3794
rect 15950 -3829 15985 -3819
rect 16195 -3889 16220 -3854
rect 16280 -3899 16315 -3889
rect 16280 -3924 16285 -3899
rect 16310 -3924 16315 -3899
rect 16280 -3934 16315 -3924
rect 16520 -3964 16545 -3929
rect 16605 -3974 16640 -3964
rect 16605 -3999 16610 -3974
rect 16635 -3999 16640 -3974
rect 16605 -4009 16640 -3999
rect 17440 -4125 17480 -3600
rect 17780 -4170 17820 -4120
rect 18120 -4125 18160 -3600
rect 19055 -3964 19080 -3929
rect 19380 -3889 19405 -3854
rect 19610 -3794 19645 -3784
rect 19610 -3819 19615 -3794
rect 19640 -3819 19645 -3794
rect 19610 -3829 19645 -3819
rect 19285 -3899 19320 -3889
rect 19285 -3924 19290 -3899
rect 19315 -3924 19320 -3899
rect 19285 -3934 19320 -3924
rect 18960 -3974 18995 -3964
rect 18960 -3999 18965 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4009 18995 -3999
rect 17780 -4190 17790 -4170
rect 17810 -4190 17820 -4170
rect 17780 -4220 17820 -4190
rect 17780 -4240 17790 -4220
rect 17810 -4240 17820 -4220
rect 17780 -4270 17820 -4240
rect 17780 -4290 17790 -4270
rect 17810 -4290 17820 -4270
rect 17780 -4300 17820 -4290
<< viali >>
rect 16495 1595 16515 1615
rect 17790 1595 17810 1615
rect 16375 1415 16395 1435
rect 16495 1415 16515 1435
rect 16615 1415 16635 1435
rect 16895 1415 16915 1435
rect 16950 1415 16970 1435
rect 17005 1415 17025 1435
rect 17060 1415 17080 1435
rect 17115 1415 17135 1435
rect 17225 1415 17245 1435
rect 17505 1415 17525 1435
rect 17570 1415 17590 1435
rect 17625 1415 17645 1435
rect 17680 1415 17700 1435
rect 17735 1415 17755 1435
rect 17790 1415 17810 1435
rect 17845 1415 17865 1435
rect 17900 1415 17920 1435
rect 17955 1415 17975 1435
rect 18010 1415 18030 1435
rect 18075 1415 18095 1435
rect 18355 1415 18375 1435
rect 18465 1415 18485 1435
rect 18520 1415 18540 1435
rect 18575 1415 18595 1435
rect 18630 1415 18650 1435
rect 18685 1415 18705 1435
rect 16440 1245 16460 1265
rect 16550 1245 16570 1265
rect 16950 1245 16970 1265
rect 17060 1245 17080 1265
rect 17170 1245 17190 1265
rect 17625 1245 17645 1265
rect 17735 1245 17755 1265
rect 17845 1245 17865 1265
rect 17955 1245 17975 1265
rect 18410 1245 18430 1265
rect 18520 1245 18540 1265
rect 18630 1245 18650 1265
rect 16980 950 17000 970
rect 17160 950 17180 970
rect 17340 950 17360 970
rect 17520 950 17540 970
rect 17700 950 17720 970
rect 17880 950 17900 970
rect 18060 950 18080 970
rect 18240 950 18260 970
rect 18420 950 18440 970
rect 18600 950 18620 970
rect 18915 950 18935 970
rect 19025 950 19045 970
rect 19085 950 19105 970
rect 16445 850 16465 870
rect 16555 850 16575 870
rect 16665 850 16685 870
rect 16490 680 16510 700
rect 16555 680 16575 700
rect 16620 680 16640 700
rect 18960 680 18980 700
rect 19010 630 19030 650
rect 17070 580 17090 600
rect 17250 580 17270 600
rect 17430 580 17450 600
rect 17610 580 17630 600
rect 17700 580 17720 600
rect 17790 580 17810 600
rect 17970 580 17990 600
rect 18150 580 18170 600
rect 18330 580 18350 600
rect 18420 580 18440 600
rect 18510 580 18530 600
rect 16430 110 16450 130
rect 16490 110 16510 130
rect 16550 110 16570 130
rect 16670 110 16690 130
rect 16790 110 16810 130
rect 16850 110 16870 130
rect 16910 110 16930 130
rect 17030 110 17050 130
rect 17150 110 17170 130
rect 17210 110 17230 130
rect 17270 110 17290 130
rect 17390 110 17410 130
rect 17510 110 17530 130
rect 17570 110 17590 130
rect 17630 110 17650 130
rect 17950 110 17970 130
rect 18010 110 18030 130
rect 18070 110 18090 130
rect 18190 110 18210 130
rect 18310 110 18330 130
rect 18370 110 18390 130
rect 18430 110 18450 130
rect 18550 110 18570 130
rect 18670 110 18690 130
rect 18730 110 18750 130
rect 18790 110 18810 130
rect 18910 110 18930 130
rect 19030 110 19050 130
rect 19090 110 19110 130
rect 19150 110 19170 130
rect 16520 -60 16540 -40
rect 16610 -60 16630 -40
rect 16730 -60 16750 -40
rect 16850 -60 16870 -40
rect 16970 -60 16990 -40
rect 17090 -60 17110 -40
rect 17210 -60 17230 -40
rect 17330 -60 17350 -40
rect 17450 -60 17470 -40
rect 17540 -60 17560 -40
rect 18040 -60 18060 -40
rect 18130 -60 18150 -40
rect 18250 -60 18270 -40
rect 18370 -60 18390 -40
rect 18490 -60 18510 -40
rect 18610 -60 18630 -40
rect 18730 -60 18750 -40
rect 18850 -60 18870 -40
rect 18970 -60 18990 -40
rect 19060 -60 19080 -40
rect 16965 -175 16985 -155
rect 17012 -175 17032 -155
rect 17095 -175 17115 -155
rect 18485 -175 18505 -155
rect 18568 -175 18588 -155
rect 18615 -175 18635 -155
rect 17030 -235 17050 -215
rect 17030 -285 17050 -265
rect 17030 -335 17050 -315
rect 17030 -385 17050 -365
rect 17030 -435 17050 -415
rect 17570 -235 17590 -215
rect 17570 -275 17590 -255
rect 17570 -315 17590 -295
rect 18010 -235 18030 -215
rect 18010 -275 18030 -255
rect 18010 -315 18030 -295
rect 17080 -495 17100 -475
rect 18500 -495 18520 -475
rect 18550 -495 18570 -475
rect 16630 -710 16650 -690
rect 16750 -710 16770 -690
rect 16870 -710 16890 -690
rect 16990 -710 17010 -690
rect 17310 -710 17330 -690
rect 17430 -710 17450 -690
rect 17550 -710 17570 -690
rect 17700 -725 17720 -705
rect 16540 -770 16560 -750
rect 16540 -820 16560 -800
rect 16540 -870 16560 -850
rect 16540 -920 16560 -900
rect 16540 -970 16560 -950
rect 17880 -725 17900 -705
rect 18030 -710 18050 -690
rect 18150 -710 18170 -690
rect 18270 -710 18290 -690
rect 18590 -710 18610 -690
rect 18710 -710 18730 -690
rect 18830 -710 18850 -690
rect 18950 -710 18970 -690
rect 19040 -730 19060 -710
rect 17120 -1030 17140 -1010
rect 18460 -1030 18480 -1010
rect 16750 -1165 16770 -1145
rect 16830 -1165 16850 -1145
rect 16910 -1165 16930 -1145
rect 16990 -1165 17010 -1145
rect 17070 -1165 17090 -1145
rect 17150 -1165 17170 -1145
rect 17230 -1165 17250 -1145
rect 17310 -1165 17330 -1145
rect 17390 -1165 17410 -1145
rect 17470 -1165 17490 -1145
rect 17550 -1165 17570 -1145
rect 17630 -1165 17650 -1145
rect 17710 -1165 17730 -1145
rect 17790 -1165 17810 -1145
rect 17870 -1165 17890 -1145
rect 17950 -1165 17970 -1145
rect 18030 -1165 18050 -1145
rect 18110 -1165 18130 -1145
rect 18190 -1165 18210 -1145
rect 18270 -1165 18290 -1145
rect 18350 -1165 18370 -1145
rect 18430 -1165 18450 -1145
rect 18510 -1165 18530 -1145
rect 18590 -1165 18610 -1145
rect 18670 -1165 18690 -1145
rect 18750 -1165 18770 -1145
rect 16710 -1250 16730 -1230
rect 18905 -1230 18925 -1210
rect 18905 -1270 18925 -1250
rect 16550 -1515 16570 -1495
rect 16605 -1515 16625 -1495
rect 16660 -1515 16680 -1495
rect 16715 -1515 16735 -1495
rect 16770 -1515 16790 -1495
rect 16830 -1515 16850 -1495
rect 17035 -1515 17055 -1495
rect 17145 -1515 17165 -1495
rect 17255 -1515 17275 -1495
rect 17310 -1515 17330 -1495
rect 17365 -1515 17385 -1495
rect 17475 -1515 17495 -1495
rect 17625 -1515 17645 -1495
rect 17735 -1515 17755 -1495
rect 17790 -1515 17810 -1495
rect 17845 -1515 17865 -1495
rect 17955 -1515 17975 -1495
rect 18105 -1515 18125 -1495
rect 18215 -1515 18235 -1495
rect 18270 -1515 18290 -1495
rect 18325 -1515 18345 -1495
rect 18435 -1515 18455 -1495
rect 18545 -1515 18565 -1495
rect 17200 -1575 17220 -1555
rect 17200 -1625 17220 -1605
rect 17420 -1575 17440 -1555
rect 17420 -1625 17440 -1605
rect 18160 -1575 18180 -1555
rect 18160 -1625 18180 -1605
rect 18380 -1575 18400 -1555
rect 18380 -1625 18400 -1605
rect 16715 -1685 16735 -1665
rect 17090 -1685 17110 -1665
rect 17200 -1685 17220 -1665
rect 17310 -1685 17330 -1665
rect 17420 -1685 17440 -1665
rect 17680 -1685 17700 -1665
rect 17790 -1685 17810 -1665
rect 17900 -1685 17920 -1665
rect 18160 -1685 18180 -1665
rect 18270 -1685 18290 -1665
rect 18380 -1685 18400 -1665
rect 18490 -1685 18510 -1665
rect 17435 -2030 17460 -2005
rect 18134 -2030 18159 -2005
rect 16490 -2930 16515 -2905
rect 16165 -3055 16190 -3030
rect 15955 -3146 15980 -3121
rect 19085 -2930 19110 -2905
rect 19410 -3027 19435 -3002
rect 19615 -3146 19640 -3121
rect 15955 -3819 15980 -3794
rect 16285 -3924 16310 -3899
rect 16610 -3999 16635 -3974
rect 19615 -3819 19640 -3794
rect 19290 -3924 19315 -3899
rect 18965 -3999 18990 -3974
rect 17790 -4290 17810 -4270
<< metal1 >>
rect 15725 -95 15765 -90
rect 15725 -125 15730 -95
rect 15760 -125 15765 -95
rect 15725 -130 15765 -125
rect 15735 -4310 15755 -130
rect 15785 -1770 15825 1755
rect 15950 135 15990 140
rect 15950 105 15955 135
rect 15985 105 15990 135
rect 15950 100 15990 105
rect 15785 -1800 15790 -1770
rect 15820 -1800 15825 -1770
rect 15785 -1810 15825 -1800
rect 15785 -1840 15790 -1810
rect 15820 -1840 15825 -1810
rect 15785 -1845 15825 -1840
rect 15820 -3115 15860 -3110
rect 15960 -3111 15980 100
rect 16040 -1710 16060 1755
rect 16030 -1715 16070 -1710
rect 16030 -1745 16035 -1715
rect 16065 -1745 16070 -1715
rect 16030 -1750 16070 -1745
rect 16115 -1895 16135 1755
rect 16950 1670 16970 1755
rect 16940 1665 16980 1670
rect 16940 1635 16945 1665
rect 16975 1635 16980 1665
rect 16940 1630 16980 1635
rect 16485 1620 16525 1625
rect 16485 1590 16490 1620
rect 16520 1590 16525 1620
rect 16485 1585 16525 1590
rect 16365 1520 16405 1525
rect 16365 1490 16370 1520
rect 16400 1490 16405 1520
rect 16365 1480 16405 1490
rect 16365 1450 16370 1480
rect 16400 1450 16405 1480
rect 16365 1440 16405 1450
rect 16365 1410 16370 1440
rect 16400 1410 16405 1440
rect 16365 1405 16405 1410
rect 16485 1520 16525 1525
rect 16485 1490 16490 1520
rect 16520 1490 16525 1520
rect 16485 1480 16525 1490
rect 16485 1450 16490 1480
rect 16520 1450 16525 1480
rect 16485 1440 16525 1450
rect 16485 1410 16490 1440
rect 16520 1410 16525 1440
rect 16485 1405 16525 1410
rect 16605 1520 16645 1525
rect 16605 1490 16610 1520
rect 16640 1490 16645 1520
rect 16605 1480 16645 1490
rect 16605 1450 16610 1480
rect 16640 1450 16645 1480
rect 16605 1440 16645 1450
rect 16605 1410 16610 1440
rect 16640 1410 16645 1440
rect 16605 1405 16645 1410
rect 16885 1520 16925 1525
rect 16885 1490 16890 1520
rect 16920 1490 16925 1520
rect 16885 1480 16925 1490
rect 16885 1450 16890 1480
rect 16920 1450 16925 1480
rect 16885 1440 16925 1450
rect 16950 1445 16970 1630
rect 17050 1620 17090 1625
rect 17050 1590 17055 1620
rect 17085 1590 17090 1620
rect 17050 1585 17090 1590
rect 16995 1520 17035 1525
rect 16995 1490 17000 1520
rect 17030 1490 17035 1520
rect 16995 1480 17035 1490
rect 16995 1450 17000 1480
rect 17030 1450 17035 1480
rect 16885 1410 16890 1440
rect 16920 1410 16925 1440
rect 16885 1405 16925 1410
rect 16945 1435 16975 1445
rect 16945 1415 16950 1435
rect 16970 1415 16975 1435
rect 16945 1405 16975 1415
rect 16995 1440 17035 1450
rect 17060 1445 17080 1585
rect 17105 1520 17145 1525
rect 17105 1490 17110 1520
rect 17140 1490 17145 1520
rect 17105 1480 17145 1490
rect 17105 1450 17110 1480
rect 17140 1450 17145 1480
rect 16995 1410 17000 1440
rect 17030 1410 17035 1440
rect 16995 1405 17035 1410
rect 17055 1435 17085 1445
rect 17055 1415 17060 1435
rect 17080 1415 17085 1435
rect 17055 1405 17085 1415
rect 17105 1440 17145 1450
rect 17105 1410 17110 1440
rect 17140 1410 17145 1440
rect 17105 1405 17145 1410
rect 17215 1520 17255 1525
rect 17215 1490 17220 1520
rect 17250 1490 17255 1520
rect 17215 1480 17255 1490
rect 17215 1450 17220 1480
rect 17250 1450 17255 1480
rect 17215 1440 17255 1450
rect 17215 1410 17220 1440
rect 17250 1410 17255 1440
rect 17215 1405 17255 1410
rect 17495 1520 17535 1525
rect 17495 1490 17500 1520
rect 17530 1490 17535 1520
rect 17495 1480 17535 1490
rect 17495 1450 17500 1480
rect 17530 1450 17535 1480
rect 17495 1440 17535 1450
rect 17495 1410 17500 1440
rect 17530 1410 17535 1440
rect 17495 1405 17535 1410
rect 17560 1520 17600 1525
rect 17560 1490 17565 1520
rect 17595 1490 17600 1520
rect 17560 1480 17600 1490
rect 17560 1450 17565 1480
rect 17595 1450 17600 1480
rect 17560 1440 17600 1450
rect 17560 1410 17565 1440
rect 17595 1410 17600 1440
rect 17560 1405 17600 1410
rect 17620 1435 17650 1755
rect 17620 1415 17625 1435
rect 17645 1415 17650 1435
rect 17620 1405 17650 1415
rect 17670 1520 17710 1525
rect 17670 1490 17675 1520
rect 17705 1490 17710 1520
rect 17670 1480 17710 1490
rect 17670 1450 17675 1480
rect 17705 1450 17710 1480
rect 17670 1440 17710 1450
rect 17670 1410 17675 1440
rect 17705 1410 17710 1440
rect 17670 1405 17710 1410
rect 17730 1435 17760 1755
rect 17780 1620 17820 1625
rect 17780 1590 17785 1620
rect 17815 1590 17820 1620
rect 17780 1585 17820 1590
rect 17730 1415 17735 1435
rect 17755 1415 17760 1435
rect 17730 1405 17760 1415
rect 17780 1520 17820 1525
rect 17780 1490 17785 1520
rect 17815 1490 17820 1520
rect 17780 1480 17820 1490
rect 17780 1450 17785 1480
rect 17815 1450 17820 1480
rect 17780 1440 17820 1450
rect 17780 1410 17785 1440
rect 17815 1410 17820 1440
rect 17780 1405 17820 1410
rect 17840 1435 17870 1755
rect 17840 1415 17845 1435
rect 17865 1415 17870 1435
rect 17840 1405 17870 1415
rect 17890 1520 17930 1525
rect 17890 1490 17895 1520
rect 17925 1490 17930 1520
rect 17890 1480 17930 1490
rect 17890 1450 17895 1480
rect 17925 1450 17930 1480
rect 17890 1440 17930 1450
rect 17890 1410 17895 1440
rect 17925 1410 17930 1440
rect 17890 1405 17930 1410
rect 17950 1435 17980 1755
rect 18630 1670 18650 1755
rect 18620 1665 18660 1670
rect 18620 1635 18625 1665
rect 18655 1635 18660 1665
rect 18620 1630 18660 1635
rect 18200 1620 18240 1625
rect 18200 1590 18205 1620
rect 18235 1590 18240 1620
rect 18200 1585 18240 1590
rect 18510 1620 18550 1625
rect 18510 1590 18515 1620
rect 18545 1590 18550 1620
rect 18510 1585 18550 1590
rect 17950 1415 17955 1435
rect 17975 1415 17980 1435
rect 17950 1405 17980 1415
rect 18000 1520 18040 1525
rect 18000 1490 18005 1520
rect 18035 1490 18040 1520
rect 18000 1480 18040 1490
rect 18000 1450 18005 1480
rect 18035 1450 18040 1480
rect 18000 1440 18040 1450
rect 18000 1410 18005 1440
rect 18035 1410 18040 1440
rect 18000 1405 18040 1410
rect 18065 1520 18105 1525
rect 18065 1490 18070 1520
rect 18100 1490 18105 1520
rect 18065 1480 18105 1490
rect 18065 1450 18070 1480
rect 18100 1450 18105 1480
rect 18065 1440 18105 1450
rect 18065 1410 18070 1440
rect 18100 1410 18105 1440
rect 18065 1405 18105 1410
rect 16430 1270 16470 1275
rect 16430 1240 16435 1270
rect 16465 1240 16470 1270
rect 16430 1235 16470 1240
rect 16540 1270 16580 1275
rect 16540 1240 16545 1270
rect 16575 1240 16580 1270
rect 16540 1235 16580 1240
rect 16940 1270 16980 1275
rect 16940 1240 16945 1270
rect 16975 1240 16980 1270
rect 16940 1235 16980 1240
rect 17050 1270 17090 1275
rect 17050 1240 17055 1270
rect 17085 1240 17090 1270
rect 17050 1235 17090 1240
rect 17160 1270 17200 1275
rect 17160 1240 17165 1270
rect 17195 1240 17200 1270
rect 17160 1235 17200 1240
rect 17615 1270 17655 1275
rect 17615 1240 17620 1270
rect 17650 1240 17655 1270
rect 17615 1235 17655 1240
rect 17725 1270 17765 1275
rect 17725 1240 17730 1270
rect 17760 1240 17765 1270
rect 17725 1235 17765 1240
rect 17835 1270 17875 1275
rect 17835 1240 17840 1270
rect 17870 1240 17875 1270
rect 17835 1235 17875 1240
rect 17945 1270 17985 1275
rect 17945 1240 17950 1270
rect 17980 1240 17985 1270
rect 17945 1235 17985 1240
rect 16440 1175 16460 1235
rect 16550 1175 16570 1235
rect 18210 1220 18230 1585
rect 18345 1520 18385 1525
rect 18345 1490 18350 1520
rect 18380 1490 18385 1520
rect 18345 1480 18385 1490
rect 18345 1450 18350 1480
rect 18380 1450 18385 1480
rect 18345 1440 18385 1450
rect 18345 1410 18350 1440
rect 18380 1410 18385 1440
rect 18345 1405 18385 1410
rect 18455 1520 18495 1525
rect 18455 1490 18460 1520
rect 18490 1490 18495 1520
rect 18455 1480 18495 1490
rect 18455 1450 18460 1480
rect 18490 1450 18495 1480
rect 18455 1440 18495 1450
rect 18520 1445 18540 1585
rect 18565 1520 18605 1525
rect 18565 1490 18570 1520
rect 18600 1490 18605 1520
rect 18565 1480 18605 1490
rect 18565 1450 18570 1480
rect 18600 1450 18605 1480
rect 18455 1410 18460 1440
rect 18490 1410 18495 1440
rect 18455 1405 18495 1410
rect 18515 1435 18545 1445
rect 18515 1415 18520 1435
rect 18540 1415 18545 1435
rect 18515 1405 18545 1415
rect 18565 1440 18605 1450
rect 18630 1445 18650 1630
rect 18675 1520 18715 1525
rect 18675 1490 18680 1520
rect 18710 1490 18715 1520
rect 18675 1480 18715 1490
rect 18675 1450 18680 1480
rect 18710 1450 18715 1480
rect 18565 1410 18570 1440
rect 18600 1410 18605 1440
rect 18565 1405 18605 1410
rect 18625 1435 18655 1445
rect 18625 1415 18630 1435
rect 18650 1415 18655 1435
rect 18625 1405 18655 1415
rect 18675 1440 18715 1450
rect 18675 1410 18680 1440
rect 18710 1410 18715 1440
rect 18675 1405 18715 1410
rect 18400 1270 18440 1275
rect 18400 1240 18405 1270
rect 18435 1240 18440 1270
rect 18400 1235 18440 1240
rect 18510 1270 18550 1275
rect 18510 1240 18515 1270
rect 18545 1240 18550 1270
rect 18510 1235 18550 1240
rect 18620 1270 18660 1275
rect 18620 1240 18625 1270
rect 18655 1240 18660 1270
rect 18620 1235 18660 1240
rect 18200 1215 18240 1220
rect 18200 1185 18205 1215
rect 18235 1185 18240 1215
rect 18200 1180 18240 1185
rect 18720 1215 18760 1220
rect 18720 1185 18725 1215
rect 18755 1185 18760 1215
rect 18720 1180 18760 1185
rect 16160 1170 16200 1175
rect 16160 1140 16165 1170
rect 16195 1140 16200 1170
rect 16160 1135 16200 1140
rect 16430 1170 16470 1175
rect 16430 1140 16435 1170
rect 16465 1140 16470 1170
rect 16430 1135 16470 1140
rect 16540 1170 16580 1175
rect 16540 1140 16545 1170
rect 16575 1140 16580 1170
rect 16540 1135 16580 1140
rect 16170 -1320 16190 1135
rect 16435 1055 16475 1060
rect 16435 1025 16440 1055
rect 16470 1025 16475 1055
rect 16435 1015 16475 1025
rect 16435 985 16440 1015
rect 16470 985 16475 1015
rect 16435 975 16475 985
rect 16435 945 16440 975
rect 16470 945 16475 975
rect 16435 940 16475 945
rect 16655 1055 16695 1060
rect 16655 1025 16660 1055
rect 16690 1025 16695 1055
rect 16655 1015 16695 1025
rect 16655 985 16660 1015
rect 16690 985 16695 1015
rect 16655 975 16695 985
rect 16655 945 16660 975
rect 16690 945 16695 975
rect 16655 940 16695 945
rect 16970 1055 17010 1060
rect 16970 1025 16975 1055
rect 17005 1025 17010 1055
rect 16970 1015 17010 1025
rect 16970 985 16975 1015
rect 17005 985 17010 1015
rect 16970 975 17010 985
rect 16970 945 16975 975
rect 17005 945 17010 975
rect 16970 940 17010 945
rect 17150 1055 17190 1060
rect 17150 1025 17155 1055
rect 17185 1025 17190 1055
rect 17150 1015 17190 1025
rect 17150 985 17155 1015
rect 17185 985 17190 1015
rect 17150 975 17190 985
rect 17150 945 17155 975
rect 17185 945 17190 975
rect 17150 940 17190 945
rect 17330 1055 17370 1060
rect 17330 1025 17335 1055
rect 17365 1025 17370 1055
rect 17330 1015 17370 1025
rect 17330 985 17335 1015
rect 17365 985 17370 1015
rect 17330 975 17370 985
rect 17330 945 17335 975
rect 17365 945 17370 975
rect 17330 940 17370 945
rect 17510 1055 17550 1060
rect 17510 1025 17515 1055
rect 17545 1025 17550 1055
rect 17510 1015 17550 1025
rect 17510 985 17515 1015
rect 17545 985 17550 1015
rect 17510 975 17550 985
rect 17510 945 17515 975
rect 17545 945 17550 975
rect 17510 940 17550 945
rect 17690 1055 17730 1060
rect 17690 1025 17695 1055
rect 17725 1025 17730 1055
rect 17690 1015 17730 1025
rect 17690 985 17695 1015
rect 17725 985 17730 1015
rect 17690 975 17730 985
rect 17690 945 17695 975
rect 17725 945 17730 975
rect 17690 940 17730 945
rect 17870 1055 17910 1060
rect 17870 1025 17875 1055
rect 17905 1025 17910 1055
rect 17870 1015 17910 1025
rect 17870 985 17875 1015
rect 17905 985 17910 1015
rect 17870 975 17910 985
rect 17870 945 17875 975
rect 17905 945 17910 975
rect 17870 940 17910 945
rect 18050 1055 18090 1060
rect 18050 1025 18055 1055
rect 18085 1025 18090 1055
rect 18050 1015 18090 1025
rect 18050 985 18055 1015
rect 18085 985 18090 1015
rect 18050 975 18090 985
rect 18050 945 18055 975
rect 18085 945 18090 975
rect 18050 940 18090 945
rect 18230 1055 18270 1060
rect 18230 1025 18235 1055
rect 18265 1025 18270 1055
rect 18230 1015 18270 1025
rect 18230 985 18235 1015
rect 18265 985 18270 1015
rect 18230 975 18270 985
rect 18230 945 18235 975
rect 18265 945 18270 975
rect 18230 940 18270 945
rect 18410 1055 18450 1060
rect 18410 1025 18415 1055
rect 18445 1025 18450 1055
rect 18410 1015 18450 1025
rect 18410 985 18415 1015
rect 18445 985 18450 1015
rect 18410 975 18450 985
rect 18410 945 18415 975
rect 18445 945 18450 975
rect 18410 940 18450 945
rect 18590 1055 18630 1060
rect 18590 1025 18595 1055
rect 18625 1025 18630 1055
rect 18590 1015 18630 1025
rect 18590 985 18595 1015
rect 18625 985 18630 1015
rect 18590 975 18630 985
rect 18590 945 18595 975
rect 18625 945 18630 975
rect 18590 940 18630 945
rect 16445 880 16465 940
rect 16665 880 16685 940
rect 16435 870 16475 880
rect 16435 850 16445 870
rect 16465 850 16475 870
rect 16435 840 16475 850
rect 16545 875 16585 880
rect 16545 845 16550 875
rect 16580 845 16585 875
rect 16545 840 16585 845
rect 16655 870 16695 880
rect 16655 850 16665 870
rect 16685 850 16695 870
rect 16655 840 16695 850
rect 16780 875 16820 880
rect 16780 845 16785 875
rect 16815 845 16820 875
rect 16780 840 16820 845
rect 16480 705 16520 710
rect 16480 675 16485 705
rect 16515 675 16520 705
rect 16480 670 16520 675
rect 16545 700 16585 710
rect 16545 680 16555 700
rect 16575 680 16585 700
rect 16545 670 16585 680
rect 16610 705 16650 710
rect 16610 675 16615 705
rect 16645 675 16650 705
rect 16610 670 16650 675
rect 16315 605 16355 610
rect 16315 575 16320 605
rect 16350 575 16355 605
rect 16260 550 16300 555
rect 16260 520 16265 550
rect 16295 520 16300 550
rect 16260 515 16300 520
rect 16205 505 16245 510
rect 16205 475 16210 505
rect 16240 475 16245 505
rect 16205 470 16245 475
rect 16215 -1220 16235 470
rect 16270 -145 16290 515
rect 16260 -150 16300 -145
rect 16260 -180 16265 -150
rect 16295 -180 16300 -150
rect 16260 -185 16300 -180
rect 16205 -1225 16245 -1220
rect 16205 -1255 16210 -1225
rect 16240 -1255 16245 -1225
rect 16205 -1260 16245 -1255
rect 16160 -1325 16200 -1320
rect 16160 -1355 16165 -1325
rect 16195 -1355 16200 -1325
rect 16160 -1360 16200 -1355
rect 16105 -1900 16145 -1895
rect 16105 -1930 16110 -1900
rect 16140 -1930 16145 -1900
rect 16105 -1935 16145 -1930
rect 16155 -1950 16195 -1945
rect 16155 -1980 16160 -1950
rect 16190 -1980 16195 -1950
rect 16155 -1985 16195 -1980
rect 16165 -3020 16185 -1985
rect 16270 -1995 16290 -185
rect 16315 -470 16355 575
rect 16555 510 16575 670
rect 16790 555 16810 840
rect 16840 705 16880 710
rect 16840 675 16845 705
rect 16875 675 16880 705
rect 16840 670 16880 675
rect 16780 550 16820 555
rect 16780 520 16785 550
rect 16815 520 16820 550
rect 16780 515 16820 520
rect 16545 505 16585 510
rect 16545 475 16550 505
rect 16580 475 16585 505
rect 16545 470 16585 475
rect 16420 270 16460 275
rect 16420 240 16425 270
rect 16455 240 16460 270
rect 16420 230 16460 240
rect 16420 200 16425 230
rect 16455 200 16460 230
rect 16420 190 16460 200
rect 16420 160 16425 190
rect 16455 160 16460 190
rect 16420 155 16460 160
rect 16540 270 16580 275
rect 16540 240 16545 270
rect 16575 240 16580 270
rect 16540 230 16580 240
rect 16540 200 16545 230
rect 16575 200 16580 230
rect 16540 190 16580 200
rect 16540 160 16545 190
rect 16575 160 16580 190
rect 16540 155 16580 160
rect 16660 270 16700 275
rect 16660 240 16665 270
rect 16695 240 16700 270
rect 16660 230 16700 240
rect 16660 200 16665 230
rect 16695 200 16700 230
rect 16660 190 16700 200
rect 16660 160 16665 190
rect 16695 160 16700 190
rect 16660 155 16700 160
rect 16780 270 16820 275
rect 16780 240 16785 270
rect 16815 240 16820 270
rect 16780 230 16820 240
rect 16780 200 16785 230
rect 16815 200 16820 230
rect 16780 190 16820 200
rect 16780 160 16785 190
rect 16815 160 16820 190
rect 16780 155 16820 160
rect 16430 140 16450 155
rect 16550 140 16570 155
rect 16670 140 16690 155
rect 16790 140 16810 155
rect 16850 140 16870 670
rect 17060 600 17100 610
rect 17060 580 17070 600
rect 17090 580 17100 600
rect 17060 570 17100 580
rect 17240 600 17280 610
rect 17240 580 17250 600
rect 17270 580 17280 600
rect 17240 570 17280 580
rect 17420 600 17460 610
rect 17420 580 17430 600
rect 17450 580 17460 600
rect 17420 570 17460 580
rect 17600 605 17640 610
rect 17600 575 17605 605
rect 17635 575 17640 605
rect 17600 570 17640 575
rect 17690 600 17730 610
rect 17690 580 17700 600
rect 17720 580 17730 600
rect 17690 570 17730 580
rect 17780 600 17820 610
rect 17780 580 17790 600
rect 17810 580 17820 600
rect 17780 570 17820 580
rect 17960 605 18000 610
rect 17960 575 17965 605
rect 17995 575 18000 605
rect 17960 570 18000 575
rect 18140 600 18180 610
rect 18140 580 18150 600
rect 18170 580 18180 600
rect 18140 570 18180 580
rect 18320 600 18360 610
rect 18320 580 18330 600
rect 18350 580 18360 600
rect 18320 570 18360 580
rect 18410 600 18450 610
rect 18410 580 18420 600
rect 18440 580 18450 600
rect 18410 570 18450 580
rect 18500 600 18540 610
rect 18500 580 18510 600
rect 18530 580 18540 600
rect 18500 570 18540 580
rect 17070 465 17090 570
rect 17250 510 17270 570
rect 17430 555 17450 570
rect 17420 550 17460 555
rect 17420 520 17425 550
rect 17455 520 17460 550
rect 17420 515 17460 520
rect 17240 505 17280 510
rect 17240 475 17245 505
rect 17275 475 17280 505
rect 17240 470 17280 475
rect 17060 460 17100 465
rect 17060 430 17065 460
rect 17095 430 17100 460
rect 17060 425 17100 430
rect 16900 270 16940 275
rect 16900 240 16905 270
rect 16935 240 16940 270
rect 16900 230 16940 240
rect 16900 200 16905 230
rect 16935 200 16940 230
rect 16900 190 16940 200
rect 16900 160 16905 190
rect 16935 160 16940 190
rect 16900 155 16940 160
rect 17020 270 17060 275
rect 17020 240 17025 270
rect 17055 240 17060 270
rect 17020 230 17060 240
rect 17020 200 17025 230
rect 17055 200 17060 230
rect 17020 190 17060 200
rect 17020 160 17025 190
rect 17055 160 17060 190
rect 17020 155 17060 160
rect 17140 270 17180 275
rect 17140 240 17145 270
rect 17175 240 17180 270
rect 17140 230 17180 240
rect 17140 200 17145 230
rect 17175 200 17180 230
rect 17140 190 17180 200
rect 17140 160 17145 190
rect 17175 160 17180 190
rect 17140 155 17180 160
rect 17260 270 17300 275
rect 17260 240 17265 270
rect 17295 240 17300 270
rect 17260 230 17300 240
rect 17260 200 17265 230
rect 17295 200 17300 230
rect 17260 190 17300 200
rect 17260 160 17265 190
rect 17295 160 17300 190
rect 17260 155 17300 160
rect 17380 270 17420 275
rect 17380 240 17385 270
rect 17415 240 17420 270
rect 17380 230 17420 240
rect 17380 200 17385 230
rect 17415 200 17420 230
rect 17380 190 17420 200
rect 17380 160 17385 190
rect 17415 160 17420 190
rect 17380 155 17420 160
rect 17500 270 17540 275
rect 17500 240 17505 270
rect 17535 240 17540 270
rect 17500 230 17540 240
rect 17500 200 17505 230
rect 17535 200 17540 230
rect 17500 190 17540 200
rect 17500 160 17505 190
rect 17535 160 17540 190
rect 17500 155 17540 160
rect 17620 270 17660 275
rect 17620 240 17625 270
rect 17655 240 17660 270
rect 17620 230 17660 240
rect 17620 200 17625 230
rect 17655 200 17660 230
rect 17620 190 17660 200
rect 17620 160 17625 190
rect 17655 160 17660 190
rect 17620 155 17660 160
rect 16910 140 16930 155
rect 17030 140 17050 155
rect 17150 140 17170 155
rect 17270 140 17290 155
rect 17390 140 17410 155
rect 17510 140 17530 155
rect 17630 140 17650 155
rect 17700 140 17720 570
rect 17790 465 17810 570
rect 18150 555 18170 570
rect 18140 550 18180 555
rect 18140 520 18145 550
rect 18175 520 18180 550
rect 18140 515 18180 520
rect 18330 510 18350 570
rect 18420 565 18440 570
rect 18320 505 18360 510
rect 18320 475 18325 505
rect 18355 475 18360 505
rect 18320 470 18360 475
rect 18510 465 18530 570
rect 17780 460 17820 465
rect 17780 430 17785 460
rect 17815 430 17820 460
rect 17780 425 17820 430
rect 18500 460 18540 465
rect 18500 430 18505 460
rect 18535 430 18540 460
rect 18500 425 18540 430
rect 18730 415 18750 1180
rect 18905 1055 18945 1060
rect 18905 1025 18910 1055
rect 18940 1025 18945 1055
rect 18905 1015 18945 1025
rect 18905 985 18910 1015
rect 18940 985 18945 1015
rect 18905 975 18945 985
rect 18905 945 18910 975
rect 18940 945 18945 975
rect 18905 940 18945 945
rect 19015 1055 19055 1060
rect 19015 1025 19020 1055
rect 19050 1025 19055 1055
rect 19015 1015 19055 1025
rect 19015 985 19020 1015
rect 19050 985 19055 1015
rect 19015 975 19055 985
rect 19015 945 19020 975
rect 19050 945 19055 975
rect 19015 940 19055 945
rect 19075 1055 19115 1060
rect 19075 1025 19080 1055
rect 19110 1025 19115 1055
rect 19075 1015 19115 1025
rect 19075 985 19080 1015
rect 19110 985 19115 1015
rect 19075 975 19115 985
rect 19075 945 19080 975
rect 19110 945 19115 975
rect 19075 940 19115 945
rect 19270 710 19290 1755
rect 19325 1170 19365 1175
rect 19325 1140 19330 1170
rect 19360 1140 19365 1170
rect 19325 1135 19365 1140
rect 18950 705 18990 710
rect 18950 675 18955 705
rect 18985 675 18990 705
rect 18950 670 18990 675
rect 19260 705 19300 710
rect 19260 675 19265 705
rect 19295 675 19300 705
rect 19260 670 19300 675
rect 19000 625 19005 655
rect 19035 625 19040 655
rect 19020 415 19040 625
rect 18000 410 18040 415
rect 18000 380 18005 410
rect 18035 380 18040 410
rect 18000 375 18040 380
rect 18720 410 18760 415
rect 18720 380 18725 410
rect 18755 380 18760 410
rect 18720 375 18760 380
rect 19010 410 19050 415
rect 19010 380 19015 410
rect 19045 380 19050 410
rect 19010 375 19050 380
rect 17940 270 17980 275
rect 17940 240 17945 270
rect 17975 240 17980 270
rect 17940 230 17980 240
rect 17940 200 17945 230
rect 17975 200 17980 230
rect 17940 190 17980 200
rect 17940 160 17945 190
rect 17975 160 17980 190
rect 17940 155 17980 160
rect 17950 140 17970 155
rect 18010 140 18030 375
rect 18060 270 18100 275
rect 18060 240 18065 270
rect 18095 240 18100 270
rect 18060 230 18100 240
rect 18060 200 18065 230
rect 18095 200 18100 230
rect 18060 190 18100 200
rect 18060 160 18065 190
rect 18095 160 18100 190
rect 18060 155 18100 160
rect 18180 270 18220 275
rect 18180 240 18185 270
rect 18215 240 18220 270
rect 18180 230 18220 240
rect 18180 200 18185 230
rect 18215 200 18220 230
rect 18180 190 18220 200
rect 18180 160 18185 190
rect 18215 160 18220 190
rect 18180 155 18220 160
rect 18300 270 18340 275
rect 18300 240 18305 270
rect 18335 240 18340 270
rect 18300 230 18340 240
rect 18300 200 18305 230
rect 18335 200 18340 230
rect 18300 190 18340 200
rect 18300 160 18305 190
rect 18335 160 18340 190
rect 18300 155 18340 160
rect 18420 270 18460 275
rect 18420 240 18425 270
rect 18455 240 18460 270
rect 18420 230 18460 240
rect 18420 200 18425 230
rect 18455 200 18460 230
rect 18420 190 18460 200
rect 18420 160 18425 190
rect 18455 160 18460 190
rect 18420 155 18460 160
rect 18540 270 18580 275
rect 18540 240 18545 270
rect 18575 240 18580 270
rect 18540 230 18580 240
rect 18540 200 18545 230
rect 18575 200 18580 230
rect 18540 190 18580 200
rect 18540 160 18545 190
rect 18575 160 18580 190
rect 18540 155 18580 160
rect 18660 270 18700 275
rect 18660 240 18665 270
rect 18695 240 18700 270
rect 18660 230 18700 240
rect 18660 200 18665 230
rect 18695 200 18700 230
rect 18660 190 18700 200
rect 18660 160 18665 190
rect 18695 160 18700 190
rect 18660 155 18700 160
rect 18780 270 18820 275
rect 18780 240 18785 270
rect 18815 240 18820 270
rect 18780 230 18820 240
rect 18780 200 18785 230
rect 18815 200 18820 230
rect 18780 190 18820 200
rect 18780 160 18785 190
rect 18815 160 18820 190
rect 18780 155 18820 160
rect 18900 270 18940 275
rect 18900 240 18905 270
rect 18935 240 18940 270
rect 18900 230 18940 240
rect 18900 200 18905 230
rect 18935 200 18940 230
rect 18900 190 18940 200
rect 18900 160 18905 190
rect 18935 160 18940 190
rect 18900 155 18940 160
rect 19020 270 19060 275
rect 19020 240 19025 270
rect 19055 240 19060 270
rect 19020 230 19060 240
rect 19020 200 19025 230
rect 19055 200 19060 230
rect 19020 190 19060 200
rect 19020 160 19025 190
rect 19055 160 19060 190
rect 19020 155 19060 160
rect 19140 270 19180 275
rect 19140 240 19145 270
rect 19175 240 19180 270
rect 19140 230 19180 240
rect 19140 200 19145 230
rect 19175 200 19180 230
rect 19140 190 19180 200
rect 19140 160 19145 190
rect 19175 160 19180 190
rect 19140 155 19180 160
rect 18070 140 18090 155
rect 18190 140 18210 155
rect 18310 140 18330 155
rect 18430 140 18450 155
rect 18550 140 18570 155
rect 18670 140 18690 155
rect 18790 140 18810 155
rect 18910 140 18930 155
rect 19030 140 19050 155
rect 19150 140 19170 155
rect 16425 130 16455 140
rect 16425 110 16430 130
rect 16450 110 16455 130
rect 16425 95 16455 110
rect 16480 135 16520 140
rect 16480 105 16485 135
rect 16515 105 16520 135
rect 16480 100 16520 105
rect 16545 130 16575 140
rect 16545 110 16550 130
rect 16570 110 16575 130
rect 16545 100 16575 110
rect 16665 130 16695 140
rect 16665 110 16670 130
rect 16690 110 16695 130
rect 16665 100 16695 110
rect 16785 130 16815 140
rect 16785 110 16790 130
rect 16810 110 16815 130
rect 16785 100 16815 110
rect 16840 135 16880 140
rect 16840 105 16845 135
rect 16875 105 16880 135
rect 16840 100 16880 105
rect 16905 130 16935 140
rect 16905 110 16910 130
rect 16930 110 16935 130
rect 16905 100 16935 110
rect 17025 130 17055 140
rect 17025 110 17030 130
rect 17050 110 17055 130
rect 17025 100 17055 110
rect 17145 130 17175 140
rect 17145 110 17150 130
rect 17170 110 17175 130
rect 17145 100 17175 110
rect 17200 135 17240 140
rect 17200 105 17205 135
rect 17235 105 17240 135
rect 17200 100 17240 105
rect 17265 130 17295 140
rect 17265 110 17270 130
rect 17290 110 17295 130
rect 17265 100 17295 110
rect 17385 130 17415 140
rect 17385 110 17390 130
rect 17410 110 17415 130
rect 17385 100 17415 110
rect 17505 130 17535 140
rect 17505 110 17510 130
rect 17530 110 17535 130
rect 17505 100 17535 110
rect 17560 135 17600 140
rect 17560 105 17565 135
rect 17595 105 17600 135
rect 17560 100 17600 105
rect 17625 130 17655 140
rect 17625 110 17630 130
rect 17650 110 17655 130
rect 17625 95 17655 110
rect 17690 135 17730 140
rect 17690 105 17695 135
rect 17725 105 17730 135
rect 17690 100 17730 105
rect 17870 135 17910 140
rect 17870 105 17875 135
rect 17905 105 17910 135
rect 17870 100 17910 105
rect 17945 130 17975 140
rect 17945 110 17950 130
rect 17970 110 17975 130
rect 16510 -40 16550 -30
rect 16510 -60 16520 -40
rect 16540 -60 16550 -40
rect 16510 -70 16550 -60
rect 16600 -35 16640 -30
rect 16600 -65 16605 -35
rect 16635 -65 16640 -35
rect 16600 -70 16640 -65
rect 16720 -40 16760 -30
rect 16720 -60 16730 -40
rect 16750 -60 16760 -40
rect 16720 -70 16760 -60
rect 16840 -40 16880 -30
rect 16840 -60 16850 -40
rect 16870 -60 16880 -40
rect 16840 -70 16880 -60
rect 16960 -35 17000 -30
rect 16960 -65 16965 -35
rect 16995 -65 17000 -35
rect 16960 -70 17000 -65
rect 17080 -40 17120 -30
rect 17080 -60 17090 -40
rect 17110 -60 17120 -40
rect 17080 -70 17120 -60
rect 17200 -40 17240 -30
rect 17200 -60 17210 -40
rect 17230 -60 17240 -40
rect 17200 -70 17240 -60
rect 17320 -35 17360 -30
rect 17320 -65 17325 -35
rect 17355 -65 17360 -35
rect 17320 -70 17360 -65
rect 17440 -40 17480 -30
rect 17440 -60 17450 -40
rect 17470 -60 17480 -40
rect 17440 -70 17480 -60
rect 17535 -40 17565 -30
rect 17535 -60 17540 -40
rect 17560 -60 17565 -40
rect 17535 -70 17565 -60
rect 16520 -90 16540 -70
rect 16730 -90 16750 -70
rect 16850 -90 16870 -70
rect 16510 -95 16550 -90
rect 16510 -125 16515 -95
rect 16545 -125 16550 -95
rect 16510 -130 16550 -125
rect 16720 -95 16760 -90
rect 16720 -125 16725 -95
rect 16755 -125 16760 -95
rect 16720 -130 16760 -125
rect 16840 -95 16880 -90
rect 16840 -125 16845 -95
rect 16875 -125 16880 -95
rect 16840 -130 16880 -125
rect 16970 -145 16990 -70
rect 17090 -90 17110 -70
rect 17210 -90 17230 -70
rect 17450 -90 17470 -70
rect 17540 -90 17560 -70
rect 17080 -95 17120 -90
rect 17080 -125 17085 -95
rect 17115 -125 17120 -95
rect 17080 -130 17120 -125
rect 17200 -95 17240 -90
rect 17200 -125 17205 -95
rect 17235 -125 17240 -95
rect 17200 -130 17240 -125
rect 17440 -95 17480 -90
rect 17440 -125 17445 -95
rect 17475 -125 17480 -95
rect 17440 -130 17480 -125
rect 17530 -95 17570 -90
rect 17530 -125 17535 -95
rect 17565 -125 17570 -95
rect 17530 -130 17570 -125
rect 17090 -145 17110 -130
rect 16960 -155 16990 -145
rect 16960 -175 16965 -155
rect 16985 -175 16990 -155
rect 16960 -185 16990 -175
rect 17007 -150 17037 -145
rect 17007 -185 17037 -180
rect 17090 -155 17120 -145
rect 17090 -175 17095 -155
rect 17115 -175 17120 -155
rect 17090 -185 17120 -175
rect 16315 -500 16320 -470
rect 16350 -500 16355 -470
rect 16315 -505 16355 -500
rect 17025 -215 17055 -205
rect 17025 -235 17030 -215
rect 17050 -235 17055 -215
rect 17025 -265 17055 -235
rect 17025 -285 17030 -265
rect 17050 -285 17055 -265
rect 17025 -315 17055 -285
rect 17025 -335 17030 -315
rect 17050 -335 17055 -315
rect 17560 -210 17600 -205
rect 17560 -240 17565 -210
rect 17595 -240 17600 -210
rect 17560 -250 17600 -240
rect 17560 -280 17565 -250
rect 17595 -280 17600 -250
rect 17560 -290 17600 -280
rect 17560 -320 17565 -290
rect 17595 -320 17600 -290
rect 17560 -325 17600 -320
rect 17025 -365 17055 -335
rect 17025 -385 17030 -365
rect 17050 -385 17055 -365
rect 17025 -415 17055 -385
rect 17025 -435 17030 -415
rect 17050 -435 17055 -415
rect 17025 -545 17055 -435
rect 17075 -470 17105 -465
rect 17075 -505 17105 -500
rect 16530 -550 16570 -545
rect 16530 -580 16535 -550
rect 16565 -580 16570 -550
rect 16530 -585 16570 -580
rect 17020 -550 17060 -545
rect 17020 -580 17025 -550
rect 17055 -580 17060 -550
rect 17020 -585 17060 -580
rect 16535 -750 16565 -585
rect 16620 -605 16660 -600
rect 16620 -635 16625 -605
rect 16655 -635 16660 -605
rect 16620 -645 16660 -635
rect 16620 -675 16625 -645
rect 16655 -675 16660 -645
rect 16620 -685 16660 -675
rect 16620 -715 16625 -685
rect 16655 -715 16660 -685
rect 16620 -720 16660 -715
rect 16740 -605 16780 -600
rect 16740 -635 16745 -605
rect 16775 -635 16780 -605
rect 16740 -645 16780 -635
rect 16740 -675 16745 -645
rect 16775 -675 16780 -645
rect 16740 -685 16780 -675
rect 16740 -715 16745 -685
rect 16775 -715 16780 -685
rect 16740 -720 16780 -715
rect 16860 -605 16900 -600
rect 16860 -635 16865 -605
rect 16895 -635 16900 -605
rect 16860 -645 16900 -635
rect 16860 -675 16865 -645
rect 16895 -675 16900 -645
rect 16860 -685 16900 -675
rect 16860 -715 16865 -685
rect 16895 -715 16900 -685
rect 16860 -720 16900 -715
rect 16980 -605 17020 -600
rect 16980 -635 16985 -605
rect 17015 -635 17020 -605
rect 16980 -645 17020 -635
rect 16980 -675 16985 -645
rect 17015 -675 17020 -645
rect 16980 -685 17020 -675
rect 16980 -715 16985 -685
rect 17015 -715 17020 -685
rect 16980 -720 17020 -715
rect 17300 -605 17340 -600
rect 17300 -635 17305 -605
rect 17335 -635 17340 -605
rect 17300 -645 17340 -635
rect 17300 -675 17305 -645
rect 17335 -675 17340 -645
rect 17300 -685 17340 -675
rect 17300 -715 17305 -685
rect 17335 -715 17340 -685
rect 17300 -720 17340 -715
rect 17420 -605 17460 -600
rect 17420 -635 17425 -605
rect 17455 -635 17460 -605
rect 17420 -645 17460 -635
rect 17420 -675 17425 -645
rect 17455 -675 17460 -645
rect 17420 -685 17460 -675
rect 17420 -715 17425 -685
rect 17455 -715 17460 -685
rect 17420 -720 17460 -715
rect 17540 -605 17580 -600
rect 17540 -635 17545 -605
rect 17575 -635 17580 -605
rect 17540 -645 17580 -635
rect 17540 -675 17545 -645
rect 17575 -675 17580 -645
rect 17540 -685 17580 -675
rect 17540 -715 17545 -685
rect 17575 -715 17580 -685
rect 17700 -695 17720 100
rect 17740 -210 17860 -205
rect 17740 -240 17745 -210
rect 17775 -240 17785 -210
rect 17815 -240 17825 -210
rect 17855 -240 17860 -210
rect 17740 -250 17860 -240
rect 17740 -280 17745 -250
rect 17775 -280 17785 -250
rect 17815 -280 17825 -250
rect 17855 -280 17860 -250
rect 17740 -290 17860 -280
rect 17740 -320 17745 -290
rect 17775 -320 17785 -290
rect 17815 -320 17825 -290
rect 17855 -320 17860 -290
rect 17540 -720 17580 -715
rect 17695 -705 17725 -695
rect 17695 -725 17700 -705
rect 17720 -725 17725 -705
rect 17695 -735 17725 -725
rect 16535 -770 16540 -750
rect 16560 -770 16565 -750
rect 16535 -800 16565 -770
rect 16535 -820 16540 -800
rect 16560 -820 16565 -800
rect 16535 -850 16565 -820
rect 16535 -870 16540 -850
rect 16560 -870 16565 -850
rect 16535 -900 16565 -870
rect 16535 -920 16540 -900
rect 16560 -920 16565 -900
rect 16535 -950 16565 -920
rect 16535 -970 16540 -950
rect 16560 -970 16565 -950
rect 16535 -980 16565 -970
rect 17110 -1005 17150 -1000
rect 17110 -1035 17115 -1005
rect 17145 -1035 17150 -1005
rect 17110 -1045 17150 -1035
rect 17110 -1075 17115 -1045
rect 17145 -1075 17150 -1045
rect 17110 -1085 17150 -1075
rect 17110 -1115 17115 -1085
rect 17145 -1115 17150 -1085
rect 17110 -1120 17150 -1115
rect 17740 -1005 17860 -320
rect 17880 -695 17900 100
rect 17945 95 17975 110
rect 18000 135 18040 140
rect 18000 105 18005 135
rect 18035 105 18040 135
rect 18000 100 18040 105
rect 18065 130 18095 140
rect 18065 110 18070 130
rect 18090 110 18095 130
rect 18065 100 18095 110
rect 18185 130 18215 140
rect 18185 110 18190 130
rect 18210 110 18215 130
rect 18185 100 18215 110
rect 18305 130 18335 140
rect 18305 110 18310 130
rect 18330 110 18335 130
rect 18305 100 18335 110
rect 18360 135 18400 140
rect 18360 105 18365 135
rect 18395 105 18400 135
rect 18360 100 18400 105
rect 18425 130 18455 140
rect 18425 110 18430 130
rect 18450 110 18455 130
rect 18425 100 18455 110
rect 18545 130 18575 140
rect 18545 110 18550 130
rect 18570 110 18575 130
rect 18545 100 18575 110
rect 18665 130 18695 140
rect 18665 110 18670 130
rect 18690 110 18695 130
rect 18665 100 18695 110
rect 18720 135 18760 140
rect 18720 105 18725 135
rect 18755 105 18760 135
rect 18720 100 18760 105
rect 18785 130 18815 140
rect 18785 110 18790 130
rect 18810 110 18815 130
rect 18785 100 18815 110
rect 18905 130 18935 140
rect 18905 110 18910 130
rect 18930 110 18935 130
rect 18905 100 18935 110
rect 19025 130 19055 140
rect 19025 110 19030 130
rect 19050 110 19055 130
rect 19025 100 19055 110
rect 19080 135 19120 140
rect 19080 105 19085 135
rect 19115 105 19120 135
rect 19080 100 19120 105
rect 19145 130 19175 140
rect 19145 110 19150 130
rect 19170 110 19175 130
rect 19145 95 19175 110
rect 18035 -40 18065 -30
rect 18035 -60 18040 -40
rect 18060 -60 18065 -40
rect 18035 -70 18065 -60
rect 18120 -40 18160 -30
rect 18120 -60 18130 -40
rect 18150 -60 18160 -40
rect 18120 -70 18160 -60
rect 18240 -35 18280 -30
rect 18240 -65 18245 -35
rect 18275 -65 18280 -35
rect 18240 -70 18280 -65
rect 18360 -40 18400 -30
rect 18360 -60 18370 -40
rect 18390 -60 18400 -40
rect 18360 -70 18400 -60
rect 18480 -40 18520 -30
rect 18480 -60 18490 -40
rect 18510 -60 18520 -40
rect 18480 -70 18520 -60
rect 18600 -35 18640 -30
rect 18600 -65 18605 -35
rect 18635 -65 18640 -35
rect 18600 -70 18640 -65
rect 18720 -40 18760 -30
rect 18720 -60 18730 -40
rect 18750 -60 18760 -40
rect 18720 -70 18760 -60
rect 18840 -40 18880 -30
rect 18840 -60 18850 -40
rect 18870 -60 18880 -40
rect 18840 -70 18880 -60
rect 18960 -35 19000 -30
rect 18960 -65 18965 -35
rect 18995 -65 19000 -35
rect 18960 -70 19000 -65
rect 19050 -40 19090 -30
rect 19050 -60 19060 -40
rect 19080 -60 19090 -40
rect 19050 -70 19090 -60
rect 18040 -90 18060 -70
rect 18130 -90 18150 -70
rect 18370 -90 18390 -70
rect 18490 -90 18510 -70
rect 18030 -95 18070 -90
rect 18030 -125 18035 -95
rect 18065 -125 18070 -95
rect 18030 -130 18070 -125
rect 18120 -95 18160 -90
rect 18120 -125 18125 -95
rect 18155 -125 18160 -95
rect 18120 -130 18160 -125
rect 18360 -95 18400 -90
rect 18360 -125 18365 -95
rect 18395 -125 18400 -95
rect 18360 -130 18400 -125
rect 18480 -95 18520 -90
rect 18480 -125 18485 -95
rect 18515 -125 18520 -95
rect 18480 -130 18520 -125
rect 18490 -145 18510 -130
rect 18610 -145 18630 -70
rect 18730 -90 18750 -70
rect 18850 -90 18870 -70
rect 19060 -90 19080 -70
rect 18720 -95 18760 -90
rect 18720 -125 18725 -95
rect 18755 -125 18760 -95
rect 18720 -130 18760 -125
rect 18840 -95 18880 -90
rect 18840 -125 18845 -95
rect 18875 -125 18880 -95
rect 18840 -130 18880 -125
rect 19050 -95 19090 -90
rect 19050 -125 19055 -95
rect 19085 -125 19090 -95
rect 19050 -130 19090 -125
rect 18480 -155 18510 -145
rect 18480 -175 18485 -155
rect 18505 -175 18510 -155
rect 18480 -185 18510 -175
rect 18563 -150 18593 -145
rect 18563 -185 18593 -180
rect 18610 -155 18640 -145
rect 18610 -175 18615 -155
rect 18635 -175 18640 -155
rect 18610 -185 18640 -175
rect 18000 -210 18040 -205
rect 18000 -240 18005 -210
rect 18035 -240 18040 -210
rect 18000 -250 18040 -240
rect 18000 -280 18005 -250
rect 18035 -280 18040 -250
rect 18000 -290 18040 -280
rect 18000 -320 18005 -290
rect 18035 -320 18040 -290
rect 18000 -325 18040 -320
rect 19335 -465 19355 1135
rect 19415 465 19435 1755
rect 19460 605 19500 610
rect 19460 575 19465 605
rect 19495 575 19500 605
rect 19405 460 19445 465
rect 19405 430 19410 460
rect 19440 430 19445 460
rect 19405 425 19445 430
rect 19415 -145 19435 425
rect 19405 -150 19445 -145
rect 19405 -180 19410 -150
rect 19440 -180 19445 -150
rect 19405 -185 19445 -180
rect 18495 -470 18525 -465
rect 18495 -505 18525 -500
rect 18545 -475 18575 -465
rect 18545 -495 18550 -475
rect 18570 -495 18575 -475
rect 18545 -505 18575 -495
rect 19325 -470 19365 -465
rect 19325 -500 19330 -470
rect 19360 -500 19365 -470
rect 19325 -505 19365 -500
rect 18550 -545 18570 -505
rect 18540 -550 18580 -545
rect 18540 -580 18545 -550
rect 18575 -580 18580 -550
rect 18540 -585 18580 -580
rect 19030 -550 19070 -545
rect 19030 -580 19035 -550
rect 19065 -580 19070 -550
rect 19030 -585 19070 -580
rect 18020 -605 18060 -600
rect 18020 -635 18025 -605
rect 18055 -635 18060 -605
rect 18020 -645 18060 -635
rect 18020 -675 18025 -645
rect 18055 -675 18060 -645
rect 18020 -685 18060 -675
rect 17875 -705 17905 -695
rect 17875 -725 17880 -705
rect 17900 -725 17905 -705
rect 18020 -715 18025 -685
rect 18055 -715 18060 -685
rect 18020 -720 18060 -715
rect 18140 -605 18180 -600
rect 18140 -635 18145 -605
rect 18175 -635 18180 -605
rect 18140 -645 18180 -635
rect 18140 -675 18145 -645
rect 18175 -675 18180 -645
rect 18140 -685 18180 -675
rect 18140 -715 18145 -685
rect 18175 -715 18180 -685
rect 18140 -720 18180 -715
rect 18260 -605 18300 -600
rect 18260 -635 18265 -605
rect 18295 -635 18300 -605
rect 18260 -645 18300 -635
rect 18260 -675 18265 -645
rect 18295 -675 18300 -645
rect 18260 -685 18300 -675
rect 18260 -715 18265 -685
rect 18295 -715 18300 -685
rect 18260 -720 18300 -715
rect 18580 -605 18620 -600
rect 18580 -635 18585 -605
rect 18615 -635 18620 -605
rect 18580 -645 18620 -635
rect 18580 -675 18585 -645
rect 18615 -675 18620 -645
rect 18580 -685 18620 -675
rect 18580 -715 18585 -685
rect 18615 -715 18620 -685
rect 18580 -720 18620 -715
rect 18700 -605 18740 -600
rect 18700 -635 18705 -605
rect 18735 -635 18740 -605
rect 18700 -645 18740 -635
rect 18700 -675 18705 -645
rect 18735 -675 18740 -645
rect 18700 -685 18740 -675
rect 18700 -715 18705 -685
rect 18735 -715 18740 -685
rect 18700 -720 18740 -715
rect 18820 -605 18860 -600
rect 18820 -635 18825 -605
rect 18855 -635 18860 -605
rect 18820 -645 18860 -635
rect 18820 -675 18825 -645
rect 18855 -675 18860 -645
rect 18820 -685 18860 -675
rect 18820 -715 18825 -685
rect 18855 -715 18860 -685
rect 18820 -720 18860 -715
rect 18940 -605 18980 -600
rect 18940 -635 18945 -605
rect 18975 -635 18980 -605
rect 18940 -645 18980 -635
rect 18940 -675 18945 -645
rect 18975 -675 18980 -645
rect 18940 -685 18980 -675
rect 18940 -715 18945 -685
rect 18975 -715 18980 -685
rect 19040 -700 19060 -585
rect 18940 -720 18980 -715
rect 19030 -710 19070 -700
rect 17875 -735 17905 -725
rect 19030 -730 19040 -710
rect 19060 -730 19070 -710
rect 19030 -740 19070 -730
rect 17740 -1035 17745 -1005
rect 17775 -1035 17785 -1005
rect 17815 -1035 17825 -1005
rect 17855 -1035 17860 -1005
rect 17740 -1045 17860 -1035
rect 17740 -1075 17745 -1045
rect 17775 -1075 17785 -1045
rect 17815 -1075 17825 -1045
rect 17855 -1075 17860 -1045
rect 17740 -1085 17860 -1075
rect 17740 -1115 17745 -1085
rect 17775 -1115 17785 -1085
rect 17815 -1115 17825 -1085
rect 17855 -1115 17860 -1085
rect 17740 -1120 17860 -1115
rect 18450 -1005 18490 -1000
rect 18450 -1035 18455 -1005
rect 18485 -1035 18490 -1005
rect 18450 -1045 18490 -1035
rect 18450 -1075 18455 -1045
rect 18485 -1075 18490 -1045
rect 18450 -1085 18490 -1075
rect 18450 -1115 18455 -1085
rect 18485 -1115 18490 -1085
rect 18450 -1120 18490 -1115
rect 16740 -1140 16780 -1135
rect 16740 -1170 16745 -1140
rect 16775 -1170 16780 -1140
rect 16740 -1175 16780 -1170
rect 16820 -1140 16860 -1135
rect 16820 -1170 16825 -1140
rect 16855 -1170 16860 -1140
rect 16820 -1175 16860 -1170
rect 16900 -1140 16940 -1135
rect 16900 -1170 16905 -1140
rect 16935 -1170 16940 -1140
rect 16900 -1175 16940 -1170
rect 16980 -1140 17020 -1135
rect 16980 -1170 16985 -1140
rect 17015 -1170 17020 -1140
rect 16980 -1175 17020 -1170
rect 17060 -1140 17100 -1135
rect 17060 -1170 17065 -1140
rect 17095 -1170 17100 -1140
rect 17060 -1175 17100 -1170
rect 17140 -1140 17180 -1135
rect 17140 -1170 17145 -1140
rect 17175 -1170 17180 -1140
rect 17140 -1175 17180 -1170
rect 17220 -1140 17260 -1135
rect 17220 -1170 17225 -1140
rect 17255 -1170 17260 -1140
rect 17220 -1175 17260 -1170
rect 17300 -1140 17340 -1135
rect 17300 -1170 17305 -1140
rect 17335 -1170 17340 -1140
rect 17300 -1175 17340 -1170
rect 17380 -1140 17420 -1135
rect 17380 -1170 17385 -1140
rect 17415 -1170 17420 -1140
rect 17380 -1175 17420 -1170
rect 17460 -1140 17500 -1135
rect 17460 -1170 17465 -1140
rect 17495 -1170 17500 -1140
rect 17460 -1175 17500 -1170
rect 17540 -1140 17580 -1135
rect 17540 -1170 17545 -1140
rect 17575 -1170 17580 -1140
rect 17540 -1175 17580 -1170
rect 17620 -1140 17660 -1135
rect 17620 -1170 17625 -1140
rect 17655 -1170 17660 -1140
rect 17620 -1175 17660 -1170
rect 17700 -1140 17740 -1135
rect 17700 -1170 17705 -1140
rect 17735 -1170 17740 -1140
rect 17700 -1175 17740 -1170
rect 17780 -1140 17820 -1135
rect 17780 -1170 17785 -1140
rect 17815 -1170 17820 -1140
rect 17780 -1175 17820 -1170
rect 17860 -1140 17900 -1135
rect 17860 -1170 17865 -1140
rect 17895 -1170 17900 -1140
rect 17860 -1175 17900 -1170
rect 17940 -1140 17980 -1135
rect 17940 -1170 17945 -1140
rect 17975 -1170 17980 -1140
rect 17940 -1175 17980 -1170
rect 18020 -1140 18060 -1135
rect 18020 -1170 18025 -1140
rect 18055 -1170 18060 -1140
rect 18020 -1175 18060 -1170
rect 18100 -1140 18140 -1135
rect 18100 -1170 18105 -1140
rect 18135 -1170 18140 -1140
rect 18100 -1175 18140 -1170
rect 18180 -1140 18220 -1135
rect 18180 -1170 18185 -1140
rect 18215 -1170 18220 -1140
rect 18180 -1175 18220 -1170
rect 18260 -1140 18300 -1135
rect 18260 -1170 18265 -1140
rect 18295 -1170 18300 -1140
rect 18260 -1175 18300 -1170
rect 18340 -1140 18380 -1135
rect 18340 -1170 18345 -1140
rect 18375 -1170 18380 -1140
rect 18340 -1175 18380 -1170
rect 18420 -1140 18460 -1135
rect 18420 -1170 18425 -1140
rect 18455 -1170 18460 -1140
rect 18420 -1175 18460 -1170
rect 18500 -1140 18540 -1135
rect 18500 -1170 18505 -1140
rect 18535 -1170 18540 -1140
rect 18500 -1175 18540 -1170
rect 18580 -1140 18620 -1135
rect 18580 -1170 18585 -1140
rect 18615 -1170 18620 -1140
rect 18580 -1175 18620 -1170
rect 18660 -1140 18700 -1135
rect 18660 -1170 18665 -1140
rect 18695 -1170 18700 -1140
rect 18660 -1175 18700 -1170
rect 18740 -1140 18780 -1135
rect 18740 -1170 18745 -1140
rect 18775 -1170 18780 -1140
rect 18740 -1175 18780 -1170
rect 18895 -1205 18935 -1200
rect 16700 -1225 16740 -1220
rect 16700 -1255 16705 -1225
rect 16735 -1255 16740 -1225
rect 16700 -1260 16740 -1255
rect 18895 -1235 18900 -1205
rect 18930 -1235 18935 -1205
rect 18895 -1245 18935 -1235
rect 18895 -1275 18900 -1245
rect 18930 -1275 18935 -1245
rect 18895 -1280 18935 -1275
rect 16595 -1325 16635 -1320
rect 16595 -1355 16600 -1325
rect 16630 -1355 16635 -1325
rect 16595 -1360 16635 -1355
rect 16705 -1325 16745 -1320
rect 16705 -1355 16710 -1325
rect 16740 -1355 16745 -1325
rect 16705 -1360 16745 -1355
rect 17300 -1325 17340 -1320
rect 17300 -1355 17305 -1325
rect 17335 -1355 17340 -1325
rect 17300 -1360 17340 -1355
rect 17780 -1325 17820 -1320
rect 17780 -1355 17785 -1325
rect 17815 -1355 17820 -1325
rect 17780 -1360 17820 -1355
rect 18260 -1325 18300 -1320
rect 18260 -1355 18265 -1325
rect 18295 -1355 18300 -1325
rect 18260 -1360 18300 -1355
rect 16540 -1410 16580 -1405
rect 16540 -1440 16545 -1410
rect 16575 -1440 16580 -1410
rect 16540 -1450 16580 -1440
rect 16540 -1480 16545 -1450
rect 16575 -1480 16580 -1450
rect 16540 -1490 16580 -1480
rect 16605 -1485 16625 -1360
rect 16650 -1410 16690 -1405
rect 16650 -1440 16655 -1410
rect 16685 -1440 16690 -1410
rect 16650 -1450 16690 -1440
rect 16650 -1480 16655 -1450
rect 16685 -1480 16690 -1450
rect 16540 -1520 16545 -1490
rect 16575 -1520 16580 -1490
rect 16540 -1525 16580 -1520
rect 16600 -1495 16630 -1485
rect 16600 -1515 16605 -1495
rect 16625 -1515 16630 -1495
rect 16600 -1525 16630 -1515
rect 16650 -1490 16690 -1480
rect 16715 -1485 16735 -1360
rect 16760 -1410 16800 -1405
rect 16760 -1440 16765 -1410
rect 16795 -1440 16800 -1410
rect 16760 -1450 16800 -1440
rect 16760 -1480 16765 -1450
rect 16795 -1480 16800 -1450
rect 16650 -1520 16655 -1490
rect 16685 -1520 16690 -1490
rect 16650 -1525 16690 -1520
rect 16710 -1495 16740 -1485
rect 16710 -1515 16715 -1495
rect 16735 -1515 16740 -1495
rect 16710 -1525 16740 -1515
rect 16760 -1490 16800 -1480
rect 16760 -1520 16765 -1490
rect 16795 -1520 16800 -1490
rect 16760 -1525 16800 -1520
rect 16820 -1410 16860 -1405
rect 16820 -1440 16825 -1410
rect 16855 -1440 16860 -1410
rect 16820 -1450 16860 -1440
rect 16820 -1480 16825 -1450
rect 16855 -1480 16860 -1450
rect 16820 -1490 16860 -1480
rect 16820 -1520 16825 -1490
rect 16855 -1520 16860 -1490
rect 16820 -1525 16860 -1520
rect 17025 -1410 17065 -1405
rect 17025 -1440 17030 -1410
rect 17060 -1440 17065 -1410
rect 17025 -1450 17065 -1440
rect 17025 -1480 17030 -1450
rect 17060 -1480 17065 -1450
rect 17025 -1490 17065 -1480
rect 17025 -1520 17030 -1490
rect 17060 -1520 17065 -1490
rect 17025 -1525 17065 -1520
rect 17135 -1410 17175 -1405
rect 17135 -1440 17140 -1410
rect 17170 -1440 17175 -1410
rect 17135 -1450 17175 -1440
rect 17135 -1480 17140 -1450
rect 17170 -1480 17175 -1450
rect 17135 -1490 17175 -1480
rect 17135 -1520 17140 -1490
rect 17170 -1520 17175 -1490
rect 17135 -1525 17175 -1520
rect 17245 -1410 17285 -1405
rect 17245 -1440 17250 -1410
rect 17280 -1440 17285 -1410
rect 17245 -1450 17285 -1440
rect 17245 -1480 17250 -1450
rect 17280 -1480 17285 -1450
rect 17245 -1490 17285 -1480
rect 17310 -1485 17330 -1360
rect 17355 -1410 17395 -1405
rect 17355 -1440 17360 -1410
rect 17390 -1440 17395 -1410
rect 17355 -1450 17395 -1440
rect 17355 -1480 17360 -1450
rect 17390 -1480 17395 -1450
rect 17245 -1520 17250 -1490
rect 17280 -1520 17285 -1490
rect 17245 -1525 17285 -1520
rect 17305 -1495 17335 -1485
rect 17305 -1515 17310 -1495
rect 17330 -1515 17335 -1495
rect 17305 -1525 17335 -1515
rect 17355 -1490 17395 -1480
rect 17355 -1520 17360 -1490
rect 17390 -1520 17395 -1490
rect 17355 -1525 17395 -1520
rect 17465 -1410 17505 -1405
rect 17465 -1440 17470 -1410
rect 17500 -1440 17505 -1410
rect 17465 -1450 17505 -1440
rect 17465 -1480 17470 -1450
rect 17500 -1480 17505 -1450
rect 17465 -1490 17505 -1480
rect 17465 -1520 17470 -1490
rect 17500 -1520 17505 -1490
rect 17465 -1525 17505 -1520
rect 17615 -1410 17655 -1405
rect 17615 -1440 17620 -1410
rect 17650 -1440 17655 -1410
rect 17615 -1450 17655 -1440
rect 17615 -1480 17620 -1450
rect 17650 -1480 17655 -1450
rect 17615 -1490 17655 -1480
rect 17615 -1520 17620 -1490
rect 17650 -1520 17655 -1490
rect 17615 -1525 17655 -1520
rect 17725 -1410 17765 -1405
rect 17725 -1440 17730 -1410
rect 17760 -1440 17765 -1410
rect 17725 -1450 17765 -1440
rect 17725 -1480 17730 -1450
rect 17760 -1480 17765 -1450
rect 17725 -1490 17765 -1480
rect 17790 -1485 17810 -1360
rect 17835 -1410 17875 -1405
rect 17835 -1440 17840 -1410
rect 17870 -1440 17875 -1410
rect 17835 -1450 17875 -1440
rect 17835 -1480 17840 -1450
rect 17870 -1480 17875 -1450
rect 17725 -1520 17730 -1490
rect 17760 -1520 17765 -1490
rect 17725 -1525 17765 -1520
rect 17785 -1495 17815 -1485
rect 17785 -1515 17790 -1495
rect 17810 -1515 17815 -1495
rect 17785 -1525 17815 -1515
rect 17835 -1490 17875 -1480
rect 17835 -1520 17840 -1490
rect 17870 -1520 17875 -1490
rect 17835 -1525 17875 -1520
rect 17945 -1410 17985 -1405
rect 17945 -1440 17950 -1410
rect 17980 -1440 17985 -1410
rect 17945 -1450 17985 -1440
rect 17945 -1480 17950 -1450
rect 17980 -1480 17985 -1450
rect 17945 -1490 17985 -1480
rect 17945 -1520 17950 -1490
rect 17980 -1520 17985 -1490
rect 17945 -1525 17985 -1520
rect 18095 -1410 18135 -1405
rect 18095 -1440 18100 -1410
rect 18130 -1440 18135 -1410
rect 18095 -1450 18135 -1440
rect 18095 -1480 18100 -1450
rect 18130 -1480 18135 -1450
rect 18095 -1490 18135 -1480
rect 18095 -1520 18100 -1490
rect 18130 -1520 18135 -1490
rect 18095 -1525 18135 -1520
rect 18205 -1410 18245 -1405
rect 18205 -1440 18210 -1410
rect 18240 -1440 18245 -1410
rect 18205 -1450 18245 -1440
rect 18205 -1480 18210 -1450
rect 18240 -1480 18245 -1450
rect 18205 -1490 18245 -1480
rect 18270 -1485 18290 -1360
rect 18315 -1410 18355 -1405
rect 18315 -1440 18320 -1410
rect 18350 -1440 18355 -1410
rect 18315 -1450 18355 -1440
rect 18315 -1480 18320 -1450
rect 18350 -1480 18355 -1450
rect 18205 -1520 18210 -1490
rect 18240 -1520 18245 -1490
rect 18205 -1525 18245 -1520
rect 18265 -1495 18295 -1485
rect 18265 -1515 18270 -1495
rect 18290 -1515 18295 -1495
rect 18265 -1525 18295 -1515
rect 18315 -1490 18355 -1480
rect 18315 -1520 18320 -1490
rect 18350 -1520 18355 -1490
rect 18315 -1525 18355 -1520
rect 18425 -1410 18465 -1405
rect 18425 -1440 18430 -1410
rect 18460 -1440 18465 -1410
rect 18425 -1450 18465 -1440
rect 18425 -1480 18430 -1450
rect 18460 -1480 18465 -1450
rect 18425 -1490 18465 -1480
rect 18425 -1520 18430 -1490
rect 18460 -1520 18465 -1490
rect 18425 -1525 18465 -1520
rect 18535 -1410 18575 -1405
rect 18535 -1440 18540 -1410
rect 18570 -1440 18575 -1410
rect 18535 -1450 18575 -1440
rect 18535 -1480 18540 -1450
rect 18570 -1480 18575 -1450
rect 18535 -1490 18575 -1480
rect 18535 -1520 18540 -1490
rect 18570 -1520 18575 -1490
rect 18535 -1525 18575 -1520
rect 17195 -1555 17225 -1545
rect 17195 -1575 17200 -1555
rect 17220 -1575 17225 -1555
rect 17195 -1605 17225 -1575
rect 17195 -1625 17200 -1605
rect 17220 -1625 17225 -1605
rect 17195 -1655 17225 -1625
rect 17415 -1555 17445 -1545
rect 17415 -1575 17420 -1555
rect 17440 -1575 17445 -1555
rect 17415 -1605 17445 -1575
rect 17415 -1625 17420 -1605
rect 17440 -1625 17445 -1605
rect 17415 -1655 17445 -1625
rect 18155 -1555 18185 -1545
rect 18155 -1575 18160 -1555
rect 18180 -1575 18185 -1555
rect 18155 -1605 18185 -1575
rect 18155 -1625 18160 -1605
rect 18180 -1625 18185 -1605
rect 18155 -1655 18185 -1625
rect 18375 -1555 18405 -1545
rect 18375 -1575 18380 -1555
rect 18400 -1575 18405 -1555
rect 18375 -1605 18405 -1575
rect 18375 -1625 18380 -1605
rect 18400 -1625 18405 -1605
rect 18375 -1655 18405 -1625
rect 16705 -1665 16745 -1655
rect 16705 -1685 16715 -1665
rect 16735 -1685 16745 -1665
rect 16705 -1695 16745 -1685
rect 17080 -1665 17120 -1655
rect 17080 -1685 17090 -1665
rect 17110 -1685 17120 -1665
rect 17080 -1695 17120 -1685
rect 17190 -1660 17230 -1655
rect 17190 -1690 17195 -1660
rect 17225 -1690 17230 -1660
rect 16715 -1895 16735 -1695
rect 17090 -1710 17110 -1695
rect 17080 -1715 17120 -1710
rect 17080 -1745 17085 -1715
rect 17115 -1745 17120 -1715
rect 17080 -1750 17120 -1745
rect 17190 -1770 17230 -1690
rect 17300 -1665 17340 -1655
rect 17300 -1685 17310 -1665
rect 17330 -1685 17340 -1665
rect 17300 -1695 17340 -1685
rect 17410 -1660 17450 -1655
rect 17410 -1690 17415 -1660
rect 17445 -1690 17450 -1660
rect 17410 -1695 17450 -1690
rect 17670 -1660 17710 -1655
rect 17670 -1690 17675 -1660
rect 17705 -1690 17710 -1660
rect 17670 -1695 17710 -1690
rect 17780 -1660 17820 -1655
rect 17780 -1690 17785 -1660
rect 17815 -1690 17820 -1660
rect 17780 -1695 17820 -1690
rect 17890 -1660 17930 -1655
rect 17890 -1690 17895 -1660
rect 17925 -1690 17930 -1660
rect 17890 -1695 17930 -1690
rect 18150 -1660 18190 -1655
rect 18150 -1690 18155 -1660
rect 18185 -1690 18190 -1660
rect 18150 -1695 18190 -1690
rect 18260 -1665 18300 -1655
rect 18260 -1685 18270 -1665
rect 18290 -1685 18300 -1665
rect 18260 -1695 18300 -1685
rect 18370 -1660 18410 -1655
rect 18370 -1690 18375 -1660
rect 18405 -1690 18410 -1660
rect 17310 -1710 17330 -1695
rect 17300 -1715 17340 -1710
rect 17300 -1745 17305 -1715
rect 17335 -1745 17340 -1715
rect 17300 -1750 17340 -1745
rect 17190 -1800 17195 -1770
rect 17225 -1800 17230 -1770
rect 17190 -1810 17230 -1800
rect 17190 -1840 17195 -1810
rect 17225 -1840 17230 -1810
rect 17190 -1845 17230 -1840
rect 17790 -1895 17810 -1695
rect 18270 -1710 18290 -1695
rect 18260 -1715 18300 -1710
rect 18260 -1745 18265 -1715
rect 18295 -1745 18300 -1715
rect 18260 -1750 18300 -1745
rect 18370 -1770 18410 -1690
rect 18480 -1665 18520 -1655
rect 18480 -1685 18490 -1665
rect 18510 -1685 18520 -1665
rect 18480 -1695 18520 -1685
rect 18490 -1710 18510 -1695
rect 18480 -1715 18520 -1710
rect 18480 -1745 18485 -1715
rect 18515 -1745 18520 -1715
rect 18480 -1750 18520 -1745
rect 18370 -1800 18375 -1770
rect 18405 -1800 18410 -1770
rect 18370 -1810 18410 -1800
rect 18370 -1840 18375 -1810
rect 18405 -1840 18410 -1810
rect 18370 -1845 18410 -1840
rect 16705 -1900 16745 -1895
rect 16705 -1930 16710 -1900
rect 16740 -1930 16745 -1900
rect 16705 -1935 16745 -1930
rect 17780 -1900 17820 -1895
rect 17780 -1930 17785 -1900
rect 17815 -1930 17820 -1900
rect 17780 -1935 17820 -1930
rect 19335 -1945 19355 -505
rect 19325 -1950 19365 -1945
rect 19325 -1980 19330 -1950
rect 19360 -1980 19365 -1950
rect 19325 -1985 19365 -1980
rect 16260 -2000 16300 -1995
rect 16260 -2030 16265 -2000
rect 16295 -2030 16300 -2000
rect 16260 -2035 16300 -2030
rect 16480 -2000 16520 -1995
rect 16480 -2030 16485 -2000
rect 16515 -2030 16520 -2000
rect 16480 -2035 16520 -2030
rect 16730 -2000 16770 -1995
rect 16730 -2030 16735 -2000
rect 16765 -2030 16770 -2000
rect 16730 -2035 16770 -2030
rect 17195 -2000 17235 -1995
rect 17195 -2030 17200 -2000
rect 17230 -2030 17235 -2000
rect 16490 -2895 16510 -2035
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 16160 -3025 16195 -3020
rect 16160 -3065 16195 -3060
rect 16740 -3100 16760 -2035
rect 17195 -2060 17235 -2030
rect 17425 -2035 17430 -2000
rect 17465 -2035 17470 -2000
rect 18124 -2035 18129 -2000
rect 18164 -2035 18169 -2000
rect 19080 -2005 19120 -2000
rect 19080 -2035 19085 -2005
rect 19115 -2035 19120 -2005
rect 17195 -2090 17200 -2060
rect 17230 -2090 17235 -2060
rect 17195 -2095 17235 -2090
rect 18830 -2060 18870 -2055
rect 18830 -2090 18835 -2060
rect 18865 -2090 18870 -2060
rect 18830 -2095 18870 -2090
rect 16945 -2615 18655 -2265
rect 16730 -3105 16770 -3100
rect 15820 -3145 15825 -3115
rect 15855 -3145 15860 -3115
rect 15820 -3150 15860 -3145
rect 15950 -3116 15985 -3111
rect 16730 -3135 16735 -3105
rect 16765 -3135 16770 -3105
rect 16730 -3140 16770 -3135
rect 15830 -4260 15850 -3150
rect 15950 -3156 15985 -3151
rect 16945 -3625 17295 -2615
rect 17625 -3105 17975 -2945
rect 17625 -3135 17785 -3105
rect 17815 -3135 17975 -3105
rect 17625 -3295 17975 -3135
rect 18305 -3105 18655 -2615
rect 18840 -3100 18860 -2095
rect 19080 -2895 19120 -2035
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19415 -2992 19435 -185
rect 19460 -2005 19500 575
rect 19545 -1895 19565 1755
rect 19610 410 19650 415
rect 19610 380 19615 410
rect 19645 380 19650 410
rect 19610 375 19650 380
rect 19535 -1900 19575 -1895
rect 19535 -1930 19540 -1900
rect 19570 -1930 19575 -1900
rect 19535 -1935 19575 -1930
rect 19460 -2035 19465 -2005
rect 19495 -2035 19500 -2005
rect 19460 -2040 19500 -2035
rect 19405 -2997 19440 -2992
rect 19405 -3037 19440 -3032
rect 18305 -3135 18620 -3105
rect 18650 -3135 18655 -3105
rect 18305 -3625 18655 -3135
rect 18830 -3105 18870 -3100
rect 18830 -3135 18835 -3105
rect 18865 -3135 18870 -3105
rect 19620 -3111 19640 375
rect 19720 -95 19760 -90
rect 19720 -125 19725 -95
rect 19755 -125 19760 -95
rect 19720 -130 19760 -125
rect 18830 -3140 18870 -3135
rect 19610 -3116 19645 -3111
rect 19610 -3156 19645 -3151
rect 15950 -3789 15985 -3784
rect 15950 -3829 15985 -3824
rect 15820 -4265 15860 -4260
rect 15820 -4295 15825 -4265
rect 15855 -4295 15860 -4265
rect 15820 -4300 15860 -4295
rect 15725 -4315 15765 -4310
rect 15725 -4345 15730 -4315
rect 15760 -4345 15765 -4315
rect 15725 -4350 15765 -4345
rect 15960 -4355 15980 -3829
rect 16280 -3894 16315 -3889
rect 16280 -3934 16315 -3929
rect 16290 -4185 16310 -3934
rect 16605 -3969 16640 -3964
rect 16945 -3975 18655 -3625
rect 19610 -3789 19645 -3784
rect 19610 -3829 19645 -3824
rect 19285 -3894 19320 -3889
rect 19285 -3934 19320 -3929
rect 18960 -3969 18995 -3964
rect 16605 -4009 16640 -4004
rect 18960 -4009 18995 -4004
rect 16615 -4185 16635 -4009
rect 16280 -4190 16320 -4185
rect 16280 -4220 16285 -4190
rect 16315 -4220 16320 -4190
rect 16280 -4225 16320 -4220
rect 16605 -4190 16645 -4185
rect 16605 -4220 16610 -4190
rect 16640 -4220 16645 -4190
rect 16605 -4225 16645 -4220
rect 17250 -4265 17300 -4255
rect 18965 -4260 18985 -4009
rect 19290 -4260 19310 -3934
rect 17250 -4295 17260 -4265
rect 17290 -4295 17300 -4265
rect 17250 -4305 17300 -4295
rect 17780 -4265 17820 -4260
rect 17780 -4295 17785 -4265
rect 17815 -4295 17820 -4265
rect 17780 -4300 17820 -4295
rect 18955 -4265 18995 -4260
rect 18955 -4295 18960 -4265
rect 18990 -4295 18995 -4265
rect 18955 -4300 18995 -4295
rect 19280 -4265 19320 -4260
rect 19280 -4295 19285 -4265
rect 19315 -4295 19320 -4265
rect 19280 -4300 19320 -4295
rect 16900 -4315 16950 -4305
rect 16900 -4345 16910 -4315
rect 16940 -4345 16950 -4315
rect 16900 -4355 16950 -4345
rect 18650 -4315 18700 -4305
rect 18650 -4345 18660 -4315
rect 18690 -4345 18700 -4315
rect 18650 -4355 18700 -4345
rect 19620 -4355 19640 -3829
rect 19730 -4310 19750 -130
rect 19775 -1770 19815 1755
rect 19775 -1800 19780 -1770
rect 19810 -1800 19815 -1770
rect 19775 -1810 19815 -1800
rect 19775 -1840 19780 -1810
rect 19810 -1840 19815 -1810
rect 19775 -1845 19815 -1840
rect 19720 -4315 19760 -4310
rect 19720 -4345 19725 -4315
rect 19755 -4345 19760 -4315
rect 19720 -4350 19760 -4345
rect 15950 -4360 15990 -4355
rect 15950 -4390 15955 -4360
rect 15985 -4390 15990 -4360
rect 15950 -4395 15990 -4390
rect 16205 -4360 16245 -4355
rect 16205 -4390 16210 -4360
rect 16240 -4390 16245 -4360
rect 16205 -4395 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4390 19395 -4360
rect 19355 -4395 19395 -4390
rect 19610 -4360 19650 -4355
rect 19610 -4390 19615 -4360
rect 19645 -4390 19650 -4360
rect 19610 -4395 19650 -4390
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4440 17995 -4410
rect 17955 -4445 17995 -4440
<< via1 >>
rect 15730 -125 15760 -95
rect 15955 105 15985 135
rect 15790 -1800 15820 -1770
rect 15790 -1840 15820 -1810
rect 16035 -1745 16065 -1715
rect 16945 1635 16975 1665
rect 16490 1615 16520 1620
rect 16490 1595 16495 1615
rect 16495 1595 16515 1615
rect 16515 1595 16520 1615
rect 16490 1590 16520 1595
rect 16370 1490 16400 1520
rect 16370 1450 16400 1480
rect 16370 1435 16400 1440
rect 16370 1415 16375 1435
rect 16375 1415 16395 1435
rect 16395 1415 16400 1435
rect 16370 1410 16400 1415
rect 16490 1490 16520 1520
rect 16490 1450 16520 1480
rect 16490 1435 16520 1440
rect 16490 1415 16495 1435
rect 16495 1415 16515 1435
rect 16515 1415 16520 1435
rect 16490 1410 16520 1415
rect 16610 1490 16640 1520
rect 16610 1450 16640 1480
rect 16610 1435 16640 1440
rect 16610 1415 16615 1435
rect 16615 1415 16635 1435
rect 16635 1415 16640 1435
rect 16610 1410 16640 1415
rect 16890 1490 16920 1520
rect 16890 1450 16920 1480
rect 17055 1590 17085 1620
rect 17000 1490 17030 1520
rect 17000 1450 17030 1480
rect 16890 1435 16920 1440
rect 16890 1415 16895 1435
rect 16895 1415 16915 1435
rect 16915 1415 16920 1435
rect 16890 1410 16920 1415
rect 17110 1490 17140 1520
rect 17110 1450 17140 1480
rect 17000 1435 17030 1440
rect 17000 1415 17005 1435
rect 17005 1415 17025 1435
rect 17025 1415 17030 1435
rect 17000 1410 17030 1415
rect 17110 1435 17140 1440
rect 17110 1415 17115 1435
rect 17115 1415 17135 1435
rect 17135 1415 17140 1435
rect 17110 1410 17140 1415
rect 17220 1490 17250 1520
rect 17220 1450 17250 1480
rect 17220 1435 17250 1440
rect 17220 1415 17225 1435
rect 17225 1415 17245 1435
rect 17245 1415 17250 1435
rect 17220 1410 17250 1415
rect 17500 1490 17530 1520
rect 17500 1450 17530 1480
rect 17500 1435 17530 1440
rect 17500 1415 17505 1435
rect 17505 1415 17525 1435
rect 17525 1415 17530 1435
rect 17500 1410 17530 1415
rect 17565 1490 17595 1520
rect 17565 1450 17595 1480
rect 17565 1435 17595 1440
rect 17565 1415 17570 1435
rect 17570 1415 17590 1435
rect 17590 1415 17595 1435
rect 17565 1410 17595 1415
rect 17675 1490 17705 1520
rect 17675 1450 17705 1480
rect 17675 1435 17705 1440
rect 17675 1415 17680 1435
rect 17680 1415 17700 1435
rect 17700 1415 17705 1435
rect 17675 1410 17705 1415
rect 17785 1615 17815 1620
rect 17785 1595 17790 1615
rect 17790 1595 17810 1615
rect 17810 1595 17815 1615
rect 17785 1590 17815 1595
rect 17785 1490 17815 1520
rect 17785 1450 17815 1480
rect 17785 1435 17815 1440
rect 17785 1415 17790 1435
rect 17790 1415 17810 1435
rect 17810 1415 17815 1435
rect 17785 1410 17815 1415
rect 17895 1490 17925 1520
rect 17895 1450 17925 1480
rect 17895 1435 17925 1440
rect 17895 1415 17900 1435
rect 17900 1415 17920 1435
rect 17920 1415 17925 1435
rect 17895 1410 17925 1415
rect 18625 1635 18655 1665
rect 18205 1590 18235 1620
rect 18515 1590 18545 1620
rect 18005 1490 18035 1520
rect 18005 1450 18035 1480
rect 18005 1435 18035 1440
rect 18005 1415 18010 1435
rect 18010 1415 18030 1435
rect 18030 1415 18035 1435
rect 18005 1410 18035 1415
rect 18070 1490 18100 1520
rect 18070 1450 18100 1480
rect 18070 1435 18100 1440
rect 18070 1415 18075 1435
rect 18075 1415 18095 1435
rect 18095 1415 18100 1435
rect 18070 1410 18100 1415
rect 16435 1265 16465 1270
rect 16435 1245 16440 1265
rect 16440 1245 16460 1265
rect 16460 1245 16465 1265
rect 16435 1240 16465 1245
rect 16545 1265 16575 1270
rect 16545 1245 16550 1265
rect 16550 1245 16570 1265
rect 16570 1245 16575 1265
rect 16545 1240 16575 1245
rect 16945 1265 16975 1270
rect 16945 1245 16950 1265
rect 16950 1245 16970 1265
rect 16970 1245 16975 1265
rect 16945 1240 16975 1245
rect 17055 1265 17085 1270
rect 17055 1245 17060 1265
rect 17060 1245 17080 1265
rect 17080 1245 17085 1265
rect 17055 1240 17085 1245
rect 17165 1265 17195 1270
rect 17165 1245 17170 1265
rect 17170 1245 17190 1265
rect 17190 1245 17195 1265
rect 17165 1240 17195 1245
rect 17620 1265 17650 1270
rect 17620 1245 17625 1265
rect 17625 1245 17645 1265
rect 17645 1245 17650 1265
rect 17620 1240 17650 1245
rect 17730 1265 17760 1270
rect 17730 1245 17735 1265
rect 17735 1245 17755 1265
rect 17755 1245 17760 1265
rect 17730 1240 17760 1245
rect 17840 1265 17870 1270
rect 17840 1245 17845 1265
rect 17845 1245 17865 1265
rect 17865 1245 17870 1265
rect 17840 1240 17870 1245
rect 17950 1265 17980 1270
rect 17950 1245 17955 1265
rect 17955 1245 17975 1265
rect 17975 1245 17980 1265
rect 17950 1240 17980 1245
rect 18350 1490 18380 1520
rect 18350 1450 18380 1480
rect 18350 1435 18380 1440
rect 18350 1415 18355 1435
rect 18355 1415 18375 1435
rect 18375 1415 18380 1435
rect 18350 1410 18380 1415
rect 18460 1490 18490 1520
rect 18460 1450 18490 1480
rect 18570 1490 18600 1520
rect 18570 1450 18600 1480
rect 18460 1435 18490 1440
rect 18460 1415 18465 1435
rect 18465 1415 18485 1435
rect 18485 1415 18490 1435
rect 18460 1410 18490 1415
rect 18680 1490 18710 1520
rect 18680 1450 18710 1480
rect 18570 1435 18600 1440
rect 18570 1415 18575 1435
rect 18575 1415 18595 1435
rect 18595 1415 18600 1435
rect 18570 1410 18600 1415
rect 18680 1435 18710 1440
rect 18680 1415 18685 1435
rect 18685 1415 18705 1435
rect 18705 1415 18710 1435
rect 18680 1410 18710 1415
rect 18405 1265 18435 1270
rect 18405 1245 18410 1265
rect 18410 1245 18430 1265
rect 18430 1245 18435 1265
rect 18405 1240 18435 1245
rect 18515 1265 18545 1270
rect 18515 1245 18520 1265
rect 18520 1245 18540 1265
rect 18540 1245 18545 1265
rect 18515 1240 18545 1245
rect 18625 1265 18655 1270
rect 18625 1245 18630 1265
rect 18630 1245 18650 1265
rect 18650 1245 18655 1265
rect 18625 1240 18655 1245
rect 18205 1185 18235 1215
rect 18725 1185 18755 1215
rect 16165 1140 16195 1170
rect 16435 1140 16465 1170
rect 16545 1140 16575 1170
rect 16440 1025 16470 1055
rect 16440 985 16470 1015
rect 16440 945 16470 975
rect 16660 1025 16690 1055
rect 16660 985 16690 1015
rect 16660 945 16690 975
rect 16975 1025 17005 1055
rect 16975 985 17005 1015
rect 16975 970 17005 975
rect 16975 950 16980 970
rect 16980 950 17000 970
rect 17000 950 17005 970
rect 16975 945 17005 950
rect 17155 1025 17185 1055
rect 17155 985 17185 1015
rect 17155 970 17185 975
rect 17155 950 17160 970
rect 17160 950 17180 970
rect 17180 950 17185 970
rect 17155 945 17185 950
rect 17335 1025 17365 1055
rect 17335 985 17365 1015
rect 17335 970 17365 975
rect 17335 950 17340 970
rect 17340 950 17360 970
rect 17360 950 17365 970
rect 17335 945 17365 950
rect 17515 1025 17545 1055
rect 17515 985 17545 1015
rect 17515 970 17545 975
rect 17515 950 17520 970
rect 17520 950 17540 970
rect 17540 950 17545 970
rect 17515 945 17545 950
rect 17695 1025 17725 1055
rect 17695 985 17725 1015
rect 17695 970 17725 975
rect 17695 950 17700 970
rect 17700 950 17720 970
rect 17720 950 17725 970
rect 17695 945 17725 950
rect 17875 1025 17905 1055
rect 17875 985 17905 1015
rect 17875 970 17905 975
rect 17875 950 17880 970
rect 17880 950 17900 970
rect 17900 950 17905 970
rect 17875 945 17905 950
rect 18055 1025 18085 1055
rect 18055 985 18085 1015
rect 18055 970 18085 975
rect 18055 950 18060 970
rect 18060 950 18080 970
rect 18080 950 18085 970
rect 18055 945 18085 950
rect 18235 1025 18265 1055
rect 18235 985 18265 1015
rect 18235 970 18265 975
rect 18235 950 18240 970
rect 18240 950 18260 970
rect 18260 950 18265 970
rect 18235 945 18265 950
rect 18415 1025 18445 1055
rect 18415 985 18445 1015
rect 18415 970 18445 975
rect 18415 950 18420 970
rect 18420 950 18440 970
rect 18440 950 18445 970
rect 18415 945 18445 950
rect 18595 1025 18625 1055
rect 18595 985 18625 1015
rect 18595 970 18625 975
rect 18595 950 18600 970
rect 18600 950 18620 970
rect 18620 950 18625 970
rect 18595 945 18625 950
rect 16550 870 16580 875
rect 16550 850 16555 870
rect 16555 850 16575 870
rect 16575 850 16580 870
rect 16550 845 16580 850
rect 16785 845 16815 875
rect 16485 700 16515 705
rect 16485 680 16490 700
rect 16490 680 16510 700
rect 16510 680 16515 700
rect 16485 675 16515 680
rect 16615 700 16645 705
rect 16615 680 16620 700
rect 16620 680 16640 700
rect 16640 680 16645 700
rect 16615 675 16645 680
rect 16320 575 16350 605
rect 16265 520 16295 550
rect 16210 475 16240 505
rect 16265 -180 16295 -150
rect 16210 -1255 16240 -1225
rect 16165 -1355 16195 -1325
rect 16110 -1930 16140 -1900
rect 16160 -1980 16190 -1950
rect 16845 675 16875 705
rect 16785 520 16815 550
rect 16550 475 16580 505
rect 16425 240 16455 270
rect 16425 200 16455 230
rect 16425 160 16455 190
rect 16545 240 16575 270
rect 16545 200 16575 230
rect 16545 160 16575 190
rect 16665 240 16695 270
rect 16665 200 16695 230
rect 16665 160 16695 190
rect 16785 240 16815 270
rect 16785 200 16815 230
rect 16785 160 16815 190
rect 17605 600 17635 605
rect 17605 580 17610 600
rect 17610 580 17630 600
rect 17630 580 17635 600
rect 17605 575 17635 580
rect 17965 600 17995 605
rect 17965 580 17970 600
rect 17970 580 17990 600
rect 17990 580 17995 600
rect 17965 575 17995 580
rect 17425 520 17455 550
rect 17245 475 17275 505
rect 17065 430 17095 460
rect 16905 240 16935 270
rect 16905 200 16935 230
rect 16905 160 16935 190
rect 17025 240 17055 270
rect 17025 200 17055 230
rect 17025 160 17055 190
rect 17145 240 17175 270
rect 17145 200 17175 230
rect 17145 160 17175 190
rect 17265 240 17295 270
rect 17265 200 17295 230
rect 17265 160 17295 190
rect 17385 240 17415 270
rect 17385 200 17415 230
rect 17385 160 17415 190
rect 17505 240 17535 270
rect 17505 200 17535 230
rect 17505 160 17535 190
rect 17625 240 17655 270
rect 17625 200 17655 230
rect 17625 160 17655 190
rect 18145 520 18175 550
rect 18325 475 18355 505
rect 17785 430 17815 460
rect 18505 430 18535 460
rect 18910 1025 18940 1055
rect 18910 985 18940 1015
rect 18910 970 18940 975
rect 18910 950 18915 970
rect 18915 950 18935 970
rect 18935 950 18940 970
rect 18910 945 18940 950
rect 19020 1025 19050 1055
rect 19020 985 19050 1015
rect 19020 970 19050 975
rect 19020 950 19025 970
rect 19025 950 19045 970
rect 19045 950 19050 970
rect 19020 945 19050 950
rect 19080 1025 19110 1055
rect 19080 985 19110 1015
rect 19080 970 19110 975
rect 19080 950 19085 970
rect 19085 950 19105 970
rect 19105 950 19110 970
rect 19080 945 19110 950
rect 19330 1140 19360 1170
rect 18955 700 18985 705
rect 18955 680 18960 700
rect 18960 680 18980 700
rect 18980 680 18985 700
rect 18955 675 18985 680
rect 19265 675 19295 705
rect 19005 650 19035 655
rect 19005 630 19010 650
rect 19010 630 19030 650
rect 19030 630 19035 650
rect 19005 625 19035 630
rect 18005 380 18035 410
rect 18725 380 18755 410
rect 19015 380 19045 410
rect 17945 240 17975 270
rect 17945 200 17975 230
rect 17945 160 17975 190
rect 18065 240 18095 270
rect 18065 200 18095 230
rect 18065 160 18095 190
rect 18185 240 18215 270
rect 18185 200 18215 230
rect 18185 160 18215 190
rect 18305 240 18335 270
rect 18305 200 18335 230
rect 18305 160 18335 190
rect 18425 240 18455 270
rect 18425 200 18455 230
rect 18425 160 18455 190
rect 18545 240 18575 270
rect 18545 200 18575 230
rect 18545 160 18575 190
rect 18665 240 18695 270
rect 18665 200 18695 230
rect 18665 160 18695 190
rect 18785 240 18815 270
rect 18785 200 18815 230
rect 18785 160 18815 190
rect 18905 240 18935 270
rect 18905 200 18935 230
rect 18905 160 18935 190
rect 19025 240 19055 270
rect 19025 200 19055 230
rect 19025 160 19055 190
rect 19145 240 19175 270
rect 19145 200 19175 230
rect 19145 160 19175 190
rect 16485 130 16515 135
rect 16485 110 16490 130
rect 16490 110 16510 130
rect 16510 110 16515 130
rect 16485 105 16515 110
rect 16845 130 16875 135
rect 16845 110 16850 130
rect 16850 110 16870 130
rect 16870 110 16875 130
rect 16845 105 16875 110
rect 17205 130 17235 135
rect 17205 110 17210 130
rect 17210 110 17230 130
rect 17230 110 17235 130
rect 17205 105 17235 110
rect 17565 130 17595 135
rect 17565 110 17570 130
rect 17570 110 17590 130
rect 17590 110 17595 130
rect 17565 105 17595 110
rect 17695 105 17725 135
rect 17875 105 17905 135
rect 16605 -40 16635 -35
rect 16605 -60 16610 -40
rect 16610 -60 16630 -40
rect 16630 -60 16635 -40
rect 16605 -65 16635 -60
rect 16965 -40 16995 -35
rect 16965 -60 16970 -40
rect 16970 -60 16990 -40
rect 16990 -60 16995 -40
rect 16965 -65 16995 -60
rect 17325 -40 17355 -35
rect 17325 -60 17330 -40
rect 17330 -60 17350 -40
rect 17350 -60 17355 -40
rect 17325 -65 17355 -60
rect 16515 -125 16545 -95
rect 16725 -125 16755 -95
rect 16845 -125 16875 -95
rect 17085 -125 17115 -95
rect 17205 -125 17235 -95
rect 17445 -125 17475 -95
rect 17535 -125 17565 -95
rect 17007 -155 17037 -150
rect 17007 -175 17012 -155
rect 17012 -175 17032 -155
rect 17032 -175 17037 -155
rect 17007 -180 17037 -175
rect 16320 -500 16350 -470
rect 17565 -215 17595 -210
rect 17565 -235 17570 -215
rect 17570 -235 17590 -215
rect 17590 -235 17595 -215
rect 17565 -240 17595 -235
rect 17565 -255 17595 -250
rect 17565 -275 17570 -255
rect 17570 -275 17590 -255
rect 17590 -275 17595 -255
rect 17565 -280 17595 -275
rect 17565 -295 17595 -290
rect 17565 -315 17570 -295
rect 17570 -315 17590 -295
rect 17590 -315 17595 -295
rect 17565 -320 17595 -315
rect 17075 -475 17105 -470
rect 17075 -495 17080 -475
rect 17080 -495 17100 -475
rect 17100 -495 17105 -475
rect 17075 -500 17105 -495
rect 16535 -580 16565 -550
rect 17025 -580 17055 -550
rect 16625 -635 16655 -605
rect 16625 -675 16655 -645
rect 16625 -690 16655 -685
rect 16625 -710 16630 -690
rect 16630 -710 16650 -690
rect 16650 -710 16655 -690
rect 16625 -715 16655 -710
rect 16745 -635 16775 -605
rect 16745 -675 16775 -645
rect 16745 -690 16775 -685
rect 16745 -710 16750 -690
rect 16750 -710 16770 -690
rect 16770 -710 16775 -690
rect 16745 -715 16775 -710
rect 16865 -635 16895 -605
rect 16865 -675 16895 -645
rect 16865 -690 16895 -685
rect 16865 -710 16870 -690
rect 16870 -710 16890 -690
rect 16890 -710 16895 -690
rect 16865 -715 16895 -710
rect 16985 -635 17015 -605
rect 16985 -675 17015 -645
rect 16985 -690 17015 -685
rect 16985 -710 16990 -690
rect 16990 -710 17010 -690
rect 17010 -710 17015 -690
rect 16985 -715 17015 -710
rect 17305 -635 17335 -605
rect 17305 -675 17335 -645
rect 17305 -690 17335 -685
rect 17305 -710 17310 -690
rect 17310 -710 17330 -690
rect 17330 -710 17335 -690
rect 17305 -715 17335 -710
rect 17425 -635 17455 -605
rect 17425 -675 17455 -645
rect 17425 -690 17455 -685
rect 17425 -710 17430 -690
rect 17430 -710 17450 -690
rect 17450 -710 17455 -690
rect 17425 -715 17455 -710
rect 17545 -635 17575 -605
rect 17545 -675 17575 -645
rect 17545 -690 17575 -685
rect 17545 -710 17550 -690
rect 17550 -710 17570 -690
rect 17570 -710 17575 -690
rect 17545 -715 17575 -710
rect 17745 -240 17775 -210
rect 17785 -240 17815 -210
rect 17825 -240 17855 -210
rect 17745 -280 17775 -250
rect 17785 -280 17815 -250
rect 17825 -280 17855 -250
rect 17745 -320 17775 -290
rect 17785 -320 17815 -290
rect 17825 -320 17855 -290
rect 17115 -1010 17145 -1005
rect 17115 -1030 17120 -1010
rect 17120 -1030 17140 -1010
rect 17140 -1030 17145 -1010
rect 17115 -1035 17145 -1030
rect 17115 -1075 17145 -1045
rect 17115 -1115 17145 -1085
rect 18005 130 18035 135
rect 18005 110 18010 130
rect 18010 110 18030 130
rect 18030 110 18035 130
rect 18005 105 18035 110
rect 18365 130 18395 135
rect 18365 110 18370 130
rect 18370 110 18390 130
rect 18390 110 18395 130
rect 18365 105 18395 110
rect 18725 130 18755 135
rect 18725 110 18730 130
rect 18730 110 18750 130
rect 18750 110 18755 130
rect 18725 105 18755 110
rect 19085 130 19115 135
rect 19085 110 19090 130
rect 19090 110 19110 130
rect 19110 110 19115 130
rect 19085 105 19115 110
rect 18245 -40 18275 -35
rect 18245 -60 18250 -40
rect 18250 -60 18270 -40
rect 18270 -60 18275 -40
rect 18245 -65 18275 -60
rect 18605 -40 18635 -35
rect 18605 -60 18610 -40
rect 18610 -60 18630 -40
rect 18630 -60 18635 -40
rect 18605 -65 18635 -60
rect 18965 -40 18995 -35
rect 18965 -60 18970 -40
rect 18970 -60 18990 -40
rect 18990 -60 18995 -40
rect 18965 -65 18995 -60
rect 18035 -125 18065 -95
rect 18125 -125 18155 -95
rect 18365 -125 18395 -95
rect 18485 -125 18515 -95
rect 18725 -125 18755 -95
rect 18845 -125 18875 -95
rect 19055 -125 19085 -95
rect 18563 -155 18593 -150
rect 18563 -175 18568 -155
rect 18568 -175 18588 -155
rect 18588 -175 18593 -155
rect 18563 -180 18593 -175
rect 18005 -215 18035 -210
rect 18005 -235 18010 -215
rect 18010 -235 18030 -215
rect 18030 -235 18035 -215
rect 18005 -240 18035 -235
rect 18005 -255 18035 -250
rect 18005 -275 18010 -255
rect 18010 -275 18030 -255
rect 18030 -275 18035 -255
rect 18005 -280 18035 -275
rect 18005 -295 18035 -290
rect 18005 -315 18010 -295
rect 18010 -315 18030 -295
rect 18030 -315 18035 -295
rect 18005 -320 18035 -315
rect 19465 575 19495 605
rect 19410 430 19440 460
rect 19410 -180 19440 -150
rect 18495 -475 18525 -470
rect 18495 -495 18500 -475
rect 18500 -495 18520 -475
rect 18520 -495 18525 -475
rect 18495 -500 18525 -495
rect 19330 -500 19360 -470
rect 18545 -580 18575 -550
rect 19035 -580 19065 -550
rect 18025 -635 18055 -605
rect 18025 -675 18055 -645
rect 18025 -690 18055 -685
rect 18025 -710 18030 -690
rect 18030 -710 18050 -690
rect 18050 -710 18055 -690
rect 18025 -715 18055 -710
rect 18145 -635 18175 -605
rect 18145 -675 18175 -645
rect 18145 -690 18175 -685
rect 18145 -710 18150 -690
rect 18150 -710 18170 -690
rect 18170 -710 18175 -690
rect 18145 -715 18175 -710
rect 18265 -635 18295 -605
rect 18265 -675 18295 -645
rect 18265 -690 18295 -685
rect 18265 -710 18270 -690
rect 18270 -710 18290 -690
rect 18290 -710 18295 -690
rect 18265 -715 18295 -710
rect 18585 -635 18615 -605
rect 18585 -675 18615 -645
rect 18585 -690 18615 -685
rect 18585 -710 18590 -690
rect 18590 -710 18610 -690
rect 18610 -710 18615 -690
rect 18585 -715 18615 -710
rect 18705 -635 18735 -605
rect 18705 -675 18735 -645
rect 18705 -690 18735 -685
rect 18705 -710 18710 -690
rect 18710 -710 18730 -690
rect 18730 -710 18735 -690
rect 18705 -715 18735 -710
rect 18825 -635 18855 -605
rect 18825 -675 18855 -645
rect 18825 -690 18855 -685
rect 18825 -710 18830 -690
rect 18830 -710 18850 -690
rect 18850 -710 18855 -690
rect 18825 -715 18855 -710
rect 18945 -635 18975 -605
rect 18945 -675 18975 -645
rect 18945 -690 18975 -685
rect 18945 -710 18950 -690
rect 18950 -710 18970 -690
rect 18970 -710 18975 -690
rect 18945 -715 18975 -710
rect 17745 -1035 17775 -1005
rect 17785 -1035 17815 -1005
rect 17825 -1035 17855 -1005
rect 17745 -1075 17775 -1045
rect 17785 -1075 17815 -1045
rect 17825 -1075 17855 -1045
rect 17745 -1115 17775 -1085
rect 17785 -1115 17815 -1085
rect 17825 -1115 17855 -1085
rect 18455 -1010 18485 -1005
rect 18455 -1030 18460 -1010
rect 18460 -1030 18480 -1010
rect 18480 -1030 18485 -1010
rect 18455 -1035 18485 -1030
rect 18455 -1075 18485 -1045
rect 18455 -1115 18485 -1085
rect 16745 -1145 16775 -1140
rect 16745 -1165 16750 -1145
rect 16750 -1165 16770 -1145
rect 16770 -1165 16775 -1145
rect 16745 -1170 16775 -1165
rect 16825 -1145 16855 -1140
rect 16825 -1165 16830 -1145
rect 16830 -1165 16850 -1145
rect 16850 -1165 16855 -1145
rect 16825 -1170 16855 -1165
rect 16905 -1145 16935 -1140
rect 16905 -1165 16910 -1145
rect 16910 -1165 16930 -1145
rect 16930 -1165 16935 -1145
rect 16905 -1170 16935 -1165
rect 16985 -1145 17015 -1140
rect 16985 -1165 16990 -1145
rect 16990 -1165 17010 -1145
rect 17010 -1165 17015 -1145
rect 16985 -1170 17015 -1165
rect 17065 -1145 17095 -1140
rect 17065 -1165 17070 -1145
rect 17070 -1165 17090 -1145
rect 17090 -1165 17095 -1145
rect 17065 -1170 17095 -1165
rect 17145 -1145 17175 -1140
rect 17145 -1165 17150 -1145
rect 17150 -1165 17170 -1145
rect 17170 -1165 17175 -1145
rect 17145 -1170 17175 -1165
rect 17225 -1145 17255 -1140
rect 17225 -1165 17230 -1145
rect 17230 -1165 17250 -1145
rect 17250 -1165 17255 -1145
rect 17225 -1170 17255 -1165
rect 17305 -1145 17335 -1140
rect 17305 -1165 17310 -1145
rect 17310 -1165 17330 -1145
rect 17330 -1165 17335 -1145
rect 17305 -1170 17335 -1165
rect 17385 -1145 17415 -1140
rect 17385 -1165 17390 -1145
rect 17390 -1165 17410 -1145
rect 17410 -1165 17415 -1145
rect 17385 -1170 17415 -1165
rect 17465 -1145 17495 -1140
rect 17465 -1165 17470 -1145
rect 17470 -1165 17490 -1145
rect 17490 -1165 17495 -1145
rect 17465 -1170 17495 -1165
rect 17545 -1145 17575 -1140
rect 17545 -1165 17550 -1145
rect 17550 -1165 17570 -1145
rect 17570 -1165 17575 -1145
rect 17545 -1170 17575 -1165
rect 17625 -1145 17655 -1140
rect 17625 -1165 17630 -1145
rect 17630 -1165 17650 -1145
rect 17650 -1165 17655 -1145
rect 17625 -1170 17655 -1165
rect 17705 -1145 17735 -1140
rect 17705 -1165 17710 -1145
rect 17710 -1165 17730 -1145
rect 17730 -1165 17735 -1145
rect 17705 -1170 17735 -1165
rect 17785 -1145 17815 -1140
rect 17785 -1165 17790 -1145
rect 17790 -1165 17810 -1145
rect 17810 -1165 17815 -1145
rect 17785 -1170 17815 -1165
rect 17865 -1145 17895 -1140
rect 17865 -1165 17870 -1145
rect 17870 -1165 17890 -1145
rect 17890 -1165 17895 -1145
rect 17865 -1170 17895 -1165
rect 17945 -1145 17975 -1140
rect 17945 -1165 17950 -1145
rect 17950 -1165 17970 -1145
rect 17970 -1165 17975 -1145
rect 17945 -1170 17975 -1165
rect 18025 -1145 18055 -1140
rect 18025 -1165 18030 -1145
rect 18030 -1165 18050 -1145
rect 18050 -1165 18055 -1145
rect 18025 -1170 18055 -1165
rect 18105 -1145 18135 -1140
rect 18105 -1165 18110 -1145
rect 18110 -1165 18130 -1145
rect 18130 -1165 18135 -1145
rect 18105 -1170 18135 -1165
rect 18185 -1145 18215 -1140
rect 18185 -1165 18190 -1145
rect 18190 -1165 18210 -1145
rect 18210 -1165 18215 -1145
rect 18185 -1170 18215 -1165
rect 18265 -1145 18295 -1140
rect 18265 -1165 18270 -1145
rect 18270 -1165 18290 -1145
rect 18290 -1165 18295 -1145
rect 18265 -1170 18295 -1165
rect 18345 -1145 18375 -1140
rect 18345 -1165 18350 -1145
rect 18350 -1165 18370 -1145
rect 18370 -1165 18375 -1145
rect 18345 -1170 18375 -1165
rect 18425 -1145 18455 -1140
rect 18425 -1165 18430 -1145
rect 18430 -1165 18450 -1145
rect 18450 -1165 18455 -1145
rect 18425 -1170 18455 -1165
rect 18505 -1145 18535 -1140
rect 18505 -1165 18510 -1145
rect 18510 -1165 18530 -1145
rect 18530 -1165 18535 -1145
rect 18505 -1170 18535 -1165
rect 18585 -1145 18615 -1140
rect 18585 -1165 18590 -1145
rect 18590 -1165 18610 -1145
rect 18610 -1165 18615 -1145
rect 18585 -1170 18615 -1165
rect 18665 -1145 18695 -1140
rect 18665 -1165 18670 -1145
rect 18670 -1165 18690 -1145
rect 18690 -1165 18695 -1145
rect 18665 -1170 18695 -1165
rect 18745 -1145 18775 -1140
rect 18745 -1165 18750 -1145
rect 18750 -1165 18770 -1145
rect 18770 -1165 18775 -1145
rect 18745 -1170 18775 -1165
rect 16705 -1230 16735 -1225
rect 16705 -1250 16710 -1230
rect 16710 -1250 16730 -1230
rect 16730 -1250 16735 -1230
rect 16705 -1255 16735 -1250
rect 18900 -1210 18930 -1205
rect 18900 -1230 18905 -1210
rect 18905 -1230 18925 -1210
rect 18925 -1230 18930 -1210
rect 18900 -1235 18930 -1230
rect 18900 -1250 18930 -1245
rect 18900 -1270 18905 -1250
rect 18905 -1270 18925 -1250
rect 18925 -1270 18930 -1250
rect 18900 -1275 18930 -1270
rect 16600 -1355 16630 -1325
rect 16710 -1355 16740 -1325
rect 17305 -1355 17335 -1325
rect 17785 -1355 17815 -1325
rect 18265 -1355 18295 -1325
rect 16545 -1440 16575 -1410
rect 16545 -1480 16575 -1450
rect 16655 -1440 16685 -1410
rect 16655 -1480 16685 -1450
rect 16545 -1495 16575 -1490
rect 16545 -1515 16550 -1495
rect 16550 -1515 16570 -1495
rect 16570 -1515 16575 -1495
rect 16545 -1520 16575 -1515
rect 16765 -1440 16795 -1410
rect 16765 -1480 16795 -1450
rect 16655 -1495 16685 -1490
rect 16655 -1515 16660 -1495
rect 16660 -1515 16680 -1495
rect 16680 -1515 16685 -1495
rect 16655 -1520 16685 -1515
rect 16765 -1495 16795 -1490
rect 16765 -1515 16770 -1495
rect 16770 -1515 16790 -1495
rect 16790 -1515 16795 -1495
rect 16765 -1520 16795 -1515
rect 16825 -1440 16855 -1410
rect 16825 -1480 16855 -1450
rect 16825 -1495 16855 -1490
rect 16825 -1515 16830 -1495
rect 16830 -1515 16850 -1495
rect 16850 -1515 16855 -1495
rect 16825 -1520 16855 -1515
rect 17030 -1440 17060 -1410
rect 17030 -1480 17060 -1450
rect 17030 -1495 17060 -1490
rect 17030 -1515 17035 -1495
rect 17035 -1515 17055 -1495
rect 17055 -1515 17060 -1495
rect 17030 -1520 17060 -1515
rect 17140 -1440 17170 -1410
rect 17140 -1480 17170 -1450
rect 17140 -1495 17170 -1490
rect 17140 -1515 17145 -1495
rect 17145 -1515 17165 -1495
rect 17165 -1515 17170 -1495
rect 17140 -1520 17170 -1515
rect 17250 -1440 17280 -1410
rect 17250 -1480 17280 -1450
rect 17360 -1440 17390 -1410
rect 17360 -1480 17390 -1450
rect 17250 -1495 17280 -1490
rect 17250 -1515 17255 -1495
rect 17255 -1515 17275 -1495
rect 17275 -1515 17280 -1495
rect 17250 -1520 17280 -1515
rect 17360 -1495 17390 -1490
rect 17360 -1515 17365 -1495
rect 17365 -1515 17385 -1495
rect 17385 -1515 17390 -1495
rect 17360 -1520 17390 -1515
rect 17470 -1440 17500 -1410
rect 17470 -1480 17500 -1450
rect 17470 -1495 17500 -1490
rect 17470 -1515 17475 -1495
rect 17475 -1515 17495 -1495
rect 17495 -1515 17500 -1495
rect 17470 -1520 17500 -1515
rect 17620 -1440 17650 -1410
rect 17620 -1480 17650 -1450
rect 17620 -1495 17650 -1490
rect 17620 -1515 17625 -1495
rect 17625 -1515 17645 -1495
rect 17645 -1515 17650 -1495
rect 17620 -1520 17650 -1515
rect 17730 -1440 17760 -1410
rect 17730 -1480 17760 -1450
rect 17840 -1440 17870 -1410
rect 17840 -1480 17870 -1450
rect 17730 -1495 17760 -1490
rect 17730 -1515 17735 -1495
rect 17735 -1515 17755 -1495
rect 17755 -1515 17760 -1495
rect 17730 -1520 17760 -1515
rect 17840 -1495 17870 -1490
rect 17840 -1515 17845 -1495
rect 17845 -1515 17865 -1495
rect 17865 -1515 17870 -1495
rect 17840 -1520 17870 -1515
rect 17950 -1440 17980 -1410
rect 17950 -1480 17980 -1450
rect 17950 -1495 17980 -1490
rect 17950 -1515 17955 -1495
rect 17955 -1515 17975 -1495
rect 17975 -1515 17980 -1495
rect 17950 -1520 17980 -1515
rect 18100 -1440 18130 -1410
rect 18100 -1480 18130 -1450
rect 18100 -1495 18130 -1490
rect 18100 -1515 18105 -1495
rect 18105 -1515 18125 -1495
rect 18125 -1515 18130 -1495
rect 18100 -1520 18130 -1515
rect 18210 -1440 18240 -1410
rect 18210 -1480 18240 -1450
rect 18320 -1440 18350 -1410
rect 18320 -1480 18350 -1450
rect 18210 -1495 18240 -1490
rect 18210 -1515 18215 -1495
rect 18215 -1515 18235 -1495
rect 18235 -1515 18240 -1495
rect 18210 -1520 18240 -1515
rect 18320 -1495 18350 -1490
rect 18320 -1515 18325 -1495
rect 18325 -1515 18345 -1495
rect 18345 -1515 18350 -1495
rect 18320 -1520 18350 -1515
rect 18430 -1440 18460 -1410
rect 18430 -1480 18460 -1450
rect 18430 -1495 18460 -1490
rect 18430 -1515 18435 -1495
rect 18435 -1515 18455 -1495
rect 18455 -1515 18460 -1495
rect 18430 -1520 18460 -1515
rect 18540 -1440 18570 -1410
rect 18540 -1480 18570 -1450
rect 18540 -1495 18570 -1490
rect 18540 -1515 18545 -1495
rect 18545 -1515 18565 -1495
rect 18565 -1515 18570 -1495
rect 18540 -1520 18570 -1515
rect 17195 -1665 17225 -1660
rect 17195 -1685 17200 -1665
rect 17200 -1685 17220 -1665
rect 17220 -1685 17225 -1665
rect 17195 -1690 17225 -1685
rect 17085 -1745 17115 -1715
rect 17415 -1665 17445 -1660
rect 17415 -1685 17420 -1665
rect 17420 -1685 17440 -1665
rect 17440 -1685 17445 -1665
rect 17415 -1690 17445 -1685
rect 17675 -1665 17705 -1660
rect 17675 -1685 17680 -1665
rect 17680 -1685 17700 -1665
rect 17700 -1685 17705 -1665
rect 17675 -1690 17705 -1685
rect 17785 -1665 17815 -1660
rect 17785 -1685 17790 -1665
rect 17790 -1685 17810 -1665
rect 17810 -1685 17815 -1665
rect 17785 -1690 17815 -1685
rect 17895 -1665 17925 -1660
rect 17895 -1685 17900 -1665
rect 17900 -1685 17920 -1665
rect 17920 -1685 17925 -1665
rect 17895 -1690 17925 -1685
rect 18155 -1665 18185 -1660
rect 18155 -1685 18160 -1665
rect 18160 -1685 18180 -1665
rect 18180 -1685 18185 -1665
rect 18155 -1690 18185 -1685
rect 18375 -1665 18405 -1660
rect 18375 -1685 18380 -1665
rect 18380 -1685 18400 -1665
rect 18400 -1685 18405 -1665
rect 18375 -1690 18405 -1685
rect 17305 -1745 17335 -1715
rect 17195 -1800 17225 -1770
rect 17195 -1840 17225 -1810
rect 18265 -1745 18295 -1715
rect 18485 -1745 18515 -1715
rect 18375 -1800 18405 -1770
rect 18375 -1840 18405 -1810
rect 16710 -1930 16740 -1900
rect 17785 -1930 17815 -1900
rect 19330 -1980 19360 -1950
rect 16265 -2030 16295 -2000
rect 16485 -2030 16515 -2000
rect 16735 -2030 16765 -2000
rect 17200 -2030 17230 -2000
rect 16485 -2905 16520 -2900
rect 16485 -2930 16490 -2905
rect 16490 -2930 16515 -2905
rect 16515 -2930 16520 -2905
rect 16485 -2935 16520 -2930
rect 16160 -3030 16195 -3025
rect 16160 -3055 16165 -3030
rect 16165 -3055 16190 -3030
rect 16190 -3055 16195 -3030
rect 16160 -3060 16195 -3055
rect 17430 -2005 17465 -2000
rect 17430 -2030 17435 -2005
rect 17435 -2030 17460 -2005
rect 17460 -2030 17465 -2005
rect 17430 -2035 17465 -2030
rect 18129 -2005 18164 -2000
rect 18129 -2030 18134 -2005
rect 18134 -2030 18159 -2005
rect 18159 -2030 18164 -2005
rect 18129 -2035 18164 -2030
rect 19085 -2035 19115 -2005
rect 17200 -2090 17230 -2060
rect 18835 -2090 18865 -2060
rect 15825 -3145 15855 -3115
rect 15950 -3121 15985 -3116
rect 15950 -3146 15955 -3121
rect 15955 -3146 15980 -3121
rect 15980 -3146 15985 -3121
rect 16735 -3135 16765 -3105
rect 15950 -3151 15985 -3146
rect 17785 -3135 17815 -3105
rect 19080 -2905 19115 -2900
rect 19080 -2930 19085 -2905
rect 19085 -2930 19110 -2905
rect 19110 -2930 19115 -2905
rect 19080 -2935 19115 -2930
rect 19615 380 19645 410
rect 19540 -1930 19570 -1900
rect 19465 -2035 19495 -2005
rect 19405 -3002 19440 -2997
rect 19405 -3027 19410 -3002
rect 19410 -3027 19435 -3002
rect 19435 -3027 19440 -3002
rect 19405 -3032 19440 -3027
rect 18620 -3135 18650 -3105
rect 18835 -3135 18865 -3105
rect 19725 -125 19755 -95
rect 19610 -3121 19645 -3116
rect 19610 -3146 19615 -3121
rect 19615 -3146 19640 -3121
rect 19640 -3146 19645 -3121
rect 19610 -3151 19645 -3146
rect 15950 -3794 15985 -3789
rect 15950 -3819 15955 -3794
rect 15955 -3819 15980 -3794
rect 15980 -3819 15985 -3794
rect 15950 -3824 15985 -3819
rect 15825 -4295 15855 -4265
rect 15730 -4345 15760 -4315
rect 16280 -3899 16315 -3894
rect 16280 -3924 16285 -3899
rect 16285 -3924 16310 -3899
rect 16310 -3924 16315 -3899
rect 16280 -3929 16315 -3924
rect 16605 -3974 16640 -3969
rect 16605 -3999 16610 -3974
rect 16610 -3999 16635 -3974
rect 16635 -3999 16640 -3974
rect 19610 -3794 19645 -3789
rect 19610 -3819 19615 -3794
rect 19615 -3819 19640 -3794
rect 19640 -3819 19645 -3794
rect 19610 -3824 19645 -3819
rect 19285 -3899 19320 -3894
rect 19285 -3924 19290 -3899
rect 19290 -3924 19315 -3899
rect 19315 -3924 19320 -3899
rect 19285 -3929 19320 -3924
rect 18960 -3974 18995 -3969
rect 16605 -4004 16640 -3999
rect 18960 -3999 18965 -3974
rect 18965 -3999 18990 -3974
rect 18990 -3999 18995 -3974
rect 18960 -4004 18995 -3999
rect 16285 -4220 16315 -4190
rect 16610 -4220 16640 -4190
rect 17260 -4295 17290 -4265
rect 17785 -4270 17815 -4265
rect 17785 -4290 17790 -4270
rect 17790 -4290 17810 -4270
rect 17810 -4290 17815 -4270
rect 17785 -4295 17815 -4290
rect 18960 -4295 18990 -4265
rect 19285 -4295 19315 -4265
rect 16910 -4345 16940 -4315
rect 18660 -4345 18690 -4315
rect 19780 -1800 19810 -1770
rect 19780 -1840 19810 -1810
rect 19725 -4345 19755 -4315
rect 15955 -4390 15985 -4360
rect 16210 -4390 16240 -4360
rect 19360 -4390 19390 -4360
rect 19615 -4390 19645 -4360
rect 17960 -4440 17990 -4410
<< metal2 >>
rect 16940 1665 16980 1670
rect 16940 1635 16945 1665
rect 16975 1635 16980 1665
rect 16940 1630 16980 1635
rect 18620 1665 18660 1670
rect 18620 1635 18625 1665
rect 18655 1635 18660 1665
rect 18620 1630 18660 1635
rect 16485 1620 16525 1625
rect 16485 1590 16490 1620
rect 16520 1615 16525 1620
rect 17050 1620 17090 1625
rect 17050 1615 17055 1620
rect 16520 1595 17055 1615
rect 16520 1590 16525 1595
rect 16485 1585 16525 1590
rect 17050 1590 17055 1595
rect 17085 1615 17090 1620
rect 17780 1620 17820 1625
rect 17780 1615 17785 1620
rect 17085 1595 17785 1615
rect 17085 1590 17090 1595
rect 17050 1585 17090 1590
rect 17780 1590 17785 1595
rect 17815 1615 17820 1620
rect 18200 1620 18240 1625
rect 18200 1615 18205 1620
rect 17815 1595 18205 1615
rect 17815 1590 17820 1595
rect 17780 1585 17820 1590
rect 18200 1590 18205 1595
rect 18235 1615 18240 1620
rect 18510 1620 18550 1625
rect 18510 1615 18515 1620
rect 18235 1595 18515 1615
rect 18235 1590 18240 1595
rect 18200 1585 18240 1590
rect 18510 1590 18515 1595
rect 18545 1590 18550 1620
rect 18510 1585 18550 1590
rect 16365 1520 18715 1525
rect 16365 1490 16370 1520
rect 16400 1490 16490 1520
rect 16520 1490 16610 1520
rect 16640 1490 16890 1520
rect 16920 1490 17000 1520
rect 17030 1490 17110 1520
rect 17140 1490 17220 1520
rect 17250 1490 17500 1520
rect 17530 1490 17565 1520
rect 17595 1490 17675 1520
rect 17705 1490 17785 1520
rect 17815 1490 17895 1520
rect 17925 1490 18005 1520
rect 18035 1490 18070 1520
rect 18100 1490 18350 1520
rect 18380 1490 18460 1520
rect 18490 1490 18570 1520
rect 18600 1490 18680 1520
rect 18710 1490 18715 1520
rect 16365 1480 18715 1490
rect 16365 1450 16370 1480
rect 16400 1450 16490 1480
rect 16520 1450 16610 1480
rect 16640 1450 16890 1480
rect 16920 1450 17000 1480
rect 17030 1450 17110 1480
rect 17140 1450 17220 1480
rect 17250 1450 17500 1480
rect 17530 1450 17565 1480
rect 17595 1450 17675 1480
rect 17705 1450 17785 1480
rect 17815 1450 17895 1480
rect 17925 1450 18005 1480
rect 18035 1450 18070 1480
rect 18100 1450 18350 1480
rect 18380 1450 18460 1480
rect 18490 1450 18570 1480
rect 18600 1450 18680 1480
rect 18710 1450 18715 1480
rect 16365 1440 18715 1450
rect 16365 1410 16370 1440
rect 16400 1410 16490 1440
rect 16520 1410 16610 1440
rect 16640 1410 16890 1440
rect 16920 1410 17000 1440
rect 17030 1410 17110 1440
rect 17140 1410 17220 1440
rect 17250 1410 17500 1440
rect 17530 1410 17565 1440
rect 17595 1410 17675 1440
rect 17705 1410 17785 1440
rect 17815 1410 17895 1440
rect 17925 1410 18005 1440
rect 18035 1410 18070 1440
rect 18100 1410 18350 1440
rect 18380 1410 18460 1440
rect 18490 1410 18570 1440
rect 18600 1410 18680 1440
rect 18710 1410 18715 1440
rect 16365 1405 18715 1410
rect 16430 1270 16470 1275
rect 16430 1240 16435 1270
rect 16465 1240 16470 1270
rect 16430 1235 16470 1240
rect 16540 1270 16580 1275
rect 16540 1240 16545 1270
rect 16575 1240 16580 1270
rect 16540 1235 16580 1240
rect 16940 1270 16980 1275
rect 16940 1240 16945 1270
rect 16975 1265 16980 1270
rect 17050 1270 17090 1275
rect 17050 1265 17055 1270
rect 16975 1245 17055 1265
rect 16975 1240 16980 1245
rect 16940 1235 16980 1240
rect 17050 1240 17055 1245
rect 17085 1265 17090 1270
rect 17160 1270 17200 1275
rect 17160 1265 17165 1270
rect 17085 1245 17165 1265
rect 17085 1240 17090 1245
rect 17050 1235 17090 1240
rect 17160 1240 17165 1245
rect 17195 1240 17200 1270
rect 17160 1235 17200 1240
rect 17615 1270 17655 1275
rect 17615 1240 17620 1270
rect 17650 1265 17655 1270
rect 17725 1270 17765 1275
rect 17725 1265 17730 1270
rect 17650 1245 17730 1265
rect 17650 1240 17655 1245
rect 17615 1235 17655 1240
rect 17725 1240 17730 1245
rect 17760 1265 17765 1270
rect 17835 1270 17875 1275
rect 17835 1265 17840 1270
rect 17760 1245 17840 1265
rect 17760 1240 17765 1245
rect 17725 1235 17765 1240
rect 17835 1240 17840 1245
rect 17870 1265 17875 1270
rect 17945 1270 17985 1275
rect 17945 1265 17950 1270
rect 17870 1245 17950 1265
rect 17870 1240 17875 1245
rect 17835 1235 17875 1240
rect 17945 1240 17950 1245
rect 17980 1240 17985 1270
rect 17945 1235 17985 1240
rect 18400 1270 18440 1275
rect 18400 1240 18405 1270
rect 18435 1265 18440 1270
rect 18510 1270 18550 1275
rect 18510 1265 18515 1270
rect 18435 1245 18515 1265
rect 18435 1240 18440 1245
rect 18400 1235 18440 1240
rect 18510 1240 18515 1245
rect 18545 1265 18550 1270
rect 18620 1270 18660 1275
rect 18620 1265 18625 1270
rect 18545 1245 18625 1265
rect 18545 1240 18550 1245
rect 18510 1235 18550 1240
rect 18620 1240 18625 1245
rect 18655 1240 18660 1270
rect 18620 1235 18660 1240
rect 18200 1215 18240 1220
rect 18200 1185 18205 1215
rect 18235 1210 18240 1215
rect 18720 1215 18760 1220
rect 18720 1210 18725 1215
rect 18235 1190 18725 1210
rect 18235 1185 18240 1190
rect 18200 1180 18240 1185
rect 18720 1185 18725 1190
rect 18755 1185 18760 1215
rect 18720 1180 18760 1185
rect 16160 1170 16200 1175
rect 16160 1140 16165 1170
rect 16195 1165 16200 1170
rect 16430 1170 16470 1175
rect 16430 1165 16435 1170
rect 16195 1145 16435 1165
rect 16195 1140 16200 1145
rect 16160 1135 16200 1140
rect 16430 1140 16435 1145
rect 16465 1140 16470 1170
rect 16430 1135 16470 1140
rect 16540 1170 16580 1175
rect 16540 1140 16545 1170
rect 16575 1165 16580 1170
rect 19325 1170 19365 1175
rect 19325 1165 19330 1170
rect 16575 1145 19330 1165
rect 16575 1140 16580 1145
rect 16540 1135 16580 1140
rect 19325 1140 19330 1145
rect 19360 1140 19365 1170
rect 19325 1135 19365 1140
rect 16435 1055 19115 1060
rect 16435 1025 16440 1055
rect 16470 1025 16660 1055
rect 16690 1025 16975 1055
rect 17005 1025 17155 1055
rect 17185 1025 17335 1055
rect 17365 1025 17515 1055
rect 17545 1025 17695 1055
rect 17725 1025 17875 1055
rect 17905 1025 18055 1055
rect 18085 1025 18235 1055
rect 18265 1025 18415 1055
rect 18445 1025 18595 1055
rect 18625 1025 18910 1055
rect 18940 1025 19020 1055
rect 19050 1025 19080 1055
rect 19110 1025 19115 1055
rect 16435 1015 19115 1025
rect 16435 985 16440 1015
rect 16470 985 16660 1015
rect 16690 985 16975 1015
rect 17005 985 17155 1015
rect 17185 985 17335 1015
rect 17365 985 17515 1015
rect 17545 985 17695 1015
rect 17725 985 17875 1015
rect 17905 985 18055 1015
rect 18085 985 18235 1015
rect 18265 985 18415 1015
rect 18445 985 18595 1015
rect 18625 985 18910 1015
rect 18940 985 19020 1015
rect 19050 985 19080 1015
rect 19110 985 19115 1015
rect 16435 975 19115 985
rect 16435 945 16440 975
rect 16470 945 16660 975
rect 16690 945 16975 975
rect 17005 945 17155 975
rect 17185 945 17335 975
rect 17365 945 17515 975
rect 17545 945 17695 975
rect 17725 945 17875 975
rect 17905 945 18055 975
rect 18085 945 18235 975
rect 18265 945 18415 975
rect 18445 945 18595 975
rect 18625 945 18910 975
rect 18940 945 19020 975
rect 19050 945 19080 975
rect 19110 945 19115 975
rect 16435 940 19115 945
rect 16545 875 16585 880
rect 16545 845 16550 875
rect 16580 870 16585 875
rect 16780 875 16820 880
rect 16780 870 16785 875
rect 16580 850 16785 870
rect 16580 845 16585 850
rect 16545 840 16585 845
rect 16780 845 16785 850
rect 16815 845 16820 875
rect 16780 840 16820 845
rect 16480 705 16520 710
rect 16480 675 16485 705
rect 16515 700 16520 705
rect 16610 705 16650 710
rect 16610 700 16615 705
rect 16515 680 16615 700
rect 16515 675 16520 680
rect 16480 670 16520 675
rect 16610 675 16615 680
rect 16645 700 16650 705
rect 16840 705 16880 710
rect 16840 700 16845 705
rect 16645 680 16845 700
rect 16645 675 16650 680
rect 16610 670 16650 675
rect 16840 675 16845 680
rect 16875 675 16880 705
rect 16840 670 16880 675
rect 18950 705 18990 710
rect 18950 675 18955 705
rect 18985 700 18990 705
rect 19260 705 19300 710
rect 19260 700 19265 705
rect 18985 680 19265 700
rect 18985 675 18990 680
rect 18950 670 18990 675
rect 19260 675 19265 680
rect 19295 675 19300 705
rect 19260 670 19300 675
rect 19000 625 19005 655
rect 19035 625 19040 655
rect 16315 605 19500 610
rect 16315 575 16320 605
rect 16350 575 17605 605
rect 17635 575 17965 605
rect 17995 575 19465 605
rect 19495 575 19500 605
rect 16315 570 19500 575
rect 16260 550 16300 555
rect 16260 520 16265 550
rect 16295 545 16300 550
rect 16780 550 16820 555
rect 16780 545 16785 550
rect 16295 525 16785 545
rect 16295 520 16300 525
rect 16260 515 16300 520
rect 16780 520 16785 525
rect 16815 545 16820 550
rect 17420 550 17460 555
rect 17420 545 17425 550
rect 16815 525 17425 545
rect 16815 520 16820 525
rect 16780 515 16820 520
rect 17420 520 17425 525
rect 17455 545 17460 550
rect 18140 550 18180 555
rect 18140 545 18145 550
rect 17455 525 18145 545
rect 17455 520 17460 525
rect 17420 515 17460 520
rect 18140 520 18145 525
rect 18175 520 18180 550
rect 18140 515 18180 520
rect 16205 505 16245 510
rect 16205 475 16210 505
rect 16240 500 16245 505
rect 16545 505 16585 510
rect 16545 500 16550 505
rect 16240 480 16550 500
rect 16240 475 16245 480
rect 16205 470 16245 475
rect 16545 475 16550 480
rect 16580 500 16585 505
rect 17240 505 17280 510
rect 17240 500 17245 505
rect 16580 480 17245 500
rect 16580 475 16585 480
rect 16545 470 16585 475
rect 17240 475 17245 480
rect 17275 500 17280 505
rect 18320 505 18360 510
rect 18320 500 18325 505
rect 17275 480 18325 500
rect 17275 475 17280 480
rect 17240 470 17280 475
rect 18320 475 18325 480
rect 18355 475 18360 505
rect 18320 470 18360 475
rect 17060 460 17100 465
rect 17060 430 17065 460
rect 17095 455 17100 460
rect 17780 460 17820 465
rect 17780 455 17785 460
rect 17095 435 17785 455
rect 17095 430 17100 435
rect 17060 425 17100 430
rect 17780 430 17785 435
rect 17815 455 17820 460
rect 18500 460 18540 465
rect 18500 455 18505 460
rect 17815 435 18505 455
rect 17815 430 17820 435
rect 17780 425 17820 430
rect 18500 430 18505 435
rect 18535 455 18540 460
rect 19405 460 19445 465
rect 19405 455 19410 460
rect 18535 435 19410 455
rect 18535 430 18540 435
rect 18500 425 18540 430
rect 19405 430 19410 435
rect 19440 430 19445 460
rect 19405 425 19445 430
rect 18000 410 18040 415
rect 18000 380 18005 410
rect 18035 405 18040 410
rect 18720 410 18760 415
rect 18720 405 18725 410
rect 18035 385 18725 405
rect 18035 380 18040 385
rect 18000 375 18040 380
rect 18720 380 18725 385
rect 18755 405 18760 410
rect 19010 410 19050 415
rect 19010 405 19015 410
rect 18755 385 19015 405
rect 18755 380 18760 385
rect 18720 375 18760 380
rect 19010 380 19015 385
rect 19045 405 19050 410
rect 19610 410 19650 415
rect 19610 405 19615 410
rect 19045 385 19615 405
rect 19045 380 19050 385
rect 19010 375 19050 380
rect 19610 380 19615 385
rect 19645 380 19650 410
rect 19610 375 19650 380
rect 16420 270 19180 275
rect 16420 240 16425 270
rect 16455 240 16545 270
rect 16575 240 16665 270
rect 16695 240 16785 270
rect 16815 240 16905 270
rect 16935 240 17025 270
rect 17055 240 17145 270
rect 17175 240 17265 270
rect 17295 240 17385 270
rect 17415 240 17505 270
rect 17535 240 17625 270
rect 17655 240 17945 270
rect 17975 240 18065 270
rect 18095 240 18185 270
rect 18215 240 18305 270
rect 18335 240 18425 270
rect 18455 240 18545 270
rect 18575 240 18665 270
rect 18695 240 18785 270
rect 18815 240 18905 270
rect 18935 240 19025 270
rect 19055 240 19145 270
rect 19175 240 19180 270
rect 16420 230 19180 240
rect 16420 200 16425 230
rect 16455 200 16545 230
rect 16575 200 16665 230
rect 16695 200 16785 230
rect 16815 200 16905 230
rect 16935 200 17025 230
rect 17055 200 17145 230
rect 17175 200 17265 230
rect 17295 200 17385 230
rect 17415 200 17505 230
rect 17535 200 17625 230
rect 17655 200 17945 230
rect 17975 200 18065 230
rect 18095 200 18185 230
rect 18215 200 18305 230
rect 18335 200 18425 230
rect 18455 200 18545 230
rect 18575 200 18665 230
rect 18695 200 18785 230
rect 18815 200 18905 230
rect 18935 200 19025 230
rect 19055 200 19145 230
rect 19175 200 19180 230
rect 16420 190 19180 200
rect 16420 160 16425 190
rect 16455 160 16545 190
rect 16575 160 16665 190
rect 16695 160 16785 190
rect 16815 160 16905 190
rect 16935 160 17025 190
rect 17055 160 17145 190
rect 17175 160 17265 190
rect 17295 160 17385 190
rect 17415 160 17505 190
rect 17535 160 17625 190
rect 17655 160 17945 190
rect 17975 160 18065 190
rect 18095 160 18185 190
rect 18215 160 18305 190
rect 18335 160 18425 190
rect 18455 160 18545 190
rect 18575 160 18665 190
rect 18695 160 18785 190
rect 18815 160 18905 190
rect 18935 160 19025 190
rect 19055 160 19145 190
rect 19175 160 19180 190
rect 16420 155 19180 160
rect 15950 135 15990 140
rect 15950 105 15955 135
rect 15985 130 15990 135
rect 16480 135 16520 140
rect 16480 130 16485 135
rect 15985 110 16485 130
rect 15985 105 15990 110
rect 15950 100 15990 105
rect 16480 105 16485 110
rect 16515 130 16520 135
rect 16840 135 16880 140
rect 16840 130 16845 135
rect 16515 110 16845 130
rect 16515 105 16520 110
rect 16480 100 16520 105
rect 16840 105 16845 110
rect 16875 130 16880 135
rect 17200 135 17240 140
rect 17200 130 17205 135
rect 16875 110 17205 130
rect 16875 105 16880 110
rect 16840 100 16880 105
rect 17200 105 17205 110
rect 17235 130 17240 135
rect 17560 135 17600 140
rect 17560 130 17565 135
rect 17235 110 17565 130
rect 17235 105 17240 110
rect 17200 100 17240 105
rect 17560 105 17565 110
rect 17595 130 17600 135
rect 17690 135 17730 140
rect 17690 130 17695 135
rect 17595 110 17695 130
rect 17595 105 17600 110
rect 17560 100 17600 105
rect 17690 105 17695 110
rect 17725 105 17730 135
rect 17690 100 17730 105
rect 17870 135 17910 140
rect 17870 105 17875 135
rect 17905 130 17910 135
rect 18000 135 18040 140
rect 18000 130 18005 135
rect 17905 110 18005 130
rect 17905 105 17910 110
rect 17870 100 17910 105
rect 18000 105 18005 110
rect 18035 130 18040 135
rect 18360 135 18400 140
rect 18360 130 18365 135
rect 18035 110 18365 130
rect 18035 105 18040 110
rect 18000 100 18040 105
rect 18360 105 18365 110
rect 18395 130 18400 135
rect 18720 135 18760 140
rect 18720 130 18725 135
rect 18395 110 18725 130
rect 18395 105 18400 110
rect 18360 100 18400 105
rect 18720 105 18725 110
rect 18755 130 18760 135
rect 19080 135 19120 140
rect 19080 130 19085 135
rect 18755 110 19085 130
rect 18755 105 18760 110
rect 18720 100 18760 105
rect 19080 105 19085 110
rect 19115 105 19120 135
rect 19080 100 19120 105
rect 16600 -35 16640 -30
rect 16600 -65 16605 -35
rect 16635 -40 16640 -35
rect 16960 -35 17000 -30
rect 16960 -40 16965 -35
rect 16635 -60 16965 -40
rect 16635 -65 16640 -60
rect 16600 -70 16640 -65
rect 16960 -65 16965 -60
rect 16995 -40 17000 -35
rect 17320 -35 17360 -30
rect 17320 -40 17325 -35
rect 16995 -60 17325 -40
rect 16995 -65 17000 -60
rect 16960 -70 17000 -65
rect 17320 -65 17325 -60
rect 17355 -65 17360 -35
rect 17320 -70 17360 -65
rect 18240 -35 18280 -30
rect 18240 -65 18245 -35
rect 18275 -40 18280 -35
rect 18600 -35 18640 -30
rect 18600 -40 18605 -35
rect 18275 -60 18605 -40
rect 18275 -65 18280 -60
rect 18240 -70 18280 -65
rect 18600 -65 18605 -60
rect 18635 -40 18640 -35
rect 18960 -35 19000 -30
rect 18960 -40 18965 -35
rect 18635 -60 18965 -40
rect 18635 -65 18640 -60
rect 18600 -70 18640 -65
rect 18960 -65 18965 -60
rect 18995 -65 19000 -35
rect 18960 -70 19000 -65
rect 15725 -95 15765 -90
rect 15725 -125 15730 -95
rect 15760 -100 15765 -95
rect 16510 -95 16550 -90
rect 16510 -100 16515 -95
rect 15760 -120 16515 -100
rect 15760 -125 15765 -120
rect 15725 -130 15765 -125
rect 16510 -125 16515 -120
rect 16545 -100 16550 -95
rect 16720 -95 16760 -90
rect 16720 -100 16725 -95
rect 16545 -120 16725 -100
rect 16545 -125 16550 -120
rect 16510 -130 16550 -125
rect 16720 -125 16725 -120
rect 16755 -100 16760 -95
rect 16840 -95 16880 -90
rect 16840 -100 16845 -95
rect 16755 -120 16845 -100
rect 16755 -125 16760 -120
rect 16720 -130 16760 -125
rect 16840 -125 16845 -120
rect 16875 -100 16880 -95
rect 17080 -95 17120 -90
rect 17080 -100 17085 -95
rect 16875 -120 17085 -100
rect 16875 -125 16880 -120
rect 16840 -130 16880 -125
rect 17080 -125 17085 -120
rect 17115 -100 17120 -95
rect 17200 -95 17240 -90
rect 17200 -100 17205 -95
rect 17115 -120 17205 -100
rect 17115 -125 17120 -120
rect 17080 -130 17120 -125
rect 17200 -125 17205 -120
rect 17235 -100 17240 -95
rect 17440 -95 17480 -90
rect 17440 -100 17445 -95
rect 17235 -120 17445 -100
rect 17235 -125 17240 -120
rect 17200 -130 17240 -125
rect 17440 -125 17445 -120
rect 17475 -100 17480 -95
rect 17530 -95 17570 -90
rect 17530 -100 17535 -95
rect 17475 -120 17535 -100
rect 17475 -125 17480 -120
rect 17440 -130 17480 -125
rect 17530 -125 17535 -120
rect 17565 -125 17570 -95
rect 17530 -130 17570 -125
rect 18030 -95 18070 -90
rect 18030 -125 18035 -95
rect 18065 -100 18070 -95
rect 18120 -95 18160 -90
rect 18120 -100 18125 -95
rect 18065 -120 18125 -100
rect 18065 -125 18070 -120
rect 18030 -130 18070 -125
rect 18120 -125 18125 -120
rect 18155 -100 18160 -95
rect 18360 -95 18400 -90
rect 18360 -100 18365 -95
rect 18155 -120 18365 -100
rect 18155 -125 18160 -120
rect 18120 -130 18160 -125
rect 18360 -125 18365 -120
rect 18395 -100 18400 -95
rect 18480 -95 18520 -90
rect 18480 -100 18485 -95
rect 18395 -120 18485 -100
rect 18395 -125 18400 -120
rect 18360 -130 18400 -125
rect 18480 -125 18485 -120
rect 18515 -100 18520 -95
rect 18720 -95 18760 -90
rect 18720 -100 18725 -95
rect 18515 -120 18725 -100
rect 18515 -125 18520 -120
rect 18480 -130 18520 -125
rect 18720 -125 18725 -120
rect 18755 -100 18760 -95
rect 18840 -95 18880 -90
rect 18840 -100 18845 -95
rect 18755 -120 18845 -100
rect 18755 -125 18760 -120
rect 18720 -130 18760 -125
rect 18840 -125 18845 -120
rect 18875 -100 18880 -95
rect 19050 -95 19090 -90
rect 19050 -100 19055 -95
rect 18875 -120 19055 -100
rect 18875 -125 18880 -120
rect 18840 -130 18880 -125
rect 19050 -125 19055 -120
rect 19085 -100 19090 -95
rect 19720 -95 19760 -90
rect 19720 -100 19725 -95
rect 19085 -120 19725 -100
rect 19085 -125 19090 -120
rect 19050 -130 19090 -125
rect 19720 -125 19725 -120
rect 19755 -125 19760 -95
rect 19720 -130 19760 -125
rect 16260 -150 16300 -145
rect 16260 -180 16265 -150
rect 16295 -155 16300 -150
rect 17007 -150 17037 -145
rect 16295 -175 17007 -155
rect 16295 -180 16300 -175
rect 16260 -185 16300 -180
rect 18563 -150 18593 -145
rect 18562 -175 18563 -155
rect 17007 -185 17037 -180
rect 19405 -150 19445 -145
rect 19405 -155 19410 -150
rect 18593 -175 19410 -155
rect 18563 -185 18593 -180
rect 19405 -180 19410 -175
rect 19440 -180 19445 -150
rect 19405 -185 19445 -180
rect 17560 -210 18040 -205
rect 17560 -240 17565 -210
rect 17595 -240 17745 -210
rect 17775 -240 17785 -210
rect 17815 -240 17825 -210
rect 17855 -240 18005 -210
rect 18035 -240 18040 -210
rect 17560 -250 18040 -240
rect 17560 -280 17565 -250
rect 17595 -280 17745 -250
rect 17775 -280 17785 -250
rect 17815 -280 17825 -250
rect 17855 -280 18005 -250
rect 18035 -280 18040 -250
rect 17560 -290 18040 -280
rect 17560 -320 17565 -290
rect 17595 -320 17745 -290
rect 17775 -320 17785 -290
rect 17815 -320 17825 -290
rect 17855 -320 18005 -290
rect 18035 -320 18040 -290
rect 17560 -325 18040 -320
rect 16315 -470 17105 -465
rect 16315 -500 16320 -470
rect 16350 -500 17075 -470
rect 16315 -505 17105 -500
rect 18495 -470 18525 -465
rect 19325 -470 19365 -465
rect 19325 -475 19330 -470
rect 18525 -495 19330 -475
rect 18495 -505 18525 -500
rect 19325 -500 19330 -495
rect 19360 -500 19365 -470
rect 19325 -505 19365 -500
rect 16530 -550 17060 -545
rect 16530 -580 16535 -550
rect 16565 -580 17025 -550
rect 17055 -580 17060 -550
rect 16530 -585 17060 -580
rect 18540 -550 18580 -545
rect 18540 -580 18545 -550
rect 18575 -555 18580 -550
rect 19030 -550 19070 -545
rect 19030 -555 19035 -550
rect 18575 -575 19035 -555
rect 18575 -580 18580 -575
rect 18540 -585 18580 -580
rect 19030 -580 19035 -575
rect 19065 -580 19070 -550
rect 19030 -585 19070 -580
rect 16620 -605 18980 -600
rect 16620 -635 16625 -605
rect 16655 -635 16745 -605
rect 16775 -635 16865 -605
rect 16895 -635 16985 -605
rect 17015 -635 17305 -605
rect 17335 -635 17425 -605
rect 17455 -635 17545 -605
rect 17575 -635 18025 -605
rect 18055 -635 18145 -605
rect 18175 -635 18265 -605
rect 18295 -635 18585 -605
rect 18615 -635 18705 -605
rect 18735 -635 18825 -605
rect 18855 -635 18945 -605
rect 18975 -635 18980 -605
rect 16620 -645 18980 -635
rect 16620 -675 16625 -645
rect 16655 -675 16745 -645
rect 16775 -675 16865 -645
rect 16895 -675 16985 -645
rect 17015 -675 17305 -645
rect 17335 -675 17425 -645
rect 17455 -675 17545 -645
rect 17575 -675 18025 -645
rect 18055 -675 18145 -645
rect 18175 -675 18265 -645
rect 18295 -675 18585 -645
rect 18615 -675 18705 -645
rect 18735 -675 18825 -645
rect 18855 -675 18945 -645
rect 18975 -675 18980 -645
rect 16620 -685 18980 -675
rect 16620 -715 16625 -685
rect 16655 -715 16745 -685
rect 16775 -715 16865 -685
rect 16895 -715 16985 -685
rect 17015 -715 17305 -685
rect 17335 -715 17425 -685
rect 17455 -715 17545 -685
rect 17575 -715 18025 -685
rect 18055 -715 18145 -685
rect 18175 -715 18265 -685
rect 18295 -715 18585 -685
rect 18615 -715 18705 -685
rect 18735 -715 18825 -685
rect 18855 -715 18945 -685
rect 18975 -715 18980 -685
rect 16620 -720 18980 -715
rect 17110 -1005 18490 -1000
rect 17110 -1035 17115 -1005
rect 17145 -1035 17745 -1005
rect 17775 -1035 17785 -1005
rect 17815 -1035 17825 -1005
rect 17855 -1035 18455 -1005
rect 18485 -1035 18490 -1005
rect 17110 -1045 18490 -1035
rect 17110 -1075 17115 -1045
rect 17145 -1075 17745 -1045
rect 17775 -1075 17785 -1045
rect 17815 -1075 17825 -1045
rect 17855 -1075 18455 -1045
rect 18485 -1075 18490 -1045
rect 17110 -1085 18490 -1075
rect 17110 -1115 17115 -1085
rect 17145 -1115 17745 -1085
rect 17775 -1115 17785 -1085
rect 17815 -1115 17825 -1085
rect 17855 -1115 18455 -1085
rect 18485 -1115 18490 -1085
rect 17110 -1120 18490 -1115
rect 16740 -1140 16780 -1135
rect 16740 -1170 16745 -1140
rect 16775 -1145 16780 -1140
rect 16820 -1140 16860 -1135
rect 16820 -1145 16825 -1140
rect 16775 -1165 16825 -1145
rect 16775 -1170 16780 -1165
rect 16740 -1175 16780 -1170
rect 16820 -1170 16825 -1165
rect 16855 -1145 16860 -1140
rect 16900 -1140 16940 -1135
rect 16900 -1145 16905 -1140
rect 16855 -1165 16905 -1145
rect 16855 -1170 16860 -1165
rect 16820 -1175 16860 -1170
rect 16900 -1170 16905 -1165
rect 16935 -1145 16940 -1140
rect 16980 -1140 17020 -1135
rect 16980 -1145 16985 -1140
rect 16935 -1165 16985 -1145
rect 16935 -1170 16940 -1165
rect 16900 -1175 16940 -1170
rect 16980 -1170 16985 -1165
rect 17015 -1145 17020 -1140
rect 17060 -1140 17100 -1135
rect 17060 -1145 17065 -1140
rect 17015 -1165 17065 -1145
rect 17015 -1170 17020 -1165
rect 16980 -1175 17020 -1170
rect 17060 -1170 17065 -1165
rect 17095 -1145 17100 -1140
rect 17140 -1140 17180 -1135
rect 17140 -1145 17145 -1140
rect 17095 -1165 17145 -1145
rect 17095 -1170 17100 -1165
rect 17060 -1175 17100 -1170
rect 17140 -1170 17145 -1165
rect 17175 -1145 17180 -1140
rect 17220 -1140 17260 -1135
rect 17220 -1145 17225 -1140
rect 17175 -1165 17225 -1145
rect 17175 -1170 17180 -1165
rect 17140 -1175 17180 -1170
rect 17220 -1170 17225 -1165
rect 17255 -1145 17260 -1140
rect 17300 -1140 17340 -1135
rect 17300 -1145 17305 -1140
rect 17255 -1165 17305 -1145
rect 17255 -1170 17260 -1165
rect 17220 -1175 17260 -1170
rect 17300 -1170 17305 -1165
rect 17335 -1145 17340 -1140
rect 17380 -1140 17420 -1135
rect 17380 -1145 17385 -1140
rect 17335 -1165 17385 -1145
rect 17335 -1170 17340 -1165
rect 17300 -1175 17340 -1170
rect 17380 -1170 17385 -1165
rect 17415 -1145 17420 -1140
rect 17460 -1140 17500 -1135
rect 17460 -1145 17465 -1140
rect 17415 -1165 17465 -1145
rect 17415 -1170 17420 -1165
rect 17380 -1175 17420 -1170
rect 17460 -1170 17465 -1165
rect 17495 -1145 17500 -1140
rect 17540 -1140 17580 -1135
rect 17540 -1145 17545 -1140
rect 17495 -1165 17545 -1145
rect 17495 -1170 17500 -1165
rect 17460 -1175 17500 -1170
rect 17540 -1170 17545 -1165
rect 17575 -1145 17580 -1140
rect 17620 -1140 17660 -1135
rect 17620 -1145 17625 -1140
rect 17575 -1165 17625 -1145
rect 17575 -1170 17580 -1165
rect 17540 -1175 17580 -1170
rect 17620 -1170 17625 -1165
rect 17655 -1145 17660 -1140
rect 17700 -1140 17740 -1135
rect 17700 -1145 17705 -1140
rect 17655 -1165 17705 -1145
rect 17655 -1170 17660 -1165
rect 17620 -1175 17660 -1170
rect 17700 -1170 17705 -1165
rect 17735 -1170 17740 -1140
rect 17700 -1175 17740 -1170
rect 17780 -1140 17820 -1135
rect 17780 -1170 17785 -1140
rect 17815 -1145 17820 -1140
rect 17860 -1140 17900 -1135
rect 17860 -1145 17865 -1140
rect 17815 -1165 17865 -1145
rect 17815 -1170 17820 -1165
rect 17780 -1175 17820 -1170
rect 17860 -1170 17865 -1165
rect 17895 -1145 17900 -1140
rect 17940 -1140 17980 -1135
rect 17940 -1145 17945 -1140
rect 17895 -1165 17945 -1145
rect 17895 -1170 17900 -1165
rect 17860 -1175 17900 -1170
rect 17940 -1170 17945 -1165
rect 17975 -1145 17980 -1140
rect 18020 -1140 18060 -1135
rect 18020 -1145 18025 -1140
rect 17975 -1165 18025 -1145
rect 17975 -1170 17980 -1165
rect 17940 -1175 17980 -1170
rect 18020 -1170 18025 -1165
rect 18055 -1145 18060 -1140
rect 18100 -1140 18140 -1135
rect 18100 -1145 18105 -1140
rect 18055 -1165 18105 -1145
rect 18055 -1170 18060 -1165
rect 18020 -1175 18060 -1170
rect 18100 -1170 18105 -1165
rect 18135 -1145 18140 -1140
rect 18180 -1140 18220 -1135
rect 18180 -1145 18185 -1140
rect 18135 -1165 18185 -1145
rect 18135 -1170 18140 -1165
rect 18100 -1175 18140 -1170
rect 18180 -1170 18185 -1165
rect 18215 -1145 18220 -1140
rect 18260 -1140 18300 -1135
rect 18260 -1145 18265 -1140
rect 18215 -1165 18265 -1145
rect 18215 -1170 18220 -1165
rect 18180 -1175 18220 -1170
rect 18260 -1170 18265 -1165
rect 18295 -1145 18300 -1140
rect 18340 -1140 18380 -1135
rect 18340 -1145 18345 -1140
rect 18295 -1165 18345 -1145
rect 18295 -1170 18300 -1165
rect 18260 -1175 18300 -1170
rect 18340 -1170 18345 -1165
rect 18375 -1145 18380 -1140
rect 18420 -1140 18460 -1135
rect 18420 -1145 18425 -1140
rect 18375 -1165 18425 -1145
rect 18375 -1170 18380 -1165
rect 18340 -1175 18380 -1170
rect 18420 -1170 18425 -1165
rect 18455 -1145 18460 -1140
rect 18500 -1140 18540 -1135
rect 18500 -1145 18505 -1140
rect 18455 -1165 18505 -1145
rect 18455 -1170 18460 -1165
rect 18420 -1175 18460 -1170
rect 18500 -1170 18505 -1165
rect 18535 -1145 18540 -1140
rect 18580 -1140 18620 -1135
rect 18580 -1145 18585 -1140
rect 18535 -1165 18585 -1145
rect 18535 -1170 18540 -1165
rect 18500 -1175 18540 -1170
rect 18580 -1170 18585 -1165
rect 18615 -1145 18620 -1140
rect 18660 -1140 18700 -1135
rect 18660 -1145 18665 -1140
rect 18615 -1165 18665 -1145
rect 18615 -1170 18620 -1165
rect 18580 -1175 18620 -1170
rect 18660 -1170 18665 -1165
rect 18695 -1145 18700 -1140
rect 18740 -1140 18780 -1135
rect 18740 -1145 18745 -1140
rect 18695 -1165 18745 -1145
rect 18695 -1170 18700 -1165
rect 18660 -1175 18700 -1170
rect 18740 -1170 18745 -1165
rect 18775 -1170 18780 -1140
rect 18740 -1175 18780 -1170
rect 18895 -1205 18935 -1200
rect 16205 -1225 16245 -1220
rect 16205 -1255 16210 -1225
rect 16240 -1230 16245 -1225
rect 16700 -1225 16740 -1220
rect 16700 -1230 16705 -1225
rect 16240 -1250 16705 -1230
rect 16240 -1255 16245 -1250
rect 16205 -1260 16245 -1255
rect 16700 -1255 16705 -1250
rect 16735 -1255 16740 -1225
rect 16700 -1260 16740 -1255
rect 18895 -1235 18900 -1205
rect 18930 -1235 18935 -1205
rect 18895 -1245 18935 -1235
rect 18895 -1275 18900 -1245
rect 18930 -1275 18935 -1245
rect 18895 -1280 18935 -1275
rect 16160 -1325 16200 -1320
rect 16160 -1355 16165 -1325
rect 16195 -1330 16200 -1325
rect 16595 -1325 16635 -1320
rect 16595 -1330 16600 -1325
rect 16195 -1350 16600 -1330
rect 16195 -1355 16200 -1350
rect 16160 -1360 16200 -1355
rect 16595 -1355 16600 -1350
rect 16630 -1330 16635 -1325
rect 16705 -1325 16745 -1320
rect 16705 -1330 16710 -1325
rect 16630 -1350 16710 -1330
rect 16630 -1355 16635 -1350
rect 16595 -1360 16635 -1355
rect 16705 -1355 16710 -1350
rect 16740 -1330 16745 -1325
rect 17300 -1325 17340 -1320
rect 17300 -1330 17305 -1325
rect 16740 -1350 17305 -1330
rect 16740 -1355 16745 -1350
rect 16705 -1360 16745 -1355
rect 17300 -1355 17305 -1350
rect 17335 -1330 17340 -1325
rect 17780 -1325 17820 -1320
rect 17780 -1330 17785 -1325
rect 17335 -1350 17785 -1330
rect 17335 -1355 17340 -1350
rect 17300 -1360 17340 -1355
rect 17780 -1355 17785 -1350
rect 17815 -1330 17820 -1325
rect 18260 -1325 18300 -1320
rect 18260 -1330 18265 -1325
rect 17815 -1350 18265 -1330
rect 17815 -1355 17820 -1350
rect 17780 -1360 17820 -1355
rect 18260 -1355 18265 -1350
rect 18295 -1355 18300 -1325
rect 18260 -1360 18300 -1355
rect 16540 -1410 18575 -1405
rect 16540 -1440 16545 -1410
rect 16575 -1440 16655 -1410
rect 16685 -1440 16765 -1410
rect 16795 -1440 16825 -1410
rect 16855 -1440 17030 -1410
rect 17060 -1440 17140 -1410
rect 17170 -1440 17250 -1410
rect 17280 -1440 17360 -1410
rect 17390 -1440 17470 -1410
rect 17500 -1440 17620 -1410
rect 17650 -1440 17730 -1410
rect 17760 -1440 17840 -1410
rect 17870 -1440 17950 -1410
rect 17980 -1440 18100 -1410
rect 18130 -1440 18210 -1410
rect 18240 -1440 18320 -1410
rect 18350 -1440 18430 -1410
rect 18460 -1440 18540 -1410
rect 18570 -1440 18575 -1410
rect 16540 -1450 18575 -1440
rect 16540 -1480 16545 -1450
rect 16575 -1480 16655 -1450
rect 16685 -1480 16765 -1450
rect 16795 -1480 16825 -1450
rect 16855 -1480 17030 -1450
rect 17060 -1480 17140 -1450
rect 17170 -1480 17250 -1450
rect 17280 -1480 17360 -1450
rect 17390 -1480 17470 -1450
rect 17500 -1480 17620 -1450
rect 17650 -1480 17730 -1450
rect 17760 -1480 17840 -1450
rect 17870 -1480 17950 -1450
rect 17980 -1480 18100 -1450
rect 18130 -1480 18210 -1450
rect 18240 -1480 18320 -1450
rect 18350 -1480 18430 -1450
rect 18460 -1480 18540 -1450
rect 18570 -1480 18575 -1450
rect 16540 -1490 18575 -1480
rect 16540 -1520 16545 -1490
rect 16575 -1520 16655 -1490
rect 16685 -1520 16765 -1490
rect 16795 -1520 16825 -1490
rect 16855 -1520 17030 -1490
rect 17060 -1520 17140 -1490
rect 17170 -1520 17250 -1490
rect 17280 -1520 17360 -1490
rect 17390 -1520 17470 -1490
rect 17500 -1520 17620 -1490
rect 17650 -1520 17730 -1490
rect 17760 -1520 17840 -1490
rect 17870 -1520 17950 -1490
rect 17980 -1520 18100 -1490
rect 18130 -1520 18210 -1490
rect 18240 -1520 18320 -1490
rect 18350 -1520 18430 -1490
rect 18460 -1520 18540 -1490
rect 18570 -1520 18575 -1490
rect 16540 -1525 18575 -1520
rect 17190 -1660 17450 -1655
rect 17190 -1690 17195 -1660
rect 17225 -1690 17415 -1660
rect 17445 -1690 17450 -1660
rect 17190 -1695 17450 -1690
rect 17670 -1660 17710 -1655
rect 17670 -1690 17675 -1660
rect 17705 -1665 17710 -1660
rect 17780 -1660 17820 -1655
rect 17780 -1665 17785 -1660
rect 17705 -1685 17785 -1665
rect 17705 -1690 17710 -1685
rect 17670 -1695 17710 -1690
rect 17780 -1690 17785 -1685
rect 17815 -1665 17820 -1660
rect 17890 -1660 17930 -1655
rect 17890 -1665 17895 -1660
rect 17815 -1685 17895 -1665
rect 17815 -1690 17820 -1685
rect 17780 -1695 17820 -1690
rect 17890 -1690 17895 -1685
rect 17925 -1690 17930 -1660
rect 17890 -1695 17930 -1690
rect 18150 -1660 18410 -1655
rect 18150 -1690 18155 -1660
rect 18185 -1690 18375 -1660
rect 18405 -1690 18410 -1660
rect 18150 -1695 18410 -1690
rect 16030 -1715 16070 -1710
rect 16030 -1745 16035 -1715
rect 16065 -1720 16070 -1715
rect 17080 -1715 17120 -1710
rect 17080 -1720 17085 -1715
rect 16065 -1740 17085 -1720
rect 16065 -1745 16070 -1740
rect 16030 -1750 16070 -1745
rect 17080 -1745 17085 -1740
rect 17115 -1720 17120 -1715
rect 17300 -1715 17340 -1710
rect 17300 -1720 17305 -1715
rect 17115 -1740 17305 -1720
rect 17115 -1745 17120 -1740
rect 17080 -1750 17120 -1745
rect 17300 -1745 17305 -1740
rect 17335 -1720 17340 -1715
rect 18260 -1715 18300 -1710
rect 18260 -1720 18265 -1715
rect 17335 -1740 18265 -1720
rect 17335 -1745 17340 -1740
rect 17300 -1750 17340 -1745
rect 18260 -1745 18265 -1740
rect 18295 -1720 18300 -1715
rect 18480 -1715 18520 -1710
rect 18480 -1720 18485 -1715
rect 18295 -1740 18485 -1720
rect 18295 -1745 18300 -1740
rect 18260 -1750 18300 -1745
rect 18480 -1745 18485 -1740
rect 18515 -1745 18520 -1715
rect 18480 -1750 18520 -1745
rect 15785 -1770 17230 -1765
rect 15785 -1800 15790 -1770
rect 15820 -1800 17195 -1770
rect 17225 -1800 17230 -1770
rect 15785 -1810 17230 -1800
rect 15785 -1840 15790 -1810
rect 15820 -1840 17195 -1810
rect 17225 -1840 17230 -1810
rect 15785 -1845 17230 -1840
rect 18370 -1770 19815 -1765
rect 18370 -1800 18375 -1770
rect 18405 -1800 19780 -1770
rect 19810 -1800 19815 -1770
rect 18370 -1810 19815 -1800
rect 18370 -1840 18375 -1810
rect 18405 -1840 19780 -1810
rect 19810 -1840 19815 -1810
rect 18370 -1845 19815 -1840
rect 16105 -1900 16145 -1895
rect 16105 -1930 16110 -1900
rect 16140 -1905 16145 -1900
rect 16705 -1900 16745 -1895
rect 16705 -1905 16710 -1900
rect 16140 -1925 16710 -1905
rect 16140 -1930 16145 -1925
rect 16105 -1935 16145 -1930
rect 16705 -1930 16710 -1925
rect 16740 -1930 16745 -1900
rect 16705 -1935 16745 -1930
rect 17780 -1900 17820 -1895
rect 17780 -1930 17785 -1900
rect 17815 -1905 17820 -1900
rect 19535 -1900 19575 -1895
rect 19535 -1905 19540 -1900
rect 17815 -1925 19540 -1905
rect 17815 -1930 17820 -1925
rect 17780 -1935 17820 -1930
rect 19535 -1930 19540 -1925
rect 19570 -1930 19575 -1900
rect 19535 -1935 19575 -1930
rect 16155 -1950 16195 -1945
rect 16155 -1980 16160 -1950
rect 16190 -1955 16195 -1950
rect 19325 -1950 19365 -1945
rect 19325 -1955 19330 -1950
rect 16190 -1975 19330 -1955
rect 16190 -1980 16195 -1975
rect 16155 -1985 16195 -1980
rect 19325 -1980 19330 -1975
rect 19360 -1980 19365 -1950
rect 19325 -1985 19365 -1980
rect 16260 -2000 16300 -1995
rect 16260 -2030 16265 -2000
rect 16295 -2005 16300 -2000
rect 16480 -2000 16520 -1995
rect 16480 -2005 16485 -2000
rect 16295 -2025 16485 -2005
rect 16295 -2030 16300 -2025
rect 16260 -2035 16300 -2030
rect 16480 -2030 16485 -2025
rect 16515 -2005 16520 -2000
rect 16730 -2000 16770 -1995
rect 16730 -2005 16735 -2000
rect 16515 -2025 16735 -2005
rect 16515 -2030 16520 -2025
rect 16480 -2035 16520 -2030
rect 16730 -2030 16735 -2025
rect 16765 -2030 16770 -2000
rect 16730 -2035 16770 -2030
rect 17195 -2000 17425 -1995
rect 17195 -2030 17200 -2000
rect 17230 -2030 17430 -2000
rect 17195 -2035 17430 -2030
rect 17465 -2035 17470 -2000
rect 18124 -2035 18129 -2000
rect 18164 -2005 19500 -2000
rect 18164 -2035 19085 -2005
rect 19115 -2035 19465 -2005
rect 19495 -2035 19500 -2005
rect 18165 -2040 19500 -2035
rect 17195 -2060 17235 -2055
rect 17195 -2090 17200 -2060
rect 17230 -2065 17235 -2060
rect 18830 -2060 18870 -2055
rect 18830 -2065 18835 -2060
rect 17230 -2085 18835 -2065
rect 17230 -2090 17235 -2085
rect 17195 -2095 17235 -2090
rect 18830 -2090 18835 -2085
rect 18865 -2090 18870 -2060
rect 18830 -2095 18870 -2090
rect 16485 -2900 16520 -2895
rect 16485 -2940 16520 -2935
rect 19080 -2900 19115 -2895
rect 19080 -2940 19115 -2935
rect 19405 -2997 19440 -2992
rect 16160 -3025 16195 -3020
rect 19405 -3037 19440 -3032
rect 16160 -3065 16195 -3060
rect 16730 -3105 16770 -3100
rect 15820 -3115 15860 -3110
rect 15960 -3111 15980 -3110
rect 15820 -3145 15825 -3115
rect 15855 -3120 15860 -3115
rect 15950 -3116 15985 -3111
rect 15855 -3140 15950 -3120
rect 15855 -3145 15860 -3140
rect 15820 -3150 15860 -3145
rect 16730 -3135 16735 -3105
rect 16765 -3110 16770 -3105
rect 17780 -3105 17820 -3100
rect 17780 -3110 17785 -3105
rect 16765 -3130 17785 -3110
rect 16765 -3135 16770 -3130
rect 16730 -3140 16770 -3135
rect 17780 -3135 17785 -3130
rect 17815 -3135 17820 -3105
rect 17780 -3140 17820 -3135
rect 18615 -3105 18655 -3100
rect 18615 -3135 18620 -3105
rect 18650 -3110 18655 -3105
rect 18830 -3105 18870 -3100
rect 18830 -3110 18835 -3105
rect 18650 -3130 18835 -3110
rect 18650 -3135 18655 -3130
rect 18615 -3140 18655 -3135
rect 18830 -3135 18835 -3130
rect 18865 -3135 18870 -3105
rect 18830 -3140 18870 -3135
rect 19610 -3116 19645 -3111
rect 15950 -3156 15985 -3151
rect 19610 -3156 19645 -3151
rect 15950 -3789 15985 -3784
rect 15950 -3829 15985 -3824
rect 19610 -3789 19645 -3784
rect 19610 -3829 19645 -3824
rect 15960 -3830 15980 -3829
rect 19620 -3830 19640 -3829
rect 16280 -3894 16315 -3889
rect 16280 -3934 16315 -3929
rect 19285 -3894 19320 -3889
rect 19285 -3934 19320 -3929
rect 16290 -3935 16310 -3934
rect 19290 -3935 19310 -3934
rect 16605 -3969 16640 -3964
rect 16605 -4009 16640 -4004
rect 18960 -3969 18995 -3964
rect 18960 -4009 18995 -4004
rect 16615 -4010 16635 -4009
rect 18965 -4010 18985 -4009
rect 16280 -4190 16320 -4185
rect 16280 -4195 16285 -4190
rect 15665 -4215 16285 -4195
rect 16280 -4220 16285 -4215
rect 16315 -4195 16320 -4190
rect 16605 -4190 16645 -4185
rect 16605 -4195 16610 -4190
rect 16315 -4215 16610 -4195
rect 16315 -4220 16320 -4215
rect 16280 -4225 16320 -4220
rect 16605 -4220 16610 -4215
rect 16640 -4220 16645 -4190
rect 16605 -4225 16645 -4220
rect 15820 -4265 15860 -4260
rect 15820 -4295 15825 -4265
rect 15855 -4270 15860 -4265
rect 17250 -4265 17300 -4255
rect 17250 -4270 17260 -4265
rect 15855 -4290 17260 -4270
rect 15855 -4295 15860 -4290
rect 15820 -4300 15860 -4295
rect 17250 -4295 17260 -4290
rect 17290 -4295 17300 -4265
rect 17250 -4305 17300 -4295
rect 17780 -4265 17820 -4260
rect 17780 -4295 17785 -4265
rect 17815 -4270 17820 -4265
rect 18955 -4265 18995 -4260
rect 18955 -4270 18960 -4265
rect 17815 -4290 18960 -4270
rect 17815 -4295 17820 -4290
rect 17780 -4300 17820 -4295
rect 18955 -4295 18960 -4290
rect 18990 -4270 18995 -4265
rect 19280 -4265 19320 -4260
rect 19280 -4270 19285 -4265
rect 18990 -4290 19285 -4270
rect 18990 -4295 18995 -4290
rect 18955 -4300 18995 -4295
rect 19280 -4295 19285 -4290
rect 19315 -4295 19320 -4265
rect 19280 -4300 19320 -4295
rect 15725 -4315 15765 -4310
rect 15725 -4345 15730 -4315
rect 15760 -4320 15765 -4315
rect 16900 -4315 16950 -4305
rect 16900 -4320 16910 -4315
rect 15760 -4340 16910 -4320
rect 15760 -4345 15765 -4340
rect 15725 -4350 15765 -4345
rect 16900 -4345 16910 -4340
rect 16940 -4345 16950 -4315
rect 16900 -4355 16950 -4345
rect 18650 -4315 18700 -4305
rect 18650 -4345 18660 -4315
rect 18690 -4320 18700 -4315
rect 19720 -4315 19760 -4310
rect 19720 -4320 19725 -4315
rect 18690 -4340 19725 -4320
rect 18690 -4345 18700 -4340
rect 18650 -4355 18700 -4345
rect 19720 -4345 19725 -4340
rect 19755 -4345 19760 -4315
rect 19720 -4350 19760 -4345
rect 15950 -4360 15990 -4355
rect 15950 -4390 15955 -4360
rect 15985 -4365 15990 -4360
rect 16205 -4360 16245 -4355
rect 16205 -4365 16210 -4360
rect 15985 -4385 16210 -4365
rect 15985 -4390 15990 -4385
rect 15950 -4395 15990 -4390
rect 16205 -4390 16210 -4385
rect 16240 -4390 16245 -4360
rect 16205 -4395 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4365 19395 -4360
rect 19610 -4360 19650 -4355
rect 19610 -4365 19615 -4360
rect 19390 -4385 19615 -4365
rect 19390 -4390 19395 -4385
rect 19355 -4395 19395 -4390
rect 19610 -4390 19615 -4385
rect 19645 -4390 19650 -4360
rect 19610 -4395 19650 -4390
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4415 17995 -4410
rect 17990 -4435 19905 -4415
rect 17990 -4440 17995 -4435
rect 17955 -4445 17995 -4440
<< via2 >>
rect 17260 -4295 17290 -4265
rect 16910 -4345 16940 -4315
rect 18660 -4345 18690 -4315
rect 16210 -4390 16240 -4360
rect 19360 -4390 19390 -4360
rect 17960 -4440 17990 -4410
<< metal3 >>
rect 17250 -4260 17300 -4255
rect 17250 -4300 17255 -4260
rect 17295 -4300 17300 -4260
rect 17250 -4305 17300 -4300
rect 16900 -4310 16950 -4305
rect 16900 -4350 16905 -4310
rect 16945 -4350 16950 -4310
rect 16900 -4355 16950 -4350
rect 18650 -4310 18700 -4305
rect 18650 -4350 18655 -4310
rect 18695 -4350 18700 -4310
rect 18650 -4355 18700 -4350
rect 16205 -4360 16245 -4355
rect 16205 -4390 16210 -4360
rect 16240 -4390 16245 -4360
rect 16205 -4520 16245 -4390
rect 19355 -4360 19395 -4355
rect 19355 -4390 19360 -4360
rect 19390 -4390 19395 -4360
rect 17955 -4410 17995 -4405
rect 17955 -4440 17960 -4410
rect 17990 -4440 17995 -4410
rect 17955 -4520 17995 -4440
rect 19355 -4520 19395 -4390
rect 15760 -4615 15990 -4520
rect 16110 -4615 16340 -4520
rect 16460 -4615 16690 -4520
rect 16810 -4615 17040 -4520
rect 15760 -4665 17040 -4615
rect 15760 -4750 15990 -4665
rect 16110 -4750 16340 -4665
rect 16460 -4750 16690 -4665
rect 16810 -4750 17040 -4665
rect 17160 -4615 17390 -4520
rect 17510 -4615 17740 -4520
rect 17860 -4615 18090 -4520
rect 18210 -4615 18440 -4520
rect 17160 -4665 18440 -4615
rect 17160 -4750 17390 -4665
rect 17510 -4750 17740 -4665
rect 17860 -4750 18090 -4665
rect 18210 -4750 18440 -4665
rect 18560 -4615 18790 -4520
rect 18910 -4615 19140 -4520
rect 19260 -4615 19490 -4520
rect 19610 -4615 19840 -4520
rect 18560 -4665 19840 -4615
rect 18560 -4750 18790 -4665
rect 18910 -4750 19140 -4665
rect 19260 -4750 19490 -4665
rect 19610 -4750 19840 -4665
rect 16200 -4870 16250 -4750
rect 17950 -4870 18000 -4750
rect 19350 -4870 19400 -4750
rect 15760 -4965 15990 -4870
rect 16110 -4965 16340 -4870
rect 16460 -4965 16690 -4870
rect 16810 -4965 17040 -4870
rect 15760 -5015 17040 -4965
rect 15760 -5100 15990 -5015
rect 16110 -5100 16340 -5015
rect 16460 -5100 16690 -5015
rect 16810 -5100 17040 -5015
rect 17160 -4965 17390 -4870
rect 17510 -4965 17740 -4870
rect 17860 -4965 18090 -4870
rect 18210 -4965 18440 -4870
rect 17160 -5015 18440 -4965
rect 17160 -5100 17390 -5015
rect 17510 -5100 17740 -5015
rect 17860 -5100 18090 -5015
rect 18210 -5100 18440 -5015
rect 18560 -4965 18790 -4870
rect 18910 -4965 19140 -4870
rect 19260 -4965 19490 -4870
rect 19610 -4965 19840 -4870
rect 18560 -5015 19840 -4965
rect 18560 -5100 18790 -5015
rect 18910 -5100 19140 -5015
rect 19260 -5100 19490 -5015
rect 19610 -5100 19840 -5015
rect 16200 -5220 16250 -5100
rect 17950 -5220 18000 -5100
rect 19350 -5220 19400 -5100
rect 15760 -5315 15990 -5220
rect 16110 -5315 16340 -5220
rect 16460 -5315 16690 -5220
rect 16810 -5315 17040 -5220
rect 15760 -5365 17040 -5315
rect 15760 -5450 15990 -5365
rect 16110 -5450 16340 -5365
rect 16460 -5450 16690 -5365
rect 16810 -5450 17040 -5365
rect 17160 -5315 17390 -5220
rect 17510 -5315 17740 -5220
rect 17860 -5315 18090 -5220
rect 18210 -5315 18440 -5220
rect 17160 -5365 18440 -5315
rect 17160 -5450 17390 -5365
rect 17510 -5450 17740 -5365
rect 17860 -5450 18090 -5365
rect 18210 -5450 18440 -5365
rect 18560 -5315 18790 -5220
rect 18910 -5315 19140 -5220
rect 19260 -5315 19490 -5220
rect 19610 -5315 19840 -5220
rect 18560 -5365 19840 -5315
rect 18560 -5450 18790 -5365
rect 18910 -5450 19140 -5365
rect 19260 -5450 19490 -5365
rect 19610 -5450 19840 -5365
rect 16200 -5570 16250 -5450
rect 17950 -5570 18000 -5450
rect 19350 -5570 19400 -5450
rect 15760 -5665 15990 -5570
rect 16110 -5665 16340 -5570
rect 16460 -5665 16690 -5570
rect 16810 -5665 17040 -5570
rect 15760 -5715 17040 -5665
rect 15760 -5800 15990 -5715
rect 16110 -5800 16340 -5715
rect 16460 -5800 16690 -5715
rect 16810 -5800 17040 -5715
rect 17160 -5665 17390 -5570
rect 17510 -5665 17740 -5570
rect 17860 -5665 18090 -5570
rect 18210 -5665 18440 -5570
rect 17160 -5715 18440 -5665
rect 17160 -5800 17390 -5715
rect 17510 -5800 17740 -5715
rect 17860 -5800 18090 -5715
rect 18210 -5800 18440 -5715
rect 18560 -5665 18790 -5570
rect 18910 -5665 19140 -5570
rect 19260 -5665 19490 -5570
rect 19610 -5665 19840 -5570
rect 18560 -5715 19840 -5665
rect 18560 -5800 18790 -5715
rect 18910 -5800 19140 -5715
rect 19260 -5800 19490 -5715
rect 19610 -5800 19840 -5715
rect 16200 -5920 16250 -5800
rect 17950 -5920 18000 -5800
rect 19350 -5920 19400 -5800
rect 15760 -6015 15990 -5920
rect 16110 -6015 16340 -5920
rect 16460 -6015 16690 -5920
rect 16810 -6015 17040 -5920
rect 15760 -6065 17040 -6015
rect 15760 -6150 15990 -6065
rect 16110 -6150 16340 -6065
rect 16460 -6150 16690 -6065
rect 16810 -6150 17040 -6065
rect 17160 -6015 17390 -5920
rect 17510 -6015 17740 -5920
rect 17860 -6015 18090 -5920
rect 18210 -6015 18440 -5920
rect 17160 -6065 18440 -6015
rect 17160 -6150 17390 -6065
rect 17510 -6150 17740 -6065
rect 17860 -6150 18090 -6065
rect 18210 -6150 18440 -6065
rect 18560 -6015 18790 -5920
rect 18910 -6015 19140 -5920
rect 19260 -6015 19490 -5920
rect 19610 -6015 19840 -5920
rect 18560 -6065 19840 -6015
rect 18560 -6150 18790 -6065
rect 18910 -6150 19140 -6065
rect 19260 -6150 19490 -6065
rect 19610 -6150 19840 -6065
<< via3 >>
rect 17255 -4265 17295 -4260
rect 17255 -4295 17260 -4265
rect 17260 -4295 17290 -4265
rect 17290 -4295 17295 -4265
rect 17255 -4300 17295 -4295
rect 16905 -4315 16945 -4310
rect 16905 -4345 16910 -4315
rect 16910 -4345 16940 -4315
rect 16940 -4345 16945 -4315
rect 16905 -4350 16945 -4345
rect 18655 -4315 18695 -4310
rect 18655 -4345 18660 -4315
rect 18660 -4345 18690 -4315
rect 18690 -4345 18695 -4315
rect 18655 -4350 18695 -4345
<< mimcap >>
rect 15775 -4620 15975 -4535
rect 15775 -4660 15855 -4620
rect 15895 -4660 15975 -4620
rect 15775 -4735 15975 -4660
rect 16125 -4620 16325 -4535
rect 16125 -4660 16205 -4620
rect 16245 -4660 16325 -4620
rect 16125 -4735 16325 -4660
rect 16475 -4620 16675 -4535
rect 16475 -4660 16555 -4620
rect 16595 -4660 16675 -4620
rect 16475 -4735 16675 -4660
rect 16825 -4620 17025 -4535
rect 16825 -4660 16905 -4620
rect 16945 -4660 17025 -4620
rect 16825 -4735 17025 -4660
rect 17175 -4620 17375 -4535
rect 17175 -4660 17255 -4620
rect 17295 -4660 17375 -4620
rect 17175 -4735 17375 -4660
rect 17525 -4620 17725 -4535
rect 17525 -4660 17605 -4620
rect 17645 -4660 17725 -4620
rect 17525 -4735 17725 -4660
rect 17875 -4620 18075 -4535
rect 17875 -4660 17955 -4620
rect 17995 -4660 18075 -4620
rect 17875 -4735 18075 -4660
rect 18225 -4620 18425 -4535
rect 18225 -4660 18305 -4620
rect 18345 -4660 18425 -4620
rect 18225 -4735 18425 -4660
rect 18575 -4620 18775 -4535
rect 18575 -4660 18655 -4620
rect 18695 -4660 18775 -4620
rect 18575 -4735 18775 -4660
rect 18925 -4620 19125 -4535
rect 18925 -4660 19005 -4620
rect 19045 -4660 19125 -4620
rect 18925 -4735 19125 -4660
rect 19275 -4620 19475 -4535
rect 19275 -4660 19355 -4620
rect 19395 -4660 19475 -4620
rect 19275 -4735 19475 -4660
rect 19625 -4620 19825 -4535
rect 19625 -4660 19705 -4620
rect 19745 -4660 19825 -4620
rect 19625 -4735 19825 -4660
rect 15775 -4970 15975 -4885
rect 15775 -5010 15855 -4970
rect 15895 -5010 15975 -4970
rect 15775 -5085 15975 -5010
rect 16125 -4970 16325 -4885
rect 16125 -5010 16205 -4970
rect 16245 -5010 16325 -4970
rect 16125 -5085 16325 -5010
rect 16475 -4970 16675 -4885
rect 16475 -5010 16555 -4970
rect 16595 -5010 16675 -4970
rect 16475 -5085 16675 -5010
rect 16825 -4970 17025 -4885
rect 16825 -5010 16905 -4970
rect 16945 -5010 17025 -4970
rect 16825 -5085 17025 -5010
rect 17175 -4970 17375 -4885
rect 17175 -5010 17255 -4970
rect 17295 -5010 17375 -4970
rect 17175 -5085 17375 -5010
rect 17525 -4970 17725 -4885
rect 17525 -5010 17605 -4970
rect 17645 -5010 17725 -4970
rect 17525 -5085 17725 -5010
rect 17875 -4970 18075 -4885
rect 17875 -5010 17955 -4970
rect 17995 -5010 18075 -4970
rect 17875 -5085 18075 -5010
rect 18225 -4970 18425 -4885
rect 18225 -5010 18305 -4970
rect 18345 -5010 18425 -4970
rect 18225 -5085 18425 -5010
rect 18575 -4970 18775 -4885
rect 18575 -5010 18655 -4970
rect 18695 -5010 18775 -4970
rect 18575 -5085 18775 -5010
rect 18925 -4970 19125 -4885
rect 18925 -5010 19005 -4970
rect 19045 -5010 19125 -4970
rect 18925 -5085 19125 -5010
rect 19275 -4970 19475 -4885
rect 19275 -5010 19355 -4970
rect 19395 -5010 19475 -4970
rect 19275 -5085 19475 -5010
rect 19625 -4970 19825 -4885
rect 19625 -5010 19705 -4970
rect 19745 -5010 19825 -4970
rect 19625 -5085 19825 -5010
rect 15775 -5320 15975 -5235
rect 15775 -5360 15855 -5320
rect 15895 -5360 15975 -5320
rect 15775 -5435 15975 -5360
rect 16125 -5320 16325 -5235
rect 16125 -5360 16205 -5320
rect 16245 -5360 16325 -5320
rect 16125 -5435 16325 -5360
rect 16475 -5320 16675 -5235
rect 16475 -5360 16555 -5320
rect 16595 -5360 16675 -5320
rect 16475 -5435 16675 -5360
rect 16825 -5320 17025 -5235
rect 16825 -5360 16905 -5320
rect 16945 -5360 17025 -5320
rect 16825 -5435 17025 -5360
rect 17175 -5320 17375 -5235
rect 17175 -5360 17255 -5320
rect 17295 -5360 17375 -5320
rect 17175 -5435 17375 -5360
rect 17525 -5320 17725 -5235
rect 17525 -5360 17605 -5320
rect 17645 -5360 17725 -5320
rect 17525 -5435 17725 -5360
rect 17875 -5320 18075 -5235
rect 17875 -5360 17955 -5320
rect 17995 -5360 18075 -5320
rect 17875 -5435 18075 -5360
rect 18225 -5320 18425 -5235
rect 18225 -5360 18305 -5320
rect 18345 -5360 18425 -5320
rect 18225 -5435 18425 -5360
rect 18575 -5320 18775 -5235
rect 18575 -5360 18655 -5320
rect 18695 -5360 18775 -5320
rect 18575 -5435 18775 -5360
rect 18925 -5320 19125 -5235
rect 18925 -5360 19005 -5320
rect 19045 -5360 19125 -5320
rect 18925 -5435 19125 -5360
rect 19275 -5320 19475 -5235
rect 19275 -5360 19355 -5320
rect 19395 -5360 19475 -5320
rect 19275 -5435 19475 -5360
rect 19625 -5320 19825 -5235
rect 19625 -5360 19705 -5320
rect 19745 -5360 19825 -5320
rect 19625 -5435 19825 -5360
rect 15775 -5670 15975 -5585
rect 15775 -5710 15855 -5670
rect 15895 -5710 15975 -5670
rect 15775 -5785 15975 -5710
rect 16125 -5670 16325 -5585
rect 16125 -5710 16205 -5670
rect 16245 -5710 16325 -5670
rect 16125 -5785 16325 -5710
rect 16475 -5670 16675 -5585
rect 16475 -5710 16555 -5670
rect 16595 -5710 16675 -5670
rect 16475 -5785 16675 -5710
rect 16825 -5670 17025 -5585
rect 16825 -5710 16905 -5670
rect 16945 -5710 17025 -5670
rect 16825 -5785 17025 -5710
rect 17175 -5670 17375 -5585
rect 17175 -5710 17255 -5670
rect 17295 -5710 17375 -5670
rect 17175 -5785 17375 -5710
rect 17525 -5670 17725 -5585
rect 17525 -5710 17605 -5670
rect 17645 -5710 17725 -5670
rect 17525 -5785 17725 -5710
rect 17875 -5670 18075 -5585
rect 17875 -5710 17955 -5670
rect 17995 -5710 18075 -5670
rect 17875 -5785 18075 -5710
rect 18225 -5670 18425 -5585
rect 18225 -5710 18305 -5670
rect 18345 -5710 18425 -5670
rect 18225 -5785 18425 -5710
rect 18575 -5670 18775 -5585
rect 18575 -5710 18655 -5670
rect 18695 -5710 18775 -5670
rect 18575 -5785 18775 -5710
rect 18925 -5670 19125 -5585
rect 18925 -5710 19005 -5670
rect 19045 -5710 19125 -5670
rect 18925 -5785 19125 -5710
rect 19275 -5670 19475 -5585
rect 19275 -5710 19355 -5670
rect 19395 -5710 19475 -5670
rect 19275 -5785 19475 -5710
rect 19625 -5670 19825 -5585
rect 19625 -5710 19705 -5670
rect 19745 -5710 19825 -5670
rect 19625 -5785 19825 -5710
rect 15775 -6020 15975 -5935
rect 15775 -6060 15855 -6020
rect 15895 -6060 15975 -6020
rect 15775 -6135 15975 -6060
rect 16125 -6020 16325 -5935
rect 16125 -6060 16205 -6020
rect 16245 -6060 16325 -6020
rect 16125 -6135 16325 -6060
rect 16475 -6020 16675 -5935
rect 16475 -6060 16555 -6020
rect 16595 -6060 16675 -6020
rect 16475 -6135 16675 -6060
rect 16825 -6020 17025 -5935
rect 16825 -6060 16905 -6020
rect 16945 -6060 17025 -6020
rect 16825 -6135 17025 -6060
rect 17175 -6020 17375 -5935
rect 17175 -6060 17255 -6020
rect 17295 -6060 17375 -6020
rect 17175 -6135 17375 -6060
rect 17525 -6020 17725 -5935
rect 17525 -6060 17605 -6020
rect 17645 -6060 17725 -6020
rect 17525 -6135 17725 -6060
rect 17875 -6020 18075 -5935
rect 17875 -6060 17955 -6020
rect 17995 -6060 18075 -6020
rect 17875 -6135 18075 -6060
rect 18225 -6020 18425 -5935
rect 18225 -6060 18305 -6020
rect 18345 -6060 18425 -6020
rect 18225 -6135 18425 -6060
rect 18575 -6020 18775 -5935
rect 18575 -6060 18655 -6020
rect 18695 -6060 18775 -6020
rect 18575 -6135 18775 -6060
rect 18925 -6020 19125 -5935
rect 18925 -6060 19005 -6020
rect 19045 -6060 19125 -6020
rect 18925 -6135 19125 -6060
rect 19275 -6020 19475 -5935
rect 19275 -6060 19355 -6020
rect 19395 -6060 19475 -6020
rect 19275 -6135 19475 -6060
rect 19625 -6020 19825 -5935
rect 19625 -6060 19705 -6020
rect 19745 -6060 19825 -6020
rect 19625 -6135 19825 -6060
<< mimcapcontact >>
rect 15855 -4660 15895 -4620
rect 16205 -4660 16245 -4620
rect 16555 -4660 16595 -4620
rect 16905 -4660 16945 -4620
rect 17255 -4660 17295 -4620
rect 17605 -4660 17645 -4620
rect 17955 -4660 17995 -4620
rect 18305 -4660 18345 -4620
rect 18655 -4660 18695 -4620
rect 19005 -4660 19045 -4620
rect 19355 -4660 19395 -4620
rect 19705 -4660 19745 -4620
rect 15855 -5010 15895 -4970
rect 16205 -5010 16245 -4970
rect 16555 -5010 16595 -4970
rect 16905 -5010 16945 -4970
rect 17255 -5010 17295 -4970
rect 17605 -5010 17645 -4970
rect 17955 -5010 17995 -4970
rect 18305 -5010 18345 -4970
rect 18655 -5010 18695 -4970
rect 19005 -5010 19045 -4970
rect 19355 -5010 19395 -4970
rect 19705 -5010 19745 -4970
rect 15855 -5360 15895 -5320
rect 16205 -5360 16245 -5320
rect 16555 -5360 16595 -5320
rect 16905 -5360 16945 -5320
rect 17255 -5360 17295 -5320
rect 17605 -5360 17645 -5320
rect 17955 -5360 17995 -5320
rect 18305 -5360 18345 -5320
rect 18655 -5360 18695 -5320
rect 19005 -5360 19045 -5320
rect 19355 -5360 19395 -5320
rect 19705 -5360 19745 -5320
rect 15855 -5710 15895 -5670
rect 16205 -5710 16245 -5670
rect 16555 -5710 16595 -5670
rect 16905 -5710 16945 -5670
rect 17255 -5710 17295 -5670
rect 17605 -5710 17645 -5670
rect 17955 -5710 17995 -5670
rect 18305 -5710 18345 -5670
rect 18655 -5710 18695 -5670
rect 19005 -5710 19045 -5670
rect 19355 -5710 19395 -5670
rect 19705 -5710 19745 -5670
rect 15855 -6060 15895 -6020
rect 16205 -6060 16245 -6020
rect 16555 -6060 16595 -6020
rect 16905 -6060 16945 -6020
rect 17255 -6060 17295 -6020
rect 17605 -6060 17645 -6020
rect 17955 -6060 17995 -6020
rect 18305 -6060 18345 -6020
rect 18655 -6060 18695 -6020
rect 19005 -6060 19045 -6020
rect 19355 -6060 19395 -6020
rect 19705 -6060 19745 -6020
<< metal4 >>
rect 17250 -4260 17300 -4255
rect 17250 -4300 17255 -4260
rect 17295 -4300 17300 -4260
rect 16900 -4310 16950 -4305
rect 16900 -4350 16905 -4310
rect 16945 -4350 16950 -4310
rect 16900 -4615 16950 -4350
rect 15850 -4620 16950 -4615
rect 15850 -4660 15855 -4620
rect 15895 -4660 16205 -4620
rect 16245 -4660 16555 -4620
rect 16595 -4660 16905 -4620
rect 16945 -4660 16950 -4620
rect 15850 -4665 16950 -4660
rect 17250 -4615 17300 -4300
rect 18650 -4310 18700 -4305
rect 18650 -4350 18655 -4310
rect 18695 -4350 18700 -4310
rect 18650 -4615 18700 -4350
rect 17250 -4620 18350 -4615
rect 17250 -4660 17255 -4620
rect 17295 -4660 17605 -4620
rect 17645 -4660 17955 -4620
rect 17995 -4660 18305 -4620
rect 18345 -4660 18350 -4620
rect 17250 -4665 18350 -4660
rect 18650 -4620 19750 -4615
rect 18650 -4660 18655 -4620
rect 18695 -4660 19005 -4620
rect 19045 -4660 19355 -4620
rect 19395 -4660 19705 -4620
rect 19745 -4660 19750 -4620
rect 18650 -4665 19750 -4660
rect 16200 -4965 16250 -4665
rect 17950 -4965 18000 -4665
rect 19350 -4965 19400 -4665
rect 15850 -4970 16950 -4965
rect 15850 -5010 15855 -4970
rect 15895 -5010 16205 -4970
rect 16245 -5010 16555 -4970
rect 16595 -5010 16905 -4970
rect 16945 -5010 16950 -4970
rect 15850 -5015 16950 -5010
rect 17250 -4970 18350 -4965
rect 17250 -5010 17255 -4970
rect 17295 -5010 17605 -4970
rect 17645 -5010 17955 -4970
rect 17995 -5010 18305 -4970
rect 18345 -5010 18350 -4970
rect 17250 -5015 18350 -5010
rect 18650 -4970 19750 -4965
rect 18650 -5010 18655 -4970
rect 18695 -5010 19005 -4970
rect 19045 -5010 19355 -4970
rect 19395 -5010 19705 -4970
rect 19745 -5010 19750 -4970
rect 18650 -5015 19750 -5010
rect 16200 -5315 16250 -5015
rect 17950 -5315 18000 -5015
rect 19350 -5315 19400 -5015
rect 15850 -5320 16950 -5315
rect 15850 -5360 15855 -5320
rect 15895 -5360 16205 -5320
rect 16245 -5360 16555 -5320
rect 16595 -5360 16905 -5320
rect 16945 -5360 16950 -5320
rect 15850 -5365 16950 -5360
rect 17250 -5320 18350 -5315
rect 17250 -5360 17255 -5320
rect 17295 -5360 17605 -5320
rect 17645 -5360 17955 -5320
rect 17995 -5360 18305 -5320
rect 18345 -5360 18350 -5320
rect 17250 -5365 18350 -5360
rect 18650 -5320 19750 -5315
rect 18650 -5360 18655 -5320
rect 18695 -5360 19005 -5320
rect 19045 -5360 19355 -5320
rect 19395 -5360 19705 -5320
rect 19745 -5360 19750 -5320
rect 18650 -5365 19750 -5360
rect 16200 -5665 16250 -5365
rect 17950 -5665 18000 -5365
rect 19350 -5665 19400 -5365
rect 15850 -5670 16950 -5665
rect 15850 -5710 15855 -5670
rect 15895 -5710 16205 -5670
rect 16245 -5710 16555 -5670
rect 16595 -5710 16905 -5670
rect 16945 -5710 16950 -5670
rect 15850 -5715 16950 -5710
rect 17250 -5670 18350 -5665
rect 17250 -5710 17255 -5670
rect 17295 -5710 17605 -5670
rect 17645 -5710 17955 -5670
rect 17995 -5710 18305 -5670
rect 18345 -5710 18350 -5670
rect 17250 -5715 18350 -5710
rect 18650 -5670 19750 -5665
rect 18650 -5710 18655 -5670
rect 18695 -5710 19005 -5670
rect 19045 -5710 19355 -5670
rect 19395 -5710 19705 -5670
rect 19745 -5710 19750 -5670
rect 18650 -5715 19750 -5710
rect 16200 -6015 16250 -5715
rect 17950 -6015 18000 -5715
rect 19350 -6015 19400 -5715
rect 15850 -6020 16950 -6015
rect 15850 -6060 15855 -6020
rect 15895 -6060 16205 -6020
rect 16245 -6060 16555 -6020
rect 16595 -6060 16905 -6020
rect 16945 -6060 16950 -6020
rect 15850 -6065 16950 -6060
rect 17250 -6020 18350 -6015
rect 17250 -6060 17255 -6020
rect 17295 -6060 17605 -6020
rect 17645 -6060 17955 -6020
rect 17995 -6060 18305 -6020
rect 18345 -6060 18350 -6020
rect 17250 -6065 18350 -6060
rect 18650 -6020 19750 -6015
rect 18650 -6060 18655 -6020
rect 18695 -6060 19005 -6020
rect 19045 -6060 19355 -6020
rect 19395 -6060 19705 -6020
rect 19745 -6060 19750 -6020
rect 18650 -6065 19750 -6060
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_8 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 18145 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_18
timestamp 1723858470
transform 1 0 16785 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_19
timestamp 1723858470
transform 1 0 17465 0 1 -2775
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_20
timestamp 1723858470
transform 1 0 18145 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_21
timestamp 1723858470
transform 1 0 18145 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_22
timestamp 1723858470
transform 1 0 17465 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23
timestamp 1723858470
transform 1 0 17465 0 1 -3455
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_24
timestamp 1723858470
transform 1 0 16785 0 1 -4135
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25
timestamp 1723858470
transform 1 0 16785 0 1 -3455
box 0 0 670 670
<< labels >>
flabel metal2 15995 -4385 15995 -4385 5 FreeSans 400 0 0 -40 cap_res1
flabel metal3 19355 -4375 19355 -4375 7 FreeSans 400 180 -40 0 cap_res2
flabel metal1 18780 -1155 18780 -1155 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal1 16170 -1295 16170 -1295 7 FreeSans 400 0 -160 0 NFET_GATE_10uA
flabel metal1 16235 -955 16235 -955 3 FreeSans 400 0 200 0 START_UP
flabel poly 18430 600 18430 600 5 FreeSans 400 0 0 -40 V_TOP
flabel metal1 16040 1745 16040 1745 7 FreeSans 240 0 -160 0 VB2_CUR_BIAS
port 11 w
flabel metal1 19415 1750 19415 1750 7 FreeSans 240 0 -160 0 ERR_AMP_REF
port 2 w
flabel metal1 19565 1750 19565 1750 3 FreeSans 240 0 160 0 VB3_CUR_BIAS
port 8 e
flabel via1 17800 1615 17800 1615 1 FreeSans 400 0 0 200 PFET_GATE_10uA
flabel metal2 18580 -585 18580 -585 3 FreeSans 400 180 200 0 V_p_2
flabel metal2 17060 -585 17060 -585 3 FreeSans 400 0 200 0 V_p_1
flabel metal2 16670 -475 16670 -475 1 FreeSans 400 0 0 80 Vin+
flabel metal2 16665 -175 16665 -175 5 FreeSans 400 0 0 -80 Vin-
flabel metal2 18930 -475 18930 -475 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal2 17570 -110 17570 -110 3 FreeSans 240 0 120 0 1st_Vout_1
flabel metal2 16620 -70 16620 -70 5 FreeSans 400 0 0 -40 V_mir1
flabel metal2 18030 -110 18030 -110 7 FreeSans 240 0 -120 0 1st_Vout_2
flabel metal2 18980 -70 18980 -70 5 FreeSans 400 0 0 -40 V_mir2
flabel metal1 15805 1755 15805 1755 1 FreeSans 240 0 0 80 V_CMFB_S2
port 10 n
flabel metal1 17750 1755 17750 1755 1 FreeSans 240 0 0 80 TAIL_CUR_MIR_BIAS
port 5 n
flabel metal1 19795 1755 19795 1755 1 FreeSans 240 0 0 80 V_CMFB_S4
port 9 n
flabel metal1 16125 1755 16125 1755 1 FreeSans 240 0 0 80 ERR_AMP_CUR_BIAS
port 7 n
flabel metal1 19280 1750 19280 1750 1 FreeSans 240 0 0 80 VB1_CUR_BIAS
port 4 n
flabel metal1 18640 1755 18640 1755 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal1 16960 1755 16960 1755 1 FreeSans 240 0 0 80 V_CMFB_S1
port 6 n
<< end >>
