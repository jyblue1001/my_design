magic
tech sky130A
timestamp 1738592334
<< psubdiff >>
rect 2570 160 2670 175
rect 2570 140 2585 160
rect 2655 140 2670 160
rect 2570 125 2670 140
<< psubdiffcont >>
rect 2585 140 2655 160
<< xpolycontact >>
rect 3020 250 3240 285
rect 3976 250 4196 285
<< xpolyres >>
rect 3240 250 3976 285
<< locali >>
rect 2900 270 2920 445
rect 1150 250 3020 270
rect 4196 250 4405 270
rect 1150 230 1170 250
rect 4385 230 4405 250
rect 1130 220 1180 230
rect 1130 190 1140 220
rect 1170 190 1180 220
rect 1130 180 1180 190
rect 2475 220 2780 230
rect 2475 185 2485 220
rect 2520 210 2610 220
rect 2520 185 2530 210
rect 2600 200 2610 210
rect 2630 210 2735 220
rect 2630 200 2640 210
rect 2600 190 2640 200
rect 2475 175 2530 185
rect 2725 185 2735 210
rect 2770 185 2780 220
rect 2725 175 2780 185
rect 4375 220 4425 230
rect 4375 190 4385 220
rect 4415 190 4425 220
rect 4375 180 4425 190
rect 2575 160 2665 170
rect 2575 140 2585 160
rect 2655 140 2665 160
rect 2575 130 2665 140
<< viali >>
rect 1140 190 1170 220
rect 2485 185 2520 220
rect 2610 200 2630 220
rect 2735 185 2770 220
rect 4385 190 4415 220
rect 2585 140 2655 160
<< metal1 >>
rect 1130 220 1180 230
rect 1130 190 1140 220
rect 1170 190 1180 220
rect 1130 180 1180 190
rect 2475 220 2530 230
rect 2475 185 2485 220
rect 2520 185 2530 220
rect 2475 175 2530 185
rect 2570 220 2670 230
rect 2570 200 2610 220
rect 2630 200 2670 220
rect 2570 160 2670 200
rect 2725 220 2780 230
rect 2725 185 2735 220
rect 2770 185 2780 220
rect 2725 175 2780 185
rect 4375 220 4425 230
rect 4375 190 4385 220
rect 4415 190 4425 220
rect 4375 180 4425 190
rect 2570 140 2585 160
rect 2655 140 2670 160
rect 2570 125 2670 140
<< via1 >>
rect 1140 190 1170 220
rect 2485 185 2520 220
rect 2735 185 2770 220
rect 4385 190 4415 220
<< metal2 >>
rect 1130 220 1180 230
rect 1130 190 1140 220
rect 1170 190 1180 220
rect 1130 180 1180 190
rect 2475 220 2530 230
rect 2475 185 2485 220
rect 2520 185 2530 220
rect 2475 175 2530 185
rect 2725 220 2780 230
rect 2725 185 2735 220
rect 2770 185 2780 220
rect 2725 175 2780 185
rect 4375 220 4425 230
rect 4375 190 4385 220
rect 4415 190 4425 220
rect 4375 180 4425 190
<< via2 >>
rect 1140 190 1170 220
rect 2485 185 2520 220
rect 2735 185 2770 220
rect 4385 190 4415 220
<< metal3 >>
rect 1130 220 1180 230
rect 1130 190 1140 220
rect 1170 190 1180 220
rect 1130 180 1180 190
rect 1135 55 1180 180
rect 2475 220 2530 230
rect 2475 185 2485 220
rect 2520 185 2530 220
rect 2475 175 2530 185
rect 2725 220 2780 230
rect 2725 185 2735 220
rect 2770 185 2780 220
rect 2725 175 2780 185
rect 4375 220 4425 230
rect 4375 190 4385 220
rect 4415 190 4425 220
rect 4375 180 4425 190
rect 4375 55 4420 180
rect 1135 -5975 2545 55
rect 2710 -5975 9720 55
<< via3 >>
rect 2485 185 2520 220
rect 2735 185 2770 220
<< mimcap >>
rect 1150 30 2530 40
rect 1150 -5 2485 30
rect 2520 -5 2530 30
rect 1150 -5960 2530 -5
rect 2725 30 9705 40
rect 2725 -5 2735 30
rect 2770 -5 9705 30
rect 2725 -5960 9705 -5
<< mimcapcontact >>
rect 2485 -5 2520 30
rect 2735 -5 2770 30
<< metal4 >>
rect 2475 220 2530 230
rect 2475 185 2485 220
rect 2520 185 2530 220
rect 2475 30 2530 185
rect 2475 -5 2485 30
rect 2520 -5 2530 30
rect 2475 -10 2530 -5
rect 2725 220 2780 230
rect 2725 185 2735 220
rect 2770 185 2780 220
rect 2725 30 2780 185
rect 2725 -5 2735 30
rect 2770 -5 2780 30
rect 2725 -10 2780 -5
<< labels >>
flabel locali 2920 445 2920 445 2 FreeSans 800 0 400 400 V_OUT
port 1 ne
flabel metal1 2620 190 2620 190 5 FreeSans 800 0 0 -400 GNDA
port 2 s
<< end >>
