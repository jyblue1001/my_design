* PEX produced on Thu Feb 20 06:38:54 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from VCO_FD_magic.ext - technology: sky130A

.subckt VCO_FD_magic V_OUT_120 VDDA GNDA V_CONT
X0 vco2_3_0.V4.t2 GNDA.t118 VDDA.t77 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X1 GNDA.t76 div120_2_0.div3_3_0.CLK.t3 div120_2_0.div3_3_0.H.t2 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X2 div120_2_0.div5_2_0.F.t1 div120_2_0.div5_2_0.E.t2 VDDA.t52 VDDA.t51 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X3 GNDA.t94 div120_2_0.div3_3_0.I.t2 div120_2_0.div3_3_0.G.t1 GNDA.t93 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X4 div120_2_0.div3_3_0.I.t0 div120_2_0.div3_3_0.CLK.t4 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X5 div120_2_0.div2.t1 a_2510_770.t3 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X6 div120_2_0.div2_4_0.C.t3 a_5110_770.t3 GNDA.t54 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X7 div120_2_0.div4.t1 div120_2_0.div2_4_2.C.t4 GNDA.t84 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X8 div120_2_0.div5_2_0.I.t2 div120_2_0.div5_2_0.Q2_b.t2 div120_2_0.div5_2_0.H.t1 GNDA.t107 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X9 vco2_3_0.V3.t1 vco2_3_0.V8.t2 V_OSC.t0 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.2
X10 VDDA.t37 div120_2_0.div8.t2 div120_2_0.div3_3_0.CLK.t1 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X11 GNDA.t74 div120_2_0.div3_3_0.CLK.t5 div120_2_0.div3_3_0.C.t2 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X12 a_5110_770.t0 div120_2_0.div4.t2 VDDA.t6 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X13 GNDA.t72 div120_2_0.div3_3_0.CLK.t6 div120_2_0.div3_3_0.H.t1 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X14 div120_2_0.div3_3_0.A.t1 div120_2_0.div3_3_0.CLK.t7 div120_2_0.div3_3_0.B.t1 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X15 GNDA.t38 div120_2_0.div4.t3 a_5110_770.t2 GNDA.t37 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X16 VDDA.t71 div120_2_0.div8.t3 div120_2_0.div2_4_0.A.t0 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X17 div120_2_0.div3_3_0.F.t1 div120_2_0.div3_3_0.CLK.t8 div120_2_0.div3_3_0.E.t0 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X18 div120_2_0.div5_2_0.A.t0 div120_2_0.div5_2_0.Q2_b.t3 GNDA.t43 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X19 div120_2_0.div5_2_0.M.t0 div120_2_0.div5_2_0.K.t2 VDDA.t35 VDDA.t34 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X20 div120_2_0.div5_2_0.K.t1 div120_2_0.div5_2_0.Q2_b.t4 div120_2_0.div5_2_0.L.t0 GNDA.t41 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X21 VDDA.t41 div120_2_0.div5_2_0.G.t3 div120_2_0.div5_2_0.J.t0 VDDA.t40 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X22 VDDA.t58 div120_2_0.div3_3_0.I.t3 div120_2_0.div24.t2 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X23 vco2_3_0.V2.t1 vco2_3_0.V8.t3 V_OSC.t1 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.2
X24 GNDA.t1 div120_2_0.div5_2_0.Q2_b.t5 div120_2_0.div5_2_0.M.t3 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X25 div120_2_0.div2_4_2.C.t2 a_3810_770.t3 GNDA.t80 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X26 VDDA.t85 V_OSC.t2 a_2510_770.t2 VDDA.t84 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X27 GNDA.t58 div120_2_0.div24.t3 div120_2_0.div5_2_0.J.t3 GNDA.t57 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X28 GNDA.t68 div120_2_0.div3_3_0.CLK.t9 div120_2_0.div3_3_0.C.t1 GNDA.t67 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X29 div120_2_0.div2.t0 div120_2_0.div2_4_1.C.t4 GNDA.t82 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X30 div120_2_0.div2_4_1.C.t0 div120_2_0.div2_4_1.A.t2 VDDA.t24 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X31 div120_2_0.div4.t0 a_3810_770.t4 VDDA.t32 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X32 VDDA.t22 vco2_3_0.V1.t1 vco2_3_0.V1.t2 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X33 div120_2_0.div2_4_0.A.t1 a_5110_770.t4 div120_2_0.div2_4_0.B.t1 GNDA.t110 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X34 div120_2_0.div5_2_0.D.t0 div120_2_0.div5_2_0.B.t2 VDDA.t83 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X35 div120_2_0.div3_3_0.CLK.t2 div120_2_0.div8.t4 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X36 GNDA.t3 div120_2_0.div5_2_0.Q2_b.t6 div120_2_0.div5_2_0.M.t2 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X37 GNDA.t52 div120_2_0.div24.t4 div120_2_0.div5_2_0.J.t2 GNDA.t51 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X38 VDDA.t12 div120_2_0.div24.t5 div120_2_0.div3_3_0.A.t0 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X39 div120_2_0.div2_4_1.C.t3 a_2510_770.t4 GNDA.t12 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X40 vco2_3_0.V7.t0 V_OSC.t3 vco2_3_0.V9.t0 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.2
X41 div120_2_0.div2_4_1.B.t0 div120_2_0.div2.t2 GNDA.t32 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X42 GNDA.t47 div120_2_0.div24.t6 div120_2_0.div5_2_0.D.t3 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X43 vco2_3_0.V4.t1 vco2_3_0.V1.t3 VDDA.t63 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X44 div120_2_0.div5_2_0.B.t0 div120_2_0.div24.t7 div120_2_0.div5_2_0.C.t0 GNDA.t104 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X45 VDDA.t30 div120_2_0.div2.t3 a_3810_770.t2 VDDA.t29 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X46 vco2_3_0.V5.t1 vco2_3_0.V9.t2 vco2_3_0.V8.t0 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.2
X47 div120_2_0.div2_4_2.C.t3 div120_2_0.div2_4_2.A.t2 VDDA.t67 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X48 a_2510_770.t0 V_OSC.t4 VDDA.t28 VDDA.t27 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X49 div120_2_0.div2_4_2.A.t0 a_3810_770.t5 div120_2_0.div2_4_2.B.t0 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X50 VDDA.t87 div120_2_0.div3_3_0.D.t2 div120_2_0.div3_3_0.E.t2 VDDA.t86 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X51 VDDA.t46 div120_2_0.div2.t4 div120_2_0.div2_4_1.A.t0 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X52 div120_2_0.div3_3_0.I.t1 div120_2_0.div3_3_0.H.t4 GNDA.t86 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X53 GNDA.t56 div120_2_0.div24.t8 div120_2_0.div5_2_0.D.t2 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X54 vco2_3_0.V2.t2 GNDA.t119 VDDA.t75 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X55 GNDA.t34 a_5110_770.t5 div120_2_0.div2_4_0.C.t2 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X56 GNDA.t14 div120_2_0.div2.t5 a_3810_770.t0 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X57 vco2_3_0.V3.t0 V_CONT.t0 GNDA.t45 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X58 VDDA.t1 div120_2_0.div5_2_0.Q2_b.t7 div120_2_0.div5_2_0.A.t2 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X59 div120_2_0.div3_3_0.D.t0 div120_2_0.div3_3_0.C.t4 GNDA.t117 GNDA.t116 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X60 div120_2_0.div3_3_0.H.t0 div120_2_0.div3_3_0.CLK.t10 GNDA.t66 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X61 vco2_3_0.V6.t0 V_OSC.t5 vco2_3_0.V9.t1 VDDA.t59 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.2
X62 div120_2_0.div3_3_0.G.t0 div120_2_0.div3_3_0.D.t3 div120_2_0.div3_3_0.F.t0 GNDA.t28 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X63 VDDA.t89 div120_2_0.div3_3_0.E.t3 div120_2_0.div3_3_0.H.t3 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X64 div120_2_0.div2_4_0.C.t0 div120_2_0.div2_4_0.A.t2 VDDA.t39 VDDA.t38 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X65 V_OUT_120.t1 div120_2_0.div5_2_0.Q2_b.t8 VDDA.t81 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X66 GNDA.t16 a_5110_770.t6 div120_2_0.div2_4_0.C.t1 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X67 GNDA.t60 a_3810_770.t6 div120_2_0.div2_4_2.C.t0 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X68 div120_2_0.div5_2_0.H.t0 div120_2_0.div24.t9 div120_2_0.div5_2_0.G.t0 GNDA.t23 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X69 div120_2_0.div5_2_0.Q2_b.t0 div120_2_0.div24.t10 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X70 div120_2_0.div5_2_0.Q2_b.t1 div120_2_0.div5_2_0.J.t4 GNDA.t10 GNDA.t9 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X71 GNDA.t40 V_CONT.t1 vco2_3_0.V1.t0 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X72 div120_2_0.div3_3_0.C.t0 div120_2_0.div3_3_0.CLK.t11 GNDA.t64 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X73 GNDA.t88 V_OSC.t6 a_2510_770.t1 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X74 vco2_3_0.V3.t2 VDDA.t94 GNDA.t48 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X75 div120_2_0.div3_3_0.B.t0 div120_2_0.div24.t11 GNDA.t22 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X76 div120_2_0.div8.t0 div120_2_0.div2_4_0.C.t4 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X77 vco2_3_0.V4.t0 vco2_3_0.V9.t3 vco2_3_0.V8.t1 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.2
X78 VDDA.t26 V_OUT_120.t2 div120_2_0.div5_2_0.K.t0 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X79 div120_2_0.div24.t1 div120_2_0.div3_3_0.I.t4 VDDA.t56 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X80 div120_2_0.div5_2_0.L.t1 V_OUT_120.t3 GNDA.t106 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X81 div120_2_0.div5_2_0.M.t1 div120_2_0.div5_2_0.Q2_b.t9 GNDA.t103 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X82 GNDA.t78 a_3810_770.t7 div120_2_0.div2_4_2.C.t1 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X83 div120_2_0.div5_2_0.A.t1 div120_2_0.div5_2_0.Q2_b.t10 VDDA.t79 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X84 div120_2_0.div8.t1 a_5110_770.t7 VDDA.t16 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X85 div120_2_0.div5_2_0.J.t1 div120_2_0.div24.t12 GNDA.t8 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X86 vco2_3_0.V7.t1 V_CONT.t2 GNDA.t101 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X87 div120_2_0.div3_3_0.C.t3 div120_2_0.div3_3_0.A.t2 VDDA.t93 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X88 GNDA.t92 a_2510_770.t5 div120_2_0.div2_4_1.C.t2 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X89 GNDA.t90 div120_2_0.div5_2_0.E.t3 div120_2_0.div5_2_0.I.t1 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X90 div120_2_0.div2_4_1.A.t1 a_2510_770.t6 div120_2_0.div2_4_1.B.t1 GNDA.t99 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X91 div120_2_0.div5_2_0.G.t1 V_OUT_120.t4 div120_2_0.div5_2_0.F.t0 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X92 VDDA.t61 div120_2_0.div5_2_0.Q2_b.t11 div120_2_0.div5_2_0.G.t2 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X93 vco2_3_0.V5.t0 V_CONT.t3 GNDA.t27 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X94 div120_2_0.div5_2_0.E.t0 div120_2_0.div5_2_0.D.t4 GNDA.t50 GNDA.t49 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X95 VDDA.t91 div120_2_0.div5_2_0.A.t3 div120_2_0.div5_2_0.B.t1 VDDA.t90 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X96 div120_2_0.div24.t0 div120_2_0.div3_3_0.I.t5 GNDA.t62 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X97 div120_2_0.div2_4_0.B.t0 div120_2_0.div8.t5 GNDA.t109 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X98 vco2_3_0.V2.t0 vco2_3_0.V1.t4 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X99 div120_2_0.div5_2_0.E.t1 div120_2_0.div24.t13 VDDA.t65 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X100 div120_2_0.div3_3_0.E.t1 div120_2_0.div3_3_0.I.t6 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X101 vco2_3_0.V6.t2 GNDA.t120 VDDA.t73 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X102 GNDA.t98 a_2510_770.t7 div120_2_0.div2_4_1.C.t1 GNDA.t97 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X103 V_OUT_120.t0 div120_2_0.div5_2_0.M.t4 GNDA.t20 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X104 VDDA.t18 div120_2_0.div4.t4 a_5110_770.t1 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X105 vco2_3_0.V6.t1 vco2_3_0.V1.t5 VDDA.t44 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=1.5
X106 vco2_3_0.V7.t2 VDDA.t95 GNDA.t111 GNDA.t100 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X107 div120_2_0.div5_2_0.D.t1 div120_2_0.div24.t14 GNDA.t96 GNDA.t95 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X108 a_3810_770.t1 div120_2_0.div2.t6 VDDA.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
X109 div120_2_0.div5_2_0.C.t1 div120_2_0.div5_2_0.A.t4 GNDA.t114 GNDA.t113 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X110 div120_2_0.div3_3_0.D.t1 div120_2_0.div3_3_0.CLK.t12 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X111 VDDA.t4 div120_2_0.div4.t5 div120_2_0.div2_4_2.A.t1 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X112 vco2_3_0.V5.t2 VDDA.t96 GNDA.t112 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.2 ps=1.8 w=0.5 l=0.15
X113 div120_2_0.div2_4_2.B.t1 div120_2_0.div4.t6 GNDA.t18 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.15
X114 GNDA.t6 div120_2_0.div8.t6 div120_2_0.div3_3_0.CLK.t0 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.15
X115 div120_2_0.div5_2_0.I.t0 V_OUT_120.t5 GNDA.t30 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.15
R0 GNDA.n274 GNDA.t26 2223.91
R1 GNDA.n273 GNDA.t44 2223.91
R2 GNDA.t100 GNDA.t87 2124.71
R3 GNDA.t42 GNDA.t61 1552.94
R4 GNDA.t49 GNDA.t23 1509.8
R5 GNDA.t9 GNDA.t105 1466.67
R6 GNDA.t29 GNDA.t51 1423.53
R7 GNDA.t69 GNDA.t116 1423.53
R8 GNDA.t67 GNDA.t70 1423.53
R9 GNDA.t15 GNDA.t110 1423.53
R10 GNDA.t77 GNDA.t24 1423.53
R11 GNDA.t99 GNDA.t97 1423.53
R12 GNDA.n55 GNDA.t42 1358.82
R13 GNDA.n211 GNDA.n22 1204.13
R14 GNDA.n53 GNDA.n31 1204.13
R15 GNDA.n260 GNDA.n259 1204.13
R16 GNDA.n54 GNDA.n43 1182.8
R17 GNDA.n56 GNDA.n55 1182.8
R18 GNDA.n268 GNDA.n267 1173.78
R19 GNDA.n273 GNDA.n272 1173.78
R20 GNDA.n275 GNDA.n274 1173.78
R21 GNDA.t41 GNDA.t2 1078.43
R22 GNDA.t104 GNDA.t55 1078.43
R23 GNDA.t61 GNDA.t85 1078.43
R24 GNDA.t5 GNDA.n53 970.588
R25 GNDA.t37 GNDA.n22 970.588
R26 GNDA.n260 GNDA.t13 970.588
R27 GNDA.t71 GNDA.n54 841.178
R28 GNDA.n53 GNDA.t35 841.178
R29 GNDA.n22 GNDA.t83 841.178
R30 GNDA.t81 GNDA.n260 841.178
R31 GNDA.n267 GNDA.t119 728.524
R32 GNDA.n272 GNDA.t118 728.524
R33 GNDA.n275 GNDA.t120 728.524
R34 GNDA.n265 GNDA.n262 686.717
R35 GNDA.n270 GNDA.n261 686.717
R36 GNDA.n278 GNDA.n277 686.717
R37 GNDA.n279 GNDA.n278 686.717
R38 GNDA.n261 GNDA.n4 686.717
R39 GNDA.n263 GNDA.n262 686.717
R40 GNDA.n268 GNDA.t39 645.653
R41 GNDA.n274 GNDA.t115 621.74
R42 GNDA.t25 GNDA.n273 621.74
R43 GNDA.t4 GNDA.n268 621.74
R44 GNDA.n55 GNDA.t113 582.354
R45 GNDA.n54 GNDA.t93 582.354
R46 GNDA.t0 GNDA.t19 474.51
R47 GNDA.t102 GNDA.t0 474.51
R48 GNDA.t2 GNDA.t102 474.51
R49 GNDA.t105 GNDA.t41 474.51
R50 GNDA.t57 GNDA.t9 474.51
R51 GNDA.t7 GNDA.t57 474.51
R52 GNDA.t51 GNDA.t7 474.51
R53 GNDA.t89 GNDA.t29 474.51
R54 GNDA.t107 GNDA.t89 474.51
R55 GNDA.t23 GNDA.t107 474.51
R56 GNDA.t46 GNDA.t49 474.51
R57 GNDA.t95 GNDA.t46 474.51
R58 GNDA.t55 GNDA.t95 474.51
R59 GNDA.t113 GNDA.t104 474.51
R60 GNDA.t85 GNDA.t75 474.51
R61 GNDA.t75 GNDA.t65 474.51
R62 GNDA.t65 GNDA.t71 474.51
R63 GNDA.t93 GNDA.t28 474.51
R64 GNDA.t28 GNDA.t69 474.51
R65 GNDA.t116 GNDA.t73 474.51
R66 GNDA.t73 GNDA.t63 474.51
R67 GNDA.t63 GNDA.t67 474.51
R68 GNDA.t70 GNDA.t21 474.51
R69 GNDA.t21 GNDA.t5 474.51
R70 GNDA.t35 GNDA.t33 474.51
R71 GNDA.t33 GNDA.t53 474.51
R72 GNDA.t53 GNDA.t15 474.51
R73 GNDA.t110 GNDA.t108 474.51
R74 GNDA.t108 GNDA.t37 474.51
R75 GNDA.t83 GNDA.t59 474.51
R76 GNDA.t59 GNDA.t79 474.51
R77 GNDA.t79 GNDA.t77 474.51
R78 GNDA.t24 GNDA.t17 474.51
R79 GNDA.t17 GNDA.t13 474.51
R80 GNDA.t91 GNDA.t81 474.51
R81 GNDA.t11 GNDA.t91 474.51
R82 GNDA.t97 GNDA.t11 474.51
R83 GNDA.t31 GNDA.t99 474.51
R84 GNDA.t87 GNDA.t31 474.51
R85 GNDA.n84 GNDA.t106 295.933
R86 GNDA.n134 GNDA.t43 295.933
R87 GNDA.n141 GNDA.t62 295.933
R88 GNDA.n265 GNDA.t40 260
R89 GNDA.n263 GNDA.t40 260
R90 GNDA.n76 GNDA.n75 256.207
R91 GNDA.n77 GNDA.n74 247.934
R92 GNDA.n91 GNDA.n69 247.934
R93 GNDA.n94 GNDA.n93 247.934
R94 GNDA.n65 GNDA.n64 247.934
R95 GNDA.n113 GNDA.n112 247.934
R96 GNDA.n119 GNDA.n59 247.934
R97 GNDA.n147 GNDA.n46 247.934
R98 GNDA.n150 GNDA.n149 247.934
R99 GNDA.n169 GNDA.n38 247.934
R100 GNDA.n172 GNDA.n171 247.934
R101 GNDA.n184 GNDA.n33 246.714
R102 GNDA.n278 GNDA.n274 241.643
R103 GNDA.n273 GNDA.n261 241.643
R104 GNDA.n268 GNDA.n262 241.643
R105 GNDA.n43 GNDA.t94 233
R106 GNDA.n56 GNDA.t114 233
R107 GNDA.n266 GNDA.t48 233
R108 GNDA.n271 GNDA.t112 233
R109 GNDA.n276 GNDA.t111 233
R110 GNDA.n29 GNDA.n28 219.133
R111 GNDA.n196 GNDA.n27 219.133
R112 GNDA.n204 GNDA.n203 219.133
R113 GNDA.n217 GNDA.n19 219.133
R114 GNDA.n17 GNDA.n16 219.133
R115 GNDA.n229 GNDA.n13 219.133
R116 GNDA.n253 GNDA.n235 219.133
R117 GNDA.n237 GNDA.n236 219.133
R118 GNDA.n241 GNDA.n240 219.133
R119 GNDA.n264 GNDA.t45 128.562
R120 GNDA.n269 GNDA.t27 127.754
R121 GNDA.n9 GNDA.t101 127.754
R122 GNDA.n157 GNDA.n43 54.4005
R123 GNDA.n127 GNDA.n56 54.4005
R124 GNDA.n75 GNDA.t20 48.0005
R125 GNDA.n75 GNDA.t1 48.0005
R126 GNDA.n74 GNDA.t103 48.0005
R127 GNDA.n74 GNDA.t3 48.0005
R128 GNDA.n69 GNDA.t10 48.0005
R129 GNDA.n69 GNDA.t58 48.0005
R130 GNDA.n93 GNDA.t8 48.0005
R131 GNDA.n93 GNDA.t52 48.0005
R132 GNDA.n64 GNDA.t30 48.0005
R133 GNDA.n64 GNDA.t90 48.0005
R134 GNDA.n112 GNDA.t50 48.0005
R135 GNDA.n112 GNDA.t47 48.0005
R136 GNDA.n59 GNDA.t96 48.0005
R137 GNDA.n59 GNDA.t56 48.0005
R138 GNDA.n46 GNDA.t86 48.0005
R139 GNDA.n46 GNDA.t76 48.0005
R140 GNDA.n149 GNDA.t66 48.0005
R141 GNDA.n149 GNDA.t72 48.0005
R142 GNDA.n38 GNDA.t117 48.0005
R143 GNDA.n38 GNDA.t74 48.0005
R144 GNDA.n171 GNDA.t64 48.0005
R145 GNDA.n171 GNDA.t68 48.0005
R146 GNDA.n33 GNDA.t22 48.0005
R147 GNDA.n33 GNDA.t6 48.0005
R148 GNDA.n28 GNDA.t36 48.0005
R149 GNDA.n28 GNDA.t34 48.0005
R150 GNDA.n27 GNDA.t54 48.0005
R151 GNDA.n27 GNDA.t16 48.0005
R152 GNDA.n203 GNDA.t109 48.0005
R153 GNDA.n203 GNDA.t38 48.0005
R154 GNDA.n19 GNDA.t84 48.0005
R155 GNDA.n19 GNDA.t60 48.0005
R156 GNDA.n16 GNDA.t80 48.0005
R157 GNDA.n16 GNDA.t78 48.0005
R158 GNDA.n13 GNDA.t18 48.0005
R159 GNDA.n13 GNDA.t14 48.0005
R160 GNDA.n235 GNDA.t82 48.0005
R161 GNDA.n235 GNDA.t92 48.0005
R162 GNDA.n236 GNDA.t12 48.0005
R163 GNDA.n236 GNDA.t98 48.0005
R164 GNDA.n240 GNDA.t32 48.0005
R165 GNDA.n240 GNDA.t88 48.0005
R166 GNDA.n271 GNDA.n270 35.6576
R167 GNDA.n290 GNDA.n4 35.6576
R168 GNDA.n277 GNDA.n276 35.6576
R169 GNDA.n280 GNDA.n279 35.6576
R170 GNDA.n266 GNDA.n265 34.3278
R171 GNDA.n263 GNDA.n0 34.3278
R172 GNDA.n292 GNDA.n291 32.0005
R173 GNDA.n292 GNDA.n2 32.0005
R174 GNDA.n296 GNDA.n2 32.0005
R175 GNDA.n297 GNDA.n296 32.0005
R176 GNDA.n298 GNDA.n297 32.0005
R177 GNDA.n284 GNDA.n7 32.0005
R178 GNDA.n285 GNDA.n284 32.0005
R179 GNDA.n286 GNDA.n285 32.0005
R180 GNDA.n286 GNDA.n5 32.0005
R181 GNDA.n290 GNDA.n5 32.0005
R182 GNDA.n79 GNDA.n78 32.0005
R183 GNDA.n79 GNDA.n72 32.0005
R184 GNDA.n83 GNDA.n72 32.0005
R185 GNDA.n86 GNDA.n85 32.0005
R186 GNDA.n86 GNDA.n70 32.0005
R187 GNDA.n90 GNDA.n70 32.0005
R188 GNDA.n95 GNDA.n92 32.0005
R189 GNDA.n99 GNDA.n67 32.0005
R190 GNDA.n100 GNDA.n99 32.0005
R191 GNDA.n101 GNDA.n100 32.0005
R192 GNDA.n105 GNDA.n104 32.0005
R193 GNDA.n106 GNDA.n105 32.0005
R194 GNDA.n106 GNDA.n62 32.0005
R195 GNDA.n110 GNDA.n62 32.0005
R196 GNDA.n111 GNDA.n110 32.0005
R197 GNDA.n114 GNDA.n111 32.0005
R198 GNDA.n118 GNDA.n60 32.0005
R199 GNDA.n121 GNDA.n120 32.0005
R200 GNDA.n121 GNDA.n57 32.0005
R201 GNDA.n125 GNDA.n57 32.0005
R202 GNDA.n126 GNDA.n125 32.0005
R203 GNDA.n128 GNDA.n51 32.0005
R204 GNDA.n132 GNDA.n51 32.0005
R205 GNDA.n133 GNDA.n132 32.0005
R206 GNDA.n135 GNDA.n133 32.0005
R207 GNDA.n139 GNDA.n49 32.0005
R208 GNDA.n140 GNDA.n139 32.0005
R209 GNDA.n142 GNDA.n47 32.0005
R210 GNDA.n146 GNDA.n47 32.0005
R211 GNDA.n151 GNDA.n148 32.0005
R212 GNDA.n155 GNDA.n44 32.0005
R213 GNDA.n156 GNDA.n155 32.0005
R214 GNDA.n158 GNDA.n41 32.0005
R215 GNDA.n162 GNDA.n41 32.0005
R216 GNDA.n163 GNDA.n162 32.0005
R217 GNDA.n164 GNDA.n163 32.0005
R218 GNDA.n164 GNDA.n39 32.0005
R219 GNDA.n168 GNDA.n39 32.0005
R220 GNDA.n173 GNDA.n170 32.0005
R221 GNDA.n177 GNDA.n36 32.0005
R222 GNDA.n178 GNDA.n177 32.0005
R223 GNDA.n179 GNDA.n178 32.0005
R224 GNDA.n179 GNDA.n34 32.0005
R225 GNDA.n183 GNDA.n34 32.0005
R226 GNDA.n186 GNDA.n185 32.0005
R227 GNDA.n190 GNDA.n189 32.0005
R228 GNDA.n191 GNDA.n190 32.0005
R229 GNDA.n195 GNDA.n194 32.0005
R230 GNDA.n197 GNDA.n25 32.0005
R231 GNDA.n201 GNDA.n25 32.0005
R232 GNDA.n202 GNDA.n201 32.0005
R233 GNDA.n205 GNDA.n202 32.0005
R234 GNDA.n209 GNDA.n23 32.0005
R235 GNDA.n210 GNDA.n209 32.0005
R236 GNDA.n212 GNDA.n20 32.0005
R237 GNDA.n216 GNDA.n20 32.0005
R238 GNDA.n219 GNDA.n218 32.0005
R239 GNDA.n223 GNDA.n222 32.0005
R240 GNDA.n224 GNDA.n223 32.0005
R241 GNDA.n224 GNDA.n14 32.0005
R242 GNDA.n228 GNDA.n14 32.0005
R243 GNDA.n231 GNDA.n230 32.0005
R244 GNDA.n231 GNDA.n10 32.0005
R245 GNDA.n258 GNDA.n11 32.0005
R246 GNDA.n254 GNDA.n11 32.0005
R247 GNDA.n252 GNDA.n251 32.0005
R248 GNDA.n248 GNDA.n247 32.0005
R249 GNDA.n247 GNDA.n246 32.0005
R250 GNDA.n246 GNDA.n239 32.0005
R251 GNDA.n242 GNDA.n239 32.0005
R252 GNDA.n78 GNDA.n77 28.8005
R253 GNDA.n134 GNDA.n49 28.8005
R254 GNDA.n148 GNDA.n147 28.8005
R255 GNDA.n185 GNDA.n184 28.8005
R256 GNDA.n205 GNDA.n204 28.8005
R257 GNDA.n229 GNDA.n228 28.8005
R258 GNDA.n242 GNDA.n241 28.8005
R259 GNDA.n298 GNDA.n0 25.6005
R260 GNDA.n84 GNDA.n83 25.6005
R261 GNDA.n92 GNDA.n91 25.6005
R262 GNDA.n101 GNDA.n65 25.6005
R263 GNDA.n119 GNDA.n118 25.6005
R264 GNDA.n170 GNDA.n169 25.6005
R265 GNDA.n194 GNDA.n29 25.6005
R266 GNDA.n218 GNDA.n217 25.6005
R267 GNDA.n253 GNDA.n252 25.6005
R268 GNDA.t115 GNDA.t100 23.9135
R269 GNDA.t26 GNDA.t25 23.9135
R270 GNDA.t44 GNDA.t4 23.9135
R271 GNDA.n281 GNDA.n8 23.6001
R272 GNDA.n150 GNDA.n44 22.4005
R273 GNDA.n186 GNDA.n31 22.4005
R274 GNDA.n211 GNDA.n210 22.4005
R275 GNDA.n259 GNDA.n10 22.4005
R276 GNDA.n94 GNDA.n67 19.2005
R277 GNDA.n114 GNDA.n113 19.2005
R278 GNDA.n141 GNDA.n140 19.2005
R279 GNDA.n157 GNDA.n156 19.2005
R280 GNDA.n172 GNDA.n36 19.2005
R281 GNDA.n197 GNDA.n196 19.2005
R282 GNDA.n222 GNDA.n17 19.2005
R283 GNDA.n248 GNDA.n237 19.2005
R284 GNDA.n127 GNDA.n126 16.0005
R285 GNDA.n128 GNDA.n127 16.0005
R286 GNDA.n291 GNDA.n290 12.8005
R287 GNDA.n280 GNDA.n7 12.8005
R288 GNDA.n95 GNDA.n94 12.8005
R289 GNDA.n113 GNDA.n60 12.8005
R290 GNDA.n142 GNDA.n141 12.8005
R291 GNDA.n158 GNDA.n157 12.8005
R292 GNDA.n173 GNDA.n172 12.8005
R293 GNDA.n196 GNDA.n195 12.8005
R294 GNDA.n219 GNDA.n17 12.8005
R295 GNDA.n251 GNDA.n237 12.8005
R296 GNDA.n241 GNDA.n8 10.7016
R297 GNDA.n77 GNDA.n76 10.4505
R298 GNDA.n151 GNDA.n150 9.6005
R299 GNDA.n189 GNDA.n31 9.6005
R300 GNDA.n212 GNDA.n211 9.6005
R301 GNDA.n259 GNDA.n258 9.6005
R302 GNDA.n243 GNDA.n242 9.3005
R303 GNDA.n244 GNDA.n239 9.3005
R304 GNDA.n246 GNDA.n245 9.3005
R305 GNDA.n247 GNDA.n238 9.3005
R306 GNDA.n249 GNDA.n248 9.3005
R307 GNDA.n251 GNDA.n250 9.3005
R308 GNDA.n252 GNDA.n234 9.3005
R309 GNDA.n255 GNDA.n254 9.3005
R310 GNDA.n256 GNDA.n11 9.3005
R311 GNDA.n258 GNDA.n257 9.3005
R312 GNDA.n233 GNDA.n10 9.3005
R313 GNDA.n232 GNDA.n231 9.3005
R314 GNDA.n230 GNDA.n12 9.3005
R315 GNDA.n228 GNDA.n227 9.3005
R316 GNDA.n226 GNDA.n14 9.3005
R317 GNDA.n225 GNDA.n224 9.3005
R318 GNDA.n223 GNDA.n15 9.3005
R319 GNDA.n222 GNDA.n221 9.3005
R320 GNDA.n220 GNDA.n219 9.3005
R321 GNDA.n218 GNDA.n18 9.3005
R322 GNDA.n216 GNDA.n215 9.3005
R323 GNDA.n214 GNDA.n20 9.3005
R324 GNDA.n213 GNDA.n212 9.3005
R325 GNDA.n210 GNDA.n21 9.3005
R326 GNDA.n209 GNDA.n208 9.3005
R327 GNDA.n207 GNDA.n23 9.3005
R328 GNDA.n206 GNDA.n205 9.3005
R329 GNDA.n202 GNDA.n24 9.3005
R330 GNDA.n201 GNDA.n200 9.3005
R331 GNDA.n199 GNDA.n25 9.3005
R332 GNDA.n198 GNDA.n197 9.3005
R333 GNDA.n195 GNDA.n26 9.3005
R334 GNDA.n194 GNDA.n193 9.3005
R335 GNDA.n192 GNDA.n191 9.3005
R336 GNDA.n190 GNDA.n30 9.3005
R337 GNDA.n189 GNDA.n188 9.3005
R338 GNDA.n187 GNDA.n186 9.3005
R339 GNDA.n185 GNDA.n32 9.3005
R340 GNDA.n78 GNDA.n73 9.3005
R341 GNDA.n80 GNDA.n79 9.3005
R342 GNDA.n81 GNDA.n72 9.3005
R343 GNDA.n83 GNDA.n82 9.3005
R344 GNDA.n85 GNDA.n71 9.3005
R345 GNDA.n87 GNDA.n86 9.3005
R346 GNDA.n88 GNDA.n70 9.3005
R347 GNDA.n90 GNDA.n89 9.3005
R348 GNDA.n92 GNDA.n68 9.3005
R349 GNDA.n96 GNDA.n95 9.3005
R350 GNDA.n97 GNDA.n67 9.3005
R351 GNDA.n99 GNDA.n98 9.3005
R352 GNDA.n100 GNDA.n66 9.3005
R353 GNDA.n102 GNDA.n101 9.3005
R354 GNDA.n104 GNDA.n103 9.3005
R355 GNDA.n105 GNDA.n63 9.3005
R356 GNDA.n107 GNDA.n106 9.3005
R357 GNDA.n108 GNDA.n62 9.3005
R358 GNDA.n110 GNDA.n109 9.3005
R359 GNDA.n111 GNDA.n61 9.3005
R360 GNDA.n115 GNDA.n114 9.3005
R361 GNDA.n116 GNDA.n60 9.3005
R362 GNDA.n118 GNDA.n117 9.3005
R363 GNDA.n120 GNDA.n58 9.3005
R364 GNDA.n122 GNDA.n121 9.3005
R365 GNDA.n123 GNDA.n57 9.3005
R366 GNDA.n125 GNDA.n124 9.3005
R367 GNDA.n126 GNDA.n52 9.3005
R368 GNDA.n129 GNDA.n128 9.3005
R369 GNDA.n130 GNDA.n51 9.3005
R370 GNDA.n132 GNDA.n131 9.3005
R371 GNDA.n133 GNDA.n50 9.3005
R372 GNDA.n136 GNDA.n135 9.3005
R373 GNDA.n137 GNDA.n49 9.3005
R374 GNDA.n139 GNDA.n138 9.3005
R375 GNDA.n140 GNDA.n48 9.3005
R376 GNDA.n143 GNDA.n142 9.3005
R377 GNDA.n144 GNDA.n47 9.3005
R378 GNDA.n146 GNDA.n145 9.3005
R379 GNDA.n148 GNDA.n45 9.3005
R380 GNDA.n152 GNDA.n151 9.3005
R381 GNDA.n153 GNDA.n44 9.3005
R382 GNDA.n155 GNDA.n154 9.3005
R383 GNDA.n156 GNDA.n42 9.3005
R384 GNDA.n159 GNDA.n158 9.3005
R385 GNDA.n160 GNDA.n41 9.3005
R386 GNDA.n162 GNDA.n161 9.3005
R387 GNDA.n163 GNDA.n40 9.3005
R388 GNDA.n165 GNDA.n164 9.3005
R389 GNDA.n166 GNDA.n39 9.3005
R390 GNDA.n168 GNDA.n167 9.3005
R391 GNDA.n170 GNDA.n37 9.3005
R392 GNDA.n174 GNDA.n173 9.3005
R393 GNDA.n175 GNDA.n36 9.3005
R394 GNDA.n177 GNDA.n176 9.3005
R395 GNDA.n178 GNDA.n35 9.3005
R396 GNDA.n180 GNDA.n179 9.3005
R397 GNDA.n181 GNDA.n34 9.3005
R398 GNDA.n183 GNDA.n182 9.3005
R399 GNDA.n282 GNDA.n7 9.3005
R400 GNDA.n284 GNDA.n283 9.3005
R401 GNDA.n285 GNDA.n6 9.3005
R402 GNDA.n287 GNDA.n286 9.3005
R403 GNDA.n288 GNDA.n5 9.3005
R404 GNDA.n290 GNDA.n289 9.3005
R405 GNDA.n291 GNDA.n3 9.3005
R406 GNDA.n293 GNDA.n292 9.3005
R407 GNDA.n294 GNDA.n2 9.3005
R408 GNDA.n296 GNDA.n295 9.3005
R409 GNDA.n297 GNDA.n1 9.3005
R410 GNDA.n299 GNDA.n298 9.3005
R411 GNDA.n281 GNDA.n280 7.49856
R412 GNDA.n300 GNDA.n0 6.86152
R413 GNDA.n85 GNDA.n84 6.4005
R414 GNDA.n91 GNDA.n90 6.4005
R415 GNDA.n104 GNDA.n65 6.4005
R416 GNDA.n120 GNDA.n119 6.4005
R417 GNDA.n169 GNDA.n168 6.4005
R418 GNDA.n191 GNDA.n29 6.4005
R419 GNDA.n217 GNDA.n216 6.4005
R420 GNDA.n254 GNDA.n253 6.4005
R421 GNDA.n269 GNDA.n4 4.49344
R422 GNDA.n270 GNDA.n269 4.49344
R423 GNDA.n279 GNDA.n9 4.49344
R424 GNDA.n277 GNDA.n9 4.49344
R425 GNDA.n267 GNDA.n266 3.8278
R426 GNDA.n272 GNDA.n271 3.8278
R427 GNDA.n276 GNDA.n275 3.8278
R428 GNDA.n135 GNDA.n134 3.2005
R429 GNDA.n147 GNDA.n146 3.2005
R430 GNDA.n184 GNDA.n183 3.2005
R431 GNDA.n204 GNDA.n23 3.2005
R432 GNDA.n230 GNDA.n229 3.2005
R433 GNDA.n264 GNDA.n263 2.8779
R434 GNDA.n265 GNDA.n264 2.8779
R435 GNDA GNDA.n300 1.23328
R436 GNDA.n76 GNDA.n73 0.442364
R437 GNDA.n300 GNDA.n299 0.206966
R438 GNDA.n282 GNDA.n281 0.193856
R439 GNDA.n243 GNDA.n8 0.193477
R440 GNDA.n80 GNDA.n73 0.15675
R441 GNDA.n81 GNDA.n80 0.15675
R442 GNDA.n82 GNDA.n81 0.15675
R443 GNDA.n82 GNDA.n71 0.15675
R444 GNDA.n87 GNDA.n71 0.15675
R445 GNDA.n88 GNDA.n87 0.15675
R446 GNDA.n89 GNDA.n88 0.15675
R447 GNDA.n89 GNDA.n68 0.15675
R448 GNDA.n96 GNDA.n68 0.15675
R449 GNDA.n97 GNDA.n96 0.15675
R450 GNDA.n98 GNDA.n97 0.15675
R451 GNDA.n98 GNDA.n66 0.15675
R452 GNDA.n102 GNDA.n66 0.15675
R453 GNDA.n103 GNDA.n102 0.15675
R454 GNDA.n103 GNDA.n63 0.15675
R455 GNDA.n107 GNDA.n63 0.15675
R456 GNDA.n108 GNDA.n107 0.15675
R457 GNDA.n109 GNDA.n108 0.15675
R458 GNDA.n109 GNDA.n61 0.15675
R459 GNDA.n115 GNDA.n61 0.15675
R460 GNDA.n116 GNDA.n115 0.15675
R461 GNDA.n117 GNDA.n116 0.15675
R462 GNDA.n117 GNDA.n58 0.15675
R463 GNDA.n122 GNDA.n58 0.15675
R464 GNDA.n123 GNDA.n122 0.15675
R465 GNDA.n124 GNDA.n123 0.15675
R466 GNDA.n124 GNDA.n52 0.15675
R467 GNDA.n129 GNDA.n52 0.15675
R468 GNDA.n130 GNDA.n129 0.15675
R469 GNDA.n131 GNDA.n130 0.15675
R470 GNDA.n131 GNDA.n50 0.15675
R471 GNDA.n136 GNDA.n50 0.15675
R472 GNDA.n137 GNDA.n136 0.15675
R473 GNDA.n138 GNDA.n137 0.15675
R474 GNDA.n138 GNDA.n48 0.15675
R475 GNDA.n143 GNDA.n48 0.15675
R476 GNDA.n144 GNDA.n143 0.15675
R477 GNDA.n145 GNDA.n144 0.15675
R478 GNDA.n145 GNDA.n45 0.15675
R479 GNDA.n152 GNDA.n45 0.15675
R480 GNDA.n153 GNDA.n152 0.15675
R481 GNDA.n154 GNDA.n153 0.15675
R482 GNDA.n154 GNDA.n42 0.15675
R483 GNDA.n159 GNDA.n42 0.15675
R484 GNDA.n160 GNDA.n159 0.15675
R485 GNDA.n161 GNDA.n160 0.15675
R486 GNDA.n161 GNDA.n40 0.15675
R487 GNDA.n165 GNDA.n40 0.15675
R488 GNDA.n166 GNDA.n165 0.15675
R489 GNDA.n167 GNDA.n166 0.15675
R490 GNDA.n167 GNDA.n37 0.15675
R491 GNDA.n174 GNDA.n37 0.15675
R492 GNDA.n175 GNDA.n174 0.15675
R493 GNDA.n176 GNDA.n175 0.15675
R494 GNDA.n176 GNDA.n35 0.15675
R495 GNDA.n180 GNDA.n35 0.15675
R496 GNDA.n181 GNDA.n180 0.15675
R497 GNDA.n182 GNDA.n181 0.15675
R498 GNDA.n182 GNDA.n32 0.15675
R499 GNDA.n187 GNDA.n32 0.15675
R500 GNDA.n188 GNDA.n187 0.15675
R501 GNDA.n188 GNDA.n30 0.15675
R502 GNDA.n192 GNDA.n30 0.15675
R503 GNDA.n193 GNDA.n192 0.15675
R504 GNDA.n193 GNDA.n26 0.15675
R505 GNDA.n198 GNDA.n26 0.15675
R506 GNDA.n199 GNDA.n198 0.15675
R507 GNDA.n200 GNDA.n199 0.15675
R508 GNDA.n200 GNDA.n24 0.15675
R509 GNDA.n206 GNDA.n24 0.15675
R510 GNDA.n207 GNDA.n206 0.15675
R511 GNDA.n208 GNDA.n207 0.15675
R512 GNDA.n208 GNDA.n21 0.15675
R513 GNDA.n213 GNDA.n21 0.15675
R514 GNDA.n214 GNDA.n213 0.15675
R515 GNDA.n215 GNDA.n214 0.15675
R516 GNDA.n215 GNDA.n18 0.15675
R517 GNDA.n220 GNDA.n18 0.15675
R518 GNDA.n221 GNDA.n220 0.15675
R519 GNDA.n221 GNDA.n15 0.15675
R520 GNDA.n225 GNDA.n15 0.15675
R521 GNDA.n226 GNDA.n225 0.15675
R522 GNDA.n227 GNDA.n226 0.15675
R523 GNDA.n227 GNDA.n12 0.15675
R524 GNDA.n232 GNDA.n12 0.15675
R525 GNDA.n233 GNDA.n232 0.15675
R526 GNDA.n257 GNDA.n233 0.15675
R527 GNDA.n257 GNDA.n256 0.15675
R528 GNDA.n256 GNDA.n255 0.15675
R529 GNDA.n255 GNDA.n234 0.15675
R530 GNDA.n250 GNDA.n234 0.15675
R531 GNDA.n250 GNDA.n249 0.15675
R532 GNDA.n249 GNDA.n238 0.15675
R533 GNDA.n245 GNDA.n238 0.15675
R534 GNDA.n245 GNDA.n244 0.15675
R535 GNDA.n244 GNDA.n243 0.15675
R536 GNDA.n283 GNDA.n282 0.15675
R537 GNDA.n283 GNDA.n6 0.15675
R538 GNDA.n287 GNDA.n6 0.15675
R539 GNDA.n288 GNDA.n287 0.15675
R540 GNDA.n289 GNDA.n288 0.15675
R541 GNDA.n289 GNDA.n3 0.15675
R542 GNDA.n293 GNDA.n3 0.15675
R543 GNDA.n294 GNDA.n293 0.15675
R544 GNDA.n295 GNDA.n294 0.15675
R545 GNDA.n295 GNDA.n1 0.15675
R546 GNDA.n299 GNDA.n1 0.15675
R547 VDDA.t60 VDDA.t64 2804.76
R548 VDDA.t25 VDDA.t9 2533.33
R549 VDDA.t47 VDDA.t86 2307.14
R550 VDDA.t36 VDDA.t15 2216.67
R551 VDDA.t31 VDDA.t17 2216.67
R552 VDDA.t29 VDDA.t13 2216.67
R553 VDDA.t49 VDDA.t55 2126.19
R554 VDDA.t78 VDDA.t90 1538.1
R555 VDDA.t40 VDDA.t33 1492.86
R556 VDDA.t53 VDDA.t88 1492.86
R557 VDDA.t72 VDDA.t84 1317.78
R558 VDDA.n47 VDDA.t34 1289.29
R559 VDDA.t82 VDDA.n146 1289.29
R560 VDDA.t57 VDDA.t0 1130.95
R561 VDDA.t11 VDDA.t68 1130.95
R562 VDDA.t5 VDDA.t70 1130.95
R563 VDDA.t3 VDDA.t7 1130.95
R564 VDDA.t27 VDDA.t45 1130.95
R565 VDDA.n147 VDDA.t92 927.381
R566 VDDA.t38 VDDA.n201 927.381
R567 VDDA.n202 VDDA.t66 927.381
R568 VDDA.t23 VDDA.n248 927.381
R569 VDDA.n265 VDDA.n264 831.25
R570 VDDA.n263 VDDA.n260 831.25
R571 VDDA.n90 VDDA.t56 726.734
R572 VDDA.n124 VDDA.t58 726.734
R573 VDDA.n247 VDDA.t14 663.801
R574 VDDA.n203 VDDA.t32 663.801
R575 VDDA.n200 VDDA.t16 663.801
R576 VDDA.n148 VDDA.t48 663.801
R577 VDDA.n145 VDDA.t65 663.801
R578 VDDA.n48 VDDA.t81 663.801
R579 VDDA.n233 VDDA.n232 647.933
R580 VDDA.n239 VDDA.n230 647.933
R581 VDDA.n219 VDDA.n16 647.933
R582 VDDA.n212 VDDA.n211 647.933
R583 VDDA.n186 VDDA.n178 647.933
R584 VDDA.n192 VDDA.n175 647.933
R585 VDDA.n164 VDDA.n27 647.933
R586 VDDA.n157 VDDA.n156 647.933
R587 VDDA.n105 VDDA.n97 647.933
R588 VDDA.n112 VDDA.n94 647.933
R589 VDDA.n130 VDDA.n87 647.933
R590 VDDA.n137 VDDA.n84 647.933
R591 VDDA.n60 VDDA.n59 647.933
R592 VDDA.n46 VDDA.n45 647.933
R593 VDDA.n72 VDDA.n38 646.715
R594 VDDA.n47 VDDA.t80 610.715
R595 VDDA.n146 VDDA.t64 610.715
R596 VDDA.n147 VDDA.t47 610.715
R597 VDDA.n201 VDDA.t15 610.715
R598 VDDA.n202 VDDA.t31 610.715
R599 VDDA.n248 VDDA.t13 610.715
R600 VDDA.n264 VDDA.n262 585
R601 VDDA.n268 VDDA.n263 585
R602 VDDA.n258 VDDA.t94 537.491
R603 VDDA.n256 VDDA.t96 537.491
R604 VDDA.n249 VDDA.t95 537.491
R605 VDDA.t34 VDDA.t25 497.62
R606 VDDA.t9 VDDA.t40 497.62
R607 VDDA.t33 VDDA.t51 497.62
R608 VDDA.t51 VDDA.t60 497.62
R609 VDDA.t90 VDDA.t82 497.62
R610 VDDA.t0 VDDA.t78 497.62
R611 VDDA.t55 VDDA.t57 497.62
R612 VDDA.t88 VDDA.t49 497.62
R613 VDDA.t86 VDDA.t53 497.62
R614 VDDA.t92 VDDA.t11 497.62
R615 VDDA.t68 VDDA.t36 497.62
R616 VDDA.t70 VDDA.t38 497.62
R617 VDDA.t17 VDDA.t5 497.62
R618 VDDA.t66 VDDA.t3 497.62
R619 VDDA.t7 VDDA.t29 497.62
R620 VDDA.t45 VDDA.t23 497.62
R621 VDDA.t84 VDDA.t27 497.62
R622 VDDA.t20 VDDA.n266 465.079
R623 VDDA.n267 VDDA.t20 465.079
R624 VDDA.t63 VDDA.n273 464.281
R625 VDDA.n275 VDDA.t63 464.281
R626 VDDA.t44 VDDA.n9 464.281
R627 VDDA.n252 VDDA.t44 464.281
R628 VDDA.n248 VDDA.n247 382.8
R629 VDDA.n203 VDDA.n202 382.8
R630 VDDA.n201 VDDA.n200 382.8
R631 VDDA.n148 VDDA.n147 382.8
R632 VDDA.n146 VDDA.n145 382.8
R633 VDDA.n48 VDDA.n47 382.8
R634 VDDA.n258 VDDA.t75 359.752
R635 VDDA.n256 VDDA.t77 359.752
R636 VDDA.n249 VDDA.t73 359.752
R637 VDDA.n279 VDDA.n5 238.367
R638 VDDA.n274 VDDA.n257 238.367
R639 VDDA.n283 VDDA.n282 238.367
R640 VDDA.n255 VDDA.n250 238.367
R641 VDDA.n270 VDDA.n260 238.367
R642 VDDA.n265 VDDA.n259 238.367
R643 VDDA.n281 VDDA.t43 219.232
R644 VDDA.t62 VDDA.n280 219.232
R645 VDDA.t19 VDDA.n271 219.232
R646 VDDA.n271 VDDA.t21 219.232
R647 VDDA.t19 VDDA.n258 185.002
R648 VDDA.t62 VDDA.n256 185.002
R649 VDDA.n249 VDDA.t43 185.002
R650 VDDA.n251 VDDA.n10 185
R651 VDDA.n254 VDDA.n253 185
R652 VDDA.n278 VDDA.n277 185
R653 VDDA.n276 VDDA.n272 185
R654 VDDA.n262 VDDA.n261 185
R655 VDDA.n269 VDDA.n268 185
R656 VDDA.n281 VDDA.t76 158.333
R657 VDDA.n280 VDDA.t74 158.333
R658 VDDA.n269 VDDA.n261 150
R659 VDDA.n278 VDDA.n272 150
R660 VDDA.n254 VDDA.n10 150
R661 VDDA.n264 VDDA.t22 123.126
R662 VDDA.t22 VDDA.n263 123.126
R663 VDDA.t43 VDDA.t59 105.556
R664 VDDA.t42 VDDA.t62 105.556
R665 VDDA.t2 VDDA.t19 105.556
R666 VDDA.n260 VDDA.n258 90.5056
R667 VDDA.n232 VDDA.t28 78.8005
R668 VDDA.n232 VDDA.t85 78.8005
R669 VDDA.n230 VDDA.t24 78.8005
R670 VDDA.n230 VDDA.t46 78.8005
R671 VDDA.n16 VDDA.t8 78.8005
R672 VDDA.n16 VDDA.t30 78.8005
R673 VDDA.n211 VDDA.t67 78.8005
R674 VDDA.n211 VDDA.t4 78.8005
R675 VDDA.n178 VDDA.t6 78.8005
R676 VDDA.n178 VDDA.t18 78.8005
R677 VDDA.n175 VDDA.t39 78.8005
R678 VDDA.n175 VDDA.t71 78.8005
R679 VDDA.n27 VDDA.t69 78.8005
R680 VDDA.n27 VDDA.t37 78.8005
R681 VDDA.n156 VDDA.t93 78.8005
R682 VDDA.n156 VDDA.t12 78.8005
R683 VDDA.n97 VDDA.t54 78.8005
R684 VDDA.n97 VDDA.t87 78.8005
R685 VDDA.n94 VDDA.t50 78.8005
R686 VDDA.n94 VDDA.t89 78.8005
R687 VDDA.n87 VDDA.t79 78.8005
R688 VDDA.n87 VDDA.t1 78.8005
R689 VDDA.n84 VDDA.t83 78.8005
R690 VDDA.n84 VDDA.t91 78.8005
R691 VDDA.n38 VDDA.t52 78.8005
R692 VDDA.n38 VDDA.t61 78.8005
R693 VDDA.n59 VDDA.t10 78.8005
R694 VDDA.n59 VDDA.t41 78.8005
R695 VDDA.n45 VDDA.t35 78.8005
R696 VDDA.n45 VDDA.t26 78.8005
R697 VDDA.n274 VDDA.n256 74.7687
R698 VDDA.n250 VDDA.n249 74.7687
R699 VDDA.n49 VDDA.n48 66.5733
R700 VDDA.n282 VDDA.n281 65.8183
R701 VDDA.n281 VDDA.n255 65.8183
R702 VDDA.n280 VDDA.n279 65.8183
R703 VDDA.n280 VDDA.n257 65.8183
R704 VDDA.n271 VDDA.n259 65.8183
R705 VDDA.n271 VDDA.n270 65.8183
R706 VDDA.n247 VDDA.n246 54.4005
R707 VDDA.n204 VDDA.n203 54.4005
R708 VDDA.n200 VDDA.n199 54.4005
R709 VDDA.n149 VDDA.n148 54.4005
R710 VDDA.n145 VDDA.n144 54.4005
R711 VDDA.n261 VDDA.n259 53.3664
R712 VDDA.n270 VDDA.n269 53.3664
R713 VDDA.n282 VDDA.n10 53.3664
R714 VDDA.n255 VDDA.n254 53.3664
R715 VDDA.n279 VDDA.n278 53.3664
R716 VDDA.n272 VDDA.n257 53.3664
R717 VDDA.n296 VDDA.n295 32.0005
R718 VDDA.n296 VDDA.n2 32.0005
R719 VDDA.n300 VDDA.n2 32.0005
R720 VDDA.n301 VDDA.n300 32.0005
R721 VDDA.n302 VDDA.n301 32.0005
R722 VDDA.n288 VDDA.n7 32.0005
R723 VDDA.n289 VDDA.n288 32.0005
R724 VDDA.n290 VDDA.n289 32.0005
R725 VDDA.n290 VDDA.n4 32.0005
R726 VDDA.n52 VDDA.n51 32.0005
R727 VDDA.n53 VDDA.n52 32.0005
R728 VDDA.n53 VDDA.n43 32.0005
R729 VDDA.n57 VDDA.n43 32.0005
R730 VDDA.n58 VDDA.n57 32.0005
R731 VDDA.n61 VDDA.n58 32.0005
R732 VDDA.n65 VDDA.n41 32.0005
R733 VDDA.n66 VDDA.n65 32.0005
R734 VDDA.n67 VDDA.n66 32.0005
R735 VDDA.n67 VDDA.n39 32.0005
R736 VDDA.n71 VDDA.n39 32.0005
R737 VDDA.n74 VDDA.n73 32.0005
R738 VDDA.n74 VDDA.n36 32.0005
R739 VDDA.n78 VDDA.n36 32.0005
R740 VDDA.n79 VDDA.n78 32.0005
R741 VDDA.n80 VDDA.n79 32.0005
R742 VDDA.n80 VDDA.n33 32.0005
R743 VDDA.n143 VDDA.n34 32.0005
R744 VDDA.n139 VDDA.n34 32.0005
R745 VDDA.n139 VDDA.n138 32.0005
R746 VDDA.n136 VDDA.n85 32.0005
R747 VDDA.n132 VDDA.n85 32.0005
R748 VDDA.n132 VDDA.n131 32.0005
R749 VDDA.n129 VDDA.n88 32.0005
R750 VDDA.n125 VDDA.n88 32.0005
R751 VDDA.n123 VDDA.n122 32.0005
R752 VDDA.n119 VDDA.n118 32.0005
R753 VDDA.n118 VDDA.n117 32.0005
R754 VDDA.n117 VDDA.n92 32.0005
R755 VDDA.n113 VDDA.n92 32.0005
R756 VDDA.n111 VDDA.n110 32.0005
R757 VDDA.n110 VDDA.n95 32.0005
R758 VDDA.n106 VDDA.n95 32.0005
R759 VDDA.n104 VDDA.n103 32.0005
R760 VDDA.n103 VDDA.n98 32.0005
R761 VDDA.n99 VDDA.n98 32.0005
R762 VDDA.n99 VDDA.n32 32.0005
R763 VDDA.n150 VDDA.n32 32.0005
R764 VDDA.n154 VDDA.n30 32.0005
R765 VDDA.n155 VDDA.n154 32.0005
R766 VDDA.n158 VDDA.n155 32.0005
R767 VDDA.n162 VDDA.n28 32.0005
R768 VDDA.n163 VDDA.n162 32.0005
R769 VDDA.n165 VDDA.n25 32.0005
R770 VDDA.n169 VDDA.n25 32.0005
R771 VDDA.n170 VDDA.n169 32.0005
R772 VDDA.n171 VDDA.n170 32.0005
R773 VDDA.n171 VDDA.n22 32.0005
R774 VDDA.n198 VDDA.n23 32.0005
R775 VDDA.n194 VDDA.n23 32.0005
R776 VDDA.n194 VDDA.n193 32.0005
R777 VDDA.n191 VDDA.n176 32.0005
R778 VDDA.n187 VDDA.n176 32.0005
R779 VDDA.n185 VDDA.n184 32.0005
R780 VDDA.n184 VDDA.n179 32.0005
R781 VDDA.n180 VDDA.n179 32.0005
R782 VDDA.n180 VDDA.n21 32.0005
R783 VDDA.n205 VDDA.n21 32.0005
R784 VDDA.n209 VDDA.n19 32.0005
R785 VDDA.n210 VDDA.n209 32.0005
R786 VDDA.n213 VDDA.n210 32.0005
R787 VDDA.n217 VDDA.n17 32.0005
R788 VDDA.n218 VDDA.n217 32.0005
R789 VDDA.n220 VDDA.n14 32.0005
R790 VDDA.n224 VDDA.n14 32.0005
R791 VDDA.n225 VDDA.n224 32.0005
R792 VDDA.n226 VDDA.n225 32.0005
R793 VDDA.n226 VDDA.n11 32.0005
R794 VDDA.n245 VDDA.n12 32.0005
R795 VDDA.n241 VDDA.n12 32.0005
R796 VDDA.n241 VDDA.n240 32.0005
R797 VDDA.n238 VDDA.n231 32.0005
R798 VDDA.n234 VDDA.n231 32.0005
R799 VDDA.n49 VDDA.n46 29.8684
R800 VDDA.n73 VDDA.n72 28.8005
R801 VDDA.n131 VDDA.n130 28.8005
R802 VDDA.n150 VDDA.n149 28.8005
R803 VDDA.n164 VDDA.n163 28.8005
R804 VDDA.n199 VDDA.n22 28.8005
R805 VDDA.n187 VDDA.n186 28.8005
R806 VDDA.n205 VDDA.n204 28.8005
R807 VDDA.n219 VDDA.n218 28.8005
R808 VDDA.n246 VDDA.n11 28.8005
R809 VDDA.n234 VDDA.n233 28.8005
R810 VDDA.n144 VDDA.n143 25.6005
R811 VDDA.n294 VDDA.n5 24.991
R812 VDDA.n284 VDDA.n283 24.991
R813 VDDA.n285 VDDA.n8 24.1919
R814 VDDA.n265 VDDA.n0 23.6611
R815 VDDA.n295 VDDA.n294 22.4005
R816 VDDA.n284 VDDA.n7 22.4005
R817 VDDA.n294 VDDA.n4 22.4005
R818 VDDA.n112 VDDA.n111 22.4005
R819 VDDA.n106 VDDA.n105 22.4005
R820 VDDA.n157 VDDA.n28 22.4005
R821 VDDA.n192 VDDA.n191 22.4005
R822 VDDA.n212 VDDA.n17 22.4005
R823 VDDA.n239 VDDA.n238 22.4005
R824 VDDA.n60 VDDA.n41 19.2005
R825 VDDA.n124 VDDA.n123 19.2005
R826 VDDA.n122 VDDA.n90 19.2005
R827 VDDA.n302 VDDA.n0 16.0005
R828 VDDA.n138 VDDA.n137 16.0005
R829 VDDA.n137 VDDA.n136 16.0005
R830 VDDA.n61 VDDA.n60 12.8005
R831 VDDA.n125 VDDA.n124 12.8005
R832 VDDA.n119 VDDA.n90 12.8005
R833 VDDA.n233 VDDA.n8 10.7016
R834 VDDA.n51 VDDA.n46 9.6005
R835 VDDA.n113 VDDA.n112 9.6005
R836 VDDA.n105 VDDA.n104 9.6005
R837 VDDA.n158 VDDA.n157 9.6005
R838 VDDA.n193 VDDA.n192 9.6005
R839 VDDA.n213 VDDA.n212 9.6005
R840 VDDA.n240 VDDA.n239 9.6005
R841 VDDA.n51 VDDA.n50 9.3005
R842 VDDA.n52 VDDA.n44 9.3005
R843 VDDA.n54 VDDA.n53 9.3005
R844 VDDA.n55 VDDA.n43 9.3005
R845 VDDA.n57 VDDA.n56 9.3005
R846 VDDA.n58 VDDA.n42 9.3005
R847 VDDA.n62 VDDA.n61 9.3005
R848 VDDA.n63 VDDA.n41 9.3005
R849 VDDA.n65 VDDA.n64 9.3005
R850 VDDA.n66 VDDA.n40 9.3005
R851 VDDA.n68 VDDA.n67 9.3005
R852 VDDA.n69 VDDA.n39 9.3005
R853 VDDA.n71 VDDA.n70 9.3005
R854 VDDA.n73 VDDA.n37 9.3005
R855 VDDA.n75 VDDA.n74 9.3005
R856 VDDA.n76 VDDA.n36 9.3005
R857 VDDA.n78 VDDA.n77 9.3005
R858 VDDA.n79 VDDA.n35 9.3005
R859 VDDA.n81 VDDA.n80 9.3005
R860 VDDA.n82 VDDA.n33 9.3005
R861 VDDA.n143 VDDA.n142 9.3005
R862 VDDA.n141 VDDA.n34 9.3005
R863 VDDA.n140 VDDA.n139 9.3005
R864 VDDA.n138 VDDA.n83 9.3005
R865 VDDA.n136 VDDA.n135 9.3005
R866 VDDA.n134 VDDA.n85 9.3005
R867 VDDA.n133 VDDA.n132 9.3005
R868 VDDA.n131 VDDA.n86 9.3005
R869 VDDA.n129 VDDA.n128 9.3005
R870 VDDA.n127 VDDA.n88 9.3005
R871 VDDA.n126 VDDA.n125 9.3005
R872 VDDA.n123 VDDA.n89 9.3005
R873 VDDA.n122 VDDA.n121 9.3005
R874 VDDA.n120 VDDA.n119 9.3005
R875 VDDA.n118 VDDA.n91 9.3005
R876 VDDA.n117 VDDA.n116 9.3005
R877 VDDA.n115 VDDA.n92 9.3005
R878 VDDA.n114 VDDA.n113 9.3005
R879 VDDA.n111 VDDA.n93 9.3005
R880 VDDA.n110 VDDA.n109 9.3005
R881 VDDA.n108 VDDA.n95 9.3005
R882 VDDA.n107 VDDA.n106 9.3005
R883 VDDA.n104 VDDA.n96 9.3005
R884 VDDA.n103 VDDA.n102 9.3005
R885 VDDA.n101 VDDA.n98 9.3005
R886 VDDA.n100 VDDA.n99 9.3005
R887 VDDA.n32 VDDA.n31 9.3005
R888 VDDA.n151 VDDA.n150 9.3005
R889 VDDA.n152 VDDA.n30 9.3005
R890 VDDA.n154 VDDA.n153 9.3005
R891 VDDA.n155 VDDA.n29 9.3005
R892 VDDA.n159 VDDA.n158 9.3005
R893 VDDA.n160 VDDA.n28 9.3005
R894 VDDA.n162 VDDA.n161 9.3005
R895 VDDA.n163 VDDA.n26 9.3005
R896 VDDA.n166 VDDA.n165 9.3005
R897 VDDA.n167 VDDA.n25 9.3005
R898 VDDA.n169 VDDA.n168 9.3005
R899 VDDA.n170 VDDA.n24 9.3005
R900 VDDA.n172 VDDA.n171 9.3005
R901 VDDA.n173 VDDA.n22 9.3005
R902 VDDA.n198 VDDA.n197 9.3005
R903 VDDA.n196 VDDA.n23 9.3005
R904 VDDA.n195 VDDA.n194 9.3005
R905 VDDA.n193 VDDA.n174 9.3005
R906 VDDA.n191 VDDA.n190 9.3005
R907 VDDA.n189 VDDA.n176 9.3005
R908 VDDA.n188 VDDA.n187 9.3005
R909 VDDA.n185 VDDA.n177 9.3005
R910 VDDA.n184 VDDA.n183 9.3005
R911 VDDA.n182 VDDA.n179 9.3005
R912 VDDA.n181 VDDA.n180 9.3005
R913 VDDA.n21 VDDA.n20 9.3005
R914 VDDA.n206 VDDA.n205 9.3005
R915 VDDA.n207 VDDA.n19 9.3005
R916 VDDA.n209 VDDA.n208 9.3005
R917 VDDA.n210 VDDA.n18 9.3005
R918 VDDA.n214 VDDA.n213 9.3005
R919 VDDA.n215 VDDA.n17 9.3005
R920 VDDA.n217 VDDA.n216 9.3005
R921 VDDA.n218 VDDA.n15 9.3005
R922 VDDA.n221 VDDA.n220 9.3005
R923 VDDA.n222 VDDA.n14 9.3005
R924 VDDA.n224 VDDA.n223 9.3005
R925 VDDA.n225 VDDA.n13 9.3005
R926 VDDA.n227 VDDA.n226 9.3005
R927 VDDA.n228 VDDA.n11 9.3005
R928 VDDA.n245 VDDA.n244 9.3005
R929 VDDA.n243 VDDA.n12 9.3005
R930 VDDA.n242 VDDA.n241 9.3005
R931 VDDA.n240 VDDA.n229 9.3005
R932 VDDA.n238 VDDA.n237 9.3005
R933 VDDA.n236 VDDA.n231 9.3005
R934 VDDA.n235 VDDA.n234 9.3005
R935 VDDA.n286 VDDA.n7 9.3005
R936 VDDA.n288 VDDA.n287 9.3005
R937 VDDA.n289 VDDA.n6 9.3005
R938 VDDA.n291 VDDA.n290 9.3005
R939 VDDA.n292 VDDA.n4 9.3005
R940 VDDA.n294 VDDA.n293 9.3005
R941 VDDA.n295 VDDA.n3 9.3005
R942 VDDA.n297 VDDA.n296 9.3005
R943 VDDA.n298 VDDA.n2 9.3005
R944 VDDA.n300 VDDA.n299 9.3005
R945 VDDA.n301 VDDA.n1 9.3005
R946 VDDA.n303 VDDA.n302 9.3005
R947 VDDA.n277 VDDA.n276 9.14336
R948 VDDA.n253 VDDA.n251 9.14336
R949 VDDA.n304 VDDA.n0 7.37301
R950 VDDA.n285 VDDA.n284 7.05969
R951 VDDA.n144 VDDA.n33 6.4005
R952 VDDA.n268 VDDA.n262 5.81868
R953 VDDA.n273 VDDA.n5 5.33286
R954 VDDA.n275 VDDA.n274 5.33286
R955 VDDA.n283 VDDA.n9 5.33286
R956 VDDA.n252 VDDA.n250 5.33286
R957 VDDA.t59 VDDA.t72 4.06033
R958 VDDA.t76 VDDA.t42 4.06033
R959 VDDA.t74 VDDA.t2 4.06033
R960 VDDA.n277 VDDA.n273 3.75335
R961 VDDA.n276 VDDA.n275 3.75335
R962 VDDA.n251 VDDA.n9 3.75335
R963 VDDA.n253 VDDA.n252 3.75335
R964 VDDA.n266 VDDA.n265 3.40194
R965 VDDA.n267 VDDA.n260 3.40194
R966 VDDA.n72 VDDA.n71 3.2005
R967 VDDA.n130 VDDA.n129 3.2005
R968 VDDA.n149 VDDA.n30 3.2005
R969 VDDA.n165 VDDA.n164 3.2005
R970 VDDA.n199 VDDA.n198 3.2005
R971 VDDA.n186 VDDA.n185 3.2005
R972 VDDA.n204 VDDA.n19 3.2005
R973 VDDA.n220 VDDA.n219 3.2005
R974 VDDA.n246 VDDA.n245 3.2005
R975 VDDA.n266 VDDA.n262 2.39444
R976 VDDA.n268 VDDA.n267 2.39444
R977 VDDA VDDA.n304 0.774519
R978 VDDA.n50 VDDA.n49 0.224489
R979 VDDA.n286 VDDA.n285 0.202927
R980 VDDA.n304 VDDA.n303 0.196483
R981 VDDA.n235 VDDA.n8 0.193477
R982 VDDA.n50 VDDA.n44 0.15675
R983 VDDA.n54 VDDA.n44 0.15675
R984 VDDA.n55 VDDA.n54 0.15675
R985 VDDA.n56 VDDA.n55 0.15675
R986 VDDA.n56 VDDA.n42 0.15675
R987 VDDA.n62 VDDA.n42 0.15675
R988 VDDA.n63 VDDA.n62 0.15675
R989 VDDA.n64 VDDA.n63 0.15675
R990 VDDA.n64 VDDA.n40 0.15675
R991 VDDA.n68 VDDA.n40 0.15675
R992 VDDA.n69 VDDA.n68 0.15675
R993 VDDA.n70 VDDA.n69 0.15675
R994 VDDA.n70 VDDA.n37 0.15675
R995 VDDA.n75 VDDA.n37 0.15675
R996 VDDA.n76 VDDA.n75 0.15675
R997 VDDA.n77 VDDA.n76 0.15675
R998 VDDA.n77 VDDA.n35 0.15675
R999 VDDA.n81 VDDA.n35 0.15675
R1000 VDDA.n82 VDDA.n81 0.15675
R1001 VDDA.n142 VDDA.n82 0.15675
R1002 VDDA.n142 VDDA.n141 0.15675
R1003 VDDA.n141 VDDA.n140 0.15675
R1004 VDDA.n140 VDDA.n83 0.15675
R1005 VDDA.n135 VDDA.n83 0.15675
R1006 VDDA.n135 VDDA.n134 0.15675
R1007 VDDA.n134 VDDA.n133 0.15675
R1008 VDDA.n133 VDDA.n86 0.15675
R1009 VDDA.n128 VDDA.n86 0.15675
R1010 VDDA.n128 VDDA.n127 0.15675
R1011 VDDA.n127 VDDA.n126 0.15675
R1012 VDDA.n126 VDDA.n89 0.15675
R1013 VDDA.n121 VDDA.n89 0.15675
R1014 VDDA.n121 VDDA.n120 0.15675
R1015 VDDA.n120 VDDA.n91 0.15675
R1016 VDDA.n116 VDDA.n91 0.15675
R1017 VDDA.n116 VDDA.n115 0.15675
R1018 VDDA.n115 VDDA.n114 0.15675
R1019 VDDA.n114 VDDA.n93 0.15675
R1020 VDDA.n109 VDDA.n93 0.15675
R1021 VDDA.n109 VDDA.n108 0.15675
R1022 VDDA.n108 VDDA.n107 0.15675
R1023 VDDA.n107 VDDA.n96 0.15675
R1024 VDDA.n102 VDDA.n96 0.15675
R1025 VDDA.n102 VDDA.n101 0.15675
R1026 VDDA.n101 VDDA.n100 0.15675
R1027 VDDA.n100 VDDA.n31 0.15675
R1028 VDDA.n151 VDDA.n31 0.15675
R1029 VDDA.n152 VDDA.n151 0.15675
R1030 VDDA.n153 VDDA.n152 0.15675
R1031 VDDA.n153 VDDA.n29 0.15675
R1032 VDDA.n159 VDDA.n29 0.15675
R1033 VDDA.n160 VDDA.n159 0.15675
R1034 VDDA.n161 VDDA.n160 0.15675
R1035 VDDA.n161 VDDA.n26 0.15675
R1036 VDDA.n166 VDDA.n26 0.15675
R1037 VDDA.n167 VDDA.n166 0.15675
R1038 VDDA.n168 VDDA.n167 0.15675
R1039 VDDA.n168 VDDA.n24 0.15675
R1040 VDDA.n172 VDDA.n24 0.15675
R1041 VDDA.n173 VDDA.n172 0.15675
R1042 VDDA.n197 VDDA.n173 0.15675
R1043 VDDA.n197 VDDA.n196 0.15675
R1044 VDDA.n196 VDDA.n195 0.15675
R1045 VDDA.n195 VDDA.n174 0.15675
R1046 VDDA.n190 VDDA.n174 0.15675
R1047 VDDA.n190 VDDA.n189 0.15675
R1048 VDDA.n189 VDDA.n188 0.15675
R1049 VDDA.n188 VDDA.n177 0.15675
R1050 VDDA.n183 VDDA.n177 0.15675
R1051 VDDA.n183 VDDA.n182 0.15675
R1052 VDDA.n182 VDDA.n181 0.15675
R1053 VDDA.n181 VDDA.n20 0.15675
R1054 VDDA.n206 VDDA.n20 0.15675
R1055 VDDA.n207 VDDA.n206 0.15675
R1056 VDDA.n208 VDDA.n207 0.15675
R1057 VDDA.n208 VDDA.n18 0.15675
R1058 VDDA.n214 VDDA.n18 0.15675
R1059 VDDA.n215 VDDA.n214 0.15675
R1060 VDDA.n216 VDDA.n215 0.15675
R1061 VDDA.n216 VDDA.n15 0.15675
R1062 VDDA.n221 VDDA.n15 0.15675
R1063 VDDA.n222 VDDA.n221 0.15675
R1064 VDDA.n223 VDDA.n222 0.15675
R1065 VDDA.n223 VDDA.n13 0.15675
R1066 VDDA.n227 VDDA.n13 0.15675
R1067 VDDA.n228 VDDA.n227 0.15675
R1068 VDDA.n244 VDDA.n228 0.15675
R1069 VDDA.n244 VDDA.n243 0.15675
R1070 VDDA.n243 VDDA.n242 0.15675
R1071 VDDA.n242 VDDA.n229 0.15675
R1072 VDDA.n237 VDDA.n229 0.15675
R1073 VDDA.n237 VDDA.n236 0.15675
R1074 VDDA.n236 VDDA.n235 0.15675
R1075 VDDA.n287 VDDA.n286 0.15675
R1076 VDDA.n287 VDDA.n6 0.15675
R1077 VDDA.n291 VDDA.n6 0.15675
R1078 VDDA.n292 VDDA.n291 0.15675
R1079 VDDA.n293 VDDA.n292 0.15675
R1080 VDDA.n293 VDDA.n3 0.15675
R1081 VDDA.n297 VDDA.n3 0.15675
R1082 VDDA.n298 VDDA.n297 0.15675
R1083 VDDA.n299 VDDA.n298 0.15675
R1084 VDDA.n299 VDDA.n1 0.15675
R1085 VDDA.n303 VDDA.n1 0.15675
R1086 vco2_3_0.V4.t2 vco2_3_0.V4.n0 708.125
R1087 vco2_3_0.V4.t2 vco2_3_0.V4.n1 708.125
R1088 vco2_3_0.V4.n1 vco2_3_0.V4.t0 410.519
R1089 vco2_3_0.V4.n0 vco2_3_0.V4.t1 305.649
R1090 vco2_3_0.V4.n1 vco2_3_0.V4.n0 21.3338
R1091 div120_2_0.div3_3_0.CLK.n3 div120_2_0.div3_3_0.CLK.n2 742.51
R1092 div120_2_0.div3_3_0.CLK.n9 div120_2_0.div3_3_0.CLK.t1 723.534
R1093 div120_2_0.div3_3_0.CLK.n8 div120_2_0.div3_3_0.CLK.t2 723.534
R1094 div120_2_0.div3_3_0.CLK.n2 div120_2_0.div3_3_0.CLK.n1 684.806
R1095 div120_2_0.div3_3_0.CLK.n7 div120_2_0.div3_3_0.CLK.n6 366.856
R1096 div120_2_0.div3_3_0.CLK.n0 div120_2_0.div3_3_0.CLK.t4 337.401
R1097 div120_2_0.div3_3_0.CLK.n0 div120_2_0.div3_3_0.CLK.t3 305.267
R1098 div120_2_0.div3_3_0.CLK.t0 div120_2_0.div3_3_0.CLK.n9 254.333
R1099 div120_2_0.div3_3_0.CLK.n4 div120_2_0.div3_3_0.CLK.n3 224.934
R1100 div120_2_0.div3_3_0.CLK.n7 div120_2_0.div3_3_0.CLK.t7 190.123
R1101 div120_2_0.div3_3_0.CLK.n8 div120_2_0.div3_3_0.CLK.n7 187.201
R1102 div120_2_0.div3_3_0.CLK.n1 div120_2_0.div3_3_0.CLK.n0 176.733
R1103 div120_2_0.div3_3_0.CLK.n5 div120_2_0.div3_3_0.CLK.n4 176.733
R1104 div120_2_0.div3_3_0.CLK.n6 div120_2_0.div3_3_0.CLK.n5 176.733
R1105 div120_2_0.div3_3_0.CLK.n3 div120_2_0.div3_3_0.CLK.t12 144.601
R1106 div120_2_0.div3_3_0.CLK.n2 div120_2_0.div3_3_0.CLK.t8 131.976
R1107 div120_2_0.div3_3_0.CLK.n0 div120_2_0.div3_3_0.CLK.t10 128.534
R1108 div120_2_0.div3_3_0.CLK.n1 div120_2_0.div3_3_0.CLK.t6 128.534
R1109 div120_2_0.div3_3_0.CLK.n4 div120_2_0.div3_3_0.CLK.t5 112.468
R1110 div120_2_0.div3_3_0.CLK.n6 div120_2_0.div3_3_0.CLK.t9 112.468
R1111 div120_2_0.div3_3_0.CLK.n5 div120_2_0.div3_3_0.CLK.t11 112.468
R1112 div120_2_0.div3_3_0.CLK.n9 div120_2_0.div3_3_0.CLK.n8 70.4005
R1113 div120_2_0.div3_3_0.H.n0 div120_2_0.div3_3_0.H.t3 723.534
R1114 div120_2_0.div3_3_0.H.n1 div120_2_0.div3_3_0.H.t4 553.534
R1115 div120_2_0.div3_3_0.H.n0 div120_2_0.div3_3_0.H.t1 254.333
R1116 div120_2_0.div3_3_0.H.n2 div120_2_0.div3_3_0.H.n1 206.333
R1117 div120_2_0.div3_3_0.H.n1 div120_2_0.div3_3_0.H.n0 70.4005
R1118 div120_2_0.div3_3_0.H.t2 div120_2_0.div3_3_0.H.n2 48.0005
R1119 div120_2_0.div3_3_0.H.n2 div120_2_0.div3_3_0.H.t0 48.0005
R1120 div120_2_0.div5_2_0.E.n0 div120_2_0.div5_2_0.E.t1 723
R1121 div120_2_0.div5_2_0.E.t2 div120_2_0.div5_2_0.E.t3 514.134
R1122 div120_2_0.div5_2_0.E.n0 div120_2_0.div5_2_0.E.t2 335.983
R1123 div120_2_0.div5_2_0.E.t0 div120_2_0.div5_2_0.E.n0 314.921
R1124 div120_2_0.div5_2_0.F.t0 div120_2_0.div5_2_0.F.t1 157.601
R1125 div120_2_0.div3_3_0.I.n0 div120_2_0.div3_3_0.I.t0 663.801
R1126 div120_2_0.div3_3_0.I.t6 div120_2_0.div3_3_0.I.t2 514.134
R1127 div120_2_0.div3_3_0.I.n0 div120_2_0.div3_3_0.I.t6 479.284
R1128 div120_2_0.div3_3_0.I.n3 div120_2_0.div3_3_0.I.n2 344.8
R1129 div120_2_0.div3_3_0.I.n1 div120_2_0.div3_3_0.I.t3 289.2
R1130 div120_2_0.div3_3_0.I.t1 div120_2_0.div3_3_0.I.n3 275.454
R1131 div120_2_0.div3_3_0.I.n2 div120_2_0.div3_3_0.I.t5 241
R1132 div120_2_0.div3_3_0.I.n1 div120_2_0.div3_3_0.I.t4 112.468
R1133 div120_2_0.div3_3_0.I.n3 div120_2_0.div3_3_0.I.n0 97.9205
R1134 div120_2_0.div3_3_0.I.n2 div120_2_0.div3_3_0.I.n1 64.2672
R1135 div120_2_0.div3_3_0.G.t0 div120_2_0.div3_3_0.G.t1 96.0005
R1136 a_2510_770.n5 a_2510_770.t2 752.333
R1137 a_2510_770.n4 a_2510_770.t0 752.333
R1138 a_2510_770.n0 a_2510_770.t3 514.134
R1139 a_2510_770.n3 a_2510_770.n2 366.856
R1140 a_2510_770.t1 a_2510_770.n5 254.333
R1141 a_2510_770.n3 a_2510_770.t6 190.123
R1142 a_2510_770.n4 a_2510_770.n3 187.201
R1143 a_2510_770.n1 a_2510_770.n0 176.733
R1144 a_2510_770.n2 a_2510_770.n1 176.733
R1145 a_2510_770.n0 a_2510_770.t5 112.468
R1146 a_2510_770.n2 a_2510_770.t7 112.468
R1147 a_2510_770.n1 a_2510_770.t4 112.468
R1148 a_2510_770.n5 a_2510_770.n4 70.4005
R1149 div120_2_0.div2.t4 div120_2_0.div2.t2 1012.2
R1150 div120_2_0.div2.n0 div120_2_0.div2.t1 663.801
R1151 div120_2_0.div2.n2 div120_2_0.div2.n1 431.401
R1152 div120_2_0.div2.t3 div120_2_0.div2.t6 401.668
R1153 div120_2_0.div2.n0 div120_2_0.div2.t4 361.692
R1154 div120_2_0.div2.n1 div120_2_0.div2.t5 353.467
R1155 div120_2_0.div2.t0 div120_2_0.div2.n2 298.921
R1156 div120_2_0.div2.n1 div120_2_0.div2.t3 257.067
R1157 div120_2_0.div2.n2 div120_2_0.div2.n0 67.2005
R1158 a_5110_770.n5 a_5110_770.t1 752.333
R1159 a_5110_770.n4 a_5110_770.t0 752.333
R1160 a_5110_770.n0 a_5110_770.t7 514.134
R1161 a_5110_770.n3 a_5110_770.n2 366.856
R1162 a_5110_770.t2 a_5110_770.n5 254.333
R1163 a_5110_770.n3 a_5110_770.t4 190.123
R1164 a_5110_770.n4 a_5110_770.n3 187.201
R1165 a_5110_770.n1 a_5110_770.n0 176.733
R1166 a_5110_770.n2 a_5110_770.n1 176.733
R1167 a_5110_770.n0 a_5110_770.t5 112.468
R1168 a_5110_770.n2 a_5110_770.t6 112.468
R1169 a_5110_770.n1 a_5110_770.t3 112.468
R1170 a_5110_770.n5 a_5110_770.n4 70.4005
R1171 div120_2_0.div2_4_0.C.n0 div120_2_0.div2_4_0.C.t0 750.201
R1172 div120_2_0.div2_4_0.C.n1 div120_2_0.div2_4_0.C.t4 349.433
R1173 div120_2_0.div2_4_0.C.n0 div120_2_0.div2_4_0.C.t1 276.733
R1174 div120_2_0.div2_4_0.C.n2 div120_2_0.div2_4_0.C.n1 206.333
R1175 div120_2_0.div2_4_0.C.n1 div120_2_0.div2_4_0.C.n0 48.0005
R1176 div120_2_0.div2_4_0.C.n2 div120_2_0.div2_4_0.C.t2 48.0005
R1177 div120_2_0.div2_4_0.C.t3 div120_2_0.div2_4_0.C.n2 48.0005
R1178 div120_2_0.div2_4_2.C.n0 div120_2_0.div2_4_2.C.t3 750.201
R1179 div120_2_0.div2_4_2.C.n1 div120_2_0.div2_4_2.C.t4 349.433
R1180 div120_2_0.div2_4_2.C.n0 div120_2_0.div2_4_2.C.t1 276.733
R1181 div120_2_0.div2_4_2.C.n2 div120_2_0.div2_4_2.C.n1 206.333
R1182 div120_2_0.div2_4_2.C.n1 div120_2_0.div2_4_2.C.n0 48.0005
R1183 div120_2_0.div2_4_2.C.t0 div120_2_0.div2_4_2.C.n2 48.0005
R1184 div120_2_0.div2_4_2.C.n2 div120_2_0.div2_4_2.C.t2 48.0005
R1185 div120_2_0.div4.t5 div120_2_0.div4.t6 1012.2
R1186 div120_2_0.div4.n0 div120_2_0.div4.t0 663.801
R1187 div120_2_0.div4.n2 div120_2_0.div4.n1 431.401
R1188 div120_2_0.div4.t4 div120_2_0.div4.t2 401.668
R1189 div120_2_0.div4.n0 div120_2_0.div4.t5 361.692
R1190 div120_2_0.div4.n1 div120_2_0.div4.t3 353.467
R1191 div120_2_0.div4.t1 div120_2_0.div4.n2 298.921
R1192 div120_2_0.div4.n1 div120_2_0.div4.t4 257.067
R1193 div120_2_0.div4.n2 div120_2_0.div4.n0 67.2005
R1194 div120_2_0.div5_2_0.Q2_b.n4 div120_2_0.div5_2_0.Q2_b.t0 777.4
R1195 div120_2_0.div5_2_0.Q2_b.t2 div120_2_0.div5_2_0.Q2_b.t11 514.134
R1196 div120_2_0.div5_2_0.Q2_b.n3 div120_2_0.div5_2_0.Q2_b.n2 364.178
R1197 div120_2_0.div5_2_0.Q2_b.n0 div120_2_0.div5_2_0.Q2_b.t8 353.467
R1198 div120_2_0.div5_2_0.Q2_b.t3 div120_2_0.div5_2_0.Q2_b.n5 353.467
R1199 div120_2_0.div5_2_0.Q2_b.n6 div120_2_0.div5_2_0.Q2_b.t3 318.702
R1200 div120_2_0.div5_2_0.Q2_b.n6 div120_2_0.div5_2_0.Q2_b.t2 307.909
R1201 div120_2_0.div5_2_0.Q2_b.n5 div120_2_0.div5_2_0.Q2_b.t10 289.2
R1202 div120_2_0.div5_2_0.Q2_b.n4 div120_2_0.div5_2_0.Q2_b.n3 257.079
R1203 div120_2_0.div5_2_0.Q2_b.t1 div120_2_0.div5_2_0.Q2_b.n7 233
R1204 div120_2_0.div5_2_0.Q2_b.n0 div120_2_0.div5_2_0.Q2_b.t5 192.8
R1205 div120_2_0.div5_2_0.Q2_b.n2 div120_2_0.div5_2_0.Q2_b.n1 176.733
R1206 div120_2_0.div5_2_0.Q2_b.n2 div120_2_0.div5_2_0.Q2_b.t6 112.468
R1207 div120_2_0.div5_2_0.Q2_b.n1 div120_2_0.div5_2_0.Q2_b.t9 112.468
R1208 div120_2_0.div5_2_0.Q2_b.n3 div120_2_0.div5_2_0.Q2_b.t4 112.468
R1209 div120_2_0.div5_2_0.Q2_b.n5 div120_2_0.div5_2_0.Q2_b.t7 112.468
R1210 div120_2_0.div5_2_0.Q2_b.n1 div120_2_0.div5_2_0.Q2_b.n0 96.4005
R1211 div120_2_0.div5_2_0.Q2_b.n7 div120_2_0.div5_2_0.Q2_b.n6 38.2642
R1212 div120_2_0.div5_2_0.Q2_b.n7 div120_2_0.div5_2_0.Q2_b.n4 21.3338
R1213 div120_2_0.div5_2_0.H.t0 div120_2_0.div5_2_0.H.t1 96.0005
R1214 div120_2_0.div5_2_0.I.t0 div120_2_0.div5_2_0.I.n0 531.067
R1215 div120_2_0.div5_2_0.I.n0 div120_2_0.div5_2_0.I.t1 48.0005
R1216 div120_2_0.div5_2_0.I.n0 div120_2_0.div5_2_0.I.t2 48.0005
R1217 vco2_3_0.V8.n1 vco2_3_0.V8.n0 412.034
R1218 vco2_3_0.V8.t1 vco2_3_0.V8.n1 372.118
R1219 vco2_3_0.V8.n1 vco2_3_0.V8.t0 247.934
R1220 vco2_3_0.V8.n0 vco2_3_0.V8.t3 186.775
R1221 vco2_3_0.V8.n0 vco2_3_0.V8.t2 126.525
R1222 V_OSC.n2 V_OSC.n0 433.8
R1223 V_OSC.t2 V_OSC.t4 401.668
R1224 V_OSC.t1 V_OSC.n3 372.118
R1225 V_OSC.n0 V_OSC.t6 353.467
R1226 V_OSC.n0 V_OSC.t2 257.067
R1227 V_OSC.n3 V_OSC.t0 247.934
R1228 V_OSC.n3 V_OSC.n2 235.156
R1229 V_OSC.n2 V_OSC.n1 200.833
R1230 V_OSC.n1 V_OSC.t5 186.775
R1231 V_OSC.n1 V_OSC.t3 126.525
R1232 vco2_3_0.V3.n0 vco2_3_0.V3.t1 284.2
R1233 vco2_3_0.V3.n0 vco2_3_0.V3.t2 233
R1234 vco2_3_0.V3.t0 vco2_3_0.V3.n0 184.191
R1235 div120_2_0.div8.t3 div120_2_0.div8.t5 1012.2
R1236 div120_2_0.div8.n0 div120_2_0.div8.t1 663.801
R1237 div120_2_0.div8.n2 div120_2_0.div8.n1 431.401
R1238 div120_2_0.div8.t2 div120_2_0.div8.t4 401.668
R1239 div120_2_0.div8.n0 div120_2_0.div8.t3 361.692
R1240 div120_2_0.div8.t0 div120_2_0.div8.n2 298.921
R1241 div120_2_0.div8.n1 div120_2_0.div8.t2 257.067
R1242 div120_2_0.div8.n1 div120_2_0.div8.t6 208.868
R1243 div120_2_0.div8.n2 div120_2_0.div8.n0 67.2005
R1244 div120_2_0.div3_3_0.C.n0 div120_2_0.div3_3_0.C.t3 721.4
R1245 div120_2_0.div3_3_0.C.n1 div120_2_0.div3_3_0.C.t4 350.349
R1246 div120_2_0.div3_3_0.C.n0 div120_2_0.div3_3_0.C.t1 276.733
R1247 div120_2_0.div3_3_0.C.n2 div120_2_0.div3_3_0.C.n1 206.333
R1248 div120_2_0.div3_3_0.C.n1 div120_2_0.div3_3_0.C.n0 48.0005
R1249 div120_2_0.div3_3_0.C.t2 div120_2_0.div3_3_0.C.n2 48.0005
R1250 div120_2_0.div3_3_0.C.n2 div120_2_0.div3_3_0.C.t0 48.0005
R1251 div120_2_0.div3_3_0.B.t0 div120_2_0.div3_3_0.B.t1 96.0005
R1252 div120_2_0.div3_3_0.A.n0 div120_2_0.div3_3_0.A.t0 713.933
R1253 div120_2_0.div3_3_0.A.n0 div120_2_0.div3_3_0.A.t2 314.233
R1254 div120_2_0.div3_3_0.A.t1 div120_2_0.div3_3_0.A.n0 308.2
R1255 div120_2_0.div2_4_0.A.n0 div120_2_0.div2_4_0.A.t0 713.933
R1256 div120_2_0.div2_4_0.A.t1 div120_2_0.div2_4_0.A.n0 337
R1257 div120_2_0.div2_4_0.A.n0 div120_2_0.div2_4_0.A.t2 314.233
R1258 div120_2_0.div3_3_0.E.n0 div120_2_0.div3_3_0.E.t1 685.134
R1259 div120_2_0.div3_3_0.E.n1 div120_2_0.div3_3_0.E.t2 663.801
R1260 div120_2_0.div3_3_0.E.n0 div120_2_0.div3_3_0.E.t3 534.268
R1261 div120_2_0.div3_3_0.E.t0 div120_2_0.div3_3_0.E.n1 362.921
R1262 div120_2_0.div3_3_0.E.n1 div120_2_0.div3_3_0.E.n0 91.7338
R1263 div120_2_0.div3_3_0.F.t0 div120_2_0.div3_3_0.F.t1 96.0005
R1264 div120_2_0.div5_2_0.A.t2 div120_2_0.div5_2_0.A.n2 755.534
R1265 div120_2_0.div5_2_0.A.n2 div120_2_0.div5_2_0.A.t1 685.134
R1266 div120_2_0.div5_2_0.A.n1 div120_2_0.div5_2_0.A.n0 389.733
R1267 div120_2_0.div5_2_0.A.n1 div120_2_0.div5_2_0.A.t0 340.2
R1268 div120_2_0.div5_2_0.A.n0 div120_2_0.div5_2_0.A.t4 321.334
R1269 div120_2_0.div5_2_0.A.n0 div120_2_0.div5_2_0.A.t3 144.601
R1270 div120_2_0.div5_2_0.A.n2 div120_2_0.div5_2_0.A.n1 19.2005
R1271 div120_2_0.div5_2_0.K.n0 div120_2_0.div5_2_0.K.t0 663.801
R1272 div120_2_0.div5_2_0.K.t1 div120_2_0.div5_2_0.K.n0 397.053
R1273 div120_2_0.div5_2_0.K.n0 div120_2_0.div5_2_0.K.t2 355.378
R1274 div120_2_0.div5_2_0.M.n0 div120_2_0.div5_2_0.M.t0 761.4
R1275 div120_2_0.div5_2_0.M.n1 div120_2_0.div5_2_0.M.t4 349.433
R1276 div120_2_0.div5_2_0.M.n0 div120_2_0.div5_2_0.M.t2 254.333
R1277 div120_2_0.div5_2_0.M.n2 div120_2_0.div5_2_0.M.n1 206.333
R1278 div120_2_0.div5_2_0.M.n1 div120_2_0.div5_2_0.M.n0 70.4005
R1279 div120_2_0.div5_2_0.M.t3 div120_2_0.div5_2_0.M.n2 48.0005
R1280 div120_2_0.div5_2_0.M.n2 div120_2_0.div5_2_0.M.t1 48.0005
R1281 div120_2_0.div5_2_0.L.t0 div120_2_0.div5_2_0.L.t1 96.0005
R1282 div120_2_0.div5_2_0.G.n0 div120_2_0.div5_2_0.G.t1 685.134
R1283 div120_2_0.div5_2_0.G.n1 div120_2_0.div5_2_0.G.t2 685.134
R1284 div120_2_0.div5_2_0.G.n0 div120_2_0.div5_2_0.G.t3 534.268
R1285 div120_2_0.div5_2_0.G.t0 div120_2_0.div5_2_0.G.n1 340.521
R1286 div120_2_0.div5_2_0.G.n1 div120_2_0.div5_2_0.G.n0 105.6
R1287 div120_2_0.div5_2_0.J.n0 div120_2_0.div5_2_0.J.t0 723.534
R1288 div120_2_0.div5_2_0.J.n1 div120_2_0.div5_2_0.J.t4 553.534
R1289 div120_2_0.div5_2_0.J.n0 div120_2_0.div5_2_0.J.t2 254.333
R1290 div120_2_0.div5_2_0.J.n2 div120_2_0.div5_2_0.J.n1 206.333
R1291 div120_2_0.div5_2_0.J.n1 div120_2_0.div5_2_0.J.n0 70.4005
R1292 div120_2_0.div5_2_0.J.n2 div120_2_0.div5_2_0.J.t3 48.0005
R1293 div120_2_0.div5_2_0.J.t1 div120_2_0.div5_2_0.J.n2 48.0005
R1294 div120_2_0.div24.n3 div120_2_0.div24.n2 919.244
R1295 div120_2_0.div24.n8 div120_2_0.div24.n7 918.702
R1296 div120_2_0.div24.t11 div120_2_0.div24.t5 819.4
R1297 div120_2_0.div24.n10 div120_2_0.div24.n9 628.734
R1298 div120_2_0.div24.n2 div120_2_0.div24.n1 520.361
R1299 div120_2_0.div24.n7 div120_2_0.div24.n6 364.178
R1300 div120_2_0.div24.n0 div120_2_0.div24.t10 337.401
R1301 div120_2_0.div24.n8 div120_2_0.div24.t11 336.25
R1302 div120_2_0.div24.n0 div120_2_0.div24.t3 305.267
R1303 div120_2_0.div24.n9 div120_2_0.div24.t0 257.534
R1304 div120_2_0.div24.n4 div120_2_0.div24.t6 192.8
R1305 div120_2_0.div24.n1 div120_2_0.div24.n0 176.733
R1306 div120_2_0.div24.n6 div120_2_0.div24.n5 176.733
R1307 div120_2_0.div24.n4 div120_2_0.div24.n3 160.667
R1308 div120_2_0.div24.n3 div120_2_0.div24.t13 144.601
R1309 div120_2_0.div24.n2 div120_2_0.div24.t9 131.976
R1310 div120_2_0.div24.n0 div120_2_0.div24.t12 128.534
R1311 div120_2_0.div24.n1 div120_2_0.div24.t4 128.534
R1312 div120_2_0.div24.n6 div120_2_0.div24.t8 112.468
R1313 div120_2_0.div24.n5 div120_2_0.div24.t14 112.468
R1314 div120_2_0.div24.n7 div120_2_0.div24.t7 112.468
R1315 div120_2_0.div24.n5 div120_2_0.div24.n4 96.4005
R1316 div120_2_0.div24.t2 div120_2_0.div24.n10 78.8005
R1317 div120_2_0.div24.n10 div120_2_0.div24.t1 78.8005
R1318 div120_2_0.div24.n9 div120_2_0.div24.n8 11.2005
R1319 vco2_3_0.V2.t2 vco2_3_0.V2.n0 708.125
R1320 vco2_3_0.V2.t2 vco2_3_0.V2.n1 708.125
R1321 vco2_3_0.V2.n1 vco2_3_0.V2.t1 410.519
R1322 vco2_3_0.V2.n0 vco2_3_0.V2.t0 305.649
R1323 vco2_3_0.V2.n1 vco2_3_0.V2.n0 21.3338
R1324 a_3810_770.n4 a_3810_770.t1 752.333
R1325 a_3810_770.t2 a_3810_770.n5 752.333
R1326 a_3810_770.n0 a_3810_770.t4 514.134
R1327 a_3810_770.n3 a_3810_770.n2 366.856
R1328 a_3810_770.n5 a_3810_770.t0 254.333
R1329 a_3810_770.n3 a_3810_770.t5 190.123
R1330 a_3810_770.n4 a_3810_770.n3 187.201
R1331 a_3810_770.n1 a_3810_770.n0 176.733
R1332 a_3810_770.n2 a_3810_770.n1 176.733
R1333 a_3810_770.n0 a_3810_770.t6 112.468
R1334 a_3810_770.n2 a_3810_770.t7 112.468
R1335 a_3810_770.n1 a_3810_770.t3 112.468
R1336 a_3810_770.n5 a_3810_770.n4 70.4005
R1337 div120_2_0.div2_4_1.C.n0 div120_2_0.div2_4_1.C.t0 750.201
R1338 div120_2_0.div2_4_1.C.n1 div120_2_0.div2_4_1.C.t4 349.433
R1339 div120_2_0.div2_4_1.C.n0 div120_2_0.div2_4_1.C.t1 276.733
R1340 div120_2_0.div2_4_1.C.n2 div120_2_0.div2_4_1.C.n1 206.333
R1341 div120_2_0.div2_4_1.C.n1 div120_2_0.div2_4_1.C.n0 48.0005
R1342 div120_2_0.div2_4_1.C.n2 div120_2_0.div2_4_1.C.t2 48.0005
R1343 div120_2_0.div2_4_1.C.t3 div120_2_0.div2_4_1.C.n2 48.0005
R1344 div120_2_0.div2_4_1.A.n0 div120_2_0.div2_4_1.A.t0 713.933
R1345 div120_2_0.div2_4_1.A.t1 div120_2_0.div2_4_1.A.n0 337
R1346 div120_2_0.div2_4_1.A.n0 div120_2_0.div2_4_1.A.t2 314.233
R1347 vco2_3_0.V1.n0 vco2_3_0.V1.t5 600.206
R1348 vco2_3_0.V1.n1 vco2_3_0.V1.n0 568.072
R1349 vco2_3_0.V1.n2 vco2_3_0.V1.n1 392.486
R1350 vco2_3_0.V1.n4 vco2_3_0.V1.t2 289.791
R1351 vco2_3_0.V1 vco2_3_0.V1.t0 266.399
R1352 vco2_3_0.V1.n5 vco2_3_0.V1.n2 168.067
R1353 vco2_3_0.V1 vco2_3_0.V1.n5 166.4
R1354 vco2_3_0.V1.n4 vco2_3_0.V1.n3 97.9242
R1355 vco2_3_0.V1.n3 vco2_3_0.V1.n2 37.7572
R1356 vco2_3_0.V1.n0 vco2_3_0.V1.t3 32.1338
R1357 vco2_3_0.V1.n1 vco2_3_0.V1.t4 32.1338
R1358 vco2_3_0.V1.n3 vco2_3_0.V1.t1 32.1338
R1359 vco2_3_0.V1.n5 vco2_3_0.V1.n4 28.3357
R1360 div120_2_0.div2_4_0.B.t0 div120_2_0.div2_4_0.B.t1 96.0005
R1361 div120_2_0.div5_2_0.B.n0 div120_2_0.div5_2_0.B.t1 663.801
R1362 div120_2_0.div5_2_0.B.n0 div120_2_0.div5_2_0.B.t2 348.851
R1363 div120_2_0.div5_2_0.B div120_2_0.div5_2_0.B.t0 282.921
R1364 div120_2_0.div5_2_0.B div120_2_0.div5_2_0.B.n0 114.133
R1365 div120_2_0.div5_2_0.D.n0 div120_2_0.div5_2_0.D.t0 761.4
R1366 div120_2_0.div5_2_0.D.n1 div120_2_0.div5_2_0.D.t4 350.349
R1367 div120_2_0.div5_2_0.D.n0 div120_2_0.div5_2_0.D.t2 254.333
R1368 div120_2_0.div5_2_0.D.n2 div120_2_0.div5_2_0.D.n1 206.333
R1369 div120_2_0.div5_2_0.D.n1 div120_2_0.div5_2_0.D.n0 70.4005
R1370 div120_2_0.div5_2_0.D.t3 div120_2_0.div5_2_0.D.n2 48.0005
R1371 div120_2_0.div5_2_0.D.n2 div120_2_0.div5_2_0.D.t1 48.0005
R1372 vco2_3_0.V9.n1 vco2_3_0.V9.n0 412.034
R1373 vco2_3_0.V9.t1 vco2_3_0.V9.n1 372.118
R1374 vco2_3_0.V9.n1 vco2_3_0.V9.t0 247.934
R1375 vco2_3_0.V9.n0 vco2_3_0.V9.t3 186.775
R1376 vco2_3_0.V9.n0 vco2_3_0.V9.t2 126.525
R1377 vco2_3_0.V7.n0 vco2_3_0.V7.t0 284.2
R1378 vco2_3_0.V7.n0 vco2_3_0.V7.t2 233
R1379 vco2_3_0.V7.t1 vco2_3_0.V7.n0 184.191
R1380 div120_2_0.div2_4_1.B.t0 div120_2_0.div2_4_1.B.t1 96.0005
R1381 div120_2_0.div5_2_0.C.t0 div120_2_0.div5_2_0.C.t1 96.0005
R1382 vco2_3_0.V5.n0 vco2_3_0.V5.t1 284.2
R1383 vco2_3_0.V5.n0 vco2_3_0.V5.t2 233
R1384 vco2_3_0.V5.t0 vco2_3_0.V5.n0 184.191
R1385 div120_2_0.div2_4_2.A.n0 div120_2_0.div2_4_2.A.t1 713.933
R1386 div120_2_0.div2_4_2.A.t0 div120_2_0.div2_4_2.A.n0 337
R1387 div120_2_0.div2_4_2.A.n0 div120_2_0.div2_4_2.A.t2 314.233
R1388 div120_2_0.div2_4_2.B.t0 div120_2_0.div2_4_2.B.t1 96.0005
R1389 div120_2_0.div3_3_0.D.n1 div120_2_0.div3_3_0.D.n0 701.467
R1390 div120_2_0.div3_3_0.D.n1 div120_2_0.div3_3_0.D.t1 694.201
R1391 div120_2_0.div3_3_0.D.n0 div120_2_0.div3_3_0.D.t3 321.334
R1392 div120_2_0.div3_3_0.D.t0 div120_2_0.div3_3_0.D.n1 314.921
R1393 div120_2_0.div3_3_0.D.n0 div120_2_0.div3_3_0.D.t2 144.601
R1394 V_CONT.n0 V_CONT.t2 1156.8
R1395 V_CONT.n1 V_CONT.n0 964
R1396 V_CONT V_CONT.n2 698.9
R1397 V_CONT.n2 V_CONT.n1 433.8
R1398 V_CONT.n2 V_CONT.t1 192.8
R1399 V_CONT.n1 V_CONT.t0 192.8
R1400 V_CONT.n0 V_CONT.t3 192.8
R1401 vco2_3_0.V6.t2 vco2_3_0.V6.n0 708.125
R1402 vco2_3_0.V6.t2 vco2_3_0.V6.n1 708.125
R1403 vco2_3_0.V6.n1 vco2_3_0.V6.t0 410.519
R1404 vco2_3_0.V6.n0 vco2_3_0.V6.t1 305.649
R1405 vco2_3_0.V6.n1 vco2_3_0.V6.n0 21.3338
R1406 V_OUT_120.n1 V_OUT_120.t4 772.196
R1407 V_OUT_120.n3 V_OUT_120.t1 751.801
R1408 V_OUT_120.n2 V_OUT_120.n1 607.465
R1409 V_OUT_120.t4 V_OUT_120.t5 514.134
R1410 V_OUT_120.n0 V_OUT_120.t3 289.2
R1411 V_OUT_120.n2 V_OUT_120.t0 233
R1412 V_OUT_120.n1 V_OUT_120.n0 208.868
R1413 V_OUT_120.n0 V_OUT_120.t2 176.733
R1414 V_OUT_120.n3 V_OUT_120.n2 40.3205
R1415 V_OUT_120 V_OUT_120.n3 38.4005
C0 VDDA div120_2_0.div5_2_0.B 0.506749f
C1 VDDA V_CONT 0.090679f
C2 vco2_3_0.V1 VDDA 2.67676f
C3 VDDA V_OUT_120 1.02478f
C4 vco2_3_0.V1 V_CONT 0.061609f
C5 V_CONT GNDA 1.52509f
C6 V_OUT_120 GNDA 1.85356f
C7 VDDA GNDA 25.15039f
C8 div120_2_0.div5_2_0.B GNDA 0.178977f
C9 vco2_3_0.V1 GNDA 1.923992f
C10 vco2_3_0.V1.t4 GNDA 0.287159f
C11 vco2_3_0.V1.t3 GNDA 0.287159f
C12 vco2_3_0.V1.t5 GNDA 0.478415f
C13 vco2_3_0.V1.n0 GNDA 0.234164f
C14 vco2_3_0.V1.n1 GNDA 0.209715f
C15 vco2_3_0.V1.n2 GNDA 0.043626f
C16 vco2_3_0.V1.t2 GNDA 0.100747f
C17 vco2_3_0.V1.t1 GNDA 0.287159f
C18 vco2_3_0.V1.n3 GNDA 0.162794f
C19 vco2_3_0.V1.n4 GNDA 0.177425f
C20 vco2_3_0.V1.n5 GNDA 0.12179f
C21 vco2_3_0.V1.t0 GNDA 0.101836f
C22 VDDA.n8 GNDA 0.036899f
C23 VDDA.t13 GNDA 0.022331f
C24 VDDA.t15 GNDA 0.022331f
C25 VDDA.t64 GNDA 0.026976f
C26 VDDA.t80 GNDA 0.030906f
C27 VDDA.t60 GNDA 0.026083f
C28 VDDA.t33 GNDA 0.015721f
C29 VDDA.t40 GNDA 0.015721f
C30 VDDA.t9 GNDA 0.023939f
C31 VDDA.t25 GNDA 0.023939f
C32 VDDA.t34 GNDA 0.014113f
C33 VDDA.n47 GNDA 0.013664f
C34 VDDA.n49 GNDA 0.029105f
C35 VDDA.n146 GNDA 0.013664f
C36 VDDA.t82 GNDA 0.014113f
C37 VDDA.t90 GNDA 0.016079f
C38 VDDA.t78 GNDA 0.016079f
C39 VDDA.t0 GNDA 0.012863f
C40 VDDA.t57 GNDA 0.012863f
C41 VDDA.t55 GNDA 0.020723f
C42 VDDA.t49 GNDA 0.020723f
C43 VDDA.t88 GNDA 0.015721f
C44 VDDA.t53 GNDA 0.015721f
C45 VDDA.t86 GNDA 0.022153f
C46 VDDA.t47 GNDA 0.023046f
C47 VDDA.t36 GNDA 0.021438f
C48 VDDA.t68 GNDA 0.012863f
C49 VDDA.t11 GNDA 0.012863f
C50 VDDA.t92 GNDA 0.011255f
C51 VDDA.n147 GNDA 0.010805f
C52 VDDA.n201 GNDA 0.010805f
C53 VDDA.t38 GNDA 0.011255f
C54 VDDA.t70 GNDA 0.012863f
C55 VDDA.t5 GNDA 0.012863f
C56 VDDA.t17 GNDA 0.021438f
C57 VDDA.t31 GNDA 0.022331f
C58 VDDA.t29 GNDA 0.021438f
C59 VDDA.t7 GNDA 0.012863f
C60 VDDA.t3 GNDA 0.012863f
C61 VDDA.t66 GNDA 0.011255f
C62 VDDA.n202 GNDA 0.010805f
C63 VDDA.n248 GNDA 0.010805f
C64 VDDA.t23 GNDA 0.011255f
C65 VDDA.t45 GNDA 0.012863f
C66 VDDA.t27 GNDA 0.012863f
C67 VDDA.t84 GNDA 0.019895f
C68 VDDA.t72 GNDA 0.067721f
C69 VDDA.t59 GNDA 0.026874f
C70 VDDA.t43 GNDA 0.082349f
C71 VDDA.n249 GNDA 0.035453f
C72 VDDA.n256 GNDA 0.035453f
C73 VDDA.n258 GNDA 0.036145f
C74 VDDA.t21 GNDA 0.161245f
C75 VDDA.n260 GNDA 0.013418f
C76 VDDA.n271 GNDA 0.107496f
C77 VDDA.t19 GNDA 0.082349f
C78 VDDA.t2 GNDA 0.026874f
C79 VDDA.t74 GNDA 0.039813f
C80 VDDA.n280 GNDA 0.092566f
C81 VDDA.t62 GNDA 0.082349f
C82 VDDA.t42 GNDA 0.026874f
C83 VDDA.t76 GNDA 0.039813f
C84 VDDA.n281 GNDA 0.092566f
C85 VDDA.n285 GNDA 0.049382f
C86 VDDA.n304 GNDA 0.010942f
.ends

