magic
tech sky130A
timestamp 1751430584
<< nwell >>
rect 2965 3260 3475 3595
rect 3605 3260 4555 3595
rect 4685 3265 5195 3595
rect 2645 2700 3050 3030
rect 3180 2595 4980 3130
rect 5110 2700 5510 3030
rect 2630 2110 4010 2440
rect 4150 2110 5530 2440
<< pwell >>
rect 20 3420 1240 3665
rect 20 3155 1210 3400
rect 215 2945 1025 3135
rect 1305 3045 2510 3530
rect 215 2735 1025 2925
rect 1470 2840 2305 3025
rect 3075 1800 3825 2095
rect 4335 1800 5085 2095
rect -45 1685 130 1725
rect 2835 1325 4065 1770
rect 4095 1325 5325 1770
rect 2935 1050 5220 1305
rect 4220 1030 4426 1031
rect 3060 730 3705 1030
rect 3730 730 4430 1030
rect 4455 730 5100 1030
<< nmos >>
rect 3170 1900 3190 1950
rect 3230 1900 3250 1950
rect 3290 1900 3310 1950
rect 3350 1900 3370 1950
rect 3410 1900 3430 1950
rect 3470 1900 3490 1950
rect 3530 1900 3550 1950
rect 3590 1900 3610 1950
rect 3650 1900 3670 1950
rect 3710 1900 3730 1950
rect 4430 1900 4450 1950
rect 4490 1900 4510 1950
rect 4550 1900 4570 1950
rect 4610 1900 4630 1950
rect 4670 1900 4690 1950
rect 4730 1900 4750 1950
rect 4790 1900 4810 1950
rect 4850 1900 4870 1950
rect 4910 1900 4930 1950
rect 4970 1900 4990 1950
rect 2930 1425 3430 1675
rect 3470 1425 3970 1675
rect 4190 1425 4690 1675
rect 4730 1425 5230 1675
rect 3060 1105 4060 1205
rect 4100 1105 5100 1205
rect 3155 830 3170 930
rect 3210 830 3225 930
rect 3265 830 3280 930
rect 3320 830 3335 930
rect 3375 830 3390 930
rect 3430 830 3445 930
rect 3485 830 3500 930
rect 3540 830 3555 930
rect 3595 830 3610 930
rect 3825 830 3840 930
rect 3880 830 3895 930
rect 3935 830 3950 930
rect 3990 830 4005 930
rect 4045 830 4060 930
rect 4100 830 4115 930
rect 4155 830 4170 930
rect 4210 830 4225 930
rect 4265 830 4280 930
rect 4320 830 4335 930
rect 4550 830 4565 930
rect 4605 830 4620 930
rect 4660 830 4675 930
rect 4715 830 4730 930
rect 4770 830 4785 930
rect 4825 830 4840 930
rect 4880 830 4895 930
rect 4935 830 4950 930
rect 4990 830 5005 930
<< pmos >>
rect 3075 3380 3090 3480
rect 3130 3380 3145 3480
rect 3185 3380 3200 3480
rect 3240 3380 3255 3480
rect 3295 3380 3310 3480
rect 3350 3380 3365 3480
rect 3715 3380 3730 3480
rect 3770 3380 3785 3480
rect 3825 3380 3840 3480
rect 3880 3380 3895 3480
rect 3935 3380 3950 3480
rect 3990 3380 4005 3480
rect 4045 3380 4060 3480
rect 4100 3380 4115 3480
rect 4155 3380 4170 3480
rect 4210 3380 4225 3480
rect 4265 3380 4280 3480
rect 4320 3380 4335 3480
rect 4375 3380 4390 3480
rect 4430 3380 4445 3480
rect 4795 3380 4810 3480
rect 4850 3380 4865 3480
rect 4905 3380 4920 3480
rect 4960 3380 4975 3480
rect 5015 3380 5030 3480
rect 5070 3380 5085 3480
rect 2755 2815 2770 2915
rect 2810 2815 2825 2915
rect 2865 2815 2880 2915
rect 2920 2815 2935 2915
rect 3290 2715 3340 3015
rect 3380 2715 3430 3015
rect 3470 2715 3520 3015
rect 3560 2715 3610 3015
rect 3650 2715 3700 3015
rect 3740 2715 3790 3015
rect 3830 2715 3880 3015
rect 3920 2715 3970 3015
rect 4010 2715 4060 3015
rect 4100 2715 4150 3015
rect 4190 2715 4240 3015
rect 4280 2715 4330 3015
rect 4370 2715 4420 3015
rect 4460 2715 4510 3015
rect 4550 2715 4600 3015
rect 4640 2715 4690 3015
rect 4730 2715 4780 3015
rect 4820 2715 4870 3015
rect 5220 2815 5235 2915
rect 5275 2815 5290 2915
rect 5330 2815 5345 2915
rect 5385 2815 5400 2915
rect 2740 2225 2760 2325
rect 2800 2225 2820 2325
rect 2860 2225 2880 2325
rect 2920 2225 2940 2325
rect 2980 2225 3000 2325
rect 3040 2225 3060 2325
rect 3100 2225 3120 2325
rect 3160 2225 3180 2325
rect 3220 2225 3240 2325
rect 3280 2225 3300 2325
rect 3340 2225 3360 2325
rect 3400 2225 3420 2325
rect 3460 2225 3480 2325
rect 3520 2225 3540 2325
rect 3580 2225 3600 2325
rect 3640 2225 3660 2325
rect 3700 2225 3720 2325
rect 3760 2225 3780 2325
rect 3820 2225 3840 2325
rect 3880 2225 3900 2325
rect 4260 2225 4280 2325
rect 4320 2225 4340 2325
rect 4380 2225 4400 2325
rect 4440 2225 4460 2325
rect 4500 2225 4520 2325
rect 4560 2225 4580 2325
rect 4620 2225 4640 2325
rect 4680 2225 4700 2325
rect 4740 2225 4760 2325
rect 4800 2225 4820 2325
rect 4860 2225 4880 2325
rect 4920 2225 4940 2325
rect 4980 2225 5000 2325
rect 5040 2225 5060 2325
rect 5100 2225 5120 2325
rect 5160 2225 5180 2325
rect 5220 2225 5240 2325
rect 5280 2225 5300 2325
rect 5340 2225 5360 2325
rect 5400 2225 5420 2325
<< ndiff >>
rect 3130 1935 3170 1950
rect 3130 1915 3140 1935
rect 3160 1915 3170 1935
rect 3130 1900 3170 1915
rect 3190 1935 3230 1950
rect 3190 1915 3200 1935
rect 3220 1915 3230 1935
rect 3190 1900 3230 1915
rect 3250 1935 3290 1950
rect 3250 1915 3260 1935
rect 3280 1915 3290 1935
rect 3250 1900 3290 1915
rect 3310 1935 3350 1950
rect 3310 1915 3320 1935
rect 3340 1915 3350 1935
rect 3310 1900 3350 1915
rect 3370 1935 3410 1950
rect 3370 1915 3380 1935
rect 3400 1915 3410 1935
rect 3370 1900 3410 1915
rect 3430 1935 3470 1950
rect 3430 1915 3440 1935
rect 3460 1915 3470 1935
rect 3430 1900 3470 1915
rect 3490 1935 3530 1950
rect 3490 1915 3500 1935
rect 3520 1915 3530 1935
rect 3490 1900 3530 1915
rect 3550 1935 3590 1950
rect 3550 1915 3560 1935
rect 3580 1915 3590 1935
rect 3550 1900 3590 1915
rect 3610 1935 3650 1950
rect 3610 1915 3620 1935
rect 3640 1915 3650 1935
rect 3610 1900 3650 1915
rect 3670 1935 3710 1950
rect 3670 1915 3680 1935
rect 3700 1915 3710 1935
rect 3670 1900 3710 1915
rect 3730 1935 3770 1950
rect 3730 1915 3740 1935
rect 3760 1915 3770 1935
rect 3730 1900 3770 1915
rect 4390 1935 4430 1950
rect 4390 1915 4400 1935
rect 4420 1915 4430 1935
rect 4390 1900 4430 1915
rect 4450 1935 4490 1950
rect 4450 1915 4460 1935
rect 4480 1915 4490 1935
rect 4450 1900 4490 1915
rect 4510 1935 4550 1950
rect 4510 1915 4520 1935
rect 4540 1915 4550 1935
rect 4510 1900 4550 1915
rect 4570 1935 4610 1950
rect 4570 1915 4580 1935
rect 4600 1915 4610 1935
rect 4570 1900 4610 1915
rect 4630 1935 4670 1950
rect 4630 1915 4640 1935
rect 4660 1915 4670 1935
rect 4630 1900 4670 1915
rect 4690 1935 4730 1950
rect 4690 1915 4700 1935
rect 4720 1915 4730 1935
rect 4690 1900 4730 1915
rect 4750 1935 4790 1950
rect 4750 1915 4760 1935
rect 4780 1915 4790 1935
rect 4750 1900 4790 1915
rect 4810 1935 4850 1950
rect 4810 1915 4820 1935
rect 4840 1915 4850 1935
rect 4810 1900 4850 1915
rect 4870 1935 4910 1950
rect 4870 1915 4880 1935
rect 4900 1915 4910 1935
rect 4870 1900 4910 1915
rect 4930 1935 4970 1950
rect 4930 1915 4940 1935
rect 4960 1915 4970 1935
rect 4930 1900 4970 1915
rect 4990 1935 5030 1950
rect 4990 1915 5000 1935
rect 5020 1915 5030 1935
rect 4990 1900 5030 1915
rect 2890 1660 2930 1675
rect 2890 1640 2900 1660
rect 2920 1640 2930 1660
rect 2890 1610 2930 1640
rect 2890 1590 2900 1610
rect 2920 1590 2930 1610
rect 2890 1560 2930 1590
rect 2890 1540 2900 1560
rect 2920 1540 2930 1560
rect 2890 1510 2930 1540
rect 2890 1490 2900 1510
rect 2920 1490 2930 1510
rect 2890 1460 2930 1490
rect 2890 1440 2900 1460
rect 2920 1440 2930 1460
rect 2890 1425 2930 1440
rect 3430 1660 3470 1675
rect 3430 1640 3440 1660
rect 3460 1640 3470 1660
rect 3430 1610 3470 1640
rect 3430 1590 3440 1610
rect 3460 1590 3470 1610
rect 3430 1560 3470 1590
rect 3430 1540 3440 1560
rect 3460 1540 3470 1560
rect 3430 1510 3470 1540
rect 3430 1490 3440 1510
rect 3460 1490 3470 1510
rect 3430 1460 3470 1490
rect 3430 1440 3440 1460
rect 3460 1440 3470 1460
rect 3430 1425 3470 1440
rect 3970 1660 4010 1675
rect 3970 1640 3980 1660
rect 4000 1640 4010 1660
rect 3970 1610 4010 1640
rect 3970 1590 3980 1610
rect 4000 1590 4010 1610
rect 3970 1560 4010 1590
rect 3970 1540 3980 1560
rect 4000 1540 4010 1560
rect 3970 1510 4010 1540
rect 3970 1490 3980 1510
rect 4000 1490 4010 1510
rect 3970 1460 4010 1490
rect 3970 1440 3980 1460
rect 4000 1440 4010 1460
rect 3970 1425 4010 1440
rect 4150 1660 4190 1675
rect 4150 1640 4160 1660
rect 4180 1640 4190 1660
rect 4150 1610 4190 1640
rect 4150 1590 4160 1610
rect 4180 1590 4190 1610
rect 4150 1560 4190 1590
rect 4150 1540 4160 1560
rect 4180 1540 4190 1560
rect 4150 1510 4190 1540
rect 4150 1490 4160 1510
rect 4180 1490 4190 1510
rect 4150 1460 4190 1490
rect 4150 1440 4160 1460
rect 4180 1440 4190 1460
rect 4150 1425 4190 1440
rect 4690 1660 4730 1675
rect 4690 1640 4700 1660
rect 4720 1640 4730 1660
rect 4690 1610 4730 1640
rect 4690 1590 4700 1610
rect 4720 1590 4730 1610
rect 4690 1560 4730 1590
rect 4690 1540 4700 1560
rect 4720 1540 4730 1560
rect 4690 1510 4730 1540
rect 4690 1490 4700 1510
rect 4720 1490 4730 1510
rect 4690 1460 4730 1490
rect 4690 1440 4700 1460
rect 4720 1440 4730 1460
rect 4690 1425 4730 1440
rect 5230 1660 5270 1675
rect 5230 1640 5240 1660
rect 5260 1640 5270 1660
rect 5230 1610 5270 1640
rect 5230 1590 5240 1610
rect 5260 1590 5270 1610
rect 5230 1560 5270 1590
rect 5230 1540 5240 1560
rect 5260 1540 5270 1560
rect 5230 1510 5270 1540
rect 5230 1490 5240 1510
rect 5260 1490 5270 1510
rect 5230 1460 5270 1490
rect 5230 1440 5240 1460
rect 5260 1440 5270 1460
rect 5230 1425 5270 1440
rect 3020 1190 3060 1205
rect 3020 1170 3030 1190
rect 3050 1170 3060 1190
rect 3020 1140 3060 1170
rect 3020 1120 3030 1140
rect 3050 1120 3060 1140
rect 3020 1105 3060 1120
rect 4060 1190 4100 1205
rect 4060 1170 4070 1190
rect 4090 1170 4100 1190
rect 4060 1140 4100 1170
rect 4060 1120 4070 1140
rect 4090 1120 4100 1140
rect 4060 1105 4100 1120
rect 5100 1190 5140 1205
rect 5100 1170 5110 1190
rect 5130 1170 5140 1190
rect 5100 1140 5140 1170
rect 5100 1120 5110 1140
rect 5130 1120 5140 1140
rect 5100 1105 5140 1120
rect 3115 915 3155 930
rect 3115 895 3125 915
rect 3145 895 3155 915
rect 3115 865 3155 895
rect 3115 845 3125 865
rect 3145 845 3155 865
rect 3115 830 3155 845
rect 3170 915 3210 930
rect 3170 895 3180 915
rect 3200 895 3210 915
rect 3170 865 3210 895
rect 3170 845 3180 865
rect 3200 845 3210 865
rect 3170 830 3210 845
rect 3225 915 3265 930
rect 3225 895 3235 915
rect 3255 895 3265 915
rect 3225 865 3265 895
rect 3225 845 3235 865
rect 3255 845 3265 865
rect 3225 830 3265 845
rect 3280 915 3320 930
rect 3280 895 3290 915
rect 3310 895 3320 915
rect 3280 865 3320 895
rect 3280 845 3290 865
rect 3310 845 3320 865
rect 3280 830 3320 845
rect 3335 915 3375 930
rect 3335 895 3345 915
rect 3365 895 3375 915
rect 3335 865 3375 895
rect 3335 845 3345 865
rect 3365 845 3375 865
rect 3335 830 3375 845
rect 3390 915 3430 930
rect 3390 895 3400 915
rect 3420 895 3430 915
rect 3390 865 3430 895
rect 3390 845 3400 865
rect 3420 845 3430 865
rect 3390 830 3430 845
rect 3445 915 3485 930
rect 3445 895 3455 915
rect 3475 895 3485 915
rect 3445 865 3485 895
rect 3445 845 3455 865
rect 3475 845 3485 865
rect 3445 830 3485 845
rect 3500 915 3540 930
rect 3500 895 3510 915
rect 3530 895 3540 915
rect 3500 865 3540 895
rect 3500 845 3510 865
rect 3530 845 3540 865
rect 3500 830 3540 845
rect 3555 915 3595 930
rect 3555 895 3565 915
rect 3585 895 3595 915
rect 3555 865 3595 895
rect 3555 845 3565 865
rect 3585 845 3595 865
rect 3555 830 3595 845
rect 3610 915 3650 930
rect 3610 895 3620 915
rect 3640 895 3650 915
rect 3610 865 3650 895
rect 3610 845 3620 865
rect 3640 845 3650 865
rect 3610 830 3650 845
rect 3785 915 3825 930
rect 3785 895 3795 915
rect 3815 895 3825 915
rect 3785 865 3825 895
rect 3785 845 3795 865
rect 3815 845 3825 865
rect 3785 830 3825 845
rect 3840 915 3880 930
rect 3840 895 3850 915
rect 3870 895 3880 915
rect 3840 865 3880 895
rect 3840 845 3850 865
rect 3870 845 3880 865
rect 3840 830 3880 845
rect 3895 915 3935 930
rect 3895 895 3905 915
rect 3925 895 3935 915
rect 3895 865 3935 895
rect 3895 845 3905 865
rect 3925 845 3935 865
rect 3895 830 3935 845
rect 3950 915 3990 930
rect 3950 895 3960 915
rect 3980 895 3990 915
rect 3950 865 3990 895
rect 3950 845 3960 865
rect 3980 845 3990 865
rect 3950 830 3990 845
rect 4005 915 4045 930
rect 4005 895 4015 915
rect 4035 895 4045 915
rect 4005 865 4045 895
rect 4005 845 4015 865
rect 4035 845 4045 865
rect 4005 830 4045 845
rect 4060 915 4100 930
rect 4060 895 4070 915
rect 4090 895 4100 915
rect 4060 865 4100 895
rect 4060 845 4070 865
rect 4090 845 4100 865
rect 4060 830 4100 845
rect 4115 915 4155 930
rect 4115 895 4125 915
rect 4145 895 4155 915
rect 4115 865 4155 895
rect 4115 845 4125 865
rect 4145 845 4155 865
rect 4115 830 4155 845
rect 4170 915 4210 930
rect 4170 895 4180 915
rect 4200 895 4210 915
rect 4170 865 4210 895
rect 4170 845 4180 865
rect 4200 845 4210 865
rect 4170 830 4210 845
rect 4225 915 4265 930
rect 4225 895 4235 915
rect 4255 895 4265 915
rect 4225 865 4265 895
rect 4225 845 4235 865
rect 4255 845 4265 865
rect 4225 830 4265 845
rect 4280 915 4320 930
rect 4280 895 4290 915
rect 4310 895 4320 915
rect 4280 865 4320 895
rect 4280 845 4290 865
rect 4310 845 4320 865
rect 4280 830 4320 845
rect 4335 915 4375 930
rect 4335 895 4345 915
rect 4365 895 4375 915
rect 4335 865 4375 895
rect 4335 845 4345 865
rect 4365 845 4375 865
rect 4335 830 4375 845
rect 4510 915 4550 930
rect 4510 895 4520 915
rect 4540 895 4550 915
rect 4510 865 4550 895
rect 4510 845 4520 865
rect 4540 845 4550 865
rect 4510 830 4550 845
rect 4565 915 4605 930
rect 4565 895 4575 915
rect 4595 895 4605 915
rect 4565 865 4605 895
rect 4565 845 4575 865
rect 4595 845 4605 865
rect 4565 830 4605 845
rect 4620 915 4660 930
rect 4620 895 4630 915
rect 4650 895 4660 915
rect 4620 865 4660 895
rect 4620 845 4630 865
rect 4650 845 4660 865
rect 4620 830 4660 845
rect 4675 915 4715 930
rect 4675 895 4685 915
rect 4705 895 4715 915
rect 4675 865 4715 895
rect 4675 845 4685 865
rect 4705 845 4715 865
rect 4675 830 4715 845
rect 4730 915 4770 930
rect 4730 895 4740 915
rect 4760 895 4770 915
rect 4730 865 4770 895
rect 4730 845 4740 865
rect 4760 845 4770 865
rect 4730 830 4770 845
rect 4785 915 4825 930
rect 4785 895 4795 915
rect 4815 895 4825 915
rect 4785 865 4825 895
rect 4785 845 4795 865
rect 4815 845 4825 865
rect 4785 830 4825 845
rect 4840 915 4880 930
rect 4840 895 4850 915
rect 4870 895 4880 915
rect 4840 865 4880 895
rect 4840 845 4850 865
rect 4870 845 4880 865
rect 4840 830 4880 845
rect 4895 915 4935 930
rect 4895 895 4905 915
rect 4925 895 4935 915
rect 4895 865 4935 895
rect 4895 845 4905 865
rect 4925 845 4935 865
rect 4895 830 4935 845
rect 4950 915 4990 930
rect 4950 895 4960 915
rect 4980 895 4990 915
rect 4950 865 4990 895
rect 4950 845 4960 865
rect 4980 845 4990 865
rect 4950 830 4990 845
rect 5005 915 5045 930
rect 5005 895 5015 915
rect 5035 895 5045 915
rect 5005 865 5045 895
rect 5005 845 5015 865
rect 5035 845 5045 865
rect 5005 830 5045 845
<< pdiff >>
rect 3035 3465 3075 3480
rect 3035 3393 3045 3465
rect 3065 3393 3075 3465
rect 3035 3380 3075 3393
rect 3090 3465 3130 3480
rect 3090 3393 3100 3465
rect 3120 3393 3130 3465
rect 3090 3380 3130 3393
rect 3145 3465 3185 3480
rect 3145 3393 3155 3465
rect 3175 3393 3185 3465
rect 3145 3380 3185 3393
rect 3200 3465 3240 3480
rect 3200 3393 3210 3465
rect 3230 3393 3240 3465
rect 3200 3380 3240 3393
rect 3255 3465 3295 3480
rect 3255 3393 3265 3465
rect 3285 3393 3295 3465
rect 3255 3380 3295 3393
rect 3310 3465 3350 3480
rect 3310 3393 3320 3465
rect 3340 3393 3350 3465
rect 3310 3380 3350 3393
rect 3365 3465 3405 3480
rect 3365 3393 3375 3465
rect 3395 3393 3405 3465
rect 3365 3380 3405 3393
rect 3675 3465 3715 3480
rect 3675 3445 3685 3465
rect 3705 3445 3715 3465
rect 3675 3415 3715 3445
rect 3675 3395 3685 3415
rect 3705 3395 3715 3415
rect 3675 3380 3715 3395
rect 3730 3465 3770 3480
rect 3730 3445 3740 3465
rect 3760 3445 3770 3465
rect 3730 3415 3770 3445
rect 3730 3395 3740 3415
rect 3760 3395 3770 3415
rect 3730 3380 3770 3395
rect 3785 3465 3825 3480
rect 3785 3445 3795 3465
rect 3815 3445 3825 3465
rect 3785 3415 3825 3445
rect 3785 3395 3795 3415
rect 3815 3395 3825 3415
rect 3785 3380 3825 3395
rect 3840 3465 3880 3480
rect 3840 3445 3850 3465
rect 3870 3445 3880 3465
rect 3840 3415 3880 3445
rect 3840 3395 3850 3415
rect 3870 3395 3880 3415
rect 3840 3380 3880 3395
rect 3895 3465 3935 3480
rect 3895 3445 3905 3465
rect 3925 3445 3935 3465
rect 3895 3415 3935 3445
rect 3895 3395 3905 3415
rect 3925 3395 3935 3415
rect 3895 3380 3935 3395
rect 3950 3465 3990 3480
rect 3950 3445 3960 3465
rect 3980 3445 3990 3465
rect 3950 3415 3990 3445
rect 3950 3395 3960 3415
rect 3980 3395 3990 3415
rect 3950 3380 3990 3395
rect 4005 3465 4045 3480
rect 4005 3445 4015 3465
rect 4035 3445 4045 3465
rect 4005 3415 4045 3445
rect 4005 3395 4015 3415
rect 4035 3395 4045 3415
rect 4005 3380 4045 3395
rect 4060 3465 4100 3480
rect 4060 3445 4070 3465
rect 4090 3445 4100 3465
rect 4060 3415 4100 3445
rect 4060 3395 4070 3415
rect 4090 3395 4100 3415
rect 4060 3380 4100 3395
rect 4115 3465 4155 3480
rect 4115 3445 4125 3465
rect 4145 3445 4155 3465
rect 4115 3415 4155 3445
rect 4115 3395 4125 3415
rect 4145 3395 4155 3415
rect 4115 3380 4155 3395
rect 4170 3465 4210 3480
rect 4170 3445 4180 3465
rect 4200 3445 4210 3465
rect 4170 3415 4210 3445
rect 4170 3395 4180 3415
rect 4200 3395 4210 3415
rect 4170 3380 4210 3395
rect 4225 3465 4265 3480
rect 4225 3445 4235 3465
rect 4255 3445 4265 3465
rect 4225 3415 4265 3445
rect 4225 3395 4235 3415
rect 4255 3395 4265 3415
rect 4225 3380 4265 3395
rect 4280 3465 4320 3480
rect 4280 3445 4290 3465
rect 4310 3445 4320 3465
rect 4280 3415 4320 3445
rect 4280 3395 4290 3415
rect 4310 3395 4320 3415
rect 4280 3380 4320 3395
rect 4335 3465 4375 3480
rect 4335 3445 4345 3465
rect 4365 3445 4375 3465
rect 4335 3415 4375 3445
rect 4335 3395 4345 3415
rect 4365 3395 4375 3415
rect 4335 3380 4375 3395
rect 4390 3465 4430 3480
rect 4390 3445 4400 3465
rect 4420 3445 4430 3465
rect 4390 3415 4430 3445
rect 4390 3395 4400 3415
rect 4420 3395 4430 3415
rect 4390 3380 4430 3395
rect 4445 3465 4485 3480
rect 4445 3445 4455 3465
rect 4475 3445 4485 3465
rect 4445 3415 4485 3445
rect 4445 3395 4455 3415
rect 4475 3395 4485 3415
rect 4445 3380 4485 3395
rect 4755 3465 4795 3480
rect 4755 3395 4765 3465
rect 4785 3395 4795 3465
rect 4755 3380 4795 3395
rect 4810 3465 4850 3480
rect 4810 3395 4820 3465
rect 4840 3395 4850 3465
rect 4810 3380 4850 3395
rect 4865 3465 4905 3480
rect 4865 3395 4875 3465
rect 4895 3395 4905 3465
rect 4865 3380 4905 3395
rect 4920 3465 4960 3480
rect 4920 3395 4930 3465
rect 4950 3395 4960 3465
rect 4920 3380 4960 3395
rect 4975 3465 5015 3480
rect 4975 3395 4985 3465
rect 5005 3395 5015 3465
rect 4975 3380 5015 3395
rect 5030 3465 5070 3480
rect 5030 3395 5040 3465
rect 5060 3395 5070 3465
rect 5030 3380 5070 3395
rect 5085 3465 5125 3480
rect 5085 3395 5095 3465
rect 5115 3395 5125 3465
rect 5085 3380 5125 3395
rect 2715 2900 2755 2915
rect 2715 2880 2725 2900
rect 2745 2880 2755 2900
rect 2715 2850 2755 2880
rect 2715 2830 2725 2850
rect 2745 2830 2755 2850
rect 2715 2815 2755 2830
rect 2770 2900 2810 2915
rect 2770 2880 2780 2900
rect 2800 2880 2810 2900
rect 2770 2850 2810 2880
rect 2770 2830 2780 2850
rect 2800 2830 2810 2850
rect 2770 2815 2810 2830
rect 2825 2900 2865 2915
rect 2825 2880 2835 2900
rect 2855 2880 2865 2900
rect 2825 2850 2865 2880
rect 2825 2830 2835 2850
rect 2855 2830 2865 2850
rect 2825 2815 2865 2830
rect 2880 2900 2920 2915
rect 2880 2880 2890 2900
rect 2910 2880 2920 2900
rect 2880 2850 2920 2880
rect 2880 2830 2890 2850
rect 2910 2830 2920 2850
rect 2880 2815 2920 2830
rect 2935 2900 2975 2915
rect 2935 2880 2945 2900
rect 2965 2880 2975 2900
rect 2935 2850 2975 2880
rect 2935 2830 2945 2850
rect 2965 2830 2975 2850
rect 2935 2815 2975 2830
rect 3250 3000 3290 3015
rect 3250 2980 3260 3000
rect 3280 2980 3290 3000
rect 3250 2950 3290 2980
rect 3250 2930 3260 2950
rect 3280 2930 3290 2950
rect 3250 2900 3290 2930
rect 3250 2880 3260 2900
rect 3280 2880 3290 2900
rect 3250 2850 3290 2880
rect 3250 2830 3260 2850
rect 3280 2830 3290 2850
rect 3250 2800 3290 2830
rect 3250 2780 3260 2800
rect 3280 2780 3290 2800
rect 3250 2750 3290 2780
rect 3250 2730 3260 2750
rect 3280 2730 3290 2750
rect 3250 2715 3290 2730
rect 3340 3000 3380 3015
rect 3340 2980 3350 3000
rect 3370 2980 3380 3000
rect 3340 2950 3380 2980
rect 3340 2930 3350 2950
rect 3370 2930 3380 2950
rect 3340 2900 3380 2930
rect 3340 2880 3350 2900
rect 3370 2880 3380 2900
rect 3340 2850 3380 2880
rect 3340 2830 3350 2850
rect 3370 2830 3380 2850
rect 3340 2800 3380 2830
rect 3340 2780 3350 2800
rect 3370 2780 3380 2800
rect 3340 2750 3380 2780
rect 3340 2730 3350 2750
rect 3370 2730 3380 2750
rect 3340 2715 3380 2730
rect 3430 3000 3470 3015
rect 3430 2980 3440 3000
rect 3460 2980 3470 3000
rect 3430 2950 3470 2980
rect 3430 2930 3440 2950
rect 3460 2930 3470 2950
rect 3430 2900 3470 2930
rect 3430 2880 3440 2900
rect 3460 2880 3470 2900
rect 3430 2850 3470 2880
rect 3430 2830 3440 2850
rect 3460 2830 3470 2850
rect 3430 2800 3470 2830
rect 3430 2780 3440 2800
rect 3460 2780 3470 2800
rect 3430 2750 3470 2780
rect 3430 2730 3440 2750
rect 3460 2730 3470 2750
rect 3430 2715 3470 2730
rect 3520 3000 3560 3015
rect 3520 2980 3530 3000
rect 3550 2980 3560 3000
rect 3520 2950 3560 2980
rect 3520 2930 3530 2950
rect 3550 2930 3560 2950
rect 3520 2900 3560 2930
rect 3520 2880 3530 2900
rect 3550 2880 3560 2900
rect 3520 2850 3560 2880
rect 3520 2830 3530 2850
rect 3550 2830 3560 2850
rect 3520 2800 3560 2830
rect 3520 2780 3530 2800
rect 3550 2780 3560 2800
rect 3520 2750 3560 2780
rect 3520 2730 3530 2750
rect 3550 2730 3560 2750
rect 3520 2715 3560 2730
rect 3610 3000 3650 3015
rect 3610 2980 3620 3000
rect 3640 2980 3650 3000
rect 3610 2950 3650 2980
rect 3610 2930 3620 2950
rect 3640 2930 3650 2950
rect 3610 2900 3650 2930
rect 3610 2880 3620 2900
rect 3640 2880 3650 2900
rect 3610 2850 3650 2880
rect 3610 2830 3620 2850
rect 3640 2830 3650 2850
rect 3610 2800 3650 2830
rect 3610 2780 3620 2800
rect 3640 2780 3650 2800
rect 3610 2750 3650 2780
rect 3610 2730 3620 2750
rect 3640 2730 3650 2750
rect 3610 2715 3650 2730
rect 3700 3000 3740 3015
rect 3700 2980 3710 3000
rect 3730 2980 3740 3000
rect 3700 2950 3740 2980
rect 3700 2930 3710 2950
rect 3730 2930 3740 2950
rect 3700 2900 3740 2930
rect 3700 2880 3710 2900
rect 3730 2880 3740 2900
rect 3700 2850 3740 2880
rect 3700 2830 3710 2850
rect 3730 2830 3740 2850
rect 3700 2800 3740 2830
rect 3700 2780 3710 2800
rect 3730 2780 3740 2800
rect 3700 2750 3740 2780
rect 3700 2730 3710 2750
rect 3730 2730 3740 2750
rect 3700 2715 3740 2730
rect 3790 3000 3830 3015
rect 3790 2980 3800 3000
rect 3820 2980 3830 3000
rect 3790 2950 3830 2980
rect 3790 2930 3800 2950
rect 3820 2930 3830 2950
rect 3790 2900 3830 2930
rect 3790 2880 3800 2900
rect 3820 2880 3830 2900
rect 3790 2850 3830 2880
rect 3790 2830 3800 2850
rect 3820 2830 3830 2850
rect 3790 2800 3830 2830
rect 3790 2780 3800 2800
rect 3820 2780 3830 2800
rect 3790 2750 3830 2780
rect 3790 2730 3800 2750
rect 3820 2730 3830 2750
rect 3790 2715 3830 2730
rect 3880 3000 3920 3015
rect 3880 2980 3890 3000
rect 3910 2980 3920 3000
rect 3880 2950 3920 2980
rect 3880 2930 3890 2950
rect 3910 2930 3920 2950
rect 3880 2900 3920 2930
rect 3880 2880 3890 2900
rect 3910 2880 3920 2900
rect 3880 2850 3920 2880
rect 3880 2830 3890 2850
rect 3910 2830 3920 2850
rect 3880 2800 3920 2830
rect 3880 2780 3890 2800
rect 3910 2780 3920 2800
rect 3880 2750 3920 2780
rect 3880 2730 3890 2750
rect 3910 2730 3920 2750
rect 3880 2715 3920 2730
rect 3970 3000 4010 3015
rect 3970 2980 3980 3000
rect 4000 2980 4010 3000
rect 3970 2950 4010 2980
rect 3970 2930 3980 2950
rect 4000 2930 4010 2950
rect 3970 2900 4010 2930
rect 3970 2880 3980 2900
rect 4000 2880 4010 2900
rect 3970 2850 4010 2880
rect 3970 2830 3980 2850
rect 4000 2830 4010 2850
rect 3970 2800 4010 2830
rect 3970 2780 3980 2800
rect 4000 2780 4010 2800
rect 3970 2750 4010 2780
rect 3970 2730 3980 2750
rect 4000 2730 4010 2750
rect 3970 2715 4010 2730
rect 4060 3000 4100 3015
rect 4060 2980 4070 3000
rect 4090 2980 4100 3000
rect 4060 2950 4100 2980
rect 4060 2930 4070 2950
rect 4090 2930 4100 2950
rect 4060 2900 4100 2930
rect 4060 2880 4070 2900
rect 4090 2880 4100 2900
rect 4060 2850 4100 2880
rect 4060 2830 4070 2850
rect 4090 2830 4100 2850
rect 4060 2800 4100 2830
rect 4060 2780 4070 2800
rect 4090 2780 4100 2800
rect 4060 2750 4100 2780
rect 4060 2730 4070 2750
rect 4090 2730 4100 2750
rect 4060 2715 4100 2730
rect 4150 3000 4190 3015
rect 4150 2980 4160 3000
rect 4180 2980 4190 3000
rect 4150 2950 4190 2980
rect 4150 2930 4160 2950
rect 4180 2930 4190 2950
rect 4150 2900 4190 2930
rect 4150 2880 4160 2900
rect 4180 2880 4190 2900
rect 4150 2850 4190 2880
rect 4150 2830 4160 2850
rect 4180 2830 4190 2850
rect 4150 2800 4190 2830
rect 4150 2780 4160 2800
rect 4180 2780 4190 2800
rect 4150 2750 4190 2780
rect 4150 2730 4160 2750
rect 4180 2730 4190 2750
rect 4150 2715 4190 2730
rect 4240 3000 4280 3015
rect 4240 2980 4250 3000
rect 4270 2980 4280 3000
rect 4240 2950 4280 2980
rect 4240 2930 4250 2950
rect 4270 2930 4280 2950
rect 4240 2900 4280 2930
rect 4240 2880 4250 2900
rect 4270 2880 4280 2900
rect 4240 2850 4280 2880
rect 4240 2830 4250 2850
rect 4270 2830 4280 2850
rect 4240 2800 4280 2830
rect 4240 2780 4250 2800
rect 4270 2780 4280 2800
rect 4240 2750 4280 2780
rect 4240 2730 4250 2750
rect 4270 2730 4280 2750
rect 4240 2715 4280 2730
rect 4330 3000 4370 3015
rect 4330 2980 4340 3000
rect 4360 2980 4370 3000
rect 4330 2950 4370 2980
rect 4330 2930 4340 2950
rect 4360 2930 4370 2950
rect 4330 2900 4370 2930
rect 4330 2880 4340 2900
rect 4360 2880 4370 2900
rect 4330 2850 4370 2880
rect 4330 2830 4340 2850
rect 4360 2830 4370 2850
rect 4330 2800 4370 2830
rect 4330 2780 4340 2800
rect 4360 2780 4370 2800
rect 4330 2750 4370 2780
rect 4330 2730 4340 2750
rect 4360 2730 4370 2750
rect 4330 2715 4370 2730
rect 4420 3000 4460 3015
rect 4420 2980 4430 3000
rect 4450 2980 4460 3000
rect 4420 2950 4460 2980
rect 4420 2930 4430 2950
rect 4450 2930 4460 2950
rect 4420 2900 4460 2930
rect 4420 2880 4430 2900
rect 4450 2880 4460 2900
rect 4420 2850 4460 2880
rect 4420 2830 4430 2850
rect 4450 2830 4460 2850
rect 4420 2800 4460 2830
rect 4420 2780 4430 2800
rect 4450 2780 4460 2800
rect 4420 2750 4460 2780
rect 4420 2730 4430 2750
rect 4450 2730 4460 2750
rect 4420 2715 4460 2730
rect 4510 3000 4550 3015
rect 4510 2980 4520 3000
rect 4540 2980 4550 3000
rect 4510 2950 4550 2980
rect 4510 2930 4520 2950
rect 4540 2930 4550 2950
rect 4510 2900 4550 2930
rect 4510 2880 4520 2900
rect 4540 2880 4550 2900
rect 4510 2850 4550 2880
rect 4510 2830 4520 2850
rect 4540 2830 4550 2850
rect 4510 2800 4550 2830
rect 4510 2780 4520 2800
rect 4540 2780 4550 2800
rect 4510 2750 4550 2780
rect 4510 2730 4520 2750
rect 4540 2730 4550 2750
rect 4510 2715 4550 2730
rect 4600 3000 4640 3015
rect 4600 2980 4610 3000
rect 4630 2980 4640 3000
rect 4600 2950 4640 2980
rect 4600 2930 4610 2950
rect 4630 2930 4640 2950
rect 4600 2900 4640 2930
rect 4600 2880 4610 2900
rect 4630 2880 4640 2900
rect 4600 2850 4640 2880
rect 4600 2830 4610 2850
rect 4630 2830 4640 2850
rect 4600 2800 4640 2830
rect 4600 2780 4610 2800
rect 4630 2780 4640 2800
rect 4600 2750 4640 2780
rect 4600 2730 4610 2750
rect 4630 2730 4640 2750
rect 4600 2715 4640 2730
rect 4690 3000 4730 3015
rect 4690 2980 4700 3000
rect 4720 2980 4730 3000
rect 4690 2950 4730 2980
rect 4690 2930 4700 2950
rect 4720 2930 4730 2950
rect 4690 2900 4730 2930
rect 4690 2880 4700 2900
rect 4720 2880 4730 2900
rect 4690 2850 4730 2880
rect 4690 2830 4700 2850
rect 4720 2830 4730 2850
rect 4690 2800 4730 2830
rect 4690 2780 4700 2800
rect 4720 2780 4730 2800
rect 4690 2750 4730 2780
rect 4690 2730 4700 2750
rect 4720 2730 4730 2750
rect 4690 2715 4730 2730
rect 4780 3000 4820 3015
rect 4780 2980 4790 3000
rect 4810 2980 4820 3000
rect 4780 2950 4820 2980
rect 4780 2930 4790 2950
rect 4810 2930 4820 2950
rect 4780 2900 4820 2930
rect 4780 2880 4790 2900
rect 4810 2880 4820 2900
rect 4780 2850 4820 2880
rect 4780 2830 4790 2850
rect 4810 2830 4820 2850
rect 4780 2800 4820 2830
rect 4780 2780 4790 2800
rect 4810 2780 4820 2800
rect 4780 2750 4820 2780
rect 4780 2730 4790 2750
rect 4810 2730 4820 2750
rect 4780 2715 4820 2730
rect 4870 3000 4910 3015
rect 4870 2980 4880 3000
rect 4900 2980 4910 3000
rect 4870 2950 4910 2980
rect 4870 2930 4880 2950
rect 4900 2930 4910 2950
rect 4870 2900 4910 2930
rect 4870 2880 4880 2900
rect 4900 2880 4910 2900
rect 4870 2850 4910 2880
rect 4870 2830 4880 2850
rect 4900 2830 4910 2850
rect 4870 2800 4910 2830
rect 4870 2780 4880 2800
rect 4900 2780 4910 2800
rect 4870 2750 4910 2780
rect 4870 2730 4880 2750
rect 4900 2730 4910 2750
rect 4870 2715 4910 2730
rect 5180 2900 5220 2915
rect 5180 2880 5190 2900
rect 5210 2880 5220 2900
rect 5180 2850 5220 2880
rect 5180 2830 5190 2850
rect 5210 2830 5220 2850
rect 5180 2815 5220 2830
rect 5235 2900 5275 2915
rect 5235 2880 5245 2900
rect 5265 2880 5275 2900
rect 5235 2850 5275 2880
rect 5235 2830 5245 2850
rect 5265 2830 5275 2850
rect 5235 2815 5275 2830
rect 5290 2900 5330 2915
rect 5290 2880 5300 2900
rect 5320 2880 5330 2900
rect 5290 2850 5330 2880
rect 5290 2830 5300 2850
rect 5320 2830 5330 2850
rect 5290 2815 5330 2830
rect 5345 2900 5385 2915
rect 5345 2880 5355 2900
rect 5375 2880 5385 2900
rect 5345 2850 5385 2880
rect 5345 2830 5355 2850
rect 5375 2830 5385 2850
rect 5345 2815 5385 2830
rect 5400 2900 5440 2915
rect 5400 2880 5410 2900
rect 5430 2880 5440 2900
rect 5400 2850 5440 2880
rect 5400 2830 5410 2850
rect 5430 2830 5440 2850
rect 5400 2815 5440 2830
rect 2700 2310 2740 2325
rect 2700 2290 2710 2310
rect 2730 2290 2740 2310
rect 2700 2260 2740 2290
rect 2700 2240 2710 2260
rect 2730 2240 2740 2260
rect 2700 2225 2740 2240
rect 2760 2310 2800 2325
rect 2760 2290 2770 2310
rect 2790 2290 2800 2310
rect 2760 2260 2800 2290
rect 2760 2240 2770 2260
rect 2790 2240 2800 2260
rect 2760 2225 2800 2240
rect 2820 2310 2860 2325
rect 2820 2290 2830 2310
rect 2850 2290 2860 2310
rect 2820 2260 2860 2290
rect 2820 2240 2830 2260
rect 2850 2240 2860 2260
rect 2820 2225 2860 2240
rect 2880 2310 2920 2325
rect 2880 2290 2890 2310
rect 2910 2290 2920 2310
rect 2880 2260 2920 2290
rect 2880 2240 2890 2260
rect 2910 2240 2920 2260
rect 2880 2225 2920 2240
rect 2940 2310 2980 2325
rect 2940 2290 2950 2310
rect 2970 2290 2980 2310
rect 2940 2260 2980 2290
rect 2940 2240 2950 2260
rect 2970 2240 2980 2260
rect 2940 2225 2980 2240
rect 3000 2310 3040 2325
rect 3000 2290 3010 2310
rect 3030 2290 3040 2310
rect 3000 2260 3040 2290
rect 3000 2240 3010 2260
rect 3030 2240 3040 2260
rect 3000 2225 3040 2240
rect 3060 2310 3100 2325
rect 3060 2290 3070 2310
rect 3090 2290 3100 2310
rect 3060 2260 3100 2290
rect 3060 2240 3070 2260
rect 3090 2240 3100 2260
rect 3060 2225 3100 2240
rect 3120 2310 3160 2325
rect 3120 2290 3130 2310
rect 3150 2290 3160 2310
rect 3120 2260 3160 2290
rect 3120 2240 3130 2260
rect 3150 2240 3160 2260
rect 3120 2225 3160 2240
rect 3180 2310 3220 2325
rect 3180 2290 3190 2310
rect 3210 2290 3220 2310
rect 3180 2260 3220 2290
rect 3180 2240 3190 2260
rect 3210 2240 3220 2260
rect 3180 2225 3220 2240
rect 3240 2310 3280 2325
rect 3240 2290 3250 2310
rect 3270 2290 3280 2310
rect 3240 2260 3280 2290
rect 3240 2240 3250 2260
rect 3270 2240 3280 2260
rect 3240 2225 3280 2240
rect 3300 2310 3340 2325
rect 3300 2290 3310 2310
rect 3330 2290 3340 2310
rect 3300 2260 3340 2290
rect 3300 2240 3310 2260
rect 3330 2240 3340 2260
rect 3300 2225 3340 2240
rect 3360 2310 3400 2325
rect 3360 2290 3370 2310
rect 3390 2290 3400 2310
rect 3360 2260 3400 2290
rect 3360 2240 3370 2260
rect 3390 2240 3400 2260
rect 3360 2225 3400 2240
rect 3420 2310 3460 2325
rect 3420 2290 3430 2310
rect 3450 2290 3460 2310
rect 3420 2260 3460 2290
rect 3420 2240 3430 2260
rect 3450 2240 3460 2260
rect 3420 2225 3460 2240
rect 3480 2310 3520 2325
rect 3480 2290 3490 2310
rect 3510 2290 3520 2310
rect 3480 2260 3520 2290
rect 3480 2240 3490 2260
rect 3510 2240 3520 2260
rect 3480 2225 3520 2240
rect 3540 2310 3580 2325
rect 3540 2290 3550 2310
rect 3570 2290 3580 2310
rect 3540 2260 3580 2290
rect 3540 2240 3550 2260
rect 3570 2240 3580 2260
rect 3540 2225 3580 2240
rect 3600 2310 3640 2325
rect 3600 2290 3610 2310
rect 3630 2290 3640 2310
rect 3600 2260 3640 2290
rect 3600 2240 3610 2260
rect 3630 2240 3640 2260
rect 3600 2225 3640 2240
rect 3660 2310 3700 2325
rect 3660 2290 3670 2310
rect 3690 2290 3700 2310
rect 3660 2260 3700 2290
rect 3660 2240 3670 2260
rect 3690 2240 3700 2260
rect 3660 2225 3700 2240
rect 3720 2310 3760 2325
rect 3720 2290 3730 2310
rect 3750 2290 3760 2310
rect 3720 2260 3760 2290
rect 3720 2240 3730 2260
rect 3750 2240 3760 2260
rect 3720 2225 3760 2240
rect 3780 2310 3820 2325
rect 3780 2290 3790 2310
rect 3810 2290 3820 2310
rect 3780 2260 3820 2290
rect 3780 2240 3790 2260
rect 3810 2240 3820 2260
rect 3780 2225 3820 2240
rect 3840 2310 3880 2325
rect 3840 2290 3850 2310
rect 3870 2290 3880 2310
rect 3840 2260 3880 2290
rect 3840 2240 3850 2260
rect 3870 2240 3880 2260
rect 3840 2225 3880 2240
rect 3900 2310 3940 2325
rect 3900 2290 3910 2310
rect 3930 2290 3940 2310
rect 3900 2260 3940 2290
rect 3900 2240 3910 2260
rect 3930 2240 3940 2260
rect 3900 2225 3940 2240
rect 4220 2310 4260 2325
rect 4220 2290 4230 2310
rect 4250 2290 4260 2310
rect 4220 2260 4260 2290
rect 4220 2240 4230 2260
rect 4250 2240 4260 2260
rect 4220 2225 4260 2240
rect 4280 2310 4320 2325
rect 4280 2290 4290 2310
rect 4310 2290 4320 2310
rect 4280 2260 4320 2290
rect 4280 2240 4290 2260
rect 4310 2240 4320 2260
rect 4280 2225 4320 2240
rect 4340 2310 4380 2325
rect 4340 2290 4350 2310
rect 4370 2290 4380 2310
rect 4340 2260 4380 2290
rect 4340 2240 4350 2260
rect 4370 2240 4380 2260
rect 4340 2225 4380 2240
rect 4400 2310 4440 2325
rect 4400 2290 4410 2310
rect 4430 2290 4440 2310
rect 4400 2260 4440 2290
rect 4400 2240 4410 2260
rect 4430 2240 4440 2260
rect 4400 2225 4440 2240
rect 4460 2310 4500 2325
rect 4460 2290 4470 2310
rect 4490 2290 4500 2310
rect 4460 2260 4500 2290
rect 4460 2240 4470 2260
rect 4490 2240 4500 2260
rect 4460 2225 4500 2240
rect 4520 2310 4560 2325
rect 4520 2290 4530 2310
rect 4550 2290 4560 2310
rect 4520 2260 4560 2290
rect 4520 2240 4530 2260
rect 4550 2240 4560 2260
rect 4520 2225 4560 2240
rect 4580 2310 4620 2325
rect 4580 2290 4590 2310
rect 4610 2290 4620 2310
rect 4580 2260 4620 2290
rect 4580 2240 4590 2260
rect 4610 2240 4620 2260
rect 4580 2225 4620 2240
rect 4640 2310 4680 2325
rect 4640 2290 4650 2310
rect 4670 2290 4680 2310
rect 4640 2260 4680 2290
rect 4640 2240 4650 2260
rect 4670 2240 4680 2260
rect 4640 2225 4680 2240
rect 4700 2310 4740 2325
rect 4700 2290 4710 2310
rect 4730 2290 4740 2310
rect 4700 2260 4740 2290
rect 4700 2240 4710 2260
rect 4730 2240 4740 2260
rect 4700 2225 4740 2240
rect 4760 2310 4800 2325
rect 4760 2290 4770 2310
rect 4790 2290 4800 2310
rect 4760 2260 4800 2290
rect 4760 2240 4770 2260
rect 4790 2240 4800 2260
rect 4760 2225 4800 2240
rect 4820 2310 4860 2325
rect 4820 2290 4830 2310
rect 4850 2290 4860 2310
rect 4820 2260 4860 2290
rect 4820 2240 4830 2260
rect 4850 2240 4860 2260
rect 4820 2225 4860 2240
rect 4880 2310 4920 2325
rect 4880 2290 4890 2310
rect 4910 2290 4920 2310
rect 4880 2260 4920 2290
rect 4880 2240 4890 2260
rect 4910 2240 4920 2260
rect 4880 2225 4920 2240
rect 4940 2310 4980 2325
rect 4940 2290 4950 2310
rect 4970 2290 4980 2310
rect 4940 2260 4980 2290
rect 4940 2240 4950 2260
rect 4970 2240 4980 2260
rect 4940 2225 4980 2240
rect 5000 2310 5040 2325
rect 5000 2290 5010 2310
rect 5030 2290 5040 2310
rect 5000 2260 5040 2290
rect 5000 2240 5010 2260
rect 5030 2240 5040 2260
rect 5000 2225 5040 2240
rect 5060 2310 5100 2325
rect 5060 2290 5070 2310
rect 5090 2290 5100 2310
rect 5060 2260 5100 2290
rect 5060 2240 5070 2260
rect 5090 2240 5100 2260
rect 5060 2225 5100 2240
rect 5120 2310 5160 2325
rect 5120 2290 5130 2310
rect 5150 2290 5160 2310
rect 5120 2260 5160 2290
rect 5120 2240 5130 2260
rect 5150 2240 5160 2260
rect 5120 2225 5160 2240
rect 5180 2310 5220 2325
rect 5180 2290 5190 2310
rect 5210 2290 5220 2310
rect 5180 2260 5220 2290
rect 5180 2240 5190 2260
rect 5210 2240 5220 2260
rect 5180 2225 5220 2240
rect 5240 2310 5280 2325
rect 5240 2290 5250 2310
rect 5270 2290 5280 2310
rect 5240 2260 5280 2290
rect 5240 2240 5250 2260
rect 5270 2240 5280 2260
rect 5240 2225 5280 2240
rect 5300 2310 5340 2325
rect 5300 2290 5310 2310
rect 5330 2290 5340 2310
rect 5300 2260 5340 2290
rect 5300 2240 5310 2260
rect 5330 2240 5340 2260
rect 5300 2225 5340 2240
rect 5360 2310 5400 2325
rect 5360 2290 5370 2310
rect 5390 2290 5400 2310
rect 5360 2260 5400 2290
rect 5360 2240 5370 2260
rect 5390 2240 5400 2260
rect 5360 2225 5400 2240
rect 5420 2310 5460 2325
rect 5420 2290 5430 2310
rect 5450 2290 5460 2310
rect 5420 2260 5460 2290
rect 5420 2240 5430 2260
rect 5450 2240 5460 2260
rect 5420 2225 5460 2240
<< ndiffc >>
rect 3140 1915 3160 1935
rect 3200 1915 3220 1935
rect 3260 1915 3280 1935
rect 3320 1915 3340 1935
rect 3380 1915 3400 1935
rect 3440 1915 3460 1935
rect 3500 1915 3520 1935
rect 3560 1915 3580 1935
rect 3620 1915 3640 1935
rect 3680 1915 3700 1935
rect 3740 1915 3760 1935
rect 4400 1915 4420 1935
rect 4460 1915 4480 1935
rect 4520 1915 4540 1935
rect 4580 1915 4600 1935
rect 4640 1915 4660 1935
rect 4700 1915 4720 1935
rect 4760 1915 4780 1935
rect 4820 1915 4840 1935
rect 4880 1915 4900 1935
rect 4940 1915 4960 1935
rect 5000 1915 5020 1935
rect 2900 1640 2920 1660
rect 2900 1590 2920 1610
rect 2900 1540 2920 1560
rect 2900 1490 2920 1510
rect 2900 1440 2920 1460
rect 3440 1640 3460 1660
rect 3440 1590 3460 1610
rect 3440 1540 3460 1560
rect 3440 1490 3460 1510
rect 3440 1440 3460 1460
rect 3980 1640 4000 1660
rect 3980 1590 4000 1610
rect 3980 1540 4000 1560
rect 3980 1490 4000 1510
rect 3980 1440 4000 1460
rect 4160 1640 4180 1660
rect 4160 1590 4180 1610
rect 4160 1540 4180 1560
rect 4160 1490 4180 1510
rect 4160 1440 4180 1460
rect 4700 1640 4720 1660
rect 4700 1590 4720 1610
rect 4700 1540 4720 1560
rect 4700 1490 4720 1510
rect 4700 1440 4720 1460
rect 5240 1640 5260 1660
rect 5240 1590 5260 1610
rect 5240 1540 5260 1560
rect 5240 1490 5260 1510
rect 5240 1440 5260 1460
rect 3030 1170 3050 1190
rect 3030 1120 3050 1140
rect 4070 1170 4090 1190
rect 4070 1120 4090 1140
rect 5110 1170 5130 1190
rect 5110 1120 5130 1140
rect 3125 895 3145 915
rect 3125 845 3145 865
rect 3180 895 3200 915
rect 3180 845 3200 865
rect 3235 895 3255 915
rect 3235 845 3255 865
rect 3290 895 3310 915
rect 3290 845 3310 865
rect 3345 895 3365 915
rect 3345 845 3365 865
rect 3400 895 3420 915
rect 3400 845 3420 865
rect 3455 895 3475 915
rect 3455 845 3475 865
rect 3510 895 3530 915
rect 3510 845 3530 865
rect 3565 895 3585 915
rect 3565 845 3585 865
rect 3620 895 3640 915
rect 3620 845 3640 865
rect 3795 895 3815 915
rect 3795 845 3815 865
rect 3850 895 3870 915
rect 3850 845 3870 865
rect 3905 895 3925 915
rect 3905 845 3925 865
rect 3960 895 3980 915
rect 3960 845 3980 865
rect 4015 895 4035 915
rect 4015 845 4035 865
rect 4070 895 4090 915
rect 4070 845 4090 865
rect 4125 895 4145 915
rect 4125 845 4145 865
rect 4180 895 4200 915
rect 4180 845 4200 865
rect 4235 895 4255 915
rect 4235 845 4255 865
rect 4290 895 4310 915
rect 4290 845 4310 865
rect 4345 895 4365 915
rect 4345 845 4365 865
rect 4520 895 4540 915
rect 4520 845 4540 865
rect 4575 895 4595 915
rect 4575 845 4595 865
rect 4630 895 4650 915
rect 4630 845 4650 865
rect 4685 895 4705 915
rect 4685 845 4705 865
rect 4740 895 4760 915
rect 4740 845 4760 865
rect 4795 895 4815 915
rect 4795 845 4815 865
rect 4850 895 4870 915
rect 4850 845 4870 865
rect 4905 895 4925 915
rect 4905 845 4925 865
rect 4960 895 4980 915
rect 4960 845 4980 865
rect 5015 895 5035 915
rect 5015 845 5035 865
<< pdiffc >>
rect 3045 3393 3065 3465
rect 3100 3393 3120 3465
rect 3155 3393 3175 3465
rect 3210 3393 3230 3465
rect 3265 3393 3285 3465
rect 3320 3393 3340 3465
rect 3375 3393 3395 3465
rect 3685 3445 3705 3465
rect 3685 3395 3705 3415
rect 3740 3445 3760 3465
rect 3740 3395 3760 3415
rect 3795 3445 3815 3465
rect 3795 3395 3815 3415
rect 3850 3445 3870 3465
rect 3850 3395 3870 3415
rect 3905 3445 3925 3465
rect 3905 3395 3925 3415
rect 3960 3445 3980 3465
rect 3960 3395 3980 3415
rect 4015 3445 4035 3465
rect 4015 3395 4035 3415
rect 4070 3445 4090 3465
rect 4070 3395 4090 3415
rect 4125 3445 4145 3465
rect 4125 3395 4145 3415
rect 4180 3445 4200 3465
rect 4180 3395 4200 3415
rect 4235 3445 4255 3465
rect 4235 3395 4255 3415
rect 4290 3445 4310 3465
rect 4290 3395 4310 3415
rect 4345 3445 4365 3465
rect 4345 3395 4365 3415
rect 4400 3445 4420 3465
rect 4400 3395 4420 3415
rect 4455 3445 4475 3465
rect 4455 3395 4475 3415
rect 4765 3395 4785 3465
rect 4820 3395 4840 3465
rect 4875 3395 4895 3465
rect 4930 3395 4950 3465
rect 4985 3395 5005 3465
rect 5040 3395 5060 3465
rect 5095 3395 5115 3465
rect 2725 2880 2745 2900
rect 2725 2830 2745 2850
rect 2780 2880 2800 2900
rect 2780 2830 2800 2850
rect 2835 2880 2855 2900
rect 2835 2830 2855 2850
rect 2890 2880 2910 2900
rect 2890 2830 2910 2850
rect 2945 2880 2965 2900
rect 2945 2830 2965 2850
rect 3260 2980 3280 3000
rect 3260 2930 3280 2950
rect 3260 2880 3280 2900
rect 3260 2830 3280 2850
rect 3260 2780 3280 2800
rect 3260 2730 3280 2750
rect 3350 2980 3370 3000
rect 3350 2930 3370 2950
rect 3350 2880 3370 2900
rect 3350 2830 3370 2850
rect 3350 2780 3370 2800
rect 3350 2730 3370 2750
rect 3440 2980 3460 3000
rect 3440 2930 3460 2950
rect 3440 2880 3460 2900
rect 3440 2830 3460 2850
rect 3440 2780 3460 2800
rect 3440 2730 3460 2750
rect 3530 2980 3550 3000
rect 3530 2930 3550 2950
rect 3530 2880 3550 2900
rect 3530 2830 3550 2850
rect 3530 2780 3550 2800
rect 3530 2730 3550 2750
rect 3620 2980 3640 3000
rect 3620 2930 3640 2950
rect 3620 2880 3640 2900
rect 3620 2830 3640 2850
rect 3620 2780 3640 2800
rect 3620 2730 3640 2750
rect 3710 2980 3730 3000
rect 3710 2930 3730 2950
rect 3710 2880 3730 2900
rect 3710 2830 3730 2850
rect 3710 2780 3730 2800
rect 3710 2730 3730 2750
rect 3800 2980 3820 3000
rect 3800 2930 3820 2950
rect 3800 2880 3820 2900
rect 3800 2830 3820 2850
rect 3800 2780 3820 2800
rect 3800 2730 3820 2750
rect 3890 2980 3910 3000
rect 3890 2930 3910 2950
rect 3890 2880 3910 2900
rect 3890 2830 3910 2850
rect 3890 2780 3910 2800
rect 3890 2730 3910 2750
rect 3980 2980 4000 3000
rect 3980 2930 4000 2950
rect 3980 2880 4000 2900
rect 3980 2830 4000 2850
rect 3980 2780 4000 2800
rect 3980 2730 4000 2750
rect 4070 2980 4090 3000
rect 4070 2930 4090 2950
rect 4070 2880 4090 2900
rect 4070 2830 4090 2850
rect 4070 2780 4090 2800
rect 4070 2730 4090 2750
rect 4160 2980 4180 3000
rect 4160 2930 4180 2950
rect 4160 2880 4180 2900
rect 4160 2830 4180 2850
rect 4160 2780 4180 2800
rect 4160 2730 4180 2750
rect 4250 2980 4270 3000
rect 4250 2930 4270 2950
rect 4250 2880 4270 2900
rect 4250 2830 4270 2850
rect 4250 2780 4270 2800
rect 4250 2730 4270 2750
rect 4340 2980 4360 3000
rect 4340 2930 4360 2950
rect 4340 2880 4360 2900
rect 4340 2830 4360 2850
rect 4340 2780 4360 2800
rect 4340 2730 4360 2750
rect 4430 2980 4450 3000
rect 4430 2930 4450 2950
rect 4430 2880 4450 2900
rect 4430 2830 4450 2850
rect 4430 2780 4450 2800
rect 4430 2730 4450 2750
rect 4520 2980 4540 3000
rect 4520 2930 4540 2950
rect 4520 2880 4540 2900
rect 4520 2830 4540 2850
rect 4520 2780 4540 2800
rect 4520 2730 4540 2750
rect 4610 2980 4630 3000
rect 4610 2930 4630 2950
rect 4610 2880 4630 2900
rect 4610 2830 4630 2850
rect 4610 2780 4630 2800
rect 4610 2730 4630 2750
rect 4700 2980 4720 3000
rect 4700 2930 4720 2950
rect 4700 2880 4720 2900
rect 4700 2830 4720 2850
rect 4700 2780 4720 2800
rect 4700 2730 4720 2750
rect 4790 2980 4810 3000
rect 4790 2930 4810 2950
rect 4790 2880 4810 2900
rect 4790 2830 4810 2850
rect 4790 2780 4810 2800
rect 4790 2730 4810 2750
rect 4880 2980 4900 3000
rect 4880 2930 4900 2950
rect 4880 2880 4900 2900
rect 4880 2830 4900 2850
rect 4880 2780 4900 2800
rect 4880 2730 4900 2750
rect 5190 2880 5210 2900
rect 5190 2830 5210 2850
rect 5245 2880 5265 2900
rect 5245 2830 5265 2850
rect 5300 2880 5320 2900
rect 5300 2830 5320 2850
rect 5355 2880 5375 2900
rect 5355 2830 5375 2850
rect 5410 2880 5430 2900
rect 5410 2830 5430 2850
rect 2710 2290 2730 2310
rect 2710 2240 2730 2260
rect 2770 2290 2790 2310
rect 2770 2240 2790 2260
rect 2830 2290 2850 2310
rect 2830 2240 2850 2260
rect 2890 2290 2910 2310
rect 2890 2240 2910 2260
rect 2950 2290 2970 2310
rect 2950 2240 2970 2260
rect 3010 2290 3030 2310
rect 3010 2240 3030 2260
rect 3070 2290 3090 2310
rect 3070 2240 3090 2260
rect 3130 2290 3150 2310
rect 3130 2240 3150 2260
rect 3190 2290 3210 2310
rect 3190 2240 3210 2260
rect 3250 2290 3270 2310
rect 3250 2240 3270 2260
rect 3310 2290 3330 2310
rect 3310 2240 3330 2260
rect 3370 2290 3390 2310
rect 3370 2240 3390 2260
rect 3430 2290 3450 2310
rect 3430 2240 3450 2260
rect 3490 2290 3510 2310
rect 3490 2240 3510 2260
rect 3550 2290 3570 2310
rect 3550 2240 3570 2260
rect 3610 2290 3630 2310
rect 3610 2240 3630 2260
rect 3670 2290 3690 2310
rect 3670 2240 3690 2260
rect 3730 2290 3750 2310
rect 3730 2240 3750 2260
rect 3790 2290 3810 2310
rect 3790 2240 3810 2260
rect 3850 2290 3870 2310
rect 3850 2240 3870 2260
rect 3910 2290 3930 2310
rect 3910 2240 3930 2260
rect 4230 2290 4250 2310
rect 4230 2240 4250 2260
rect 4290 2290 4310 2310
rect 4290 2240 4310 2260
rect 4350 2290 4370 2310
rect 4350 2240 4370 2260
rect 4410 2290 4430 2310
rect 4410 2240 4430 2260
rect 4470 2290 4490 2310
rect 4470 2240 4490 2260
rect 4530 2290 4550 2310
rect 4530 2240 4550 2260
rect 4590 2290 4610 2310
rect 4590 2240 4610 2260
rect 4650 2290 4670 2310
rect 4650 2240 4670 2260
rect 4710 2290 4730 2310
rect 4710 2240 4730 2260
rect 4770 2290 4790 2310
rect 4770 2240 4790 2260
rect 4830 2290 4850 2310
rect 4830 2240 4850 2260
rect 4890 2290 4910 2310
rect 4890 2240 4910 2260
rect 4950 2290 4970 2310
rect 4950 2240 4970 2260
rect 5010 2290 5030 2310
rect 5010 2240 5030 2260
rect 5070 2290 5090 2310
rect 5070 2240 5090 2260
rect 5130 2290 5150 2310
rect 5130 2240 5150 2260
rect 5190 2290 5210 2310
rect 5190 2240 5210 2260
rect 5250 2290 5270 2310
rect 5250 2240 5270 2260
rect 5310 2290 5330 2310
rect 5310 2240 5330 2260
rect 5370 2290 5390 2310
rect 5370 2240 5390 2260
rect 5430 2290 5450 2310
rect 5430 2240 5450 2260
<< psubdiff >>
rect 25 3640 590 3660
rect 670 3640 1235 3660
rect 25 3580 45 3640
rect 1215 3580 1235 3640
rect 25 3445 45 3500
rect 1215 3445 1235 3500
rect 25 3425 590 3445
rect 670 3425 1235 3445
rect 1310 3505 1845 3525
rect 1925 3505 2505 3525
rect 25 3375 575 3395
rect 655 3375 1205 3395
rect 25 3315 45 3375
rect 1185 3315 1205 3375
rect 25 3180 45 3235
rect 1185 3180 1205 3235
rect 25 3160 575 3180
rect 655 3160 1205 3180
rect 1310 3325 1330 3505
rect 2485 3325 2505 3505
rect 220 3110 575 3130
rect 655 3110 1020 3130
rect 220 3080 240 3110
rect 1000 3080 1020 3110
rect 220 2970 240 3000
rect 1310 3070 1330 3245
rect 2485 3070 2505 3245
rect 1310 3050 1845 3070
rect 1925 3050 2505 3070
rect 1000 2970 1020 3000
rect 220 2950 575 2970
rect 655 2950 1020 2970
rect 1475 3000 1845 3020
rect 1925 3000 2300 3020
rect 1475 2970 1495 3000
rect 220 2900 575 2920
rect 655 2900 1020 2920
rect 220 2870 240 2900
rect 1000 2870 1020 2900
rect 220 2760 240 2790
rect 2280 2970 2300 3000
rect 1475 2865 1495 2890
rect 2280 2865 2300 2890
rect 1475 2845 1845 2865
rect 1925 2845 2300 2865
rect 1000 2760 1020 2790
rect 220 2740 575 2760
rect 655 2740 1020 2760
rect 3080 2070 3410 2090
rect 3490 2070 3820 2090
rect 3080 1965 3100 2070
rect 3800 1965 3820 2070
rect 3080 1825 3100 1885
rect 3800 1825 3820 1885
rect 3080 1805 3410 1825
rect 3490 1805 3820 1825
rect 4340 2070 4670 2090
rect 4750 2070 5080 2090
rect 4340 1965 4360 2070
rect 5060 1965 5080 2070
rect 4340 1825 4360 1885
rect 5060 1825 5080 1885
rect 4340 1805 5080 1825
rect 2840 1745 3410 1765
rect 3490 1745 4060 1765
rect -50 1715 100 1730
rect -50 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 100 1715
rect -50 1680 100 1695
rect 2840 1590 2860 1745
rect 2840 1350 2860 1510
rect 4040 1590 4060 1745
rect 4040 1350 4060 1510
rect 2840 1330 3410 1350
rect 3490 1330 4060 1350
rect 4100 1745 4670 1765
rect 4750 1745 5320 1765
rect 4100 1590 4120 1745
rect 4100 1350 4120 1510
rect 5300 1590 5320 1745
rect 5300 1350 5320 1510
rect 4100 1330 4670 1350
rect 4750 1330 5320 1350
rect 2940 1280 4040 1300
rect 4120 1280 5215 1300
rect 2940 1195 2960 1280
rect 2940 1075 2960 1115
rect 5195 1195 5215 1280
rect 5195 1075 5215 1115
rect 2940 1055 4040 1075
rect 4120 1055 5215 1075
rect 3065 1005 3345 1025
rect 3425 1005 3700 1025
rect 3065 920 3085 1005
rect 3065 755 3085 840
rect 3680 920 3700 1005
rect 3680 755 3700 840
rect 3065 735 3345 755
rect 3425 735 3700 755
rect 3735 1005 4040 1025
rect 4120 1005 4425 1025
rect 3735 920 3755 1005
rect 3735 755 3755 840
rect 4405 920 4425 1005
rect 4405 755 4425 840
rect 3735 735 4040 755
rect 4120 735 4425 755
rect 4460 1005 4735 1025
rect 4815 1005 5095 1025
rect 4460 920 4480 1005
rect 4460 755 4480 840
rect 5075 920 5095 1005
rect 5075 755 5095 840
rect 4460 735 4735 755
rect 4815 735 5095 755
<< nsubdiff >>
rect 2985 3555 3180 3575
rect 3260 3555 3455 3575
rect 2985 3470 3005 3555
rect 2985 3305 3005 3390
rect 3435 3470 3455 3555
rect 3435 3305 3455 3390
rect 2985 3285 3180 3305
rect 3260 3285 3455 3305
rect 3625 3555 4040 3575
rect 4120 3555 4535 3575
rect 3625 3470 3645 3555
rect 3625 3305 3645 3390
rect 4515 3470 4535 3555
rect 4515 3305 4535 3390
rect 3625 3285 4040 3305
rect 4120 3285 4535 3305
rect 4705 3555 4900 3575
rect 4980 3555 5175 3575
rect 4705 3470 4725 3555
rect 4705 3305 4725 3390
rect 5155 3470 5175 3555
rect 5155 3305 5175 3390
rect 4705 3285 4900 3305
rect 4965 3285 5175 3305
rect 3200 3090 4040 3110
rect 4120 3090 4960 3110
rect 2665 2990 2805 3010
rect 2885 2990 3025 3010
rect 2665 2905 2685 2990
rect 2665 2740 2685 2825
rect 3005 2905 3025 2990
rect 3005 2740 3025 2825
rect 2665 2720 2805 2740
rect 2885 2720 3025 2740
rect 3200 2905 3220 3090
rect 3200 2635 3220 2825
rect 4940 2905 4960 3090
rect 4940 2635 4960 2825
rect 5130 2990 5270 3010
rect 5350 2990 5490 3010
rect 5130 2905 5150 2990
rect 5130 2740 5150 2825
rect 5470 2905 5490 2990
rect 5470 2740 5490 2825
rect 5130 2720 5270 2740
rect 5350 2720 5490 2740
rect 3200 2615 4040 2635
rect 4120 2615 4960 2635
rect 2650 2400 3280 2420
rect 3360 2400 3990 2420
rect 2650 2315 2670 2400
rect 2650 2150 2670 2235
rect 3970 2315 3990 2400
rect 3970 2150 3990 2235
rect 2650 2130 3280 2150
rect 3360 2130 3990 2150
rect 4170 2400 4800 2420
rect 4880 2400 5510 2420
rect 4170 2315 4190 2400
rect 4170 2150 4190 2235
rect 5490 2315 5510 2400
rect 5490 2150 5510 2235
rect 4170 2130 4800 2150
rect 4880 2130 5510 2150
<< psubdiffcont >>
rect 590 3640 670 3660
rect 25 3500 45 3580
rect 1215 3500 1235 3580
rect 590 3425 670 3445
rect 1845 3505 1925 3525
rect 575 3375 655 3395
rect 25 3235 45 3315
rect 1185 3235 1205 3315
rect 575 3160 655 3180
rect 1310 3245 1330 3325
rect 575 3110 655 3130
rect 220 3000 240 3080
rect 1000 3000 1020 3080
rect 2485 3245 2505 3325
rect 1845 3050 1925 3070
rect 575 2950 655 2970
rect 1845 3000 1925 3020
rect 575 2900 655 2920
rect 220 2790 240 2870
rect 1000 2790 1020 2870
rect 1475 2890 1495 2970
rect 2280 2890 2300 2970
rect 1845 2845 1925 2865
rect 575 2740 655 2760
rect 3410 2070 3490 2090
rect 3080 1885 3100 1965
rect 3800 1885 3820 1965
rect 3410 1805 3490 1825
rect 4670 2070 4750 2090
rect 4340 1885 4360 1965
rect 5060 1885 5080 1965
rect 3410 1745 3490 1765
rect -35 1695 -15 1715
rect 15 1695 35 1715
rect 65 1695 85 1715
rect 2840 1510 2860 1590
rect 4040 1510 4060 1590
rect 3410 1330 3490 1350
rect 4670 1745 4750 1765
rect 4100 1510 4120 1590
rect 5300 1510 5320 1590
rect 4670 1330 4750 1350
rect 4040 1280 4120 1300
rect 2940 1115 2960 1195
rect 5195 1115 5215 1195
rect 4040 1055 4120 1075
rect 3345 1005 3425 1025
rect 3065 840 3085 920
rect 3680 840 3700 920
rect 3345 735 3425 755
rect 4040 1005 4120 1025
rect 3735 840 3755 920
rect 4405 840 4425 920
rect 4040 735 4120 755
rect 4735 1005 4815 1025
rect 4460 840 4480 920
rect 5075 840 5095 920
rect 4735 735 4815 755
<< nsubdiffcont >>
rect 3180 3555 3260 3575
rect 2985 3390 3005 3470
rect 3435 3390 3455 3470
rect 3180 3285 3260 3305
rect 4040 3555 4120 3575
rect 3625 3390 3645 3470
rect 4515 3390 4535 3470
rect 4040 3285 4120 3305
rect 4900 3555 4980 3575
rect 4705 3390 4725 3470
rect 5155 3390 5175 3470
rect 4900 3285 4965 3305
rect 4040 3090 4120 3110
rect 2805 2990 2885 3010
rect 2665 2825 2685 2905
rect 3005 2825 3025 2905
rect 2805 2720 2885 2740
rect 3200 2825 3220 2905
rect 4940 2825 4960 2905
rect 5270 2990 5350 3010
rect 5130 2825 5150 2905
rect 5470 2825 5490 2905
rect 5270 2720 5350 2740
rect 4040 2615 4120 2635
rect 3280 2400 3360 2420
rect 2650 2235 2670 2315
rect 3970 2235 3990 2315
rect 3280 2130 3360 2150
rect 4800 2400 4880 2420
rect 4170 2235 4190 2315
rect 5490 2235 5510 2315
rect 4800 2130 4880 2150
<< poly >>
rect 3035 3525 3075 3535
rect 3035 3505 3045 3525
rect 3065 3510 3075 3525
rect 3205 3525 3235 3535
rect 3065 3505 3090 3510
rect 3205 3505 3210 3525
rect 3230 3505 3235 3525
rect 3365 3525 3405 3535
rect 3365 3505 3375 3525
rect 3395 3505 3405 3525
rect 3035 3495 3090 3505
rect 3075 3480 3090 3495
rect 3130 3490 3310 3505
rect 3130 3480 3145 3490
rect 3185 3480 3200 3490
rect 3240 3480 3255 3490
rect 3295 3480 3310 3490
rect 3350 3490 3405 3505
rect 3350 3480 3365 3490
rect 3075 3365 3090 3380
rect 3130 3365 3145 3380
rect 3185 3365 3200 3380
rect 3240 3365 3255 3380
rect 3295 3365 3310 3380
rect 3350 3365 3365 3380
rect 3675 3525 3715 3535
rect 3675 3505 3685 3525
rect 3705 3510 3715 3525
rect 4065 3525 4095 3535
rect 3705 3505 3730 3510
rect 4065 3505 4070 3525
rect 4090 3505 4095 3525
rect 4445 3525 4485 3535
rect 4445 3510 4455 3525
rect 4265 3505 4390 3510
rect 3675 3495 3730 3505
rect 3715 3480 3730 3495
rect 3770 3490 4390 3505
rect 3770 3480 3785 3490
rect 3825 3480 3840 3490
rect 3880 3480 3895 3490
rect 3935 3480 3950 3490
rect 3990 3480 4005 3490
rect 4045 3480 4060 3490
rect 4100 3480 4115 3490
rect 4155 3480 4170 3490
rect 4210 3480 4225 3490
rect 4265 3480 4280 3490
rect 4320 3480 4335 3490
rect 4375 3480 4390 3490
rect 4430 3505 4455 3510
rect 4475 3505 4485 3525
rect 4430 3495 4485 3505
rect 4430 3480 4445 3495
rect 3715 3365 3730 3380
rect 3770 3365 3785 3380
rect 3825 3365 3840 3380
rect 3880 3365 3895 3380
rect 3935 3365 3950 3380
rect 3990 3365 4005 3380
rect 4045 3365 4060 3380
rect 4100 3365 4115 3380
rect 4155 3365 4170 3380
rect 4210 3365 4225 3380
rect 4265 3365 4280 3380
rect 4320 3365 4335 3380
rect 4375 3365 4390 3380
rect 4430 3365 4445 3380
rect 4755 3525 4795 3535
rect 4755 3505 4765 3525
rect 4785 3510 4795 3525
rect 4925 3525 4955 3535
rect 4785 3505 4810 3510
rect 4925 3505 4930 3525
rect 4950 3505 4955 3525
rect 5085 3525 5125 3535
rect 5085 3510 5095 3525
rect 5070 3505 5095 3510
rect 5115 3505 5125 3525
rect 4755 3495 4810 3505
rect 4795 3480 4810 3495
rect 4850 3490 5030 3505
rect 4850 3480 4865 3490
rect 4905 3480 4920 3490
rect 4960 3480 4975 3490
rect 5015 3480 5030 3490
rect 5070 3495 5125 3505
rect 5070 3480 5085 3495
rect 4795 3365 4810 3380
rect 4850 3365 4865 3380
rect 4905 3365 4920 3380
rect 4960 3365 4975 3380
rect 5015 3365 5030 3380
rect 5070 3365 5085 3380
rect 2720 2960 2750 2970
rect 2720 2940 2725 2960
rect 2745 2940 2750 2960
rect 2940 2960 2970 2970
rect 2940 2940 2945 2960
rect 2965 2940 2970 2960
rect 2720 2925 2770 2940
rect 2755 2915 2770 2925
rect 2810 2915 2825 2930
rect 2865 2915 2880 2930
rect 2920 2925 2970 2940
rect 2920 2915 2935 2925
rect 2755 2800 2770 2815
rect 2810 2805 2825 2815
rect 2865 2805 2880 2815
rect 2810 2790 2880 2805
rect 2920 2800 2935 2815
rect 2825 2770 2835 2790
rect 2855 2770 2865 2790
rect 2825 2760 2865 2770
rect 3250 3060 3290 3070
rect 3250 3040 3260 3060
rect 3280 3045 3290 3060
rect 4870 3060 4910 3070
rect 4870 3045 4880 3060
rect 3280 3040 3340 3045
rect 3250 3030 3340 3040
rect 4820 3040 4880 3045
rect 4900 3040 4910 3060
rect 4820 3030 4910 3040
rect 3290 3015 3340 3030
rect 3380 3015 3430 3030
rect 3470 3015 3520 3030
rect 3560 3015 3610 3030
rect 3650 3015 3700 3030
rect 3740 3015 3790 3030
rect 3830 3015 3880 3030
rect 3920 3015 3970 3030
rect 4010 3015 4060 3030
rect 4100 3015 4150 3030
rect 4190 3015 4240 3030
rect 4280 3015 4330 3030
rect 4370 3015 4420 3030
rect 4460 3015 4510 3030
rect 4550 3015 4600 3030
rect 4640 3015 4690 3030
rect 4730 3015 4780 3030
rect 4820 3015 4870 3030
rect 3290 2700 3340 2715
rect 3380 2705 3430 2715
rect 3470 2705 3520 2715
rect 3560 2705 3610 2715
rect 3650 2705 3700 2715
rect 3740 2705 3790 2715
rect 3830 2705 3880 2715
rect 3920 2705 3970 2715
rect 4010 2705 4060 2715
rect 4100 2705 4150 2715
rect 4190 2705 4240 2715
rect 4280 2705 4330 2715
rect 4370 2705 4420 2715
rect 4460 2705 4510 2715
rect 4550 2705 4600 2715
rect 4640 2705 4690 2715
rect 4730 2705 4780 2715
rect 3380 2690 4780 2705
rect 4820 2700 4870 2715
rect 3970 2670 3980 2690
rect 4000 2670 4010 2690
rect 3970 2660 4010 2670
rect 4690 2670 4700 2690
rect 4720 2670 4730 2690
rect 4690 2660 4730 2670
rect 5185 2960 5215 2970
rect 5185 2940 5190 2960
rect 5210 2945 5215 2960
rect 5405 2960 5435 2970
rect 5405 2945 5410 2960
rect 5210 2940 5235 2945
rect 5185 2930 5235 2940
rect 5385 2940 5410 2945
rect 5430 2940 5435 2960
rect 5385 2930 5435 2940
rect 5220 2915 5235 2930
rect 5275 2915 5290 2930
rect 5330 2915 5345 2930
rect 5385 2915 5400 2930
rect 5220 2800 5235 2815
rect 5275 2805 5290 2815
rect 5330 2805 5345 2815
rect 5275 2790 5345 2805
rect 5385 2800 5400 2815
rect 5290 2770 5300 2790
rect 5320 2770 5330 2790
rect 5290 2760 5330 2770
rect 2740 2325 2760 2340
rect 2800 2325 2820 2340
rect 2860 2325 2880 2340
rect 2920 2325 2940 2340
rect 2980 2325 3000 2340
rect 3040 2325 3060 2340
rect 3100 2325 3120 2340
rect 3160 2325 3180 2340
rect 3220 2325 3240 2340
rect 3280 2325 3300 2340
rect 3340 2325 3360 2340
rect 3400 2325 3420 2340
rect 3460 2325 3480 2340
rect 3520 2325 3540 2340
rect 3580 2325 3600 2340
rect 3640 2325 3660 2340
rect 3700 2325 3720 2340
rect 3760 2325 3780 2340
rect 3820 2325 3840 2340
rect 3880 2325 3900 2340
rect 2740 2215 2760 2225
rect 2705 2200 2760 2215
rect 2800 2210 2820 2225
rect 2860 2215 2880 2225
rect 2920 2215 2940 2225
rect 2980 2215 3000 2225
rect 3040 2215 3060 2225
rect 2790 2200 2830 2210
rect 2860 2200 3060 2215
rect 3100 2215 3120 2225
rect 3160 2215 3180 2225
rect 3100 2200 3180 2215
rect 3220 2215 3240 2225
rect 3280 2215 3300 2225
rect 3340 2215 3360 2225
rect 3400 2215 3420 2225
rect 3220 2200 3420 2215
rect 3460 2215 3480 2225
rect 3520 2215 3540 2225
rect 3460 2200 3540 2215
rect 3580 2215 3600 2225
rect 3640 2215 3660 2225
rect 3700 2215 3720 2225
rect 3760 2215 3780 2225
rect 3580 2200 3780 2215
rect 3820 2210 3840 2225
rect 3880 2215 3900 2225
rect 3815 2200 3845 2210
rect 3880 2200 3935 2215
rect 2705 2180 2710 2200
rect 2730 2180 2735 2200
rect 2705 2170 2735 2180
rect 2790 2180 2800 2200
rect 2820 2180 2830 2200
rect 2790 2170 2830 2180
rect 2880 2180 2890 2200
rect 2910 2180 2920 2200
rect 2880 2170 2920 2180
rect 3120 2180 3130 2200
rect 3150 2180 3160 2200
rect 3120 2170 3160 2180
rect 3240 2180 3250 2200
rect 3270 2180 3280 2200
rect 3240 2170 3280 2180
rect 3480 2180 3490 2200
rect 3510 2180 3520 2200
rect 3480 2170 3520 2180
rect 3600 2180 3610 2200
rect 3630 2180 3640 2200
rect 3600 2170 3640 2180
rect 3815 2180 3820 2200
rect 3840 2180 3845 2200
rect 3815 2170 3845 2180
rect 3905 2180 3910 2200
rect 3930 2180 3935 2200
rect 3905 2170 3935 2180
rect 4260 2325 4280 2340
rect 4320 2325 4340 2340
rect 4380 2325 4400 2340
rect 4440 2325 4460 2340
rect 4500 2325 4520 2340
rect 4560 2325 4580 2340
rect 4620 2325 4640 2340
rect 4680 2325 4700 2340
rect 4740 2325 4760 2340
rect 4800 2325 4820 2340
rect 4860 2325 4880 2340
rect 4920 2325 4940 2340
rect 4980 2325 5000 2340
rect 5040 2325 5060 2340
rect 5100 2325 5120 2340
rect 5160 2325 5180 2340
rect 5220 2325 5240 2340
rect 5280 2325 5300 2340
rect 5340 2325 5360 2340
rect 5400 2325 5420 2340
rect 4260 2215 4280 2225
rect 4225 2200 4280 2215
rect 4320 2210 4340 2225
rect 4380 2215 4400 2225
rect 4440 2215 4460 2225
rect 4500 2215 4520 2225
rect 4560 2215 4580 2225
rect 4315 2200 4345 2210
rect 4380 2200 4580 2215
rect 4620 2215 4640 2225
rect 4680 2215 4700 2225
rect 4620 2200 4700 2215
rect 4740 2215 4760 2225
rect 4800 2215 4820 2225
rect 4860 2215 4880 2225
rect 4920 2215 4940 2225
rect 4740 2200 4940 2215
rect 4980 2215 5000 2225
rect 5040 2215 5060 2225
rect 4980 2200 5060 2215
rect 5100 2215 5120 2225
rect 5160 2215 5180 2225
rect 5220 2215 5240 2225
rect 5280 2215 5300 2225
rect 5100 2200 5300 2215
rect 5340 2210 5360 2225
rect 5400 2215 5420 2225
rect 5330 2200 5370 2210
rect 5400 2200 5455 2215
rect 4225 2180 4230 2200
rect 4250 2180 4255 2200
rect 4225 2170 4255 2180
rect 4315 2180 4320 2200
rect 4340 2180 4345 2200
rect 4315 2170 4345 2180
rect 4520 2180 4530 2200
rect 4550 2180 4560 2200
rect 4520 2170 4560 2180
rect 4640 2180 4650 2200
rect 4670 2180 4680 2200
rect 4640 2170 4680 2180
rect 4880 2180 4890 2200
rect 4910 2180 4920 2200
rect 4880 2170 4920 2180
rect 5000 2180 5010 2200
rect 5030 2180 5040 2200
rect 5000 2170 5040 2180
rect 5240 2180 5250 2200
rect 5270 2180 5280 2200
rect 5240 2170 5280 2180
rect 5330 2180 5340 2200
rect 5360 2180 5370 2200
rect 5330 2170 5370 2180
rect 5425 2180 5430 2200
rect 5450 2180 5455 2200
rect 5425 2170 5455 2180
rect 3190 2040 3230 2050
rect 3190 2020 3200 2040
rect 3220 2020 3230 2040
rect 3190 2005 3230 2020
rect 3190 1990 3730 2005
rect 3170 1950 3190 1965
rect 3230 1950 3250 1990
rect 3290 1950 3310 1990
rect 3350 1950 3370 1965
rect 3410 1950 3430 1965
rect 3470 1950 3490 1990
rect 3530 1950 3550 1990
rect 3590 1950 3610 1965
rect 3650 1950 3670 1965
rect 3710 1950 3730 1990
rect 3170 1885 3190 1900
rect 3230 1885 3250 1900
rect 3290 1885 3310 1900
rect 3130 1875 3190 1885
rect 3130 1855 3140 1875
rect 3160 1860 3190 1875
rect 3350 1860 3370 1900
rect 3410 1860 3430 1900
rect 3470 1885 3490 1900
rect 3530 1885 3550 1900
rect 3590 1860 3610 1900
rect 3650 1860 3670 1900
rect 3710 1885 3730 1900
rect 3160 1855 3670 1860
rect 3130 1845 3670 1855
rect 4930 2040 4970 2050
rect 4930 2020 4940 2040
rect 4960 2020 4970 2040
rect 4930 2005 4970 2020
rect 4430 1990 4970 2005
rect 4430 1950 4450 1990
rect 4490 1950 4510 1965
rect 4550 1950 4570 1965
rect 4610 1950 4630 1990
rect 4670 1950 4690 1990
rect 4730 1950 4750 1965
rect 4790 1950 4810 1965
rect 4850 1950 4870 1990
rect 4910 1950 4930 1990
rect 4970 1950 4990 1965
rect 4430 1885 4450 1900
rect 4490 1860 4510 1900
rect 4550 1860 4570 1900
rect 4610 1885 4630 1900
rect 4670 1885 4690 1900
rect 4730 1860 4750 1900
rect 4790 1860 4810 1900
rect 4850 1885 4870 1900
rect 4910 1885 4930 1900
rect 4970 1885 4990 1900
rect 4970 1875 5030 1885
rect 4970 1860 5000 1875
rect 4490 1855 5000 1860
rect 5020 1855 5030 1875
rect 4490 1845 5030 1855
rect 2980 1715 3020 1725
rect 2980 1695 2990 1715
rect 3010 1695 3020 1715
rect 2980 1690 3020 1695
rect 3100 1715 3140 1725
rect 3100 1695 3110 1715
rect 3130 1695 3140 1715
rect 3100 1690 3140 1695
rect 3220 1715 3260 1725
rect 3220 1695 3230 1715
rect 3250 1695 3260 1715
rect 3220 1690 3260 1695
rect 3340 1715 3380 1725
rect 3340 1695 3350 1715
rect 3370 1695 3380 1715
rect 3340 1690 3380 1695
rect 3580 1715 3620 1725
rect 3580 1695 3590 1715
rect 3610 1695 3620 1715
rect 3580 1690 3620 1695
rect 3700 1715 3740 1725
rect 3700 1695 3710 1715
rect 3730 1695 3740 1715
rect 3700 1690 3740 1695
rect 3820 1715 3860 1725
rect 3820 1695 3830 1715
rect 3850 1695 3860 1715
rect 3820 1690 3860 1695
rect 2930 1675 3430 1690
rect 3470 1675 3970 1690
rect 2930 1410 3430 1425
rect 3470 1410 3970 1425
rect 4300 1715 4340 1725
rect 4300 1695 4310 1715
rect 4330 1695 4340 1715
rect 4300 1690 4340 1695
rect 4420 1715 4460 1725
rect 4420 1695 4430 1715
rect 4450 1695 4460 1715
rect 4420 1690 4460 1695
rect 4540 1715 4580 1725
rect 4540 1695 4550 1715
rect 4570 1695 4580 1715
rect 4540 1690 4580 1695
rect 4780 1715 4820 1725
rect 4780 1695 4790 1715
rect 4810 1695 4820 1715
rect 4780 1690 4820 1695
rect 4900 1715 4940 1725
rect 4900 1695 4910 1715
rect 4930 1695 4940 1715
rect 4900 1690 4940 1695
rect 5020 1715 5060 1725
rect 5020 1695 5030 1715
rect 5050 1695 5060 1715
rect 5020 1690 5060 1695
rect 5140 1715 5180 1725
rect 5140 1695 5150 1715
rect 5170 1695 5180 1715
rect 5140 1690 5180 1695
rect 4190 1675 4690 1690
rect 4730 1675 5230 1690
rect 4190 1410 4690 1425
rect 4730 1410 5230 1425
rect 3100 1250 3140 1260
rect 3100 1230 3110 1250
rect 3130 1230 3140 1250
rect 3100 1220 3140 1230
rect 3180 1250 3220 1260
rect 3180 1230 3190 1250
rect 3210 1230 3220 1250
rect 3180 1220 3220 1230
rect 3260 1250 3300 1260
rect 3260 1230 3270 1250
rect 3290 1230 3300 1250
rect 3260 1220 3300 1230
rect 3340 1250 3380 1260
rect 3340 1230 3350 1250
rect 3370 1230 3380 1250
rect 3340 1220 3380 1230
rect 3420 1250 3460 1260
rect 3420 1230 3430 1250
rect 3450 1230 3460 1250
rect 3420 1220 3460 1230
rect 3500 1250 3540 1260
rect 3500 1230 3510 1250
rect 3530 1230 3540 1250
rect 3500 1220 3540 1230
rect 3580 1250 3620 1260
rect 3580 1230 3590 1250
rect 3610 1230 3620 1250
rect 3580 1220 3620 1230
rect 3660 1250 3700 1260
rect 3660 1230 3670 1250
rect 3690 1230 3700 1250
rect 3660 1220 3700 1230
rect 3740 1250 3780 1260
rect 3740 1230 3750 1250
rect 3770 1230 3780 1250
rect 3740 1220 3780 1230
rect 3820 1250 3860 1260
rect 3820 1230 3830 1250
rect 3850 1230 3860 1250
rect 3820 1220 3860 1230
rect 3900 1250 3940 1260
rect 3900 1230 3910 1250
rect 3930 1230 3940 1250
rect 3900 1220 3940 1230
rect 3980 1250 4020 1260
rect 3980 1230 3990 1250
rect 4010 1230 4020 1250
rect 3980 1220 4020 1230
rect 4140 1250 4180 1260
rect 4140 1230 4150 1250
rect 4170 1230 4180 1250
rect 4140 1220 4180 1230
rect 4220 1250 4260 1260
rect 4220 1230 4230 1250
rect 4250 1230 4260 1250
rect 4220 1220 4260 1230
rect 4300 1250 4340 1260
rect 4300 1230 4310 1250
rect 4330 1230 4340 1250
rect 4300 1220 4340 1230
rect 4380 1250 4420 1260
rect 4380 1230 4390 1250
rect 4410 1230 4420 1250
rect 4380 1220 4420 1230
rect 4460 1250 4500 1260
rect 4460 1230 4470 1250
rect 4490 1230 4500 1250
rect 4460 1220 4500 1230
rect 4540 1250 4580 1260
rect 4540 1230 4550 1250
rect 4570 1230 4580 1250
rect 4540 1220 4580 1230
rect 4620 1250 4660 1260
rect 4620 1230 4630 1250
rect 4650 1230 4660 1250
rect 4620 1220 4660 1230
rect 4700 1250 4740 1260
rect 4700 1230 4710 1250
rect 4730 1230 4740 1250
rect 4700 1220 4740 1230
rect 4780 1250 4820 1260
rect 4780 1230 4790 1250
rect 4810 1230 4820 1250
rect 4780 1220 4820 1230
rect 4860 1250 4900 1260
rect 4860 1230 4870 1250
rect 4890 1230 4900 1250
rect 4860 1220 4900 1230
rect 4940 1250 4980 1260
rect 4940 1230 4950 1250
rect 4970 1230 4980 1250
rect 4940 1220 4980 1230
rect 5020 1250 5060 1260
rect 5020 1230 5030 1250
rect 5050 1230 5060 1250
rect 5020 1220 5060 1230
rect 3060 1205 4060 1220
rect 4100 1205 5100 1220
rect 3060 1090 4060 1105
rect 4100 1090 5100 1105
rect 3395 975 3425 985
rect 3395 955 3400 975
rect 3420 955 3425 975
rect 3155 930 3170 945
rect 3210 940 3555 955
rect 3210 930 3225 940
rect 3265 930 3280 940
rect 3320 930 3335 940
rect 3375 930 3390 940
rect 3430 930 3445 940
rect 3485 930 3500 940
rect 3540 930 3555 940
rect 3595 930 3610 945
rect 3155 820 3170 830
rect 3120 805 3170 820
rect 3210 815 3225 830
rect 3265 815 3280 830
rect 3320 815 3335 830
rect 3375 815 3390 830
rect 3430 815 3445 830
rect 3485 815 3500 830
rect 3540 815 3555 830
rect 3595 820 3610 830
rect 3595 805 3645 820
rect 3120 785 3125 805
rect 3145 785 3150 805
rect 3120 775 3150 785
rect 3615 785 3620 805
rect 3640 785 3645 805
rect 3615 775 3645 785
rect 4065 975 4095 985
rect 4065 955 4070 975
rect 4090 955 4095 975
rect 3825 930 3840 945
rect 3880 940 4280 955
rect 3880 930 3895 940
rect 3935 930 3950 940
rect 3990 930 4005 940
rect 4045 930 4060 940
rect 4100 930 4115 940
rect 4155 930 4170 940
rect 4210 930 4225 940
rect 4265 930 4280 940
rect 4320 930 4335 945
rect 3825 820 3840 830
rect 3790 805 3840 820
rect 3880 815 3895 830
rect 3935 815 3950 830
rect 3990 815 4005 830
rect 4045 815 4060 830
rect 4100 815 4115 830
rect 4155 815 4170 830
rect 4210 815 4225 830
rect 4265 815 4280 830
rect 4320 820 4335 830
rect 3865 805 3905 815
rect 4320 805 4370 820
rect 3790 785 3795 805
rect 3815 785 3820 805
rect 3790 775 3820 785
rect 3865 785 3875 805
rect 3895 785 3905 805
rect 3865 775 3905 785
rect 4340 785 4345 805
rect 4365 785 4370 805
rect 4340 775 4370 785
rect 4735 975 4765 985
rect 4735 955 4740 975
rect 4760 955 4765 975
rect 4550 930 4565 945
rect 4605 940 4950 955
rect 4605 930 4620 940
rect 4660 930 4675 940
rect 4715 930 4730 940
rect 4770 930 4785 940
rect 4825 930 4840 940
rect 4880 930 4895 940
rect 4935 930 4950 940
rect 4990 930 5005 945
rect 4550 820 4565 830
rect 4515 805 4565 820
rect 4605 815 4620 830
rect 4660 815 4675 830
rect 4715 815 4730 830
rect 4770 815 4785 830
rect 4825 815 4840 830
rect 4880 815 4895 830
rect 4935 815 4950 830
rect 4990 820 5005 830
rect 4990 805 5040 820
rect 4515 785 4520 805
rect 4540 785 4545 805
rect 4515 775 4545 785
rect 5010 785 5015 805
rect 5035 785 5040 805
rect 5010 775 5040 785
<< polycont >>
rect 3045 3505 3065 3525
rect 3210 3505 3230 3525
rect 3375 3505 3395 3525
rect 3685 3505 3705 3525
rect 4070 3505 4090 3525
rect 4455 3505 4475 3525
rect 4765 3505 4785 3525
rect 4930 3505 4950 3525
rect 5095 3505 5115 3525
rect 2725 2940 2745 2960
rect 2945 2940 2965 2960
rect 2835 2770 2855 2790
rect 3260 3040 3280 3060
rect 4880 3040 4900 3060
rect 3980 2670 4000 2690
rect 4700 2670 4720 2690
rect 5190 2940 5210 2960
rect 5410 2940 5430 2960
rect 5300 2770 5320 2790
rect 2710 2180 2730 2200
rect 2800 2180 2820 2200
rect 2890 2180 2910 2200
rect 3130 2180 3150 2200
rect 3250 2180 3270 2200
rect 3490 2180 3510 2200
rect 3610 2180 3630 2200
rect 3820 2180 3840 2200
rect 3910 2180 3930 2200
rect 4230 2180 4250 2200
rect 4320 2180 4340 2200
rect 4530 2180 4550 2200
rect 4650 2180 4670 2200
rect 4890 2180 4910 2200
rect 5010 2180 5030 2200
rect 5250 2180 5270 2200
rect 5340 2180 5360 2200
rect 5430 2180 5450 2200
rect 3200 2020 3220 2040
rect 3140 1855 3160 1875
rect 4940 2020 4960 2040
rect 5000 1855 5020 1875
rect 2990 1695 3010 1715
rect 3110 1695 3130 1715
rect 3230 1695 3250 1715
rect 3350 1695 3370 1715
rect 3590 1695 3610 1715
rect 3710 1695 3730 1715
rect 3830 1695 3850 1715
rect 4310 1695 4330 1715
rect 4430 1695 4450 1715
rect 4550 1695 4570 1715
rect 4790 1695 4810 1715
rect 4910 1695 4930 1715
rect 5030 1695 5050 1715
rect 5150 1695 5170 1715
rect 3110 1230 3130 1250
rect 3190 1230 3210 1250
rect 3270 1230 3290 1250
rect 3350 1230 3370 1250
rect 3430 1230 3450 1250
rect 3510 1230 3530 1250
rect 3590 1230 3610 1250
rect 3670 1230 3690 1250
rect 3750 1230 3770 1250
rect 3830 1230 3850 1250
rect 3910 1230 3930 1250
rect 3990 1230 4010 1250
rect 4150 1230 4170 1250
rect 4230 1230 4250 1250
rect 4310 1230 4330 1250
rect 4390 1230 4410 1250
rect 4470 1230 4490 1250
rect 4550 1230 4570 1250
rect 4630 1230 4650 1250
rect 4710 1230 4730 1250
rect 4790 1230 4810 1250
rect 4870 1230 4890 1250
rect 4950 1230 4970 1250
rect 5030 1230 5050 1250
rect 3400 955 3420 975
rect 3125 785 3145 805
rect 3620 785 3640 805
rect 4070 955 4090 975
rect 3795 785 3815 805
rect 3875 785 3895 805
rect 4345 785 4365 805
rect 4740 955 4760 975
rect 4520 785 4540 805
rect 5015 785 5035 805
<< xpolycontact >>
rect 111 3555 331 3590
rect 945 3555 1165 3590
rect 111 3495 331 3530
rect 945 3495 1165 3530
rect 111 3290 331 3325
rect 915 3290 1135 3325
rect 111 3230 331 3265
rect 915 3230 1135 3265
rect 1396 3420 1616 3455
rect 2200 3420 2420 3455
rect 1396 3360 1616 3395
rect 2200 3360 2420 3395
rect 1396 3300 1616 3335
rect 2200 3300 2420 3335
rect 306 3025 525 3060
rect 714 3025 934 3060
rect 1396 3240 1616 3275
rect 2200 3240 2420 3275
rect 1396 3180 1616 3215
rect 2200 3180 2420 3215
rect 1396 3120 1616 3155
rect 2200 3120 2420 3155
rect 306 2815 525 2850
rect 714 2815 934 2850
rect 1561 2915 1781 2950
rect 1995 2915 2215 2950
<< ppolyres >>
rect 525 3025 714 3060
rect 525 2815 714 2850
<< xpolyres >>
rect 331 3555 945 3590
rect 331 3495 945 3530
rect 331 3290 915 3325
rect 331 3230 915 3265
rect 1616 3420 2200 3455
rect 1616 3360 2200 3395
rect 1616 3300 2200 3335
rect 1616 3240 2200 3275
rect 1616 3180 2200 3215
rect 1616 3120 2200 3155
rect 1781 2915 1995 2950
<< locali >>
rect 4445 3815 4475 3845
rect 945 3765 975 3795
rect 1645 3765 1675 3795
rect 5145 3765 5175 3795
rect 2695 3710 2725 3740
rect 3395 3710 3425 3740
rect 25 3640 590 3660
rect 670 3640 1235 3660
rect 25 3580 45 3640
rect 66 3585 111 3590
rect 66 3560 76 3585
rect 101 3560 111 3585
rect 66 3555 111 3560
rect 1130 3530 1165 3555
rect 25 3445 45 3500
rect 66 3525 111 3530
rect 66 3500 76 3525
rect 101 3500 111 3525
rect 66 3495 111 3500
rect 1215 3580 1235 3640
rect 2985 3555 3180 3575
rect 3260 3555 3455 3575
rect 1215 3445 1235 3500
rect 25 3425 590 3445
rect 670 3425 1235 3445
rect 1310 3505 1845 3525
rect 1925 3505 2505 3525
rect 615 3395 635 3425
rect 25 3375 575 3395
rect 655 3375 1205 3395
rect 25 3315 45 3375
rect 66 3320 111 3325
rect 66 3295 76 3320
rect 101 3295 111 3320
rect 66 3290 111 3295
rect 1100 3265 1135 3290
rect 25 3180 45 3235
rect 66 3260 111 3265
rect 66 3235 76 3260
rect 101 3235 111 3260
rect 66 3230 111 3235
rect 1185 3315 1205 3375
rect 1310 3325 1330 3505
rect 1351 3450 1396 3455
rect 1351 3425 1361 3450
rect 1386 3425 1396 3450
rect 1351 3420 1396 3425
rect 2420 3420 2460 3455
rect 1351 3390 1396 3395
rect 1351 3365 1361 3390
rect 1386 3365 1396 3390
rect 1351 3360 1396 3365
rect 2385 3335 2420 3360
rect 1205 3285 1225 3295
rect 1215 3265 1225 3285
rect 1205 3255 1225 3265
rect 1290 3285 1310 3295
rect 1290 3265 1300 3285
rect 1290 3255 1310 3265
rect 595 3190 635 3200
rect 595 3180 605 3190
rect 625 3180 635 3190
rect 1185 3180 1205 3235
rect 25 3160 575 3180
rect 655 3160 1205 3180
rect 605 3130 625 3160
rect 220 3110 575 3130
rect 655 3110 1020 3130
rect 220 3080 240 3110
rect 1000 3080 1020 3110
rect 261 3055 306 3060
rect 261 3030 271 3055
rect 296 3030 306 3055
rect 261 3025 306 3030
rect 934 3055 979 3060
rect 934 3030 944 3055
rect 969 3030 979 3055
rect 934 3025 979 3030
rect 220 2970 240 3000
rect 1310 3070 1330 3245
rect 1356 3300 1396 3335
rect 1356 3155 1376 3300
rect 2440 3275 2460 3420
rect 2420 3240 2460 3275
rect 2485 3325 2505 3505
rect 2985 3470 3005 3555
rect 3045 3535 3065 3555
rect 3375 3535 3395 3555
rect 3035 3525 3075 3535
rect 3035 3505 3045 3525
rect 3065 3505 3075 3525
rect 3035 3495 3075 3505
rect 3145 3525 3185 3535
rect 3145 3505 3155 3525
rect 3175 3505 3185 3525
rect 3145 3495 3185 3505
rect 3205 3525 3235 3535
rect 3205 3505 3210 3525
rect 3230 3505 3235 3525
rect 3205 3495 3235 3505
rect 3255 3525 3295 3535
rect 3255 3505 3265 3525
rect 3285 3505 3295 3525
rect 3255 3495 3295 3505
rect 3315 3525 3345 3535
rect 3315 3505 3320 3525
rect 3340 3505 3345 3525
rect 3315 3495 3345 3505
rect 3365 3525 3405 3535
rect 3365 3505 3375 3525
rect 3395 3505 3405 3525
rect 3365 3495 3405 3505
rect 3045 3475 3065 3495
rect 3155 3475 3175 3495
rect 3265 3475 3285 3495
rect 3320 3475 3340 3495
rect 3375 3475 3395 3495
rect 2985 3305 3005 3390
rect 3040 3465 3070 3475
rect 3040 3393 3045 3465
rect 3065 3393 3070 3465
rect 3040 3385 3070 3393
rect 3095 3465 3125 3475
rect 3095 3393 3100 3465
rect 3120 3393 3125 3465
rect 3095 3385 3125 3393
rect 3150 3465 3180 3475
rect 3150 3393 3155 3465
rect 3175 3393 3180 3465
rect 3150 3385 3180 3393
rect 3205 3465 3235 3475
rect 3205 3393 3210 3465
rect 3230 3393 3235 3465
rect 3205 3385 3235 3393
rect 3260 3465 3290 3475
rect 3260 3393 3265 3465
rect 3285 3393 3290 3465
rect 3260 3385 3290 3393
rect 3315 3465 3345 3475
rect 3315 3393 3320 3465
rect 3340 3393 3345 3465
rect 3315 3385 3345 3393
rect 3370 3465 3400 3475
rect 3370 3393 3375 3465
rect 3395 3393 3400 3465
rect 3370 3385 3400 3393
rect 3435 3470 3455 3555
rect 3100 3365 3120 3385
rect 3210 3365 3230 3385
rect 3320 3365 3340 3385
rect 3090 3355 3130 3365
rect 3090 3335 3100 3355
rect 3120 3335 3130 3355
rect 3090 3325 3130 3335
rect 3200 3355 3240 3365
rect 3200 3335 3210 3355
rect 3230 3335 3240 3355
rect 3200 3325 3240 3335
rect 3310 3355 3350 3365
rect 3310 3335 3320 3355
rect 3340 3335 3350 3355
rect 3310 3325 3350 3335
rect 3435 3305 3455 3390
rect 2985 3285 3180 3305
rect 3260 3285 3455 3305
rect 3625 3555 4040 3575
rect 4120 3555 4535 3575
rect 3625 3470 3645 3555
rect 3685 3535 3705 3555
rect 4455 3535 4475 3555
rect 3675 3525 3715 3535
rect 3675 3505 3685 3525
rect 3705 3505 3715 3525
rect 3675 3495 3715 3505
rect 3785 3525 3825 3535
rect 3785 3505 3795 3525
rect 3815 3505 3825 3525
rect 3785 3495 3825 3505
rect 3895 3525 3935 3535
rect 3895 3505 3905 3525
rect 3925 3505 3935 3525
rect 3895 3495 3935 3505
rect 4005 3525 4045 3535
rect 4005 3505 4015 3525
rect 4035 3505 4045 3525
rect 4005 3495 4045 3505
rect 4065 3525 4095 3535
rect 4065 3505 4070 3525
rect 4090 3505 4095 3525
rect 4065 3495 4095 3505
rect 4115 3525 4155 3535
rect 4115 3505 4125 3525
rect 4145 3505 4155 3525
rect 4115 3495 4155 3505
rect 4225 3525 4265 3535
rect 4225 3505 4235 3525
rect 4255 3505 4265 3525
rect 4225 3495 4265 3505
rect 4335 3525 4375 3535
rect 4335 3505 4345 3525
rect 4365 3505 4375 3525
rect 4335 3495 4375 3505
rect 4395 3525 4425 3535
rect 4395 3505 4400 3525
rect 4420 3505 4425 3525
rect 4395 3495 4425 3505
rect 4445 3525 4485 3535
rect 4445 3505 4455 3525
rect 4475 3505 4485 3525
rect 4445 3495 4485 3505
rect 3685 3475 3705 3495
rect 3795 3475 3815 3495
rect 3905 3475 3925 3495
rect 4015 3475 4035 3495
rect 4125 3475 4145 3495
rect 4235 3475 4255 3495
rect 4345 3475 4365 3495
rect 4400 3475 4420 3495
rect 4455 3475 4475 3495
rect 3625 3305 3645 3390
rect 3680 3465 3710 3475
rect 3680 3445 3685 3465
rect 3705 3445 3710 3465
rect 3680 3415 3710 3445
rect 3680 3395 3685 3415
rect 3705 3395 3710 3415
rect 3680 3385 3710 3395
rect 3735 3465 3765 3475
rect 3735 3445 3740 3465
rect 3760 3445 3765 3465
rect 3735 3415 3765 3445
rect 3735 3395 3740 3415
rect 3760 3395 3765 3415
rect 3735 3385 3765 3395
rect 3790 3465 3820 3475
rect 3790 3445 3795 3465
rect 3815 3445 3820 3465
rect 3790 3415 3820 3445
rect 3790 3395 3795 3415
rect 3815 3395 3820 3415
rect 3790 3385 3820 3395
rect 3845 3465 3875 3475
rect 3845 3445 3850 3465
rect 3870 3445 3875 3465
rect 3845 3415 3875 3445
rect 3845 3395 3850 3415
rect 3870 3395 3875 3415
rect 3845 3385 3875 3395
rect 3900 3465 3930 3475
rect 3900 3445 3905 3465
rect 3925 3445 3930 3465
rect 3900 3415 3930 3445
rect 3900 3395 3905 3415
rect 3925 3395 3930 3415
rect 3900 3385 3930 3395
rect 3955 3465 3985 3475
rect 3955 3445 3960 3465
rect 3980 3445 3985 3465
rect 3955 3415 3985 3445
rect 3955 3395 3960 3415
rect 3980 3395 3985 3415
rect 3955 3385 3985 3395
rect 4010 3465 4040 3475
rect 4010 3445 4015 3465
rect 4035 3445 4040 3465
rect 4010 3415 4040 3445
rect 4010 3395 4015 3415
rect 4035 3395 4040 3415
rect 4010 3385 4040 3395
rect 4065 3465 4095 3475
rect 4065 3445 4070 3465
rect 4090 3445 4095 3465
rect 4065 3415 4095 3445
rect 4065 3395 4070 3415
rect 4090 3395 4095 3415
rect 4065 3385 4095 3395
rect 4120 3465 4150 3475
rect 4120 3445 4125 3465
rect 4145 3445 4150 3465
rect 4120 3415 4150 3445
rect 4120 3395 4125 3415
rect 4145 3395 4150 3415
rect 4120 3385 4150 3395
rect 4175 3465 4205 3475
rect 4175 3445 4180 3465
rect 4200 3445 4205 3465
rect 4175 3415 4205 3445
rect 4175 3395 4180 3415
rect 4200 3395 4205 3415
rect 4175 3385 4205 3395
rect 4230 3465 4260 3475
rect 4230 3445 4235 3465
rect 4255 3445 4260 3465
rect 4230 3415 4260 3445
rect 4230 3395 4235 3415
rect 4255 3395 4260 3415
rect 4230 3385 4260 3395
rect 4285 3465 4315 3475
rect 4285 3445 4290 3465
rect 4310 3445 4315 3465
rect 4285 3415 4315 3445
rect 4285 3395 4290 3415
rect 4310 3395 4315 3415
rect 4285 3385 4315 3395
rect 4340 3465 4370 3475
rect 4340 3445 4345 3465
rect 4365 3445 4370 3465
rect 4340 3415 4370 3445
rect 4340 3395 4345 3415
rect 4365 3395 4370 3415
rect 4340 3385 4370 3395
rect 4395 3465 4425 3475
rect 4395 3445 4400 3465
rect 4420 3445 4425 3465
rect 4395 3415 4425 3445
rect 4395 3395 4400 3415
rect 4420 3395 4425 3415
rect 4395 3385 4425 3395
rect 4450 3465 4480 3475
rect 4450 3445 4455 3465
rect 4475 3445 4480 3465
rect 4450 3415 4480 3445
rect 4450 3395 4455 3415
rect 4475 3395 4480 3415
rect 4450 3385 4480 3395
rect 4515 3470 4535 3555
rect 3740 3365 3760 3385
rect 3850 3365 3870 3385
rect 3960 3365 3980 3385
rect 4070 3365 4090 3385
rect 4180 3365 4200 3385
rect 4290 3365 4310 3385
rect 4400 3365 4420 3385
rect 3730 3355 3770 3365
rect 3730 3335 3740 3355
rect 3760 3335 3770 3355
rect 3730 3325 3770 3335
rect 3840 3355 3880 3365
rect 3840 3335 3850 3355
rect 3870 3335 3880 3355
rect 3840 3325 3880 3335
rect 3950 3355 3990 3365
rect 3950 3335 3960 3355
rect 3980 3335 3990 3355
rect 3950 3325 3990 3335
rect 4060 3355 4100 3365
rect 4060 3335 4070 3355
rect 4090 3335 4100 3355
rect 4060 3325 4100 3335
rect 4170 3355 4210 3365
rect 4170 3335 4180 3355
rect 4200 3335 4210 3355
rect 4170 3325 4210 3335
rect 4280 3355 4320 3365
rect 4280 3335 4290 3355
rect 4310 3335 4320 3355
rect 4280 3325 4320 3335
rect 4390 3355 4430 3365
rect 4390 3335 4400 3355
rect 4420 3335 4430 3355
rect 4390 3325 4430 3335
rect 4515 3305 4535 3390
rect 3625 3285 4040 3305
rect 4120 3285 4535 3305
rect 4705 3555 4900 3575
rect 4980 3555 5175 3575
rect 4705 3470 4725 3555
rect 4765 3535 4785 3555
rect 5095 3535 5115 3555
rect 4755 3525 4795 3535
rect 4755 3505 4765 3525
rect 4785 3505 4795 3525
rect 4755 3495 4795 3505
rect 4865 3525 4905 3535
rect 4865 3505 4875 3525
rect 4895 3505 4905 3525
rect 4865 3495 4905 3505
rect 4925 3525 4955 3535
rect 4925 3505 4930 3525
rect 4950 3505 4955 3525
rect 4925 3495 4955 3505
rect 4975 3525 5015 3535
rect 4975 3505 4985 3525
rect 5005 3505 5015 3525
rect 4975 3495 5015 3505
rect 5085 3525 5125 3535
rect 5085 3505 5095 3525
rect 5115 3505 5125 3525
rect 5085 3495 5125 3505
rect 4765 3475 4785 3495
rect 4875 3475 4895 3495
rect 4985 3475 5005 3495
rect 5095 3475 5115 3495
rect 4705 3305 4725 3390
rect 4760 3465 4790 3475
rect 4760 3395 4765 3465
rect 4785 3395 4790 3465
rect 4760 3385 4790 3395
rect 4815 3465 4845 3475
rect 4815 3395 4820 3465
rect 4840 3395 4845 3465
rect 4815 3385 4845 3395
rect 4870 3465 4900 3475
rect 4870 3395 4875 3465
rect 4895 3395 4900 3465
rect 4870 3385 4900 3395
rect 4925 3465 4955 3475
rect 4925 3395 4930 3465
rect 4950 3395 4955 3465
rect 4925 3385 4955 3395
rect 4980 3465 5010 3475
rect 4980 3395 4985 3465
rect 5005 3395 5010 3465
rect 4980 3385 5010 3395
rect 5035 3465 5065 3475
rect 5035 3395 5040 3465
rect 5060 3395 5065 3465
rect 5035 3385 5065 3395
rect 5090 3465 5120 3475
rect 5090 3395 5095 3465
rect 5115 3395 5120 3465
rect 5090 3385 5120 3395
rect 5155 3470 5175 3555
rect 4820 3365 4840 3385
rect 4930 3365 4950 3385
rect 5040 3365 5060 3385
rect 4810 3355 4850 3365
rect 4810 3335 4820 3355
rect 4840 3335 4850 3355
rect 4810 3325 4850 3335
rect 4920 3355 4960 3365
rect 4920 3335 4930 3355
rect 4950 3335 4960 3355
rect 4920 3325 4960 3335
rect 5030 3355 5070 3365
rect 5030 3335 5040 3355
rect 5060 3335 5070 3355
rect 5030 3325 5070 3335
rect 5155 3305 5175 3390
rect 4705 3285 4900 3305
rect 4965 3285 5175 3305
rect 1396 3215 1431 3240
rect 2420 3210 2465 3215
rect 2420 3185 2430 3210
rect 2455 3185 2465 3210
rect 2420 3180 2465 3185
rect 1356 3120 1396 3155
rect 2420 3150 2465 3160
rect 2420 3125 2430 3150
rect 2455 3125 2465 3150
rect 2420 3115 2465 3125
rect 2485 3070 2505 3245
rect 1310 3050 1845 3070
rect 1925 3050 2505 3070
rect 3200 3090 4040 3110
rect 4120 3090 4960 3110
rect 1875 3020 1895 3050
rect 2825 3020 2865 3030
rect 1000 2970 1020 3000
rect 220 2950 575 2970
rect 655 2950 1020 2970
rect 1475 3000 1845 3020
rect 1925 3000 2300 3020
rect 2825 3010 2835 3020
rect 2855 3010 2865 3020
rect 1475 2970 1495 3000
rect 605 2920 625 2950
rect 220 2900 575 2920
rect 655 2900 1020 2920
rect 220 2870 240 2900
rect 1000 2870 1020 2900
rect 261 2845 306 2850
rect 261 2820 271 2845
rect 296 2820 306 2845
rect 261 2815 306 2820
rect 934 2845 979 2850
rect 934 2820 944 2845
rect 969 2820 979 2845
rect 934 2815 979 2820
rect 220 2760 240 2790
rect 2280 2970 2300 3000
rect 1516 2945 1561 2950
rect 1516 2920 1526 2945
rect 1551 2920 1561 2945
rect 1516 2915 1561 2920
rect 2215 2945 2260 2950
rect 2215 2920 2225 2945
rect 2250 2920 2260 2945
rect 2215 2915 2260 2920
rect 1475 2865 1495 2890
rect 2280 2865 2300 2890
rect 1475 2845 1845 2865
rect 1925 2845 2300 2865
rect 2665 2990 2805 3010
rect 2885 2990 3025 3010
rect 2665 2905 2685 2990
rect 2725 2970 2745 2990
rect 2945 2970 2965 2990
rect 1000 2760 1020 2790
rect 220 2740 575 2760
rect 655 2740 1020 2760
rect 2665 2740 2685 2825
rect 2720 2960 2750 2970
rect 2720 2940 2725 2960
rect 2745 2940 2750 2960
rect 2720 2900 2750 2940
rect 2825 2960 2865 2970
rect 2825 2940 2835 2960
rect 2855 2940 2865 2960
rect 2825 2930 2865 2940
rect 2940 2960 2970 2970
rect 2940 2940 2945 2960
rect 2965 2940 2970 2960
rect 2835 2910 2855 2930
rect 2720 2880 2725 2900
rect 2745 2880 2750 2900
rect 2720 2850 2750 2880
rect 2720 2830 2725 2850
rect 2745 2830 2750 2850
rect 2720 2820 2750 2830
rect 2775 2900 2805 2910
rect 2775 2880 2780 2900
rect 2800 2880 2805 2900
rect 2775 2850 2805 2880
rect 2775 2830 2780 2850
rect 2800 2830 2805 2850
rect 2775 2820 2805 2830
rect 2830 2900 2860 2910
rect 2830 2880 2835 2900
rect 2855 2880 2860 2900
rect 2830 2850 2860 2880
rect 2830 2830 2835 2850
rect 2855 2830 2860 2850
rect 2830 2820 2860 2830
rect 2885 2900 2915 2910
rect 2885 2880 2890 2900
rect 2910 2880 2915 2900
rect 2885 2850 2915 2880
rect 2885 2830 2890 2850
rect 2910 2830 2915 2850
rect 2885 2820 2915 2830
rect 2940 2900 2970 2940
rect 2940 2880 2945 2900
rect 2965 2880 2970 2900
rect 2940 2850 2970 2880
rect 2940 2830 2945 2850
rect 2965 2830 2970 2850
rect 2940 2820 2970 2830
rect 3005 2905 3025 2990
rect 2780 2800 2800 2820
rect 2890 2800 2910 2820
rect 2760 2790 2800 2800
rect 2760 2770 2770 2790
rect 2790 2770 2800 2790
rect 2760 2760 2800 2770
rect 2825 2790 2865 2800
rect 2825 2770 2835 2790
rect 2855 2770 2865 2790
rect 2825 2760 2865 2770
rect 2890 2790 2930 2800
rect 2890 2770 2900 2790
rect 2920 2770 2930 2790
rect 2890 2760 2930 2770
rect 3005 2740 3025 2825
rect 2665 2720 2805 2740
rect 2885 2720 3025 2740
rect 3200 2905 3220 3090
rect 3260 3070 3280 3090
rect 4880 3070 4900 3090
rect 3250 3060 3290 3070
rect 3250 3040 3260 3060
rect 3280 3040 3290 3060
rect 3250 3030 3290 3040
rect 3430 3060 3470 3070
rect 3430 3040 3440 3060
rect 3460 3040 3470 3060
rect 3430 3030 3470 3040
rect 3610 3060 3650 3070
rect 3610 3040 3620 3060
rect 3640 3040 3650 3060
rect 3610 3030 3650 3040
rect 3790 3060 3830 3070
rect 3790 3040 3800 3060
rect 3820 3040 3830 3060
rect 3790 3030 3830 3040
rect 3970 3060 4010 3070
rect 3970 3040 3980 3060
rect 4000 3040 4010 3060
rect 3970 3030 4010 3040
rect 4150 3060 4190 3070
rect 4150 3040 4160 3060
rect 4180 3040 4190 3060
rect 4150 3030 4190 3040
rect 4330 3060 4370 3070
rect 4330 3040 4340 3060
rect 4360 3040 4370 3060
rect 4330 3030 4370 3040
rect 4510 3060 4550 3070
rect 4510 3040 4520 3060
rect 4540 3040 4550 3060
rect 4510 3030 4550 3040
rect 4690 3060 4730 3070
rect 4690 3040 4700 3060
rect 4720 3040 4730 3060
rect 4690 3030 4730 3040
rect 4870 3060 4910 3070
rect 4870 3040 4880 3060
rect 4900 3040 4910 3060
rect 4870 3030 4910 3040
rect 3260 3010 3280 3030
rect 3440 3010 3460 3030
rect 3620 3010 3640 3030
rect 3800 3010 3820 3030
rect 3980 3010 4000 3030
rect 4160 3010 4180 3030
rect 4340 3010 4360 3030
rect 4520 3010 4540 3030
rect 4700 3010 4720 3030
rect 4880 3010 4900 3030
rect 650 2055 775 2700
rect 1330 2055 1455 2700
rect 2010 2055 2135 2700
rect 3200 2635 3220 2825
rect 3255 3000 3285 3010
rect 3255 2980 3260 3000
rect 3280 2980 3285 3000
rect 3255 2950 3285 2980
rect 3255 2930 3260 2950
rect 3280 2930 3285 2950
rect 3255 2900 3285 2930
rect 3255 2880 3260 2900
rect 3280 2880 3285 2900
rect 3255 2850 3285 2880
rect 3255 2830 3260 2850
rect 3280 2830 3285 2850
rect 3255 2800 3285 2830
rect 3255 2780 3260 2800
rect 3280 2780 3285 2800
rect 3255 2750 3285 2780
rect 3255 2730 3260 2750
rect 3280 2730 3285 2750
rect 3255 2720 3285 2730
rect 3345 3000 3375 3010
rect 3345 2980 3350 3000
rect 3370 2980 3375 3000
rect 3345 2950 3375 2980
rect 3345 2930 3350 2950
rect 3370 2930 3375 2950
rect 3345 2900 3375 2930
rect 3345 2880 3350 2900
rect 3370 2880 3375 2900
rect 3345 2850 3375 2880
rect 3345 2830 3350 2850
rect 3370 2830 3375 2850
rect 3345 2800 3375 2830
rect 3345 2780 3350 2800
rect 3370 2780 3375 2800
rect 3345 2750 3375 2780
rect 3345 2730 3350 2750
rect 3370 2730 3375 2750
rect 3345 2720 3375 2730
rect 3435 3000 3465 3010
rect 3435 2980 3440 3000
rect 3460 2980 3465 3000
rect 3435 2950 3465 2980
rect 3435 2930 3440 2950
rect 3460 2930 3465 2950
rect 3435 2900 3465 2930
rect 3435 2880 3440 2900
rect 3460 2880 3465 2900
rect 3435 2850 3465 2880
rect 3435 2830 3440 2850
rect 3460 2830 3465 2850
rect 3435 2800 3465 2830
rect 3435 2780 3440 2800
rect 3460 2780 3465 2800
rect 3435 2750 3465 2780
rect 3435 2730 3440 2750
rect 3460 2730 3465 2750
rect 3435 2720 3465 2730
rect 3525 3000 3555 3010
rect 3525 2980 3530 3000
rect 3550 2980 3555 3000
rect 3525 2950 3555 2980
rect 3525 2930 3530 2950
rect 3550 2930 3555 2950
rect 3525 2900 3555 2930
rect 3525 2880 3530 2900
rect 3550 2880 3555 2900
rect 3525 2850 3555 2880
rect 3525 2830 3530 2850
rect 3550 2830 3555 2850
rect 3525 2800 3555 2830
rect 3525 2780 3530 2800
rect 3550 2780 3555 2800
rect 3525 2750 3555 2780
rect 3525 2730 3530 2750
rect 3550 2730 3555 2750
rect 3525 2720 3555 2730
rect 3615 3000 3645 3010
rect 3615 2980 3620 3000
rect 3640 2980 3645 3000
rect 3615 2950 3645 2980
rect 3615 2930 3620 2950
rect 3640 2930 3645 2950
rect 3615 2900 3645 2930
rect 3615 2880 3620 2900
rect 3640 2880 3645 2900
rect 3615 2850 3645 2880
rect 3615 2830 3620 2850
rect 3640 2830 3645 2850
rect 3615 2800 3645 2830
rect 3615 2780 3620 2800
rect 3640 2780 3645 2800
rect 3615 2750 3645 2780
rect 3615 2730 3620 2750
rect 3640 2730 3645 2750
rect 3615 2720 3645 2730
rect 3705 3000 3735 3010
rect 3705 2980 3710 3000
rect 3730 2980 3735 3000
rect 3705 2950 3735 2980
rect 3705 2930 3710 2950
rect 3730 2930 3735 2950
rect 3705 2900 3735 2930
rect 3705 2880 3710 2900
rect 3730 2880 3735 2900
rect 3705 2850 3735 2880
rect 3705 2830 3710 2850
rect 3730 2830 3735 2850
rect 3705 2800 3735 2830
rect 3705 2780 3710 2800
rect 3730 2780 3735 2800
rect 3705 2750 3735 2780
rect 3705 2730 3710 2750
rect 3730 2730 3735 2750
rect 3705 2720 3735 2730
rect 3795 3000 3825 3010
rect 3795 2980 3800 3000
rect 3820 2980 3825 3000
rect 3795 2950 3825 2980
rect 3795 2930 3800 2950
rect 3820 2930 3825 2950
rect 3795 2900 3825 2930
rect 3795 2880 3800 2900
rect 3820 2880 3825 2900
rect 3795 2850 3825 2880
rect 3795 2830 3800 2850
rect 3820 2830 3825 2850
rect 3795 2800 3825 2830
rect 3795 2780 3800 2800
rect 3820 2780 3825 2800
rect 3795 2750 3825 2780
rect 3795 2730 3800 2750
rect 3820 2730 3825 2750
rect 3795 2720 3825 2730
rect 3885 3000 3915 3010
rect 3885 2980 3890 3000
rect 3910 2980 3915 3000
rect 3885 2950 3915 2980
rect 3885 2930 3890 2950
rect 3910 2930 3915 2950
rect 3885 2900 3915 2930
rect 3885 2880 3890 2900
rect 3910 2880 3915 2900
rect 3885 2850 3915 2880
rect 3885 2830 3890 2850
rect 3910 2830 3915 2850
rect 3885 2800 3915 2830
rect 3885 2780 3890 2800
rect 3910 2780 3915 2800
rect 3885 2750 3915 2780
rect 3885 2730 3890 2750
rect 3910 2730 3915 2750
rect 3885 2720 3915 2730
rect 3975 3000 4005 3010
rect 3975 2980 3980 3000
rect 4000 2980 4005 3000
rect 3975 2950 4005 2980
rect 3975 2930 3980 2950
rect 4000 2930 4005 2950
rect 3975 2900 4005 2930
rect 3975 2880 3980 2900
rect 4000 2880 4005 2900
rect 3975 2850 4005 2880
rect 3975 2830 3980 2850
rect 4000 2830 4005 2850
rect 3975 2800 4005 2830
rect 3975 2780 3980 2800
rect 4000 2780 4005 2800
rect 3975 2750 4005 2780
rect 3975 2730 3980 2750
rect 4000 2730 4005 2750
rect 3975 2720 4005 2730
rect 4065 3000 4095 3010
rect 4065 2980 4070 3000
rect 4090 2980 4095 3000
rect 4065 2950 4095 2980
rect 4065 2930 4070 2950
rect 4090 2930 4095 2950
rect 4065 2900 4095 2930
rect 4065 2880 4070 2900
rect 4090 2880 4095 2900
rect 4065 2850 4095 2880
rect 4065 2830 4070 2850
rect 4090 2830 4095 2850
rect 4065 2800 4095 2830
rect 4065 2780 4070 2800
rect 4090 2780 4095 2800
rect 4065 2750 4095 2780
rect 4065 2730 4070 2750
rect 4090 2730 4095 2750
rect 4065 2720 4095 2730
rect 4155 3000 4185 3010
rect 4155 2980 4160 3000
rect 4180 2980 4185 3000
rect 4155 2950 4185 2980
rect 4155 2930 4160 2950
rect 4180 2930 4185 2950
rect 4155 2900 4185 2930
rect 4155 2880 4160 2900
rect 4180 2880 4185 2900
rect 4155 2850 4185 2880
rect 4155 2830 4160 2850
rect 4180 2830 4185 2850
rect 4155 2800 4185 2830
rect 4155 2780 4160 2800
rect 4180 2780 4185 2800
rect 4155 2750 4185 2780
rect 4155 2730 4160 2750
rect 4180 2730 4185 2750
rect 4155 2720 4185 2730
rect 4245 3000 4275 3010
rect 4245 2980 4250 3000
rect 4270 2980 4275 3000
rect 4245 2950 4275 2980
rect 4245 2930 4250 2950
rect 4270 2930 4275 2950
rect 4245 2900 4275 2930
rect 4245 2880 4250 2900
rect 4270 2880 4275 2900
rect 4245 2850 4275 2880
rect 4245 2830 4250 2850
rect 4270 2830 4275 2850
rect 4245 2800 4275 2830
rect 4245 2780 4250 2800
rect 4270 2780 4275 2800
rect 4245 2750 4275 2780
rect 4245 2730 4250 2750
rect 4270 2730 4275 2750
rect 4245 2720 4275 2730
rect 4335 3000 4365 3010
rect 4335 2980 4340 3000
rect 4360 2980 4365 3000
rect 4335 2950 4365 2980
rect 4335 2930 4340 2950
rect 4360 2930 4365 2950
rect 4335 2900 4365 2930
rect 4335 2880 4340 2900
rect 4360 2880 4365 2900
rect 4335 2850 4365 2880
rect 4335 2830 4340 2850
rect 4360 2830 4365 2850
rect 4335 2800 4365 2830
rect 4335 2780 4340 2800
rect 4360 2780 4365 2800
rect 4335 2750 4365 2780
rect 4335 2730 4340 2750
rect 4360 2730 4365 2750
rect 4335 2720 4365 2730
rect 4425 3000 4455 3010
rect 4425 2980 4430 3000
rect 4450 2980 4455 3000
rect 4425 2950 4455 2980
rect 4425 2930 4430 2950
rect 4450 2930 4455 2950
rect 4425 2900 4455 2930
rect 4425 2880 4430 2900
rect 4450 2880 4455 2900
rect 4425 2850 4455 2880
rect 4425 2830 4430 2850
rect 4450 2830 4455 2850
rect 4425 2800 4455 2830
rect 4425 2780 4430 2800
rect 4450 2780 4455 2800
rect 4425 2750 4455 2780
rect 4425 2730 4430 2750
rect 4450 2730 4455 2750
rect 4425 2720 4455 2730
rect 4515 3000 4545 3010
rect 4515 2980 4520 3000
rect 4540 2980 4545 3000
rect 4515 2950 4545 2980
rect 4515 2930 4520 2950
rect 4540 2930 4545 2950
rect 4515 2900 4545 2930
rect 4515 2880 4520 2900
rect 4540 2880 4545 2900
rect 4515 2850 4545 2880
rect 4515 2830 4520 2850
rect 4540 2830 4545 2850
rect 4515 2800 4545 2830
rect 4515 2780 4520 2800
rect 4540 2780 4545 2800
rect 4515 2750 4545 2780
rect 4515 2730 4520 2750
rect 4540 2730 4545 2750
rect 4515 2720 4545 2730
rect 4605 3000 4635 3010
rect 4605 2980 4610 3000
rect 4630 2980 4635 3000
rect 4605 2950 4635 2980
rect 4605 2930 4610 2950
rect 4630 2930 4635 2950
rect 4605 2900 4635 2930
rect 4605 2880 4610 2900
rect 4630 2880 4635 2900
rect 4605 2850 4635 2880
rect 4605 2830 4610 2850
rect 4630 2830 4635 2850
rect 4605 2800 4635 2830
rect 4605 2780 4610 2800
rect 4630 2780 4635 2800
rect 4605 2750 4635 2780
rect 4605 2730 4610 2750
rect 4630 2730 4635 2750
rect 4605 2720 4635 2730
rect 4695 3000 4725 3010
rect 4695 2980 4700 3000
rect 4720 2980 4725 3000
rect 4695 2950 4725 2980
rect 4695 2930 4700 2950
rect 4720 2930 4725 2950
rect 4695 2900 4725 2930
rect 4695 2880 4700 2900
rect 4720 2880 4725 2900
rect 4695 2850 4725 2880
rect 4695 2830 4700 2850
rect 4720 2830 4725 2850
rect 4695 2800 4725 2830
rect 4695 2780 4700 2800
rect 4720 2780 4725 2800
rect 4695 2750 4725 2780
rect 4695 2730 4700 2750
rect 4720 2730 4725 2750
rect 4695 2720 4725 2730
rect 4785 3000 4815 3010
rect 4785 2980 4790 3000
rect 4810 2980 4815 3000
rect 4785 2950 4815 2980
rect 4785 2930 4790 2950
rect 4810 2930 4815 2950
rect 4785 2900 4815 2930
rect 4785 2880 4790 2900
rect 4810 2880 4815 2900
rect 4785 2850 4815 2880
rect 4785 2830 4790 2850
rect 4810 2830 4815 2850
rect 4785 2800 4815 2830
rect 4785 2780 4790 2800
rect 4810 2780 4815 2800
rect 4785 2750 4815 2780
rect 4785 2730 4790 2750
rect 4810 2730 4815 2750
rect 4785 2720 4815 2730
rect 4875 3000 4905 3010
rect 4875 2980 4880 3000
rect 4900 2980 4905 3000
rect 4875 2950 4905 2980
rect 4875 2930 4880 2950
rect 4900 2930 4905 2950
rect 4875 2900 4905 2930
rect 4875 2880 4880 2900
rect 4900 2880 4905 2900
rect 4875 2850 4905 2880
rect 4875 2830 4880 2850
rect 4900 2830 4905 2850
rect 4875 2800 4905 2830
rect 4875 2780 4880 2800
rect 4900 2780 4905 2800
rect 4875 2750 4905 2780
rect 4875 2730 4880 2750
rect 4900 2730 4905 2750
rect 4875 2720 4905 2730
rect 4940 2905 4960 3090
rect 5290 3020 5330 3040
rect 5290 3010 5300 3020
rect 5320 3010 5330 3020
rect 3350 2700 3370 2720
rect 3530 2700 3550 2720
rect 3710 2700 3730 2720
rect 3890 2700 3910 2720
rect 4070 2700 4090 2720
rect 4250 2700 4270 2720
rect 4430 2700 4450 2720
rect 4610 2700 4630 2720
rect 4790 2700 4810 2720
rect 3340 2690 3380 2700
rect 3340 2670 3350 2690
rect 3370 2670 3380 2690
rect 3340 2660 3380 2670
rect 3520 2690 3560 2700
rect 3520 2670 3530 2690
rect 3550 2670 3560 2690
rect 3520 2660 3560 2670
rect 3700 2690 3740 2700
rect 3700 2670 3710 2690
rect 3730 2670 3740 2690
rect 3700 2660 3740 2670
rect 3880 2690 3920 2700
rect 3880 2670 3890 2690
rect 3910 2670 3920 2690
rect 3880 2660 3920 2670
rect 3970 2690 4010 2700
rect 3970 2670 3980 2690
rect 4000 2670 4010 2690
rect 3970 2660 4010 2670
rect 4060 2690 4100 2700
rect 4060 2670 4070 2690
rect 4090 2670 4100 2690
rect 4060 2660 4100 2670
rect 4240 2690 4280 2700
rect 4240 2670 4250 2690
rect 4270 2670 4280 2690
rect 4240 2660 4280 2670
rect 4420 2690 4460 2700
rect 4420 2670 4430 2690
rect 4450 2670 4460 2690
rect 4420 2660 4460 2670
rect 4600 2690 4640 2700
rect 4600 2670 4610 2690
rect 4630 2670 4640 2690
rect 4600 2660 4640 2670
rect 4690 2690 4730 2700
rect 4690 2670 4700 2690
rect 4720 2670 4730 2690
rect 4690 2660 4730 2670
rect 4780 2690 4820 2700
rect 4780 2670 4790 2690
rect 4810 2670 4820 2690
rect 4780 2660 4820 2670
rect 4940 2635 4960 2825
rect 5130 2990 5270 3010
rect 5350 2990 5490 3010
rect 5130 2905 5150 2990
rect 5190 2970 5210 2990
rect 5410 2970 5430 2990
rect 5185 2960 5215 2970
rect 5185 2940 5190 2960
rect 5210 2940 5215 2960
rect 5185 2930 5215 2940
rect 5290 2960 5330 2970
rect 5290 2940 5300 2960
rect 5320 2940 5330 2960
rect 5290 2930 5330 2940
rect 5405 2960 5435 2970
rect 5405 2940 5410 2960
rect 5430 2940 5435 2960
rect 5405 2930 5435 2940
rect 5190 2910 5210 2930
rect 5300 2910 5320 2930
rect 5410 2910 5430 2930
rect 5130 2740 5150 2825
rect 5185 2900 5215 2910
rect 5185 2880 5190 2900
rect 5210 2880 5215 2900
rect 5185 2850 5215 2880
rect 5185 2830 5190 2850
rect 5210 2830 5215 2850
rect 5185 2820 5215 2830
rect 5240 2900 5270 2910
rect 5240 2880 5245 2900
rect 5265 2880 5270 2900
rect 5240 2850 5270 2880
rect 5240 2830 5245 2850
rect 5265 2830 5270 2850
rect 5240 2820 5270 2830
rect 5295 2900 5325 2910
rect 5295 2880 5300 2900
rect 5320 2880 5325 2900
rect 5295 2850 5325 2880
rect 5295 2830 5300 2850
rect 5320 2830 5325 2850
rect 5295 2820 5325 2830
rect 5350 2900 5380 2910
rect 5350 2880 5355 2900
rect 5375 2880 5380 2900
rect 5350 2850 5380 2880
rect 5350 2830 5355 2850
rect 5375 2830 5380 2850
rect 5350 2820 5380 2830
rect 5405 2900 5435 2910
rect 5405 2880 5410 2900
rect 5430 2880 5435 2900
rect 5405 2850 5435 2880
rect 5405 2830 5410 2850
rect 5430 2830 5435 2850
rect 5405 2820 5435 2830
rect 5470 2905 5490 2990
rect 5245 2800 5265 2820
rect 5355 2800 5375 2820
rect 5225 2790 5265 2800
rect 5225 2770 5235 2790
rect 5255 2770 5265 2790
rect 5225 2760 5265 2770
rect 5290 2790 5330 2800
rect 5290 2770 5300 2790
rect 5320 2770 5330 2790
rect 5290 2760 5330 2770
rect 5355 2790 5395 2800
rect 5355 2770 5365 2790
rect 5385 2770 5395 2790
rect 5355 2760 5395 2770
rect 5470 2740 5490 2825
rect 5130 2720 5270 2740
rect 5350 2720 5490 2740
rect 3200 2615 4040 2635
rect 4120 2615 4960 2635
rect 3300 2430 3340 2440
rect 3300 2420 3310 2430
rect 3330 2420 3340 2430
rect 4340 2430 4380 2440
rect 4340 2420 4350 2430
rect 2650 2400 3280 2420
rect 3360 2400 3990 2420
rect 2650 2315 2670 2400
rect 2760 2370 2800 2380
rect 2760 2350 2770 2370
rect 2790 2350 2800 2370
rect 2760 2340 2800 2350
rect 2825 2370 2855 2380
rect 2825 2350 2830 2370
rect 2850 2350 2855 2370
rect 2825 2340 2855 2350
rect 2945 2370 2975 2380
rect 2945 2350 2950 2370
rect 2970 2350 2975 2370
rect 2945 2340 2975 2350
rect 3065 2370 3095 2380
rect 3065 2350 3070 2370
rect 3090 2350 3095 2370
rect 3065 2340 3095 2350
rect 3120 2370 3160 2380
rect 3120 2350 3130 2370
rect 3150 2350 3160 2370
rect 3120 2340 3160 2350
rect 3185 2370 3215 2380
rect 3185 2350 3190 2370
rect 3210 2350 3215 2370
rect 3185 2340 3215 2350
rect 3305 2370 3335 2380
rect 3305 2350 3310 2370
rect 3330 2350 3335 2370
rect 3305 2340 3335 2350
rect 3425 2370 3455 2380
rect 3425 2350 3430 2370
rect 3450 2350 3455 2370
rect 3425 2340 3455 2350
rect 3480 2370 3520 2380
rect 3480 2350 3490 2370
rect 3510 2350 3520 2370
rect 3480 2340 3520 2350
rect 3545 2370 3575 2380
rect 3545 2350 3550 2370
rect 3570 2350 3575 2370
rect 3545 2340 3575 2350
rect 3665 2370 3695 2380
rect 3665 2350 3670 2370
rect 3690 2350 3695 2370
rect 3665 2340 3695 2350
rect 3785 2370 3815 2380
rect 3785 2350 3790 2370
rect 3810 2350 3815 2370
rect 3785 2340 3815 2350
rect 3840 2370 3880 2380
rect 3840 2350 3850 2370
rect 3870 2350 3880 2370
rect 3840 2340 3880 2350
rect 2770 2320 2790 2340
rect 2830 2320 2850 2340
rect 2950 2320 2970 2340
rect 3070 2320 3090 2340
rect 3130 2320 3150 2340
rect 3190 2320 3210 2340
rect 3310 2320 3330 2340
rect 3430 2320 3450 2340
rect 3490 2320 3510 2340
rect 3550 2320 3570 2340
rect 3670 2320 3690 2340
rect 3790 2320 3810 2340
rect 3850 2320 3870 2340
rect 2650 2150 2670 2235
rect 2705 2310 2735 2320
rect 2705 2290 2710 2310
rect 2730 2290 2735 2310
rect 2705 2260 2735 2290
rect 2705 2240 2710 2260
rect 2730 2240 2735 2260
rect 2705 2200 2735 2240
rect 2765 2310 2795 2320
rect 2765 2290 2770 2310
rect 2790 2290 2795 2310
rect 2765 2260 2795 2290
rect 2765 2240 2770 2260
rect 2790 2240 2795 2260
rect 2765 2230 2795 2240
rect 2825 2310 2855 2320
rect 2825 2290 2830 2310
rect 2850 2290 2855 2310
rect 2825 2260 2855 2290
rect 2825 2240 2830 2260
rect 2850 2240 2855 2260
rect 2825 2230 2855 2240
rect 2885 2310 2915 2320
rect 2885 2290 2890 2310
rect 2910 2290 2915 2310
rect 2885 2260 2915 2290
rect 2885 2240 2890 2260
rect 2910 2240 2915 2260
rect 2885 2230 2915 2240
rect 2945 2310 2975 2320
rect 2945 2290 2950 2310
rect 2970 2290 2975 2310
rect 2945 2260 2975 2290
rect 2945 2240 2950 2260
rect 2970 2240 2975 2260
rect 2945 2230 2975 2240
rect 3005 2310 3035 2320
rect 3005 2290 3010 2310
rect 3030 2290 3035 2310
rect 3005 2260 3035 2290
rect 3005 2240 3010 2260
rect 3030 2240 3035 2260
rect 3005 2230 3035 2240
rect 3065 2310 3095 2320
rect 3065 2290 3070 2310
rect 3090 2290 3095 2310
rect 3065 2260 3095 2290
rect 3065 2240 3070 2260
rect 3090 2240 3095 2260
rect 3065 2230 3095 2240
rect 3125 2310 3155 2320
rect 3125 2290 3130 2310
rect 3150 2290 3155 2310
rect 3125 2260 3155 2290
rect 3125 2240 3130 2260
rect 3150 2240 3155 2260
rect 3125 2230 3155 2240
rect 3185 2310 3215 2320
rect 3185 2290 3190 2310
rect 3210 2290 3215 2310
rect 3185 2260 3215 2290
rect 3185 2240 3190 2260
rect 3210 2240 3215 2260
rect 3185 2230 3215 2240
rect 3245 2310 3275 2320
rect 3245 2290 3250 2310
rect 3270 2290 3275 2310
rect 3245 2260 3275 2290
rect 3245 2240 3250 2260
rect 3270 2240 3275 2260
rect 3245 2230 3275 2240
rect 3305 2310 3335 2320
rect 3305 2290 3310 2310
rect 3330 2290 3335 2310
rect 3305 2260 3335 2290
rect 3305 2240 3310 2260
rect 3330 2240 3335 2260
rect 3305 2230 3335 2240
rect 3365 2310 3395 2320
rect 3365 2290 3370 2310
rect 3390 2290 3395 2310
rect 3365 2260 3395 2290
rect 3365 2240 3370 2260
rect 3390 2240 3395 2260
rect 3365 2230 3395 2240
rect 3425 2310 3455 2320
rect 3425 2290 3430 2310
rect 3450 2290 3455 2310
rect 3425 2260 3455 2290
rect 3425 2240 3430 2260
rect 3450 2240 3455 2260
rect 3425 2230 3455 2240
rect 3485 2310 3515 2320
rect 3485 2290 3490 2310
rect 3510 2290 3515 2310
rect 3485 2260 3515 2290
rect 3485 2240 3490 2260
rect 3510 2240 3515 2260
rect 3485 2230 3515 2240
rect 3545 2310 3575 2320
rect 3545 2290 3550 2310
rect 3570 2290 3575 2310
rect 3545 2260 3575 2290
rect 3545 2240 3550 2260
rect 3570 2240 3575 2260
rect 3545 2230 3575 2240
rect 3605 2310 3635 2320
rect 3605 2290 3610 2310
rect 3630 2290 3635 2310
rect 3605 2260 3635 2290
rect 3605 2240 3610 2260
rect 3630 2240 3635 2260
rect 3605 2230 3635 2240
rect 3665 2310 3695 2320
rect 3665 2290 3670 2310
rect 3690 2290 3695 2310
rect 3665 2260 3695 2290
rect 3665 2240 3670 2260
rect 3690 2240 3695 2260
rect 3665 2230 3695 2240
rect 3725 2310 3755 2320
rect 3725 2290 3730 2310
rect 3750 2290 3755 2310
rect 3725 2260 3755 2290
rect 3725 2240 3730 2260
rect 3750 2240 3755 2260
rect 3725 2230 3755 2240
rect 3785 2310 3815 2320
rect 3785 2290 3790 2310
rect 3810 2290 3815 2310
rect 3785 2260 3815 2290
rect 3785 2240 3790 2260
rect 3810 2240 3815 2260
rect 3785 2230 3815 2240
rect 3845 2310 3875 2320
rect 3845 2290 3850 2310
rect 3870 2290 3875 2310
rect 3845 2260 3875 2290
rect 3845 2240 3850 2260
rect 3870 2240 3875 2260
rect 3845 2230 3875 2240
rect 3905 2310 3935 2320
rect 3905 2290 3910 2310
rect 3930 2290 3935 2310
rect 3905 2260 3935 2290
rect 3905 2240 3910 2260
rect 3930 2240 3935 2260
rect 2890 2210 2910 2230
rect 3010 2210 3030 2230
rect 3250 2210 3270 2230
rect 3370 2210 3390 2230
rect 3610 2210 3630 2230
rect 3730 2210 3750 2230
rect 2705 2180 2710 2200
rect 2730 2180 2735 2200
rect 2705 2170 2735 2180
rect 2790 2200 2830 2210
rect 2790 2180 2800 2200
rect 2820 2180 2830 2200
rect 2790 2170 2830 2180
rect 2880 2200 2920 2210
rect 2880 2180 2890 2200
rect 2910 2180 2920 2200
rect 2880 2170 2920 2180
rect 3000 2200 3040 2210
rect 3000 2180 3010 2200
rect 3030 2180 3040 2200
rect 3000 2170 3040 2180
rect 3120 2200 3160 2210
rect 3120 2180 3130 2200
rect 3150 2180 3160 2200
rect 3120 2170 3160 2180
rect 3240 2200 3280 2210
rect 3240 2180 3250 2200
rect 3270 2180 3280 2200
rect 3240 2170 3280 2180
rect 3360 2200 3400 2210
rect 3360 2180 3370 2200
rect 3390 2180 3400 2200
rect 3360 2170 3400 2180
rect 3480 2200 3520 2210
rect 3480 2180 3490 2200
rect 3510 2180 3520 2200
rect 3480 2170 3520 2180
rect 3600 2200 3640 2210
rect 3600 2180 3610 2200
rect 3630 2180 3640 2200
rect 3600 2170 3640 2180
rect 3720 2200 3760 2210
rect 3720 2180 3730 2200
rect 3750 2180 3760 2200
rect 3720 2170 3760 2180
rect 3815 2200 3845 2210
rect 3815 2180 3820 2200
rect 3840 2180 3845 2200
rect 3815 2170 3845 2180
rect 3905 2200 3935 2240
rect 3905 2180 3910 2200
rect 3930 2180 3935 2200
rect 3905 2170 3935 2180
rect 3970 2315 3990 2400
rect 2710 2150 2730 2170
rect 3910 2150 3930 2170
rect 3970 2150 3990 2235
rect 2650 2130 3280 2150
rect 3360 2130 3990 2150
rect 4170 2410 4350 2420
rect 4370 2420 4380 2430
rect 4460 2430 4500 2440
rect 4460 2420 4470 2430
rect 4370 2410 4470 2420
rect 4490 2420 4500 2430
rect 4580 2430 4620 2440
rect 4580 2420 4590 2430
rect 4490 2410 4590 2420
rect 4610 2420 4620 2430
rect 4700 2430 4740 2440
rect 4700 2420 4710 2430
rect 4610 2410 4710 2420
rect 4730 2420 4740 2430
rect 4820 2430 4860 2440
rect 4820 2420 4830 2430
rect 4850 2420 4860 2430
rect 4940 2430 4980 2440
rect 4940 2420 4950 2430
rect 4730 2410 4800 2420
rect 4880 2410 4950 2420
rect 4970 2420 4980 2430
rect 5060 2430 5100 2440
rect 5060 2420 5070 2430
rect 4970 2410 5070 2420
rect 5090 2420 5100 2430
rect 5180 2430 5220 2440
rect 5180 2420 5190 2430
rect 5090 2410 5190 2420
rect 5210 2420 5220 2430
rect 5300 2430 5340 2440
rect 5300 2420 5310 2430
rect 5210 2410 5310 2420
rect 5330 2420 5340 2430
rect 5330 2410 5510 2420
rect 4170 2400 4800 2410
rect 4880 2400 5510 2410
rect 4170 2315 4190 2400
rect 4280 2370 4320 2380
rect 4280 2350 4290 2370
rect 4310 2350 4320 2370
rect 4280 2340 4320 2350
rect 4345 2370 4375 2380
rect 4345 2350 4350 2370
rect 4370 2350 4375 2370
rect 4345 2340 4375 2350
rect 4465 2370 4495 2380
rect 4465 2350 4470 2370
rect 4490 2350 4495 2370
rect 4465 2340 4495 2350
rect 4585 2370 4615 2380
rect 4585 2350 4590 2370
rect 4610 2350 4615 2370
rect 4585 2340 4615 2350
rect 4640 2370 4680 2380
rect 4640 2350 4650 2370
rect 4670 2350 4680 2370
rect 4640 2340 4680 2350
rect 4705 2370 4735 2380
rect 4705 2350 4710 2370
rect 4730 2350 4735 2370
rect 4705 2340 4735 2350
rect 4825 2370 4855 2380
rect 4825 2350 4830 2370
rect 4850 2350 4855 2370
rect 4825 2340 4855 2350
rect 4945 2370 4975 2380
rect 4945 2350 4950 2370
rect 4970 2350 4975 2370
rect 4945 2340 4975 2350
rect 5000 2370 5040 2380
rect 5000 2350 5010 2370
rect 5030 2350 5040 2370
rect 5000 2340 5040 2350
rect 5065 2370 5095 2380
rect 5065 2350 5070 2370
rect 5090 2350 5095 2370
rect 5065 2340 5095 2350
rect 5185 2370 5215 2380
rect 5185 2350 5190 2370
rect 5210 2350 5215 2370
rect 5185 2340 5215 2350
rect 5305 2370 5335 2380
rect 5305 2350 5310 2370
rect 5330 2350 5335 2370
rect 5305 2340 5335 2350
rect 5360 2370 5400 2380
rect 5360 2350 5370 2370
rect 5390 2350 5400 2370
rect 5360 2340 5400 2350
rect 4290 2320 4310 2340
rect 4350 2320 4370 2340
rect 4470 2320 4490 2340
rect 4590 2320 4610 2340
rect 4650 2320 4670 2340
rect 4710 2320 4730 2340
rect 4830 2320 4850 2340
rect 4950 2320 4970 2340
rect 5010 2320 5030 2340
rect 5070 2320 5090 2340
rect 5190 2320 5210 2340
rect 5310 2320 5330 2340
rect 5370 2320 5390 2340
rect 4170 2150 4190 2235
rect 4225 2310 4255 2320
rect 4225 2290 4230 2310
rect 4250 2290 4255 2310
rect 4225 2260 4255 2290
rect 4225 2240 4230 2260
rect 4250 2240 4255 2260
rect 4225 2200 4255 2240
rect 4285 2310 4315 2320
rect 4285 2290 4290 2310
rect 4310 2290 4315 2310
rect 4285 2260 4315 2290
rect 4285 2240 4290 2260
rect 4310 2240 4315 2260
rect 4285 2230 4315 2240
rect 4345 2310 4375 2320
rect 4345 2290 4350 2310
rect 4370 2290 4375 2310
rect 4345 2260 4375 2290
rect 4345 2240 4350 2260
rect 4370 2240 4375 2260
rect 4345 2230 4375 2240
rect 4405 2310 4435 2320
rect 4405 2290 4410 2310
rect 4430 2290 4435 2310
rect 4405 2260 4435 2290
rect 4405 2240 4410 2260
rect 4430 2240 4435 2260
rect 4405 2230 4435 2240
rect 4465 2310 4495 2320
rect 4465 2290 4470 2310
rect 4490 2290 4495 2310
rect 4465 2260 4495 2290
rect 4465 2240 4470 2260
rect 4490 2240 4495 2260
rect 4465 2230 4495 2240
rect 4525 2310 4555 2320
rect 4525 2290 4530 2310
rect 4550 2290 4555 2310
rect 4525 2260 4555 2290
rect 4525 2240 4530 2260
rect 4550 2240 4555 2260
rect 4525 2230 4555 2240
rect 4585 2310 4615 2320
rect 4585 2290 4590 2310
rect 4610 2290 4615 2310
rect 4585 2260 4615 2290
rect 4585 2240 4590 2260
rect 4610 2240 4615 2260
rect 4585 2230 4615 2240
rect 4645 2310 4675 2320
rect 4645 2290 4650 2310
rect 4670 2290 4675 2310
rect 4645 2260 4675 2290
rect 4645 2240 4650 2260
rect 4670 2240 4675 2260
rect 4645 2230 4675 2240
rect 4705 2310 4735 2320
rect 4705 2290 4710 2310
rect 4730 2290 4735 2310
rect 4705 2260 4735 2290
rect 4705 2240 4710 2260
rect 4730 2240 4735 2260
rect 4705 2230 4735 2240
rect 4765 2310 4795 2320
rect 4765 2290 4770 2310
rect 4790 2290 4795 2310
rect 4765 2260 4795 2290
rect 4765 2240 4770 2260
rect 4790 2240 4795 2260
rect 4765 2230 4795 2240
rect 4825 2310 4855 2320
rect 4825 2290 4830 2310
rect 4850 2290 4855 2310
rect 4825 2260 4855 2290
rect 4825 2240 4830 2260
rect 4850 2240 4855 2260
rect 4825 2230 4855 2240
rect 4885 2310 4915 2320
rect 4885 2290 4890 2310
rect 4910 2290 4915 2310
rect 4885 2260 4915 2290
rect 4885 2240 4890 2260
rect 4910 2240 4915 2260
rect 4885 2230 4915 2240
rect 4945 2310 4975 2320
rect 4945 2290 4950 2310
rect 4970 2290 4975 2310
rect 4945 2260 4975 2290
rect 4945 2240 4950 2260
rect 4970 2240 4975 2260
rect 4945 2230 4975 2240
rect 5005 2310 5035 2320
rect 5005 2290 5010 2310
rect 5030 2290 5035 2310
rect 5005 2260 5035 2290
rect 5005 2240 5010 2260
rect 5030 2240 5035 2260
rect 5005 2230 5035 2240
rect 5065 2310 5095 2320
rect 5065 2290 5070 2310
rect 5090 2290 5095 2310
rect 5065 2260 5095 2290
rect 5065 2240 5070 2260
rect 5090 2240 5095 2260
rect 5065 2230 5095 2240
rect 5125 2310 5155 2320
rect 5125 2290 5130 2310
rect 5150 2290 5155 2310
rect 5125 2260 5155 2290
rect 5125 2240 5130 2260
rect 5150 2240 5155 2260
rect 5125 2230 5155 2240
rect 5185 2310 5215 2320
rect 5185 2290 5190 2310
rect 5210 2290 5215 2310
rect 5185 2260 5215 2290
rect 5185 2240 5190 2260
rect 5210 2240 5215 2260
rect 5185 2230 5215 2240
rect 5245 2310 5275 2320
rect 5245 2290 5250 2310
rect 5270 2290 5275 2310
rect 5245 2260 5275 2290
rect 5245 2240 5250 2260
rect 5270 2240 5275 2260
rect 5245 2230 5275 2240
rect 5305 2310 5335 2320
rect 5305 2290 5310 2310
rect 5330 2290 5335 2310
rect 5305 2260 5335 2290
rect 5305 2240 5310 2260
rect 5330 2240 5335 2260
rect 5305 2230 5335 2240
rect 5365 2310 5395 2320
rect 5365 2290 5370 2310
rect 5390 2290 5395 2310
rect 5365 2260 5395 2290
rect 5365 2240 5370 2260
rect 5390 2240 5395 2260
rect 5365 2230 5395 2240
rect 5425 2310 5455 2320
rect 5425 2290 5430 2310
rect 5450 2290 5455 2310
rect 5425 2260 5455 2290
rect 5425 2240 5430 2260
rect 5450 2240 5455 2260
rect 4410 2210 4430 2230
rect 4530 2210 4550 2230
rect 4770 2210 4790 2230
rect 4890 2210 4910 2230
rect 5130 2210 5150 2230
rect 5250 2210 5270 2230
rect 4225 2180 4230 2200
rect 4250 2180 4255 2200
rect 4225 2170 4255 2180
rect 4315 2200 4345 2210
rect 4315 2180 4320 2200
rect 4340 2180 4345 2200
rect 4315 2170 4345 2180
rect 4400 2200 4440 2210
rect 4400 2180 4410 2200
rect 4430 2180 4440 2200
rect 4400 2170 4440 2180
rect 4520 2200 4560 2210
rect 4520 2180 4530 2200
rect 4550 2180 4560 2200
rect 4520 2170 4560 2180
rect 4640 2200 4680 2210
rect 4640 2180 4650 2200
rect 4670 2180 4680 2200
rect 4640 2170 4680 2180
rect 4760 2200 4800 2210
rect 4760 2180 4770 2200
rect 4790 2180 4800 2200
rect 4760 2170 4800 2180
rect 4880 2200 4920 2210
rect 4880 2180 4890 2200
rect 4910 2180 4920 2200
rect 4880 2170 4920 2180
rect 5000 2200 5040 2210
rect 5000 2180 5010 2200
rect 5030 2180 5040 2200
rect 5000 2170 5040 2180
rect 5120 2200 5160 2210
rect 5120 2180 5130 2200
rect 5150 2180 5160 2200
rect 5120 2170 5160 2180
rect 5240 2200 5280 2210
rect 5240 2180 5250 2200
rect 5270 2180 5280 2200
rect 5240 2170 5280 2180
rect 5330 2200 5370 2210
rect 5330 2180 5340 2200
rect 5360 2180 5370 2200
rect 5330 2170 5370 2180
rect 5425 2200 5455 2240
rect 5425 2180 5430 2200
rect 5450 2180 5455 2200
rect 5425 2170 5455 2180
rect 5490 2315 5510 2400
rect 4230 2150 4250 2170
rect 5430 2150 5450 2170
rect 5490 2150 5510 2235
rect 4170 2130 4800 2150
rect 4880 2130 5510 2150
rect 125 2015 2135 2055
rect -45 1715 130 1725
rect -45 1695 -35 1715
rect -15 1695 15 1715
rect 35 1695 65 1715
rect 85 1695 130 1715
rect -45 1685 130 1695
rect 650 1375 775 2015
rect 1330 1375 1455 2015
rect 2010 1375 2135 2015
rect 3080 2070 3410 2090
rect 3490 2070 3820 2090
rect 3080 1965 3100 2070
rect 3190 2040 3230 2050
rect 3190 2020 3200 2040
rect 3220 2020 3230 2040
rect 3190 2010 3230 2020
rect 3130 1995 3170 2005
rect 3130 1975 3140 1995
rect 3160 1975 3170 1995
rect 3130 1965 3170 1975
rect 3255 1995 3285 2005
rect 3255 1975 3260 1995
rect 3280 1975 3285 1995
rect 3255 1965 3285 1975
rect 3370 1995 3410 2005
rect 3370 1975 3380 1995
rect 3400 1975 3410 1995
rect 3370 1965 3410 1975
rect 3495 1995 3525 2005
rect 3495 1975 3500 1995
rect 3520 1975 3525 1995
rect 3495 1965 3525 1975
rect 3610 1995 3650 2005
rect 3610 1975 3620 1995
rect 3640 1975 3650 1995
rect 3610 1965 3650 1975
rect 3735 1995 3765 2005
rect 3735 1975 3740 1995
rect 3760 1975 3765 1995
rect 3735 1965 3765 1975
rect 3800 1965 3820 2070
rect 3140 1945 3160 1965
rect 3260 1945 3280 1965
rect 3380 1945 3400 1965
rect 3500 1945 3520 1965
rect 3620 1945 3640 1965
rect 3740 1945 3760 1965
rect 3135 1935 3165 1945
rect 3135 1915 3140 1935
rect 3160 1915 3165 1935
rect 3135 1905 3165 1915
rect 3195 1935 3225 1945
rect 3195 1915 3200 1935
rect 3220 1915 3225 1935
rect 3195 1905 3225 1915
rect 3255 1935 3285 1945
rect 3255 1915 3260 1935
rect 3280 1915 3285 1935
rect 3255 1905 3285 1915
rect 3315 1935 3345 1945
rect 3315 1915 3320 1935
rect 3340 1915 3345 1935
rect 3315 1905 3345 1915
rect 3375 1935 3405 1945
rect 3375 1915 3380 1935
rect 3400 1915 3405 1935
rect 3375 1905 3405 1915
rect 3435 1935 3465 1945
rect 3435 1915 3440 1935
rect 3460 1915 3465 1935
rect 3435 1905 3465 1915
rect 3495 1935 3525 1945
rect 3495 1915 3500 1935
rect 3520 1915 3525 1935
rect 3495 1905 3525 1915
rect 3555 1935 3585 1945
rect 3555 1915 3560 1935
rect 3580 1915 3585 1935
rect 3555 1905 3585 1915
rect 3615 1935 3645 1945
rect 3615 1915 3620 1935
rect 3640 1915 3645 1935
rect 3615 1905 3645 1915
rect 3675 1935 3705 1945
rect 3675 1915 3680 1935
rect 3700 1915 3705 1935
rect 3675 1905 3705 1915
rect 3735 1935 3765 1945
rect 3735 1915 3740 1935
rect 3760 1915 3765 1935
rect 3735 1905 3765 1915
rect 3790 1905 3800 1945
rect 4340 2070 4670 2090
rect 4750 2070 5080 2090
rect 4340 1965 4360 2070
rect 4930 2040 4970 2050
rect 4930 2020 4940 2040
rect 4960 2020 4970 2040
rect 4930 2010 4970 2020
rect 4395 1995 4425 2005
rect 4395 1975 4400 1995
rect 4420 1975 4425 1995
rect 4395 1965 4425 1975
rect 4510 1995 4550 2005
rect 4510 1975 4520 1995
rect 4540 1975 4550 1995
rect 4510 1965 4550 1975
rect 4635 1995 4665 2005
rect 4635 1975 4640 1995
rect 4660 1975 4665 1995
rect 4635 1965 4665 1975
rect 4750 1995 4790 2005
rect 4750 1975 4760 1995
rect 4780 1975 4790 1995
rect 4750 1965 4790 1975
rect 4875 1995 4905 2005
rect 4875 1975 4880 1995
rect 4900 1975 4905 1995
rect 4875 1965 4905 1975
rect 4990 1995 5030 2005
rect 4990 1975 5000 1995
rect 5020 1975 5030 1995
rect 4990 1965 5030 1975
rect 5060 1965 5080 2070
rect 3200 1885 3220 1905
rect 3320 1885 3340 1905
rect 3440 1885 3460 1905
rect 3560 1885 3580 1905
rect 3680 1885 3700 1905
rect 3820 1905 3830 1945
rect 4330 1905 4340 1945
rect 4400 1945 4420 1965
rect 4520 1945 4540 1965
rect 4640 1945 4660 1965
rect 4760 1945 4780 1965
rect 4880 1945 4900 1965
rect 5000 1945 5020 1965
rect 3080 1825 3100 1885
rect 3130 1875 3170 1885
rect 3130 1855 3140 1875
rect 3160 1855 3170 1875
rect 3130 1845 3170 1855
rect 3195 1875 3225 1885
rect 3195 1855 3200 1875
rect 3220 1855 3225 1875
rect 3195 1845 3225 1855
rect 3315 1875 3345 1885
rect 3315 1855 3320 1875
rect 3340 1855 3345 1875
rect 3315 1845 3345 1855
rect 3435 1875 3465 1885
rect 3435 1855 3440 1875
rect 3460 1855 3465 1875
rect 3435 1845 3465 1855
rect 3555 1875 3585 1885
rect 3555 1855 3560 1875
rect 3580 1855 3585 1875
rect 3555 1845 3585 1855
rect 3675 1875 3705 1885
rect 3675 1855 3680 1875
rect 3700 1855 3705 1875
rect 3675 1845 3705 1855
rect 3800 1825 3820 1885
rect 3080 1805 3410 1825
rect 3490 1805 3820 1825
rect 4360 1905 4370 1945
rect 4395 1935 4425 1945
rect 4395 1915 4400 1935
rect 4420 1915 4425 1935
rect 4395 1905 4425 1915
rect 4455 1935 4485 1945
rect 4455 1915 4460 1935
rect 4480 1915 4485 1935
rect 4455 1905 4485 1915
rect 4515 1935 4545 1945
rect 4515 1915 4520 1935
rect 4540 1915 4545 1935
rect 4515 1905 4545 1915
rect 4575 1935 4605 1945
rect 4575 1915 4580 1935
rect 4600 1915 4605 1935
rect 4575 1905 4605 1915
rect 4635 1935 4665 1945
rect 4635 1915 4640 1935
rect 4660 1915 4665 1935
rect 4635 1905 4665 1915
rect 4695 1935 4725 1945
rect 4695 1915 4700 1935
rect 4720 1915 4725 1935
rect 4695 1905 4725 1915
rect 4755 1935 4785 1945
rect 4755 1915 4760 1935
rect 4780 1915 4785 1935
rect 4755 1905 4785 1915
rect 4815 1935 4845 1945
rect 4815 1915 4820 1935
rect 4840 1915 4845 1935
rect 4815 1905 4845 1915
rect 4875 1935 4905 1945
rect 4875 1915 4880 1935
rect 4900 1915 4905 1935
rect 4875 1905 4905 1915
rect 4935 1935 4965 1945
rect 4935 1915 4940 1935
rect 4960 1915 4965 1935
rect 4935 1905 4965 1915
rect 4995 1935 5025 1945
rect 4995 1915 5000 1935
rect 5020 1915 5025 1935
rect 4995 1905 5025 1915
rect 4460 1885 4480 1905
rect 4580 1885 4600 1905
rect 4700 1885 4720 1905
rect 4820 1885 4840 1905
rect 4940 1885 4960 1905
rect 4340 1825 4360 1885
rect 4455 1875 4485 1885
rect 4455 1855 4460 1875
rect 4480 1855 4485 1875
rect 4455 1845 4485 1855
rect 4575 1875 4605 1885
rect 4575 1855 4580 1875
rect 4600 1855 4605 1875
rect 4575 1845 4605 1855
rect 4695 1875 4725 1885
rect 4695 1855 4700 1875
rect 4720 1855 4725 1875
rect 4695 1845 4725 1855
rect 4815 1875 4845 1885
rect 4815 1855 4820 1875
rect 4840 1855 4845 1875
rect 4815 1845 4845 1855
rect 4935 1875 4965 1885
rect 4935 1855 4940 1875
rect 4960 1855 4965 1875
rect 4935 1845 4965 1855
rect 4990 1875 5030 1885
rect 4990 1855 5000 1875
rect 5020 1855 5030 1875
rect 4990 1845 5030 1855
rect 5060 1825 5080 1885
rect 4340 1805 5080 1825
rect 4930 1785 4970 1805
rect 125 1335 2135 1375
rect 650 690 775 1335
rect 1330 690 1455 1335
rect 2010 695 2135 1335
rect 2840 1745 3410 1765
rect 3490 1745 4060 1765
rect 2840 1590 2860 1745
rect 2980 1715 3020 1725
rect 2890 1700 2930 1710
rect 2890 1680 2900 1700
rect 2920 1680 2930 1700
rect 2980 1695 2990 1715
rect 3010 1695 3020 1715
rect 2980 1685 3020 1695
rect 3100 1715 3140 1725
rect 3100 1695 3110 1715
rect 3130 1695 3140 1715
rect 3100 1685 3140 1695
rect 3220 1715 3260 1725
rect 3220 1695 3230 1715
rect 3250 1695 3260 1715
rect 3220 1685 3260 1695
rect 3340 1715 3380 1725
rect 3340 1695 3350 1715
rect 3370 1695 3380 1715
rect 3340 1685 3380 1695
rect 3580 1715 3620 1725
rect 3580 1695 3590 1715
rect 3610 1695 3620 1715
rect 3580 1685 3620 1695
rect 3700 1715 3740 1725
rect 3700 1695 3710 1715
rect 3730 1695 3740 1715
rect 3700 1685 3740 1695
rect 3820 1715 3860 1725
rect 3820 1695 3830 1715
rect 3850 1695 3860 1715
rect 3820 1685 3860 1695
rect 3970 1700 4010 1710
rect 2890 1670 2930 1680
rect 3970 1680 3980 1700
rect 4000 1680 4010 1700
rect 3970 1670 4010 1680
rect 2840 1350 2860 1510
rect 2895 1660 2925 1670
rect 2895 1640 2900 1660
rect 2920 1640 2925 1660
rect 2895 1610 2925 1640
rect 2895 1590 2900 1610
rect 2920 1590 2925 1610
rect 2895 1560 2925 1590
rect 2895 1540 2900 1560
rect 2920 1540 2925 1560
rect 2895 1510 2925 1540
rect 2895 1490 2900 1510
rect 2920 1490 2925 1510
rect 2895 1460 2925 1490
rect 2895 1440 2900 1460
rect 2920 1440 2925 1460
rect 2895 1430 2925 1440
rect 3435 1660 3465 1670
rect 3435 1640 3440 1660
rect 3460 1640 3465 1660
rect 3435 1610 3465 1640
rect 3435 1590 3440 1610
rect 3460 1590 3465 1610
rect 3435 1560 3465 1590
rect 3435 1540 3440 1560
rect 3460 1540 3465 1560
rect 3435 1510 3465 1540
rect 3435 1490 3440 1510
rect 3460 1490 3465 1510
rect 3435 1460 3465 1490
rect 3435 1440 3440 1460
rect 3460 1440 3465 1460
rect 3435 1430 3465 1440
rect 3975 1660 4005 1670
rect 3975 1640 3980 1660
rect 4000 1640 4005 1660
rect 3975 1610 4005 1640
rect 3975 1590 3980 1610
rect 4000 1590 4005 1610
rect 3975 1560 4005 1590
rect 3975 1540 3980 1560
rect 4000 1540 4005 1560
rect 3975 1510 4005 1540
rect 3975 1490 3980 1510
rect 4000 1490 4005 1510
rect 3975 1460 4005 1490
rect 3975 1440 3980 1460
rect 4000 1440 4005 1460
rect 3975 1430 4005 1440
rect 4040 1590 4060 1745
rect 3440 1410 3460 1430
rect 3430 1400 3470 1410
rect 3430 1380 3440 1400
rect 3460 1380 3470 1400
rect 3430 1370 3470 1380
rect 3440 1350 3460 1370
rect 4040 1350 4060 1510
rect 2840 1330 3410 1350
rect 3490 1330 4060 1350
rect 4100 1745 4670 1765
rect 4750 1745 5320 1765
rect 4100 1590 4120 1745
rect 4300 1715 4340 1725
rect 4150 1700 4190 1710
rect 4150 1680 4160 1700
rect 4180 1680 4190 1700
rect 4300 1695 4310 1715
rect 4330 1695 4340 1715
rect 4300 1685 4340 1695
rect 4420 1715 4460 1725
rect 4420 1695 4430 1715
rect 4450 1695 4460 1715
rect 4420 1685 4460 1695
rect 4540 1715 4580 1725
rect 4540 1695 4550 1715
rect 4570 1695 4580 1715
rect 4540 1685 4580 1695
rect 4780 1715 4820 1725
rect 4780 1695 4790 1715
rect 4810 1695 4820 1715
rect 4780 1685 4820 1695
rect 4900 1715 4940 1725
rect 4900 1695 4910 1715
rect 4930 1695 4940 1715
rect 4900 1685 4940 1695
rect 5020 1715 5060 1725
rect 5020 1695 5030 1715
rect 5050 1695 5060 1715
rect 5020 1685 5060 1695
rect 5140 1715 5180 1725
rect 5140 1695 5150 1715
rect 5170 1695 5180 1715
rect 5140 1685 5180 1695
rect 5230 1700 5270 1710
rect 4150 1670 4190 1680
rect 5230 1680 5240 1700
rect 5260 1680 5270 1700
rect 5230 1670 5270 1680
rect 4100 1350 4120 1510
rect 4155 1660 4185 1670
rect 4155 1640 4160 1660
rect 4180 1640 4185 1660
rect 4155 1610 4185 1640
rect 4155 1590 4160 1610
rect 4180 1590 4185 1610
rect 4155 1560 4185 1590
rect 4155 1540 4160 1560
rect 4180 1540 4185 1560
rect 4155 1510 4185 1540
rect 4155 1490 4160 1510
rect 4180 1490 4185 1510
rect 4155 1460 4185 1490
rect 4155 1440 4160 1460
rect 4180 1440 4185 1460
rect 4155 1430 4185 1440
rect 4695 1660 4725 1670
rect 4695 1640 4700 1660
rect 4720 1640 4725 1660
rect 4695 1610 4725 1640
rect 4695 1590 4700 1610
rect 4720 1590 4725 1610
rect 4695 1560 4725 1590
rect 4695 1540 4700 1560
rect 4720 1540 4725 1560
rect 4695 1510 4725 1540
rect 4695 1490 4700 1510
rect 4720 1490 4725 1510
rect 4695 1460 4725 1490
rect 4695 1440 4700 1460
rect 4720 1440 4725 1460
rect 4695 1430 4725 1440
rect 5235 1660 5265 1670
rect 5235 1640 5240 1660
rect 5260 1640 5265 1660
rect 5235 1610 5265 1640
rect 5235 1590 5240 1610
rect 5260 1590 5265 1610
rect 5235 1560 5265 1590
rect 5235 1540 5240 1560
rect 5260 1540 5265 1560
rect 5235 1510 5265 1540
rect 5235 1490 5240 1510
rect 5260 1490 5265 1510
rect 5235 1460 5265 1490
rect 5235 1440 5240 1460
rect 5260 1440 5265 1460
rect 5235 1430 5265 1440
rect 5300 1590 5320 1745
rect 4700 1410 4720 1430
rect 4690 1400 4730 1410
rect 4690 1380 4700 1400
rect 4720 1380 4730 1400
rect 4690 1370 4730 1380
rect 4700 1350 4720 1370
rect 5300 1350 5320 1510
rect 4100 1330 4670 1350
rect 4750 1330 5320 1350
rect 2940 1280 4040 1300
rect 4120 1280 5215 1300
rect 2940 1195 2960 1280
rect 3020 1250 3060 1260
rect 3020 1230 3030 1250
rect 3050 1230 3060 1250
rect 3020 1220 3060 1230
rect 3100 1250 3140 1260
rect 3100 1230 3110 1250
rect 3130 1230 3140 1250
rect 3100 1220 3140 1230
rect 3180 1250 3220 1260
rect 3180 1230 3190 1250
rect 3210 1230 3220 1250
rect 3180 1220 3220 1230
rect 3260 1250 3300 1260
rect 3260 1230 3270 1250
rect 3290 1230 3300 1250
rect 3260 1220 3300 1230
rect 3340 1250 3380 1260
rect 3340 1230 3350 1250
rect 3370 1230 3380 1250
rect 3340 1220 3380 1230
rect 3420 1250 3460 1260
rect 3420 1230 3430 1250
rect 3450 1230 3460 1250
rect 3420 1220 3460 1230
rect 3500 1250 3540 1260
rect 3500 1230 3510 1250
rect 3530 1230 3540 1250
rect 3500 1220 3540 1230
rect 3580 1250 3620 1260
rect 3580 1230 3590 1250
rect 3610 1230 3620 1250
rect 3580 1220 3620 1230
rect 3660 1250 3700 1260
rect 3660 1230 3670 1250
rect 3690 1230 3700 1250
rect 3660 1220 3700 1230
rect 3740 1250 3780 1260
rect 3740 1230 3750 1250
rect 3770 1230 3780 1250
rect 3740 1220 3780 1230
rect 3820 1250 3860 1260
rect 3820 1230 3830 1250
rect 3850 1230 3860 1250
rect 3820 1220 3860 1230
rect 3900 1250 3940 1260
rect 3900 1230 3910 1250
rect 3930 1230 3940 1250
rect 3900 1220 3940 1230
rect 3980 1250 4020 1260
rect 3980 1230 3990 1250
rect 4010 1230 4020 1250
rect 3980 1220 4020 1230
rect 4060 1250 4100 1260
rect 4060 1230 4070 1250
rect 4090 1230 4100 1250
rect 4060 1220 4100 1230
rect 4140 1250 4180 1260
rect 4140 1230 4150 1250
rect 4170 1230 4180 1250
rect 4140 1220 4180 1230
rect 4220 1250 4260 1260
rect 4220 1230 4230 1250
rect 4250 1230 4260 1250
rect 4220 1220 4260 1230
rect 4300 1250 4340 1260
rect 4300 1230 4310 1250
rect 4330 1230 4340 1250
rect 4300 1220 4340 1230
rect 4380 1250 4420 1260
rect 4380 1230 4390 1250
rect 4410 1230 4420 1250
rect 4380 1220 4420 1230
rect 4460 1250 4500 1260
rect 4460 1230 4470 1250
rect 4490 1230 4500 1250
rect 4460 1220 4500 1230
rect 4540 1250 4580 1260
rect 4540 1230 4550 1250
rect 4570 1230 4580 1250
rect 4540 1220 4580 1230
rect 4620 1250 4660 1260
rect 4620 1230 4630 1250
rect 4650 1230 4660 1250
rect 4620 1220 4660 1230
rect 4700 1250 4740 1260
rect 4700 1230 4710 1250
rect 4730 1230 4740 1250
rect 4700 1220 4740 1230
rect 4780 1250 4820 1260
rect 4780 1230 4790 1250
rect 4810 1230 4820 1250
rect 4780 1220 4820 1230
rect 4860 1250 4900 1260
rect 4860 1230 4870 1250
rect 4890 1230 4900 1250
rect 4860 1220 4900 1230
rect 4940 1250 4980 1260
rect 4940 1230 4950 1250
rect 4970 1230 4980 1250
rect 4940 1220 4980 1230
rect 5020 1250 5060 1260
rect 5020 1230 5030 1250
rect 5050 1230 5060 1250
rect 5020 1220 5060 1230
rect 3030 1200 3050 1220
rect 4070 1200 4090 1220
rect 3025 1190 3055 1200
rect 3025 1175 3030 1190
rect 2980 1170 3030 1175
rect 3050 1170 3055 1190
rect 2980 1165 3055 1170
rect 2980 1145 2990 1165
rect 3010 1145 3055 1165
rect 2980 1140 3055 1145
rect 2980 1135 3030 1140
rect 2940 1075 2960 1115
rect 3025 1120 3030 1135
rect 3050 1120 3055 1140
rect 3025 1110 3055 1120
rect 4065 1190 4095 1200
rect 4065 1170 4070 1190
rect 4090 1170 4095 1190
rect 4065 1140 4095 1170
rect 4065 1120 4070 1140
rect 4090 1120 4095 1140
rect 4065 1110 4095 1120
rect 5105 1190 5135 1200
rect 5105 1170 5110 1190
rect 5130 1175 5135 1190
rect 5195 1195 5215 1280
rect 5130 1170 5175 1175
rect 5105 1165 5175 1170
rect 5105 1145 5145 1165
rect 5165 1145 5175 1165
rect 5105 1140 5175 1145
rect 5105 1120 5110 1140
rect 5130 1135 5175 1140
rect 5130 1120 5135 1135
rect 5105 1110 5135 1120
rect 5195 1075 5215 1115
rect 2940 1055 4040 1075
rect 4120 1055 5215 1075
rect 3065 1005 3345 1025
rect 3425 1005 3700 1025
rect 3065 920 3085 1005
rect 3225 975 3265 985
rect 3225 955 3235 975
rect 3255 955 3265 975
rect 3225 945 3265 955
rect 3335 975 3375 985
rect 3335 955 3345 975
rect 3365 955 3375 975
rect 3335 945 3375 955
rect 3395 975 3425 985
rect 3395 955 3400 975
rect 3420 955 3425 975
rect 3395 945 3425 955
rect 3445 975 3485 985
rect 3445 955 3455 975
rect 3475 955 3485 975
rect 3445 945 3485 955
rect 3235 925 3255 945
rect 3345 925 3365 945
rect 3455 925 3475 945
rect 3065 755 3085 840
rect 3120 915 3150 925
rect 3120 895 3125 915
rect 3145 895 3150 915
rect 3120 865 3150 895
rect 3120 845 3125 865
rect 3145 845 3150 865
rect 3120 805 3150 845
rect 3175 915 3205 925
rect 3175 895 3180 915
rect 3200 895 3205 915
rect 3175 865 3205 895
rect 3175 845 3180 865
rect 3200 845 3205 865
rect 3175 835 3205 845
rect 3230 915 3260 925
rect 3230 895 3235 915
rect 3255 895 3260 915
rect 3230 865 3260 895
rect 3230 845 3235 865
rect 3255 845 3260 865
rect 3230 835 3260 845
rect 3285 915 3315 925
rect 3285 895 3290 915
rect 3310 895 3315 915
rect 3285 865 3315 895
rect 3285 845 3290 865
rect 3310 845 3315 865
rect 3285 835 3315 845
rect 3340 915 3370 925
rect 3340 895 3345 915
rect 3365 895 3370 915
rect 3340 865 3370 895
rect 3340 845 3345 865
rect 3365 845 3370 865
rect 3340 835 3370 845
rect 3395 915 3425 925
rect 3395 895 3400 915
rect 3420 895 3425 915
rect 3395 865 3425 895
rect 3395 845 3400 865
rect 3420 845 3425 865
rect 3395 835 3425 845
rect 3450 915 3480 925
rect 3450 895 3455 915
rect 3475 895 3480 915
rect 3450 865 3480 895
rect 3450 845 3455 865
rect 3475 845 3480 865
rect 3450 835 3480 845
rect 3505 915 3535 925
rect 3505 895 3510 915
rect 3530 895 3535 915
rect 3505 865 3535 895
rect 3505 845 3510 865
rect 3530 845 3535 865
rect 3505 835 3535 845
rect 3560 915 3590 925
rect 3560 895 3565 915
rect 3585 895 3590 915
rect 3560 865 3590 895
rect 3560 845 3565 865
rect 3585 845 3590 865
rect 3560 835 3590 845
rect 3615 915 3645 925
rect 3615 895 3620 915
rect 3640 895 3645 915
rect 3615 865 3645 895
rect 3615 845 3620 865
rect 3640 845 3645 865
rect 3180 815 3200 835
rect 3290 815 3310 835
rect 3400 815 3420 835
rect 3510 815 3530 835
rect 3120 785 3125 805
rect 3145 785 3150 805
rect 3120 775 3150 785
rect 3170 805 3210 815
rect 3170 785 3180 805
rect 3200 785 3210 805
rect 3170 775 3210 785
rect 3280 805 3320 815
rect 3280 785 3290 805
rect 3310 785 3320 805
rect 3280 775 3320 785
rect 3390 805 3430 815
rect 3390 785 3400 805
rect 3420 785 3430 805
rect 3390 775 3430 785
rect 3500 805 3540 815
rect 3500 785 3510 805
rect 3530 785 3540 805
rect 3500 775 3540 785
rect 3615 805 3645 845
rect 3615 785 3620 805
rect 3640 785 3645 805
rect 3615 775 3645 785
rect 3680 920 3700 1005
rect 3125 755 3145 775
rect 3620 755 3640 775
rect 3680 755 3700 840
rect 3065 735 3345 755
rect 3425 735 3700 755
rect 3735 1005 4040 1025
rect 4120 1005 4425 1025
rect 3735 920 3755 1005
rect 3895 975 3935 985
rect 3895 955 3905 975
rect 3925 955 3935 975
rect 3895 945 3935 955
rect 4005 975 4045 985
rect 4005 955 4015 975
rect 4035 955 4045 975
rect 4005 945 4045 955
rect 4065 975 4095 985
rect 4065 955 4070 975
rect 4090 955 4095 975
rect 4065 945 4095 955
rect 4115 975 4155 985
rect 4115 955 4125 975
rect 4145 955 4155 975
rect 4115 945 4155 955
rect 4225 975 4265 985
rect 4225 955 4235 975
rect 4255 955 4265 975
rect 4225 945 4265 955
rect 3905 925 3925 945
rect 4015 925 4035 945
rect 4125 925 4145 945
rect 4235 925 4255 945
rect 3735 755 3755 840
rect 3790 915 3820 925
rect 3790 895 3795 915
rect 3815 895 3820 915
rect 3790 865 3820 895
rect 3790 845 3795 865
rect 3815 845 3820 865
rect 3790 805 3820 845
rect 3845 915 3875 925
rect 3845 895 3850 915
rect 3870 895 3875 915
rect 3845 865 3875 895
rect 3845 845 3850 865
rect 3870 845 3875 865
rect 3845 835 3875 845
rect 3900 915 3930 925
rect 3900 895 3905 915
rect 3925 895 3930 915
rect 3900 865 3930 895
rect 3900 845 3905 865
rect 3925 845 3930 865
rect 3900 835 3930 845
rect 3955 915 3985 925
rect 3955 895 3960 915
rect 3980 895 3985 915
rect 3955 865 3985 895
rect 3955 845 3960 865
rect 3980 845 3985 865
rect 3955 835 3985 845
rect 4010 915 4040 925
rect 4010 895 4015 915
rect 4035 895 4040 915
rect 4010 865 4040 895
rect 4010 845 4015 865
rect 4035 845 4040 865
rect 4010 835 4040 845
rect 4065 915 4095 925
rect 4065 895 4070 915
rect 4090 895 4095 915
rect 4065 865 4095 895
rect 4065 845 4070 865
rect 4090 845 4095 865
rect 4065 835 4095 845
rect 4120 915 4150 925
rect 4120 895 4125 915
rect 4145 895 4150 915
rect 4120 865 4150 895
rect 4120 845 4125 865
rect 4145 845 4150 865
rect 4120 835 4150 845
rect 4175 915 4205 925
rect 4175 895 4180 915
rect 4200 895 4205 915
rect 4175 865 4205 895
rect 4175 845 4180 865
rect 4200 845 4205 865
rect 4175 835 4205 845
rect 4230 915 4260 925
rect 4230 895 4235 915
rect 4255 895 4260 915
rect 4230 865 4260 895
rect 4230 845 4235 865
rect 4255 845 4260 865
rect 4230 835 4260 845
rect 4285 915 4315 925
rect 4285 895 4290 915
rect 4310 895 4315 915
rect 4285 865 4315 895
rect 4285 845 4290 865
rect 4310 845 4315 865
rect 4285 835 4315 845
rect 4340 915 4370 925
rect 4340 895 4345 915
rect 4365 895 4370 915
rect 4340 865 4370 895
rect 4340 845 4345 865
rect 4365 845 4370 865
rect 3790 785 3795 805
rect 3815 785 3820 805
rect 3790 775 3820 785
rect 3850 815 3870 835
rect 3960 815 3980 835
rect 4070 815 4090 835
rect 4180 815 4200 835
rect 4290 815 4310 835
rect 3850 805 3905 815
rect 3850 785 3875 805
rect 3895 785 3905 805
rect 3850 775 3905 785
rect 3950 805 3990 815
rect 3950 785 3960 805
rect 3980 785 3990 805
rect 3950 775 3990 785
rect 4060 805 4100 815
rect 4060 785 4070 805
rect 4090 785 4100 805
rect 4060 775 4100 785
rect 4170 805 4210 815
rect 4170 785 4180 805
rect 4200 785 4210 805
rect 4170 775 4210 785
rect 4280 805 4320 815
rect 4280 785 4290 805
rect 4310 785 4320 805
rect 4280 775 4320 785
rect 4340 805 4370 845
rect 4340 785 4345 805
rect 4365 785 4370 805
rect 4340 775 4370 785
rect 4405 920 4425 1005
rect 3795 755 3815 775
rect 4345 755 4365 775
rect 4405 755 4425 840
rect 3735 735 4040 755
rect 4120 735 4425 755
rect 4460 1005 4735 1025
rect 4815 1005 5095 1025
rect 4460 920 4480 1005
rect 4675 975 4715 985
rect 4675 955 4685 975
rect 4705 955 4715 975
rect 4675 945 4715 955
rect 4735 975 4765 985
rect 4735 955 4740 975
rect 4760 955 4765 975
rect 4735 945 4765 955
rect 4785 975 4825 985
rect 4785 955 4795 975
rect 4815 955 4825 975
rect 4785 945 4825 955
rect 4895 975 4935 985
rect 4895 955 4905 975
rect 4925 955 4935 975
rect 4895 945 4935 955
rect 4685 925 4705 945
rect 4795 925 4815 945
rect 4905 925 4925 945
rect 4460 755 4480 840
rect 4515 915 4545 925
rect 4515 895 4520 915
rect 4540 895 4545 915
rect 4515 865 4545 895
rect 4515 845 4520 865
rect 4540 845 4545 865
rect 4515 805 4545 845
rect 4570 915 4600 925
rect 4570 895 4575 915
rect 4595 895 4600 915
rect 4570 865 4600 895
rect 4570 845 4575 865
rect 4595 845 4600 865
rect 4570 835 4600 845
rect 4625 915 4655 925
rect 4625 895 4630 915
rect 4650 895 4655 915
rect 4625 865 4655 895
rect 4625 845 4630 865
rect 4650 845 4655 865
rect 4625 835 4655 845
rect 4680 915 4710 925
rect 4680 895 4685 915
rect 4705 895 4710 915
rect 4680 865 4710 895
rect 4680 845 4685 865
rect 4705 845 4710 865
rect 4680 835 4710 845
rect 4735 915 4765 925
rect 4735 895 4740 915
rect 4760 895 4765 915
rect 4735 865 4765 895
rect 4735 845 4740 865
rect 4760 845 4765 865
rect 4735 835 4765 845
rect 4790 915 4820 925
rect 4790 895 4795 915
rect 4815 895 4820 915
rect 4790 865 4820 895
rect 4790 845 4795 865
rect 4815 845 4820 865
rect 4790 835 4820 845
rect 4845 915 4875 925
rect 4845 895 4850 915
rect 4870 895 4875 915
rect 4845 865 4875 895
rect 4845 845 4850 865
rect 4870 845 4875 865
rect 4845 835 4875 845
rect 4900 915 4930 925
rect 4900 895 4905 915
rect 4925 895 4930 915
rect 4900 865 4930 895
rect 4900 845 4905 865
rect 4925 845 4930 865
rect 4900 835 4930 845
rect 4955 915 4985 925
rect 4955 895 4960 915
rect 4980 895 4985 915
rect 4955 865 4985 895
rect 4955 845 4960 865
rect 4980 845 4985 865
rect 4955 835 4985 845
rect 5010 915 5040 925
rect 5010 895 5015 915
rect 5035 895 5040 915
rect 5010 865 5040 895
rect 5010 845 5015 865
rect 5035 845 5040 865
rect 4630 815 4650 835
rect 4740 815 4760 835
rect 4850 815 4870 835
rect 4960 815 4980 835
rect 4515 785 4520 805
rect 4540 785 4545 805
rect 4515 775 4545 785
rect 4620 805 4660 815
rect 4620 785 4630 805
rect 4650 785 4660 805
rect 4620 775 4660 785
rect 4730 805 4770 815
rect 4730 785 4740 805
rect 4760 785 4770 805
rect 4730 775 4770 785
rect 4840 805 4880 815
rect 4840 785 4850 805
rect 4870 785 4880 805
rect 4840 775 4880 785
rect 4950 805 4990 815
rect 4950 785 4960 805
rect 4980 785 4990 805
rect 4950 775 4990 785
rect 5010 805 5040 845
rect 5010 785 5015 805
rect 5035 785 5040 805
rect 5010 775 5040 785
rect 5075 920 5095 1005
rect 4520 755 4540 775
rect 5015 755 5035 775
rect 5075 755 5095 840
rect 4460 735 4735 755
rect 4815 735 5095 755
rect 3285 725 3315 735
rect 3505 725 3535 735
rect 4625 725 4655 735
rect 4845 725 4875 735
<< viali >>
rect 76 3560 101 3585
rect 76 3500 101 3525
rect 76 3295 101 3320
rect 76 3235 101 3260
rect 1361 3425 1386 3450
rect 1361 3365 1386 3390
rect 1195 3265 1205 3285
rect 1205 3265 1215 3285
rect 1300 3265 1310 3285
rect 1310 3265 1320 3285
rect 605 3180 625 3190
rect 605 3170 625 3180
rect 271 3030 296 3055
rect 944 3030 969 3055
rect 3045 3505 3065 3525
rect 3155 3505 3175 3525
rect 3210 3505 3230 3525
rect 3265 3505 3285 3525
rect 3320 3505 3340 3525
rect 3375 3505 3395 3525
rect 3100 3335 3120 3355
rect 3210 3335 3230 3355
rect 3320 3335 3340 3355
rect 3685 3505 3705 3525
rect 3795 3505 3815 3525
rect 3905 3505 3925 3525
rect 4015 3505 4035 3525
rect 4070 3505 4090 3525
rect 4125 3505 4145 3525
rect 4235 3505 4255 3525
rect 4345 3505 4365 3525
rect 4400 3505 4420 3525
rect 4455 3505 4475 3525
rect 3740 3335 3760 3355
rect 3850 3335 3870 3355
rect 3960 3335 3980 3355
rect 4070 3335 4090 3355
rect 4180 3335 4200 3355
rect 4290 3335 4310 3355
rect 4400 3335 4420 3355
rect 4765 3505 4785 3525
rect 4875 3505 4895 3525
rect 4930 3505 4950 3525
rect 4985 3505 5005 3525
rect 5095 3505 5115 3525
rect 4820 3335 4840 3355
rect 4930 3335 4950 3355
rect 5040 3335 5060 3355
rect 2430 3185 2455 3210
rect 2430 3125 2455 3150
rect 2835 3010 2855 3020
rect 271 2820 296 2845
rect 944 2820 969 2845
rect 1526 2920 1551 2945
rect 2225 2920 2250 2945
rect 2835 3000 2855 3010
rect 2835 2940 2855 2960
rect 2770 2770 2790 2790
rect 2835 2770 2855 2790
rect 2900 2770 2920 2790
rect 3260 3040 3280 3060
rect 3440 3040 3460 3060
rect 3620 3040 3640 3060
rect 3800 3040 3820 3060
rect 3980 3040 4000 3060
rect 4160 3040 4180 3060
rect 4340 3040 4360 3060
rect 4520 3040 4540 3060
rect 4700 3040 4720 3060
rect 4880 3040 4900 3060
rect 5300 3010 5320 3020
rect 3350 2670 3370 2690
rect 3530 2670 3550 2690
rect 3710 2670 3730 2690
rect 3890 2670 3910 2690
rect 3980 2670 4000 2690
rect 4070 2670 4090 2690
rect 4250 2670 4270 2690
rect 4430 2670 4450 2690
rect 4610 2670 4630 2690
rect 4700 2670 4720 2690
rect 4790 2670 4810 2690
rect 5300 3000 5320 3010
rect 5300 2940 5320 2960
rect 5235 2770 5255 2790
rect 5300 2770 5320 2790
rect 5365 2770 5385 2790
rect 3310 2420 3330 2430
rect 3310 2410 3330 2420
rect 2770 2350 2790 2370
rect 2830 2350 2850 2370
rect 2950 2350 2970 2370
rect 3070 2350 3090 2370
rect 3130 2350 3150 2370
rect 3190 2350 3210 2370
rect 3310 2350 3330 2370
rect 3430 2350 3450 2370
rect 3490 2350 3510 2370
rect 3550 2350 3570 2370
rect 3670 2350 3690 2370
rect 3790 2350 3810 2370
rect 3850 2350 3870 2370
rect 2800 2180 2820 2200
rect 2890 2180 2910 2200
rect 3010 2180 3030 2200
rect 3130 2180 3150 2200
rect 3250 2180 3270 2200
rect 3370 2180 3390 2200
rect 3490 2180 3510 2200
rect 3610 2180 3630 2200
rect 3730 2180 3750 2200
rect 3820 2180 3840 2200
rect 4350 2410 4370 2430
rect 4470 2410 4490 2430
rect 4590 2410 4610 2430
rect 4710 2410 4730 2430
rect 4830 2420 4850 2430
rect 4830 2410 4850 2420
rect 4950 2410 4970 2430
rect 5070 2410 5090 2430
rect 5190 2410 5210 2430
rect 5310 2410 5330 2430
rect 4290 2350 4310 2370
rect 4350 2350 4370 2370
rect 4470 2350 4490 2370
rect 4590 2350 4610 2370
rect 4650 2350 4670 2370
rect 4710 2350 4730 2370
rect 4830 2350 4850 2370
rect 4950 2350 4970 2370
rect 5010 2350 5030 2370
rect 5070 2350 5090 2370
rect 5190 2350 5210 2370
rect 5310 2350 5330 2370
rect 5370 2350 5390 2370
rect 4320 2180 4340 2200
rect 4410 2180 4430 2200
rect 4530 2180 4550 2200
rect 4650 2180 4670 2200
rect 4770 2180 4790 2200
rect 4890 2180 4910 2200
rect 5010 2180 5030 2200
rect 5130 2180 5150 2200
rect 5250 2180 5270 2200
rect 5340 2180 5360 2200
rect -35 1695 -15 1715
rect 3200 2020 3220 2040
rect 3140 1975 3160 1995
rect 3260 1975 3280 1995
rect 3380 1975 3400 1995
rect 3500 1975 3520 1995
rect 3620 1975 3640 1995
rect 3740 1975 3760 1995
rect 4940 2020 4960 2040
rect 4400 1975 4420 1995
rect 4520 1975 4540 1995
rect 4640 1975 4660 1995
rect 4760 1975 4780 1995
rect 4880 1975 4900 1995
rect 5000 1975 5020 1995
rect 3800 1915 3820 1935
rect 4340 1915 4360 1935
rect 3140 1855 3160 1875
rect 3200 1855 3220 1875
rect 3320 1855 3340 1875
rect 3440 1855 3460 1875
rect 3560 1855 3580 1875
rect 3680 1855 3700 1875
rect 4460 1855 4480 1875
rect 4580 1855 4600 1875
rect 4700 1855 4720 1875
rect 4820 1855 4840 1875
rect 4940 1855 4960 1875
rect 5000 1855 5020 1875
rect 2900 1680 2920 1700
rect 2990 1695 3010 1715
rect 3110 1695 3130 1715
rect 3230 1695 3250 1715
rect 3350 1695 3370 1715
rect 3590 1695 3610 1715
rect 3710 1695 3730 1715
rect 3830 1695 3850 1715
rect 3980 1680 4000 1700
rect 3440 1380 3460 1400
rect 4160 1680 4180 1700
rect 4310 1695 4330 1715
rect 4430 1695 4450 1715
rect 4550 1695 4570 1715
rect 4790 1695 4810 1715
rect 4910 1695 4930 1715
rect 5030 1695 5050 1715
rect 5150 1695 5170 1715
rect 5240 1680 5260 1700
rect 4700 1380 4720 1400
rect 4070 1280 4090 1300
rect 3030 1230 3050 1250
rect 3110 1230 3130 1250
rect 3190 1230 3210 1250
rect 3270 1230 3290 1250
rect 3350 1230 3370 1250
rect 3430 1230 3450 1250
rect 3510 1230 3530 1250
rect 3590 1230 3610 1250
rect 3670 1230 3690 1250
rect 3750 1230 3770 1250
rect 3830 1230 3850 1250
rect 3910 1230 3930 1250
rect 3990 1230 4010 1250
rect 4070 1230 4090 1250
rect 4150 1230 4170 1250
rect 4230 1230 4250 1250
rect 4310 1230 4330 1250
rect 4390 1230 4410 1250
rect 4470 1230 4490 1250
rect 4550 1230 4570 1250
rect 4630 1230 4650 1250
rect 4710 1230 4730 1250
rect 4790 1230 4810 1250
rect 4870 1230 4890 1250
rect 4950 1230 4970 1250
rect 5030 1230 5050 1250
rect 2990 1145 3010 1165
rect 5145 1145 5165 1165
rect 3235 955 3255 975
rect 3345 955 3365 975
rect 3400 955 3420 975
rect 3455 955 3475 975
rect 3180 785 3200 805
rect 3290 785 3310 805
rect 3400 785 3420 805
rect 3510 785 3530 805
rect 3680 870 3700 890
rect 3905 955 3925 975
rect 4015 955 4035 975
rect 4070 955 4090 975
rect 4125 955 4145 975
rect 4235 955 4255 975
rect 3735 870 3755 890
rect 3875 785 3895 805
rect 3960 785 3980 805
rect 4070 785 4090 805
rect 4180 785 4200 805
rect 4290 785 4310 805
rect 4405 870 4425 890
rect 4685 955 4705 975
rect 4740 955 4760 975
rect 4795 955 4815 975
rect 4905 955 4925 975
rect 4460 870 4480 890
rect 4630 785 4650 805
rect 4740 785 4760 805
rect 4850 785 4870 805
rect 4960 785 4980 805
rect 5075 870 5095 890
<< metal1 >>
rect 1350 3875 1390 3880
rect 1350 3845 1355 3875
rect 1385 3845 1390 3875
rect 1350 3840 1390 3845
rect 4440 3845 4480 3850
rect -15 3795 25 3800
rect -15 3765 -10 3795
rect 20 3765 25 3795
rect -15 3760 25 3765
rect 940 3795 980 3800
rect 940 3765 945 3795
rect 975 3765 980 3795
rect 940 3760 980 3765
rect -60 3740 -20 3745
rect -60 3710 -55 3740
rect -25 3710 -20 3740
rect -60 3705 -20 3710
rect -50 3060 -30 3705
rect -60 3055 -20 3060
rect -60 3025 -55 3055
rect -25 3025 -20 3055
rect -60 3020 -20 3025
rect -5 2855 15 3760
rect 1255 3690 1295 3695
rect 1255 3660 1260 3690
rect 1290 3660 1295 3690
rect 1255 3655 1295 3660
rect 70 3640 110 3645
rect 70 3610 75 3640
rect 105 3610 110 3640
rect 70 3605 110 3610
rect 75 3590 100 3605
rect 66 3555 71 3590
rect 106 3555 111 3590
rect 66 3495 71 3530
rect 106 3495 111 3530
rect 1265 3380 1285 3655
rect 1360 3455 1380 3840
rect 4440 3815 4445 3845
rect 4475 3815 4480 3845
rect 4440 3810 4480 3815
rect 1635 3795 1685 3805
rect 1635 3765 1645 3795
rect 1675 3765 1685 3795
rect 2510 3800 2550 3805
rect 2510 3770 2515 3800
rect 2545 3770 2550 3800
rect 2510 3765 2550 3770
rect 4655 3795 4695 3800
rect 4655 3765 4660 3795
rect 4690 3765 4695 3795
rect 1635 3755 1685 3765
rect 1351 3420 1356 3455
rect 1391 3420 1396 3455
rect 1361 3395 1381 3420
rect 70 3375 110 3380
rect 70 3345 75 3375
rect 105 3345 110 3375
rect 70 3340 110 3345
rect 1255 3375 1295 3380
rect 1255 3345 1260 3375
rect 1290 3345 1295 3375
rect 1351 3360 1356 3395
rect 1391 3360 1396 3395
rect 1255 3340 1295 3345
rect 75 3325 100 3340
rect 66 3290 71 3325
rect 106 3290 111 3325
rect 1185 3290 1225 3295
rect 66 3230 71 3265
rect 106 3230 111 3265
rect 1185 3260 1190 3290
rect 1220 3260 1225 3290
rect 1185 3255 1225 3260
rect 1290 3290 1330 3295
rect 1290 3260 1295 3290
rect 1325 3260 1330 3290
rect 1290 3255 1330 3260
rect 595 3195 635 3200
rect 595 3165 600 3195
rect 630 3165 635 3195
rect 2420 3180 2425 3215
rect 2460 3180 2465 3215
rect 595 3160 635 3165
rect 2420 3155 2465 3160
rect 2420 3120 2425 3155
rect 2460 3120 2465 3155
rect 2420 3115 2465 3120
rect 261 3025 266 3060
rect 301 3025 306 3060
rect 934 3025 939 3060
rect 974 3025 979 3060
rect 1210 3055 1250 3060
rect 1210 3025 1215 3055
rect 1245 3025 1250 3055
rect 1210 3020 1250 3025
rect 1105 2950 1145 2955
rect 1105 2920 1110 2950
rect 1140 2920 1145 2950
rect 1105 2915 1145 2920
rect -15 2850 25 2855
rect -15 2820 -10 2850
rect 20 2820 25 2850
rect -15 2815 25 2820
rect 261 2815 266 2850
rect 301 2815 306 2850
rect 934 2815 939 2850
rect 974 2815 979 2850
rect 1115 2550 1135 2915
rect 1220 2805 1240 3020
rect 2430 2950 2450 3115
rect 1516 2915 1521 2950
rect 1556 2915 1561 2950
rect 2215 2915 2220 2950
rect 2255 2915 2260 2950
rect 2420 2945 2460 2950
rect 2420 2915 2425 2945
rect 2455 2915 2460 2945
rect 2420 2910 2460 2915
rect 1210 2800 1250 2805
rect 1210 2770 1215 2800
rect 1245 2770 1250 2800
rect 1210 2765 1250 2770
rect 2375 2800 2415 2805
rect 2375 2770 2380 2800
rect 2410 2770 2415 2800
rect 2375 2765 2415 2770
rect 2330 2640 2370 2645
rect 2330 2610 2335 2640
rect 2365 2610 2370 2640
rect 2330 2605 2370 2610
rect 2275 2595 2315 2600
rect 2275 2565 2280 2595
rect 2310 2565 2315 2595
rect 2275 2560 2315 2565
rect 275 2200 1985 2550
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1715 -70 1720
rect -45 1720 -5 1725
rect -45 1715 -40 1720
rect -75 1695 -40 1715
rect -75 1690 -70 1695
rect -110 1685 -70 1690
rect -45 1690 -40 1695
rect -10 1690 -5 1720
rect -45 1685 -5 1690
rect 275 1190 625 2200
rect 952 1710 1302 1870
rect 952 1680 1270 1710
rect 1297 1680 1302 1710
rect 952 1520 1302 1680
rect 1635 1190 1985 2200
rect 275 840 1985 1190
rect 2285 1175 2305 2560
rect 2340 2050 2360 2605
rect 2385 2505 2405 2765
rect 2430 2700 2450 2910
rect 2465 2845 2505 2850
rect 2465 2815 2470 2845
rect 2500 2815 2505 2845
rect 2465 2810 2505 2815
rect 2420 2695 2460 2700
rect 2420 2665 2425 2695
rect 2455 2665 2460 2695
rect 2420 2660 2460 2665
rect 2375 2500 2415 2505
rect 2375 2470 2380 2500
rect 2410 2470 2415 2500
rect 2375 2465 2415 2470
rect 2330 2045 2370 2050
rect 2330 2015 2335 2045
rect 2365 2015 2370 2045
rect 2330 2010 2370 2015
rect 2340 1715 2360 2010
rect 2430 1885 2450 2660
rect 2475 2380 2495 2810
rect 2465 2375 2505 2380
rect 2465 2345 2470 2375
rect 2500 2345 2505 2375
rect 2465 2340 2505 2345
rect 2520 2150 2540 3765
rect 4655 3760 4695 3765
rect 5135 3795 5185 3805
rect 5135 3765 5145 3795
rect 5175 3765 5185 3795
rect 2690 3740 2730 3745
rect 2690 3710 2695 3740
rect 2725 3710 2730 3740
rect 2690 3705 2730 3710
rect 3385 3740 3435 3750
rect 3385 3710 3395 3740
rect 3425 3710 3435 3740
rect 3385 3700 3435 3710
rect 4610 3740 4650 3745
rect 4610 3710 4615 3740
rect 4645 3710 4650 3740
rect 4610 3705 4650 3710
rect 4390 3690 4430 3695
rect 4390 3660 4395 3690
rect 4425 3660 4430 3690
rect 4390 3655 4430 3660
rect 2555 3640 2595 3645
rect 2555 3610 2560 3640
rect 2590 3610 2595 3640
rect 2555 3605 2595 3610
rect 3310 3635 3350 3640
rect 3310 3605 3315 3635
rect 3345 3605 3350 3635
rect 2565 3260 2585 3605
rect 3310 3600 3350 3605
rect 3200 3590 3240 3595
rect 3200 3560 3205 3590
rect 3235 3560 3240 3590
rect 3200 3555 3240 3560
rect 3210 3535 3230 3555
rect 3320 3535 3340 3600
rect 4060 3590 4100 3595
rect 4060 3560 4065 3590
rect 4095 3560 4100 3590
rect 4060 3555 4100 3560
rect 4070 3535 4090 3555
rect 4400 3535 4420 3655
rect 4565 3590 4605 3595
rect 4565 3560 4570 3590
rect 4600 3560 4605 3590
rect 4565 3555 4605 3560
rect 3035 3530 3075 3535
rect 3035 3500 3040 3530
rect 3070 3500 3075 3530
rect 3035 3495 3075 3500
rect 3145 3530 3185 3535
rect 3145 3500 3150 3530
rect 3180 3500 3185 3530
rect 3145 3495 3185 3500
rect 3205 3525 3235 3535
rect 3205 3505 3210 3525
rect 3230 3505 3235 3525
rect 3205 3495 3235 3505
rect 3255 3530 3295 3535
rect 3255 3500 3260 3530
rect 3290 3500 3295 3530
rect 3255 3495 3295 3500
rect 3315 3525 3345 3535
rect 3315 3505 3320 3525
rect 3340 3505 3345 3525
rect 3315 3495 3345 3505
rect 3365 3530 3405 3535
rect 3365 3500 3370 3530
rect 3400 3500 3405 3530
rect 3365 3495 3405 3500
rect 3675 3530 3715 3535
rect 3675 3500 3680 3530
rect 3710 3500 3715 3530
rect 3675 3495 3715 3500
rect 3785 3530 3825 3535
rect 3785 3500 3790 3530
rect 3820 3500 3825 3530
rect 3785 3495 3825 3500
rect 3895 3530 3935 3535
rect 3895 3500 3900 3530
rect 3930 3500 3935 3530
rect 3895 3495 3935 3500
rect 4005 3530 4045 3535
rect 4005 3500 4010 3530
rect 4040 3500 4045 3530
rect 4005 3495 4045 3500
rect 4065 3525 4095 3535
rect 4065 3505 4070 3525
rect 4090 3505 4095 3525
rect 4065 3495 4095 3505
rect 4115 3530 4155 3535
rect 4115 3500 4120 3530
rect 4150 3500 4155 3530
rect 4115 3495 4155 3500
rect 4225 3530 4265 3535
rect 4225 3500 4230 3530
rect 4260 3500 4265 3530
rect 4225 3495 4265 3500
rect 4335 3530 4375 3535
rect 4335 3500 4340 3530
rect 4370 3500 4375 3530
rect 4335 3495 4375 3500
rect 4395 3525 4425 3535
rect 4395 3505 4400 3525
rect 4420 3505 4425 3525
rect 4395 3495 4425 3505
rect 4445 3530 4485 3535
rect 4445 3500 4450 3530
rect 4480 3500 4485 3530
rect 4445 3495 4485 3500
rect 3090 3360 3130 3365
rect 3090 3330 3095 3360
rect 3125 3330 3130 3360
rect 3090 3325 3130 3330
rect 3200 3360 3240 3365
rect 3200 3330 3205 3360
rect 3235 3330 3240 3360
rect 3200 3325 3240 3330
rect 3310 3360 3350 3365
rect 3310 3330 3315 3360
rect 3345 3330 3350 3360
rect 3310 3325 3350 3330
rect 3730 3355 3770 3365
rect 3730 3335 3740 3355
rect 3760 3335 3770 3355
rect 3730 3325 3770 3335
rect 3840 3360 3880 3365
rect 3840 3330 3845 3360
rect 3875 3330 3880 3360
rect 3840 3325 3880 3330
rect 3950 3360 3990 3365
rect 3950 3330 3955 3360
rect 3985 3330 3990 3360
rect 3950 3325 3990 3330
rect 4060 3360 4100 3365
rect 4060 3330 4065 3360
rect 4095 3330 4100 3360
rect 4060 3325 4100 3330
rect 4170 3360 4210 3365
rect 4170 3330 4175 3360
rect 4205 3330 4210 3360
rect 4170 3325 4210 3330
rect 4280 3360 4320 3365
rect 4280 3330 4285 3360
rect 4315 3330 4320 3360
rect 4280 3325 4320 3330
rect 4390 3355 4430 3365
rect 4390 3335 4400 3355
rect 4420 3335 4430 3355
rect 4390 3325 4430 3335
rect 2555 3255 2595 3260
rect 2555 3225 2560 3255
rect 2590 3225 2595 3255
rect 2555 3220 2595 3225
rect 2610 3255 2650 3260
rect 2610 3225 2615 3255
rect 2645 3225 2650 3255
rect 2610 3220 2650 3225
rect 2555 3165 2595 3170
rect 2555 3135 2560 3165
rect 2590 3135 2595 3165
rect 2555 3130 2595 3135
rect 2510 2145 2550 2150
rect 2510 2115 2515 2145
rect 2545 2115 2550 2145
rect 2510 2110 2550 2115
rect 2420 1880 2460 1885
rect 2420 1850 2425 1880
rect 2455 1850 2460 1880
rect 2420 1845 2460 1850
rect 2330 1710 2370 1715
rect 2330 1680 2335 1710
rect 2365 1680 2370 1710
rect 2330 1675 2370 1680
rect 2275 1170 2315 1175
rect 2275 1140 2280 1170
rect 2310 1140 2315 1170
rect 2275 1135 2315 1140
rect 2565 715 2585 3130
rect 2620 2555 2640 3220
rect 3060 3210 3100 3215
rect 3060 3180 3065 3210
rect 3095 3180 3100 3210
rect 3060 3175 3100 3180
rect 2825 3025 2865 3030
rect 2825 2995 2830 3025
rect 2860 2995 2865 3025
rect 2825 2990 2865 2995
rect 3070 2970 3090 3175
rect 3740 3170 3760 3325
rect 3730 3165 3770 3170
rect 3730 3135 3735 3165
rect 3765 3135 3770 3165
rect 3730 3130 3770 3135
rect 4070 3130 4090 3325
rect 4400 3165 4420 3325
rect 4575 3320 4595 3555
rect 4565 3315 4605 3320
rect 4565 3285 4570 3315
rect 4600 3285 4605 3315
rect 4565 3280 4605 3285
rect 4620 3265 4640 3705
rect 4610 3260 4650 3265
rect 4610 3230 4615 3260
rect 4645 3230 4650 3260
rect 4610 3225 4650 3230
rect 4665 3210 4685 3760
rect 5135 3755 5185 3765
rect 4920 3590 4960 3595
rect 4920 3560 4925 3590
rect 4955 3560 4960 3590
rect 4920 3555 4960 3560
rect 4930 3535 4950 3555
rect 4755 3530 4795 3535
rect 4755 3500 4760 3530
rect 4790 3500 4795 3530
rect 4755 3495 4795 3500
rect 4865 3530 4905 3535
rect 4865 3500 4870 3530
rect 4900 3500 4905 3530
rect 4865 3495 4905 3500
rect 4925 3525 4955 3535
rect 4925 3505 4930 3525
rect 4950 3505 4955 3525
rect 4925 3495 4955 3505
rect 4975 3530 5015 3535
rect 4975 3500 4980 3530
rect 5010 3500 5015 3530
rect 4975 3495 5015 3500
rect 5085 3530 5125 3535
rect 5085 3500 5090 3530
rect 5120 3500 5125 3530
rect 5085 3495 5125 3500
rect 4810 3360 4850 3365
rect 4810 3330 4815 3360
rect 4845 3330 4850 3360
rect 4810 3325 4850 3330
rect 4920 3360 4960 3365
rect 4920 3330 4925 3360
rect 4955 3330 4960 3360
rect 4920 3325 4960 3330
rect 5030 3360 5070 3365
rect 5030 3330 5035 3360
rect 5065 3330 5070 3360
rect 5030 3325 5070 3330
rect 4970 3305 5010 3310
rect 4970 3275 4975 3305
rect 5005 3275 5010 3305
rect 4970 3270 5010 3275
rect 4655 3205 4695 3210
rect 4655 3175 4660 3205
rect 4690 3175 4695 3205
rect 4655 3170 4695 3175
rect 4390 3160 4430 3165
rect 4390 3130 4395 3160
rect 4425 3130 4430 3160
rect 4060 3125 4100 3130
rect 4390 3125 4430 3130
rect 4060 3095 4065 3125
rect 4095 3095 4100 3125
rect 4060 3090 4100 3095
rect 3250 3065 3290 3070
rect 3250 3035 3255 3065
rect 3285 3035 3290 3065
rect 3250 3030 3290 3035
rect 3430 3065 3470 3070
rect 3430 3035 3435 3065
rect 3465 3035 3470 3065
rect 3430 3030 3470 3035
rect 3610 3065 3650 3070
rect 3610 3035 3615 3065
rect 3645 3035 3650 3065
rect 3610 3030 3650 3035
rect 3790 3065 3830 3070
rect 3790 3035 3795 3065
rect 3825 3035 3830 3065
rect 3790 3030 3830 3035
rect 3970 3065 4010 3070
rect 3970 3035 3975 3065
rect 4005 3035 4010 3065
rect 3970 3030 4010 3035
rect 4150 3065 4190 3070
rect 4150 3035 4155 3065
rect 4185 3035 4190 3065
rect 4150 3030 4190 3035
rect 4330 3065 4370 3070
rect 4330 3035 4335 3065
rect 4365 3035 4370 3065
rect 4330 3030 4370 3035
rect 4510 3065 4550 3070
rect 4510 3035 4515 3065
rect 4545 3035 4550 3065
rect 4510 3030 4550 3035
rect 4690 3065 4730 3070
rect 4690 3035 4695 3065
rect 4725 3035 4730 3065
rect 4690 3030 4730 3035
rect 4870 3065 4910 3070
rect 4870 3035 4875 3065
rect 4905 3035 4910 3065
rect 4870 3030 4910 3035
rect 2825 2965 2865 2970
rect 2825 2935 2830 2965
rect 2860 2935 2865 2965
rect 2825 2930 2865 2935
rect 3060 2965 3100 2970
rect 3060 2935 3065 2965
rect 3095 2935 3100 2965
rect 3060 2930 3100 2935
rect 2760 2795 2800 2800
rect 2760 2765 2765 2795
rect 2795 2765 2800 2795
rect 2760 2760 2800 2765
rect 2825 2790 2865 2800
rect 2825 2770 2835 2790
rect 2855 2770 2865 2790
rect 2825 2760 2865 2770
rect 2890 2795 2930 2800
rect 2890 2765 2895 2795
rect 2925 2765 2930 2795
rect 2890 2760 2930 2765
rect 2835 2600 2855 2760
rect 3070 2645 3090 2930
rect 3120 2795 3160 2800
rect 3120 2765 3125 2795
rect 3155 2765 3160 2795
rect 3120 2760 3160 2765
rect 3060 2640 3100 2645
rect 3060 2610 3065 2640
rect 3095 2610 3100 2640
rect 3060 2605 3100 2610
rect 2825 2595 2865 2600
rect 2825 2565 2830 2595
rect 2860 2565 2865 2595
rect 2825 2560 2865 2565
rect 2610 2550 2650 2555
rect 2610 2520 2615 2550
rect 2645 2520 2650 2550
rect 2610 2515 2650 2520
rect 2820 2435 2860 2440
rect 2820 2405 2825 2435
rect 2855 2405 2860 2435
rect 2820 2400 2860 2405
rect 2940 2435 2980 2440
rect 2940 2405 2945 2435
rect 2975 2405 2980 2435
rect 2940 2400 2980 2405
rect 3060 2435 3100 2440
rect 3060 2405 3065 2435
rect 3095 2405 3100 2435
rect 3060 2400 3100 2405
rect 2830 2380 2850 2400
rect 2950 2380 2970 2400
rect 3070 2380 3090 2400
rect 3130 2380 3150 2760
rect 3340 2690 3380 2700
rect 3340 2670 3350 2690
rect 3370 2670 3380 2690
rect 3340 2660 3380 2670
rect 3520 2690 3560 2700
rect 3520 2670 3530 2690
rect 3550 2670 3560 2690
rect 3520 2660 3560 2670
rect 3700 2690 3740 2700
rect 3700 2670 3710 2690
rect 3730 2670 3740 2690
rect 3700 2660 3740 2670
rect 3880 2695 3920 2700
rect 3880 2665 3885 2695
rect 3915 2665 3920 2695
rect 3880 2660 3920 2665
rect 3970 2690 4010 2700
rect 3970 2670 3980 2690
rect 4000 2670 4010 2690
rect 3970 2660 4010 2670
rect 4060 2690 4100 2700
rect 4060 2670 4070 2690
rect 4090 2670 4100 2690
rect 4060 2660 4100 2670
rect 4240 2695 4280 2700
rect 4240 2665 4245 2695
rect 4275 2665 4280 2695
rect 4240 2660 4280 2665
rect 4420 2690 4460 2700
rect 4420 2670 4430 2690
rect 4450 2670 4460 2690
rect 4420 2660 4460 2670
rect 4600 2690 4640 2700
rect 4600 2670 4610 2690
rect 4630 2670 4640 2690
rect 4600 2660 4640 2670
rect 4690 2690 4730 2700
rect 4690 2670 4700 2690
rect 4720 2670 4730 2690
rect 4690 2660 4730 2670
rect 4780 2690 4820 2700
rect 4780 2670 4790 2690
rect 4810 2670 4820 2690
rect 4780 2660 4820 2670
rect 3350 2555 3370 2660
rect 3530 2600 3550 2660
rect 3710 2645 3730 2660
rect 3700 2640 3740 2645
rect 3700 2610 3705 2640
rect 3735 2610 3740 2640
rect 3700 2605 3740 2610
rect 3520 2595 3560 2600
rect 3520 2565 3525 2595
rect 3555 2565 3560 2595
rect 3520 2560 3560 2565
rect 3340 2550 3380 2555
rect 3340 2520 3345 2550
rect 3375 2520 3380 2550
rect 3340 2515 3380 2520
rect 3180 2435 3220 2440
rect 3180 2405 3185 2435
rect 3215 2405 3220 2435
rect 3180 2400 3220 2405
rect 3300 2435 3340 2440
rect 3300 2405 3305 2435
rect 3335 2405 3340 2435
rect 3300 2400 3340 2405
rect 3420 2435 3460 2440
rect 3420 2405 3425 2435
rect 3455 2405 3460 2435
rect 3420 2400 3460 2405
rect 3540 2435 3580 2440
rect 3540 2405 3545 2435
rect 3575 2405 3580 2435
rect 3540 2400 3580 2405
rect 3660 2435 3700 2440
rect 3660 2405 3665 2435
rect 3695 2405 3700 2435
rect 3660 2400 3700 2405
rect 3780 2435 3820 2440
rect 3780 2405 3785 2435
rect 3815 2405 3820 2435
rect 3780 2400 3820 2405
rect 3190 2380 3210 2400
rect 3310 2380 3330 2400
rect 3430 2380 3450 2400
rect 3550 2380 3570 2400
rect 3670 2380 3690 2400
rect 3790 2380 3810 2400
rect 3980 2380 4000 2660
rect 4070 2555 4090 2660
rect 4430 2645 4450 2660
rect 4420 2640 4460 2645
rect 4420 2610 4425 2640
rect 4455 2610 4460 2640
rect 4420 2605 4460 2610
rect 4610 2600 4630 2660
rect 4700 2600 4720 2660
rect 4600 2595 4640 2600
rect 4600 2565 4605 2595
rect 4635 2565 4640 2595
rect 4600 2560 4640 2565
rect 4690 2595 4730 2600
rect 4690 2565 4695 2595
rect 4725 2565 4730 2595
rect 4690 2560 4730 2565
rect 4790 2555 4810 2660
rect 4060 2550 4100 2555
rect 4060 2520 4065 2550
rect 4095 2520 4100 2550
rect 4060 2515 4100 2520
rect 4780 2550 4820 2555
rect 4780 2520 4785 2550
rect 4815 2520 4820 2550
rect 4780 2515 4820 2520
rect 4980 2505 5000 3270
rect 5060 3260 5100 3265
rect 5060 3230 5065 3260
rect 5095 3230 5100 3260
rect 5060 3225 5100 3230
rect 5015 3205 5055 3210
rect 5015 3175 5020 3205
rect 5050 3175 5055 3205
rect 5015 3170 5055 3175
rect 5025 2600 5045 3170
rect 5070 2655 5090 3225
rect 5615 3160 5655 3165
rect 5615 3130 5620 3160
rect 5650 3130 5655 3160
rect 5615 3125 5655 3130
rect 5290 3025 5330 3040
rect 5290 2995 5295 3025
rect 5325 2995 5330 3025
rect 5290 2990 5330 2995
rect 5300 2970 5320 2990
rect 5290 2965 5330 2970
rect 5290 2935 5295 2965
rect 5325 2935 5330 2965
rect 5290 2930 5330 2935
rect 5225 2795 5265 2800
rect 5225 2765 5230 2795
rect 5260 2765 5265 2795
rect 5225 2760 5265 2765
rect 5290 2790 5330 2800
rect 5290 2770 5300 2790
rect 5320 2770 5330 2790
rect 5290 2760 5330 2770
rect 5355 2795 5395 2800
rect 5355 2765 5360 2795
rect 5390 2765 5395 2795
rect 5355 2760 5395 2765
rect 5060 2650 5100 2655
rect 5060 2620 5065 2650
rect 5095 2620 5100 2650
rect 5060 2615 5100 2620
rect 5015 2595 5055 2600
rect 5015 2565 5020 2595
rect 5050 2565 5055 2595
rect 5015 2560 5055 2565
rect 5300 2505 5320 2760
rect 5525 2650 5565 2655
rect 5525 2620 5530 2650
rect 5560 2620 5565 2650
rect 5525 2615 5565 2620
rect 4280 2500 4320 2505
rect 4280 2470 4285 2500
rect 4315 2470 4320 2500
rect 4280 2465 4320 2470
rect 4970 2500 5010 2505
rect 4970 2470 4975 2500
rect 5005 2470 5010 2500
rect 4970 2465 5010 2470
rect 5290 2500 5330 2505
rect 5290 2470 5295 2500
rect 5325 2470 5330 2500
rect 5290 2465 5330 2470
rect 4290 2380 4310 2465
rect 4340 2435 4380 2440
rect 4340 2405 4345 2435
rect 4375 2405 4380 2435
rect 4340 2400 4380 2405
rect 4460 2435 4500 2440
rect 4460 2405 4465 2435
rect 4495 2405 4500 2435
rect 4460 2400 4500 2405
rect 4580 2435 4620 2440
rect 4580 2405 4585 2435
rect 4615 2405 4620 2435
rect 4580 2400 4620 2405
rect 4700 2435 4740 2440
rect 4700 2405 4705 2435
rect 4735 2405 4740 2435
rect 4700 2400 4740 2405
rect 4820 2435 4860 2440
rect 4820 2405 4825 2435
rect 4855 2405 4860 2435
rect 4820 2400 4860 2405
rect 4940 2435 4980 2440
rect 4940 2405 4945 2435
rect 4975 2405 4980 2435
rect 4940 2400 4980 2405
rect 5060 2435 5100 2440
rect 5060 2405 5065 2435
rect 5095 2405 5100 2435
rect 5060 2400 5100 2405
rect 5180 2435 5220 2440
rect 5180 2405 5185 2435
rect 5215 2405 5220 2435
rect 5180 2400 5220 2405
rect 5300 2435 5340 2440
rect 5300 2405 5305 2435
rect 5335 2405 5340 2435
rect 5300 2400 5340 2405
rect 4350 2380 4370 2400
rect 4470 2380 4490 2400
rect 4590 2380 4610 2400
rect 4710 2380 4730 2400
rect 4830 2380 4850 2400
rect 4950 2380 4970 2400
rect 5070 2380 5090 2400
rect 5190 2380 5210 2400
rect 5310 2380 5330 2400
rect 2760 2375 2800 2380
rect 2760 2345 2765 2375
rect 2795 2345 2800 2375
rect 2760 2340 2800 2345
rect 2825 2370 2855 2380
rect 2825 2350 2830 2370
rect 2850 2350 2855 2370
rect 2825 2340 2855 2350
rect 2945 2370 2975 2380
rect 2945 2350 2950 2370
rect 2970 2350 2975 2370
rect 2945 2340 2975 2350
rect 3065 2370 3095 2380
rect 3065 2350 3070 2370
rect 3090 2350 3095 2370
rect 3065 2340 3095 2350
rect 3120 2375 3160 2380
rect 3120 2345 3125 2375
rect 3155 2345 3160 2375
rect 3120 2340 3160 2345
rect 3185 2370 3215 2380
rect 3185 2350 3190 2370
rect 3210 2350 3215 2370
rect 3185 2340 3215 2350
rect 3305 2370 3335 2380
rect 3305 2350 3310 2370
rect 3330 2350 3335 2370
rect 3305 2340 3335 2350
rect 3425 2370 3455 2380
rect 3425 2350 3430 2370
rect 3450 2350 3455 2370
rect 3425 2340 3455 2350
rect 3480 2375 3520 2380
rect 3480 2345 3485 2375
rect 3515 2345 3520 2375
rect 3480 2340 3520 2345
rect 3545 2370 3575 2380
rect 3545 2350 3550 2370
rect 3570 2350 3575 2370
rect 3545 2340 3575 2350
rect 3665 2370 3695 2380
rect 3665 2350 3670 2370
rect 3690 2350 3695 2370
rect 3665 2340 3695 2350
rect 3785 2370 3815 2380
rect 3785 2350 3790 2370
rect 3810 2350 3815 2370
rect 3785 2340 3815 2350
rect 3840 2375 3880 2380
rect 3840 2345 3845 2375
rect 3875 2345 3880 2375
rect 3840 2340 3880 2345
rect 3970 2375 4010 2380
rect 3970 2345 3975 2375
rect 4005 2345 4010 2375
rect 3970 2340 4010 2345
rect 4150 2375 4190 2380
rect 4150 2345 4155 2375
rect 4185 2345 4190 2375
rect 4150 2340 4190 2345
rect 4280 2375 4320 2380
rect 4280 2345 4285 2375
rect 4315 2345 4320 2375
rect 4280 2340 4320 2345
rect 4345 2370 4375 2380
rect 4345 2350 4350 2370
rect 4370 2350 4375 2370
rect 4345 2340 4375 2350
rect 4465 2370 4495 2380
rect 4465 2350 4470 2370
rect 4490 2350 4495 2370
rect 4465 2340 4495 2350
rect 4585 2370 4615 2380
rect 4585 2350 4590 2370
rect 4610 2350 4615 2370
rect 4585 2340 4615 2350
rect 4640 2375 4680 2380
rect 4640 2345 4645 2375
rect 4675 2345 4680 2375
rect 4640 2340 4680 2345
rect 4705 2370 4735 2380
rect 4705 2350 4710 2370
rect 4730 2350 4735 2370
rect 4705 2340 4735 2350
rect 4825 2370 4855 2380
rect 4825 2350 4830 2370
rect 4850 2350 4855 2370
rect 4825 2340 4855 2350
rect 4945 2370 4975 2380
rect 4945 2350 4950 2370
rect 4970 2350 4975 2370
rect 4945 2340 4975 2350
rect 5000 2375 5040 2380
rect 5000 2345 5005 2375
rect 5035 2345 5040 2375
rect 5000 2340 5040 2345
rect 5065 2370 5095 2380
rect 5065 2350 5070 2370
rect 5090 2350 5095 2370
rect 5065 2340 5095 2350
rect 5185 2370 5215 2380
rect 5185 2350 5190 2370
rect 5210 2350 5215 2370
rect 5185 2340 5215 2350
rect 5305 2370 5335 2380
rect 5305 2350 5310 2370
rect 5330 2350 5335 2370
rect 5305 2340 5335 2350
rect 5360 2375 5400 2380
rect 5360 2345 5365 2375
rect 5395 2345 5400 2375
rect 5360 2340 5400 2345
rect 2790 2200 2830 2210
rect 2790 2180 2800 2200
rect 2820 2180 2830 2200
rect 2790 2170 2830 2180
rect 2880 2205 2920 2210
rect 2880 2175 2885 2205
rect 2915 2175 2920 2205
rect 2880 2170 2920 2175
rect 3000 2200 3040 2210
rect 3000 2180 3010 2200
rect 3030 2180 3040 2200
rect 3000 2170 3040 2180
rect 3120 2200 3160 2210
rect 3120 2180 3130 2200
rect 3150 2180 3160 2200
rect 3120 2170 3160 2180
rect 3240 2205 3280 2210
rect 3240 2175 3245 2205
rect 3275 2175 3280 2205
rect 3240 2170 3280 2175
rect 3360 2200 3400 2210
rect 3360 2180 3370 2200
rect 3390 2180 3400 2200
rect 3360 2170 3400 2180
rect 3480 2200 3520 2210
rect 3480 2180 3490 2200
rect 3510 2180 3520 2200
rect 3480 2170 3520 2180
rect 3600 2205 3640 2210
rect 3600 2175 3605 2205
rect 3635 2175 3640 2205
rect 3600 2170 3640 2175
rect 3720 2200 3760 2210
rect 3720 2180 3730 2200
rect 3750 2180 3760 2200
rect 3720 2170 3760 2180
rect 3815 2200 3845 2210
rect 3815 2180 3820 2200
rect 3840 2180 3845 2200
rect 3815 2170 3845 2180
rect 2800 2150 2820 2170
rect 3010 2150 3030 2170
rect 3130 2150 3150 2170
rect 2790 2145 2830 2150
rect 2790 2115 2795 2145
rect 2825 2115 2830 2145
rect 2790 2110 2830 2115
rect 3000 2145 3040 2150
rect 3000 2115 3005 2145
rect 3035 2115 3040 2145
rect 3000 2110 3040 2115
rect 3120 2145 3160 2150
rect 3120 2115 3125 2145
rect 3155 2115 3160 2145
rect 3120 2110 3160 2115
rect 3260 2065 3280 2170
rect 3370 2150 3390 2170
rect 3490 2150 3510 2170
rect 3730 2150 3750 2170
rect 3820 2150 3840 2170
rect 3360 2145 3400 2150
rect 3360 2115 3365 2145
rect 3395 2115 3400 2145
rect 3360 2110 3400 2115
rect 3480 2145 3520 2150
rect 3480 2115 3485 2145
rect 3515 2115 3520 2145
rect 3480 2110 3520 2115
rect 3720 2145 3760 2150
rect 3720 2115 3725 2145
rect 3755 2115 3760 2145
rect 3720 2110 3760 2115
rect 3810 2145 3850 2150
rect 3810 2115 3815 2145
rect 3845 2115 3850 2145
rect 3810 2110 3850 2115
rect 3250 2060 3290 2065
rect 3190 2045 3230 2050
rect 3190 2015 3195 2045
rect 3225 2015 3230 2045
rect 3250 2030 3255 2060
rect 3285 2030 3290 2060
rect 3250 2025 3290 2030
rect 3190 2010 3230 2015
rect 3260 2005 3280 2025
rect 3370 2005 3390 2110
rect 3490 2060 3530 2065
rect 3490 2030 3495 2060
rect 3525 2030 3530 2060
rect 3490 2025 3530 2030
rect 3730 2060 3770 2065
rect 3730 2030 3735 2060
rect 3765 2030 3770 2060
rect 3730 2025 3770 2030
rect 3500 2005 3520 2025
rect 3740 2005 3760 2025
rect 3130 2000 3170 2005
rect 3130 1970 3135 2000
rect 3165 1970 3170 2000
rect 3130 1965 3170 1970
rect 3255 1995 3285 2005
rect 3255 1975 3260 1995
rect 3280 1975 3285 1995
rect 3255 1965 3285 1975
rect 3370 2000 3410 2005
rect 3370 1970 3375 2000
rect 3405 1970 3410 2000
rect 3370 1965 3410 1970
rect 3495 1995 3525 2005
rect 3495 1975 3500 1995
rect 3520 1975 3525 1995
rect 3495 1965 3525 1975
rect 3610 2000 3650 2005
rect 3610 1970 3615 2000
rect 3645 1970 3650 2000
rect 3610 1965 3650 1970
rect 3735 1995 3765 2005
rect 3735 1975 3740 1995
rect 3760 1975 3765 1995
rect 3735 1965 3765 1975
rect 3790 1940 3830 1945
rect 3790 1910 3795 1940
rect 3825 1910 3830 1940
rect 3790 1905 3830 1910
rect 3130 1880 3170 1885
rect 3130 1850 3135 1880
rect 3165 1850 3170 1880
rect 3130 1845 3170 1850
rect 3195 1875 3225 1885
rect 3195 1855 3200 1875
rect 3220 1855 3225 1875
rect 3195 1845 3225 1855
rect 3315 1875 3345 1885
rect 3315 1855 3320 1875
rect 3340 1855 3345 1875
rect 3315 1845 3345 1855
rect 3435 1875 3465 1885
rect 3435 1855 3440 1875
rect 3460 1855 3465 1875
rect 3435 1845 3465 1855
rect 3555 1875 3585 1885
rect 3555 1855 3560 1875
rect 3580 1855 3585 1875
rect 3555 1845 3585 1855
rect 3675 1875 3705 1885
rect 3675 1855 3680 1875
rect 3700 1855 3705 1875
rect 3675 1845 3705 1855
rect 3200 1825 3220 1845
rect 3320 1825 3340 1845
rect 3440 1825 3460 1845
rect 3560 1825 3580 1845
rect 3680 1825 3700 1845
rect 2890 1820 2930 1825
rect 2890 1790 2895 1820
rect 2925 1790 2930 1820
rect 2890 1785 2930 1790
rect 3190 1820 3230 1825
rect 3190 1790 3195 1820
rect 3225 1790 3230 1820
rect 3190 1785 3230 1790
rect 3310 1820 3350 1825
rect 3310 1790 3315 1820
rect 3345 1790 3350 1820
rect 3310 1785 3350 1790
rect 3430 1820 3470 1825
rect 3430 1790 3435 1820
rect 3465 1790 3470 1820
rect 3430 1785 3470 1790
rect 3550 1820 3590 1825
rect 3550 1790 3555 1820
rect 3585 1790 3590 1820
rect 3550 1785 3590 1790
rect 3670 1820 3710 1825
rect 3670 1790 3675 1820
rect 3705 1790 3710 1820
rect 3670 1785 3710 1790
rect 2900 1710 2920 1785
rect 2980 1720 3020 1725
rect 2890 1700 2930 1710
rect 2890 1680 2900 1700
rect 2920 1680 2930 1700
rect 2980 1690 2985 1720
rect 3015 1690 3020 1720
rect 2980 1685 3020 1690
rect 3100 1720 3140 1725
rect 3100 1690 3105 1720
rect 3135 1690 3140 1720
rect 3100 1685 3140 1690
rect 3220 1720 3260 1725
rect 3220 1690 3225 1720
rect 3255 1690 3260 1720
rect 3220 1685 3260 1690
rect 3340 1720 3380 1725
rect 3340 1690 3345 1720
rect 3375 1690 3380 1720
rect 3340 1685 3380 1690
rect 3580 1720 3620 1725
rect 3580 1690 3585 1720
rect 3615 1690 3620 1720
rect 3580 1685 3620 1690
rect 3700 1720 3740 1725
rect 3700 1690 3705 1720
rect 3735 1690 3740 1720
rect 3700 1685 3740 1690
rect 3820 1720 3860 1725
rect 3820 1690 3825 1720
rect 3855 1690 3860 1720
rect 3980 1710 4000 2340
rect 4060 1940 4100 1945
rect 4060 1910 4065 1940
rect 4095 1910 4100 1940
rect 4060 1905 4100 1910
rect 3820 1685 3860 1690
rect 3970 1700 4010 1710
rect 2890 1670 2930 1680
rect 3970 1680 3980 1700
rect 4000 1680 4010 1700
rect 3970 1670 4010 1680
rect 4070 1410 4090 1905
rect 4160 1710 4180 2340
rect 4315 2200 4345 2210
rect 4315 2180 4320 2200
rect 4340 2180 4345 2200
rect 4315 2170 4345 2180
rect 4400 2200 4440 2210
rect 4400 2180 4410 2200
rect 4430 2180 4440 2200
rect 4400 2170 4440 2180
rect 4520 2205 4560 2210
rect 4520 2175 4525 2205
rect 4555 2175 4560 2205
rect 4520 2170 4560 2175
rect 4640 2200 4680 2210
rect 4640 2180 4650 2200
rect 4670 2180 4680 2200
rect 4640 2170 4680 2180
rect 4760 2200 4800 2210
rect 4760 2180 4770 2200
rect 4790 2180 4800 2200
rect 4760 2170 4800 2180
rect 4880 2205 4920 2210
rect 4880 2175 4885 2205
rect 4915 2175 4920 2205
rect 4880 2170 4920 2175
rect 5000 2200 5040 2210
rect 5000 2180 5010 2200
rect 5030 2180 5040 2200
rect 5000 2170 5040 2180
rect 5120 2200 5160 2210
rect 5120 2180 5130 2200
rect 5150 2180 5160 2200
rect 5120 2170 5160 2180
rect 5240 2205 5280 2210
rect 5240 2175 5245 2205
rect 5275 2175 5280 2205
rect 5240 2170 5280 2175
rect 5330 2200 5370 2210
rect 5330 2180 5340 2200
rect 5360 2180 5370 2200
rect 5330 2170 5370 2180
rect 4320 2150 4340 2170
rect 4410 2150 4430 2170
rect 4650 2150 4670 2170
rect 4770 2150 4790 2170
rect 4310 2145 4350 2150
rect 4310 2115 4315 2145
rect 4345 2115 4350 2145
rect 4310 2110 4350 2115
rect 4400 2145 4440 2150
rect 4400 2115 4405 2145
rect 4435 2115 4440 2145
rect 4400 2110 4440 2115
rect 4640 2145 4680 2150
rect 4640 2115 4645 2145
rect 4675 2115 4680 2145
rect 4640 2110 4680 2115
rect 4760 2145 4800 2150
rect 4760 2115 4765 2145
rect 4795 2115 4800 2145
rect 4760 2110 4800 2115
rect 4390 2060 4430 2065
rect 4390 2030 4395 2060
rect 4425 2030 4430 2060
rect 4390 2025 4430 2030
rect 4630 2060 4670 2065
rect 4630 2030 4635 2060
rect 4665 2030 4670 2060
rect 4630 2025 4670 2030
rect 4400 2005 4420 2025
rect 4640 2005 4660 2025
rect 4760 2005 4780 2110
rect 4880 2065 4900 2170
rect 5010 2150 5030 2170
rect 5130 2150 5150 2170
rect 5340 2150 5360 2170
rect 5535 2150 5555 2615
rect 5570 2550 5610 2555
rect 5570 2520 5575 2550
rect 5605 2520 5610 2550
rect 5570 2515 5610 2520
rect 5000 2145 5040 2150
rect 5000 2115 5005 2145
rect 5035 2115 5040 2145
rect 5000 2110 5040 2115
rect 5120 2145 5160 2150
rect 5120 2115 5125 2145
rect 5155 2115 5160 2145
rect 5120 2110 5160 2115
rect 5330 2145 5370 2150
rect 5330 2115 5335 2145
rect 5365 2115 5370 2145
rect 5330 2110 5370 2115
rect 5525 2145 5565 2150
rect 5525 2115 5530 2145
rect 5560 2115 5565 2145
rect 5525 2110 5565 2115
rect 4870 2060 4910 2065
rect 4870 2030 4875 2060
rect 4905 2030 4910 2060
rect 5580 2050 5600 2515
rect 4870 2025 4910 2030
rect 4930 2045 4970 2050
rect 4880 2005 4900 2025
rect 4930 2015 4935 2045
rect 4965 2015 4970 2045
rect 4930 2010 4970 2015
rect 5570 2045 5610 2050
rect 5570 2015 5575 2045
rect 5605 2015 5610 2045
rect 5570 2010 5610 2015
rect 4395 1995 4425 2005
rect 4395 1975 4400 1995
rect 4420 1975 4425 1995
rect 4395 1965 4425 1975
rect 4510 2000 4550 2005
rect 4510 1970 4515 2000
rect 4545 1970 4550 2000
rect 4510 1965 4550 1970
rect 4635 1995 4665 2005
rect 4635 1975 4640 1995
rect 4660 1975 4665 1995
rect 4635 1965 4665 1975
rect 4750 2000 4790 2005
rect 4750 1970 4755 2000
rect 4785 1970 4790 2000
rect 4750 1965 4790 1970
rect 4875 1995 4905 2005
rect 4875 1975 4880 1995
rect 4900 1975 4905 1995
rect 4875 1965 4905 1975
rect 4990 2000 5030 2005
rect 4990 1970 4995 2000
rect 5025 1970 5030 2000
rect 4990 1965 5030 1970
rect 4330 1940 4370 1945
rect 4330 1910 4335 1940
rect 4365 1910 4370 1940
rect 4330 1905 4370 1910
rect 5625 1885 5645 3125
rect 4455 1875 4485 1885
rect 4455 1855 4460 1875
rect 4480 1855 4485 1875
rect 4455 1845 4485 1855
rect 4575 1875 4605 1885
rect 4575 1855 4580 1875
rect 4600 1855 4605 1875
rect 4575 1845 4605 1855
rect 4695 1875 4725 1885
rect 4695 1855 4700 1875
rect 4720 1855 4725 1875
rect 4695 1845 4725 1855
rect 4815 1875 4845 1885
rect 4815 1855 4820 1875
rect 4840 1855 4845 1875
rect 4815 1845 4845 1855
rect 4935 1875 4965 1885
rect 4935 1855 4940 1875
rect 4960 1855 4965 1875
rect 4935 1845 4965 1855
rect 4990 1880 5030 1885
rect 4990 1850 4995 1880
rect 5025 1850 5030 1880
rect 4990 1845 5030 1850
rect 5615 1880 5655 1885
rect 5615 1850 5620 1880
rect 5650 1850 5655 1880
rect 5615 1845 5655 1850
rect 4460 1825 4480 1845
rect 4580 1825 4600 1845
rect 4700 1825 4720 1845
rect 4820 1825 4840 1845
rect 4940 1825 4960 1845
rect 4450 1820 4490 1825
rect 4450 1790 4455 1820
rect 4485 1790 4490 1820
rect 4450 1785 4490 1790
rect 4570 1820 4610 1825
rect 4570 1790 4575 1820
rect 4605 1790 4610 1820
rect 4570 1785 4610 1790
rect 4690 1820 4730 1825
rect 4690 1790 4695 1820
rect 4725 1790 4730 1820
rect 4690 1785 4730 1790
rect 4810 1820 4850 1825
rect 4810 1790 4815 1820
rect 4845 1790 4850 1820
rect 4810 1785 4850 1790
rect 4930 1820 4970 1825
rect 4930 1790 4935 1820
rect 4965 1790 4970 1820
rect 4930 1785 4970 1790
rect 5230 1820 5270 1825
rect 5230 1790 5235 1820
rect 5265 1790 5270 1820
rect 5230 1785 5270 1790
rect 4300 1720 4340 1725
rect 4150 1700 4190 1710
rect 4150 1680 4160 1700
rect 4180 1680 4190 1700
rect 4300 1690 4305 1720
rect 4335 1690 4340 1720
rect 4300 1685 4340 1690
rect 4420 1720 4460 1725
rect 4420 1690 4425 1720
rect 4455 1690 4460 1720
rect 4420 1685 4460 1690
rect 4540 1720 4580 1725
rect 4540 1690 4545 1720
rect 4575 1690 4580 1720
rect 4540 1685 4580 1690
rect 4780 1720 4820 1725
rect 4780 1690 4785 1720
rect 4815 1690 4820 1720
rect 4780 1685 4820 1690
rect 4900 1720 4940 1725
rect 4900 1690 4905 1720
rect 4935 1690 4940 1720
rect 4900 1685 4940 1690
rect 5020 1720 5060 1725
rect 5020 1690 5025 1720
rect 5055 1690 5060 1720
rect 5020 1685 5060 1690
rect 5140 1720 5180 1725
rect 5140 1690 5145 1720
rect 5175 1690 5180 1720
rect 5240 1710 5260 1785
rect 5140 1685 5180 1690
rect 5230 1700 5270 1710
rect 4150 1670 4190 1680
rect 5230 1680 5240 1700
rect 5260 1680 5270 1700
rect 5230 1670 5270 1680
rect 3430 1405 3470 1410
rect 3430 1375 3435 1405
rect 3465 1375 3470 1405
rect 3430 1370 3470 1375
rect 4060 1405 4100 1410
rect 4060 1375 4065 1405
rect 4095 1375 4100 1405
rect 4060 1370 4100 1375
rect 4690 1405 4730 1410
rect 4690 1375 4695 1405
rect 4725 1375 4730 1405
rect 4690 1370 4730 1375
rect 4070 1315 4090 1370
rect 4060 1310 4100 1315
rect 4060 1280 4065 1310
rect 4095 1280 4100 1310
rect 4060 1275 4100 1280
rect 3020 1255 3060 1260
rect 3020 1225 3025 1255
rect 3055 1225 3060 1255
rect 3020 1220 3060 1225
rect 3100 1255 3140 1260
rect 3100 1225 3105 1255
rect 3135 1225 3140 1255
rect 3100 1220 3140 1225
rect 3180 1255 3220 1260
rect 3180 1225 3185 1255
rect 3215 1225 3220 1255
rect 3180 1220 3220 1225
rect 3260 1255 3300 1260
rect 3260 1225 3265 1255
rect 3295 1225 3300 1255
rect 3260 1220 3300 1225
rect 3340 1255 3380 1260
rect 3340 1225 3345 1255
rect 3375 1225 3380 1255
rect 3340 1220 3380 1225
rect 3420 1255 3460 1260
rect 3420 1225 3425 1255
rect 3455 1225 3460 1255
rect 3420 1220 3460 1225
rect 3500 1255 3540 1260
rect 3500 1225 3505 1255
rect 3535 1225 3540 1255
rect 3500 1220 3540 1225
rect 3580 1255 3620 1260
rect 3580 1225 3585 1255
rect 3615 1225 3620 1255
rect 3580 1220 3620 1225
rect 3660 1255 3700 1260
rect 3660 1225 3665 1255
rect 3695 1225 3700 1255
rect 3660 1220 3700 1225
rect 3740 1255 3780 1260
rect 3740 1225 3745 1255
rect 3775 1225 3780 1255
rect 3740 1220 3780 1225
rect 3820 1255 3860 1260
rect 3820 1225 3825 1255
rect 3855 1225 3860 1255
rect 3820 1220 3860 1225
rect 3900 1255 3940 1260
rect 3900 1225 3905 1255
rect 3935 1225 3940 1255
rect 3900 1220 3940 1225
rect 3980 1255 4020 1260
rect 3980 1225 3985 1255
rect 4015 1225 4020 1255
rect 3980 1220 4020 1225
rect 4060 1255 4100 1260
rect 4060 1225 4065 1255
rect 4095 1225 4100 1255
rect 4060 1220 4100 1225
rect 4140 1255 4180 1260
rect 4140 1225 4145 1255
rect 4175 1225 4180 1255
rect 4140 1220 4180 1225
rect 4220 1255 4260 1260
rect 4220 1225 4225 1255
rect 4255 1225 4260 1255
rect 4220 1220 4260 1225
rect 4300 1255 4340 1260
rect 4300 1225 4305 1255
rect 4335 1225 4340 1255
rect 4300 1220 4340 1225
rect 4380 1255 4420 1260
rect 4380 1225 4385 1255
rect 4415 1225 4420 1255
rect 4380 1220 4420 1225
rect 4460 1255 4500 1260
rect 4460 1225 4465 1255
rect 4495 1225 4500 1255
rect 4460 1220 4500 1225
rect 4540 1255 4580 1260
rect 4540 1225 4545 1255
rect 4575 1225 4580 1255
rect 4540 1220 4580 1225
rect 4620 1255 4660 1260
rect 4620 1225 4625 1255
rect 4655 1225 4660 1255
rect 4620 1220 4660 1225
rect 4700 1255 4740 1260
rect 4700 1225 4705 1255
rect 4735 1225 4740 1255
rect 4700 1220 4740 1225
rect 4780 1255 4820 1260
rect 4780 1225 4785 1255
rect 4815 1225 4820 1255
rect 4780 1220 4820 1225
rect 4860 1255 4900 1260
rect 4860 1225 4865 1255
rect 4895 1225 4900 1255
rect 4860 1220 4900 1225
rect 4940 1255 4980 1260
rect 4940 1225 4945 1255
rect 4975 1225 4980 1255
rect 4940 1220 4980 1225
rect 5020 1255 5060 1260
rect 5020 1225 5025 1255
rect 5055 1225 5060 1255
rect 5020 1220 5060 1225
rect 2980 1170 3020 1175
rect 2980 1140 2985 1170
rect 3015 1140 3020 1170
rect 2980 1135 3020 1140
rect 5135 1170 5175 1175
rect 5135 1140 5140 1170
rect 5170 1140 5175 1170
rect 5135 1135 5175 1140
rect 3390 1050 3430 1055
rect 3390 1020 3395 1050
rect 3425 1020 3430 1050
rect 3390 1015 3430 1020
rect 4060 1050 4100 1055
rect 4060 1020 4065 1050
rect 4095 1020 4100 1050
rect 4060 1015 4100 1020
rect 4730 1050 4770 1055
rect 4730 1020 4735 1050
rect 4765 1020 4770 1050
rect 4730 1015 4770 1020
rect 3400 985 3420 1015
rect 4070 985 4090 1015
rect 4740 985 4760 1015
rect 3225 980 3265 985
rect 3225 950 3230 980
rect 3260 950 3265 980
rect 3225 945 3265 950
rect 3335 980 3375 985
rect 3335 950 3340 980
rect 3370 950 3375 980
rect 3335 945 3375 950
rect 3395 975 3425 985
rect 3395 955 3400 975
rect 3420 955 3425 975
rect 3395 945 3425 955
rect 3445 980 3485 985
rect 3445 950 3450 980
rect 3480 950 3485 980
rect 3445 945 3485 950
rect 3895 980 3935 985
rect 3895 950 3900 980
rect 3930 950 3935 980
rect 3895 945 3935 950
rect 4005 980 4045 985
rect 4005 950 4010 980
rect 4040 950 4045 980
rect 4005 945 4045 950
rect 4065 975 4095 985
rect 4065 955 4070 975
rect 4090 955 4095 975
rect 4065 945 4095 955
rect 4115 980 4155 985
rect 4115 950 4120 980
rect 4150 950 4155 980
rect 4115 945 4155 950
rect 4225 980 4265 985
rect 4225 950 4230 980
rect 4260 950 4265 980
rect 4225 945 4265 950
rect 4675 980 4715 985
rect 4675 950 4680 980
rect 4710 950 4715 980
rect 4675 945 4715 950
rect 4735 975 4765 985
rect 4735 955 4740 975
rect 4760 955 4765 975
rect 4735 945 4765 955
rect 4785 980 4825 985
rect 4785 950 4790 980
rect 4820 950 4825 980
rect 4785 945 4825 950
rect 4895 980 4935 985
rect 4895 950 4900 980
rect 4930 950 4935 980
rect 4895 945 4935 950
rect 3670 895 3710 900
rect 3670 865 3675 895
rect 3705 865 3710 895
rect 3670 860 3710 865
rect 3725 895 3765 900
rect 3725 865 3730 895
rect 3760 865 3765 895
rect 3725 860 3765 865
rect 4395 895 4435 900
rect 4395 865 4400 895
rect 4430 865 4435 895
rect 4395 860 4435 865
rect 4450 895 4490 900
rect 4450 865 4455 895
rect 4485 865 4490 895
rect 4450 860 4490 865
rect 5065 895 5105 900
rect 5065 865 5070 895
rect 5100 865 5105 895
rect 5065 860 5105 865
rect 3170 810 3210 815
rect 3170 780 3175 810
rect 3205 780 3210 810
rect 3170 775 3210 780
rect 3280 805 3320 815
rect 3280 785 3290 805
rect 3310 785 3320 805
rect 3280 775 3320 785
rect 3390 810 3430 815
rect 3390 780 3395 810
rect 3425 780 3430 810
rect 3390 775 3430 780
rect 3500 805 3540 815
rect 3500 785 3510 805
rect 3530 785 3540 805
rect 3500 775 3540 785
rect 3865 805 3905 815
rect 3865 785 3875 805
rect 3895 785 3905 805
rect 3865 775 3905 785
rect 3950 805 3990 815
rect 3950 785 3960 805
rect 3980 785 3990 805
rect 3950 775 3990 785
rect 4060 810 4100 815
rect 4060 780 4065 810
rect 4095 780 4100 810
rect 4060 775 4100 780
rect 4170 810 4210 815
rect 4170 780 4175 810
rect 4205 780 4210 810
rect 4170 775 4210 780
rect 4280 810 4320 815
rect 4280 780 4285 810
rect 4315 780 4320 810
rect 4280 775 4320 780
rect 4620 805 4660 815
rect 4620 785 4630 805
rect 4650 785 4660 805
rect 4620 775 4660 785
rect 4730 810 4770 815
rect 4730 780 4735 810
rect 4765 780 4770 810
rect 4730 775 4770 780
rect 4840 805 4880 815
rect 4840 785 4850 805
rect 4870 785 4880 805
rect 4840 775 4880 785
rect 4950 810 4990 815
rect 4950 780 4955 810
rect 4985 780 4990 810
rect 4950 775 4990 780
rect 2555 710 2595 715
rect 2555 680 2560 710
rect 2590 680 2595 710
rect 2555 675 2595 680
rect 3180 350 3200 775
rect 3290 760 3310 775
rect 3510 760 3530 775
rect 3280 755 3320 760
rect 3280 725 3285 755
rect 3315 725 3320 755
rect 3280 720 3320 725
rect 3500 755 3540 760
rect 3500 725 3505 755
rect 3535 725 3540 755
rect 3500 720 3540 725
rect 3875 715 3895 775
rect 3865 710 3905 715
rect 3865 680 3870 710
rect 3900 680 3905 710
rect 3865 675 3905 680
rect 3960 350 3980 775
rect 4060 755 4100 760
rect 4060 725 4065 755
rect 4095 725 4100 755
rect 4060 720 4100 725
rect 4070 350 4090 720
rect 4180 350 4200 775
rect 4630 760 4650 775
rect 4850 760 4870 775
rect 4620 755 4660 760
rect 4620 725 4625 755
rect 4655 725 4660 755
rect 4620 720 4660 725
rect 4840 755 4880 760
rect 4840 725 4845 755
rect 4875 725 4880 755
rect 4840 720 4880 725
rect 4960 350 4980 775
<< via1 >>
rect 1355 3845 1385 3875
rect -10 3765 20 3795
rect 945 3765 975 3795
rect -55 3710 -25 3740
rect -55 3025 -25 3055
rect 1260 3660 1290 3690
rect 75 3610 105 3640
rect 71 3585 106 3590
rect 71 3560 76 3585
rect 76 3560 101 3585
rect 101 3560 106 3585
rect 71 3555 106 3560
rect 71 3525 106 3530
rect 71 3500 76 3525
rect 76 3500 101 3525
rect 101 3500 106 3525
rect 71 3495 106 3500
rect 4445 3815 4475 3845
rect 1645 3765 1675 3795
rect 2515 3770 2545 3800
rect 4660 3765 4690 3795
rect 1356 3450 1391 3455
rect 1356 3425 1361 3450
rect 1361 3425 1386 3450
rect 1386 3425 1391 3450
rect 1356 3420 1391 3425
rect 75 3345 105 3375
rect 1260 3345 1290 3375
rect 1356 3390 1391 3395
rect 1356 3365 1361 3390
rect 1361 3365 1386 3390
rect 1386 3365 1391 3390
rect 1356 3360 1391 3365
rect 71 3320 106 3325
rect 71 3295 76 3320
rect 76 3295 101 3320
rect 101 3295 106 3320
rect 71 3290 106 3295
rect 71 3260 106 3265
rect 71 3235 76 3260
rect 76 3235 101 3260
rect 101 3235 106 3260
rect 71 3230 106 3235
rect 1190 3285 1220 3290
rect 1190 3265 1195 3285
rect 1195 3265 1215 3285
rect 1215 3265 1220 3285
rect 1190 3260 1220 3265
rect 1295 3285 1325 3290
rect 1295 3265 1300 3285
rect 1300 3265 1320 3285
rect 1320 3265 1325 3285
rect 1295 3260 1325 3265
rect 600 3190 630 3195
rect 600 3170 605 3190
rect 605 3170 625 3190
rect 625 3170 630 3190
rect 600 3165 630 3170
rect 2425 3210 2460 3215
rect 2425 3185 2430 3210
rect 2430 3185 2455 3210
rect 2455 3185 2460 3210
rect 2425 3180 2460 3185
rect 2425 3150 2460 3155
rect 2425 3125 2430 3150
rect 2430 3125 2455 3150
rect 2455 3125 2460 3150
rect 2425 3120 2460 3125
rect 266 3055 301 3060
rect 266 3030 271 3055
rect 271 3030 296 3055
rect 296 3030 301 3055
rect 266 3025 301 3030
rect 939 3055 974 3060
rect 939 3030 944 3055
rect 944 3030 969 3055
rect 969 3030 974 3055
rect 939 3025 974 3030
rect 1215 3025 1245 3055
rect 1110 2920 1140 2950
rect -10 2820 20 2850
rect 266 2845 301 2850
rect 266 2820 271 2845
rect 271 2820 296 2845
rect 296 2820 301 2845
rect 266 2815 301 2820
rect 939 2845 974 2850
rect 939 2820 944 2845
rect 944 2820 969 2845
rect 969 2820 974 2845
rect 939 2815 974 2820
rect 1521 2945 1556 2950
rect 1521 2920 1526 2945
rect 1526 2920 1551 2945
rect 1551 2920 1556 2945
rect 1521 2915 1556 2920
rect 2220 2945 2255 2950
rect 2220 2920 2225 2945
rect 2225 2920 2250 2945
rect 2250 2920 2255 2945
rect 2220 2915 2255 2920
rect 2425 2915 2455 2945
rect 1215 2770 1245 2800
rect 2380 2770 2410 2800
rect 2335 2610 2365 2640
rect 2280 2565 2310 2595
rect -105 1690 -75 1720
rect -40 1715 -10 1720
rect -40 1695 -35 1715
rect -35 1695 -15 1715
rect -15 1695 -10 1715
rect -40 1690 -10 1695
rect 1270 1680 1297 1710
rect 2470 2815 2500 2845
rect 2425 2665 2455 2695
rect 2380 2470 2410 2500
rect 2335 2015 2365 2045
rect 2470 2345 2500 2375
rect 5145 3765 5175 3795
rect 2695 3710 2725 3740
rect 3395 3710 3425 3740
rect 4615 3710 4645 3740
rect 4395 3660 4425 3690
rect 2560 3610 2590 3640
rect 3315 3605 3345 3635
rect 3205 3560 3235 3590
rect 4065 3560 4095 3590
rect 4570 3560 4600 3590
rect 3040 3525 3070 3530
rect 3040 3505 3045 3525
rect 3045 3505 3065 3525
rect 3065 3505 3070 3525
rect 3040 3500 3070 3505
rect 3150 3525 3180 3530
rect 3150 3505 3155 3525
rect 3155 3505 3175 3525
rect 3175 3505 3180 3525
rect 3150 3500 3180 3505
rect 3260 3525 3290 3530
rect 3260 3505 3265 3525
rect 3265 3505 3285 3525
rect 3285 3505 3290 3525
rect 3260 3500 3290 3505
rect 3370 3525 3400 3530
rect 3370 3505 3375 3525
rect 3375 3505 3395 3525
rect 3395 3505 3400 3525
rect 3370 3500 3400 3505
rect 3680 3525 3710 3530
rect 3680 3505 3685 3525
rect 3685 3505 3705 3525
rect 3705 3505 3710 3525
rect 3680 3500 3710 3505
rect 3790 3525 3820 3530
rect 3790 3505 3795 3525
rect 3795 3505 3815 3525
rect 3815 3505 3820 3525
rect 3790 3500 3820 3505
rect 3900 3525 3930 3530
rect 3900 3505 3905 3525
rect 3905 3505 3925 3525
rect 3925 3505 3930 3525
rect 3900 3500 3930 3505
rect 4010 3525 4040 3530
rect 4010 3505 4015 3525
rect 4015 3505 4035 3525
rect 4035 3505 4040 3525
rect 4010 3500 4040 3505
rect 4120 3525 4150 3530
rect 4120 3505 4125 3525
rect 4125 3505 4145 3525
rect 4145 3505 4150 3525
rect 4120 3500 4150 3505
rect 4230 3525 4260 3530
rect 4230 3505 4235 3525
rect 4235 3505 4255 3525
rect 4255 3505 4260 3525
rect 4230 3500 4260 3505
rect 4340 3525 4370 3530
rect 4340 3505 4345 3525
rect 4345 3505 4365 3525
rect 4365 3505 4370 3525
rect 4340 3500 4370 3505
rect 4450 3525 4480 3530
rect 4450 3505 4455 3525
rect 4455 3505 4475 3525
rect 4475 3505 4480 3525
rect 4450 3500 4480 3505
rect 3095 3355 3125 3360
rect 3095 3335 3100 3355
rect 3100 3335 3120 3355
rect 3120 3335 3125 3355
rect 3095 3330 3125 3335
rect 3205 3355 3235 3360
rect 3205 3335 3210 3355
rect 3210 3335 3230 3355
rect 3230 3335 3235 3355
rect 3205 3330 3235 3335
rect 3315 3355 3345 3360
rect 3315 3335 3320 3355
rect 3320 3335 3340 3355
rect 3340 3335 3345 3355
rect 3315 3330 3345 3335
rect 3845 3355 3875 3360
rect 3845 3335 3850 3355
rect 3850 3335 3870 3355
rect 3870 3335 3875 3355
rect 3845 3330 3875 3335
rect 3955 3355 3985 3360
rect 3955 3335 3960 3355
rect 3960 3335 3980 3355
rect 3980 3335 3985 3355
rect 3955 3330 3985 3335
rect 4065 3355 4095 3360
rect 4065 3335 4070 3355
rect 4070 3335 4090 3355
rect 4090 3335 4095 3355
rect 4065 3330 4095 3335
rect 4175 3355 4205 3360
rect 4175 3335 4180 3355
rect 4180 3335 4200 3355
rect 4200 3335 4205 3355
rect 4175 3330 4205 3335
rect 4285 3355 4315 3360
rect 4285 3335 4290 3355
rect 4290 3335 4310 3355
rect 4310 3335 4315 3355
rect 4285 3330 4315 3335
rect 2560 3225 2590 3255
rect 2615 3225 2645 3255
rect 2560 3135 2590 3165
rect 2515 2115 2545 2145
rect 2425 1850 2455 1880
rect 2335 1680 2365 1710
rect 2280 1140 2310 1170
rect 3065 3180 3095 3210
rect 2830 3020 2860 3025
rect 2830 3000 2835 3020
rect 2835 3000 2855 3020
rect 2855 3000 2860 3020
rect 2830 2995 2860 3000
rect 3735 3135 3765 3165
rect 4570 3285 4600 3315
rect 4615 3230 4645 3260
rect 4925 3560 4955 3590
rect 4760 3525 4790 3530
rect 4760 3505 4765 3525
rect 4765 3505 4785 3525
rect 4785 3505 4790 3525
rect 4760 3500 4790 3505
rect 4870 3525 4900 3530
rect 4870 3505 4875 3525
rect 4875 3505 4895 3525
rect 4895 3505 4900 3525
rect 4870 3500 4900 3505
rect 4980 3525 5010 3530
rect 4980 3505 4985 3525
rect 4985 3505 5005 3525
rect 5005 3505 5010 3525
rect 4980 3500 5010 3505
rect 5090 3525 5120 3530
rect 5090 3505 5095 3525
rect 5095 3505 5115 3525
rect 5115 3505 5120 3525
rect 5090 3500 5120 3505
rect 4815 3355 4845 3360
rect 4815 3335 4820 3355
rect 4820 3335 4840 3355
rect 4840 3335 4845 3355
rect 4815 3330 4845 3335
rect 4925 3355 4955 3360
rect 4925 3335 4930 3355
rect 4930 3335 4950 3355
rect 4950 3335 4955 3355
rect 4925 3330 4955 3335
rect 5035 3355 5065 3360
rect 5035 3335 5040 3355
rect 5040 3335 5060 3355
rect 5060 3335 5065 3355
rect 5035 3330 5065 3335
rect 4975 3275 5005 3305
rect 4660 3175 4690 3205
rect 4395 3130 4425 3160
rect 4065 3095 4095 3125
rect 3255 3060 3285 3065
rect 3255 3040 3260 3060
rect 3260 3040 3280 3060
rect 3280 3040 3285 3060
rect 3255 3035 3285 3040
rect 3435 3060 3465 3065
rect 3435 3040 3440 3060
rect 3440 3040 3460 3060
rect 3460 3040 3465 3060
rect 3435 3035 3465 3040
rect 3615 3060 3645 3065
rect 3615 3040 3620 3060
rect 3620 3040 3640 3060
rect 3640 3040 3645 3060
rect 3615 3035 3645 3040
rect 3795 3060 3825 3065
rect 3795 3040 3800 3060
rect 3800 3040 3820 3060
rect 3820 3040 3825 3060
rect 3795 3035 3825 3040
rect 3975 3060 4005 3065
rect 3975 3040 3980 3060
rect 3980 3040 4000 3060
rect 4000 3040 4005 3060
rect 3975 3035 4005 3040
rect 4155 3060 4185 3065
rect 4155 3040 4160 3060
rect 4160 3040 4180 3060
rect 4180 3040 4185 3060
rect 4155 3035 4185 3040
rect 4335 3060 4365 3065
rect 4335 3040 4340 3060
rect 4340 3040 4360 3060
rect 4360 3040 4365 3060
rect 4335 3035 4365 3040
rect 4515 3060 4545 3065
rect 4515 3040 4520 3060
rect 4520 3040 4540 3060
rect 4540 3040 4545 3060
rect 4515 3035 4545 3040
rect 4695 3060 4725 3065
rect 4695 3040 4700 3060
rect 4700 3040 4720 3060
rect 4720 3040 4725 3060
rect 4695 3035 4725 3040
rect 4875 3060 4905 3065
rect 4875 3040 4880 3060
rect 4880 3040 4900 3060
rect 4900 3040 4905 3060
rect 4875 3035 4905 3040
rect 2830 2960 2860 2965
rect 2830 2940 2835 2960
rect 2835 2940 2855 2960
rect 2855 2940 2860 2960
rect 2830 2935 2860 2940
rect 3065 2935 3095 2965
rect 2765 2790 2795 2795
rect 2765 2770 2770 2790
rect 2770 2770 2790 2790
rect 2790 2770 2795 2790
rect 2765 2765 2795 2770
rect 2895 2790 2925 2795
rect 2895 2770 2900 2790
rect 2900 2770 2920 2790
rect 2920 2770 2925 2790
rect 2895 2765 2925 2770
rect 3125 2765 3155 2795
rect 3065 2610 3095 2640
rect 2830 2565 2860 2595
rect 2615 2520 2645 2550
rect 2825 2405 2855 2435
rect 2945 2405 2975 2435
rect 3065 2405 3095 2435
rect 3885 2690 3915 2695
rect 3885 2670 3890 2690
rect 3890 2670 3910 2690
rect 3910 2670 3915 2690
rect 3885 2665 3915 2670
rect 4245 2690 4275 2695
rect 4245 2670 4250 2690
rect 4250 2670 4270 2690
rect 4270 2670 4275 2690
rect 4245 2665 4275 2670
rect 3705 2610 3735 2640
rect 3525 2565 3555 2595
rect 3345 2520 3375 2550
rect 3185 2405 3215 2435
rect 3305 2430 3335 2435
rect 3305 2410 3310 2430
rect 3310 2410 3330 2430
rect 3330 2410 3335 2430
rect 3305 2405 3335 2410
rect 3425 2405 3455 2435
rect 3545 2405 3575 2435
rect 3665 2405 3695 2435
rect 3785 2405 3815 2435
rect 4425 2610 4455 2640
rect 4605 2565 4635 2595
rect 4695 2565 4725 2595
rect 4065 2520 4095 2550
rect 4785 2520 4815 2550
rect 5065 3230 5095 3260
rect 5020 3175 5050 3205
rect 5620 3130 5650 3160
rect 5295 3020 5325 3025
rect 5295 3000 5300 3020
rect 5300 3000 5320 3020
rect 5320 3000 5325 3020
rect 5295 2995 5325 3000
rect 5295 2960 5325 2965
rect 5295 2940 5300 2960
rect 5300 2940 5320 2960
rect 5320 2940 5325 2960
rect 5295 2935 5325 2940
rect 5230 2790 5260 2795
rect 5230 2770 5235 2790
rect 5235 2770 5255 2790
rect 5255 2770 5260 2790
rect 5230 2765 5260 2770
rect 5360 2790 5390 2795
rect 5360 2770 5365 2790
rect 5365 2770 5385 2790
rect 5385 2770 5390 2790
rect 5360 2765 5390 2770
rect 5065 2620 5095 2650
rect 5020 2565 5050 2595
rect 5530 2620 5560 2650
rect 4285 2470 4315 2500
rect 4975 2470 5005 2500
rect 5295 2470 5325 2500
rect 4345 2430 4375 2435
rect 4345 2410 4350 2430
rect 4350 2410 4370 2430
rect 4370 2410 4375 2430
rect 4345 2405 4375 2410
rect 4465 2430 4495 2435
rect 4465 2410 4470 2430
rect 4470 2410 4490 2430
rect 4490 2410 4495 2430
rect 4465 2405 4495 2410
rect 4585 2430 4615 2435
rect 4585 2410 4590 2430
rect 4590 2410 4610 2430
rect 4610 2410 4615 2430
rect 4585 2405 4615 2410
rect 4705 2430 4735 2435
rect 4705 2410 4710 2430
rect 4710 2410 4730 2430
rect 4730 2410 4735 2430
rect 4705 2405 4735 2410
rect 4825 2430 4855 2435
rect 4825 2410 4830 2430
rect 4830 2410 4850 2430
rect 4850 2410 4855 2430
rect 4825 2405 4855 2410
rect 4945 2430 4975 2435
rect 4945 2410 4950 2430
rect 4950 2410 4970 2430
rect 4970 2410 4975 2430
rect 4945 2405 4975 2410
rect 5065 2430 5095 2435
rect 5065 2410 5070 2430
rect 5070 2410 5090 2430
rect 5090 2410 5095 2430
rect 5065 2405 5095 2410
rect 5185 2430 5215 2435
rect 5185 2410 5190 2430
rect 5190 2410 5210 2430
rect 5210 2410 5215 2430
rect 5185 2405 5215 2410
rect 5305 2430 5335 2435
rect 5305 2410 5310 2430
rect 5310 2410 5330 2430
rect 5330 2410 5335 2430
rect 5305 2405 5335 2410
rect 2765 2370 2795 2375
rect 2765 2350 2770 2370
rect 2770 2350 2790 2370
rect 2790 2350 2795 2370
rect 2765 2345 2795 2350
rect 3125 2370 3155 2375
rect 3125 2350 3130 2370
rect 3130 2350 3150 2370
rect 3150 2350 3155 2370
rect 3125 2345 3155 2350
rect 3485 2370 3515 2375
rect 3485 2350 3490 2370
rect 3490 2350 3510 2370
rect 3510 2350 3515 2370
rect 3485 2345 3515 2350
rect 3845 2370 3875 2375
rect 3845 2350 3850 2370
rect 3850 2350 3870 2370
rect 3870 2350 3875 2370
rect 3845 2345 3875 2350
rect 3975 2345 4005 2375
rect 4155 2345 4185 2375
rect 4285 2370 4315 2375
rect 4285 2350 4290 2370
rect 4290 2350 4310 2370
rect 4310 2350 4315 2370
rect 4285 2345 4315 2350
rect 4645 2370 4675 2375
rect 4645 2350 4650 2370
rect 4650 2350 4670 2370
rect 4670 2350 4675 2370
rect 4645 2345 4675 2350
rect 5005 2370 5035 2375
rect 5005 2350 5010 2370
rect 5010 2350 5030 2370
rect 5030 2350 5035 2370
rect 5005 2345 5035 2350
rect 5365 2370 5395 2375
rect 5365 2350 5370 2370
rect 5370 2350 5390 2370
rect 5390 2350 5395 2370
rect 5365 2345 5395 2350
rect 2885 2200 2915 2205
rect 2885 2180 2890 2200
rect 2890 2180 2910 2200
rect 2910 2180 2915 2200
rect 2885 2175 2915 2180
rect 3245 2200 3275 2205
rect 3245 2180 3250 2200
rect 3250 2180 3270 2200
rect 3270 2180 3275 2200
rect 3245 2175 3275 2180
rect 3605 2200 3635 2205
rect 3605 2180 3610 2200
rect 3610 2180 3630 2200
rect 3630 2180 3635 2200
rect 3605 2175 3635 2180
rect 2795 2115 2825 2145
rect 3005 2115 3035 2145
rect 3125 2115 3155 2145
rect 3365 2115 3395 2145
rect 3485 2115 3515 2145
rect 3725 2115 3755 2145
rect 3815 2115 3845 2145
rect 3195 2040 3225 2045
rect 3195 2020 3200 2040
rect 3200 2020 3220 2040
rect 3220 2020 3225 2040
rect 3195 2015 3225 2020
rect 3255 2030 3285 2060
rect 3495 2030 3525 2060
rect 3735 2030 3765 2060
rect 3135 1995 3165 2000
rect 3135 1975 3140 1995
rect 3140 1975 3160 1995
rect 3160 1975 3165 1995
rect 3135 1970 3165 1975
rect 3375 1995 3405 2000
rect 3375 1975 3380 1995
rect 3380 1975 3400 1995
rect 3400 1975 3405 1995
rect 3375 1970 3405 1975
rect 3615 1995 3645 2000
rect 3615 1975 3620 1995
rect 3620 1975 3640 1995
rect 3640 1975 3645 1995
rect 3615 1970 3645 1975
rect 3795 1935 3825 1940
rect 3795 1915 3800 1935
rect 3800 1915 3820 1935
rect 3820 1915 3825 1935
rect 3795 1910 3825 1915
rect 3135 1875 3165 1880
rect 3135 1855 3140 1875
rect 3140 1855 3160 1875
rect 3160 1855 3165 1875
rect 3135 1850 3165 1855
rect 2895 1790 2925 1820
rect 3195 1790 3225 1820
rect 3315 1790 3345 1820
rect 3435 1790 3465 1820
rect 3555 1790 3585 1820
rect 3675 1790 3705 1820
rect 2985 1715 3015 1720
rect 2985 1695 2990 1715
rect 2990 1695 3010 1715
rect 3010 1695 3015 1715
rect 2985 1690 3015 1695
rect 3105 1715 3135 1720
rect 3105 1695 3110 1715
rect 3110 1695 3130 1715
rect 3130 1695 3135 1715
rect 3105 1690 3135 1695
rect 3225 1715 3255 1720
rect 3225 1695 3230 1715
rect 3230 1695 3250 1715
rect 3250 1695 3255 1715
rect 3225 1690 3255 1695
rect 3345 1715 3375 1720
rect 3345 1695 3350 1715
rect 3350 1695 3370 1715
rect 3370 1695 3375 1715
rect 3345 1690 3375 1695
rect 3585 1715 3615 1720
rect 3585 1695 3590 1715
rect 3590 1695 3610 1715
rect 3610 1695 3615 1715
rect 3585 1690 3615 1695
rect 3705 1715 3735 1720
rect 3705 1695 3710 1715
rect 3710 1695 3730 1715
rect 3730 1695 3735 1715
rect 3705 1690 3735 1695
rect 3825 1715 3855 1720
rect 3825 1695 3830 1715
rect 3830 1695 3850 1715
rect 3850 1695 3855 1715
rect 3825 1690 3855 1695
rect 4065 1910 4095 1940
rect 4525 2200 4555 2205
rect 4525 2180 4530 2200
rect 4530 2180 4550 2200
rect 4550 2180 4555 2200
rect 4525 2175 4555 2180
rect 4885 2200 4915 2205
rect 4885 2180 4890 2200
rect 4890 2180 4910 2200
rect 4910 2180 4915 2200
rect 4885 2175 4915 2180
rect 5245 2200 5275 2205
rect 5245 2180 5250 2200
rect 5250 2180 5270 2200
rect 5270 2180 5275 2200
rect 5245 2175 5275 2180
rect 4315 2115 4345 2145
rect 4405 2115 4435 2145
rect 4645 2115 4675 2145
rect 4765 2115 4795 2145
rect 4395 2030 4425 2060
rect 4635 2030 4665 2060
rect 5575 2520 5605 2550
rect 5005 2115 5035 2145
rect 5125 2115 5155 2145
rect 5335 2115 5365 2145
rect 5530 2115 5560 2145
rect 4875 2030 4905 2060
rect 4935 2040 4965 2045
rect 4935 2020 4940 2040
rect 4940 2020 4960 2040
rect 4960 2020 4965 2040
rect 4935 2015 4965 2020
rect 5575 2015 5605 2045
rect 4515 1995 4545 2000
rect 4515 1975 4520 1995
rect 4520 1975 4540 1995
rect 4540 1975 4545 1995
rect 4515 1970 4545 1975
rect 4755 1995 4785 2000
rect 4755 1975 4760 1995
rect 4760 1975 4780 1995
rect 4780 1975 4785 1995
rect 4755 1970 4785 1975
rect 4995 1995 5025 2000
rect 4995 1975 5000 1995
rect 5000 1975 5020 1995
rect 5020 1975 5025 1995
rect 4995 1970 5025 1975
rect 4335 1935 4365 1940
rect 4335 1915 4340 1935
rect 4340 1915 4360 1935
rect 4360 1915 4365 1935
rect 4335 1910 4365 1915
rect 4995 1875 5025 1880
rect 4995 1855 5000 1875
rect 5000 1855 5020 1875
rect 5020 1855 5025 1875
rect 4995 1850 5025 1855
rect 5620 1850 5650 1880
rect 4455 1790 4485 1820
rect 4575 1790 4605 1820
rect 4695 1790 4725 1820
rect 4815 1790 4845 1820
rect 4935 1790 4965 1820
rect 5235 1790 5265 1820
rect 4305 1715 4335 1720
rect 4305 1695 4310 1715
rect 4310 1695 4330 1715
rect 4330 1695 4335 1715
rect 4305 1690 4335 1695
rect 4425 1715 4455 1720
rect 4425 1695 4430 1715
rect 4430 1695 4450 1715
rect 4450 1695 4455 1715
rect 4425 1690 4455 1695
rect 4545 1715 4575 1720
rect 4545 1695 4550 1715
rect 4550 1695 4570 1715
rect 4570 1695 4575 1715
rect 4545 1690 4575 1695
rect 4785 1715 4815 1720
rect 4785 1695 4790 1715
rect 4790 1695 4810 1715
rect 4810 1695 4815 1715
rect 4785 1690 4815 1695
rect 4905 1715 4935 1720
rect 4905 1695 4910 1715
rect 4910 1695 4930 1715
rect 4930 1695 4935 1715
rect 4905 1690 4935 1695
rect 5025 1715 5055 1720
rect 5025 1695 5030 1715
rect 5030 1695 5050 1715
rect 5050 1695 5055 1715
rect 5025 1690 5055 1695
rect 5145 1715 5175 1720
rect 5145 1695 5150 1715
rect 5150 1695 5170 1715
rect 5170 1695 5175 1715
rect 5145 1690 5175 1695
rect 3435 1400 3465 1405
rect 3435 1380 3440 1400
rect 3440 1380 3460 1400
rect 3460 1380 3465 1400
rect 3435 1375 3465 1380
rect 4065 1375 4095 1405
rect 4695 1400 4725 1405
rect 4695 1380 4700 1400
rect 4700 1380 4720 1400
rect 4720 1380 4725 1400
rect 4695 1375 4725 1380
rect 4065 1300 4095 1310
rect 4065 1280 4070 1300
rect 4070 1280 4090 1300
rect 4090 1280 4095 1300
rect 3025 1250 3055 1255
rect 3025 1230 3030 1250
rect 3030 1230 3050 1250
rect 3050 1230 3055 1250
rect 3025 1225 3055 1230
rect 3105 1250 3135 1255
rect 3105 1230 3110 1250
rect 3110 1230 3130 1250
rect 3130 1230 3135 1250
rect 3105 1225 3135 1230
rect 3185 1250 3215 1255
rect 3185 1230 3190 1250
rect 3190 1230 3210 1250
rect 3210 1230 3215 1250
rect 3185 1225 3215 1230
rect 3265 1250 3295 1255
rect 3265 1230 3270 1250
rect 3270 1230 3290 1250
rect 3290 1230 3295 1250
rect 3265 1225 3295 1230
rect 3345 1250 3375 1255
rect 3345 1230 3350 1250
rect 3350 1230 3370 1250
rect 3370 1230 3375 1250
rect 3345 1225 3375 1230
rect 3425 1250 3455 1255
rect 3425 1230 3430 1250
rect 3430 1230 3450 1250
rect 3450 1230 3455 1250
rect 3425 1225 3455 1230
rect 3505 1250 3535 1255
rect 3505 1230 3510 1250
rect 3510 1230 3530 1250
rect 3530 1230 3535 1250
rect 3505 1225 3535 1230
rect 3585 1250 3615 1255
rect 3585 1230 3590 1250
rect 3590 1230 3610 1250
rect 3610 1230 3615 1250
rect 3585 1225 3615 1230
rect 3665 1250 3695 1255
rect 3665 1230 3670 1250
rect 3670 1230 3690 1250
rect 3690 1230 3695 1250
rect 3665 1225 3695 1230
rect 3745 1250 3775 1255
rect 3745 1230 3750 1250
rect 3750 1230 3770 1250
rect 3770 1230 3775 1250
rect 3745 1225 3775 1230
rect 3825 1250 3855 1255
rect 3825 1230 3830 1250
rect 3830 1230 3850 1250
rect 3850 1230 3855 1250
rect 3825 1225 3855 1230
rect 3905 1250 3935 1255
rect 3905 1230 3910 1250
rect 3910 1230 3930 1250
rect 3930 1230 3935 1250
rect 3905 1225 3935 1230
rect 3985 1250 4015 1255
rect 3985 1230 3990 1250
rect 3990 1230 4010 1250
rect 4010 1230 4015 1250
rect 3985 1225 4015 1230
rect 4065 1250 4095 1255
rect 4065 1230 4070 1250
rect 4070 1230 4090 1250
rect 4090 1230 4095 1250
rect 4065 1225 4095 1230
rect 4145 1250 4175 1255
rect 4145 1230 4150 1250
rect 4150 1230 4170 1250
rect 4170 1230 4175 1250
rect 4145 1225 4175 1230
rect 4225 1250 4255 1255
rect 4225 1230 4230 1250
rect 4230 1230 4250 1250
rect 4250 1230 4255 1250
rect 4225 1225 4255 1230
rect 4305 1250 4335 1255
rect 4305 1230 4310 1250
rect 4310 1230 4330 1250
rect 4330 1230 4335 1250
rect 4305 1225 4335 1230
rect 4385 1250 4415 1255
rect 4385 1230 4390 1250
rect 4390 1230 4410 1250
rect 4410 1230 4415 1250
rect 4385 1225 4415 1230
rect 4465 1250 4495 1255
rect 4465 1230 4470 1250
rect 4470 1230 4490 1250
rect 4490 1230 4495 1250
rect 4465 1225 4495 1230
rect 4545 1250 4575 1255
rect 4545 1230 4550 1250
rect 4550 1230 4570 1250
rect 4570 1230 4575 1250
rect 4545 1225 4575 1230
rect 4625 1250 4655 1255
rect 4625 1230 4630 1250
rect 4630 1230 4650 1250
rect 4650 1230 4655 1250
rect 4625 1225 4655 1230
rect 4705 1250 4735 1255
rect 4705 1230 4710 1250
rect 4710 1230 4730 1250
rect 4730 1230 4735 1250
rect 4705 1225 4735 1230
rect 4785 1250 4815 1255
rect 4785 1230 4790 1250
rect 4790 1230 4810 1250
rect 4810 1230 4815 1250
rect 4785 1225 4815 1230
rect 4865 1250 4895 1255
rect 4865 1230 4870 1250
rect 4870 1230 4890 1250
rect 4890 1230 4895 1250
rect 4865 1225 4895 1230
rect 4945 1250 4975 1255
rect 4945 1230 4950 1250
rect 4950 1230 4970 1250
rect 4970 1230 4975 1250
rect 4945 1225 4975 1230
rect 5025 1250 5055 1255
rect 5025 1230 5030 1250
rect 5030 1230 5050 1250
rect 5050 1230 5055 1250
rect 5025 1225 5055 1230
rect 2985 1165 3015 1170
rect 2985 1145 2990 1165
rect 2990 1145 3010 1165
rect 3010 1145 3015 1165
rect 2985 1140 3015 1145
rect 5140 1165 5170 1170
rect 5140 1145 5145 1165
rect 5145 1145 5165 1165
rect 5165 1145 5170 1165
rect 5140 1140 5170 1145
rect 3395 1020 3425 1050
rect 4065 1020 4095 1050
rect 4735 1020 4765 1050
rect 3230 975 3260 980
rect 3230 955 3235 975
rect 3235 955 3255 975
rect 3255 955 3260 975
rect 3230 950 3260 955
rect 3340 975 3370 980
rect 3340 955 3345 975
rect 3345 955 3365 975
rect 3365 955 3370 975
rect 3340 950 3370 955
rect 3450 975 3480 980
rect 3450 955 3455 975
rect 3455 955 3475 975
rect 3475 955 3480 975
rect 3450 950 3480 955
rect 3900 975 3930 980
rect 3900 955 3905 975
rect 3905 955 3925 975
rect 3925 955 3930 975
rect 3900 950 3930 955
rect 4010 975 4040 980
rect 4010 955 4015 975
rect 4015 955 4035 975
rect 4035 955 4040 975
rect 4010 950 4040 955
rect 4120 975 4150 980
rect 4120 955 4125 975
rect 4125 955 4145 975
rect 4145 955 4150 975
rect 4120 950 4150 955
rect 4230 975 4260 980
rect 4230 955 4235 975
rect 4235 955 4255 975
rect 4255 955 4260 975
rect 4230 950 4260 955
rect 4680 975 4710 980
rect 4680 955 4685 975
rect 4685 955 4705 975
rect 4705 955 4710 975
rect 4680 950 4710 955
rect 4790 975 4820 980
rect 4790 955 4795 975
rect 4795 955 4815 975
rect 4815 955 4820 975
rect 4790 950 4820 955
rect 4900 975 4930 980
rect 4900 955 4905 975
rect 4905 955 4925 975
rect 4925 955 4930 975
rect 4900 950 4930 955
rect 3675 890 3705 895
rect 3675 870 3680 890
rect 3680 870 3700 890
rect 3700 870 3705 890
rect 3675 865 3705 870
rect 3730 890 3760 895
rect 3730 870 3735 890
rect 3735 870 3755 890
rect 3755 870 3760 890
rect 3730 865 3760 870
rect 4400 890 4430 895
rect 4400 870 4405 890
rect 4405 870 4425 890
rect 4425 870 4430 890
rect 4400 865 4430 870
rect 4455 890 4485 895
rect 4455 870 4460 890
rect 4460 870 4480 890
rect 4480 870 4485 890
rect 4455 865 4485 870
rect 5070 890 5100 895
rect 5070 870 5075 890
rect 5075 870 5095 890
rect 5095 870 5100 890
rect 5070 865 5100 870
rect 3175 805 3205 810
rect 3175 785 3180 805
rect 3180 785 3200 805
rect 3200 785 3205 805
rect 3175 780 3205 785
rect 3395 805 3425 810
rect 3395 785 3400 805
rect 3400 785 3420 805
rect 3420 785 3425 805
rect 3395 780 3425 785
rect 4065 805 4095 810
rect 4065 785 4070 805
rect 4070 785 4090 805
rect 4090 785 4095 805
rect 4065 780 4095 785
rect 4175 805 4205 810
rect 4175 785 4180 805
rect 4180 785 4200 805
rect 4200 785 4205 805
rect 4175 780 4205 785
rect 4285 805 4315 810
rect 4285 785 4290 805
rect 4290 785 4310 805
rect 4310 785 4315 805
rect 4285 780 4315 785
rect 4735 805 4765 810
rect 4735 785 4740 805
rect 4740 785 4760 805
rect 4760 785 4765 805
rect 4735 780 4765 785
rect 4955 805 4985 810
rect 4955 785 4960 805
rect 4960 785 4980 805
rect 4980 785 4985 805
rect 4955 780 4985 785
rect 2560 680 2590 710
rect 3285 725 3315 755
rect 3505 725 3535 755
rect 3870 680 3900 710
rect 4065 725 4095 755
rect 4625 725 4655 755
rect 4845 725 4875 755
<< metal2 >>
rect -195 5340 -155 5345
rect -195 5310 -190 5340
rect -160 5310 -155 5340
rect -195 5305 -155 5310
rect 5750 5340 5790 5345
rect 5750 5310 5755 5340
rect 5785 5310 5790 5340
rect 5750 5305 5790 5310
rect -110 3875 -70 3880
rect -110 3845 -105 3875
rect -75 3870 -70 3875
rect 1350 3875 1390 3880
rect 1350 3870 1355 3875
rect -75 3850 1355 3870
rect -75 3845 -70 3850
rect -110 3840 -70 3845
rect 1350 3845 1355 3850
rect 1385 3845 1390 3875
rect 1350 3840 1390 3845
rect 4440 3845 4480 3850
rect 4440 3815 4445 3845
rect 4475 3840 4480 3845
rect 5750 3845 5790 3850
rect 5750 3840 5755 3845
rect 4475 3820 5755 3840
rect 4475 3815 4480 3820
rect 4440 3810 4480 3815
rect 5750 3815 5755 3820
rect 5785 3815 5790 3845
rect 5750 3810 5790 3815
rect -15 3795 25 3800
rect -15 3765 -10 3795
rect 20 3790 25 3795
rect 940 3795 980 3800
rect 940 3790 945 3795
rect 20 3770 945 3790
rect 20 3765 25 3770
rect -15 3760 25 3765
rect 940 3765 945 3770
rect 975 3765 980 3795
rect 940 3760 980 3765
rect 1635 3795 1685 3805
rect 2510 3800 2550 3805
rect 2510 3795 2515 3800
rect 1635 3765 1645 3795
rect 1675 3775 2515 3795
rect 1675 3765 1685 3775
rect 2510 3770 2515 3775
rect 2545 3770 2550 3800
rect 2510 3765 2550 3770
rect 4655 3795 4695 3800
rect 4655 3765 4660 3795
rect 4690 3790 4695 3795
rect 5135 3795 5185 3805
rect 5135 3790 5145 3795
rect 4690 3770 5145 3790
rect 4690 3765 4695 3770
rect 1635 3755 1685 3765
rect 4655 3760 4695 3765
rect 5135 3765 5145 3770
rect 5175 3765 5185 3795
rect 5135 3755 5185 3765
rect -60 3740 -20 3745
rect -60 3710 -55 3740
rect -25 3735 -20 3740
rect 2690 3740 2730 3745
rect 2690 3735 2695 3740
rect -25 3715 2695 3735
rect -25 3710 -20 3715
rect -60 3705 -20 3710
rect 2690 3710 2695 3715
rect 2725 3710 2730 3740
rect 2690 3705 2730 3710
rect 3385 3740 3435 3750
rect 3385 3710 3395 3740
rect 3425 3735 3435 3740
rect 4610 3740 4650 3745
rect 4610 3735 4615 3740
rect 3425 3715 4615 3735
rect 3425 3710 3435 3715
rect 3385 3700 3435 3710
rect 4610 3710 4615 3715
rect 4645 3710 4650 3740
rect 4610 3705 4650 3710
rect 1255 3690 1295 3695
rect 1255 3660 1260 3690
rect 1290 3685 1295 3690
rect 4390 3690 4430 3695
rect 4390 3685 4395 3690
rect 1290 3665 4395 3685
rect 1290 3660 1295 3665
rect 1255 3655 1295 3660
rect 4390 3660 4395 3665
rect 4425 3660 4430 3690
rect 4390 3655 4430 3660
rect 70 3640 110 3645
rect 70 3610 75 3640
rect 105 3635 110 3640
rect 2555 3640 2595 3645
rect 2555 3635 2560 3640
rect 105 3615 2560 3635
rect 105 3610 110 3615
rect 70 3605 110 3610
rect 2555 3610 2560 3615
rect 2590 3610 2595 3640
rect 2555 3605 2595 3610
rect 3310 3635 3350 3640
rect 3310 3605 3315 3635
rect 3345 3630 3350 3635
rect 3345 3610 6100 3630
rect 3345 3605 3350 3610
rect 3310 3600 3350 3605
rect 3200 3590 3240 3595
rect 66 3555 71 3590
rect 106 3555 111 3590
rect 3200 3560 3205 3590
rect 3235 3585 3240 3590
rect 4060 3590 4100 3595
rect 4060 3585 4065 3590
rect 3235 3565 4065 3585
rect 3235 3560 3240 3565
rect 3200 3555 3240 3560
rect 4060 3560 4065 3565
rect 4095 3585 4100 3590
rect 4565 3590 4605 3595
rect 4565 3585 4570 3590
rect 4095 3565 4570 3585
rect 4095 3560 4100 3565
rect 4060 3555 4100 3560
rect 4565 3560 4570 3565
rect 4600 3585 4605 3590
rect 4920 3590 4960 3595
rect 4920 3585 4925 3590
rect 4600 3565 4925 3585
rect 4600 3560 4605 3565
rect 4565 3555 4605 3560
rect 4920 3560 4925 3565
rect 4955 3560 4960 3590
rect 4920 3555 4960 3560
rect 3035 3530 3075 3535
rect -110 3525 -70 3530
rect -110 3495 -105 3525
rect -75 3520 -70 3525
rect 66 3520 71 3530
rect -75 3500 71 3520
rect -75 3495 -70 3500
rect 66 3495 71 3500
rect 106 3495 111 3530
rect 3035 3500 3040 3530
rect 3070 3525 3075 3530
rect 3145 3530 3185 3535
rect 3145 3525 3150 3530
rect 3070 3505 3150 3525
rect 3070 3500 3075 3505
rect 3035 3495 3075 3500
rect 3145 3500 3150 3505
rect 3180 3525 3185 3530
rect 3255 3530 3295 3535
rect 3255 3525 3260 3530
rect 3180 3505 3260 3525
rect 3180 3500 3185 3505
rect 3145 3495 3185 3500
rect 3255 3500 3260 3505
rect 3290 3525 3295 3530
rect 3365 3530 3405 3535
rect 3365 3525 3370 3530
rect 3290 3505 3370 3525
rect 3290 3500 3295 3505
rect 3255 3495 3295 3500
rect 3365 3500 3370 3505
rect 3400 3525 3405 3530
rect 3675 3530 3715 3535
rect 3675 3525 3680 3530
rect 3400 3505 3680 3525
rect 3400 3500 3405 3505
rect 3365 3495 3405 3500
rect 3675 3500 3680 3505
rect 3710 3525 3715 3530
rect 3785 3530 3825 3535
rect 3785 3525 3790 3530
rect 3710 3505 3790 3525
rect 3710 3500 3715 3505
rect 3675 3495 3715 3500
rect 3785 3500 3790 3505
rect 3820 3525 3825 3530
rect 3895 3530 3935 3535
rect 3895 3525 3900 3530
rect 3820 3505 3900 3525
rect 3820 3500 3825 3505
rect 3785 3495 3825 3500
rect 3895 3500 3900 3505
rect 3930 3525 3935 3530
rect 4005 3530 4045 3535
rect 4005 3525 4010 3530
rect 3930 3505 4010 3525
rect 3930 3500 3935 3505
rect 3895 3495 3935 3500
rect 4005 3500 4010 3505
rect 4040 3525 4045 3530
rect 4115 3530 4155 3535
rect 4115 3525 4120 3530
rect 4040 3505 4120 3525
rect 4040 3500 4045 3505
rect 4005 3495 4045 3500
rect 4115 3500 4120 3505
rect 4150 3525 4155 3530
rect 4225 3530 4265 3535
rect 4225 3525 4230 3530
rect 4150 3505 4230 3525
rect 4150 3500 4155 3505
rect 4115 3495 4155 3500
rect 4225 3500 4230 3505
rect 4260 3525 4265 3530
rect 4335 3530 4375 3535
rect 4335 3525 4340 3530
rect 4260 3505 4340 3525
rect 4260 3500 4265 3505
rect 4225 3495 4265 3500
rect 4335 3500 4340 3505
rect 4370 3525 4375 3530
rect 4445 3530 4485 3535
rect 4445 3525 4450 3530
rect 4370 3505 4450 3525
rect 4370 3500 4375 3505
rect 4335 3495 4375 3500
rect 4445 3500 4450 3505
rect 4480 3525 4485 3530
rect 4755 3530 4795 3535
rect 4755 3525 4760 3530
rect 4480 3505 4760 3525
rect 4480 3500 4485 3505
rect 4445 3495 4485 3500
rect 4755 3500 4760 3505
rect 4790 3525 4795 3530
rect 4865 3530 4905 3535
rect 4865 3525 4870 3530
rect 4790 3505 4870 3525
rect 4790 3500 4795 3505
rect 4755 3495 4795 3500
rect 4865 3500 4870 3505
rect 4900 3525 4905 3530
rect 4975 3530 5015 3535
rect 4975 3525 4980 3530
rect 4900 3505 4980 3525
rect 4900 3500 4905 3505
rect 4865 3495 4905 3500
rect 4975 3500 4980 3505
rect 5010 3525 5015 3530
rect 5085 3530 5125 3535
rect 5085 3525 5090 3530
rect 5010 3505 5090 3525
rect 5010 3500 5015 3505
rect 4975 3495 5015 3500
rect 5085 3500 5090 3505
rect 5120 3525 5125 3530
rect 5750 3530 5790 3535
rect 5750 3525 5755 3530
rect 5120 3505 5755 3525
rect 5120 3500 5125 3505
rect 5085 3495 5125 3500
rect 5750 3500 5755 3505
rect 5785 3500 5790 3530
rect 5750 3495 5790 3500
rect -110 3490 -70 3495
rect 1351 3420 1356 3455
rect 1391 3420 1396 3455
rect 70 3375 110 3380
rect 70 3345 75 3375
rect 105 3370 110 3375
rect 1255 3375 1295 3380
rect 1255 3370 1260 3375
rect 105 3350 1260 3370
rect 105 3345 110 3350
rect 70 3340 110 3345
rect 1255 3345 1260 3350
rect 1290 3345 1295 3375
rect 1351 3360 1356 3395
rect 1391 3360 1396 3395
rect 3090 3360 3130 3365
rect 1255 3340 1295 3345
rect 3090 3330 3095 3360
rect 3125 3355 3130 3360
rect 3200 3360 3240 3365
rect 3200 3355 3205 3360
rect 3125 3335 3205 3355
rect 3125 3330 3130 3335
rect 3090 3325 3130 3330
rect 3200 3330 3205 3335
rect 3235 3355 3240 3360
rect 3310 3360 3350 3365
rect 3310 3355 3315 3360
rect 3235 3335 3315 3355
rect 3235 3330 3240 3335
rect 3200 3325 3240 3330
rect 3310 3330 3315 3335
rect 3345 3330 3350 3360
rect 3310 3325 3350 3330
rect 3840 3360 3880 3365
rect 3840 3330 3845 3360
rect 3875 3355 3880 3360
rect 3950 3360 3990 3365
rect 3950 3355 3955 3360
rect 3875 3335 3955 3355
rect 3875 3330 3880 3335
rect 3840 3325 3880 3330
rect 3950 3330 3955 3335
rect 3985 3355 3990 3360
rect 4060 3360 4100 3365
rect 4060 3355 4065 3360
rect 3985 3335 4065 3355
rect 3985 3330 3990 3335
rect 3950 3325 3990 3330
rect 4060 3330 4065 3335
rect 4095 3355 4100 3360
rect 4170 3360 4210 3365
rect 4170 3355 4175 3360
rect 4095 3335 4175 3355
rect 4095 3330 4100 3335
rect 4060 3325 4100 3330
rect 4170 3330 4175 3335
rect 4205 3355 4210 3360
rect 4280 3360 4320 3365
rect 4280 3355 4285 3360
rect 4205 3335 4285 3355
rect 4205 3330 4210 3335
rect 4170 3325 4210 3330
rect 4280 3330 4285 3335
rect 4315 3330 4320 3360
rect 4280 3325 4320 3330
rect 4810 3360 4850 3365
rect 4810 3330 4815 3360
rect 4845 3355 4850 3360
rect 4920 3360 4960 3365
rect 4920 3355 4925 3360
rect 4845 3335 4925 3355
rect 4845 3330 4850 3335
rect 4810 3325 4850 3330
rect 4920 3330 4925 3335
rect 4955 3355 4960 3360
rect 5030 3360 5070 3365
rect 5030 3355 5035 3360
rect 4955 3335 5035 3355
rect 4955 3330 4960 3335
rect 4920 3325 4960 3330
rect 5030 3330 5035 3335
rect 5065 3355 5070 3360
rect 5065 3335 6100 3355
rect 5065 3330 5070 3335
rect 5030 3325 5070 3330
rect 66 3290 71 3325
rect 106 3290 111 3325
rect 4565 3315 4605 3320
rect 1185 3290 1225 3295
rect -110 3260 -70 3265
rect -110 3230 -105 3260
rect -75 3255 -70 3260
rect 66 3255 71 3265
rect -75 3235 71 3255
rect -75 3230 -70 3235
rect 66 3230 71 3235
rect 106 3230 111 3265
rect 1185 3260 1190 3290
rect 1220 3285 1225 3290
rect 1290 3290 1330 3295
rect 1290 3285 1295 3290
rect 1220 3265 1295 3285
rect 1220 3260 1225 3265
rect 1185 3255 1225 3260
rect 1290 3260 1295 3265
rect 1325 3260 1330 3290
rect 4565 3285 4570 3315
rect 4600 3310 4605 3315
rect 4600 3305 5010 3310
rect 4600 3290 4975 3305
rect 4600 3285 4605 3290
rect 4565 3280 4605 3285
rect 4970 3275 4975 3290
rect 5005 3275 5010 3305
rect 4970 3270 5010 3275
rect 4610 3260 4650 3265
rect 1290 3255 1330 3260
rect 2555 3255 2595 3260
rect -110 3225 -70 3230
rect 2555 3225 2560 3255
rect 2590 3250 2595 3255
rect 2610 3255 2650 3260
rect 2610 3250 2615 3255
rect 2590 3230 2615 3250
rect 2590 3225 2595 3230
rect 2555 3220 2595 3225
rect 2610 3225 2615 3230
rect 2645 3225 2650 3255
rect 4610 3230 4615 3260
rect 4645 3255 4650 3260
rect 5060 3260 5100 3265
rect 5060 3255 5065 3260
rect 4645 3235 5065 3255
rect 4645 3230 4650 3235
rect 4610 3225 4650 3230
rect 5060 3230 5065 3235
rect 5095 3230 5100 3260
rect 5060 3225 5100 3230
rect 2610 3220 2650 3225
rect -110 3195 -70 3200
rect -110 3165 -105 3195
rect -75 3190 -70 3195
rect 595 3195 635 3200
rect 595 3190 600 3195
rect -75 3170 600 3190
rect -75 3165 -70 3170
rect -110 3160 -70 3165
rect 595 3165 600 3170
rect 630 3165 635 3195
rect 2420 3180 2425 3215
rect 2460 3205 2465 3215
rect 3060 3210 3100 3215
rect 3060 3205 3065 3210
rect 2460 3185 3065 3205
rect 2460 3180 2465 3185
rect 3060 3180 3065 3185
rect 3095 3180 3100 3210
rect 3060 3175 3100 3180
rect 4655 3205 4695 3210
rect 4655 3175 4660 3205
rect 4690 3200 4695 3205
rect 5015 3205 5055 3210
rect 5015 3200 5020 3205
rect 4690 3180 5020 3200
rect 4690 3175 4695 3180
rect 4655 3170 4695 3175
rect 5015 3175 5020 3180
rect 5050 3175 5055 3205
rect 5015 3170 5055 3175
rect 595 3160 635 3165
rect 2555 3165 2595 3170
rect 2420 3155 2465 3160
rect 2420 3120 2425 3155
rect 2460 3120 2465 3155
rect 2555 3135 2560 3165
rect 2590 3160 2595 3165
rect 3730 3165 3770 3170
rect 3730 3160 3735 3165
rect 2590 3140 3735 3160
rect 2590 3135 2595 3140
rect 2555 3130 2595 3135
rect 3730 3135 3735 3140
rect 3765 3135 3770 3165
rect 3730 3130 3770 3135
rect 4390 3160 4430 3165
rect 4390 3130 4395 3160
rect 4425 3155 4430 3160
rect 5615 3160 5655 3165
rect 5615 3155 5620 3160
rect 4425 3135 5620 3155
rect 4425 3130 4430 3135
rect 2420 3115 2465 3120
rect 4060 3125 4100 3130
rect 4390 3125 4430 3130
rect 5615 3130 5620 3135
rect 5650 3130 5655 3160
rect 5615 3125 5655 3130
rect 4060 3095 4065 3125
rect 4095 3110 4100 3125
rect 4095 3095 6100 3110
rect 4060 3090 6100 3095
rect 3250 3065 3290 3070
rect -60 3055 -20 3060
rect -60 3025 -55 3055
rect -25 3050 -20 3055
rect 261 3050 266 3060
rect -25 3030 266 3050
rect -25 3025 -20 3030
rect 261 3025 266 3030
rect 301 3025 306 3060
rect 934 3025 939 3060
rect 974 3050 979 3060
rect 1210 3055 1250 3060
rect 1210 3050 1215 3055
rect 974 3030 1215 3050
rect 974 3025 979 3030
rect 1210 3025 1215 3030
rect 1245 3025 1250 3055
rect 3250 3050 3255 3065
rect -60 3020 -20 3025
rect 1210 3020 1250 3025
rect 2825 3035 3255 3050
rect 3285 3060 3290 3065
rect 3430 3065 3470 3070
rect 3430 3060 3435 3065
rect 3285 3040 3435 3060
rect 3285 3035 3290 3040
rect 2825 3030 3290 3035
rect 3430 3035 3435 3040
rect 3465 3060 3470 3065
rect 3610 3065 3650 3070
rect 3610 3060 3615 3065
rect 3465 3040 3615 3060
rect 3465 3035 3470 3040
rect 3430 3030 3470 3035
rect 3610 3035 3615 3040
rect 3645 3060 3650 3065
rect 3790 3065 3830 3070
rect 3790 3060 3795 3065
rect 3645 3040 3795 3060
rect 3645 3035 3650 3040
rect 3610 3030 3650 3035
rect 3790 3035 3795 3040
rect 3825 3060 3830 3065
rect 3970 3065 4010 3070
rect 3970 3060 3975 3065
rect 3825 3040 3975 3060
rect 3825 3035 3830 3040
rect 3790 3030 3830 3035
rect 3970 3035 3975 3040
rect 4005 3060 4010 3065
rect 4150 3065 4190 3070
rect 4150 3060 4155 3065
rect 4005 3040 4155 3060
rect 4005 3035 4010 3040
rect 3970 3030 4010 3035
rect 4150 3035 4155 3040
rect 4185 3060 4190 3065
rect 4330 3065 4370 3070
rect 4330 3060 4335 3065
rect 4185 3040 4335 3060
rect 4185 3035 4190 3040
rect 4150 3030 4190 3035
rect 4330 3035 4335 3040
rect 4365 3060 4370 3065
rect 4510 3065 4550 3070
rect 4510 3060 4515 3065
rect 4365 3040 4515 3060
rect 4365 3035 4370 3040
rect 4330 3030 4370 3035
rect 4510 3035 4515 3040
rect 4545 3060 4550 3065
rect 4690 3065 4730 3070
rect 4690 3060 4695 3065
rect 4545 3040 4695 3060
rect 4545 3035 4550 3040
rect 4510 3030 4550 3035
rect 4690 3035 4695 3040
rect 4725 3060 4730 3065
rect 4870 3065 4910 3070
rect 4870 3060 4875 3065
rect 4725 3040 4875 3060
rect 4725 3035 4730 3040
rect 4690 3030 4730 3035
rect 4870 3035 4875 3040
rect 4905 3060 4910 3065
rect 5750 3065 5790 3070
rect 5750 3060 5755 3065
rect 4905 3040 5755 3060
rect 4905 3035 4910 3040
rect 4870 3030 4910 3035
rect 2825 3025 2865 3030
rect 2825 2995 2830 3025
rect 2860 2995 2865 3025
rect 2825 2990 2865 2995
rect 5290 3025 5330 3040
rect 5750 3035 5755 3040
rect 5785 3035 5790 3065
rect 5750 3030 5790 3035
rect 5290 2995 5295 3025
rect 5325 2995 5330 3025
rect 5290 2990 5330 2995
rect 2825 2965 2865 2970
rect 1105 2950 1145 2955
rect 1105 2920 1110 2950
rect 1140 2945 1145 2950
rect 1516 2945 1521 2950
rect 1140 2925 1521 2945
rect 1140 2920 1145 2925
rect 1105 2915 1145 2920
rect 1516 2915 1521 2925
rect 1556 2915 1561 2950
rect 2215 2915 2220 2950
rect 2255 2940 2260 2950
rect 2420 2945 2460 2950
rect 2420 2940 2425 2945
rect 2255 2920 2425 2940
rect 2255 2915 2260 2920
rect 2420 2915 2425 2920
rect 2455 2915 2460 2945
rect 2825 2935 2830 2965
rect 2860 2960 2865 2965
rect 3060 2965 3100 2970
rect 3060 2960 3065 2965
rect 2860 2940 3065 2960
rect 2860 2935 2865 2940
rect 2825 2930 2865 2935
rect 3060 2935 3065 2940
rect 3095 2935 3100 2965
rect 3060 2930 3100 2935
rect 5290 2965 5330 2970
rect 5290 2935 5295 2965
rect 5325 2935 5330 2965
rect 5290 2930 5330 2935
rect 2420 2910 2460 2915
rect -15 2850 25 2855
rect -15 2820 -10 2850
rect 20 2840 25 2850
rect 261 2840 266 2850
rect 20 2820 266 2840
rect -15 2815 25 2820
rect 261 2815 266 2820
rect 301 2815 306 2850
rect 934 2815 939 2850
rect 974 2840 979 2850
rect 2465 2845 2505 2850
rect 2465 2840 2470 2845
rect 974 2820 2470 2840
rect 974 2815 979 2820
rect 2465 2815 2470 2820
rect 2500 2815 2505 2845
rect 2465 2810 2505 2815
rect 1210 2800 1250 2805
rect 1210 2770 1215 2800
rect 1245 2795 1250 2800
rect 2375 2800 2415 2805
rect 2375 2795 2380 2800
rect 1245 2775 2380 2795
rect 1245 2770 1250 2775
rect 1210 2765 1250 2770
rect 2375 2770 2380 2775
rect 2410 2770 2415 2800
rect 2375 2765 2415 2770
rect 2760 2795 2800 2800
rect 2760 2765 2765 2795
rect 2795 2790 2800 2795
rect 2890 2795 2930 2800
rect 2890 2790 2895 2795
rect 2795 2770 2895 2790
rect 2795 2765 2800 2770
rect 2760 2760 2800 2765
rect 2890 2765 2895 2770
rect 2925 2790 2930 2795
rect 3120 2795 3160 2800
rect 3120 2790 3125 2795
rect 2925 2770 3125 2790
rect 2925 2765 2930 2770
rect 2890 2760 2930 2765
rect 3120 2765 3125 2770
rect 3155 2765 3160 2795
rect 3120 2760 3160 2765
rect 5225 2795 5265 2800
rect 5225 2765 5230 2795
rect 5260 2790 5265 2795
rect 5355 2795 5395 2800
rect 5355 2790 5360 2795
rect 5260 2770 5360 2790
rect 5260 2765 5265 2770
rect 5225 2760 5265 2765
rect 5355 2765 5360 2770
rect 5390 2790 5395 2795
rect 5390 2770 6100 2790
rect 5390 2765 5395 2770
rect 5355 2760 5395 2765
rect 2420 2695 2460 2700
rect 2420 2665 2425 2695
rect 2455 2690 2460 2695
rect 3880 2695 3920 2700
rect 3880 2690 3885 2695
rect 2455 2670 3885 2690
rect 2455 2665 2460 2670
rect 2420 2660 2460 2665
rect 3880 2665 3885 2670
rect 3915 2690 3920 2695
rect 4240 2695 4280 2700
rect 4240 2690 4245 2695
rect 3915 2670 4245 2690
rect 3915 2665 3920 2670
rect 3880 2660 3920 2665
rect 4240 2665 4245 2670
rect 4275 2665 4280 2695
rect 4240 2660 4280 2665
rect 5060 2650 5100 2655
rect 2330 2640 2370 2645
rect 2330 2610 2335 2640
rect 2365 2635 2370 2640
rect 3060 2640 3100 2645
rect 3060 2635 3065 2640
rect 2365 2615 3065 2635
rect 2365 2610 2370 2615
rect 2330 2605 2370 2610
rect 3060 2610 3065 2615
rect 3095 2635 3100 2640
rect 3700 2640 3740 2645
rect 3700 2635 3705 2640
rect 3095 2615 3705 2635
rect 3095 2610 3100 2615
rect 3060 2605 3100 2610
rect 3700 2610 3705 2615
rect 3735 2635 3740 2640
rect 4420 2640 4460 2645
rect 4420 2635 4425 2640
rect 3735 2615 4425 2635
rect 3735 2610 3740 2615
rect 3700 2605 3740 2610
rect 4420 2610 4425 2615
rect 4455 2610 4460 2640
rect 5060 2620 5065 2650
rect 5095 2645 5100 2650
rect 5525 2650 5565 2655
rect 5525 2645 5530 2650
rect 5095 2625 5530 2645
rect 5095 2620 5100 2625
rect 5060 2615 5100 2620
rect 5525 2620 5530 2625
rect 5560 2620 5565 2650
rect 5525 2615 5565 2620
rect 4420 2605 4460 2610
rect 2275 2595 2315 2600
rect 2275 2565 2280 2595
rect 2310 2590 2315 2595
rect 2825 2595 2865 2600
rect 2825 2590 2830 2595
rect 2310 2570 2830 2590
rect 2310 2565 2315 2570
rect 2275 2560 2315 2565
rect 2825 2565 2830 2570
rect 2860 2590 2865 2595
rect 3520 2595 3560 2600
rect 3520 2590 3525 2595
rect 2860 2570 3525 2590
rect 2860 2565 2865 2570
rect 2825 2560 2865 2565
rect 3520 2565 3525 2570
rect 3555 2590 3560 2595
rect 4600 2595 4640 2600
rect 4600 2590 4605 2595
rect 3555 2570 4605 2590
rect 3555 2565 3560 2570
rect 3520 2560 3560 2565
rect 4600 2565 4605 2570
rect 4635 2565 4640 2595
rect 4600 2560 4640 2565
rect 4690 2595 4730 2600
rect 4690 2565 4695 2595
rect 4725 2590 4730 2595
rect 5015 2595 5055 2600
rect 5015 2590 5020 2595
rect 4725 2570 5020 2590
rect 4725 2565 4730 2570
rect 4690 2560 4730 2565
rect 5015 2565 5020 2570
rect 5050 2565 5055 2595
rect 5015 2560 5055 2565
rect 2610 2550 2650 2555
rect 2610 2520 2615 2550
rect 2645 2545 2650 2550
rect 3340 2550 3380 2555
rect 3340 2545 3345 2550
rect 2645 2525 3345 2545
rect 2645 2520 2650 2525
rect 2610 2515 2650 2520
rect 3340 2520 3345 2525
rect 3375 2545 3380 2550
rect 4060 2550 4100 2555
rect 4060 2545 4065 2550
rect 3375 2525 4065 2545
rect 3375 2520 3380 2525
rect 3340 2515 3380 2520
rect 4060 2520 4065 2525
rect 4095 2545 4100 2550
rect 4780 2550 4820 2555
rect 4780 2545 4785 2550
rect 4095 2525 4785 2545
rect 4095 2520 4100 2525
rect 4060 2515 4100 2520
rect 4780 2520 4785 2525
rect 4815 2545 4820 2550
rect 5570 2550 5610 2555
rect 5570 2545 5575 2550
rect 4815 2525 5575 2545
rect 4815 2520 4820 2525
rect 4780 2515 4820 2520
rect 5570 2520 5575 2525
rect 5605 2520 5610 2550
rect 5570 2515 5610 2520
rect 2375 2500 2415 2505
rect 2375 2470 2380 2500
rect 2410 2495 2415 2500
rect 4280 2500 4320 2505
rect 4280 2495 4285 2500
rect 2410 2475 4285 2495
rect 2410 2470 2415 2475
rect 2375 2465 2415 2470
rect 4280 2470 4285 2475
rect 4315 2495 4320 2500
rect 4970 2500 5010 2505
rect 4970 2495 4975 2500
rect 4315 2475 4975 2495
rect 4315 2470 4320 2475
rect 4280 2465 4320 2470
rect 4970 2470 4975 2475
rect 5005 2495 5010 2500
rect 5290 2500 5330 2505
rect 5290 2495 5295 2500
rect 5005 2475 5295 2495
rect 5005 2470 5010 2475
rect 4970 2465 5010 2470
rect 5290 2470 5295 2475
rect 5325 2470 5330 2500
rect 5290 2465 5330 2470
rect 2820 2435 2860 2440
rect 2820 2405 2825 2435
rect 2855 2430 2860 2435
rect 2940 2435 2980 2440
rect 2940 2430 2945 2435
rect 2855 2410 2945 2430
rect 2855 2405 2860 2410
rect 2820 2400 2860 2405
rect 2940 2405 2945 2410
rect 2975 2430 2980 2435
rect 3060 2435 3100 2440
rect 3060 2430 3065 2435
rect 2975 2410 3065 2430
rect 2975 2405 2980 2410
rect 2940 2400 2980 2405
rect 3060 2405 3065 2410
rect 3095 2430 3100 2435
rect 3180 2435 3220 2440
rect 3180 2430 3185 2435
rect 3095 2410 3185 2430
rect 3095 2405 3100 2410
rect 3060 2400 3100 2405
rect 3180 2405 3185 2410
rect 3215 2430 3220 2435
rect 3300 2435 3340 2440
rect 3300 2430 3305 2435
rect 3215 2410 3305 2430
rect 3215 2405 3220 2410
rect 3180 2400 3220 2405
rect 3300 2405 3305 2410
rect 3335 2430 3340 2435
rect 3420 2435 3460 2440
rect 3420 2430 3425 2435
rect 3335 2410 3425 2430
rect 3335 2405 3340 2410
rect 3300 2400 3340 2405
rect 3420 2405 3425 2410
rect 3455 2430 3460 2435
rect 3540 2435 3580 2440
rect 3540 2430 3545 2435
rect 3455 2410 3545 2430
rect 3455 2405 3460 2410
rect 3420 2400 3460 2405
rect 3540 2405 3545 2410
rect 3575 2430 3580 2435
rect 3660 2435 3700 2440
rect 3660 2430 3665 2435
rect 3575 2410 3665 2430
rect 3575 2405 3580 2410
rect 3540 2400 3580 2405
rect 3660 2405 3665 2410
rect 3695 2430 3700 2435
rect 3780 2435 3820 2440
rect 3780 2430 3785 2435
rect 3695 2410 3785 2430
rect 3695 2405 3700 2410
rect 3660 2400 3700 2405
rect 3780 2405 3785 2410
rect 3815 2430 3820 2435
rect 4340 2435 4380 2440
rect 4340 2430 4345 2435
rect 3815 2410 4345 2430
rect 3815 2405 3820 2410
rect 3780 2400 3820 2405
rect 4340 2405 4345 2410
rect 4375 2430 4380 2435
rect 4460 2435 4500 2440
rect 4460 2430 4465 2435
rect 4375 2410 4465 2430
rect 4375 2405 4380 2410
rect 4340 2400 4380 2405
rect 4460 2405 4465 2410
rect 4495 2430 4500 2435
rect 4580 2435 4620 2440
rect 4580 2430 4585 2435
rect 4495 2410 4585 2430
rect 4495 2405 4500 2410
rect 4460 2400 4500 2405
rect 4580 2405 4585 2410
rect 4615 2430 4620 2435
rect 4700 2435 4740 2440
rect 4700 2430 4705 2435
rect 4615 2410 4705 2430
rect 4615 2405 4620 2410
rect 4580 2400 4620 2405
rect 4700 2405 4705 2410
rect 4735 2430 4740 2435
rect 4820 2435 4860 2440
rect 4820 2430 4825 2435
rect 4735 2410 4825 2430
rect 4735 2405 4740 2410
rect 4700 2400 4740 2405
rect 4820 2405 4825 2410
rect 4855 2430 4860 2435
rect 4940 2435 4980 2440
rect 4940 2430 4945 2435
rect 4855 2410 4945 2430
rect 4855 2405 4860 2410
rect 4820 2400 4860 2405
rect 4940 2405 4945 2410
rect 4975 2430 4980 2435
rect 5060 2435 5100 2440
rect 5060 2430 5065 2435
rect 4975 2410 5065 2430
rect 4975 2405 4980 2410
rect 4940 2400 4980 2405
rect 5060 2405 5065 2410
rect 5095 2430 5100 2435
rect 5180 2435 5220 2440
rect 5180 2430 5185 2435
rect 5095 2410 5185 2430
rect 5095 2405 5100 2410
rect 5060 2400 5100 2405
rect 5180 2405 5185 2410
rect 5215 2430 5220 2435
rect 5300 2435 5340 2440
rect 5300 2430 5305 2435
rect 5215 2410 5305 2430
rect 5215 2405 5220 2410
rect 5180 2400 5220 2405
rect 5300 2405 5305 2410
rect 5335 2430 5340 2435
rect 5750 2435 5790 2440
rect 5750 2430 5755 2435
rect 5335 2410 5755 2430
rect 5335 2405 5340 2410
rect 5300 2400 5340 2405
rect 5750 2405 5755 2410
rect 5785 2405 5790 2435
rect 5750 2400 5790 2405
rect 2465 2375 2505 2380
rect 2465 2345 2470 2375
rect 2500 2370 2505 2375
rect 2760 2375 2800 2380
rect 2760 2370 2765 2375
rect 2500 2350 2765 2370
rect 2500 2345 2505 2350
rect 2465 2340 2505 2345
rect 2760 2345 2765 2350
rect 2795 2370 2800 2375
rect 3120 2375 3160 2380
rect 3120 2370 3125 2375
rect 2795 2350 3125 2370
rect 2795 2345 2800 2350
rect 2760 2340 2800 2345
rect 3120 2345 3125 2350
rect 3155 2370 3160 2375
rect 3480 2375 3520 2380
rect 3480 2370 3485 2375
rect 3155 2350 3485 2370
rect 3155 2345 3160 2350
rect 3120 2340 3160 2345
rect 3480 2345 3485 2350
rect 3515 2370 3520 2375
rect 3840 2375 3880 2380
rect 3840 2370 3845 2375
rect 3515 2350 3845 2370
rect 3515 2345 3520 2350
rect 3480 2340 3520 2345
rect 3840 2345 3845 2350
rect 3875 2370 3880 2375
rect 3970 2375 4010 2380
rect 3970 2370 3975 2375
rect 3875 2350 3975 2370
rect 3875 2345 3880 2350
rect 3840 2340 3880 2345
rect 3970 2345 3975 2350
rect 4005 2345 4010 2375
rect 3970 2340 4010 2345
rect 4150 2375 4190 2380
rect 4150 2345 4155 2375
rect 4185 2370 4190 2375
rect 4280 2375 4320 2380
rect 4280 2370 4285 2375
rect 4185 2350 4285 2370
rect 4185 2345 4190 2350
rect 4150 2340 4190 2345
rect 4280 2345 4285 2350
rect 4315 2370 4320 2375
rect 4640 2375 4680 2380
rect 4640 2370 4645 2375
rect 4315 2350 4645 2370
rect 4315 2345 4320 2350
rect 4280 2340 4320 2345
rect 4640 2345 4645 2350
rect 4675 2370 4680 2375
rect 5000 2375 5040 2380
rect 5000 2370 5005 2375
rect 4675 2350 5005 2370
rect 4675 2345 4680 2350
rect 4640 2340 4680 2345
rect 5000 2345 5005 2350
rect 5035 2370 5040 2375
rect 5360 2375 5400 2380
rect 5360 2370 5365 2375
rect 5035 2350 5365 2370
rect 5035 2345 5040 2350
rect 5000 2340 5040 2345
rect 5360 2345 5365 2350
rect 5395 2345 5400 2375
rect 5360 2340 5400 2345
rect 2880 2205 2920 2210
rect 2880 2175 2885 2205
rect 2915 2200 2920 2205
rect 3000 2200 3040 2210
rect 3240 2205 3280 2210
rect 3240 2200 3245 2205
rect 2915 2180 3245 2200
rect 2915 2175 2920 2180
rect 2880 2170 2920 2175
rect 3000 2170 3040 2180
rect 3240 2175 3245 2180
rect 3275 2200 3280 2205
rect 3360 2200 3400 2210
rect 3600 2205 3640 2210
rect 3600 2200 3605 2205
rect 3275 2180 3605 2200
rect 3275 2175 3280 2180
rect 3240 2170 3280 2175
rect 3360 2170 3400 2180
rect 3600 2175 3605 2180
rect 3635 2175 3640 2205
rect 3600 2170 3640 2175
rect 3720 2170 3760 2210
rect 4400 2170 4440 2210
rect 4520 2205 4560 2210
rect 4520 2175 4525 2205
rect 4555 2200 4560 2205
rect 4760 2200 4800 2210
rect 4880 2205 4920 2210
rect 4880 2200 4885 2205
rect 4555 2180 4885 2200
rect 4555 2175 4560 2180
rect 4520 2170 4560 2175
rect 4760 2170 4800 2180
rect 4880 2175 4885 2180
rect 4915 2200 4920 2205
rect 5120 2200 5160 2210
rect 5240 2205 5280 2210
rect 5240 2200 5245 2205
rect 4915 2180 5245 2200
rect 4915 2175 4920 2180
rect 4880 2170 4920 2175
rect 5120 2170 5160 2180
rect 5240 2175 5245 2180
rect 5275 2175 5280 2205
rect 5240 2170 5280 2175
rect 2510 2145 2550 2150
rect 2510 2115 2515 2145
rect 2545 2140 2550 2145
rect 2790 2145 2830 2150
rect 2790 2140 2795 2145
rect 2545 2120 2795 2140
rect 2545 2115 2550 2120
rect 2510 2110 2550 2115
rect 2790 2115 2795 2120
rect 2825 2140 2830 2145
rect 3000 2145 3040 2150
rect 3000 2140 3005 2145
rect 2825 2120 3005 2140
rect 2825 2115 2830 2120
rect 2790 2110 2830 2115
rect 3000 2115 3005 2120
rect 3035 2140 3040 2145
rect 3120 2145 3160 2150
rect 3120 2140 3125 2145
rect 3035 2120 3125 2140
rect 3035 2115 3040 2120
rect 3000 2110 3040 2115
rect 3120 2115 3125 2120
rect 3155 2140 3160 2145
rect 3360 2145 3400 2150
rect 3360 2140 3365 2145
rect 3155 2120 3365 2140
rect 3155 2115 3160 2120
rect 3120 2110 3160 2115
rect 3360 2115 3365 2120
rect 3395 2140 3400 2145
rect 3480 2145 3520 2150
rect 3480 2140 3485 2145
rect 3395 2120 3485 2140
rect 3395 2115 3400 2120
rect 3360 2110 3400 2115
rect 3480 2115 3485 2120
rect 3515 2140 3520 2145
rect 3720 2145 3760 2150
rect 3720 2140 3725 2145
rect 3515 2120 3725 2140
rect 3515 2115 3520 2120
rect 3480 2110 3520 2115
rect 3720 2115 3725 2120
rect 3755 2140 3760 2145
rect 3810 2145 3850 2150
rect 3810 2140 3815 2145
rect 3755 2120 3815 2140
rect 3755 2115 3760 2120
rect 3720 2110 3760 2115
rect 3810 2115 3815 2120
rect 3845 2115 3850 2145
rect 3810 2110 3850 2115
rect 4310 2145 4350 2150
rect 4310 2115 4315 2145
rect 4345 2140 4350 2145
rect 4400 2145 4440 2150
rect 4400 2140 4405 2145
rect 4345 2120 4405 2140
rect 4345 2115 4350 2120
rect 4310 2110 4350 2115
rect 4400 2115 4405 2120
rect 4435 2140 4440 2145
rect 4640 2145 4680 2150
rect 4640 2140 4645 2145
rect 4435 2120 4645 2140
rect 4435 2115 4440 2120
rect 4400 2110 4440 2115
rect 4640 2115 4645 2120
rect 4675 2140 4680 2145
rect 4760 2145 4800 2150
rect 4760 2140 4765 2145
rect 4675 2120 4765 2140
rect 4675 2115 4680 2120
rect 4640 2110 4680 2115
rect 4760 2115 4765 2120
rect 4795 2140 4800 2145
rect 5000 2145 5040 2150
rect 5000 2140 5005 2145
rect 4795 2120 5005 2140
rect 4795 2115 4800 2120
rect 4760 2110 4800 2115
rect 5000 2115 5005 2120
rect 5035 2140 5040 2145
rect 5120 2145 5160 2150
rect 5120 2140 5125 2145
rect 5035 2120 5125 2140
rect 5035 2115 5040 2120
rect 5000 2110 5040 2115
rect 5120 2115 5125 2120
rect 5155 2140 5160 2145
rect 5330 2145 5370 2150
rect 5330 2140 5335 2145
rect 5155 2120 5335 2140
rect 5155 2115 5160 2120
rect 5120 2110 5160 2115
rect 5330 2115 5335 2120
rect 5365 2140 5370 2145
rect 5525 2145 5565 2150
rect 5525 2140 5530 2145
rect 5365 2120 5530 2140
rect 5365 2115 5370 2120
rect 5330 2110 5370 2115
rect 5525 2115 5530 2120
rect 5560 2115 5565 2145
rect 5525 2110 5565 2115
rect 3250 2060 3290 2065
rect 2330 2045 2370 2050
rect 2330 2015 2335 2045
rect 2365 2040 2370 2045
rect 3190 2045 3230 2050
rect 3190 2040 3195 2045
rect 2365 2020 3195 2040
rect 2365 2015 2370 2020
rect 2330 2010 2370 2015
rect 3190 2015 3195 2020
rect 3225 2015 3230 2045
rect 3250 2030 3255 2060
rect 3285 2055 3290 2060
rect 3490 2060 3530 2065
rect 3490 2055 3495 2060
rect 3285 2035 3495 2055
rect 3285 2030 3290 2035
rect 3250 2025 3290 2030
rect 3490 2030 3495 2035
rect 3525 2055 3530 2060
rect 3730 2060 3770 2065
rect 3730 2055 3735 2060
rect 3525 2035 3735 2055
rect 3525 2030 3530 2035
rect 3490 2025 3530 2030
rect 3730 2030 3735 2035
rect 3765 2030 3770 2060
rect 3730 2025 3770 2030
rect 4390 2060 4430 2065
rect 4390 2030 4395 2060
rect 4425 2055 4430 2060
rect 4630 2060 4670 2065
rect 4630 2055 4635 2060
rect 4425 2035 4635 2055
rect 4425 2030 4430 2035
rect 4390 2025 4430 2030
rect 4630 2030 4635 2035
rect 4665 2055 4670 2060
rect 4870 2060 4910 2065
rect 4870 2055 4875 2060
rect 4665 2035 4875 2055
rect 4665 2030 4670 2035
rect 4630 2025 4670 2030
rect 4870 2030 4875 2035
rect 4905 2030 4910 2060
rect 4870 2025 4910 2030
rect 4930 2045 4970 2050
rect 3190 2010 3230 2015
rect 4930 2015 4935 2045
rect 4965 2040 4970 2045
rect 5570 2045 5610 2050
rect 5570 2040 5575 2045
rect 4965 2020 5575 2040
rect 4965 2015 4970 2020
rect 4930 2010 4970 2015
rect 5570 2015 5575 2020
rect 5605 2040 5610 2045
rect 5605 2020 6100 2040
rect 5605 2015 5610 2020
rect 5570 2010 5610 2015
rect 3130 2000 3170 2005
rect 3130 1970 3135 2000
rect 3165 1995 3170 2000
rect 3370 2000 3410 2005
rect 3370 1995 3375 2000
rect 3165 1975 3375 1995
rect 3165 1970 3170 1975
rect 3130 1965 3170 1970
rect 3370 1970 3375 1975
rect 3405 1995 3410 2000
rect 3610 2000 3650 2005
rect 3610 1995 3615 2000
rect 3405 1975 3615 1995
rect 3405 1970 3410 1975
rect 3370 1965 3410 1970
rect 3610 1970 3615 1975
rect 3645 1970 3650 2000
rect 3610 1965 3650 1970
rect 4510 2000 4550 2005
rect 4510 1970 4515 2000
rect 4545 1995 4550 2000
rect 4750 2000 4790 2005
rect 4750 1995 4755 2000
rect 4545 1975 4755 1995
rect 4545 1970 4550 1975
rect 4510 1965 4550 1970
rect 4750 1970 4755 1975
rect 4785 1995 4790 2000
rect 4990 2000 5030 2005
rect 4990 1995 4995 2000
rect 4785 1975 4995 1995
rect 4785 1970 4790 1975
rect 4750 1965 4790 1970
rect 4990 1970 4995 1975
rect 5025 1970 5030 2000
rect 4990 1965 5030 1970
rect 3790 1940 3830 1945
rect 3790 1910 3795 1940
rect 3825 1935 3830 1940
rect 4060 1940 4100 1945
rect 4060 1935 4065 1940
rect 3825 1915 4065 1935
rect 3825 1910 3830 1915
rect 3790 1905 3830 1910
rect 4060 1910 4065 1915
rect 4095 1935 4100 1940
rect 4330 1940 4370 1945
rect 4330 1935 4335 1940
rect 4095 1915 4335 1935
rect 4095 1910 4100 1915
rect 4060 1905 4100 1910
rect 4330 1910 4335 1915
rect 4365 1910 4370 1940
rect 4330 1905 4370 1910
rect 2420 1880 2460 1885
rect 2420 1850 2425 1880
rect 2455 1875 2460 1880
rect 3130 1880 3170 1885
rect 3130 1875 3135 1880
rect 2455 1855 3135 1875
rect 2455 1850 2460 1855
rect 2420 1845 2460 1850
rect 3130 1850 3135 1855
rect 3165 1850 3170 1880
rect 3130 1845 3170 1850
rect 4990 1880 5030 1885
rect 4990 1850 4995 1880
rect 5025 1875 5030 1880
rect 5615 1880 5655 1885
rect 5615 1875 5620 1880
rect 5025 1855 5620 1875
rect 5025 1850 5030 1855
rect 4990 1845 5030 1850
rect 5615 1850 5620 1855
rect 5650 1850 5655 1880
rect 5615 1845 5655 1850
rect 2890 1820 2930 1825
rect 2890 1790 2895 1820
rect 2925 1815 2930 1820
rect 3190 1820 3230 1825
rect 3190 1815 3195 1820
rect 2925 1795 3195 1815
rect 2925 1790 2930 1795
rect 2890 1785 2930 1790
rect 3190 1790 3195 1795
rect 3225 1815 3230 1820
rect 3310 1820 3350 1825
rect 3310 1815 3315 1820
rect 3225 1795 3315 1815
rect 3225 1790 3230 1795
rect 3190 1785 3230 1790
rect 3310 1790 3315 1795
rect 3345 1815 3350 1820
rect 3430 1820 3470 1825
rect 3430 1815 3435 1820
rect 3345 1795 3435 1815
rect 3345 1790 3350 1795
rect 3310 1785 3350 1790
rect 3430 1790 3435 1795
rect 3465 1815 3470 1820
rect 3550 1820 3590 1825
rect 3550 1815 3555 1820
rect 3465 1795 3555 1815
rect 3465 1790 3470 1795
rect 3430 1785 3470 1790
rect 3550 1790 3555 1795
rect 3585 1815 3590 1820
rect 3670 1820 3710 1825
rect 3670 1815 3675 1820
rect 3585 1795 3675 1815
rect 3585 1790 3590 1795
rect 3550 1785 3590 1790
rect 3670 1790 3675 1795
rect 3705 1790 3710 1820
rect 3670 1785 3710 1790
rect 4450 1820 4490 1825
rect 4450 1790 4455 1820
rect 4485 1815 4490 1820
rect 4570 1820 4610 1825
rect 4570 1815 4575 1820
rect 4485 1795 4575 1815
rect 4485 1790 4490 1795
rect 4450 1785 4490 1790
rect 4570 1790 4575 1795
rect 4605 1815 4610 1820
rect 4690 1820 4730 1825
rect 4690 1815 4695 1820
rect 4605 1795 4695 1815
rect 4605 1790 4610 1795
rect 4570 1785 4610 1790
rect 4690 1790 4695 1795
rect 4725 1815 4730 1820
rect 4810 1820 4850 1825
rect 4810 1815 4815 1820
rect 4725 1795 4815 1815
rect 4725 1790 4730 1795
rect 4690 1785 4730 1790
rect 4810 1790 4815 1795
rect 4845 1815 4850 1820
rect 4930 1820 4970 1825
rect 4930 1815 4935 1820
rect 4845 1795 4935 1815
rect 4845 1790 4850 1795
rect 4810 1785 4850 1790
rect 4930 1790 4935 1795
rect 4965 1815 4970 1820
rect 5230 1820 5270 1825
rect 5230 1815 5235 1820
rect 4965 1795 5235 1815
rect 4965 1790 4970 1795
rect 4930 1785 4970 1790
rect 5230 1790 5235 1795
rect 5265 1790 5270 1820
rect 5230 1785 5270 1790
rect -110 1720 -70 1725
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 1685 -70 1690
rect -45 1720 -5 1725
rect -45 1690 -40 1720
rect -10 1690 -5 1720
rect 2980 1720 3020 1725
rect -45 1685 -5 1690
rect 1262 1710 1302 1715
rect 1262 1680 1270 1710
rect 1297 1705 1302 1710
rect 2330 1710 2370 1715
rect 2330 1705 2335 1710
rect 1297 1685 2335 1705
rect 1297 1680 1302 1685
rect 1262 1675 1302 1680
rect 2330 1680 2335 1685
rect 2365 1680 2370 1710
rect 2980 1690 2985 1720
rect 3015 1715 3020 1720
rect 3100 1720 3140 1725
rect 3100 1715 3105 1720
rect 3015 1695 3105 1715
rect 3015 1690 3020 1695
rect 2980 1685 3020 1690
rect 3100 1690 3105 1695
rect 3135 1715 3140 1720
rect 3220 1720 3260 1725
rect 3220 1715 3225 1720
rect 3135 1695 3225 1715
rect 3135 1690 3140 1695
rect 3100 1685 3140 1690
rect 3220 1690 3225 1695
rect 3255 1715 3260 1720
rect 3340 1720 3380 1725
rect 3340 1715 3345 1720
rect 3255 1695 3345 1715
rect 3255 1690 3260 1695
rect 3220 1685 3260 1690
rect 3340 1690 3345 1695
rect 3375 1715 3380 1720
rect 3580 1720 3620 1725
rect 3580 1715 3585 1720
rect 3375 1695 3585 1715
rect 3375 1690 3380 1695
rect 3340 1685 3380 1690
rect 3580 1690 3585 1695
rect 3615 1715 3620 1720
rect 3700 1720 3740 1725
rect 3700 1715 3705 1720
rect 3615 1695 3705 1715
rect 3615 1690 3620 1695
rect 3580 1685 3620 1690
rect 3700 1690 3705 1695
rect 3735 1715 3740 1720
rect 3820 1720 3860 1725
rect 3820 1715 3825 1720
rect 3735 1695 3825 1715
rect 3735 1690 3740 1695
rect 3700 1685 3740 1690
rect 3820 1690 3825 1695
rect 3855 1715 3860 1720
rect 4300 1720 4340 1725
rect 4300 1715 4305 1720
rect 3855 1695 4305 1715
rect 3855 1690 3860 1695
rect 3820 1685 3860 1690
rect 4300 1690 4305 1695
rect 4335 1715 4340 1720
rect 4420 1720 4460 1725
rect 4420 1715 4425 1720
rect 4335 1695 4425 1715
rect 4335 1690 4340 1695
rect 4300 1685 4340 1690
rect 4420 1690 4425 1695
rect 4455 1715 4460 1720
rect 4540 1720 4580 1725
rect 4540 1715 4545 1720
rect 4455 1695 4545 1715
rect 4455 1690 4460 1695
rect 4420 1685 4460 1690
rect 4540 1690 4545 1695
rect 4575 1715 4580 1720
rect 4780 1720 4820 1725
rect 4780 1715 4785 1720
rect 4575 1695 4785 1715
rect 4575 1690 4580 1695
rect 4540 1685 4580 1690
rect 4780 1690 4785 1695
rect 4815 1715 4820 1720
rect 4900 1720 4940 1725
rect 4900 1715 4905 1720
rect 4815 1695 4905 1715
rect 4815 1690 4820 1695
rect 4780 1685 4820 1690
rect 4900 1690 4905 1695
rect 4935 1715 4940 1720
rect 5020 1720 5060 1725
rect 5020 1715 5025 1720
rect 4935 1695 5025 1715
rect 4935 1690 4940 1695
rect 4900 1685 4940 1690
rect 5020 1690 5025 1695
rect 5055 1715 5060 1720
rect 5140 1720 5180 1725
rect 5140 1715 5145 1720
rect 5055 1695 5145 1715
rect 5055 1690 5060 1695
rect 5020 1685 5060 1690
rect 5140 1690 5145 1695
rect 5175 1715 5180 1720
rect 5750 1720 5790 1725
rect 5750 1715 5755 1720
rect 5175 1695 5755 1715
rect 5175 1690 5180 1695
rect 5140 1685 5180 1690
rect 5750 1690 5755 1695
rect 5785 1690 5790 1720
rect 5750 1685 5790 1690
rect 2330 1675 2370 1680
rect 3430 1405 3470 1410
rect 3430 1375 3435 1405
rect 3465 1400 3470 1405
rect 4060 1405 4100 1410
rect 4060 1400 4065 1405
rect 3465 1380 4065 1400
rect 3465 1375 3470 1380
rect 3430 1370 3470 1375
rect 4060 1375 4065 1380
rect 4095 1400 4100 1405
rect 4690 1405 4730 1410
rect 4690 1400 4695 1405
rect 4095 1380 4695 1400
rect 4095 1375 4100 1380
rect 4060 1370 4100 1375
rect 4690 1375 4695 1380
rect 4725 1400 4730 1405
rect 5665 1405 5705 1410
rect 5665 1400 5670 1405
rect 4725 1380 5670 1400
rect 4725 1375 4730 1380
rect 4690 1370 4730 1375
rect 5665 1375 5670 1380
rect 5700 1375 5705 1405
rect 5665 1370 5705 1375
rect 4060 1310 4100 1315
rect 4060 1280 4065 1310
rect 4095 1280 4100 1310
rect 4060 1275 4100 1280
rect 3020 1255 3060 1260
rect 3020 1225 3025 1255
rect 3055 1250 3060 1255
rect 3100 1255 3140 1260
rect 3100 1250 3105 1255
rect 3055 1230 3105 1250
rect 3055 1225 3060 1230
rect 3020 1220 3060 1225
rect 3100 1225 3105 1230
rect 3135 1250 3140 1255
rect 3180 1255 3220 1260
rect 3180 1250 3185 1255
rect 3135 1230 3185 1250
rect 3135 1225 3140 1230
rect 3100 1220 3140 1225
rect 3180 1225 3185 1230
rect 3215 1250 3220 1255
rect 3260 1255 3300 1260
rect 3260 1250 3265 1255
rect 3215 1230 3265 1250
rect 3215 1225 3220 1230
rect 3180 1220 3220 1225
rect 3260 1225 3265 1230
rect 3295 1250 3300 1255
rect 3340 1255 3380 1260
rect 3340 1250 3345 1255
rect 3295 1230 3345 1250
rect 3295 1225 3300 1230
rect 3260 1220 3300 1225
rect 3340 1225 3345 1230
rect 3375 1250 3380 1255
rect 3420 1255 3460 1260
rect 3420 1250 3425 1255
rect 3375 1230 3425 1250
rect 3375 1225 3380 1230
rect 3340 1220 3380 1225
rect 3420 1225 3425 1230
rect 3455 1250 3460 1255
rect 3500 1255 3540 1260
rect 3500 1250 3505 1255
rect 3455 1230 3505 1250
rect 3455 1225 3460 1230
rect 3420 1220 3460 1225
rect 3500 1225 3505 1230
rect 3535 1250 3540 1255
rect 3580 1255 3620 1260
rect 3580 1250 3585 1255
rect 3535 1230 3585 1250
rect 3535 1225 3540 1230
rect 3500 1220 3540 1225
rect 3580 1225 3585 1230
rect 3615 1250 3620 1255
rect 3660 1255 3700 1260
rect 3660 1250 3665 1255
rect 3615 1230 3665 1250
rect 3615 1225 3620 1230
rect 3580 1220 3620 1225
rect 3660 1225 3665 1230
rect 3695 1250 3700 1255
rect 3740 1255 3780 1260
rect 3740 1250 3745 1255
rect 3695 1230 3745 1250
rect 3695 1225 3700 1230
rect 3660 1220 3700 1225
rect 3740 1225 3745 1230
rect 3775 1250 3780 1255
rect 3820 1255 3860 1260
rect 3820 1250 3825 1255
rect 3775 1230 3825 1250
rect 3775 1225 3780 1230
rect 3740 1220 3780 1225
rect 3820 1225 3825 1230
rect 3855 1250 3860 1255
rect 3900 1255 3940 1260
rect 3900 1250 3905 1255
rect 3855 1230 3905 1250
rect 3855 1225 3860 1230
rect 3820 1220 3860 1225
rect 3900 1225 3905 1230
rect 3935 1250 3940 1255
rect 3980 1255 4020 1260
rect 3980 1250 3985 1255
rect 3935 1230 3985 1250
rect 3935 1225 3940 1230
rect 3900 1220 3940 1225
rect 3980 1225 3985 1230
rect 4015 1225 4020 1255
rect 3980 1220 4020 1225
rect 4060 1255 4100 1260
rect 4060 1225 4065 1255
rect 4095 1250 4100 1255
rect 4140 1255 4180 1260
rect 4140 1250 4145 1255
rect 4095 1230 4145 1250
rect 4095 1225 4100 1230
rect 4060 1220 4100 1225
rect 4140 1225 4145 1230
rect 4175 1250 4180 1255
rect 4220 1255 4260 1260
rect 4220 1250 4225 1255
rect 4175 1230 4225 1250
rect 4175 1225 4180 1230
rect 4140 1220 4180 1225
rect 4220 1225 4225 1230
rect 4255 1250 4260 1255
rect 4300 1255 4340 1260
rect 4300 1250 4305 1255
rect 4255 1230 4305 1250
rect 4255 1225 4260 1230
rect 4220 1220 4260 1225
rect 4300 1225 4305 1230
rect 4335 1250 4340 1255
rect 4380 1255 4420 1260
rect 4380 1250 4385 1255
rect 4335 1230 4385 1250
rect 4335 1225 4340 1230
rect 4300 1220 4340 1225
rect 4380 1225 4385 1230
rect 4415 1250 4420 1255
rect 4460 1255 4500 1260
rect 4460 1250 4465 1255
rect 4415 1230 4465 1250
rect 4415 1225 4420 1230
rect 4380 1220 4420 1225
rect 4460 1225 4465 1230
rect 4495 1250 4500 1255
rect 4540 1255 4580 1260
rect 4540 1250 4545 1255
rect 4495 1230 4545 1250
rect 4495 1225 4500 1230
rect 4460 1220 4500 1225
rect 4540 1225 4545 1230
rect 4575 1250 4580 1255
rect 4620 1255 4660 1260
rect 4620 1250 4625 1255
rect 4575 1230 4625 1250
rect 4575 1225 4580 1230
rect 4540 1220 4580 1225
rect 4620 1225 4625 1230
rect 4655 1250 4660 1255
rect 4700 1255 4740 1260
rect 4700 1250 4705 1255
rect 4655 1230 4705 1250
rect 4655 1225 4660 1230
rect 4620 1220 4660 1225
rect 4700 1225 4705 1230
rect 4735 1250 4740 1255
rect 4780 1255 4820 1260
rect 4780 1250 4785 1255
rect 4735 1230 4785 1250
rect 4735 1225 4740 1230
rect 4700 1220 4740 1225
rect 4780 1225 4785 1230
rect 4815 1250 4820 1255
rect 4860 1255 4900 1260
rect 4860 1250 4865 1255
rect 4815 1230 4865 1250
rect 4815 1225 4820 1230
rect 4780 1220 4820 1225
rect 4860 1225 4865 1230
rect 4895 1250 4900 1255
rect 4940 1255 4980 1260
rect 4940 1250 4945 1255
rect 4895 1230 4945 1250
rect 4895 1225 4900 1230
rect 4860 1220 4900 1225
rect 4940 1225 4945 1230
rect 4975 1250 4980 1255
rect 5020 1255 5060 1260
rect 5020 1250 5025 1255
rect 4975 1230 5025 1250
rect 4975 1225 4980 1230
rect 4940 1220 4980 1225
rect 5020 1225 5025 1230
rect 5055 1225 5060 1255
rect 5020 1220 5060 1225
rect 2275 1170 2315 1175
rect 2275 1140 2280 1170
rect 2310 1165 2315 1170
rect 2980 1170 3020 1175
rect 2980 1165 2985 1170
rect 2310 1145 2985 1165
rect 2310 1140 2315 1145
rect 2275 1135 2315 1140
rect 2980 1140 2985 1145
rect 3015 1140 3020 1170
rect 2980 1135 3020 1140
rect 5135 1170 5175 1175
rect 5135 1140 5140 1170
rect 5170 1165 5175 1170
rect 5665 1170 5705 1175
rect 5665 1165 5670 1170
rect 5170 1145 5670 1165
rect 5170 1140 5175 1145
rect 5135 1135 5175 1140
rect 5665 1140 5670 1145
rect 5700 1140 5705 1170
rect 5665 1135 5705 1140
rect 3390 1050 3430 1055
rect 3390 1020 3395 1050
rect 3425 1045 3430 1050
rect 4060 1050 4100 1055
rect 4060 1045 4065 1050
rect 3425 1025 4065 1045
rect 3425 1020 3430 1025
rect 3390 1015 3430 1020
rect 4060 1020 4065 1025
rect 4095 1045 4100 1050
rect 4730 1050 4770 1055
rect 4730 1045 4735 1050
rect 4095 1025 4735 1045
rect 4095 1020 4100 1025
rect 4060 1015 4100 1020
rect 4730 1020 4735 1025
rect 4765 1020 4770 1050
rect 4730 1015 4770 1020
rect 3225 980 3265 985
rect 3225 950 3230 980
rect 3260 975 3265 980
rect 3335 980 3375 985
rect 3335 975 3340 980
rect 3260 955 3340 975
rect 3260 950 3265 955
rect 3225 945 3265 950
rect 3335 950 3340 955
rect 3370 975 3375 980
rect 3445 980 3485 985
rect 3445 975 3450 980
rect 3370 955 3450 975
rect 3370 950 3375 955
rect 3335 945 3375 950
rect 3445 950 3450 955
rect 3480 975 3485 980
rect 3895 980 3935 985
rect 3895 975 3900 980
rect 3480 955 3900 975
rect 3480 950 3485 955
rect 3445 945 3485 950
rect 3895 950 3900 955
rect 3930 975 3935 980
rect 4005 980 4045 985
rect 4005 975 4010 980
rect 3930 955 4010 975
rect 3930 950 3935 955
rect 3895 945 3935 950
rect 4005 950 4010 955
rect 4040 975 4045 980
rect 4115 980 4155 985
rect 4115 975 4120 980
rect 4040 955 4120 975
rect 4040 950 4045 955
rect 4005 945 4045 950
rect 4115 950 4120 955
rect 4150 975 4155 980
rect 4225 980 4265 985
rect 4225 975 4230 980
rect 4150 955 4230 975
rect 4150 950 4155 955
rect 4115 945 4155 950
rect 4225 950 4230 955
rect 4260 975 4265 980
rect 4675 980 4715 985
rect 4675 975 4680 980
rect 4260 955 4680 975
rect 4260 950 4265 955
rect 4225 945 4265 950
rect 4675 950 4680 955
rect 4710 975 4715 980
rect 4785 980 4825 985
rect 4785 975 4790 980
rect 4710 955 4790 975
rect 4710 950 4715 955
rect 4675 945 4715 950
rect 4785 950 4790 955
rect 4820 975 4825 980
rect 4895 980 4935 985
rect 4895 975 4900 980
rect 4820 955 4900 975
rect 4820 950 4825 955
rect 4785 945 4825 950
rect 4895 950 4900 955
rect 4930 975 4935 980
rect 5665 980 5705 985
rect 5665 975 5670 980
rect 4930 955 5670 975
rect 4930 950 4935 955
rect 4895 945 4935 950
rect 5665 950 5670 955
rect 5700 950 5705 980
rect 5665 945 5705 950
rect 3670 895 3710 900
rect 3670 865 3675 895
rect 3705 890 3710 895
rect 3725 895 3765 900
rect 3725 890 3730 895
rect 3705 870 3730 890
rect 3705 865 3710 870
rect 3670 860 3710 865
rect 3725 865 3730 870
rect 3760 865 3765 895
rect 3725 860 3765 865
rect 4395 895 4435 900
rect 4395 865 4400 895
rect 4430 890 4435 895
rect 4450 895 4490 900
rect 4450 890 4455 895
rect 4430 870 4455 890
rect 4430 865 4435 870
rect 4395 860 4435 865
rect 4450 865 4455 870
rect 4485 865 4490 895
rect 4450 860 4490 865
rect 5065 895 5105 900
rect 5065 865 5070 895
rect 5100 890 5105 895
rect 5665 895 5705 900
rect 5665 890 5670 895
rect 5100 870 5670 890
rect 5100 865 5105 870
rect 5065 860 5105 865
rect 5665 865 5670 870
rect 5700 865 5705 895
rect 5665 860 5705 865
rect 3170 810 3210 815
rect 3170 780 3175 810
rect 3205 805 3210 810
rect 3390 810 3430 815
rect 3390 805 3395 810
rect 3205 785 3395 805
rect 3205 780 3210 785
rect 3170 775 3210 780
rect 3390 780 3395 785
rect 3425 780 3430 810
rect 3390 775 3430 780
rect 4060 810 4100 815
rect 4060 780 4065 810
rect 4095 805 4100 810
rect 4170 810 4210 815
rect 4170 805 4175 810
rect 4095 785 4175 805
rect 4095 780 4100 785
rect 4060 775 4100 780
rect 4170 780 4175 785
rect 4205 805 4210 810
rect 4280 810 4320 815
rect 4280 805 4285 810
rect 4205 785 4285 805
rect 4205 780 4210 785
rect 4170 775 4210 780
rect 4280 780 4285 785
rect 4315 780 4320 810
rect 4280 775 4320 780
rect 4730 810 4770 815
rect 4730 780 4735 810
rect 4765 805 4770 810
rect 4950 810 4990 815
rect 4950 805 4955 810
rect 4765 785 4955 805
rect 4765 780 4770 785
rect 4730 775 4770 780
rect 4950 780 4955 785
rect 4985 780 4990 810
rect 4950 775 4990 780
rect 3280 755 3320 760
rect 3280 725 3285 755
rect 3315 750 3320 755
rect 3500 755 3540 760
rect 3500 750 3505 755
rect 3315 730 3505 750
rect 3315 725 3320 730
rect 3280 720 3320 725
rect 3500 725 3505 730
rect 3535 750 3540 755
rect 4060 755 4100 760
rect 4060 750 4065 755
rect 3535 730 4065 750
rect 3535 725 3540 730
rect 3500 720 3540 725
rect 4060 725 4065 730
rect 4095 750 4100 755
rect 4620 755 4660 760
rect 4620 750 4625 755
rect 4095 730 4625 750
rect 4095 725 4100 730
rect 4060 720 4100 725
rect 4620 725 4625 730
rect 4655 750 4660 755
rect 4840 755 4880 760
rect 4840 750 4845 755
rect 4655 730 4845 750
rect 4655 725 4660 730
rect 4620 720 4660 725
rect 4840 725 4845 730
rect 4875 725 4880 755
rect 4840 720 4880 725
rect 2555 710 2595 715
rect 2555 680 2560 710
rect 2590 705 2595 710
rect 3865 710 3905 715
rect 3865 705 3870 710
rect 2590 685 3870 705
rect 2590 680 2595 685
rect 2555 675 2595 680
rect 3865 680 3870 685
rect 3900 680 3905 710
rect 3865 675 3905 680
rect -195 575 -155 580
rect -195 545 -190 575
rect -160 545 -155 575
rect -195 540 -155 545
<< via2 >>
rect -190 5310 -160 5340
rect 5755 5310 5785 5340
rect -105 3845 -75 3875
rect 4445 3815 4475 3845
rect 5755 3815 5785 3845
rect 945 3765 975 3795
rect 1645 3765 1675 3795
rect 5145 3765 5175 3795
rect 2695 3710 2725 3740
rect 3395 3710 3425 3740
rect -105 3495 -75 3525
rect 5755 3500 5785 3530
rect -105 3230 -75 3260
rect -105 3165 -75 3195
rect 5755 3035 5785 3065
rect 5755 2405 5785 2435
rect -105 1690 -75 1720
rect 5755 1690 5785 1720
rect 5670 1375 5700 1405
rect 5670 1140 5700 1170
rect 5670 950 5700 980
rect 5670 865 5700 895
rect -190 545 -160 575
<< metal3 >>
rect -200 5345 -150 5350
rect -200 5305 -195 5345
rect -155 5305 -150 5345
rect -200 5300 -150 5305
rect 5745 5345 5795 5350
rect 5745 5305 5750 5345
rect 5790 5305 5795 5345
rect 5745 5300 5795 5305
rect -195 585 -155 5300
rect -115 5260 -65 5265
rect -115 5220 -110 5260
rect -70 5220 -65 5260
rect -115 5215 -65 5220
rect 5660 5260 5710 5265
rect 5660 5220 5665 5260
rect 5705 5220 5710 5260
rect 5660 5215 5710 5220
rect -110 3875 -70 5215
rect 145 5120 375 5205
rect 495 5120 725 5205
rect 845 5120 1075 5205
rect 1195 5120 1425 5205
rect 1545 5120 1775 5205
rect 145 5070 1775 5120
rect 145 4975 375 5070
rect 495 4975 725 5070
rect 845 4975 1075 5070
rect 1195 4975 1425 5070
rect 1545 4975 1775 5070
rect 1895 5120 2125 5205
rect 2245 5120 2475 5205
rect 2595 5120 2825 5205
rect 2945 5120 3175 5205
rect 3295 5120 3525 5205
rect 1895 5070 3525 5120
rect 1895 4975 2125 5070
rect 2245 4975 2475 5070
rect 2595 4975 2825 5070
rect 2945 4975 3175 5070
rect 3295 4975 3525 5070
rect 3645 5120 3875 5205
rect 3995 5120 4225 5205
rect 4345 5120 4575 5205
rect 4695 5120 4925 5205
rect 5045 5120 5275 5205
rect 3645 5070 5275 5120
rect 3645 4975 3875 5070
rect 3995 4975 4225 5070
rect 4345 4975 4575 5070
rect 4695 4975 4925 5070
rect 5045 4975 5275 5070
rect 935 4855 985 4975
rect 2685 4855 2735 4975
rect 4435 4855 4485 4975
rect 145 4770 375 4855
rect 495 4770 725 4855
rect 845 4770 1075 4855
rect 1195 4770 1425 4855
rect 1545 4770 1775 4855
rect 145 4720 1775 4770
rect 145 4625 375 4720
rect 495 4625 725 4720
rect 845 4625 1075 4720
rect 1195 4625 1425 4720
rect 1545 4625 1775 4720
rect 1895 4770 2125 4855
rect 2245 4770 2475 4855
rect 2595 4770 2825 4855
rect 2945 4770 3175 4855
rect 3295 4770 3525 4855
rect 1895 4720 3525 4770
rect 1895 4625 2125 4720
rect 2245 4625 2475 4720
rect 2595 4625 2825 4720
rect 2945 4625 3175 4720
rect 3295 4625 3525 4720
rect 3645 4770 3875 4855
rect 3995 4770 4225 4855
rect 4345 4770 4575 4855
rect 4695 4770 4925 4855
rect 5045 4770 5275 4855
rect 3645 4720 5275 4770
rect 3645 4625 3875 4720
rect 3995 4625 4225 4720
rect 4345 4625 4575 4720
rect 4695 4625 4925 4720
rect 5045 4625 5275 4720
rect 935 4505 985 4625
rect 2685 4505 2735 4625
rect 4435 4505 4485 4625
rect 145 4420 375 4505
rect 495 4420 725 4505
rect 845 4420 1075 4505
rect 1195 4420 1425 4505
rect 1545 4420 1775 4505
rect 145 4370 1775 4420
rect 145 4275 375 4370
rect 495 4275 725 4370
rect 845 4275 1075 4370
rect 1195 4275 1425 4370
rect 1545 4275 1775 4370
rect 1895 4420 2125 4505
rect 2245 4420 2475 4505
rect 2595 4420 2825 4505
rect 2945 4420 3175 4505
rect 3295 4420 3525 4505
rect 1895 4370 3525 4420
rect 1895 4275 2125 4370
rect 2245 4275 2475 4370
rect 2595 4275 2825 4370
rect 2945 4275 3175 4370
rect 3295 4275 3525 4370
rect 3645 4420 3875 4505
rect 3995 4420 4225 4505
rect 4345 4420 4575 4505
rect 4695 4420 4925 4505
rect 5045 4420 5275 4505
rect 3645 4370 5275 4420
rect 3645 4275 3875 4370
rect 3995 4275 4225 4370
rect 4345 4275 4575 4370
rect 4695 4275 4925 4370
rect 5045 4275 5275 4370
rect 935 4155 985 4275
rect 2685 4155 2735 4275
rect 4435 4155 4485 4275
rect 145 4070 375 4155
rect 495 4070 725 4155
rect 845 4070 1075 4155
rect 1195 4070 1425 4155
rect 1545 4070 1775 4155
rect 145 4020 1775 4070
rect 145 3925 375 4020
rect 495 3925 725 4020
rect 845 3925 1075 4020
rect 1195 3925 1425 4020
rect 1545 3925 1775 4020
rect 1895 4070 2125 4155
rect 2245 4070 2475 4155
rect 2595 4070 2825 4155
rect 2945 4070 3175 4155
rect 3295 4070 3525 4155
rect 1895 4020 3525 4070
rect 1895 3925 2125 4020
rect 2245 3925 2475 4020
rect 2595 3925 2825 4020
rect 2945 3925 3175 4020
rect 3295 3925 3525 4020
rect 3645 4070 3875 4155
rect 3995 4070 4225 4155
rect 4345 4070 4575 4155
rect 4695 4070 4925 4155
rect 5045 4070 5275 4155
rect 3645 4020 5275 4070
rect 3645 3925 3875 4020
rect 3995 3925 4225 4020
rect 4345 3925 4575 4020
rect 4695 3925 4925 4020
rect 5045 3925 5275 4020
rect -110 3845 -105 3875
rect -75 3845 -70 3875
rect -110 3525 -70 3845
rect 940 3795 980 3925
rect 940 3765 945 3795
rect 975 3765 980 3795
rect 940 3760 980 3765
rect 1635 3800 1685 3805
rect 1635 3760 1640 3800
rect 1680 3760 1685 3800
rect 1635 3755 1685 3760
rect 2690 3740 2730 3925
rect 4440 3845 4480 3925
rect 4440 3815 4445 3845
rect 4475 3815 4480 3845
rect 4440 3810 4480 3815
rect 5135 3800 5185 3805
rect 5135 3760 5140 3800
rect 5180 3760 5185 3800
rect 5135 3755 5185 3760
rect 2690 3710 2695 3740
rect 2725 3710 2730 3740
rect 2690 3705 2730 3710
rect 3385 3745 3435 3750
rect 3385 3705 3390 3745
rect 3430 3705 3435 3745
rect 3385 3700 3435 3705
rect -110 3495 -105 3525
rect -75 3495 -70 3525
rect -110 3260 -70 3495
rect -110 3230 -105 3260
rect -75 3230 -70 3260
rect -110 3195 -70 3230
rect -110 3165 -105 3195
rect -75 3165 -70 3195
rect -110 1720 -70 3165
rect -110 1690 -105 1720
rect -75 1690 -70 1720
rect -110 665 -70 1690
rect 5665 1405 5705 5215
rect 5665 1375 5670 1405
rect 5700 1375 5705 1405
rect 5665 1170 5705 1375
rect 5665 1140 5670 1170
rect 5700 1140 5705 1170
rect 5665 980 5705 1140
rect 5665 950 5670 980
rect 5700 950 5705 980
rect 5665 895 5705 950
rect 5665 865 5670 895
rect 5700 865 5705 895
rect 5665 665 5705 865
rect 5750 3845 5790 5300
rect 5750 3815 5755 3845
rect 5785 3815 5790 3845
rect 5750 3530 5790 3815
rect 5750 3500 5755 3530
rect 5785 3500 5790 3530
rect 5750 3065 5790 3500
rect 5750 3035 5755 3065
rect 5785 3035 5790 3065
rect 5750 2435 5790 3035
rect 5750 2405 5755 2435
rect 5785 2405 5790 2435
rect 5750 1720 5790 2405
rect 5750 1690 5755 1720
rect 5785 1690 5790 1720
rect -115 660 -65 665
rect -115 620 -110 660
rect -70 620 -65 660
rect -115 615 -65 620
rect 5660 660 5710 665
rect 5660 620 5665 660
rect 5705 620 5710 660
rect 5660 615 5710 620
rect 5750 585 5790 1690
rect -200 580 -150 585
rect -200 540 -195 580
rect -155 540 -150 580
rect -200 535 -150 540
rect 5745 580 5795 585
rect 5745 540 5750 580
rect 5790 540 5795 580
rect 5745 535 5795 540
<< via3 >>
rect -195 5340 -155 5345
rect -195 5310 -190 5340
rect -190 5310 -160 5340
rect -160 5310 -155 5340
rect -195 5305 -155 5310
rect 5750 5340 5790 5345
rect 5750 5310 5755 5340
rect 5755 5310 5785 5340
rect 5785 5310 5790 5340
rect 5750 5305 5790 5310
rect -110 5220 -70 5260
rect 5665 5220 5705 5260
rect 1640 3795 1680 3800
rect 1640 3765 1645 3795
rect 1645 3765 1675 3795
rect 1675 3765 1680 3795
rect 1640 3760 1680 3765
rect 5140 3795 5180 3800
rect 5140 3765 5145 3795
rect 5145 3765 5175 3795
rect 5175 3765 5180 3795
rect 5140 3760 5180 3765
rect 3390 3740 3430 3745
rect 3390 3710 3395 3740
rect 3395 3710 3425 3740
rect 3425 3710 3430 3740
rect 3390 3705 3430 3710
rect -110 620 -70 660
rect 5665 620 5705 660
rect -195 575 -155 580
rect -195 545 -190 575
rect -190 545 -160 575
rect -160 545 -155 575
rect -195 540 -155 545
rect 5750 540 5790 580
<< mimcap >>
rect 160 5115 360 5190
rect 160 5075 240 5115
rect 280 5075 360 5115
rect 160 4990 360 5075
rect 510 5115 710 5190
rect 510 5075 590 5115
rect 630 5075 710 5115
rect 510 4990 710 5075
rect 860 5115 1060 5190
rect 860 5075 940 5115
rect 980 5075 1060 5115
rect 860 4990 1060 5075
rect 1210 5115 1410 5190
rect 1210 5075 1290 5115
rect 1330 5075 1410 5115
rect 1210 4990 1410 5075
rect 1560 5115 1760 5190
rect 1560 5075 1640 5115
rect 1680 5075 1760 5115
rect 1560 4990 1760 5075
rect 1910 5115 2110 5190
rect 1910 5075 1990 5115
rect 2030 5075 2110 5115
rect 1910 4990 2110 5075
rect 2260 5115 2460 5190
rect 2260 5075 2340 5115
rect 2380 5075 2460 5115
rect 2260 4990 2460 5075
rect 2610 5115 2810 5190
rect 2610 5075 2690 5115
rect 2730 5075 2810 5115
rect 2610 4990 2810 5075
rect 2960 5115 3160 5190
rect 2960 5075 3040 5115
rect 3080 5075 3160 5115
rect 2960 4990 3160 5075
rect 3310 5115 3510 5190
rect 3310 5075 3390 5115
rect 3430 5075 3510 5115
rect 3310 4990 3510 5075
rect 3660 5115 3860 5190
rect 3660 5075 3740 5115
rect 3780 5075 3860 5115
rect 3660 4990 3860 5075
rect 4010 5115 4210 5190
rect 4010 5075 4090 5115
rect 4130 5075 4210 5115
rect 4010 4990 4210 5075
rect 4360 5115 4560 5190
rect 4360 5075 4440 5115
rect 4480 5075 4560 5115
rect 4360 4990 4560 5075
rect 4710 5115 4910 5190
rect 4710 5075 4790 5115
rect 4830 5075 4910 5115
rect 4710 4990 4910 5075
rect 5060 5115 5260 5190
rect 5060 5075 5140 5115
rect 5180 5075 5260 5115
rect 5060 4990 5260 5075
rect 160 4765 360 4840
rect 160 4725 240 4765
rect 280 4725 360 4765
rect 160 4640 360 4725
rect 510 4765 710 4840
rect 510 4725 590 4765
rect 630 4725 710 4765
rect 510 4640 710 4725
rect 860 4765 1060 4840
rect 860 4725 940 4765
rect 980 4725 1060 4765
rect 860 4640 1060 4725
rect 1210 4765 1410 4840
rect 1210 4725 1290 4765
rect 1330 4725 1410 4765
rect 1210 4640 1410 4725
rect 1560 4765 1760 4840
rect 1560 4725 1640 4765
rect 1680 4725 1760 4765
rect 1560 4640 1760 4725
rect 1910 4765 2110 4840
rect 1910 4725 1990 4765
rect 2030 4725 2110 4765
rect 1910 4640 2110 4725
rect 2260 4765 2460 4840
rect 2260 4725 2340 4765
rect 2380 4725 2460 4765
rect 2260 4640 2460 4725
rect 2610 4765 2810 4840
rect 2610 4725 2690 4765
rect 2730 4725 2810 4765
rect 2610 4640 2810 4725
rect 2960 4765 3160 4840
rect 2960 4725 3040 4765
rect 3080 4725 3160 4765
rect 2960 4640 3160 4725
rect 3310 4765 3510 4840
rect 3310 4725 3390 4765
rect 3430 4725 3510 4765
rect 3310 4640 3510 4725
rect 3660 4765 3860 4840
rect 3660 4725 3740 4765
rect 3780 4725 3860 4765
rect 3660 4640 3860 4725
rect 4010 4765 4210 4840
rect 4010 4725 4090 4765
rect 4130 4725 4210 4765
rect 4010 4640 4210 4725
rect 4360 4765 4560 4840
rect 4360 4725 4440 4765
rect 4480 4725 4560 4765
rect 4360 4640 4560 4725
rect 4710 4765 4910 4840
rect 4710 4725 4790 4765
rect 4830 4725 4910 4765
rect 4710 4640 4910 4725
rect 5060 4765 5260 4840
rect 5060 4725 5140 4765
rect 5180 4725 5260 4765
rect 5060 4640 5260 4725
rect 160 4415 360 4490
rect 160 4375 240 4415
rect 280 4375 360 4415
rect 160 4290 360 4375
rect 510 4415 710 4490
rect 510 4375 590 4415
rect 630 4375 710 4415
rect 510 4290 710 4375
rect 860 4415 1060 4490
rect 860 4375 940 4415
rect 980 4375 1060 4415
rect 860 4290 1060 4375
rect 1210 4415 1410 4490
rect 1210 4375 1290 4415
rect 1330 4375 1410 4415
rect 1210 4290 1410 4375
rect 1560 4415 1760 4490
rect 1560 4375 1640 4415
rect 1680 4375 1760 4415
rect 1560 4290 1760 4375
rect 1910 4415 2110 4490
rect 1910 4375 1990 4415
rect 2030 4375 2110 4415
rect 1910 4290 2110 4375
rect 2260 4415 2460 4490
rect 2260 4375 2340 4415
rect 2380 4375 2460 4415
rect 2260 4290 2460 4375
rect 2610 4415 2810 4490
rect 2610 4375 2690 4415
rect 2730 4375 2810 4415
rect 2610 4290 2810 4375
rect 2960 4415 3160 4490
rect 2960 4375 3040 4415
rect 3080 4375 3160 4415
rect 2960 4290 3160 4375
rect 3310 4415 3510 4490
rect 3310 4375 3390 4415
rect 3430 4375 3510 4415
rect 3310 4290 3510 4375
rect 3660 4415 3860 4490
rect 3660 4375 3740 4415
rect 3780 4375 3860 4415
rect 3660 4290 3860 4375
rect 4010 4415 4210 4490
rect 4010 4375 4090 4415
rect 4130 4375 4210 4415
rect 4010 4290 4210 4375
rect 4360 4415 4560 4490
rect 4360 4375 4440 4415
rect 4480 4375 4560 4415
rect 4360 4290 4560 4375
rect 4710 4415 4910 4490
rect 4710 4375 4790 4415
rect 4830 4375 4910 4415
rect 4710 4290 4910 4375
rect 5060 4415 5260 4490
rect 5060 4375 5140 4415
rect 5180 4375 5260 4415
rect 5060 4290 5260 4375
rect 160 4065 360 4140
rect 160 4025 240 4065
rect 280 4025 360 4065
rect 160 3940 360 4025
rect 510 4065 710 4140
rect 510 4025 590 4065
rect 630 4025 710 4065
rect 510 3940 710 4025
rect 860 4065 1060 4140
rect 860 4025 940 4065
rect 980 4025 1060 4065
rect 860 3940 1060 4025
rect 1210 4065 1410 4140
rect 1210 4025 1290 4065
rect 1330 4025 1410 4065
rect 1210 3940 1410 4025
rect 1560 4065 1760 4140
rect 1560 4025 1640 4065
rect 1680 4025 1760 4065
rect 1560 3940 1760 4025
rect 1910 4065 2110 4140
rect 1910 4025 1990 4065
rect 2030 4025 2110 4065
rect 1910 3940 2110 4025
rect 2260 4065 2460 4140
rect 2260 4025 2340 4065
rect 2380 4025 2460 4065
rect 2260 3940 2460 4025
rect 2610 4065 2810 4140
rect 2610 4025 2690 4065
rect 2730 4025 2810 4065
rect 2610 3940 2810 4025
rect 2960 4065 3160 4140
rect 2960 4025 3040 4065
rect 3080 4025 3160 4065
rect 2960 3940 3160 4025
rect 3310 4065 3510 4140
rect 3310 4025 3390 4065
rect 3430 4025 3510 4065
rect 3310 3940 3510 4025
rect 3660 4065 3860 4140
rect 3660 4025 3740 4065
rect 3780 4025 3860 4065
rect 3660 3940 3860 4025
rect 4010 4065 4210 4140
rect 4010 4025 4090 4065
rect 4130 4025 4210 4065
rect 4010 3940 4210 4025
rect 4360 4065 4560 4140
rect 4360 4025 4440 4065
rect 4480 4025 4560 4065
rect 4360 3940 4560 4025
rect 4710 4065 4910 4140
rect 4710 4025 4790 4065
rect 4830 4025 4910 4065
rect 4710 3940 4910 4025
rect 5060 4065 5260 4140
rect 5060 4025 5140 4065
rect 5180 4025 5260 4065
rect 5060 3940 5260 4025
<< mimcapcontact >>
rect 240 5075 280 5115
rect 590 5075 630 5115
rect 940 5075 980 5115
rect 1290 5075 1330 5115
rect 1640 5075 1680 5115
rect 1990 5075 2030 5115
rect 2340 5075 2380 5115
rect 2690 5075 2730 5115
rect 3040 5075 3080 5115
rect 3390 5075 3430 5115
rect 3740 5075 3780 5115
rect 4090 5075 4130 5115
rect 4440 5075 4480 5115
rect 4790 5075 4830 5115
rect 5140 5075 5180 5115
rect 240 4725 280 4765
rect 590 4725 630 4765
rect 940 4725 980 4765
rect 1290 4725 1330 4765
rect 1640 4725 1680 4765
rect 1990 4725 2030 4765
rect 2340 4725 2380 4765
rect 2690 4725 2730 4765
rect 3040 4725 3080 4765
rect 3390 4725 3430 4765
rect 3740 4725 3780 4765
rect 4090 4725 4130 4765
rect 4440 4725 4480 4765
rect 4790 4725 4830 4765
rect 5140 4725 5180 4765
rect 240 4375 280 4415
rect 590 4375 630 4415
rect 940 4375 980 4415
rect 1290 4375 1330 4415
rect 1640 4375 1680 4415
rect 1990 4375 2030 4415
rect 2340 4375 2380 4415
rect 2690 4375 2730 4415
rect 3040 4375 3080 4415
rect 3390 4375 3430 4415
rect 3740 4375 3780 4415
rect 4090 4375 4130 4415
rect 4440 4375 4480 4415
rect 4790 4375 4830 4415
rect 5140 4375 5180 4415
rect 240 4025 280 4065
rect 590 4025 630 4065
rect 940 4025 980 4065
rect 1290 4025 1330 4065
rect 1640 4025 1680 4065
rect 1990 4025 2030 4065
rect 2340 4025 2380 4065
rect 2690 4025 2730 4065
rect 3040 4025 3080 4065
rect 3390 4025 3430 4065
rect 3740 4025 3780 4065
rect 4090 4025 4130 4065
rect 4440 4025 4480 4065
rect 4790 4025 4830 4065
rect 5140 4025 5180 4065
<< metal4 >>
rect -200 5345 5795 5350
rect -200 5305 -195 5345
rect -155 5305 5750 5345
rect 5790 5305 5795 5345
rect -200 5300 5795 5305
rect -115 5260 5710 5265
rect -115 5220 -110 5260
rect -70 5220 5665 5260
rect 5705 5220 5710 5260
rect -115 5215 5710 5220
rect 235 5115 1685 5120
rect 235 5075 240 5115
rect 280 5075 590 5115
rect 630 5075 940 5115
rect 980 5075 1290 5115
rect 1330 5075 1640 5115
rect 1680 5075 1685 5115
rect 235 5070 1685 5075
rect 1985 5115 3435 5120
rect 1985 5075 1990 5115
rect 2030 5075 2340 5115
rect 2380 5075 2690 5115
rect 2730 5075 3040 5115
rect 3080 5075 3390 5115
rect 3430 5075 3435 5115
rect 1985 5070 3435 5075
rect 3735 5115 5185 5120
rect 3735 5075 3740 5115
rect 3780 5075 4090 5115
rect 4130 5075 4440 5115
rect 4480 5075 4790 5115
rect 4830 5075 5140 5115
rect 5180 5075 5185 5115
rect 3735 5070 5185 5075
rect 935 4770 985 5070
rect 2685 4770 2735 5070
rect 4435 4770 4485 5070
rect 235 4765 1685 4770
rect 235 4725 240 4765
rect 280 4725 590 4765
rect 630 4725 940 4765
rect 980 4725 1290 4765
rect 1330 4725 1640 4765
rect 1680 4725 1685 4765
rect 235 4720 1685 4725
rect 1985 4765 3435 4770
rect 1985 4725 1990 4765
rect 2030 4725 2340 4765
rect 2380 4725 2690 4765
rect 2730 4725 3040 4765
rect 3080 4725 3390 4765
rect 3430 4725 3435 4765
rect 1985 4720 3435 4725
rect 3735 4765 5185 4770
rect 3735 4725 3740 4765
rect 3780 4725 4090 4765
rect 4130 4725 4440 4765
rect 4480 4725 4790 4765
rect 4830 4725 5140 4765
rect 5180 4725 5185 4765
rect 3735 4720 5185 4725
rect 935 4420 985 4720
rect 2685 4420 2735 4720
rect 4435 4420 4485 4720
rect 235 4415 1685 4420
rect 235 4375 240 4415
rect 280 4375 590 4415
rect 630 4375 940 4415
rect 980 4375 1290 4415
rect 1330 4375 1640 4415
rect 1680 4375 1685 4415
rect 235 4370 1685 4375
rect 1985 4415 3435 4420
rect 1985 4375 1990 4415
rect 2030 4375 2340 4415
rect 2380 4375 2690 4415
rect 2730 4375 3040 4415
rect 3080 4375 3390 4415
rect 3430 4375 3435 4415
rect 1985 4370 3435 4375
rect 3735 4415 5185 4420
rect 3735 4375 3740 4415
rect 3780 4375 4090 4415
rect 4130 4375 4440 4415
rect 4480 4375 4790 4415
rect 4830 4375 5140 4415
rect 5180 4375 5185 4415
rect 3735 4370 5185 4375
rect 935 4070 985 4370
rect 2685 4070 2735 4370
rect 4435 4070 4485 4370
rect 235 4065 1685 4070
rect 235 4025 240 4065
rect 280 4025 590 4065
rect 630 4025 940 4065
rect 980 4025 1290 4065
rect 1330 4025 1640 4065
rect 1680 4025 1685 4065
rect 235 4020 1685 4025
rect 1985 4065 3435 4070
rect 1985 4025 1990 4065
rect 2030 4025 2340 4065
rect 2380 4025 2690 4065
rect 2730 4025 3040 4065
rect 3080 4025 3390 4065
rect 3430 4025 3435 4065
rect 1985 4020 3435 4025
rect 3735 4065 5185 4070
rect 3735 4025 3740 4065
rect 3780 4025 4090 4065
rect 4130 4025 4440 4065
rect 4480 4025 4790 4065
rect 4830 4025 5140 4065
rect 5180 4025 5185 4065
rect 3735 4020 5185 4025
rect 1635 3800 1685 4020
rect 1635 3760 1640 3800
rect 1680 3760 1685 3800
rect 1635 3755 1685 3760
rect 3385 3745 3435 4020
rect 5135 3800 5185 4020
rect 5135 3760 5140 3800
rect 5180 3760 5185 3800
rect 5135 3755 5185 3760
rect 3385 3705 3390 3745
rect 3430 3705 3435 3745
rect 3385 3700 3435 3705
rect -115 660 5710 665
rect -115 620 -110 660
rect -70 620 5665 660
rect 5705 620 5710 660
rect -115 615 5710 620
rect -200 580 5795 585
rect -200 540 -195 580
rect -155 540 5750 580
rect 5790 540 5795 580
rect -200 535 5795 540
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_9 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 1475 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_10
timestamp 1723858470
transform 1 0 1475 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_11
timestamp 1723858470
transform 1 0 1475 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_12
timestamp 1723858470
transform 1 0 115 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_13
timestamp 1723858470
transform 1 0 115 0 1 1360
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_14
timestamp 1723858470
transform 1 0 115 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_15
timestamp 1723858470
transform 1 0 795 0 1 680
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_16
timestamp 1723858470
transform 1 0 795 0 1 2040
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_17
timestamp 1723858470
transform 1 0 795 0 1 1360
box 0 0 670 670
<< labels >>
flabel metal2 455 3790 455 3790 1 FreeSans 400 0 0 40 cap_res1
flabel metal3 2730 3725 2730 3725 3 FreeSans 400 0 40 0 cap_res2
flabel metal1 1985 2370 1985 2370 3 FreeSans 400 0 40 0 Vbe2
flabel poly 4710 2690 4710 2690 5 FreeSans 400 0 0 -40 V_TOP
flabel metal1 5060 1240 5060 1240 3 FreeSans 400 0 200 0 START_UP_NFET1
flabel metal2 5210 1875 5210 1875 1 FreeSans 400 0 0 80 V_CUR_REF_REG
flabel metal2 5260 2170 5260 2170 5 FreeSans 400 0 0 -40 V_mir2
flabel metal1 2585 995 2585 995 3 FreeSans 400 0 40 0 NFET_GATE_10uA
flabel metal1 4080 350 4080 350 5 FreeSans 400 0 0 -200 VB2_CUR_BIAS
port 5 s
flabel metal2 6100 3100 6100 3100 3 FreeSans 400 0 200 0 TAIL_CUR_MIR_BIAS
port 9 e
flabel metal2 6100 3620 6100 3620 3 FreeSans 400 0 200 0 V_CMFB_S1
port 10 e
flabel metal2 6100 2030 6100 2030 3 FreeSans 400 0 200 0 ERR_AMP_REF
port 3 e
flabel metal3 5790 4750 5790 4750 3 FreeSans 400 0 200 0 VDDA
port 4 e
flabel metal3 5705 4525 5705 4525 3 FreeSans 400 0 200 0 GNDA
port 2 e
flabel metal2 2950 1875 2950 1875 1 FreeSans 400 0 0 80 Vin+
flabel metal2 2945 2020 2945 2020 5 FreeSans 400 0 0 -80 Vin-
flabel metal1 2305 1455 2305 1455 3 FreeSans 400 0 200 0 START_UP
flabel metal2 4310 2130 4310 2130 7 FreeSans 240 0 -120 0 1st_Vout_2
flabel metal2 4450 1785 4450 1785 7 FreeSans 400 0 -200 0 V_p_2
flabel metal2 3710 1785 3710 1785 3 FreeSans 400 0 200 0 V_p_1
flabel metal2 2900 2170 2900 2170 5 FreeSans 400 0 0 -40 V_mir1
flabel metal2 3850 2130 3850 2130 3 FreeSans 240 0 120 0 1st_Vout_1
flabel metal2 6100 2780 6100 2780 3 FreeSans 400 0 200 0 VB1_CUR_BIAS
port 1 e
flabel metal2 6100 3345 6100 3345 3 FreeSans 400 0 200 0 V_CMFB_S3
port 12 e
flabel metal1 3960 385 3960 385 7 FreeSans 400 0 -200 0 ERR_AMP_CUR_BIAS
port 7 w
flabel metal1 4200 385 4200 385 3 FreeSans 400 0 200 0 VB3_CUR_BIAS
port 6 e
flabel metal1 4970 350 4970 350 5 FreeSans 400 0 0 -200 V_CMFB_S4
port 11 s
flabel metal1 3190 350 3190 350 5 FreeSans 400 0 0 -200 V_CMFB_S2
port 8 s
flabel via1 4080 3585 4080 3585 1 FreeSans 400 0 0 200 PFET_GATE_10uA
<< end >>
