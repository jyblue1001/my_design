* NGSPICE file created from charge_pump_full_4.ext - technology: sky130A

.subckt A a_540_n9930# a_2200_n8070# w_240_n9000# a_n80_n8330# a_380_n8130#
X0 w_240_n9000# a_380_n8130# a_n80_n8330# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X1 w_240_n9000# a_380_n8130# a_n80_n8330# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X2 w_240_n9000# a_1630_n9420# a_2200_n8070# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X3 w_240_n9000# a_1630_n9420# a_2200_n8070# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X4 a_1630_n9420# a_1050_n9420# a_380_n8130# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X5 a_1050_n9420# a_760_n9420# a_540_n9930# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X6 a_1340_n9420# a_1050_n9420# a_540_n9930# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X7 a_1630_n9420# a_1340_n9420# a_380_n8130# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X8 a_540_n9930# I_IN a_n80_n8330# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X9 a_n80_n8330# a_380_n8130# w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X10 a_1340_n9420# a_1050_n9420# w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X11 a_2200_n8070# a_1630_n9420# w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X12 a_1050_n9420# a_760_n9420# w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X13 a_760_n9420# UP_PFD a_540_n9930# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X14 I_IN I_IN a_540_n9930# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X15 a_2790_n9420# a_2210_n9420# a_540_n9930# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X16 a_n80_n8330# I_IN a_540_n9930# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X17 a_2200_n8070# a_2790_n9420# a_540_n9930# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X18 a_2200_n8070# a_1630_n9420# w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X19 a_760_n9420# UP_PFD w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X20 a_1630_n9420# a_1050_n9420# w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X21 a_2790_n9420# a_2500_n9420# I_IN a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X22 a_n80_n8330# I_IN a_540_n9930# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X23 w_240_n9000# a_380_n8130# a_n80_n8330# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X24 w_240_n9000# a_380_n8130# a_n80_n8330# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X25 w_240_n9000# a_1630_n9420# a_2200_n8070# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X26 a_2500_n9420# a_2210_n9420# a_540_n9930# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X27 a_2790_n9420# a_2500_n9420# sky130_fd_pr__cap_mim_m3_1 l=2.6 w=2.6
X28 a_2210_n9420# w_240_n9000# a_1790_n9420# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X29 a_2790_n9420# a_2210_n9420# I_IN w_240_n9000# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X30 a_2210_n9420# a_540_n9930# a_1790_n9420# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X31 a_2500_n9420# a_2210_n9420# w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X32 a_1630_n9420# a_1340_n9420# sky130_fd_pr__cap_mim_m3_1 l=6 w=4.2
X33 a_540_n9930# I_IN I_IN a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X34 a_540_n9930# a_2790_n9420# a_2200_n8070# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X35 a_540_n9930# a_2790_n9420# a_2200_n8070# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X36 a_n80_n8330# a_380_n8130# w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X37 a_540_n9930# DOWN_PFD a_1790_n9420# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X38 a_540_n9930# I_IN a_n80_n8330# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X39 a_2200_n8070# a_1630_n9420# w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X40 w_240_n9000# DOWN_PFD a_1790_n9420# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X41 a_n80_n8330# a_380_n8130# w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X42 I_IN I_IN a_540_n9930# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X43 a_n80_n8330# a_380_n8130# w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
X44 w_240_n9000# a_1630_n9420# a_2200_n8070# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X45 a_2200_n8070# a_1630_n9420# w_240_n9000# w_240_n9000# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.6
X46 a_540_n9930# I_IN I_IN a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.6
X47 a_2200_n8070# a_2790_n9420# a_540_n9930# a_540_n9930# sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.6
.ends

.subckt B a_4510_n8940# a_5700_n9470# a_4510_n8350# w_5530_n8860# a_4510_n7380#
X0 a_4510_n8350# p_right a_5700_n9470# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X1 w_5530_n8860# p_bias v_common_p w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X2 p_left a_4510_n7380# v_common_p w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X3 a_4510_n8350# n_right w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 n_right a_4510_n8940# v_common_n a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X5 v_common_p p_bias w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X6 a_5700_n9470# p_right a_4510_n8350# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X7 p_right p_left a_5700_n9470# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X8 p_bias n_bias a_5700_n9470# sky130_fd_pr__res_xhigh_po_2p85 l=0.51
X9 v_common_p p_bias w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X10 w_5530_n8860# n_right a_4510_n8350# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X11 v_common_n a_4510_n8940# n_right a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X12 w_5530_n8860# p_bias p_bias w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X13 a_5700_n9470# p_left p_right a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X14 a_4510_n8350# a_8196_n10872# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X15 n_right n_left w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X16 p_left p_left a_5700_n9470# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0.125 ps=1 w=0.5 l=0.15
X17 n_left a_4510_n7380# v_common_n a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X18 w_5530_n8860# p_bias p_bias w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X19 a_4510_n8350# n_right w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X20 v_common_n n_bias a_5700_n9470# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X21 w_5530_n8860# n_left n_right w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X22 a_5700_n9470# n_bias n_bias a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=1.25 ps=6 w=2.5 l=0.5
X23 v_common_p a_4510_n7380# p_left w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X24 w_5530_n8860# n_right a_4510_n8350# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X25 a_5700_n9470# p_left p_left a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.25 ps=2 w=0.5 l=0.15
X26 a_4510_n8350# a_5270_n10872# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X27 p_bias p_bias w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X28 a_4510_n8350# p_right a_5700_n9470# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X29 n_right a_8196_n10872# a_5700_n9470# sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X30 n_left n_left w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X31 p_right a_4510_n8940# v_common_p w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X32 p_bias p_bias w_5530_n8860# w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X33 a_5270_n10872# p_right a_5700_n9470# sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X34 w_5530_n8860# p_bias v_common_p w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X35 v_common_p a_4510_n8940# p_right w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X36 w_5530_n8860# n_left n_left w_5530_n8860# sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X37 a_5700_n9470# p_right a_4510_n8350# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X38 n_bias n_bias a_5700_n9470# a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=1.25 pd=6 as=0.625 ps=3 w=2.5 l=0.5
X39 a_5700_n9470# n_bias v_common_n a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X40 v_common_n a_4510_n7380# n_left a_5700_n9470# sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
.ends

**.subckt charge_pump_full_4
XA_0 GDDA V_OUT VDDA x A_0/a_380_n8130# A
XB_0 V_OUT GDDA A_0/a_380_n8130# VDDA x B
**.ends

