magic
tech sky130A
timestamp 1752163061
<< nwell >>
rect -30 2305 310 2695
rect 440 2305 780 2525
rect 910 2305 1250 2695
rect 1378 2305 1718 2695
rect -1145 1730 -265 2120
rect -100 1730 780 2120
rect 910 1730 1790 2120
rect 1955 1730 2835 2120
rect 160 1465 1530 1550
rect 160 1460 1525 1465
rect -1115 815 -295 1455
rect -65 1135 755 1225
rect 935 1135 1755 1225
rect 1985 815 2805 1455
rect -1115 400 -295 640
rect 1985 400 2805 640
<< nmos >>
rect 535 830 550 880
rect 590 830 605 880
rect 645 830 660 880
rect 700 830 715 880
rect 755 830 770 880
rect 810 830 825 880
rect 865 830 880 880
rect 920 830 935 880
rect 975 830 990 880
rect 1030 830 1045 880
rect 1085 830 1100 880
rect 1140 830 1155 880
rect 15 455 30 605
rect 70 455 85 605
rect 125 455 140 605
rect 180 455 195 605
rect 235 455 250 605
rect 290 455 305 605
rect 345 455 360 605
rect 400 455 415 605
rect 455 455 470 605
rect 510 455 525 605
rect 565 455 580 605
rect 620 455 635 605
rect 1055 455 1070 605
rect 1110 455 1125 605
rect 1165 455 1180 605
rect 1220 455 1235 605
rect 1275 455 1290 605
rect 1330 455 1345 605
rect 1385 455 1400 605
rect 1440 455 1455 605
rect 1495 455 1510 605
rect 1550 455 1565 605
rect 1605 455 1620 605
rect 1660 455 1675 605
rect -1015 -70 -1000 230
rect -960 -70 -945 230
rect -905 -70 -890 230
rect -850 -70 -835 230
rect -795 -70 -780 230
rect -740 -70 -725 230
rect -685 -70 -670 230
rect -630 -70 -615 230
rect -575 -70 -560 230
rect -520 -70 -505 230
rect -465 -70 -450 230
rect -410 -70 -395 230
rect 15 -20 30 130
rect 70 -20 85 130
rect 125 -20 140 130
rect 180 -20 195 130
rect 235 -20 250 130
rect 290 -20 305 130
rect 345 -20 360 130
rect 400 -20 415 130
rect 455 -20 470 130
rect 510 -20 525 130
rect 565 -20 580 130
rect 620 -20 635 130
rect 755 -20 770 130
rect 810 -20 825 130
rect 865 -20 880 130
rect 920 -20 935 130
rect 1055 -20 1070 130
rect 1110 -20 1125 130
rect 1165 -20 1180 130
rect 1220 -20 1235 130
rect 1275 -20 1290 130
rect 1330 -20 1345 130
rect 1385 -20 1400 130
rect 1440 -20 1455 130
rect 1495 -20 1510 130
rect 1550 -20 1565 130
rect 1605 -20 1620 130
rect 1660 -20 1675 130
rect 2085 -70 2100 230
rect 2140 -70 2155 230
rect 2195 -70 2210 230
rect 2250 -70 2265 230
rect 2305 -70 2320 230
rect 2360 -70 2375 230
rect 2415 -70 2430 230
rect 2470 -70 2485 230
rect 2525 -70 2540 230
rect 2580 -70 2595 230
rect 2635 -70 2650 230
rect 2690 -70 2705 230
rect -985 -1055 -925 -355
rect -885 -1055 -825 -355
rect -785 -1055 -725 -355
rect -685 -1055 -625 -355
rect -585 -1055 -525 -355
rect -485 -1055 -425 -355
rect 200 -655 215 -405
rect 255 -655 270 -405
rect 310 -655 325 -405
rect 365 -655 380 -405
rect 420 -655 435 -405
rect 475 -655 490 -405
rect 530 -655 545 -405
rect 585 -655 600 -405
rect 640 -655 655 -405
rect 695 -655 710 -405
rect 750 -655 765 -405
rect 805 -655 820 -405
rect 860 -655 875 -405
rect 915 -655 930 -405
rect 970 -655 985 -405
rect 1025 -655 1040 -405
rect 1080 -655 1095 -405
rect 1135 -655 1150 -405
rect 1190 -655 1205 -405
rect 1245 -655 1260 -405
rect 1300 -655 1315 -405
rect 1355 -655 1370 -405
rect 1410 -655 1425 -405
rect 705 -920 995 -820
rect 2115 -1055 2175 -355
rect 2215 -1055 2275 -355
rect 2315 -1055 2375 -355
rect 2415 -1055 2475 -355
rect 2515 -1055 2575 -355
rect 2615 -1055 2675 -355
<< pmos >>
rect 70 2325 90 2675
rect 130 2325 150 2675
rect 190 2325 210 2675
rect 540 2325 560 2505
rect 600 2325 620 2505
rect 660 2325 680 2505
rect 1010 2325 1030 2675
rect 1070 2325 1090 2675
rect 1130 2325 1150 2675
rect 1478 2325 1498 2675
rect 1538 2325 1558 2675
rect 1598 2325 1618 2675
rect -1045 1750 -1025 2100
rect -985 1750 -965 2100
rect -925 1750 -905 2100
rect -865 1750 -845 2100
rect -805 1750 -785 2100
rect -745 1750 -725 2100
rect -685 1750 -665 2100
rect -625 1750 -605 2100
rect -565 1750 -545 2100
rect -505 1750 -485 2100
rect -445 1750 -425 2100
rect -385 1750 -365 2100
rect 0 1750 20 2100
rect 60 1750 80 2100
rect 120 1750 140 2100
rect 180 1750 200 2100
rect 240 1750 260 2100
rect 300 1750 320 2100
rect 360 1750 380 2100
rect 420 1750 440 2100
rect 480 1750 500 2100
rect 540 1750 560 2100
rect 600 1750 620 2100
rect 660 1750 680 2100
rect 1010 1750 1030 2100
rect 1070 1750 1090 2100
rect 1130 1750 1150 2100
rect 1190 1750 1210 2100
rect 1250 1750 1270 2100
rect 1310 1750 1330 2100
rect 1370 1750 1390 2100
rect 1430 1750 1450 2100
rect 1490 1750 1510 2100
rect 1550 1750 1570 2100
rect 1610 1750 1630 2100
rect 1670 1750 1690 2100
rect 2055 1750 2075 2100
rect 2115 1750 2135 2100
rect 2175 1750 2195 2100
rect 2235 1750 2255 2100
rect 2295 1750 2315 2100
rect 2355 1750 2375 2100
rect 2415 1750 2435 2100
rect 2475 1750 2495 2100
rect 2535 1750 2555 2100
rect 2595 1750 2615 2100
rect 2655 1750 2675 2100
rect 2715 1750 2735 2100
rect 260 1480 275 1530
rect 315 1480 330 1530
rect 370 1480 385 1530
rect 425 1480 440 1530
rect 480 1480 495 1530
rect 535 1480 550 1530
rect 590 1480 605 1530
rect 645 1480 660 1530
rect 700 1480 715 1530
rect 755 1480 770 1530
rect 810 1480 825 1530
rect 865 1480 880 1530
rect 920 1480 935 1530
rect 975 1480 990 1530
rect 1030 1480 1045 1530
rect 1085 1480 1100 1530
rect 1140 1480 1155 1530
rect 1195 1480 1210 1530
rect 1250 1480 1265 1530
rect 1305 1480 1320 1530
rect 1360 1480 1375 1530
rect 1415 1480 1430 1530
rect -1015 835 -1000 1435
rect -960 835 -945 1435
rect -905 835 -890 1435
rect -850 835 -835 1435
rect -795 835 -780 1435
rect -740 835 -725 1435
rect -685 835 -670 1435
rect -630 835 -615 1435
rect -575 835 -560 1435
rect -520 835 -505 1435
rect -465 835 -450 1435
rect -410 835 -395 1435
rect 35 1155 50 1205
rect 90 1155 105 1205
rect 145 1155 160 1205
rect 200 1155 215 1205
rect 255 1155 270 1205
rect 310 1155 325 1205
rect 365 1155 380 1205
rect 420 1155 435 1205
rect 475 1155 490 1205
rect 530 1155 545 1205
rect 585 1155 600 1205
rect 640 1155 655 1205
rect 1035 1155 1050 1205
rect 1090 1155 1105 1205
rect 1145 1155 1160 1205
rect 1200 1155 1215 1205
rect 1255 1155 1270 1205
rect 1310 1155 1325 1205
rect 1365 1155 1380 1205
rect 1420 1155 1435 1205
rect 1475 1155 1490 1205
rect 1530 1155 1545 1205
rect 1585 1155 1600 1205
rect 1640 1155 1655 1205
rect 2085 835 2100 1435
rect 2140 835 2155 1435
rect 2195 835 2210 1435
rect 2250 835 2265 1435
rect 2305 835 2320 1435
rect 2360 835 2375 1435
rect 2415 835 2430 1435
rect 2470 835 2485 1435
rect 2525 835 2540 1435
rect 2580 835 2595 1435
rect 2635 835 2650 1435
rect 2690 835 2705 1435
rect -1015 420 -1000 620
rect -960 420 -945 620
rect -905 420 -890 620
rect -850 420 -835 620
rect -795 420 -780 620
rect -740 420 -725 620
rect -685 420 -670 620
rect -630 420 -615 620
rect -575 420 -560 620
rect -520 420 -505 620
rect -465 420 -450 620
rect -410 420 -395 620
rect 2085 420 2100 620
rect 2140 420 2155 620
rect 2195 420 2210 620
rect 2250 420 2265 620
rect 2305 420 2320 620
rect 2360 420 2375 620
rect 2415 420 2430 620
rect 2470 420 2485 620
rect 2525 420 2540 620
rect 2580 420 2595 620
rect 2635 420 2650 620
rect 2690 420 2705 620
<< ndiff >>
rect 495 865 535 880
rect 495 845 505 865
rect 525 845 535 865
rect 495 830 535 845
rect 550 865 590 880
rect 550 845 560 865
rect 580 845 590 865
rect 550 830 590 845
rect 605 865 645 880
rect 605 845 615 865
rect 635 845 645 865
rect 605 830 645 845
rect 660 865 700 880
rect 660 845 670 865
rect 690 845 700 865
rect 660 830 700 845
rect 715 865 755 880
rect 715 845 725 865
rect 745 845 755 865
rect 715 830 755 845
rect 770 865 810 880
rect 770 845 780 865
rect 800 845 810 865
rect 770 830 810 845
rect 825 865 865 880
rect 825 845 835 865
rect 855 845 865 865
rect 825 830 865 845
rect 880 865 920 880
rect 880 845 890 865
rect 910 845 920 865
rect 880 830 920 845
rect 935 865 975 880
rect 935 845 945 865
rect 965 845 975 865
rect 935 830 975 845
rect 990 865 1030 880
rect 990 845 1000 865
rect 1020 845 1030 865
rect 990 830 1030 845
rect 1045 865 1085 880
rect 1045 845 1055 865
rect 1075 845 1085 865
rect 1045 830 1085 845
rect 1100 865 1140 880
rect 1100 845 1110 865
rect 1130 845 1140 865
rect 1100 830 1140 845
rect 1155 865 1195 880
rect 1155 845 1165 865
rect 1185 845 1195 865
rect 1155 830 1195 845
rect -25 590 15 605
rect -25 570 -15 590
rect 5 570 15 590
rect -25 540 15 570
rect -25 520 -15 540
rect 5 520 15 540
rect -25 490 15 520
rect -25 470 -15 490
rect 5 470 15 490
rect -25 455 15 470
rect 30 590 70 605
rect 30 570 40 590
rect 60 570 70 590
rect 30 540 70 570
rect 30 520 40 540
rect 60 520 70 540
rect 30 490 70 520
rect 30 470 40 490
rect 60 470 70 490
rect 30 455 70 470
rect 85 590 125 605
rect 85 570 95 590
rect 115 570 125 590
rect 85 540 125 570
rect 85 520 95 540
rect 115 520 125 540
rect 85 490 125 520
rect 85 470 95 490
rect 115 470 125 490
rect 85 455 125 470
rect 140 590 180 605
rect 140 570 150 590
rect 170 570 180 590
rect 140 540 180 570
rect 140 520 150 540
rect 170 520 180 540
rect 140 490 180 520
rect 140 470 150 490
rect 170 470 180 490
rect 140 455 180 470
rect 195 590 235 605
rect 195 570 205 590
rect 225 570 235 590
rect 195 540 235 570
rect 195 520 205 540
rect 225 520 235 540
rect 195 490 235 520
rect 195 470 205 490
rect 225 470 235 490
rect 195 455 235 470
rect 250 590 290 605
rect 250 570 260 590
rect 280 570 290 590
rect 250 540 290 570
rect 250 520 260 540
rect 280 520 290 540
rect 250 490 290 520
rect 250 470 260 490
rect 280 470 290 490
rect 250 455 290 470
rect 305 590 345 605
rect 305 570 315 590
rect 335 570 345 590
rect 305 540 345 570
rect 305 520 315 540
rect 335 520 345 540
rect 305 490 345 520
rect 305 470 315 490
rect 335 470 345 490
rect 305 455 345 470
rect 360 590 400 605
rect 360 570 370 590
rect 390 570 400 590
rect 360 540 400 570
rect 360 520 370 540
rect 390 520 400 540
rect 360 490 400 520
rect 360 470 370 490
rect 390 470 400 490
rect 360 455 400 470
rect 415 590 455 605
rect 415 570 425 590
rect 445 570 455 590
rect 415 540 455 570
rect 415 520 425 540
rect 445 520 455 540
rect 415 490 455 520
rect 415 470 425 490
rect 445 470 455 490
rect 415 455 455 470
rect 470 590 510 605
rect 470 570 480 590
rect 500 570 510 590
rect 470 540 510 570
rect 470 520 480 540
rect 500 520 510 540
rect 470 490 510 520
rect 470 470 480 490
rect 500 470 510 490
rect 470 455 510 470
rect 525 590 565 605
rect 525 570 535 590
rect 555 570 565 590
rect 525 540 565 570
rect 525 520 535 540
rect 555 520 565 540
rect 525 490 565 520
rect 525 470 535 490
rect 555 470 565 490
rect 525 455 565 470
rect 580 590 620 605
rect 580 570 590 590
rect 610 570 620 590
rect 580 540 620 570
rect 580 520 590 540
rect 610 520 620 540
rect 580 490 620 520
rect 580 470 590 490
rect 610 470 620 490
rect 580 455 620 470
rect 635 590 675 605
rect 635 570 645 590
rect 665 570 675 590
rect 635 540 675 570
rect 635 520 645 540
rect 665 520 675 540
rect 635 490 675 520
rect 635 470 645 490
rect 665 470 675 490
rect 635 455 675 470
rect 1015 590 1055 605
rect 1015 570 1025 590
rect 1045 570 1055 590
rect 1015 540 1055 570
rect 1015 520 1025 540
rect 1045 520 1055 540
rect 1015 490 1055 520
rect 1015 470 1025 490
rect 1045 470 1055 490
rect 1015 455 1055 470
rect 1070 590 1110 605
rect 1070 570 1080 590
rect 1100 570 1110 590
rect 1070 540 1110 570
rect 1070 520 1080 540
rect 1100 520 1110 540
rect 1070 490 1110 520
rect 1070 470 1080 490
rect 1100 470 1110 490
rect 1070 455 1110 470
rect 1125 590 1165 605
rect 1125 570 1135 590
rect 1155 570 1165 590
rect 1125 540 1165 570
rect 1125 520 1135 540
rect 1155 520 1165 540
rect 1125 490 1165 520
rect 1125 470 1135 490
rect 1155 470 1165 490
rect 1125 455 1165 470
rect 1180 590 1220 605
rect 1180 570 1190 590
rect 1210 570 1220 590
rect 1180 540 1220 570
rect 1180 520 1190 540
rect 1210 520 1220 540
rect 1180 490 1220 520
rect 1180 470 1190 490
rect 1210 470 1220 490
rect 1180 455 1220 470
rect 1235 590 1275 605
rect 1235 570 1245 590
rect 1265 570 1275 590
rect 1235 540 1275 570
rect 1235 520 1245 540
rect 1265 520 1275 540
rect 1235 490 1275 520
rect 1235 470 1245 490
rect 1265 470 1275 490
rect 1235 455 1275 470
rect 1290 590 1330 605
rect 1290 570 1300 590
rect 1320 570 1330 590
rect 1290 540 1330 570
rect 1290 520 1300 540
rect 1320 520 1330 540
rect 1290 490 1330 520
rect 1290 470 1300 490
rect 1320 470 1330 490
rect 1290 455 1330 470
rect 1345 590 1385 605
rect 1345 570 1355 590
rect 1375 570 1385 590
rect 1345 540 1385 570
rect 1345 520 1355 540
rect 1375 520 1385 540
rect 1345 490 1385 520
rect 1345 470 1355 490
rect 1375 470 1385 490
rect 1345 455 1385 470
rect 1400 590 1440 605
rect 1400 570 1410 590
rect 1430 570 1440 590
rect 1400 540 1440 570
rect 1400 520 1410 540
rect 1430 520 1440 540
rect 1400 490 1440 520
rect 1400 470 1410 490
rect 1430 470 1440 490
rect 1400 455 1440 470
rect 1455 590 1495 605
rect 1455 570 1465 590
rect 1485 570 1495 590
rect 1455 540 1495 570
rect 1455 520 1465 540
rect 1485 520 1495 540
rect 1455 490 1495 520
rect 1455 470 1465 490
rect 1485 470 1495 490
rect 1455 455 1495 470
rect 1510 590 1550 605
rect 1510 570 1520 590
rect 1540 570 1550 590
rect 1510 540 1550 570
rect 1510 520 1520 540
rect 1540 520 1550 540
rect 1510 490 1550 520
rect 1510 470 1520 490
rect 1540 470 1550 490
rect 1510 455 1550 470
rect 1565 590 1605 605
rect 1565 570 1575 590
rect 1595 570 1605 590
rect 1565 540 1605 570
rect 1565 520 1575 540
rect 1595 520 1605 540
rect 1565 490 1605 520
rect 1565 470 1575 490
rect 1595 470 1605 490
rect 1565 455 1605 470
rect 1620 590 1660 605
rect 1620 570 1630 590
rect 1650 570 1660 590
rect 1620 540 1660 570
rect 1620 520 1630 540
rect 1650 520 1660 540
rect 1620 490 1660 520
rect 1620 470 1630 490
rect 1650 470 1660 490
rect 1620 455 1660 470
rect 1675 590 1715 605
rect 1675 570 1685 590
rect 1705 570 1715 590
rect 1675 540 1715 570
rect 1675 520 1685 540
rect 1705 520 1715 540
rect 1675 490 1715 520
rect 1675 470 1685 490
rect 1705 470 1715 490
rect 1675 455 1715 470
rect -1055 215 -1015 230
rect -1055 195 -1045 215
rect -1025 195 -1015 215
rect -1055 165 -1015 195
rect -1055 145 -1045 165
rect -1025 145 -1015 165
rect -1055 115 -1015 145
rect -1055 95 -1045 115
rect -1025 95 -1015 115
rect -1055 65 -1015 95
rect -1055 45 -1045 65
rect -1025 45 -1015 65
rect -1055 15 -1015 45
rect -1055 -5 -1045 15
rect -1025 -5 -1015 15
rect -1055 -35 -1015 -5
rect -1055 -55 -1045 -35
rect -1025 -55 -1015 -35
rect -1055 -70 -1015 -55
rect -1000 215 -960 230
rect -1000 195 -990 215
rect -970 195 -960 215
rect -1000 165 -960 195
rect -1000 145 -990 165
rect -970 145 -960 165
rect -1000 115 -960 145
rect -1000 95 -990 115
rect -970 95 -960 115
rect -1000 65 -960 95
rect -1000 45 -990 65
rect -970 45 -960 65
rect -1000 15 -960 45
rect -1000 -5 -990 15
rect -970 -5 -960 15
rect -1000 -35 -960 -5
rect -1000 -55 -990 -35
rect -970 -55 -960 -35
rect -1000 -70 -960 -55
rect -945 215 -905 230
rect -945 195 -935 215
rect -915 195 -905 215
rect -945 165 -905 195
rect -945 145 -935 165
rect -915 145 -905 165
rect -945 115 -905 145
rect -945 95 -935 115
rect -915 95 -905 115
rect -945 65 -905 95
rect -945 45 -935 65
rect -915 45 -905 65
rect -945 15 -905 45
rect -945 -5 -935 15
rect -915 -5 -905 15
rect -945 -35 -905 -5
rect -945 -55 -935 -35
rect -915 -55 -905 -35
rect -945 -70 -905 -55
rect -890 215 -850 230
rect -890 195 -880 215
rect -860 195 -850 215
rect -890 165 -850 195
rect -890 145 -880 165
rect -860 145 -850 165
rect -890 115 -850 145
rect -890 95 -880 115
rect -860 95 -850 115
rect -890 65 -850 95
rect -890 45 -880 65
rect -860 45 -850 65
rect -890 15 -850 45
rect -890 -5 -880 15
rect -860 -5 -850 15
rect -890 -35 -850 -5
rect -890 -55 -880 -35
rect -860 -55 -850 -35
rect -890 -70 -850 -55
rect -835 215 -795 230
rect -835 195 -825 215
rect -805 195 -795 215
rect -835 165 -795 195
rect -835 145 -825 165
rect -805 145 -795 165
rect -835 115 -795 145
rect -835 95 -825 115
rect -805 95 -795 115
rect -835 65 -795 95
rect -835 45 -825 65
rect -805 45 -795 65
rect -835 15 -795 45
rect -835 -5 -825 15
rect -805 -5 -795 15
rect -835 -35 -795 -5
rect -835 -55 -825 -35
rect -805 -55 -795 -35
rect -835 -70 -795 -55
rect -780 215 -740 230
rect -780 195 -770 215
rect -750 195 -740 215
rect -780 165 -740 195
rect -780 145 -770 165
rect -750 145 -740 165
rect -780 115 -740 145
rect -780 95 -770 115
rect -750 95 -740 115
rect -780 65 -740 95
rect -780 45 -770 65
rect -750 45 -740 65
rect -780 15 -740 45
rect -780 -5 -770 15
rect -750 -5 -740 15
rect -780 -35 -740 -5
rect -780 -55 -770 -35
rect -750 -55 -740 -35
rect -780 -70 -740 -55
rect -725 215 -685 230
rect -725 195 -715 215
rect -695 195 -685 215
rect -725 165 -685 195
rect -725 145 -715 165
rect -695 145 -685 165
rect -725 115 -685 145
rect -725 95 -715 115
rect -695 95 -685 115
rect -725 65 -685 95
rect -725 45 -715 65
rect -695 45 -685 65
rect -725 15 -685 45
rect -725 -5 -715 15
rect -695 -5 -685 15
rect -725 -35 -685 -5
rect -725 -55 -715 -35
rect -695 -55 -685 -35
rect -725 -70 -685 -55
rect -670 215 -630 230
rect -670 195 -660 215
rect -640 195 -630 215
rect -670 165 -630 195
rect -670 145 -660 165
rect -640 145 -630 165
rect -670 115 -630 145
rect -670 95 -660 115
rect -640 95 -630 115
rect -670 65 -630 95
rect -670 45 -660 65
rect -640 45 -630 65
rect -670 15 -630 45
rect -670 -5 -660 15
rect -640 -5 -630 15
rect -670 -35 -630 -5
rect -670 -55 -660 -35
rect -640 -55 -630 -35
rect -670 -70 -630 -55
rect -615 215 -575 230
rect -615 195 -605 215
rect -585 195 -575 215
rect -615 165 -575 195
rect -615 145 -605 165
rect -585 145 -575 165
rect -615 115 -575 145
rect -615 95 -605 115
rect -585 95 -575 115
rect -615 65 -575 95
rect -615 45 -605 65
rect -585 45 -575 65
rect -615 15 -575 45
rect -615 -5 -605 15
rect -585 -5 -575 15
rect -615 -35 -575 -5
rect -615 -55 -605 -35
rect -585 -55 -575 -35
rect -615 -70 -575 -55
rect -560 215 -520 230
rect -560 195 -550 215
rect -530 195 -520 215
rect -560 165 -520 195
rect -560 145 -550 165
rect -530 145 -520 165
rect -560 115 -520 145
rect -560 95 -550 115
rect -530 95 -520 115
rect -560 65 -520 95
rect -560 45 -550 65
rect -530 45 -520 65
rect -560 15 -520 45
rect -560 -5 -550 15
rect -530 -5 -520 15
rect -560 -35 -520 -5
rect -560 -55 -550 -35
rect -530 -55 -520 -35
rect -560 -70 -520 -55
rect -505 215 -465 230
rect -505 195 -495 215
rect -475 195 -465 215
rect -505 165 -465 195
rect -505 145 -495 165
rect -475 145 -465 165
rect -505 115 -465 145
rect -505 95 -495 115
rect -475 95 -465 115
rect -505 65 -465 95
rect -505 45 -495 65
rect -475 45 -465 65
rect -505 15 -465 45
rect -505 -5 -495 15
rect -475 -5 -465 15
rect -505 -35 -465 -5
rect -505 -55 -495 -35
rect -475 -55 -465 -35
rect -505 -70 -465 -55
rect -450 215 -410 230
rect -450 195 -440 215
rect -420 195 -410 215
rect -450 165 -410 195
rect -450 145 -440 165
rect -420 145 -410 165
rect -450 115 -410 145
rect -450 95 -440 115
rect -420 95 -410 115
rect -450 65 -410 95
rect -450 45 -440 65
rect -420 45 -410 65
rect -450 15 -410 45
rect -450 -5 -440 15
rect -420 -5 -410 15
rect -450 -35 -410 -5
rect -450 -55 -440 -35
rect -420 -55 -410 -35
rect -450 -70 -410 -55
rect -395 215 -355 230
rect -395 195 -385 215
rect -365 195 -355 215
rect -395 165 -355 195
rect 2045 215 2085 230
rect 2045 195 2055 215
rect 2075 195 2085 215
rect -395 145 -385 165
rect -365 145 -355 165
rect -395 115 -355 145
rect 2045 165 2085 195
rect 2045 145 2055 165
rect 2075 145 2085 165
rect -395 95 -385 115
rect -365 95 -355 115
rect -395 65 -355 95
rect -395 45 -385 65
rect -365 45 -355 65
rect -395 15 -355 45
rect -395 -5 -385 15
rect -365 -5 -355 15
rect -395 -35 -355 -5
rect -25 115 15 130
rect -25 95 -15 115
rect 5 95 15 115
rect -25 65 15 95
rect -25 45 -15 65
rect 5 45 15 65
rect -25 15 15 45
rect -25 -5 -15 15
rect 5 -5 15 15
rect -25 -20 15 -5
rect 30 115 70 130
rect 30 95 40 115
rect 60 95 70 115
rect 30 65 70 95
rect 30 45 40 65
rect 60 45 70 65
rect 30 15 70 45
rect 30 -5 40 15
rect 60 -5 70 15
rect 30 -20 70 -5
rect 85 115 125 130
rect 85 95 95 115
rect 115 95 125 115
rect 85 65 125 95
rect 85 45 95 65
rect 115 45 125 65
rect 85 15 125 45
rect 85 -5 95 15
rect 115 -5 125 15
rect 85 -20 125 -5
rect 140 115 180 130
rect 140 95 150 115
rect 170 95 180 115
rect 140 65 180 95
rect 140 45 150 65
rect 170 45 180 65
rect 140 15 180 45
rect 140 -5 150 15
rect 170 -5 180 15
rect 140 -20 180 -5
rect 195 115 235 130
rect 195 95 205 115
rect 225 95 235 115
rect 195 65 235 95
rect 195 45 205 65
rect 225 45 235 65
rect 195 15 235 45
rect 195 -5 205 15
rect 225 -5 235 15
rect 195 -20 235 -5
rect 250 115 290 130
rect 250 95 260 115
rect 280 95 290 115
rect 250 65 290 95
rect 250 45 260 65
rect 280 45 290 65
rect 250 15 290 45
rect 250 -5 260 15
rect 280 -5 290 15
rect 250 -20 290 -5
rect 305 115 345 130
rect 305 95 315 115
rect 335 95 345 115
rect 305 65 345 95
rect 305 45 315 65
rect 335 45 345 65
rect 305 15 345 45
rect 305 -5 315 15
rect 335 -5 345 15
rect 305 -20 345 -5
rect 360 115 400 130
rect 360 95 370 115
rect 390 95 400 115
rect 360 65 400 95
rect 360 45 370 65
rect 390 45 400 65
rect 360 15 400 45
rect 360 -5 370 15
rect 390 -5 400 15
rect 360 -20 400 -5
rect 415 115 455 130
rect 415 95 425 115
rect 445 95 455 115
rect 415 65 455 95
rect 415 45 425 65
rect 445 45 455 65
rect 415 15 455 45
rect 415 -5 425 15
rect 445 -5 455 15
rect 415 -20 455 -5
rect 470 115 510 130
rect 470 95 480 115
rect 500 95 510 115
rect 470 65 510 95
rect 470 45 480 65
rect 500 45 510 65
rect 470 15 510 45
rect 470 -5 480 15
rect 500 -5 510 15
rect 470 -20 510 -5
rect 525 115 565 130
rect 525 95 535 115
rect 555 95 565 115
rect 525 65 565 95
rect 525 45 535 65
rect 555 45 565 65
rect 525 15 565 45
rect 525 -5 535 15
rect 555 -5 565 15
rect 525 -20 565 -5
rect 580 115 620 130
rect 580 95 590 115
rect 610 95 620 115
rect 580 65 620 95
rect 580 45 590 65
rect 610 45 620 65
rect 580 15 620 45
rect 580 -5 590 15
rect 610 -5 620 15
rect 580 -20 620 -5
rect 635 115 675 130
rect 715 115 755 130
rect 635 95 645 115
rect 665 95 675 115
rect 715 95 725 115
rect 745 95 755 115
rect 635 65 675 95
rect 715 65 755 95
rect 635 45 645 65
rect 665 45 675 65
rect 715 45 725 65
rect 745 45 755 65
rect 635 15 675 45
rect 715 15 755 45
rect 635 -5 645 15
rect 665 -5 675 15
rect 715 -5 725 15
rect 745 -5 755 15
rect 635 -20 675 -5
rect 715 -20 755 -5
rect 770 115 810 130
rect 770 95 780 115
rect 800 95 810 115
rect 770 65 810 95
rect 770 45 780 65
rect 800 45 810 65
rect 770 15 810 45
rect 770 -5 780 15
rect 800 -5 810 15
rect 770 -20 810 -5
rect 825 115 865 130
rect 825 95 835 115
rect 855 95 865 115
rect 825 65 865 95
rect 825 45 835 65
rect 855 45 865 65
rect 825 15 865 45
rect 825 -5 835 15
rect 855 -5 865 15
rect 825 -20 865 -5
rect 880 115 920 130
rect 880 95 890 115
rect 910 95 920 115
rect 880 65 920 95
rect 880 45 890 65
rect 910 45 920 65
rect 880 15 920 45
rect 880 -5 890 15
rect 910 -5 920 15
rect 880 -20 920 -5
rect 935 115 975 130
rect 1015 115 1055 130
rect 935 95 945 115
rect 965 95 975 115
rect 1015 95 1025 115
rect 1045 95 1055 115
rect 935 65 975 95
rect 1015 65 1055 95
rect 935 45 945 65
rect 965 45 975 65
rect 1015 45 1025 65
rect 1045 45 1055 65
rect 935 15 975 45
rect 1015 15 1055 45
rect 935 -5 945 15
rect 965 -5 975 15
rect 1015 -5 1025 15
rect 1045 -5 1055 15
rect 935 -20 975 -5
rect 1015 -20 1055 -5
rect 1070 115 1110 130
rect 1070 95 1080 115
rect 1100 95 1110 115
rect 1070 65 1110 95
rect 1070 45 1080 65
rect 1100 45 1110 65
rect 1070 15 1110 45
rect 1070 -5 1080 15
rect 1100 -5 1110 15
rect 1070 -20 1110 -5
rect 1125 115 1165 130
rect 1125 95 1135 115
rect 1155 95 1165 115
rect 1125 65 1165 95
rect 1125 45 1135 65
rect 1155 45 1165 65
rect 1125 15 1165 45
rect 1125 -5 1135 15
rect 1155 -5 1165 15
rect 1125 -20 1165 -5
rect 1180 115 1220 130
rect 1180 95 1190 115
rect 1210 95 1220 115
rect 1180 65 1220 95
rect 1180 45 1190 65
rect 1210 45 1220 65
rect 1180 15 1220 45
rect 1180 -5 1190 15
rect 1210 -5 1220 15
rect 1180 -20 1220 -5
rect 1235 115 1275 130
rect 1235 95 1245 115
rect 1265 95 1275 115
rect 1235 65 1275 95
rect 1235 45 1245 65
rect 1265 45 1275 65
rect 1235 15 1275 45
rect 1235 -5 1245 15
rect 1265 -5 1275 15
rect 1235 -20 1275 -5
rect 1290 115 1330 130
rect 1290 95 1300 115
rect 1320 95 1330 115
rect 1290 65 1330 95
rect 1290 45 1300 65
rect 1320 45 1330 65
rect 1290 15 1330 45
rect 1290 -5 1300 15
rect 1320 -5 1330 15
rect 1290 -20 1330 -5
rect 1345 115 1385 130
rect 1345 95 1355 115
rect 1375 95 1385 115
rect 1345 65 1385 95
rect 1345 45 1355 65
rect 1375 45 1385 65
rect 1345 15 1385 45
rect 1345 -5 1355 15
rect 1375 -5 1385 15
rect 1345 -20 1385 -5
rect 1400 115 1440 130
rect 1400 95 1410 115
rect 1430 95 1440 115
rect 1400 65 1440 95
rect 1400 45 1410 65
rect 1430 45 1440 65
rect 1400 15 1440 45
rect 1400 -5 1410 15
rect 1430 -5 1440 15
rect 1400 -20 1440 -5
rect 1455 115 1495 130
rect 1455 95 1465 115
rect 1485 95 1495 115
rect 1455 65 1495 95
rect 1455 45 1465 65
rect 1485 45 1495 65
rect 1455 15 1495 45
rect 1455 -5 1465 15
rect 1485 -5 1495 15
rect 1455 -20 1495 -5
rect 1510 115 1550 130
rect 1510 95 1520 115
rect 1540 95 1550 115
rect 1510 65 1550 95
rect 1510 45 1520 65
rect 1540 45 1550 65
rect 1510 15 1550 45
rect 1510 -5 1520 15
rect 1540 -5 1550 15
rect 1510 -20 1550 -5
rect 1565 115 1605 130
rect 1565 95 1575 115
rect 1595 95 1605 115
rect 1565 65 1605 95
rect 1565 45 1575 65
rect 1595 45 1605 65
rect 1565 15 1605 45
rect 1565 -5 1575 15
rect 1595 -5 1605 15
rect 1565 -20 1605 -5
rect 1620 115 1660 130
rect 1620 95 1630 115
rect 1650 95 1660 115
rect 1620 65 1660 95
rect 1620 45 1630 65
rect 1650 45 1660 65
rect 1620 15 1660 45
rect 1620 -5 1630 15
rect 1650 -5 1660 15
rect 1620 -20 1660 -5
rect 1675 115 1715 130
rect 1675 95 1685 115
rect 1705 95 1715 115
rect 1675 65 1715 95
rect 1675 45 1685 65
rect 1705 45 1715 65
rect 1675 15 1715 45
rect 1675 -5 1685 15
rect 1705 -5 1715 15
rect 1675 -20 1715 -5
rect 2045 115 2085 145
rect 2045 95 2055 115
rect 2075 95 2085 115
rect 2045 65 2085 95
rect 2045 45 2055 65
rect 2075 45 2085 65
rect 2045 15 2085 45
rect 2045 -5 2055 15
rect 2075 -5 2085 15
rect 2045 -35 2085 -5
rect -395 -55 -385 -35
rect -365 -55 -355 -35
rect -395 -70 -355 -55
rect 2045 -55 2055 -35
rect 2075 -55 2085 -35
rect 2045 -70 2085 -55
rect 2100 215 2140 230
rect 2100 195 2110 215
rect 2130 195 2140 215
rect 2100 165 2140 195
rect 2100 145 2110 165
rect 2130 145 2140 165
rect 2100 115 2140 145
rect 2100 95 2110 115
rect 2130 95 2140 115
rect 2100 65 2140 95
rect 2100 45 2110 65
rect 2130 45 2140 65
rect 2100 15 2140 45
rect 2100 -5 2110 15
rect 2130 -5 2140 15
rect 2100 -35 2140 -5
rect 2100 -55 2110 -35
rect 2130 -55 2140 -35
rect 2100 -70 2140 -55
rect 2155 215 2195 230
rect 2155 195 2165 215
rect 2185 195 2195 215
rect 2155 165 2195 195
rect 2155 145 2165 165
rect 2185 145 2195 165
rect 2155 115 2195 145
rect 2155 95 2165 115
rect 2185 95 2195 115
rect 2155 65 2195 95
rect 2155 45 2165 65
rect 2185 45 2195 65
rect 2155 15 2195 45
rect 2155 -5 2165 15
rect 2185 -5 2195 15
rect 2155 -35 2195 -5
rect 2155 -55 2165 -35
rect 2185 -55 2195 -35
rect 2155 -70 2195 -55
rect 2210 215 2250 230
rect 2210 195 2220 215
rect 2240 195 2250 215
rect 2210 165 2250 195
rect 2210 145 2220 165
rect 2240 145 2250 165
rect 2210 115 2250 145
rect 2210 95 2220 115
rect 2240 95 2250 115
rect 2210 65 2250 95
rect 2210 45 2220 65
rect 2240 45 2250 65
rect 2210 15 2250 45
rect 2210 -5 2220 15
rect 2240 -5 2250 15
rect 2210 -35 2250 -5
rect 2210 -55 2220 -35
rect 2240 -55 2250 -35
rect 2210 -70 2250 -55
rect 2265 215 2305 230
rect 2265 195 2275 215
rect 2295 195 2305 215
rect 2265 165 2305 195
rect 2265 145 2275 165
rect 2295 145 2305 165
rect 2265 115 2305 145
rect 2265 95 2275 115
rect 2295 95 2305 115
rect 2265 65 2305 95
rect 2265 45 2275 65
rect 2295 45 2305 65
rect 2265 15 2305 45
rect 2265 -5 2275 15
rect 2295 -5 2305 15
rect 2265 -35 2305 -5
rect 2265 -55 2275 -35
rect 2295 -55 2305 -35
rect 2265 -70 2305 -55
rect 2320 215 2360 230
rect 2320 195 2330 215
rect 2350 195 2360 215
rect 2320 165 2360 195
rect 2320 145 2330 165
rect 2350 145 2360 165
rect 2320 115 2360 145
rect 2320 95 2330 115
rect 2350 95 2360 115
rect 2320 65 2360 95
rect 2320 45 2330 65
rect 2350 45 2360 65
rect 2320 15 2360 45
rect 2320 -5 2330 15
rect 2350 -5 2360 15
rect 2320 -35 2360 -5
rect 2320 -55 2330 -35
rect 2350 -55 2360 -35
rect 2320 -70 2360 -55
rect 2375 215 2415 230
rect 2375 195 2385 215
rect 2405 195 2415 215
rect 2375 165 2415 195
rect 2375 145 2385 165
rect 2405 145 2415 165
rect 2375 115 2415 145
rect 2375 95 2385 115
rect 2405 95 2415 115
rect 2375 65 2415 95
rect 2375 45 2385 65
rect 2405 45 2415 65
rect 2375 15 2415 45
rect 2375 -5 2385 15
rect 2405 -5 2415 15
rect 2375 -35 2415 -5
rect 2375 -55 2385 -35
rect 2405 -55 2415 -35
rect 2375 -70 2415 -55
rect 2430 215 2470 230
rect 2430 195 2440 215
rect 2460 195 2470 215
rect 2430 165 2470 195
rect 2430 145 2440 165
rect 2460 145 2470 165
rect 2430 115 2470 145
rect 2430 95 2440 115
rect 2460 95 2470 115
rect 2430 65 2470 95
rect 2430 45 2440 65
rect 2460 45 2470 65
rect 2430 15 2470 45
rect 2430 -5 2440 15
rect 2460 -5 2470 15
rect 2430 -35 2470 -5
rect 2430 -55 2440 -35
rect 2460 -55 2470 -35
rect 2430 -70 2470 -55
rect 2485 215 2525 230
rect 2485 195 2495 215
rect 2515 195 2525 215
rect 2485 165 2525 195
rect 2485 145 2495 165
rect 2515 145 2525 165
rect 2485 115 2525 145
rect 2485 95 2495 115
rect 2515 95 2525 115
rect 2485 65 2525 95
rect 2485 45 2495 65
rect 2515 45 2525 65
rect 2485 15 2525 45
rect 2485 -5 2495 15
rect 2515 -5 2525 15
rect 2485 -35 2525 -5
rect 2485 -55 2495 -35
rect 2515 -55 2525 -35
rect 2485 -70 2525 -55
rect 2540 215 2580 230
rect 2540 195 2550 215
rect 2570 195 2580 215
rect 2540 165 2580 195
rect 2540 145 2550 165
rect 2570 145 2580 165
rect 2540 115 2580 145
rect 2540 95 2550 115
rect 2570 95 2580 115
rect 2540 65 2580 95
rect 2540 45 2550 65
rect 2570 45 2580 65
rect 2540 15 2580 45
rect 2540 -5 2550 15
rect 2570 -5 2580 15
rect 2540 -35 2580 -5
rect 2540 -55 2550 -35
rect 2570 -55 2580 -35
rect 2540 -70 2580 -55
rect 2595 215 2635 230
rect 2595 195 2605 215
rect 2625 195 2635 215
rect 2595 165 2635 195
rect 2595 145 2605 165
rect 2625 145 2635 165
rect 2595 115 2635 145
rect 2595 95 2605 115
rect 2625 95 2635 115
rect 2595 65 2635 95
rect 2595 45 2605 65
rect 2625 45 2635 65
rect 2595 15 2635 45
rect 2595 -5 2605 15
rect 2625 -5 2635 15
rect 2595 -35 2635 -5
rect 2595 -55 2605 -35
rect 2625 -55 2635 -35
rect 2595 -70 2635 -55
rect 2650 215 2690 230
rect 2650 195 2660 215
rect 2680 195 2690 215
rect 2650 165 2690 195
rect 2650 145 2660 165
rect 2680 145 2690 165
rect 2650 115 2690 145
rect 2650 95 2660 115
rect 2680 95 2690 115
rect 2650 65 2690 95
rect 2650 45 2660 65
rect 2680 45 2690 65
rect 2650 15 2690 45
rect 2650 -5 2660 15
rect 2680 -5 2690 15
rect 2650 -35 2690 -5
rect 2650 -55 2660 -35
rect 2680 -55 2690 -35
rect 2650 -70 2690 -55
rect 2705 215 2745 230
rect 2705 195 2715 215
rect 2735 195 2745 215
rect 2705 165 2745 195
rect 2705 145 2715 165
rect 2735 145 2745 165
rect 2705 115 2745 145
rect 2705 95 2715 115
rect 2735 95 2745 115
rect 2705 65 2745 95
rect 2705 45 2715 65
rect 2735 45 2745 65
rect 2705 15 2745 45
rect 2705 -5 2715 15
rect 2735 -5 2745 15
rect 2705 -35 2745 -5
rect 2705 -55 2715 -35
rect 2735 -55 2745 -35
rect 2705 -70 2745 -55
rect -1025 -370 -985 -355
rect -1025 -390 -1015 -370
rect -995 -390 -985 -370
rect -1025 -420 -985 -390
rect -1025 -440 -1015 -420
rect -995 -440 -985 -420
rect -1025 -470 -985 -440
rect -1025 -490 -1015 -470
rect -995 -490 -985 -470
rect -1025 -520 -985 -490
rect -1025 -540 -1015 -520
rect -995 -540 -985 -520
rect -1025 -570 -985 -540
rect -1025 -590 -1015 -570
rect -995 -590 -985 -570
rect -1025 -620 -985 -590
rect -1025 -640 -1015 -620
rect -995 -640 -985 -620
rect -1025 -670 -985 -640
rect -1025 -690 -1015 -670
rect -995 -690 -985 -670
rect -1025 -720 -985 -690
rect -1025 -740 -1015 -720
rect -995 -740 -985 -720
rect -1025 -770 -985 -740
rect -1025 -790 -1015 -770
rect -995 -790 -985 -770
rect -1025 -820 -985 -790
rect -1025 -840 -1015 -820
rect -995 -840 -985 -820
rect -1025 -870 -985 -840
rect -1025 -890 -1015 -870
rect -995 -890 -985 -870
rect -1025 -920 -985 -890
rect -1025 -940 -1015 -920
rect -995 -940 -985 -920
rect -1025 -970 -985 -940
rect -1025 -990 -1015 -970
rect -995 -990 -985 -970
rect -1025 -1020 -985 -990
rect -1025 -1040 -1015 -1020
rect -995 -1040 -985 -1020
rect -1025 -1055 -985 -1040
rect -925 -370 -885 -355
rect -925 -390 -915 -370
rect -895 -390 -885 -370
rect -925 -420 -885 -390
rect -925 -440 -915 -420
rect -895 -440 -885 -420
rect -925 -470 -885 -440
rect -925 -490 -915 -470
rect -895 -490 -885 -470
rect -925 -520 -885 -490
rect -925 -540 -915 -520
rect -895 -540 -885 -520
rect -925 -570 -885 -540
rect -925 -590 -915 -570
rect -895 -590 -885 -570
rect -925 -620 -885 -590
rect -925 -640 -915 -620
rect -895 -640 -885 -620
rect -925 -670 -885 -640
rect -925 -690 -915 -670
rect -895 -690 -885 -670
rect -925 -720 -885 -690
rect -925 -740 -915 -720
rect -895 -740 -885 -720
rect -925 -770 -885 -740
rect -925 -790 -915 -770
rect -895 -790 -885 -770
rect -925 -820 -885 -790
rect -925 -840 -915 -820
rect -895 -840 -885 -820
rect -925 -870 -885 -840
rect -925 -890 -915 -870
rect -895 -890 -885 -870
rect -925 -920 -885 -890
rect -925 -940 -915 -920
rect -895 -940 -885 -920
rect -925 -970 -885 -940
rect -925 -990 -915 -970
rect -895 -990 -885 -970
rect -925 -1020 -885 -990
rect -925 -1040 -915 -1020
rect -895 -1040 -885 -1020
rect -925 -1055 -885 -1040
rect -825 -370 -785 -355
rect -825 -390 -815 -370
rect -795 -390 -785 -370
rect -825 -420 -785 -390
rect -825 -440 -815 -420
rect -795 -440 -785 -420
rect -825 -470 -785 -440
rect -825 -490 -815 -470
rect -795 -490 -785 -470
rect -825 -520 -785 -490
rect -825 -540 -815 -520
rect -795 -540 -785 -520
rect -825 -570 -785 -540
rect -825 -590 -815 -570
rect -795 -590 -785 -570
rect -825 -620 -785 -590
rect -825 -640 -815 -620
rect -795 -640 -785 -620
rect -825 -670 -785 -640
rect -825 -690 -815 -670
rect -795 -690 -785 -670
rect -825 -720 -785 -690
rect -825 -740 -815 -720
rect -795 -740 -785 -720
rect -825 -770 -785 -740
rect -825 -790 -815 -770
rect -795 -790 -785 -770
rect -825 -820 -785 -790
rect -825 -840 -815 -820
rect -795 -840 -785 -820
rect -825 -870 -785 -840
rect -825 -890 -815 -870
rect -795 -890 -785 -870
rect -825 -920 -785 -890
rect -825 -940 -815 -920
rect -795 -940 -785 -920
rect -825 -970 -785 -940
rect -825 -990 -815 -970
rect -795 -990 -785 -970
rect -825 -1020 -785 -990
rect -825 -1040 -815 -1020
rect -795 -1040 -785 -1020
rect -825 -1055 -785 -1040
rect -725 -370 -685 -355
rect -725 -390 -715 -370
rect -695 -390 -685 -370
rect -725 -420 -685 -390
rect -725 -440 -715 -420
rect -695 -440 -685 -420
rect -725 -470 -685 -440
rect -725 -490 -715 -470
rect -695 -490 -685 -470
rect -725 -520 -685 -490
rect -725 -540 -715 -520
rect -695 -540 -685 -520
rect -725 -570 -685 -540
rect -725 -590 -715 -570
rect -695 -590 -685 -570
rect -725 -620 -685 -590
rect -725 -640 -715 -620
rect -695 -640 -685 -620
rect -725 -670 -685 -640
rect -725 -690 -715 -670
rect -695 -690 -685 -670
rect -725 -720 -685 -690
rect -725 -740 -715 -720
rect -695 -740 -685 -720
rect -725 -770 -685 -740
rect -725 -790 -715 -770
rect -695 -790 -685 -770
rect -725 -820 -685 -790
rect -725 -840 -715 -820
rect -695 -840 -685 -820
rect -725 -870 -685 -840
rect -725 -890 -715 -870
rect -695 -890 -685 -870
rect -725 -920 -685 -890
rect -725 -940 -715 -920
rect -695 -940 -685 -920
rect -725 -970 -685 -940
rect -725 -990 -715 -970
rect -695 -990 -685 -970
rect -725 -1020 -685 -990
rect -725 -1040 -715 -1020
rect -695 -1040 -685 -1020
rect -725 -1055 -685 -1040
rect -625 -370 -585 -355
rect -625 -390 -615 -370
rect -595 -390 -585 -370
rect -625 -420 -585 -390
rect -625 -440 -615 -420
rect -595 -440 -585 -420
rect -625 -470 -585 -440
rect -625 -490 -615 -470
rect -595 -490 -585 -470
rect -625 -520 -585 -490
rect -625 -540 -615 -520
rect -595 -540 -585 -520
rect -625 -570 -585 -540
rect -625 -590 -615 -570
rect -595 -590 -585 -570
rect -625 -620 -585 -590
rect -625 -640 -615 -620
rect -595 -640 -585 -620
rect -625 -670 -585 -640
rect -625 -690 -615 -670
rect -595 -690 -585 -670
rect -625 -720 -585 -690
rect -625 -740 -615 -720
rect -595 -740 -585 -720
rect -625 -770 -585 -740
rect -625 -790 -615 -770
rect -595 -790 -585 -770
rect -625 -820 -585 -790
rect -625 -840 -615 -820
rect -595 -840 -585 -820
rect -625 -870 -585 -840
rect -625 -890 -615 -870
rect -595 -890 -585 -870
rect -625 -920 -585 -890
rect -625 -940 -615 -920
rect -595 -940 -585 -920
rect -625 -970 -585 -940
rect -625 -990 -615 -970
rect -595 -990 -585 -970
rect -625 -1020 -585 -990
rect -625 -1040 -615 -1020
rect -595 -1040 -585 -1020
rect -625 -1055 -585 -1040
rect -525 -370 -485 -355
rect -525 -390 -515 -370
rect -495 -390 -485 -370
rect -525 -420 -485 -390
rect -525 -440 -515 -420
rect -495 -440 -485 -420
rect -525 -470 -485 -440
rect -525 -490 -515 -470
rect -495 -490 -485 -470
rect -525 -520 -485 -490
rect -525 -540 -515 -520
rect -495 -540 -485 -520
rect -525 -570 -485 -540
rect -525 -590 -515 -570
rect -495 -590 -485 -570
rect -525 -620 -485 -590
rect -525 -640 -515 -620
rect -495 -640 -485 -620
rect -525 -670 -485 -640
rect -525 -690 -515 -670
rect -495 -690 -485 -670
rect -525 -720 -485 -690
rect -525 -740 -515 -720
rect -495 -740 -485 -720
rect -525 -770 -485 -740
rect -525 -790 -515 -770
rect -495 -790 -485 -770
rect -525 -820 -485 -790
rect -525 -840 -515 -820
rect -495 -840 -485 -820
rect -525 -870 -485 -840
rect -525 -890 -515 -870
rect -495 -890 -485 -870
rect -525 -920 -485 -890
rect -525 -940 -515 -920
rect -495 -940 -485 -920
rect -525 -970 -485 -940
rect -525 -990 -515 -970
rect -495 -990 -485 -970
rect -525 -1020 -485 -990
rect -525 -1040 -515 -1020
rect -495 -1040 -485 -1020
rect -525 -1055 -485 -1040
rect -425 -370 -385 -355
rect -425 -390 -415 -370
rect -395 -390 -385 -370
rect 2075 -370 2115 -355
rect -425 -420 -385 -390
rect 2075 -390 2085 -370
rect 2105 -390 2115 -370
rect -425 -440 -415 -420
rect -395 -440 -385 -420
rect -425 -470 -385 -440
rect -425 -490 -415 -470
rect -395 -490 -385 -470
rect -425 -520 -385 -490
rect -425 -540 -415 -520
rect -395 -540 -385 -520
rect -425 -570 -385 -540
rect -425 -590 -415 -570
rect -395 -590 -385 -570
rect -425 -620 -385 -590
rect -425 -640 -415 -620
rect -395 -640 -385 -620
rect -425 -670 -385 -640
rect 160 -420 200 -405
rect 160 -440 170 -420
rect 190 -440 200 -420
rect 160 -470 200 -440
rect 160 -490 170 -470
rect 190 -490 200 -470
rect 160 -520 200 -490
rect 160 -540 170 -520
rect 190 -540 200 -520
rect 160 -570 200 -540
rect 160 -590 170 -570
rect 190 -590 200 -570
rect 160 -620 200 -590
rect 160 -640 170 -620
rect 190 -640 200 -620
rect 160 -655 200 -640
rect 215 -420 255 -405
rect 215 -440 225 -420
rect 245 -440 255 -420
rect 215 -470 255 -440
rect 215 -490 225 -470
rect 245 -490 255 -470
rect 215 -520 255 -490
rect 215 -540 225 -520
rect 245 -540 255 -520
rect 215 -570 255 -540
rect 215 -590 225 -570
rect 245 -590 255 -570
rect 215 -620 255 -590
rect 215 -640 225 -620
rect 245 -640 255 -620
rect 215 -655 255 -640
rect 270 -420 310 -405
rect 270 -440 280 -420
rect 300 -440 310 -420
rect 270 -470 310 -440
rect 270 -490 280 -470
rect 300 -490 310 -470
rect 270 -520 310 -490
rect 270 -540 280 -520
rect 300 -540 310 -520
rect 270 -570 310 -540
rect 270 -590 280 -570
rect 300 -590 310 -570
rect 270 -620 310 -590
rect 270 -640 280 -620
rect 300 -640 310 -620
rect 270 -655 310 -640
rect 325 -420 365 -405
rect 325 -440 335 -420
rect 355 -440 365 -420
rect 325 -470 365 -440
rect 325 -490 335 -470
rect 355 -490 365 -470
rect 325 -520 365 -490
rect 325 -540 335 -520
rect 355 -540 365 -520
rect 325 -570 365 -540
rect 325 -590 335 -570
rect 355 -590 365 -570
rect 325 -620 365 -590
rect 325 -640 335 -620
rect 355 -640 365 -620
rect 325 -655 365 -640
rect 380 -420 420 -405
rect 380 -440 390 -420
rect 410 -440 420 -420
rect 380 -470 420 -440
rect 380 -490 390 -470
rect 410 -490 420 -470
rect 380 -520 420 -490
rect 380 -540 390 -520
rect 410 -540 420 -520
rect 380 -570 420 -540
rect 380 -590 390 -570
rect 410 -590 420 -570
rect 380 -620 420 -590
rect 380 -640 390 -620
rect 410 -640 420 -620
rect 380 -655 420 -640
rect 435 -420 475 -405
rect 435 -440 445 -420
rect 465 -440 475 -420
rect 435 -470 475 -440
rect 435 -490 445 -470
rect 465 -490 475 -470
rect 435 -520 475 -490
rect 435 -540 445 -520
rect 465 -540 475 -520
rect 435 -570 475 -540
rect 435 -590 445 -570
rect 465 -590 475 -570
rect 435 -620 475 -590
rect 435 -640 445 -620
rect 465 -640 475 -620
rect 435 -655 475 -640
rect 490 -420 530 -405
rect 490 -440 500 -420
rect 520 -440 530 -420
rect 490 -470 530 -440
rect 490 -490 500 -470
rect 520 -490 530 -470
rect 490 -520 530 -490
rect 490 -540 500 -520
rect 520 -540 530 -520
rect 490 -570 530 -540
rect 490 -590 500 -570
rect 520 -590 530 -570
rect 490 -620 530 -590
rect 490 -640 500 -620
rect 520 -640 530 -620
rect 490 -655 530 -640
rect 545 -420 585 -405
rect 545 -440 555 -420
rect 575 -440 585 -420
rect 545 -470 585 -440
rect 545 -490 555 -470
rect 575 -490 585 -470
rect 545 -520 585 -490
rect 545 -540 555 -520
rect 575 -540 585 -520
rect 545 -570 585 -540
rect 545 -590 555 -570
rect 575 -590 585 -570
rect 545 -620 585 -590
rect 545 -640 555 -620
rect 575 -640 585 -620
rect 545 -655 585 -640
rect 600 -420 640 -405
rect 600 -440 610 -420
rect 630 -440 640 -420
rect 600 -470 640 -440
rect 600 -490 610 -470
rect 630 -490 640 -470
rect 600 -520 640 -490
rect 600 -540 610 -520
rect 630 -540 640 -520
rect 600 -570 640 -540
rect 600 -590 610 -570
rect 630 -590 640 -570
rect 600 -620 640 -590
rect 600 -640 610 -620
rect 630 -640 640 -620
rect 600 -655 640 -640
rect 655 -420 695 -405
rect 655 -440 665 -420
rect 685 -440 695 -420
rect 655 -470 695 -440
rect 655 -490 665 -470
rect 685 -490 695 -470
rect 655 -520 695 -490
rect 655 -540 665 -520
rect 685 -540 695 -520
rect 655 -570 695 -540
rect 655 -590 665 -570
rect 685 -590 695 -570
rect 655 -620 695 -590
rect 655 -640 665 -620
rect 685 -640 695 -620
rect 655 -655 695 -640
rect 710 -420 750 -405
rect 710 -440 720 -420
rect 740 -440 750 -420
rect 710 -470 750 -440
rect 710 -490 720 -470
rect 740 -490 750 -470
rect 710 -520 750 -490
rect 710 -540 720 -520
rect 740 -540 750 -520
rect 710 -570 750 -540
rect 710 -590 720 -570
rect 740 -590 750 -570
rect 710 -620 750 -590
rect 710 -640 720 -620
rect 740 -640 750 -620
rect 710 -655 750 -640
rect 765 -420 805 -405
rect 765 -440 775 -420
rect 795 -440 805 -420
rect 765 -470 805 -440
rect 765 -490 775 -470
rect 795 -490 805 -470
rect 765 -520 805 -490
rect 765 -540 775 -520
rect 795 -540 805 -520
rect 765 -570 805 -540
rect 765 -590 775 -570
rect 795 -590 805 -570
rect 765 -620 805 -590
rect 765 -640 775 -620
rect 795 -640 805 -620
rect 765 -655 805 -640
rect 820 -420 860 -405
rect 820 -440 830 -420
rect 850 -440 860 -420
rect 820 -470 860 -440
rect 820 -490 830 -470
rect 850 -490 860 -470
rect 820 -520 860 -490
rect 820 -540 830 -520
rect 850 -540 860 -520
rect 820 -570 860 -540
rect 820 -590 830 -570
rect 850 -590 860 -570
rect 820 -620 860 -590
rect 820 -640 830 -620
rect 850 -640 860 -620
rect 820 -655 860 -640
rect 875 -420 915 -405
rect 875 -440 885 -420
rect 905 -440 915 -420
rect 875 -470 915 -440
rect 875 -490 885 -470
rect 905 -490 915 -470
rect 875 -520 915 -490
rect 875 -540 885 -520
rect 905 -540 915 -520
rect 875 -570 915 -540
rect 875 -590 885 -570
rect 905 -590 915 -570
rect 875 -620 915 -590
rect 875 -640 885 -620
rect 905 -640 915 -620
rect 875 -655 915 -640
rect 930 -420 970 -405
rect 930 -440 940 -420
rect 960 -440 970 -420
rect 930 -470 970 -440
rect 930 -490 940 -470
rect 960 -490 970 -470
rect 930 -520 970 -490
rect 930 -540 940 -520
rect 960 -540 970 -520
rect 930 -570 970 -540
rect 930 -590 940 -570
rect 960 -590 970 -570
rect 930 -620 970 -590
rect 930 -640 940 -620
rect 960 -640 970 -620
rect 930 -655 970 -640
rect 985 -420 1025 -405
rect 985 -440 995 -420
rect 1015 -440 1025 -420
rect 985 -470 1025 -440
rect 985 -490 995 -470
rect 1015 -490 1025 -470
rect 985 -520 1025 -490
rect 985 -540 995 -520
rect 1015 -540 1025 -520
rect 985 -570 1025 -540
rect 985 -590 995 -570
rect 1015 -590 1025 -570
rect 985 -620 1025 -590
rect 985 -640 995 -620
rect 1015 -640 1025 -620
rect 985 -655 1025 -640
rect 1040 -420 1080 -405
rect 1040 -440 1050 -420
rect 1070 -440 1080 -420
rect 1040 -470 1080 -440
rect 1040 -490 1050 -470
rect 1070 -490 1080 -470
rect 1040 -520 1080 -490
rect 1040 -540 1050 -520
rect 1070 -540 1080 -520
rect 1040 -570 1080 -540
rect 1040 -590 1050 -570
rect 1070 -590 1080 -570
rect 1040 -620 1080 -590
rect 1040 -640 1050 -620
rect 1070 -640 1080 -620
rect 1040 -655 1080 -640
rect 1095 -420 1135 -405
rect 1095 -440 1105 -420
rect 1125 -440 1135 -420
rect 1095 -470 1135 -440
rect 1095 -490 1105 -470
rect 1125 -490 1135 -470
rect 1095 -520 1135 -490
rect 1095 -540 1105 -520
rect 1125 -540 1135 -520
rect 1095 -570 1135 -540
rect 1095 -590 1105 -570
rect 1125 -590 1135 -570
rect 1095 -620 1135 -590
rect 1095 -640 1105 -620
rect 1125 -640 1135 -620
rect 1095 -655 1135 -640
rect 1150 -420 1190 -405
rect 1150 -440 1160 -420
rect 1180 -440 1190 -420
rect 1150 -470 1190 -440
rect 1150 -490 1160 -470
rect 1180 -490 1190 -470
rect 1150 -520 1190 -490
rect 1150 -540 1160 -520
rect 1180 -540 1190 -520
rect 1150 -570 1190 -540
rect 1150 -590 1160 -570
rect 1180 -590 1190 -570
rect 1150 -620 1190 -590
rect 1150 -640 1160 -620
rect 1180 -640 1190 -620
rect 1150 -655 1190 -640
rect 1205 -420 1245 -405
rect 1205 -440 1215 -420
rect 1235 -440 1245 -420
rect 1205 -470 1245 -440
rect 1205 -490 1215 -470
rect 1235 -490 1245 -470
rect 1205 -520 1245 -490
rect 1205 -540 1215 -520
rect 1235 -540 1245 -520
rect 1205 -570 1245 -540
rect 1205 -590 1215 -570
rect 1235 -590 1245 -570
rect 1205 -620 1245 -590
rect 1205 -640 1215 -620
rect 1235 -640 1245 -620
rect 1205 -655 1245 -640
rect 1260 -420 1300 -405
rect 1260 -440 1270 -420
rect 1290 -440 1300 -420
rect 1260 -470 1300 -440
rect 1260 -490 1270 -470
rect 1290 -490 1300 -470
rect 1260 -520 1300 -490
rect 1260 -540 1270 -520
rect 1290 -540 1300 -520
rect 1260 -570 1300 -540
rect 1260 -590 1270 -570
rect 1290 -590 1300 -570
rect 1260 -620 1300 -590
rect 1260 -640 1270 -620
rect 1290 -640 1300 -620
rect 1260 -655 1300 -640
rect 1315 -420 1355 -405
rect 1315 -440 1325 -420
rect 1345 -440 1355 -420
rect 1315 -470 1355 -440
rect 1315 -490 1325 -470
rect 1345 -490 1355 -470
rect 1315 -520 1355 -490
rect 1315 -540 1325 -520
rect 1345 -540 1355 -520
rect 1315 -570 1355 -540
rect 1315 -590 1325 -570
rect 1345 -590 1355 -570
rect 1315 -620 1355 -590
rect 1315 -640 1325 -620
rect 1345 -640 1355 -620
rect 1315 -655 1355 -640
rect 1370 -420 1410 -405
rect 1370 -440 1380 -420
rect 1400 -440 1410 -420
rect 1370 -470 1410 -440
rect 1370 -490 1380 -470
rect 1400 -490 1410 -470
rect 1370 -520 1410 -490
rect 1370 -540 1380 -520
rect 1400 -540 1410 -520
rect 1370 -570 1410 -540
rect 1370 -590 1380 -570
rect 1400 -590 1410 -570
rect 1370 -620 1410 -590
rect 1370 -640 1380 -620
rect 1400 -640 1410 -620
rect 1370 -655 1410 -640
rect 1425 -420 1465 -405
rect 1425 -440 1435 -420
rect 1455 -440 1465 -420
rect 1425 -470 1465 -440
rect 1425 -490 1435 -470
rect 1455 -490 1465 -470
rect 1425 -520 1465 -490
rect 1425 -540 1435 -520
rect 1455 -540 1465 -520
rect 1425 -570 1465 -540
rect 1425 -590 1435 -570
rect 1455 -590 1465 -570
rect 1425 -620 1465 -590
rect 1425 -640 1435 -620
rect 1455 -640 1465 -620
rect 1425 -655 1465 -640
rect 2075 -420 2115 -390
rect 2075 -440 2085 -420
rect 2105 -440 2115 -420
rect 2075 -470 2115 -440
rect 2075 -490 2085 -470
rect 2105 -490 2115 -470
rect 2075 -520 2115 -490
rect 2075 -540 2085 -520
rect 2105 -540 2115 -520
rect 2075 -570 2115 -540
rect 2075 -590 2085 -570
rect 2105 -590 2115 -570
rect 2075 -620 2115 -590
rect 2075 -640 2085 -620
rect 2105 -640 2115 -620
rect 2075 -670 2115 -640
rect -425 -690 -415 -670
rect -395 -690 -385 -670
rect -425 -720 -385 -690
rect 2075 -690 2085 -670
rect 2105 -690 2115 -670
rect -425 -740 -415 -720
rect -395 -740 -385 -720
rect -425 -770 -385 -740
rect 2075 -720 2115 -690
rect 2075 -740 2085 -720
rect 2105 -740 2115 -720
rect -425 -790 -415 -770
rect -395 -790 -385 -770
rect -425 -820 -385 -790
rect 2075 -770 2115 -740
rect 2075 -790 2085 -770
rect 2105 -790 2115 -770
rect 2075 -820 2115 -790
rect -425 -840 -415 -820
rect -395 -840 -385 -820
rect -425 -870 -385 -840
rect -425 -890 -415 -870
rect -395 -890 -385 -870
rect -425 -920 -385 -890
rect 665 -835 705 -820
rect 665 -855 675 -835
rect 695 -855 705 -835
rect 665 -885 705 -855
rect 665 -905 675 -885
rect 695 -905 705 -885
rect 665 -920 705 -905
rect 995 -835 1035 -820
rect 995 -855 1005 -835
rect 1025 -855 1035 -835
rect 995 -885 1035 -855
rect 995 -905 1005 -885
rect 1025 -905 1035 -885
rect 995 -920 1035 -905
rect 2075 -840 2085 -820
rect 2105 -840 2115 -820
rect 2075 -870 2115 -840
rect 2075 -890 2085 -870
rect 2105 -890 2115 -870
rect 2075 -920 2115 -890
rect -425 -940 -415 -920
rect -395 -940 -385 -920
rect -425 -970 -385 -940
rect -425 -990 -415 -970
rect -395 -990 -385 -970
rect -425 -1020 -385 -990
rect -425 -1040 -415 -1020
rect -395 -1040 -385 -1020
rect -425 -1055 -385 -1040
rect 2075 -940 2085 -920
rect 2105 -940 2115 -920
rect 2075 -970 2115 -940
rect 2075 -990 2085 -970
rect 2105 -990 2115 -970
rect 2075 -1020 2115 -990
rect 2075 -1040 2085 -1020
rect 2105 -1040 2115 -1020
rect 2075 -1055 2115 -1040
rect 2175 -370 2215 -355
rect 2175 -390 2185 -370
rect 2205 -390 2215 -370
rect 2175 -420 2215 -390
rect 2175 -440 2185 -420
rect 2205 -440 2215 -420
rect 2175 -470 2215 -440
rect 2175 -490 2185 -470
rect 2205 -490 2215 -470
rect 2175 -520 2215 -490
rect 2175 -540 2185 -520
rect 2205 -540 2215 -520
rect 2175 -570 2215 -540
rect 2175 -590 2185 -570
rect 2205 -590 2215 -570
rect 2175 -620 2215 -590
rect 2175 -640 2185 -620
rect 2205 -640 2215 -620
rect 2175 -670 2215 -640
rect 2175 -690 2185 -670
rect 2205 -690 2215 -670
rect 2175 -720 2215 -690
rect 2175 -740 2185 -720
rect 2205 -740 2215 -720
rect 2175 -770 2215 -740
rect 2175 -790 2185 -770
rect 2205 -790 2215 -770
rect 2175 -820 2215 -790
rect 2175 -840 2185 -820
rect 2205 -840 2215 -820
rect 2175 -870 2215 -840
rect 2175 -890 2185 -870
rect 2205 -890 2215 -870
rect 2175 -920 2215 -890
rect 2175 -940 2185 -920
rect 2205 -940 2215 -920
rect 2175 -970 2215 -940
rect 2175 -990 2185 -970
rect 2205 -990 2215 -970
rect 2175 -1020 2215 -990
rect 2175 -1040 2185 -1020
rect 2205 -1040 2215 -1020
rect 2175 -1055 2215 -1040
rect 2275 -370 2315 -355
rect 2275 -390 2285 -370
rect 2305 -390 2315 -370
rect 2275 -420 2315 -390
rect 2275 -440 2285 -420
rect 2305 -440 2315 -420
rect 2275 -470 2315 -440
rect 2275 -490 2285 -470
rect 2305 -490 2315 -470
rect 2275 -520 2315 -490
rect 2275 -540 2285 -520
rect 2305 -540 2315 -520
rect 2275 -570 2315 -540
rect 2275 -590 2285 -570
rect 2305 -590 2315 -570
rect 2275 -620 2315 -590
rect 2275 -640 2285 -620
rect 2305 -640 2315 -620
rect 2275 -670 2315 -640
rect 2275 -690 2285 -670
rect 2305 -690 2315 -670
rect 2275 -720 2315 -690
rect 2275 -740 2285 -720
rect 2305 -740 2315 -720
rect 2275 -770 2315 -740
rect 2275 -790 2285 -770
rect 2305 -790 2315 -770
rect 2275 -820 2315 -790
rect 2275 -840 2285 -820
rect 2305 -840 2315 -820
rect 2275 -870 2315 -840
rect 2275 -890 2285 -870
rect 2305 -890 2315 -870
rect 2275 -920 2315 -890
rect 2275 -940 2285 -920
rect 2305 -940 2315 -920
rect 2275 -970 2315 -940
rect 2275 -990 2285 -970
rect 2305 -990 2315 -970
rect 2275 -1020 2315 -990
rect 2275 -1040 2285 -1020
rect 2305 -1040 2315 -1020
rect 2275 -1055 2315 -1040
rect 2375 -370 2415 -355
rect 2375 -390 2385 -370
rect 2405 -390 2415 -370
rect 2375 -420 2415 -390
rect 2375 -440 2385 -420
rect 2405 -440 2415 -420
rect 2375 -470 2415 -440
rect 2375 -490 2385 -470
rect 2405 -490 2415 -470
rect 2375 -520 2415 -490
rect 2375 -540 2385 -520
rect 2405 -540 2415 -520
rect 2375 -570 2415 -540
rect 2375 -590 2385 -570
rect 2405 -590 2415 -570
rect 2375 -620 2415 -590
rect 2375 -640 2385 -620
rect 2405 -640 2415 -620
rect 2375 -670 2415 -640
rect 2375 -690 2385 -670
rect 2405 -690 2415 -670
rect 2375 -720 2415 -690
rect 2375 -740 2385 -720
rect 2405 -740 2415 -720
rect 2375 -770 2415 -740
rect 2375 -790 2385 -770
rect 2405 -790 2415 -770
rect 2375 -820 2415 -790
rect 2375 -840 2385 -820
rect 2405 -840 2415 -820
rect 2375 -870 2415 -840
rect 2375 -890 2385 -870
rect 2405 -890 2415 -870
rect 2375 -920 2415 -890
rect 2375 -940 2385 -920
rect 2405 -940 2415 -920
rect 2375 -970 2415 -940
rect 2375 -990 2385 -970
rect 2405 -990 2415 -970
rect 2375 -1020 2415 -990
rect 2375 -1040 2385 -1020
rect 2405 -1040 2415 -1020
rect 2375 -1055 2415 -1040
rect 2475 -370 2515 -355
rect 2475 -390 2485 -370
rect 2505 -390 2515 -370
rect 2475 -420 2515 -390
rect 2475 -440 2485 -420
rect 2505 -440 2515 -420
rect 2475 -470 2515 -440
rect 2475 -490 2485 -470
rect 2505 -490 2515 -470
rect 2475 -520 2515 -490
rect 2475 -540 2485 -520
rect 2505 -540 2515 -520
rect 2475 -570 2515 -540
rect 2475 -590 2485 -570
rect 2505 -590 2515 -570
rect 2475 -620 2515 -590
rect 2475 -640 2485 -620
rect 2505 -640 2515 -620
rect 2475 -670 2515 -640
rect 2475 -690 2485 -670
rect 2505 -690 2515 -670
rect 2475 -720 2515 -690
rect 2475 -740 2485 -720
rect 2505 -740 2515 -720
rect 2475 -770 2515 -740
rect 2475 -790 2485 -770
rect 2505 -790 2515 -770
rect 2475 -820 2515 -790
rect 2475 -840 2485 -820
rect 2505 -840 2515 -820
rect 2475 -870 2515 -840
rect 2475 -890 2485 -870
rect 2505 -890 2515 -870
rect 2475 -920 2515 -890
rect 2475 -940 2485 -920
rect 2505 -940 2515 -920
rect 2475 -970 2515 -940
rect 2475 -990 2485 -970
rect 2505 -990 2515 -970
rect 2475 -1020 2515 -990
rect 2475 -1040 2485 -1020
rect 2505 -1040 2515 -1020
rect 2475 -1055 2515 -1040
rect 2575 -370 2615 -355
rect 2575 -390 2585 -370
rect 2605 -390 2615 -370
rect 2575 -420 2615 -390
rect 2575 -440 2585 -420
rect 2605 -440 2615 -420
rect 2575 -470 2615 -440
rect 2575 -490 2585 -470
rect 2605 -490 2615 -470
rect 2575 -520 2615 -490
rect 2575 -540 2585 -520
rect 2605 -540 2615 -520
rect 2575 -570 2615 -540
rect 2575 -590 2585 -570
rect 2605 -590 2615 -570
rect 2575 -620 2615 -590
rect 2575 -640 2585 -620
rect 2605 -640 2615 -620
rect 2575 -670 2615 -640
rect 2575 -690 2585 -670
rect 2605 -690 2615 -670
rect 2575 -720 2615 -690
rect 2575 -740 2585 -720
rect 2605 -740 2615 -720
rect 2575 -770 2615 -740
rect 2575 -790 2585 -770
rect 2605 -790 2615 -770
rect 2575 -820 2615 -790
rect 2575 -840 2585 -820
rect 2605 -840 2615 -820
rect 2575 -870 2615 -840
rect 2575 -890 2585 -870
rect 2605 -890 2615 -870
rect 2575 -920 2615 -890
rect 2575 -940 2585 -920
rect 2605 -940 2615 -920
rect 2575 -970 2615 -940
rect 2575 -990 2585 -970
rect 2605 -990 2615 -970
rect 2575 -1020 2615 -990
rect 2575 -1040 2585 -1020
rect 2605 -1040 2615 -1020
rect 2575 -1055 2615 -1040
rect 2675 -370 2715 -355
rect 2675 -390 2685 -370
rect 2705 -390 2715 -370
rect 2675 -420 2715 -390
rect 2675 -440 2685 -420
rect 2705 -440 2715 -420
rect 2675 -470 2715 -440
rect 2675 -490 2685 -470
rect 2705 -490 2715 -470
rect 2675 -520 2715 -490
rect 2675 -540 2685 -520
rect 2705 -540 2715 -520
rect 2675 -570 2715 -540
rect 2675 -590 2685 -570
rect 2705 -590 2715 -570
rect 2675 -620 2715 -590
rect 2675 -640 2685 -620
rect 2705 -640 2715 -620
rect 2675 -670 2715 -640
rect 2675 -690 2685 -670
rect 2705 -690 2715 -670
rect 2675 -720 2715 -690
rect 2675 -740 2685 -720
rect 2705 -740 2715 -720
rect 2675 -770 2715 -740
rect 2675 -790 2685 -770
rect 2705 -790 2715 -770
rect 2675 -820 2715 -790
rect 2675 -840 2685 -820
rect 2705 -840 2715 -820
rect 2675 -870 2715 -840
rect 2675 -890 2685 -870
rect 2705 -890 2715 -870
rect 2675 -920 2715 -890
rect 2675 -940 2685 -920
rect 2705 -940 2715 -920
rect 2675 -970 2715 -940
rect 2675 -990 2685 -970
rect 2705 -990 2715 -970
rect 2675 -1020 2715 -990
rect 2675 -1040 2685 -1020
rect 2705 -1040 2715 -1020
rect 2675 -1055 2715 -1040
<< pdiff >>
rect 30 2660 70 2675
rect 30 2640 40 2660
rect 60 2640 70 2660
rect 30 2610 70 2640
rect 30 2590 40 2610
rect 60 2590 70 2610
rect 30 2560 70 2590
rect 30 2540 40 2560
rect 60 2540 70 2560
rect 30 2510 70 2540
rect 30 2490 40 2510
rect 60 2490 70 2510
rect 30 2460 70 2490
rect 30 2440 40 2460
rect 60 2440 70 2460
rect 30 2410 70 2440
rect 30 2390 40 2410
rect 60 2390 70 2410
rect 30 2360 70 2390
rect 30 2340 40 2360
rect 60 2340 70 2360
rect 30 2325 70 2340
rect 90 2660 130 2675
rect 90 2640 100 2660
rect 120 2640 130 2660
rect 90 2610 130 2640
rect 90 2590 100 2610
rect 120 2590 130 2610
rect 90 2560 130 2590
rect 90 2540 100 2560
rect 120 2540 130 2560
rect 90 2510 130 2540
rect 90 2490 100 2510
rect 120 2490 130 2510
rect 90 2460 130 2490
rect 90 2440 100 2460
rect 120 2440 130 2460
rect 90 2410 130 2440
rect 90 2390 100 2410
rect 120 2390 130 2410
rect 90 2360 130 2390
rect 90 2340 100 2360
rect 120 2340 130 2360
rect 90 2325 130 2340
rect 150 2660 190 2675
rect 150 2640 160 2660
rect 180 2640 190 2660
rect 150 2610 190 2640
rect 150 2590 160 2610
rect 180 2590 190 2610
rect 150 2560 190 2590
rect 150 2540 160 2560
rect 180 2540 190 2560
rect 150 2510 190 2540
rect 150 2490 160 2510
rect 180 2490 190 2510
rect 150 2460 190 2490
rect 150 2440 160 2460
rect 180 2440 190 2460
rect 150 2410 190 2440
rect 150 2390 160 2410
rect 180 2390 190 2410
rect 150 2360 190 2390
rect 150 2340 160 2360
rect 180 2340 190 2360
rect 150 2325 190 2340
rect 210 2660 250 2675
rect 210 2640 220 2660
rect 240 2640 250 2660
rect 210 2610 250 2640
rect 210 2590 220 2610
rect 240 2590 250 2610
rect 210 2560 250 2590
rect 970 2660 1010 2675
rect 970 2640 980 2660
rect 1000 2640 1010 2660
rect 970 2610 1010 2640
rect 970 2590 980 2610
rect 1000 2590 1010 2610
rect 970 2560 1010 2590
rect 210 2540 220 2560
rect 240 2540 250 2560
rect 210 2510 250 2540
rect 970 2540 980 2560
rect 1000 2540 1010 2560
rect 210 2490 220 2510
rect 240 2490 250 2510
rect 970 2510 1010 2540
rect 210 2460 250 2490
rect 210 2440 220 2460
rect 240 2440 250 2460
rect 210 2410 250 2440
rect 210 2390 220 2410
rect 240 2390 250 2410
rect 210 2360 250 2390
rect 210 2340 220 2360
rect 240 2340 250 2360
rect 210 2325 250 2340
rect 500 2360 540 2505
rect 500 2340 510 2360
rect 530 2340 540 2360
rect 500 2325 540 2340
rect 560 2360 600 2505
rect 560 2340 570 2360
rect 590 2340 600 2360
rect 560 2325 600 2340
rect 620 2360 660 2505
rect 620 2340 630 2360
rect 650 2340 660 2360
rect 620 2325 660 2340
rect 680 2360 720 2505
rect 680 2340 690 2360
rect 710 2340 720 2360
rect 680 2325 720 2340
rect 970 2490 980 2510
rect 1000 2490 1010 2510
rect 970 2460 1010 2490
rect 970 2440 980 2460
rect 1000 2440 1010 2460
rect 970 2410 1010 2440
rect 970 2390 980 2410
rect 1000 2390 1010 2410
rect 970 2360 1010 2390
rect 970 2340 980 2360
rect 1000 2340 1010 2360
rect 970 2325 1010 2340
rect 1030 2660 1070 2675
rect 1030 2640 1040 2660
rect 1060 2640 1070 2660
rect 1030 2610 1070 2640
rect 1030 2590 1040 2610
rect 1060 2590 1070 2610
rect 1030 2560 1070 2590
rect 1030 2540 1040 2560
rect 1060 2540 1070 2560
rect 1030 2510 1070 2540
rect 1030 2490 1040 2510
rect 1060 2490 1070 2510
rect 1030 2460 1070 2490
rect 1030 2440 1040 2460
rect 1060 2440 1070 2460
rect 1030 2410 1070 2440
rect 1030 2390 1040 2410
rect 1060 2390 1070 2410
rect 1030 2360 1070 2390
rect 1030 2340 1040 2360
rect 1060 2340 1070 2360
rect 1030 2325 1070 2340
rect 1090 2660 1130 2675
rect 1090 2640 1100 2660
rect 1120 2640 1130 2660
rect 1090 2610 1130 2640
rect 1090 2590 1100 2610
rect 1120 2590 1130 2610
rect 1090 2560 1130 2590
rect 1090 2540 1100 2560
rect 1120 2540 1130 2560
rect 1090 2510 1130 2540
rect 1090 2490 1100 2510
rect 1120 2490 1130 2510
rect 1090 2460 1130 2490
rect 1090 2440 1100 2460
rect 1120 2440 1130 2460
rect 1090 2410 1130 2440
rect 1090 2390 1100 2410
rect 1120 2390 1130 2410
rect 1090 2360 1130 2390
rect 1090 2340 1100 2360
rect 1120 2340 1130 2360
rect 1090 2325 1130 2340
rect 1150 2660 1190 2675
rect 1150 2640 1160 2660
rect 1180 2640 1190 2660
rect 1150 2610 1190 2640
rect 1150 2590 1160 2610
rect 1180 2590 1190 2610
rect 1150 2560 1190 2590
rect 1150 2540 1160 2560
rect 1180 2540 1190 2560
rect 1150 2510 1190 2540
rect 1150 2490 1160 2510
rect 1180 2490 1190 2510
rect 1150 2460 1190 2490
rect 1150 2440 1160 2460
rect 1180 2440 1190 2460
rect 1150 2410 1190 2440
rect 1150 2390 1160 2410
rect 1180 2390 1190 2410
rect 1150 2360 1190 2390
rect 1150 2340 1160 2360
rect 1180 2340 1190 2360
rect 1150 2325 1190 2340
rect 1438 2660 1478 2675
rect 1438 2640 1448 2660
rect 1468 2640 1478 2660
rect 1438 2610 1478 2640
rect 1438 2590 1448 2610
rect 1468 2590 1478 2610
rect 1438 2560 1478 2590
rect 1438 2540 1448 2560
rect 1468 2540 1478 2560
rect 1438 2510 1478 2540
rect 1438 2490 1448 2510
rect 1468 2490 1478 2510
rect 1438 2460 1478 2490
rect 1438 2440 1448 2460
rect 1468 2440 1478 2460
rect 1438 2410 1478 2440
rect 1438 2390 1448 2410
rect 1468 2390 1478 2410
rect 1438 2360 1478 2390
rect 1438 2340 1448 2360
rect 1468 2340 1478 2360
rect 1438 2325 1478 2340
rect 1498 2660 1538 2675
rect 1498 2640 1508 2660
rect 1528 2640 1538 2660
rect 1498 2610 1538 2640
rect 1498 2590 1508 2610
rect 1528 2590 1538 2610
rect 1498 2560 1538 2590
rect 1498 2540 1508 2560
rect 1528 2540 1538 2560
rect 1498 2510 1538 2540
rect 1498 2490 1508 2510
rect 1528 2490 1538 2510
rect 1498 2460 1538 2490
rect 1498 2440 1508 2460
rect 1528 2440 1538 2460
rect 1498 2410 1538 2440
rect 1498 2390 1508 2410
rect 1528 2390 1538 2410
rect 1498 2360 1538 2390
rect 1498 2340 1508 2360
rect 1528 2340 1538 2360
rect 1498 2325 1538 2340
rect 1558 2660 1598 2675
rect 1558 2640 1568 2660
rect 1588 2640 1598 2660
rect 1558 2610 1598 2640
rect 1558 2590 1568 2610
rect 1588 2590 1598 2610
rect 1558 2560 1598 2590
rect 1558 2540 1568 2560
rect 1588 2540 1598 2560
rect 1558 2510 1598 2540
rect 1558 2490 1568 2510
rect 1588 2490 1598 2510
rect 1558 2460 1598 2490
rect 1558 2440 1568 2460
rect 1588 2440 1598 2460
rect 1558 2410 1598 2440
rect 1558 2390 1568 2410
rect 1588 2390 1598 2410
rect 1558 2360 1598 2390
rect 1558 2340 1568 2360
rect 1588 2340 1598 2360
rect 1558 2325 1598 2340
rect 1618 2660 1658 2675
rect 1618 2640 1628 2660
rect 1648 2640 1658 2660
rect 1618 2610 1658 2640
rect 1618 2590 1628 2610
rect 1648 2590 1658 2610
rect 1618 2560 1658 2590
rect 1618 2540 1628 2560
rect 1648 2540 1658 2560
rect 1618 2510 1658 2540
rect 1618 2490 1628 2510
rect 1648 2490 1658 2510
rect 1618 2460 1658 2490
rect 1618 2440 1628 2460
rect 1648 2440 1658 2460
rect 1618 2410 1658 2440
rect 1618 2390 1628 2410
rect 1648 2390 1658 2410
rect 1618 2360 1658 2390
rect 1618 2340 1628 2360
rect 1648 2340 1658 2360
rect 1618 2325 1658 2340
rect -1085 2085 -1045 2100
rect -1085 2065 -1075 2085
rect -1055 2065 -1045 2085
rect -1085 2035 -1045 2065
rect -1085 2015 -1075 2035
rect -1055 2015 -1045 2035
rect -1085 1985 -1045 2015
rect -1085 1965 -1075 1985
rect -1055 1965 -1045 1985
rect -1085 1935 -1045 1965
rect -1085 1915 -1075 1935
rect -1055 1915 -1045 1935
rect -1085 1885 -1045 1915
rect -1085 1865 -1075 1885
rect -1055 1865 -1045 1885
rect -1085 1835 -1045 1865
rect -1085 1815 -1075 1835
rect -1055 1815 -1045 1835
rect -1085 1785 -1045 1815
rect -1085 1765 -1075 1785
rect -1055 1765 -1045 1785
rect -1085 1750 -1045 1765
rect -1025 2085 -985 2100
rect -1025 2065 -1015 2085
rect -995 2065 -985 2085
rect -1025 2035 -985 2065
rect -1025 2015 -1015 2035
rect -995 2015 -985 2035
rect -1025 1985 -985 2015
rect -1025 1965 -1015 1985
rect -995 1965 -985 1985
rect -1025 1935 -985 1965
rect -1025 1915 -1015 1935
rect -995 1915 -985 1935
rect -1025 1885 -985 1915
rect -1025 1865 -1015 1885
rect -995 1865 -985 1885
rect -1025 1835 -985 1865
rect -1025 1815 -1015 1835
rect -995 1815 -985 1835
rect -1025 1785 -985 1815
rect -1025 1765 -1015 1785
rect -995 1765 -985 1785
rect -1025 1750 -985 1765
rect -965 2085 -925 2100
rect -965 2065 -955 2085
rect -935 2065 -925 2085
rect -965 2035 -925 2065
rect -965 2015 -955 2035
rect -935 2015 -925 2035
rect -965 1985 -925 2015
rect -965 1965 -955 1985
rect -935 1965 -925 1985
rect -965 1935 -925 1965
rect -965 1915 -955 1935
rect -935 1915 -925 1935
rect -965 1885 -925 1915
rect -965 1865 -955 1885
rect -935 1865 -925 1885
rect -965 1835 -925 1865
rect -965 1815 -955 1835
rect -935 1815 -925 1835
rect -965 1785 -925 1815
rect -965 1765 -955 1785
rect -935 1765 -925 1785
rect -965 1750 -925 1765
rect -905 2085 -865 2100
rect -905 2065 -895 2085
rect -875 2065 -865 2085
rect -905 2035 -865 2065
rect -905 2015 -895 2035
rect -875 2015 -865 2035
rect -905 1985 -865 2015
rect -905 1965 -895 1985
rect -875 1965 -865 1985
rect -905 1935 -865 1965
rect -905 1915 -895 1935
rect -875 1915 -865 1935
rect -905 1885 -865 1915
rect -905 1865 -895 1885
rect -875 1865 -865 1885
rect -905 1835 -865 1865
rect -905 1815 -895 1835
rect -875 1815 -865 1835
rect -905 1785 -865 1815
rect -905 1765 -895 1785
rect -875 1765 -865 1785
rect -905 1750 -865 1765
rect -845 2085 -805 2100
rect -845 2065 -835 2085
rect -815 2065 -805 2085
rect -845 2035 -805 2065
rect -845 2015 -835 2035
rect -815 2015 -805 2035
rect -845 1985 -805 2015
rect -845 1965 -835 1985
rect -815 1965 -805 1985
rect -845 1935 -805 1965
rect -845 1915 -835 1935
rect -815 1915 -805 1935
rect -845 1885 -805 1915
rect -845 1865 -835 1885
rect -815 1865 -805 1885
rect -845 1835 -805 1865
rect -845 1815 -835 1835
rect -815 1815 -805 1835
rect -845 1785 -805 1815
rect -845 1765 -835 1785
rect -815 1765 -805 1785
rect -845 1750 -805 1765
rect -785 2085 -745 2100
rect -785 2065 -775 2085
rect -755 2065 -745 2085
rect -785 2035 -745 2065
rect -785 2015 -775 2035
rect -755 2015 -745 2035
rect -785 1985 -745 2015
rect -785 1965 -775 1985
rect -755 1965 -745 1985
rect -785 1935 -745 1965
rect -785 1915 -775 1935
rect -755 1915 -745 1935
rect -785 1885 -745 1915
rect -785 1865 -775 1885
rect -755 1865 -745 1885
rect -785 1835 -745 1865
rect -785 1815 -775 1835
rect -755 1815 -745 1835
rect -785 1785 -745 1815
rect -785 1765 -775 1785
rect -755 1765 -745 1785
rect -785 1750 -745 1765
rect -725 2085 -685 2100
rect -725 2065 -715 2085
rect -695 2065 -685 2085
rect -725 2035 -685 2065
rect -725 2015 -715 2035
rect -695 2015 -685 2035
rect -725 1985 -685 2015
rect -725 1965 -715 1985
rect -695 1965 -685 1985
rect -725 1935 -685 1965
rect -725 1915 -715 1935
rect -695 1915 -685 1935
rect -725 1885 -685 1915
rect -725 1865 -715 1885
rect -695 1865 -685 1885
rect -725 1835 -685 1865
rect -725 1815 -715 1835
rect -695 1815 -685 1835
rect -725 1785 -685 1815
rect -725 1765 -715 1785
rect -695 1765 -685 1785
rect -725 1750 -685 1765
rect -665 2085 -625 2100
rect -665 2065 -655 2085
rect -635 2065 -625 2085
rect -665 2035 -625 2065
rect -665 2015 -655 2035
rect -635 2015 -625 2035
rect -665 1985 -625 2015
rect -665 1965 -655 1985
rect -635 1965 -625 1985
rect -665 1935 -625 1965
rect -665 1915 -655 1935
rect -635 1915 -625 1935
rect -665 1885 -625 1915
rect -665 1865 -655 1885
rect -635 1865 -625 1885
rect -665 1835 -625 1865
rect -665 1815 -655 1835
rect -635 1815 -625 1835
rect -665 1785 -625 1815
rect -665 1765 -655 1785
rect -635 1765 -625 1785
rect -665 1750 -625 1765
rect -605 2085 -565 2100
rect -605 2065 -595 2085
rect -575 2065 -565 2085
rect -605 2035 -565 2065
rect -605 2015 -595 2035
rect -575 2015 -565 2035
rect -605 1985 -565 2015
rect -605 1965 -595 1985
rect -575 1965 -565 1985
rect -605 1935 -565 1965
rect -605 1915 -595 1935
rect -575 1915 -565 1935
rect -605 1885 -565 1915
rect -605 1865 -595 1885
rect -575 1865 -565 1885
rect -605 1835 -565 1865
rect -605 1815 -595 1835
rect -575 1815 -565 1835
rect -605 1785 -565 1815
rect -605 1765 -595 1785
rect -575 1765 -565 1785
rect -605 1750 -565 1765
rect -545 2085 -505 2100
rect -545 2065 -535 2085
rect -515 2065 -505 2085
rect -545 2035 -505 2065
rect -545 2015 -535 2035
rect -515 2015 -505 2035
rect -545 1985 -505 2015
rect -545 1965 -535 1985
rect -515 1965 -505 1985
rect -545 1935 -505 1965
rect -545 1915 -535 1935
rect -515 1915 -505 1935
rect -545 1885 -505 1915
rect -545 1865 -535 1885
rect -515 1865 -505 1885
rect -545 1835 -505 1865
rect -545 1815 -535 1835
rect -515 1815 -505 1835
rect -545 1785 -505 1815
rect -545 1765 -535 1785
rect -515 1765 -505 1785
rect -545 1750 -505 1765
rect -485 2085 -445 2100
rect -485 2065 -475 2085
rect -455 2065 -445 2085
rect -485 2035 -445 2065
rect -485 2015 -475 2035
rect -455 2015 -445 2035
rect -485 1985 -445 2015
rect -485 1965 -475 1985
rect -455 1965 -445 1985
rect -485 1935 -445 1965
rect -485 1915 -475 1935
rect -455 1915 -445 1935
rect -485 1885 -445 1915
rect -485 1865 -475 1885
rect -455 1865 -445 1885
rect -485 1835 -445 1865
rect -485 1815 -475 1835
rect -455 1815 -445 1835
rect -485 1785 -445 1815
rect -485 1765 -475 1785
rect -455 1765 -445 1785
rect -485 1750 -445 1765
rect -425 2085 -385 2100
rect -425 2065 -415 2085
rect -395 2065 -385 2085
rect -425 2035 -385 2065
rect -425 2015 -415 2035
rect -395 2015 -385 2035
rect -425 1985 -385 2015
rect -425 1965 -415 1985
rect -395 1965 -385 1985
rect -425 1935 -385 1965
rect -425 1915 -415 1935
rect -395 1915 -385 1935
rect -425 1885 -385 1915
rect -425 1865 -415 1885
rect -395 1865 -385 1885
rect -425 1835 -385 1865
rect -425 1815 -415 1835
rect -395 1815 -385 1835
rect -425 1785 -385 1815
rect -425 1765 -415 1785
rect -395 1765 -385 1785
rect -425 1750 -385 1765
rect -365 2085 -325 2100
rect -365 2065 -355 2085
rect -335 2065 -325 2085
rect -365 2035 -325 2065
rect -365 2015 -355 2035
rect -335 2015 -325 2035
rect -365 1985 -325 2015
rect -365 1965 -355 1985
rect -335 1965 -325 1985
rect -365 1935 -325 1965
rect -365 1915 -355 1935
rect -335 1915 -325 1935
rect -365 1885 -325 1915
rect -365 1865 -355 1885
rect -335 1865 -325 1885
rect -365 1835 -325 1865
rect -365 1815 -355 1835
rect -335 1815 -325 1835
rect -365 1785 -325 1815
rect -365 1765 -355 1785
rect -335 1765 -325 1785
rect -365 1750 -325 1765
rect -40 2085 0 2100
rect -40 2065 -30 2085
rect -10 2065 0 2085
rect -40 2035 0 2065
rect -40 2015 -30 2035
rect -10 2015 0 2035
rect -40 1985 0 2015
rect -40 1965 -30 1985
rect -10 1965 0 1985
rect -40 1935 0 1965
rect -40 1915 -30 1935
rect -10 1915 0 1935
rect -40 1885 0 1915
rect -40 1865 -30 1885
rect -10 1865 0 1885
rect -40 1835 0 1865
rect -40 1815 -30 1835
rect -10 1815 0 1835
rect -40 1785 0 1815
rect -40 1765 -30 1785
rect -10 1765 0 1785
rect -40 1750 0 1765
rect 20 2085 60 2100
rect 20 2065 30 2085
rect 50 2065 60 2085
rect 20 2035 60 2065
rect 20 2015 30 2035
rect 50 2015 60 2035
rect 20 1985 60 2015
rect 20 1965 30 1985
rect 50 1965 60 1985
rect 20 1935 60 1965
rect 20 1915 30 1935
rect 50 1915 60 1935
rect 20 1885 60 1915
rect 20 1865 30 1885
rect 50 1865 60 1885
rect 20 1835 60 1865
rect 20 1815 30 1835
rect 50 1815 60 1835
rect 20 1785 60 1815
rect 20 1765 30 1785
rect 50 1765 60 1785
rect 20 1750 60 1765
rect 80 2085 120 2100
rect 80 2065 90 2085
rect 110 2065 120 2085
rect 80 2035 120 2065
rect 80 2015 90 2035
rect 110 2015 120 2035
rect 80 1985 120 2015
rect 80 1965 90 1985
rect 110 1965 120 1985
rect 80 1935 120 1965
rect 80 1915 90 1935
rect 110 1915 120 1935
rect 80 1885 120 1915
rect 80 1865 90 1885
rect 110 1865 120 1885
rect 80 1835 120 1865
rect 80 1815 90 1835
rect 110 1815 120 1835
rect 80 1785 120 1815
rect 80 1765 90 1785
rect 110 1765 120 1785
rect 80 1750 120 1765
rect 140 2085 180 2100
rect 140 2065 150 2085
rect 170 2065 180 2085
rect 140 2035 180 2065
rect 140 2015 150 2035
rect 170 2015 180 2035
rect 140 1985 180 2015
rect 140 1965 150 1985
rect 170 1965 180 1985
rect 140 1935 180 1965
rect 140 1915 150 1935
rect 170 1915 180 1935
rect 140 1885 180 1915
rect 140 1865 150 1885
rect 170 1865 180 1885
rect 140 1835 180 1865
rect 140 1815 150 1835
rect 170 1815 180 1835
rect 140 1785 180 1815
rect 140 1765 150 1785
rect 170 1765 180 1785
rect 140 1750 180 1765
rect 200 2085 240 2100
rect 200 2065 210 2085
rect 230 2065 240 2085
rect 200 2035 240 2065
rect 200 2015 210 2035
rect 230 2015 240 2035
rect 200 1985 240 2015
rect 200 1965 210 1985
rect 230 1965 240 1985
rect 200 1935 240 1965
rect 200 1915 210 1935
rect 230 1915 240 1935
rect 200 1885 240 1915
rect 200 1865 210 1885
rect 230 1865 240 1885
rect 200 1835 240 1865
rect 200 1815 210 1835
rect 230 1815 240 1835
rect 200 1785 240 1815
rect 200 1765 210 1785
rect 230 1765 240 1785
rect 200 1750 240 1765
rect 260 2085 300 2100
rect 260 2065 270 2085
rect 290 2065 300 2085
rect 260 2035 300 2065
rect 260 2015 270 2035
rect 290 2015 300 2035
rect 260 1985 300 2015
rect 260 1965 270 1985
rect 290 1965 300 1985
rect 260 1935 300 1965
rect 260 1915 270 1935
rect 290 1915 300 1935
rect 260 1885 300 1915
rect 260 1865 270 1885
rect 290 1865 300 1885
rect 260 1835 300 1865
rect 260 1815 270 1835
rect 290 1815 300 1835
rect 260 1785 300 1815
rect 260 1765 270 1785
rect 290 1765 300 1785
rect 260 1750 300 1765
rect 320 2085 360 2100
rect 320 2065 330 2085
rect 350 2065 360 2085
rect 320 2035 360 2065
rect 320 2015 330 2035
rect 350 2015 360 2035
rect 320 1985 360 2015
rect 320 1965 330 1985
rect 350 1965 360 1985
rect 320 1935 360 1965
rect 320 1915 330 1935
rect 350 1915 360 1935
rect 320 1885 360 1915
rect 320 1865 330 1885
rect 350 1865 360 1885
rect 320 1835 360 1865
rect 320 1815 330 1835
rect 350 1815 360 1835
rect 320 1785 360 1815
rect 320 1765 330 1785
rect 350 1765 360 1785
rect 320 1750 360 1765
rect 380 2085 420 2100
rect 380 2065 390 2085
rect 410 2065 420 2085
rect 380 2035 420 2065
rect 380 2015 390 2035
rect 410 2015 420 2035
rect 380 1985 420 2015
rect 380 1965 390 1985
rect 410 1965 420 1985
rect 380 1935 420 1965
rect 380 1915 390 1935
rect 410 1915 420 1935
rect 380 1885 420 1915
rect 380 1865 390 1885
rect 410 1865 420 1885
rect 380 1835 420 1865
rect 380 1815 390 1835
rect 410 1815 420 1835
rect 380 1785 420 1815
rect 380 1765 390 1785
rect 410 1765 420 1785
rect 380 1750 420 1765
rect 440 2085 480 2100
rect 440 2065 450 2085
rect 470 2065 480 2085
rect 440 2035 480 2065
rect 440 2015 450 2035
rect 470 2015 480 2035
rect 440 1985 480 2015
rect 440 1965 450 1985
rect 470 1965 480 1985
rect 440 1935 480 1965
rect 440 1915 450 1935
rect 470 1915 480 1935
rect 440 1885 480 1915
rect 440 1865 450 1885
rect 470 1865 480 1885
rect 440 1835 480 1865
rect 440 1815 450 1835
rect 470 1815 480 1835
rect 440 1785 480 1815
rect 440 1765 450 1785
rect 470 1765 480 1785
rect 440 1750 480 1765
rect 500 2085 540 2100
rect 500 2065 510 2085
rect 530 2065 540 2085
rect 500 2035 540 2065
rect 500 2015 510 2035
rect 530 2015 540 2035
rect 500 1985 540 2015
rect 500 1965 510 1985
rect 530 1965 540 1985
rect 500 1935 540 1965
rect 500 1915 510 1935
rect 530 1915 540 1935
rect 500 1885 540 1915
rect 500 1865 510 1885
rect 530 1865 540 1885
rect 500 1835 540 1865
rect 500 1815 510 1835
rect 530 1815 540 1835
rect 500 1785 540 1815
rect 500 1765 510 1785
rect 530 1765 540 1785
rect 500 1750 540 1765
rect 560 2085 600 2100
rect 560 2065 570 2085
rect 590 2065 600 2085
rect 560 2035 600 2065
rect 560 2015 570 2035
rect 590 2015 600 2035
rect 560 1985 600 2015
rect 560 1965 570 1985
rect 590 1965 600 1985
rect 560 1935 600 1965
rect 560 1915 570 1935
rect 590 1915 600 1935
rect 560 1885 600 1915
rect 560 1865 570 1885
rect 590 1865 600 1885
rect 560 1835 600 1865
rect 560 1815 570 1835
rect 590 1815 600 1835
rect 560 1785 600 1815
rect 560 1765 570 1785
rect 590 1765 600 1785
rect 560 1750 600 1765
rect 620 2085 660 2100
rect 620 2065 630 2085
rect 650 2065 660 2085
rect 620 2035 660 2065
rect 620 2015 630 2035
rect 650 2015 660 2035
rect 620 1985 660 2015
rect 620 1965 630 1985
rect 650 1965 660 1985
rect 620 1935 660 1965
rect 620 1915 630 1935
rect 650 1915 660 1935
rect 620 1885 660 1915
rect 620 1865 630 1885
rect 650 1865 660 1885
rect 620 1835 660 1865
rect 620 1815 630 1835
rect 650 1815 660 1835
rect 620 1785 660 1815
rect 620 1765 630 1785
rect 650 1765 660 1785
rect 620 1750 660 1765
rect 680 2085 720 2100
rect 680 2065 690 2085
rect 710 2065 720 2085
rect 680 2035 720 2065
rect 680 2015 690 2035
rect 710 2015 720 2035
rect 680 1985 720 2015
rect 680 1965 690 1985
rect 710 1965 720 1985
rect 680 1935 720 1965
rect 680 1915 690 1935
rect 710 1915 720 1935
rect 680 1885 720 1915
rect 680 1865 690 1885
rect 710 1865 720 1885
rect 680 1835 720 1865
rect 680 1815 690 1835
rect 710 1815 720 1835
rect 680 1785 720 1815
rect 680 1765 690 1785
rect 710 1765 720 1785
rect 680 1750 720 1765
rect 970 2085 1010 2100
rect 970 2065 980 2085
rect 1000 2065 1010 2085
rect 970 2035 1010 2065
rect 970 2015 980 2035
rect 1000 2015 1010 2035
rect 970 1985 1010 2015
rect 970 1965 980 1985
rect 1000 1965 1010 1985
rect 970 1935 1010 1965
rect 970 1915 980 1935
rect 1000 1915 1010 1935
rect 970 1885 1010 1915
rect 970 1865 980 1885
rect 1000 1865 1010 1885
rect 970 1835 1010 1865
rect 970 1815 980 1835
rect 1000 1815 1010 1835
rect 970 1785 1010 1815
rect 970 1765 980 1785
rect 1000 1765 1010 1785
rect 970 1750 1010 1765
rect 1030 2085 1070 2100
rect 1030 2065 1040 2085
rect 1060 2065 1070 2085
rect 1030 2035 1070 2065
rect 1030 2015 1040 2035
rect 1060 2015 1070 2035
rect 1030 1985 1070 2015
rect 1030 1965 1040 1985
rect 1060 1965 1070 1985
rect 1030 1935 1070 1965
rect 1030 1915 1040 1935
rect 1060 1915 1070 1935
rect 1030 1885 1070 1915
rect 1030 1865 1040 1885
rect 1060 1865 1070 1885
rect 1030 1835 1070 1865
rect 1030 1815 1040 1835
rect 1060 1815 1070 1835
rect 1030 1785 1070 1815
rect 1030 1765 1040 1785
rect 1060 1765 1070 1785
rect 1030 1750 1070 1765
rect 1090 2085 1130 2100
rect 1090 2065 1100 2085
rect 1120 2065 1130 2085
rect 1090 2035 1130 2065
rect 1090 2015 1100 2035
rect 1120 2015 1130 2035
rect 1090 1985 1130 2015
rect 1090 1965 1100 1985
rect 1120 1965 1130 1985
rect 1090 1935 1130 1965
rect 1090 1915 1100 1935
rect 1120 1915 1130 1935
rect 1090 1885 1130 1915
rect 1090 1865 1100 1885
rect 1120 1865 1130 1885
rect 1090 1835 1130 1865
rect 1090 1815 1100 1835
rect 1120 1815 1130 1835
rect 1090 1785 1130 1815
rect 1090 1765 1100 1785
rect 1120 1765 1130 1785
rect 1090 1750 1130 1765
rect 1150 2085 1190 2100
rect 1150 2065 1160 2085
rect 1180 2065 1190 2085
rect 1150 2035 1190 2065
rect 1150 2015 1160 2035
rect 1180 2015 1190 2035
rect 1150 1985 1190 2015
rect 1150 1965 1160 1985
rect 1180 1965 1190 1985
rect 1150 1935 1190 1965
rect 1150 1915 1160 1935
rect 1180 1915 1190 1935
rect 1150 1885 1190 1915
rect 1150 1865 1160 1885
rect 1180 1865 1190 1885
rect 1150 1835 1190 1865
rect 1150 1815 1160 1835
rect 1180 1815 1190 1835
rect 1150 1785 1190 1815
rect 1150 1765 1160 1785
rect 1180 1765 1190 1785
rect 1150 1750 1190 1765
rect 1210 2085 1250 2100
rect 1210 2065 1220 2085
rect 1240 2065 1250 2085
rect 1210 2035 1250 2065
rect 1210 2015 1220 2035
rect 1240 2015 1250 2035
rect 1210 1985 1250 2015
rect 1210 1965 1220 1985
rect 1240 1965 1250 1985
rect 1210 1935 1250 1965
rect 1210 1915 1220 1935
rect 1240 1915 1250 1935
rect 1210 1885 1250 1915
rect 1210 1865 1220 1885
rect 1240 1865 1250 1885
rect 1210 1835 1250 1865
rect 1210 1815 1220 1835
rect 1240 1815 1250 1835
rect 1210 1785 1250 1815
rect 1210 1765 1220 1785
rect 1240 1765 1250 1785
rect 1210 1750 1250 1765
rect 1270 2085 1310 2100
rect 1270 2065 1280 2085
rect 1300 2065 1310 2085
rect 1270 2035 1310 2065
rect 1270 2015 1280 2035
rect 1300 2015 1310 2035
rect 1270 1985 1310 2015
rect 1270 1965 1280 1985
rect 1300 1965 1310 1985
rect 1270 1935 1310 1965
rect 1270 1915 1280 1935
rect 1300 1915 1310 1935
rect 1270 1885 1310 1915
rect 1270 1865 1280 1885
rect 1300 1865 1310 1885
rect 1270 1835 1310 1865
rect 1270 1815 1280 1835
rect 1300 1815 1310 1835
rect 1270 1785 1310 1815
rect 1270 1765 1280 1785
rect 1300 1765 1310 1785
rect 1270 1750 1310 1765
rect 1330 2085 1370 2100
rect 1330 2065 1340 2085
rect 1360 2065 1370 2085
rect 1330 2035 1370 2065
rect 1330 2015 1340 2035
rect 1360 2015 1370 2035
rect 1330 1985 1370 2015
rect 1330 1965 1340 1985
rect 1360 1965 1370 1985
rect 1330 1935 1370 1965
rect 1330 1915 1340 1935
rect 1360 1915 1370 1935
rect 1330 1885 1370 1915
rect 1330 1865 1340 1885
rect 1360 1865 1370 1885
rect 1330 1835 1370 1865
rect 1330 1815 1340 1835
rect 1360 1815 1370 1835
rect 1330 1785 1370 1815
rect 1330 1765 1340 1785
rect 1360 1765 1370 1785
rect 1330 1750 1370 1765
rect 1390 2085 1430 2100
rect 1390 2065 1400 2085
rect 1420 2065 1430 2085
rect 1390 2035 1430 2065
rect 1390 2015 1400 2035
rect 1420 2015 1430 2035
rect 1390 1985 1430 2015
rect 1390 1965 1400 1985
rect 1420 1965 1430 1985
rect 1390 1935 1430 1965
rect 1390 1915 1400 1935
rect 1420 1915 1430 1935
rect 1390 1885 1430 1915
rect 1390 1865 1400 1885
rect 1420 1865 1430 1885
rect 1390 1835 1430 1865
rect 1390 1815 1400 1835
rect 1420 1815 1430 1835
rect 1390 1785 1430 1815
rect 1390 1765 1400 1785
rect 1420 1765 1430 1785
rect 1390 1750 1430 1765
rect 1450 2085 1490 2100
rect 1450 2065 1460 2085
rect 1480 2065 1490 2085
rect 1450 2035 1490 2065
rect 1450 2015 1460 2035
rect 1480 2015 1490 2035
rect 1450 1985 1490 2015
rect 1450 1965 1460 1985
rect 1480 1965 1490 1985
rect 1450 1935 1490 1965
rect 1450 1915 1460 1935
rect 1480 1915 1490 1935
rect 1450 1885 1490 1915
rect 1450 1865 1460 1885
rect 1480 1865 1490 1885
rect 1450 1835 1490 1865
rect 1450 1815 1460 1835
rect 1480 1815 1490 1835
rect 1450 1785 1490 1815
rect 1450 1765 1460 1785
rect 1480 1765 1490 1785
rect 1450 1750 1490 1765
rect 1510 2085 1550 2100
rect 1510 2065 1520 2085
rect 1540 2065 1550 2085
rect 1510 2035 1550 2065
rect 1510 2015 1520 2035
rect 1540 2015 1550 2035
rect 1510 1985 1550 2015
rect 1510 1965 1520 1985
rect 1540 1965 1550 1985
rect 1510 1935 1550 1965
rect 1510 1915 1520 1935
rect 1540 1915 1550 1935
rect 1510 1885 1550 1915
rect 1510 1865 1520 1885
rect 1540 1865 1550 1885
rect 1510 1835 1550 1865
rect 1510 1815 1520 1835
rect 1540 1815 1550 1835
rect 1510 1785 1550 1815
rect 1510 1765 1520 1785
rect 1540 1765 1550 1785
rect 1510 1750 1550 1765
rect 1570 2085 1610 2100
rect 1570 2065 1580 2085
rect 1600 2065 1610 2085
rect 1570 2035 1610 2065
rect 1570 2015 1580 2035
rect 1600 2015 1610 2035
rect 1570 1985 1610 2015
rect 1570 1965 1580 1985
rect 1600 1965 1610 1985
rect 1570 1935 1610 1965
rect 1570 1915 1580 1935
rect 1600 1915 1610 1935
rect 1570 1885 1610 1915
rect 1570 1865 1580 1885
rect 1600 1865 1610 1885
rect 1570 1835 1610 1865
rect 1570 1815 1580 1835
rect 1600 1815 1610 1835
rect 1570 1785 1610 1815
rect 1570 1765 1580 1785
rect 1600 1765 1610 1785
rect 1570 1750 1610 1765
rect 1630 2085 1670 2100
rect 1630 2065 1640 2085
rect 1660 2065 1670 2085
rect 1630 2035 1670 2065
rect 1630 2015 1640 2035
rect 1660 2015 1670 2035
rect 1630 1985 1670 2015
rect 1630 1965 1640 1985
rect 1660 1965 1670 1985
rect 1630 1935 1670 1965
rect 1630 1915 1640 1935
rect 1660 1915 1670 1935
rect 1630 1885 1670 1915
rect 1630 1865 1640 1885
rect 1660 1865 1670 1885
rect 1630 1835 1670 1865
rect 1630 1815 1640 1835
rect 1660 1815 1670 1835
rect 1630 1785 1670 1815
rect 1630 1765 1640 1785
rect 1660 1765 1670 1785
rect 1630 1750 1670 1765
rect 1690 2085 1730 2100
rect 1690 2065 1700 2085
rect 1720 2065 1730 2085
rect 1690 2035 1730 2065
rect 1690 2015 1700 2035
rect 1720 2015 1730 2035
rect 1690 1985 1730 2015
rect 1690 1965 1700 1985
rect 1720 1965 1730 1985
rect 1690 1935 1730 1965
rect 1690 1915 1700 1935
rect 1720 1915 1730 1935
rect 1690 1885 1730 1915
rect 1690 1865 1700 1885
rect 1720 1865 1730 1885
rect 1690 1835 1730 1865
rect 1690 1815 1700 1835
rect 1720 1815 1730 1835
rect 1690 1785 1730 1815
rect 1690 1765 1700 1785
rect 1720 1765 1730 1785
rect 1690 1750 1730 1765
rect 2015 2085 2055 2100
rect 2015 2065 2025 2085
rect 2045 2065 2055 2085
rect 2015 2035 2055 2065
rect 2015 2015 2025 2035
rect 2045 2015 2055 2035
rect 2015 1985 2055 2015
rect 2015 1965 2025 1985
rect 2045 1965 2055 1985
rect 2015 1935 2055 1965
rect 2015 1915 2025 1935
rect 2045 1915 2055 1935
rect 2015 1885 2055 1915
rect 2015 1865 2025 1885
rect 2045 1865 2055 1885
rect 2015 1835 2055 1865
rect 2015 1815 2025 1835
rect 2045 1815 2055 1835
rect 2015 1785 2055 1815
rect 2015 1765 2025 1785
rect 2045 1765 2055 1785
rect 2015 1750 2055 1765
rect 2075 2085 2115 2100
rect 2075 2065 2085 2085
rect 2105 2065 2115 2085
rect 2075 2035 2115 2065
rect 2075 2015 2085 2035
rect 2105 2015 2115 2035
rect 2075 1985 2115 2015
rect 2075 1965 2085 1985
rect 2105 1965 2115 1985
rect 2075 1935 2115 1965
rect 2075 1915 2085 1935
rect 2105 1915 2115 1935
rect 2075 1885 2115 1915
rect 2075 1865 2085 1885
rect 2105 1865 2115 1885
rect 2075 1835 2115 1865
rect 2075 1815 2085 1835
rect 2105 1815 2115 1835
rect 2075 1785 2115 1815
rect 2075 1765 2085 1785
rect 2105 1765 2115 1785
rect 2075 1750 2115 1765
rect 2135 2085 2175 2100
rect 2135 2065 2145 2085
rect 2165 2065 2175 2085
rect 2135 2035 2175 2065
rect 2135 2015 2145 2035
rect 2165 2015 2175 2035
rect 2135 1985 2175 2015
rect 2135 1965 2145 1985
rect 2165 1965 2175 1985
rect 2135 1935 2175 1965
rect 2135 1915 2145 1935
rect 2165 1915 2175 1935
rect 2135 1885 2175 1915
rect 2135 1865 2145 1885
rect 2165 1865 2175 1885
rect 2135 1835 2175 1865
rect 2135 1815 2145 1835
rect 2165 1815 2175 1835
rect 2135 1785 2175 1815
rect 2135 1765 2145 1785
rect 2165 1765 2175 1785
rect 2135 1750 2175 1765
rect 2195 2085 2235 2100
rect 2195 2065 2205 2085
rect 2225 2065 2235 2085
rect 2195 2035 2235 2065
rect 2195 2015 2205 2035
rect 2225 2015 2235 2035
rect 2195 1985 2235 2015
rect 2195 1965 2205 1985
rect 2225 1965 2235 1985
rect 2195 1935 2235 1965
rect 2195 1915 2205 1935
rect 2225 1915 2235 1935
rect 2195 1885 2235 1915
rect 2195 1865 2205 1885
rect 2225 1865 2235 1885
rect 2195 1835 2235 1865
rect 2195 1815 2205 1835
rect 2225 1815 2235 1835
rect 2195 1785 2235 1815
rect 2195 1765 2205 1785
rect 2225 1765 2235 1785
rect 2195 1750 2235 1765
rect 2255 2085 2295 2100
rect 2255 2065 2265 2085
rect 2285 2065 2295 2085
rect 2255 2035 2295 2065
rect 2255 2015 2265 2035
rect 2285 2015 2295 2035
rect 2255 1985 2295 2015
rect 2255 1965 2265 1985
rect 2285 1965 2295 1985
rect 2255 1935 2295 1965
rect 2255 1915 2265 1935
rect 2285 1915 2295 1935
rect 2255 1885 2295 1915
rect 2255 1865 2265 1885
rect 2285 1865 2295 1885
rect 2255 1835 2295 1865
rect 2255 1815 2265 1835
rect 2285 1815 2295 1835
rect 2255 1785 2295 1815
rect 2255 1765 2265 1785
rect 2285 1765 2295 1785
rect 2255 1750 2295 1765
rect 2315 2085 2355 2100
rect 2315 2065 2325 2085
rect 2345 2065 2355 2085
rect 2315 2035 2355 2065
rect 2315 2015 2325 2035
rect 2345 2015 2355 2035
rect 2315 1985 2355 2015
rect 2315 1965 2325 1985
rect 2345 1965 2355 1985
rect 2315 1935 2355 1965
rect 2315 1915 2325 1935
rect 2345 1915 2355 1935
rect 2315 1885 2355 1915
rect 2315 1865 2325 1885
rect 2345 1865 2355 1885
rect 2315 1835 2355 1865
rect 2315 1815 2325 1835
rect 2345 1815 2355 1835
rect 2315 1785 2355 1815
rect 2315 1765 2325 1785
rect 2345 1765 2355 1785
rect 2315 1750 2355 1765
rect 2375 2085 2415 2100
rect 2375 2065 2385 2085
rect 2405 2065 2415 2085
rect 2375 2035 2415 2065
rect 2375 2015 2385 2035
rect 2405 2015 2415 2035
rect 2375 1985 2415 2015
rect 2375 1965 2385 1985
rect 2405 1965 2415 1985
rect 2375 1935 2415 1965
rect 2375 1915 2385 1935
rect 2405 1915 2415 1935
rect 2375 1885 2415 1915
rect 2375 1865 2385 1885
rect 2405 1865 2415 1885
rect 2375 1835 2415 1865
rect 2375 1815 2385 1835
rect 2405 1815 2415 1835
rect 2375 1785 2415 1815
rect 2375 1765 2385 1785
rect 2405 1765 2415 1785
rect 2375 1750 2415 1765
rect 2435 2085 2475 2100
rect 2435 2065 2445 2085
rect 2465 2065 2475 2085
rect 2435 2035 2475 2065
rect 2435 2015 2445 2035
rect 2465 2015 2475 2035
rect 2435 1985 2475 2015
rect 2435 1965 2445 1985
rect 2465 1965 2475 1985
rect 2435 1935 2475 1965
rect 2435 1915 2445 1935
rect 2465 1915 2475 1935
rect 2435 1885 2475 1915
rect 2435 1865 2445 1885
rect 2465 1865 2475 1885
rect 2435 1835 2475 1865
rect 2435 1815 2445 1835
rect 2465 1815 2475 1835
rect 2435 1785 2475 1815
rect 2435 1765 2445 1785
rect 2465 1765 2475 1785
rect 2435 1750 2475 1765
rect 2495 2085 2535 2100
rect 2495 2065 2505 2085
rect 2525 2065 2535 2085
rect 2495 2035 2535 2065
rect 2495 2015 2505 2035
rect 2525 2015 2535 2035
rect 2495 1985 2535 2015
rect 2495 1965 2505 1985
rect 2525 1965 2535 1985
rect 2495 1935 2535 1965
rect 2495 1915 2505 1935
rect 2525 1915 2535 1935
rect 2495 1885 2535 1915
rect 2495 1865 2505 1885
rect 2525 1865 2535 1885
rect 2495 1835 2535 1865
rect 2495 1815 2505 1835
rect 2525 1815 2535 1835
rect 2495 1785 2535 1815
rect 2495 1765 2505 1785
rect 2525 1765 2535 1785
rect 2495 1750 2535 1765
rect 2555 2085 2595 2100
rect 2555 2065 2565 2085
rect 2585 2065 2595 2085
rect 2555 2035 2595 2065
rect 2555 2015 2565 2035
rect 2585 2015 2595 2035
rect 2555 1985 2595 2015
rect 2555 1965 2565 1985
rect 2585 1965 2595 1985
rect 2555 1935 2595 1965
rect 2555 1915 2565 1935
rect 2585 1915 2595 1935
rect 2555 1885 2595 1915
rect 2555 1865 2565 1885
rect 2585 1865 2595 1885
rect 2555 1835 2595 1865
rect 2555 1815 2565 1835
rect 2585 1815 2595 1835
rect 2555 1785 2595 1815
rect 2555 1765 2565 1785
rect 2585 1765 2595 1785
rect 2555 1750 2595 1765
rect 2615 2085 2655 2100
rect 2615 2065 2625 2085
rect 2645 2065 2655 2085
rect 2615 2035 2655 2065
rect 2615 2015 2625 2035
rect 2645 2015 2655 2035
rect 2615 1985 2655 2015
rect 2615 1965 2625 1985
rect 2645 1965 2655 1985
rect 2615 1935 2655 1965
rect 2615 1915 2625 1935
rect 2645 1915 2655 1935
rect 2615 1885 2655 1915
rect 2615 1865 2625 1885
rect 2645 1865 2655 1885
rect 2615 1835 2655 1865
rect 2615 1815 2625 1835
rect 2645 1815 2655 1835
rect 2615 1785 2655 1815
rect 2615 1765 2625 1785
rect 2645 1765 2655 1785
rect 2615 1750 2655 1765
rect 2675 2085 2715 2100
rect 2675 2065 2685 2085
rect 2705 2065 2715 2085
rect 2675 2035 2715 2065
rect 2675 2015 2685 2035
rect 2705 2015 2715 2035
rect 2675 1985 2715 2015
rect 2675 1965 2685 1985
rect 2705 1965 2715 1985
rect 2675 1935 2715 1965
rect 2675 1915 2685 1935
rect 2705 1915 2715 1935
rect 2675 1885 2715 1915
rect 2675 1865 2685 1885
rect 2705 1865 2715 1885
rect 2675 1835 2715 1865
rect 2675 1815 2685 1835
rect 2705 1815 2715 1835
rect 2675 1785 2715 1815
rect 2675 1765 2685 1785
rect 2705 1765 2715 1785
rect 2675 1750 2715 1765
rect 2735 2085 2775 2100
rect 2735 2065 2745 2085
rect 2765 2065 2775 2085
rect 2735 2035 2775 2065
rect 2735 2015 2745 2035
rect 2765 2015 2775 2035
rect 2735 1985 2775 2015
rect 2735 1965 2745 1985
rect 2765 1965 2775 1985
rect 2735 1935 2775 1965
rect 2735 1915 2745 1935
rect 2765 1915 2775 1935
rect 2735 1885 2775 1915
rect 2735 1865 2745 1885
rect 2765 1865 2775 1885
rect 2735 1835 2775 1865
rect 2735 1815 2745 1835
rect 2765 1815 2775 1835
rect 2735 1785 2775 1815
rect 2735 1765 2745 1785
rect 2765 1765 2775 1785
rect 2735 1750 2775 1765
rect 220 1515 260 1530
rect 220 1495 230 1515
rect 250 1495 260 1515
rect 220 1480 260 1495
rect 275 1515 315 1530
rect 275 1495 285 1515
rect 305 1495 315 1515
rect 275 1480 315 1495
rect 330 1515 370 1530
rect 330 1495 340 1515
rect 360 1495 370 1515
rect 330 1480 370 1495
rect 385 1515 425 1530
rect 385 1495 395 1515
rect 415 1495 425 1515
rect 385 1480 425 1495
rect 440 1515 480 1530
rect 440 1495 450 1515
rect 470 1495 480 1515
rect 440 1480 480 1495
rect 495 1515 535 1530
rect 495 1495 505 1515
rect 525 1495 535 1515
rect 495 1480 535 1495
rect 550 1515 590 1530
rect 550 1495 560 1515
rect 580 1495 590 1515
rect 550 1480 590 1495
rect 605 1515 645 1530
rect 605 1495 615 1515
rect 635 1495 645 1515
rect 605 1480 645 1495
rect 660 1515 700 1530
rect 660 1495 670 1515
rect 690 1495 700 1515
rect 660 1480 700 1495
rect 715 1515 755 1530
rect 715 1495 725 1515
rect 745 1495 755 1515
rect 715 1480 755 1495
rect 770 1515 810 1530
rect 770 1495 780 1515
rect 800 1495 810 1515
rect 770 1480 810 1495
rect 825 1515 865 1530
rect 825 1495 835 1515
rect 855 1495 865 1515
rect 825 1480 865 1495
rect 880 1515 920 1530
rect 880 1495 890 1515
rect 910 1495 920 1515
rect 880 1480 920 1495
rect 935 1515 975 1530
rect 935 1495 945 1515
rect 965 1495 975 1515
rect 935 1480 975 1495
rect 990 1515 1030 1530
rect 990 1495 1000 1515
rect 1020 1495 1030 1515
rect 990 1480 1030 1495
rect 1045 1515 1085 1530
rect 1045 1495 1055 1515
rect 1075 1495 1085 1515
rect 1045 1480 1085 1495
rect 1100 1515 1140 1530
rect 1100 1495 1110 1515
rect 1130 1495 1140 1515
rect 1100 1480 1140 1495
rect 1155 1515 1195 1530
rect 1155 1495 1165 1515
rect 1185 1495 1195 1515
rect 1155 1480 1195 1495
rect 1210 1515 1250 1530
rect 1210 1495 1220 1515
rect 1240 1495 1250 1515
rect 1210 1480 1250 1495
rect 1265 1515 1305 1530
rect 1265 1495 1275 1515
rect 1295 1495 1305 1515
rect 1265 1480 1305 1495
rect 1320 1515 1360 1530
rect 1320 1495 1330 1515
rect 1350 1495 1360 1515
rect 1320 1480 1360 1495
rect 1375 1515 1415 1530
rect 1375 1495 1385 1515
rect 1405 1495 1415 1515
rect 1375 1480 1415 1495
rect 1430 1515 1470 1530
rect 1430 1495 1440 1515
rect 1460 1495 1470 1515
rect 1430 1480 1470 1495
rect -1055 1420 -1015 1435
rect -1055 1400 -1045 1420
rect -1025 1400 -1015 1420
rect -1055 1370 -1015 1400
rect -1055 1350 -1045 1370
rect -1025 1350 -1015 1370
rect -1055 1320 -1015 1350
rect -1055 1300 -1045 1320
rect -1025 1300 -1015 1320
rect -1055 1270 -1015 1300
rect -1055 1250 -1045 1270
rect -1025 1250 -1015 1270
rect -1055 1220 -1015 1250
rect -1055 1200 -1045 1220
rect -1025 1200 -1015 1220
rect -1055 1170 -1015 1200
rect -1055 1150 -1045 1170
rect -1025 1150 -1015 1170
rect -1055 1120 -1015 1150
rect -1055 1100 -1045 1120
rect -1025 1100 -1015 1120
rect -1055 1070 -1015 1100
rect -1055 1050 -1045 1070
rect -1025 1050 -1015 1070
rect -1055 1020 -1015 1050
rect -1055 1000 -1045 1020
rect -1025 1000 -1015 1020
rect -1055 970 -1015 1000
rect -1055 950 -1045 970
rect -1025 950 -1015 970
rect -1055 920 -1015 950
rect -1055 900 -1045 920
rect -1025 900 -1015 920
rect -1055 870 -1015 900
rect -1055 850 -1045 870
rect -1025 850 -1015 870
rect -1055 835 -1015 850
rect -1000 1420 -960 1435
rect -1000 1400 -990 1420
rect -970 1400 -960 1420
rect -1000 1370 -960 1400
rect -1000 1350 -990 1370
rect -970 1350 -960 1370
rect -1000 1320 -960 1350
rect -1000 1300 -990 1320
rect -970 1300 -960 1320
rect -1000 1270 -960 1300
rect -1000 1250 -990 1270
rect -970 1250 -960 1270
rect -1000 1220 -960 1250
rect -1000 1200 -990 1220
rect -970 1200 -960 1220
rect -1000 1170 -960 1200
rect -1000 1150 -990 1170
rect -970 1150 -960 1170
rect -1000 1120 -960 1150
rect -1000 1100 -990 1120
rect -970 1100 -960 1120
rect -1000 1070 -960 1100
rect -1000 1050 -990 1070
rect -970 1050 -960 1070
rect -1000 1020 -960 1050
rect -1000 1000 -990 1020
rect -970 1000 -960 1020
rect -1000 970 -960 1000
rect -1000 950 -990 970
rect -970 950 -960 970
rect -1000 920 -960 950
rect -1000 900 -990 920
rect -970 900 -960 920
rect -1000 870 -960 900
rect -1000 850 -990 870
rect -970 850 -960 870
rect -1000 835 -960 850
rect -945 1420 -905 1435
rect -945 1400 -935 1420
rect -915 1400 -905 1420
rect -945 1370 -905 1400
rect -945 1350 -935 1370
rect -915 1350 -905 1370
rect -945 1320 -905 1350
rect -945 1300 -935 1320
rect -915 1300 -905 1320
rect -945 1270 -905 1300
rect -945 1250 -935 1270
rect -915 1250 -905 1270
rect -945 1220 -905 1250
rect -945 1200 -935 1220
rect -915 1200 -905 1220
rect -945 1170 -905 1200
rect -945 1150 -935 1170
rect -915 1150 -905 1170
rect -945 1120 -905 1150
rect -945 1100 -935 1120
rect -915 1100 -905 1120
rect -945 1070 -905 1100
rect -945 1050 -935 1070
rect -915 1050 -905 1070
rect -945 1020 -905 1050
rect -945 1000 -935 1020
rect -915 1000 -905 1020
rect -945 970 -905 1000
rect -945 950 -935 970
rect -915 950 -905 970
rect -945 920 -905 950
rect -945 900 -935 920
rect -915 900 -905 920
rect -945 870 -905 900
rect -945 850 -935 870
rect -915 850 -905 870
rect -945 835 -905 850
rect -890 1420 -850 1435
rect -890 1400 -880 1420
rect -860 1400 -850 1420
rect -890 1370 -850 1400
rect -890 1350 -880 1370
rect -860 1350 -850 1370
rect -890 1320 -850 1350
rect -890 1300 -880 1320
rect -860 1300 -850 1320
rect -890 1270 -850 1300
rect -890 1250 -880 1270
rect -860 1250 -850 1270
rect -890 1220 -850 1250
rect -890 1200 -880 1220
rect -860 1200 -850 1220
rect -890 1170 -850 1200
rect -890 1150 -880 1170
rect -860 1150 -850 1170
rect -890 1120 -850 1150
rect -890 1100 -880 1120
rect -860 1100 -850 1120
rect -890 1070 -850 1100
rect -890 1050 -880 1070
rect -860 1050 -850 1070
rect -890 1020 -850 1050
rect -890 1000 -880 1020
rect -860 1000 -850 1020
rect -890 970 -850 1000
rect -890 950 -880 970
rect -860 950 -850 970
rect -890 920 -850 950
rect -890 900 -880 920
rect -860 900 -850 920
rect -890 870 -850 900
rect -890 850 -880 870
rect -860 850 -850 870
rect -890 835 -850 850
rect -835 1420 -795 1435
rect -835 1400 -825 1420
rect -805 1400 -795 1420
rect -835 1370 -795 1400
rect -835 1350 -825 1370
rect -805 1350 -795 1370
rect -835 1320 -795 1350
rect -835 1300 -825 1320
rect -805 1300 -795 1320
rect -835 1270 -795 1300
rect -835 1250 -825 1270
rect -805 1250 -795 1270
rect -835 1220 -795 1250
rect -835 1200 -825 1220
rect -805 1200 -795 1220
rect -835 1170 -795 1200
rect -835 1150 -825 1170
rect -805 1150 -795 1170
rect -835 1120 -795 1150
rect -835 1100 -825 1120
rect -805 1100 -795 1120
rect -835 1070 -795 1100
rect -835 1050 -825 1070
rect -805 1050 -795 1070
rect -835 1020 -795 1050
rect -835 1000 -825 1020
rect -805 1000 -795 1020
rect -835 970 -795 1000
rect -835 950 -825 970
rect -805 950 -795 970
rect -835 920 -795 950
rect -835 900 -825 920
rect -805 900 -795 920
rect -835 870 -795 900
rect -835 850 -825 870
rect -805 850 -795 870
rect -835 835 -795 850
rect -780 1420 -740 1435
rect -780 1400 -770 1420
rect -750 1400 -740 1420
rect -780 1370 -740 1400
rect -780 1350 -770 1370
rect -750 1350 -740 1370
rect -780 1320 -740 1350
rect -780 1300 -770 1320
rect -750 1300 -740 1320
rect -780 1270 -740 1300
rect -780 1250 -770 1270
rect -750 1250 -740 1270
rect -780 1220 -740 1250
rect -780 1200 -770 1220
rect -750 1200 -740 1220
rect -780 1170 -740 1200
rect -780 1150 -770 1170
rect -750 1150 -740 1170
rect -780 1120 -740 1150
rect -780 1100 -770 1120
rect -750 1100 -740 1120
rect -780 1070 -740 1100
rect -780 1050 -770 1070
rect -750 1050 -740 1070
rect -780 1020 -740 1050
rect -780 1000 -770 1020
rect -750 1000 -740 1020
rect -780 970 -740 1000
rect -780 950 -770 970
rect -750 950 -740 970
rect -780 920 -740 950
rect -780 900 -770 920
rect -750 900 -740 920
rect -780 870 -740 900
rect -780 850 -770 870
rect -750 850 -740 870
rect -780 835 -740 850
rect -725 1420 -685 1435
rect -725 1400 -715 1420
rect -695 1400 -685 1420
rect -725 1370 -685 1400
rect -725 1350 -715 1370
rect -695 1350 -685 1370
rect -725 1320 -685 1350
rect -725 1300 -715 1320
rect -695 1300 -685 1320
rect -725 1270 -685 1300
rect -725 1250 -715 1270
rect -695 1250 -685 1270
rect -725 1220 -685 1250
rect -725 1200 -715 1220
rect -695 1200 -685 1220
rect -725 1170 -685 1200
rect -725 1150 -715 1170
rect -695 1150 -685 1170
rect -725 1120 -685 1150
rect -725 1100 -715 1120
rect -695 1100 -685 1120
rect -725 1070 -685 1100
rect -725 1050 -715 1070
rect -695 1050 -685 1070
rect -725 1020 -685 1050
rect -725 1000 -715 1020
rect -695 1000 -685 1020
rect -725 970 -685 1000
rect -725 950 -715 970
rect -695 950 -685 970
rect -725 920 -685 950
rect -725 900 -715 920
rect -695 900 -685 920
rect -725 870 -685 900
rect -725 850 -715 870
rect -695 850 -685 870
rect -725 835 -685 850
rect -670 1420 -630 1435
rect -670 1400 -660 1420
rect -640 1400 -630 1420
rect -670 1370 -630 1400
rect -670 1350 -660 1370
rect -640 1350 -630 1370
rect -670 1320 -630 1350
rect -670 1300 -660 1320
rect -640 1300 -630 1320
rect -670 1270 -630 1300
rect -670 1250 -660 1270
rect -640 1250 -630 1270
rect -670 1220 -630 1250
rect -670 1200 -660 1220
rect -640 1200 -630 1220
rect -670 1170 -630 1200
rect -670 1150 -660 1170
rect -640 1150 -630 1170
rect -670 1120 -630 1150
rect -670 1100 -660 1120
rect -640 1100 -630 1120
rect -670 1070 -630 1100
rect -670 1050 -660 1070
rect -640 1050 -630 1070
rect -670 1020 -630 1050
rect -670 1000 -660 1020
rect -640 1000 -630 1020
rect -670 970 -630 1000
rect -670 950 -660 970
rect -640 950 -630 970
rect -670 920 -630 950
rect -670 900 -660 920
rect -640 900 -630 920
rect -670 870 -630 900
rect -670 850 -660 870
rect -640 850 -630 870
rect -670 835 -630 850
rect -615 1420 -575 1435
rect -615 1400 -605 1420
rect -585 1400 -575 1420
rect -615 1370 -575 1400
rect -615 1350 -605 1370
rect -585 1350 -575 1370
rect -615 1320 -575 1350
rect -615 1300 -605 1320
rect -585 1300 -575 1320
rect -615 1270 -575 1300
rect -615 1250 -605 1270
rect -585 1250 -575 1270
rect -615 1220 -575 1250
rect -615 1200 -605 1220
rect -585 1200 -575 1220
rect -615 1170 -575 1200
rect -615 1150 -605 1170
rect -585 1150 -575 1170
rect -615 1120 -575 1150
rect -615 1100 -605 1120
rect -585 1100 -575 1120
rect -615 1070 -575 1100
rect -615 1050 -605 1070
rect -585 1050 -575 1070
rect -615 1020 -575 1050
rect -615 1000 -605 1020
rect -585 1000 -575 1020
rect -615 970 -575 1000
rect -615 950 -605 970
rect -585 950 -575 970
rect -615 920 -575 950
rect -615 900 -605 920
rect -585 900 -575 920
rect -615 870 -575 900
rect -615 850 -605 870
rect -585 850 -575 870
rect -615 835 -575 850
rect -560 1420 -520 1435
rect -560 1400 -550 1420
rect -530 1400 -520 1420
rect -560 1370 -520 1400
rect -560 1350 -550 1370
rect -530 1350 -520 1370
rect -560 1320 -520 1350
rect -560 1300 -550 1320
rect -530 1300 -520 1320
rect -560 1270 -520 1300
rect -560 1250 -550 1270
rect -530 1250 -520 1270
rect -560 1220 -520 1250
rect -560 1200 -550 1220
rect -530 1200 -520 1220
rect -560 1170 -520 1200
rect -560 1150 -550 1170
rect -530 1150 -520 1170
rect -560 1120 -520 1150
rect -560 1100 -550 1120
rect -530 1100 -520 1120
rect -560 1070 -520 1100
rect -560 1050 -550 1070
rect -530 1050 -520 1070
rect -560 1020 -520 1050
rect -560 1000 -550 1020
rect -530 1000 -520 1020
rect -560 970 -520 1000
rect -560 950 -550 970
rect -530 950 -520 970
rect -560 920 -520 950
rect -560 900 -550 920
rect -530 900 -520 920
rect -560 870 -520 900
rect -560 850 -550 870
rect -530 850 -520 870
rect -560 835 -520 850
rect -505 1420 -465 1435
rect -505 1400 -495 1420
rect -475 1400 -465 1420
rect -505 1370 -465 1400
rect -505 1350 -495 1370
rect -475 1350 -465 1370
rect -505 1320 -465 1350
rect -505 1300 -495 1320
rect -475 1300 -465 1320
rect -505 1270 -465 1300
rect -505 1250 -495 1270
rect -475 1250 -465 1270
rect -505 1220 -465 1250
rect -505 1200 -495 1220
rect -475 1200 -465 1220
rect -505 1170 -465 1200
rect -505 1150 -495 1170
rect -475 1150 -465 1170
rect -505 1120 -465 1150
rect -505 1100 -495 1120
rect -475 1100 -465 1120
rect -505 1070 -465 1100
rect -505 1050 -495 1070
rect -475 1050 -465 1070
rect -505 1020 -465 1050
rect -505 1000 -495 1020
rect -475 1000 -465 1020
rect -505 970 -465 1000
rect -505 950 -495 970
rect -475 950 -465 970
rect -505 920 -465 950
rect -505 900 -495 920
rect -475 900 -465 920
rect -505 870 -465 900
rect -505 850 -495 870
rect -475 850 -465 870
rect -505 835 -465 850
rect -450 1420 -410 1435
rect -450 1400 -440 1420
rect -420 1400 -410 1420
rect -450 1370 -410 1400
rect -450 1350 -440 1370
rect -420 1350 -410 1370
rect -450 1320 -410 1350
rect -450 1300 -440 1320
rect -420 1300 -410 1320
rect -450 1270 -410 1300
rect -450 1250 -440 1270
rect -420 1250 -410 1270
rect -450 1220 -410 1250
rect -450 1200 -440 1220
rect -420 1200 -410 1220
rect -450 1170 -410 1200
rect -450 1150 -440 1170
rect -420 1150 -410 1170
rect -450 1120 -410 1150
rect -450 1100 -440 1120
rect -420 1100 -410 1120
rect -450 1070 -410 1100
rect -450 1050 -440 1070
rect -420 1050 -410 1070
rect -450 1020 -410 1050
rect -450 1000 -440 1020
rect -420 1000 -410 1020
rect -450 970 -410 1000
rect -450 950 -440 970
rect -420 950 -410 970
rect -450 920 -410 950
rect -450 900 -440 920
rect -420 900 -410 920
rect -450 870 -410 900
rect -450 850 -440 870
rect -420 850 -410 870
rect -450 835 -410 850
rect -395 1420 -355 1435
rect 2045 1420 2085 1435
rect -395 1400 -385 1420
rect -365 1400 -355 1420
rect -395 1370 -355 1400
rect -395 1350 -385 1370
rect -365 1350 -355 1370
rect -395 1320 -355 1350
rect -395 1300 -385 1320
rect -365 1300 -355 1320
rect -395 1270 -355 1300
rect -395 1250 -385 1270
rect -365 1250 -355 1270
rect 2045 1400 2055 1420
rect 2075 1400 2085 1420
rect 2045 1370 2085 1400
rect 2045 1350 2055 1370
rect 2075 1350 2085 1370
rect 2045 1320 2085 1350
rect 2045 1300 2055 1320
rect 2075 1300 2085 1320
rect 2045 1270 2085 1300
rect -395 1220 -355 1250
rect 2045 1250 2055 1270
rect 2075 1250 2085 1270
rect -395 1200 -385 1220
rect -365 1200 -355 1220
rect 2045 1220 2085 1250
rect -395 1170 -355 1200
rect -395 1150 -385 1170
rect -365 1150 -355 1170
rect -5 1190 35 1205
rect -5 1170 5 1190
rect 25 1170 35 1190
rect -5 1155 35 1170
rect 50 1190 90 1205
rect 50 1170 60 1190
rect 80 1170 90 1190
rect 50 1155 90 1170
rect 105 1190 145 1205
rect 105 1170 115 1190
rect 135 1170 145 1190
rect 105 1155 145 1170
rect 160 1190 200 1205
rect 160 1170 170 1190
rect 190 1170 200 1190
rect 160 1155 200 1170
rect 215 1190 255 1205
rect 215 1170 225 1190
rect 245 1170 255 1190
rect 215 1155 255 1170
rect 270 1190 310 1205
rect 270 1170 280 1190
rect 300 1170 310 1190
rect 270 1155 310 1170
rect 325 1190 365 1205
rect 325 1170 335 1190
rect 355 1170 365 1190
rect 325 1155 365 1170
rect 380 1190 420 1205
rect 380 1170 390 1190
rect 410 1170 420 1190
rect 380 1155 420 1170
rect 435 1190 475 1205
rect 435 1170 445 1190
rect 465 1170 475 1190
rect 435 1155 475 1170
rect 490 1190 530 1205
rect 490 1170 500 1190
rect 520 1170 530 1190
rect 490 1155 530 1170
rect 545 1190 585 1205
rect 545 1170 555 1190
rect 575 1170 585 1190
rect 545 1155 585 1170
rect 600 1190 640 1205
rect 600 1170 610 1190
rect 630 1170 640 1190
rect 600 1155 640 1170
rect 655 1190 695 1205
rect 655 1170 665 1190
rect 685 1170 695 1190
rect 655 1155 695 1170
rect 995 1190 1035 1205
rect 995 1170 1005 1190
rect 1025 1170 1035 1190
rect 995 1155 1035 1170
rect 1050 1190 1090 1205
rect 1050 1170 1060 1190
rect 1080 1170 1090 1190
rect 1050 1155 1090 1170
rect 1105 1190 1145 1205
rect 1105 1170 1115 1190
rect 1135 1170 1145 1190
rect 1105 1155 1145 1170
rect 1160 1190 1200 1205
rect 1160 1170 1170 1190
rect 1190 1170 1200 1190
rect 1160 1155 1200 1170
rect 1215 1190 1255 1205
rect 1215 1170 1225 1190
rect 1245 1170 1255 1190
rect 1215 1155 1255 1170
rect 1270 1190 1310 1205
rect 1270 1170 1280 1190
rect 1300 1170 1310 1190
rect 1270 1155 1310 1170
rect 1325 1190 1365 1205
rect 1325 1170 1335 1190
rect 1355 1170 1365 1190
rect 1325 1155 1365 1170
rect 1380 1190 1420 1205
rect 1380 1170 1390 1190
rect 1410 1170 1420 1190
rect 1380 1155 1420 1170
rect 1435 1190 1475 1205
rect 1435 1170 1445 1190
rect 1465 1170 1475 1190
rect 1435 1155 1475 1170
rect 1490 1190 1530 1205
rect 1490 1170 1500 1190
rect 1520 1170 1530 1190
rect 1490 1155 1530 1170
rect 1545 1190 1585 1205
rect 1545 1170 1555 1190
rect 1575 1170 1585 1190
rect 1545 1155 1585 1170
rect 1600 1190 1640 1205
rect 1600 1170 1610 1190
rect 1630 1170 1640 1190
rect 1600 1155 1640 1170
rect 1655 1190 1695 1205
rect 1655 1170 1665 1190
rect 1685 1170 1695 1190
rect 1655 1155 1695 1170
rect 2045 1200 2055 1220
rect 2075 1200 2085 1220
rect 2045 1170 2085 1200
rect -395 1120 -355 1150
rect -395 1100 -385 1120
rect -365 1100 -355 1120
rect 2045 1150 2055 1170
rect 2075 1150 2085 1170
rect 2045 1120 2085 1150
rect 2045 1100 2055 1120
rect 2075 1100 2085 1120
rect -395 1070 -355 1100
rect -395 1050 -385 1070
rect -365 1050 -355 1070
rect -395 1020 -355 1050
rect -395 1000 -385 1020
rect -365 1000 -355 1020
rect -395 970 -355 1000
rect -395 950 -385 970
rect -365 950 -355 970
rect -395 920 -355 950
rect 2045 1070 2085 1100
rect 2045 1050 2055 1070
rect 2075 1050 2085 1070
rect 2045 1020 2085 1050
rect 2045 1000 2055 1020
rect 2075 1000 2085 1020
rect 2045 970 2085 1000
rect 2045 950 2055 970
rect 2075 950 2085 970
rect -395 900 -385 920
rect -365 900 -355 920
rect 2045 920 2085 950
rect -395 870 -355 900
rect 2045 900 2055 920
rect 2075 900 2085 920
rect -395 850 -385 870
rect -365 850 -355 870
rect -395 835 -355 850
rect 2045 870 2085 900
rect 2045 850 2055 870
rect 2075 850 2085 870
rect 2045 835 2085 850
rect 2100 1420 2140 1435
rect 2100 1400 2110 1420
rect 2130 1400 2140 1420
rect 2100 1370 2140 1400
rect 2100 1350 2110 1370
rect 2130 1350 2140 1370
rect 2100 1320 2140 1350
rect 2100 1300 2110 1320
rect 2130 1300 2140 1320
rect 2100 1270 2140 1300
rect 2100 1250 2110 1270
rect 2130 1250 2140 1270
rect 2100 1220 2140 1250
rect 2100 1200 2110 1220
rect 2130 1200 2140 1220
rect 2100 1170 2140 1200
rect 2100 1150 2110 1170
rect 2130 1150 2140 1170
rect 2100 1120 2140 1150
rect 2100 1100 2110 1120
rect 2130 1100 2140 1120
rect 2100 1070 2140 1100
rect 2100 1050 2110 1070
rect 2130 1050 2140 1070
rect 2100 1020 2140 1050
rect 2100 1000 2110 1020
rect 2130 1000 2140 1020
rect 2100 970 2140 1000
rect 2100 950 2110 970
rect 2130 950 2140 970
rect 2100 920 2140 950
rect 2100 900 2110 920
rect 2130 900 2140 920
rect 2100 870 2140 900
rect 2100 850 2110 870
rect 2130 850 2140 870
rect 2100 835 2140 850
rect 2155 1420 2195 1435
rect 2155 1400 2165 1420
rect 2185 1400 2195 1420
rect 2155 1370 2195 1400
rect 2155 1350 2165 1370
rect 2185 1350 2195 1370
rect 2155 1320 2195 1350
rect 2155 1300 2165 1320
rect 2185 1300 2195 1320
rect 2155 1270 2195 1300
rect 2155 1250 2165 1270
rect 2185 1250 2195 1270
rect 2155 1220 2195 1250
rect 2155 1200 2165 1220
rect 2185 1200 2195 1220
rect 2155 1170 2195 1200
rect 2155 1150 2165 1170
rect 2185 1150 2195 1170
rect 2155 1120 2195 1150
rect 2155 1100 2165 1120
rect 2185 1100 2195 1120
rect 2155 1070 2195 1100
rect 2155 1050 2165 1070
rect 2185 1050 2195 1070
rect 2155 1020 2195 1050
rect 2155 1000 2165 1020
rect 2185 1000 2195 1020
rect 2155 970 2195 1000
rect 2155 950 2165 970
rect 2185 950 2195 970
rect 2155 920 2195 950
rect 2155 900 2165 920
rect 2185 900 2195 920
rect 2155 870 2195 900
rect 2155 850 2165 870
rect 2185 850 2195 870
rect 2155 835 2195 850
rect 2210 1420 2250 1435
rect 2210 1400 2220 1420
rect 2240 1400 2250 1420
rect 2210 1370 2250 1400
rect 2210 1350 2220 1370
rect 2240 1350 2250 1370
rect 2210 1320 2250 1350
rect 2210 1300 2220 1320
rect 2240 1300 2250 1320
rect 2210 1270 2250 1300
rect 2210 1250 2220 1270
rect 2240 1250 2250 1270
rect 2210 1220 2250 1250
rect 2210 1200 2220 1220
rect 2240 1200 2250 1220
rect 2210 1170 2250 1200
rect 2210 1150 2220 1170
rect 2240 1150 2250 1170
rect 2210 1120 2250 1150
rect 2210 1100 2220 1120
rect 2240 1100 2250 1120
rect 2210 1070 2250 1100
rect 2210 1050 2220 1070
rect 2240 1050 2250 1070
rect 2210 1020 2250 1050
rect 2210 1000 2220 1020
rect 2240 1000 2250 1020
rect 2210 970 2250 1000
rect 2210 950 2220 970
rect 2240 950 2250 970
rect 2210 920 2250 950
rect 2210 900 2220 920
rect 2240 900 2250 920
rect 2210 870 2250 900
rect 2210 850 2220 870
rect 2240 850 2250 870
rect 2210 835 2250 850
rect 2265 1420 2305 1435
rect 2265 1400 2275 1420
rect 2295 1400 2305 1420
rect 2265 1370 2305 1400
rect 2265 1350 2275 1370
rect 2295 1350 2305 1370
rect 2265 1320 2305 1350
rect 2265 1300 2275 1320
rect 2295 1300 2305 1320
rect 2265 1270 2305 1300
rect 2265 1250 2275 1270
rect 2295 1250 2305 1270
rect 2265 1220 2305 1250
rect 2265 1200 2275 1220
rect 2295 1200 2305 1220
rect 2265 1170 2305 1200
rect 2265 1150 2275 1170
rect 2295 1150 2305 1170
rect 2265 1120 2305 1150
rect 2265 1100 2275 1120
rect 2295 1100 2305 1120
rect 2265 1070 2305 1100
rect 2265 1050 2275 1070
rect 2295 1050 2305 1070
rect 2265 1020 2305 1050
rect 2265 1000 2275 1020
rect 2295 1000 2305 1020
rect 2265 970 2305 1000
rect 2265 950 2275 970
rect 2295 950 2305 970
rect 2265 920 2305 950
rect 2265 900 2275 920
rect 2295 900 2305 920
rect 2265 870 2305 900
rect 2265 850 2275 870
rect 2295 850 2305 870
rect 2265 835 2305 850
rect 2320 1420 2360 1435
rect 2320 1400 2330 1420
rect 2350 1400 2360 1420
rect 2320 1370 2360 1400
rect 2320 1350 2330 1370
rect 2350 1350 2360 1370
rect 2320 1320 2360 1350
rect 2320 1300 2330 1320
rect 2350 1300 2360 1320
rect 2320 1270 2360 1300
rect 2320 1250 2330 1270
rect 2350 1250 2360 1270
rect 2320 1220 2360 1250
rect 2320 1200 2330 1220
rect 2350 1200 2360 1220
rect 2320 1170 2360 1200
rect 2320 1150 2330 1170
rect 2350 1150 2360 1170
rect 2320 1120 2360 1150
rect 2320 1100 2330 1120
rect 2350 1100 2360 1120
rect 2320 1070 2360 1100
rect 2320 1050 2330 1070
rect 2350 1050 2360 1070
rect 2320 1020 2360 1050
rect 2320 1000 2330 1020
rect 2350 1000 2360 1020
rect 2320 970 2360 1000
rect 2320 950 2330 970
rect 2350 950 2360 970
rect 2320 920 2360 950
rect 2320 900 2330 920
rect 2350 900 2360 920
rect 2320 870 2360 900
rect 2320 850 2330 870
rect 2350 850 2360 870
rect 2320 835 2360 850
rect 2375 1420 2415 1435
rect 2375 1400 2385 1420
rect 2405 1400 2415 1420
rect 2375 1370 2415 1400
rect 2375 1350 2385 1370
rect 2405 1350 2415 1370
rect 2375 1320 2415 1350
rect 2375 1300 2385 1320
rect 2405 1300 2415 1320
rect 2375 1270 2415 1300
rect 2375 1250 2385 1270
rect 2405 1250 2415 1270
rect 2375 1220 2415 1250
rect 2375 1200 2385 1220
rect 2405 1200 2415 1220
rect 2375 1170 2415 1200
rect 2375 1150 2385 1170
rect 2405 1150 2415 1170
rect 2375 1120 2415 1150
rect 2375 1100 2385 1120
rect 2405 1100 2415 1120
rect 2375 1070 2415 1100
rect 2375 1050 2385 1070
rect 2405 1050 2415 1070
rect 2375 1020 2415 1050
rect 2375 1000 2385 1020
rect 2405 1000 2415 1020
rect 2375 970 2415 1000
rect 2375 950 2385 970
rect 2405 950 2415 970
rect 2375 920 2415 950
rect 2375 900 2385 920
rect 2405 900 2415 920
rect 2375 870 2415 900
rect 2375 850 2385 870
rect 2405 850 2415 870
rect 2375 835 2415 850
rect 2430 1420 2470 1435
rect 2430 1400 2440 1420
rect 2460 1400 2470 1420
rect 2430 1370 2470 1400
rect 2430 1350 2440 1370
rect 2460 1350 2470 1370
rect 2430 1320 2470 1350
rect 2430 1300 2440 1320
rect 2460 1300 2470 1320
rect 2430 1270 2470 1300
rect 2430 1250 2440 1270
rect 2460 1250 2470 1270
rect 2430 1220 2470 1250
rect 2430 1200 2440 1220
rect 2460 1200 2470 1220
rect 2430 1170 2470 1200
rect 2430 1150 2440 1170
rect 2460 1150 2470 1170
rect 2430 1120 2470 1150
rect 2430 1100 2440 1120
rect 2460 1100 2470 1120
rect 2430 1070 2470 1100
rect 2430 1050 2440 1070
rect 2460 1050 2470 1070
rect 2430 1020 2470 1050
rect 2430 1000 2440 1020
rect 2460 1000 2470 1020
rect 2430 970 2470 1000
rect 2430 950 2440 970
rect 2460 950 2470 970
rect 2430 920 2470 950
rect 2430 900 2440 920
rect 2460 900 2470 920
rect 2430 870 2470 900
rect 2430 850 2440 870
rect 2460 850 2470 870
rect 2430 835 2470 850
rect 2485 1420 2525 1435
rect 2485 1400 2495 1420
rect 2515 1400 2525 1420
rect 2485 1370 2525 1400
rect 2485 1350 2495 1370
rect 2515 1350 2525 1370
rect 2485 1320 2525 1350
rect 2485 1300 2495 1320
rect 2515 1300 2525 1320
rect 2485 1270 2525 1300
rect 2485 1250 2495 1270
rect 2515 1250 2525 1270
rect 2485 1220 2525 1250
rect 2485 1200 2495 1220
rect 2515 1200 2525 1220
rect 2485 1170 2525 1200
rect 2485 1150 2495 1170
rect 2515 1150 2525 1170
rect 2485 1120 2525 1150
rect 2485 1100 2495 1120
rect 2515 1100 2525 1120
rect 2485 1070 2525 1100
rect 2485 1050 2495 1070
rect 2515 1050 2525 1070
rect 2485 1020 2525 1050
rect 2485 1000 2495 1020
rect 2515 1000 2525 1020
rect 2485 970 2525 1000
rect 2485 950 2495 970
rect 2515 950 2525 970
rect 2485 920 2525 950
rect 2485 900 2495 920
rect 2515 900 2525 920
rect 2485 870 2525 900
rect 2485 850 2495 870
rect 2515 850 2525 870
rect 2485 835 2525 850
rect 2540 1420 2580 1435
rect 2540 1400 2550 1420
rect 2570 1400 2580 1420
rect 2540 1370 2580 1400
rect 2540 1350 2550 1370
rect 2570 1350 2580 1370
rect 2540 1320 2580 1350
rect 2540 1300 2550 1320
rect 2570 1300 2580 1320
rect 2540 1270 2580 1300
rect 2540 1250 2550 1270
rect 2570 1250 2580 1270
rect 2540 1220 2580 1250
rect 2540 1200 2550 1220
rect 2570 1200 2580 1220
rect 2540 1170 2580 1200
rect 2540 1150 2550 1170
rect 2570 1150 2580 1170
rect 2540 1120 2580 1150
rect 2540 1100 2550 1120
rect 2570 1100 2580 1120
rect 2540 1070 2580 1100
rect 2540 1050 2550 1070
rect 2570 1050 2580 1070
rect 2540 1020 2580 1050
rect 2540 1000 2550 1020
rect 2570 1000 2580 1020
rect 2540 970 2580 1000
rect 2540 950 2550 970
rect 2570 950 2580 970
rect 2540 920 2580 950
rect 2540 900 2550 920
rect 2570 900 2580 920
rect 2540 870 2580 900
rect 2540 850 2550 870
rect 2570 850 2580 870
rect 2540 835 2580 850
rect 2595 1420 2635 1435
rect 2595 1400 2605 1420
rect 2625 1400 2635 1420
rect 2595 1370 2635 1400
rect 2595 1350 2605 1370
rect 2625 1350 2635 1370
rect 2595 1320 2635 1350
rect 2595 1300 2605 1320
rect 2625 1300 2635 1320
rect 2595 1270 2635 1300
rect 2595 1250 2605 1270
rect 2625 1250 2635 1270
rect 2595 1220 2635 1250
rect 2595 1200 2605 1220
rect 2625 1200 2635 1220
rect 2595 1170 2635 1200
rect 2595 1150 2605 1170
rect 2625 1150 2635 1170
rect 2595 1120 2635 1150
rect 2595 1100 2605 1120
rect 2625 1100 2635 1120
rect 2595 1070 2635 1100
rect 2595 1050 2605 1070
rect 2625 1050 2635 1070
rect 2595 1020 2635 1050
rect 2595 1000 2605 1020
rect 2625 1000 2635 1020
rect 2595 970 2635 1000
rect 2595 950 2605 970
rect 2625 950 2635 970
rect 2595 920 2635 950
rect 2595 900 2605 920
rect 2625 900 2635 920
rect 2595 870 2635 900
rect 2595 850 2605 870
rect 2625 850 2635 870
rect 2595 835 2635 850
rect 2650 1420 2690 1435
rect 2650 1400 2660 1420
rect 2680 1400 2690 1420
rect 2650 1370 2690 1400
rect 2650 1350 2660 1370
rect 2680 1350 2690 1370
rect 2650 1320 2690 1350
rect 2650 1300 2660 1320
rect 2680 1300 2690 1320
rect 2650 1270 2690 1300
rect 2650 1250 2660 1270
rect 2680 1250 2690 1270
rect 2650 1220 2690 1250
rect 2650 1200 2660 1220
rect 2680 1200 2690 1220
rect 2650 1170 2690 1200
rect 2650 1150 2660 1170
rect 2680 1150 2690 1170
rect 2650 1120 2690 1150
rect 2650 1100 2660 1120
rect 2680 1100 2690 1120
rect 2650 1070 2690 1100
rect 2650 1050 2660 1070
rect 2680 1050 2690 1070
rect 2650 1020 2690 1050
rect 2650 1000 2660 1020
rect 2680 1000 2690 1020
rect 2650 970 2690 1000
rect 2650 950 2660 970
rect 2680 950 2690 970
rect 2650 920 2690 950
rect 2650 900 2660 920
rect 2680 900 2690 920
rect 2650 870 2690 900
rect 2650 850 2660 870
rect 2680 850 2690 870
rect 2650 835 2690 850
rect 2705 1420 2745 1435
rect 2705 1400 2715 1420
rect 2735 1400 2745 1420
rect 2705 1370 2745 1400
rect 2705 1350 2715 1370
rect 2735 1350 2745 1370
rect 2705 1320 2745 1350
rect 2705 1300 2715 1320
rect 2735 1300 2745 1320
rect 2705 1270 2745 1300
rect 2705 1250 2715 1270
rect 2735 1250 2745 1270
rect 2705 1220 2745 1250
rect 2705 1200 2715 1220
rect 2735 1200 2745 1220
rect 2705 1170 2745 1200
rect 2705 1150 2715 1170
rect 2735 1150 2745 1170
rect 2705 1120 2745 1150
rect 2705 1100 2715 1120
rect 2735 1100 2745 1120
rect 2705 1070 2745 1100
rect 2705 1050 2715 1070
rect 2735 1050 2745 1070
rect 2705 1020 2745 1050
rect 2705 1000 2715 1020
rect 2735 1000 2745 1020
rect 2705 970 2745 1000
rect 2705 950 2715 970
rect 2735 950 2745 970
rect 2705 920 2745 950
rect 2705 900 2715 920
rect 2735 900 2745 920
rect 2705 870 2745 900
rect 2705 850 2715 870
rect 2735 850 2745 870
rect 2705 835 2745 850
rect -1055 605 -1015 620
rect -1055 585 -1045 605
rect -1025 585 -1015 605
rect -1055 555 -1015 585
rect -1055 535 -1045 555
rect -1025 535 -1015 555
rect -1055 505 -1015 535
rect -1055 485 -1045 505
rect -1025 485 -1015 505
rect -1055 455 -1015 485
rect -1055 435 -1045 455
rect -1025 435 -1015 455
rect -1055 420 -1015 435
rect -1000 605 -960 620
rect -1000 585 -990 605
rect -970 585 -960 605
rect -1000 555 -960 585
rect -1000 535 -990 555
rect -970 535 -960 555
rect -1000 505 -960 535
rect -1000 485 -990 505
rect -970 485 -960 505
rect -1000 455 -960 485
rect -1000 435 -990 455
rect -970 435 -960 455
rect -1000 420 -960 435
rect -945 605 -905 620
rect -945 585 -935 605
rect -915 585 -905 605
rect -945 555 -905 585
rect -945 535 -935 555
rect -915 535 -905 555
rect -945 505 -905 535
rect -945 485 -935 505
rect -915 485 -905 505
rect -945 455 -905 485
rect -945 435 -935 455
rect -915 435 -905 455
rect -945 420 -905 435
rect -890 605 -850 620
rect -890 585 -880 605
rect -860 585 -850 605
rect -890 555 -850 585
rect -890 535 -880 555
rect -860 535 -850 555
rect -890 505 -850 535
rect -890 485 -880 505
rect -860 485 -850 505
rect -890 455 -850 485
rect -890 435 -880 455
rect -860 435 -850 455
rect -890 420 -850 435
rect -835 605 -795 620
rect -835 585 -825 605
rect -805 585 -795 605
rect -835 555 -795 585
rect -835 535 -825 555
rect -805 535 -795 555
rect -835 505 -795 535
rect -835 485 -825 505
rect -805 485 -795 505
rect -835 455 -795 485
rect -835 435 -825 455
rect -805 435 -795 455
rect -835 420 -795 435
rect -780 605 -740 620
rect -780 585 -770 605
rect -750 585 -740 605
rect -780 555 -740 585
rect -780 535 -770 555
rect -750 535 -740 555
rect -780 505 -740 535
rect -780 485 -770 505
rect -750 485 -740 505
rect -780 455 -740 485
rect -780 435 -770 455
rect -750 435 -740 455
rect -780 420 -740 435
rect -725 605 -685 620
rect -725 585 -715 605
rect -695 585 -685 605
rect -725 555 -685 585
rect -725 535 -715 555
rect -695 535 -685 555
rect -725 505 -685 535
rect -725 485 -715 505
rect -695 485 -685 505
rect -725 455 -685 485
rect -725 435 -715 455
rect -695 435 -685 455
rect -725 420 -685 435
rect -670 605 -630 620
rect -670 585 -660 605
rect -640 585 -630 605
rect -670 555 -630 585
rect -670 535 -660 555
rect -640 535 -630 555
rect -670 505 -630 535
rect -670 485 -660 505
rect -640 485 -630 505
rect -670 455 -630 485
rect -670 435 -660 455
rect -640 435 -630 455
rect -670 420 -630 435
rect -615 605 -575 620
rect -615 585 -605 605
rect -585 585 -575 605
rect -615 555 -575 585
rect -615 535 -605 555
rect -585 535 -575 555
rect -615 505 -575 535
rect -615 485 -605 505
rect -585 485 -575 505
rect -615 455 -575 485
rect -615 435 -605 455
rect -585 435 -575 455
rect -615 420 -575 435
rect -560 605 -520 620
rect -560 585 -550 605
rect -530 585 -520 605
rect -560 555 -520 585
rect -560 535 -550 555
rect -530 535 -520 555
rect -560 505 -520 535
rect -560 485 -550 505
rect -530 485 -520 505
rect -560 455 -520 485
rect -560 435 -550 455
rect -530 435 -520 455
rect -560 420 -520 435
rect -505 605 -465 620
rect -505 585 -495 605
rect -475 585 -465 605
rect -505 555 -465 585
rect -505 535 -495 555
rect -475 535 -465 555
rect -505 505 -465 535
rect -505 485 -495 505
rect -475 485 -465 505
rect -505 455 -465 485
rect -505 435 -495 455
rect -475 435 -465 455
rect -505 420 -465 435
rect -450 605 -410 620
rect -450 585 -440 605
rect -420 585 -410 605
rect -450 555 -410 585
rect -450 535 -440 555
rect -420 535 -410 555
rect -450 505 -410 535
rect -450 485 -440 505
rect -420 485 -410 505
rect -450 455 -410 485
rect -450 435 -440 455
rect -420 435 -410 455
rect -450 420 -410 435
rect -395 605 -355 620
rect 2045 605 2085 620
rect -395 585 -385 605
rect -365 585 -355 605
rect -395 555 -355 585
rect -395 535 -385 555
rect -365 535 -355 555
rect -395 505 -355 535
rect -395 485 -385 505
rect -365 485 -355 505
rect -395 455 -355 485
rect 2045 585 2055 605
rect 2075 585 2085 605
rect 2045 555 2085 585
rect 2045 535 2055 555
rect 2075 535 2085 555
rect 2045 505 2085 535
rect 2045 485 2055 505
rect 2075 485 2085 505
rect 2045 455 2085 485
rect -395 435 -385 455
rect -365 435 -355 455
rect -395 420 -355 435
rect 2045 435 2055 455
rect 2075 435 2085 455
rect 2045 420 2085 435
rect 2100 605 2140 620
rect 2100 585 2110 605
rect 2130 585 2140 605
rect 2100 555 2140 585
rect 2100 535 2110 555
rect 2130 535 2140 555
rect 2100 505 2140 535
rect 2100 485 2110 505
rect 2130 485 2140 505
rect 2100 455 2140 485
rect 2100 435 2110 455
rect 2130 435 2140 455
rect 2100 420 2140 435
rect 2155 605 2195 620
rect 2155 585 2165 605
rect 2185 585 2195 605
rect 2155 555 2195 585
rect 2155 535 2165 555
rect 2185 535 2195 555
rect 2155 505 2195 535
rect 2155 485 2165 505
rect 2185 485 2195 505
rect 2155 455 2195 485
rect 2155 435 2165 455
rect 2185 435 2195 455
rect 2155 420 2195 435
rect 2210 605 2250 620
rect 2210 585 2220 605
rect 2240 585 2250 605
rect 2210 555 2250 585
rect 2210 535 2220 555
rect 2240 535 2250 555
rect 2210 505 2250 535
rect 2210 485 2220 505
rect 2240 485 2250 505
rect 2210 455 2250 485
rect 2210 435 2220 455
rect 2240 435 2250 455
rect 2210 420 2250 435
rect 2265 605 2305 620
rect 2265 585 2275 605
rect 2295 585 2305 605
rect 2265 555 2305 585
rect 2265 535 2275 555
rect 2295 535 2305 555
rect 2265 505 2305 535
rect 2265 485 2275 505
rect 2295 485 2305 505
rect 2265 455 2305 485
rect 2265 435 2275 455
rect 2295 435 2305 455
rect 2265 420 2305 435
rect 2320 605 2360 620
rect 2320 585 2330 605
rect 2350 585 2360 605
rect 2320 555 2360 585
rect 2320 535 2330 555
rect 2350 535 2360 555
rect 2320 505 2360 535
rect 2320 485 2330 505
rect 2350 485 2360 505
rect 2320 455 2360 485
rect 2320 435 2330 455
rect 2350 435 2360 455
rect 2320 420 2360 435
rect 2375 605 2415 620
rect 2375 585 2385 605
rect 2405 585 2415 605
rect 2375 555 2415 585
rect 2375 535 2385 555
rect 2405 535 2415 555
rect 2375 505 2415 535
rect 2375 485 2385 505
rect 2405 485 2415 505
rect 2375 455 2415 485
rect 2375 435 2385 455
rect 2405 435 2415 455
rect 2375 420 2415 435
rect 2430 605 2470 620
rect 2430 585 2440 605
rect 2460 585 2470 605
rect 2430 555 2470 585
rect 2430 535 2440 555
rect 2460 535 2470 555
rect 2430 505 2470 535
rect 2430 485 2440 505
rect 2460 485 2470 505
rect 2430 455 2470 485
rect 2430 435 2440 455
rect 2460 435 2470 455
rect 2430 420 2470 435
rect 2485 605 2525 620
rect 2485 585 2495 605
rect 2515 585 2525 605
rect 2485 555 2525 585
rect 2485 535 2495 555
rect 2515 535 2525 555
rect 2485 505 2525 535
rect 2485 485 2495 505
rect 2515 485 2525 505
rect 2485 455 2525 485
rect 2485 435 2495 455
rect 2515 435 2525 455
rect 2485 420 2525 435
rect 2540 605 2580 620
rect 2540 585 2550 605
rect 2570 585 2580 605
rect 2540 555 2580 585
rect 2540 535 2550 555
rect 2570 535 2580 555
rect 2540 505 2580 535
rect 2540 485 2550 505
rect 2570 485 2580 505
rect 2540 455 2580 485
rect 2540 435 2550 455
rect 2570 435 2580 455
rect 2540 420 2580 435
rect 2595 605 2635 620
rect 2595 585 2605 605
rect 2625 585 2635 605
rect 2595 555 2635 585
rect 2595 535 2605 555
rect 2625 535 2635 555
rect 2595 505 2635 535
rect 2595 485 2605 505
rect 2625 485 2635 505
rect 2595 455 2635 485
rect 2595 435 2605 455
rect 2625 435 2635 455
rect 2595 420 2635 435
rect 2650 605 2690 620
rect 2650 585 2660 605
rect 2680 585 2690 605
rect 2650 555 2690 585
rect 2650 535 2660 555
rect 2680 535 2690 555
rect 2650 505 2690 535
rect 2650 485 2660 505
rect 2680 485 2690 505
rect 2650 455 2690 485
rect 2650 435 2660 455
rect 2680 435 2690 455
rect 2650 420 2690 435
rect 2705 605 2745 620
rect 2705 585 2715 605
rect 2735 585 2745 605
rect 2705 555 2745 585
rect 2705 535 2715 555
rect 2735 535 2745 555
rect 2705 505 2745 535
rect 2705 485 2715 505
rect 2735 485 2745 505
rect 2705 455 2745 485
rect 2705 435 2715 455
rect 2735 435 2745 455
rect 2705 420 2745 435
<< ndiffc >>
rect 505 845 525 865
rect 560 845 580 865
rect 615 845 635 865
rect 670 845 690 865
rect 725 845 745 865
rect 780 845 800 865
rect 835 845 855 865
rect 890 845 910 865
rect 945 845 965 865
rect 1000 845 1020 865
rect 1055 845 1075 865
rect 1110 845 1130 865
rect 1165 845 1185 865
rect -15 570 5 590
rect -15 520 5 540
rect -15 470 5 490
rect 40 570 60 590
rect 40 520 60 540
rect 40 470 60 490
rect 95 570 115 590
rect 95 520 115 540
rect 95 470 115 490
rect 150 570 170 590
rect 150 520 170 540
rect 150 470 170 490
rect 205 570 225 590
rect 205 520 225 540
rect 205 470 225 490
rect 260 570 280 590
rect 260 520 280 540
rect 260 470 280 490
rect 315 570 335 590
rect 315 520 335 540
rect 315 470 335 490
rect 370 570 390 590
rect 370 520 390 540
rect 370 470 390 490
rect 425 570 445 590
rect 425 520 445 540
rect 425 470 445 490
rect 480 570 500 590
rect 480 520 500 540
rect 480 470 500 490
rect 535 570 555 590
rect 535 520 555 540
rect 535 470 555 490
rect 590 570 610 590
rect 590 520 610 540
rect 590 470 610 490
rect 645 570 665 590
rect 645 520 665 540
rect 645 470 665 490
rect 1025 570 1045 590
rect 1025 520 1045 540
rect 1025 470 1045 490
rect 1080 570 1100 590
rect 1080 520 1100 540
rect 1080 470 1100 490
rect 1135 570 1155 590
rect 1135 520 1155 540
rect 1135 470 1155 490
rect 1190 570 1210 590
rect 1190 520 1210 540
rect 1190 470 1210 490
rect 1245 570 1265 590
rect 1245 520 1265 540
rect 1245 470 1265 490
rect 1300 570 1320 590
rect 1300 520 1320 540
rect 1300 470 1320 490
rect 1355 570 1375 590
rect 1355 520 1375 540
rect 1355 470 1375 490
rect 1410 570 1430 590
rect 1410 520 1430 540
rect 1410 470 1430 490
rect 1465 570 1485 590
rect 1465 520 1485 540
rect 1465 470 1485 490
rect 1520 570 1540 590
rect 1520 520 1540 540
rect 1520 470 1540 490
rect 1575 570 1595 590
rect 1575 520 1595 540
rect 1575 470 1595 490
rect 1630 570 1650 590
rect 1630 520 1650 540
rect 1630 470 1650 490
rect 1685 570 1705 590
rect 1685 520 1705 540
rect 1685 470 1705 490
rect -1045 195 -1025 215
rect -1045 145 -1025 165
rect -1045 95 -1025 115
rect -1045 45 -1025 65
rect -1045 -5 -1025 15
rect -1045 -55 -1025 -35
rect -990 195 -970 215
rect -990 145 -970 165
rect -990 95 -970 115
rect -990 45 -970 65
rect -990 -5 -970 15
rect -990 -55 -970 -35
rect -935 195 -915 215
rect -935 145 -915 165
rect -935 95 -915 115
rect -935 45 -915 65
rect -935 -5 -915 15
rect -935 -55 -915 -35
rect -880 195 -860 215
rect -880 145 -860 165
rect -880 95 -860 115
rect -880 45 -860 65
rect -880 -5 -860 15
rect -880 -55 -860 -35
rect -825 195 -805 215
rect -825 145 -805 165
rect -825 95 -805 115
rect -825 45 -805 65
rect -825 -5 -805 15
rect -825 -55 -805 -35
rect -770 195 -750 215
rect -770 145 -750 165
rect -770 95 -750 115
rect -770 45 -750 65
rect -770 -5 -750 15
rect -770 -55 -750 -35
rect -715 195 -695 215
rect -715 145 -695 165
rect -715 95 -695 115
rect -715 45 -695 65
rect -715 -5 -695 15
rect -715 -55 -695 -35
rect -660 195 -640 215
rect -660 145 -640 165
rect -660 95 -640 115
rect -660 45 -640 65
rect -660 -5 -640 15
rect -660 -55 -640 -35
rect -605 195 -585 215
rect -605 145 -585 165
rect -605 95 -585 115
rect -605 45 -585 65
rect -605 -5 -585 15
rect -605 -55 -585 -35
rect -550 195 -530 215
rect -550 145 -530 165
rect -550 95 -530 115
rect -550 45 -530 65
rect -550 -5 -530 15
rect -550 -55 -530 -35
rect -495 195 -475 215
rect -495 145 -475 165
rect -495 95 -475 115
rect -495 45 -475 65
rect -495 -5 -475 15
rect -495 -55 -475 -35
rect -440 195 -420 215
rect -440 145 -420 165
rect -440 95 -420 115
rect -440 45 -420 65
rect -440 -5 -420 15
rect -440 -55 -420 -35
rect -385 195 -365 215
rect 2055 195 2075 215
rect -385 145 -365 165
rect 2055 145 2075 165
rect -385 95 -365 115
rect -385 45 -365 65
rect -385 -5 -365 15
rect -15 95 5 115
rect -15 45 5 65
rect -15 -5 5 15
rect 40 95 60 115
rect 40 45 60 65
rect 40 -5 60 15
rect 95 95 115 115
rect 95 45 115 65
rect 95 -5 115 15
rect 150 95 170 115
rect 150 45 170 65
rect 150 -5 170 15
rect 205 95 225 115
rect 205 45 225 65
rect 205 -5 225 15
rect 260 95 280 115
rect 260 45 280 65
rect 260 -5 280 15
rect 315 95 335 115
rect 315 45 335 65
rect 315 -5 335 15
rect 370 95 390 115
rect 370 45 390 65
rect 370 -5 390 15
rect 425 95 445 115
rect 425 45 445 65
rect 425 -5 445 15
rect 480 95 500 115
rect 480 45 500 65
rect 480 -5 500 15
rect 535 95 555 115
rect 535 45 555 65
rect 535 -5 555 15
rect 590 95 610 115
rect 590 45 610 65
rect 590 -5 610 15
rect 645 95 665 115
rect 725 95 745 115
rect 645 45 665 65
rect 725 45 745 65
rect 645 -5 665 15
rect 725 -5 745 15
rect 780 95 800 115
rect 780 45 800 65
rect 780 -5 800 15
rect 835 95 855 115
rect 835 45 855 65
rect 835 -5 855 15
rect 890 95 910 115
rect 890 45 910 65
rect 890 -5 910 15
rect 945 95 965 115
rect 1025 95 1045 115
rect 945 45 965 65
rect 1025 45 1045 65
rect 945 -5 965 15
rect 1025 -5 1045 15
rect 1080 95 1100 115
rect 1080 45 1100 65
rect 1080 -5 1100 15
rect 1135 95 1155 115
rect 1135 45 1155 65
rect 1135 -5 1155 15
rect 1190 95 1210 115
rect 1190 45 1210 65
rect 1190 -5 1210 15
rect 1245 95 1265 115
rect 1245 45 1265 65
rect 1245 -5 1265 15
rect 1300 95 1320 115
rect 1300 45 1320 65
rect 1300 -5 1320 15
rect 1355 95 1375 115
rect 1355 45 1375 65
rect 1355 -5 1375 15
rect 1410 95 1430 115
rect 1410 45 1430 65
rect 1410 -5 1430 15
rect 1465 95 1485 115
rect 1465 45 1485 65
rect 1465 -5 1485 15
rect 1520 95 1540 115
rect 1520 45 1540 65
rect 1520 -5 1540 15
rect 1575 95 1595 115
rect 1575 45 1595 65
rect 1575 -5 1595 15
rect 1630 95 1650 115
rect 1630 45 1650 65
rect 1630 -5 1650 15
rect 1685 95 1705 115
rect 1685 45 1705 65
rect 1685 -5 1705 15
rect 2055 95 2075 115
rect 2055 45 2075 65
rect 2055 -5 2075 15
rect -385 -55 -365 -35
rect 2055 -55 2075 -35
rect 2110 195 2130 215
rect 2110 145 2130 165
rect 2110 95 2130 115
rect 2110 45 2130 65
rect 2110 -5 2130 15
rect 2110 -55 2130 -35
rect 2165 195 2185 215
rect 2165 145 2185 165
rect 2165 95 2185 115
rect 2165 45 2185 65
rect 2165 -5 2185 15
rect 2165 -55 2185 -35
rect 2220 195 2240 215
rect 2220 145 2240 165
rect 2220 95 2240 115
rect 2220 45 2240 65
rect 2220 -5 2240 15
rect 2220 -55 2240 -35
rect 2275 195 2295 215
rect 2275 145 2295 165
rect 2275 95 2295 115
rect 2275 45 2295 65
rect 2275 -5 2295 15
rect 2275 -55 2295 -35
rect 2330 195 2350 215
rect 2330 145 2350 165
rect 2330 95 2350 115
rect 2330 45 2350 65
rect 2330 -5 2350 15
rect 2330 -55 2350 -35
rect 2385 195 2405 215
rect 2385 145 2405 165
rect 2385 95 2405 115
rect 2385 45 2405 65
rect 2385 -5 2405 15
rect 2385 -55 2405 -35
rect 2440 195 2460 215
rect 2440 145 2460 165
rect 2440 95 2460 115
rect 2440 45 2460 65
rect 2440 -5 2460 15
rect 2440 -55 2460 -35
rect 2495 195 2515 215
rect 2495 145 2515 165
rect 2495 95 2515 115
rect 2495 45 2515 65
rect 2495 -5 2515 15
rect 2495 -55 2515 -35
rect 2550 195 2570 215
rect 2550 145 2570 165
rect 2550 95 2570 115
rect 2550 45 2570 65
rect 2550 -5 2570 15
rect 2550 -55 2570 -35
rect 2605 195 2625 215
rect 2605 145 2625 165
rect 2605 95 2625 115
rect 2605 45 2625 65
rect 2605 -5 2625 15
rect 2605 -55 2625 -35
rect 2660 195 2680 215
rect 2660 145 2680 165
rect 2660 95 2680 115
rect 2660 45 2680 65
rect 2660 -5 2680 15
rect 2660 -55 2680 -35
rect 2715 195 2735 215
rect 2715 145 2735 165
rect 2715 95 2735 115
rect 2715 45 2735 65
rect 2715 -5 2735 15
rect 2715 -55 2735 -35
rect -1015 -390 -995 -370
rect -1015 -440 -995 -420
rect -1015 -490 -995 -470
rect -1015 -540 -995 -520
rect -1015 -590 -995 -570
rect -1015 -640 -995 -620
rect -1015 -690 -995 -670
rect -1015 -740 -995 -720
rect -1015 -790 -995 -770
rect -1015 -840 -995 -820
rect -1015 -890 -995 -870
rect -1015 -940 -995 -920
rect -1015 -990 -995 -970
rect -1015 -1040 -995 -1020
rect -915 -390 -895 -370
rect -915 -440 -895 -420
rect -915 -490 -895 -470
rect -915 -540 -895 -520
rect -915 -590 -895 -570
rect -915 -640 -895 -620
rect -915 -690 -895 -670
rect -915 -740 -895 -720
rect -915 -790 -895 -770
rect -915 -840 -895 -820
rect -915 -890 -895 -870
rect -915 -940 -895 -920
rect -915 -990 -895 -970
rect -915 -1040 -895 -1020
rect -815 -390 -795 -370
rect -815 -440 -795 -420
rect -815 -490 -795 -470
rect -815 -540 -795 -520
rect -815 -590 -795 -570
rect -815 -640 -795 -620
rect -815 -690 -795 -670
rect -815 -740 -795 -720
rect -815 -790 -795 -770
rect -815 -840 -795 -820
rect -815 -890 -795 -870
rect -815 -940 -795 -920
rect -815 -990 -795 -970
rect -815 -1040 -795 -1020
rect -715 -390 -695 -370
rect -715 -440 -695 -420
rect -715 -490 -695 -470
rect -715 -540 -695 -520
rect -715 -590 -695 -570
rect -715 -640 -695 -620
rect -715 -690 -695 -670
rect -715 -740 -695 -720
rect -715 -790 -695 -770
rect -715 -840 -695 -820
rect -715 -890 -695 -870
rect -715 -940 -695 -920
rect -715 -990 -695 -970
rect -715 -1040 -695 -1020
rect -615 -390 -595 -370
rect -615 -440 -595 -420
rect -615 -490 -595 -470
rect -615 -540 -595 -520
rect -615 -590 -595 -570
rect -615 -640 -595 -620
rect -615 -690 -595 -670
rect -615 -740 -595 -720
rect -615 -790 -595 -770
rect -615 -840 -595 -820
rect -615 -890 -595 -870
rect -615 -940 -595 -920
rect -615 -990 -595 -970
rect -615 -1040 -595 -1020
rect -515 -390 -495 -370
rect -515 -440 -495 -420
rect -515 -490 -495 -470
rect -515 -540 -495 -520
rect -515 -590 -495 -570
rect -515 -640 -495 -620
rect -515 -690 -495 -670
rect -515 -740 -495 -720
rect -515 -790 -495 -770
rect -515 -840 -495 -820
rect -515 -890 -495 -870
rect -515 -940 -495 -920
rect -515 -990 -495 -970
rect -515 -1040 -495 -1020
rect -415 -390 -395 -370
rect 2085 -390 2105 -370
rect -415 -440 -395 -420
rect -415 -490 -395 -470
rect -415 -540 -395 -520
rect -415 -590 -395 -570
rect -415 -640 -395 -620
rect 170 -440 190 -420
rect 170 -490 190 -470
rect 170 -540 190 -520
rect 170 -590 190 -570
rect 170 -640 190 -620
rect 225 -440 245 -420
rect 225 -490 245 -470
rect 225 -540 245 -520
rect 225 -590 245 -570
rect 225 -640 245 -620
rect 280 -440 300 -420
rect 280 -490 300 -470
rect 280 -540 300 -520
rect 280 -590 300 -570
rect 280 -640 300 -620
rect 335 -440 355 -420
rect 335 -490 355 -470
rect 335 -540 355 -520
rect 335 -590 355 -570
rect 335 -640 355 -620
rect 390 -440 410 -420
rect 390 -490 410 -470
rect 390 -540 410 -520
rect 390 -590 410 -570
rect 390 -640 410 -620
rect 445 -440 465 -420
rect 445 -490 465 -470
rect 445 -540 465 -520
rect 445 -590 465 -570
rect 445 -640 465 -620
rect 500 -440 520 -420
rect 500 -490 520 -470
rect 500 -540 520 -520
rect 500 -590 520 -570
rect 500 -640 520 -620
rect 555 -440 575 -420
rect 555 -490 575 -470
rect 555 -540 575 -520
rect 555 -590 575 -570
rect 555 -640 575 -620
rect 610 -440 630 -420
rect 610 -490 630 -470
rect 610 -540 630 -520
rect 610 -590 630 -570
rect 610 -640 630 -620
rect 665 -440 685 -420
rect 665 -490 685 -470
rect 665 -540 685 -520
rect 665 -590 685 -570
rect 665 -640 685 -620
rect 720 -440 740 -420
rect 720 -490 740 -470
rect 720 -540 740 -520
rect 720 -590 740 -570
rect 720 -640 740 -620
rect 775 -440 795 -420
rect 775 -490 795 -470
rect 775 -540 795 -520
rect 775 -590 795 -570
rect 775 -640 795 -620
rect 830 -440 850 -420
rect 830 -490 850 -470
rect 830 -540 850 -520
rect 830 -590 850 -570
rect 830 -640 850 -620
rect 885 -440 905 -420
rect 885 -490 905 -470
rect 885 -540 905 -520
rect 885 -590 905 -570
rect 885 -640 905 -620
rect 940 -440 960 -420
rect 940 -490 960 -470
rect 940 -540 960 -520
rect 940 -590 960 -570
rect 940 -640 960 -620
rect 995 -440 1015 -420
rect 995 -490 1015 -470
rect 995 -540 1015 -520
rect 995 -590 1015 -570
rect 995 -640 1015 -620
rect 1050 -440 1070 -420
rect 1050 -490 1070 -470
rect 1050 -540 1070 -520
rect 1050 -590 1070 -570
rect 1050 -640 1070 -620
rect 1105 -440 1125 -420
rect 1105 -490 1125 -470
rect 1105 -540 1125 -520
rect 1105 -590 1125 -570
rect 1105 -640 1125 -620
rect 1160 -440 1180 -420
rect 1160 -490 1180 -470
rect 1160 -540 1180 -520
rect 1160 -590 1180 -570
rect 1160 -640 1180 -620
rect 1215 -440 1235 -420
rect 1215 -490 1235 -470
rect 1215 -540 1235 -520
rect 1215 -590 1235 -570
rect 1215 -640 1235 -620
rect 1270 -440 1290 -420
rect 1270 -490 1290 -470
rect 1270 -540 1290 -520
rect 1270 -590 1290 -570
rect 1270 -640 1290 -620
rect 1325 -440 1345 -420
rect 1325 -490 1345 -470
rect 1325 -540 1345 -520
rect 1325 -590 1345 -570
rect 1325 -640 1345 -620
rect 1380 -440 1400 -420
rect 1380 -490 1400 -470
rect 1380 -540 1400 -520
rect 1380 -590 1400 -570
rect 1380 -640 1400 -620
rect 1435 -440 1455 -420
rect 1435 -490 1455 -470
rect 1435 -540 1455 -520
rect 1435 -590 1455 -570
rect 1435 -640 1455 -620
rect 2085 -440 2105 -420
rect 2085 -490 2105 -470
rect 2085 -540 2105 -520
rect 2085 -590 2105 -570
rect 2085 -640 2105 -620
rect -415 -690 -395 -670
rect 2085 -690 2105 -670
rect -415 -740 -395 -720
rect 2085 -740 2105 -720
rect -415 -790 -395 -770
rect 2085 -790 2105 -770
rect -415 -840 -395 -820
rect -415 -890 -395 -870
rect 675 -855 695 -835
rect 675 -905 695 -885
rect 1005 -855 1025 -835
rect 1005 -905 1025 -885
rect 2085 -840 2105 -820
rect 2085 -890 2105 -870
rect -415 -940 -395 -920
rect -415 -990 -395 -970
rect -415 -1040 -395 -1020
rect 2085 -940 2105 -920
rect 2085 -990 2105 -970
rect 2085 -1040 2105 -1020
rect 2185 -390 2205 -370
rect 2185 -440 2205 -420
rect 2185 -490 2205 -470
rect 2185 -540 2205 -520
rect 2185 -590 2205 -570
rect 2185 -640 2205 -620
rect 2185 -690 2205 -670
rect 2185 -740 2205 -720
rect 2185 -790 2205 -770
rect 2185 -840 2205 -820
rect 2185 -890 2205 -870
rect 2185 -940 2205 -920
rect 2185 -990 2205 -970
rect 2185 -1040 2205 -1020
rect 2285 -390 2305 -370
rect 2285 -440 2305 -420
rect 2285 -490 2305 -470
rect 2285 -540 2305 -520
rect 2285 -590 2305 -570
rect 2285 -640 2305 -620
rect 2285 -690 2305 -670
rect 2285 -740 2305 -720
rect 2285 -790 2305 -770
rect 2285 -840 2305 -820
rect 2285 -890 2305 -870
rect 2285 -940 2305 -920
rect 2285 -990 2305 -970
rect 2285 -1040 2305 -1020
rect 2385 -390 2405 -370
rect 2385 -440 2405 -420
rect 2385 -490 2405 -470
rect 2385 -540 2405 -520
rect 2385 -590 2405 -570
rect 2385 -640 2405 -620
rect 2385 -690 2405 -670
rect 2385 -740 2405 -720
rect 2385 -790 2405 -770
rect 2385 -840 2405 -820
rect 2385 -890 2405 -870
rect 2385 -940 2405 -920
rect 2385 -990 2405 -970
rect 2385 -1040 2405 -1020
rect 2485 -390 2505 -370
rect 2485 -440 2505 -420
rect 2485 -490 2505 -470
rect 2485 -540 2505 -520
rect 2485 -590 2505 -570
rect 2485 -640 2505 -620
rect 2485 -690 2505 -670
rect 2485 -740 2505 -720
rect 2485 -790 2505 -770
rect 2485 -840 2505 -820
rect 2485 -890 2505 -870
rect 2485 -940 2505 -920
rect 2485 -990 2505 -970
rect 2485 -1040 2505 -1020
rect 2585 -390 2605 -370
rect 2585 -440 2605 -420
rect 2585 -490 2605 -470
rect 2585 -540 2605 -520
rect 2585 -590 2605 -570
rect 2585 -640 2605 -620
rect 2585 -690 2605 -670
rect 2585 -740 2605 -720
rect 2585 -790 2605 -770
rect 2585 -840 2605 -820
rect 2585 -890 2605 -870
rect 2585 -940 2605 -920
rect 2585 -990 2605 -970
rect 2585 -1040 2605 -1020
rect 2685 -390 2705 -370
rect 2685 -440 2705 -420
rect 2685 -490 2705 -470
rect 2685 -540 2705 -520
rect 2685 -590 2705 -570
rect 2685 -640 2705 -620
rect 2685 -690 2705 -670
rect 2685 -740 2705 -720
rect 2685 -790 2705 -770
rect 2685 -840 2705 -820
rect 2685 -890 2705 -870
rect 2685 -940 2705 -920
rect 2685 -990 2705 -970
rect 2685 -1040 2705 -1020
<< pdiffc >>
rect 40 2640 60 2660
rect 40 2590 60 2610
rect 40 2540 60 2560
rect 40 2490 60 2510
rect 40 2440 60 2460
rect 40 2390 60 2410
rect 40 2340 60 2360
rect 100 2640 120 2660
rect 100 2590 120 2610
rect 100 2540 120 2560
rect 100 2490 120 2510
rect 100 2440 120 2460
rect 100 2390 120 2410
rect 100 2340 120 2360
rect 160 2640 180 2660
rect 160 2590 180 2610
rect 160 2540 180 2560
rect 160 2490 180 2510
rect 160 2440 180 2460
rect 160 2390 180 2410
rect 160 2340 180 2360
rect 220 2640 240 2660
rect 220 2590 240 2610
rect 980 2640 1000 2660
rect 980 2590 1000 2610
rect 220 2540 240 2560
rect 980 2540 1000 2560
rect 220 2490 240 2510
rect 220 2440 240 2460
rect 220 2390 240 2410
rect 220 2340 240 2360
rect 510 2340 530 2360
rect 570 2340 590 2360
rect 630 2340 650 2360
rect 690 2340 710 2360
rect 980 2490 1000 2510
rect 980 2440 1000 2460
rect 980 2390 1000 2410
rect 980 2340 1000 2360
rect 1040 2640 1060 2660
rect 1040 2590 1060 2610
rect 1040 2540 1060 2560
rect 1040 2490 1060 2510
rect 1040 2440 1060 2460
rect 1040 2390 1060 2410
rect 1040 2340 1060 2360
rect 1100 2640 1120 2660
rect 1100 2590 1120 2610
rect 1100 2540 1120 2560
rect 1100 2490 1120 2510
rect 1100 2440 1120 2460
rect 1100 2390 1120 2410
rect 1100 2340 1120 2360
rect 1160 2640 1180 2660
rect 1160 2590 1180 2610
rect 1160 2540 1180 2560
rect 1160 2490 1180 2510
rect 1160 2440 1180 2460
rect 1160 2390 1180 2410
rect 1160 2340 1180 2360
rect 1448 2640 1468 2660
rect 1448 2590 1468 2610
rect 1448 2540 1468 2560
rect 1448 2490 1468 2510
rect 1448 2440 1468 2460
rect 1448 2390 1468 2410
rect 1448 2340 1468 2360
rect 1508 2640 1528 2660
rect 1508 2590 1528 2610
rect 1508 2540 1528 2560
rect 1508 2490 1528 2510
rect 1508 2440 1528 2460
rect 1508 2390 1528 2410
rect 1508 2340 1528 2360
rect 1568 2640 1588 2660
rect 1568 2590 1588 2610
rect 1568 2540 1588 2560
rect 1568 2490 1588 2510
rect 1568 2440 1588 2460
rect 1568 2390 1588 2410
rect 1568 2340 1588 2360
rect 1628 2640 1648 2660
rect 1628 2590 1648 2610
rect 1628 2540 1648 2560
rect 1628 2490 1648 2510
rect 1628 2440 1648 2460
rect 1628 2390 1648 2410
rect 1628 2340 1648 2360
rect -1075 2065 -1055 2085
rect -1075 2015 -1055 2035
rect -1075 1965 -1055 1985
rect -1075 1915 -1055 1935
rect -1075 1865 -1055 1885
rect -1075 1815 -1055 1835
rect -1075 1765 -1055 1785
rect -1015 2065 -995 2085
rect -1015 2015 -995 2035
rect -1015 1965 -995 1985
rect -1015 1915 -995 1935
rect -1015 1865 -995 1885
rect -1015 1815 -995 1835
rect -1015 1765 -995 1785
rect -955 2065 -935 2085
rect -955 2015 -935 2035
rect -955 1965 -935 1985
rect -955 1915 -935 1935
rect -955 1865 -935 1885
rect -955 1815 -935 1835
rect -955 1765 -935 1785
rect -895 2065 -875 2085
rect -895 2015 -875 2035
rect -895 1965 -875 1985
rect -895 1915 -875 1935
rect -895 1865 -875 1885
rect -895 1815 -875 1835
rect -895 1765 -875 1785
rect -835 2065 -815 2085
rect -835 2015 -815 2035
rect -835 1965 -815 1985
rect -835 1915 -815 1935
rect -835 1865 -815 1885
rect -835 1815 -815 1835
rect -835 1765 -815 1785
rect -775 2065 -755 2085
rect -775 2015 -755 2035
rect -775 1965 -755 1985
rect -775 1915 -755 1935
rect -775 1865 -755 1885
rect -775 1815 -755 1835
rect -775 1765 -755 1785
rect -715 2065 -695 2085
rect -715 2015 -695 2035
rect -715 1965 -695 1985
rect -715 1915 -695 1935
rect -715 1865 -695 1885
rect -715 1815 -695 1835
rect -715 1765 -695 1785
rect -655 2065 -635 2085
rect -655 2015 -635 2035
rect -655 1965 -635 1985
rect -655 1915 -635 1935
rect -655 1865 -635 1885
rect -655 1815 -635 1835
rect -655 1765 -635 1785
rect -595 2065 -575 2085
rect -595 2015 -575 2035
rect -595 1965 -575 1985
rect -595 1915 -575 1935
rect -595 1865 -575 1885
rect -595 1815 -575 1835
rect -595 1765 -575 1785
rect -535 2065 -515 2085
rect -535 2015 -515 2035
rect -535 1965 -515 1985
rect -535 1915 -515 1935
rect -535 1865 -515 1885
rect -535 1815 -515 1835
rect -535 1765 -515 1785
rect -475 2065 -455 2085
rect -475 2015 -455 2035
rect -475 1965 -455 1985
rect -475 1915 -455 1935
rect -475 1865 -455 1885
rect -475 1815 -455 1835
rect -475 1765 -455 1785
rect -415 2065 -395 2085
rect -415 2015 -395 2035
rect -415 1965 -395 1985
rect -415 1915 -395 1935
rect -415 1865 -395 1885
rect -415 1815 -395 1835
rect -415 1765 -395 1785
rect -355 2065 -335 2085
rect -355 2015 -335 2035
rect -355 1965 -335 1985
rect -355 1915 -335 1935
rect -355 1865 -335 1885
rect -355 1815 -335 1835
rect -355 1765 -335 1785
rect -30 2065 -10 2085
rect -30 2015 -10 2035
rect -30 1965 -10 1985
rect -30 1915 -10 1935
rect -30 1865 -10 1885
rect -30 1815 -10 1835
rect -30 1765 -10 1785
rect 30 2065 50 2085
rect 30 2015 50 2035
rect 30 1965 50 1985
rect 30 1915 50 1935
rect 30 1865 50 1885
rect 30 1815 50 1835
rect 30 1765 50 1785
rect 90 2065 110 2085
rect 90 2015 110 2035
rect 90 1965 110 1985
rect 90 1915 110 1935
rect 90 1865 110 1885
rect 90 1815 110 1835
rect 90 1765 110 1785
rect 150 2065 170 2085
rect 150 2015 170 2035
rect 150 1965 170 1985
rect 150 1915 170 1935
rect 150 1865 170 1885
rect 150 1815 170 1835
rect 150 1765 170 1785
rect 210 2065 230 2085
rect 210 2015 230 2035
rect 210 1965 230 1985
rect 210 1915 230 1935
rect 210 1865 230 1885
rect 210 1815 230 1835
rect 210 1765 230 1785
rect 270 2065 290 2085
rect 270 2015 290 2035
rect 270 1965 290 1985
rect 270 1915 290 1935
rect 270 1865 290 1885
rect 270 1815 290 1835
rect 270 1765 290 1785
rect 330 2065 350 2085
rect 330 2015 350 2035
rect 330 1965 350 1985
rect 330 1915 350 1935
rect 330 1865 350 1885
rect 330 1815 350 1835
rect 330 1765 350 1785
rect 390 2065 410 2085
rect 390 2015 410 2035
rect 390 1965 410 1985
rect 390 1915 410 1935
rect 390 1865 410 1885
rect 390 1815 410 1835
rect 390 1765 410 1785
rect 450 2065 470 2085
rect 450 2015 470 2035
rect 450 1965 470 1985
rect 450 1915 470 1935
rect 450 1865 470 1885
rect 450 1815 470 1835
rect 450 1765 470 1785
rect 510 2065 530 2085
rect 510 2015 530 2035
rect 510 1965 530 1985
rect 510 1915 530 1935
rect 510 1865 530 1885
rect 510 1815 530 1835
rect 510 1765 530 1785
rect 570 2065 590 2085
rect 570 2015 590 2035
rect 570 1965 590 1985
rect 570 1915 590 1935
rect 570 1865 590 1885
rect 570 1815 590 1835
rect 570 1765 590 1785
rect 630 2065 650 2085
rect 630 2015 650 2035
rect 630 1965 650 1985
rect 630 1915 650 1935
rect 630 1865 650 1885
rect 630 1815 650 1835
rect 630 1765 650 1785
rect 690 2065 710 2085
rect 690 2015 710 2035
rect 690 1965 710 1985
rect 690 1915 710 1935
rect 690 1865 710 1885
rect 690 1815 710 1835
rect 690 1765 710 1785
rect 980 2065 1000 2085
rect 980 2015 1000 2035
rect 980 1965 1000 1985
rect 980 1915 1000 1935
rect 980 1865 1000 1885
rect 980 1815 1000 1835
rect 980 1765 1000 1785
rect 1040 2065 1060 2085
rect 1040 2015 1060 2035
rect 1040 1965 1060 1985
rect 1040 1915 1060 1935
rect 1040 1865 1060 1885
rect 1040 1815 1060 1835
rect 1040 1765 1060 1785
rect 1100 2065 1120 2085
rect 1100 2015 1120 2035
rect 1100 1965 1120 1985
rect 1100 1915 1120 1935
rect 1100 1865 1120 1885
rect 1100 1815 1120 1835
rect 1100 1765 1120 1785
rect 1160 2065 1180 2085
rect 1160 2015 1180 2035
rect 1160 1965 1180 1985
rect 1160 1915 1180 1935
rect 1160 1865 1180 1885
rect 1160 1815 1180 1835
rect 1160 1765 1180 1785
rect 1220 2065 1240 2085
rect 1220 2015 1240 2035
rect 1220 1965 1240 1985
rect 1220 1915 1240 1935
rect 1220 1865 1240 1885
rect 1220 1815 1240 1835
rect 1220 1765 1240 1785
rect 1280 2065 1300 2085
rect 1280 2015 1300 2035
rect 1280 1965 1300 1985
rect 1280 1915 1300 1935
rect 1280 1865 1300 1885
rect 1280 1815 1300 1835
rect 1280 1765 1300 1785
rect 1340 2065 1360 2085
rect 1340 2015 1360 2035
rect 1340 1965 1360 1985
rect 1340 1915 1360 1935
rect 1340 1865 1360 1885
rect 1340 1815 1360 1835
rect 1340 1765 1360 1785
rect 1400 2065 1420 2085
rect 1400 2015 1420 2035
rect 1400 1965 1420 1985
rect 1400 1915 1420 1935
rect 1400 1865 1420 1885
rect 1400 1815 1420 1835
rect 1400 1765 1420 1785
rect 1460 2065 1480 2085
rect 1460 2015 1480 2035
rect 1460 1965 1480 1985
rect 1460 1915 1480 1935
rect 1460 1865 1480 1885
rect 1460 1815 1480 1835
rect 1460 1765 1480 1785
rect 1520 2065 1540 2085
rect 1520 2015 1540 2035
rect 1520 1965 1540 1985
rect 1520 1915 1540 1935
rect 1520 1865 1540 1885
rect 1520 1815 1540 1835
rect 1520 1765 1540 1785
rect 1580 2065 1600 2085
rect 1580 2015 1600 2035
rect 1580 1965 1600 1985
rect 1580 1915 1600 1935
rect 1580 1865 1600 1885
rect 1580 1815 1600 1835
rect 1580 1765 1600 1785
rect 1640 2065 1660 2085
rect 1640 2015 1660 2035
rect 1640 1965 1660 1985
rect 1640 1915 1660 1935
rect 1640 1865 1660 1885
rect 1640 1815 1660 1835
rect 1640 1765 1660 1785
rect 1700 2065 1720 2085
rect 1700 2015 1720 2035
rect 1700 1965 1720 1985
rect 1700 1915 1720 1935
rect 1700 1865 1720 1885
rect 1700 1815 1720 1835
rect 1700 1765 1720 1785
rect 2025 2065 2045 2085
rect 2025 2015 2045 2035
rect 2025 1965 2045 1985
rect 2025 1915 2045 1935
rect 2025 1865 2045 1885
rect 2025 1815 2045 1835
rect 2025 1765 2045 1785
rect 2085 2065 2105 2085
rect 2085 2015 2105 2035
rect 2085 1965 2105 1985
rect 2085 1915 2105 1935
rect 2085 1865 2105 1885
rect 2085 1815 2105 1835
rect 2085 1765 2105 1785
rect 2145 2065 2165 2085
rect 2145 2015 2165 2035
rect 2145 1965 2165 1985
rect 2145 1915 2165 1935
rect 2145 1865 2165 1885
rect 2145 1815 2165 1835
rect 2145 1765 2165 1785
rect 2205 2065 2225 2085
rect 2205 2015 2225 2035
rect 2205 1965 2225 1985
rect 2205 1915 2225 1935
rect 2205 1865 2225 1885
rect 2205 1815 2225 1835
rect 2205 1765 2225 1785
rect 2265 2065 2285 2085
rect 2265 2015 2285 2035
rect 2265 1965 2285 1985
rect 2265 1915 2285 1935
rect 2265 1865 2285 1885
rect 2265 1815 2285 1835
rect 2265 1765 2285 1785
rect 2325 2065 2345 2085
rect 2325 2015 2345 2035
rect 2325 1965 2345 1985
rect 2325 1915 2345 1935
rect 2325 1865 2345 1885
rect 2325 1815 2345 1835
rect 2325 1765 2345 1785
rect 2385 2065 2405 2085
rect 2385 2015 2405 2035
rect 2385 1965 2405 1985
rect 2385 1915 2405 1935
rect 2385 1865 2405 1885
rect 2385 1815 2405 1835
rect 2385 1765 2405 1785
rect 2445 2065 2465 2085
rect 2445 2015 2465 2035
rect 2445 1965 2465 1985
rect 2445 1915 2465 1935
rect 2445 1865 2465 1885
rect 2445 1815 2465 1835
rect 2445 1765 2465 1785
rect 2505 2065 2525 2085
rect 2505 2015 2525 2035
rect 2505 1965 2525 1985
rect 2505 1915 2525 1935
rect 2505 1865 2525 1885
rect 2505 1815 2525 1835
rect 2505 1765 2525 1785
rect 2565 2065 2585 2085
rect 2565 2015 2585 2035
rect 2565 1965 2585 1985
rect 2565 1915 2585 1935
rect 2565 1865 2585 1885
rect 2565 1815 2585 1835
rect 2565 1765 2585 1785
rect 2625 2065 2645 2085
rect 2625 2015 2645 2035
rect 2625 1965 2645 1985
rect 2625 1915 2645 1935
rect 2625 1865 2645 1885
rect 2625 1815 2645 1835
rect 2625 1765 2645 1785
rect 2685 2065 2705 2085
rect 2685 2015 2705 2035
rect 2685 1965 2705 1985
rect 2685 1915 2705 1935
rect 2685 1865 2705 1885
rect 2685 1815 2705 1835
rect 2685 1765 2705 1785
rect 2745 2065 2765 2085
rect 2745 2015 2765 2035
rect 2745 1965 2765 1985
rect 2745 1915 2765 1935
rect 2745 1865 2765 1885
rect 2745 1815 2765 1835
rect 2745 1765 2765 1785
rect 230 1495 250 1515
rect 285 1495 305 1515
rect 340 1495 360 1515
rect 395 1495 415 1515
rect 450 1495 470 1515
rect 505 1495 525 1515
rect 560 1495 580 1515
rect 615 1495 635 1515
rect 670 1495 690 1515
rect 725 1495 745 1515
rect 780 1495 800 1515
rect 835 1495 855 1515
rect 890 1495 910 1515
rect 945 1495 965 1515
rect 1000 1495 1020 1515
rect 1055 1495 1075 1515
rect 1110 1495 1130 1515
rect 1165 1495 1185 1515
rect 1220 1495 1240 1515
rect 1275 1495 1295 1515
rect 1330 1495 1350 1515
rect 1385 1495 1405 1515
rect 1440 1495 1460 1515
rect -1045 1400 -1025 1420
rect -1045 1350 -1025 1370
rect -1045 1300 -1025 1320
rect -1045 1250 -1025 1270
rect -1045 1200 -1025 1220
rect -1045 1150 -1025 1170
rect -1045 1100 -1025 1120
rect -1045 1050 -1025 1070
rect -1045 1000 -1025 1020
rect -1045 950 -1025 970
rect -1045 900 -1025 920
rect -1045 850 -1025 870
rect -990 1400 -970 1420
rect -990 1350 -970 1370
rect -990 1300 -970 1320
rect -990 1250 -970 1270
rect -990 1200 -970 1220
rect -990 1150 -970 1170
rect -990 1100 -970 1120
rect -990 1050 -970 1070
rect -990 1000 -970 1020
rect -990 950 -970 970
rect -990 900 -970 920
rect -990 850 -970 870
rect -935 1400 -915 1420
rect -935 1350 -915 1370
rect -935 1300 -915 1320
rect -935 1250 -915 1270
rect -935 1200 -915 1220
rect -935 1150 -915 1170
rect -935 1100 -915 1120
rect -935 1050 -915 1070
rect -935 1000 -915 1020
rect -935 950 -915 970
rect -935 900 -915 920
rect -935 850 -915 870
rect -880 1400 -860 1420
rect -880 1350 -860 1370
rect -880 1300 -860 1320
rect -880 1250 -860 1270
rect -880 1200 -860 1220
rect -880 1150 -860 1170
rect -880 1100 -860 1120
rect -880 1050 -860 1070
rect -880 1000 -860 1020
rect -880 950 -860 970
rect -880 900 -860 920
rect -880 850 -860 870
rect -825 1400 -805 1420
rect -825 1350 -805 1370
rect -825 1300 -805 1320
rect -825 1250 -805 1270
rect -825 1200 -805 1220
rect -825 1150 -805 1170
rect -825 1100 -805 1120
rect -825 1050 -805 1070
rect -825 1000 -805 1020
rect -825 950 -805 970
rect -825 900 -805 920
rect -825 850 -805 870
rect -770 1400 -750 1420
rect -770 1350 -750 1370
rect -770 1300 -750 1320
rect -770 1250 -750 1270
rect -770 1200 -750 1220
rect -770 1150 -750 1170
rect -770 1100 -750 1120
rect -770 1050 -750 1070
rect -770 1000 -750 1020
rect -770 950 -750 970
rect -770 900 -750 920
rect -770 850 -750 870
rect -715 1400 -695 1420
rect -715 1350 -695 1370
rect -715 1300 -695 1320
rect -715 1250 -695 1270
rect -715 1200 -695 1220
rect -715 1150 -695 1170
rect -715 1100 -695 1120
rect -715 1050 -695 1070
rect -715 1000 -695 1020
rect -715 950 -695 970
rect -715 900 -695 920
rect -715 850 -695 870
rect -660 1400 -640 1420
rect -660 1350 -640 1370
rect -660 1300 -640 1320
rect -660 1250 -640 1270
rect -660 1200 -640 1220
rect -660 1150 -640 1170
rect -660 1100 -640 1120
rect -660 1050 -640 1070
rect -660 1000 -640 1020
rect -660 950 -640 970
rect -660 900 -640 920
rect -660 850 -640 870
rect -605 1400 -585 1420
rect -605 1350 -585 1370
rect -605 1300 -585 1320
rect -605 1250 -585 1270
rect -605 1200 -585 1220
rect -605 1150 -585 1170
rect -605 1100 -585 1120
rect -605 1050 -585 1070
rect -605 1000 -585 1020
rect -605 950 -585 970
rect -605 900 -585 920
rect -605 850 -585 870
rect -550 1400 -530 1420
rect -550 1350 -530 1370
rect -550 1300 -530 1320
rect -550 1250 -530 1270
rect -550 1200 -530 1220
rect -550 1150 -530 1170
rect -550 1100 -530 1120
rect -550 1050 -530 1070
rect -550 1000 -530 1020
rect -550 950 -530 970
rect -550 900 -530 920
rect -550 850 -530 870
rect -495 1400 -475 1420
rect -495 1350 -475 1370
rect -495 1300 -475 1320
rect -495 1250 -475 1270
rect -495 1200 -475 1220
rect -495 1150 -475 1170
rect -495 1100 -475 1120
rect -495 1050 -475 1070
rect -495 1000 -475 1020
rect -495 950 -475 970
rect -495 900 -475 920
rect -495 850 -475 870
rect -440 1400 -420 1420
rect -440 1350 -420 1370
rect -440 1300 -420 1320
rect -440 1250 -420 1270
rect -440 1200 -420 1220
rect -440 1150 -420 1170
rect -440 1100 -420 1120
rect -440 1050 -420 1070
rect -440 1000 -420 1020
rect -440 950 -420 970
rect -440 900 -420 920
rect -440 850 -420 870
rect -385 1400 -365 1420
rect -385 1350 -365 1370
rect -385 1300 -365 1320
rect -385 1250 -365 1270
rect 2055 1400 2075 1420
rect 2055 1350 2075 1370
rect 2055 1300 2075 1320
rect 2055 1250 2075 1270
rect -385 1200 -365 1220
rect -385 1150 -365 1170
rect 5 1170 25 1190
rect 60 1170 80 1190
rect 115 1170 135 1190
rect 170 1170 190 1190
rect 225 1170 245 1190
rect 280 1170 300 1190
rect 335 1170 355 1190
rect 390 1170 410 1190
rect 445 1170 465 1190
rect 500 1170 520 1190
rect 555 1170 575 1190
rect 610 1170 630 1190
rect 665 1170 685 1190
rect 1005 1170 1025 1190
rect 1060 1170 1080 1190
rect 1115 1170 1135 1190
rect 1170 1170 1190 1190
rect 1225 1170 1245 1190
rect 1280 1170 1300 1190
rect 1335 1170 1355 1190
rect 1390 1170 1410 1190
rect 1445 1170 1465 1190
rect 1500 1170 1520 1190
rect 1555 1170 1575 1190
rect 1610 1170 1630 1190
rect 1665 1170 1685 1190
rect 2055 1200 2075 1220
rect -385 1100 -365 1120
rect 2055 1150 2075 1170
rect 2055 1100 2075 1120
rect -385 1050 -365 1070
rect -385 1000 -365 1020
rect -385 950 -365 970
rect 2055 1050 2075 1070
rect 2055 1000 2075 1020
rect 2055 950 2075 970
rect -385 900 -365 920
rect 2055 900 2075 920
rect -385 850 -365 870
rect 2055 850 2075 870
rect 2110 1400 2130 1420
rect 2110 1350 2130 1370
rect 2110 1300 2130 1320
rect 2110 1250 2130 1270
rect 2110 1200 2130 1220
rect 2110 1150 2130 1170
rect 2110 1100 2130 1120
rect 2110 1050 2130 1070
rect 2110 1000 2130 1020
rect 2110 950 2130 970
rect 2110 900 2130 920
rect 2110 850 2130 870
rect 2165 1400 2185 1420
rect 2165 1350 2185 1370
rect 2165 1300 2185 1320
rect 2165 1250 2185 1270
rect 2165 1200 2185 1220
rect 2165 1150 2185 1170
rect 2165 1100 2185 1120
rect 2165 1050 2185 1070
rect 2165 1000 2185 1020
rect 2165 950 2185 970
rect 2165 900 2185 920
rect 2165 850 2185 870
rect 2220 1400 2240 1420
rect 2220 1350 2240 1370
rect 2220 1300 2240 1320
rect 2220 1250 2240 1270
rect 2220 1200 2240 1220
rect 2220 1150 2240 1170
rect 2220 1100 2240 1120
rect 2220 1050 2240 1070
rect 2220 1000 2240 1020
rect 2220 950 2240 970
rect 2220 900 2240 920
rect 2220 850 2240 870
rect 2275 1400 2295 1420
rect 2275 1350 2295 1370
rect 2275 1300 2295 1320
rect 2275 1250 2295 1270
rect 2275 1200 2295 1220
rect 2275 1150 2295 1170
rect 2275 1100 2295 1120
rect 2275 1050 2295 1070
rect 2275 1000 2295 1020
rect 2275 950 2295 970
rect 2275 900 2295 920
rect 2275 850 2295 870
rect 2330 1400 2350 1420
rect 2330 1350 2350 1370
rect 2330 1300 2350 1320
rect 2330 1250 2350 1270
rect 2330 1200 2350 1220
rect 2330 1150 2350 1170
rect 2330 1100 2350 1120
rect 2330 1050 2350 1070
rect 2330 1000 2350 1020
rect 2330 950 2350 970
rect 2330 900 2350 920
rect 2330 850 2350 870
rect 2385 1400 2405 1420
rect 2385 1350 2405 1370
rect 2385 1300 2405 1320
rect 2385 1250 2405 1270
rect 2385 1200 2405 1220
rect 2385 1150 2405 1170
rect 2385 1100 2405 1120
rect 2385 1050 2405 1070
rect 2385 1000 2405 1020
rect 2385 950 2405 970
rect 2385 900 2405 920
rect 2385 850 2405 870
rect 2440 1400 2460 1420
rect 2440 1350 2460 1370
rect 2440 1300 2460 1320
rect 2440 1250 2460 1270
rect 2440 1200 2460 1220
rect 2440 1150 2460 1170
rect 2440 1100 2460 1120
rect 2440 1050 2460 1070
rect 2440 1000 2460 1020
rect 2440 950 2460 970
rect 2440 900 2460 920
rect 2440 850 2460 870
rect 2495 1400 2515 1420
rect 2495 1350 2515 1370
rect 2495 1300 2515 1320
rect 2495 1250 2515 1270
rect 2495 1200 2515 1220
rect 2495 1150 2515 1170
rect 2495 1100 2515 1120
rect 2495 1050 2515 1070
rect 2495 1000 2515 1020
rect 2495 950 2515 970
rect 2495 900 2515 920
rect 2495 850 2515 870
rect 2550 1400 2570 1420
rect 2550 1350 2570 1370
rect 2550 1300 2570 1320
rect 2550 1250 2570 1270
rect 2550 1200 2570 1220
rect 2550 1150 2570 1170
rect 2550 1100 2570 1120
rect 2550 1050 2570 1070
rect 2550 1000 2570 1020
rect 2550 950 2570 970
rect 2550 900 2570 920
rect 2550 850 2570 870
rect 2605 1400 2625 1420
rect 2605 1350 2625 1370
rect 2605 1300 2625 1320
rect 2605 1250 2625 1270
rect 2605 1200 2625 1220
rect 2605 1150 2625 1170
rect 2605 1100 2625 1120
rect 2605 1050 2625 1070
rect 2605 1000 2625 1020
rect 2605 950 2625 970
rect 2605 900 2625 920
rect 2605 850 2625 870
rect 2660 1400 2680 1420
rect 2660 1350 2680 1370
rect 2660 1300 2680 1320
rect 2660 1250 2680 1270
rect 2660 1200 2680 1220
rect 2660 1150 2680 1170
rect 2660 1100 2680 1120
rect 2660 1050 2680 1070
rect 2660 1000 2680 1020
rect 2660 950 2680 970
rect 2660 900 2680 920
rect 2660 850 2680 870
rect 2715 1400 2735 1420
rect 2715 1350 2735 1370
rect 2715 1300 2735 1320
rect 2715 1250 2735 1270
rect 2715 1200 2735 1220
rect 2715 1150 2735 1170
rect 2715 1100 2735 1120
rect 2715 1050 2735 1070
rect 2715 1000 2735 1020
rect 2715 950 2735 970
rect 2715 900 2735 920
rect 2715 850 2735 870
rect -1045 585 -1025 605
rect -1045 535 -1025 555
rect -1045 485 -1025 505
rect -1045 435 -1025 455
rect -990 585 -970 605
rect -990 535 -970 555
rect -990 485 -970 505
rect -990 435 -970 455
rect -935 585 -915 605
rect -935 535 -915 555
rect -935 485 -915 505
rect -935 435 -915 455
rect -880 585 -860 605
rect -880 535 -860 555
rect -880 485 -860 505
rect -880 435 -860 455
rect -825 585 -805 605
rect -825 535 -805 555
rect -825 485 -805 505
rect -825 435 -805 455
rect -770 585 -750 605
rect -770 535 -750 555
rect -770 485 -750 505
rect -770 435 -750 455
rect -715 585 -695 605
rect -715 535 -695 555
rect -715 485 -695 505
rect -715 435 -695 455
rect -660 585 -640 605
rect -660 535 -640 555
rect -660 485 -640 505
rect -660 435 -640 455
rect -605 585 -585 605
rect -605 535 -585 555
rect -605 485 -585 505
rect -605 435 -585 455
rect -550 585 -530 605
rect -550 535 -530 555
rect -550 485 -530 505
rect -550 435 -530 455
rect -495 585 -475 605
rect -495 535 -475 555
rect -495 485 -475 505
rect -495 435 -475 455
rect -440 585 -420 605
rect -440 535 -420 555
rect -440 485 -420 505
rect -440 435 -420 455
rect -385 585 -365 605
rect -385 535 -365 555
rect -385 485 -365 505
rect 2055 585 2075 605
rect 2055 535 2075 555
rect 2055 485 2075 505
rect -385 435 -365 455
rect 2055 435 2075 455
rect 2110 585 2130 605
rect 2110 535 2130 555
rect 2110 485 2130 505
rect 2110 435 2130 455
rect 2165 585 2185 605
rect 2165 535 2185 555
rect 2165 485 2185 505
rect 2165 435 2185 455
rect 2220 585 2240 605
rect 2220 535 2240 555
rect 2220 485 2240 505
rect 2220 435 2240 455
rect 2275 585 2295 605
rect 2275 535 2295 555
rect 2275 485 2295 505
rect 2275 435 2295 455
rect 2330 585 2350 605
rect 2330 535 2350 555
rect 2330 485 2350 505
rect 2330 435 2350 455
rect 2385 585 2405 605
rect 2385 535 2405 555
rect 2385 485 2405 505
rect 2385 435 2405 455
rect 2440 585 2460 605
rect 2440 535 2460 555
rect 2440 485 2460 505
rect 2440 435 2460 455
rect 2495 585 2515 605
rect 2495 535 2515 555
rect 2495 485 2515 505
rect 2495 435 2515 455
rect 2550 585 2570 605
rect 2550 535 2570 555
rect 2550 485 2570 505
rect 2550 435 2570 455
rect 2605 585 2625 605
rect 2605 535 2625 555
rect 2605 485 2625 505
rect 2605 435 2625 455
rect 2660 585 2680 605
rect 2660 535 2680 555
rect 2660 485 2680 505
rect 2660 435 2680 455
rect 2715 585 2735 605
rect 2715 535 2735 555
rect 2715 485 2735 505
rect 2715 435 2735 455
<< psubdiff >>
rect 455 865 495 880
rect 455 845 465 865
rect 485 845 495 865
rect 455 830 495 845
rect 1195 865 1235 880
rect 1195 845 1205 865
rect 1225 845 1235 865
rect 1195 830 1235 845
rect -65 590 -25 605
rect -65 570 -55 590
rect -35 570 -25 590
rect -65 540 -25 570
rect -65 520 -55 540
rect -35 520 -25 540
rect -65 490 -25 520
rect -65 470 -55 490
rect -35 470 -25 490
rect -65 455 -25 470
rect 675 590 715 605
rect 675 570 685 590
rect 705 570 715 590
rect 675 540 715 570
rect 675 520 685 540
rect 705 520 715 540
rect 675 490 715 520
rect 675 470 685 490
rect 705 470 715 490
rect 675 455 715 470
rect 975 590 1015 605
rect 975 570 985 590
rect 1005 570 1015 590
rect 975 540 1015 570
rect 975 520 985 540
rect 1005 520 1015 540
rect 975 490 1015 520
rect 975 470 985 490
rect 1005 470 1015 490
rect 975 455 1015 470
rect 1715 590 1755 605
rect 1715 570 1725 590
rect 1745 570 1755 590
rect 1715 540 1755 570
rect 1715 520 1725 540
rect 1745 520 1755 540
rect 1715 490 1755 520
rect 1715 470 1725 490
rect 1745 470 1755 490
rect 1715 455 1755 470
rect -1095 215 -1055 230
rect -1095 195 -1085 215
rect -1065 195 -1055 215
rect -1095 165 -1055 195
rect -1095 145 -1085 165
rect -1065 145 -1055 165
rect -1095 115 -1055 145
rect -1095 95 -1085 115
rect -1065 95 -1055 115
rect -1095 65 -1055 95
rect -1095 45 -1085 65
rect -1065 45 -1055 65
rect -1095 15 -1055 45
rect -1095 -5 -1085 15
rect -1065 -5 -1055 15
rect -1095 -35 -1055 -5
rect -1095 -55 -1085 -35
rect -1065 -55 -1055 -35
rect -1095 -70 -1055 -55
rect -355 215 -315 230
rect -355 195 -345 215
rect -325 195 -315 215
rect -355 165 -315 195
rect 2005 215 2045 230
rect 2005 195 2015 215
rect 2035 195 2045 215
rect -355 145 -345 165
rect -325 145 -315 165
rect -355 115 -315 145
rect 2005 165 2045 195
rect 2005 145 2015 165
rect 2035 145 2045 165
rect -355 95 -345 115
rect -325 95 -315 115
rect -355 65 -315 95
rect -355 45 -345 65
rect -325 45 -315 65
rect -355 15 -315 45
rect -355 -5 -345 15
rect -325 -5 -315 15
rect -355 -35 -315 -5
rect -65 115 -25 130
rect -65 95 -55 115
rect -35 95 -25 115
rect -65 65 -25 95
rect -65 45 -55 65
rect -35 45 -25 65
rect -65 15 -25 45
rect -65 -5 -55 15
rect -35 -5 -25 15
rect -65 -20 -25 -5
rect 675 115 715 130
rect 675 95 685 115
rect 705 95 715 115
rect 675 65 715 95
rect 675 45 685 65
rect 705 45 715 65
rect 675 15 715 45
rect 675 -5 685 15
rect 705 -5 715 15
rect 675 -20 715 -5
rect 975 115 1015 130
rect 975 95 985 115
rect 1005 95 1015 115
rect 975 65 1015 95
rect 975 45 985 65
rect 1005 45 1015 65
rect 975 15 1015 45
rect 975 -5 985 15
rect 1005 -5 1015 15
rect 975 -20 1015 -5
rect 1715 115 1755 130
rect 1715 95 1725 115
rect 1745 95 1755 115
rect 1715 65 1755 95
rect 1715 45 1725 65
rect 1745 45 1755 65
rect 1715 15 1755 45
rect 1715 -5 1725 15
rect 1745 -5 1755 15
rect 1715 -20 1755 -5
rect 2005 115 2045 145
rect 2005 95 2015 115
rect 2035 95 2045 115
rect 2005 65 2045 95
rect 2005 45 2015 65
rect 2035 45 2045 65
rect 2005 15 2045 45
rect 2005 -5 2015 15
rect 2035 -5 2045 15
rect 2005 -35 2045 -5
rect -355 -55 -345 -35
rect -325 -55 -315 -35
rect -355 -70 -315 -55
rect 2005 -55 2015 -35
rect 2035 -55 2045 -35
rect 2005 -70 2045 -55
rect 2745 215 2785 230
rect 2745 195 2755 215
rect 2775 195 2785 215
rect 2745 165 2785 195
rect 2745 145 2755 165
rect 2775 145 2785 165
rect 2745 115 2785 145
rect 2745 95 2755 115
rect 2775 95 2785 115
rect 2745 65 2785 95
rect 2745 45 2755 65
rect 2775 45 2785 65
rect 2745 15 2785 45
rect 2745 -5 2755 15
rect 2775 -5 2785 15
rect 2745 -35 2785 -5
rect 2745 -55 2755 -35
rect 2775 -55 2785 -35
rect 2745 -70 2785 -55
rect -1065 -370 -1025 -355
rect -1065 -390 -1055 -370
rect -1035 -390 -1025 -370
rect -1065 -420 -1025 -390
rect -1065 -440 -1055 -420
rect -1035 -440 -1025 -420
rect -1065 -470 -1025 -440
rect -1065 -490 -1055 -470
rect -1035 -490 -1025 -470
rect -1065 -520 -1025 -490
rect -1065 -540 -1055 -520
rect -1035 -540 -1025 -520
rect -1065 -570 -1025 -540
rect -1065 -590 -1055 -570
rect -1035 -590 -1025 -570
rect -1065 -620 -1025 -590
rect -1065 -640 -1055 -620
rect -1035 -640 -1025 -620
rect -1065 -670 -1025 -640
rect -1065 -690 -1055 -670
rect -1035 -690 -1025 -670
rect -1065 -720 -1025 -690
rect -1065 -740 -1055 -720
rect -1035 -740 -1025 -720
rect -1065 -770 -1025 -740
rect -1065 -790 -1055 -770
rect -1035 -790 -1025 -770
rect -1065 -820 -1025 -790
rect -1065 -840 -1055 -820
rect -1035 -840 -1025 -820
rect -1065 -870 -1025 -840
rect -1065 -890 -1055 -870
rect -1035 -890 -1025 -870
rect -1065 -920 -1025 -890
rect -1065 -940 -1055 -920
rect -1035 -940 -1025 -920
rect -1065 -970 -1025 -940
rect -1065 -990 -1055 -970
rect -1035 -990 -1025 -970
rect -1065 -1020 -1025 -990
rect -1065 -1040 -1055 -1020
rect -1035 -1040 -1025 -1020
rect -1065 -1055 -1025 -1040
rect -385 -370 -345 -355
rect -385 -390 -375 -370
rect -355 -390 -345 -370
rect 2035 -370 2075 -355
rect -385 -420 -345 -390
rect 2035 -390 2045 -370
rect 2065 -390 2075 -370
rect -385 -440 -375 -420
rect -355 -440 -345 -420
rect -385 -470 -345 -440
rect -385 -490 -375 -470
rect -355 -490 -345 -470
rect -385 -520 -345 -490
rect -385 -540 -375 -520
rect -355 -540 -345 -520
rect -385 -570 -345 -540
rect -385 -590 -375 -570
rect -355 -590 -345 -570
rect -385 -620 -345 -590
rect -385 -640 -375 -620
rect -355 -640 -345 -620
rect -385 -670 -345 -640
rect 120 -420 160 -405
rect 120 -440 130 -420
rect 150 -440 160 -420
rect 120 -470 160 -440
rect 120 -490 130 -470
rect 150 -490 160 -470
rect 120 -520 160 -490
rect 120 -540 130 -520
rect 150 -540 160 -520
rect 120 -570 160 -540
rect 120 -590 130 -570
rect 150 -590 160 -570
rect 120 -620 160 -590
rect 120 -640 130 -620
rect 150 -640 160 -620
rect 120 -655 160 -640
rect 1465 -420 1505 -405
rect 1465 -440 1475 -420
rect 1495 -440 1505 -420
rect 1465 -470 1505 -440
rect 1465 -490 1475 -470
rect 1495 -490 1505 -470
rect 1465 -520 1505 -490
rect 1465 -540 1475 -520
rect 1495 -540 1505 -520
rect 1465 -570 1505 -540
rect 1465 -590 1475 -570
rect 1495 -590 1505 -570
rect 1465 -620 1505 -590
rect 1465 -640 1475 -620
rect 1495 -640 1505 -620
rect 1465 -655 1505 -640
rect 2035 -420 2075 -390
rect 2035 -440 2045 -420
rect 2065 -440 2075 -420
rect 2035 -470 2075 -440
rect 2035 -490 2045 -470
rect 2065 -490 2075 -470
rect 2035 -520 2075 -490
rect 2035 -540 2045 -520
rect 2065 -540 2075 -520
rect 2035 -570 2075 -540
rect 2035 -590 2045 -570
rect 2065 -590 2075 -570
rect 2035 -620 2075 -590
rect 2035 -640 2045 -620
rect 2065 -640 2075 -620
rect 2035 -670 2075 -640
rect -385 -690 -375 -670
rect -355 -690 -345 -670
rect -385 -720 -345 -690
rect 2035 -690 2045 -670
rect 2065 -690 2075 -670
rect -385 -740 -375 -720
rect -355 -740 -345 -720
rect -385 -770 -345 -740
rect 2035 -720 2075 -690
rect 2035 -740 2045 -720
rect 2065 -740 2075 -720
rect -385 -790 -375 -770
rect -355 -790 -345 -770
rect -385 -820 -345 -790
rect 2035 -770 2075 -740
rect 2035 -790 2045 -770
rect 2065 -790 2075 -770
rect 2035 -820 2075 -790
rect -385 -840 -375 -820
rect -355 -840 -345 -820
rect -385 -870 -345 -840
rect -385 -890 -375 -870
rect -355 -890 -345 -870
rect -385 -920 -345 -890
rect 2035 -840 2045 -820
rect 2065 -840 2075 -820
rect 2035 -870 2075 -840
rect 2035 -890 2045 -870
rect 2065 -890 2075 -870
rect 2035 -920 2075 -890
rect -385 -940 -375 -920
rect -355 -940 -345 -920
rect -385 -970 -345 -940
rect -385 -990 -375 -970
rect -355 -990 -345 -970
rect -385 -1020 -345 -990
rect -385 -1040 -375 -1020
rect -355 -1040 -345 -1020
rect -385 -1055 -345 -1040
rect 2035 -940 2045 -920
rect 2065 -940 2075 -920
rect 2035 -970 2075 -940
rect 2035 -990 2045 -970
rect 2065 -990 2075 -970
rect 2035 -1020 2075 -990
rect 2035 -1040 2045 -1020
rect 2065 -1040 2075 -1020
rect 2035 -1055 2075 -1040
rect 2715 -370 2755 -355
rect 2715 -390 2725 -370
rect 2745 -390 2755 -370
rect 2715 -420 2755 -390
rect 2715 -440 2725 -420
rect 2745 -440 2755 -420
rect 2715 -470 2755 -440
rect 2715 -490 2725 -470
rect 2745 -490 2755 -470
rect 2715 -520 2755 -490
rect 2715 -540 2725 -520
rect 2745 -540 2755 -520
rect 2715 -570 2755 -540
rect 2715 -590 2725 -570
rect 2745 -590 2755 -570
rect 2715 -620 2755 -590
rect 2715 -640 2725 -620
rect 2745 -640 2755 -620
rect 2715 -670 2755 -640
rect 2715 -690 2725 -670
rect 2745 -690 2755 -670
rect 2715 -720 2755 -690
rect 2715 -740 2725 -720
rect 2745 -740 2755 -720
rect 2715 -770 2755 -740
rect 2715 -790 2725 -770
rect 2745 -790 2755 -770
rect 2715 -820 2755 -790
rect 2715 -840 2725 -820
rect 2745 -840 2755 -820
rect 2715 -870 2755 -840
rect 2715 -890 2725 -870
rect 2745 -890 2755 -870
rect 2715 -920 2755 -890
rect 2715 -940 2725 -920
rect 2745 -940 2755 -920
rect 2715 -970 2755 -940
rect 2715 -990 2725 -970
rect 2745 -990 2755 -970
rect 2715 -1020 2755 -990
rect 2715 -1040 2725 -1020
rect 2745 -1040 2755 -1020
rect 2715 -1055 2755 -1040
<< nsubdiff >>
rect -10 2660 30 2675
rect -10 2640 0 2660
rect 20 2640 30 2660
rect -10 2610 30 2640
rect -10 2590 0 2610
rect 20 2590 30 2610
rect -10 2560 30 2590
rect -10 2540 0 2560
rect 20 2540 30 2560
rect -10 2510 30 2540
rect -10 2490 0 2510
rect 20 2490 30 2510
rect -10 2460 30 2490
rect -10 2440 0 2460
rect 20 2440 30 2460
rect -10 2410 30 2440
rect -10 2390 0 2410
rect 20 2390 30 2410
rect -10 2360 30 2390
rect -10 2340 0 2360
rect 20 2340 30 2360
rect -10 2325 30 2340
rect 250 2660 290 2675
rect 250 2640 260 2660
rect 280 2640 290 2660
rect 250 2610 290 2640
rect 250 2590 260 2610
rect 280 2590 290 2610
rect 250 2560 290 2590
rect 930 2660 970 2675
rect 930 2640 940 2660
rect 960 2640 970 2660
rect 930 2610 970 2640
rect 930 2590 940 2610
rect 960 2590 970 2610
rect 930 2560 970 2590
rect 250 2540 260 2560
rect 280 2540 290 2560
rect 250 2510 290 2540
rect 930 2540 940 2560
rect 960 2540 970 2560
rect 250 2490 260 2510
rect 280 2490 290 2510
rect 930 2510 970 2540
rect 250 2460 290 2490
rect 250 2440 260 2460
rect 280 2440 290 2460
rect 250 2410 290 2440
rect 250 2390 260 2410
rect 280 2390 290 2410
rect 250 2360 290 2390
rect 250 2340 260 2360
rect 280 2340 290 2360
rect 250 2325 290 2340
rect 460 2360 500 2505
rect 460 2340 470 2360
rect 490 2340 500 2360
rect 460 2325 500 2340
rect 720 2360 760 2505
rect 720 2340 730 2360
rect 750 2340 760 2360
rect 720 2325 760 2340
rect 930 2490 940 2510
rect 960 2490 970 2510
rect 930 2460 970 2490
rect 930 2440 940 2460
rect 960 2440 970 2460
rect 930 2410 970 2440
rect 930 2390 940 2410
rect 960 2390 970 2410
rect 930 2360 970 2390
rect 930 2340 940 2360
rect 960 2340 970 2360
rect 930 2325 970 2340
rect 1190 2660 1230 2675
rect 1190 2640 1200 2660
rect 1220 2640 1230 2660
rect 1190 2610 1230 2640
rect 1190 2590 1200 2610
rect 1220 2590 1230 2610
rect 1190 2560 1230 2590
rect 1190 2540 1200 2560
rect 1220 2540 1230 2560
rect 1190 2510 1230 2540
rect 1190 2490 1200 2510
rect 1220 2490 1230 2510
rect 1190 2460 1230 2490
rect 1190 2440 1200 2460
rect 1220 2440 1230 2460
rect 1190 2410 1230 2440
rect 1190 2390 1200 2410
rect 1220 2390 1230 2410
rect 1190 2360 1230 2390
rect 1190 2340 1200 2360
rect 1220 2340 1230 2360
rect 1190 2325 1230 2340
rect 1398 2660 1438 2675
rect 1398 2640 1408 2660
rect 1428 2640 1438 2660
rect 1398 2610 1438 2640
rect 1398 2590 1408 2610
rect 1428 2590 1438 2610
rect 1398 2560 1438 2590
rect 1398 2540 1408 2560
rect 1428 2540 1438 2560
rect 1398 2510 1438 2540
rect 1398 2490 1408 2510
rect 1428 2490 1438 2510
rect 1398 2460 1438 2490
rect 1398 2440 1408 2460
rect 1428 2440 1438 2460
rect 1398 2410 1438 2440
rect 1398 2390 1408 2410
rect 1428 2390 1438 2410
rect 1398 2360 1438 2390
rect 1398 2340 1408 2360
rect 1428 2340 1438 2360
rect 1398 2325 1438 2340
rect 1658 2660 1698 2675
rect 1658 2640 1668 2660
rect 1688 2640 1698 2660
rect 1658 2610 1698 2640
rect 1658 2590 1668 2610
rect 1688 2590 1698 2610
rect 1658 2560 1698 2590
rect 1658 2540 1668 2560
rect 1688 2540 1698 2560
rect 1658 2510 1698 2540
rect 1658 2490 1668 2510
rect 1688 2490 1698 2510
rect 1658 2460 1698 2490
rect 1658 2440 1668 2460
rect 1688 2440 1698 2460
rect 1658 2410 1698 2440
rect 1658 2390 1668 2410
rect 1688 2390 1698 2410
rect 1658 2360 1698 2390
rect 1658 2340 1668 2360
rect 1688 2340 1698 2360
rect 1658 2325 1698 2340
rect -1125 2085 -1085 2100
rect -1125 2065 -1115 2085
rect -1095 2065 -1085 2085
rect -1125 2035 -1085 2065
rect -1125 2015 -1115 2035
rect -1095 2015 -1085 2035
rect -1125 1985 -1085 2015
rect -1125 1965 -1115 1985
rect -1095 1965 -1085 1985
rect -1125 1935 -1085 1965
rect -1125 1915 -1115 1935
rect -1095 1915 -1085 1935
rect -1125 1885 -1085 1915
rect -1125 1865 -1115 1885
rect -1095 1865 -1085 1885
rect -1125 1835 -1085 1865
rect -1125 1815 -1115 1835
rect -1095 1815 -1085 1835
rect -1125 1785 -1085 1815
rect -1125 1765 -1115 1785
rect -1095 1765 -1085 1785
rect -1125 1750 -1085 1765
rect -325 2085 -285 2100
rect -325 2065 -315 2085
rect -295 2065 -285 2085
rect -325 2035 -285 2065
rect -325 2015 -315 2035
rect -295 2015 -285 2035
rect -325 1985 -285 2015
rect -325 1965 -315 1985
rect -295 1965 -285 1985
rect -325 1935 -285 1965
rect -325 1915 -315 1935
rect -295 1915 -285 1935
rect -325 1885 -285 1915
rect -325 1865 -315 1885
rect -295 1865 -285 1885
rect -325 1835 -285 1865
rect -325 1815 -315 1835
rect -295 1815 -285 1835
rect -325 1785 -285 1815
rect -325 1765 -315 1785
rect -295 1765 -285 1785
rect -325 1750 -285 1765
rect -80 2085 -40 2100
rect -80 2065 -70 2085
rect -50 2065 -40 2085
rect -80 2035 -40 2065
rect -80 2015 -70 2035
rect -50 2015 -40 2035
rect -80 1985 -40 2015
rect -80 1965 -70 1985
rect -50 1965 -40 1985
rect -80 1935 -40 1965
rect -80 1915 -70 1935
rect -50 1915 -40 1935
rect -80 1885 -40 1915
rect -80 1865 -70 1885
rect -50 1865 -40 1885
rect -80 1835 -40 1865
rect -80 1815 -70 1835
rect -50 1815 -40 1835
rect -80 1785 -40 1815
rect -80 1765 -70 1785
rect -50 1765 -40 1785
rect -80 1750 -40 1765
rect 720 2085 760 2100
rect 720 2065 730 2085
rect 750 2065 760 2085
rect 720 2035 760 2065
rect 720 2015 730 2035
rect 750 2015 760 2035
rect 720 1985 760 2015
rect 720 1965 730 1985
rect 750 1965 760 1985
rect 720 1935 760 1965
rect 720 1915 730 1935
rect 750 1915 760 1935
rect 720 1885 760 1915
rect 720 1865 730 1885
rect 750 1865 760 1885
rect 720 1835 760 1865
rect 720 1815 730 1835
rect 750 1815 760 1835
rect 720 1785 760 1815
rect 720 1765 730 1785
rect 750 1765 760 1785
rect 720 1750 760 1765
rect 930 2085 970 2100
rect 930 2065 940 2085
rect 960 2065 970 2085
rect 930 2035 970 2065
rect 930 2015 940 2035
rect 960 2015 970 2035
rect 930 1985 970 2015
rect 930 1965 940 1985
rect 960 1965 970 1985
rect 930 1935 970 1965
rect 930 1915 940 1935
rect 960 1915 970 1935
rect 930 1885 970 1915
rect 930 1865 940 1885
rect 960 1865 970 1885
rect 930 1835 970 1865
rect 930 1815 940 1835
rect 960 1815 970 1835
rect 930 1785 970 1815
rect 930 1765 940 1785
rect 960 1765 970 1785
rect 930 1750 970 1765
rect 1730 2085 1770 2100
rect 1730 2065 1740 2085
rect 1760 2065 1770 2085
rect 1730 2035 1770 2065
rect 1730 2015 1740 2035
rect 1760 2015 1770 2035
rect 1730 1985 1770 2015
rect 1730 1965 1740 1985
rect 1760 1965 1770 1985
rect 1730 1935 1770 1965
rect 1730 1915 1740 1935
rect 1760 1915 1770 1935
rect 1730 1885 1770 1915
rect 1730 1865 1740 1885
rect 1760 1865 1770 1885
rect 1730 1835 1770 1865
rect 1730 1815 1740 1835
rect 1760 1815 1770 1835
rect 1730 1785 1770 1815
rect 1730 1765 1740 1785
rect 1760 1765 1770 1785
rect 1730 1750 1770 1765
rect 1975 2085 2015 2100
rect 1975 2065 1985 2085
rect 2005 2065 2015 2085
rect 1975 2035 2015 2065
rect 1975 2015 1985 2035
rect 2005 2015 2015 2035
rect 1975 1985 2015 2015
rect 1975 1965 1985 1985
rect 2005 1965 2015 1985
rect 1975 1935 2015 1965
rect 1975 1915 1985 1935
rect 2005 1915 2015 1935
rect 1975 1885 2015 1915
rect 1975 1865 1985 1885
rect 2005 1865 2015 1885
rect 1975 1835 2015 1865
rect 1975 1815 1985 1835
rect 2005 1815 2015 1835
rect 1975 1785 2015 1815
rect 1975 1765 1985 1785
rect 2005 1765 2015 1785
rect 1975 1750 2015 1765
rect 2775 2085 2815 2100
rect 2775 2065 2785 2085
rect 2805 2065 2815 2085
rect 2775 2035 2815 2065
rect 2775 2015 2785 2035
rect 2805 2015 2815 2035
rect 2775 1985 2815 2015
rect 2775 1965 2785 1985
rect 2805 1965 2815 1985
rect 2775 1935 2815 1965
rect 2775 1915 2785 1935
rect 2805 1915 2815 1935
rect 2775 1885 2815 1915
rect 2775 1865 2785 1885
rect 2805 1865 2815 1885
rect 2775 1835 2815 1865
rect 2775 1815 2785 1835
rect 2805 1815 2815 1835
rect 2775 1785 2815 1815
rect 2775 1765 2785 1785
rect 2805 1765 2815 1785
rect 2775 1750 2815 1765
rect 180 1515 220 1530
rect 180 1495 190 1515
rect 210 1495 220 1515
rect 180 1480 220 1495
rect 1470 1515 1510 1530
rect 1470 1495 1480 1515
rect 1500 1495 1510 1515
rect 1470 1480 1510 1495
rect -1095 1420 -1055 1435
rect -1095 1400 -1085 1420
rect -1065 1400 -1055 1420
rect -1095 1370 -1055 1400
rect -1095 1350 -1085 1370
rect -1065 1350 -1055 1370
rect -1095 1320 -1055 1350
rect -1095 1300 -1085 1320
rect -1065 1300 -1055 1320
rect -1095 1270 -1055 1300
rect -1095 1250 -1085 1270
rect -1065 1250 -1055 1270
rect -1095 1220 -1055 1250
rect -1095 1200 -1085 1220
rect -1065 1200 -1055 1220
rect -1095 1170 -1055 1200
rect -1095 1150 -1085 1170
rect -1065 1150 -1055 1170
rect -1095 1120 -1055 1150
rect -1095 1100 -1085 1120
rect -1065 1100 -1055 1120
rect -1095 1070 -1055 1100
rect -1095 1050 -1085 1070
rect -1065 1050 -1055 1070
rect -1095 1020 -1055 1050
rect -1095 1000 -1085 1020
rect -1065 1000 -1055 1020
rect -1095 970 -1055 1000
rect -1095 950 -1085 970
rect -1065 950 -1055 970
rect -1095 920 -1055 950
rect -1095 900 -1085 920
rect -1065 900 -1055 920
rect -1095 870 -1055 900
rect -1095 850 -1085 870
rect -1065 850 -1055 870
rect -1095 835 -1055 850
rect -355 1420 -315 1435
rect 2005 1420 2045 1435
rect -355 1400 -345 1420
rect -325 1400 -315 1420
rect -355 1370 -315 1400
rect -355 1350 -345 1370
rect -325 1350 -315 1370
rect -355 1320 -315 1350
rect -355 1300 -345 1320
rect -325 1300 -315 1320
rect -355 1270 -315 1300
rect -355 1250 -345 1270
rect -325 1250 -315 1270
rect 2005 1400 2015 1420
rect 2035 1400 2045 1420
rect 2005 1370 2045 1400
rect 2005 1350 2015 1370
rect 2035 1350 2045 1370
rect 2005 1320 2045 1350
rect 2005 1300 2015 1320
rect 2035 1300 2045 1320
rect 2005 1270 2045 1300
rect -355 1220 -315 1250
rect 2005 1250 2015 1270
rect 2035 1250 2045 1270
rect -355 1200 -345 1220
rect -325 1200 -315 1220
rect 2005 1220 2045 1250
rect -355 1170 -315 1200
rect -355 1150 -345 1170
rect -325 1150 -315 1170
rect -45 1190 -5 1205
rect -45 1170 -35 1190
rect -15 1170 -5 1190
rect -45 1155 -5 1170
rect 695 1190 735 1205
rect 695 1170 705 1190
rect 725 1170 735 1190
rect 695 1155 735 1170
rect 955 1190 995 1205
rect 955 1170 965 1190
rect 985 1170 995 1190
rect 955 1155 995 1170
rect 1695 1190 1735 1205
rect 1695 1170 1705 1190
rect 1725 1170 1735 1190
rect 1695 1155 1735 1170
rect 2005 1200 2015 1220
rect 2035 1200 2045 1220
rect 2005 1170 2045 1200
rect -355 1120 -315 1150
rect -355 1100 -345 1120
rect -325 1100 -315 1120
rect 2005 1150 2015 1170
rect 2035 1150 2045 1170
rect 2005 1120 2045 1150
rect 2005 1100 2015 1120
rect 2035 1100 2045 1120
rect -355 1070 -315 1100
rect -355 1050 -345 1070
rect -325 1050 -315 1070
rect -355 1020 -315 1050
rect -355 1000 -345 1020
rect -325 1000 -315 1020
rect -355 970 -315 1000
rect -355 950 -345 970
rect -325 950 -315 970
rect -355 920 -315 950
rect 2005 1070 2045 1100
rect 2005 1050 2015 1070
rect 2035 1050 2045 1070
rect 2005 1020 2045 1050
rect 2005 1000 2015 1020
rect 2035 1000 2045 1020
rect 2005 970 2045 1000
rect 2005 950 2015 970
rect 2035 950 2045 970
rect -355 900 -345 920
rect -325 900 -315 920
rect 2005 920 2045 950
rect -355 870 -315 900
rect 2005 900 2015 920
rect 2035 900 2045 920
rect -355 850 -345 870
rect -325 850 -315 870
rect -355 835 -315 850
rect 2005 870 2045 900
rect 2005 850 2015 870
rect 2035 850 2045 870
rect 2005 835 2045 850
rect 2745 1420 2785 1435
rect 2745 1400 2755 1420
rect 2775 1400 2785 1420
rect 2745 1370 2785 1400
rect 2745 1350 2755 1370
rect 2775 1350 2785 1370
rect 2745 1320 2785 1350
rect 2745 1300 2755 1320
rect 2775 1300 2785 1320
rect 2745 1270 2785 1300
rect 2745 1250 2755 1270
rect 2775 1250 2785 1270
rect 2745 1220 2785 1250
rect 2745 1200 2755 1220
rect 2775 1200 2785 1220
rect 2745 1170 2785 1200
rect 2745 1150 2755 1170
rect 2775 1150 2785 1170
rect 2745 1120 2785 1150
rect 2745 1100 2755 1120
rect 2775 1100 2785 1120
rect 2745 1070 2785 1100
rect 2745 1050 2755 1070
rect 2775 1050 2785 1070
rect 2745 1020 2785 1050
rect 2745 1000 2755 1020
rect 2775 1000 2785 1020
rect 2745 970 2785 1000
rect 2745 950 2755 970
rect 2775 950 2785 970
rect 2745 920 2785 950
rect 2745 900 2755 920
rect 2775 900 2785 920
rect 2745 870 2785 900
rect 2745 850 2755 870
rect 2775 850 2785 870
rect 2745 835 2785 850
rect -1095 605 -1055 620
rect -1095 585 -1085 605
rect -1065 585 -1055 605
rect -1095 555 -1055 585
rect -1095 535 -1085 555
rect -1065 535 -1055 555
rect -1095 505 -1055 535
rect -1095 485 -1085 505
rect -1065 485 -1055 505
rect -1095 455 -1055 485
rect -1095 435 -1085 455
rect -1065 435 -1055 455
rect -1095 420 -1055 435
rect -355 605 -315 620
rect 2005 605 2045 620
rect -355 585 -345 605
rect -325 585 -315 605
rect -355 555 -315 585
rect -355 535 -345 555
rect -325 535 -315 555
rect -355 505 -315 535
rect -355 485 -345 505
rect -325 485 -315 505
rect -355 455 -315 485
rect 2005 585 2015 605
rect 2035 585 2045 605
rect 2005 555 2045 585
rect 2005 535 2015 555
rect 2035 535 2045 555
rect 2005 505 2045 535
rect 2005 485 2015 505
rect 2035 485 2045 505
rect 2005 455 2045 485
rect -355 435 -345 455
rect -325 435 -315 455
rect -355 420 -315 435
rect 2005 435 2015 455
rect 2035 435 2045 455
rect 2005 420 2045 435
rect 2745 605 2785 620
rect 2745 585 2755 605
rect 2775 585 2785 605
rect 2745 555 2785 585
rect 2745 535 2755 555
rect 2775 535 2785 555
rect 2745 505 2785 535
rect 2745 485 2755 505
rect 2775 485 2785 505
rect 2745 455 2785 485
rect 2745 435 2755 455
rect 2775 435 2785 455
rect 2745 420 2785 435
<< psubdiffcont >>
rect 465 845 485 865
rect 1205 845 1225 865
rect -55 570 -35 590
rect -55 520 -35 540
rect -55 470 -35 490
rect 685 570 705 590
rect 685 520 705 540
rect 685 470 705 490
rect 985 570 1005 590
rect 985 520 1005 540
rect 985 470 1005 490
rect 1725 570 1745 590
rect 1725 520 1745 540
rect 1725 470 1745 490
rect -1085 195 -1065 215
rect -1085 145 -1065 165
rect -1085 95 -1065 115
rect -1085 45 -1065 65
rect -1085 -5 -1065 15
rect -1085 -55 -1065 -35
rect -345 195 -325 215
rect 2015 195 2035 215
rect -345 145 -325 165
rect 2015 145 2035 165
rect -345 95 -325 115
rect -345 45 -325 65
rect -345 -5 -325 15
rect -55 95 -35 115
rect -55 45 -35 65
rect -55 -5 -35 15
rect 685 95 705 115
rect 685 45 705 65
rect 685 -5 705 15
rect 985 95 1005 115
rect 985 45 1005 65
rect 985 -5 1005 15
rect 1725 95 1745 115
rect 1725 45 1745 65
rect 1725 -5 1745 15
rect 2015 95 2035 115
rect 2015 45 2035 65
rect 2015 -5 2035 15
rect -345 -55 -325 -35
rect 2015 -55 2035 -35
rect 2755 195 2775 215
rect 2755 145 2775 165
rect 2755 95 2775 115
rect 2755 45 2775 65
rect 2755 -5 2775 15
rect 2755 -55 2775 -35
rect -1055 -390 -1035 -370
rect -1055 -440 -1035 -420
rect -1055 -490 -1035 -470
rect -1055 -540 -1035 -520
rect -1055 -590 -1035 -570
rect -1055 -640 -1035 -620
rect -1055 -690 -1035 -670
rect -1055 -740 -1035 -720
rect -1055 -790 -1035 -770
rect -1055 -840 -1035 -820
rect -1055 -890 -1035 -870
rect -1055 -940 -1035 -920
rect -1055 -990 -1035 -970
rect -1055 -1040 -1035 -1020
rect -375 -390 -355 -370
rect 2045 -390 2065 -370
rect -375 -440 -355 -420
rect -375 -490 -355 -470
rect -375 -540 -355 -520
rect -375 -590 -355 -570
rect -375 -640 -355 -620
rect 130 -440 150 -420
rect 130 -490 150 -470
rect 130 -540 150 -520
rect 130 -590 150 -570
rect 130 -640 150 -620
rect 1475 -440 1495 -420
rect 1475 -490 1495 -470
rect 1475 -540 1495 -520
rect 1475 -590 1495 -570
rect 1475 -640 1495 -620
rect 2045 -440 2065 -420
rect 2045 -490 2065 -470
rect 2045 -540 2065 -520
rect 2045 -590 2065 -570
rect 2045 -640 2065 -620
rect -375 -690 -355 -670
rect 2045 -690 2065 -670
rect -375 -740 -355 -720
rect 2045 -740 2065 -720
rect -375 -790 -355 -770
rect 2045 -790 2065 -770
rect -375 -840 -355 -820
rect -375 -890 -355 -870
rect 2045 -840 2065 -820
rect 2045 -890 2065 -870
rect -375 -940 -355 -920
rect -375 -990 -355 -970
rect -375 -1040 -355 -1020
rect 2045 -940 2065 -920
rect 2045 -990 2065 -970
rect 2045 -1040 2065 -1020
rect 2725 -390 2745 -370
rect 2725 -440 2745 -420
rect 2725 -490 2745 -470
rect 2725 -540 2745 -520
rect 2725 -590 2745 -570
rect 2725 -640 2745 -620
rect 2725 -690 2745 -670
rect 2725 -740 2745 -720
rect 2725 -790 2745 -770
rect 2725 -840 2745 -820
rect 2725 -890 2745 -870
rect 2725 -940 2745 -920
rect 2725 -990 2745 -970
rect 2725 -1040 2745 -1020
<< nsubdiffcont >>
rect 0 2640 20 2660
rect 0 2590 20 2610
rect 0 2540 20 2560
rect 0 2490 20 2510
rect 0 2440 20 2460
rect 0 2390 20 2410
rect 0 2340 20 2360
rect 260 2640 280 2660
rect 260 2590 280 2610
rect 940 2640 960 2660
rect 940 2590 960 2610
rect 260 2540 280 2560
rect 940 2540 960 2560
rect 260 2490 280 2510
rect 260 2440 280 2460
rect 260 2390 280 2410
rect 260 2340 280 2360
rect 470 2340 490 2360
rect 730 2340 750 2360
rect 940 2490 960 2510
rect 940 2440 960 2460
rect 940 2390 960 2410
rect 940 2340 960 2360
rect 1200 2640 1220 2660
rect 1200 2590 1220 2610
rect 1200 2540 1220 2560
rect 1200 2490 1220 2510
rect 1200 2440 1220 2460
rect 1200 2390 1220 2410
rect 1200 2340 1220 2360
rect 1408 2640 1428 2660
rect 1408 2590 1428 2610
rect 1408 2540 1428 2560
rect 1408 2490 1428 2510
rect 1408 2440 1428 2460
rect 1408 2390 1428 2410
rect 1408 2340 1428 2360
rect 1668 2640 1688 2660
rect 1668 2590 1688 2610
rect 1668 2540 1688 2560
rect 1668 2490 1688 2510
rect 1668 2440 1688 2460
rect 1668 2390 1688 2410
rect 1668 2340 1688 2360
rect -1115 2065 -1095 2085
rect -1115 2015 -1095 2035
rect -1115 1965 -1095 1985
rect -1115 1915 -1095 1935
rect -1115 1865 -1095 1885
rect -1115 1815 -1095 1835
rect -1115 1765 -1095 1785
rect -315 2065 -295 2085
rect -315 2015 -295 2035
rect -315 1965 -295 1985
rect -315 1915 -295 1935
rect -315 1865 -295 1885
rect -315 1815 -295 1835
rect -315 1765 -295 1785
rect -70 2065 -50 2085
rect -70 2015 -50 2035
rect -70 1965 -50 1985
rect -70 1915 -50 1935
rect -70 1865 -50 1885
rect -70 1815 -50 1835
rect -70 1765 -50 1785
rect 730 2065 750 2085
rect 730 2015 750 2035
rect 730 1965 750 1985
rect 730 1915 750 1935
rect 730 1865 750 1885
rect 730 1815 750 1835
rect 730 1765 750 1785
rect 940 2065 960 2085
rect 940 2015 960 2035
rect 940 1965 960 1985
rect 940 1915 960 1935
rect 940 1865 960 1885
rect 940 1815 960 1835
rect 940 1765 960 1785
rect 1740 2065 1760 2085
rect 1740 2015 1760 2035
rect 1740 1965 1760 1985
rect 1740 1915 1760 1935
rect 1740 1865 1760 1885
rect 1740 1815 1760 1835
rect 1740 1765 1760 1785
rect 1985 2065 2005 2085
rect 1985 2015 2005 2035
rect 1985 1965 2005 1985
rect 1985 1915 2005 1935
rect 1985 1865 2005 1885
rect 1985 1815 2005 1835
rect 1985 1765 2005 1785
rect 2785 2065 2805 2085
rect 2785 2015 2805 2035
rect 2785 1965 2805 1985
rect 2785 1915 2805 1935
rect 2785 1865 2805 1885
rect 2785 1815 2805 1835
rect 2785 1765 2805 1785
rect 190 1495 210 1515
rect 1480 1495 1500 1515
rect -1085 1400 -1065 1420
rect -1085 1350 -1065 1370
rect -1085 1300 -1065 1320
rect -1085 1250 -1065 1270
rect -1085 1200 -1065 1220
rect -1085 1150 -1065 1170
rect -1085 1100 -1065 1120
rect -1085 1050 -1065 1070
rect -1085 1000 -1065 1020
rect -1085 950 -1065 970
rect -1085 900 -1065 920
rect -1085 850 -1065 870
rect -345 1400 -325 1420
rect -345 1350 -325 1370
rect -345 1300 -325 1320
rect -345 1250 -325 1270
rect 2015 1400 2035 1420
rect 2015 1350 2035 1370
rect 2015 1300 2035 1320
rect 2015 1250 2035 1270
rect -345 1200 -325 1220
rect -345 1150 -325 1170
rect -35 1170 -15 1190
rect 705 1170 725 1190
rect 965 1170 985 1190
rect 1705 1170 1725 1190
rect 2015 1200 2035 1220
rect -345 1100 -325 1120
rect 2015 1150 2035 1170
rect 2015 1100 2035 1120
rect -345 1050 -325 1070
rect -345 1000 -325 1020
rect -345 950 -325 970
rect 2015 1050 2035 1070
rect 2015 1000 2035 1020
rect 2015 950 2035 970
rect -345 900 -325 920
rect 2015 900 2035 920
rect -345 850 -325 870
rect 2015 850 2035 870
rect 2755 1400 2775 1420
rect 2755 1350 2775 1370
rect 2755 1300 2775 1320
rect 2755 1250 2775 1270
rect 2755 1200 2775 1220
rect 2755 1150 2775 1170
rect 2755 1100 2775 1120
rect 2755 1050 2775 1070
rect 2755 1000 2775 1020
rect 2755 950 2775 970
rect 2755 900 2775 920
rect 2755 850 2775 870
rect -1085 585 -1065 605
rect -1085 535 -1065 555
rect -1085 485 -1065 505
rect -1085 435 -1065 455
rect -345 585 -325 605
rect -345 535 -325 555
rect -345 485 -325 505
rect 2015 585 2035 605
rect 2015 535 2035 555
rect 2015 485 2035 505
rect -345 435 -325 455
rect 2015 435 2035 455
rect 2755 585 2775 605
rect 2755 535 2775 555
rect 2755 485 2775 505
rect 2755 435 2775 455
<< poly >>
rect 30 2720 70 2730
rect 30 2700 40 2720
rect 60 2705 70 2720
rect 210 2720 250 2730
rect 210 2705 220 2720
rect 60 2700 90 2705
rect 30 2690 90 2700
rect 190 2700 220 2705
rect 240 2700 250 2720
rect 190 2690 250 2700
rect 970 2720 1010 2730
rect 970 2700 980 2720
rect 1000 2705 1010 2720
rect 1150 2720 1190 2730
rect 1150 2705 1160 2720
rect 1000 2700 1030 2705
rect 970 2690 1030 2700
rect 1130 2700 1160 2705
rect 1180 2700 1190 2720
rect 1130 2690 1190 2700
rect 1438 2720 1478 2730
rect 1438 2700 1448 2720
rect 1468 2705 1478 2720
rect 1618 2720 1658 2730
rect 1618 2705 1628 2720
rect 1468 2700 1498 2705
rect 1438 2690 1498 2700
rect 1598 2700 1628 2705
rect 1648 2700 1658 2720
rect 1598 2690 1658 2700
rect 70 2675 90 2690
rect 130 2675 150 2690
rect 190 2675 210 2690
rect 1010 2675 1030 2690
rect 1070 2675 1090 2690
rect 1130 2675 1150 2690
rect 1478 2675 1498 2690
rect 1538 2675 1558 2690
rect 1598 2675 1618 2690
rect 500 2550 540 2560
rect 500 2530 510 2550
rect 530 2535 540 2550
rect 680 2550 720 2560
rect 680 2535 690 2550
rect 530 2530 560 2535
rect 500 2520 560 2530
rect 660 2530 690 2535
rect 710 2530 720 2550
rect 660 2520 720 2530
rect 540 2505 560 2520
rect 600 2505 620 2520
rect 660 2505 680 2520
rect 70 2310 90 2325
rect 130 2310 150 2325
rect 190 2310 210 2325
rect 540 2310 560 2325
rect 600 2310 620 2325
rect 660 2310 680 2325
rect 1010 2310 1030 2325
rect 1070 2310 1090 2325
rect 1130 2310 1150 2325
rect 1478 2310 1498 2325
rect 1538 2310 1558 2325
rect 1598 2310 1618 2325
rect 130 2300 169 2310
rect 130 2295 144 2300
rect 139 2280 144 2295
rect 164 2280 169 2300
rect 600 2300 639 2310
rect 600 2295 614 2300
rect 139 2270 169 2280
rect 609 2280 614 2295
rect 634 2280 639 2300
rect 609 2270 639 2280
rect 1051 2300 1090 2310
rect 1051 2280 1056 2300
rect 1076 2295 1090 2300
rect 1519 2300 1558 2310
rect 1076 2280 1081 2295
rect 1051 2270 1081 2280
rect 1519 2280 1524 2300
rect 1544 2295 1558 2300
rect 1544 2280 1549 2295
rect 1519 2270 1549 2280
rect -1085 2145 -1045 2155
rect -1085 2125 -1075 2145
rect -1055 2130 -1045 2145
rect -365 2145 -325 2155
rect -365 2130 -355 2145
rect -1055 2125 -1025 2130
rect -1085 2115 -1025 2125
rect -385 2125 -355 2130
rect -335 2125 -325 2145
rect -385 2115 -325 2125
rect -40 2145 0 2155
rect -40 2125 -30 2145
rect -10 2130 0 2145
rect 680 2145 720 2155
rect 680 2130 690 2145
rect -10 2125 20 2130
rect -40 2115 20 2125
rect 660 2125 690 2130
rect 710 2125 720 2145
rect 660 2115 720 2125
rect 970 2145 1010 2155
rect 970 2125 980 2145
rect 1000 2130 1010 2145
rect 1690 2145 1730 2155
rect 1690 2130 1700 2145
rect 1000 2125 1030 2130
rect 970 2115 1030 2125
rect 1670 2125 1700 2130
rect 1720 2125 1730 2145
rect 1670 2115 1730 2125
rect 2015 2145 2055 2155
rect 2015 2125 2025 2145
rect 2045 2130 2055 2145
rect 2735 2145 2775 2155
rect 2735 2130 2745 2145
rect 2045 2125 2075 2130
rect 2015 2115 2075 2125
rect 2715 2125 2745 2130
rect 2765 2125 2775 2145
rect 2715 2115 2775 2125
rect -1045 2100 -1025 2115
rect -985 2100 -965 2115
rect -925 2100 -905 2115
rect -865 2100 -845 2115
rect -805 2100 -785 2115
rect -745 2100 -725 2115
rect -685 2100 -665 2115
rect -625 2100 -605 2115
rect -565 2100 -545 2115
rect -505 2100 -485 2115
rect -445 2100 -425 2115
rect -385 2100 -365 2115
rect 0 2100 20 2115
rect 60 2100 80 2115
rect 120 2100 140 2115
rect 180 2100 200 2115
rect 240 2100 260 2115
rect 300 2100 320 2115
rect 360 2100 380 2115
rect 420 2100 440 2115
rect 480 2100 500 2115
rect 540 2100 560 2115
rect 600 2100 620 2115
rect 660 2100 680 2115
rect 1010 2100 1030 2115
rect 1070 2100 1090 2115
rect 1130 2100 1150 2115
rect 1190 2100 1210 2115
rect 1250 2100 1270 2115
rect 1310 2100 1330 2115
rect 1370 2100 1390 2115
rect 1430 2100 1450 2115
rect 1490 2100 1510 2115
rect 1550 2100 1570 2115
rect 1610 2100 1630 2115
rect 1670 2100 1690 2115
rect 2055 2100 2075 2115
rect 2115 2100 2135 2115
rect 2175 2100 2195 2115
rect 2235 2100 2255 2115
rect 2295 2100 2315 2115
rect 2355 2100 2375 2115
rect 2415 2100 2435 2115
rect 2475 2100 2495 2115
rect 2535 2100 2555 2115
rect 2595 2100 2615 2115
rect 2655 2100 2675 2115
rect 2715 2100 2735 2115
rect -1045 1735 -1025 1750
rect -985 1740 -965 1750
rect -925 1740 -905 1750
rect -865 1740 -845 1750
rect -805 1740 -785 1750
rect -745 1740 -725 1750
rect -685 1740 -665 1750
rect -625 1740 -605 1750
rect -565 1740 -545 1750
rect -505 1740 -485 1750
rect -445 1740 -425 1750
rect -985 1725 -425 1740
rect -385 1735 -365 1750
rect 0 1735 20 1750
rect 60 1740 80 1750
rect 120 1740 140 1750
rect 180 1740 200 1750
rect 240 1740 260 1750
rect 300 1740 320 1750
rect 360 1740 380 1750
rect 420 1740 440 1750
rect 480 1740 500 1750
rect 540 1740 560 1750
rect 600 1740 620 1750
rect 60 1725 620 1740
rect 660 1735 680 1750
rect 1010 1735 1030 1750
rect 1070 1740 1090 1750
rect 1130 1740 1150 1750
rect 1190 1740 1210 1750
rect 1250 1740 1270 1750
rect 1310 1740 1330 1750
rect 1370 1740 1390 1750
rect 1430 1740 1450 1750
rect 1490 1740 1510 1750
rect 1550 1740 1570 1750
rect 1610 1740 1630 1750
rect 1070 1725 1630 1740
rect 1670 1735 1690 1750
rect 2055 1735 2075 1750
rect 2115 1740 2135 1750
rect 2175 1740 2195 1750
rect 2235 1740 2255 1750
rect 2295 1740 2315 1750
rect 2355 1740 2375 1750
rect 2415 1740 2435 1750
rect 2475 1740 2495 1750
rect 2535 1740 2555 1750
rect 2595 1740 2615 1750
rect 2655 1740 2675 1750
rect 2115 1725 2675 1740
rect 2715 1735 2735 1750
rect -720 1720 -690 1725
rect -720 1700 -715 1720
rect -695 1700 -690 1720
rect -720 1690 -690 1700
rect 325 1720 355 1725
rect 325 1700 330 1720
rect 350 1700 355 1720
rect 325 1690 355 1700
rect 1335 1720 1365 1725
rect 1335 1700 1340 1720
rect 1360 1700 1365 1720
rect 1335 1690 1365 1700
rect 2380 1720 2410 1725
rect 2380 1700 2385 1720
rect 2405 1700 2410 1720
rect 2380 1690 2410 1700
rect 220 1575 260 1585
rect 220 1555 230 1575
rect 250 1560 260 1575
rect 1430 1575 1470 1585
rect 1430 1560 1440 1575
rect 250 1555 275 1560
rect 220 1545 275 1555
rect 1415 1555 1440 1560
rect 1460 1555 1470 1575
rect 1415 1545 1470 1555
rect 260 1530 275 1545
rect 315 1530 330 1545
rect 370 1530 385 1545
rect 425 1530 440 1545
rect 480 1530 495 1545
rect 535 1530 550 1545
rect 590 1530 605 1545
rect 645 1530 660 1545
rect 700 1530 715 1545
rect 755 1530 770 1545
rect 810 1530 825 1545
rect 865 1530 880 1545
rect 920 1530 935 1545
rect 975 1530 990 1545
rect 1030 1530 1045 1545
rect 1085 1530 1100 1545
rect 1140 1530 1155 1545
rect 1195 1530 1210 1545
rect 1250 1530 1265 1545
rect 1305 1530 1320 1545
rect 1360 1530 1375 1545
rect 1415 1530 1430 1545
rect -1055 1480 -1015 1490
rect -1055 1460 -1045 1480
rect -1025 1465 -1015 1480
rect -395 1480 -355 1490
rect 2045 1480 2085 1490
rect -395 1465 -385 1480
rect -1025 1460 -1000 1465
rect -1055 1450 -1000 1460
rect -410 1460 -385 1465
rect -365 1460 -355 1480
rect 260 1465 275 1480
rect 315 1470 330 1480
rect 370 1470 385 1480
rect 425 1470 440 1480
rect 480 1470 495 1480
rect 535 1470 550 1480
rect 590 1470 605 1480
rect 645 1470 660 1480
rect 700 1470 715 1480
rect 755 1470 770 1480
rect 810 1470 825 1480
rect 865 1470 880 1480
rect 920 1470 935 1480
rect 975 1470 990 1480
rect 1030 1470 1045 1480
rect 1085 1470 1100 1480
rect 1140 1470 1155 1480
rect 1195 1470 1210 1480
rect 1250 1470 1265 1480
rect 1305 1470 1320 1480
rect 1360 1470 1375 1480
rect -410 1450 -355 1460
rect 315 1455 1375 1470
rect 1415 1455 1430 1480
rect 2045 1460 2055 1480
rect 2075 1465 2085 1480
rect 2705 1480 2745 1490
rect 2705 1465 2715 1480
rect 2075 1460 2100 1465
rect 885 1450 915 1455
rect 2045 1450 2100 1460
rect 2690 1460 2715 1465
rect 2735 1460 2745 1480
rect 2690 1450 2745 1460
rect -1015 1435 -1000 1450
rect -960 1435 -945 1450
rect -905 1435 -890 1450
rect -850 1435 -835 1450
rect -795 1435 -780 1450
rect -740 1435 -725 1450
rect -685 1435 -670 1450
rect -630 1435 -615 1450
rect -575 1435 -560 1450
rect -520 1435 -505 1450
rect -465 1435 -450 1450
rect -410 1435 -395 1450
rect 885 1430 890 1450
rect 910 1430 915 1450
rect 2085 1435 2100 1450
rect 2140 1435 2155 1450
rect 2195 1435 2210 1450
rect 2250 1435 2265 1450
rect 2305 1435 2320 1450
rect 2360 1435 2375 1450
rect 2415 1435 2430 1450
rect 2470 1435 2485 1450
rect 2525 1435 2540 1450
rect 2580 1435 2595 1450
rect 2635 1435 2650 1450
rect 2690 1435 2705 1450
rect 885 1420 915 1430
rect 71 1250 101 1260
rect 71 1230 76 1250
rect 96 1235 101 1250
rect 275 1250 305 1260
rect 96 1230 105 1235
rect 275 1230 280 1250
rect 300 1230 305 1250
rect 495 1250 525 1260
rect 495 1230 500 1250
rect 520 1230 525 1250
rect 1071 1250 1101 1260
rect 1071 1230 1076 1250
rect 1096 1235 1101 1250
rect 1275 1250 1305 1260
rect 1096 1230 1105 1235
rect 1275 1230 1280 1250
rect 1300 1230 1305 1250
rect 1495 1250 1525 1260
rect 1495 1230 1500 1250
rect 1520 1230 1525 1250
rect 71 1220 105 1230
rect 35 1205 50 1220
rect 90 1205 105 1220
rect 145 1205 160 1220
rect 200 1205 215 1220
rect 255 1215 325 1230
rect 255 1205 270 1215
rect 310 1205 325 1215
rect 365 1205 380 1220
rect 420 1205 435 1220
rect 475 1215 545 1230
rect 1071 1220 1105 1230
rect 475 1205 490 1215
rect 530 1205 545 1215
rect 585 1205 600 1220
rect 640 1205 655 1220
rect 1035 1205 1050 1220
rect 1090 1205 1105 1220
rect 1145 1205 1160 1220
rect 1200 1205 1215 1220
rect 1255 1215 1325 1230
rect 1255 1205 1270 1215
rect 1310 1205 1325 1215
rect 1365 1205 1380 1220
rect 1420 1205 1435 1220
rect 1475 1215 1545 1230
rect 1475 1205 1490 1215
rect 1530 1205 1545 1215
rect 1585 1205 1600 1220
rect 1640 1205 1655 1220
rect 35 1145 50 1155
rect -5 1130 50 1145
rect 90 1140 105 1155
rect 145 1145 160 1155
rect 200 1145 215 1155
rect 145 1141 215 1145
rect 145 1131 234 1141
rect 255 1140 270 1155
rect 310 1140 325 1155
rect 365 1145 380 1155
rect 420 1145 435 1155
rect 365 1141 435 1145
rect 145 1130 209 1131
rect -5 1110 0 1130
rect 20 1110 25 1130
rect -5 1100 25 1110
rect 204 1111 209 1130
rect 229 1111 234 1131
rect 365 1131 454 1141
rect 475 1140 490 1155
rect 530 1140 545 1155
rect 585 1141 600 1155
rect 365 1125 429 1131
rect 204 1101 234 1111
rect 424 1111 429 1125
rect 449 1111 454 1131
rect 424 1101 454 1111
rect 566 1131 600 1141
rect 566 1111 571 1131
rect 591 1125 600 1131
rect 640 1145 655 1155
rect 1035 1145 1050 1155
rect 640 1130 695 1145
rect 591 1111 596 1125
rect 566 1101 596 1111
rect 665 1110 670 1130
rect 690 1110 695 1130
rect 665 1100 695 1110
rect 995 1130 1050 1145
rect 1090 1140 1105 1155
rect 1145 1145 1160 1155
rect 1200 1145 1215 1155
rect 1145 1141 1215 1145
rect 1145 1131 1234 1141
rect 1255 1140 1270 1155
rect 1310 1140 1325 1155
rect 1365 1145 1380 1155
rect 1420 1145 1435 1155
rect 1365 1141 1435 1145
rect 1145 1130 1209 1131
rect 995 1110 1000 1130
rect 1020 1110 1025 1130
rect 995 1100 1025 1110
rect 1204 1111 1209 1130
rect 1229 1111 1234 1131
rect 1365 1131 1454 1141
rect 1475 1140 1490 1155
rect 1530 1140 1545 1155
rect 1585 1141 1600 1155
rect 1365 1125 1429 1131
rect 1204 1101 1234 1111
rect 1424 1111 1429 1125
rect 1449 1111 1454 1131
rect 1424 1101 1454 1111
rect 1566 1131 1600 1141
rect 1566 1111 1571 1131
rect 1591 1125 1600 1131
rect 1640 1145 1655 1155
rect 1640 1130 1695 1145
rect 1591 1111 1596 1125
rect 1566 1101 1596 1111
rect 1665 1110 1670 1130
rect 1690 1110 1695 1130
rect 1665 1100 1695 1110
rect 660 925 700 935
rect 660 905 670 925
rect 690 905 700 925
rect 880 925 920 935
rect 880 905 890 925
rect 910 905 920 925
rect 535 880 550 895
rect 590 890 1100 905
rect 590 880 605 890
rect 645 880 660 890
rect 700 880 715 890
rect 755 880 770 890
rect 810 880 825 890
rect 865 880 880 890
rect 920 880 935 890
rect 975 880 990 890
rect 1030 880 1045 890
rect 1085 880 1100 890
rect 1140 880 1155 895
rect -1015 820 -1000 835
rect -960 825 -945 835
rect -905 825 -890 835
rect -850 825 -835 835
rect -795 825 -780 835
rect -740 825 -725 835
rect -685 825 -670 835
rect -630 825 -615 835
rect -575 825 -560 835
rect -520 825 -505 835
rect -465 825 -450 835
rect -960 810 -450 825
rect -410 820 -395 835
rect 535 815 550 830
rect 590 815 605 830
rect 645 815 660 830
rect 700 815 715 830
rect 755 815 770 830
rect 810 815 825 830
rect 865 815 880 830
rect 920 815 935 830
rect 975 815 990 830
rect 1030 815 1045 830
rect 1085 815 1100 830
rect 1140 815 1155 830
rect 2085 820 2100 835
rect 2140 825 2155 835
rect 2195 825 2210 835
rect 2250 825 2265 835
rect 2305 825 2320 835
rect 2360 825 2375 835
rect 2415 825 2430 835
rect 2470 825 2485 835
rect 2525 825 2540 835
rect 2580 825 2595 835
rect 2635 825 2650 835
rect -720 800 -690 810
rect -720 780 -715 800
rect -695 780 -690 800
rect -720 770 -690 780
rect 495 805 550 815
rect 495 785 505 805
rect 525 800 550 805
rect 1140 805 1195 815
rect 2140 810 2650 825
rect 2690 820 2705 835
rect 1140 800 1165 805
rect 525 785 535 800
rect 495 775 535 785
rect 1155 785 1165 800
rect 1185 785 1195 805
rect 1155 775 1195 785
rect 2380 800 2410 810
rect 2380 780 2385 800
rect 2405 780 2410 800
rect 2380 770 2410 780
rect -1065 665 -1025 675
rect -1065 645 -1055 665
rect -1035 650 -1025 665
rect -385 665 -345 675
rect 2035 665 2075 675
rect -385 650 -375 665
rect -1035 645 -1000 650
rect -1065 635 -1000 645
rect -410 645 -375 650
rect -355 645 -345 665
rect -410 635 -345 645
rect 310 655 340 665
rect 310 635 315 655
rect 335 635 340 655
rect -1015 620 -1000 635
rect -960 620 -945 635
rect -905 620 -890 635
rect -850 620 -835 635
rect -795 620 -780 635
rect -740 620 -725 635
rect -685 620 -670 635
rect -630 620 -615 635
rect -575 620 -560 635
rect -520 620 -505 635
rect -465 620 -450 635
rect -410 620 -395 635
rect 310 630 340 635
rect 1350 655 1380 665
rect 1350 635 1355 655
rect 1375 635 1380 655
rect 2035 645 2045 665
rect 2065 650 2075 665
rect 2715 665 2755 675
rect 2715 650 2725 665
rect 2065 645 2100 650
rect 2035 635 2100 645
rect 2690 645 2725 650
rect 2745 645 2755 665
rect 2690 635 2755 645
rect 1350 630 1380 635
rect 15 605 30 620
rect 70 615 580 630
rect 70 605 85 615
rect 125 605 140 615
rect 180 605 195 615
rect 235 605 250 615
rect 290 605 305 615
rect 345 605 360 615
rect 400 605 415 615
rect 455 605 470 615
rect 510 605 525 615
rect 565 605 580 615
rect 620 605 635 620
rect 1055 605 1070 620
rect 1110 615 1620 630
rect 2085 620 2100 635
rect 2140 620 2155 635
rect 2195 620 2210 635
rect 2250 620 2265 635
rect 2305 620 2320 635
rect 2360 620 2375 635
rect 2415 620 2430 635
rect 2470 620 2485 635
rect 2525 620 2540 635
rect 2580 620 2595 635
rect 2635 620 2650 635
rect 2690 620 2705 635
rect 1110 605 1125 615
rect 1165 605 1180 615
rect 1220 605 1235 615
rect 1275 605 1290 615
rect 1330 605 1345 615
rect 1385 605 1400 615
rect 1440 605 1455 615
rect 1495 605 1510 615
rect 1550 605 1565 615
rect 1605 605 1620 615
rect 1660 605 1675 620
rect 15 440 30 455
rect 70 440 85 455
rect 125 440 140 455
rect 180 440 195 455
rect 235 440 250 455
rect 290 440 305 455
rect 345 440 360 455
rect 400 440 415 455
rect 455 440 470 455
rect 510 440 525 455
rect 565 440 580 455
rect 620 440 635 455
rect 1055 440 1070 455
rect 1110 440 1125 455
rect 1165 440 1180 455
rect 1220 440 1235 455
rect 1275 440 1290 455
rect 1330 440 1345 455
rect 1385 440 1400 455
rect 1440 440 1455 455
rect 1495 440 1510 455
rect 1550 440 1565 455
rect 1605 440 1620 455
rect 1660 440 1675 455
rect -25 430 30 440
rect -1015 405 -1000 420
rect -960 410 -945 420
rect -905 410 -890 420
rect -850 410 -835 420
rect -795 410 -780 420
rect -740 410 -725 420
rect -685 410 -670 420
rect -630 410 -615 420
rect -575 410 -560 420
rect -520 410 -505 420
rect -465 410 -450 420
rect -960 395 -450 410
rect -410 405 -395 420
rect -25 410 -15 430
rect 5 425 30 430
rect 620 430 675 440
rect 620 425 645 430
rect 5 410 15 425
rect -25 400 15 410
rect 635 410 645 425
rect 665 410 675 430
rect 635 400 675 410
rect 1015 430 1070 440
rect 1015 410 1025 430
rect 1045 425 1070 430
rect 1660 430 1715 440
rect 1660 425 1685 430
rect 1045 410 1055 425
rect 1015 400 1055 410
rect 1675 410 1685 425
rect 1705 410 1715 430
rect 1675 400 1715 410
rect 2085 405 2100 420
rect 2140 410 2155 420
rect 2195 410 2210 420
rect 2250 410 2265 420
rect 2305 410 2320 420
rect 2360 410 2375 420
rect 2415 410 2430 420
rect 2470 410 2485 420
rect 2525 410 2540 420
rect 2580 410 2595 420
rect 2635 410 2650 420
rect 2140 395 2650 410
rect 2690 405 2705 420
rect -665 390 -635 395
rect -665 370 -660 390
rect -640 370 -635 390
rect -665 360 -635 370
rect 2325 390 2355 395
rect 2325 370 2330 390
rect 2350 370 2355 390
rect 2325 360 2355 370
rect -665 280 -635 290
rect -665 260 -660 280
rect -640 260 -635 280
rect -665 255 -635 260
rect 2325 280 2355 290
rect 2325 260 2330 280
rect 2350 260 2355 280
rect 2325 255 2355 260
rect -1015 230 -1000 245
rect -960 240 -450 255
rect -960 230 -945 240
rect -905 230 -890 240
rect -850 230 -835 240
rect -795 230 -780 240
rect -740 230 -725 240
rect -685 230 -670 240
rect -630 230 -615 240
rect -575 230 -560 240
rect -520 230 -505 240
rect -465 230 -450 240
rect -410 230 -395 245
rect 2085 230 2100 245
rect 2140 240 2650 255
rect 2140 230 2155 240
rect 2195 230 2210 240
rect 2250 230 2265 240
rect 2305 230 2320 240
rect 2360 230 2375 240
rect 2415 230 2430 240
rect 2470 230 2485 240
rect 2525 230 2540 240
rect 2580 230 2595 240
rect 2635 230 2650 240
rect 2690 230 2705 245
rect 310 175 340 185
rect 310 155 315 175
rect 335 155 340 175
rect 795 175 825 185
rect 795 155 800 175
rect 820 155 825 175
rect 15 130 30 145
rect 70 140 580 155
rect 795 145 825 155
rect 848 175 878 185
rect 848 155 853 175
rect 873 155 878 175
rect 1350 175 1380 185
rect 1350 155 1355 175
rect 1375 155 1380 175
rect 848 145 880 155
rect 70 130 85 140
rect 125 130 140 140
rect 180 130 195 140
rect 235 130 250 140
rect 290 130 305 140
rect 345 130 360 140
rect 400 130 415 140
rect 455 130 470 140
rect 510 130 525 140
rect 565 130 580 140
rect 620 130 635 145
rect 755 130 770 145
rect 810 130 825 145
rect 865 130 880 145
rect 920 130 935 145
rect 1055 130 1070 145
rect 1110 140 1620 155
rect 1110 130 1125 140
rect 1165 130 1180 140
rect 1220 130 1235 140
rect 1275 130 1290 140
rect 1330 130 1345 140
rect 1385 130 1400 140
rect 1440 130 1455 140
rect 1495 130 1510 140
rect 1550 130 1565 140
rect 1605 130 1620 140
rect 1660 130 1675 145
rect 15 -35 30 -20
rect 70 -35 85 -20
rect 125 -35 140 -20
rect 180 -35 195 -20
rect 235 -35 250 -20
rect 290 -35 305 -20
rect 345 -35 360 -20
rect 400 -35 415 -20
rect 455 -35 470 -20
rect 510 -35 525 -20
rect 565 -35 580 -20
rect 620 -35 635 -20
rect 755 -35 770 -20
rect 810 -35 825 -20
rect 865 -35 880 -20
rect 920 -35 935 -20
rect 1055 -35 1070 -20
rect 1110 -35 1125 -20
rect 1165 -35 1180 -20
rect 1220 -35 1235 -20
rect 1275 -35 1290 -20
rect 1330 -35 1345 -20
rect 1385 -35 1400 -20
rect 1440 -35 1455 -20
rect 1495 -35 1510 -20
rect 1550 -35 1565 -20
rect 1605 -35 1620 -20
rect 1660 -35 1675 -20
rect -20 -45 30 -35
rect -20 -65 -15 -45
rect 5 -50 30 -45
rect 620 -45 770 -35
rect 620 -50 685 -45
rect 5 -65 10 -50
rect -1015 -85 -1000 -70
rect -960 -85 -945 -70
rect -905 -85 -890 -70
rect -850 -85 -835 -70
rect -795 -85 -780 -70
rect -740 -85 -725 -70
rect -685 -85 -670 -70
rect -630 -85 -615 -70
rect -575 -85 -560 -70
rect -520 -85 -505 -70
rect -465 -85 -450 -70
rect -410 -85 -395 -70
rect -20 -75 10 -65
rect 680 -65 685 -50
rect 705 -50 770 -45
rect 920 -45 1070 -35
rect 920 -50 985 -45
rect 705 -65 710 -50
rect 680 -75 710 -65
rect 980 -65 985 -50
rect 1005 -50 1070 -45
rect 1660 -45 1710 -35
rect 1660 -50 1685 -45
rect 1005 -65 1010 -50
rect 980 -75 1010 -65
rect 1680 -65 1685 -50
rect 1705 -65 1710 -45
rect 1680 -75 1710 -65
rect 2085 -85 2100 -70
rect 2140 -85 2155 -70
rect 2195 -85 2210 -70
rect 2250 -85 2265 -70
rect 2305 -85 2320 -70
rect 2360 -85 2375 -70
rect 2415 -85 2430 -70
rect 2470 -85 2485 -70
rect 2525 -85 2540 -70
rect 2580 -85 2595 -70
rect 2635 -85 2650 -70
rect 2690 -85 2705 -70
rect -1065 -95 -1000 -85
rect -1065 -115 -1055 -95
rect -1035 -100 -1000 -95
rect -410 -95 -345 -85
rect -410 -100 -375 -95
rect -1035 -115 -1025 -100
rect -1065 -125 -1025 -115
rect -385 -115 -375 -100
rect -355 -115 -345 -95
rect -385 -125 -345 -115
rect 2035 -95 2100 -85
rect 2035 -115 2045 -95
rect 2065 -100 2100 -95
rect 2690 -95 2755 -85
rect 2690 -100 2725 -95
rect 2065 -115 2075 -100
rect 2035 -125 2075 -115
rect 2715 -115 2725 -100
rect 2745 -115 2755 -95
rect 2715 -125 2755 -115
rect -625 -305 -585 -295
rect -625 -325 -615 -305
rect -595 -325 -585 -305
rect -625 -330 -585 -325
rect 2275 -305 2315 -295
rect 2275 -325 2285 -305
rect 2305 -325 2315 -305
rect 2275 -330 2315 -325
rect -985 -355 -925 -340
rect -885 -345 -525 -330
rect -885 -355 -825 -345
rect -785 -355 -725 -345
rect -685 -355 -625 -345
rect -585 -355 -525 -345
rect -485 -355 -425 -340
rect 770 -355 800 -345
rect 770 -375 775 -355
rect 795 -375 800 -355
rect 770 -380 800 -375
rect 1336 -355 1366 -345
rect 2115 -355 2175 -340
rect 2215 -345 2575 -330
rect 2215 -355 2275 -345
rect 2315 -355 2375 -345
rect 2415 -355 2475 -345
rect 2515 -355 2575 -345
rect 2615 -355 2675 -340
rect 1336 -375 1341 -355
rect 1361 -370 1366 -355
rect 1361 -375 1370 -370
rect 200 -405 215 -390
rect 255 -395 1315 -380
rect 1336 -385 1370 -375
rect 255 -405 270 -395
rect 310 -405 325 -395
rect 365 -405 380 -395
rect 420 -405 435 -395
rect 475 -405 490 -395
rect 530 -405 545 -395
rect 585 -405 600 -395
rect 640 -405 655 -395
rect 695 -405 710 -395
rect 750 -405 765 -395
rect 805 -405 820 -395
rect 860 -405 875 -395
rect 915 -405 930 -395
rect 970 -405 985 -395
rect 1025 -405 1040 -395
rect 1080 -405 1095 -395
rect 1135 -405 1150 -395
rect 1190 -405 1205 -395
rect 1245 -405 1260 -395
rect 1300 -405 1315 -395
rect 1355 -405 1370 -385
rect 1410 -405 1425 -390
rect 200 -670 215 -655
rect 255 -670 270 -655
rect 310 -670 325 -655
rect 365 -670 380 -655
rect 420 -670 435 -655
rect 475 -670 490 -655
rect 530 -670 545 -655
rect 585 -670 600 -655
rect 640 -670 655 -655
rect 695 -670 710 -655
rect 750 -670 765 -655
rect 805 -670 820 -655
rect 860 -670 875 -655
rect 915 -670 930 -655
rect 970 -670 985 -655
rect 1025 -670 1040 -655
rect 1080 -670 1095 -655
rect 1135 -670 1150 -655
rect 1190 -670 1205 -655
rect 1245 -670 1260 -655
rect 1300 -670 1315 -655
rect 1355 -670 1370 -655
rect 1410 -670 1425 -655
rect 150 -680 215 -670
rect 150 -700 160 -680
rect 180 -685 215 -680
rect 1410 -680 1465 -670
rect 1410 -685 1435 -680
rect 180 -700 190 -685
rect 150 -710 190 -700
rect 1425 -700 1435 -685
rect 1455 -700 1465 -680
rect 1425 -710 1465 -700
rect 710 -775 750 -765
rect 710 -795 720 -775
rect 740 -795 750 -775
rect 710 -805 750 -795
rect 825 -775 865 -765
rect 825 -795 835 -775
rect 855 -795 865 -775
rect 825 -805 865 -795
rect 950 -775 990 -765
rect 950 -795 960 -775
rect 980 -795 990 -775
rect 950 -805 990 -795
rect 705 -820 995 -805
rect 705 -935 995 -920
rect -985 -1070 -925 -1055
rect -885 -1070 -825 -1055
rect -785 -1070 -725 -1055
rect -685 -1070 -625 -1055
rect -585 -1070 -525 -1055
rect -485 -1070 -425 -1055
rect 2115 -1070 2175 -1055
rect 2215 -1070 2275 -1055
rect 2315 -1070 2375 -1055
rect 2415 -1070 2475 -1055
rect 2515 -1070 2575 -1055
rect 2615 -1070 2675 -1055
rect -1025 -1080 -925 -1070
rect -1025 -1100 -1015 -1080
rect -995 -1085 -925 -1080
rect -485 -1080 -385 -1070
rect -485 -1085 -415 -1080
rect -995 -1100 -985 -1085
rect -1025 -1110 -985 -1100
rect -425 -1100 -415 -1085
rect -395 -1100 -385 -1080
rect -425 -1110 -385 -1100
rect 2075 -1080 2175 -1070
rect 2075 -1100 2085 -1080
rect 2105 -1085 2175 -1080
rect 2615 -1080 2715 -1070
rect 2615 -1085 2685 -1080
rect 2105 -1100 2115 -1085
rect 2075 -1110 2115 -1100
rect 2675 -1100 2685 -1085
rect 2705 -1100 2715 -1080
rect 2675 -1110 2715 -1100
<< polycont >>
rect 40 2700 60 2720
rect 220 2700 240 2720
rect 980 2700 1000 2720
rect 1160 2700 1180 2720
rect 1448 2700 1468 2720
rect 1628 2700 1648 2720
rect 510 2530 530 2550
rect 690 2530 710 2550
rect 144 2280 164 2300
rect 614 2280 634 2300
rect 1056 2280 1076 2300
rect 1524 2280 1544 2300
rect -1075 2125 -1055 2145
rect -355 2125 -335 2145
rect -30 2125 -10 2145
rect 690 2125 710 2145
rect 980 2125 1000 2145
rect 1700 2125 1720 2145
rect 2025 2125 2045 2145
rect 2745 2125 2765 2145
rect -715 1700 -695 1720
rect 330 1700 350 1720
rect 1340 1700 1360 1720
rect 2385 1700 2405 1720
rect 230 1555 250 1575
rect 1440 1555 1460 1575
rect -1045 1460 -1025 1480
rect -385 1460 -365 1480
rect 2055 1460 2075 1480
rect 2715 1460 2735 1480
rect 890 1430 910 1450
rect 76 1230 96 1250
rect 280 1230 300 1250
rect 500 1230 520 1250
rect 1076 1230 1096 1250
rect 1280 1230 1300 1250
rect 1500 1230 1520 1250
rect 0 1110 20 1130
rect 209 1111 229 1131
rect 429 1111 449 1131
rect 571 1111 591 1131
rect 670 1110 690 1130
rect 1000 1110 1020 1130
rect 1209 1111 1229 1131
rect 1429 1111 1449 1131
rect 1571 1111 1591 1131
rect 1670 1110 1690 1130
rect 670 905 690 925
rect 890 905 910 925
rect -715 780 -695 800
rect 505 785 525 805
rect 1165 785 1185 805
rect 2385 780 2405 800
rect -1055 645 -1035 665
rect -375 645 -355 665
rect 315 635 335 655
rect 1355 635 1375 655
rect 2045 645 2065 665
rect 2725 645 2745 665
rect -15 410 5 430
rect 645 410 665 430
rect 1025 410 1045 430
rect 1685 410 1705 430
rect -660 370 -640 390
rect 2330 370 2350 390
rect -660 260 -640 280
rect 2330 260 2350 280
rect 315 155 335 175
rect 800 155 820 175
rect 853 155 873 175
rect 1355 155 1375 175
rect -15 -65 5 -45
rect 685 -65 705 -45
rect 985 -65 1005 -45
rect 1685 -65 1705 -45
rect -1055 -115 -1035 -95
rect -375 -115 -355 -95
rect 2045 -115 2065 -95
rect 2725 -115 2745 -95
rect -615 -325 -595 -305
rect 2285 -325 2305 -305
rect 775 -375 795 -355
rect 1341 -375 1361 -355
rect 160 -700 180 -680
rect 1435 -700 1455 -680
rect 720 -795 740 -775
rect 835 -795 855 -775
rect 960 -795 980 -775
rect -1015 -1100 -995 -1080
rect -415 -1100 -395 -1080
rect 2085 -1100 2105 -1080
rect 2685 -1100 2705 -1080
<< xpolycontact >>
rect -1501 1170 -1360 1390
rect -1501 825 -1360 1045
rect 3050 1170 3191 1390
rect 3050 825 3191 1045
rect -1410 297 -1375 517
rect -1410 -85 -1375 138
rect -1350 297 -1315 517
rect -1350 -85 -1315 138
rect -1290 297 -1255 517
rect -1290 -85 -1255 138
rect -1230 297 -1195 517
rect 2885 297 2920 517
rect -1230 -85 -1195 138
rect 2885 -85 2920 138
rect 2945 297 2980 517
rect 2945 -85 2980 138
rect 3005 297 3040 517
rect 3005 -85 3040 138
rect 3065 297 3100 517
rect 3065 -85 3100 138
rect -1210 -638 -1175 -415
rect -1210 -1105 -1175 -885
rect -1150 -638 -1115 -415
rect -1150 -1105 -1115 -885
rect 2805 -638 2840 -415
rect 2805 -1105 2840 -885
rect 2865 -638 2900 -415
rect 2865 -1105 2900 -885
<< ppolyres >>
rect -1501 1045 -1360 1170
rect 3050 1045 3191 1170
<< xpolyres >>
rect -1410 138 -1375 297
rect -1350 138 -1315 297
rect -1290 138 -1255 297
rect -1230 138 -1195 297
rect 2885 138 2920 297
rect 2945 138 2980 297
rect 3005 138 3040 297
rect 3065 138 3100 297
rect -1210 -885 -1175 -638
rect -1150 -885 -1115 -638
rect 2805 -885 2840 -638
rect 2865 -885 2900 -638
<< locali >>
rect 30 2720 70 2730
rect 30 2700 40 2720
rect 60 2700 70 2720
rect 30 2690 70 2700
rect 150 2720 190 2730
rect 150 2700 160 2720
rect 180 2700 190 2720
rect 150 2690 190 2700
rect 210 2720 250 2730
rect 210 2700 220 2720
rect 240 2700 250 2720
rect 210 2690 250 2700
rect 970 2720 1010 2730
rect 970 2700 980 2720
rect 1000 2700 1010 2720
rect 970 2690 1010 2700
rect 1035 2720 1065 2730
rect 1035 2700 1040 2720
rect 1060 2700 1065 2720
rect 1035 2690 1065 2700
rect 1090 2720 1130 2730
rect 1090 2700 1100 2720
rect 1120 2700 1130 2720
rect 1090 2690 1130 2700
rect 1150 2720 1190 2730
rect 1150 2700 1160 2720
rect 1180 2700 1190 2720
rect 1150 2690 1190 2700
rect 1438 2720 1478 2730
rect 1438 2700 1448 2720
rect 1468 2700 1478 2720
rect 1438 2690 1478 2700
rect 1498 2720 1538 2730
rect 1498 2700 1508 2720
rect 1528 2700 1538 2720
rect 1498 2690 1538 2700
rect 1618 2720 1658 2730
rect 1618 2700 1628 2720
rect 1648 2700 1658 2720
rect 1618 2690 1658 2700
rect 40 2670 60 2690
rect 160 2670 180 2690
rect 220 2670 240 2690
rect 980 2670 1000 2690
rect 1040 2670 1060 2690
rect 1100 2670 1120 2690
rect 1160 2670 1180 2690
rect 1448 2670 1468 2690
rect 1508 2670 1528 2690
rect 1628 2670 1648 2690
rect -5 2660 65 2670
rect -5 2640 0 2660
rect 20 2640 40 2660
rect 60 2640 65 2660
rect -5 2610 65 2640
rect -5 2590 0 2610
rect 20 2590 40 2610
rect 60 2590 65 2610
rect -5 2560 65 2590
rect -5 2540 0 2560
rect 20 2540 40 2560
rect 60 2540 65 2560
rect -5 2510 65 2540
rect -5 2490 0 2510
rect 20 2490 40 2510
rect 60 2490 65 2510
rect -5 2460 65 2490
rect -5 2440 0 2460
rect 20 2440 40 2460
rect 60 2440 65 2460
rect -5 2410 65 2440
rect -5 2390 0 2410
rect 20 2390 40 2410
rect 60 2390 65 2410
rect -5 2360 65 2390
rect -5 2340 0 2360
rect 20 2340 40 2360
rect 60 2340 65 2360
rect -5 2330 65 2340
rect 95 2660 125 2670
rect 95 2640 100 2660
rect 120 2640 125 2660
rect 95 2610 125 2640
rect 95 2590 100 2610
rect 120 2590 125 2610
rect 95 2560 125 2590
rect 95 2540 100 2560
rect 120 2540 125 2560
rect 95 2510 125 2540
rect 95 2490 100 2510
rect 120 2490 125 2510
rect 95 2460 125 2490
rect 95 2440 100 2460
rect 120 2440 125 2460
rect 95 2410 125 2440
rect 95 2390 100 2410
rect 120 2390 125 2410
rect 95 2360 125 2390
rect 95 2340 100 2360
rect 120 2340 125 2360
rect 95 2330 125 2340
rect 155 2660 185 2670
rect 155 2640 160 2660
rect 180 2640 185 2660
rect 155 2610 185 2640
rect 155 2590 160 2610
rect 180 2590 185 2610
rect 155 2560 185 2590
rect 155 2540 160 2560
rect 180 2540 185 2560
rect 155 2510 185 2540
rect 155 2490 160 2510
rect 180 2490 185 2510
rect 155 2460 185 2490
rect 155 2440 160 2460
rect 180 2440 185 2460
rect 155 2410 185 2440
rect 155 2390 160 2410
rect 180 2390 185 2410
rect 155 2360 185 2390
rect 155 2340 160 2360
rect 180 2340 185 2360
rect 155 2330 185 2340
rect 215 2660 285 2670
rect 215 2640 220 2660
rect 240 2640 260 2660
rect 280 2640 285 2660
rect 215 2610 285 2640
rect 215 2590 220 2610
rect 240 2590 260 2610
rect 280 2590 285 2610
rect 215 2560 285 2590
rect 935 2660 1005 2670
rect 935 2640 940 2660
rect 960 2640 980 2660
rect 1000 2640 1005 2660
rect 935 2610 1005 2640
rect 935 2590 940 2610
rect 960 2590 980 2610
rect 1000 2590 1005 2610
rect 935 2560 1005 2590
rect 215 2540 220 2560
rect 240 2540 260 2560
rect 280 2540 285 2560
rect 215 2510 285 2540
rect 500 2550 540 2560
rect 500 2530 510 2550
rect 530 2530 540 2550
rect 500 2520 540 2530
rect 560 2550 600 2560
rect 560 2530 570 2550
rect 590 2530 600 2550
rect 560 2520 600 2530
rect 625 2550 655 2560
rect 625 2530 630 2550
rect 650 2530 655 2550
rect 625 2520 655 2530
rect 680 2550 720 2560
rect 680 2530 690 2550
rect 710 2530 720 2550
rect 680 2520 720 2530
rect 935 2540 940 2560
rect 960 2540 980 2560
rect 1000 2540 1005 2560
rect 215 2490 220 2510
rect 240 2490 260 2510
rect 280 2490 285 2510
rect 510 2500 530 2520
rect 570 2500 590 2520
rect 630 2500 650 2520
rect 690 2500 710 2520
rect 935 2510 1005 2540
rect 215 2460 285 2490
rect 215 2440 220 2460
rect 240 2440 260 2460
rect 280 2440 285 2460
rect 215 2410 285 2440
rect 215 2390 220 2410
rect 240 2390 260 2410
rect 280 2390 285 2410
rect 215 2360 285 2390
rect 215 2340 220 2360
rect 240 2340 260 2360
rect 280 2340 285 2360
rect 215 2330 285 2340
rect 465 2360 535 2500
rect 465 2340 470 2360
rect 490 2340 510 2360
rect 530 2340 535 2360
rect 465 2330 535 2340
rect 565 2360 595 2500
rect 565 2340 570 2360
rect 590 2340 595 2360
rect 565 2330 595 2340
rect 625 2360 655 2500
rect 625 2340 630 2360
rect 650 2340 655 2360
rect 625 2330 655 2340
rect 685 2360 755 2500
rect 685 2340 690 2360
rect 710 2340 730 2360
rect 750 2340 755 2360
rect 685 2330 755 2340
rect 935 2490 940 2510
rect 960 2490 980 2510
rect 1000 2490 1005 2510
rect 935 2460 1005 2490
rect 935 2440 940 2460
rect 960 2440 980 2460
rect 1000 2440 1005 2460
rect 935 2410 1005 2440
rect 935 2390 940 2410
rect 960 2390 980 2410
rect 1000 2390 1005 2410
rect 935 2360 1005 2390
rect 935 2340 940 2360
rect 960 2340 980 2360
rect 1000 2340 1005 2360
rect 935 2330 1005 2340
rect 1035 2660 1065 2670
rect 1035 2640 1040 2660
rect 1060 2640 1065 2660
rect 1035 2610 1065 2640
rect 1035 2590 1040 2610
rect 1060 2590 1065 2610
rect 1035 2560 1065 2590
rect 1035 2540 1040 2560
rect 1060 2540 1065 2560
rect 1035 2510 1065 2540
rect 1035 2490 1040 2510
rect 1060 2490 1065 2510
rect 1035 2460 1065 2490
rect 1035 2440 1040 2460
rect 1060 2440 1065 2460
rect 1035 2410 1065 2440
rect 1035 2390 1040 2410
rect 1060 2390 1065 2410
rect 1035 2360 1065 2390
rect 1035 2340 1040 2360
rect 1060 2340 1065 2360
rect 1035 2330 1065 2340
rect 1095 2660 1125 2670
rect 1095 2640 1100 2660
rect 1120 2640 1125 2660
rect 1095 2610 1125 2640
rect 1095 2590 1100 2610
rect 1120 2590 1125 2610
rect 1095 2560 1125 2590
rect 1095 2540 1100 2560
rect 1120 2540 1125 2560
rect 1095 2510 1125 2540
rect 1095 2490 1100 2510
rect 1120 2490 1125 2510
rect 1095 2460 1125 2490
rect 1095 2440 1100 2460
rect 1120 2440 1125 2460
rect 1095 2410 1125 2440
rect 1095 2390 1100 2410
rect 1120 2390 1125 2410
rect 1095 2360 1125 2390
rect 1095 2340 1100 2360
rect 1120 2340 1125 2360
rect 1095 2330 1125 2340
rect 1155 2660 1225 2670
rect 1155 2640 1160 2660
rect 1180 2640 1200 2660
rect 1220 2640 1225 2660
rect 1155 2610 1225 2640
rect 1155 2590 1160 2610
rect 1180 2590 1200 2610
rect 1220 2590 1225 2610
rect 1155 2560 1225 2590
rect 1155 2540 1160 2560
rect 1180 2540 1200 2560
rect 1220 2540 1225 2560
rect 1155 2510 1225 2540
rect 1155 2490 1160 2510
rect 1180 2490 1200 2510
rect 1220 2490 1225 2510
rect 1155 2460 1225 2490
rect 1155 2440 1160 2460
rect 1180 2440 1200 2460
rect 1220 2440 1225 2460
rect 1155 2410 1225 2440
rect 1155 2390 1160 2410
rect 1180 2390 1200 2410
rect 1220 2390 1225 2410
rect 1155 2360 1225 2390
rect 1155 2340 1160 2360
rect 1180 2340 1200 2360
rect 1220 2340 1225 2360
rect 1155 2330 1225 2340
rect 1403 2660 1473 2670
rect 1403 2640 1408 2660
rect 1428 2640 1448 2660
rect 1468 2640 1473 2660
rect 1403 2610 1473 2640
rect 1403 2590 1408 2610
rect 1428 2590 1448 2610
rect 1468 2590 1473 2610
rect 1403 2560 1473 2590
rect 1403 2540 1408 2560
rect 1428 2540 1448 2560
rect 1468 2540 1473 2560
rect 1403 2510 1473 2540
rect 1403 2490 1408 2510
rect 1428 2490 1448 2510
rect 1468 2490 1473 2510
rect 1403 2460 1473 2490
rect 1403 2440 1408 2460
rect 1428 2440 1448 2460
rect 1468 2440 1473 2460
rect 1403 2410 1473 2440
rect 1403 2390 1408 2410
rect 1428 2390 1448 2410
rect 1468 2390 1473 2410
rect 1403 2360 1473 2390
rect 1403 2340 1408 2360
rect 1428 2340 1448 2360
rect 1468 2340 1473 2360
rect 1403 2330 1473 2340
rect 1503 2660 1533 2670
rect 1503 2640 1508 2660
rect 1528 2640 1533 2660
rect 1503 2610 1533 2640
rect 1503 2590 1508 2610
rect 1528 2590 1533 2610
rect 1503 2560 1533 2590
rect 1503 2540 1508 2560
rect 1528 2540 1533 2560
rect 1503 2510 1533 2540
rect 1503 2490 1508 2510
rect 1528 2490 1533 2510
rect 1503 2460 1533 2490
rect 1503 2440 1508 2460
rect 1528 2440 1533 2460
rect 1503 2410 1533 2440
rect 1503 2390 1508 2410
rect 1528 2390 1533 2410
rect 1503 2360 1533 2390
rect 1503 2340 1508 2360
rect 1528 2340 1533 2360
rect 1503 2330 1533 2340
rect 1563 2660 1593 2670
rect 1563 2640 1568 2660
rect 1588 2640 1593 2660
rect 1563 2610 1593 2640
rect 1563 2590 1568 2610
rect 1588 2590 1593 2610
rect 1563 2560 1593 2590
rect 1563 2540 1568 2560
rect 1588 2540 1593 2560
rect 1563 2510 1593 2540
rect 1563 2490 1568 2510
rect 1588 2490 1593 2510
rect 1563 2460 1593 2490
rect 1563 2440 1568 2460
rect 1588 2440 1593 2460
rect 1563 2410 1593 2440
rect 1563 2390 1568 2410
rect 1588 2390 1593 2410
rect 1563 2360 1593 2390
rect 1563 2340 1568 2360
rect 1588 2340 1593 2360
rect 1563 2330 1593 2340
rect 1623 2660 1693 2670
rect 1623 2640 1628 2660
rect 1648 2640 1668 2660
rect 1688 2640 1693 2660
rect 1623 2610 1693 2640
rect 1623 2590 1628 2610
rect 1648 2590 1668 2610
rect 1688 2590 1693 2610
rect 1623 2560 1693 2590
rect 1623 2540 1628 2560
rect 1648 2540 1668 2560
rect 1688 2540 1693 2560
rect 1623 2510 1693 2540
rect 1623 2490 1628 2510
rect 1648 2490 1668 2510
rect 1688 2490 1693 2510
rect 1623 2460 1693 2490
rect 1623 2440 1628 2460
rect 1648 2440 1668 2460
rect 1688 2440 1693 2460
rect 1623 2410 1693 2440
rect 1623 2390 1628 2410
rect 1648 2390 1668 2410
rect 1688 2390 1693 2410
rect 1623 2360 1693 2390
rect 1623 2340 1628 2360
rect 1648 2340 1668 2360
rect 1688 2340 1693 2360
rect 1623 2330 1693 2340
rect 95 2310 115 2330
rect 1573 2310 1593 2330
rect 75 2300 115 2310
rect 75 2280 85 2300
rect 105 2280 115 2300
rect 75 2270 115 2280
rect 139 2300 169 2310
rect 139 2280 144 2300
rect 164 2280 169 2300
rect 139 2270 169 2280
rect 609 2300 639 2310
rect 609 2280 614 2300
rect 634 2280 639 2300
rect 609 2270 639 2280
rect 1051 2300 1081 2310
rect 1051 2280 1056 2300
rect 1076 2280 1081 2300
rect 1051 2270 1081 2280
rect 1519 2300 1549 2310
rect 1519 2280 1524 2300
rect 1544 2280 1549 2300
rect 1519 2270 1549 2280
rect 1573 2300 1613 2310
rect 1573 2280 1583 2300
rect 1603 2280 1613 2300
rect 1573 2270 1613 2280
rect -1085 2145 -1045 2155
rect -1085 2125 -1075 2145
rect -1055 2125 -1045 2145
rect -1085 2115 -1045 2125
rect -965 2145 -925 2155
rect -965 2125 -955 2145
rect -935 2125 -925 2145
rect -965 2115 -925 2125
rect -845 2145 -805 2155
rect -845 2125 -835 2145
rect -815 2125 -805 2145
rect -845 2115 -805 2125
rect -725 2145 -685 2155
rect -725 2125 -715 2145
rect -695 2125 -685 2145
rect -725 2115 -685 2125
rect -605 2145 -565 2155
rect -605 2125 -595 2145
rect -575 2125 -565 2145
rect -605 2115 -565 2125
rect -485 2145 -445 2155
rect -485 2125 -475 2145
rect -455 2125 -445 2145
rect -485 2115 -445 2125
rect -365 2145 -325 2155
rect -365 2125 -355 2145
rect -335 2125 -325 2145
rect -365 2115 -325 2125
rect -40 2145 0 2155
rect -40 2125 -30 2145
rect -10 2125 0 2145
rect -40 2115 0 2125
rect 80 2145 120 2155
rect 80 2125 90 2145
rect 110 2125 120 2145
rect 80 2115 120 2125
rect 200 2145 240 2155
rect 200 2125 210 2145
rect 230 2125 240 2145
rect 200 2115 240 2125
rect 320 2145 360 2155
rect 320 2125 330 2145
rect 350 2125 360 2145
rect 320 2115 360 2125
rect 440 2145 480 2155
rect 440 2125 450 2145
rect 470 2125 480 2145
rect 440 2115 480 2125
rect 560 2145 600 2155
rect 560 2125 570 2145
rect 590 2125 600 2145
rect 560 2115 600 2125
rect 680 2145 720 2155
rect 680 2125 690 2145
rect 710 2125 720 2145
rect 680 2115 720 2125
rect 970 2145 1010 2155
rect 970 2125 980 2145
rect 1000 2125 1010 2145
rect 970 2115 1010 2125
rect 1090 2145 1130 2155
rect 1090 2125 1100 2145
rect 1120 2125 1130 2145
rect 1090 2115 1130 2125
rect 1210 2145 1250 2155
rect 1210 2125 1220 2145
rect 1240 2125 1250 2145
rect 1210 2115 1250 2125
rect 1330 2145 1370 2155
rect 1330 2125 1340 2145
rect 1360 2125 1370 2145
rect 1330 2115 1370 2125
rect 1450 2145 1490 2155
rect 1450 2125 1460 2145
rect 1480 2125 1490 2145
rect 1450 2115 1490 2125
rect 1570 2145 1610 2155
rect 1570 2125 1580 2145
rect 1600 2125 1610 2145
rect 1570 2115 1610 2125
rect 1690 2145 1730 2155
rect 1690 2125 1700 2145
rect 1720 2125 1730 2145
rect 1690 2115 1730 2125
rect 2015 2145 2055 2155
rect 2015 2125 2025 2145
rect 2045 2125 2055 2145
rect 2015 2115 2055 2125
rect 2135 2145 2175 2155
rect 2135 2125 2145 2145
rect 2165 2125 2175 2145
rect 2135 2115 2175 2125
rect 2255 2145 2295 2155
rect 2255 2125 2265 2145
rect 2285 2125 2295 2145
rect 2255 2115 2295 2125
rect 2375 2145 2415 2155
rect 2375 2125 2385 2145
rect 2405 2125 2415 2145
rect 2375 2115 2415 2125
rect 2495 2145 2535 2155
rect 2495 2125 2505 2145
rect 2525 2125 2535 2145
rect 2495 2115 2535 2125
rect 2615 2145 2655 2155
rect 2615 2125 2625 2145
rect 2645 2125 2655 2145
rect 2615 2115 2655 2125
rect 2735 2145 2775 2155
rect 2735 2125 2745 2145
rect 2765 2125 2775 2145
rect 2735 2115 2775 2125
rect -1075 2095 -1055 2115
rect -955 2095 -935 2115
rect -835 2095 -815 2115
rect -715 2095 -695 2115
rect -595 2095 -575 2115
rect -475 2095 -455 2115
rect -355 2095 -335 2115
rect -30 2095 -10 2115
rect 90 2095 110 2115
rect 210 2095 230 2115
rect 330 2095 350 2115
rect 450 2095 470 2115
rect 570 2095 590 2115
rect 690 2095 710 2115
rect 980 2095 1000 2115
rect 1100 2095 1120 2115
rect 1220 2095 1240 2115
rect 1340 2095 1360 2115
rect 1460 2095 1480 2115
rect 1580 2095 1600 2115
rect 1700 2095 1720 2115
rect 2025 2095 2045 2115
rect 2145 2095 2165 2115
rect 2265 2095 2285 2115
rect 2385 2095 2405 2115
rect 2505 2095 2525 2115
rect 2625 2095 2645 2115
rect 2745 2095 2765 2115
rect -1120 2085 -1050 2095
rect -1120 2065 -1115 2085
rect -1095 2065 -1075 2085
rect -1055 2065 -1050 2085
rect -1120 2035 -1050 2065
rect -1120 2015 -1115 2035
rect -1095 2015 -1075 2035
rect -1055 2015 -1050 2035
rect -1120 1985 -1050 2015
rect -1120 1965 -1115 1985
rect -1095 1965 -1075 1985
rect -1055 1965 -1050 1985
rect -1120 1935 -1050 1965
rect -1120 1915 -1115 1935
rect -1095 1915 -1075 1935
rect -1055 1915 -1050 1935
rect -1120 1885 -1050 1915
rect -1120 1865 -1115 1885
rect -1095 1865 -1075 1885
rect -1055 1865 -1050 1885
rect -1120 1835 -1050 1865
rect -1120 1815 -1115 1835
rect -1095 1815 -1075 1835
rect -1055 1815 -1050 1835
rect -1120 1785 -1050 1815
rect -1120 1765 -1115 1785
rect -1095 1765 -1075 1785
rect -1055 1765 -1050 1785
rect -1120 1755 -1050 1765
rect -1020 2085 -990 2095
rect -1020 2065 -1015 2085
rect -995 2065 -990 2085
rect -1020 2035 -990 2065
rect -1020 2015 -1015 2035
rect -995 2015 -990 2035
rect -1020 1985 -990 2015
rect -1020 1965 -1015 1985
rect -995 1965 -990 1985
rect -1020 1935 -990 1965
rect -1020 1915 -1015 1935
rect -995 1915 -990 1935
rect -1020 1885 -990 1915
rect -1020 1865 -1015 1885
rect -995 1865 -990 1885
rect -1020 1835 -990 1865
rect -1020 1815 -1015 1835
rect -995 1815 -990 1835
rect -1020 1785 -990 1815
rect -1020 1765 -1015 1785
rect -995 1765 -990 1785
rect -1020 1755 -990 1765
rect -960 2085 -930 2095
rect -960 2065 -955 2085
rect -935 2065 -930 2085
rect -960 2035 -930 2065
rect -960 2015 -955 2035
rect -935 2015 -930 2035
rect -960 1985 -930 2015
rect -960 1965 -955 1985
rect -935 1965 -930 1985
rect -960 1935 -930 1965
rect -960 1915 -955 1935
rect -935 1915 -930 1935
rect -960 1885 -930 1915
rect -960 1865 -955 1885
rect -935 1865 -930 1885
rect -960 1835 -930 1865
rect -960 1815 -955 1835
rect -935 1815 -930 1835
rect -960 1785 -930 1815
rect -960 1765 -955 1785
rect -935 1765 -930 1785
rect -960 1755 -930 1765
rect -900 2085 -870 2095
rect -900 2065 -895 2085
rect -875 2065 -870 2085
rect -900 2035 -870 2065
rect -900 2015 -895 2035
rect -875 2015 -870 2035
rect -900 1985 -870 2015
rect -900 1965 -895 1985
rect -875 1965 -870 1985
rect -900 1935 -870 1965
rect -900 1915 -895 1935
rect -875 1915 -870 1935
rect -900 1885 -870 1915
rect -900 1865 -895 1885
rect -875 1865 -870 1885
rect -900 1835 -870 1865
rect -900 1815 -895 1835
rect -875 1815 -870 1835
rect -900 1785 -870 1815
rect -900 1765 -895 1785
rect -875 1765 -870 1785
rect -900 1755 -870 1765
rect -840 2085 -810 2095
rect -840 2065 -835 2085
rect -815 2065 -810 2085
rect -840 2035 -810 2065
rect -840 2015 -835 2035
rect -815 2015 -810 2035
rect -840 1985 -810 2015
rect -840 1965 -835 1985
rect -815 1965 -810 1985
rect -840 1935 -810 1965
rect -840 1915 -835 1935
rect -815 1915 -810 1935
rect -840 1885 -810 1915
rect -840 1865 -835 1885
rect -815 1865 -810 1885
rect -840 1835 -810 1865
rect -840 1815 -835 1835
rect -815 1815 -810 1835
rect -840 1785 -810 1815
rect -840 1765 -835 1785
rect -815 1765 -810 1785
rect -840 1755 -810 1765
rect -780 2085 -750 2095
rect -780 2065 -775 2085
rect -755 2065 -750 2085
rect -780 2035 -750 2065
rect -780 2015 -775 2035
rect -755 2015 -750 2035
rect -780 1985 -750 2015
rect -780 1965 -775 1985
rect -755 1965 -750 1985
rect -780 1935 -750 1965
rect -780 1915 -775 1935
rect -755 1915 -750 1935
rect -780 1885 -750 1915
rect -780 1865 -775 1885
rect -755 1865 -750 1885
rect -780 1835 -750 1865
rect -780 1815 -775 1835
rect -755 1815 -750 1835
rect -780 1785 -750 1815
rect -780 1765 -775 1785
rect -755 1765 -750 1785
rect -780 1755 -750 1765
rect -720 2085 -690 2095
rect -720 2065 -715 2085
rect -695 2065 -690 2085
rect -720 2035 -690 2065
rect -720 2015 -715 2035
rect -695 2015 -690 2035
rect -720 1985 -690 2015
rect -720 1965 -715 1985
rect -695 1965 -690 1985
rect -720 1935 -690 1965
rect -720 1915 -715 1935
rect -695 1915 -690 1935
rect -720 1885 -690 1915
rect -720 1865 -715 1885
rect -695 1865 -690 1885
rect -720 1835 -690 1865
rect -720 1815 -715 1835
rect -695 1815 -690 1835
rect -720 1785 -690 1815
rect -720 1765 -715 1785
rect -695 1765 -690 1785
rect -720 1755 -690 1765
rect -660 2085 -630 2095
rect -660 2065 -655 2085
rect -635 2065 -630 2085
rect -660 2035 -630 2065
rect -660 2015 -655 2035
rect -635 2015 -630 2035
rect -660 1985 -630 2015
rect -660 1965 -655 1985
rect -635 1965 -630 1985
rect -660 1935 -630 1965
rect -660 1915 -655 1935
rect -635 1915 -630 1935
rect -660 1885 -630 1915
rect -660 1865 -655 1885
rect -635 1865 -630 1885
rect -660 1835 -630 1865
rect -660 1815 -655 1835
rect -635 1815 -630 1835
rect -660 1785 -630 1815
rect -660 1765 -655 1785
rect -635 1765 -630 1785
rect -660 1755 -630 1765
rect -600 2085 -570 2095
rect -600 2065 -595 2085
rect -575 2065 -570 2085
rect -600 2035 -570 2065
rect -600 2015 -595 2035
rect -575 2015 -570 2035
rect -600 1985 -570 2015
rect -600 1965 -595 1985
rect -575 1965 -570 1985
rect -600 1935 -570 1965
rect -600 1915 -595 1935
rect -575 1915 -570 1935
rect -600 1885 -570 1915
rect -600 1865 -595 1885
rect -575 1865 -570 1885
rect -600 1835 -570 1865
rect -600 1815 -595 1835
rect -575 1815 -570 1835
rect -600 1785 -570 1815
rect -600 1765 -595 1785
rect -575 1765 -570 1785
rect -600 1755 -570 1765
rect -540 2085 -510 2095
rect -540 2065 -535 2085
rect -515 2065 -510 2085
rect -540 2035 -510 2065
rect -540 2015 -535 2035
rect -515 2015 -510 2035
rect -540 1985 -510 2015
rect -540 1965 -535 1985
rect -515 1965 -510 1985
rect -540 1935 -510 1965
rect -540 1915 -535 1935
rect -515 1915 -510 1935
rect -540 1885 -510 1915
rect -540 1865 -535 1885
rect -515 1865 -510 1885
rect -540 1835 -510 1865
rect -540 1815 -535 1835
rect -515 1815 -510 1835
rect -540 1785 -510 1815
rect -540 1765 -535 1785
rect -515 1765 -510 1785
rect -540 1755 -510 1765
rect -480 2085 -450 2095
rect -480 2065 -475 2085
rect -455 2065 -450 2085
rect -480 2035 -450 2065
rect -480 2015 -475 2035
rect -455 2015 -450 2035
rect -480 1985 -450 2015
rect -480 1965 -475 1985
rect -455 1965 -450 1985
rect -480 1935 -450 1965
rect -480 1915 -475 1935
rect -455 1915 -450 1935
rect -480 1885 -450 1915
rect -480 1865 -475 1885
rect -455 1865 -450 1885
rect -480 1835 -450 1865
rect -480 1815 -475 1835
rect -455 1815 -450 1835
rect -480 1785 -450 1815
rect -480 1765 -475 1785
rect -455 1765 -450 1785
rect -480 1755 -450 1765
rect -420 2085 -390 2095
rect -420 2065 -415 2085
rect -395 2065 -390 2085
rect -420 2035 -390 2065
rect -420 2015 -415 2035
rect -395 2015 -390 2035
rect -420 1985 -390 2015
rect -420 1965 -415 1985
rect -395 1965 -390 1985
rect -420 1935 -390 1965
rect -420 1915 -415 1935
rect -395 1915 -390 1935
rect -420 1885 -390 1915
rect -420 1865 -415 1885
rect -395 1865 -390 1885
rect -420 1835 -390 1865
rect -420 1815 -415 1835
rect -395 1815 -390 1835
rect -420 1785 -390 1815
rect -420 1765 -415 1785
rect -395 1765 -390 1785
rect -420 1755 -390 1765
rect -360 2085 -290 2095
rect -360 2065 -355 2085
rect -335 2065 -315 2085
rect -295 2065 -290 2085
rect -360 2035 -290 2065
rect -360 2015 -355 2035
rect -335 2015 -315 2035
rect -295 2015 -290 2035
rect -360 1985 -290 2015
rect -360 1965 -355 1985
rect -335 1965 -315 1985
rect -295 1965 -290 1985
rect -360 1935 -290 1965
rect -360 1915 -355 1935
rect -335 1915 -315 1935
rect -295 1915 -290 1935
rect -360 1885 -290 1915
rect -360 1865 -355 1885
rect -335 1865 -315 1885
rect -295 1865 -290 1885
rect -360 1835 -290 1865
rect -360 1815 -355 1835
rect -335 1815 -315 1835
rect -295 1815 -290 1835
rect -360 1785 -290 1815
rect -360 1765 -355 1785
rect -335 1765 -315 1785
rect -295 1765 -290 1785
rect -360 1755 -290 1765
rect -75 2085 -5 2095
rect -75 2065 -70 2085
rect -50 2065 -30 2085
rect -10 2065 -5 2085
rect -75 2035 -5 2065
rect -75 2015 -70 2035
rect -50 2015 -30 2035
rect -10 2015 -5 2035
rect -75 1985 -5 2015
rect -75 1965 -70 1985
rect -50 1965 -30 1985
rect -10 1965 -5 1985
rect -75 1935 -5 1965
rect -75 1915 -70 1935
rect -50 1915 -30 1935
rect -10 1915 -5 1935
rect -75 1885 -5 1915
rect -75 1865 -70 1885
rect -50 1865 -30 1885
rect -10 1865 -5 1885
rect -75 1835 -5 1865
rect -75 1815 -70 1835
rect -50 1815 -30 1835
rect -10 1815 -5 1835
rect -75 1785 -5 1815
rect -75 1765 -70 1785
rect -50 1765 -30 1785
rect -10 1765 -5 1785
rect -75 1755 -5 1765
rect 25 2085 55 2095
rect 25 2065 30 2085
rect 50 2065 55 2085
rect 25 2035 55 2065
rect 25 2015 30 2035
rect 50 2015 55 2035
rect 25 1985 55 2015
rect 25 1965 30 1985
rect 50 1965 55 1985
rect 25 1935 55 1965
rect 25 1915 30 1935
rect 50 1915 55 1935
rect 25 1885 55 1915
rect 25 1865 30 1885
rect 50 1865 55 1885
rect 25 1835 55 1865
rect 25 1815 30 1835
rect 50 1815 55 1835
rect 25 1785 55 1815
rect 25 1765 30 1785
rect 50 1765 55 1785
rect 25 1755 55 1765
rect 85 2085 115 2095
rect 85 2065 90 2085
rect 110 2065 115 2085
rect 85 2035 115 2065
rect 85 2015 90 2035
rect 110 2015 115 2035
rect 85 1985 115 2015
rect 85 1965 90 1985
rect 110 1965 115 1985
rect 85 1935 115 1965
rect 85 1915 90 1935
rect 110 1915 115 1935
rect 85 1885 115 1915
rect 85 1865 90 1885
rect 110 1865 115 1885
rect 85 1835 115 1865
rect 85 1815 90 1835
rect 110 1815 115 1835
rect 85 1785 115 1815
rect 85 1765 90 1785
rect 110 1765 115 1785
rect 85 1755 115 1765
rect 145 2085 175 2095
rect 145 2065 150 2085
rect 170 2065 175 2085
rect 145 2035 175 2065
rect 145 2015 150 2035
rect 170 2015 175 2035
rect 145 1985 175 2015
rect 145 1965 150 1985
rect 170 1965 175 1985
rect 145 1935 175 1965
rect 145 1915 150 1935
rect 170 1915 175 1935
rect 145 1885 175 1915
rect 145 1865 150 1885
rect 170 1865 175 1885
rect 145 1835 175 1865
rect 145 1815 150 1835
rect 170 1815 175 1835
rect 145 1785 175 1815
rect 145 1765 150 1785
rect 170 1765 175 1785
rect 145 1755 175 1765
rect 205 2085 235 2095
rect 205 2065 210 2085
rect 230 2065 235 2085
rect 205 2035 235 2065
rect 205 2015 210 2035
rect 230 2015 235 2035
rect 205 1985 235 2015
rect 205 1965 210 1985
rect 230 1965 235 1985
rect 205 1935 235 1965
rect 205 1915 210 1935
rect 230 1915 235 1935
rect 205 1885 235 1915
rect 205 1865 210 1885
rect 230 1865 235 1885
rect 205 1835 235 1865
rect 205 1815 210 1835
rect 230 1815 235 1835
rect 205 1785 235 1815
rect 205 1765 210 1785
rect 230 1765 235 1785
rect 205 1755 235 1765
rect 265 2085 295 2095
rect 265 2065 270 2085
rect 290 2065 295 2085
rect 265 2035 295 2065
rect 265 2015 270 2035
rect 290 2015 295 2035
rect 265 1985 295 2015
rect 265 1965 270 1985
rect 290 1965 295 1985
rect 265 1935 295 1965
rect 265 1915 270 1935
rect 290 1915 295 1935
rect 265 1885 295 1915
rect 265 1865 270 1885
rect 290 1865 295 1885
rect 265 1835 295 1865
rect 265 1815 270 1835
rect 290 1815 295 1835
rect 265 1785 295 1815
rect 265 1765 270 1785
rect 290 1765 295 1785
rect 265 1755 295 1765
rect 325 2085 355 2095
rect 325 2065 330 2085
rect 350 2065 355 2085
rect 325 2035 355 2065
rect 325 2015 330 2035
rect 350 2015 355 2035
rect 325 1985 355 2015
rect 325 1965 330 1985
rect 350 1965 355 1985
rect 325 1935 355 1965
rect 325 1915 330 1935
rect 350 1915 355 1935
rect 325 1885 355 1915
rect 325 1865 330 1885
rect 350 1865 355 1885
rect 325 1835 355 1865
rect 325 1815 330 1835
rect 350 1815 355 1835
rect 325 1785 355 1815
rect 325 1765 330 1785
rect 350 1765 355 1785
rect 325 1755 355 1765
rect 385 2085 415 2095
rect 385 2065 390 2085
rect 410 2065 415 2085
rect 385 2035 415 2065
rect 385 2015 390 2035
rect 410 2015 415 2035
rect 385 1985 415 2015
rect 385 1965 390 1985
rect 410 1965 415 1985
rect 385 1935 415 1965
rect 385 1915 390 1935
rect 410 1915 415 1935
rect 385 1885 415 1915
rect 385 1865 390 1885
rect 410 1865 415 1885
rect 385 1835 415 1865
rect 385 1815 390 1835
rect 410 1815 415 1835
rect 385 1785 415 1815
rect 385 1765 390 1785
rect 410 1765 415 1785
rect 385 1755 415 1765
rect 445 2085 475 2095
rect 445 2065 450 2085
rect 470 2065 475 2085
rect 445 2035 475 2065
rect 445 2015 450 2035
rect 470 2015 475 2035
rect 445 1985 475 2015
rect 445 1965 450 1985
rect 470 1965 475 1985
rect 445 1935 475 1965
rect 445 1915 450 1935
rect 470 1915 475 1935
rect 445 1885 475 1915
rect 445 1865 450 1885
rect 470 1865 475 1885
rect 445 1835 475 1865
rect 445 1815 450 1835
rect 470 1815 475 1835
rect 445 1785 475 1815
rect 445 1765 450 1785
rect 470 1765 475 1785
rect 445 1755 475 1765
rect 505 2085 535 2095
rect 505 2065 510 2085
rect 530 2065 535 2085
rect 505 2035 535 2065
rect 505 2015 510 2035
rect 530 2015 535 2035
rect 505 1985 535 2015
rect 505 1965 510 1985
rect 530 1965 535 1985
rect 505 1935 535 1965
rect 505 1915 510 1935
rect 530 1915 535 1935
rect 505 1885 535 1915
rect 505 1865 510 1885
rect 530 1865 535 1885
rect 505 1835 535 1865
rect 505 1815 510 1835
rect 530 1815 535 1835
rect 505 1785 535 1815
rect 505 1765 510 1785
rect 530 1765 535 1785
rect 505 1755 535 1765
rect 565 2085 595 2095
rect 565 2065 570 2085
rect 590 2065 595 2085
rect 565 2035 595 2065
rect 565 2015 570 2035
rect 590 2015 595 2035
rect 565 1985 595 2015
rect 565 1965 570 1985
rect 590 1965 595 1985
rect 565 1935 595 1965
rect 565 1915 570 1935
rect 590 1915 595 1935
rect 565 1885 595 1915
rect 565 1865 570 1885
rect 590 1865 595 1885
rect 565 1835 595 1865
rect 565 1815 570 1835
rect 590 1815 595 1835
rect 565 1785 595 1815
rect 565 1765 570 1785
rect 590 1765 595 1785
rect 565 1755 595 1765
rect 625 2085 655 2095
rect 625 2065 630 2085
rect 650 2065 655 2085
rect 625 2035 655 2065
rect 625 2015 630 2035
rect 650 2015 655 2035
rect 625 1985 655 2015
rect 625 1965 630 1985
rect 650 1965 655 1985
rect 625 1935 655 1965
rect 625 1915 630 1935
rect 650 1915 655 1935
rect 625 1885 655 1915
rect 625 1865 630 1885
rect 650 1865 655 1885
rect 625 1835 655 1865
rect 625 1815 630 1835
rect 650 1815 655 1835
rect 625 1785 655 1815
rect 625 1765 630 1785
rect 650 1765 655 1785
rect 625 1755 655 1765
rect 685 2085 755 2095
rect 685 2065 690 2085
rect 710 2065 730 2085
rect 750 2065 755 2085
rect 685 2035 755 2065
rect 685 2015 690 2035
rect 710 2015 730 2035
rect 750 2015 755 2035
rect 685 1985 755 2015
rect 685 1965 690 1985
rect 710 1965 730 1985
rect 750 1965 755 1985
rect 685 1935 755 1965
rect 685 1915 690 1935
rect 710 1915 730 1935
rect 750 1915 755 1935
rect 685 1885 755 1915
rect 685 1865 690 1885
rect 710 1865 730 1885
rect 750 1865 755 1885
rect 685 1835 755 1865
rect 685 1815 690 1835
rect 710 1815 730 1835
rect 750 1815 755 1835
rect 685 1785 755 1815
rect 685 1765 690 1785
rect 710 1765 730 1785
rect 750 1765 755 1785
rect 685 1755 755 1765
rect 935 2085 1005 2095
rect 935 2065 940 2085
rect 960 2065 980 2085
rect 1000 2065 1005 2085
rect 935 2035 1005 2065
rect 935 2015 940 2035
rect 960 2015 980 2035
rect 1000 2015 1005 2035
rect 935 1985 1005 2015
rect 935 1965 940 1985
rect 960 1965 980 1985
rect 1000 1965 1005 1985
rect 935 1935 1005 1965
rect 935 1915 940 1935
rect 960 1915 980 1935
rect 1000 1915 1005 1935
rect 935 1885 1005 1915
rect 935 1865 940 1885
rect 960 1865 980 1885
rect 1000 1865 1005 1885
rect 935 1835 1005 1865
rect 935 1815 940 1835
rect 960 1815 980 1835
rect 1000 1815 1005 1835
rect 935 1785 1005 1815
rect 935 1765 940 1785
rect 960 1765 980 1785
rect 1000 1765 1005 1785
rect 935 1755 1005 1765
rect 1035 2085 1065 2095
rect 1035 2065 1040 2085
rect 1060 2065 1065 2085
rect 1035 2035 1065 2065
rect 1035 2015 1040 2035
rect 1060 2015 1065 2035
rect 1035 1985 1065 2015
rect 1035 1965 1040 1985
rect 1060 1965 1065 1985
rect 1035 1935 1065 1965
rect 1035 1915 1040 1935
rect 1060 1915 1065 1935
rect 1035 1885 1065 1915
rect 1035 1865 1040 1885
rect 1060 1865 1065 1885
rect 1035 1835 1065 1865
rect 1035 1815 1040 1835
rect 1060 1815 1065 1835
rect 1035 1785 1065 1815
rect 1035 1765 1040 1785
rect 1060 1765 1065 1785
rect 1035 1755 1065 1765
rect 1095 2085 1125 2095
rect 1095 2065 1100 2085
rect 1120 2065 1125 2085
rect 1095 2035 1125 2065
rect 1095 2015 1100 2035
rect 1120 2015 1125 2035
rect 1095 1985 1125 2015
rect 1095 1965 1100 1985
rect 1120 1965 1125 1985
rect 1095 1935 1125 1965
rect 1095 1915 1100 1935
rect 1120 1915 1125 1935
rect 1095 1885 1125 1915
rect 1095 1865 1100 1885
rect 1120 1865 1125 1885
rect 1095 1835 1125 1865
rect 1095 1815 1100 1835
rect 1120 1815 1125 1835
rect 1095 1785 1125 1815
rect 1095 1765 1100 1785
rect 1120 1765 1125 1785
rect 1095 1755 1125 1765
rect 1155 2085 1185 2095
rect 1155 2065 1160 2085
rect 1180 2065 1185 2085
rect 1155 2035 1185 2065
rect 1155 2015 1160 2035
rect 1180 2015 1185 2035
rect 1155 1985 1185 2015
rect 1155 1965 1160 1985
rect 1180 1965 1185 1985
rect 1155 1935 1185 1965
rect 1155 1915 1160 1935
rect 1180 1915 1185 1935
rect 1155 1885 1185 1915
rect 1155 1865 1160 1885
rect 1180 1865 1185 1885
rect 1155 1835 1185 1865
rect 1155 1815 1160 1835
rect 1180 1815 1185 1835
rect 1155 1785 1185 1815
rect 1155 1765 1160 1785
rect 1180 1765 1185 1785
rect 1155 1755 1185 1765
rect 1215 2085 1245 2095
rect 1215 2065 1220 2085
rect 1240 2065 1245 2085
rect 1215 2035 1245 2065
rect 1215 2015 1220 2035
rect 1240 2015 1245 2035
rect 1215 1985 1245 2015
rect 1215 1965 1220 1985
rect 1240 1965 1245 1985
rect 1215 1935 1245 1965
rect 1215 1915 1220 1935
rect 1240 1915 1245 1935
rect 1215 1885 1245 1915
rect 1215 1865 1220 1885
rect 1240 1865 1245 1885
rect 1215 1835 1245 1865
rect 1215 1815 1220 1835
rect 1240 1815 1245 1835
rect 1215 1785 1245 1815
rect 1215 1765 1220 1785
rect 1240 1765 1245 1785
rect 1215 1755 1245 1765
rect 1275 2085 1305 2095
rect 1275 2065 1280 2085
rect 1300 2065 1305 2085
rect 1275 2035 1305 2065
rect 1275 2015 1280 2035
rect 1300 2015 1305 2035
rect 1275 1985 1305 2015
rect 1275 1965 1280 1985
rect 1300 1965 1305 1985
rect 1275 1935 1305 1965
rect 1275 1915 1280 1935
rect 1300 1915 1305 1935
rect 1275 1885 1305 1915
rect 1275 1865 1280 1885
rect 1300 1865 1305 1885
rect 1275 1835 1305 1865
rect 1275 1815 1280 1835
rect 1300 1815 1305 1835
rect 1275 1785 1305 1815
rect 1275 1765 1280 1785
rect 1300 1765 1305 1785
rect 1275 1755 1305 1765
rect 1335 2085 1365 2095
rect 1335 2065 1340 2085
rect 1360 2065 1365 2085
rect 1335 2035 1365 2065
rect 1335 2015 1340 2035
rect 1360 2015 1365 2035
rect 1335 1985 1365 2015
rect 1335 1965 1340 1985
rect 1360 1965 1365 1985
rect 1335 1935 1365 1965
rect 1335 1915 1340 1935
rect 1360 1915 1365 1935
rect 1335 1885 1365 1915
rect 1335 1865 1340 1885
rect 1360 1865 1365 1885
rect 1335 1835 1365 1865
rect 1335 1815 1340 1835
rect 1360 1815 1365 1835
rect 1335 1785 1365 1815
rect 1335 1765 1340 1785
rect 1360 1765 1365 1785
rect 1335 1755 1365 1765
rect 1395 2085 1425 2095
rect 1395 2065 1400 2085
rect 1420 2065 1425 2085
rect 1395 2035 1425 2065
rect 1395 2015 1400 2035
rect 1420 2015 1425 2035
rect 1395 1985 1425 2015
rect 1395 1965 1400 1985
rect 1420 1965 1425 1985
rect 1395 1935 1425 1965
rect 1395 1915 1400 1935
rect 1420 1915 1425 1935
rect 1395 1885 1425 1915
rect 1395 1865 1400 1885
rect 1420 1865 1425 1885
rect 1395 1835 1425 1865
rect 1395 1815 1400 1835
rect 1420 1815 1425 1835
rect 1395 1785 1425 1815
rect 1395 1765 1400 1785
rect 1420 1765 1425 1785
rect 1395 1755 1425 1765
rect 1455 2085 1485 2095
rect 1455 2065 1460 2085
rect 1480 2065 1485 2085
rect 1455 2035 1485 2065
rect 1455 2015 1460 2035
rect 1480 2015 1485 2035
rect 1455 1985 1485 2015
rect 1455 1965 1460 1985
rect 1480 1965 1485 1985
rect 1455 1935 1485 1965
rect 1455 1915 1460 1935
rect 1480 1915 1485 1935
rect 1455 1885 1485 1915
rect 1455 1865 1460 1885
rect 1480 1865 1485 1885
rect 1455 1835 1485 1865
rect 1455 1815 1460 1835
rect 1480 1815 1485 1835
rect 1455 1785 1485 1815
rect 1455 1765 1460 1785
rect 1480 1765 1485 1785
rect 1455 1755 1485 1765
rect 1515 2085 1545 2095
rect 1515 2065 1520 2085
rect 1540 2065 1545 2085
rect 1515 2035 1545 2065
rect 1515 2015 1520 2035
rect 1540 2015 1545 2035
rect 1515 1985 1545 2015
rect 1515 1965 1520 1985
rect 1540 1965 1545 1985
rect 1515 1935 1545 1965
rect 1515 1915 1520 1935
rect 1540 1915 1545 1935
rect 1515 1885 1545 1915
rect 1515 1865 1520 1885
rect 1540 1865 1545 1885
rect 1515 1835 1545 1865
rect 1515 1815 1520 1835
rect 1540 1815 1545 1835
rect 1515 1785 1545 1815
rect 1515 1765 1520 1785
rect 1540 1765 1545 1785
rect 1515 1755 1545 1765
rect 1575 2085 1605 2095
rect 1575 2065 1580 2085
rect 1600 2065 1605 2085
rect 1575 2035 1605 2065
rect 1575 2015 1580 2035
rect 1600 2015 1605 2035
rect 1575 1985 1605 2015
rect 1575 1965 1580 1985
rect 1600 1965 1605 1985
rect 1575 1935 1605 1965
rect 1575 1915 1580 1935
rect 1600 1915 1605 1935
rect 1575 1885 1605 1915
rect 1575 1865 1580 1885
rect 1600 1865 1605 1885
rect 1575 1835 1605 1865
rect 1575 1815 1580 1835
rect 1600 1815 1605 1835
rect 1575 1785 1605 1815
rect 1575 1765 1580 1785
rect 1600 1765 1605 1785
rect 1575 1755 1605 1765
rect 1635 2085 1665 2095
rect 1635 2065 1640 2085
rect 1660 2065 1665 2085
rect 1635 2035 1665 2065
rect 1635 2015 1640 2035
rect 1660 2015 1665 2035
rect 1635 1985 1665 2015
rect 1635 1965 1640 1985
rect 1660 1965 1665 1985
rect 1635 1935 1665 1965
rect 1635 1915 1640 1935
rect 1660 1915 1665 1935
rect 1635 1885 1665 1915
rect 1635 1865 1640 1885
rect 1660 1865 1665 1885
rect 1635 1835 1665 1865
rect 1635 1815 1640 1835
rect 1660 1815 1665 1835
rect 1635 1785 1665 1815
rect 1635 1765 1640 1785
rect 1660 1765 1665 1785
rect 1635 1755 1665 1765
rect 1695 2085 1765 2095
rect 1695 2065 1700 2085
rect 1720 2065 1740 2085
rect 1760 2065 1765 2085
rect 1695 2035 1765 2065
rect 1695 2015 1700 2035
rect 1720 2015 1740 2035
rect 1760 2015 1765 2035
rect 1695 1985 1765 2015
rect 1695 1965 1700 1985
rect 1720 1965 1740 1985
rect 1760 1965 1765 1985
rect 1695 1935 1765 1965
rect 1695 1915 1700 1935
rect 1720 1915 1740 1935
rect 1760 1915 1765 1935
rect 1695 1885 1765 1915
rect 1695 1865 1700 1885
rect 1720 1865 1740 1885
rect 1760 1865 1765 1885
rect 1695 1835 1765 1865
rect 1695 1815 1700 1835
rect 1720 1815 1740 1835
rect 1760 1815 1765 1835
rect 1695 1785 1765 1815
rect 1695 1765 1700 1785
rect 1720 1765 1740 1785
rect 1760 1765 1765 1785
rect 1695 1755 1765 1765
rect 1980 2085 2050 2095
rect 1980 2065 1985 2085
rect 2005 2065 2025 2085
rect 2045 2065 2050 2085
rect 1980 2035 2050 2065
rect 1980 2015 1985 2035
rect 2005 2015 2025 2035
rect 2045 2015 2050 2035
rect 1980 1985 2050 2015
rect 1980 1965 1985 1985
rect 2005 1965 2025 1985
rect 2045 1965 2050 1985
rect 1980 1935 2050 1965
rect 1980 1915 1985 1935
rect 2005 1915 2025 1935
rect 2045 1915 2050 1935
rect 1980 1885 2050 1915
rect 1980 1865 1985 1885
rect 2005 1865 2025 1885
rect 2045 1865 2050 1885
rect 1980 1835 2050 1865
rect 1980 1815 1985 1835
rect 2005 1815 2025 1835
rect 2045 1815 2050 1835
rect 1980 1785 2050 1815
rect 1980 1765 1985 1785
rect 2005 1765 2025 1785
rect 2045 1765 2050 1785
rect 1980 1755 2050 1765
rect 2080 2085 2110 2095
rect 2080 2065 2085 2085
rect 2105 2065 2110 2085
rect 2080 2035 2110 2065
rect 2080 2015 2085 2035
rect 2105 2015 2110 2035
rect 2080 1985 2110 2015
rect 2080 1965 2085 1985
rect 2105 1965 2110 1985
rect 2080 1935 2110 1965
rect 2080 1915 2085 1935
rect 2105 1915 2110 1935
rect 2080 1885 2110 1915
rect 2080 1865 2085 1885
rect 2105 1865 2110 1885
rect 2080 1835 2110 1865
rect 2080 1815 2085 1835
rect 2105 1815 2110 1835
rect 2080 1785 2110 1815
rect 2080 1765 2085 1785
rect 2105 1765 2110 1785
rect 2080 1755 2110 1765
rect 2140 2085 2170 2095
rect 2140 2065 2145 2085
rect 2165 2065 2170 2085
rect 2140 2035 2170 2065
rect 2140 2015 2145 2035
rect 2165 2015 2170 2035
rect 2140 1985 2170 2015
rect 2140 1965 2145 1985
rect 2165 1965 2170 1985
rect 2140 1935 2170 1965
rect 2140 1915 2145 1935
rect 2165 1915 2170 1935
rect 2140 1885 2170 1915
rect 2140 1865 2145 1885
rect 2165 1865 2170 1885
rect 2140 1835 2170 1865
rect 2140 1815 2145 1835
rect 2165 1815 2170 1835
rect 2140 1785 2170 1815
rect 2140 1765 2145 1785
rect 2165 1765 2170 1785
rect 2140 1755 2170 1765
rect 2200 2085 2230 2095
rect 2200 2065 2205 2085
rect 2225 2065 2230 2085
rect 2200 2035 2230 2065
rect 2200 2015 2205 2035
rect 2225 2015 2230 2035
rect 2200 1985 2230 2015
rect 2200 1965 2205 1985
rect 2225 1965 2230 1985
rect 2200 1935 2230 1965
rect 2200 1915 2205 1935
rect 2225 1915 2230 1935
rect 2200 1885 2230 1915
rect 2200 1865 2205 1885
rect 2225 1865 2230 1885
rect 2200 1835 2230 1865
rect 2200 1815 2205 1835
rect 2225 1815 2230 1835
rect 2200 1785 2230 1815
rect 2200 1765 2205 1785
rect 2225 1765 2230 1785
rect 2200 1755 2230 1765
rect 2260 2085 2290 2095
rect 2260 2065 2265 2085
rect 2285 2065 2290 2085
rect 2260 2035 2290 2065
rect 2260 2015 2265 2035
rect 2285 2015 2290 2035
rect 2260 1985 2290 2015
rect 2260 1965 2265 1985
rect 2285 1965 2290 1985
rect 2260 1935 2290 1965
rect 2260 1915 2265 1935
rect 2285 1915 2290 1935
rect 2260 1885 2290 1915
rect 2260 1865 2265 1885
rect 2285 1865 2290 1885
rect 2260 1835 2290 1865
rect 2260 1815 2265 1835
rect 2285 1815 2290 1835
rect 2260 1785 2290 1815
rect 2260 1765 2265 1785
rect 2285 1765 2290 1785
rect 2260 1755 2290 1765
rect 2320 2085 2350 2095
rect 2320 2065 2325 2085
rect 2345 2065 2350 2085
rect 2320 2035 2350 2065
rect 2320 2015 2325 2035
rect 2345 2015 2350 2035
rect 2320 1985 2350 2015
rect 2320 1965 2325 1985
rect 2345 1965 2350 1985
rect 2320 1935 2350 1965
rect 2320 1915 2325 1935
rect 2345 1915 2350 1935
rect 2320 1885 2350 1915
rect 2320 1865 2325 1885
rect 2345 1865 2350 1885
rect 2320 1835 2350 1865
rect 2320 1815 2325 1835
rect 2345 1815 2350 1835
rect 2320 1785 2350 1815
rect 2320 1765 2325 1785
rect 2345 1765 2350 1785
rect 2320 1755 2350 1765
rect 2380 2085 2410 2095
rect 2380 2065 2385 2085
rect 2405 2065 2410 2085
rect 2380 2035 2410 2065
rect 2380 2015 2385 2035
rect 2405 2015 2410 2035
rect 2380 1985 2410 2015
rect 2380 1965 2385 1985
rect 2405 1965 2410 1985
rect 2380 1935 2410 1965
rect 2380 1915 2385 1935
rect 2405 1915 2410 1935
rect 2380 1885 2410 1915
rect 2380 1865 2385 1885
rect 2405 1865 2410 1885
rect 2380 1835 2410 1865
rect 2380 1815 2385 1835
rect 2405 1815 2410 1835
rect 2380 1785 2410 1815
rect 2380 1765 2385 1785
rect 2405 1765 2410 1785
rect 2380 1755 2410 1765
rect 2440 2085 2470 2095
rect 2440 2065 2445 2085
rect 2465 2065 2470 2085
rect 2440 2035 2470 2065
rect 2440 2015 2445 2035
rect 2465 2015 2470 2035
rect 2440 1985 2470 2015
rect 2440 1965 2445 1985
rect 2465 1965 2470 1985
rect 2440 1935 2470 1965
rect 2440 1915 2445 1935
rect 2465 1915 2470 1935
rect 2440 1885 2470 1915
rect 2440 1865 2445 1885
rect 2465 1865 2470 1885
rect 2440 1835 2470 1865
rect 2440 1815 2445 1835
rect 2465 1815 2470 1835
rect 2440 1785 2470 1815
rect 2440 1765 2445 1785
rect 2465 1765 2470 1785
rect 2440 1755 2470 1765
rect 2500 2085 2530 2095
rect 2500 2065 2505 2085
rect 2525 2065 2530 2085
rect 2500 2035 2530 2065
rect 2500 2015 2505 2035
rect 2525 2015 2530 2035
rect 2500 1985 2530 2015
rect 2500 1965 2505 1985
rect 2525 1965 2530 1985
rect 2500 1935 2530 1965
rect 2500 1915 2505 1935
rect 2525 1915 2530 1935
rect 2500 1885 2530 1915
rect 2500 1865 2505 1885
rect 2525 1865 2530 1885
rect 2500 1835 2530 1865
rect 2500 1815 2505 1835
rect 2525 1815 2530 1835
rect 2500 1785 2530 1815
rect 2500 1765 2505 1785
rect 2525 1765 2530 1785
rect 2500 1755 2530 1765
rect 2560 2085 2590 2095
rect 2560 2065 2565 2085
rect 2585 2065 2590 2085
rect 2560 2035 2590 2065
rect 2560 2015 2565 2035
rect 2585 2015 2590 2035
rect 2560 1985 2590 2015
rect 2560 1965 2565 1985
rect 2585 1965 2590 1985
rect 2560 1935 2590 1965
rect 2560 1915 2565 1935
rect 2585 1915 2590 1935
rect 2560 1885 2590 1915
rect 2560 1865 2565 1885
rect 2585 1865 2590 1885
rect 2560 1835 2590 1865
rect 2560 1815 2565 1835
rect 2585 1815 2590 1835
rect 2560 1785 2590 1815
rect 2560 1765 2565 1785
rect 2585 1765 2590 1785
rect 2560 1755 2590 1765
rect 2620 2085 2650 2095
rect 2620 2065 2625 2085
rect 2645 2065 2650 2085
rect 2620 2035 2650 2065
rect 2620 2015 2625 2035
rect 2645 2015 2650 2035
rect 2620 1985 2650 2015
rect 2620 1965 2625 1985
rect 2645 1965 2650 1985
rect 2620 1935 2650 1965
rect 2620 1915 2625 1935
rect 2645 1915 2650 1935
rect 2620 1885 2650 1915
rect 2620 1865 2625 1885
rect 2645 1865 2650 1885
rect 2620 1835 2650 1865
rect 2620 1815 2625 1835
rect 2645 1815 2650 1835
rect 2620 1785 2650 1815
rect 2620 1765 2625 1785
rect 2645 1765 2650 1785
rect 2620 1755 2650 1765
rect 2680 2085 2710 2095
rect 2680 2065 2685 2085
rect 2705 2065 2710 2085
rect 2680 2035 2710 2065
rect 2680 2015 2685 2035
rect 2705 2015 2710 2035
rect 2680 1985 2710 2015
rect 2680 1965 2685 1985
rect 2705 1965 2710 1985
rect 2680 1935 2710 1965
rect 2680 1915 2685 1935
rect 2705 1915 2710 1935
rect 2680 1885 2710 1915
rect 2680 1865 2685 1885
rect 2705 1865 2710 1885
rect 2680 1835 2710 1865
rect 2680 1815 2685 1835
rect 2705 1815 2710 1835
rect 2680 1785 2710 1815
rect 2680 1765 2685 1785
rect 2705 1765 2710 1785
rect 2680 1755 2710 1765
rect 2740 2085 2810 2095
rect 2740 2065 2745 2085
rect 2765 2065 2785 2085
rect 2805 2065 2810 2085
rect 2740 2035 2810 2065
rect 2740 2015 2745 2035
rect 2765 2015 2785 2035
rect 2805 2015 2810 2035
rect 2740 1985 2810 2015
rect 2740 1965 2745 1985
rect 2765 1965 2785 1985
rect 2805 1965 2810 1985
rect 2740 1935 2810 1965
rect 2740 1915 2745 1935
rect 2765 1915 2785 1935
rect 2805 1915 2810 1935
rect 2740 1885 2810 1915
rect 2740 1865 2745 1885
rect 2765 1865 2785 1885
rect 2805 1865 2810 1885
rect 2740 1835 2810 1865
rect 2740 1815 2745 1835
rect 2765 1815 2785 1835
rect 2805 1815 2810 1835
rect 2740 1785 2810 1815
rect 2740 1765 2745 1785
rect 2765 1765 2785 1785
rect 2805 1765 2810 1785
rect 2740 1755 2810 1765
rect -1015 1730 -995 1755
rect -895 1730 -875 1755
rect -775 1730 -755 1755
rect -655 1730 -635 1755
rect -535 1730 -515 1755
rect -415 1730 -395 1755
rect 30 1730 50 1755
rect 150 1730 170 1755
rect 270 1730 290 1755
rect 390 1730 410 1755
rect 510 1730 530 1755
rect 630 1730 650 1755
rect 1040 1730 1060 1755
rect 1160 1730 1180 1755
rect 1280 1730 1300 1755
rect 1400 1730 1420 1755
rect 1520 1730 1540 1755
rect 1640 1730 1660 1755
rect 2085 1730 2105 1755
rect 2205 1730 2225 1755
rect 2325 1730 2345 1755
rect 2445 1730 2465 1755
rect 2565 1730 2585 1755
rect 2685 1730 2705 1755
rect -1025 1720 -985 1730
rect -1025 1700 -1015 1720
rect -995 1700 -985 1720
rect -1025 1690 -985 1700
rect -905 1720 -865 1730
rect -905 1700 -895 1720
rect -875 1700 -865 1720
rect -905 1690 -865 1700
rect -785 1720 -745 1730
rect -785 1700 -775 1720
rect -755 1700 -745 1720
rect -785 1690 -745 1700
rect -720 1720 -690 1730
rect -720 1700 -715 1720
rect -695 1700 -690 1720
rect -720 1690 -690 1700
rect -665 1720 -625 1730
rect -665 1700 -655 1720
rect -635 1700 -625 1720
rect -665 1690 -625 1700
rect -545 1720 -505 1730
rect -545 1700 -535 1720
rect -515 1700 -505 1720
rect -545 1690 -505 1700
rect -425 1720 -385 1730
rect -425 1700 -415 1720
rect -395 1700 -385 1720
rect -425 1690 -385 1700
rect 20 1720 60 1730
rect 20 1700 30 1720
rect 50 1700 60 1720
rect 20 1690 60 1700
rect 140 1720 180 1730
rect 140 1700 150 1720
rect 170 1700 180 1720
rect 140 1690 180 1700
rect 260 1720 300 1730
rect 260 1700 270 1720
rect 290 1700 300 1720
rect 260 1690 300 1700
rect 325 1720 355 1730
rect 325 1700 330 1720
rect 350 1700 355 1720
rect 325 1690 355 1700
rect 380 1720 420 1730
rect 380 1700 390 1720
rect 410 1700 420 1720
rect 380 1690 420 1700
rect 500 1720 540 1730
rect 500 1700 510 1720
rect 530 1700 540 1720
rect 500 1690 540 1700
rect 620 1720 660 1730
rect 620 1700 630 1720
rect 650 1700 660 1720
rect 620 1690 660 1700
rect 1030 1720 1070 1730
rect 1030 1700 1040 1720
rect 1060 1700 1070 1720
rect 1030 1690 1070 1700
rect 1150 1720 1190 1730
rect 1150 1700 1160 1720
rect 1180 1700 1190 1720
rect 1150 1690 1190 1700
rect 1270 1720 1310 1730
rect 1270 1700 1280 1720
rect 1300 1700 1310 1720
rect 1270 1690 1310 1700
rect 1335 1720 1365 1730
rect 1335 1700 1340 1720
rect 1360 1700 1365 1720
rect 1335 1690 1365 1700
rect 1390 1720 1430 1730
rect 1390 1700 1400 1720
rect 1420 1700 1430 1720
rect 1390 1690 1430 1700
rect 1510 1720 1550 1730
rect 1510 1700 1520 1720
rect 1540 1700 1550 1720
rect 1510 1690 1550 1700
rect 1630 1720 1670 1730
rect 1630 1700 1640 1720
rect 1660 1700 1670 1720
rect 1630 1690 1670 1700
rect 2075 1720 2115 1730
rect 2075 1700 2085 1720
rect 2105 1700 2115 1720
rect 2075 1690 2115 1700
rect 2195 1720 2235 1730
rect 2195 1700 2205 1720
rect 2225 1700 2235 1720
rect 2195 1690 2235 1700
rect 2315 1720 2355 1730
rect 2315 1700 2325 1720
rect 2345 1700 2355 1720
rect 2315 1690 2355 1700
rect 2380 1720 2410 1730
rect 2380 1700 2385 1720
rect 2405 1700 2410 1720
rect 2380 1690 2410 1700
rect 2435 1720 2475 1730
rect 2435 1700 2445 1720
rect 2465 1700 2475 1720
rect 2435 1690 2475 1700
rect 2555 1720 2595 1730
rect 2555 1700 2565 1720
rect 2585 1700 2595 1720
rect 2555 1690 2595 1700
rect 2675 1720 2715 1730
rect 2675 1700 2685 1720
rect 2705 1700 2715 1720
rect 2675 1690 2715 1700
rect 220 1575 260 1585
rect 220 1555 230 1575
rect 250 1555 260 1575
rect 220 1545 260 1555
rect 330 1575 370 1585
rect 330 1555 340 1575
rect 360 1555 370 1575
rect 330 1545 370 1555
rect 440 1575 480 1585
rect 440 1555 450 1575
rect 470 1555 480 1575
rect 440 1545 480 1555
rect 550 1575 590 1585
rect 550 1555 560 1575
rect 580 1555 590 1575
rect 550 1545 590 1555
rect 660 1575 700 1585
rect 660 1555 670 1575
rect 690 1555 700 1575
rect 660 1545 700 1555
rect 770 1575 810 1585
rect 770 1555 780 1575
rect 800 1555 810 1575
rect 770 1545 810 1555
rect 880 1575 920 1585
rect 880 1555 890 1575
rect 910 1555 920 1575
rect 880 1545 920 1555
rect 990 1575 1030 1585
rect 990 1555 1000 1575
rect 1020 1555 1030 1575
rect 990 1545 1030 1555
rect 1100 1575 1140 1585
rect 1100 1555 1110 1575
rect 1130 1555 1140 1575
rect 1100 1545 1140 1555
rect 1210 1575 1250 1585
rect 1210 1555 1220 1575
rect 1240 1555 1250 1575
rect 1210 1545 1250 1555
rect 1320 1575 1360 1585
rect 1320 1555 1330 1575
rect 1350 1555 1360 1575
rect 1320 1545 1360 1555
rect 1430 1575 1470 1585
rect 1430 1555 1440 1575
rect 1460 1555 1470 1575
rect 1430 1545 1470 1555
rect 230 1525 250 1545
rect 340 1525 360 1545
rect 450 1525 470 1545
rect 560 1525 580 1545
rect 670 1525 690 1545
rect 780 1525 800 1545
rect 890 1525 910 1545
rect 1000 1525 1020 1545
rect 1110 1525 1130 1545
rect 1220 1525 1240 1545
rect 1330 1525 1350 1545
rect 1440 1525 1460 1545
rect 185 1515 255 1525
rect 185 1495 190 1515
rect 210 1495 230 1515
rect 250 1495 255 1515
rect -1055 1480 -1015 1490
rect -1055 1460 -1045 1480
rect -1025 1460 -1015 1480
rect -1055 1450 -1015 1460
rect -945 1480 -905 1490
rect -945 1460 -935 1480
rect -915 1460 -905 1480
rect -945 1450 -905 1460
rect -835 1480 -795 1490
rect -835 1460 -825 1480
rect -805 1460 -795 1480
rect -835 1450 -795 1460
rect -725 1480 -685 1490
rect -725 1460 -715 1480
rect -695 1460 -685 1480
rect -725 1450 -685 1460
rect -615 1480 -575 1490
rect -615 1460 -605 1480
rect -585 1460 -575 1480
rect -615 1450 -575 1460
rect -505 1480 -465 1490
rect -505 1460 -495 1480
rect -475 1460 -465 1480
rect -505 1450 -465 1460
rect -395 1480 -355 1490
rect 185 1485 255 1495
rect 280 1515 310 1525
rect 280 1495 285 1515
rect 305 1495 310 1515
rect 280 1485 310 1495
rect 335 1515 365 1525
rect 335 1495 340 1515
rect 360 1495 365 1515
rect 335 1485 365 1495
rect 390 1515 420 1525
rect 390 1495 395 1515
rect 415 1495 420 1515
rect 390 1485 420 1495
rect 445 1515 475 1525
rect 445 1495 450 1515
rect 470 1495 475 1515
rect 445 1485 475 1495
rect 500 1515 530 1525
rect 500 1495 505 1515
rect 525 1495 530 1515
rect 500 1485 530 1495
rect 555 1515 585 1525
rect 555 1495 560 1515
rect 580 1495 585 1515
rect 555 1485 585 1495
rect 610 1515 640 1525
rect 610 1495 615 1515
rect 635 1495 640 1515
rect 610 1485 640 1495
rect 665 1515 695 1525
rect 665 1495 670 1515
rect 690 1495 695 1515
rect 665 1485 695 1495
rect 720 1515 750 1525
rect 720 1495 725 1515
rect 745 1495 750 1515
rect 720 1485 750 1495
rect 775 1515 805 1525
rect 775 1495 780 1515
rect 800 1495 805 1515
rect 775 1485 805 1495
rect 830 1515 860 1525
rect 830 1495 835 1515
rect 855 1495 860 1515
rect 830 1485 860 1495
rect 885 1515 915 1525
rect 885 1495 890 1515
rect 910 1495 915 1515
rect 885 1485 915 1495
rect 940 1515 970 1525
rect 940 1495 945 1515
rect 965 1495 970 1515
rect 940 1485 970 1495
rect 995 1515 1025 1525
rect 995 1495 1000 1515
rect 1020 1495 1025 1515
rect 995 1485 1025 1495
rect 1050 1515 1080 1525
rect 1050 1495 1055 1515
rect 1075 1495 1080 1515
rect 1050 1485 1080 1495
rect 1105 1515 1135 1525
rect 1105 1495 1110 1515
rect 1130 1495 1135 1515
rect 1105 1485 1135 1495
rect 1160 1515 1190 1525
rect 1160 1495 1165 1515
rect 1185 1495 1190 1515
rect 1160 1485 1190 1495
rect 1215 1515 1245 1525
rect 1215 1495 1220 1515
rect 1240 1495 1245 1515
rect 1215 1485 1245 1495
rect 1270 1515 1300 1525
rect 1270 1495 1275 1515
rect 1295 1495 1300 1515
rect 1270 1485 1300 1495
rect 1325 1515 1355 1525
rect 1325 1495 1330 1515
rect 1350 1495 1355 1515
rect 1325 1485 1355 1495
rect 1380 1515 1410 1525
rect 1380 1495 1385 1515
rect 1405 1495 1410 1515
rect 1380 1485 1410 1495
rect 1435 1515 1505 1525
rect 1435 1495 1440 1515
rect 1460 1495 1480 1515
rect 1500 1495 1505 1515
rect 1435 1485 1505 1495
rect -395 1460 -385 1480
rect -365 1460 -355 1480
rect 285 1460 305 1485
rect 395 1460 415 1485
rect 505 1460 525 1485
rect 615 1460 635 1485
rect 725 1460 745 1485
rect 835 1460 855 1485
rect 945 1460 965 1485
rect 1055 1460 1075 1485
rect 1165 1460 1185 1485
rect 1275 1460 1295 1485
rect 1385 1460 1405 1485
rect 2045 1480 2085 1490
rect 2045 1460 2055 1480
rect 2075 1460 2085 1480
rect -395 1450 -355 1460
rect 275 1450 315 1460
rect -1045 1430 -1025 1450
rect -935 1430 -915 1450
rect -825 1430 -805 1450
rect -715 1430 -695 1450
rect -605 1430 -585 1450
rect -495 1430 -475 1450
rect -385 1430 -365 1450
rect 275 1430 285 1450
rect 305 1430 315 1450
rect -1501 1420 -1360 1430
rect -1501 1400 -1495 1420
rect -1475 1400 -1440 1420
rect -1420 1400 -1385 1420
rect -1365 1400 -1360 1420
rect -1501 1390 -1360 1400
rect -1090 1420 -1020 1430
rect -1090 1400 -1085 1420
rect -1065 1400 -1045 1420
rect -1025 1400 -1020 1420
rect -1090 1370 -1020 1400
rect -1090 1350 -1085 1370
rect -1065 1350 -1045 1370
rect -1025 1350 -1020 1370
rect -1090 1320 -1020 1350
rect -1090 1300 -1085 1320
rect -1065 1300 -1045 1320
rect -1025 1300 -1020 1320
rect -1090 1270 -1020 1300
rect -1090 1250 -1085 1270
rect -1065 1250 -1045 1270
rect -1025 1250 -1020 1270
rect -1090 1220 -1020 1250
rect -1090 1200 -1085 1220
rect -1065 1200 -1045 1220
rect -1025 1200 -1020 1220
rect -1090 1170 -1020 1200
rect -1090 1150 -1085 1170
rect -1065 1150 -1045 1170
rect -1025 1150 -1020 1170
rect -1090 1120 -1020 1150
rect -1090 1100 -1085 1120
rect -1065 1100 -1045 1120
rect -1025 1100 -1020 1120
rect -1090 1070 -1020 1100
rect -1090 1050 -1085 1070
rect -1065 1050 -1045 1070
rect -1025 1050 -1020 1070
rect -1090 1020 -1020 1050
rect -1090 1000 -1085 1020
rect -1065 1000 -1045 1020
rect -1025 1000 -1020 1020
rect -1090 970 -1020 1000
rect -1090 950 -1085 970
rect -1065 950 -1045 970
rect -1025 950 -1020 970
rect -1090 920 -1020 950
rect -1090 900 -1085 920
rect -1065 900 -1045 920
rect -1025 900 -1020 920
rect -1090 870 -1020 900
rect -1090 850 -1085 870
rect -1065 850 -1045 870
rect -1025 850 -1020 870
rect -1090 840 -1020 850
rect -995 1420 -965 1430
rect -995 1400 -990 1420
rect -970 1400 -965 1420
rect -995 1370 -965 1400
rect -995 1350 -990 1370
rect -970 1350 -965 1370
rect -995 1320 -965 1350
rect -995 1300 -990 1320
rect -970 1300 -965 1320
rect -995 1270 -965 1300
rect -995 1250 -990 1270
rect -970 1250 -965 1270
rect -995 1220 -965 1250
rect -995 1200 -990 1220
rect -970 1200 -965 1220
rect -995 1170 -965 1200
rect -995 1150 -990 1170
rect -970 1150 -965 1170
rect -995 1120 -965 1150
rect -995 1100 -990 1120
rect -970 1100 -965 1120
rect -995 1070 -965 1100
rect -995 1050 -990 1070
rect -970 1050 -965 1070
rect -995 1020 -965 1050
rect -995 1000 -990 1020
rect -970 1000 -965 1020
rect -995 970 -965 1000
rect -995 950 -990 970
rect -970 950 -965 970
rect -995 920 -965 950
rect -995 900 -990 920
rect -970 900 -965 920
rect -995 870 -965 900
rect -995 850 -990 870
rect -970 850 -965 870
rect -995 840 -965 850
rect -940 1420 -910 1430
rect -940 1400 -935 1420
rect -915 1400 -910 1420
rect -940 1370 -910 1400
rect -940 1350 -935 1370
rect -915 1350 -910 1370
rect -940 1320 -910 1350
rect -940 1300 -935 1320
rect -915 1300 -910 1320
rect -940 1270 -910 1300
rect -940 1250 -935 1270
rect -915 1250 -910 1270
rect -940 1220 -910 1250
rect -940 1200 -935 1220
rect -915 1200 -910 1220
rect -940 1170 -910 1200
rect -940 1150 -935 1170
rect -915 1150 -910 1170
rect -940 1120 -910 1150
rect -940 1100 -935 1120
rect -915 1100 -910 1120
rect -940 1070 -910 1100
rect -940 1050 -935 1070
rect -915 1050 -910 1070
rect -940 1020 -910 1050
rect -940 1000 -935 1020
rect -915 1000 -910 1020
rect -940 970 -910 1000
rect -940 950 -935 970
rect -915 950 -910 970
rect -940 920 -910 950
rect -940 900 -935 920
rect -915 900 -910 920
rect -940 870 -910 900
rect -940 850 -935 870
rect -915 850 -910 870
rect -940 840 -910 850
rect -885 1420 -855 1430
rect -885 1400 -880 1420
rect -860 1400 -855 1420
rect -885 1370 -855 1400
rect -885 1350 -880 1370
rect -860 1350 -855 1370
rect -885 1320 -855 1350
rect -885 1300 -880 1320
rect -860 1300 -855 1320
rect -885 1270 -855 1300
rect -885 1250 -880 1270
rect -860 1250 -855 1270
rect -885 1220 -855 1250
rect -885 1200 -880 1220
rect -860 1200 -855 1220
rect -885 1170 -855 1200
rect -885 1150 -880 1170
rect -860 1150 -855 1170
rect -885 1120 -855 1150
rect -885 1100 -880 1120
rect -860 1100 -855 1120
rect -885 1070 -855 1100
rect -885 1050 -880 1070
rect -860 1050 -855 1070
rect -885 1020 -855 1050
rect -885 1000 -880 1020
rect -860 1000 -855 1020
rect -885 970 -855 1000
rect -885 950 -880 970
rect -860 950 -855 970
rect -885 920 -855 950
rect -885 900 -880 920
rect -860 900 -855 920
rect -885 870 -855 900
rect -885 850 -880 870
rect -860 850 -855 870
rect -885 840 -855 850
rect -830 1420 -800 1430
rect -830 1400 -825 1420
rect -805 1400 -800 1420
rect -830 1370 -800 1400
rect -830 1350 -825 1370
rect -805 1350 -800 1370
rect -830 1320 -800 1350
rect -830 1300 -825 1320
rect -805 1300 -800 1320
rect -830 1270 -800 1300
rect -830 1250 -825 1270
rect -805 1250 -800 1270
rect -830 1220 -800 1250
rect -830 1200 -825 1220
rect -805 1200 -800 1220
rect -830 1170 -800 1200
rect -830 1150 -825 1170
rect -805 1150 -800 1170
rect -830 1120 -800 1150
rect -830 1100 -825 1120
rect -805 1100 -800 1120
rect -830 1070 -800 1100
rect -830 1050 -825 1070
rect -805 1050 -800 1070
rect -830 1020 -800 1050
rect -830 1000 -825 1020
rect -805 1000 -800 1020
rect -830 970 -800 1000
rect -830 950 -825 970
rect -805 950 -800 970
rect -830 920 -800 950
rect -830 900 -825 920
rect -805 900 -800 920
rect -830 870 -800 900
rect -830 850 -825 870
rect -805 850 -800 870
rect -830 840 -800 850
rect -775 1420 -745 1430
rect -775 1400 -770 1420
rect -750 1400 -745 1420
rect -775 1370 -745 1400
rect -775 1350 -770 1370
rect -750 1350 -745 1370
rect -775 1320 -745 1350
rect -775 1300 -770 1320
rect -750 1300 -745 1320
rect -775 1270 -745 1300
rect -775 1250 -770 1270
rect -750 1250 -745 1270
rect -775 1220 -745 1250
rect -775 1200 -770 1220
rect -750 1200 -745 1220
rect -775 1170 -745 1200
rect -775 1150 -770 1170
rect -750 1150 -745 1170
rect -775 1120 -745 1150
rect -775 1100 -770 1120
rect -750 1100 -745 1120
rect -775 1070 -745 1100
rect -775 1050 -770 1070
rect -750 1050 -745 1070
rect -775 1020 -745 1050
rect -775 1000 -770 1020
rect -750 1000 -745 1020
rect -775 970 -745 1000
rect -775 950 -770 970
rect -750 950 -745 970
rect -775 920 -745 950
rect -775 900 -770 920
rect -750 900 -745 920
rect -775 870 -745 900
rect -775 850 -770 870
rect -750 850 -745 870
rect -775 840 -745 850
rect -720 1420 -690 1430
rect -720 1400 -715 1420
rect -695 1400 -690 1420
rect -720 1370 -690 1400
rect -720 1350 -715 1370
rect -695 1350 -690 1370
rect -720 1320 -690 1350
rect -720 1300 -715 1320
rect -695 1300 -690 1320
rect -720 1270 -690 1300
rect -720 1250 -715 1270
rect -695 1250 -690 1270
rect -720 1220 -690 1250
rect -720 1200 -715 1220
rect -695 1200 -690 1220
rect -720 1170 -690 1200
rect -720 1150 -715 1170
rect -695 1150 -690 1170
rect -720 1120 -690 1150
rect -720 1100 -715 1120
rect -695 1100 -690 1120
rect -720 1070 -690 1100
rect -720 1050 -715 1070
rect -695 1050 -690 1070
rect -720 1020 -690 1050
rect -720 1000 -715 1020
rect -695 1000 -690 1020
rect -720 970 -690 1000
rect -720 950 -715 970
rect -695 950 -690 970
rect -720 920 -690 950
rect -720 900 -715 920
rect -695 900 -690 920
rect -720 870 -690 900
rect -720 850 -715 870
rect -695 850 -690 870
rect -720 840 -690 850
rect -665 1420 -635 1430
rect -665 1400 -660 1420
rect -640 1400 -635 1420
rect -665 1370 -635 1400
rect -665 1350 -660 1370
rect -640 1350 -635 1370
rect -665 1320 -635 1350
rect -665 1300 -660 1320
rect -640 1300 -635 1320
rect -665 1270 -635 1300
rect -665 1250 -660 1270
rect -640 1250 -635 1270
rect -665 1220 -635 1250
rect -665 1200 -660 1220
rect -640 1200 -635 1220
rect -665 1170 -635 1200
rect -665 1150 -660 1170
rect -640 1150 -635 1170
rect -665 1120 -635 1150
rect -665 1100 -660 1120
rect -640 1100 -635 1120
rect -665 1070 -635 1100
rect -665 1050 -660 1070
rect -640 1050 -635 1070
rect -665 1020 -635 1050
rect -665 1000 -660 1020
rect -640 1000 -635 1020
rect -665 970 -635 1000
rect -665 950 -660 970
rect -640 950 -635 970
rect -665 920 -635 950
rect -665 900 -660 920
rect -640 900 -635 920
rect -665 870 -635 900
rect -665 850 -660 870
rect -640 850 -635 870
rect -665 840 -635 850
rect -610 1420 -580 1430
rect -610 1400 -605 1420
rect -585 1400 -580 1420
rect -610 1370 -580 1400
rect -610 1350 -605 1370
rect -585 1350 -580 1370
rect -610 1320 -580 1350
rect -610 1300 -605 1320
rect -585 1300 -580 1320
rect -610 1270 -580 1300
rect -610 1250 -605 1270
rect -585 1250 -580 1270
rect -610 1220 -580 1250
rect -610 1200 -605 1220
rect -585 1200 -580 1220
rect -610 1170 -580 1200
rect -610 1150 -605 1170
rect -585 1150 -580 1170
rect -610 1120 -580 1150
rect -610 1100 -605 1120
rect -585 1100 -580 1120
rect -610 1070 -580 1100
rect -610 1050 -605 1070
rect -585 1050 -580 1070
rect -610 1020 -580 1050
rect -610 1000 -605 1020
rect -585 1000 -580 1020
rect -610 970 -580 1000
rect -610 950 -605 970
rect -585 950 -580 970
rect -610 920 -580 950
rect -610 900 -605 920
rect -585 900 -580 920
rect -610 870 -580 900
rect -610 850 -605 870
rect -585 850 -580 870
rect -610 840 -580 850
rect -555 1420 -525 1430
rect -555 1400 -550 1420
rect -530 1400 -525 1420
rect -555 1370 -525 1400
rect -555 1350 -550 1370
rect -530 1350 -525 1370
rect -555 1320 -525 1350
rect -555 1300 -550 1320
rect -530 1300 -525 1320
rect -555 1270 -525 1300
rect -555 1250 -550 1270
rect -530 1250 -525 1270
rect -555 1220 -525 1250
rect -555 1200 -550 1220
rect -530 1200 -525 1220
rect -555 1170 -525 1200
rect -555 1150 -550 1170
rect -530 1150 -525 1170
rect -555 1120 -525 1150
rect -555 1100 -550 1120
rect -530 1100 -525 1120
rect -555 1070 -525 1100
rect -555 1050 -550 1070
rect -530 1050 -525 1070
rect -555 1020 -525 1050
rect -555 1000 -550 1020
rect -530 1000 -525 1020
rect -555 970 -525 1000
rect -555 950 -550 970
rect -530 950 -525 970
rect -555 920 -525 950
rect -555 900 -550 920
rect -530 900 -525 920
rect -555 870 -525 900
rect -555 850 -550 870
rect -530 850 -525 870
rect -555 840 -525 850
rect -500 1420 -470 1430
rect -500 1400 -495 1420
rect -475 1400 -470 1420
rect -500 1370 -470 1400
rect -500 1350 -495 1370
rect -475 1350 -470 1370
rect -500 1320 -470 1350
rect -500 1300 -495 1320
rect -475 1300 -470 1320
rect -500 1270 -470 1300
rect -500 1250 -495 1270
rect -475 1250 -470 1270
rect -500 1220 -470 1250
rect -500 1200 -495 1220
rect -475 1200 -470 1220
rect -500 1170 -470 1200
rect -500 1150 -495 1170
rect -475 1150 -470 1170
rect -500 1120 -470 1150
rect -500 1100 -495 1120
rect -475 1100 -470 1120
rect -500 1070 -470 1100
rect -500 1050 -495 1070
rect -475 1050 -470 1070
rect -500 1020 -470 1050
rect -500 1000 -495 1020
rect -475 1000 -470 1020
rect -500 970 -470 1000
rect -500 950 -495 970
rect -475 950 -470 970
rect -500 920 -470 950
rect -500 900 -495 920
rect -475 900 -470 920
rect -500 870 -470 900
rect -500 850 -495 870
rect -475 850 -470 870
rect -500 840 -470 850
rect -445 1420 -415 1430
rect -445 1400 -440 1420
rect -420 1400 -415 1420
rect -445 1370 -415 1400
rect -445 1350 -440 1370
rect -420 1350 -415 1370
rect -445 1320 -415 1350
rect -445 1300 -440 1320
rect -420 1300 -415 1320
rect -445 1270 -415 1300
rect -445 1250 -440 1270
rect -420 1250 -415 1270
rect -445 1220 -415 1250
rect -445 1200 -440 1220
rect -420 1200 -415 1220
rect -445 1170 -415 1200
rect -445 1150 -440 1170
rect -420 1150 -415 1170
rect -445 1120 -415 1150
rect -445 1100 -440 1120
rect -420 1100 -415 1120
rect -445 1070 -415 1100
rect -445 1050 -440 1070
rect -420 1050 -415 1070
rect -445 1020 -415 1050
rect -445 1000 -440 1020
rect -420 1000 -415 1020
rect -445 970 -415 1000
rect -445 950 -440 970
rect -420 950 -415 970
rect -445 920 -415 950
rect -445 900 -440 920
rect -420 900 -415 920
rect -445 870 -415 900
rect -445 850 -440 870
rect -420 850 -415 870
rect -445 840 -415 850
rect -390 1420 -320 1430
rect 275 1420 315 1430
rect 385 1450 425 1460
rect 385 1430 395 1450
rect 415 1430 425 1450
rect 385 1420 425 1430
rect 495 1450 535 1460
rect 495 1430 505 1450
rect 525 1430 535 1450
rect 495 1420 535 1430
rect 605 1450 645 1460
rect 605 1430 615 1450
rect 635 1430 645 1450
rect 605 1420 645 1430
rect 715 1450 755 1460
rect 715 1430 725 1450
rect 745 1430 755 1450
rect 715 1420 755 1430
rect 825 1450 865 1460
rect 825 1430 835 1450
rect 855 1430 865 1450
rect 825 1420 865 1430
rect 885 1450 915 1460
rect 885 1430 890 1450
rect 910 1430 915 1450
rect 885 1420 915 1430
rect 935 1450 975 1460
rect 935 1430 945 1450
rect 965 1430 975 1450
rect 935 1420 975 1430
rect 1045 1450 1085 1460
rect 1045 1430 1055 1450
rect 1075 1430 1085 1450
rect 1045 1420 1085 1430
rect 1155 1450 1195 1460
rect 1155 1430 1165 1450
rect 1185 1430 1195 1450
rect 1155 1420 1195 1430
rect 1265 1450 1305 1460
rect 1265 1430 1275 1450
rect 1295 1430 1305 1450
rect 1265 1420 1305 1430
rect 1375 1450 1415 1460
rect 2045 1450 2085 1460
rect 2155 1480 2195 1490
rect 2155 1460 2165 1480
rect 2185 1460 2195 1480
rect 2155 1450 2195 1460
rect 2265 1480 2305 1490
rect 2265 1460 2275 1480
rect 2295 1460 2305 1480
rect 2265 1450 2305 1460
rect 2375 1480 2415 1490
rect 2375 1460 2385 1480
rect 2405 1460 2415 1480
rect 2375 1450 2415 1460
rect 2485 1480 2525 1490
rect 2485 1460 2495 1480
rect 2515 1460 2525 1480
rect 2485 1450 2525 1460
rect 2595 1480 2635 1490
rect 2595 1460 2605 1480
rect 2625 1460 2635 1480
rect 2595 1450 2635 1460
rect 2705 1480 2745 1490
rect 2705 1460 2715 1480
rect 2735 1460 2745 1480
rect 2705 1450 2745 1460
rect 1375 1430 1385 1450
rect 1405 1430 1415 1450
rect 2055 1430 2075 1450
rect 2165 1430 2185 1450
rect 2275 1430 2295 1450
rect 2385 1430 2405 1450
rect 2495 1430 2515 1450
rect 2605 1430 2625 1450
rect 2715 1430 2735 1450
rect 1375 1420 1415 1430
rect 2010 1420 2080 1430
rect -390 1400 -385 1420
rect -365 1400 -345 1420
rect -325 1400 -320 1420
rect -390 1370 -320 1400
rect -390 1350 -385 1370
rect -365 1350 -345 1370
rect -325 1350 -320 1370
rect -390 1320 -320 1350
rect -390 1300 -385 1320
rect -365 1300 -345 1320
rect -325 1300 -320 1320
rect -390 1270 -320 1300
rect -390 1250 -385 1270
rect -365 1250 -345 1270
rect -325 1250 -320 1270
rect 2010 1400 2015 1420
rect 2035 1400 2055 1420
rect 2075 1400 2080 1420
rect 2010 1370 2080 1400
rect 2010 1350 2015 1370
rect 2035 1350 2055 1370
rect 2075 1350 2080 1370
rect 2010 1320 2080 1350
rect 2010 1300 2015 1320
rect 2035 1300 2055 1320
rect 2075 1300 2080 1320
rect 2010 1270 2080 1300
rect -390 1220 -320 1250
rect 71 1250 101 1260
rect 71 1230 76 1250
rect 96 1230 101 1250
rect 71 1220 101 1230
rect 120 1250 150 1260
rect 120 1230 125 1250
rect 145 1230 150 1250
rect 120 1220 150 1230
rect 220 1250 250 1260
rect 220 1230 225 1250
rect 245 1230 250 1250
rect 220 1220 250 1230
rect 275 1250 305 1260
rect 275 1230 280 1250
rect 300 1230 305 1250
rect 275 1220 305 1230
rect 330 1250 360 1260
rect 330 1230 335 1250
rect 355 1230 360 1250
rect 330 1220 360 1230
rect 440 1250 470 1260
rect 440 1230 445 1250
rect 465 1230 470 1250
rect 440 1220 470 1230
rect 495 1250 525 1260
rect 495 1230 500 1250
rect 520 1230 525 1250
rect 495 1220 525 1230
rect 550 1250 580 1260
rect 550 1230 555 1250
rect 575 1230 580 1250
rect 550 1220 580 1230
rect 1071 1250 1101 1260
rect 1071 1230 1076 1250
rect 1096 1230 1101 1250
rect 1071 1220 1101 1230
rect 1120 1250 1150 1260
rect 1120 1230 1125 1250
rect 1145 1230 1150 1250
rect 1120 1220 1150 1230
rect 1220 1250 1250 1260
rect 1220 1230 1225 1250
rect 1245 1230 1250 1250
rect 1220 1220 1250 1230
rect 1275 1250 1305 1260
rect 1275 1230 1280 1250
rect 1300 1230 1305 1250
rect 1275 1220 1305 1230
rect 1330 1250 1360 1260
rect 1330 1230 1335 1250
rect 1355 1230 1360 1250
rect 1330 1220 1360 1230
rect 1440 1250 1470 1260
rect 1440 1230 1445 1250
rect 1465 1230 1470 1250
rect 1440 1220 1470 1230
rect 1495 1250 1525 1260
rect 1495 1230 1500 1250
rect 1520 1230 1525 1250
rect 1495 1220 1525 1230
rect 1550 1250 1580 1260
rect 1550 1230 1555 1250
rect 1575 1230 1580 1250
rect 1550 1220 1580 1230
rect 2010 1250 2015 1270
rect 2035 1250 2055 1270
rect 2075 1250 2080 1270
rect 2010 1220 2080 1250
rect -390 1200 -385 1220
rect -365 1200 -345 1220
rect -325 1200 -320 1220
rect 120 1200 140 1220
rect 225 1200 245 1220
rect 335 1200 355 1220
rect 445 1200 465 1220
rect 555 1200 575 1220
rect 1120 1200 1140 1220
rect 1225 1200 1245 1220
rect 1335 1200 1355 1220
rect 1445 1200 1465 1220
rect 1555 1200 1575 1220
rect 2010 1200 2015 1220
rect 2035 1200 2055 1220
rect 2075 1200 2080 1220
rect -390 1170 -320 1200
rect -390 1150 -385 1170
rect -365 1150 -345 1170
rect -325 1150 -320 1170
rect -45 1190 30 1200
rect -45 1170 -35 1190
rect -15 1170 5 1190
rect 25 1170 30 1190
rect -45 1160 30 1170
rect 55 1190 85 1200
rect 55 1170 60 1190
rect 80 1170 85 1190
rect 55 1160 85 1170
rect 110 1190 140 1200
rect 110 1170 115 1190
rect 135 1170 140 1190
rect 110 1160 140 1170
rect 165 1190 195 1200
rect 165 1170 170 1190
rect 190 1170 195 1190
rect 165 1160 195 1170
rect 220 1190 250 1200
rect 220 1170 225 1190
rect 245 1170 250 1190
rect 220 1160 250 1170
rect 275 1190 305 1200
rect 275 1170 280 1190
rect 300 1170 305 1190
rect 275 1160 305 1170
rect 330 1190 360 1200
rect 330 1170 335 1190
rect 355 1170 360 1190
rect 330 1160 360 1170
rect 385 1190 415 1200
rect 385 1170 390 1190
rect 410 1170 415 1190
rect 385 1160 415 1170
rect 440 1190 470 1200
rect 440 1170 445 1190
rect 465 1170 470 1190
rect 440 1160 470 1170
rect 495 1190 525 1200
rect 495 1170 500 1190
rect 520 1170 525 1190
rect 495 1160 525 1170
rect 550 1190 580 1200
rect 550 1170 555 1190
rect 575 1170 580 1190
rect 550 1160 580 1170
rect 605 1190 635 1200
rect 605 1170 610 1190
rect 630 1170 635 1190
rect 605 1160 635 1170
rect 660 1190 730 1200
rect 660 1170 665 1190
rect 685 1170 705 1190
rect 725 1170 730 1190
rect 660 1160 730 1170
rect 960 1190 1030 1200
rect 960 1170 965 1190
rect 985 1170 1005 1190
rect 1025 1170 1030 1190
rect 960 1160 1030 1170
rect 1055 1190 1085 1200
rect 1055 1170 1060 1190
rect 1080 1170 1085 1190
rect 1055 1160 1085 1170
rect 1110 1190 1140 1200
rect 1110 1170 1115 1190
rect 1135 1170 1140 1190
rect 1110 1160 1140 1170
rect 1165 1190 1195 1200
rect 1165 1170 1170 1190
rect 1190 1170 1195 1190
rect 1165 1160 1195 1170
rect 1220 1190 1250 1200
rect 1220 1170 1225 1190
rect 1245 1170 1250 1190
rect 1220 1160 1250 1170
rect 1275 1190 1305 1200
rect 1275 1170 1280 1190
rect 1300 1170 1305 1190
rect 1275 1160 1305 1170
rect 1330 1190 1360 1200
rect 1330 1170 1335 1190
rect 1355 1170 1360 1190
rect 1330 1160 1360 1170
rect 1385 1190 1415 1200
rect 1385 1170 1390 1190
rect 1410 1170 1415 1190
rect 1385 1160 1415 1170
rect 1440 1190 1470 1200
rect 1440 1170 1445 1190
rect 1465 1170 1470 1190
rect 1440 1160 1470 1170
rect 1495 1190 1525 1200
rect 1495 1170 1500 1190
rect 1520 1170 1525 1190
rect 1495 1160 1525 1170
rect 1550 1190 1580 1200
rect 1550 1170 1555 1190
rect 1575 1170 1580 1190
rect 1550 1160 1580 1170
rect 1605 1190 1635 1200
rect 1605 1170 1610 1190
rect 1630 1170 1635 1190
rect 1605 1160 1635 1170
rect 1660 1190 1735 1200
rect 1660 1170 1665 1190
rect 1685 1170 1705 1190
rect 1725 1170 1735 1190
rect 1660 1160 1735 1170
rect 2010 1170 2080 1200
rect -390 1120 -320 1150
rect -390 1100 -385 1120
rect -365 1100 -345 1120
rect -325 1100 -320 1120
rect -5 1130 25 1160
rect 60 1135 80 1160
rect 165 1135 185 1160
rect -5 1110 0 1130
rect 20 1110 25 1130
rect -5 1100 25 1110
rect 50 1125 90 1135
rect 50 1105 60 1125
rect 80 1105 90 1125
rect -390 1070 -320 1100
rect 50 1095 90 1105
rect 145 1125 185 1135
rect 145 1105 155 1125
rect 175 1105 185 1125
rect 145 1095 185 1105
rect 204 1131 234 1141
rect 280 1135 300 1160
rect 385 1135 405 1160
rect 204 1111 209 1131
rect 229 1111 234 1131
rect 204 1101 234 1111
rect 270 1125 310 1135
rect 270 1105 280 1125
rect 300 1105 310 1125
rect 270 1095 310 1105
rect 365 1125 405 1135
rect 365 1105 375 1125
rect 395 1105 405 1125
rect 365 1095 405 1105
rect 424 1131 454 1141
rect 500 1135 520 1160
rect 424 1111 429 1131
rect 449 1111 454 1131
rect 424 1101 454 1111
rect 490 1125 530 1135
rect 490 1105 500 1125
rect 520 1105 530 1125
rect 490 1095 530 1105
rect 566 1131 596 1141
rect 566 1111 571 1131
rect 591 1111 596 1131
rect 566 1101 596 1111
rect 615 1135 635 1160
rect 615 1125 645 1135
rect 615 1105 620 1125
rect 640 1105 645 1125
rect 615 1095 645 1105
rect 665 1130 695 1160
rect 665 1110 670 1130
rect 690 1110 695 1130
rect 665 1100 695 1110
rect 995 1130 1025 1160
rect 1060 1135 1080 1160
rect 1165 1135 1185 1160
rect 995 1110 1000 1130
rect 1020 1110 1025 1130
rect 995 1100 1025 1110
rect 1050 1125 1090 1135
rect 1050 1105 1060 1125
rect 1080 1105 1090 1125
rect 1050 1095 1090 1105
rect 1145 1125 1185 1135
rect 1145 1105 1155 1125
rect 1175 1105 1185 1125
rect 1145 1095 1185 1105
rect 1204 1131 1234 1141
rect 1280 1135 1300 1160
rect 1385 1135 1405 1160
rect 1204 1111 1209 1131
rect 1229 1111 1234 1131
rect 1204 1101 1234 1111
rect 1270 1125 1310 1135
rect 1270 1105 1280 1125
rect 1300 1105 1310 1125
rect 1270 1095 1310 1105
rect 1365 1125 1405 1135
rect 1365 1105 1375 1125
rect 1395 1105 1405 1125
rect 1365 1095 1405 1105
rect 1424 1131 1454 1141
rect 1500 1135 1520 1160
rect 1424 1111 1429 1131
rect 1449 1111 1454 1131
rect 1424 1101 1454 1111
rect 1490 1125 1530 1135
rect 1490 1105 1500 1125
rect 1520 1105 1530 1125
rect 1490 1095 1530 1105
rect 1566 1131 1596 1141
rect 1566 1111 1571 1131
rect 1591 1111 1596 1131
rect 1566 1101 1596 1111
rect 1615 1135 1635 1160
rect 1615 1125 1645 1135
rect 1615 1105 1620 1125
rect 1640 1105 1645 1125
rect 1615 1095 1645 1105
rect 1665 1130 1695 1160
rect 1665 1110 1670 1130
rect 1690 1110 1695 1130
rect 1665 1100 1695 1110
rect 2010 1150 2015 1170
rect 2035 1150 2055 1170
rect 2075 1150 2080 1170
rect 2010 1120 2080 1150
rect 2010 1100 2015 1120
rect 2035 1100 2055 1120
rect 2075 1100 2080 1120
rect -390 1050 -385 1070
rect -365 1050 -345 1070
rect -325 1050 -320 1070
rect -390 1020 -320 1050
rect -390 1000 -385 1020
rect -365 1000 -345 1020
rect -325 1000 -320 1020
rect -390 970 -320 1000
rect -390 950 -385 970
rect -365 950 -345 970
rect -325 950 -320 970
rect -390 920 -320 950
rect 2010 1070 2080 1100
rect 2010 1050 2015 1070
rect 2035 1050 2055 1070
rect 2075 1050 2080 1070
rect 2010 1020 2080 1050
rect 2010 1000 2015 1020
rect 2035 1000 2055 1020
rect 2075 1000 2080 1020
rect 2010 970 2080 1000
rect 2010 950 2015 970
rect 2035 950 2055 970
rect 2075 950 2080 970
rect -390 900 -385 920
rect -365 900 -345 920
rect -325 900 -320 920
rect -390 870 -320 900
rect 550 925 590 935
rect 550 905 560 925
rect 580 905 590 925
rect 550 895 590 905
rect 660 925 700 935
rect 660 905 670 925
rect 690 905 700 925
rect 660 895 700 905
rect 770 925 810 935
rect 770 905 780 925
rect 800 905 810 925
rect 770 895 810 905
rect 880 925 920 935
rect 880 905 890 925
rect 910 905 920 925
rect 880 895 920 905
rect 990 925 1030 935
rect 990 905 1000 925
rect 1020 905 1030 925
rect 990 895 1030 905
rect 1100 925 1140 935
rect 1100 905 1110 925
rect 1130 905 1140 925
rect 1100 895 1140 905
rect 2010 920 2080 950
rect 2010 900 2015 920
rect 2035 900 2055 920
rect 2075 900 2080 920
rect 560 875 580 895
rect 670 875 690 895
rect 780 875 800 895
rect 890 875 910 895
rect 1000 875 1020 895
rect 1110 875 1130 895
rect -390 850 -385 870
rect -365 850 -345 870
rect -325 850 -320 870
rect -390 840 -320 850
rect 460 865 530 875
rect 460 845 465 865
rect 485 845 505 865
rect 525 845 530 865
rect -1501 815 -1360 825
rect -990 815 -970 840
rect -880 815 -860 840
rect -770 815 -750 840
rect -660 815 -640 840
rect -550 815 -530 840
rect -440 815 -420 840
rect 460 835 530 845
rect 555 865 585 875
rect 555 845 560 865
rect 580 845 585 865
rect 555 835 585 845
rect 610 865 640 875
rect 610 845 615 865
rect 635 845 640 865
rect 610 835 640 845
rect 665 865 695 875
rect 665 845 670 865
rect 690 845 695 865
rect 665 835 695 845
rect 720 865 750 875
rect 720 845 725 865
rect 745 845 750 865
rect 720 835 750 845
rect 775 865 805 875
rect 775 845 780 865
rect 800 845 805 865
rect 775 835 805 845
rect 830 865 860 875
rect 830 845 835 865
rect 855 845 860 865
rect 830 835 860 845
rect 885 865 915 875
rect 885 845 890 865
rect 910 845 915 865
rect 885 835 915 845
rect 940 865 970 875
rect 940 845 945 865
rect 965 845 970 865
rect 940 835 970 845
rect 995 865 1025 875
rect 995 845 1000 865
rect 1020 845 1025 865
rect 995 835 1025 845
rect 1050 865 1080 875
rect 1050 845 1055 865
rect 1075 845 1080 865
rect 1050 835 1080 845
rect 1105 865 1135 875
rect 1105 845 1110 865
rect 1130 845 1135 865
rect 1105 835 1135 845
rect 1160 865 1230 875
rect 1160 845 1165 865
rect 1185 845 1205 865
rect 1225 845 1230 865
rect 1160 835 1230 845
rect 2010 870 2080 900
rect 2010 850 2015 870
rect 2035 850 2055 870
rect 2075 850 2080 870
rect 2010 840 2080 850
rect 2105 1420 2135 1430
rect 2105 1400 2110 1420
rect 2130 1400 2135 1420
rect 2105 1370 2135 1400
rect 2105 1350 2110 1370
rect 2130 1350 2135 1370
rect 2105 1320 2135 1350
rect 2105 1300 2110 1320
rect 2130 1300 2135 1320
rect 2105 1270 2135 1300
rect 2105 1250 2110 1270
rect 2130 1250 2135 1270
rect 2105 1220 2135 1250
rect 2105 1200 2110 1220
rect 2130 1200 2135 1220
rect 2105 1170 2135 1200
rect 2105 1150 2110 1170
rect 2130 1150 2135 1170
rect 2105 1120 2135 1150
rect 2105 1100 2110 1120
rect 2130 1100 2135 1120
rect 2105 1070 2135 1100
rect 2105 1050 2110 1070
rect 2130 1050 2135 1070
rect 2105 1020 2135 1050
rect 2105 1000 2110 1020
rect 2130 1000 2135 1020
rect 2105 970 2135 1000
rect 2105 950 2110 970
rect 2130 950 2135 970
rect 2105 920 2135 950
rect 2105 900 2110 920
rect 2130 900 2135 920
rect 2105 870 2135 900
rect 2105 850 2110 870
rect 2130 850 2135 870
rect 2105 840 2135 850
rect 2160 1420 2190 1430
rect 2160 1400 2165 1420
rect 2185 1400 2190 1420
rect 2160 1370 2190 1400
rect 2160 1350 2165 1370
rect 2185 1350 2190 1370
rect 2160 1320 2190 1350
rect 2160 1300 2165 1320
rect 2185 1300 2190 1320
rect 2160 1270 2190 1300
rect 2160 1250 2165 1270
rect 2185 1250 2190 1270
rect 2160 1220 2190 1250
rect 2160 1200 2165 1220
rect 2185 1200 2190 1220
rect 2160 1170 2190 1200
rect 2160 1150 2165 1170
rect 2185 1150 2190 1170
rect 2160 1120 2190 1150
rect 2160 1100 2165 1120
rect 2185 1100 2190 1120
rect 2160 1070 2190 1100
rect 2160 1050 2165 1070
rect 2185 1050 2190 1070
rect 2160 1020 2190 1050
rect 2160 1000 2165 1020
rect 2185 1000 2190 1020
rect 2160 970 2190 1000
rect 2160 950 2165 970
rect 2185 950 2190 970
rect 2160 920 2190 950
rect 2160 900 2165 920
rect 2185 900 2190 920
rect 2160 870 2190 900
rect 2160 850 2165 870
rect 2185 850 2190 870
rect 2160 840 2190 850
rect 2215 1420 2245 1430
rect 2215 1400 2220 1420
rect 2240 1400 2245 1420
rect 2215 1370 2245 1400
rect 2215 1350 2220 1370
rect 2240 1350 2245 1370
rect 2215 1320 2245 1350
rect 2215 1300 2220 1320
rect 2240 1300 2245 1320
rect 2215 1270 2245 1300
rect 2215 1250 2220 1270
rect 2240 1250 2245 1270
rect 2215 1220 2245 1250
rect 2215 1200 2220 1220
rect 2240 1200 2245 1220
rect 2215 1170 2245 1200
rect 2215 1150 2220 1170
rect 2240 1150 2245 1170
rect 2215 1120 2245 1150
rect 2215 1100 2220 1120
rect 2240 1100 2245 1120
rect 2215 1070 2245 1100
rect 2215 1050 2220 1070
rect 2240 1050 2245 1070
rect 2215 1020 2245 1050
rect 2215 1000 2220 1020
rect 2240 1000 2245 1020
rect 2215 970 2245 1000
rect 2215 950 2220 970
rect 2240 950 2245 970
rect 2215 920 2245 950
rect 2215 900 2220 920
rect 2240 900 2245 920
rect 2215 870 2245 900
rect 2215 850 2220 870
rect 2240 850 2245 870
rect 2215 840 2245 850
rect 2270 1420 2300 1430
rect 2270 1400 2275 1420
rect 2295 1400 2300 1420
rect 2270 1370 2300 1400
rect 2270 1350 2275 1370
rect 2295 1350 2300 1370
rect 2270 1320 2300 1350
rect 2270 1300 2275 1320
rect 2295 1300 2300 1320
rect 2270 1270 2300 1300
rect 2270 1250 2275 1270
rect 2295 1250 2300 1270
rect 2270 1220 2300 1250
rect 2270 1200 2275 1220
rect 2295 1200 2300 1220
rect 2270 1170 2300 1200
rect 2270 1150 2275 1170
rect 2295 1150 2300 1170
rect 2270 1120 2300 1150
rect 2270 1100 2275 1120
rect 2295 1100 2300 1120
rect 2270 1070 2300 1100
rect 2270 1050 2275 1070
rect 2295 1050 2300 1070
rect 2270 1020 2300 1050
rect 2270 1000 2275 1020
rect 2295 1000 2300 1020
rect 2270 970 2300 1000
rect 2270 950 2275 970
rect 2295 950 2300 970
rect 2270 920 2300 950
rect 2270 900 2275 920
rect 2295 900 2300 920
rect 2270 870 2300 900
rect 2270 850 2275 870
rect 2295 850 2300 870
rect 2270 840 2300 850
rect 2325 1420 2355 1430
rect 2325 1400 2330 1420
rect 2350 1400 2355 1420
rect 2325 1370 2355 1400
rect 2325 1350 2330 1370
rect 2350 1350 2355 1370
rect 2325 1320 2355 1350
rect 2325 1300 2330 1320
rect 2350 1300 2355 1320
rect 2325 1270 2355 1300
rect 2325 1250 2330 1270
rect 2350 1250 2355 1270
rect 2325 1220 2355 1250
rect 2325 1200 2330 1220
rect 2350 1200 2355 1220
rect 2325 1170 2355 1200
rect 2325 1150 2330 1170
rect 2350 1150 2355 1170
rect 2325 1120 2355 1150
rect 2325 1100 2330 1120
rect 2350 1100 2355 1120
rect 2325 1070 2355 1100
rect 2325 1050 2330 1070
rect 2350 1050 2355 1070
rect 2325 1020 2355 1050
rect 2325 1000 2330 1020
rect 2350 1000 2355 1020
rect 2325 970 2355 1000
rect 2325 950 2330 970
rect 2350 950 2355 970
rect 2325 920 2355 950
rect 2325 900 2330 920
rect 2350 900 2355 920
rect 2325 870 2355 900
rect 2325 850 2330 870
rect 2350 850 2355 870
rect 2325 840 2355 850
rect 2380 1420 2410 1430
rect 2380 1400 2385 1420
rect 2405 1400 2410 1420
rect 2380 1370 2410 1400
rect 2380 1350 2385 1370
rect 2405 1350 2410 1370
rect 2380 1320 2410 1350
rect 2380 1300 2385 1320
rect 2405 1300 2410 1320
rect 2380 1270 2410 1300
rect 2380 1250 2385 1270
rect 2405 1250 2410 1270
rect 2380 1220 2410 1250
rect 2380 1200 2385 1220
rect 2405 1200 2410 1220
rect 2380 1170 2410 1200
rect 2380 1150 2385 1170
rect 2405 1150 2410 1170
rect 2380 1120 2410 1150
rect 2380 1100 2385 1120
rect 2405 1100 2410 1120
rect 2380 1070 2410 1100
rect 2380 1050 2385 1070
rect 2405 1050 2410 1070
rect 2380 1020 2410 1050
rect 2380 1000 2385 1020
rect 2405 1000 2410 1020
rect 2380 970 2410 1000
rect 2380 950 2385 970
rect 2405 950 2410 970
rect 2380 920 2410 950
rect 2380 900 2385 920
rect 2405 900 2410 920
rect 2380 870 2410 900
rect 2380 850 2385 870
rect 2405 850 2410 870
rect 2380 840 2410 850
rect 2435 1420 2465 1430
rect 2435 1400 2440 1420
rect 2460 1400 2465 1420
rect 2435 1370 2465 1400
rect 2435 1350 2440 1370
rect 2460 1350 2465 1370
rect 2435 1320 2465 1350
rect 2435 1300 2440 1320
rect 2460 1300 2465 1320
rect 2435 1270 2465 1300
rect 2435 1250 2440 1270
rect 2460 1250 2465 1270
rect 2435 1220 2465 1250
rect 2435 1200 2440 1220
rect 2460 1200 2465 1220
rect 2435 1170 2465 1200
rect 2435 1150 2440 1170
rect 2460 1150 2465 1170
rect 2435 1120 2465 1150
rect 2435 1100 2440 1120
rect 2460 1100 2465 1120
rect 2435 1070 2465 1100
rect 2435 1050 2440 1070
rect 2460 1050 2465 1070
rect 2435 1020 2465 1050
rect 2435 1000 2440 1020
rect 2460 1000 2465 1020
rect 2435 970 2465 1000
rect 2435 950 2440 970
rect 2460 950 2465 970
rect 2435 920 2465 950
rect 2435 900 2440 920
rect 2460 900 2465 920
rect 2435 870 2465 900
rect 2435 850 2440 870
rect 2460 850 2465 870
rect 2435 840 2465 850
rect 2490 1420 2520 1430
rect 2490 1400 2495 1420
rect 2515 1400 2520 1420
rect 2490 1370 2520 1400
rect 2490 1350 2495 1370
rect 2515 1350 2520 1370
rect 2490 1320 2520 1350
rect 2490 1300 2495 1320
rect 2515 1300 2520 1320
rect 2490 1270 2520 1300
rect 2490 1250 2495 1270
rect 2515 1250 2520 1270
rect 2490 1220 2520 1250
rect 2490 1200 2495 1220
rect 2515 1200 2520 1220
rect 2490 1170 2520 1200
rect 2490 1150 2495 1170
rect 2515 1150 2520 1170
rect 2490 1120 2520 1150
rect 2490 1100 2495 1120
rect 2515 1100 2520 1120
rect 2490 1070 2520 1100
rect 2490 1050 2495 1070
rect 2515 1050 2520 1070
rect 2490 1020 2520 1050
rect 2490 1000 2495 1020
rect 2515 1000 2520 1020
rect 2490 970 2520 1000
rect 2490 950 2495 970
rect 2515 950 2520 970
rect 2490 920 2520 950
rect 2490 900 2495 920
rect 2515 900 2520 920
rect 2490 870 2520 900
rect 2490 850 2495 870
rect 2515 850 2520 870
rect 2490 840 2520 850
rect 2545 1420 2575 1430
rect 2545 1400 2550 1420
rect 2570 1400 2575 1420
rect 2545 1370 2575 1400
rect 2545 1350 2550 1370
rect 2570 1350 2575 1370
rect 2545 1320 2575 1350
rect 2545 1300 2550 1320
rect 2570 1300 2575 1320
rect 2545 1270 2575 1300
rect 2545 1250 2550 1270
rect 2570 1250 2575 1270
rect 2545 1220 2575 1250
rect 2545 1200 2550 1220
rect 2570 1200 2575 1220
rect 2545 1170 2575 1200
rect 2545 1150 2550 1170
rect 2570 1150 2575 1170
rect 2545 1120 2575 1150
rect 2545 1100 2550 1120
rect 2570 1100 2575 1120
rect 2545 1070 2575 1100
rect 2545 1050 2550 1070
rect 2570 1050 2575 1070
rect 2545 1020 2575 1050
rect 2545 1000 2550 1020
rect 2570 1000 2575 1020
rect 2545 970 2575 1000
rect 2545 950 2550 970
rect 2570 950 2575 970
rect 2545 920 2575 950
rect 2545 900 2550 920
rect 2570 900 2575 920
rect 2545 870 2575 900
rect 2545 850 2550 870
rect 2570 850 2575 870
rect 2545 840 2575 850
rect 2600 1420 2630 1430
rect 2600 1400 2605 1420
rect 2625 1400 2630 1420
rect 2600 1370 2630 1400
rect 2600 1350 2605 1370
rect 2625 1350 2630 1370
rect 2600 1320 2630 1350
rect 2600 1300 2605 1320
rect 2625 1300 2630 1320
rect 2600 1270 2630 1300
rect 2600 1250 2605 1270
rect 2625 1250 2630 1270
rect 2600 1220 2630 1250
rect 2600 1200 2605 1220
rect 2625 1200 2630 1220
rect 2600 1170 2630 1200
rect 2600 1150 2605 1170
rect 2625 1150 2630 1170
rect 2600 1120 2630 1150
rect 2600 1100 2605 1120
rect 2625 1100 2630 1120
rect 2600 1070 2630 1100
rect 2600 1050 2605 1070
rect 2625 1050 2630 1070
rect 2600 1020 2630 1050
rect 2600 1000 2605 1020
rect 2625 1000 2630 1020
rect 2600 970 2630 1000
rect 2600 950 2605 970
rect 2625 950 2630 970
rect 2600 920 2630 950
rect 2600 900 2605 920
rect 2625 900 2630 920
rect 2600 870 2630 900
rect 2600 850 2605 870
rect 2625 850 2630 870
rect 2600 840 2630 850
rect 2655 1420 2685 1430
rect 2655 1400 2660 1420
rect 2680 1400 2685 1420
rect 2655 1370 2685 1400
rect 2655 1350 2660 1370
rect 2680 1350 2685 1370
rect 2655 1320 2685 1350
rect 2655 1300 2660 1320
rect 2680 1300 2685 1320
rect 2655 1270 2685 1300
rect 2655 1250 2660 1270
rect 2680 1250 2685 1270
rect 2655 1220 2685 1250
rect 2655 1200 2660 1220
rect 2680 1200 2685 1220
rect 2655 1170 2685 1200
rect 2655 1150 2660 1170
rect 2680 1150 2685 1170
rect 2655 1120 2685 1150
rect 2655 1100 2660 1120
rect 2680 1100 2685 1120
rect 2655 1070 2685 1100
rect 2655 1050 2660 1070
rect 2680 1050 2685 1070
rect 2655 1020 2685 1050
rect 2655 1000 2660 1020
rect 2680 1000 2685 1020
rect 2655 970 2685 1000
rect 2655 950 2660 970
rect 2680 950 2685 970
rect 2655 920 2685 950
rect 2655 900 2660 920
rect 2680 900 2685 920
rect 2655 870 2685 900
rect 2655 850 2660 870
rect 2680 850 2685 870
rect 2655 840 2685 850
rect 2710 1420 2780 1430
rect 2710 1400 2715 1420
rect 2735 1400 2755 1420
rect 2775 1400 2780 1420
rect 2710 1370 2780 1400
rect 2710 1350 2715 1370
rect 2735 1350 2755 1370
rect 2775 1350 2780 1370
rect 2710 1320 2780 1350
rect 2710 1300 2715 1320
rect 2735 1300 2755 1320
rect 2775 1300 2780 1320
rect 2710 1270 2780 1300
rect 2710 1250 2715 1270
rect 2735 1250 2755 1270
rect 2775 1250 2780 1270
rect 2710 1220 2780 1250
rect 2710 1200 2715 1220
rect 2735 1200 2755 1220
rect 2775 1200 2780 1220
rect 2710 1170 2780 1200
rect 3050 1420 3191 1430
rect 3050 1400 3055 1420
rect 3075 1400 3110 1420
rect 3130 1400 3165 1420
rect 3185 1400 3191 1420
rect 3050 1390 3191 1400
rect 2710 1150 2715 1170
rect 2735 1150 2755 1170
rect 2775 1150 2780 1170
rect 2710 1120 2780 1150
rect 2710 1100 2715 1120
rect 2735 1100 2755 1120
rect 2775 1100 2780 1120
rect 2710 1070 2780 1100
rect 2710 1050 2715 1070
rect 2735 1050 2755 1070
rect 2775 1050 2780 1070
rect 2710 1020 2780 1050
rect 2710 1000 2715 1020
rect 2735 1000 2755 1020
rect 2775 1000 2780 1020
rect 2710 970 2780 1000
rect 2710 950 2715 970
rect 2735 950 2755 970
rect 2775 950 2780 970
rect 2710 920 2780 950
rect 2710 900 2715 920
rect 2735 900 2755 920
rect 2775 900 2780 920
rect 2710 870 2780 900
rect 2710 850 2715 870
rect 2735 850 2755 870
rect 2775 850 2780 870
rect 2710 840 2780 850
rect 505 815 525 835
rect 615 815 635 835
rect 725 815 745 835
rect 835 815 855 835
rect 945 815 965 835
rect 1055 815 1075 835
rect 1165 815 1185 835
rect 2110 815 2130 840
rect 2220 815 2240 840
rect 2330 815 2350 840
rect 2440 815 2460 840
rect 2550 815 2570 840
rect 2660 815 2680 840
rect 3050 815 3191 825
rect -1501 795 -1495 815
rect -1475 795 -1440 815
rect -1420 795 -1385 815
rect -1365 795 -1360 815
rect -1501 785 -1360 795
rect -1000 805 -960 815
rect -1000 785 -990 805
rect -970 785 -960 805
rect -1000 775 -960 785
rect -890 805 -850 815
rect -890 785 -880 805
rect -860 785 -850 805
rect -890 775 -850 785
rect -780 805 -740 815
rect -780 785 -770 805
rect -750 785 -740 805
rect -780 775 -740 785
rect -720 800 -690 810
rect -720 780 -715 800
rect -695 780 -690 800
rect -720 770 -690 780
rect -670 805 -630 815
rect -670 785 -660 805
rect -640 785 -630 805
rect -670 775 -630 785
rect -560 805 -520 815
rect -560 785 -550 805
rect -530 785 -520 805
rect -560 775 -520 785
rect -450 805 -410 815
rect -450 785 -440 805
rect -420 785 -410 805
rect -450 775 -410 785
rect 495 805 535 815
rect 495 785 505 805
rect 525 785 535 805
rect 495 775 535 785
rect 605 805 645 815
rect 605 785 615 805
rect 635 785 645 805
rect 605 775 645 785
rect 715 805 755 815
rect 715 785 725 805
rect 745 785 755 805
rect 715 775 755 785
rect 825 805 865 815
rect 825 785 835 805
rect 855 785 865 805
rect 825 775 865 785
rect 935 805 975 815
rect 935 785 945 805
rect 965 785 975 805
rect 935 775 975 785
rect 1045 805 1085 815
rect 1045 785 1055 805
rect 1075 785 1085 805
rect 1045 775 1085 785
rect 1155 805 1195 815
rect 1155 785 1165 805
rect 1185 785 1195 805
rect 1155 775 1195 785
rect 2100 805 2140 815
rect 2100 785 2110 805
rect 2130 785 2140 805
rect 2100 775 2140 785
rect 2210 805 2250 815
rect 2210 785 2220 805
rect 2240 785 2250 805
rect 2210 775 2250 785
rect 2320 805 2360 815
rect 2320 785 2330 805
rect 2350 785 2360 805
rect 2320 775 2360 785
rect 2380 800 2410 810
rect 2380 780 2385 800
rect 2405 780 2410 800
rect 2380 770 2410 780
rect 2430 805 2470 815
rect 2430 785 2440 805
rect 2460 785 2470 805
rect 2430 775 2470 785
rect 2540 805 2580 815
rect 2540 785 2550 805
rect 2570 785 2580 805
rect 2540 775 2580 785
rect 2650 805 2690 815
rect 2650 785 2660 805
rect 2680 785 2690 805
rect 3050 795 3055 815
rect 3075 795 3110 815
rect 3130 795 3165 815
rect 3185 795 3191 815
rect 3050 785 3191 795
rect 2650 775 2690 785
rect -1065 665 -1025 675
rect -1065 645 -1055 665
rect -1035 645 -1025 665
rect -1065 635 -1025 645
rect -1000 665 -960 675
rect -1000 645 -990 665
rect -970 645 -960 665
rect -1000 635 -960 645
rect -890 665 -850 675
rect -890 645 -880 665
rect -860 645 -850 665
rect -890 635 -850 645
rect -780 665 -740 675
rect -780 645 -770 665
rect -750 645 -740 665
rect -780 635 -740 645
rect -670 665 -630 675
rect -670 645 -660 665
rect -640 645 -630 665
rect -670 635 -630 645
rect -560 665 -520 675
rect -560 645 -550 665
rect -530 645 -520 665
rect -560 635 -520 645
rect -450 665 -410 675
rect -450 645 -440 665
rect -420 645 -410 665
rect -450 635 -410 645
rect -385 665 -345 675
rect 2035 665 2075 675
rect -385 645 -375 665
rect -355 645 -345 665
rect -385 635 -345 645
rect 30 655 70 665
rect 30 635 40 655
rect 60 635 70 655
rect -1045 615 -1025 635
rect -990 615 -970 635
rect -880 615 -860 635
rect -770 615 -750 635
rect -660 615 -640 635
rect -550 615 -530 635
rect -440 615 -420 635
rect -385 615 -365 635
rect 30 625 70 635
rect 140 655 180 665
rect 140 635 150 655
rect 170 635 180 655
rect 140 625 180 635
rect 250 655 290 665
rect 250 635 260 655
rect 280 635 290 655
rect 250 625 290 635
rect 310 655 340 665
rect 310 635 315 655
rect 335 635 340 655
rect 310 625 340 635
rect 360 655 400 665
rect 360 635 370 655
rect 390 635 400 655
rect 360 625 400 635
rect 470 655 510 665
rect 470 635 480 655
rect 500 635 510 655
rect 470 625 510 635
rect 580 655 620 665
rect 580 635 590 655
rect 610 635 620 655
rect 580 625 620 635
rect 1070 655 1110 665
rect 1070 635 1080 655
rect 1100 635 1110 655
rect 1070 625 1110 635
rect 1180 655 1220 665
rect 1180 635 1190 655
rect 1210 635 1220 655
rect 1180 625 1220 635
rect 1290 655 1330 665
rect 1290 635 1300 655
rect 1320 635 1330 655
rect 1290 625 1330 635
rect 1350 655 1380 665
rect 1350 635 1355 655
rect 1375 635 1380 655
rect 1350 625 1380 635
rect 1400 655 1440 665
rect 1400 635 1410 655
rect 1430 635 1440 655
rect 1400 625 1440 635
rect 1510 655 1550 665
rect 1510 635 1520 655
rect 1540 635 1550 655
rect 1510 625 1550 635
rect 1620 655 1660 665
rect 1620 635 1630 655
rect 1650 635 1660 655
rect 2035 645 2045 665
rect 2065 645 2075 665
rect 2035 635 2075 645
rect 2100 665 2140 675
rect 2100 645 2110 665
rect 2130 645 2140 665
rect 2100 635 2140 645
rect 2210 665 2250 675
rect 2210 645 2220 665
rect 2240 645 2250 665
rect 2210 635 2250 645
rect 2320 665 2360 675
rect 2320 645 2330 665
rect 2350 645 2360 665
rect 2320 635 2360 645
rect 2430 665 2470 675
rect 2430 645 2440 665
rect 2460 645 2470 665
rect 2430 635 2470 645
rect 2540 665 2580 675
rect 2540 645 2550 665
rect 2570 645 2580 665
rect 2540 635 2580 645
rect 2650 665 2690 675
rect 2650 645 2660 665
rect 2680 645 2690 665
rect 2650 635 2690 645
rect 2715 665 2755 675
rect 2715 645 2725 665
rect 2745 645 2755 665
rect 2715 635 2755 645
rect 1620 625 1660 635
rect -1090 605 -1020 615
rect -1090 585 -1085 605
rect -1065 585 -1045 605
rect -1025 585 -1020 605
rect -1410 537 -1195 572
rect -1410 517 -1375 537
rect -1230 517 -1195 537
rect -1315 467 -1290 517
rect -1090 555 -1020 585
rect -1090 535 -1085 555
rect -1065 535 -1045 555
rect -1025 535 -1020 555
rect -1090 505 -1020 535
rect -1090 485 -1085 505
rect -1065 485 -1045 505
rect -1025 485 -1020 505
rect -1090 455 -1020 485
rect -1090 435 -1085 455
rect -1065 435 -1045 455
rect -1025 435 -1020 455
rect -1090 425 -1020 435
rect -995 605 -965 615
rect -995 585 -990 605
rect -970 585 -965 605
rect -995 555 -965 585
rect -995 535 -990 555
rect -970 535 -965 555
rect -995 505 -965 535
rect -995 485 -990 505
rect -970 485 -965 505
rect -995 455 -965 485
rect -995 435 -990 455
rect -970 435 -965 455
rect -995 425 -965 435
rect -940 605 -910 615
rect -940 585 -935 605
rect -915 585 -910 605
rect -940 555 -910 585
rect -940 535 -935 555
rect -915 535 -910 555
rect -940 505 -910 535
rect -940 485 -935 505
rect -915 485 -910 505
rect -940 455 -910 485
rect -940 435 -935 455
rect -915 435 -910 455
rect -940 425 -910 435
rect -885 605 -855 615
rect -885 585 -880 605
rect -860 585 -855 605
rect -885 555 -855 585
rect -885 535 -880 555
rect -860 535 -855 555
rect -885 505 -855 535
rect -885 485 -880 505
rect -860 485 -855 505
rect -885 455 -855 485
rect -885 435 -880 455
rect -860 435 -855 455
rect -885 425 -855 435
rect -830 605 -800 615
rect -830 585 -825 605
rect -805 585 -800 605
rect -830 555 -800 585
rect -830 535 -825 555
rect -805 535 -800 555
rect -830 505 -800 535
rect -830 485 -825 505
rect -805 485 -800 505
rect -830 455 -800 485
rect -830 435 -825 455
rect -805 435 -800 455
rect -830 425 -800 435
rect -775 605 -745 615
rect -775 585 -770 605
rect -750 585 -745 605
rect -775 555 -745 585
rect -775 535 -770 555
rect -750 535 -745 555
rect -775 505 -745 535
rect -775 485 -770 505
rect -750 485 -745 505
rect -775 455 -745 485
rect -775 435 -770 455
rect -750 435 -745 455
rect -775 425 -745 435
rect -720 605 -690 615
rect -720 585 -715 605
rect -695 585 -690 605
rect -720 555 -690 585
rect -720 535 -715 555
rect -695 535 -690 555
rect -720 505 -690 535
rect -720 485 -715 505
rect -695 485 -690 505
rect -720 455 -690 485
rect -720 435 -715 455
rect -695 435 -690 455
rect -720 425 -690 435
rect -665 605 -635 615
rect -665 585 -660 605
rect -640 585 -635 605
rect -665 555 -635 585
rect -665 535 -660 555
rect -640 535 -635 555
rect -665 505 -635 535
rect -665 485 -660 505
rect -640 485 -635 505
rect -665 455 -635 485
rect -665 435 -660 455
rect -640 435 -635 455
rect -665 425 -635 435
rect -610 605 -580 615
rect -610 585 -605 605
rect -585 585 -580 605
rect -610 555 -580 585
rect -610 535 -605 555
rect -585 535 -580 555
rect -610 505 -580 535
rect -610 485 -605 505
rect -585 485 -580 505
rect -610 455 -580 485
rect -610 435 -605 455
rect -585 435 -580 455
rect -610 425 -580 435
rect -555 605 -525 615
rect -555 585 -550 605
rect -530 585 -525 605
rect -555 555 -525 585
rect -555 535 -550 555
rect -530 535 -525 555
rect -555 505 -525 535
rect -555 485 -550 505
rect -530 485 -525 505
rect -555 455 -525 485
rect -555 435 -550 455
rect -530 435 -525 455
rect -555 425 -525 435
rect -500 605 -470 615
rect -500 585 -495 605
rect -475 585 -470 605
rect -500 555 -470 585
rect -500 535 -495 555
rect -475 535 -470 555
rect -500 505 -470 535
rect -500 485 -495 505
rect -475 485 -470 505
rect -500 455 -470 485
rect -500 435 -495 455
rect -475 435 -470 455
rect -500 425 -470 435
rect -445 605 -415 615
rect -445 585 -440 605
rect -420 585 -415 605
rect -445 555 -415 585
rect -445 535 -440 555
rect -420 535 -415 555
rect -445 505 -415 535
rect -445 485 -440 505
rect -420 485 -415 505
rect -445 455 -415 485
rect -445 435 -440 455
rect -420 435 -415 455
rect -445 425 -415 435
rect -390 605 -320 615
rect -390 585 -385 605
rect -365 585 -345 605
rect -325 585 -320 605
rect 40 600 60 625
rect 150 600 170 625
rect 260 600 280 625
rect 370 600 390 625
rect 480 600 500 625
rect 590 600 610 625
rect 1080 600 1100 625
rect 1190 600 1210 625
rect 1300 600 1320 625
rect 1410 600 1430 625
rect 1520 600 1540 625
rect 1630 600 1650 625
rect 2055 615 2075 635
rect 2110 615 2130 635
rect 2220 615 2240 635
rect 2330 615 2350 635
rect 2440 615 2460 635
rect 2550 615 2570 635
rect 2660 615 2680 635
rect 2715 615 2735 635
rect 2010 605 2080 615
rect -390 555 -320 585
rect -390 535 -385 555
rect -365 535 -345 555
rect -325 535 -320 555
rect -390 505 -320 535
rect -390 485 -385 505
rect -365 485 -345 505
rect -325 485 -320 505
rect -390 455 -320 485
rect -60 590 10 600
rect -60 570 -55 590
rect -35 570 -15 590
rect 5 570 10 590
rect -60 540 10 570
rect -60 520 -55 540
rect -35 520 -15 540
rect 5 520 10 540
rect -60 490 10 520
rect -60 470 -55 490
rect -35 470 -15 490
rect 5 470 10 490
rect -60 460 10 470
rect 35 590 65 600
rect 35 570 40 590
rect 60 570 65 590
rect 35 540 65 570
rect 35 520 40 540
rect 60 520 65 540
rect 35 490 65 520
rect 35 470 40 490
rect 60 470 65 490
rect 35 460 65 470
rect 90 590 120 600
rect 90 570 95 590
rect 115 570 120 590
rect 90 540 120 570
rect 90 520 95 540
rect 115 520 120 540
rect 90 490 120 520
rect 90 470 95 490
rect 115 470 120 490
rect 90 460 120 470
rect 145 590 175 600
rect 145 570 150 590
rect 170 570 175 590
rect 145 540 175 570
rect 145 520 150 540
rect 170 520 175 540
rect 145 490 175 520
rect 145 470 150 490
rect 170 470 175 490
rect 145 460 175 470
rect 200 590 230 600
rect 200 570 205 590
rect 225 570 230 590
rect 200 540 230 570
rect 200 520 205 540
rect 225 520 230 540
rect 200 490 230 520
rect 200 470 205 490
rect 225 470 230 490
rect 200 460 230 470
rect 255 590 285 600
rect 255 570 260 590
rect 280 570 285 590
rect 255 540 285 570
rect 255 520 260 540
rect 280 520 285 540
rect 255 490 285 520
rect 255 470 260 490
rect 280 470 285 490
rect 255 460 285 470
rect 310 590 340 600
rect 310 570 315 590
rect 335 570 340 590
rect 310 540 340 570
rect 310 520 315 540
rect 335 520 340 540
rect 310 490 340 520
rect 310 470 315 490
rect 335 470 340 490
rect 310 460 340 470
rect 365 590 395 600
rect 365 570 370 590
rect 390 570 395 590
rect 365 540 395 570
rect 365 520 370 540
rect 390 520 395 540
rect 365 490 395 520
rect 365 470 370 490
rect 390 470 395 490
rect 365 460 395 470
rect 420 590 450 600
rect 420 570 425 590
rect 445 570 450 590
rect 420 540 450 570
rect 420 520 425 540
rect 445 520 450 540
rect 420 490 450 520
rect 420 470 425 490
rect 445 470 450 490
rect 420 460 450 470
rect 475 590 505 600
rect 475 570 480 590
rect 500 570 505 590
rect 475 540 505 570
rect 475 520 480 540
rect 500 520 505 540
rect 475 490 505 520
rect 475 470 480 490
rect 500 470 505 490
rect 475 460 505 470
rect 530 590 560 600
rect 530 570 535 590
rect 555 570 560 590
rect 530 540 560 570
rect 530 520 535 540
rect 555 520 560 540
rect 530 490 560 520
rect 530 470 535 490
rect 555 470 560 490
rect 530 460 560 470
rect 585 590 615 600
rect 585 570 590 590
rect 610 570 615 590
rect 585 540 615 570
rect 585 520 590 540
rect 610 520 615 540
rect 585 490 615 520
rect 585 470 590 490
rect 610 470 615 490
rect 585 460 615 470
rect 640 590 710 600
rect 640 570 645 590
rect 665 570 685 590
rect 705 570 710 590
rect 640 540 710 570
rect 640 520 645 540
rect 665 520 685 540
rect 705 520 710 540
rect 640 490 710 520
rect 640 470 645 490
rect 665 470 685 490
rect 705 470 710 490
rect 640 460 710 470
rect 980 590 1050 600
rect 980 570 985 590
rect 1005 570 1025 590
rect 1045 570 1050 590
rect 980 540 1050 570
rect 980 520 985 540
rect 1005 520 1025 540
rect 1045 520 1050 540
rect 980 490 1050 520
rect 980 470 985 490
rect 1005 470 1025 490
rect 1045 470 1050 490
rect 980 460 1050 470
rect 1075 590 1105 600
rect 1075 570 1080 590
rect 1100 570 1105 590
rect 1075 540 1105 570
rect 1075 520 1080 540
rect 1100 520 1105 540
rect 1075 490 1105 520
rect 1075 470 1080 490
rect 1100 470 1105 490
rect 1075 460 1105 470
rect 1130 590 1160 600
rect 1130 570 1135 590
rect 1155 570 1160 590
rect 1130 540 1160 570
rect 1130 520 1135 540
rect 1155 520 1160 540
rect 1130 490 1160 520
rect 1130 470 1135 490
rect 1155 470 1160 490
rect 1130 460 1160 470
rect 1185 590 1215 600
rect 1185 570 1190 590
rect 1210 570 1215 590
rect 1185 540 1215 570
rect 1185 520 1190 540
rect 1210 520 1215 540
rect 1185 490 1215 520
rect 1185 470 1190 490
rect 1210 470 1215 490
rect 1185 460 1215 470
rect 1240 590 1270 600
rect 1240 570 1245 590
rect 1265 570 1270 590
rect 1240 540 1270 570
rect 1240 520 1245 540
rect 1265 520 1270 540
rect 1240 490 1270 520
rect 1240 470 1245 490
rect 1265 470 1270 490
rect 1240 460 1270 470
rect 1295 590 1325 600
rect 1295 570 1300 590
rect 1320 570 1325 590
rect 1295 540 1325 570
rect 1295 520 1300 540
rect 1320 520 1325 540
rect 1295 490 1325 520
rect 1295 470 1300 490
rect 1320 470 1325 490
rect 1295 460 1325 470
rect 1350 590 1380 600
rect 1350 570 1355 590
rect 1375 570 1380 590
rect 1350 540 1380 570
rect 1350 520 1355 540
rect 1375 520 1380 540
rect 1350 490 1380 520
rect 1350 470 1355 490
rect 1375 470 1380 490
rect 1350 460 1380 470
rect 1405 590 1435 600
rect 1405 570 1410 590
rect 1430 570 1435 590
rect 1405 540 1435 570
rect 1405 520 1410 540
rect 1430 520 1435 540
rect 1405 490 1435 520
rect 1405 470 1410 490
rect 1430 470 1435 490
rect 1405 460 1435 470
rect 1460 590 1490 600
rect 1460 570 1465 590
rect 1485 570 1490 590
rect 1460 540 1490 570
rect 1460 520 1465 540
rect 1485 520 1490 540
rect 1460 490 1490 520
rect 1460 470 1465 490
rect 1485 470 1490 490
rect 1460 460 1490 470
rect 1515 590 1545 600
rect 1515 570 1520 590
rect 1540 570 1545 590
rect 1515 540 1545 570
rect 1515 520 1520 540
rect 1540 520 1545 540
rect 1515 490 1545 520
rect 1515 470 1520 490
rect 1540 470 1545 490
rect 1515 460 1545 470
rect 1570 590 1600 600
rect 1570 570 1575 590
rect 1595 570 1600 590
rect 1570 540 1600 570
rect 1570 520 1575 540
rect 1595 520 1600 540
rect 1570 490 1600 520
rect 1570 470 1575 490
rect 1595 470 1600 490
rect 1570 460 1600 470
rect 1625 590 1655 600
rect 1625 570 1630 590
rect 1650 570 1655 590
rect 1625 540 1655 570
rect 1625 520 1630 540
rect 1650 520 1655 540
rect 1625 490 1655 520
rect 1625 470 1630 490
rect 1650 470 1655 490
rect 1625 460 1655 470
rect 1680 590 1750 600
rect 1680 570 1685 590
rect 1705 570 1725 590
rect 1745 570 1750 590
rect 1680 540 1750 570
rect 1680 520 1685 540
rect 1705 520 1725 540
rect 1745 520 1750 540
rect 1680 490 1750 520
rect 1680 470 1685 490
rect 1705 470 1725 490
rect 1745 470 1750 490
rect 1680 460 1750 470
rect 2010 585 2015 605
rect 2035 585 2055 605
rect 2075 585 2080 605
rect 2010 555 2080 585
rect 2010 535 2015 555
rect 2035 535 2055 555
rect 2075 535 2080 555
rect 2010 505 2080 535
rect 2010 485 2015 505
rect 2035 485 2055 505
rect 2075 485 2080 505
rect -390 435 -385 455
rect -365 435 -345 455
rect -325 435 -320 455
rect -15 440 5 460
rect 95 440 115 460
rect 205 440 225 460
rect 315 440 335 460
rect 425 440 445 460
rect 535 440 555 460
rect 645 440 665 460
rect 1025 440 1045 460
rect 1135 440 1155 460
rect 1245 440 1265 460
rect 1355 440 1375 460
rect 1465 440 1485 460
rect 1575 440 1595 460
rect 1685 440 1705 460
rect 2010 455 2080 485
rect -390 425 -320 435
rect -25 430 15 440
rect -935 400 -915 425
rect -825 400 -805 425
rect -715 400 -695 425
rect -605 400 -585 425
rect -495 400 -475 425
rect -25 410 -15 430
rect 5 410 15 430
rect -25 400 15 410
rect 85 430 125 440
rect 85 410 95 430
rect 115 410 125 430
rect 85 400 125 410
rect 195 430 235 440
rect 195 410 205 430
rect 225 410 235 430
rect 195 400 235 410
rect 305 430 345 440
rect 305 410 315 430
rect 335 410 345 430
rect 305 400 345 410
rect 415 430 455 440
rect 415 410 425 430
rect 445 410 455 430
rect 415 400 455 410
rect 525 430 565 440
rect 525 410 535 430
rect 555 410 565 430
rect 525 400 565 410
rect 635 430 675 440
rect 635 410 645 430
rect 665 410 675 430
rect 635 400 675 410
rect 1015 430 1055 440
rect 1015 410 1025 430
rect 1045 410 1055 430
rect 1015 400 1055 410
rect 1125 430 1165 440
rect 1125 410 1135 430
rect 1155 410 1165 430
rect 1125 400 1165 410
rect 1235 430 1275 440
rect 1235 410 1245 430
rect 1265 410 1275 430
rect 1235 400 1275 410
rect 1345 430 1385 440
rect 1345 410 1355 430
rect 1375 410 1385 430
rect 1345 400 1385 410
rect 1455 430 1495 440
rect 1455 410 1465 430
rect 1485 410 1495 430
rect 1455 400 1495 410
rect 1565 430 1605 440
rect 1565 410 1575 430
rect 1595 410 1605 430
rect 1565 400 1605 410
rect 1675 430 1715 440
rect 1675 410 1685 430
rect 1705 410 1715 430
rect 2010 435 2015 455
rect 2035 435 2055 455
rect 2075 435 2080 455
rect 2010 425 2080 435
rect 2105 605 2135 615
rect 2105 585 2110 605
rect 2130 585 2135 605
rect 2105 555 2135 585
rect 2105 535 2110 555
rect 2130 535 2135 555
rect 2105 505 2135 535
rect 2105 485 2110 505
rect 2130 485 2135 505
rect 2105 455 2135 485
rect 2105 435 2110 455
rect 2130 435 2135 455
rect 2105 425 2135 435
rect 2160 605 2190 615
rect 2160 585 2165 605
rect 2185 585 2190 605
rect 2160 555 2190 585
rect 2160 535 2165 555
rect 2185 535 2190 555
rect 2160 505 2190 535
rect 2160 485 2165 505
rect 2185 485 2190 505
rect 2160 455 2190 485
rect 2160 435 2165 455
rect 2185 435 2190 455
rect 2160 425 2190 435
rect 2215 605 2245 615
rect 2215 585 2220 605
rect 2240 585 2245 605
rect 2215 555 2245 585
rect 2215 535 2220 555
rect 2240 535 2245 555
rect 2215 505 2245 535
rect 2215 485 2220 505
rect 2240 485 2245 505
rect 2215 455 2245 485
rect 2215 435 2220 455
rect 2240 435 2245 455
rect 2215 425 2245 435
rect 2270 605 2300 615
rect 2270 585 2275 605
rect 2295 585 2300 605
rect 2270 555 2300 585
rect 2270 535 2275 555
rect 2295 535 2300 555
rect 2270 505 2300 535
rect 2270 485 2275 505
rect 2295 485 2300 505
rect 2270 455 2300 485
rect 2270 435 2275 455
rect 2295 435 2300 455
rect 2270 425 2300 435
rect 2325 605 2355 615
rect 2325 585 2330 605
rect 2350 585 2355 605
rect 2325 555 2355 585
rect 2325 535 2330 555
rect 2350 535 2355 555
rect 2325 505 2355 535
rect 2325 485 2330 505
rect 2350 485 2355 505
rect 2325 455 2355 485
rect 2325 435 2330 455
rect 2350 435 2355 455
rect 2325 425 2355 435
rect 2380 605 2410 615
rect 2380 585 2385 605
rect 2405 585 2410 605
rect 2380 555 2410 585
rect 2380 535 2385 555
rect 2405 535 2410 555
rect 2380 505 2410 535
rect 2380 485 2385 505
rect 2405 485 2410 505
rect 2380 455 2410 485
rect 2380 435 2385 455
rect 2405 435 2410 455
rect 2380 425 2410 435
rect 2435 605 2465 615
rect 2435 585 2440 605
rect 2460 585 2465 605
rect 2435 555 2465 585
rect 2435 535 2440 555
rect 2460 535 2465 555
rect 2435 505 2465 535
rect 2435 485 2440 505
rect 2460 485 2465 505
rect 2435 455 2465 485
rect 2435 435 2440 455
rect 2460 435 2465 455
rect 2435 425 2465 435
rect 2490 605 2520 615
rect 2490 585 2495 605
rect 2515 585 2520 605
rect 2490 555 2520 585
rect 2490 535 2495 555
rect 2515 535 2520 555
rect 2490 505 2520 535
rect 2490 485 2495 505
rect 2515 485 2520 505
rect 2490 455 2520 485
rect 2490 435 2495 455
rect 2515 435 2520 455
rect 2490 425 2520 435
rect 2545 605 2575 615
rect 2545 585 2550 605
rect 2570 585 2575 605
rect 2545 555 2575 585
rect 2545 535 2550 555
rect 2570 535 2575 555
rect 2545 505 2575 535
rect 2545 485 2550 505
rect 2570 485 2575 505
rect 2545 455 2575 485
rect 2545 435 2550 455
rect 2570 435 2575 455
rect 2545 425 2575 435
rect 2600 605 2630 615
rect 2600 585 2605 605
rect 2625 585 2630 605
rect 2600 555 2630 585
rect 2600 535 2605 555
rect 2625 535 2630 555
rect 2600 505 2630 535
rect 2600 485 2605 505
rect 2625 485 2630 505
rect 2600 455 2630 485
rect 2600 435 2605 455
rect 2625 435 2630 455
rect 2600 425 2630 435
rect 2655 605 2685 615
rect 2655 585 2660 605
rect 2680 585 2685 605
rect 2655 555 2685 585
rect 2655 535 2660 555
rect 2680 535 2685 555
rect 2655 505 2685 535
rect 2655 485 2660 505
rect 2680 485 2685 505
rect 2655 455 2685 485
rect 2655 435 2660 455
rect 2680 435 2685 455
rect 2655 425 2685 435
rect 2710 605 2780 615
rect 2710 585 2715 605
rect 2735 585 2755 605
rect 2775 585 2780 605
rect 2710 555 2780 585
rect 2710 535 2715 555
rect 2735 535 2755 555
rect 2775 535 2780 555
rect 2710 505 2780 535
rect 2710 485 2715 505
rect 2735 485 2755 505
rect 2775 485 2780 505
rect 2710 455 2780 485
rect 2710 435 2715 455
rect 2735 435 2755 455
rect 2775 435 2780 455
rect 2710 425 2780 435
rect 2885 537 3100 572
rect 2885 517 2920 537
rect 3065 517 3100 537
rect 1675 400 1715 410
rect 2165 400 2185 425
rect 2275 400 2295 425
rect 2385 400 2405 425
rect 2495 400 2515 425
rect 2605 400 2625 425
rect -945 390 -905 400
rect -945 370 -935 390
rect -915 370 -905 390
rect -945 360 -905 370
rect -835 390 -795 400
rect -835 370 -825 390
rect -805 370 -795 390
rect -835 360 -795 370
rect -725 390 -685 400
rect -725 370 -715 390
rect -695 370 -685 390
rect -725 360 -685 370
rect -665 390 -635 400
rect -665 370 -660 390
rect -640 370 -635 390
rect -665 360 -635 370
rect -615 390 -575 400
rect -615 370 -605 390
rect -585 370 -575 390
rect -615 360 -575 370
rect -505 390 -465 400
rect -505 370 -495 390
rect -475 370 -465 390
rect -505 360 -465 370
rect 2155 390 2195 400
rect 2155 370 2165 390
rect 2185 370 2195 390
rect 2155 360 2195 370
rect 2265 390 2305 400
rect 2265 370 2275 390
rect 2295 370 2305 390
rect 2265 360 2305 370
rect 2325 390 2355 400
rect 2325 370 2330 390
rect 2350 370 2355 390
rect 2325 360 2355 370
rect 2375 390 2415 400
rect 2375 370 2385 390
rect 2405 370 2415 390
rect 2375 360 2415 370
rect 2485 390 2525 400
rect 2485 370 2495 390
rect 2515 370 2525 390
rect 2485 360 2525 370
rect 2595 390 2635 400
rect 2595 370 2605 390
rect 2625 370 2635 390
rect 2595 360 2635 370
rect 2980 467 3005 517
rect -945 280 -905 290
rect -945 260 -935 280
rect -915 260 -905 280
rect -945 250 -905 260
rect -835 280 -795 290
rect -835 260 -825 280
rect -805 260 -795 280
rect -835 250 -795 260
rect -725 280 -685 290
rect -725 260 -715 280
rect -695 260 -685 280
rect -725 250 -685 260
rect -665 280 -635 290
rect -665 260 -660 280
rect -640 260 -635 280
rect -665 250 -635 260
rect -615 280 -575 290
rect -615 260 -605 280
rect -585 260 -575 280
rect -615 250 -575 260
rect -505 280 -465 290
rect -505 260 -495 280
rect -475 260 -465 280
rect -505 250 -465 260
rect 2155 280 2195 290
rect 2155 260 2165 280
rect 2185 260 2195 280
rect 2155 250 2195 260
rect 2265 280 2305 290
rect 2265 260 2275 280
rect 2295 260 2305 280
rect 2265 250 2305 260
rect 2325 280 2355 290
rect 2325 260 2330 280
rect 2350 260 2355 280
rect 2325 250 2355 260
rect 2375 280 2415 290
rect 2375 260 2385 280
rect 2405 260 2415 280
rect 2375 250 2415 260
rect 2485 280 2525 290
rect 2485 260 2495 280
rect 2515 260 2525 280
rect 2485 250 2525 260
rect 2595 280 2635 290
rect 2595 260 2605 280
rect 2625 260 2635 280
rect 2595 250 2635 260
rect -935 225 -915 250
rect -825 225 -805 250
rect -715 225 -695 250
rect -605 225 -585 250
rect -495 225 -475 250
rect 30 225 70 235
rect -1090 215 -1020 225
rect -1090 195 -1085 215
rect -1065 195 -1045 215
rect -1025 195 -1020 215
rect -1090 165 -1020 195
rect -1090 145 -1085 165
rect -1065 145 -1045 165
rect -1025 145 -1020 165
rect -1410 -93 -1375 -85
rect -1410 -113 -1405 -93
rect -1380 -113 -1375 -93
rect -1410 -120 -1375 -113
rect -1350 -93 -1315 -85
rect -1350 -113 -1345 -93
rect -1320 -113 -1315 -93
rect -1350 -120 -1315 -113
rect -1290 -93 -1255 -85
rect -1290 -113 -1285 -93
rect -1260 -113 -1255 -93
rect -1290 -120 -1255 -113
rect -1090 115 -1020 145
rect -1090 95 -1085 115
rect -1065 95 -1045 115
rect -1025 95 -1020 115
rect -1090 65 -1020 95
rect -1090 45 -1085 65
rect -1065 45 -1045 65
rect -1025 45 -1020 65
rect -1090 15 -1020 45
rect -1090 -5 -1085 15
rect -1065 -5 -1045 15
rect -1025 -5 -1020 15
rect -1090 -35 -1020 -5
rect -1090 -55 -1085 -35
rect -1065 -55 -1045 -35
rect -1025 -55 -1020 -35
rect -1090 -65 -1020 -55
rect -995 215 -965 225
rect -995 195 -990 215
rect -970 195 -965 215
rect -995 165 -965 195
rect -995 145 -990 165
rect -970 145 -965 165
rect -995 115 -965 145
rect -995 95 -990 115
rect -970 95 -965 115
rect -995 65 -965 95
rect -995 45 -990 65
rect -970 45 -965 65
rect -995 15 -965 45
rect -995 -5 -990 15
rect -970 -5 -965 15
rect -995 -35 -965 -5
rect -995 -55 -990 -35
rect -970 -55 -965 -35
rect -995 -65 -965 -55
rect -940 215 -910 225
rect -940 195 -935 215
rect -915 195 -910 215
rect -940 165 -910 195
rect -940 145 -935 165
rect -915 145 -910 165
rect -940 115 -910 145
rect -940 95 -935 115
rect -915 95 -910 115
rect -940 65 -910 95
rect -940 45 -935 65
rect -915 45 -910 65
rect -940 15 -910 45
rect -940 -5 -935 15
rect -915 -5 -910 15
rect -940 -35 -910 -5
rect -940 -55 -935 -35
rect -915 -55 -910 -35
rect -940 -65 -910 -55
rect -885 215 -855 225
rect -885 195 -880 215
rect -860 195 -855 215
rect -885 165 -855 195
rect -885 145 -880 165
rect -860 145 -855 165
rect -885 115 -855 145
rect -885 95 -880 115
rect -860 95 -855 115
rect -885 65 -855 95
rect -885 45 -880 65
rect -860 45 -855 65
rect -885 15 -855 45
rect -885 -5 -880 15
rect -860 -5 -855 15
rect -885 -35 -855 -5
rect -885 -55 -880 -35
rect -860 -55 -855 -35
rect -885 -65 -855 -55
rect -830 215 -800 225
rect -830 195 -825 215
rect -805 195 -800 215
rect -830 165 -800 195
rect -830 145 -825 165
rect -805 145 -800 165
rect -830 115 -800 145
rect -830 95 -825 115
rect -805 95 -800 115
rect -830 65 -800 95
rect -830 45 -825 65
rect -805 45 -800 65
rect -830 15 -800 45
rect -830 -5 -825 15
rect -805 -5 -800 15
rect -830 -35 -800 -5
rect -830 -55 -825 -35
rect -805 -55 -800 -35
rect -830 -65 -800 -55
rect -775 215 -745 225
rect -775 195 -770 215
rect -750 195 -745 215
rect -775 165 -745 195
rect -775 145 -770 165
rect -750 145 -745 165
rect -775 115 -745 145
rect -775 95 -770 115
rect -750 95 -745 115
rect -775 65 -745 95
rect -775 45 -770 65
rect -750 45 -745 65
rect -775 15 -745 45
rect -775 -5 -770 15
rect -750 -5 -745 15
rect -775 -35 -745 -5
rect -775 -55 -770 -35
rect -750 -55 -745 -35
rect -775 -65 -745 -55
rect -720 215 -690 225
rect -720 195 -715 215
rect -695 195 -690 215
rect -720 165 -690 195
rect -720 145 -715 165
rect -695 145 -690 165
rect -720 115 -690 145
rect -720 95 -715 115
rect -695 95 -690 115
rect -720 65 -690 95
rect -720 45 -715 65
rect -695 45 -690 65
rect -720 15 -690 45
rect -720 -5 -715 15
rect -695 -5 -690 15
rect -720 -35 -690 -5
rect -720 -55 -715 -35
rect -695 -55 -690 -35
rect -720 -65 -690 -55
rect -665 215 -635 225
rect -665 195 -660 215
rect -640 195 -635 215
rect -665 165 -635 195
rect -665 145 -660 165
rect -640 145 -635 165
rect -665 115 -635 145
rect -665 95 -660 115
rect -640 95 -635 115
rect -665 65 -635 95
rect -665 45 -660 65
rect -640 45 -635 65
rect -665 15 -635 45
rect -665 -5 -660 15
rect -640 -5 -635 15
rect -665 -35 -635 -5
rect -665 -55 -660 -35
rect -640 -55 -635 -35
rect -665 -65 -635 -55
rect -610 215 -580 225
rect -610 195 -605 215
rect -585 195 -580 215
rect -610 165 -580 195
rect -610 145 -605 165
rect -585 145 -580 165
rect -610 115 -580 145
rect -610 95 -605 115
rect -585 95 -580 115
rect -610 65 -580 95
rect -610 45 -605 65
rect -585 45 -580 65
rect -610 15 -580 45
rect -610 -5 -605 15
rect -585 -5 -580 15
rect -610 -35 -580 -5
rect -610 -55 -605 -35
rect -585 -55 -580 -35
rect -610 -65 -580 -55
rect -555 215 -525 225
rect -555 195 -550 215
rect -530 195 -525 215
rect -555 165 -525 195
rect -555 145 -550 165
rect -530 145 -525 165
rect -555 115 -525 145
rect -555 95 -550 115
rect -530 95 -525 115
rect -555 65 -525 95
rect -555 45 -550 65
rect -530 45 -525 65
rect -555 15 -525 45
rect -555 -5 -550 15
rect -530 -5 -525 15
rect -555 -35 -525 -5
rect -555 -55 -550 -35
rect -530 -55 -525 -35
rect -555 -65 -525 -55
rect -500 215 -470 225
rect -500 195 -495 215
rect -475 195 -470 215
rect -500 165 -470 195
rect -500 145 -495 165
rect -475 145 -470 165
rect -500 115 -470 145
rect -500 95 -495 115
rect -475 95 -470 115
rect -500 65 -470 95
rect -500 45 -495 65
rect -475 45 -470 65
rect -500 15 -470 45
rect -500 -5 -495 15
rect -475 -5 -470 15
rect -500 -35 -470 -5
rect -500 -55 -495 -35
rect -475 -55 -470 -35
rect -500 -65 -470 -55
rect -445 215 -415 225
rect -445 195 -440 215
rect -420 195 -415 215
rect -445 165 -415 195
rect -445 145 -440 165
rect -420 145 -415 165
rect -445 115 -415 145
rect -445 95 -440 115
rect -420 95 -415 115
rect -445 65 -415 95
rect -445 45 -440 65
rect -420 45 -415 65
rect -445 15 -415 45
rect -445 -5 -440 15
rect -420 -5 -415 15
rect -445 -35 -415 -5
rect -445 -55 -440 -35
rect -420 -55 -415 -35
rect -445 -65 -415 -55
rect -390 215 -320 225
rect -390 195 -385 215
rect -365 195 -345 215
rect -325 195 -320 215
rect 30 205 40 225
rect 60 205 70 225
rect 30 195 70 205
rect 140 225 180 235
rect 140 205 150 225
rect 170 205 180 225
rect 140 195 180 205
rect 250 225 290 235
rect 250 205 260 225
rect 280 205 290 225
rect 310 205 340 245
rect 360 225 400 235
rect 360 205 370 225
rect 390 205 400 225
rect 250 195 290 205
rect 360 195 400 205
rect 470 225 510 235
rect 470 205 480 225
rect 500 205 510 225
rect 470 195 510 205
rect 580 225 620 235
rect 580 205 590 225
rect 610 205 620 225
rect 580 195 620 205
rect 1070 225 1110 235
rect 1070 205 1080 225
rect 1100 205 1110 225
rect 1070 195 1110 205
rect 1180 225 1220 235
rect 1180 205 1190 225
rect 1210 205 1220 225
rect 1180 195 1220 205
rect 1290 225 1330 235
rect 1290 205 1300 225
rect 1320 205 1330 225
rect 1350 205 1380 245
rect 1400 225 1440 235
rect 1400 205 1410 225
rect 1430 205 1440 225
rect 1290 195 1330 205
rect 1400 195 1440 205
rect 1510 225 1550 235
rect 1510 205 1520 225
rect 1540 205 1550 225
rect 1510 195 1550 205
rect 1620 225 1660 235
rect 2165 225 2185 250
rect 2275 225 2295 250
rect 2385 225 2405 250
rect 2495 225 2515 250
rect 2605 225 2625 250
rect 1620 205 1630 225
rect 1650 205 1660 225
rect 1620 195 1660 205
rect 2010 215 2080 225
rect 2010 195 2015 215
rect 2035 195 2055 215
rect 2075 195 2080 215
rect -390 165 -320 195
rect -390 145 -385 165
rect -365 145 -345 165
rect -325 145 -320 165
rect -390 115 -320 145
rect 40 125 60 195
rect 150 125 170 195
rect 260 125 280 195
rect 310 175 340 185
rect 310 155 315 175
rect 335 155 340 175
rect 310 145 340 155
rect 370 125 390 195
rect 480 125 500 195
rect 590 125 610 195
rect 795 175 825 185
rect 795 155 800 175
rect 820 155 825 175
rect 795 145 825 155
rect 848 175 878 185
rect 848 155 853 175
rect 873 155 878 175
rect 848 145 878 155
rect 895 175 925 185
rect 895 155 900 175
rect 920 155 925 175
rect 895 145 925 155
rect 895 125 915 145
rect 1080 125 1100 195
rect 1190 125 1210 195
rect 1300 125 1320 195
rect 1350 175 1380 185
rect 1350 155 1355 175
rect 1375 155 1380 175
rect 1350 145 1380 155
rect 1410 125 1430 195
rect 1520 125 1540 195
rect 1630 125 1650 195
rect 2010 165 2080 195
rect 2010 145 2015 165
rect 2035 145 2055 165
rect 2075 145 2080 165
rect -390 95 -385 115
rect -365 95 -345 115
rect -325 95 -320 115
rect -390 65 -320 95
rect -390 45 -385 65
rect -365 45 -345 65
rect -325 45 -320 65
rect -390 15 -320 45
rect -390 -5 -385 15
rect -365 -5 -345 15
rect -325 -5 -320 15
rect -390 -35 -320 -5
rect -60 115 10 125
rect -60 95 -55 115
rect -35 95 -15 115
rect 5 95 10 115
rect -60 65 10 95
rect -60 45 -55 65
rect -35 45 -15 65
rect 5 45 10 65
rect -60 15 10 45
rect -60 -5 -55 15
rect -35 -5 -15 15
rect 5 -5 10 15
rect -60 -15 10 -5
rect 35 115 65 125
rect 35 95 40 115
rect 60 95 65 115
rect 35 65 65 95
rect 35 45 40 65
rect 60 45 65 65
rect 35 15 65 45
rect 35 -5 40 15
rect 60 -5 65 15
rect 35 -15 65 -5
rect 90 115 120 125
rect 90 95 95 115
rect 115 95 120 115
rect 90 65 120 95
rect 90 45 95 65
rect 115 45 120 65
rect 90 15 120 45
rect 90 -5 95 15
rect 115 -5 120 15
rect 90 -15 120 -5
rect 145 115 175 125
rect 145 95 150 115
rect 170 95 175 115
rect 145 65 175 95
rect 145 45 150 65
rect 170 45 175 65
rect 145 15 175 45
rect 145 -5 150 15
rect 170 -5 175 15
rect 145 -15 175 -5
rect 200 115 230 125
rect 200 95 205 115
rect 225 95 230 115
rect 200 65 230 95
rect 200 45 205 65
rect 225 45 230 65
rect 200 15 230 45
rect 200 -5 205 15
rect 225 -5 230 15
rect 200 -15 230 -5
rect 255 115 285 125
rect 255 95 260 115
rect 280 95 285 115
rect 255 65 285 95
rect 255 45 260 65
rect 280 45 285 65
rect 255 15 285 45
rect 255 -5 260 15
rect 280 -5 285 15
rect 255 -15 285 -5
rect 310 115 340 125
rect 310 95 315 115
rect 335 95 340 115
rect 310 65 340 95
rect 310 45 315 65
rect 335 45 340 65
rect 310 15 340 45
rect 310 -5 315 15
rect 335 -5 340 15
rect 310 -15 340 -5
rect 365 115 395 125
rect 365 95 370 115
rect 390 95 395 115
rect 365 65 395 95
rect 365 45 370 65
rect 390 45 395 65
rect 365 15 395 45
rect 365 -5 370 15
rect 390 -5 395 15
rect 365 -15 395 -5
rect 420 115 450 125
rect 420 95 425 115
rect 445 95 450 115
rect 420 65 450 95
rect 420 45 425 65
rect 445 45 450 65
rect 420 15 450 45
rect 420 -5 425 15
rect 445 -5 450 15
rect 420 -15 450 -5
rect 475 115 505 125
rect 475 95 480 115
rect 500 95 505 115
rect 475 65 505 95
rect 475 45 480 65
rect 500 45 505 65
rect 475 15 505 45
rect 475 -5 480 15
rect 500 -5 505 15
rect 475 -15 505 -5
rect 530 115 560 125
rect 530 95 535 115
rect 555 95 560 115
rect 530 65 560 95
rect 530 45 535 65
rect 555 45 560 65
rect 530 15 560 45
rect 530 -5 535 15
rect 555 -5 560 15
rect 530 -15 560 -5
rect 585 115 615 125
rect 585 95 590 115
rect 610 95 615 115
rect 585 65 615 95
rect 585 45 590 65
rect 610 45 615 65
rect 585 15 615 45
rect 585 -5 590 15
rect 610 -5 615 15
rect 585 -15 615 -5
rect 640 115 750 125
rect 640 95 645 115
rect 665 95 685 115
rect 705 95 725 115
rect 745 95 750 115
rect 640 65 750 95
rect 640 45 645 65
rect 665 45 685 65
rect 705 45 725 65
rect 745 45 750 65
rect 640 15 750 45
rect 640 -5 645 15
rect 665 -5 685 15
rect 705 -5 725 15
rect 745 -5 750 15
rect 640 -15 750 -5
rect 775 115 805 125
rect 775 95 780 115
rect 800 95 805 115
rect 775 65 805 95
rect 775 45 780 65
rect 800 45 805 65
rect 775 15 805 45
rect 775 -5 780 15
rect 800 -5 805 15
rect 775 -15 805 -5
rect 830 115 860 125
rect 830 95 835 115
rect 855 95 860 115
rect 830 65 860 95
rect 830 45 835 65
rect 855 45 860 65
rect 830 15 860 45
rect 830 -5 835 15
rect 855 -5 860 15
rect 830 -15 860 -5
rect 885 115 915 125
rect 885 95 890 115
rect 910 95 915 115
rect 885 65 915 95
rect 885 45 890 65
rect 910 45 915 65
rect 885 15 915 45
rect 885 -5 890 15
rect 910 -5 915 15
rect 885 -15 915 -5
rect 940 115 1050 125
rect 940 95 945 115
rect 965 95 985 115
rect 1005 95 1025 115
rect 1045 95 1050 115
rect 940 65 1050 95
rect 940 45 945 65
rect 965 45 985 65
rect 1005 45 1025 65
rect 1045 45 1050 65
rect 940 15 1050 45
rect 940 -5 945 15
rect 965 -5 985 15
rect 1005 -5 1025 15
rect 1045 -5 1050 15
rect 940 -15 1050 -5
rect 1075 115 1105 125
rect 1075 95 1080 115
rect 1100 95 1105 115
rect 1075 65 1105 95
rect 1075 45 1080 65
rect 1100 45 1105 65
rect 1075 15 1105 45
rect 1075 -5 1080 15
rect 1100 -5 1105 15
rect 1075 -15 1105 -5
rect 1130 115 1160 125
rect 1130 95 1135 115
rect 1155 95 1160 115
rect 1130 65 1160 95
rect 1130 45 1135 65
rect 1155 45 1160 65
rect 1130 15 1160 45
rect 1130 -5 1135 15
rect 1155 -5 1160 15
rect 1130 -15 1160 -5
rect 1185 115 1215 125
rect 1185 95 1190 115
rect 1210 95 1215 115
rect 1185 65 1215 95
rect 1185 45 1190 65
rect 1210 45 1215 65
rect 1185 15 1215 45
rect 1185 -5 1190 15
rect 1210 -5 1215 15
rect 1185 -15 1215 -5
rect 1240 115 1270 125
rect 1240 95 1245 115
rect 1265 95 1270 115
rect 1240 65 1270 95
rect 1240 45 1245 65
rect 1265 45 1270 65
rect 1240 15 1270 45
rect 1240 -5 1245 15
rect 1265 -5 1270 15
rect 1240 -15 1270 -5
rect 1295 115 1325 125
rect 1295 95 1300 115
rect 1320 95 1325 115
rect 1295 65 1325 95
rect 1295 45 1300 65
rect 1320 45 1325 65
rect 1295 15 1325 45
rect 1295 -5 1300 15
rect 1320 -5 1325 15
rect 1295 -15 1325 -5
rect 1350 115 1380 125
rect 1350 95 1355 115
rect 1375 95 1380 115
rect 1350 65 1380 95
rect 1350 45 1355 65
rect 1375 45 1380 65
rect 1350 15 1380 45
rect 1350 -5 1355 15
rect 1375 -5 1380 15
rect 1350 -15 1380 -5
rect 1405 115 1435 125
rect 1405 95 1410 115
rect 1430 95 1435 115
rect 1405 65 1435 95
rect 1405 45 1410 65
rect 1430 45 1435 65
rect 1405 15 1435 45
rect 1405 -5 1410 15
rect 1430 -5 1435 15
rect 1405 -15 1435 -5
rect 1460 115 1490 125
rect 1460 95 1465 115
rect 1485 95 1490 115
rect 1460 65 1490 95
rect 1460 45 1465 65
rect 1485 45 1490 65
rect 1460 15 1490 45
rect 1460 -5 1465 15
rect 1485 -5 1490 15
rect 1460 -15 1490 -5
rect 1515 115 1545 125
rect 1515 95 1520 115
rect 1540 95 1545 115
rect 1515 65 1545 95
rect 1515 45 1520 65
rect 1540 45 1545 65
rect 1515 15 1545 45
rect 1515 -5 1520 15
rect 1540 -5 1545 15
rect 1515 -15 1545 -5
rect 1570 115 1600 125
rect 1570 95 1575 115
rect 1595 95 1600 115
rect 1570 65 1600 95
rect 1570 45 1575 65
rect 1595 45 1600 65
rect 1570 15 1600 45
rect 1570 -5 1575 15
rect 1595 -5 1600 15
rect 1570 -15 1600 -5
rect 1625 115 1655 125
rect 1625 95 1630 115
rect 1650 95 1655 115
rect 1625 65 1655 95
rect 1625 45 1630 65
rect 1650 45 1655 65
rect 1625 15 1655 45
rect 1625 -5 1630 15
rect 1650 -5 1655 15
rect 1625 -15 1655 -5
rect 1680 115 1755 125
rect 1680 95 1685 115
rect 1705 95 1725 115
rect 1745 95 1755 115
rect 1680 65 1755 95
rect 1680 45 1685 65
rect 1705 45 1725 65
rect 1745 45 1755 65
rect 1680 15 1755 45
rect 1680 -5 1685 15
rect 1705 -5 1725 15
rect 1745 -5 1755 15
rect 1680 -15 1755 -5
rect 2010 115 2080 145
rect 2010 95 2015 115
rect 2035 95 2055 115
rect 2075 95 2080 115
rect 2010 65 2080 95
rect 2010 45 2015 65
rect 2035 45 2055 65
rect 2075 45 2080 65
rect 2010 15 2080 45
rect 2010 -5 2015 15
rect 2035 -5 2055 15
rect 2075 -5 2080 15
rect -15 -35 5 -15
rect 95 -35 115 -15
rect 205 -35 225 -15
rect 315 -35 335 -15
rect 425 -35 445 -15
rect 535 -35 555 -15
rect 685 -35 705 -15
rect 780 -35 800 -15
rect 835 -35 855 -15
rect 890 -35 910 -15
rect 985 -35 1005 -15
rect 1135 -35 1155 -15
rect 1245 -35 1265 -15
rect 1355 -35 1375 -15
rect 1465 -35 1485 -15
rect 1575 -35 1595 -15
rect 1685 -35 1705 -15
rect 2010 -35 2080 -5
rect -390 -55 -385 -35
rect -365 -55 -345 -35
rect -325 -55 -320 -35
rect -390 -65 -320 -55
rect -20 -45 10 -35
rect -20 -65 -15 -45
rect 5 -65 10 -45
rect -1045 -85 -1025 -65
rect -990 -85 -970 -65
rect -880 -85 -860 -65
rect -770 -85 -750 -65
rect -660 -85 -640 -65
rect -550 -85 -530 -65
rect -440 -85 -420 -65
rect -385 -85 -365 -65
rect -20 -75 10 -65
rect 85 -45 125 -35
rect 85 -65 95 -45
rect 115 -65 125 -45
rect 85 -75 125 -65
rect 195 -45 235 -35
rect 195 -65 205 -45
rect 225 -65 235 -45
rect 195 -75 235 -65
rect 305 -45 345 -35
rect 305 -65 315 -45
rect 335 -65 345 -45
rect 305 -75 345 -65
rect 415 -45 455 -35
rect 415 -65 425 -45
rect 445 -65 455 -45
rect 415 -75 455 -65
rect 525 -45 565 -35
rect 525 -65 535 -45
rect 555 -65 565 -45
rect 525 -75 565 -65
rect 680 -45 710 -35
rect 680 -65 685 -45
rect 705 -65 710 -45
rect 680 -75 710 -65
rect 775 -45 805 -35
rect 775 -65 780 -45
rect 800 -65 805 -45
rect 775 -75 805 -65
rect 830 -45 860 -35
rect 830 -65 835 -45
rect 855 -65 860 -45
rect 830 -75 860 -65
rect 885 -45 915 -35
rect 885 -65 890 -45
rect 910 -65 915 -45
rect 885 -75 915 -65
rect 980 -45 1010 -35
rect 980 -65 985 -45
rect 1005 -65 1010 -45
rect 980 -75 1010 -65
rect 1125 -45 1165 -35
rect 1125 -65 1135 -45
rect 1155 -65 1165 -45
rect 1125 -75 1165 -65
rect 1235 -45 1275 -35
rect 1235 -65 1245 -45
rect 1265 -65 1275 -45
rect 1235 -75 1275 -65
rect 1345 -45 1385 -35
rect 1345 -65 1355 -45
rect 1375 -65 1385 -45
rect 1345 -75 1385 -65
rect 1455 -45 1495 -35
rect 1455 -65 1465 -45
rect 1485 -65 1495 -45
rect 1455 -75 1495 -65
rect 1565 -45 1605 -35
rect 1565 -65 1575 -45
rect 1595 -65 1605 -45
rect 1565 -75 1605 -65
rect 1680 -45 1710 -35
rect 1680 -65 1685 -45
rect 1705 -65 1710 -45
rect 2010 -55 2015 -35
rect 2035 -55 2055 -35
rect 2075 -55 2080 -35
rect 2010 -65 2080 -55
rect 2105 215 2135 225
rect 2105 195 2110 215
rect 2130 195 2135 215
rect 2105 165 2135 195
rect 2105 145 2110 165
rect 2130 145 2135 165
rect 2105 115 2135 145
rect 2105 95 2110 115
rect 2130 95 2135 115
rect 2105 65 2135 95
rect 2105 45 2110 65
rect 2130 45 2135 65
rect 2105 15 2135 45
rect 2105 -5 2110 15
rect 2130 -5 2135 15
rect 2105 -35 2135 -5
rect 2105 -55 2110 -35
rect 2130 -55 2135 -35
rect 2105 -65 2135 -55
rect 2160 215 2190 225
rect 2160 195 2165 215
rect 2185 195 2190 215
rect 2160 165 2190 195
rect 2160 145 2165 165
rect 2185 145 2190 165
rect 2160 115 2190 145
rect 2160 95 2165 115
rect 2185 95 2190 115
rect 2160 65 2190 95
rect 2160 45 2165 65
rect 2185 45 2190 65
rect 2160 15 2190 45
rect 2160 -5 2165 15
rect 2185 -5 2190 15
rect 2160 -35 2190 -5
rect 2160 -55 2165 -35
rect 2185 -55 2190 -35
rect 2160 -65 2190 -55
rect 2215 215 2245 225
rect 2215 195 2220 215
rect 2240 195 2245 215
rect 2215 165 2245 195
rect 2215 145 2220 165
rect 2240 145 2245 165
rect 2215 115 2245 145
rect 2215 95 2220 115
rect 2240 95 2245 115
rect 2215 65 2245 95
rect 2215 45 2220 65
rect 2240 45 2245 65
rect 2215 15 2245 45
rect 2215 -5 2220 15
rect 2240 -5 2245 15
rect 2215 -35 2245 -5
rect 2215 -55 2220 -35
rect 2240 -55 2245 -35
rect 2215 -65 2245 -55
rect 2270 215 2300 225
rect 2270 195 2275 215
rect 2295 195 2300 215
rect 2270 165 2300 195
rect 2270 145 2275 165
rect 2295 145 2300 165
rect 2270 115 2300 145
rect 2270 95 2275 115
rect 2295 95 2300 115
rect 2270 65 2300 95
rect 2270 45 2275 65
rect 2295 45 2300 65
rect 2270 15 2300 45
rect 2270 -5 2275 15
rect 2295 -5 2300 15
rect 2270 -35 2300 -5
rect 2270 -55 2275 -35
rect 2295 -55 2300 -35
rect 2270 -65 2300 -55
rect 2325 215 2355 225
rect 2325 195 2330 215
rect 2350 195 2355 215
rect 2325 165 2355 195
rect 2325 145 2330 165
rect 2350 145 2355 165
rect 2325 115 2355 145
rect 2325 95 2330 115
rect 2350 95 2355 115
rect 2325 65 2355 95
rect 2325 45 2330 65
rect 2350 45 2355 65
rect 2325 15 2355 45
rect 2325 -5 2330 15
rect 2350 -5 2355 15
rect 2325 -35 2355 -5
rect 2325 -55 2330 -35
rect 2350 -55 2355 -35
rect 2325 -65 2355 -55
rect 2380 215 2410 225
rect 2380 195 2385 215
rect 2405 195 2410 215
rect 2380 165 2410 195
rect 2380 145 2385 165
rect 2405 145 2410 165
rect 2380 115 2410 145
rect 2380 95 2385 115
rect 2405 95 2410 115
rect 2380 65 2410 95
rect 2380 45 2385 65
rect 2405 45 2410 65
rect 2380 15 2410 45
rect 2380 -5 2385 15
rect 2405 -5 2410 15
rect 2380 -35 2410 -5
rect 2380 -55 2385 -35
rect 2405 -55 2410 -35
rect 2380 -65 2410 -55
rect 2435 215 2465 225
rect 2435 195 2440 215
rect 2460 195 2465 215
rect 2435 165 2465 195
rect 2435 145 2440 165
rect 2460 145 2465 165
rect 2435 115 2465 145
rect 2435 95 2440 115
rect 2460 95 2465 115
rect 2435 65 2465 95
rect 2435 45 2440 65
rect 2460 45 2465 65
rect 2435 15 2465 45
rect 2435 -5 2440 15
rect 2460 -5 2465 15
rect 2435 -35 2465 -5
rect 2435 -55 2440 -35
rect 2460 -55 2465 -35
rect 2435 -65 2465 -55
rect 2490 215 2520 225
rect 2490 195 2495 215
rect 2515 195 2520 215
rect 2490 165 2520 195
rect 2490 145 2495 165
rect 2515 145 2520 165
rect 2490 115 2520 145
rect 2490 95 2495 115
rect 2515 95 2520 115
rect 2490 65 2520 95
rect 2490 45 2495 65
rect 2515 45 2520 65
rect 2490 15 2520 45
rect 2490 -5 2495 15
rect 2515 -5 2520 15
rect 2490 -35 2520 -5
rect 2490 -55 2495 -35
rect 2515 -55 2520 -35
rect 2490 -65 2520 -55
rect 2545 215 2575 225
rect 2545 195 2550 215
rect 2570 195 2575 215
rect 2545 165 2575 195
rect 2545 145 2550 165
rect 2570 145 2575 165
rect 2545 115 2575 145
rect 2545 95 2550 115
rect 2570 95 2575 115
rect 2545 65 2575 95
rect 2545 45 2550 65
rect 2570 45 2575 65
rect 2545 15 2575 45
rect 2545 -5 2550 15
rect 2570 -5 2575 15
rect 2545 -35 2575 -5
rect 2545 -55 2550 -35
rect 2570 -55 2575 -35
rect 2545 -65 2575 -55
rect 2600 215 2630 225
rect 2600 195 2605 215
rect 2625 195 2630 215
rect 2600 165 2630 195
rect 2600 145 2605 165
rect 2625 145 2630 165
rect 2600 115 2630 145
rect 2600 95 2605 115
rect 2625 95 2630 115
rect 2600 65 2630 95
rect 2600 45 2605 65
rect 2625 45 2630 65
rect 2600 15 2630 45
rect 2600 -5 2605 15
rect 2625 -5 2630 15
rect 2600 -35 2630 -5
rect 2600 -55 2605 -35
rect 2625 -55 2630 -35
rect 2600 -65 2630 -55
rect 2655 215 2685 225
rect 2655 195 2660 215
rect 2680 195 2685 215
rect 2655 165 2685 195
rect 2655 145 2660 165
rect 2680 145 2685 165
rect 2655 115 2685 145
rect 2655 95 2660 115
rect 2680 95 2685 115
rect 2655 65 2685 95
rect 2655 45 2660 65
rect 2680 45 2685 65
rect 2655 15 2685 45
rect 2655 -5 2660 15
rect 2680 -5 2685 15
rect 2655 -35 2685 -5
rect 2655 -55 2660 -35
rect 2680 -55 2685 -35
rect 2655 -65 2685 -55
rect 2710 215 2780 225
rect 2710 195 2715 215
rect 2735 195 2755 215
rect 2775 195 2780 215
rect 2710 165 2780 195
rect 2710 145 2715 165
rect 2735 145 2755 165
rect 2775 145 2780 165
rect 2710 115 2780 145
rect 2710 95 2715 115
rect 2735 95 2755 115
rect 2775 95 2780 115
rect 2710 65 2780 95
rect 2710 45 2715 65
rect 2735 45 2755 65
rect 2775 45 2780 65
rect 2710 15 2780 45
rect 2710 -5 2715 15
rect 2735 -5 2755 15
rect 2775 -5 2780 15
rect 2710 -35 2780 -5
rect 2710 -55 2715 -35
rect 2735 -55 2755 -35
rect 2775 -55 2780 -35
rect 2710 -65 2780 -55
rect 1680 -75 1710 -65
rect 2055 -85 2075 -65
rect 2110 -85 2130 -65
rect 2220 -85 2240 -65
rect 2330 -85 2350 -65
rect 2440 -85 2460 -65
rect 2550 -85 2570 -65
rect 2660 -85 2680 -65
rect 2715 -85 2735 -65
rect -1230 -93 -1195 -85
rect -1230 -113 -1225 -93
rect -1200 -113 -1195 -93
rect -1230 -120 -1195 -113
rect -1065 -95 -1025 -85
rect -1065 -115 -1055 -95
rect -1035 -115 -1025 -95
rect -1065 -125 -1025 -115
rect -1000 -95 -960 -85
rect -1000 -115 -990 -95
rect -970 -115 -960 -95
rect -1000 -125 -960 -115
rect -890 -95 -850 -85
rect -890 -115 -880 -95
rect -860 -115 -850 -95
rect -890 -125 -850 -115
rect -780 -95 -740 -85
rect -780 -115 -770 -95
rect -750 -115 -740 -95
rect -780 -125 -740 -115
rect -670 -95 -630 -85
rect -670 -115 -660 -95
rect -640 -115 -630 -95
rect -670 -125 -630 -115
rect -560 -95 -520 -85
rect -560 -115 -550 -95
rect -530 -115 -520 -95
rect -560 -125 -520 -115
rect -450 -95 -410 -85
rect -450 -115 -440 -95
rect -420 -115 -410 -95
rect -450 -125 -410 -115
rect -385 -95 -345 -85
rect -385 -115 -375 -95
rect -355 -115 -345 -95
rect -385 -125 -345 -115
rect 2035 -95 2075 -85
rect 2035 -115 2045 -95
rect 2065 -115 2075 -95
rect 2035 -125 2075 -115
rect 2100 -95 2140 -85
rect 2100 -115 2110 -95
rect 2130 -115 2140 -95
rect 2100 -125 2140 -115
rect 2210 -95 2250 -85
rect 2210 -115 2220 -95
rect 2240 -115 2250 -95
rect 2210 -125 2250 -115
rect 2320 -95 2360 -85
rect 2320 -115 2330 -95
rect 2350 -115 2360 -95
rect 2320 -125 2360 -115
rect 2430 -95 2470 -85
rect 2430 -115 2440 -95
rect 2460 -115 2470 -95
rect 2430 -125 2470 -115
rect 2540 -95 2580 -85
rect 2540 -115 2550 -95
rect 2570 -115 2580 -95
rect 2540 -125 2580 -115
rect 2650 -95 2690 -85
rect 2650 -115 2660 -95
rect 2680 -115 2690 -95
rect 2650 -125 2690 -115
rect 2715 -95 2755 -85
rect 2715 -115 2725 -95
rect 2745 -115 2755 -95
rect 2715 -125 2755 -115
rect 2885 -93 2920 -85
rect 2885 -113 2890 -93
rect 2915 -113 2920 -93
rect 2885 -120 2920 -113
rect 2945 -93 2980 -85
rect 2945 -113 2950 -93
rect 2975 -113 2980 -93
rect 2945 -120 2980 -113
rect 3005 -93 3040 -85
rect 3005 -113 3010 -93
rect 3035 -113 3040 -93
rect 3005 -120 3040 -113
rect 3065 -93 3100 -85
rect 3065 -113 3070 -93
rect 3095 -113 3100 -93
rect 3065 -120 3100 -113
rect -925 -305 -885 -295
rect -925 -325 -915 -305
rect -895 -325 -885 -305
rect -925 -335 -885 -325
rect -725 -305 -685 -295
rect -725 -325 -715 -305
rect -695 -325 -685 -305
rect -725 -335 -685 -325
rect -625 -305 -585 -295
rect -625 -325 -615 -305
rect -595 -325 -585 -305
rect -625 -335 -585 -325
rect -525 -305 -485 -295
rect -525 -325 -515 -305
rect -495 -325 -485 -305
rect -525 -335 -485 -325
rect 2175 -305 2215 -295
rect 2175 -325 2185 -305
rect 2205 -325 2215 -305
rect 2175 -335 2215 -325
rect 2275 -305 2315 -295
rect 2275 -325 2285 -305
rect 2305 -325 2315 -305
rect 2275 -335 2315 -325
rect 2375 -305 2415 -295
rect 2375 -325 2385 -305
rect 2405 -325 2415 -305
rect 2375 -335 2415 -325
rect 2575 -305 2615 -295
rect 2575 -325 2585 -305
rect 2605 -325 2615 -305
rect 2575 -335 2615 -325
rect -915 -360 -895 -335
rect -715 -360 -695 -335
rect -515 -360 -495 -335
rect 270 -355 310 -345
rect -1060 -370 -990 -360
rect -1210 -387 -1175 -380
rect -1210 -407 -1205 -387
rect -1180 -407 -1175 -387
rect -1210 -415 -1175 -407
rect -1150 -387 -1115 -380
rect -1150 -407 -1145 -387
rect -1120 -407 -1115 -387
rect -1150 -415 -1115 -407
rect -1060 -390 -1055 -370
rect -1035 -390 -1015 -370
rect -995 -390 -990 -370
rect -1060 -420 -990 -390
rect -1060 -440 -1055 -420
rect -1035 -440 -1015 -420
rect -995 -440 -990 -420
rect -1060 -470 -990 -440
rect -1060 -490 -1055 -470
rect -1035 -490 -1015 -470
rect -995 -490 -990 -470
rect -1060 -520 -990 -490
rect -1060 -540 -1055 -520
rect -1035 -540 -1015 -520
rect -995 -540 -990 -520
rect -1060 -570 -990 -540
rect -1060 -590 -1055 -570
rect -1035 -590 -1015 -570
rect -995 -590 -990 -570
rect -1060 -620 -990 -590
rect -1060 -640 -1055 -620
rect -1035 -640 -1015 -620
rect -995 -640 -990 -620
rect -1060 -670 -990 -640
rect -1060 -690 -1055 -670
rect -1035 -690 -1015 -670
rect -995 -690 -990 -670
rect -1060 -720 -990 -690
rect -1060 -740 -1055 -720
rect -1035 -740 -1015 -720
rect -995 -740 -990 -720
rect -1060 -770 -990 -740
rect -1060 -790 -1055 -770
rect -1035 -790 -1015 -770
rect -995 -790 -990 -770
rect -1060 -820 -990 -790
rect -1060 -840 -1055 -820
rect -1035 -840 -1015 -820
rect -995 -840 -990 -820
rect -1060 -870 -990 -840
rect -1175 -1105 -1150 -1055
rect -1060 -890 -1055 -870
rect -1035 -890 -1015 -870
rect -995 -890 -990 -870
rect -1060 -920 -990 -890
rect -1060 -940 -1055 -920
rect -1035 -940 -1015 -920
rect -995 -940 -990 -920
rect -1060 -970 -990 -940
rect -1060 -990 -1055 -970
rect -1035 -990 -1015 -970
rect -995 -990 -990 -970
rect -1060 -1020 -990 -990
rect -1060 -1040 -1055 -1020
rect -1035 -1040 -1015 -1020
rect -995 -1040 -990 -1020
rect -1060 -1050 -990 -1040
rect -920 -370 -890 -360
rect -920 -390 -915 -370
rect -895 -390 -890 -370
rect -920 -420 -890 -390
rect -920 -440 -915 -420
rect -895 -440 -890 -420
rect -920 -470 -890 -440
rect -920 -490 -915 -470
rect -895 -490 -890 -470
rect -920 -520 -890 -490
rect -920 -540 -915 -520
rect -895 -540 -890 -520
rect -920 -570 -890 -540
rect -920 -590 -915 -570
rect -895 -590 -890 -570
rect -920 -620 -890 -590
rect -920 -640 -915 -620
rect -895 -640 -890 -620
rect -920 -670 -890 -640
rect -920 -690 -915 -670
rect -895 -690 -890 -670
rect -920 -720 -890 -690
rect -920 -740 -915 -720
rect -895 -740 -890 -720
rect -920 -770 -890 -740
rect -920 -790 -915 -770
rect -895 -790 -890 -770
rect -920 -820 -890 -790
rect -920 -840 -915 -820
rect -895 -840 -890 -820
rect -920 -870 -890 -840
rect -920 -890 -915 -870
rect -895 -890 -890 -870
rect -920 -920 -890 -890
rect -920 -940 -915 -920
rect -895 -940 -890 -920
rect -920 -970 -890 -940
rect -920 -990 -915 -970
rect -895 -990 -890 -970
rect -920 -1020 -890 -990
rect -920 -1040 -915 -1020
rect -895 -1040 -890 -1020
rect -920 -1050 -890 -1040
rect -820 -370 -790 -360
rect -820 -390 -815 -370
rect -795 -390 -790 -370
rect -820 -420 -790 -390
rect -820 -440 -815 -420
rect -795 -440 -790 -420
rect -820 -470 -790 -440
rect -820 -490 -815 -470
rect -795 -490 -790 -470
rect -820 -520 -790 -490
rect -820 -540 -815 -520
rect -795 -540 -790 -520
rect -820 -570 -790 -540
rect -820 -590 -815 -570
rect -795 -590 -790 -570
rect -820 -620 -790 -590
rect -820 -640 -815 -620
rect -795 -640 -790 -620
rect -820 -670 -790 -640
rect -820 -690 -815 -670
rect -795 -690 -790 -670
rect -820 -720 -790 -690
rect -820 -740 -815 -720
rect -795 -740 -790 -720
rect -820 -770 -790 -740
rect -820 -790 -815 -770
rect -795 -790 -790 -770
rect -820 -820 -790 -790
rect -820 -840 -815 -820
rect -795 -840 -790 -820
rect -820 -870 -790 -840
rect -820 -890 -815 -870
rect -795 -890 -790 -870
rect -820 -920 -790 -890
rect -820 -940 -815 -920
rect -795 -940 -790 -920
rect -820 -970 -790 -940
rect -820 -990 -815 -970
rect -795 -990 -790 -970
rect -820 -1020 -790 -990
rect -820 -1040 -815 -1020
rect -795 -1040 -790 -1020
rect -820 -1050 -790 -1040
rect -720 -370 -690 -360
rect -720 -390 -715 -370
rect -695 -390 -690 -370
rect -720 -420 -690 -390
rect -720 -440 -715 -420
rect -695 -440 -690 -420
rect -720 -470 -690 -440
rect -720 -490 -715 -470
rect -695 -490 -690 -470
rect -720 -520 -690 -490
rect -720 -540 -715 -520
rect -695 -540 -690 -520
rect -720 -570 -690 -540
rect -720 -590 -715 -570
rect -695 -590 -690 -570
rect -720 -620 -690 -590
rect -720 -640 -715 -620
rect -695 -640 -690 -620
rect -720 -670 -690 -640
rect -720 -690 -715 -670
rect -695 -690 -690 -670
rect -720 -720 -690 -690
rect -720 -740 -715 -720
rect -695 -740 -690 -720
rect -720 -770 -690 -740
rect -720 -790 -715 -770
rect -695 -790 -690 -770
rect -720 -820 -690 -790
rect -720 -840 -715 -820
rect -695 -840 -690 -820
rect -720 -870 -690 -840
rect -720 -890 -715 -870
rect -695 -890 -690 -870
rect -720 -920 -690 -890
rect -720 -940 -715 -920
rect -695 -940 -690 -920
rect -720 -970 -690 -940
rect -720 -990 -715 -970
rect -695 -990 -690 -970
rect -720 -1020 -690 -990
rect -720 -1040 -715 -1020
rect -695 -1040 -690 -1020
rect -720 -1050 -690 -1040
rect -620 -370 -590 -360
rect -620 -390 -615 -370
rect -595 -390 -590 -370
rect -620 -420 -590 -390
rect -620 -440 -615 -420
rect -595 -440 -590 -420
rect -620 -470 -590 -440
rect -620 -490 -615 -470
rect -595 -490 -590 -470
rect -620 -520 -590 -490
rect -620 -540 -615 -520
rect -595 -540 -590 -520
rect -620 -570 -590 -540
rect -620 -590 -615 -570
rect -595 -590 -590 -570
rect -620 -620 -590 -590
rect -620 -640 -615 -620
rect -595 -640 -590 -620
rect -620 -670 -590 -640
rect -620 -690 -615 -670
rect -595 -690 -590 -670
rect -620 -720 -590 -690
rect -620 -740 -615 -720
rect -595 -740 -590 -720
rect -620 -770 -590 -740
rect -620 -790 -615 -770
rect -595 -790 -590 -770
rect -620 -820 -590 -790
rect -620 -840 -615 -820
rect -595 -840 -590 -820
rect -620 -870 -590 -840
rect -620 -890 -615 -870
rect -595 -890 -590 -870
rect -620 -920 -590 -890
rect -620 -940 -615 -920
rect -595 -940 -590 -920
rect -620 -970 -590 -940
rect -620 -990 -615 -970
rect -595 -990 -590 -970
rect -620 -1020 -590 -990
rect -620 -1040 -615 -1020
rect -595 -1040 -590 -1020
rect -620 -1050 -590 -1040
rect -520 -370 -490 -360
rect -520 -390 -515 -370
rect -495 -390 -490 -370
rect -520 -420 -490 -390
rect -520 -440 -515 -420
rect -495 -440 -490 -420
rect -520 -470 -490 -440
rect -520 -490 -515 -470
rect -495 -490 -490 -470
rect -520 -520 -490 -490
rect -520 -540 -515 -520
rect -495 -540 -490 -520
rect -520 -570 -490 -540
rect -520 -590 -515 -570
rect -495 -590 -490 -570
rect -520 -620 -490 -590
rect -520 -640 -515 -620
rect -495 -640 -490 -620
rect -520 -670 -490 -640
rect -520 -690 -515 -670
rect -495 -690 -490 -670
rect -520 -720 -490 -690
rect -520 -740 -515 -720
rect -495 -740 -490 -720
rect -520 -770 -490 -740
rect -520 -790 -515 -770
rect -495 -790 -490 -770
rect -520 -820 -490 -790
rect -520 -840 -515 -820
rect -495 -840 -490 -820
rect -520 -870 -490 -840
rect -520 -890 -515 -870
rect -495 -890 -490 -870
rect -520 -920 -490 -890
rect -520 -940 -515 -920
rect -495 -940 -490 -920
rect -520 -970 -490 -940
rect -520 -990 -515 -970
rect -495 -990 -490 -970
rect -520 -1020 -490 -990
rect -520 -1040 -515 -1020
rect -495 -1040 -490 -1020
rect -520 -1050 -490 -1040
rect -420 -370 -350 -360
rect -420 -390 -415 -370
rect -395 -390 -375 -370
rect -355 -390 -350 -370
rect 270 -375 280 -355
rect 300 -375 310 -355
rect 270 -385 310 -375
rect 380 -355 420 -345
rect 380 -375 390 -355
rect 410 -375 420 -355
rect 380 -385 420 -375
rect 490 -355 530 -345
rect 490 -375 500 -355
rect 520 -375 530 -355
rect 490 -385 530 -375
rect 600 -355 640 -345
rect 600 -375 610 -355
rect 630 -375 640 -355
rect 600 -385 640 -375
rect 710 -355 750 -345
rect 710 -375 720 -355
rect 740 -375 750 -355
rect 710 -385 750 -375
rect 770 -355 800 -345
rect 770 -375 775 -355
rect 795 -375 800 -355
rect 770 -385 800 -375
rect 820 -355 860 -345
rect 820 -375 830 -355
rect 850 -375 860 -355
rect 820 -385 860 -375
rect 930 -355 970 -345
rect 930 -375 940 -355
rect 960 -375 970 -355
rect 930 -385 970 -375
rect 1040 -355 1080 -345
rect 1040 -375 1050 -355
rect 1070 -375 1080 -355
rect 1040 -385 1080 -375
rect 1150 -355 1190 -345
rect 1150 -375 1160 -355
rect 1180 -375 1190 -355
rect 1150 -385 1190 -375
rect 1260 -355 1300 -345
rect 1260 -375 1270 -355
rect 1290 -375 1300 -355
rect 1260 -385 1300 -375
rect 1336 -355 1366 -345
rect 1336 -375 1341 -355
rect 1361 -375 1366 -355
rect 1336 -385 1366 -375
rect 1385 -355 1425 -345
rect 1385 -375 1395 -355
rect 1415 -375 1425 -355
rect 2185 -360 2205 -335
rect 2385 -360 2405 -335
rect 2585 -360 2605 -335
rect 1385 -385 1425 -375
rect 2040 -370 2110 -360
rect -420 -420 -350 -390
rect 280 -410 300 -385
rect 390 -410 410 -385
rect 500 -410 520 -385
rect 610 -410 630 -385
rect 720 -410 740 -385
rect 830 -410 850 -385
rect 940 -410 960 -385
rect 1050 -410 1070 -385
rect 1160 -410 1180 -385
rect 1270 -410 1290 -385
rect 1385 -410 1405 -385
rect 2040 -390 2045 -370
rect 2065 -390 2085 -370
rect 2105 -390 2110 -370
rect -420 -440 -415 -420
rect -395 -440 -375 -420
rect -355 -440 -350 -420
rect -420 -470 -350 -440
rect -420 -490 -415 -470
rect -395 -490 -375 -470
rect -355 -490 -350 -470
rect -420 -520 -350 -490
rect -420 -540 -415 -520
rect -395 -540 -375 -520
rect -355 -540 -350 -520
rect -420 -570 -350 -540
rect -420 -590 -415 -570
rect -395 -590 -375 -570
rect -355 -590 -350 -570
rect -420 -620 -350 -590
rect -420 -640 -415 -620
rect -395 -640 -375 -620
rect -355 -640 -350 -620
rect -420 -670 -350 -640
rect 125 -420 195 -410
rect 125 -440 130 -420
rect 150 -440 170 -420
rect 190 -440 195 -420
rect 125 -470 195 -440
rect 125 -490 130 -470
rect 150 -490 170 -470
rect 190 -490 195 -470
rect 125 -520 195 -490
rect 125 -540 130 -520
rect 150 -540 170 -520
rect 190 -540 195 -520
rect 125 -570 195 -540
rect 125 -590 130 -570
rect 150 -590 170 -570
rect 190 -590 195 -570
rect 125 -620 195 -590
rect 125 -640 130 -620
rect 150 -640 170 -620
rect 190 -640 195 -620
rect 125 -650 195 -640
rect 220 -420 250 -410
rect 220 -440 225 -420
rect 245 -440 250 -420
rect 220 -470 250 -440
rect 220 -490 225 -470
rect 245 -490 250 -470
rect 220 -520 250 -490
rect 220 -540 225 -520
rect 245 -540 250 -520
rect 220 -570 250 -540
rect 220 -590 225 -570
rect 245 -590 250 -570
rect 220 -620 250 -590
rect 220 -640 225 -620
rect 245 -640 250 -620
rect 220 -650 250 -640
rect 275 -420 305 -410
rect 275 -440 280 -420
rect 300 -440 305 -420
rect 275 -470 305 -440
rect 275 -490 280 -470
rect 300 -490 305 -470
rect 275 -520 305 -490
rect 275 -540 280 -520
rect 300 -540 305 -520
rect 275 -570 305 -540
rect 275 -590 280 -570
rect 300 -590 305 -570
rect 275 -620 305 -590
rect 275 -640 280 -620
rect 300 -640 305 -620
rect 275 -650 305 -640
rect 330 -420 360 -410
rect 330 -440 335 -420
rect 355 -440 360 -420
rect 330 -470 360 -440
rect 330 -490 335 -470
rect 355 -490 360 -470
rect 330 -520 360 -490
rect 330 -540 335 -520
rect 355 -540 360 -520
rect 330 -570 360 -540
rect 330 -590 335 -570
rect 355 -590 360 -570
rect 330 -620 360 -590
rect 330 -640 335 -620
rect 355 -640 360 -620
rect 330 -650 360 -640
rect 385 -420 415 -410
rect 385 -440 390 -420
rect 410 -440 415 -420
rect 385 -470 415 -440
rect 385 -490 390 -470
rect 410 -490 415 -470
rect 385 -520 415 -490
rect 385 -540 390 -520
rect 410 -540 415 -520
rect 385 -570 415 -540
rect 385 -590 390 -570
rect 410 -590 415 -570
rect 385 -620 415 -590
rect 385 -640 390 -620
rect 410 -640 415 -620
rect 385 -650 415 -640
rect 440 -420 470 -410
rect 440 -440 445 -420
rect 465 -440 470 -420
rect 440 -470 470 -440
rect 440 -490 445 -470
rect 465 -490 470 -470
rect 440 -520 470 -490
rect 440 -540 445 -520
rect 465 -540 470 -520
rect 440 -570 470 -540
rect 440 -590 445 -570
rect 465 -590 470 -570
rect 440 -620 470 -590
rect 440 -640 445 -620
rect 465 -640 470 -620
rect 440 -650 470 -640
rect 495 -420 525 -410
rect 495 -440 500 -420
rect 520 -440 525 -420
rect 495 -470 525 -440
rect 495 -490 500 -470
rect 520 -490 525 -470
rect 495 -520 525 -490
rect 495 -540 500 -520
rect 520 -540 525 -520
rect 495 -570 525 -540
rect 495 -590 500 -570
rect 520 -590 525 -570
rect 495 -620 525 -590
rect 495 -640 500 -620
rect 520 -640 525 -620
rect 495 -650 525 -640
rect 550 -420 580 -410
rect 550 -440 555 -420
rect 575 -440 580 -420
rect 550 -470 580 -440
rect 550 -490 555 -470
rect 575 -490 580 -470
rect 550 -520 580 -490
rect 550 -540 555 -520
rect 575 -540 580 -520
rect 550 -570 580 -540
rect 550 -590 555 -570
rect 575 -590 580 -570
rect 550 -620 580 -590
rect 550 -640 555 -620
rect 575 -640 580 -620
rect 550 -650 580 -640
rect 605 -420 635 -410
rect 605 -440 610 -420
rect 630 -440 635 -420
rect 605 -470 635 -440
rect 605 -490 610 -470
rect 630 -490 635 -470
rect 605 -520 635 -490
rect 605 -540 610 -520
rect 630 -540 635 -520
rect 605 -570 635 -540
rect 605 -590 610 -570
rect 630 -590 635 -570
rect 605 -620 635 -590
rect 605 -640 610 -620
rect 630 -640 635 -620
rect 605 -650 635 -640
rect 660 -420 690 -410
rect 660 -440 665 -420
rect 685 -440 690 -420
rect 660 -470 690 -440
rect 660 -490 665 -470
rect 685 -490 690 -470
rect 660 -520 690 -490
rect 660 -540 665 -520
rect 685 -540 690 -520
rect 660 -570 690 -540
rect 660 -590 665 -570
rect 685 -590 690 -570
rect 660 -620 690 -590
rect 660 -640 665 -620
rect 685 -640 690 -620
rect 660 -650 690 -640
rect 715 -420 745 -410
rect 715 -440 720 -420
rect 740 -440 745 -420
rect 715 -470 745 -440
rect 715 -490 720 -470
rect 740 -490 745 -470
rect 715 -520 745 -490
rect 715 -540 720 -520
rect 740 -540 745 -520
rect 715 -570 745 -540
rect 715 -590 720 -570
rect 740 -590 745 -570
rect 715 -620 745 -590
rect 715 -640 720 -620
rect 740 -640 745 -620
rect 715 -650 745 -640
rect 770 -420 800 -410
rect 770 -440 775 -420
rect 795 -440 800 -420
rect 770 -470 800 -440
rect 770 -490 775 -470
rect 795 -490 800 -470
rect 770 -520 800 -490
rect 770 -540 775 -520
rect 795 -540 800 -520
rect 770 -570 800 -540
rect 770 -590 775 -570
rect 795 -590 800 -570
rect 770 -620 800 -590
rect 770 -640 775 -620
rect 795 -640 800 -620
rect 770 -650 800 -640
rect 825 -420 855 -410
rect 825 -440 830 -420
rect 850 -440 855 -420
rect 825 -470 855 -440
rect 825 -490 830 -470
rect 850 -490 855 -470
rect 825 -520 855 -490
rect 825 -540 830 -520
rect 850 -540 855 -520
rect 825 -570 855 -540
rect 825 -590 830 -570
rect 850 -590 855 -570
rect 825 -620 855 -590
rect 825 -640 830 -620
rect 850 -640 855 -620
rect 825 -650 855 -640
rect 880 -420 910 -410
rect 880 -440 885 -420
rect 905 -440 910 -420
rect 880 -470 910 -440
rect 880 -490 885 -470
rect 905 -490 910 -470
rect 880 -520 910 -490
rect 880 -540 885 -520
rect 905 -540 910 -520
rect 880 -570 910 -540
rect 880 -590 885 -570
rect 905 -590 910 -570
rect 880 -620 910 -590
rect 880 -640 885 -620
rect 905 -640 910 -620
rect 880 -650 910 -640
rect 935 -420 965 -410
rect 935 -440 940 -420
rect 960 -440 965 -420
rect 935 -470 965 -440
rect 935 -490 940 -470
rect 960 -490 965 -470
rect 935 -520 965 -490
rect 935 -540 940 -520
rect 960 -540 965 -520
rect 935 -570 965 -540
rect 935 -590 940 -570
rect 960 -590 965 -570
rect 935 -620 965 -590
rect 935 -640 940 -620
rect 960 -640 965 -620
rect 935 -650 965 -640
rect 990 -420 1020 -410
rect 990 -440 995 -420
rect 1015 -440 1020 -420
rect 990 -470 1020 -440
rect 990 -490 995 -470
rect 1015 -490 1020 -470
rect 990 -520 1020 -490
rect 990 -540 995 -520
rect 1015 -540 1020 -520
rect 990 -570 1020 -540
rect 990 -590 995 -570
rect 1015 -590 1020 -570
rect 990 -620 1020 -590
rect 990 -640 995 -620
rect 1015 -640 1020 -620
rect 990 -650 1020 -640
rect 1045 -420 1075 -410
rect 1045 -440 1050 -420
rect 1070 -440 1075 -420
rect 1045 -470 1075 -440
rect 1045 -490 1050 -470
rect 1070 -490 1075 -470
rect 1045 -520 1075 -490
rect 1045 -540 1050 -520
rect 1070 -540 1075 -520
rect 1045 -570 1075 -540
rect 1045 -590 1050 -570
rect 1070 -590 1075 -570
rect 1045 -620 1075 -590
rect 1045 -640 1050 -620
rect 1070 -640 1075 -620
rect 1045 -650 1075 -640
rect 1100 -420 1130 -410
rect 1100 -440 1105 -420
rect 1125 -440 1130 -420
rect 1100 -470 1130 -440
rect 1100 -490 1105 -470
rect 1125 -490 1130 -470
rect 1100 -520 1130 -490
rect 1100 -540 1105 -520
rect 1125 -540 1130 -520
rect 1100 -570 1130 -540
rect 1100 -590 1105 -570
rect 1125 -590 1130 -570
rect 1100 -620 1130 -590
rect 1100 -640 1105 -620
rect 1125 -640 1130 -620
rect 1100 -650 1130 -640
rect 1155 -420 1185 -410
rect 1155 -440 1160 -420
rect 1180 -440 1185 -420
rect 1155 -470 1185 -440
rect 1155 -490 1160 -470
rect 1180 -490 1185 -470
rect 1155 -520 1185 -490
rect 1155 -540 1160 -520
rect 1180 -540 1185 -520
rect 1155 -570 1185 -540
rect 1155 -590 1160 -570
rect 1180 -590 1185 -570
rect 1155 -620 1185 -590
rect 1155 -640 1160 -620
rect 1180 -640 1185 -620
rect 1155 -650 1185 -640
rect 1210 -420 1240 -410
rect 1210 -440 1215 -420
rect 1235 -440 1240 -420
rect 1210 -470 1240 -440
rect 1210 -490 1215 -470
rect 1235 -490 1240 -470
rect 1210 -520 1240 -490
rect 1210 -540 1215 -520
rect 1235 -540 1240 -520
rect 1210 -570 1240 -540
rect 1210 -590 1215 -570
rect 1235 -590 1240 -570
rect 1210 -620 1240 -590
rect 1210 -640 1215 -620
rect 1235 -640 1240 -620
rect 1210 -650 1240 -640
rect 1265 -420 1295 -410
rect 1265 -440 1270 -420
rect 1290 -440 1295 -420
rect 1265 -470 1295 -440
rect 1265 -490 1270 -470
rect 1290 -490 1295 -470
rect 1265 -520 1295 -490
rect 1265 -540 1270 -520
rect 1290 -540 1295 -520
rect 1265 -570 1295 -540
rect 1265 -590 1270 -570
rect 1290 -590 1295 -570
rect 1265 -620 1295 -590
rect 1265 -640 1270 -620
rect 1290 -640 1295 -620
rect 1265 -650 1295 -640
rect 1320 -420 1350 -410
rect 1320 -440 1325 -420
rect 1345 -440 1350 -420
rect 1320 -470 1350 -440
rect 1320 -490 1325 -470
rect 1345 -490 1350 -470
rect 1320 -520 1350 -490
rect 1320 -540 1325 -520
rect 1345 -540 1350 -520
rect 1320 -570 1350 -540
rect 1320 -590 1325 -570
rect 1345 -590 1350 -570
rect 1320 -620 1350 -590
rect 1320 -640 1325 -620
rect 1345 -640 1350 -620
rect 1320 -650 1350 -640
rect 1375 -420 1405 -410
rect 1375 -440 1380 -420
rect 1400 -440 1405 -420
rect 1375 -470 1405 -440
rect 1375 -490 1380 -470
rect 1400 -490 1405 -470
rect 1375 -520 1405 -490
rect 1375 -540 1380 -520
rect 1400 -540 1405 -520
rect 1375 -570 1405 -540
rect 1375 -590 1380 -570
rect 1400 -590 1405 -570
rect 1375 -620 1405 -590
rect 1375 -640 1380 -620
rect 1400 -640 1405 -620
rect 1375 -650 1405 -640
rect 1430 -420 1500 -410
rect 1430 -440 1435 -420
rect 1455 -440 1475 -420
rect 1495 -440 1500 -420
rect 1430 -470 1500 -440
rect 1430 -490 1435 -470
rect 1455 -490 1475 -470
rect 1495 -490 1500 -470
rect 1430 -520 1500 -490
rect 1430 -540 1435 -520
rect 1455 -540 1475 -520
rect 1495 -540 1500 -520
rect 1430 -570 1500 -540
rect 1430 -590 1435 -570
rect 1455 -590 1475 -570
rect 1495 -590 1500 -570
rect 1430 -620 1500 -590
rect 1430 -640 1435 -620
rect 1455 -640 1475 -620
rect 1495 -640 1500 -620
rect 1430 -650 1500 -640
rect 2040 -420 2110 -390
rect 2040 -440 2045 -420
rect 2065 -440 2085 -420
rect 2105 -440 2110 -420
rect 2040 -470 2110 -440
rect 2040 -490 2045 -470
rect 2065 -490 2085 -470
rect 2105 -490 2110 -470
rect 2040 -520 2110 -490
rect 2040 -540 2045 -520
rect 2065 -540 2085 -520
rect 2105 -540 2110 -520
rect 2040 -570 2110 -540
rect 2040 -590 2045 -570
rect 2065 -590 2085 -570
rect 2105 -590 2110 -570
rect 2040 -620 2110 -590
rect 2040 -640 2045 -620
rect 2065 -640 2085 -620
rect 2105 -640 2110 -620
rect 170 -670 190 -650
rect 225 -670 245 -650
rect 335 -670 355 -650
rect 445 -670 465 -650
rect 555 -670 575 -650
rect 665 -670 685 -650
rect 775 -670 795 -650
rect 885 -670 905 -650
rect 995 -670 1015 -650
rect 1105 -670 1125 -650
rect 1215 -670 1235 -650
rect 1325 -670 1345 -650
rect 1435 -670 1455 -650
rect 2040 -670 2110 -640
rect -420 -690 -415 -670
rect -395 -690 -375 -670
rect -355 -690 -350 -670
rect -420 -720 -350 -690
rect 150 -680 190 -670
rect 150 -700 160 -680
rect 180 -700 190 -680
rect 150 -710 190 -700
rect 215 -680 255 -670
rect 215 -700 225 -680
rect 245 -700 255 -680
rect 215 -710 255 -700
rect 325 -680 365 -670
rect 325 -700 335 -680
rect 355 -700 365 -680
rect 325 -710 365 -700
rect 435 -680 475 -670
rect 435 -700 445 -680
rect 465 -700 475 -680
rect 435 -710 475 -700
rect 545 -680 585 -670
rect 545 -700 555 -680
rect 575 -700 585 -680
rect 545 -710 585 -700
rect 655 -680 695 -670
rect 655 -700 665 -680
rect 685 -700 695 -680
rect 655 -710 695 -700
rect 765 -680 805 -670
rect 765 -700 775 -680
rect 795 -700 805 -680
rect 765 -710 805 -700
rect 875 -680 915 -670
rect 875 -700 885 -680
rect 905 -700 915 -680
rect 875 -710 915 -700
rect 985 -680 1025 -670
rect 985 -700 995 -680
rect 1015 -700 1025 -680
rect 985 -710 1025 -700
rect 1095 -680 1135 -670
rect 1095 -700 1105 -680
rect 1125 -700 1135 -680
rect 1095 -710 1135 -700
rect 1205 -680 1245 -670
rect 1205 -700 1215 -680
rect 1235 -700 1245 -680
rect 1205 -710 1245 -700
rect 1315 -680 1355 -670
rect 1315 -700 1325 -680
rect 1345 -700 1355 -680
rect 1315 -710 1355 -700
rect 1425 -680 1465 -670
rect 1425 -700 1435 -680
rect 1455 -700 1465 -680
rect 1425 -710 1465 -700
rect 2040 -690 2045 -670
rect 2065 -690 2085 -670
rect 2105 -690 2110 -670
rect -420 -740 -415 -720
rect -395 -740 -375 -720
rect -355 -740 -350 -720
rect 2040 -720 2110 -690
rect -420 -770 -350 -740
rect 1010 -740 1050 -730
rect 1010 -760 1020 -740
rect 1040 -760 1050 -740
rect -420 -790 -415 -770
rect -395 -790 -375 -770
rect -355 -790 -350 -770
rect -420 -820 -350 -790
rect -420 -840 -415 -820
rect -395 -840 -375 -820
rect -355 -840 -350 -820
rect -420 -870 -350 -840
rect -420 -890 -415 -870
rect -395 -890 -375 -870
rect -355 -890 -350 -870
rect -420 -920 -350 -890
rect 670 -775 750 -765
rect 670 -795 720 -775
rect 740 -795 750 -775
rect 670 -805 750 -795
rect 825 -775 865 -765
rect 825 -795 835 -775
rect 855 -795 865 -775
rect 825 -805 865 -795
rect 950 -775 990 -765
rect 950 -795 960 -775
rect 980 -795 990 -775
rect 950 -805 990 -795
rect 1010 -770 1050 -760
rect 2040 -740 2045 -720
rect 2065 -740 2085 -720
rect 2105 -740 2110 -720
rect 2040 -770 2110 -740
rect 670 -835 700 -805
rect 1010 -825 1030 -770
rect 670 -855 675 -835
rect 695 -855 700 -835
rect 670 -885 700 -855
rect 670 -905 675 -885
rect 695 -905 700 -885
rect 670 -915 700 -905
rect 1000 -835 1030 -825
rect 1000 -855 1005 -835
rect 1025 -855 1030 -835
rect 1000 -885 1030 -855
rect 1000 -905 1005 -885
rect 1025 -905 1030 -885
rect 1000 -915 1030 -905
rect 2040 -790 2045 -770
rect 2065 -790 2085 -770
rect 2105 -790 2110 -770
rect 2040 -820 2110 -790
rect 2040 -840 2045 -820
rect 2065 -840 2085 -820
rect 2105 -840 2110 -820
rect 2040 -870 2110 -840
rect 2040 -890 2045 -870
rect 2065 -890 2085 -870
rect 2105 -890 2110 -870
rect -420 -940 -415 -920
rect -395 -940 -375 -920
rect -355 -940 -350 -920
rect -420 -970 -350 -940
rect -420 -990 -415 -970
rect -395 -990 -375 -970
rect -355 -990 -350 -970
rect -420 -1020 -350 -990
rect -420 -1040 -415 -1020
rect -395 -1040 -375 -1020
rect -355 -1040 -350 -1020
rect -420 -1050 -350 -1040
rect 2040 -920 2110 -890
rect 2040 -940 2045 -920
rect 2065 -940 2085 -920
rect 2105 -940 2110 -920
rect 2040 -970 2110 -940
rect 2040 -990 2045 -970
rect 2065 -990 2085 -970
rect 2105 -990 2110 -970
rect 2040 -1020 2110 -990
rect 2040 -1040 2045 -1020
rect 2065 -1040 2085 -1020
rect 2105 -1040 2110 -1020
rect 2040 -1050 2110 -1040
rect 2180 -370 2210 -360
rect 2180 -390 2185 -370
rect 2205 -390 2210 -370
rect 2180 -420 2210 -390
rect 2180 -440 2185 -420
rect 2205 -440 2210 -420
rect 2180 -470 2210 -440
rect 2180 -490 2185 -470
rect 2205 -490 2210 -470
rect 2180 -520 2210 -490
rect 2180 -540 2185 -520
rect 2205 -540 2210 -520
rect 2180 -570 2210 -540
rect 2180 -590 2185 -570
rect 2205 -590 2210 -570
rect 2180 -620 2210 -590
rect 2180 -640 2185 -620
rect 2205 -640 2210 -620
rect 2180 -670 2210 -640
rect 2180 -690 2185 -670
rect 2205 -690 2210 -670
rect 2180 -720 2210 -690
rect 2180 -740 2185 -720
rect 2205 -740 2210 -720
rect 2180 -770 2210 -740
rect 2180 -790 2185 -770
rect 2205 -790 2210 -770
rect 2180 -820 2210 -790
rect 2180 -840 2185 -820
rect 2205 -840 2210 -820
rect 2180 -870 2210 -840
rect 2180 -890 2185 -870
rect 2205 -890 2210 -870
rect 2180 -920 2210 -890
rect 2180 -940 2185 -920
rect 2205 -940 2210 -920
rect 2180 -970 2210 -940
rect 2180 -990 2185 -970
rect 2205 -990 2210 -970
rect 2180 -1020 2210 -990
rect 2180 -1040 2185 -1020
rect 2205 -1040 2210 -1020
rect 2180 -1050 2210 -1040
rect 2280 -370 2310 -360
rect 2280 -390 2285 -370
rect 2305 -390 2310 -370
rect 2280 -420 2310 -390
rect 2280 -440 2285 -420
rect 2305 -440 2310 -420
rect 2280 -470 2310 -440
rect 2280 -490 2285 -470
rect 2305 -490 2310 -470
rect 2280 -520 2310 -490
rect 2280 -540 2285 -520
rect 2305 -540 2310 -520
rect 2280 -570 2310 -540
rect 2280 -590 2285 -570
rect 2305 -590 2310 -570
rect 2280 -620 2310 -590
rect 2280 -640 2285 -620
rect 2305 -640 2310 -620
rect 2280 -670 2310 -640
rect 2280 -690 2285 -670
rect 2305 -690 2310 -670
rect 2280 -720 2310 -690
rect 2280 -740 2285 -720
rect 2305 -740 2310 -720
rect 2280 -770 2310 -740
rect 2280 -790 2285 -770
rect 2305 -790 2310 -770
rect 2280 -820 2310 -790
rect 2280 -840 2285 -820
rect 2305 -840 2310 -820
rect 2280 -870 2310 -840
rect 2280 -890 2285 -870
rect 2305 -890 2310 -870
rect 2280 -920 2310 -890
rect 2280 -940 2285 -920
rect 2305 -940 2310 -920
rect 2280 -970 2310 -940
rect 2280 -990 2285 -970
rect 2305 -990 2310 -970
rect 2280 -1020 2310 -990
rect 2280 -1040 2285 -1020
rect 2305 -1040 2310 -1020
rect 2280 -1050 2310 -1040
rect 2380 -370 2410 -360
rect 2380 -390 2385 -370
rect 2405 -390 2410 -370
rect 2380 -420 2410 -390
rect 2380 -440 2385 -420
rect 2405 -440 2410 -420
rect 2380 -470 2410 -440
rect 2380 -490 2385 -470
rect 2405 -490 2410 -470
rect 2380 -520 2410 -490
rect 2380 -540 2385 -520
rect 2405 -540 2410 -520
rect 2380 -570 2410 -540
rect 2380 -590 2385 -570
rect 2405 -590 2410 -570
rect 2380 -620 2410 -590
rect 2380 -640 2385 -620
rect 2405 -640 2410 -620
rect 2380 -670 2410 -640
rect 2380 -690 2385 -670
rect 2405 -690 2410 -670
rect 2380 -720 2410 -690
rect 2380 -740 2385 -720
rect 2405 -740 2410 -720
rect 2380 -770 2410 -740
rect 2380 -790 2385 -770
rect 2405 -790 2410 -770
rect 2380 -820 2410 -790
rect 2380 -840 2385 -820
rect 2405 -840 2410 -820
rect 2380 -870 2410 -840
rect 2380 -890 2385 -870
rect 2405 -890 2410 -870
rect 2380 -920 2410 -890
rect 2380 -940 2385 -920
rect 2405 -940 2410 -920
rect 2380 -970 2410 -940
rect 2380 -990 2385 -970
rect 2405 -990 2410 -970
rect 2380 -1020 2410 -990
rect 2380 -1040 2385 -1020
rect 2405 -1040 2410 -1020
rect 2380 -1050 2410 -1040
rect 2480 -370 2510 -360
rect 2480 -390 2485 -370
rect 2505 -390 2510 -370
rect 2480 -420 2510 -390
rect 2480 -440 2485 -420
rect 2505 -440 2510 -420
rect 2480 -470 2510 -440
rect 2480 -490 2485 -470
rect 2505 -490 2510 -470
rect 2480 -520 2510 -490
rect 2480 -540 2485 -520
rect 2505 -540 2510 -520
rect 2480 -570 2510 -540
rect 2480 -590 2485 -570
rect 2505 -590 2510 -570
rect 2480 -620 2510 -590
rect 2480 -640 2485 -620
rect 2505 -640 2510 -620
rect 2480 -670 2510 -640
rect 2480 -690 2485 -670
rect 2505 -690 2510 -670
rect 2480 -720 2510 -690
rect 2480 -740 2485 -720
rect 2505 -740 2510 -720
rect 2480 -770 2510 -740
rect 2480 -790 2485 -770
rect 2505 -790 2510 -770
rect 2480 -820 2510 -790
rect 2480 -840 2485 -820
rect 2505 -840 2510 -820
rect 2480 -870 2510 -840
rect 2480 -890 2485 -870
rect 2505 -890 2510 -870
rect 2480 -920 2510 -890
rect 2480 -940 2485 -920
rect 2505 -940 2510 -920
rect 2480 -970 2510 -940
rect 2480 -990 2485 -970
rect 2505 -990 2510 -970
rect 2480 -1020 2510 -990
rect 2480 -1040 2485 -1020
rect 2505 -1040 2510 -1020
rect 2480 -1050 2510 -1040
rect 2580 -370 2610 -360
rect 2580 -390 2585 -370
rect 2605 -390 2610 -370
rect 2580 -420 2610 -390
rect 2580 -440 2585 -420
rect 2605 -440 2610 -420
rect 2580 -470 2610 -440
rect 2580 -490 2585 -470
rect 2605 -490 2610 -470
rect 2580 -520 2610 -490
rect 2580 -540 2585 -520
rect 2605 -540 2610 -520
rect 2580 -570 2610 -540
rect 2580 -590 2585 -570
rect 2605 -590 2610 -570
rect 2580 -620 2610 -590
rect 2580 -640 2585 -620
rect 2605 -640 2610 -620
rect 2580 -670 2610 -640
rect 2580 -690 2585 -670
rect 2605 -690 2610 -670
rect 2580 -720 2610 -690
rect 2580 -740 2585 -720
rect 2605 -740 2610 -720
rect 2580 -770 2610 -740
rect 2580 -790 2585 -770
rect 2605 -790 2610 -770
rect 2580 -820 2610 -790
rect 2580 -840 2585 -820
rect 2605 -840 2610 -820
rect 2580 -870 2610 -840
rect 2580 -890 2585 -870
rect 2605 -890 2610 -870
rect 2580 -920 2610 -890
rect 2580 -940 2585 -920
rect 2605 -940 2610 -920
rect 2580 -970 2610 -940
rect 2580 -990 2585 -970
rect 2605 -990 2610 -970
rect 2580 -1020 2610 -990
rect 2580 -1040 2585 -1020
rect 2605 -1040 2610 -1020
rect 2580 -1050 2610 -1040
rect 2680 -370 2750 -360
rect 2680 -390 2685 -370
rect 2705 -390 2725 -370
rect 2745 -390 2750 -370
rect 2680 -420 2750 -390
rect 2680 -440 2685 -420
rect 2705 -440 2725 -420
rect 2745 -440 2750 -420
rect 2680 -470 2750 -440
rect 2680 -490 2685 -470
rect 2705 -490 2725 -470
rect 2745 -490 2750 -470
rect 2680 -520 2750 -490
rect 2680 -540 2685 -520
rect 2705 -540 2725 -520
rect 2745 -540 2750 -520
rect 2680 -570 2750 -540
rect 2680 -590 2685 -570
rect 2705 -590 2725 -570
rect 2745 -590 2750 -570
rect 2680 -620 2750 -590
rect 2680 -640 2685 -620
rect 2705 -640 2725 -620
rect 2745 -640 2750 -620
rect 2805 -387 2840 -380
rect 2805 -407 2810 -387
rect 2835 -407 2840 -387
rect 2805 -415 2840 -407
rect 2865 -387 2900 -380
rect 2865 -407 2870 -387
rect 2895 -407 2900 -387
rect 2865 -415 2900 -407
rect 2680 -670 2750 -640
rect 2680 -690 2685 -670
rect 2705 -690 2725 -670
rect 2745 -690 2750 -670
rect 2680 -720 2750 -690
rect 2680 -740 2685 -720
rect 2705 -740 2725 -720
rect 2745 -740 2750 -720
rect 2680 -770 2750 -740
rect 2680 -790 2685 -770
rect 2705 -790 2725 -770
rect 2745 -790 2750 -770
rect 2680 -820 2750 -790
rect 2680 -840 2685 -820
rect 2705 -840 2725 -820
rect 2745 -840 2750 -820
rect 2680 -870 2750 -840
rect 2680 -890 2685 -870
rect 2705 -890 2725 -870
rect 2745 -890 2750 -870
rect 2680 -920 2750 -890
rect 2680 -940 2685 -920
rect 2705 -940 2725 -920
rect 2745 -940 2750 -920
rect 2680 -970 2750 -940
rect 2680 -990 2685 -970
rect 2705 -990 2725 -970
rect 2745 -990 2750 -970
rect 2680 -1020 2750 -990
rect 2680 -1040 2685 -1020
rect 2705 -1040 2725 -1020
rect 2745 -1040 2750 -1020
rect 2680 -1050 2750 -1040
rect -1015 -1070 -995 -1050
rect -815 -1070 -795 -1050
rect -615 -1070 -595 -1050
rect -415 -1070 -395 -1050
rect 2085 -1070 2105 -1050
rect 2285 -1070 2305 -1050
rect 2485 -1070 2505 -1050
rect 2685 -1070 2705 -1050
rect -1025 -1080 -985 -1070
rect -1025 -1100 -1015 -1080
rect -995 -1100 -985 -1080
rect -1025 -1110 -985 -1100
rect -825 -1080 -785 -1070
rect -825 -1100 -815 -1080
rect -795 -1100 -785 -1080
rect -825 -1110 -785 -1100
rect -625 -1080 -585 -1070
rect -625 -1100 -615 -1080
rect -595 -1100 -585 -1080
rect -625 -1110 -585 -1100
rect -425 -1080 -385 -1070
rect -425 -1100 -415 -1080
rect -395 -1100 -385 -1080
rect -425 -1110 -385 -1100
rect 2075 -1080 2115 -1070
rect 2075 -1100 2085 -1080
rect 2105 -1100 2115 -1080
rect 2075 -1110 2115 -1100
rect 2275 -1080 2315 -1070
rect 2275 -1100 2285 -1080
rect 2305 -1100 2315 -1080
rect 2275 -1110 2315 -1100
rect 2475 -1080 2515 -1070
rect 2475 -1100 2485 -1080
rect 2505 -1100 2515 -1080
rect 2475 -1110 2515 -1100
rect 2675 -1080 2715 -1070
rect 2675 -1100 2685 -1080
rect 2705 -1100 2715 -1080
rect 2675 -1110 2715 -1100
rect 2840 -1105 2865 -1055
<< viali >>
rect 40 2700 60 2720
rect 160 2700 180 2720
rect 220 2700 240 2720
rect 980 2700 1000 2720
rect 1040 2700 1060 2720
rect 1100 2700 1120 2720
rect 1160 2700 1180 2720
rect 1448 2700 1468 2720
rect 1508 2700 1528 2720
rect 1628 2700 1648 2720
rect 510 2530 530 2550
rect 570 2530 590 2550
rect 630 2530 650 2550
rect 690 2530 710 2550
rect 85 2280 105 2300
rect 144 2280 164 2300
rect 614 2280 634 2300
rect 1056 2280 1076 2300
rect 1524 2280 1544 2300
rect 1583 2280 1603 2300
rect -1075 2125 -1055 2145
rect -955 2125 -935 2145
rect -835 2125 -815 2145
rect -715 2125 -695 2145
rect -595 2125 -575 2145
rect -475 2125 -455 2145
rect -355 2125 -335 2145
rect -30 2125 -10 2145
rect 90 2125 110 2145
rect 210 2125 230 2145
rect 330 2125 350 2145
rect 450 2125 470 2145
rect 570 2125 590 2145
rect 690 2125 710 2145
rect 980 2125 1000 2145
rect 1100 2125 1120 2145
rect 1220 2125 1240 2145
rect 1340 2125 1360 2145
rect 1460 2125 1480 2145
rect 1580 2125 1600 2145
rect 1700 2125 1720 2145
rect 2025 2125 2045 2145
rect 2145 2125 2165 2145
rect 2265 2125 2285 2145
rect 2385 2125 2405 2145
rect 2505 2125 2525 2145
rect 2625 2125 2645 2145
rect 2745 2125 2765 2145
rect -1015 1700 -995 1720
rect -895 1700 -875 1720
rect -775 1700 -755 1720
rect -715 1700 -695 1720
rect -655 1700 -635 1720
rect -535 1700 -515 1720
rect -415 1700 -395 1720
rect 30 1700 50 1720
rect 150 1700 170 1720
rect 270 1700 290 1720
rect 330 1700 350 1720
rect 390 1700 410 1720
rect 510 1700 530 1720
rect 630 1700 650 1720
rect 1040 1700 1060 1720
rect 1160 1700 1180 1720
rect 1280 1700 1300 1720
rect 1340 1700 1360 1720
rect 1400 1700 1420 1720
rect 1520 1700 1540 1720
rect 1640 1700 1660 1720
rect 2085 1700 2105 1720
rect 2205 1700 2225 1720
rect 2325 1700 2345 1720
rect 2385 1700 2405 1720
rect 2445 1700 2465 1720
rect 2565 1700 2585 1720
rect 2685 1700 2705 1720
rect 230 1555 250 1575
rect 340 1555 360 1575
rect 450 1555 470 1575
rect 560 1555 580 1575
rect 670 1555 690 1575
rect 780 1555 800 1575
rect 890 1555 910 1575
rect 1000 1555 1020 1575
rect 1110 1555 1130 1575
rect 1220 1555 1240 1575
rect 1330 1555 1350 1575
rect 1440 1555 1460 1575
rect -1045 1460 -1025 1480
rect -935 1460 -915 1480
rect -825 1460 -805 1480
rect -715 1460 -695 1480
rect -605 1460 -585 1480
rect -495 1460 -475 1480
rect -385 1460 -365 1480
rect 2055 1460 2075 1480
rect 285 1430 305 1450
rect -1495 1400 -1475 1420
rect -1440 1400 -1420 1420
rect -1385 1400 -1365 1420
rect 395 1430 415 1450
rect 505 1430 525 1450
rect 615 1430 635 1450
rect 725 1430 745 1450
rect 835 1430 855 1450
rect 890 1430 910 1450
rect 945 1430 965 1450
rect 1055 1430 1075 1450
rect 1165 1430 1185 1450
rect 1275 1430 1295 1450
rect 2165 1460 2185 1480
rect 2275 1460 2295 1480
rect 2385 1460 2405 1480
rect 2495 1460 2515 1480
rect 2605 1460 2625 1480
rect 2715 1460 2735 1480
rect 1385 1430 1405 1450
rect 76 1230 96 1250
rect 125 1230 145 1250
rect 225 1230 245 1250
rect 280 1230 300 1250
rect 335 1230 355 1250
rect 445 1230 465 1250
rect 500 1230 520 1250
rect 555 1230 575 1250
rect 1076 1230 1096 1250
rect 1125 1230 1145 1250
rect 1225 1230 1245 1250
rect 1280 1230 1300 1250
rect 1335 1230 1355 1250
rect 1445 1230 1465 1250
rect 1500 1230 1520 1250
rect 1555 1230 1575 1250
rect -35 1170 -15 1190
rect 1705 1170 1725 1190
rect 60 1105 80 1125
rect 155 1105 175 1125
rect 209 1111 229 1131
rect 280 1105 300 1125
rect 375 1105 395 1125
rect 429 1111 449 1131
rect 500 1105 520 1125
rect 571 1111 591 1131
rect 620 1105 640 1125
rect 1060 1105 1080 1125
rect 1155 1105 1175 1125
rect 1209 1111 1229 1131
rect 1280 1105 1300 1125
rect 1375 1105 1395 1125
rect 1429 1111 1449 1131
rect 1500 1105 1520 1125
rect 1571 1111 1591 1131
rect 1620 1105 1640 1125
rect 560 905 580 925
rect 670 905 690 925
rect 780 905 800 925
rect 890 905 910 925
rect 1000 905 1020 925
rect 1110 905 1130 925
rect 3055 1400 3075 1420
rect 3110 1400 3130 1420
rect 3165 1400 3185 1420
rect -1495 795 -1475 815
rect -1440 795 -1420 815
rect -1385 795 -1365 815
rect -990 785 -970 805
rect -880 785 -860 805
rect -770 785 -750 805
rect -715 780 -695 800
rect -660 785 -640 805
rect -550 785 -530 805
rect -440 785 -420 805
rect 505 785 525 805
rect 615 785 635 805
rect 725 785 745 805
rect 835 785 855 805
rect 945 785 965 805
rect 1055 785 1075 805
rect 1165 785 1185 805
rect 2110 785 2130 805
rect 2220 785 2240 805
rect 2330 785 2350 805
rect 2385 780 2405 800
rect 2440 785 2460 805
rect 2550 785 2570 805
rect 2660 785 2680 805
rect 3055 795 3075 815
rect 3110 795 3130 815
rect 3165 795 3185 815
rect -1055 645 -1035 665
rect -990 645 -970 665
rect -880 645 -860 665
rect -770 645 -750 665
rect -660 645 -640 665
rect -550 645 -530 665
rect -440 645 -420 665
rect -375 645 -355 665
rect 40 635 60 655
rect 150 635 170 655
rect 260 635 280 655
rect 315 635 335 655
rect 370 635 390 655
rect 480 635 500 655
rect 590 635 610 655
rect 1080 635 1100 655
rect 1190 635 1210 655
rect 1300 635 1320 655
rect 1355 635 1375 655
rect 1410 635 1430 655
rect 1520 635 1540 655
rect 1630 635 1650 655
rect 2045 645 2065 665
rect 2110 645 2130 665
rect 2220 645 2240 665
rect 2330 645 2350 665
rect 2440 645 2460 665
rect 2550 645 2570 665
rect 2660 645 2680 665
rect 2725 645 2745 665
rect -15 410 5 430
rect 95 410 115 430
rect 205 410 225 430
rect 315 410 335 430
rect 425 410 445 430
rect 535 410 555 430
rect 645 410 665 430
rect 1025 410 1045 430
rect 1135 410 1155 430
rect 1245 410 1265 430
rect 1355 410 1375 430
rect 1465 410 1485 430
rect 1575 410 1595 430
rect 1685 410 1705 430
rect -935 370 -915 390
rect -825 370 -805 390
rect -715 370 -695 390
rect -660 370 -640 390
rect -605 370 -585 390
rect -495 370 -475 390
rect 2165 370 2185 390
rect 2275 370 2295 390
rect 2330 370 2350 390
rect 2385 370 2405 390
rect 2495 370 2515 390
rect 2605 370 2625 390
rect -935 260 -915 280
rect -825 260 -805 280
rect -715 260 -695 280
rect -660 260 -640 280
rect -605 260 -585 280
rect -495 260 -475 280
rect 2165 260 2185 280
rect 2275 260 2295 280
rect 2330 260 2350 280
rect 2385 260 2405 280
rect 2495 260 2515 280
rect 2605 260 2625 280
rect -1405 -113 -1380 -93
rect -1345 -113 -1320 -93
rect -1285 -113 -1260 -93
rect 40 205 60 225
rect 150 205 170 225
rect 260 205 280 225
rect 370 205 390 225
rect 480 205 500 225
rect 590 205 610 225
rect 1080 205 1100 225
rect 1190 205 1210 225
rect 1300 205 1320 225
rect 1410 205 1430 225
rect 1520 205 1540 225
rect 1630 205 1650 225
rect 315 155 335 175
rect 800 155 820 175
rect 853 155 873 175
rect 900 155 920 175
rect 1355 155 1375 175
rect -15 -65 5 -45
rect 95 -65 115 -45
rect 205 -65 225 -45
rect 315 -65 335 -45
rect 425 -65 445 -45
rect 535 -65 555 -45
rect 685 -65 705 -45
rect 780 -65 800 -45
rect 835 -65 855 -45
rect 890 -65 910 -45
rect 985 -65 1005 -45
rect 1135 -65 1155 -45
rect 1245 -65 1265 -45
rect 1355 -65 1375 -45
rect 1465 -65 1485 -45
rect 1575 -65 1595 -45
rect 1685 -65 1705 -45
rect -1225 -113 -1200 -93
rect -1055 -115 -1035 -95
rect -990 -115 -970 -95
rect -880 -115 -860 -95
rect -770 -115 -750 -95
rect -660 -115 -640 -95
rect -550 -115 -530 -95
rect -440 -115 -420 -95
rect -375 -115 -355 -95
rect 2045 -115 2065 -95
rect 2110 -115 2130 -95
rect 2220 -115 2240 -95
rect 2330 -115 2350 -95
rect 2440 -115 2460 -95
rect 2550 -115 2570 -95
rect 2660 -115 2680 -95
rect 2725 -115 2745 -95
rect 2890 -113 2915 -93
rect 2950 -113 2975 -93
rect 3010 -113 3035 -93
rect 3070 -113 3095 -93
rect -915 -325 -895 -305
rect -715 -325 -695 -305
rect -615 -325 -595 -305
rect -515 -325 -495 -305
rect 2185 -325 2205 -305
rect 2285 -325 2305 -305
rect 2385 -325 2405 -305
rect 2585 -325 2605 -305
rect -1205 -407 -1180 -387
rect -1145 -407 -1120 -387
rect 280 -375 300 -355
rect 390 -375 410 -355
rect 500 -375 520 -355
rect 610 -375 630 -355
rect 720 -375 740 -355
rect 775 -375 795 -355
rect 830 -375 850 -355
rect 940 -375 960 -355
rect 1050 -375 1070 -355
rect 1160 -375 1180 -355
rect 1270 -375 1290 -355
rect 1341 -375 1361 -355
rect 1395 -375 1415 -355
rect 160 -700 180 -680
rect 225 -700 245 -680
rect 335 -700 355 -680
rect 445 -700 465 -680
rect 555 -700 575 -680
rect 665 -700 685 -680
rect 775 -700 795 -680
rect 885 -700 905 -680
rect 995 -700 1015 -680
rect 1105 -700 1125 -680
rect 1215 -700 1235 -680
rect 1325 -700 1345 -680
rect 1435 -700 1455 -680
rect 1020 -760 1040 -740
rect 720 -795 740 -775
rect 835 -795 855 -775
rect 960 -795 980 -775
rect 2810 -407 2835 -387
rect 2870 -407 2895 -387
rect -1015 -1100 -995 -1080
rect -815 -1100 -795 -1080
rect -615 -1100 -595 -1080
rect -415 -1100 -395 -1080
rect 2085 -1100 2105 -1080
rect 2285 -1100 2305 -1080
rect 2485 -1100 2505 -1080
rect 2685 -1100 2705 -1080
<< metal1 >>
rect 825 4275 865 4280
rect 825 4245 830 4275
rect 860 4245 865 4275
rect 825 4240 865 4245
rect 150 2780 190 2785
rect 150 2750 155 2780
rect 185 2750 190 2780
rect 150 2745 190 2750
rect 620 2780 660 2785
rect 620 2750 625 2780
rect 655 2750 660 2780
rect 620 2745 660 2750
rect 160 2730 180 2745
rect 30 2725 70 2730
rect 30 2695 35 2725
rect 65 2695 70 2725
rect 30 2690 70 2695
rect 150 2725 190 2730
rect 150 2695 155 2725
rect 185 2695 190 2725
rect 150 2690 190 2695
rect 210 2725 250 2730
rect 210 2695 215 2725
rect 245 2695 250 2725
rect 210 2690 250 2695
rect 630 2560 650 2745
rect 835 2730 855 4240
rect 1030 2780 1070 2785
rect 1030 2750 1035 2780
rect 1065 2750 1070 2780
rect 1030 2745 1070 2750
rect 1498 2780 1538 2785
rect 1498 2750 1503 2780
rect 1533 2750 1538 2780
rect 1498 2745 1538 2750
rect 1040 2730 1060 2745
rect 1508 2730 1528 2745
rect 825 2725 865 2730
rect 825 2695 830 2725
rect 860 2695 865 2725
rect 825 2690 865 2695
rect 970 2725 1010 2730
rect 970 2695 975 2725
rect 1005 2695 1010 2725
rect 970 2690 1010 2695
rect 1035 2720 1065 2730
rect 1035 2700 1040 2720
rect 1060 2700 1065 2720
rect 1035 2690 1065 2700
rect 1090 2725 1130 2730
rect 1090 2695 1095 2725
rect 1125 2695 1130 2725
rect 1090 2690 1130 2695
rect 1150 2725 1190 2730
rect 1150 2695 1155 2725
rect 1185 2695 1190 2725
rect 1150 2690 1190 2695
rect 1438 2725 1478 2730
rect 1438 2695 1443 2725
rect 1473 2695 1478 2725
rect 1438 2690 1478 2695
rect 1498 2725 1538 2730
rect 1498 2695 1503 2725
rect 1533 2695 1538 2725
rect 1498 2690 1538 2695
rect 1618 2725 1658 2730
rect 1618 2695 1623 2725
rect 1653 2695 1658 2725
rect 1618 2690 1658 2695
rect 835 2560 855 2690
rect 500 2555 540 2560
rect 500 2525 505 2555
rect 535 2525 540 2555
rect 500 2520 540 2525
rect 560 2555 600 2560
rect 560 2525 565 2555
rect 595 2525 600 2555
rect 560 2520 600 2525
rect 625 2550 655 2560
rect 625 2530 630 2550
rect 650 2530 655 2550
rect 625 2520 655 2530
rect 680 2555 720 2560
rect 680 2525 685 2555
rect 715 2525 720 2555
rect 680 2520 720 2525
rect 825 2555 865 2560
rect 825 2525 830 2555
rect 860 2525 865 2555
rect 825 2520 865 2525
rect 75 2305 115 2310
rect 75 2275 80 2305
rect 110 2275 115 2305
rect 75 2270 115 2275
rect 139 2305 169 2310
rect 139 2270 169 2275
rect 609 2305 639 2310
rect 609 2270 639 2275
rect 770 2305 810 2310
rect 770 2275 775 2305
rect 805 2275 810 2305
rect 770 2270 810 2275
rect -725 2205 -685 2210
rect -725 2175 -720 2205
rect -690 2175 -685 2205
rect -725 2170 -685 2175
rect -155 2205 -115 2210
rect -155 2175 -150 2205
rect -120 2175 -115 2205
rect -155 2170 -115 2175
rect -715 2155 -695 2170
rect -1085 2150 -1045 2155
rect -1085 2120 -1080 2150
rect -1050 2120 -1045 2150
rect -1085 2115 -1045 2120
rect -965 2150 -925 2155
rect -965 2120 -960 2150
rect -930 2120 -925 2150
rect -965 2115 -925 2120
rect -845 2150 -805 2155
rect -845 2120 -840 2150
rect -810 2120 -805 2150
rect -845 2115 -805 2120
rect -725 2150 -685 2155
rect -725 2120 -720 2150
rect -690 2120 -685 2150
rect -725 2115 -685 2120
rect -605 2150 -565 2155
rect -605 2120 -600 2150
rect -570 2120 -565 2150
rect -605 2115 -565 2120
rect -485 2150 -445 2155
rect -485 2120 -480 2150
rect -450 2120 -445 2150
rect -485 2115 -445 2120
rect -365 2150 -325 2155
rect -365 2120 -360 2150
rect -330 2120 -325 2150
rect -365 2115 -325 2120
rect -200 2150 -160 2155
rect -200 2120 -195 2150
rect -165 2120 -160 2150
rect -200 2115 -160 2120
rect -190 1730 -170 2115
rect -1025 1725 -985 1730
rect -1025 1695 -1020 1725
rect -990 1695 -985 1725
rect -1025 1690 -985 1695
rect -905 1725 -865 1730
rect -905 1695 -900 1725
rect -870 1695 -865 1725
rect -905 1690 -865 1695
rect -785 1725 -745 1730
rect -785 1695 -780 1725
rect -750 1695 -745 1725
rect -785 1690 -745 1695
rect -720 1720 -690 1730
rect -720 1700 -715 1720
rect -695 1700 -690 1720
rect -720 1690 -690 1700
rect -665 1725 -625 1730
rect -665 1695 -660 1725
rect -630 1695 -625 1725
rect -665 1690 -625 1695
rect -545 1725 -505 1730
rect -545 1695 -540 1725
rect -510 1695 -505 1725
rect -545 1690 -505 1695
rect -425 1725 -385 1730
rect -425 1695 -420 1725
rect -390 1695 -385 1725
rect -425 1690 -385 1695
rect -200 1725 -160 1730
rect -200 1695 -195 1725
rect -165 1695 -160 1725
rect -200 1690 -160 1695
rect -715 1630 -695 1690
rect -290 1670 -250 1675
rect -290 1640 -285 1670
rect -255 1640 -250 1670
rect -290 1635 -250 1640
rect -725 1625 -685 1630
rect -725 1595 -720 1625
rect -690 1595 -685 1625
rect -725 1590 -685 1595
rect -1450 1540 -1410 1545
rect -1450 1510 -1445 1540
rect -1415 1510 -1410 1540
rect -1450 1505 -1410 1510
rect -1440 1430 -1420 1505
rect -1055 1485 -1015 1490
rect -1055 1455 -1050 1485
rect -1020 1455 -1015 1485
rect -1055 1450 -1015 1455
rect -945 1485 -905 1490
rect -945 1455 -940 1485
rect -910 1455 -905 1485
rect -945 1450 -905 1455
rect -835 1485 -795 1490
rect -835 1455 -830 1485
rect -800 1455 -795 1485
rect -835 1450 -795 1455
rect -725 1485 -685 1490
rect -725 1455 -720 1485
rect -690 1455 -685 1485
rect -725 1450 -685 1455
rect -615 1485 -575 1490
rect -615 1455 -610 1485
rect -580 1455 -575 1485
rect -615 1450 -575 1455
rect -505 1485 -465 1490
rect -505 1455 -500 1485
rect -470 1455 -465 1485
rect -505 1450 -465 1455
rect -395 1485 -355 1490
rect -395 1455 -390 1485
rect -360 1455 -355 1485
rect -395 1450 -355 1455
rect -1501 1420 -1360 1430
rect -1501 1400 -1495 1420
rect -1475 1400 -1440 1420
rect -1420 1400 -1385 1420
rect -1365 1400 -1360 1420
rect -1501 1390 -1360 1400
rect -1501 815 -1360 825
rect -1501 795 -1495 815
rect -1475 795 -1440 815
rect -1420 795 -1385 815
rect -1365 795 -1360 815
rect -1501 785 -1360 795
rect -1000 810 -960 815
rect -1540 760 -1500 765
rect -1540 730 -1535 760
rect -1505 730 -1500 760
rect -1540 725 -1500 730
rect -1530 360 -1510 725
rect -1440 720 -1420 785
rect -1000 780 -995 810
rect -965 780 -960 810
rect -1000 775 -960 780
rect -890 810 -850 815
rect -890 780 -885 810
rect -855 780 -850 810
rect -890 775 -850 780
rect -780 810 -740 815
rect -670 810 -630 815
rect -780 780 -775 810
rect -745 780 -740 810
rect -780 775 -740 780
rect -720 800 -690 810
rect -720 780 -715 800
rect -695 780 -690 800
rect -880 760 -860 775
rect -720 770 -690 780
rect -670 780 -665 810
rect -635 780 -630 810
rect -670 775 -630 780
rect -560 810 -520 815
rect -560 780 -555 810
rect -525 780 -520 810
rect -560 775 -520 780
rect -450 810 -410 815
rect -450 780 -445 810
rect -415 780 -410 810
rect -450 775 -410 780
rect -890 730 -885 760
rect -855 730 -850 760
rect -715 720 -695 770
rect -450 730 -445 760
rect -415 730 -410 760
rect -1450 715 -1410 720
rect -1450 685 -1445 715
rect -1415 685 -1410 715
rect -1450 680 -1410 685
rect -725 715 -685 720
rect -725 685 -720 715
rect -690 685 -685 715
rect -725 680 -685 685
rect -440 675 -420 730
rect -280 720 -260 1635
rect -145 1490 -125 2170
rect -40 2150 0 2155
rect -40 2120 -35 2150
rect -5 2120 0 2150
rect -40 2115 0 2120
rect 80 2150 120 2155
rect 80 2120 85 2150
rect 115 2120 120 2150
rect 80 2115 120 2120
rect 200 2150 240 2155
rect 200 2120 205 2150
rect 235 2120 240 2150
rect 200 2115 240 2120
rect 320 2150 360 2155
rect 320 2120 325 2150
rect 355 2120 360 2150
rect 320 2115 360 2120
rect 440 2150 480 2155
rect 440 2120 445 2150
rect 475 2120 480 2150
rect 440 2115 480 2120
rect 560 2150 600 2155
rect 560 2120 565 2150
rect 595 2120 600 2150
rect 560 2115 600 2120
rect 680 2150 720 2155
rect 680 2120 685 2150
rect 715 2120 720 2150
rect 680 2115 720 2120
rect 20 1725 60 1730
rect 20 1695 25 1725
rect 55 1695 60 1725
rect 20 1690 60 1695
rect 140 1725 180 1730
rect 140 1695 145 1725
rect 175 1695 180 1725
rect 140 1690 180 1695
rect 260 1725 300 1730
rect 260 1695 265 1725
rect 295 1695 300 1725
rect 260 1690 300 1695
rect 325 1720 355 1730
rect 325 1700 330 1720
rect 350 1700 355 1720
rect 325 1690 355 1700
rect 380 1725 420 1730
rect 380 1695 385 1725
rect 415 1695 420 1725
rect 380 1690 420 1695
rect 500 1725 540 1730
rect 500 1695 505 1725
rect 535 1695 540 1725
rect 500 1690 540 1695
rect 620 1725 660 1730
rect 620 1695 625 1725
rect 655 1695 660 1725
rect 620 1690 660 1695
rect 30 1675 50 1690
rect 330 1675 350 1690
rect 790 1675 810 2270
rect 835 2210 855 2520
rect 1051 2300 1081 2310
rect 1051 2280 1056 2300
rect 1076 2280 1081 2300
rect 1051 2270 1081 2280
rect 1519 2305 1549 2310
rect 1519 2270 1549 2275
rect 1573 2300 1613 2310
rect 1573 2280 1583 2300
rect 1603 2280 1613 2300
rect 1573 2270 1613 2280
rect 880 2260 920 2265
rect 880 2230 885 2260
rect 915 2230 920 2260
rect 1055 2255 1075 2270
rect 1583 2255 1603 2270
rect 880 2225 920 2230
rect 1045 2250 1085 2255
rect 825 2205 865 2210
rect 825 2175 830 2205
rect 860 2175 865 2205
rect 825 2170 865 2175
rect 20 1670 60 1675
rect 20 1640 25 1670
rect 55 1640 60 1670
rect 20 1635 60 1640
rect 320 1670 360 1675
rect 320 1640 325 1670
rect 355 1640 360 1670
rect 320 1635 360 1640
rect 780 1670 820 1675
rect 780 1640 785 1670
rect 815 1640 820 1670
rect 780 1635 820 1640
rect 880 1630 900 2225
rect 1045 2220 1050 2250
rect 1080 2220 1085 2250
rect 1045 2215 1085 2220
rect 1573 2250 1613 2255
rect 1573 2220 1578 2250
rect 1608 2220 1613 2250
rect 1573 2215 1613 2220
rect 1805 2205 1845 2210
rect 1805 2175 1810 2205
rect 1840 2175 1845 2205
rect 1805 2170 1845 2175
rect 2375 2205 2415 2210
rect 2375 2175 2380 2205
rect 2410 2175 2415 2205
rect 2375 2170 2415 2175
rect 970 2150 1010 2155
rect 970 2120 975 2150
rect 1005 2120 1010 2150
rect 970 2115 1010 2120
rect 1090 2150 1130 2155
rect 1090 2120 1095 2150
rect 1125 2120 1130 2150
rect 1090 2115 1130 2120
rect 1210 2150 1250 2155
rect 1210 2120 1215 2150
rect 1245 2120 1250 2150
rect 1210 2115 1250 2120
rect 1330 2150 1370 2155
rect 1330 2120 1335 2150
rect 1365 2120 1370 2150
rect 1330 2115 1370 2120
rect 1450 2150 1490 2155
rect 1450 2120 1455 2150
rect 1485 2120 1490 2150
rect 1450 2115 1490 2120
rect 1570 2150 1610 2155
rect 1570 2120 1575 2150
rect 1605 2120 1610 2150
rect 1570 2115 1610 2120
rect 1690 2150 1730 2155
rect 1690 2120 1695 2150
rect 1725 2120 1730 2150
rect 1690 2115 1730 2120
rect 1030 1725 1070 1730
rect 1030 1695 1035 1725
rect 1065 1695 1070 1725
rect 1030 1690 1070 1695
rect 1150 1725 1190 1730
rect 1150 1695 1155 1725
rect 1185 1695 1190 1725
rect 1150 1690 1190 1695
rect 1270 1725 1310 1730
rect 1270 1695 1275 1725
rect 1305 1695 1310 1725
rect 1270 1690 1310 1695
rect 1335 1720 1365 1730
rect 1335 1700 1340 1720
rect 1360 1700 1365 1720
rect 1335 1690 1365 1700
rect 1390 1725 1430 1730
rect 1390 1695 1395 1725
rect 1425 1695 1430 1725
rect 1390 1690 1430 1695
rect 1510 1725 1550 1730
rect 1510 1695 1515 1725
rect 1545 1695 1550 1725
rect 1510 1690 1550 1695
rect 1630 1725 1670 1730
rect 1630 1695 1635 1725
rect 1665 1695 1670 1725
rect 1630 1690 1670 1695
rect 1340 1675 1360 1690
rect 1640 1675 1660 1690
rect 1330 1670 1370 1675
rect 1330 1640 1335 1670
rect 1365 1640 1370 1670
rect 1330 1635 1370 1640
rect 1630 1670 1670 1675
rect 1630 1640 1635 1670
rect 1665 1640 1670 1670
rect 1630 1635 1670 1640
rect 870 1600 875 1630
rect 905 1600 910 1630
rect 1815 1585 1835 2170
rect 2385 2155 2405 2170
rect 1850 2150 1890 2155
rect 1850 2120 1855 2150
rect 1885 2120 1890 2150
rect 1850 2115 1890 2120
rect 2015 2150 2055 2155
rect 2015 2120 2020 2150
rect 2050 2120 2055 2150
rect 2015 2115 2055 2120
rect 2135 2150 2175 2155
rect 2135 2120 2140 2150
rect 2170 2120 2175 2150
rect 2135 2115 2175 2120
rect 2255 2150 2295 2155
rect 2255 2120 2260 2150
rect 2290 2120 2295 2150
rect 2255 2115 2295 2120
rect 2375 2150 2415 2155
rect 2375 2120 2380 2150
rect 2410 2120 2415 2150
rect 2375 2115 2415 2120
rect 2495 2150 2535 2155
rect 2495 2120 2500 2150
rect 2530 2120 2535 2150
rect 2495 2115 2535 2120
rect 2615 2150 2655 2155
rect 2615 2120 2620 2150
rect 2650 2120 2655 2150
rect 2615 2115 2655 2120
rect 2735 2150 2775 2155
rect 2735 2120 2740 2150
rect 2770 2120 2775 2150
rect 2735 2115 2775 2120
rect 1860 1730 1880 2115
rect 1850 1725 1890 1730
rect 1850 1695 1855 1725
rect 1885 1695 1890 1725
rect 1850 1690 1890 1695
rect 2075 1725 2115 1730
rect 2075 1695 2080 1725
rect 2110 1695 2115 1725
rect 2075 1690 2115 1695
rect 2195 1725 2235 1730
rect 2195 1695 2200 1725
rect 2230 1695 2235 1725
rect 2195 1690 2235 1695
rect 2315 1725 2355 1730
rect 2315 1695 2320 1725
rect 2350 1695 2355 1725
rect 2315 1690 2355 1695
rect 2380 1720 2410 1730
rect 2380 1700 2385 1720
rect 2405 1700 2410 1720
rect 2380 1690 2410 1700
rect 2435 1725 2475 1730
rect 2435 1695 2440 1725
rect 2470 1695 2475 1725
rect 2435 1690 2475 1695
rect 2555 1725 2595 1730
rect 2555 1695 2560 1725
rect 2590 1695 2595 1725
rect 2555 1690 2595 1695
rect 2675 1725 2715 1730
rect 2675 1695 2680 1725
rect 2710 1695 2715 1725
rect 2675 1690 2715 1695
rect 1940 1670 1980 1675
rect 1940 1640 1945 1670
rect 1975 1640 1980 1670
rect 1940 1635 1980 1640
rect 220 1580 260 1585
rect 220 1550 225 1580
rect 255 1550 260 1580
rect 220 1545 260 1550
rect 330 1580 370 1585
rect 330 1550 335 1580
rect 365 1550 370 1580
rect 330 1545 370 1550
rect 440 1580 480 1585
rect 440 1550 445 1580
rect 475 1550 480 1580
rect 440 1545 480 1550
rect 550 1580 590 1585
rect 550 1550 555 1580
rect 585 1550 590 1580
rect 550 1545 590 1550
rect 660 1580 700 1585
rect 660 1550 665 1580
rect 695 1550 700 1580
rect 660 1545 700 1550
rect 770 1580 810 1585
rect 770 1550 775 1580
rect 805 1550 810 1580
rect 770 1545 810 1550
rect 880 1580 920 1585
rect 880 1550 885 1580
rect 915 1550 920 1580
rect 880 1545 920 1550
rect 990 1580 1030 1585
rect 990 1550 995 1580
rect 1025 1550 1030 1580
rect 990 1545 1030 1550
rect 1100 1580 1140 1585
rect 1100 1550 1105 1580
rect 1135 1550 1140 1580
rect 1100 1545 1140 1550
rect 1210 1580 1250 1585
rect 1210 1550 1215 1580
rect 1245 1550 1250 1580
rect 1210 1545 1250 1550
rect 1320 1580 1360 1585
rect 1320 1550 1325 1580
rect 1355 1550 1360 1580
rect 1320 1545 1360 1550
rect 1430 1580 1470 1585
rect 1430 1550 1435 1580
rect 1465 1550 1470 1580
rect 1430 1545 1470 1550
rect 1805 1580 1845 1585
rect 1805 1550 1810 1580
rect 1840 1550 1845 1580
rect 1805 1545 1845 1550
rect 1815 1490 1835 1545
rect -155 1485 -115 1490
rect -155 1455 -150 1485
rect -120 1455 -115 1485
rect 1805 1485 1845 1490
rect -155 1450 -115 1455
rect 275 1455 315 1460
rect -245 1255 -205 1260
rect -245 1225 -240 1255
rect -210 1225 -205 1255
rect -245 1220 -205 1225
rect -290 715 -250 720
rect -290 685 -285 715
rect -255 685 -250 715
rect -290 680 -250 685
rect -1065 670 -1025 675
rect -1065 640 -1060 670
rect -1030 640 -1025 670
rect -1065 635 -1025 640
rect -1000 670 -960 675
rect -1000 640 -995 670
rect -965 640 -960 670
rect -1000 635 -960 640
rect -890 670 -850 675
rect -890 640 -885 670
rect -855 640 -850 670
rect -890 635 -850 640
rect -780 670 -740 675
rect -780 640 -775 670
rect -745 640 -740 670
rect -780 635 -740 640
rect -670 670 -630 675
rect -670 640 -665 670
rect -635 640 -630 670
rect -670 635 -630 640
rect -560 670 -520 675
rect -560 640 -555 670
rect -525 640 -520 670
rect -560 635 -520 640
rect -450 670 -410 675
rect -450 640 -445 670
rect -415 640 -410 670
rect -450 635 -410 640
rect -385 670 -345 675
rect -385 640 -380 670
rect -350 640 -345 670
rect -385 635 -345 640
rect -1190 395 -1150 400
rect -1190 365 -1185 395
rect -1155 365 -1150 395
rect -1190 360 -1150 365
rect -945 395 -905 400
rect -945 365 -940 395
rect -910 365 -905 395
rect -945 360 -905 365
rect -835 395 -795 400
rect -835 365 -830 395
rect -800 365 -795 395
rect -835 360 -795 365
rect -725 395 -685 400
rect -725 365 -720 395
rect -690 365 -685 395
rect -725 360 -685 365
rect -665 390 -635 400
rect -665 370 -660 390
rect -640 370 -635 390
rect -665 360 -635 370
rect -615 395 -575 400
rect -615 365 -610 395
rect -580 365 -575 395
rect -615 360 -575 365
rect -505 395 -465 400
rect -505 365 -500 395
rect -470 365 -465 395
rect -505 360 -465 365
rect -1545 350 -1495 360
rect -1545 320 -1535 350
rect -1505 320 -1495 350
rect -1545 310 -1495 320
rect -1530 -295 -1510 310
rect -1410 -120 -1406 -85
rect -1379 -120 -1375 -85
rect -1350 -120 -1346 -85
rect -1319 -120 -1315 -85
rect -1290 -120 -1286 -85
rect -1259 -120 -1255 -85
rect -1230 -120 -1226 -85
rect -1199 -120 -1195 -85
rect -1405 -185 -1380 -120
rect -1290 -145 -1255 -120
rect -1180 -140 -1160 360
rect -660 345 -640 360
rect -280 345 -260 680
rect -670 340 -630 345
rect -670 310 -665 340
rect -635 310 -630 340
rect -670 305 -630 310
rect -290 340 -250 345
rect -290 310 -285 340
rect -255 310 -250 340
rect -290 305 -250 310
rect -660 290 -640 305
rect -1145 285 -1105 290
rect -1145 255 -1140 285
rect -1110 255 -1105 285
rect -1145 250 -1105 255
rect -945 285 -905 290
rect -945 255 -940 285
rect -910 255 -905 285
rect -945 250 -905 255
rect -835 285 -795 290
rect -835 255 -830 285
rect -800 255 -795 285
rect -835 250 -795 255
rect -725 285 -685 290
rect -725 255 -720 285
rect -690 255 -685 285
rect -725 250 -685 255
rect -665 280 -635 290
rect -665 260 -660 280
rect -640 260 -635 280
rect -665 250 -635 260
rect -615 285 -575 290
rect -615 255 -610 285
rect -580 255 -575 285
rect -615 250 -575 255
rect -505 285 -465 290
rect -505 255 -500 285
rect -470 255 -465 285
rect -505 250 -465 255
rect -1135 -85 -1115 250
rect -1145 -90 -1105 -85
rect -1145 -120 -1140 -90
rect -1110 -120 -1105 -90
rect -1145 -125 -1105 -120
rect -1065 -95 -1025 -85
rect -1065 -115 -1055 -95
rect -1035 -115 -1025 -95
rect -1065 -125 -1025 -115
rect -1000 -90 -960 -85
rect -1000 -120 -995 -90
rect -965 -120 -960 -90
rect -1000 -125 -960 -120
rect -890 -90 -850 -85
rect -890 -120 -885 -90
rect -855 -120 -850 -90
rect -890 -125 -850 -120
rect -780 -90 -740 -85
rect -780 -120 -775 -90
rect -745 -120 -740 -90
rect -780 -125 -740 -120
rect -670 -90 -630 -85
rect -670 -120 -665 -90
rect -635 -120 -630 -90
rect -670 -125 -630 -120
rect -560 -90 -520 -85
rect -560 -120 -555 -90
rect -525 -120 -520 -90
rect -560 -125 -520 -120
rect -450 -90 -410 -85
rect -450 -120 -445 -90
rect -415 -120 -410 -90
rect -450 -125 -410 -120
rect -385 -95 -345 -85
rect -385 -115 -375 -95
rect -355 -115 -345 -95
rect -385 -125 -345 -115
rect -1055 -140 -1035 -125
rect -375 -140 -355 -125
rect -1290 -180 -1255 -175
rect -1190 -145 -1150 -140
rect -1190 -175 -1185 -145
rect -1155 -175 -1150 -145
rect -1190 -180 -1150 -175
rect -1065 -145 -1025 -140
rect -1065 -175 -1060 -145
rect -1030 -175 -1025 -145
rect -1065 -180 -1025 -175
rect -385 -145 -345 -140
rect -385 -175 -380 -145
rect -350 -175 -345 -145
rect -385 -180 -345 -175
rect -1410 -190 -1375 -185
rect -235 -190 -215 1220
rect -145 1200 -125 1450
rect 275 1425 280 1455
rect 310 1425 315 1455
rect 275 1420 315 1425
rect 385 1450 425 1460
rect 385 1430 395 1450
rect 415 1430 425 1450
rect 385 1420 425 1430
rect 495 1455 535 1460
rect 495 1425 500 1455
rect 530 1425 535 1455
rect 495 1420 535 1425
rect 605 1450 645 1460
rect 605 1430 615 1450
rect 635 1430 645 1450
rect 605 1420 645 1430
rect 715 1455 755 1460
rect 715 1425 720 1455
rect 750 1425 755 1455
rect 715 1420 755 1425
rect 825 1450 865 1460
rect 825 1430 835 1450
rect 855 1430 865 1450
rect 825 1420 865 1430
rect 885 1450 915 1460
rect 885 1430 890 1450
rect 910 1430 915 1450
rect 885 1420 915 1430
rect 935 1455 975 1460
rect 935 1425 940 1455
rect 970 1425 975 1455
rect 935 1420 975 1425
rect 1045 1450 1085 1460
rect 1045 1430 1055 1450
rect 1075 1430 1085 1450
rect 1045 1420 1085 1430
rect 1155 1455 1195 1460
rect 1155 1425 1160 1455
rect 1190 1425 1195 1455
rect 1155 1420 1195 1425
rect 1265 1450 1305 1460
rect 1265 1430 1275 1450
rect 1295 1430 1305 1450
rect 1265 1420 1305 1430
rect 1375 1455 1415 1460
rect 1375 1425 1380 1455
rect 1410 1425 1415 1455
rect 1805 1455 1810 1485
rect 1840 1455 1845 1485
rect 1805 1450 1845 1455
rect 1375 1420 1415 1425
rect 395 1405 415 1420
rect 615 1405 635 1420
rect 835 1405 855 1420
rect 385 1400 425 1405
rect 385 1370 390 1400
rect 420 1370 425 1400
rect 385 1365 425 1370
rect 585 1400 645 1405
rect 585 1370 610 1400
rect 640 1370 645 1400
rect 585 1365 645 1370
rect 825 1400 865 1405
rect 825 1370 830 1400
rect 860 1370 865 1400
rect 825 1365 865 1370
rect 585 1315 605 1365
rect 115 1310 155 1315
rect 115 1280 120 1310
rect 150 1280 155 1310
rect 115 1275 155 1280
rect 215 1310 255 1315
rect 215 1280 220 1310
rect 250 1280 255 1310
rect 215 1275 255 1280
rect 325 1310 365 1315
rect 325 1280 330 1310
rect 360 1280 365 1310
rect 325 1275 365 1280
rect 435 1310 475 1315
rect 435 1280 440 1310
rect 470 1280 475 1310
rect 435 1275 475 1280
rect 545 1310 605 1315
rect 545 1280 550 1310
rect 580 1280 605 1310
rect 545 1275 605 1280
rect 120 1260 140 1275
rect 225 1260 245 1275
rect 335 1260 355 1275
rect 445 1260 465 1275
rect 555 1260 575 1275
rect 71 1255 101 1260
rect 71 1220 101 1225
rect 120 1250 150 1260
rect 120 1230 125 1250
rect 145 1230 150 1250
rect 120 1220 150 1230
rect 220 1250 250 1260
rect 220 1230 225 1250
rect 245 1230 250 1250
rect 220 1220 250 1230
rect 275 1255 305 1260
rect 275 1220 305 1225
rect 330 1250 360 1260
rect 330 1230 335 1250
rect 355 1230 360 1250
rect 330 1220 360 1230
rect 440 1250 470 1260
rect 440 1230 445 1250
rect 465 1230 470 1250
rect 440 1220 470 1230
rect 495 1255 525 1260
rect 495 1220 525 1225
rect 550 1250 580 1260
rect 550 1230 555 1250
rect 575 1230 580 1250
rect 550 1220 580 1230
rect -155 1195 -115 1200
rect -155 1165 -150 1195
rect -120 1165 -115 1195
rect -155 1160 -115 1165
rect -45 1195 -5 1200
rect -45 1165 -40 1195
rect -10 1165 -5 1195
rect -45 1160 -5 1165
rect -200 770 -160 775
rect -200 740 -195 770
rect -165 740 -160 770
rect -200 735 -160 740
rect -190 -140 -170 735
rect -145 675 -125 1160
rect 204 1136 234 1141
rect 50 1125 90 1135
rect 50 1105 60 1125
rect 80 1105 90 1125
rect 50 1095 90 1105
rect 145 1125 185 1135
rect 145 1105 155 1125
rect 175 1105 185 1125
rect 145 1095 185 1105
rect 424 1136 454 1141
rect 204 1101 234 1106
rect 270 1125 310 1135
rect 270 1105 280 1125
rect 300 1105 310 1125
rect 270 1095 310 1105
rect 365 1125 405 1135
rect 365 1105 375 1125
rect 395 1105 405 1125
rect 365 1095 405 1105
rect 566 1136 596 1141
rect 424 1101 454 1106
rect 490 1125 530 1135
rect 490 1105 500 1125
rect 520 1105 530 1125
rect 490 1095 530 1105
rect 566 1101 596 1106
rect 615 1125 645 1135
rect 615 1105 620 1125
rect 640 1105 645 1125
rect 615 1095 645 1105
rect 60 1080 80 1095
rect 165 1080 185 1095
rect 280 1080 300 1095
rect 385 1080 405 1095
rect 500 1080 520 1095
rect 615 1080 635 1095
rect 890 1080 910 1420
rect 1055 1405 1075 1420
rect 1045 1400 1085 1405
rect 1045 1370 1050 1400
rect 1080 1370 1085 1400
rect 1045 1365 1085 1370
rect 1155 1315 1175 1420
rect 1275 1405 1295 1420
rect 1265 1400 1305 1405
rect 1265 1370 1270 1400
rect 1300 1370 1305 1400
rect 1265 1365 1305 1370
rect 1115 1310 1175 1315
rect 1115 1280 1120 1310
rect 1150 1280 1175 1310
rect 1115 1275 1175 1280
rect 1215 1310 1255 1315
rect 1215 1280 1220 1310
rect 1250 1280 1255 1310
rect 1215 1275 1255 1280
rect 1325 1310 1365 1315
rect 1325 1280 1330 1310
rect 1360 1280 1365 1310
rect 1325 1275 1365 1280
rect 1435 1310 1475 1315
rect 1435 1280 1440 1310
rect 1470 1280 1475 1310
rect 1435 1275 1475 1280
rect 1545 1310 1585 1315
rect 1545 1280 1550 1310
rect 1580 1280 1585 1310
rect 1545 1275 1585 1280
rect 1120 1260 1140 1275
rect 1225 1260 1245 1275
rect 1335 1260 1355 1275
rect 1445 1260 1465 1275
rect 1555 1260 1575 1275
rect 1071 1255 1101 1260
rect 1071 1220 1101 1225
rect 1120 1250 1150 1260
rect 1120 1230 1125 1250
rect 1145 1230 1150 1250
rect 1120 1220 1150 1230
rect 1220 1250 1250 1260
rect 1220 1230 1225 1250
rect 1245 1230 1250 1250
rect 1220 1220 1250 1230
rect 1275 1255 1305 1260
rect 1275 1220 1305 1225
rect 1330 1250 1360 1260
rect 1330 1230 1335 1250
rect 1355 1230 1360 1250
rect 1330 1220 1360 1230
rect 1440 1250 1470 1260
rect 1440 1230 1445 1250
rect 1465 1230 1470 1250
rect 1440 1220 1470 1230
rect 1495 1255 1525 1260
rect 1495 1220 1525 1225
rect 1550 1250 1580 1260
rect 1550 1230 1555 1250
rect 1575 1230 1580 1250
rect 1550 1220 1580 1230
rect 1815 1200 1835 1450
rect 1895 1255 1935 1260
rect 1895 1225 1900 1255
rect 1930 1225 1935 1255
rect 1895 1220 1935 1225
rect 1695 1195 1735 1200
rect 1695 1165 1700 1195
rect 1730 1165 1735 1195
rect 1695 1160 1735 1165
rect 1805 1195 1845 1200
rect 1805 1165 1810 1195
rect 1840 1165 1845 1195
rect 1805 1160 1845 1165
rect 1204 1136 1234 1141
rect 1050 1125 1090 1135
rect 1050 1105 1060 1125
rect 1080 1105 1090 1125
rect 1050 1095 1090 1105
rect 1145 1125 1185 1135
rect 1145 1105 1155 1125
rect 1175 1105 1185 1125
rect 1145 1095 1185 1105
rect 1424 1136 1454 1141
rect 1204 1101 1234 1106
rect 1270 1125 1310 1135
rect 1270 1105 1280 1125
rect 1300 1105 1310 1125
rect 1270 1095 1310 1105
rect 1365 1125 1405 1135
rect 1365 1105 1375 1125
rect 1395 1105 1405 1125
rect 1365 1095 1405 1105
rect 1566 1136 1596 1141
rect 1424 1101 1454 1106
rect 1490 1125 1530 1135
rect 1490 1105 1500 1125
rect 1520 1105 1530 1125
rect 1490 1095 1530 1105
rect 1566 1101 1596 1106
rect 1615 1125 1645 1135
rect 1615 1105 1620 1125
rect 1640 1105 1645 1125
rect 1615 1095 1645 1105
rect 1060 1080 1080 1095
rect 50 1075 90 1080
rect 50 1045 55 1075
rect 85 1045 90 1075
rect 50 1040 90 1045
rect 160 1075 200 1080
rect 160 1045 165 1075
rect 195 1045 200 1075
rect 160 1040 200 1045
rect 270 1075 310 1080
rect 270 1045 275 1075
rect 305 1045 310 1075
rect 270 1040 310 1045
rect 380 1075 420 1080
rect 380 1045 385 1075
rect 415 1045 420 1075
rect 380 1040 420 1045
rect 490 1075 530 1080
rect 490 1045 495 1075
rect 525 1045 530 1075
rect 490 1040 530 1045
rect 600 1075 640 1080
rect 600 1045 605 1075
rect 635 1045 640 1075
rect 600 1040 640 1045
rect 880 1075 920 1080
rect 880 1045 885 1075
rect 915 1045 920 1075
rect 880 1040 920 1045
rect 1050 1075 1090 1080
rect 1050 1045 1055 1075
rect 1085 1045 1090 1075
rect 1050 1040 1090 1045
rect 550 1020 590 1025
rect 550 990 555 1020
rect 585 990 590 1020
rect 1060 990 1080 1040
rect 1165 1035 1185 1095
rect 1280 1080 1300 1095
rect 1270 1075 1310 1080
rect 1270 1045 1275 1075
rect 1305 1045 1310 1075
rect 1270 1040 1310 1045
rect 1385 1035 1405 1095
rect 1500 1080 1520 1095
rect 1490 1075 1530 1080
rect 1490 1045 1495 1075
rect 1525 1045 1530 1075
rect 1490 1040 1530 1045
rect 1615 1035 1635 1095
rect 1160 1030 1200 1035
rect 1160 1000 1165 1030
rect 1195 1000 1200 1030
rect 1160 995 1200 1000
rect 1380 1030 1420 1035
rect 1380 1000 1385 1030
rect 1415 1000 1420 1030
rect 1380 995 1420 1000
rect 1600 1030 1640 1035
rect 1600 1000 1605 1030
rect 1635 1000 1640 1030
rect 1600 995 1640 1000
rect 550 985 590 990
rect 660 985 700 990
rect 560 935 580 985
rect 660 955 665 985
rect 695 955 700 985
rect 660 950 700 955
rect 880 985 920 990
rect 880 955 885 985
rect 915 955 920 985
rect 880 950 920 955
rect 1040 985 1080 990
rect 1040 955 1045 985
rect 1075 955 1080 985
rect 1040 950 1080 955
rect 1100 985 1140 990
rect 1100 955 1105 985
rect 1135 955 1140 985
rect 1100 950 1140 955
rect 670 935 690 950
rect 890 935 910 950
rect 1110 935 1130 950
rect 550 930 590 935
rect 550 900 555 930
rect 585 900 590 930
rect 550 895 590 900
rect 660 925 700 935
rect 660 905 670 925
rect 690 905 700 925
rect 660 895 700 905
rect 770 930 810 935
rect 770 900 775 930
rect 805 900 810 930
rect 770 895 810 900
rect 880 925 920 935
rect 880 905 890 925
rect 910 905 920 925
rect 880 895 920 905
rect 990 930 1030 935
rect 990 900 995 930
rect 1025 900 1030 930
rect 990 895 1030 900
rect 1100 925 1140 935
rect 1100 905 1110 925
rect 1130 905 1140 925
rect 1100 895 1140 905
rect 1760 930 1800 935
rect 1760 900 1765 930
rect 1795 900 1800 930
rect 1760 895 1800 900
rect 495 810 535 815
rect 495 780 500 810
rect 530 780 535 810
rect 495 775 535 780
rect 605 810 645 815
rect 605 780 610 810
rect 640 780 645 810
rect 605 775 645 780
rect 715 810 755 815
rect 715 780 720 810
rect 750 780 755 810
rect 715 775 755 780
rect 825 810 865 815
rect 825 780 830 810
rect 860 780 865 810
rect 825 775 865 780
rect 935 810 975 815
rect 935 780 940 810
rect 970 780 975 810
rect 935 775 975 780
rect 1045 810 1085 815
rect 1045 780 1050 810
rect 1080 780 1085 810
rect 1045 775 1085 780
rect 1155 810 1195 815
rect 1155 780 1160 810
rect 1190 780 1195 810
rect 1155 775 1195 780
rect 30 715 70 720
rect 30 685 35 715
rect 65 685 70 715
rect 30 680 70 685
rect 140 715 180 720
rect 140 685 145 715
rect 175 685 180 715
rect 140 680 180 685
rect 250 715 290 720
rect 250 685 255 715
rect 285 685 290 715
rect 250 680 290 685
rect 360 715 400 720
rect 360 685 365 715
rect 395 685 400 715
rect 360 680 400 685
rect 470 715 510 720
rect 470 685 475 715
rect 505 685 510 715
rect 470 680 510 685
rect 580 715 620 720
rect 580 685 585 715
rect 615 685 620 715
rect 580 680 620 685
rect 1070 715 1110 720
rect 1070 685 1075 715
rect 1105 685 1110 715
rect 1070 680 1110 685
rect 1180 715 1220 720
rect 1180 685 1185 715
rect 1215 685 1220 715
rect 1180 680 1220 685
rect 1290 715 1330 720
rect 1290 685 1295 715
rect 1325 685 1330 715
rect 1290 680 1330 685
rect 1400 715 1440 720
rect 1400 685 1405 715
rect 1435 685 1440 715
rect 1400 680 1440 685
rect 1510 715 1550 720
rect 1510 685 1515 715
rect 1545 685 1550 715
rect 1510 680 1550 685
rect 1620 715 1660 720
rect 1620 685 1625 715
rect 1655 685 1660 715
rect 1620 680 1660 685
rect -155 670 -115 675
rect -155 640 -150 670
rect -120 640 -115 670
rect 40 665 60 680
rect 150 665 170 680
rect 260 665 280 680
rect 370 665 390 680
rect 480 665 500 680
rect 590 665 610 680
rect 1080 665 1100 680
rect 1190 665 1210 680
rect 1300 665 1320 680
rect 1410 665 1430 680
rect 1520 665 1540 680
rect 1630 665 1650 680
rect -155 635 -115 640
rect -100 660 -60 665
rect -145 -85 -125 635
rect -100 630 -95 660
rect -65 630 -60 660
rect -100 625 -60 630
rect 30 655 70 665
rect 30 635 40 655
rect 60 635 70 655
rect 30 625 70 635
rect 140 655 180 665
rect 140 635 150 655
rect 170 635 180 655
rect 140 625 180 635
rect 250 655 290 665
rect 250 635 260 655
rect 280 635 290 655
rect 250 625 290 635
rect 310 660 340 665
rect 310 625 340 630
rect 360 655 400 665
rect 360 635 370 655
rect 390 635 400 655
rect 360 625 400 635
rect 470 655 510 665
rect 470 635 480 655
rect 500 635 510 655
rect 470 625 510 635
rect 580 655 620 665
rect 580 635 590 655
rect 610 635 620 655
rect 580 625 620 635
rect 1070 655 1110 665
rect 1070 635 1080 655
rect 1100 635 1110 655
rect 1070 625 1110 635
rect 1180 655 1220 665
rect 1180 635 1190 655
rect 1210 635 1220 655
rect 1180 625 1220 635
rect 1290 655 1330 665
rect 1290 635 1300 655
rect 1320 635 1330 655
rect 1290 625 1330 635
rect 1350 660 1380 665
rect 1350 625 1380 630
rect 1400 655 1440 665
rect 1400 635 1410 655
rect 1430 635 1440 655
rect 1400 625 1440 635
rect 1510 655 1550 665
rect 1510 635 1520 655
rect 1540 635 1550 655
rect 1510 625 1550 635
rect 1620 655 1660 665
rect 1620 635 1630 655
rect 1650 635 1660 655
rect 1620 625 1660 635
rect -155 -90 -115 -85
rect -155 -120 -150 -90
rect -120 -120 -115 -90
rect -155 -125 -115 -120
rect -200 -145 -160 -140
rect -200 -175 -195 -145
rect -165 -175 -160 -145
rect -1410 -225 -1375 -220
rect -245 -220 -240 -190
rect -210 -220 -205 -190
rect -245 -225 -205 -220
rect -1210 -240 -1175 -235
rect -1210 -275 -1175 -270
rect -625 -240 -585 -235
rect -625 -270 -620 -240
rect -590 -270 -585 -240
rect -625 -275 -585 -270
rect -1540 -300 -1500 -295
rect -1540 -330 -1535 -300
rect -1505 -330 -1500 -300
rect -1540 -335 -1500 -330
rect -1205 -380 -1180 -275
rect -615 -295 -595 -275
rect -1150 -300 -1115 -295
rect -1150 -335 -1115 -330
rect -925 -300 -885 -295
rect -925 -330 -920 -300
rect -890 -330 -885 -300
rect -925 -335 -885 -330
rect -725 -300 -685 -295
rect -725 -330 -720 -300
rect -690 -330 -685 -300
rect -725 -335 -685 -330
rect -625 -305 -585 -295
rect -625 -325 -615 -305
rect -595 -325 -585 -305
rect -625 -335 -585 -325
rect -525 -300 -485 -295
rect -525 -330 -520 -300
rect -490 -330 -485 -300
rect -525 -335 -485 -330
rect -1145 -380 -1120 -335
rect -1210 -415 -1206 -380
rect -1179 -415 -1175 -380
rect -1150 -415 -1146 -380
rect -1119 -415 -1115 -380
rect -190 -1070 -170 -175
rect -100 -765 -80 625
rect -25 435 15 440
rect -25 405 -20 435
rect 10 405 15 435
rect -25 400 15 405
rect 85 430 125 440
rect 85 410 95 430
rect 115 410 125 430
rect 85 400 125 410
rect 195 430 235 440
rect 195 410 205 430
rect 225 410 235 430
rect 195 400 235 410
rect 305 430 345 440
rect 305 410 315 430
rect 335 410 345 430
rect 305 400 345 410
rect 415 430 455 440
rect 415 410 425 430
rect 445 410 455 430
rect 415 400 455 410
rect 525 430 565 440
rect 525 410 535 430
rect 555 410 565 430
rect 525 400 565 410
rect 635 435 675 440
rect 635 405 640 435
rect 670 405 675 435
rect 635 400 675 405
rect 1015 435 1055 440
rect 1015 405 1020 435
rect 1050 405 1055 435
rect 1015 400 1055 405
rect 1125 430 1165 440
rect 1125 410 1135 430
rect 1155 410 1165 430
rect 1125 400 1165 410
rect 1235 430 1275 440
rect 1235 410 1245 430
rect 1265 410 1275 430
rect 1235 400 1275 410
rect 1345 430 1385 440
rect 1345 410 1355 430
rect 1375 410 1385 430
rect 1345 400 1385 410
rect 1455 430 1495 440
rect 1455 410 1465 430
rect 1485 410 1495 430
rect 1455 400 1495 410
rect 1565 430 1605 440
rect 1565 410 1575 430
rect 1595 410 1605 430
rect 1565 400 1605 410
rect 1675 435 1715 440
rect 1675 405 1680 435
rect 1710 405 1715 435
rect 1675 400 1715 405
rect 95 380 115 400
rect 205 380 225 400
rect 315 380 335 400
rect 425 380 445 400
rect 535 380 555 400
rect 1135 380 1155 400
rect 1245 380 1265 400
rect 1355 380 1375 400
rect 1465 380 1485 400
rect 1575 380 1595 400
rect 85 375 125 380
rect 85 345 90 375
rect 120 345 125 375
rect 85 340 125 345
rect 195 375 235 380
rect 195 345 200 375
rect 230 345 235 375
rect 195 340 235 345
rect 305 375 345 380
rect 305 345 310 375
rect 340 345 345 375
rect 305 340 345 345
rect 415 375 455 380
rect 415 345 420 375
rect 450 345 455 375
rect 415 340 455 345
rect 525 375 565 380
rect 525 345 530 375
rect 560 345 565 375
rect 525 340 565 345
rect 1125 375 1165 380
rect 1125 345 1130 375
rect 1160 345 1165 375
rect 1125 340 1165 345
rect 1235 375 1275 380
rect 1235 345 1240 375
rect 1270 345 1275 375
rect 1235 340 1275 345
rect 1345 375 1385 380
rect 1345 345 1350 375
rect 1380 345 1385 375
rect 1345 340 1385 345
rect 1455 375 1495 380
rect 1455 345 1460 375
rect 1490 345 1495 375
rect 1455 340 1495 345
rect 1565 375 1605 380
rect 1565 345 1570 375
rect 1600 345 1605 375
rect 1565 340 1605 345
rect 315 245 335 340
rect 310 240 340 245
rect 30 230 70 235
rect 30 200 35 230
rect 65 200 70 230
rect 30 195 70 200
rect 140 230 180 235
rect 140 200 145 230
rect 175 200 180 230
rect 140 195 180 200
rect 250 230 290 235
rect 250 200 255 230
rect 285 200 290 230
rect 310 205 340 210
rect 360 230 400 235
rect 250 195 290 200
rect 360 200 365 230
rect 395 200 400 230
rect 360 195 400 200
rect 470 230 510 235
rect 470 200 475 230
rect 505 200 510 230
rect 470 195 510 200
rect 580 230 620 235
rect 580 200 585 230
rect 615 200 620 230
rect 580 195 620 200
rect 905 185 925 275
rect 1355 245 1375 340
rect 1350 240 1380 245
rect 1070 230 1110 235
rect 1070 200 1075 230
rect 1105 200 1110 230
rect 1070 195 1110 200
rect 1180 230 1220 235
rect 1180 200 1185 230
rect 1215 200 1220 230
rect 1180 195 1220 200
rect 1290 230 1330 235
rect 1290 200 1295 230
rect 1325 200 1330 230
rect 1350 205 1380 210
rect 1400 230 1440 235
rect 1290 195 1330 200
rect 1400 200 1405 230
rect 1435 200 1440 230
rect 1400 195 1440 200
rect 1510 230 1550 235
rect 1510 200 1515 230
rect 1545 200 1550 230
rect 1510 195 1550 200
rect 1620 230 1660 235
rect 1620 200 1625 230
rect 1655 200 1660 230
rect 1620 195 1660 200
rect 310 180 340 185
rect 310 145 340 150
rect 795 180 825 185
rect 795 145 825 150
rect 848 180 878 185
rect 848 145 878 150
rect 895 175 925 185
rect 895 155 900 175
rect 920 155 925 175
rect 895 145 925 155
rect 1350 180 1380 185
rect 1350 145 1380 150
rect -20 -45 10 -35
rect -20 -65 -15 -45
rect 5 -65 10 -45
rect -20 -75 10 -65
rect 85 -40 125 -35
rect 85 -70 90 -40
rect 120 -70 125 -40
rect 85 -75 125 -70
rect 195 -40 235 -35
rect 195 -70 200 -40
rect 230 -70 235 -40
rect 195 -75 235 -70
rect 305 -40 345 -35
rect 305 -70 310 -40
rect 340 -70 345 -40
rect 305 -75 345 -70
rect 415 -40 455 -35
rect 415 -70 420 -40
rect 450 -70 455 -40
rect 415 -75 455 -70
rect 525 -40 565 -35
rect 525 -70 530 -40
rect 560 -70 565 -40
rect 525 -75 565 -70
rect 680 -45 710 -35
rect 680 -65 685 -45
rect 705 -65 710 -45
rect 680 -75 710 -65
rect 775 -45 805 -35
rect 775 -65 780 -45
rect 800 -65 805 -45
rect 775 -75 805 -65
rect 830 -45 860 -35
rect 830 -65 835 -45
rect 855 -65 860 -45
rect 830 -75 860 -65
rect 885 -45 915 -35
rect 885 -65 890 -45
rect 910 -65 915 -45
rect 885 -75 915 -65
rect 980 -45 1010 -35
rect 980 -65 985 -45
rect 1005 -65 1010 -45
rect 980 -75 1010 -65
rect 1125 -40 1170 -35
rect 1125 -70 1130 -40
rect 1160 -70 1170 -40
rect 1125 -75 1170 -70
rect 1235 -40 1275 -35
rect 1235 -70 1240 -40
rect 1270 -70 1275 -40
rect 1235 -75 1275 -70
rect 1345 -40 1385 -35
rect 1345 -70 1350 -40
rect 1380 -70 1385 -40
rect 1345 -75 1385 -70
rect 1455 -40 1495 -35
rect 1455 -70 1460 -40
rect 1490 -70 1495 -40
rect 1455 -75 1495 -70
rect 1565 -40 1605 -35
rect 1565 -70 1570 -40
rect 1600 -70 1605 -40
rect 1565 -75 1605 -70
rect 1680 -45 1710 -35
rect 1680 -65 1685 -45
rect 1705 -65 1710 -45
rect 1680 -75 1710 -65
rect -15 -135 5 -75
rect 685 -135 705 -75
rect 780 -90 800 -75
rect 760 -95 800 -90
rect 760 -125 765 -95
rect 795 -125 800 -95
rect 760 -130 800 -125
rect -25 -140 15 -135
rect -25 -170 -20 -140
rect 10 -170 15 -140
rect -25 -175 15 -170
rect 675 -140 715 -135
rect 675 -170 680 -140
rect 710 -170 715 -140
rect 675 -175 715 -170
rect 75 -195 115 -190
rect 75 -225 80 -195
rect 110 -225 115 -195
rect 75 -230 115 -225
rect 710 -195 750 -190
rect 710 -225 715 -195
rect 745 -225 750 -195
rect 710 -230 750 -225
rect 85 -720 105 -230
rect 270 -295 310 -290
rect 270 -325 275 -295
rect 305 -325 310 -295
rect 270 -330 310 -325
rect 280 -345 300 -330
rect 720 -345 740 -230
rect 775 -345 795 -130
rect 835 -290 855 -75
rect 890 -90 910 -75
rect 890 -95 930 -90
rect 890 -125 895 -95
rect 925 -125 930 -95
rect 890 -130 930 -125
rect 985 -135 1005 -75
rect 975 -140 1015 -135
rect 975 -170 980 -140
rect 1010 -170 1015 -140
rect 975 -175 1015 -170
rect 825 -295 865 -290
rect 825 -325 830 -295
rect 860 -325 865 -295
rect 825 -330 865 -325
rect 1150 -345 1170 -75
rect 1685 -135 1705 -75
rect 1675 -140 1715 -135
rect 1675 -170 1680 -140
rect 1710 -170 1715 -140
rect 1675 -175 1715 -170
rect 1770 -290 1790 895
rect 1815 675 1835 1160
rect 1850 770 1890 775
rect 1850 740 1855 770
rect 1885 740 1890 770
rect 1850 735 1890 740
rect 1805 670 1845 675
rect 1805 640 1810 670
rect 1840 640 1845 670
rect 1805 635 1845 640
rect 1815 -85 1835 635
rect 1860 440 1880 735
rect 1850 435 1890 440
rect 1850 405 1855 435
rect 1885 405 1890 435
rect 1850 400 1890 405
rect 1805 -90 1845 -85
rect 1805 -120 1810 -90
rect 1840 -120 1845 -90
rect 1805 -125 1845 -120
rect 1860 -140 1880 400
rect 1850 -145 1890 -140
rect 1850 -175 1855 -145
rect 1885 -175 1890 -145
rect 1330 -295 1370 -290
rect 1330 -325 1335 -295
rect 1365 -325 1370 -295
rect 1330 -330 1370 -325
rect 1760 -295 1800 -290
rect 1760 -325 1765 -295
rect 1795 -325 1800 -295
rect 1760 -330 1800 -325
rect 1340 -345 1360 -330
rect 270 -355 310 -345
rect 270 -375 280 -355
rect 300 -375 310 -355
rect 270 -385 310 -375
rect 380 -350 420 -345
rect 380 -380 385 -350
rect 415 -380 420 -350
rect 380 -385 420 -380
rect 490 -350 530 -345
rect 490 -380 495 -350
rect 525 -380 530 -350
rect 490 -385 530 -380
rect 600 -350 640 -345
rect 600 -380 605 -350
rect 635 -380 640 -350
rect 600 -385 640 -380
rect 710 -350 750 -345
rect 710 -380 715 -350
rect 745 -380 750 -350
rect 710 -385 750 -380
rect 770 -355 800 -345
rect 770 -375 775 -355
rect 795 -375 800 -355
rect 770 -385 800 -375
rect 820 -350 860 -345
rect 820 -380 825 -350
rect 855 -380 860 -350
rect 820 -385 860 -380
rect 930 -350 970 -345
rect 930 -380 935 -350
rect 965 -380 970 -350
rect 930 -385 970 -380
rect 1040 -350 1080 -345
rect 1040 -380 1045 -350
rect 1075 -380 1080 -350
rect 1040 -385 1080 -380
rect 1150 -350 1190 -345
rect 1150 -380 1155 -350
rect 1185 -380 1190 -350
rect 1150 -385 1190 -380
rect 1260 -350 1300 -345
rect 1260 -380 1265 -350
rect 1295 -380 1300 -350
rect 1260 -385 1300 -380
rect 1336 -355 1366 -345
rect 1336 -375 1341 -355
rect 1361 -375 1366 -355
rect 1336 -385 1366 -375
rect 1385 -350 1425 -345
rect 1385 -380 1390 -350
rect 1420 -380 1425 -350
rect 1385 -385 1425 -380
rect 1860 -670 1880 -175
rect 1905 -190 1925 1220
rect 1950 720 1970 1635
rect 2385 1630 2405 1690
rect 2375 1625 2415 1630
rect 2375 1595 2380 1625
rect 2410 1595 2415 1625
rect 2375 1590 2415 1595
rect 3100 1490 3140 1495
rect 2045 1485 2085 1490
rect 2045 1455 2050 1485
rect 2080 1455 2085 1485
rect 2045 1450 2085 1455
rect 2155 1485 2195 1490
rect 2155 1455 2160 1485
rect 2190 1455 2195 1485
rect 2155 1450 2195 1455
rect 2265 1485 2305 1490
rect 2265 1455 2270 1485
rect 2300 1455 2305 1485
rect 2265 1450 2305 1455
rect 2375 1485 2415 1490
rect 2375 1455 2380 1485
rect 2410 1455 2415 1485
rect 2375 1450 2415 1455
rect 2485 1485 2525 1490
rect 2485 1455 2490 1485
rect 2520 1455 2525 1485
rect 2485 1450 2525 1455
rect 2595 1485 2635 1490
rect 2595 1455 2600 1485
rect 2630 1455 2635 1485
rect 2595 1450 2635 1455
rect 2705 1485 2745 1490
rect 2705 1455 2710 1485
rect 2740 1455 2745 1485
rect 3100 1460 3105 1490
rect 3135 1460 3140 1490
rect 3100 1455 3140 1460
rect 2705 1450 2745 1455
rect 3110 1430 3130 1455
rect 3050 1420 3191 1430
rect 3050 1400 3055 1420
rect 3075 1400 3110 1420
rect 3130 1400 3165 1420
rect 3185 1400 3191 1420
rect 3050 1390 3191 1400
rect 3050 815 3191 825
rect 2100 810 2140 815
rect 2100 780 2105 810
rect 2135 780 2140 810
rect 2100 775 2140 780
rect 2210 810 2250 815
rect 2210 780 2215 810
rect 2245 780 2250 810
rect 2210 775 2250 780
rect 2320 810 2360 815
rect 2430 810 2470 815
rect 2320 780 2325 810
rect 2355 780 2360 810
rect 2320 775 2360 780
rect 2380 800 2410 810
rect 2380 780 2385 800
rect 2405 780 2410 800
rect 2380 770 2410 780
rect 2430 780 2435 810
rect 2465 780 2470 810
rect 2430 775 2470 780
rect 2540 810 2580 815
rect 2540 780 2545 810
rect 2575 780 2580 810
rect 2540 775 2580 780
rect 2650 810 2690 815
rect 2650 780 2655 810
rect 2685 780 2690 810
rect 3050 795 3055 815
rect 3075 795 3110 815
rect 3130 795 3165 815
rect 3185 795 3191 815
rect 3050 785 3191 795
rect 2650 775 2690 780
rect 2100 730 2105 760
rect 2135 730 2140 760
rect 1940 715 1980 720
rect 1940 685 1945 715
rect 1975 685 1980 715
rect 1940 680 1980 685
rect 1950 345 1970 680
rect 2110 675 2130 730
rect 2385 720 2405 770
rect 2550 760 2570 775
rect 2540 730 2545 760
rect 2575 730 2580 760
rect 3110 720 3130 785
rect 3190 760 3230 765
rect 3190 730 3195 760
rect 3225 730 3230 760
rect 3190 725 3230 730
rect 2375 715 2415 720
rect 2375 685 2380 715
rect 2410 685 2415 715
rect 2375 680 2415 685
rect 3100 715 3140 720
rect 3100 685 3105 715
rect 3135 685 3140 715
rect 3100 680 3140 685
rect 2035 670 2075 675
rect 2035 640 2040 670
rect 2070 640 2075 670
rect 2035 635 2075 640
rect 2100 670 2140 675
rect 2100 640 2105 670
rect 2135 640 2140 670
rect 2100 635 2140 640
rect 2210 670 2250 675
rect 2210 640 2215 670
rect 2245 640 2250 670
rect 2210 635 2250 640
rect 2320 670 2360 675
rect 2320 640 2325 670
rect 2355 640 2360 670
rect 2320 635 2360 640
rect 2430 670 2470 675
rect 2430 640 2435 670
rect 2465 640 2470 670
rect 2430 635 2470 640
rect 2540 670 2580 675
rect 2540 640 2545 670
rect 2575 640 2580 670
rect 2540 635 2580 640
rect 2650 670 2690 675
rect 2650 640 2655 670
rect 2685 640 2690 670
rect 2650 635 2690 640
rect 2715 670 2755 675
rect 2715 640 2720 670
rect 2750 640 2755 670
rect 2715 635 2755 640
rect 2155 395 2195 400
rect 2155 365 2160 395
rect 2190 365 2195 395
rect 2155 360 2195 365
rect 2265 395 2305 400
rect 2265 365 2270 395
rect 2300 365 2305 395
rect 2265 360 2305 365
rect 2325 390 2355 400
rect 2325 370 2330 390
rect 2350 370 2355 390
rect 2325 360 2355 370
rect 2375 395 2415 400
rect 2375 365 2380 395
rect 2410 365 2415 395
rect 2375 360 2415 365
rect 2485 395 2525 400
rect 2485 365 2490 395
rect 2520 365 2525 395
rect 2485 360 2525 365
rect 2595 395 2635 400
rect 2595 365 2600 395
rect 2630 365 2635 395
rect 2595 360 2635 365
rect 2840 395 2880 400
rect 2840 365 2845 395
rect 2875 365 2880 395
rect 2840 360 2880 365
rect 3200 360 3220 725
rect 2330 345 2350 360
rect 1940 340 1980 345
rect 1940 310 1945 340
rect 1975 310 1980 340
rect 1940 305 1980 310
rect 2320 340 2360 345
rect 2320 310 2325 340
rect 2355 310 2360 340
rect 2320 305 2360 310
rect 2330 290 2350 305
rect 2155 285 2195 290
rect 2155 255 2160 285
rect 2190 255 2195 285
rect 2155 250 2195 255
rect 2265 285 2305 290
rect 2265 255 2270 285
rect 2300 255 2305 285
rect 2265 250 2305 255
rect 2325 280 2355 290
rect 2325 260 2330 280
rect 2350 260 2355 280
rect 2325 250 2355 260
rect 2375 285 2415 290
rect 2375 255 2380 285
rect 2410 255 2415 285
rect 2375 250 2415 255
rect 2485 285 2525 290
rect 2485 255 2490 285
rect 2520 255 2525 285
rect 2485 250 2525 255
rect 2595 285 2635 290
rect 2595 255 2600 285
rect 2630 255 2635 285
rect 2595 250 2635 255
rect 2795 285 2835 290
rect 2795 255 2800 285
rect 2830 255 2835 285
rect 2795 250 2835 255
rect 2805 -85 2825 250
rect 2035 -95 2075 -85
rect 2035 -115 2045 -95
rect 2065 -115 2075 -95
rect 2035 -125 2075 -115
rect 2100 -90 2140 -85
rect 2100 -120 2105 -90
rect 2135 -120 2140 -90
rect 2100 -125 2140 -120
rect 2210 -90 2250 -85
rect 2210 -120 2215 -90
rect 2245 -120 2250 -90
rect 2210 -125 2250 -120
rect 2320 -90 2360 -85
rect 2320 -120 2325 -90
rect 2355 -120 2360 -90
rect 2320 -125 2360 -120
rect 2430 -90 2470 -85
rect 2430 -120 2435 -90
rect 2465 -120 2470 -90
rect 2430 -125 2470 -120
rect 2540 -90 2580 -85
rect 2540 -120 2545 -90
rect 2575 -120 2580 -90
rect 2540 -125 2580 -120
rect 2650 -90 2690 -85
rect 2650 -120 2655 -90
rect 2685 -120 2690 -90
rect 2650 -125 2690 -120
rect 2715 -95 2755 -85
rect 2715 -115 2725 -95
rect 2745 -115 2755 -95
rect 2715 -125 2755 -115
rect 2795 -90 2835 -85
rect 2795 -120 2800 -90
rect 2830 -120 2835 -90
rect 2795 -125 2835 -120
rect 2045 -140 2065 -125
rect 2725 -140 2745 -125
rect 2850 -140 2870 360
rect 3185 350 3235 360
rect 3185 320 3195 350
rect 3225 320 3235 350
rect 3185 310 3235 320
rect 2885 -120 2889 -85
rect 2916 -120 2920 -85
rect 2945 -120 2949 -85
rect 2976 -120 2980 -85
rect 3005 -120 3009 -85
rect 3036 -120 3040 -85
rect 3065 -120 3069 -85
rect 3096 -120 3100 -85
rect 2035 -145 2075 -140
rect 2035 -175 2040 -145
rect 2070 -175 2075 -145
rect 2035 -180 2075 -175
rect 2715 -145 2755 -140
rect 2715 -175 2720 -145
rect 2750 -175 2755 -145
rect 2715 -180 2755 -175
rect 2840 -145 2880 -140
rect 2840 -175 2845 -145
rect 2875 -175 2880 -145
rect 2840 -180 2880 -175
rect 2945 -145 2980 -120
rect 2945 -180 2980 -175
rect 3070 -185 3095 -120
rect 3065 -190 3100 -185
rect 1895 -220 1900 -190
rect 1930 -220 1935 -190
rect 1895 -225 1935 -220
rect 3065 -225 3100 -220
rect 2275 -240 2315 -235
rect 2275 -270 2280 -240
rect 2310 -270 2315 -240
rect 2275 -275 2315 -270
rect 2865 -240 2900 -235
rect 2865 -275 2900 -270
rect 2285 -295 2305 -275
rect 2175 -300 2215 -295
rect 2175 -330 2180 -300
rect 2210 -330 2215 -300
rect 2175 -335 2215 -330
rect 2275 -305 2315 -295
rect 2275 -325 2285 -305
rect 2305 -325 2315 -305
rect 2275 -335 2315 -325
rect 2375 -300 2415 -295
rect 2375 -330 2380 -300
rect 2410 -330 2415 -300
rect 2375 -335 2415 -330
rect 2575 -300 2615 -295
rect 2575 -330 2580 -300
rect 2610 -330 2615 -300
rect 2575 -335 2615 -330
rect 2805 -300 2840 -295
rect 2805 -335 2840 -330
rect 2810 -380 2835 -335
rect 2870 -380 2895 -275
rect 3200 -295 3220 310
rect 3190 -300 3230 -295
rect 3190 -330 3195 -300
rect 3225 -330 3230 -300
rect 3190 -335 3230 -330
rect 2805 -415 2809 -380
rect 2836 -415 2840 -380
rect 2865 -415 2869 -380
rect 2896 -415 2900 -380
rect 150 -675 190 -670
rect 150 -705 155 -675
rect 185 -705 190 -675
rect 150 -710 190 -705
rect 215 -675 255 -670
rect 215 -705 220 -675
rect 250 -705 255 -675
rect 215 -710 255 -705
rect 325 -675 365 -670
rect 325 -705 330 -675
rect 360 -705 365 -675
rect 325 -710 365 -705
rect 435 -675 475 -670
rect 435 -705 440 -675
rect 470 -705 475 -675
rect 435 -710 475 -705
rect 545 -675 585 -670
rect 545 -705 550 -675
rect 580 -705 585 -675
rect 545 -710 585 -705
rect 655 -675 695 -670
rect 655 -705 660 -675
rect 690 -705 695 -675
rect 655 -710 695 -705
rect 765 -675 805 -670
rect 765 -705 770 -675
rect 800 -705 805 -675
rect 765 -710 805 -705
rect 875 -675 915 -670
rect 875 -705 880 -675
rect 910 -705 915 -675
rect 875 -710 915 -705
rect 985 -675 1025 -670
rect 985 -705 990 -675
rect 1020 -705 1025 -675
rect 985 -710 1025 -705
rect 1095 -675 1135 -670
rect 1095 -705 1100 -675
rect 1130 -705 1135 -675
rect 1095 -710 1135 -705
rect 1205 -675 1245 -670
rect 1205 -705 1210 -675
rect 1240 -705 1245 -675
rect 1205 -710 1245 -705
rect 1315 -675 1355 -670
rect 1315 -705 1320 -675
rect 1350 -705 1355 -675
rect 1315 -710 1355 -705
rect 1425 -675 1465 -670
rect 1425 -705 1430 -675
rect 1460 -705 1465 -675
rect 1425 -710 1465 -705
rect 1850 -675 1890 -670
rect 1850 -705 1855 -675
rect 1885 -705 1890 -675
rect 1850 -710 1890 -705
rect 75 -725 115 -720
rect 75 -755 80 -725
rect 110 -755 115 -725
rect 75 -760 115 -755
rect 1010 -735 1050 -730
rect 1010 -765 1015 -735
rect 1045 -765 1050 -735
rect -110 -770 -70 -765
rect -110 -800 -105 -770
rect -75 -800 -70 -770
rect -110 -805 -70 -800
rect 710 -770 750 -765
rect 710 -800 715 -770
rect 745 -800 750 -770
rect 710 -805 750 -800
rect 825 -770 865 -765
rect 825 -800 830 -770
rect 860 -800 865 -770
rect 825 -805 865 -800
rect 950 -770 990 -765
rect 1010 -770 1050 -765
rect 950 -800 955 -770
rect 985 -800 990 -770
rect 950 -805 990 -800
rect 1860 -1070 1880 -710
rect -1025 -1075 -985 -1070
rect -1025 -1105 -1020 -1075
rect -990 -1105 -985 -1075
rect -1025 -1110 -985 -1105
rect -825 -1075 -785 -1070
rect -825 -1105 -820 -1075
rect -790 -1105 -785 -1075
rect -825 -1110 -785 -1105
rect -625 -1075 -585 -1070
rect -625 -1105 -620 -1075
rect -590 -1105 -585 -1075
rect -625 -1110 -585 -1105
rect -425 -1075 -385 -1070
rect -425 -1105 -420 -1075
rect -390 -1105 -385 -1075
rect -425 -1110 -385 -1105
rect -200 -1075 -160 -1070
rect -200 -1105 -195 -1075
rect -165 -1105 -160 -1075
rect -200 -1110 -160 -1105
rect 825 -1075 865 -1070
rect 825 -1105 830 -1075
rect 860 -1105 865 -1075
rect 825 -1110 865 -1105
rect 1850 -1075 1890 -1070
rect 1850 -1105 1855 -1075
rect 1885 -1105 1890 -1075
rect 1850 -1110 1890 -1105
rect 2075 -1075 2115 -1070
rect 2075 -1105 2080 -1075
rect 2110 -1105 2115 -1075
rect 2075 -1110 2115 -1105
rect 2275 -1075 2315 -1070
rect 2275 -1105 2280 -1075
rect 2310 -1105 2315 -1075
rect 2275 -1110 2315 -1105
rect 2475 -1075 2515 -1070
rect 2475 -1105 2480 -1075
rect 2510 -1105 2515 -1075
rect 2475 -1110 2515 -1105
rect 2675 -1075 2715 -1070
rect 2675 -1105 2680 -1075
rect 2710 -1105 2715 -1075
rect 2675 -1110 2715 -1105
rect 835 -2420 855 -1110
rect 825 -2425 865 -2420
rect 825 -2455 830 -2425
rect 860 -2455 865 -2425
rect 825 -2460 865 -2455
<< via1 >>
rect 830 4245 860 4275
rect 155 2750 185 2780
rect 625 2750 655 2780
rect 35 2720 65 2725
rect 35 2700 40 2720
rect 40 2700 60 2720
rect 60 2700 65 2720
rect 35 2695 65 2700
rect 155 2720 185 2725
rect 155 2700 160 2720
rect 160 2700 180 2720
rect 180 2700 185 2720
rect 155 2695 185 2700
rect 215 2720 245 2725
rect 215 2700 220 2720
rect 220 2700 240 2720
rect 240 2700 245 2720
rect 215 2695 245 2700
rect 1035 2750 1065 2780
rect 1503 2750 1533 2780
rect 830 2695 860 2725
rect 975 2720 1005 2725
rect 975 2700 980 2720
rect 980 2700 1000 2720
rect 1000 2700 1005 2720
rect 975 2695 1005 2700
rect 1095 2720 1125 2725
rect 1095 2700 1100 2720
rect 1100 2700 1120 2720
rect 1120 2700 1125 2720
rect 1095 2695 1125 2700
rect 1155 2720 1185 2725
rect 1155 2700 1160 2720
rect 1160 2700 1180 2720
rect 1180 2700 1185 2720
rect 1155 2695 1185 2700
rect 1443 2720 1473 2725
rect 1443 2700 1448 2720
rect 1448 2700 1468 2720
rect 1468 2700 1473 2720
rect 1443 2695 1473 2700
rect 1503 2720 1533 2725
rect 1503 2700 1508 2720
rect 1508 2700 1528 2720
rect 1528 2700 1533 2720
rect 1503 2695 1533 2700
rect 1623 2720 1653 2725
rect 1623 2700 1628 2720
rect 1628 2700 1648 2720
rect 1648 2700 1653 2720
rect 1623 2695 1653 2700
rect 505 2550 535 2555
rect 505 2530 510 2550
rect 510 2530 530 2550
rect 530 2530 535 2550
rect 505 2525 535 2530
rect 565 2550 595 2555
rect 565 2530 570 2550
rect 570 2530 590 2550
rect 590 2530 595 2550
rect 565 2525 595 2530
rect 685 2550 715 2555
rect 685 2530 690 2550
rect 690 2530 710 2550
rect 710 2530 715 2550
rect 685 2525 715 2530
rect 830 2525 860 2555
rect 80 2300 110 2305
rect 80 2280 85 2300
rect 85 2280 105 2300
rect 105 2280 110 2300
rect 80 2275 110 2280
rect 139 2300 169 2305
rect 139 2280 144 2300
rect 144 2280 164 2300
rect 164 2280 169 2300
rect 139 2275 169 2280
rect 609 2300 639 2305
rect 609 2280 614 2300
rect 614 2280 634 2300
rect 634 2280 639 2300
rect 609 2275 639 2280
rect 775 2275 805 2305
rect -720 2175 -690 2205
rect -150 2175 -120 2205
rect -1080 2145 -1050 2150
rect -1080 2125 -1075 2145
rect -1075 2125 -1055 2145
rect -1055 2125 -1050 2145
rect -1080 2120 -1050 2125
rect -960 2145 -930 2150
rect -960 2125 -955 2145
rect -955 2125 -935 2145
rect -935 2125 -930 2145
rect -960 2120 -930 2125
rect -840 2145 -810 2150
rect -840 2125 -835 2145
rect -835 2125 -815 2145
rect -815 2125 -810 2145
rect -840 2120 -810 2125
rect -720 2145 -690 2150
rect -720 2125 -715 2145
rect -715 2125 -695 2145
rect -695 2125 -690 2145
rect -720 2120 -690 2125
rect -600 2145 -570 2150
rect -600 2125 -595 2145
rect -595 2125 -575 2145
rect -575 2125 -570 2145
rect -600 2120 -570 2125
rect -480 2145 -450 2150
rect -480 2125 -475 2145
rect -475 2125 -455 2145
rect -455 2125 -450 2145
rect -480 2120 -450 2125
rect -360 2145 -330 2150
rect -360 2125 -355 2145
rect -355 2125 -335 2145
rect -335 2125 -330 2145
rect -360 2120 -330 2125
rect -195 2120 -165 2150
rect -1020 1720 -990 1725
rect -1020 1700 -1015 1720
rect -1015 1700 -995 1720
rect -995 1700 -990 1720
rect -1020 1695 -990 1700
rect -900 1720 -870 1725
rect -900 1700 -895 1720
rect -895 1700 -875 1720
rect -875 1700 -870 1720
rect -900 1695 -870 1700
rect -780 1720 -750 1725
rect -780 1700 -775 1720
rect -775 1700 -755 1720
rect -755 1700 -750 1720
rect -780 1695 -750 1700
rect -660 1720 -630 1725
rect -660 1700 -655 1720
rect -655 1700 -635 1720
rect -635 1700 -630 1720
rect -660 1695 -630 1700
rect -540 1720 -510 1725
rect -540 1700 -535 1720
rect -535 1700 -515 1720
rect -515 1700 -510 1720
rect -540 1695 -510 1700
rect -420 1720 -390 1725
rect -420 1700 -415 1720
rect -415 1700 -395 1720
rect -395 1700 -390 1720
rect -420 1695 -390 1700
rect -195 1695 -165 1725
rect -285 1640 -255 1670
rect -720 1595 -690 1625
rect -1445 1510 -1415 1540
rect -1050 1480 -1020 1485
rect -1050 1460 -1045 1480
rect -1045 1460 -1025 1480
rect -1025 1460 -1020 1480
rect -1050 1455 -1020 1460
rect -940 1480 -910 1485
rect -940 1460 -935 1480
rect -935 1460 -915 1480
rect -915 1460 -910 1480
rect -940 1455 -910 1460
rect -830 1480 -800 1485
rect -830 1460 -825 1480
rect -825 1460 -805 1480
rect -805 1460 -800 1480
rect -830 1455 -800 1460
rect -720 1480 -690 1485
rect -720 1460 -715 1480
rect -715 1460 -695 1480
rect -695 1460 -690 1480
rect -720 1455 -690 1460
rect -610 1480 -580 1485
rect -610 1460 -605 1480
rect -605 1460 -585 1480
rect -585 1460 -580 1480
rect -610 1455 -580 1460
rect -500 1480 -470 1485
rect -500 1460 -495 1480
rect -495 1460 -475 1480
rect -475 1460 -470 1480
rect -500 1455 -470 1460
rect -390 1480 -360 1485
rect -390 1460 -385 1480
rect -385 1460 -365 1480
rect -365 1460 -360 1480
rect -390 1455 -360 1460
rect -1535 730 -1505 760
rect -995 805 -965 810
rect -995 785 -990 805
rect -990 785 -970 805
rect -970 785 -965 805
rect -995 780 -965 785
rect -885 805 -855 810
rect -885 785 -880 805
rect -880 785 -860 805
rect -860 785 -855 805
rect -885 780 -855 785
rect -775 805 -745 810
rect -775 785 -770 805
rect -770 785 -750 805
rect -750 785 -745 805
rect -775 780 -745 785
rect -665 805 -635 810
rect -665 785 -660 805
rect -660 785 -640 805
rect -640 785 -635 805
rect -665 780 -635 785
rect -555 805 -525 810
rect -555 785 -550 805
rect -550 785 -530 805
rect -530 785 -525 805
rect -555 780 -525 785
rect -445 805 -415 810
rect -445 785 -440 805
rect -440 785 -420 805
rect -420 785 -415 805
rect -445 780 -415 785
rect -885 730 -855 760
rect -445 730 -415 760
rect -1445 685 -1415 715
rect -720 685 -690 715
rect -35 2145 -5 2150
rect -35 2125 -30 2145
rect -30 2125 -10 2145
rect -10 2125 -5 2145
rect -35 2120 -5 2125
rect 85 2145 115 2150
rect 85 2125 90 2145
rect 90 2125 110 2145
rect 110 2125 115 2145
rect 85 2120 115 2125
rect 205 2145 235 2150
rect 205 2125 210 2145
rect 210 2125 230 2145
rect 230 2125 235 2145
rect 205 2120 235 2125
rect 325 2145 355 2150
rect 325 2125 330 2145
rect 330 2125 350 2145
rect 350 2125 355 2145
rect 325 2120 355 2125
rect 445 2145 475 2150
rect 445 2125 450 2145
rect 450 2125 470 2145
rect 470 2125 475 2145
rect 445 2120 475 2125
rect 565 2145 595 2150
rect 565 2125 570 2145
rect 570 2125 590 2145
rect 590 2125 595 2145
rect 565 2120 595 2125
rect 685 2145 715 2150
rect 685 2125 690 2145
rect 690 2125 710 2145
rect 710 2125 715 2145
rect 685 2120 715 2125
rect 25 1720 55 1725
rect 25 1700 30 1720
rect 30 1700 50 1720
rect 50 1700 55 1720
rect 25 1695 55 1700
rect 145 1720 175 1725
rect 145 1700 150 1720
rect 150 1700 170 1720
rect 170 1700 175 1720
rect 145 1695 175 1700
rect 265 1720 295 1725
rect 265 1700 270 1720
rect 270 1700 290 1720
rect 290 1700 295 1720
rect 265 1695 295 1700
rect 385 1720 415 1725
rect 385 1700 390 1720
rect 390 1700 410 1720
rect 410 1700 415 1720
rect 385 1695 415 1700
rect 505 1720 535 1725
rect 505 1700 510 1720
rect 510 1700 530 1720
rect 530 1700 535 1720
rect 505 1695 535 1700
rect 625 1720 655 1725
rect 625 1700 630 1720
rect 630 1700 650 1720
rect 650 1700 655 1720
rect 625 1695 655 1700
rect 1519 2300 1549 2305
rect 1519 2280 1524 2300
rect 1524 2280 1544 2300
rect 1544 2280 1549 2300
rect 1519 2275 1549 2280
rect 885 2230 915 2260
rect 830 2175 860 2205
rect 25 1640 55 1670
rect 325 1640 355 1670
rect 785 1640 815 1670
rect 1050 2220 1080 2250
rect 1578 2220 1608 2250
rect 1810 2175 1840 2205
rect 2380 2175 2410 2205
rect 975 2145 1005 2150
rect 975 2125 980 2145
rect 980 2125 1000 2145
rect 1000 2125 1005 2145
rect 975 2120 1005 2125
rect 1095 2145 1125 2150
rect 1095 2125 1100 2145
rect 1100 2125 1120 2145
rect 1120 2125 1125 2145
rect 1095 2120 1125 2125
rect 1215 2145 1245 2150
rect 1215 2125 1220 2145
rect 1220 2125 1240 2145
rect 1240 2125 1245 2145
rect 1215 2120 1245 2125
rect 1335 2145 1365 2150
rect 1335 2125 1340 2145
rect 1340 2125 1360 2145
rect 1360 2125 1365 2145
rect 1335 2120 1365 2125
rect 1455 2145 1485 2150
rect 1455 2125 1460 2145
rect 1460 2125 1480 2145
rect 1480 2125 1485 2145
rect 1455 2120 1485 2125
rect 1575 2145 1605 2150
rect 1575 2125 1580 2145
rect 1580 2125 1600 2145
rect 1600 2125 1605 2145
rect 1575 2120 1605 2125
rect 1695 2145 1725 2150
rect 1695 2125 1700 2145
rect 1700 2125 1720 2145
rect 1720 2125 1725 2145
rect 1695 2120 1725 2125
rect 1035 1720 1065 1725
rect 1035 1700 1040 1720
rect 1040 1700 1060 1720
rect 1060 1700 1065 1720
rect 1035 1695 1065 1700
rect 1155 1720 1185 1725
rect 1155 1700 1160 1720
rect 1160 1700 1180 1720
rect 1180 1700 1185 1720
rect 1155 1695 1185 1700
rect 1275 1720 1305 1725
rect 1275 1700 1280 1720
rect 1280 1700 1300 1720
rect 1300 1700 1305 1720
rect 1275 1695 1305 1700
rect 1395 1720 1425 1725
rect 1395 1700 1400 1720
rect 1400 1700 1420 1720
rect 1420 1700 1425 1720
rect 1395 1695 1425 1700
rect 1515 1720 1545 1725
rect 1515 1700 1520 1720
rect 1520 1700 1540 1720
rect 1540 1700 1545 1720
rect 1515 1695 1545 1700
rect 1635 1720 1665 1725
rect 1635 1700 1640 1720
rect 1640 1700 1660 1720
rect 1660 1700 1665 1720
rect 1635 1695 1665 1700
rect 1335 1640 1365 1670
rect 1635 1640 1665 1670
rect 875 1600 905 1630
rect 1855 2120 1885 2150
rect 2020 2145 2050 2150
rect 2020 2125 2025 2145
rect 2025 2125 2045 2145
rect 2045 2125 2050 2145
rect 2020 2120 2050 2125
rect 2140 2145 2170 2150
rect 2140 2125 2145 2145
rect 2145 2125 2165 2145
rect 2165 2125 2170 2145
rect 2140 2120 2170 2125
rect 2260 2145 2290 2150
rect 2260 2125 2265 2145
rect 2265 2125 2285 2145
rect 2285 2125 2290 2145
rect 2260 2120 2290 2125
rect 2380 2145 2410 2150
rect 2380 2125 2385 2145
rect 2385 2125 2405 2145
rect 2405 2125 2410 2145
rect 2380 2120 2410 2125
rect 2500 2145 2530 2150
rect 2500 2125 2505 2145
rect 2505 2125 2525 2145
rect 2525 2125 2530 2145
rect 2500 2120 2530 2125
rect 2620 2145 2650 2150
rect 2620 2125 2625 2145
rect 2625 2125 2645 2145
rect 2645 2125 2650 2145
rect 2620 2120 2650 2125
rect 2740 2145 2770 2150
rect 2740 2125 2745 2145
rect 2745 2125 2765 2145
rect 2765 2125 2770 2145
rect 2740 2120 2770 2125
rect 1855 1695 1885 1725
rect 2080 1720 2110 1725
rect 2080 1700 2085 1720
rect 2085 1700 2105 1720
rect 2105 1700 2110 1720
rect 2080 1695 2110 1700
rect 2200 1720 2230 1725
rect 2200 1700 2205 1720
rect 2205 1700 2225 1720
rect 2225 1700 2230 1720
rect 2200 1695 2230 1700
rect 2320 1720 2350 1725
rect 2320 1700 2325 1720
rect 2325 1700 2345 1720
rect 2345 1700 2350 1720
rect 2320 1695 2350 1700
rect 2440 1720 2470 1725
rect 2440 1700 2445 1720
rect 2445 1700 2465 1720
rect 2465 1700 2470 1720
rect 2440 1695 2470 1700
rect 2560 1720 2590 1725
rect 2560 1700 2565 1720
rect 2565 1700 2585 1720
rect 2585 1700 2590 1720
rect 2560 1695 2590 1700
rect 2680 1720 2710 1725
rect 2680 1700 2685 1720
rect 2685 1700 2705 1720
rect 2705 1700 2710 1720
rect 2680 1695 2710 1700
rect 1945 1640 1975 1670
rect 225 1575 255 1580
rect 225 1555 230 1575
rect 230 1555 250 1575
rect 250 1555 255 1575
rect 225 1550 255 1555
rect 335 1575 365 1580
rect 335 1555 340 1575
rect 340 1555 360 1575
rect 360 1555 365 1575
rect 335 1550 365 1555
rect 445 1575 475 1580
rect 445 1555 450 1575
rect 450 1555 470 1575
rect 470 1555 475 1575
rect 445 1550 475 1555
rect 555 1575 585 1580
rect 555 1555 560 1575
rect 560 1555 580 1575
rect 580 1555 585 1575
rect 555 1550 585 1555
rect 665 1575 695 1580
rect 665 1555 670 1575
rect 670 1555 690 1575
rect 690 1555 695 1575
rect 665 1550 695 1555
rect 775 1575 805 1580
rect 775 1555 780 1575
rect 780 1555 800 1575
rect 800 1555 805 1575
rect 775 1550 805 1555
rect 885 1575 915 1580
rect 885 1555 890 1575
rect 890 1555 910 1575
rect 910 1555 915 1575
rect 885 1550 915 1555
rect 995 1575 1025 1580
rect 995 1555 1000 1575
rect 1000 1555 1020 1575
rect 1020 1555 1025 1575
rect 995 1550 1025 1555
rect 1105 1575 1135 1580
rect 1105 1555 1110 1575
rect 1110 1555 1130 1575
rect 1130 1555 1135 1575
rect 1105 1550 1135 1555
rect 1215 1575 1245 1580
rect 1215 1555 1220 1575
rect 1220 1555 1240 1575
rect 1240 1555 1245 1575
rect 1215 1550 1245 1555
rect 1325 1575 1355 1580
rect 1325 1555 1330 1575
rect 1330 1555 1350 1575
rect 1350 1555 1355 1575
rect 1325 1550 1355 1555
rect 1435 1575 1465 1580
rect 1435 1555 1440 1575
rect 1440 1555 1460 1575
rect 1460 1555 1465 1575
rect 1435 1550 1465 1555
rect 1810 1550 1840 1580
rect -150 1455 -120 1485
rect -240 1225 -210 1255
rect -285 685 -255 715
rect -1060 665 -1030 670
rect -1060 645 -1055 665
rect -1055 645 -1035 665
rect -1035 645 -1030 665
rect -1060 640 -1030 645
rect -995 665 -965 670
rect -995 645 -990 665
rect -990 645 -970 665
rect -970 645 -965 665
rect -995 640 -965 645
rect -885 665 -855 670
rect -885 645 -880 665
rect -880 645 -860 665
rect -860 645 -855 665
rect -885 640 -855 645
rect -775 665 -745 670
rect -775 645 -770 665
rect -770 645 -750 665
rect -750 645 -745 665
rect -775 640 -745 645
rect -665 665 -635 670
rect -665 645 -660 665
rect -660 645 -640 665
rect -640 645 -635 665
rect -665 640 -635 645
rect -555 665 -525 670
rect -555 645 -550 665
rect -550 645 -530 665
rect -530 645 -525 665
rect -555 640 -525 645
rect -445 665 -415 670
rect -445 645 -440 665
rect -440 645 -420 665
rect -420 645 -415 665
rect -445 640 -415 645
rect -380 665 -350 670
rect -380 645 -375 665
rect -375 645 -355 665
rect -355 645 -350 665
rect -380 640 -350 645
rect -1185 365 -1155 395
rect -940 390 -910 395
rect -940 370 -935 390
rect -935 370 -915 390
rect -915 370 -910 390
rect -940 365 -910 370
rect -830 390 -800 395
rect -830 370 -825 390
rect -825 370 -805 390
rect -805 370 -800 390
rect -830 365 -800 370
rect -720 390 -690 395
rect -720 370 -715 390
rect -715 370 -695 390
rect -695 370 -690 390
rect -720 365 -690 370
rect -610 390 -580 395
rect -610 370 -605 390
rect -605 370 -585 390
rect -585 370 -580 390
rect -610 365 -580 370
rect -500 390 -470 395
rect -500 370 -495 390
rect -495 370 -475 390
rect -475 370 -470 390
rect -500 365 -470 370
rect -1535 320 -1505 350
rect -1406 -93 -1379 -85
rect -1406 -113 -1405 -93
rect -1405 -113 -1380 -93
rect -1380 -113 -1379 -93
rect -1406 -120 -1379 -113
rect -1346 -93 -1319 -85
rect -1346 -113 -1345 -93
rect -1345 -113 -1320 -93
rect -1320 -113 -1319 -93
rect -1346 -120 -1319 -113
rect -1286 -93 -1259 -85
rect -1286 -113 -1285 -93
rect -1285 -113 -1260 -93
rect -1260 -113 -1259 -93
rect -1286 -120 -1259 -113
rect -1226 -93 -1199 -85
rect -1226 -113 -1225 -93
rect -1225 -113 -1200 -93
rect -1200 -113 -1199 -93
rect -1226 -120 -1199 -113
rect -665 310 -635 340
rect -285 310 -255 340
rect -1140 255 -1110 285
rect -940 280 -910 285
rect -940 260 -935 280
rect -935 260 -915 280
rect -915 260 -910 280
rect -940 255 -910 260
rect -830 280 -800 285
rect -830 260 -825 280
rect -825 260 -805 280
rect -805 260 -800 280
rect -830 255 -800 260
rect -720 280 -690 285
rect -720 260 -715 280
rect -715 260 -695 280
rect -695 260 -690 280
rect -720 255 -690 260
rect -610 280 -580 285
rect -610 260 -605 280
rect -605 260 -585 280
rect -585 260 -580 280
rect -610 255 -580 260
rect -500 280 -470 285
rect -500 260 -495 280
rect -495 260 -475 280
rect -475 260 -470 280
rect -500 255 -470 260
rect -1140 -120 -1110 -90
rect -995 -95 -965 -90
rect -995 -115 -990 -95
rect -990 -115 -970 -95
rect -970 -115 -965 -95
rect -995 -120 -965 -115
rect -885 -95 -855 -90
rect -885 -115 -880 -95
rect -880 -115 -860 -95
rect -860 -115 -855 -95
rect -885 -120 -855 -115
rect -775 -95 -745 -90
rect -775 -115 -770 -95
rect -770 -115 -750 -95
rect -750 -115 -745 -95
rect -775 -120 -745 -115
rect -665 -95 -635 -90
rect -665 -115 -660 -95
rect -660 -115 -640 -95
rect -640 -115 -635 -95
rect -665 -120 -635 -115
rect -555 -95 -525 -90
rect -555 -115 -550 -95
rect -550 -115 -530 -95
rect -530 -115 -525 -95
rect -555 -120 -525 -115
rect -445 -95 -415 -90
rect -445 -115 -440 -95
rect -440 -115 -420 -95
rect -420 -115 -415 -95
rect -445 -120 -415 -115
rect -1290 -175 -1255 -145
rect -1185 -175 -1155 -145
rect -1060 -175 -1030 -145
rect -380 -175 -350 -145
rect 280 1450 310 1455
rect 280 1430 285 1450
rect 285 1430 305 1450
rect 305 1430 310 1450
rect 280 1425 310 1430
rect 500 1450 530 1455
rect 500 1430 505 1450
rect 505 1430 525 1450
rect 525 1430 530 1450
rect 500 1425 530 1430
rect 720 1450 750 1455
rect 720 1430 725 1450
rect 725 1430 745 1450
rect 745 1430 750 1450
rect 720 1425 750 1430
rect 940 1450 970 1455
rect 940 1430 945 1450
rect 945 1430 965 1450
rect 965 1430 970 1450
rect 940 1425 970 1430
rect 1160 1450 1190 1455
rect 1160 1430 1165 1450
rect 1165 1430 1185 1450
rect 1185 1430 1190 1450
rect 1160 1425 1190 1430
rect 1380 1450 1410 1455
rect 1380 1430 1385 1450
rect 1385 1430 1405 1450
rect 1405 1430 1410 1450
rect 1380 1425 1410 1430
rect 1810 1455 1840 1485
rect 390 1370 420 1400
rect 610 1370 640 1400
rect 830 1370 860 1400
rect 120 1280 150 1310
rect 220 1280 250 1310
rect 330 1280 360 1310
rect 440 1280 470 1310
rect 550 1280 580 1310
rect 71 1250 101 1255
rect 71 1230 76 1250
rect 76 1230 96 1250
rect 96 1230 101 1250
rect 71 1225 101 1230
rect 275 1250 305 1255
rect 275 1230 280 1250
rect 280 1230 300 1250
rect 300 1230 305 1250
rect 275 1225 305 1230
rect 495 1250 525 1255
rect 495 1230 500 1250
rect 500 1230 520 1250
rect 520 1230 525 1250
rect 495 1225 525 1230
rect -150 1165 -120 1195
rect -40 1190 -10 1195
rect -40 1170 -35 1190
rect -35 1170 -15 1190
rect -15 1170 -10 1190
rect -40 1165 -10 1170
rect -195 740 -165 770
rect 204 1131 234 1136
rect 204 1111 209 1131
rect 209 1111 229 1131
rect 229 1111 234 1131
rect 204 1106 234 1111
rect 424 1131 454 1136
rect 424 1111 429 1131
rect 429 1111 449 1131
rect 449 1111 454 1131
rect 424 1106 454 1111
rect 566 1131 596 1136
rect 566 1111 571 1131
rect 571 1111 591 1131
rect 591 1111 596 1131
rect 566 1106 596 1111
rect 1050 1370 1080 1400
rect 1270 1370 1300 1400
rect 1120 1280 1150 1310
rect 1220 1280 1250 1310
rect 1330 1280 1360 1310
rect 1440 1280 1470 1310
rect 1550 1280 1580 1310
rect 1071 1250 1101 1255
rect 1071 1230 1076 1250
rect 1076 1230 1096 1250
rect 1096 1230 1101 1250
rect 1071 1225 1101 1230
rect 1275 1250 1305 1255
rect 1275 1230 1280 1250
rect 1280 1230 1300 1250
rect 1300 1230 1305 1250
rect 1275 1225 1305 1230
rect 1495 1250 1525 1255
rect 1495 1230 1500 1250
rect 1500 1230 1520 1250
rect 1520 1230 1525 1250
rect 1495 1225 1525 1230
rect 1900 1225 1930 1255
rect 1700 1190 1730 1195
rect 1700 1170 1705 1190
rect 1705 1170 1725 1190
rect 1725 1170 1730 1190
rect 1700 1165 1730 1170
rect 1810 1165 1840 1195
rect 1204 1131 1234 1136
rect 1204 1111 1209 1131
rect 1209 1111 1229 1131
rect 1229 1111 1234 1131
rect 1204 1106 1234 1111
rect 1424 1131 1454 1136
rect 1424 1111 1429 1131
rect 1429 1111 1449 1131
rect 1449 1111 1454 1131
rect 1424 1106 1454 1111
rect 1566 1131 1596 1136
rect 1566 1111 1571 1131
rect 1571 1111 1591 1131
rect 1591 1111 1596 1131
rect 1566 1106 1596 1111
rect 55 1045 85 1075
rect 165 1045 195 1075
rect 275 1045 305 1075
rect 385 1045 415 1075
rect 495 1045 525 1075
rect 605 1045 635 1075
rect 885 1045 915 1075
rect 1055 1045 1085 1075
rect 555 990 585 1020
rect 1275 1045 1305 1075
rect 1495 1045 1525 1075
rect 1165 1000 1195 1030
rect 1385 1000 1415 1030
rect 1605 1000 1635 1030
rect 665 955 695 985
rect 885 955 915 985
rect 1045 955 1075 985
rect 1105 955 1135 985
rect 555 925 585 930
rect 555 905 560 925
rect 560 905 580 925
rect 580 905 585 925
rect 555 900 585 905
rect 775 925 805 930
rect 775 905 780 925
rect 780 905 800 925
rect 800 905 805 925
rect 775 900 805 905
rect 995 925 1025 930
rect 995 905 1000 925
rect 1000 905 1020 925
rect 1020 905 1025 925
rect 995 900 1025 905
rect 1765 900 1795 930
rect 500 805 530 810
rect 500 785 505 805
rect 505 785 525 805
rect 525 785 530 805
rect 500 780 530 785
rect 610 805 640 810
rect 610 785 615 805
rect 615 785 635 805
rect 635 785 640 805
rect 610 780 640 785
rect 720 805 750 810
rect 720 785 725 805
rect 725 785 745 805
rect 745 785 750 805
rect 720 780 750 785
rect 830 805 860 810
rect 830 785 835 805
rect 835 785 855 805
rect 855 785 860 805
rect 830 780 860 785
rect 940 805 970 810
rect 940 785 945 805
rect 945 785 965 805
rect 965 785 970 805
rect 940 780 970 785
rect 1050 805 1080 810
rect 1050 785 1055 805
rect 1055 785 1075 805
rect 1075 785 1080 805
rect 1050 780 1080 785
rect 1160 805 1190 810
rect 1160 785 1165 805
rect 1165 785 1185 805
rect 1185 785 1190 805
rect 1160 780 1190 785
rect 35 685 65 715
rect 145 685 175 715
rect 255 685 285 715
rect 365 685 395 715
rect 475 685 505 715
rect 585 685 615 715
rect 1075 685 1105 715
rect 1185 685 1215 715
rect 1295 685 1325 715
rect 1405 685 1435 715
rect 1515 685 1545 715
rect 1625 685 1655 715
rect -150 640 -120 670
rect -95 630 -65 660
rect 310 655 340 660
rect 310 635 315 655
rect 315 635 335 655
rect 335 635 340 655
rect 310 630 340 635
rect 1350 655 1380 660
rect 1350 635 1355 655
rect 1355 635 1375 655
rect 1375 635 1380 655
rect 1350 630 1380 635
rect -150 -120 -120 -90
rect -195 -175 -165 -145
rect -1410 -220 -1375 -190
rect -240 -220 -210 -190
rect -1210 -270 -1175 -240
rect -620 -270 -590 -240
rect -1535 -330 -1505 -300
rect -1150 -330 -1115 -300
rect -920 -305 -890 -300
rect -920 -325 -915 -305
rect -915 -325 -895 -305
rect -895 -325 -890 -305
rect -920 -330 -890 -325
rect -720 -305 -690 -300
rect -720 -325 -715 -305
rect -715 -325 -695 -305
rect -695 -325 -690 -305
rect -720 -330 -690 -325
rect -520 -305 -490 -300
rect -520 -325 -515 -305
rect -515 -325 -495 -305
rect -495 -325 -490 -305
rect -520 -330 -490 -325
rect -1206 -387 -1179 -380
rect -1206 -407 -1205 -387
rect -1205 -407 -1180 -387
rect -1180 -407 -1179 -387
rect -1206 -415 -1179 -407
rect -1146 -387 -1119 -380
rect -1146 -407 -1145 -387
rect -1145 -407 -1120 -387
rect -1120 -407 -1119 -387
rect -1146 -415 -1119 -407
rect -20 430 10 435
rect -20 410 -15 430
rect -15 410 5 430
rect 5 410 10 430
rect -20 405 10 410
rect 640 430 670 435
rect 640 410 645 430
rect 645 410 665 430
rect 665 410 670 430
rect 640 405 670 410
rect 1020 430 1050 435
rect 1020 410 1025 430
rect 1025 410 1045 430
rect 1045 410 1050 430
rect 1020 405 1050 410
rect 1680 430 1710 435
rect 1680 410 1685 430
rect 1685 410 1705 430
rect 1705 410 1710 430
rect 1680 405 1710 410
rect 90 345 120 375
rect 200 345 230 375
rect 310 345 340 375
rect 420 345 450 375
rect 530 345 560 375
rect 1130 345 1160 375
rect 1240 345 1270 375
rect 1350 345 1380 375
rect 1460 345 1490 375
rect 1570 345 1600 375
rect 35 225 65 230
rect 35 205 40 225
rect 40 205 60 225
rect 60 205 65 225
rect 35 200 65 205
rect 145 225 175 230
rect 145 205 150 225
rect 150 205 170 225
rect 170 205 175 225
rect 145 200 175 205
rect 255 225 285 230
rect 255 205 260 225
rect 260 205 280 225
rect 280 205 285 225
rect 255 200 285 205
rect 310 210 340 240
rect 365 225 395 230
rect 365 205 370 225
rect 370 205 390 225
rect 390 205 395 225
rect 365 200 395 205
rect 475 225 505 230
rect 475 205 480 225
rect 480 205 500 225
rect 500 205 505 225
rect 475 200 505 205
rect 585 225 615 230
rect 585 205 590 225
rect 590 205 610 225
rect 610 205 615 225
rect 585 200 615 205
rect 1075 225 1105 230
rect 1075 205 1080 225
rect 1080 205 1100 225
rect 1100 205 1105 225
rect 1075 200 1105 205
rect 1185 225 1215 230
rect 1185 205 1190 225
rect 1190 205 1210 225
rect 1210 205 1215 225
rect 1185 200 1215 205
rect 1295 225 1325 230
rect 1295 205 1300 225
rect 1300 205 1320 225
rect 1320 205 1325 225
rect 1295 200 1325 205
rect 1350 210 1380 240
rect 1405 225 1435 230
rect 1405 205 1410 225
rect 1410 205 1430 225
rect 1430 205 1435 225
rect 1405 200 1435 205
rect 1515 225 1545 230
rect 1515 205 1520 225
rect 1520 205 1540 225
rect 1540 205 1545 225
rect 1515 200 1545 205
rect 1625 225 1655 230
rect 1625 205 1630 225
rect 1630 205 1650 225
rect 1650 205 1655 225
rect 1625 200 1655 205
rect 310 175 340 180
rect 310 155 315 175
rect 315 155 335 175
rect 335 155 340 175
rect 310 150 340 155
rect 795 175 825 180
rect 795 155 800 175
rect 800 155 820 175
rect 820 155 825 175
rect 795 150 825 155
rect 848 175 878 180
rect 848 155 853 175
rect 853 155 873 175
rect 873 155 878 175
rect 848 150 878 155
rect 1350 175 1380 180
rect 1350 155 1355 175
rect 1355 155 1375 175
rect 1375 155 1380 175
rect 1350 150 1380 155
rect 90 -45 120 -40
rect 90 -65 95 -45
rect 95 -65 115 -45
rect 115 -65 120 -45
rect 90 -70 120 -65
rect 200 -45 230 -40
rect 200 -65 205 -45
rect 205 -65 225 -45
rect 225 -65 230 -45
rect 200 -70 230 -65
rect 310 -45 340 -40
rect 310 -65 315 -45
rect 315 -65 335 -45
rect 335 -65 340 -45
rect 310 -70 340 -65
rect 420 -45 450 -40
rect 420 -65 425 -45
rect 425 -65 445 -45
rect 445 -65 450 -45
rect 420 -70 450 -65
rect 530 -45 560 -40
rect 530 -65 535 -45
rect 535 -65 555 -45
rect 555 -65 560 -45
rect 530 -70 560 -65
rect 1130 -45 1160 -40
rect 1130 -65 1135 -45
rect 1135 -65 1155 -45
rect 1155 -65 1160 -45
rect 1130 -70 1160 -65
rect 1240 -45 1270 -40
rect 1240 -65 1245 -45
rect 1245 -65 1265 -45
rect 1265 -65 1270 -45
rect 1240 -70 1270 -65
rect 1350 -45 1380 -40
rect 1350 -65 1355 -45
rect 1355 -65 1375 -45
rect 1375 -65 1380 -45
rect 1350 -70 1380 -65
rect 1460 -45 1490 -40
rect 1460 -65 1465 -45
rect 1465 -65 1485 -45
rect 1485 -65 1490 -45
rect 1460 -70 1490 -65
rect 1570 -45 1600 -40
rect 1570 -65 1575 -45
rect 1575 -65 1595 -45
rect 1595 -65 1600 -45
rect 1570 -70 1600 -65
rect 765 -125 795 -95
rect -20 -170 10 -140
rect 680 -170 710 -140
rect 80 -225 110 -195
rect 715 -225 745 -195
rect 275 -325 305 -295
rect 895 -125 925 -95
rect 980 -170 1010 -140
rect 830 -325 860 -295
rect 1680 -170 1710 -140
rect 1855 740 1885 770
rect 1810 640 1840 670
rect 1855 405 1885 435
rect 1810 -120 1840 -90
rect 1855 -175 1885 -145
rect 1335 -325 1365 -295
rect 1765 -325 1795 -295
rect 385 -355 415 -350
rect 385 -375 390 -355
rect 390 -375 410 -355
rect 410 -375 415 -355
rect 385 -380 415 -375
rect 495 -355 525 -350
rect 495 -375 500 -355
rect 500 -375 520 -355
rect 520 -375 525 -355
rect 495 -380 525 -375
rect 605 -355 635 -350
rect 605 -375 610 -355
rect 610 -375 630 -355
rect 630 -375 635 -355
rect 605 -380 635 -375
rect 715 -355 745 -350
rect 715 -375 720 -355
rect 720 -375 740 -355
rect 740 -375 745 -355
rect 715 -380 745 -375
rect 825 -355 855 -350
rect 825 -375 830 -355
rect 830 -375 850 -355
rect 850 -375 855 -355
rect 825 -380 855 -375
rect 935 -355 965 -350
rect 935 -375 940 -355
rect 940 -375 960 -355
rect 960 -375 965 -355
rect 935 -380 965 -375
rect 1045 -355 1075 -350
rect 1045 -375 1050 -355
rect 1050 -375 1070 -355
rect 1070 -375 1075 -355
rect 1045 -380 1075 -375
rect 1155 -355 1185 -350
rect 1155 -375 1160 -355
rect 1160 -375 1180 -355
rect 1180 -375 1185 -355
rect 1155 -380 1185 -375
rect 1265 -355 1295 -350
rect 1265 -375 1270 -355
rect 1270 -375 1290 -355
rect 1290 -375 1295 -355
rect 1265 -380 1295 -375
rect 1390 -355 1420 -350
rect 1390 -375 1395 -355
rect 1395 -375 1415 -355
rect 1415 -375 1420 -355
rect 1390 -380 1420 -375
rect 2380 1595 2410 1625
rect 2050 1480 2080 1485
rect 2050 1460 2055 1480
rect 2055 1460 2075 1480
rect 2075 1460 2080 1480
rect 2050 1455 2080 1460
rect 2160 1480 2190 1485
rect 2160 1460 2165 1480
rect 2165 1460 2185 1480
rect 2185 1460 2190 1480
rect 2160 1455 2190 1460
rect 2270 1480 2300 1485
rect 2270 1460 2275 1480
rect 2275 1460 2295 1480
rect 2295 1460 2300 1480
rect 2270 1455 2300 1460
rect 2380 1480 2410 1485
rect 2380 1460 2385 1480
rect 2385 1460 2405 1480
rect 2405 1460 2410 1480
rect 2380 1455 2410 1460
rect 2490 1480 2520 1485
rect 2490 1460 2495 1480
rect 2495 1460 2515 1480
rect 2515 1460 2520 1480
rect 2490 1455 2520 1460
rect 2600 1480 2630 1485
rect 2600 1460 2605 1480
rect 2605 1460 2625 1480
rect 2625 1460 2630 1480
rect 2600 1455 2630 1460
rect 2710 1480 2740 1485
rect 2710 1460 2715 1480
rect 2715 1460 2735 1480
rect 2735 1460 2740 1480
rect 2710 1455 2740 1460
rect 3105 1460 3135 1490
rect 2105 805 2135 810
rect 2105 785 2110 805
rect 2110 785 2130 805
rect 2130 785 2135 805
rect 2105 780 2135 785
rect 2215 805 2245 810
rect 2215 785 2220 805
rect 2220 785 2240 805
rect 2240 785 2245 805
rect 2215 780 2245 785
rect 2325 805 2355 810
rect 2325 785 2330 805
rect 2330 785 2350 805
rect 2350 785 2355 805
rect 2325 780 2355 785
rect 2435 805 2465 810
rect 2435 785 2440 805
rect 2440 785 2460 805
rect 2460 785 2465 805
rect 2435 780 2465 785
rect 2545 805 2575 810
rect 2545 785 2550 805
rect 2550 785 2570 805
rect 2570 785 2575 805
rect 2545 780 2575 785
rect 2655 805 2685 810
rect 2655 785 2660 805
rect 2660 785 2680 805
rect 2680 785 2685 805
rect 2655 780 2685 785
rect 2105 730 2135 760
rect 1945 685 1975 715
rect 2545 730 2575 760
rect 3195 730 3225 760
rect 2380 685 2410 715
rect 3105 685 3135 715
rect 2040 665 2070 670
rect 2040 645 2045 665
rect 2045 645 2065 665
rect 2065 645 2070 665
rect 2040 640 2070 645
rect 2105 665 2135 670
rect 2105 645 2110 665
rect 2110 645 2130 665
rect 2130 645 2135 665
rect 2105 640 2135 645
rect 2215 665 2245 670
rect 2215 645 2220 665
rect 2220 645 2240 665
rect 2240 645 2245 665
rect 2215 640 2245 645
rect 2325 665 2355 670
rect 2325 645 2330 665
rect 2330 645 2350 665
rect 2350 645 2355 665
rect 2325 640 2355 645
rect 2435 665 2465 670
rect 2435 645 2440 665
rect 2440 645 2460 665
rect 2460 645 2465 665
rect 2435 640 2465 645
rect 2545 665 2575 670
rect 2545 645 2550 665
rect 2550 645 2570 665
rect 2570 645 2575 665
rect 2545 640 2575 645
rect 2655 665 2685 670
rect 2655 645 2660 665
rect 2660 645 2680 665
rect 2680 645 2685 665
rect 2655 640 2685 645
rect 2720 665 2750 670
rect 2720 645 2725 665
rect 2725 645 2745 665
rect 2745 645 2750 665
rect 2720 640 2750 645
rect 2160 390 2190 395
rect 2160 370 2165 390
rect 2165 370 2185 390
rect 2185 370 2190 390
rect 2160 365 2190 370
rect 2270 390 2300 395
rect 2270 370 2275 390
rect 2275 370 2295 390
rect 2295 370 2300 390
rect 2270 365 2300 370
rect 2380 390 2410 395
rect 2380 370 2385 390
rect 2385 370 2405 390
rect 2405 370 2410 390
rect 2380 365 2410 370
rect 2490 390 2520 395
rect 2490 370 2495 390
rect 2495 370 2515 390
rect 2515 370 2520 390
rect 2490 365 2520 370
rect 2600 390 2630 395
rect 2600 370 2605 390
rect 2605 370 2625 390
rect 2625 370 2630 390
rect 2600 365 2630 370
rect 2845 365 2875 395
rect 1945 310 1975 340
rect 2325 310 2355 340
rect 2160 280 2190 285
rect 2160 260 2165 280
rect 2165 260 2185 280
rect 2185 260 2190 280
rect 2160 255 2190 260
rect 2270 280 2300 285
rect 2270 260 2275 280
rect 2275 260 2295 280
rect 2295 260 2300 280
rect 2270 255 2300 260
rect 2380 280 2410 285
rect 2380 260 2385 280
rect 2385 260 2405 280
rect 2405 260 2410 280
rect 2380 255 2410 260
rect 2490 280 2520 285
rect 2490 260 2495 280
rect 2495 260 2515 280
rect 2515 260 2520 280
rect 2490 255 2520 260
rect 2600 280 2630 285
rect 2600 260 2605 280
rect 2605 260 2625 280
rect 2625 260 2630 280
rect 2600 255 2630 260
rect 2800 255 2830 285
rect 2105 -95 2135 -90
rect 2105 -115 2110 -95
rect 2110 -115 2130 -95
rect 2130 -115 2135 -95
rect 2105 -120 2135 -115
rect 2215 -95 2245 -90
rect 2215 -115 2220 -95
rect 2220 -115 2240 -95
rect 2240 -115 2245 -95
rect 2215 -120 2245 -115
rect 2325 -95 2355 -90
rect 2325 -115 2330 -95
rect 2330 -115 2350 -95
rect 2350 -115 2355 -95
rect 2325 -120 2355 -115
rect 2435 -95 2465 -90
rect 2435 -115 2440 -95
rect 2440 -115 2460 -95
rect 2460 -115 2465 -95
rect 2435 -120 2465 -115
rect 2545 -95 2575 -90
rect 2545 -115 2550 -95
rect 2550 -115 2570 -95
rect 2570 -115 2575 -95
rect 2545 -120 2575 -115
rect 2655 -95 2685 -90
rect 2655 -115 2660 -95
rect 2660 -115 2680 -95
rect 2680 -115 2685 -95
rect 2655 -120 2685 -115
rect 2800 -120 2830 -90
rect 3195 320 3225 350
rect 2889 -93 2916 -85
rect 2889 -113 2890 -93
rect 2890 -113 2915 -93
rect 2915 -113 2916 -93
rect 2889 -120 2916 -113
rect 2949 -93 2976 -85
rect 2949 -113 2950 -93
rect 2950 -113 2975 -93
rect 2975 -113 2976 -93
rect 2949 -120 2976 -113
rect 3009 -93 3036 -85
rect 3009 -113 3010 -93
rect 3010 -113 3035 -93
rect 3035 -113 3036 -93
rect 3009 -120 3036 -113
rect 3069 -93 3096 -85
rect 3069 -113 3070 -93
rect 3070 -113 3095 -93
rect 3095 -113 3096 -93
rect 3069 -120 3096 -113
rect 2040 -175 2070 -145
rect 2720 -175 2750 -145
rect 2845 -175 2875 -145
rect 2945 -175 2980 -145
rect 1900 -220 1930 -190
rect 3065 -220 3100 -190
rect 2280 -270 2310 -240
rect 2865 -270 2900 -240
rect 2180 -305 2210 -300
rect 2180 -325 2185 -305
rect 2185 -325 2205 -305
rect 2205 -325 2210 -305
rect 2180 -330 2210 -325
rect 2380 -305 2410 -300
rect 2380 -325 2385 -305
rect 2385 -325 2405 -305
rect 2405 -325 2410 -305
rect 2380 -330 2410 -325
rect 2580 -305 2610 -300
rect 2580 -325 2585 -305
rect 2585 -325 2605 -305
rect 2605 -325 2610 -305
rect 2580 -330 2610 -325
rect 2805 -330 2840 -300
rect 3195 -330 3225 -300
rect 2809 -387 2836 -380
rect 2809 -407 2810 -387
rect 2810 -407 2835 -387
rect 2835 -407 2836 -387
rect 2809 -415 2836 -407
rect 2869 -387 2896 -380
rect 2869 -407 2870 -387
rect 2870 -407 2895 -387
rect 2895 -407 2896 -387
rect 2869 -415 2896 -407
rect 155 -680 185 -675
rect 155 -700 160 -680
rect 160 -700 180 -680
rect 180 -700 185 -680
rect 155 -705 185 -700
rect 220 -680 250 -675
rect 220 -700 225 -680
rect 225 -700 245 -680
rect 245 -700 250 -680
rect 220 -705 250 -700
rect 330 -680 360 -675
rect 330 -700 335 -680
rect 335 -700 355 -680
rect 355 -700 360 -680
rect 330 -705 360 -700
rect 440 -680 470 -675
rect 440 -700 445 -680
rect 445 -700 465 -680
rect 465 -700 470 -680
rect 440 -705 470 -700
rect 550 -680 580 -675
rect 550 -700 555 -680
rect 555 -700 575 -680
rect 575 -700 580 -680
rect 550 -705 580 -700
rect 660 -680 690 -675
rect 660 -700 665 -680
rect 665 -700 685 -680
rect 685 -700 690 -680
rect 660 -705 690 -700
rect 770 -680 800 -675
rect 770 -700 775 -680
rect 775 -700 795 -680
rect 795 -700 800 -680
rect 770 -705 800 -700
rect 880 -680 910 -675
rect 880 -700 885 -680
rect 885 -700 905 -680
rect 905 -700 910 -680
rect 880 -705 910 -700
rect 990 -680 1020 -675
rect 990 -700 995 -680
rect 995 -700 1015 -680
rect 1015 -700 1020 -680
rect 990 -705 1020 -700
rect 1100 -680 1130 -675
rect 1100 -700 1105 -680
rect 1105 -700 1125 -680
rect 1125 -700 1130 -680
rect 1100 -705 1130 -700
rect 1210 -680 1240 -675
rect 1210 -700 1215 -680
rect 1215 -700 1235 -680
rect 1235 -700 1240 -680
rect 1210 -705 1240 -700
rect 1320 -680 1350 -675
rect 1320 -700 1325 -680
rect 1325 -700 1345 -680
rect 1345 -700 1350 -680
rect 1320 -705 1350 -700
rect 1430 -680 1460 -675
rect 1430 -700 1435 -680
rect 1435 -700 1455 -680
rect 1455 -700 1460 -680
rect 1430 -705 1460 -700
rect 1855 -705 1885 -675
rect 80 -755 110 -725
rect 1015 -740 1045 -735
rect 1015 -760 1020 -740
rect 1020 -760 1040 -740
rect 1040 -760 1045 -740
rect 1015 -765 1045 -760
rect -105 -800 -75 -770
rect 715 -775 745 -770
rect 715 -795 720 -775
rect 720 -795 740 -775
rect 740 -795 745 -775
rect 715 -800 745 -795
rect 830 -775 860 -770
rect 830 -795 835 -775
rect 835 -795 855 -775
rect 855 -795 860 -775
rect 830 -800 860 -795
rect 955 -775 985 -770
rect 955 -795 960 -775
rect 960 -795 980 -775
rect 980 -795 985 -775
rect 955 -800 985 -795
rect -1020 -1080 -990 -1075
rect -1020 -1100 -1015 -1080
rect -1015 -1100 -995 -1080
rect -995 -1100 -990 -1080
rect -1020 -1105 -990 -1100
rect -820 -1080 -790 -1075
rect -820 -1100 -815 -1080
rect -815 -1100 -795 -1080
rect -795 -1100 -790 -1080
rect -820 -1105 -790 -1100
rect -620 -1080 -590 -1075
rect -620 -1100 -615 -1080
rect -615 -1100 -595 -1080
rect -595 -1100 -590 -1080
rect -620 -1105 -590 -1100
rect -420 -1080 -390 -1075
rect -420 -1100 -415 -1080
rect -415 -1100 -395 -1080
rect -395 -1100 -390 -1080
rect -420 -1105 -390 -1100
rect -195 -1105 -165 -1075
rect 830 -1105 860 -1075
rect 1855 -1105 1885 -1075
rect 2080 -1080 2110 -1075
rect 2080 -1100 2085 -1080
rect 2085 -1100 2105 -1080
rect 2105 -1100 2110 -1080
rect 2080 -1105 2110 -1100
rect 2280 -1080 2310 -1075
rect 2280 -1100 2285 -1080
rect 2285 -1100 2305 -1080
rect 2305 -1100 2310 -1080
rect 2280 -1105 2310 -1100
rect 2480 -1080 2510 -1075
rect 2480 -1100 2485 -1080
rect 2485 -1100 2505 -1080
rect 2505 -1100 2510 -1080
rect 2480 -1105 2510 -1100
rect 2680 -1080 2710 -1075
rect 2680 -1100 2685 -1080
rect 2685 -1100 2705 -1080
rect 2705 -1100 2710 -1080
rect 2680 -1105 2710 -1100
rect 830 -2455 860 -2425
<< metal2 >>
rect 825 4275 865 4280
rect 825 4245 830 4275
rect 860 4245 865 4275
rect 825 4240 865 4245
rect 150 2780 190 2785
rect 150 2750 155 2780
rect 185 2775 190 2780
rect 620 2780 660 2785
rect 620 2775 625 2780
rect 185 2755 625 2775
rect 185 2750 190 2755
rect 150 2745 190 2750
rect 620 2750 625 2755
rect 655 2750 660 2780
rect 620 2745 660 2750
rect 1030 2780 1070 2785
rect 1030 2750 1035 2780
rect 1065 2775 1070 2780
rect 1498 2780 1538 2785
rect 1498 2775 1503 2780
rect 1065 2755 1503 2775
rect 1065 2750 1070 2755
rect 1030 2745 1070 2750
rect 1498 2750 1503 2755
rect 1533 2750 1538 2780
rect 1498 2745 1538 2750
rect 30 2725 70 2730
rect 30 2695 35 2725
rect 65 2720 70 2725
rect 150 2725 190 2730
rect 150 2720 155 2725
rect 65 2700 155 2720
rect 65 2695 70 2700
rect 30 2690 70 2695
rect 150 2695 155 2700
rect 185 2720 190 2725
rect 210 2725 250 2730
rect 210 2720 215 2725
rect 185 2700 215 2720
rect 185 2695 190 2700
rect 150 2690 190 2695
rect 210 2695 215 2700
rect 245 2695 250 2725
rect 210 2690 250 2695
rect 825 2725 865 2730
rect 825 2695 830 2725
rect 860 2720 865 2725
rect 970 2725 1010 2730
rect 970 2720 975 2725
rect 860 2700 975 2720
rect 860 2695 865 2700
rect 825 2690 865 2695
rect 970 2695 975 2700
rect 1005 2720 1010 2725
rect 1090 2725 1130 2730
rect 1090 2720 1095 2725
rect 1005 2700 1095 2720
rect 1005 2695 1010 2700
rect 970 2690 1010 2695
rect 1090 2695 1095 2700
rect 1125 2720 1130 2725
rect 1150 2725 1190 2730
rect 1150 2720 1155 2725
rect 1125 2700 1155 2720
rect 1125 2695 1130 2700
rect 1090 2690 1130 2695
rect 1150 2695 1155 2700
rect 1185 2695 1190 2725
rect 1150 2690 1190 2695
rect 1438 2725 1478 2730
rect 1438 2695 1443 2725
rect 1473 2720 1478 2725
rect 1498 2725 1538 2730
rect 1498 2720 1503 2725
rect 1473 2700 1503 2720
rect 1473 2695 1478 2700
rect 1438 2690 1478 2695
rect 1498 2695 1503 2700
rect 1533 2720 1538 2725
rect 1618 2725 1658 2730
rect 1618 2720 1623 2725
rect 1533 2700 1623 2720
rect 1533 2695 1538 2700
rect 1498 2690 1538 2695
rect 1618 2695 1623 2700
rect 1653 2695 1658 2725
rect 1618 2690 1658 2695
rect 500 2555 540 2560
rect 500 2525 505 2555
rect 535 2550 540 2555
rect 560 2555 600 2560
rect 560 2550 565 2555
rect 535 2530 565 2550
rect 535 2525 540 2530
rect 500 2520 540 2525
rect 560 2525 565 2530
rect 595 2550 600 2555
rect 680 2555 720 2560
rect 680 2550 685 2555
rect 595 2530 685 2550
rect 595 2525 600 2530
rect 560 2520 600 2525
rect 680 2525 685 2530
rect 715 2550 720 2555
rect 825 2555 865 2560
rect 825 2550 830 2555
rect 715 2530 830 2550
rect 715 2525 720 2530
rect 680 2520 720 2525
rect 825 2525 830 2530
rect 860 2525 865 2555
rect 825 2520 865 2525
rect 75 2305 115 2310
rect 75 2275 80 2305
rect 110 2300 115 2305
rect 139 2305 169 2310
rect 110 2280 139 2300
rect 110 2275 115 2280
rect 75 2270 115 2275
rect 609 2305 639 2310
rect 169 2280 609 2300
rect 139 2270 169 2275
rect 770 2305 810 2310
rect 770 2300 775 2305
rect 639 2280 775 2300
rect 609 2270 639 2275
rect 770 2275 775 2280
rect 805 2300 810 2305
rect 1519 2305 1549 2310
rect 805 2280 1519 2300
rect 805 2275 810 2280
rect 770 2270 810 2275
rect 1519 2270 1549 2275
rect 880 2260 920 2265
rect 880 2230 885 2260
rect 915 2245 920 2260
rect 1045 2250 1085 2255
rect 1045 2245 1050 2250
rect 915 2230 1050 2245
rect 880 2225 1050 2230
rect 1045 2220 1050 2225
rect 1080 2245 1085 2250
rect 1573 2250 1613 2255
rect 1573 2245 1578 2250
rect 1080 2225 1578 2245
rect 1080 2220 1085 2225
rect 1045 2215 1085 2220
rect 1573 2220 1578 2225
rect 1608 2220 1613 2250
rect 1573 2215 1613 2220
rect -725 2205 -685 2210
rect -725 2175 -720 2205
rect -690 2200 -685 2205
rect -155 2205 -115 2210
rect -155 2200 -150 2205
rect -690 2180 -150 2200
rect -690 2175 -685 2180
rect -725 2170 -685 2175
rect -155 2175 -150 2180
rect -120 2200 -115 2205
rect 825 2205 865 2210
rect 825 2200 830 2205
rect -120 2180 830 2200
rect -120 2175 -115 2180
rect -155 2170 -115 2175
rect 825 2175 830 2180
rect 860 2200 865 2205
rect 1805 2205 1845 2210
rect 1805 2200 1810 2205
rect 860 2180 1810 2200
rect 860 2175 865 2180
rect 825 2170 865 2175
rect 1805 2175 1810 2180
rect 1840 2200 1845 2205
rect 2375 2205 2415 2210
rect 2375 2200 2380 2205
rect 1840 2180 2380 2200
rect 1840 2175 1845 2180
rect 1805 2170 1845 2175
rect 2375 2175 2380 2180
rect 2410 2175 2415 2205
rect 2375 2170 2415 2175
rect -1085 2150 -1045 2155
rect -1085 2120 -1080 2150
rect -1050 2145 -1045 2150
rect -965 2150 -925 2155
rect -965 2145 -960 2150
rect -1050 2125 -960 2145
rect -1050 2120 -1045 2125
rect -1085 2115 -1045 2120
rect -965 2120 -960 2125
rect -930 2145 -925 2150
rect -845 2150 -805 2155
rect -845 2145 -840 2150
rect -930 2125 -840 2145
rect -930 2120 -925 2125
rect -965 2115 -925 2120
rect -845 2120 -840 2125
rect -810 2145 -805 2150
rect -725 2150 -685 2155
rect -725 2145 -720 2150
rect -810 2125 -720 2145
rect -810 2120 -805 2125
rect -845 2115 -805 2120
rect -725 2120 -720 2125
rect -690 2145 -685 2150
rect -605 2150 -565 2155
rect -605 2145 -600 2150
rect -690 2125 -600 2145
rect -690 2120 -685 2125
rect -725 2115 -685 2120
rect -605 2120 -600 2125
rect -570 2145 -565 2150
rect -485 2150 -445 2155
rect -485 2145 -480 2150
rect -570 2125 -480 2145
rect -570 2120 -565 2125
rect -605 2115 -565 2120
rect -485 2120 -480 2125
rect -450 2145 -445 2150
rect -365 2150 -325 2155
rect -365 2145 -360 2150
rect -450 2125 -360 2145
rect -450 2120 -445 2125
rect -485 2115 -445 2120
rect -365 2120 -360 2125
rect -330 2120 -325 2150
rect -365 2115 -325 2120
rect -200 2150 -160 2155
rect -200 2120 -195 2150
rect -165 2145 -160 2150
rect -40 2150 0 2155
rect -40 2145 -35 2150
rect -165 2125 -35 2145
rect -165 2120 -160 2125
rect -200 2115 -160 2120
rect -40 2120 -35 2125
rect -5 2145 0 2150
rect 80 2150 120 2155
rect 80 2145 85 2150
rect -5 2125 85 2145
rect -5 2120 0 2125
rect -40 2115 0 2120
rect 80 2120 85 2125
rect 115 2145 120 2150
rect 200 2150 240 2155
rect 200 2145 205 2150
rect 115 2125 205 2145
rect 115 2120 120 2125
rect 80 2115 120 2120
rect 200 2120 205 2125
rect 235 2145 240 2150
rect 320 2150 360 2155
rect 320 2145 325 2150
rect 235 2125 325 2145
rect 235 2120 240 2125
rect 200 2115 240 2120
rect 320 2120 325 2125
rect 355 2145 360 2150
rect 440 2150 480 2155
rect 440 2145 445 2150
rect 355 2125 445 2145
rect 355 2120 360 2125
rect 320 2115 360 2120
rect 440 2120 445 2125
rect 475 2145 480 2150
rect 560 2150 600 2155
rect 560 2145 565 2150
rect 475 2125 565 2145
rect 475 2120 480 2125
rect 440 2115 480 2120
rect 560 2120 565 2125
rect 595 2145 600 2150
rect 680 2150 720 2155
rect 680 2145 685 2150
rect 595 2125 685 2145
rect 595 2120 600 2125
rect 560 2115 600 2120
rect 680 2120 685 2125
rect 715 2120 720 2150
rect 680 2115 720 2120
rect 970 2150 1010 2155
rect 970 2120 975 2150
rect 1005 2145 1010 2150
rect 1090 2150 1130 2155
rect 1090 2145 1095 2150
rect 1005 2125 1095 2145
rect 1005 2120 1010 2125
rect 970 2115 1010 2120
rect 1090 2120 1095 2125
rect 1125 2145 1130 2150
rect 1210 2150 1250 2155
rect 1210 2145 1215 2150
rect 1125 2125 1215 2145
rect 1125 2120 1130 2125
rect 1090 2115 1130 2120
rect 1210 2120 1215 2125
rect 1245 2145 1250 2150
rect 1330 2150 1370 2155
rect 1330 2145 1335 2150
rect 1245 2125 1335 2145
rect 1245 2120 1250 2125
rect 1210 2115 1250 2120
rect 1330 2120 1335 2125
rect 1365 2145 1370 2150
rect 1450 2150 1490 2155
rect 1450 2145 1455 2150
rect 1365 2125 1455 2145
rect 1365 2120 1370 2125
rect 1330 2115 1370 2120
rect 1450 2120 1455 2125
rect 1485 2145 1490 2150
rect 1570 2150 1610 2155
rect 1570 2145 1575 2150
rect 1485 2125 1575 2145
rect 1485 2120 1490 2125
rect 1450 2115 1490 2120
rect 1570 2120 1575 2125
rect 1605 2145 1610 2150
rect 1690 2150 1730 2155
rect 1690 2145 1695 2150
rect 1605 2125 1695 2145
rect 1605 2120 1610 2125
rect 1570 2115 1610 2120
rect 1690 2120 1695 2125
rect 1725 2145 1730 2150
rect 1850 2150 1890 2155
rect 1850 2145 1855 2150
rect 1725 2125 1855 2145
rect 1725 2120 1730 2125
rect 1690 2115 1730 2120
rect 1850 2120 1855 2125
rect 1885 2120 1890 2150
rect 1850 2115 1890 2120
rect 2015 2150 2055 2155
rect 2015 2120 2020 2150
rect 2050 2145 2055 2150
rect 2135 2150 2175 2155
rect 2135 2145 2140 2150
rect 2050 2125 2140 2145
rect 2050 2120 2055 2125
rect 2015 2115 2055 2120
rect 2135 2120 2140 2125
rect 2170 2145 2175 2150
rect 2255 2150 2295 2155
rect 2255 2145 2260 2150
rect 2170 2125 2260 2145
rect 2170 2120 2175 2125
rect 2135 2115 2175 2120
rect 2255 2120 2260 2125
rect 2290 2145 2295 2150
rect 2375 2150 2415 2155
rect 2375 2145 2380 2150
rect 2290 2125 2380 2145
rect 2290 2120 2295 2125
rect 2255 2115 2295 2120
rect 2375 2120 2380 2125
rect 2410 2145 2415 2150
rect 2495 2150 2535 2155
rect 2495 2145 2500 2150
rect 2410 2125 2500 2145
rect 2410 2120 2415 2125
rect 2375 2115 2415 2120
rect 2495 2120 2500 2125
rect 2530 2145 2535 2150
rect 2615 2150 2655 2155
rect 2615 2145 2620 2150
rect 2530 2125 2620 2145
rect 2530 2120 2535 2125
rect 2495 2115 2535 2120
rect 2615 2120 2620 2125
rect 2650 2145 2655 2150
rect 2735 2150 2775 2155
rect 2735 2145 2740 2150
rect 2650 2125 2740 2145
rect 2650 2120 2655 2125
rect 2615 2115 2655 2120
rect 2735 2120 2740 2125
rect 2770 2120 2775 2150
rect 2735 2115 2775 2120
rect -1025 1725 -985 1730
rect -1025 1695 -1020 1725
rect -990 1720 -985 1725
rect -905 1725 -865 1730
rect -905 1720 -900 1725
rect -990 1700 -900 1720
rect -990 1695 -985 1700
rect -1025 1690 -985 1695
rect -905 1695 -900 1700
rect -870 1720 -865 1725
rect -785 1725 -745 1730
rect -785 1720 -780 1725
rect -870 1700 -780 1720
rect -870 1695 -865 1700
rect -905 1690 -865 1695
rect -785 1695 -780 1700
rect -750 1720 -745 1725
rect -665 1725 -625 1730
rect -665 1720 -660 1725
rect -750 1700 -660 1720
rect -750 1695 -745 1700
rect -785 1690 -745 1695
rect -665 1695 -660 1700
rect -630 1720 -625 1725
rect -545 1725 -505 1730
rect -545 1720 -540 1725
rect -630 1700 -540 1720
rect -630 1695 -625 1700
rect -665 1690 -625 1695
rect -545 1695 -540 1700
rect -510 1720 -505 1725
rect -425 1725 -385 1730
rect -425 1720 -420 1725
rect -510 1700 -420 1720
rect -510 1695 -505 1700
rect -545 1690 -505 1695
rect -425 1695 -420 1700
rect -390 1720 -385 1725
rect -200 1725 -160 1730
rect -200 1720 -195 1725
rect -390 1700 -195 1720
rect -390 1695 -385 1700
rect -425 1690 -385 1695
rect -200 1695 -195 1700
rect -165 1695 -160 1725
rect -200 1690 -160 1695
rect 20 1725 60 1730
rect 20 1695 25 1725
rect 55 1720 60 1725
rect 140 1725 180 1730
rect 140 1720 145 1725
rect 55 1700 145 1720
rect 55 1695 60 1700
rect 20 1690 60 1695
rect 140 1695 145 1700
rect 175 1720 180 1725
rect 260 1725 300 1730
rect 260 1720 265 1725
rect 175 1700 265 1720
rect 175 1695 180 1700
rect 140 1690 180 1695
rect 260 1695 265 1700
rect 295 1720 300 1725
rect 380 1725 420 1730
rect 380 1720 385 1725
rect 295 1700 385 1720
rect 295 1695 300 1700
rect 260 1690 300 1695
rect 380 1695 385 1700
rect 415 1720 420 1725
rect 500 1725 540 1730
rect 500 1720 505 1725
rect 415 1700 505 1720
rect 415 1695 420 1700
rect 380 1690 420 1695
rect 500 1695 505 1700
rect 535 1720 540 1725
rect 620 1725 660 1730
rect 620 1720 625 1725
rect 535 1700 625 1720
rect 535 1695 540 1700
rect 500 1690 540 1695
rect 620 1695 625 1700
rect 655 1695 660 1725
rect 620 1690 660 1695
rect 1030 1725 1070 1730
rect 1030 1695 1035 1725
rect 1065 1720 1070 1725
rect 1150 1725 1190 1730
rect 1150 1720 1155 1725
rect 1065 1700 1155 1720
rect 1065 1695 1070 1700
rect 1030 1690 1070 1695
rect 1150 1695 1155 1700
rect 1185 1720 1190 1725
rect 1270 1725 1310 1730
rect 1270 1720 1275 1725
rect 1185 1700 1275 1720
rect 1185 1695 1190 1700
rect 1150 1690 1190 1695
rect 1270 1695 1275 1700
rect 1305 1720 1310 1725
rect 1390 1725 1430 1730
rect 1390 1720 1395 1725
rect 1305 1700 1395 1720
rect 1305 1695 1310 1700
rect 1270 1690 1310 1695
rect 1390 1695 1395 1700
rect 1425 1720 1430 1725
rect 1510 1725 1550 1730
rect 1510 1720 1515 1725
rect 1425 1700 1515 1720
rect 1425 1695 1430 1700
rect 1390 1690 1430 1695
rect 1510 1695 1515 1700
rect 1545 1720 1550 1725
rect 1630 1725 1670 1730
rect 1630 1720 1635 1725
rect 1545 1700 1635 1720
rect 1545 1695 1550 1700
rect 1510 1690 1550 1695
rect 1630 1695 1635 1700
rect 1665 1695 1670 1725
rect 1630 1690 1670 1695
rect 1850 1725 1890 1730
rect 1850 1695 1855 1725
rect 1885 1720 1890 1725
rect 2075 1725 2115 1730
rect 2075 1720 2080 1725
rect 1885 1700 2080 1720
rect 1885 1695 1890 1700
rect 1850 1690 1890 1695
rect 2075 1695 2080 1700
rect 2110 1720 2115 1725
rect 2195 1725 2235 1730
rect 2195 1720 2200 1725
rect 2110 1700 2200 1720
rect 2110 1695 2115 1700
rect 2075 1690 2115 1695
rect 2195 1695 2200 1700
rect 2230 1720 2235 1725
rect 2315 1725 2355 1730
rect 2315 1720 2320 1725
rect 2230 1700 2320 1720
rect 2230 1695 2235 1700
rect 2195 1690 2235 1695
rect 2315 1695 2320 1700
rect 2350 1720 2355 1725
rect 2435 1725 2475 1730
rect 2435 1720 2440 1725
rect 2350 1700 2440 1720
rect 2350 1695 2355 1700
rect 2315 1690 2355 1695
rect 2435 1695 2440 1700
rect 2470 1720 2475 1725
rect 2555 1725 2595 1730
rect 2555 1720 2560 1725
rect 2470 1700 2560 1720
rect 2470 1695 2475 1700
rect 2435 1690 2475 1695
rect 2555 1695 2560 1700
rect 2590 1720 2595 1725
rect 2675 1725 2715 1730
rect 2675 1720 2680 1725
rect 2590 1700 2680 1720
rect 2590 1695 2595 1700
rect 2555 1690 2595 1695
rect 2675 1695 2680 1700
rect 2710 1695 2715 1725
rect 2675 1690 2715 1695
rect -290 1670 -250 1675
rect -290 1640 -285 1670
rect -255 1665 -250 1670
rect 20 1670 60 1675
rect 20 1665 25 1670
rect -255 1645 25 1665
rect -255 1640 -250 1645
rect -290 1635 -250 1640
rect 20 1640 25 1645
rect 55 1640 60 1670
rect 20 1635 60 1640
rect 320 1670 360 1675
rect 320 1640 325 1670
rect 355 1665 360 1670
rect 780 1670 820 1675
rect 780 1665 785 1670
rect 355 1645 785 1665
rect 355 1640 360 1645
rect 320 1635 360 1640
rect 780 1640 785 1645
rect 815 1665 820 1670
rect 1330 1670 1370 1675
rect 1330 1665 1335 1670
rect 815 1645 1335 1665
rect 815 1640 820 1645
rect 780 1635 820 1640
rect 1330 1640 1335 1645
rect 1365 1640 1370 1670
rect 1330 1635 1370 1640
rect 1630 1670 1670 1675
rect 1630 1640 1635 1670
rect 1665 1665 1670 1670
rect 1940 1670 1980 1675
rect 1940 1665 1945 1670
rect 1665 1645 1945 1665
rect 1665 1640 1670 1645
rect 1630 1635 1670 1640
rect 1940 1640 1945 1645
rect 1975 1640 1980 1670
rect 1940 1635 1980 1640
rect -725 1625 -685 1630
rect -725 1595 -720 1625
rect -690 1620 -685 1625
rect 870 1620 875 1630
rect -690 1600 875 1620
rect 905 1620 910 1630
rect 2375 1625 2415 1630
rect 2375 1620 2380 1625
rect 905 1600 2380 1620
rect -690 1595 -685 1600
rect -725 1590 -685 1595
rect 2375 1595 2380 1600
rect 2410 1595 2415 1625
rect 2375 1590 2415 1595
rect 220 1580 260 1585
rect 220 1550 225 1580
rect 255 1575 260 1580
rect 330 1580 370 1585
rect 330 1575 335 1580
rect 255 1555 335 1575
rect 255 1550 260 1555
rect 220 1545 260 1550
rect 330 1550 335 1555
rect 365 1575 370 1580
rect 440 1580 480 1585
rect 440 1575 445 1580
rect 365 1555 445 1575
rect 365 1550 370 1555
rect 330 1545 370 1550
rect 440 1550 445 1555
rect 475 1575 480 1580
rect 550 1580 590 1585
rect 550 1575 555 1580
rect 475 1555 555 1575
rect 475 1550 480 1555
rect 440 1545 480 1550
rect 550 1550 555 1555
rect 585 1575 590 1580
rect 660 1580 700 1585
rect 660 1575 665 1580
rect 585 1555 665 1575
rect 585 1550 590 1555
rect 550 1545 590 1550
rect 660 1550 665 1555
rect 695 1575 700 1580
rect 770 1580 810 1585
rect 770 1575 775 1580
rect 695 1555 775 1575
rect 695 1550 700 1555
rect 660 1545 700 1550
rect 770 1550 775 1555
rect 805 1575 810 1580
rect 880 1580 920 1585
rect 880 1575 885 1580
rect 805 1555 885 1575
rect 805 1550 810 1555
rect 770 1545 810 1550
rect 880 1550 885 1555
rect 915 1575 920 1580
rect 990 1580 1030 1585
rect 990 1575 995 1580
rect 915 1555 995 1575
rect 915 1550 920 1555
rect 880 1545 920 1550
rect 990 1550 995 1555
rect 1025 1575 1030 1580
rect 1100 1580 1140 1585
rect 1100 1575 1105 1580
rect 1025 1555 1105 1575
rect 1025 1550 1030 1555
rect 990 1545 1030 1550
rect 1100 1550 1105 1555
rect 1135 1575 1140 1580
rect 1210 1580 1250 1585
rect 1210 1575 1215 1580
rect 1135 1555 1215 1575
rect 1135 1550 1140 1555
rect 1100 1545 1140 1550
rect 1210 1550 1215 1555
rect 1245 1575 1250 1580
rect 1320 1580 1360 1585
rect 1320 1575 1325 1580
rect 1245 1555 1325 1575
rect 1245 1550 1250 1555
rect 1210 1545 1250 1550
rect 1320 1550 1325 1555
rect 1355 1575 1360 1580
rect 1430 1580 1470 1585
rect 1430 1575 1435 1580
rect 1355 1555 1435 1575
rect 1355 1550 1360 1555
rect 1320 1545 1360 1550
rect 1430 1550 1435 1555
rect 1465 1575 1470 1580
rect 1805 1580 1845 1585
rect 1805 1575 1810 1580
rect 1465 1555 1810 1575
rect 1465 1550 1470 1555
rect 1430 1545 1470 1550
rect 1805 1550 1810 1555
rect 1840 1550 1845 1580
rect 1805 1545 1845 1550
rect -1450 1540 -1410 1545
rect -1450 1510 -1445 1540
rect -1415 1510 -1410 1540
rect -1450 1505 -1410 1510
rect 3100 1490 3140 1495
rect -1055 1485 -1015 1490
rect -1055 1455 -1050 1485
rect -1020 1480 -1015 1485
rect -945 1485 -905 1490
rect -945 1480 -940 1485
rect -1020 1460 -940 1480
rect -1020 1455 -1015 1460
rect -1055 1450 -1015 1455
rect -945 1455 -940 1460
rect -910 1480 -905 1485
rect -835 1485 -795 1490
rect -835 1480 -830 1485
rect -910 1460 -830 1480
rect -910 1455 -905 1460
rect -945 1450 -905 1455
rect -835 1455 -830 1460
rect -800 1480 -795 1485
rect -725 1485 -685 1490
rect -725 1480 -720 1485
rect -800 1460 -720 1480
rect -800 1455 -795 1460
rect -835 1450 -795 1455
rect -725 1455 -720 1460
rect -690 1480 -685 1485
rect -615 1485 -575 1490
rect -615 1480 -610 1485
rect -690 1460 -610 1480
rect -690 1455 -685 1460
rect -725 1450 -685 1455
rect -615 1455 -610 1460
rect -580 1480 -575 1485
rect -505 1485 -465 1490
rect -505 1480 -500 1485
rect -580 1460 -500 1480
rect -580 1455 -575 1460
rect -615 1450 -575 1455
rect -505 1455 -500 1460
rect -470 1480 -465 1485
rect -395 1485 -355 1490
rect -395 1480 -390 1485
rect -470 1460 -390 1480
rect -470 1455 -465 1460
rect -505 1450 -465 1455
rect -395 1455 -390 1460
rect -360 1480 -355 1485
rect -155 1485 -115 1490
rect -155 1480 -150 1485
rect -360 1460 -150 1480
rect -360 1455 -355 1460
rect -395 1450 -355 1455
rect -155 1455 -150 1460
rect -120 1455 -115 1485
rect 1805 1485 1845 1490
rect -155 1450 -115 1455
rect 275 1455 315 1460
rect 275 1425 280 1455
rect 310 1450 315 1455
rect 495 1455 535 1460
rect 495 1450 500 1455
rect 310 1430 500 1450
rect 310 1425 315 1430
rect 275 1420 315 1425
rect 495 1425 500 1430
rect 530 1450 535 1455
rect 715 1455 755 1460
rect 715 1450 720 1455
rect 530 1430 720 1450
rect 530 1425 535 1430
rect 495 1420 535 1425
rect 715 1425 720 1430
rect 750 1450 755 1455
rect 935 1455 975 1460
rect 935 1450 940 1455
rect 750 1430 940 1450
rect 750 1425 755 1430
rect 715 1420 755 1425
rect 935 1425 940 1430
rect 970 1450 975 1455
rect 1155 1455 1195 1460
rect 1155 1450 1160 1455
rect 970 1430 1160 1450
rect 970 1425 975 1430
rect 935 1420 975 1425
rect 1155 1425 1160 1430
rect 1190 1450 1195 1455
rect 1375 1455 1415 1460
rect 1375 1450 1380 1455
rect 1190 1430 1380 1450
rect 1190 1425 1195 1430
rect 1155 1420 1195 1425
rect 1375 1425 1380 1430
rect 1410 1425 1415 1455
rect 1805 1455 1810 1485
rect 1840 1480 1845 1485
rect 2045 1485 2085 1490
rect 2045 1480 2050 1485
rect 1840 1460 2050 1480
rect 1840 1455 1845 1460
rect 1805 1450 1845 1455
rect 2045 1455 2050 1460
rect 2080 1480 2085 1485
rect 2155 1485 2195 1490
rect 2155 1480 2160 1485
rect 2080 1460 2160 1480
rect 2080 1455 2085 1460
rect 2045 1450 2085 1455
rect 2155 1455 2160 1460
rect 2190 1480 2195 1485
rect 2265 1485 2305 1490
rect 2265 1480 2270 1485
rect 2190 1460 2270 1480
rect 2190 1455 2195 1460
rect 2155 1450 2195 1455
rect 2265 1455 2270 1460
rect 2300 1480 2305 1485
rect 2375 1485 2415 1490
rect 2375 1480 2380 1485
rect 2300 1460 2380 1480
rect 2300 1455 2305 1460
rect 2265 1450 2305 1455
rect 2375 1455 2380 1460
rect 2410 1480 2415 1485
rect 2485 1485 2525 1490
rect 2485 1480 2490 1485
rect 2410 1460 2490 1480
rect 2410 1455 2415 1460
rect 2375 1450 2415 1455
rect 2485 1455 2490 1460
rect 2520 1480 2525 1485
rect 2595 1485 2635 1490
rect 2595 1480 2600 1485
rect 2520 1460 2600 1480
rect 2520 1455 2525 1460
rect 2485 1450 2525 1455
rect 2595 1455 2600 1460
rect 2630 1480 2635 1485
rect 2705 1485 2745 1490
rect 2705 1480 2710 1485
rect 2630 1460 2710 1480
rect 2630 1455 2635 1460
rect 2595 1450 2635 1455
rect 2705 1455 2710 1460
rect 2740 1455 2745 1485
rect 3100 1460 3105 1490
rect 3135 1460 3140 1490
rect 3100 1455 3140 1460
rect 2705 1450 2745 1455
rect 1375 1420 1415 1425
rect 385 1400 425 1405
rect 385 1370 390 1400
rect 420 1395 425 1400
rect 605 1400 645 1405
rect 605 1395 610 1400
rect 420 1375 610 1395
rect 420 1370 425 1375
rect 385 1365 425 1370
rect 605 1370 610 1375
rect 640 1395 645 1400
rect 825 1400 865 1405
rect 825 1395 830 1400
rect 640 1375 830 1395
rect 640 1370 645 1375
rect 605 1365 645 1370
rect 825 1370 830 1375
rect 860 1395 865 1400
rect 1045 1400 1085 1405
rect 1045 1395 1050 1400
rect 860 1375 1050 1395
rect 860 1370 865 1375
rect 825 1365 865 1370
rect 1045 1370 1050 1375
rect 1080 1395 1085 1400
rect 1265 1400 1305 1405
rect 1265 1395 1270 1400
rect 1080 1375 1270 1395
rect 1080 1370 1085 1375
rect 1045 1365 1085 1370
rect 1265 1370 1270 1375
rect 1300 1370 1305 1400
rect 1265 1365 1305 1370
rect 115 1310 155 1315
rect 115 1280 120 1310
rect 150 1305 155 1310
rect 215 1310 255 1315
rect 215 1305 220 1310
rect 150 1285 220 1305
rect 150 1280 155 1285
rect 115 1275 155 1280
rect 215 1280 220 1285
rect 250 1305 255 1310
rect 325 1310 365 1315
rect 325 1305 330 1310
rect 250 1285 330 1305
rect 250 1280 255 1285
rect 215 1275 255 1280
rect 325 1280 330 1285
rect 360 1305 365 1310
rect 435 1310 475 1315
rect 435 1305 440 1310
rect 360 1285 440 1305
rect 360 1280 365 1285
rect 325 1275 365 1280
rect 435 1280 440 1285
rect 470 1305 475 1310
rect 545 1310 585 1315
rect 545 1305 550 1310
rect 470 1285 550 1305
rect 470 1280 475 1285
rect 435 1275 475 1280
rect 545 1280 550 1285
rect 580 1280 585 1310
rect 545 1275 585 1280
rect 1115 1310 1155 1315
rect 1115 1280 1120 1310
rect 1150 1305 1155 1310
rect 1215 1310 1255 1315
rect 1215 1305 1220 1310
rect 1150 1285 1220 1305
rect 1150 1280 1155 1285
rect 1115 1275 1155 1280
rect 1215 1280 1220 1285
rect 1250 1305 1255 1310
rect 1325 1310 1365 1315
rect 1325 1305 1330 1310
rect 1250 1285 1330 1305
rect 1250 1280 1255 1285
rect 1215 1275 1255 1280
rect 1325 1280 1330 1285
rect 1360 1305 1365 1310
rect 1435 1310 1475 1315
rect 1435 1305 1440 1310
rect 1360 1285 1440 1305
rect 1360 1280 1365 1285
rect 1325 1275 1365 1280
rect 1435 1280 1440 1285
rect 1470 1305 1475 1310
rect 1545 1310 1585 1315
rect 1545 1305 1550 1310
rect 1470 1285 1550 1305
rect 1470 1280 1475 1285
rect 1435 1275 1475 1280
rect 1545 1280 1550 1285
rect 1580 1280 1585 1310
rect 1545 1275 1585 1280
rect -245 1255 -205 1260
rect -245 1225 -240 1255
rect -210 1250 -205 1255
rect 71 1255 101 1260
rect -210 1230 71 1250
rect -210 1225 -205 1230
rect -245 1220 -205 1225
rect 275 1255 305 1260
rect 101 1230 275 1250
rect 71 1220 101 1225
rect 495 1255 525 1260
rect 305 1230 495 1250
rect 275 1220 305 1225
rect 1071 1255 1101 1260
rect 525 1230 1071 1250
rect 495 1220 525 1225
rect 1275 1255 1305 1260
rect 1101 1230 1275 1250
rect 1071 1220 1101 1225
rect 1495 1255 1525 1260
rect 1305 1230 1495 1250
rect 1275 1220 1305 1225
rect 1895 1255 1935 1260
rect 1895 1250 1900 1255
rect 1525 1230 1900 1250
rect 1495 1220 1525 1225
rect 1895 1225 1900 1230
rect 1930 1225 1935 1255
rect 1895 1220 1935 1225
rect -155 1195 -115 1200
rect -155 1165 -150 1195
rect -120 1190 -115 1195
rect -45 1195 -5 1200
rect -45 1190 -40 1195
rect -120 1170 -40 1190
rect -120 1165 -115 1170
rect -155 1160 -115 1165
rect -45 1165 -40 1170
rect -10 1165 -5 1195
rect -45 1160 -5 1165
rect 1695 1195 1735 1200
rect 1695 1165 1700 1195
rect 1730 1190 1735 1195
rect 1805 1195 1845 1200
rect 1805 1190 1810 1195
rect 1730 1170 1810 1190
rect 1730 1165 1735 1170
rect 1695 1160 1735 1165
rect 1805 1165 1810 1170
rect 1840 1165 1845 1195
rect 1805 1160 1845 1165
rect 204 1136 234 1141
rect -90 1110 204 1130
rect 424 1136 454 1141
rect 234 1110 424 1130
rect 204 1101 234 1106
rect 566 1136 596 1141
rect 454 1110 566 1130
rect 424 1101 454 1106
rect 1204 1136 1234 1141
rect 596 1110 1204 1130
rect 566 1101 596 1106
rect 1424 1136 1454 1141
rect 1234 1110 1424 1130
rect 1204 1101 1234 1106
rect 1566 1136 1596 1141
rect 1454 1110 1566 1130
rect 1424 1101 1454 1106
rect 1566 1101 1596 1106
rect 50 1075 90 1080
rect 50 1045 55 1075
rect 85 1070 90 1075
rect 160 1075 200 1080
rect 160 1070 165 1075
rect 85 1050 165 1070
rect 85 1045 90 1050
rect 50 1040 90 1045
rect 160 1045 165 1050
rect 195 1070 200 1075
rect 270 1075 310 1080
rect 270 1070 275 1075
rect 195 1050 275 1070
rect 195 1045 200 1050
rect 160 1040 200 1045
rect 270 1045 275 1050
rect 305 1070 310 1075
rect 380 1075 420 1080
rect 380 1070 385 1075
rect 305 1050 385 1070
rect 305 1045 310 1050
rect 270 1040 310 1045
rect 380 1045 385 1050
rect 415 1070 420 1075
rect 490 1075 530 1080
rect 490 1070 495 1075
rect 415 1050 495 1070
rect 415 1045 420 1050
rect 380 1040 420 1045
rect 490 1045 495 1050
rect 525 1070 530 1075
rect 600 1075 640 1080
rect 600 1070 605 1075
rect 525 1050 605 1070
rect 525 1045 530 1050
rect 490 1040 530 1045
rect 600 1045 605 1050
rect 635 1070 640 1075
rect 880 1075 920 1080
rect 880 1070 885 1075
rect 635 1050 885 1070
rect 635 1045 640 1050
rect 600 1040 640 1045
rect 880 1045 885 1050
rect 915 1045 920 1075
rect 880 1040 920 1045
rect 1050 1075 1090 1080
rect 1050 1045 1055 1075
rect 1085 1070 1090 1075
rect 1270 1075 1310 1080
rect 1270 1070 1275 1075
rect 1085 1050 1275 1070
rect 1085 1045 1090 1050
rect 1050 1040 1090 1045
rect 1270 1045 1275 1050
rect 1305 1070 1310 1075
rect 1490 1075 1530 1080
rect 1490 1070 1495 1075
rect 1305 1050 1495 1070
rect 1305 1045 1310 1050
rect 1270 1040 1310 1045
rect 1490 1045 1495 1050
rect 1525 1045 1530 1075
rect 1490 1040 1530 1045
rect 1160 1030 1200 1035
rect 1160 1025 1165 1030
rect 550 1020 1165 1025
rect 550 990 555 1020
rect 585 1005 1165 1020
rect 585 990 590 1005
rect 1160 1000 1165 1005
rect 1195 1025 1200 1030
rect 1380 1030 1420 1035
rect 1380 1025 1385 1030
rect 1195 1005 1385 1025
rect 1195 1000 1200 1005
rect 1160 995 1200 1000
rect 1380 1000 1385 1005
rect 1415 1025 1420 1030
rect 1600 1030 1640 1035
rect 1600 1025 1605 1030
rect 1415 1005 1605 1025
rect 1415 1000 1420 1005
rect 1380 995 1420 1000
rect 1600 1000 1605 1005
rect 1635 1000 1640 1030
rect 1600 995 1640 1000
rect 550 985 590 990
rect 660 985 700 990
rect 660 955 665 985
rect 695 980 700 985
rect 880 985 920 990
rect 880 980 885 985
rect 695 960 885 980
rect 695 955 700 960
rect 660 950 700 955
rect 880 955 885 960
rect 915 980 920 985
rect 1040 985 1080 990
rect 1040 980 1045 985
rect 915 960 1045 980
rect 915 955 920 960
rect 880 950 920 955
rect 1040 955 1045 960
rect 1075 980 1080 985
rect 1100 985 1140 990
rect 1100 980 1105 985
rect 1075 960 1105 980
rect 1075 955 1080 960
rect 1040 950 1080 955
rect 1100 955 1105 960
rect 1135 955 1140 985
rect 1100 950 1140 955
rect 550 930 590 935
rect 550 900 555 930
rect 585 925 590 930
rect 770 930 810 935
rect 770 925 775 930
rect 585 905 775 925
rect 585 900 590 905
rect 550 895 590 900
rect 770 900 775 905
rect 805 925 810 930
rect 990 930 1030 935
rect 990 925 995 930
rect 805 905 995 925
rect 805 900 810 905
rect 770 895 810 900
rect 990 900 995 905
rect 1025 925 1030 930
rect 1760 930 1800 935
rect 1760 925 1765 930
rect 1025 905 1765 925
rect 1025 900 1030 905
rect 990 895 1030 900
rect 1760 900 1765 905
rect 1795 900 1800 930
rect 1760 895 1800 900
rect -1000 810 -960 815
rect -1000 780 -995 810
rect -965 805 -960 810
rect -890 810 -850 815
rect -890 805 -885 810
rect -965 785 -885 805
rect -965 780 -960 785
rect -1000 775 -960 780
rect -890 780 -885 785
rect -855 805 -850 810
rect -780 810 -740 815
rect -780 805 -775 810
rect -855 785 -775 805
rect -855 780 -850 785
rect -890 775 -850 780
rect -780 780 -775 785
rect -745 805 -740 810
rect -670 810 -630 815
rect -670 805 -665 810
rect -745 785 -665 805
rect -745 780 -740 785
rect -780 775 -740 780
rect -670 780 -665 785
rect -635 805 -630 810
rect -560 810 -520 815
rect -560 805 -555 810
rect -635 785 -555 805
rect -635 780 -630 785
rect -670 775 -630 780
rect -560 780 -555 785
rect -525 805 -520 810
rect -450 810 -410 815
rect -450 805 -445 810
rect -525 785 -445 805
rect -525 780 -520 785
rect -560 775 -520 780
rect -450 780 -445 785
rect -415 780 -410 810
rect 495 810 535 815
rect 495 795 500 810
rect -450 775 -410 780
rect -200 780 500 795
rect 530 805 535 810
rect 605 810 645 815
rect 605 805 610 810
rect 530 785 610 805
rect 530 780 535 785
rect -200 775 535 780
rect 605 780 610 785
rect 640 805 645 810
rect 715 810 755 815
rect 715 805 720 810
rect 640 785 720 805
rect 640 780 645 785
rect 605 775 645 780
rect 715 780 720 785
rect 750 805 755 810
rect 825 810 865 815
rect 825 805 830 810
rect 750 785 830 805
rect 750 780 755 785
rect 715 775 755 780
rect 825 780 830 785
rect 860 805 865 810
rect 935 810 975 815
rect 935 805 940 810
rect 860 785 940 805
rect 860 780 865 785
rect 825 775 865 780
rect 935 780 940 785
rect 970 805 975 810
rect 1045 810 1085 815
rect 1045 805 1050 810
rect 970 785 1050 805
rect 970 780 975 785
rect 935 775 975 780
rect 1045 780 1050 785
rect 1080 805 1085 810
rect 1155 810 1195 815
rect 1155 805 1160 810
rect 1080 785 1160 805
rect 1080 780 1085 785
rect 1045 775 1085 780
rect 1155 780 1160 785
rect 1190 780 1195 810
rect 1155 775 1195 780
rect 2100 810 2140 815
rect 2100 780 2105 810
rect 2135 805 2140 810
rect 2210 810 2250 815
rect 2210 805 2215 810
rect 2135 785 2215 805
rect 2135 780 2140 785
rect 2100 775 2140 780
rect 2210 780 2215 785
rect 2245 805 2250 810
rect 2320 810 2360 815
rect 2320 805 2325 810
rect 2245 785 2325 805
rect 2245 780 2250 785
rect 2210 775 2250 780
rect 2320 780 2325 785
rect 2355 805 2360 810
rect 2430 810 2470 815
rect 2430 805 2435 810
rect 2355 785 2435 805
rect 2355 780 2360 785
rect 2320 775 2360 780
rect 2430 780 2435 785
rect 2465 805 2470 810
rect 2540 810 2580 815
rect 2540 805 2545 810
rect 2465 785 2545 805
rect 2465 780 2470 785
rect 2430 775 2470 780
rect 2540 780 2545 785
rect 2575 805 2580 810
rect 2650 810 2690 815
rect 2650 805 2655 810
rect 2575 785 2655 805
rect 2575 780 2580 785
rect 2540 775 2580 780
rect 2650 780 2655 785
rect 2685 780 2690 810
rect 2650 775 2690 780
rect -200 770 -160 775
rect -1540 760 -1500 765
rect -1540 730 -1535 760
rect -1505 755 -1500 760
rect -890 755 -885 760
rect -1505 735 -885 755
rect -1505 730 -1500 735
rect -890 730 -885 735
rect -855 730 -850 760
rect -450 730 -445 760
rect -415 755 -410 760
rect -200 755 -195 770
rect -415 740 -195 755
rect -165 740 -160 770
rect -415 735 -160 740
rect 1850 770 1890 775
rect 1850 740 1855 770
rect 1885 755 1890 770
rect 3190 760 3230 765
rect 2100 755 2105 760
rect 1885 740 2105 755
rect 1850 735 2105 740
rect -415 730 -410 735
rect 2100 730 2105 735
rect 2135 730 2140 760
rect 2540 730 2545 760
rect 2575 755 2580 760
rect 3190 755 3195 760
rect 2575 735 3195 755
rect 2575 730 2580 735
rect 3190 730 3195 735
rect 3225 730 3230 760
rect -1540 725 -1500 730
rect 3190 725 3230 730
rect -1450 715 -1410 720
rect -1450 685 -1445 715
rect -1415 710 -1410 715
rect -725 715 -685 720
rect -725 710 -720 715
rect -1415 690 -720 710
rect -1415 685 -1410 690
rect -1450 680 -1410 685
rect -725 685 -720 690
rect -690 710 -685 715
rect -290 715 -250 720
rect -290 710 -285 715
rect -690 690 -285 710
rect -690 685 -685 690
rect -725 680 -685 685
rect -290 685 -285 690
rect -255 710 -250 715
rect 30 715 70 720
rect 30 710 35 715
rect -255 690 35 710
rect -255 685 -250 690
rect -290 680 -250 685
rect 30 685 35 690
rect 65 710 70 715
rect 140 715 180 720
rect 140 710 145 715
rect 65 690 145 710
rect 65 685 70 690
rect 30 680 70 685
rect 140 685 145 690
rect 175 710 180 715
rect 250 715 290 720
rect 250 710 255 715
rect 175 690 255 710
rect 175 685 180 690
rect 140 680 180 685
rect 250 685 255 690
rect 285 710 290 715
rect 360 715 400 720
rect 360 710 365 715
rect 285 690 365 710
rect 285 685 290 690
rect 250 680 290 685
rect 360 685 365 690
rect 395 710 400 715
rect 470 715 510 720
rect 470 710 475 715
rect 395 690 475 710
rect 395 685 400 690
rect 360 680 400 685
rect 470 685 475 690
rect 505 710 510 715
rect 580 715 620 720
rect 580 710 585 715
rect 505 690 585 710
rect 505 685 510 690
rect 470 680 510 685
rect 580 685 585 690
rect 615 685 620 715
rect 580 680 620 685
rect 1070 715 1110 720
rect 1070 685 1075 715
rect 1105 710 1110 715
rect 1180 715 1220 720
rect 1180 710 1185 715
rect 1105 690 1185 710
rect 1105 685 1110 690
rect 1070 680 1110 685
rect 1180 685 1185 690
rect 1215 710 1220 715
rect 1290 715 1330 720
rect 1290 710 1295 715
rect 1215 690 1295 710
rect 1215 685 1220 690
rect 1180 680 1220 685
rect 1290 685 1295 690
rect 1325 710 1330 715
rect 1400 715 1440 720
rect 1400 710 1405 715
rect 1325 690 1405 710
rect 1325 685 1330 690
rect 1290 680 1330 685
rect 1400 685 1405 690
rect 1435 710 1440 715
rect 1510 715 1550 720
rect 1510 710 1515 715
rect 1435 690 1515 710
rect 1435 685 1440 690
rect 1400 680 1440 685
rect 1510 685 1515 690
rect 1545 710 1550 715
rect 1620 715 1660 720
rect 1620 710 1625 715
rect 1545 690 1625 710
rect 1545 685 1550 690
rect 1510 680 1550 685
rect 1620 685 1625 690
rect 1655 710 1660 715
rect 1940 715 1980 720
rect 1940 710 1945 715
rect 1655 690 1945 710
rect 1655 685 1660 690
rect 1620 680 1660 685
rect 1940 685 1945 690
rect 1975 710 1980 715
rect 2375 715 2415 720
rect 2375 710 2380 715
rect 1975 690 2380 710
rect 1975 685 1980 690
rect 1940 680 1980 685
rect 2375 685 2380 690
rect 2410 710 2415 715
rect 3100 715 3140 720
rect 3100 710 3105 715
rect 2410 690 3105 710
rect 2410 685 2415 690
rect 2375 680 2415 685
rect 3100 685 3105 690
rect 3135 685 3140 715
rect 3100 680 3140 685
rect -1065 670 -1025 675
rect -1065 640 -1060 670
rect -1030 640 -1025 670
rect -1065 635 -1025 640
rect -1000 670 -960 675
rect -1000 640 -995 670
rect -965 665 -960 670
rect -890 670 -850 675
rect -890 665 -885 670
rect -965 645 -885 665
rect -965 640 -960 645
rect -1000 635 -960 640
rect -890 640 -885 645
rect -855 665 -850 670
rect -780 670 -740 675
rect -780 665 -775 670
rect -855 645 -775 665
rect -855 640 -850 645
rect -890 635 -850 640
rect -780 640 -775 645
rect -745 665 -740 670
rect -670 670 -630 675
rect -670 665 -665 670
rect -745 645 -665 665
rect -745 640 -740 645
rect -780 635 -740 640
rect -670 640 -665 645
rect -635 665 -630 670
rect -560 670 -520 675
rect -560 665 -555 670
rect -635 645 -555 665
rect -635 640 -630 645
rect -670 635 -630 640
rect -560 640 -555 645
rect -525 665 -520 670
rect -450 670 -410 675
rect -450 665 -445 670
rect -525 645 -445 665
rect -525 640 -520 645
rect -560 635 -520 640
rect -450 640 -445 645
rect -415 640 -410 670
rect -450 635 -410 640
rect -385 670 -345 675
rect -385 640 -380 670
rect -350 665 -345 670
rect -155 670 -115 675
rect -155 665 -150 670
rect -350 645 -150 665
rect -350 640 -345 645
rect -385 635 -345 640
rect -155 640 -150 645
rect -120 640 -115 670
rect 1805 670 1845 675
rect -155 635 -115 640
rect -100 660 -60 665
rect -100 630 -95 660
rect -65 655 -60 660
rect 310 660 340 665
rect -65 635 310 655
rect -65 630 -60 635
rect -100 625 -60 630
rect 1350 660 1380 665
rect 340 635 1350 655
rect 310 625 340 630
rect 1805 640 1810 670
rect 1840 665 1845 670
rect 2035 670 2075 675
rect 2035 665 2040 670
rect 1840 645 2040 665
rect 1840 640 1845 645
rect 1805 635 1845 640
rect 2035 640 2040 645
rect 2070 640 2075 670
rect 2035 635 2075 640
rect 2100 670 2140 675
rect 2100 640 2105 670
rect 2135 665 2140 670
rect 2210 670 2250 675
rect 2210 665 2215 670
rect 2135 645 2215 665
rect 2135 640 2140 645
rect 2100 635 2140 640
rect 2210 640 2215 645
rect 2245 665 2250 670
rect 2320 670 2360 675
rect 2320 665 2325 670
rect 2245 645 2325 665
rect 2245 640 2250 645
rect 2210 635 2250 640
rect 2320 640 2325 645
rect 2355 665 2360 670
rect 2430 670 2470 675
rect 2430 665 2435 670
rect 2355 645 2435 665
rect 2355 640 2360 645
rect 2320 635 2360 640
rect 2430 640 2435 645
rect 2465 665 2470 670
rect 2540 670 2580 675
rect 2540 665 2545 670
rect 2465 645 2545 665
rect 2465 640 2470 645
rect 2430 635 2470 640
rect 2540 640 2545 645
rect 2575 665 2580 670
rect 2650 670 2690 675
rect 2650 665 2655 670
rect 2575 645 2655 665
rect 2575 640 2580 645
rect 2540 635 2580 640
rect 2650 640 2655 645
rect 2685 640 2690 670
rect 2650 635 2690 640
rect 2715 670 2755 675
rect 2715 640 2720 670
rect 2750 640 2755 670
rect 2715 635 2755 640
rect 1350 625 1380 630
rect -25 435 15 440
rect -25 405 -20 435
rect 10 430 15 435
rect 635 435 675 440
rect 635 430 640 435
rect 10 410 640 430
rect 10 405 15 410
rect -25 400 15 405
rect 635 405 640 410
rect 670 430 675 435
rect 1015 435 1055 440
rect 1015 430 1020 435
rect 670 410 1020 430
rect 670 405 675 410
rect 635 400 675 405
rect 1015 405 1020 410
rect 1050 430 1055 435
rect 1675 435 1715 440
rect 1675 430 1680 435
rect 1050 410 1680 430
rect 1050 405 1055 410
rect 1015 400 1055 405
rect 1675 405 1680 410
rect 1710 430 1715 435
rect 1850 435 1890 440
rect 1850 430 1855 435
rect 1710 410 1855 430
rect 1710 405 1715 410
rect 1675 400 1715 405
rect 1850 405 1855 410
rect 1885 405 1890 435
rect 1850 400 1890 405
rect -1190 395 -1150 400
rect -1190 365 -1185 395
rect -1155 390 -1150 395
rect -945 395 -905 400
rect -945 390 -940 395
rect -1155 370 -940 390
rect -1155 365 -1150 370
rect -1190 360 -1150 365
rect -945 365 -940 370
rect -910 390 -905 395
rect -835 395 -795 400
rect -835 390 -830 395
rect -910 370 -830 390
rect -910 365 -905 370
rect -945 360 -905 365
rect -835 365 -830 370
rect -800 390 -795 395
rect -725 395 -685 400
rect -725 390 -720 395
rect -800 370 -720 390
rect -800 365 -795 370
rect -835 360 -795 365
rect -725 365 -720 370
rect -690 390 -685 395
rect -615 395 -575 400
rect -615 390 -610 395
rect -690 370 -610 390
rect -690 365 -685 370
rect -725 360 -685 365
rect -615 365 -610 370
rect -580 390 -575 395
rect -505 395 -465 400
rect -505 390 -500 395
rect -580 370 -500 390
rect -580 365 -575 370
rect -615 360 -575 365
rect -505 365 -500 370
rect -470 365 -465 395
rect 2155 395 2195 400
rect -505 360 -465 365
rect 85 375 125 380
rect -1545 350 -1495 360
rect -1545 320 -1535 350
rect -1505 320 -1495 350
rect 85 345 90 375
rect 120 370 125 375
rect 195 375 235 380
rect 195 370 200 375
rect 120 350 200 370
rect 120 345 125 350
rect -1545 310 -1495 320
rect -670 340 -630 345
rect -670 310 -665 340
rect -635 335 -630 340
rect -290 340 -250 345
rect 85 340 125 345
rect 195 345 200 350
rect 230 370 235 375
rect 305 375 345 380
rect 305 370 310 375
rect 230 350 310 370
rect 230 345 235 350
rect 195 340 235 345
rect 305 345 310 350
rect 340 370 345 375
rect 415 375 455 380
rect 415 370 420 375
rect 340 350 420 370
rect 340 345 345 350
rect 305 340 345 345
rect 415 345 420 350
rect 450 370 455 375
rect 525 375 565 380
rect 525 370 530 375
rect 450 350 530 370
rect 450 345 455 350
rect 415 340 455 345
rect 525 345 530 350
rect 560 345 565 375
rect 525 340 565 345
rect 1125 375 1165 380
rect 1125 345 1130 375
rect 1160 370 1165 375
rect 1235 375 1275 380
rect 1235 370 1240 375
rect 1160 350 1240 370
rect 1160 345 1165 350
rect 1125 340 1165 345
rect 1235 345 1240 350
rect 1270 370 1275 375
rect 1345 375 1385 380
rect 1345 370 1350 375
rect 1270 350 1350 370
rect 1270 345 1275 350
rect 1235 340 1275 345
rect 1345 345 1350 350
rect 1380 370 1385 375
rect 1455 375 1495 380
rect 1455 370 1460 375
rect 1380 350 1460 370
rect 1380 345 1385 350
rect 1345 340 1385 345
rect 1455 345 1460 350
rect 1490 370 1495 375
rect 1565 375 1605 380
rect 1565 370 1570 375
rect 1490 350 1570 370
rect 1490 345 1495 350
rect 1455 340 1495 345
rect 1565 345 1570 350
rect 1600 345 1605 375
rect 2155 365 2160 395
rect 2190 390 2195 395
rect 2265 395 2305 400
rect 2265 390 2270 395
rect 2190 370 2270 390
rect 2190 365 2195 370
rect 2155 360 2195 365
rect 2265 365 2270 370
rect 2300 390 2305 395
rect 2375 395 2415 400
rect 2375 390 2380 395
rect 2300 370 2380 390
rect 2300 365 2305 370
rect 2265 360 2305 365
rect 2375 365 2380 370
rect 2410 390 2415 395
rect 2485 395 2525 400
rect 2485 390 2490 395
rect 2410 370 2490 390
rect 2410 365 2415 370
rect 2375 360 2415 365
rect 2485 365 2490 370
rect 2520 390 2525 395
rect 2595 395 2635 400
rect 2595 390 2600 395
rect 2520 370 2600 390
rect 2520 365 2525 370
rect 2485 360 2525 365
rect 2595 365 2600 370
rect 2630 390 2635 395
rect 2840 395 2880 400
rect 2840 390 2845 395
rect 2630 370 2845 390
rect 2630 365 2635 370
rect 2595 360 2635 365
rect 2840 365 2845 370
rect 2875 365 2880 395
rect 2840 360 2880 365
rect 3185 350 3235 360
rect 1565 340 1605 345
rect 1940 340 1980 345
rect -290 335 -285 340
rect -635 315 -285 335
rect -635 310 -630 315
rect -670 305 -630 310
rect -290 310 -285 315
rect -255 310 -250 340
rect -290 305 -250 310
rect 1940 310 1945 340
rect 1975 335 1980 340
rect 2320 340 2360 345
rect 2320 335 2325 340
rect 1975 315 2325 335
rect 1975 310 1980 315
rect 1940 305 1980 310
rect 2320 310 2325 315
rect 2355 310 2360 340
rect 3185 320 3195 350
rect 3225 320 3235 350
rect 3185 310 3235 320
rect 2320 305 2360 310
rect -1145 285 -1105 290
rect -1145 255 -1140 285
rect -1110 280 -1105 285
rect -945 285 -905 290
rect -945 280 -940 285
rect -1110 260 -940 280
rect -1110 255 -1105 260
rect -1145 250 -1105 255
rect -945 255 -940 260
rect -910 280 -905 285
rect -835 285 -795 290
rect -835 280 -830 285
rect -910 260 -830 280
rect -910 255 -905 260
rect -945 250 -905 255
rect -835 255 -830 260
rect -800 280 -795 285
rect -725 285 -685 290
rect -725 280 -720 285
rect -800 260 -720 280
rect -800 255 -795 260
rect -835 250 -795 255
rect -725 255 -720 260
rect -690 280 -685 285
rect -615 285 -575 290
rect -615 280 -610 285
rect -690 260 -610 280
rect -690 255 -685 260
rect -725 250 -685 255
rect -615 255 -610 260
rect -580 280 -575 285
rect -505 285 -465 290
rect -505 280 -500 285
rect -580 260 -500 280
rect -580 255 -575 260
rect -615 250 -575 255
rect -505 255 -500 260
rect -470 255 -465 285
rect -505 250 -465 255
rect 2155 285 2195 290
rect 2155 255 2160 285
rect 2190 280 2195 285
rect 2265 285 2305 290
rect 2265 280 2270 285
rect 2190 260 2270 280
rect 2190 255 2195 260
rect 2155 250 2195 255
rect 2265 255 2270 260
rect 2300 280 2305 285
rect 2375 285 2415 290
rect 2375 280 2380 285
rect 2300 260 2380 280
rect 2300 255 2305 260
rect 2265 250 2305 255
rect 2375 255 2380 260
rect 2410 280 2415 285
rect 2485 285 2525 290
rect 2485 280 2490 285
rect 2410 260 2490 280
rect 2410 255 2415 260
rect 2375 250 2415 255
rect 2485 255 2490 260
rect 2520 280 2525 285
rect 2595 285 2635 290
rect 2595 280 2600 285
rect 2520 260 2600 280
rect 2520 255 2525 260
rect 2485 250 2525 255
rect 2595 255 2600 260
rect 2630 280 2635 285
rect 2795 285 2835 290
rect 2795 280 2800 285
rect 2630 260 2800 280
rect 2630 255 2635 260
rect 2595 250 2635 255
rect 2795 255 2800 260
rect 2830 255 2835 285
rect 2795 250 2835 255
rect 310 240 340 245
rect 30 230 70 235
rect 30 200 35 230
rect 65 225 70 230
rect 140 230 180 235
rect 140 225 145 230
rect 65 205 145 225
rect 65 200 70 205
rect 30 195 70 200
rect 140 200 145 205
rect 175 225 180 230
rect 250 230 290 235
rect 250 225 255 230
rect 175 205 255 225
rect 175 200 180 205
rect 140 195 180 200
rect 250 200 255 205
rect 285 225 290 230
rect 285 210 310 225
rect 1350 240 1380 245
rect 360 230 400 235
rect 360 225 365 230
rect 340 210 365 225
rect 285 205 365 210
rect 285 200 290 205
rect 250 195 290 200
rect 360 200 365 205
rect 395 225 400 230
rect 470 230 510 235
rect 470 225 475 230
rect 395 205 475 225
rect 395 200 400 205
rect 360 195 400 200
rect 470 200 475 205
rect 505 225 510 230
rect 580 230 620 235
rect 580 225 585 230
rect 505 205 585 225
rect 505 200 510 205
rect 470 195 510 200
rect 580 200 585 205
rect 615 200 620 230
rect 580 195 620 200
rect 1070 230 1110 235
rect 1070 200 1075 230
rect 1105 225 1110 230
rect 1180 230 1220 235
rect 1180 225 1185 230
rect 1105 205 1185 225
rect 1105 200 1110 205
rect 1070 195 1110 200
rect 1180 200 1185 205
rect 1215 225 1220 230
rect 1290 230 1330 235
rect 1290 225 1295 230
rect 1215 205 1295 225
rect 1215 200 1220 205
rect 1180 195 1220 200
rect 1290 200 1295 205
rect 1325 225 1330 230
rect 1325 210 1350 225
rect 1400 230 1440 235
rect 1400 225 1405 230
rect 1380 210 1405 225
rect 1325 205 1405 210
rect 1325 200 1330 205
rect 1290 195 1330 200
rect 1400 200 1405 205
rect 1435 225 1440 230
rect 1510 230 1550 235
rect 1510 225 1515 230
rect 1435 205 1515 225
rect 1435 200 1440 205
rect 1400 195 1440 200
rect 1510 200 1515 205
rect 1545 225 1550 230
rect 1620 230 1660 235
rect 1620 225 1625 230
rect 1545 205 1625 225
rect 1545 200 1550 205
rect 1510 195 1550 200
rect 1620 200 1625 205
rect 1655 200 1660 230
rect 1620 195 1660 200
rect 310 180 340 185
rect -25 155 310 175
rect 795 180 825 185
rect 340 155 795 175
rect 310 145 340 150
rect 795 145 825 150
rect 848 180 878 185
rect 1350 180 1380 185
rect 878 155 1350 175
rect 848 145 878 150
rect 1380 155 1715 175
rect 1350 145 1380 150
rect 85 -40 125 -35
rect -30 -65 10 -45
rect 85 -70 90 -40
rect 120 -45 125 -40
rect 195 -40 235 -35
rect 195 -45 200 -40
rect 120 -65 200 -45
rect 120 -70 125 -65
rect 85 -75 125 -70
rect 195 -70 200 -65
rect 230 -45 235 -40
rect 305 -40 345 -35
rect 305 -45 310 -40
rect 230 -65 310 -45
rect 230 -70 235 -65
rect 195 -75 235 -70
rect 305 -70 310 -65
rect 340 -45 345 -40
rect 415 -40 455 -35
rect 415 -45 420 -40
rect 340 -65 420 -45
rect 340 -70 345 -65
rect 305 -75 345 -70
rect 415 -70 420 -65
rect 450 -45 455 -40
rect 525 -40 565 -35
rect 525 -45 530 -40
rect 450 -65 530 -45
rect 450 -70 455 -65
rect 415 -75 455 -70
rect 525 -70 530 -65
rect 560 -45 565 -40
rect 1125 -40 1165 -35
rect 1125 -45 1130 -40
rect 560 -65 1130 -45
rect 560 -70 565 -65
rect 525 -75 565 -70
rect 1125 -70 1130 -65
rect 1160 -45 1165 -40
rect 1235 -40 1275 -35
rect 1235 -45 1240 -40
rect 1160 -65 1240 -45
rect 1160 -70 1165 -65
rect 1125 -75 1165 -70
rect 1235 -70 1240 -65
rect 1270 -45 1275 -40
rect 1345 -40 1385 -35
rect 1345 -45 1350 -40
rect 1270 -65 1350 -45
rect 1270 -70 1275 -65
rect 1235 -75 1275 -70
rect 1345 -70 1350 -65
rect 1380 -45 1385 -40
rect 1455 -40 1495 -35
rect 1455 -45 1460 -40
rect 1380 -65 1460 -45
rect 1380 -70 1385 -65
rect 1345 -75 1385 -70
rect 1455 -70 1460 -65
rect 1490 -45 1495 -40
rect 1565 -40 1605 -35
rect 1565 -45 1570 -40
rect 1490 -65 1570 -45
rect 1490 -70 1495 -65
rect 1455 -75 1495 -70
rect 1565 -70 1570 -65
rect 1600 -70 1605 -40
rect 1565 -75 1605 -70
rect -1410 -120 -1406 -85
rect -1379 -120 -1346 -85
rect -1319 -120 -1315 -85
rect -1290 -120 -1286 -85
rect -1259 -120 -1255 -85
rect -1230 -120 -1226 -85
rect -1199 -95 -1195 -85
rect -1145 -90 -1105 -85
rect -1145 -95 -1140 -90
rect -1199 -115 -1140 -95
rect -1199 -120 -1195 -115
rect -1145 -120 -1140 -115
rect -1110 -120 -1105 -90
rect -1145 -125 -1105 -120
rect -1000 -90 -960 -85
rect -1000 -120 -995 -90
rect -965 -95 -960 -90
rect -890 -90 -850 -85
rect -890 -95 -885 -90
rect -965 -115 -885 -95
rect -965 -120 -960 -115
rect -1000 -125 -960 -120
rect -890 -120 -885 -115
rect -855 -95 -850 -90
rect -780 -90 -740 -85
rect -780 -95 -775 -90
rect -855 -115 -775 -95
rect -855 -120 -850 -115
rect -890 -125 -850 -120
rect -780 -120 -775 -115
rect -745 -95 -740 -90
rect -670 -90 -630 -85
rect -670 -95 -665 -90
rect -745 -115 -665 -95
rect -745 -120 -740 -115
rect -780 -125 -740 -120
rect -670 -120 -665 -115
rect -635 -95 -630 -90
rect -560 -90 -520 -85
rect -560 -95 -555 -90
rect -635 -115 -555 -95
rect -635 -120 -630 -115
rect -670 -125 -630 -120
rect -560 -120 -555 -115
rect -525 -95 -520 -90
rect -450 -90 -410 -85
rect -450 -95 -445 -90
rect -525 -115 -445 -95
rect -525 -120 -520 -115
rect -560 -125 -520 -120
rect -450 -120 -445 -115
rect -415 -95 -410 -90
rect -155 -90 -115 -85
rect 1805 -90 1845 -85
rect -155 -95 -150 -90
rect -415 -115 -150 -95
rect -415 -120 -410 -115
rect -450 -125 -410 -120
rect -155 -120 -150 -115
rect -120 -120 -115 -90
rect -155 -125 -115 -120
rect 760 -95 800 -90
rect 760 -125 765 -95
rect 795 -100 800 -95
rect 890 -95 930 -90
rect 890 -100 895 -95
rect 795 -120 895 -100
rect 795 -125 800 -120
rect 760 -130 800 -125
rect 890 -125 895 -120
rect 925 -125 930 -95
rect 1805 -120 1810 -90
rect 1840 -95 1845 -90
rect 2100 -90 2140 -85
rect 2100 -95 2105 -90
rect 1840 -115 2105 -95
rect 1840 -120 1845 -115
rect 1805 -125 1845 -120
rect 2100 -120 2105 -115
rect 2135 -95 2140 -90
rect 2210 -90 2250 -85
rect 2210 -95 2215 -90
rect 2135 -115 2215 -95
rect 2135 -120 2140 -115
rect 2100 -125 2140 -120
rect 2210 -120 2215 -115
rect 2245 -95 2250 -90
rect 2320 -90 2360 -85
rect 2320 -95 2325 -90
rect 2245 -115 2325 -95
rect 2245 -120 2250 -115
rect 2210 -125 2250 -120
rect 2320 -120 2325 -115
rect 2355 -95 2360 -90
rect 2430 -90 2470 -85
rect 2430 -95 2435 -90
rect 2355 -115 2435 -95
rect 2355 -120 2360 -115
rect 2320 -125 2360 -120
rect 2430 -120 2435 -115
rect 2465 -95 2470 -90
rect 2540 -90 2580 -85
rect 2540 -95 2545 -90
rect 2465 -115 2545 -95
rect 2465 -120 2470 -115
rect 2430 -125 2470 -120
rect 2540 -120 2545 -115
rect 2575 -95 2580 -90
rect 2650 -90 2690 -85
rect 2650 -95 2655 -90
rect 2575 -115 2655 -95
rect 2575 -120 2580 -115
rect 2540 -125 2580 -120
rect 2650 -120 2655 -115
rect 2685 -120 2690 -90
rect 2650 -125 2690 -120
rect 2795 -90 2835 -85
rect 2795 -120 2800 -90
rect 2830 -95 2835 -90
rect 2885 -95 2889 -85
rect 2830 -115 2889 -95
rect 2830 -120 2835 -115
rect 2885 -120 2889 -115
rect 2916 -120 2920 -85
rect 2945 -120 2949 -85
rect 2976 -120 2980 -85
rect 3005 -120 3009 -85
rect 3036 -120 3069 -85
rect 3096 -120 3100 -85
rect 2795 -125 2835 -120
rect 890 -130 930 -125
rect -25 -140 15 -135
rect -1290 -145 -1255 -140
rect -1190 -145 -1150 -140
rect -1190 -150 -1185 -145
rect -1255 -170 -1185 -150
rect -1290 -180 -1255 -175
rect -1190 -175 -1185 -170
rect -1155 -175 -1150 -145
rect -1190 -180 -1150 -175
rect -1065 -145 -1025 -140
rect -1065 -175 -1060 -145
rect -1030 -150 -1025 -145
rect -385 -145 -345 -140
rect -385 -150 -380 -145
rect -1030 -170 -380 -150
rect -1030 -175 -1025 -170
rect -1065 -180 -1025 -175
rect -385 -175 -380 -170
rect -350 -150 -345 -145
rect -200 -145 -160 -140
rect -200 -150 -195 -145
rect -350 -170 -195 -150
rect -350 -175 -345 -170
rect -200 -175 -195 -170
rect -165 -175 -160 -145
rect -25 -170 -20 -140
rect 10 -145 15 -140
rect 675 -140 715 -135
rect 675 -145 680 -140
rect 10 -165 680 -145
rect 10 -170 15 -165
rect -25 -175 15 -170
rect 675 -170 680 -165
rect 710 -145 715 -140
rect 975 -140 1015 -135
rect 975 -145 980 -140
rect 710 -165 980 -145
rect 710 -170 715 -165
rect 675 -175 715 -170
rect 975 -170 980 -165
rect 1010 -145 1015 -140
rect 1675 -140 1715 -135
rect 1675 -145 1680 -140
rect 1010 -165 1680 -145
rect 1010 -170 1015 -165
rect 975 -175 1015 -170
rect 1675 -170 1680 -165
rect 1710 -145 1715 -140
rect 1850 -145 1890 -140
rect 1710 -165 1855 -145
rect 1710 -170 1715 -165
rect 1675 -175 1715 -170
rect 1850 -175 1855 -165
rect 1885 -150 1890 -145
rect 2035 -145 2075 -140
rect 2035 -150 2040 -145
rect 1885 -170 2040 -150
rect 1885 -175 1890 -170
rect 2035 -175 2040 -170
rect 2070 -150 2075 -145
rect 2715 -145 2755 -140
rect 2715 -150 2720 -145
rect 2070 -170 2720 -150
rect 2070 -175 2075 -170
rect -385 -180 -345 -175
rect 2035 -180 2075 -175
rect 2715 -175 2720 -170
rect 2750 -175 2755 -145
rect 2715 -180 2755 -175
rect 2840 -145 2880 -140
rect 2840 -175 2845 -145
rect 2875 -150 2880 -145
rect 2945 -145 2980 -140
rect 2875 -170 2945 -150
rect 2875 -175 2880 -170
rect 2840 -180 2880 -175
rect 2945 -180 2980 -175
rect -1410 -190 -1375 -185
rect 3065 -190 3100 -185
rect -245 -195 -240 -190
rect -1375 -215 -240 -195
rect -1410 -225 -1375 -220
rect -245 -220 -240 -215
rect -210 -220 -205 -190
rect -245 -225 -205 -220
rect 75 -195 115 -190
rect 75 -225 80 -195
rect 110 -200 115 -195
rect 710 -195 750 -190
rect 710 -200 715 -195
rect 110 -220 715 -200
rect 110 -225 115 -220
rect 75 -230 115 -225
rect 710 -225 715 -220
rect 745 -225 750 -195
rect 1895 -220 1900 -190
rect 1930 -195 1935 -190
rect 1930 -215 3065 -195
rect 1930 -220 1935 -215
rect 1895 -225 1935 -220
rect 3065 -225 3100 -220
rect 710 -230 750 -225
rect -1210 -240 -1175 -235
rect -625 -240 -585 -235
rect -625 -245 -620 -240
rect -1175 -265 -620 -245
rect -1210 -275 -1175 -270
rect -625 -270 -620 -265
rect -590 -245 -585 -240
rect 2275 -240 2315 -235
rect 2275 -245 2280 -240
rect -590 -265 2280 -245
rect -590 -270 -585 -265
rect -625 -275 -585 -270
rect 2275 -270 2280 -265
rect 2310 -245 2315 -240
rect 2865 -240 2900 -235
rect 2310 -265 2865 -245
rect 2310 -270 2315 -265
rect 2275 -275 2315 -270
rect 2865 -275 2900 -270
rect 270 -295 310 -290
rect -1540 -300 -1500 -295
rect -1540 -330 -1535 -300
rect -1505 -305 -1500 -300
rect -1150 -300 -1115 -295
rect -1505 -325 -1150 -305
rect -1505 -330 -1500 -325
rect -1540 -335 -1500 -330
rect -925 -300 -885 -295
rect -925 -305 -920 -300
rect -1115 -325 -920 -305
rect -1150 -335 -1115 -330
rect -925 -330 -920 -325
rect -890 -305 -885 -300
rect -725 -300 -685 -295
rect -725 -305 -720 -300
rect -890 -325 -720 -305
rect -890 -330 -885 -325
rect -925 -335 -885 -330
rect -725 -330 -720 -325
rect -690 -305 -685 -300
rect -525 -300 -485 -295
rect -525 -305 -520 -300
rect -690 -325 -520 -305
rect -690 -330 -685 -325
rect -725 -335 -685 -330
rect -525 -330 -520 -325
rect -490 -330 -485 -300
rect 270 -325 275 -295
rect 305 -300 310 -295
rect 825 -295 865 -290
rect 825 -300 830 -295
rect 305 -320 830 -300
rect 305 -325 310 -320
rect 270 -330 310 -325
rect 825 -325 830 -320
rect 860 -325 865 -295
rect 825 -330 865 -325
rect 1330 -295 1370 -290
rect 1330 -325 1335 -295
rect 1365 -300 1370 -295
rect 1760 -295 1800 -290
rect 1760 -300 1765 -295
rect 1365 -320 1765 -300
rect 1365 -325 1370 -320
rect 1330 -330 1370 -325
rect 1760 -325 1765 -320
rect 1795 -325 1800 -295
rect 1760 -330 1800 -325
rect 2175 -300 2215 -295
rect 2175 -330 2180 -300
rect 2210 -305 2215 -300
rect 2375 -300 2415 -295
rect 2375 -305 2380 -300
rect 2210 -325 2380 -305
rect 2210 -330 2215 -325
rect -525 -335 -485 -330
rect 2175 -335 2215 -330
rect 2375 -330 2380 -325
rect 2410 -305 2415 -300
rect 2575 -300 2615 -295
rect 2575 -305 2580 -300
rect 2410 -325 2580 -305
rect 2410 -330 2415 -325
rect 2375 -335 2415 -330
rect 2575 -330 2580 -325
rect 2610 -305 2615 -300
rect 2805 -300 2840 -295
rect 2610 -325 2805 -305
rect 2610 -330 2615 -325
rect 2575 -335 2615 -330
rect 3190 -300 3230 -295
rect 3190 -305 3195 -300
rect 2840 -325 3195 -305
rect 2805 -335 2840 -330
rect 3190 -330 3195 -325
rect 3225 -330 3230 -300
rect 3190 -335 3230 -330
rect 380 -350 420 -345
rect 380 -380 385 -350
rect 415 -355 420 -350
rect 490 -350 530 -345
rect 490 -355 495 -350
rect 415 -375 495 -355
rect 415 -380 420 -375
rect -1210 -415 -1206 -380
rect -1179 -415 -1175 -380
rect -1150 -415 -1146 -380
rect -1119 -415 -1115 -380
rect 380 -385 420 -380
rect 490 -380 495 -375
rect 525 -355 530 -350
rect 600 -350 640 -345
rect 600 -355 605 -350
rect 525 -375 605 -355
rect 525 -380 530 -375
rect 490 -385 530 -380
rect 600 -380 605 -375
rect 635 -355 640 -350
rect 710 -350 750 -345
rect 710 -355 715 -350
rect 635 -375 715 -355
rect 635 -380 640 -375
rect 600 -385 640 -380
rect 710 -380 715 -375
rect 745 -355 750 -350
rect 820 -350 860 -345
rect 820 -355 825 -350
rect 745 -375 825 -355
rect 745 -380 750 -375
rect 710 -385 750 -380
rect 820 -380 825 -375
rect 855 -355 860 -350
rect 930 -350 970 -345
rect 930 -355 935 -350
rect 855 -375 935 -355
rect 855 -380 860 -375
rect 820 -385 860 -380
rect 930 -380 935 -375
rect 965 -355 970 -350
rect 1040 -350 1080 -345
rect 1040 -355 1045 -350
rect 965 -375 1045 -355
rect 965 -380 970 -375
rect 930 -385 970 -380
rect 1040 -380 1045 -375
rect 1075 -355 1080 -350
rect 1150 -350 1190 -345
rect 1150 -355 1155 -350
rect 1075 -375 1155 -355
rect 1075 -380 1080 -375
rect 1040 -385 1080 -380
rect 1150 -380 1155 -375
rect 1185 -355 1190 -350
rect 1260 -350 1300 -345
rect 1260 -355 1265 -350
rect 1185 -375 1265 -355
rect 1185 -380 1190 -375
rect 1150 -385 1190 -380
rect 1260 -380 1265 -375
rect 1295 -355 1300 -350
rect 1385 -350 1425 -345
rect 1385 -355 1390 -350
rect 1295 -375 1390 -355
rect 1295 -380 1300 -375
rect 1260 -385 1300 -380
rect 1385 -380 1390 -375
rect 1420 -380 1425 -350
rect 1385 -385 1425 -380
rect 2805 -415 2809 -380
rect 2836 -415 2840 -380
rect 2865 -415 2869 -380
rect 2896 -415 2900 -380
rect 150 -675 190 -670
rect 150 -705 155 -675
rect 185 -680 190 -675
rect 215 -675 255 -670
rect 215 -680 220 -675
rect 185 -700 220 -680
rect 185 -705 190 -700
rect 150 -710 190 -705
rect 215 -705 220 -700
rect 250 -680 255 -675
rect 325 -675 365 -670
rect 325 -680 330 -675
rect 250 -700 330 -680
rect 250 -705 255 -700
rect 215 -710 255 -705
rect 325 -705 330 -700
rect 360 -680 365 -675
rect 435 -675 475 -670
rect 435 -680 440 -675
rect 360 -700 440 -680
rect 360 -705 365 -700
rect 325 -710 365 -705
rect 435 -705 440 -700
rect 470 -680 475 -675
rect 545 -675 585 -670
rect 545 -680 550 -675
rect 470 -700 550 -680
rect 470 -705 475 -700
rect 435 -710 475 -705
rect 545 -705 550 -700
rect 580 -680 585 -675
rect 655 -675 695 -670
rect 655 -680 660 -675
rect 580 -700 660 -680
rect 580 -705 585 -700
rect 545 -710 585 -705
rect 655 -705 660 -700
rect 690 -680 695 -675
rect 765 -675 805 -670
rect 765 -680 770 -675
rect 690 -700 770 -680
rect 690 -705 695 -700
rect 655 -710 695 -705
rect 765 -705 770 -700
rect 800 -680 805 -675
rect 875 -675 915 -670
rect 875 -680 880 -675
rect 800 -700 880 -680
rect 800 -705 805 -700
rect 765 -710 805 -705
rect 875 -705 880 -700
rect 910 -680 915 -675
rect 985 -675 1025 -670
rect 985 -680 990 -675
rect 910 -700 990 -680
rect 910 -705 915 -700
rect 875 -710 915 -705
rect 985 -705 990 -700
rect 1020 -680 1025 -675
rect 1095 -675 1135 -670
rect 1095 -680 1100 -675
rect 1020 -700 1100 -680
rect 1020 -705 1025 -700
rect 985 -710 1025 -705
rect 1095 -705 1100 -700
rect 1130 -680 1135 -675
rect 1205 -675 1245 -670
rect 1205 -680 1210 -675
rect 1130 -700 1210 -680
rect 1130 -705 1135 -700
rect 1095 -710 1135 -705
rect 1205 -705 1210 -700
rect 1240 -680 1245 -675
rect 1315 -675 1355 -670
rect 1315 -680 1320 -675
rect 1240 -700 1320 -680
rect 1240 -705 1245 -700
rect 1205 -710 1245 -705
rect 1315 -705 1320 -700
rect 1350 -680 1355 -675
rect 1425 -675 1465 -670
rect 1425 -680 1430 -675
rect 1350 -700 1430 -680
rect 1350 -705 1355 -700
rect 1315 -710 1355 -705
rect 1425 -705 1430 -700
rect 1460 -680 1465 -675
rect 1850 -675 1890 -670
rect 1850 -680 1855 -675
rect 1460 -700 1855 -680
rect 1460 -705 1465 -700
rect 1425 -710 1465 -705
rect 1850 -705 1855 -700
rect 1885 -705 1890 -675
rect 1850 -710 1890 -705
rect 75 -725 115 -720
rect 75 -755 80 -725
rect 110 -730 115 -725
rect 110 -735 1050 -730
rect 110 -750 1015 -735
rect 110 -755 115 -750
rect 75 -760 115 -755
rect 1010 -765 1015 -750
rect 1045 -765 1050 -735
rect -110 -770 -70 -765
rect -110 -800 -105 -770
rect -75 -775 -70 -770
rect 710 -770 750 -765
rect 710 -775 715 -770
rect -75 -795 715 -775
rect -75 -800 -70 -795
rect -110 -805 -70 -800
rect 710 -800 715 -795
rect 745 -775 750 -770
rect 825 -770 865 -765
rect 825 -775 830 -770
rect 745 -795 830 -775
rect 745 -800 750 -795
rect 710 -805 750 -800
rect 825 -800 830 -795
rect 860 -775 865 -770
rect 950 -770 990 -765
rect 1010 -770 1050 -765
rect 950 -775 955 -770
rect 860 -795 955 -775
rect 860 -800 865 -795
rect 825 -805 865 -800
rect 950 -800 955 -795
rect 985 -800 990 -770
rect 950 -805 990 -800
rect -1025 -1075 -985 -1070
rect -1025 -1105 -1020 -1075
rect -990 -1080 -985 -1075
rect -825 -1075 -785 -1070
rect -825 -1080 -820 -1075
rect -990 -1100 -820 -1080
rect -990 -1105 -985 -1100
rect -1025 -1110 -985 -1105
rect -825 -1105 -820 -1100
rect -790 -1080 -785 -1075
rect -625 -1075 -585 -1070
rect -625 -1080 -620 -1075
rect -790 -1100 -620 -1080
rect -790 -1105 -785 -1100
rect -825 -1110 -785 -1105
rect -625 -1105 -620 -1100
rect -590 -1080 -585 -1075
rect -425 -1075 -385 -1070
rect -425 -1080 -420 -1075
rect -590 -1100 -420 -1080
rect -590 -1105 -585 -1100
rect -625 -1110 -585 -1105
rect -425 -1105 -420 -1100
rect -390 -1080 -385 -1075
rect -200 -1075 -160 -1070
rect -200 -1080 -195 -1075
rect -390 -1100 -195 -1080
rect -390 -1105 -385 -1100
rect -425 -1110 -385 -1105
rect -200 -1105 -195 -1100
rect -165 -1080 -160 -1075
rect 825 -1075 865 -1070
rect 825 -1080 830 -1075
rect -165 -1100 830 -1080
rect -165 -1105 -160 -1100
rect -200 -1110 -160 -1105
rect 825 -1105 830 -1100
rect 860 -1080 865 -1075
rect 1850 -1075 1890 -1070
rect 1850 -1080 1855 -1075
rect 860 -1100 1855 -1080
rect 860 -1105 865 -1100
rect 825 -1110 865 -1105
rect 1850 -1105 1855 -1100
rect 1885 -1080 1890 -1075
rect 2075 -1075 2115 -1070
rect 2075 -1080 2080 -1075
rect 1885 -1100 2080 -1080
rect 1885 -1105 1890 -1100
rect 1850 -1110 1890 -1105
rect 2075 -1105 2080 -1100
rect 2110 -1080 2115 -1075
rect 2275 -1075 2315 -1070
rect 2275 -1080 2280 -1075
rect 2110 -1100 2280 -1080
rect 2110 -1105 2115 -1100
rect 2075 -1110 2115 -1105
rect 2275 -1105 2280 -1100
rect 2310 -1080 2315 -1075
rect 2475 -1075 2515 -1070
rect 2475 -1080 2480 -1075
rect 2310 -1100 2480 -1080
rect 2310 -1105 2315 -1100
rect 2275 -1110 2315 -1105
rect 2475 -1105 2480 -1100
rect 2510 -1080 2515 -1075
rect 2675 -1075 2715 -1070
rect 2675 -1080 2680 -1075
rect 2510 -1100 2680 -1080
rect 2510 -1105 2515 -1100
rect 2475 -1110 2515 -1105
rect 2675 -1105 2680 -1100
rect 2710 -1105 2715 -1075
rect 2675 -1110 2715 -1105
rect 825 -2425 865 -2420
rect 825 -2455 830 -2425
rect 860 -2455 865 -2425
rect 825 -2460 865 -2455
<< via2 >>
rect 830 4245 860 4275
rect -1445 1510 -1415 1540
rect 3105 1460 3135 1490
rect -1535 320 -1505 350
rect 3195 320 3225 350
rect 830 -2455 860 -2425
<< metal3 >>
rect 820 4280 870 4285
rect 820 4240 825 4280
rect 865 4240 870 4280
rect 820 4235 870 4240
rect -3295 3860 -3065 3945
rect -2945 3860 -2715 3945
rect -2595 3860 -2365 3945
rect -3295 3810 -2365 3860
rect -3295 3715 -3065 3810
rect -2945 3715 -2715 3810
rect -2595 3715 -2365 3810
rect -2245 3715 -2015 3945
rect -1895 3715 -1665 3945
rect -1545 3715 -1315 3945
rect -1195 3715 -965 3945
rect -845 3715 -615 3945
rect -495 3715 -265 3945
rect -145 3715 85 3945
rect 205 3715 435 3945
rect 555 3715 785 3945
rect 905 3715 1135 3945
rect 1255 3715 1485 3945
rect 1605 3715 1835 3945
rect 1955 3715 2185 3945
rect 2305 3715 2535 3945
rect 2655 3715 2885 3945
rect 3005 3715 3235 3945
rect 3355 3715 3585 3945
rect 3705 3715 3935 3945
rect 4055 3860 4285 3945
rect 4405 3860 4635 3945
rect 4755 3860 4985 3945
rect 4055 3810 4985 3860
rect 4055 3715 4285 3810
rect 4405 3715 4635 3810
rect 4755 3715 4985 3810
rect -2505 3595 -2455 3715
rect -2155 3595 -2105 3715
rect -1805 3595 -1755 3715
rect -1455 3595 -1405 3715
rect -1105 3595 -1055 3715
rect -755 3595 -705 3715
rect -405 3595 -355 3715
rect -55 3595 -5 3715
rect 295 3595 345 3715
rect 645 3595 695 3715
rect 995 3595 1045 3715
rect 1345 3595 1395 3715
rect 1695 3595 1745 3715
rect 2045 3595 2095 3715
rect 2395 3595 2445 3715
rect 2745 3595 2795 3715
rect 3095 3595 3145 3715
rect 3445 3595 3495 3715
rect 3795 3595 3845 3715
rect 4145 3595 4195 3715
rect -3295 3510 -3065 3595
rect -2945 3510 -2715 3595
rect -2595 3510 -2365 3595
rect -2245 3510 -2015 3595
rect -1895 3510 -1665 3595
rect -1545 3510 -1315 3595
rect -1195 3510 -965 3595
rect -845 3510 -615 3595
rect -495 3510 -265 3595
rect -145 3510 85 3595
rect 205 3510 435 3595
rect 555 3510 785 3595
rect -3295 3460 785 3510
rect -3295 3365 -3065 3460
rect -2945 3365 -2715 3460
rect -2595 3365 -2365 3460
rect -2245 3365 -2015 3460
rect -1895 3365 -1665 3460
rect -1545 3365 -1315 3460
rect -1195 3365 -965 3460
rect -845 3365 -615 3460
rect -495 3365 -265 3460
rect -145 3365 85 3460
rect 205 3365 435 3460
rect 555 3365 785 3460
rect 905 3510 1135 3595
rect 1255 3510 1485 3595
rect 1605 3510 1835 3595
rect 1955 3510 2185 3595
rect 2305 3510 2535 3595
rect 2655 3510 2885 3595
rect 3005 3510 3235 3595
rect 3355 3510 3585 3595
rect 3705 3510 3935 3595
rect 4055 3510 4285 3595
rect 4405 3510 4635 3595
rect 4755 3510 4985 3595
rect 905 3460 4985 3510
rect 905 3365 1135 3460
rect 1255 3365 1485 3460
rect 1605 3365 1835 3460
rect 1955 3365 2185 3460
rect 2305 3365 2535 3460
rect 2655 3365 2885 3460
rect 3005 3365 3235 3460
rect 3355 3365 3585 3460
rect 3705 3365 3935 3460
rect 4055 3365 4285 3460
rect 4405 3365 4635 3460
rect 4755 3365 4985 3460
rect -2505 3245 -2455 3365
rect -1805 3245 -1755 3365
rect -1455 3245 -1405 3365
rect -1105 3245 -1055 3365
rect -755 3245 -705 3365
rect -405 3245 -355 3365
rect -55 3245 -5 3365
rect 295 3245 345 3365
rect 645 3245 695 3365
rect 995 3245 1045 3365
rect 1345 3245 1395 3365
rect 1695 3245 1745 3365
rect 2045 3245 2095 3365
rect 2395 3245 2445 3365
rect 2745 3245 2795 3365
rect 3095 3245 3145 3365
rect 3445 3245 3495 3365
rect 4145 3245 4195 3365
rect -3295 3160 -3065 3245
rect -2945 3160 -2715 3245
rect -2595 3160 -2365 3245
rect -2245 3160 -2015 3245
rect -3295 3110 -2015 3160
rect -3295 3015 -3065 3110
rect -2945 3015 -2715 3110
rect -2595 3015 -2365 3110
rect -2245 3015 -2015 3110
rect -1895 3015 -1665 3245
rect -1545 3015 -1315 3245
rect -1195 3015 -965 3245
rect -845 3015 -615 3245
rect -495 3015 -265 3245
rect -145 3015 85 3245
rect 205 3015 435 3245
rect 555 3015 785 3245
rect 905 3015 1135 3245
rect 1255 3015 1485 3245
rect 1605 3015 1835 3245
rect 1955 3015 2185 3245
rect 2305 3015 2535 3245
rect 2655 3015 2885 3245
rect 3005 3015 3235 3245
rect 3355 3015 3585 3245
rect 3705 3160 3935 3245
rect 4055 3160 4285 3245
rect 4405 3160 4635 3245
rect 4755 3160 4985 3245
rect 3705 3110 4985 3160
rect 3705 3015 3935 3110
rect 4055 3015 4285 3110
rect 4405 3015 4635 3110
rect 4755 3015 4985 3110
rect -2505 2895 -2455 3015
rect -1805 2895 -1755 3015
rect -1455 2895 -1405 3015
rect -1105 2895 -1055 3015
rect -755 2895 -705 3015
rect 2395 2895 2445 3015
rect 2745 2895 2795 3015
rect 3095 2895 3145 3015
rect 3445 2895 3495 3015
rect 4145 2895 4195 3015
rect -3295 2810 -3065 2895
rect -2945 2810 -2715 2895
rect -2595 2810 -2365 2895
rect -2245 2810 -2015 2895
rect -3295 2760 -2015 2810
rect -3295 2665 -3065 2760
rect -2945 2665 -2715 2760
rect -2595 2665 -2365 2760
rect -2245 2665 -2015 2760
rect -1895 2665 -1665 2895
rect -1545 2665 -1315 2895
rect -1195 2665 -965 2895
rect -845 2665 -615 2895
rect 2305 2665 2535 2895
rect 2655 2665 2885 2895
rect 3005 2665 3235 2895
rect 3355 2665 3585 2895
rect 3705 2810 3935 2895
rect 4055 2810 4285 2895
rect 4405 2810 4635 2895
rect 4755 2810 4985 2895
rect 3705 2760 4985 2810
rect 3705 2665 3935 2760
rect 4055 2665 4285 2760
rect 4405 2665 4635 2760
rect 4755 2665 4985 2760
rect -2505 2545 -2455 2665
rect -1455 2545 -1405 2665
rect -1105 2545 -1055 2665
rect -755 2545 -705 2665
rect 2395 2545 2445 2665
rect 2745 2545 2795 2665
rect 3095 2545 3145 2665
rect 4145 2545 4195 2665
rect -3295 2460 -3065 2545
rect -2945 2460 -2715 2545
rect -2595 2460 -2365 2545
rect -2245 2460 -2015 2545
rect -1895 2460 -1665 2545
rect -3295 2410 -1665 2460
rect -3295 2315 -3065 2410
rect -2945 2315 -2715 2410
rect -2595 2315 -2365 2410
rect -2245 2315 -2015 2410
rect -1895 2315 -1665 2410
rect -1545 2315 -1315 2545
rect -1195 2315 -965 2545
rect -845 2315 -615 2545
rect 2305 2315 2535 2545
rect 2655 2315 2885 2545
rect 3005 2315 3235 2545
rect 3355 2460 3585 2545
rect 3705 2460 3935 2545
rect 4055 2460 4285 2545
rect 4405 2460 4635 2545
rect 4755 2460 4985 2545
rect 3355 2410 4985 2460
rect 3355 2315 3585 2410
rect 3705 2315 3935 2410
rect 4055 2315 4285 2410
rect 4405 2315 4635 2410
rect 4755 2315 4985 2410
rect -2505 2195 -2455 2315
rect -3295 2110 -3065 2195
rect -2945 2110 -2715 2195
rect -2595 2110 -2365 2195
rect -2245 2110 -2015 2195
rect -1895 2110 -1665 2195
rect -3295 2060 -1665 2110
rect -3295 1965 -3065 2060
rect -2945 1965 -2715 2060
rect -2595 1965 -2365 2060
rect -2245 1965 -2015 2060
rect -1895 1965 -1665 2060
rect -2505 1845 -2455 1965
rect -3295 1760 -3065 1845
rect -2945 1760 -2715 1845
rect -2595 1760 -2365 1845
rect -2245 1760 -2015 1845
rect -1895 1760 -1665 1845
rect -3295 1710 -1665 1760
rect -3295 1615 -3065 1710
rect -2945 1615 -2715 1710
rect -2595 1615 -2365 1710
rect -2245 1615 -2015 1710
rect -1895 1615 -1665 1710
rect -2505 1495 -2455 1615
rect -1450 1540 -1410 2315
rect -1450 1510 -1445 1540
rect -1415 1510 -1410 1540
rect -1450 1505 -1410 1510
rect -3295 1410 -3065 1495
rect -2945 1410 -2715 1495
rect -2595 1410 -2365 1495
rect -2245 1410 -2015 1495
rect -1895 1410 -1665 1495
rect 3100 1490 3140 2315
rect 4145 2195 4195 2315
rect 3355 2110 3585 2195
rect 3705 2110 3935 2195
rect 4055 2110 4285 2195
rect 4405 2110 4635 2195
rect 4755 2110 4985 2195
rect 3355 2060 4985 2110
rect 3355 1965 3585 2060
rect 3705 1965 3935 2060
rect 4055 1965 4285 2060
rect 4405 1965 4635 2060
rect 4755 1965 4985 2060
rect 4145 1845 4195 1965
rect 3355 1760 3585 1845
rect 3705 1760 3935 1845
rect 4055 1760 4285 1845
rect 4405 1760 4635 1845
rect 4755 1760 4985 1845
rect 3355 1710 4985 1760
rect 3355 1615 3585 1710
rect 3705 1615 3935 1710
rect 4055 1615 4285 1710
rect 4405 1615 4635 1710
rect 4755 1615 4985 1710
rect 4145 1495 4195 1615
rect 3100 1460 3105 1490
rect 3135 1460 3140 1490
rect 3100 1455 3140 1460
rect -3295 1360 -1665 1410
rect -3295 1265 -3065 1360
rect -2945 1265 -2715 1360
rect -2595 1265 -2365 1360
rect -2245 1265 -2015 1360
rect -1895 1265 -1665 1360
rect 3355 1410 3585 1495
rect 3705 1410 3935 1495
rect 4055 1410 4285 1495
rect 4405 1410 4635 1495
rect 4755 1410 4985 1495
rect 3355 1360 4985 1410
rect 3355 1265 3585 1360
rect 3705 1265 3935 1360
rect 4055 1265 4285 1360
rect 4405 1265 4635 1360
rect 4755 1265 4985 1360
rect -2505 1145 -2455 1265
rect 4145 1145 4195 1265
rect -3295 1060 -3065 1145
rect -2945 1060 -2715 1145
rect -2595 1060 -2365 1145
rect -2245 1060 -2015 1145
rect -1895 1060 -1665 1145
rect -3295 1010 -1665 1060
rect -3295 915 -3065 1010
rect -2945 915 -2715 1010
rect -2595 915 -2365 1010
rect -2245 915 -2015 1010
rect -1895 915 -1665 1010
rect 3355 1060 3585 1145
rect 3705 1060 3935 1145
rect 4055 1060 4285 1145
rect 4405 1060 4635 1145
rect 4755 1060 4985 1145
rect 3355 1010 4985 1060
rect 3355 915 3585 1010
rect 3705 915 3935 1010
rect 4055 915 4285 1010
rect 4405 915 4635 1010
rect 4755 915 4985 1010
rect -2505 795 -2455 915
rect 4145 795 4195 915
rect -3295 710 -3065 795
rect -2945 710 -2715 795
rect -2595 710 -2365 795
rect -2245 710 -2015 795
rect -1895 710 -1665 795
rect -3295 660 -1665 710
rect -3295 565 -3065 660
rect -2945 565 -2715 660
rect -2595 565 -2365 660
rect -2245 565 -2015 660
rect -1895 565 -1665 660
rect 3355 710 3585 795
rect 3705 710 3935 795
rect 4055 710 4285 795
rect 4405 710 4635 795
rect 4755 710 4985 795
rect 3355 660 4985 710
rect 3355 565 3585 660
rect 3705 565 3935 660
rect 4055 565 4285 660
rect 4405 565 4635 660
rect 4755 565 4985 660
rect -2505 445 -2455 565
rect 4145 445 4195 565
rect -3295 360 -3065 445
rect -2945 360 -2715 445
rect -2595 360 -2365 445
rect -2245 360 -2015 445
rect -1895 360 -1665 445
rect 3355 360 3585 445
rect 3705 360 3935 445
rect 4055 360 4285 445
rect 4405 360 4635 445
rect 4755 360 4985 445
rect -3295 310 -1665 360
rect -1545 355 -1495 360
rect -1545 315 -1540 355
rect -1500 315 -1495 355
rect -1545 310 -1495 315
rect 3185 355 3235 360
rect 3185 315 3190 355
rect 3230 315 3235 355
rect 3185 310 3235 315
rect 3355 310 4985 360
rect -3295 215 -3065 310
rect -2945 215 -2715 310
rect -2595 215 -2365 310
rect -2245 215 -2015 310
rect -1895 215 -1665 310
rect 3355 215 3585 310
rect 3705 215 3935 310
rect 4055 215 4285 310
rect 4405 215 4635 310
rect 4755 215 4985 310
rect -2505 95 -2455 215
rect 4145 95 4195 215
rect -3295 10 -3065 95
rect -2945 10 -2715 95
rect -2595 10 -2365 95
rect -2245 10 -2015 95
rect -1895 10 -1665 95
rect -3295 -40 -1665 10
rect -3295 -135 -3065 -40
rect -2945 -135 -2715 -40
rect -2595 -135 -2365 -40
rect -2245 -135 -2015 -40
rect -1895 -135 -1665 -40
rect 3355 10 3585 95
rect 3705 10 3935 95
rect 4055 10 4285 95
rect 4405 10 4635 95
rect 4755 10 4985 95
rect 3355 -40 4985 10
rect 3355 -135 3585 -40
rect 3705 -135 3935 -40
rect 4055 -135 4285 -40
rect 4405 -135 4635 -40
rect 4755 -135 4985 -40
rect -2505 -255 -2455 -135
rect 4145 -255 4195 -135
rect -3295 -340 -3065 -255
rect -2945 -340 -2715 -255
rect -2595 -340 -2365 -255
rect -2245 -340 -2015 -255
rect -1895 -340 -1665 -255
rect -3295 -390 -1665 -340
rect -3295 -485 -3065 -390
rect -2945 -485 -2715 -390
rect -2595 -485 -2365 -390
rect -2245 -485 -2015 -390
rect -1895 -485 -1665 -390
rect 3355 -340 3585 -255
rect 3705 -340 3935 -255
rect 4055 -340 4285 -255
rect 4405 -340 4635 -255
rect 4755 -340 4985 -255
rect 3355 -390 4985 -340
rect 3355 -485 3585 -390
rect 3705 -485 3935 -390
rect 4055 -485 4285 -390
rect 4405 -485 4635 -390
rect 4755 -485 4985 -390
rect -2505 -605 -2455 -485
rect 4145 -605 4195 -485
rect -3295 -690 -3065 -605
rect -2945 -690 -2715 -605
rect -2595 -690 -2365 -605
rect -2245 -690 -2015 -605
rect -1895 -690 -1665 -605
rect -3295 -740 -1665 -690
rect -3295 -835 -3065 -740
rect -2945 -835 -2715 -740
rect -2595 -835 -2365 -740
rect -2245 -835 -2015 -740
rect -1895 -835 -1665 -740
rect 3355 -690 3585 -605
rect 3705 -690 3935 -605
rect 4055 -690 4285 -605
rect 4405 -690 4635 -605
rect 4755 -690 4985 -605
rect 3355 -740 4985 -690
rect 3355 -835 3585 -740
rect 3705 -835 3935 -740
rect 4055 -835 4285 -740
rect 4405 -835 4635 -740
rect 4755 -835 4985 -740
rect -2505 -955 -2455 -835
rect 4145 -955 4195 -835
rect -3295 -1040 -3065 -955
rect -2945 -1040 -2715 -955
rect -2595 -1040 -2365 -955
rect -2245 -1040 -2015 -955
rect -1895 -1040 -1665 -955
rect -3295 -1090 -1665 -1040
rect -3295 -1185 -3065 -1090
rect -2945 -1185 -2715 -1090
rect -2595 -1185 -2365 -1090
rect -2245 -1185 -2015 -1090
rect -1895 -1185 -1665 -1090
rect 3355 -1040 3585 -955
rect 3705 -1040 3935 -955
rect 4055 -1040 4285 -955
rect 4405 -1040 4635 -955
rect 4755 -1040 4985 -955
rect 3355 -1090 4985 -1040
rect 3355 -1185 3585 -1090
rect 3705 -1185 3935 -1090
rect 4055 -1185 4285 -1090
rect 4405 -1185 4635 -1090
rect 4755 -1185 4985 -1090
rect -2505 -1305 -2455 -1185
rect 4145 -1305 4195 -1185
rect -3295 -1390 -3065 -1305
rect -2945 -1390 -2715 -1305
rect -2595 -1390 -2365 -1305
rect -2245 -1390 -2015 -1305
rect -1895 -1390 -1665 -1305
rect -3295 -1440 -1665 -1390
rect -3295 -1535 -3065 -1440
rect -2945 -1535 -2715 -1440
rect -2595 -1535 -2365 -1440
rect -2245 -1535 -2015 -1440
rect -1895 -1535 -1665 -1440
rect -1545 -1535 -1315 -1305
rect -1195 -1535 -965 -1305
rect -845 -1535 -615 -1305
rect -495 -1535 -265 -1305
rect -145 -1535 85 -1305
rect 205 -1535 435 -1305
rect 555 -1535 785 -1305
rect 905 -1535 1135 -1305
rect 1255 -1535 1485 -1305
rect 1605 -1535 1835 -1305
rect 1955 -1535 2185 -1305
rect 2305 -1535 2535 -1305
rect 2655 -1535 2885 -1305
rect 3005 -1535 3235 -1305
rect 3355 -1390 3585 -1305
rect 3705 -1390 3935 -1305
rect 4055 -1390 4285 -1305
rect 4405 -1390 4635 -1305
rect 4755 -1390 4985 -1305
rect 3355 -1440 4985 -1390
rect 3355 -1535 3585 -1440
rect 3705 -1535 3935 -1440
rect 4055 -1535 4285 -1440
rect 4405 -1535 4635 -1440
rect 4755 -1535 4985 -1440
rect -2505 -1655 -2455 -1535
rect -1455 -1655 -1405 -1535
rect -1105 -1655 -1055 -1535
rect -755 -1655 -705 -1535
rect -405 -1655 -355 -1535
rect -55 -1655 -5 -1535
rect 295 -1655 345 -1535
rect 645 -1655 695 -1535
rect 995 -1655 1045 -1535
rect 1345 -1655 1395 -1535
rect 1695 -1655 1745 -1535
rect 2045 -1655 2095 -1535
rect 2395 -1655 2445 -1535
rect 2745 -1655 2795 -1535
rect 3095 -1655 3145 -1535
rect 4145 -1655 4195 -1535
rect -3295 -1740 -3065 -1655
rect -2945 -1740 -2715 -1655
rect -2595 -1740 -2365 -1655
rect -2245 -1740 -2015 -1655
rect -1895 -1740 -1665 -1655
rect -1545 -1740 -1315 -1655
rect -1195 -1740 -965 -1655
rect -845 -1740 -615 -1655
rect -495 -1740 -265 -1655
rect -145 -1740 85 -1655
rect 205 -1740 435 -1655
rect 555 -1740 785 -1655
rect -3295 -1790 785 -1740
rect -3295 -1885 -3065 -1790
rect -2945 -1885 -2715 -1790
rect -2595 -1885 -2365 -1790
rect -2245 -1885 -2015 -1790
rect -1895 -1885 -1665 -1790
rect -1545 -1885 -1315 -1790
rect -1195 -1885 -965 -1790
rect -845 -1885 -615 -1790
rect -495 -1885 -265 -1790
rect -145 -1885 85 -1790
rect 205 -1885 435 -1790
rect 555 -1885 785 -1790
rect 905 -1740 1135 -1655
rect 1255 -1740 1485 -1655
rect 1605 -1740 1835 -1655
rect 1955 -1740 2185 -1655
rect 2305 -1740 2535 -1655
rect 2655 -1740 2885 -1655
rect 3005 -1740 3235 -1655
rect 3355 -1740 3585 -1655
rect 3705 -1740 3935 -1655
rect 4055 -1740 4285 -1655
rect 4405 -1740 4635 -1655
rect 4755 -1740 4985 -1655
rect 905 -1790 4985 -1740
rect 905 -1885 1135 -1790
rect 1255 -1885 1485 -1790
rect 1605 -1885 1835 -1790
rect 1955 -1885 2185 -1790
rect 2305 -1885 2535 -1790
rect 2655 -1885 2885 -1790
rect 3005 -1885 3235 -1790
rect 3355 -1885 3585 -1790
rect 3705 -1885 3935 -1790
rect 4055 -1885 4285 -1790
rect 4405 -1885 4635 -1790
rect 4755 -1885 4985 -1790
rect -2505 -2005 -2455 -1885
rect -2155 -2005 -2105 -1885
rect -1805 -2005 -1755 -1885
rect -1455 -2005 -1405 -1885
rect -1105 -2005 -1055 -1885
rect -755 -2005 -705 -1885
rect -405 -2005 -355 -1885
rect -55 -2005 -5 -1885
rect 295 -2005 345 -1885
rect 645 -2005 695 -1885
rect 995 -2005 1045 -1885
rect 1345 -2005 1395 -1885
rect 1695 -2005 1745 -1885
rect 2045 -2005 2095 -1885
rect 2395 -2005 2445 -1885
rect 2745 -2005 2795 -1885
rect 3095 -2005 3145 -1885
rect 3445 -2005 3495 -1885
rect 3795 -2005 3845 -1885
rect 4145 -2005 4195 -1885
rect -3295 -2090 -3065 -2005
rect -2945 -2090 -2715 -2005
rect -2595 -2090 -2365 -2005
rect -3295 -2140 -2365 -2090
rect -3295 -2235 -3065 -2140
rect -2945 -2235 -2715 -2140
rect -2595 -2235 -2365 -2140
rect -2245 -2235 -2015 -2005
rect -1895 -2235 -1665 -2005
rect -1545 -2235 -1315 -2005
rect -1195 -2235 -965 -2005
rect -845 -2235 -615 -2005
rect -495 -2235 -265 -2005
rect -145 -2235 85 -2005
rect 205 -2235 435 -2005
rect 555 -2235 785 -2005
rect 905 -2235 1135 -2005
rect 1255 -2235 1485 -2005
rect 1605 -2235 1835 -2005
rect 1955 -2235 2185 -2005
rect 2305 -2235 2535 -2005
rect 2655 -2235 2885 -2005
rect 3005 -2235 3235 -2005
rect 3355 -2235 3585 -2005
rect 3705 -2235 3935 -2005
rect 4055 -2090 4285 -2005
rect 4405 -2090 4635 -2005
rect 4755 -2090 4985 -2005
rect 4055 -2140 4985 -2090
rect 4055 -2235 4285 -2140
rect 4405 -2235 4635 -2140
rect 4755 -2235 4985 -2140
rect 820 -2420 870 -2415
rect 820 -2460 825 -2420
rect 865 -2460 870 -2420
rect 820 -2465 870 -2460
<< via3 >>
rect 825 4275 865 4280
rect 825 4245 830 4275
rect 830 4245 860 4275
rect 860 4245 865 4275
rect 825 4240 865 4245
rect -1540 350 -1500 355
rect -1540 320 -1535 350
rect -1535 320 -1505 350
rect -1505 320 -1500 350
rect -1540 315 -1500 320
rect 3190 350 3230 355
rect 3190 320 3195 350
rect 3195 320 3225 350
rect 3225 320 3230 350
rect 3190 315 3230 320
rect 825 -2425 865 -2420
rect 825 -2455 830 -2425
rect 830 -2455 860 -2425
rect 860 -2455 865 -2425
rect 825 -2460 865 -2455
<< mimcap >>
rect -3280 3855 -3080 3930
rect -3280 3815 -3200 3855
rect -3160 3815 -3080 3855
rect -3280 3730 -3080 3815
rect -2930 3855 -2730 3930
rect -2930 3815 -2850 3855
rect -2810 3815 -2730 3855
rect -2930 3730 -2730 3815
rect -2580 3855 -2380 3930
rect -2580 3815 -2500 3855
rect -2460 3815 -2380 3855
rect -2580 3730 -2380 3815
rect -2230 3855 -2030 3930
rect -2230 3815 -2150 3855
rect -2110 3815 -2030 3855
rect -2230 3730 -2030 3815
rect -1880 3855 -1680 3930
rect -1880 3815 -1800 3855
rect -1760 3815 -1680 3855
rect -1880 3730 -1680 3815
rect -1530 3855 -1330 3930
rect -1530 3815 -1450 3855
rect -1410 3815 -1330 3855
rect -1530 3730 -1330 3815
rect -1180 3855 -980 3930
rect -1180 3815 -1100 3855
rect -1060 3815 -980 3855
rect -1180 3730 -980 3815
rect -830 3855 -630 3930
rect -830 3815 -750 3855
rect -710 3815 -630 3855
rect -830 3730 -630 3815
rect -480 3855 -280 3930
rect -480 3815 -400 3855
rect -360 3815 -280 3855
rect -480 3730 -280 3815
rect -130 3855 70 3930
rect -130 3815 -50 3855
rect -10 3815 70 3855
rect -130 3730 70 3815
rect 220 3855 420 3930
rect 220 3815 300 3855
rect 340 3815 420 3855
rect 220 3730 420 3815
rect 570 3855 770 3930
rect 570 3815 650 3855
rect 690 3815 770 3855
rect 570 3730 770 3815
rect 920 3855 1120 3930
rect 920 3815 1000 3855
rect 1040 3815 1120 3855
rect 920 3730 1120 3815
rect 1270 3855 1470 3930
rect 1270 3815 1350 3855
rect 1390 3815 1470 3855
rect 1270 3730 1470 3815
rect 1620 3855 1820 3930
rect 1620 3815 1700 3855
rect 1740 3815 1820 3855
rect 1620 3730 1820 3815
rect 1970 3855 2170 3930
rect 1970 3815 2050 3855
rect 2090 3815 2170 3855
rect 1970 3730 2170 3815
rect 2320 3855 2520 3930
rect 2320 3815 2400 3855
rect 2440 3815 2520 3855
rect 2320 3730 2520 3815
rect 2670 3855 2870 3930
rect 2670 3815 2750 3855
rect 2790 3815 2870 3855
rect 2670 3730 2870 3815
rect 3020 3855 3220 3930
rect 3020 3815 3100 3855
rect 3140 3815 3220 3855
rect 3020 3730 3220 3815
rect 3370 3855 3570 3930
rect 3370 3815 3450 3855
rect 3490 3815 3570 3855
rect 3370 3730 3570 3815
rect 3720 3855 3920 3930
rect 3720 3815 3800 3855
rect 3840 3815 3920 3855
rect 3720 3730 3920 3815
rect 4070 3855 4270 3930
rect 4070 3815 4150 3855
rect 4190 3815 4270 3855
rect 4070 3730 4270 3815
rect 4420 3855 4620 3930
rect 4420 3815 4500 3855
rect 4540 3815 4620 3855
rect 4420 3730 4620 3815
rect 4770 3855 4970 3930
rect 4770 3815 4850 3855
rect 4890 3815 4970 3855
rect 4770 3730 4970 3815
rect -3280 3505 -3080 3580
rect -3280 3465 -3200 3505
rect -3160 3465 -3080 3505
rect -3280 3380 -3080 3465
rect -2930 3505 -2730 3580
rect -2930 3465 -2850 3505
rect -2810 3465 -2730 3505
rect -2930 3380 -2730 3465
rect -2580 3505 -2380 3580
rect -2580 3465 -2500 3505
rect -2460 3465 -2380 3505
rect -2580 3380 -2380 3465
rect -2230 3505 -2030 3580
rect -2230 3465 -2150 3505
rect -2110 3465 -2030 3505
rect -2230 3380 -2030 3465
rect -1880 3505 -1680 3580
rect -1880 3465 -1800 3505
rect -1760 3465 -1680 3505
rect -1880 3380 -1680 3465
rect -1530 3505 -1330 3580
rect -1530 3465 -1450 3505
rect -1410 3465 -1330 3505
rect -1530 3380 -1330 3465
rect -1180 3505 -980 3580
rect -1180 3465 -1100 3505
rect -1060 3465 -980 3505
rect -1180 3380 -980 3465
rect -830 3505 -630 3580
rect -830 3465 -750 3505
rect -710 3465 -630 3505
rect -830 3380 -630 3465
rect -480 3505 -280 3580
rect -480 3465 -400 3505
rect -360 3465 -280 3505
rect -480 3380 -280 3465
rect -130 3505 70 3580
rect -130 3465 -50 3505
rect -10 3465 70 3505
rect -130 3380 70 3465
rect 220 3505 420 3580
rect 220 3465 300 3505
rect 340 3465 420 3505
rect 220 3380 420 3465
rect 570 3505 770 3580
rect 570 3465 650 3505
rect 690 3465 770 3505
rect 570 3380 770 3465
rect 920 3505 1120 3580
rect 920 3465 1000 3505
rect 1040 3465 1120 3505
rect 920 3380 1120 3465
rect 1270 3505 1470 3580
rect 1270 3465 1350 3505
rect 1390 3465 1470 3505
rect 1270 3380 1470 3465
rect 1620 3505 1820 3580
rect 1620 3465 1700 3505
rect 1740 3465 1820 3505
rect 1620 3380 1820 3465
rect 1970 3505 2170 3580
rect 1970 3465 2050 3505
rect 2090 3465 2170 3505
rect 1970 3380 2170 3465
rect 2320 3505 2520 3580
rect 2320 3465 2400 3505
rect 2440 3465 2520 3505
rect 2320 3380 2520 3465
rect 2670 3505 2870 3580
rect 2670 3465 2750 3505
rect 2790 3465 2870 3505
rect 2670 3380 2870 3465
rect 3020 3505 3220 3580
rect 3020 3465 3100 3505
rect 3140 3465 3220 3505
rect 3020 3380 3220 3465
rect 3370 3505 3570 3580
rect 3370 3465 3450 3505
rect 3490 3465 3570 3505
rect 3370 3380 3570 3465
rect 3720 3505 3920 3580
rect 3720 3465 3800 3505
rect 3840 3465 3920 3505
rect 3720 3380 3920 3465
rect 4070 3505 4270 3580
rect 4070 3465 4150 3505
rect 4190 3465 4270 3505
rect 4070 3380 4270 3465
rect 4420 3505 4620 3580
rect 4420 3465 4500 3505
rect 4540 3465 4620 3505
rect 4420 3380 4620 3465
rect 4770 3505 4970 3580
rect 4770 3465 4850 3505
rect 4890 3465 4970 3505
rect 4770 3380 4970 3465
rect -3280 3155 -3080 3230
rect -3280 3115 -3200 3155
rect -3160 3115 -3080 3155
rect -3280 3030 -3080 3115
rect -2930 3155 -2730 3230
rect -2930 3115 -2850 3155
rect -2810 3115 -2730 3155
rect -2930 3030 -2730 3115
rect -2580 3155 -2380 3230
rect -2580 3115 -2500 3155
rect -2460 3115 -2380 3155
rect -2580 3030 -2380 3115
rect -2230 3155 -2030 3230
rect -2230 3115 -2150 3155
rect -2110 3115 -2030 3155
rect -2230 3030 -2030 3115
rect -1880 3155 -1680 3230
rect -1880 3115 -1800 3155
rect -1760 3115 -1680 3155
rect -1880 3030 -1680 3115
rect -1530 3155 -1330 3230
rect -1530 3115 -1450 3155
rect -1410 3115 -1330 3155
rect -1530 3030 -1330 3115
rect -1180 3155 -980 3230
rect -1180 3115 -1100 3155
rect -1060 3115 -980 3155
rect -1180 3030 -980 3115
rect -830 3155 -630 3230
rect -830 3115 -750 3155
rect -710 3115 -630 3155
rect -830 3030 -630 3115
rect -480 3155 -280 3230
rect -480 3115 -400 3155
rect -360 3115 -280 3155
rect -480 3030 -280 3115
rect -130 3145 70 3230
rect -130 3105 -50 3145
rect -10 3105 70 3145
rect -130 3030 70 3105
rect 220 3145 420 3230
rect 220 3105 300 3145
rect 340 3105 420 3145
rect 220 3030 420 3105
rect 570 3145 770 3230
rect 570 3105 650 3145
rect 690 3105 770 3145
rect 570 3030 770 3105
rect 920 3145 1120 3230
rect 920 3105 1000 3145
rect 1040 3105 1120 3145
rect 920 3030 1120 3105
rect 1270 3145 1470 3230
rect 1270 3105 1350 3145
rect 1390 3105 1470 3145
rect 1270 3030 1470 3105
rect 1620 3145 1820 3230
rect 1620 3105 1700 3145
rect 1740 3105 1820 3145
rect 1620 3030 1820 3105
rect 1970 3155 2170 3230
rect 1970 3115 2050 3155
rect 2090 3115 2170 3155
rect 1970 3030 2170 3115
rect 2320 3155 2520 3230
rect 2320 3115 2400 3155
rect 2440 3115 2520 3155
rect 2320 3030 2520 3115
rect 2670 3155 2870 3230
rect 2670 3115 2750 3155
rect 2790 3115 2870 3155
rect 2670 3030 2870 3115
rect 3020 3155 3220 3230
rect 3020 3115 3100 3155
rect 3140 3115 3220 3155
rect 3020 3030 3220 3115
rect 3370 3155 3570 3230
rect 3370 3115 3450 3155
rect 3490 3115 3570 3155
rect 3370 3030 3570 3115
rect 3720 3155 3920 3230
rect 3720 3115 3800 3155
rect 3840 3115 3920 3155
rect 3720 3030 3920 3115
rect 4070 3155 4270 3230
rect 4070 3115 4150 3155
rect 4190 3115 4270 3155
rect 4070 3030 4270 3115
rect 4420 3155 4620 3230
rect 4420 3115 4500 3155
rect 4540 3115 4620 3155
rect 4420 3030 4620 3115
rect 4770 3155 4970 3230
rect 4770 3115 4850 3155
rect 4890 3115 4970 3155
rect 4770 3030 4970 3115
rect -3280 2805 -3080 2880
rect -3280 2765 -3200 2805
rect -3160 2765 -3080 2805
rect -3280 2680 -3080 2765
rect -2930 2805 -2730 2880
rect -2930 2765 -2850 2805
rect -2810 2765 -2730 2805
rect -2930 2680 -2730 2765
rect -2580 2805 -2380 2880
rect -2580 2765 -2500 2805
rect -2460 2765 -2380 2805
rect -2580 2680 -2380 2765
rect -2230 2805 -2030 2880
rect -2230 2765 -2150 2805
rect -2110 2765 -2030 2805
rect -2230 2680 -2030 2765
rect -1880 2805 -1680 2880
rect -1880 2765 -1800 2805
rect -1760 2765 -1680 2805
rect -1880 2680 -1680 2765
rect -1530 2805 -1330 2880
rect -1530 2765 -1450 2805
rect -1410 2765 -1330 2805
rect -1530 2680 -1330 2765
rect -1180 2805 -980 2880
rect -1180 2765 -1100 2805
rect -1060 2765 -980 2805
rect -1180 2680 -980 2765
rect -830 2805 -630 2880
rect -830 2765 -750 2805
rect -710 2765 -630 2805
rect -830 2680 -630 2765
rect 2320 2805 2520 2880
rect 2320 2765 2400 2805
rect 2440 2765 2520 2805
rect 2320 2680 2520 2765
rect 2670 2805 2870 2880
rect 2670 2765 2750 2805
rect 2790 2765 2870 2805
rect 2670 2680 2870 2765
rect 3020 2805 3220 2880
rect 3020 2765 3100 2805
rect 3140 2765 3220 2805
rect 3020 2680 3220 2765
rect 3370 2805 3570 2880
rect 3370 2765 3450 2805
rect 3490 2765 3570 2805
rect 3370 2680 3570 2765
rect 3720 2805 3920 2880
rect 3720 2765 3800 2805
rect 3840 2765 3920 2805
rect 3720 2680 3920 2765
rect 4070 2805 4270 2880
rect 4070 2765 4150 2805
rect 4190 2765 4270 2805
rect 4070 2680 4270 2765
rect 4420 2805 4620 2880
rect 4420 2765 4500 2805
rect 4540 2765 4620 2805
rect 4420 2680 4620 2765
rect 4770 2805 4970 2880
rect 4770 2765 4850 2805
rect 4890 2765 4970 2805
rect 4770 2680 4970 2765
rect -3280 2455 -3080 2530
rect -3280 2415 -3200 2455
rect -3160 2415 -3080 2455
rect -3280 2330 -3080 2415
rect -2930 2455 -2730 2530
rect -2930 2415 -2850 2455
rect -2810 2415 -2730 2455
rect -2930 2330 -2730 2415
rect -2580 2455 -2380 2530
rect -2580 2415 -2500 2455
rect -2460 2415 -2380 2455
rect -2580 2330 -2380 2415
rect -2230 2455 -2030 2530
rect -2230 2415 -2150 2455
rect -2110 2415 -2030 2455
rect -2230 2330 -2030 2415
rect -1880 2455 -1680 2530
rect -1880 2415 -1800 2455
rect -1760 2415 -1680 2455
rect -1880 2330 -1680 2415
rect -1530 2455 -1330 2530
rect -1530 2415 -1450 2455
rect -1410 2415 -1330 2455
rect -1530 2330 -1330 2415
rect -1180 2455 -980 2530
rect -1180 2415 -1100 2455
rect -1060 2415 -980 2455
rect -1180 2330 -980 2415
rect -830 2455 -630 2530
rect -830 2415 -750 2455
rect -710 2415 -630 2455
rect -830 2330 -630 2415
rect 2320 2455 2520 2530
rect 2320 2415 2400 2455
rect 2440 2415 2520 2455
rect 2320 2330 2520 2415
rect 2670 2455 2870 2530
rect 2670 2415 2750 2455
rect 2790 2415 2870 2455
rect 2670 2330 2870 2415
rect 3020 2455 3220 2530
rect 3020 2415 3100 2455
rect 3140 2415 3220 2455
rect 3020 2330 3220 2415
rect 3370 2455 3570 2530
rect 3370 2415 3450 2455
rect 3490 2415 3570 2455
rect 3370 2330 3570 2415
rect 3720 2455 3920 2530
rect 3720 2415 3800 2455
rect 3840 2415 3920 2455
rect 3720 2330 3920 2415
rect 4070 2455 4270 2530
rect 4070 2415 4150 2455
rect 4190 2415 4270 2455
rect 4070 2330 4270 2415
rect 4420 2455 4620 2530
rect 4420 2415 4500 2455
rect 4540 2415 4620 2455
rect 4420 2330 4620 2415
rect 4770 2455 4970 2530
rect 4770 2415 4850 2455
rect 4890 2415 4970 2455
rect 4770 2330 4970 2415
rect -3280 2105 -3080 2180
rect -3280 2065 -3200 2105
rect -3160 2065 -3080 2105
rect -3280 1980 -3080 2065
rect -2930 2105 -2730 2180
rect -2930 2065 -2850 2105
rect -2810 2065 -2730 2105
rect -2930 1980 -2730 2065
rect -2580 2105 -2380 2180
rect -2580 2065 -2500 2105
rect -2460 2065 -2380 2105
rect -2580 1980 -2380 2065
rect -2230 2105 -2030 2180
rect -2230 2065 -2150 2105
rect -2110 2065 -2030 2105
rect -2230 1980 -2030 2065
rect -1880 2105 -1680 2180
rect -1880 2065 -1800 2105
rect -1760 2065 -1680 2105
rect -1880 1980 -1680 2065
rect 3370 2105 3570 2180
rect 3370 2065 3450 2105
rect 3490 2065 3570 2105
rect 3370 1980 3570 2065
rect 3720 2105 3920 2180
rect 3720 2065 3800 2105
rect 3840 2065 3920 2105
rect 3720 1980 3920 2065
rect 4070 2105 4270 2180
rect 4070 2065 4150 2105
rect 4190 2065 4270 2105
rect 4070 1980 4270 2065
rect 4420 2105 4620 2180
rect 4420 2065 4500 2105
rect 4540 2065 4620 2105
rect 4420 1980 4620 2065
rect 4770 2105 4970 2180
rect 4770 2065 4850 2105
rect 4890 2065 4970 2105
rect 4770 1980 4970 2065
rect -3280 1755 -3080 1830
rect -3280 1715 -3200 1755
rect -3160 1715 -3080 1755
rect -3280 1630 -3080 1715
rect -2930 1755 -2730 1830
rect -2930 1715 -2850 1755
rect -2810 1715 -2730 1755
rect -2930 1630 -2730 1715
rect -2580 1755 -2380 1830
rect -2580 1715 -2500 1755
rect -2460 1715 -2380 1755
rect -2580 1630 -2380 1715
rect -2230 1755 -2030 1830
rect -2230 1715 -2150 1755
rect -2110 1715 -2030 1755
rect -2230 1630 -2030 1715
rect -1880 1755 -1680 1830
rect -1880 1715 -1800 1755
rect -1760 1715 -1680 1755
rect -1880 1630 -1680 1715
rect 3370 1755 3570 1830
rect 3370 1715 3450 1755
rect 3490 1715 3570 1755
rect 3370 1630 3570 1715
rect 3720 1755 3920 1830
rect 3720 1715 3800 1755
rect 3840 1715 3920 1755
rect 3720 1630 3920 1715
rect 4070 1755 4270 1830
rect 4070 1715 4150 1755
rect 4190 1715 4270 1755
rect 4070 1630 4270 1715
rect 4420 1755 4620 1830
rect 4420 1715 4500 1755
rect 4540 1715 4620 1755
rect 4420 1630 4620 1715
rect 4770 1755 4970 1830
rect 4770 1715 4850 1755
rect 4890 1715 4970 1755
rect 4770 1630 4970 1715
rect -3280 1405 -3080 1480
rect -3280 1365 -3200 1405
rect -3160 1365 -3080 1405
rect -3280 1280 -3080 1365
rect -2930 1405 -2730 1480
rect -2930 1365 -2850 1405
rect -2810 1365 -2730 1405
rect -2930 1280 -2730 1365
rect -2580 1405 -2380 1480
rect -2580 1365 -2500 1405
rect -2460 1365 -2380 1405
rect -2580 1280 -2380 1365
rect -2230 1405 -2030 1480
rect -2230 1365 -2150 1405
rect -2110 1365 -2030 1405
rect -2230 1280 -2030 1365
rect -1880 1405 -1680 1480
rect -1880 1365 -1800 1405
rect -1760 1365 -1680 1405
rect -1880 1280 -1680 1365
rect 3370 1405 3570 1480
rect 3370 1365 3450 1405
rect 3490 1365 3570 1405
rect 3370 1280 3570 1365
rect 3720 1405 3920 1480
rect 3720 1365 3800 1405
rect 3840 1365 3920 1405
rect 3720 1280 3920 1365
rect 4070 1405 4270 1480
rect 4070 1365 4150 1405
rect 4190 1365 4270 1405
rect 4070 1280 4270 1365
rect 4420 1405 4620 1480
rect 4420 1365 4500 1405
rect 4540 1365 4620 1405
rect 4420 1280 4620 1365
rect 4770 1405 4970 1480
rect 4770 1365 4850 1405
rect 4890 1365 4970 1405
rect 4770 1280 4970 1365
rect -3280 1055 -3080 1130
rect -3280 1015 -3200 1055
rect -3160 1015 -3080 1055
rect -3280 930 -3080 1015
rect -2930 1055 -2730 1130
rect -2930 1015 -2850 1055
rect -2810 1015 -2730 1055
rect -2930 930 -2730 1015
rect -2580 1055 -2380 1130
rect -2580 1015 -2500 1055
rect -2460 1015 -2380 1055
rect -2580 930 -2380 1015
rect -2230 1055 -2030 1130
rect -2230 1015 -2150 1055
rect -2110 1015 -2030 1055
rect -2230 930 -2030 1015
rect -1880 1055 -1680 1130
rect -1880 1015 -1800 1055
rect -1760 1015 -1680 1055
rect -1880 930 -1680 1015
rect 3370 1055 3570 1130
rect 3370 1015 3450 1055
rect 3490 1015 3570 1055
rect 3370 930 3570 1015
rect 3720 1055 3920 1130
rect 3720 1015 3800 1055
rect 3840 1015 3920 1055
rect 3720 930 3920 1015
rect 4070 1055 4270 1130
rect 4070 1015 4150 1055
rect 4190 1015 4270 1055
rect 4070 930 4270 1015
rect 4420 1055 4620 1130
rect 4420 1015 4500 1055
rect 4540 1015 4620 1055
rect 4420 930 4620 1015
rect 4770 1055 4970 1130
rect 4770 1015 4850 1055
rect 4890 1015 4970 1055
rect 4770 930 4970 1015
rect -3280 705 -3080 780
rect -3280 665 -3200 705
rect -3160 665 -3080 705
rect -3280 580 -3080 665
rect -2930 705 -2730 780
rect -2930 665 -2850 705
rect -2810 665 -2730 705
rect -2930 580 -2730 665
rect -2580 705 -2380 780
rect -2580 665 -2500 705
rect -2460 665 -2380 705
rect -2580 580 -2380 665
rect -2230 705 -2030 780
rect -2230 665 -2150 705
rect -2110 665 -2030 705
rect -2230 580 -2030 665
rect -1880 705 -1680 780
rect -1880 665 -1800 705
rect -1760 665 -1680 705
rect -1880 580 -1680 665
rect 3370 705 3570 780
rect 3370 665 3450 705
rect 3490 665 3570 705
rect 3370 580 3570 665
rect 3720 705 3920 780
rect 3720 665 3800 705
rect 3840 665 3920 705
rect 3720 580 3920 665
rect 4070 705 4270 780
rect 4070 665 4150 705
rect 4190 665 4270 705
rect 4070 580 4270 665
rect 4420 705 4620 780
rect 4420 665 4500 705
rect 4540 665 4620 705
rect 4420 580 4620 665
rect 4770 705 4970 780
rect 4770 665 4850 705
rect 4890 665 4970 705
rect 4770 580 4970 665
rect -3280 355 -3080 430
rect -3280 315 -3200 355
rect -3160 315 -3080 355
rect -3280 230 -3080 315
rect -2930 355 -2730 430
rect -2930 315 -2850 355
rect -2810 315 -2730 355
rect -2930 230 -2730 315
rect -2580 355 -2380 430
rect -2580 315 -2500 355
rect -2460 315 -2380 355
rect -2580 230 -2380 315
rect -2230 355 -2030 430
rect -2230 315 -2150 355
rect -2110 315 -2030 355
rect -2230 230 -2030 315
rect -1880 355 -1680 430
rect -1880 315 -1800 355
rect -1760 315 -1680 355
rect -1880 230 -1680 315
rect 3370 355 3570 430
rect 3370 315 3450 355
rect 3490 315 3570 355
rect 3370 230 3570 315
rect 3720 355 3920 430
rect 3720 315 3800 355
rect 3840 315 3920 355
rect 3720 230 3920 315
rect 4070 355 4270 430
rect 4070 315 4150 355
rect 4190 315 4270 355
rect 4070 230 4270 315
rect 4420 355 4620 430
rect 4420 315 4500 355
rect 4540 315 4620 355
rect 4420 230 4620 315
rect 4770 355 4970 430
rect 4770 315 4850 355
rect 4890 315 4970 355
rect 4770 230 4970 315
rect -3280 5 -3080 80
rect -3280 -35 -3200 5
rect -3160 -35 -3080 5
rect -3280 -120 -3080 -35
rect -2930 5 -2730 80
rect -2930 -35 -2850 5
rect -2810 -35 -2730 5
rect -2930 -120 -2730 -35
rect -2580 5 -2380 80
rect -2580 -35 -2500 5
rect -2460 -35 -2380 5
rect -2580 -120 -2380 -35
rect -2230 5 -2030 80
rect -2230 -35 -2150 5
rect -2110 -35 -2030 5
rect -2230 -120 -2030 -35
rect -1880 5 -1680 80
rect -1880 -35 -1800 5
rect -1760 -35 -1680 5
rect -1880 -120 -1680 -35
rect 3370 5 3570 80
rect 3370 -35 3450 5
rect 3490 -35 3570 5
rect 3370 -120 3570 -35
rect 3720 5 3920 80
rect 3720 -35 3800 5
rect 3840 -35 3920 5
rect 3720 -120 3920 -35
rect 4070 5 4270 80
rect 4070 -35 4150 5
rect 4190 -35 4270 5
rect 4070 -120 4270 -35
rect 4420 5 4620 80
rect 4420 -35 4500 5
rect 4540 -35 4620 5
rect 4420 -120 4620 -35
rect 4770 5 4970 80
rect 4770 -35 4850 5
rect 4890 -35 4970 5
rect 4770 -120 4970 -35
rect -3280 -345 -3080 -270
rect -3280 -385 -3200 -345
rect -3160 -385 -3080 -345
rect -3280 -470 -3080 -385
rect -2930 -345 -2730 -270
rect -2930 -385 -2850 -345
rect -2810 -385 -2730 -345
rect -2930 -470 -2730 -385
rect -2580 -345 -2380 -270
rect -2580 -385 -2500 -345
rect -2460 -385 -2380 -345
rect -2580 -470 -2380 -385
rect -2230 -345 -2030 -270
rect -2230 -385 -2150 -345
rect -2110 -385 -2030 -345
rect -2230 -470 -2030 -385
rect -1880 -345 -1680 -270
rect -1880 -385 -1800 -345
rect -1760 -385 -1680 -345
rect -1880 -470 -1680 -385
rect 3370 -345 3570 -270
rect 3370 -385 3450 -345
rect 3490 -385 3570 -345
rect 3370 -470 3570 -385
rect 3720 -345 3920 -270
rect 3720 -385 3800 -345
rect 3840 -385 3920 -345
rect 3720 -470 3920 -385
rect 4070 -345 4270 -270
rect 4070 -385 4150 -345
rect 4190 -385 4270 -345
rect 4070 -470 4270 -385
rect 4420 -345 4620 -270
rect 4420 -385 4500 -345
rect 4540 -385 4620 -345
rect 4420 -470 4620 -385
rect 4770 -345 4970 -270
rect 4770 -385 4850 -345
rect 4890 -385 4970 -345
rect 4770 -470 4970 -385
rect -3280 -695 -3080 -620
rect -3280 -735 -3200 -695
rect -3160 -735 -3080 -695
rect -3280 -820 -3080 -735
rect -2930 -695 -2730 -620
rect -2930 -735 -2850 -695
rect -2810 -735 -2730 -695
rect -2930 -820 -2730 -735
rect -2580 -695 -2380 -620
rect -2580 -735 -2500 -695
rect -2460 -735 -2380 -695
rect -2580 -820 -2380 -735
rect -2230 -695 -2030 -620
rect -2230 -735 -2150 -695
rect -2110 -735 -2030 -695
rect -2230 -820 -2030 -735
rect -1880 -695 -1680 -620
rect -1880 -735 -1800 -695
rect -1760 -735 -1680 -695
rect -1880 -820 -1680 -735
rect 3370 -695 3570 -620
rect 3370 -735 3450 -695
rect 3490 -735 3570 -695
rect 3370 -820 3570 -735
rect 3720 -695 3920 -620
rect 3720 -735 3800 -695
rect 3840 -735 3920 -695
rect 3720 -820 3920 -735
rect 4070 -695 4270 -620
rect 4070 -735 4150 -695
rect 4190 -735 4270 -695
rect 4070 -820 4270 -735
rect 4420 -695 4620 -620
rect 4420 -735 4500 -695
rect 4540 -735 4620 -695
rect 4420 -820 4620 -735
rect 4770 -695 4970 -620
rect 4770 -735 4850 -695
rect 4890 -735 4970 -695
rect 4770 -820 4970 -735
rect -3280 -1045 -3080 -970
rect -3280 -1085 -3200 -1045
rect -3160 -1085 -3080 -1045
rect -3280 -1170 -3080 -1085
rect -2930 -1045 -2730 -970
rect -2930 -1085 -2850 -1045
rect -2810 -1085 -2730 -1045
rect -2930 -1170 -2730 -1085
rect -2580 -1045 -2380 -970
rect -2580 -1085 -2500 -1045
rect -2460 -1085 -2380 -1045
rect -2580 -1170 -2380 -1085
rect -2230 -1045 -2030 -970
rect -2230 -1085 -2150 -1045
rect -2110 -1085 -2030 -1045
rect -2230 -1170 -2030 -1085
rect -1880 -1045 -1680 -970
rect -1880 -1085 -1800 -1045
rect -1760 -1085 -1680 -1045
rect -1880 -1170 -1680 -1085
rect 3370 -1045 3570 -970
rect 3370 -1085 3450 -1045
rect 3490 -1085 3570 -1045
rect 3370 -1170 3570 -1085
rect 3720 -1045 3920 -970
rect 3720 -1085 3800 -1045
rect 3840 -1085 3920 -1045
rect 3720 -1170 3920 -1085
rect 4070 -1045 4270 -970
rect 4070 -1085 4150 -1045
rect 4190 -1085 4270 -1045
rect 4070 -1170 4270 -1085
rect 4420 -1045 4620 -970
rect 4420 -1085 4500 -1045
rect 4540 -1085 4620 -1045
rect 4420 -1170 4620 -1085
rect 4770 -1045 4970 -970
rect 4770 -1085 4850 -1045
rect 4890 -1085 4970 -1045
rect 4770 -1170 4970 -1085
rect -3280 -1395 -3080 -1320
rect -3280 -1435 -3200 -1395
rect -3160 -1435 -3080 -1395
rect -3280 -1520 -3080 -1435
rect -2930 -1395 -2730 -1320
rect -2930 -1435 -2850 -1395
rect -2810 -1435 -2730 -1395
rect -2930 -1520 -2730 -1435
rect -2580 -1395 -2380 -1320
rect -2580 -1435 -2500 -1395
rect -2460 -1435 -2380 -1395
rect -2580 -1520 -2380 -1435
rect -2230 -1395 -2030 -1320
rect -2230 -1435 -2150 -1395
rect -2110 -1435 -2030 -1395
rect -2230 -1520 -2030 -1435
rect -1880 -1395 -1680 -1320
rect -1880 -1435 -1800 -1395
rect -1760 -1435 -1680 -1395
rect -1880 -1520 -1680 -1435
rect -1530 -1395 -1330 -1320
rect -1530 -1435 -1450 -1395
rect -1410 -1435 -1330 -1395
rect -1530 -1520 -1330 -1435
rect -1180 -1395 -980 -1320
rect -1180 -1435 -1100 -1395
rect -1060 -1435 -980 -1395
rect -1180 -1520 -980 -1435
rect -830 -1395 -630 -1320
rect -830 -1435 -750 -1395
rect -710 -1435 -630 -1395
rect -830 -1520 -630 -1435
rect -480 -1395 -280 -1320
rect -480 -1435 -400 -1395
rect -360 -1435 -280 -1395
rect -480 -1520 -280 -1435
rect -130 -1395 70 -1320
rect -130 -1435 -50 -1395
rect -10 -1435 70 -1395
rect -130 -1520 70 -1435
rect 220 -1395 420 -1320
rect 220 -1435 300 -1395
rect 340 -1435 420 -1395
rect 220 -1520 420 -1435
rect 570 -1395 770 -1320
rect 570 -1435 650 -1395
rect 690 -1435 770 -1395
rect 570 -1520 770 -1435
rect 920 -1395 1120 -1320
rect 920 -1435 1000 -1395
rect 1040 -1435 1120 -1395
rect 920 -1520 1120 -1435
rect 1270 -1395 1470 -1320
rect 1270 -1435 1350 -1395
rect 1390 -1435 1470 -1395
rect 1270 -1520 1470 -1435
rect 1620 -1395 1820 -1320
rect 1620 -1435 1700 -1395
rect 1740 -1435 1820 -1395
rect 1620 -1520 1820 -1435
rect 1970 -1395 2170 -1320
rect 1970 -1435 2050 -1395
rect 2090 -1435 2170 -1395
rect 1970 -1520 2170 -1435
rect 2320 -1395 2520 -1320
rect 2320 -1435 2400 -1395
rect 2440 -1435 2520 -1395
rect 2320 -1520 2520 -1435
rect 2670 -1395 2870 -1320
rect 2670 -1435 2750 -1395
rect 2790 -1435 2870 -1395
rect 2670 -1520 2870 -1435
rect 3020 -1395 3220 -1320
rect 3020 -1435 3100 -1395
rect 3140 -1435 3220 -1395
rect 3020 -1520 3220 -1435
rect 3370 -1395 3570 -1320
rect 3370 -1435 3450 -1395
rect 3490 -1435 3570 -1395
rect 3370 -1520 3570 -1435
rect 3720 -1395 3920 -1320
rect 3720 -1435 3800 -1395
rect 3840 -1435 3920 -1395
rect 3720 -1520 3920 -1435
rect 4070 -1395 4270 -1320
rect 4070 -1435 4150 -1395
rect 4190 -1435 4270 -1395
rect 4070 -1520 4270 -1435
rect 4420 -1395 4620 -1320
rect 4420 -1435 4500 -1395
rect 4540 -1435 4620 -1395
rect 4420 -1520 4620 -1435
rect 4770 -1395 4970 -1320
rect 4770 -1435 4850 -1395
rect 4890 -1435 4970 -1395
rect 4770 -1520 4970 -1435
rect -3280 -1745 -3080 -1670
rect -3280 -1785 -3200 -1745
rect -3160 -1785 -3080 -1745
rect -3280 -1870 -3080 -1785
rect -2930 -1745 -2730 -1670
rect -2930 -1785 -2850 -1745
rect -2810 -1785 -2730 -1745
rect -2930 -1870 -2730 -1785
rect -2580 -1745 -2380 -1670
rect -2580 -1785 -2500 -1745
rect -2460 -1785 -2380 -1745
rect -2580 -1870 -2380 -1785
rect -2230 -1745 -2030 -1670
rect -2230 -1785 -2150 -1745
rect -2110 -1785 -2030 -1745
rect -2230 -1870 -2030 -1785
rect -1880 -1745 -1680 -1670
rect -1880 -1785 -1800 -1745
rect -1760 -1785 -1680 -1745
rect -1880 -1870 -1680 -1785
rect -1530 -1745 -1330 -1670
rect -1530 -1785 -1450 -1745
rect -1410 -1785 -1330 -1745
rect -1530 -1870 -1330 -1785
rect -1180 -1745 -980 -1670
rect -1180 -1785 -1100 -1745
rect -1060 -1785 -980 -1745
rect -1180 -1870 -980 -1785
rect -830 -1745 -630 -1670
rect -830 -1785 -750 -1745
rect -710 -1785 -630 -1745
rect -830 -1870 -630 -1785
rect -480 -1745 -280 -1670
rect -480 -1785 -400 -1745
rect -360 -1785 -280 -1745
rect -480 -1870 -280 -1785
rect -130 -1745 70 -1670
rect -130 -1785 -50 -1745
rect -10 -1785 70 -1745
rect -130 -1870 70 -1785
rect 220 -1745 420 -1670
rect 220 -1785 300 -1745
rect 340 -1785 420 -1745
rect 220 -1870 420 -1785
rect 570 -1745 770 -1670
rect 570 -1785 650 -1745
rect 690 -1785 770 -1745
rect 570 -1870 770 -1785
rect 920 -1745 1120 -1670
rect 920 -1785 1000 -1745
rect 1040 -1785 1120 -1745
rect 920 -1870 1120 -1785
rect 1270 -1745 1470 -1670
rect 1270 -1785 1350 -1745
rect 1390 -1785 1470 -1745
rect 1270 -1870 1470 -1785
rect 1620 -1745 1820 -1670
rect 1620 -1785 1700 -1745
rect 1740 -1785 1820 -1745
rect 1620 -1870 1820 -1785
rect 1970 -1745 2170 -1670
rect 1970 -1785 2050 -1745
rect 2090 -1785 2170 -1745
rect 1970 -1870 2170 -1785
rect 2320 -1745 2520 -1670
rect 2320 -1785 2400 -1745
rect 2440 -1785 2520 -1745
rect 2320 -1870 2520 -1785
rect 2670 -1745 2870 -1670
rect 2670 -1785 2750 -1745
rect 2790 -1785 2870 -1745
rect 2670 -1870 2870 -1785
rect 3020 -1745 3220 -1670
rect 3020 -1785 3100 -1745
rect 3140 -1785 3220 -1745
rect 3020 -1870 3220 -1785
rect 3370 -1745 3570 -1670
rect 3370 -1785 3450 -1745
rect 3490 -1785 3570 -1745
rect 3370 -1870 3570 -1785
rect 3720 -1745 3920 -1670
rect 3720 -1785 3800 -1745
rect 3840 -1785 3920 -1745
rect 3720 -1870 3920 -1785
rect 4070 -1745 4270 -1670
rect 4070 -1785 4150 -1745
rect 4190 -1785 4270 -1745
rect 4070 -1870 4270 -1785
rect 4420 -1745 4620 -1670
rect 4420 -1785 4500 -1745
rect 4540 -1785 4620 -1745
rect 4420 -1870 4620 -1785
rect 4770 -1745 4970 -1670
rect 4770 -1785 4850 -1745
rect 4890 -1785 4970 -1745
rect 4770 -1870 4970 -1785
rect -3280 -2095 -3080 -2020
rect -3280 -2135 -3200 -2095
rect -3160 -2135 -3080 -2095
rect -3280 -2220 -3080 -2135
rect -2930 -2095 -2730 -2020
rect -2930 -2135 -2850 -2095
rect -2810 -2135 -2730 -2095
rect -2930 -2220 -2730 -2135
rect -2580 -2095 -2380 -2020
rect -2580 -2135 -2500 -2095
rect -2460 -2135 -2380 -2095
rect -2580 -2220 -2380 -2135
rect -2230 -2095 -2030 -2020
rect -2230 -2135 -2150 -2095
rect -2110 -2135 -2030 -2095
rect -2230 -2220 -2030 -2135
rect -1880 -2095 -1680 -2020
rect -1880 -2135 -1800 -2095
rect -1760 -2135 -1680 -2095
rect -1880 -2220 -1680 -2135
rect -1530 -2095 -1330 -2020
rect -1530 -2135 -1450 -2095
rect -1410 -2135 -1330 -2095
rect -1530 -2220 -1330 -2135
rect -1180 -2095 -980 -2020
rect -1180 -2135 -1100 -2095
rect -1060 -2135 -980 -2095
rect -1180 -2220 -980 -2135
rect -830 -2095 -630 -2020
rect -830 -2135 -750 -2095
rect -710 -2135 -630 -2095
rect -830 -2220 -630 -2135
rect -480 -2095 -280 -2020
rect -480 -2135 -400 -2095
rect -360 -2135 -280 -2095
rect -480 -2220 -280 -2135
rect -130 -2095 70 -2020
rect -130 -2135 -50 -2095
rect -10 -2135 70 -2095
rect -130 -2220 70 -2135
rect 220 -2095 420 -2020
rect 220 -2135 300 -2095
rect 340 -2135 420 -2095
rect 220 -2220 420 -2135
rect 570 -2095 770 -2020
rect 570 -2135 650 -2095
rect 690 -2135 770 -2095
rect 570 -2220 770 -2135
rect 920 -2095 1120 -2020
rect 920 -2135 1000 -2095
rect 1040 -2135 1120 -2095
rect 920 -2220 1120 -2135
rect 1270 -2095 1470 -2020
rect 1270 -2135 1350 -2095
rect 1390 -2135 1470 -2095
rect 1270 -2220 1470 -2135
rect 1620 -2095 1820 -2020
rect 1620 -2135 1700 -2095
rect 1740 -2135 1820 -2095
rect 1620 -2220 1820 -2135
rect 1970 -2095 2170 -2020
rect 1970 -2135 2050 -2095
rect 2090 -2135 2170 -2095
rect 1970 -2220 2170 -2135
rect 2320 -2095 2520 -2020
rect 2320 -2135 2400 -2095
rect 2440 -2135 2520 -2095
rect 2320 -2220 2520 -2135
rect 2670 -2095 2870 -2020
rect 2670 -2135 2750 -2095
rect 2790 -2135 2870 -2095
rect 2670 -2220 2870 -2135
rect 3020 -2095 3220 -2020
rect 3020 -2135 3100 -2095
rect 3140 -2135 3220 -2095
rect 3020 -2220 3220 -2135
rect 3370 -2095 3570 -2020
rect 3370 -2135 3450 -2095
rect 3490 -2135 3570 -2095
rect 3370 -2220 3570 -2135
rect 3720 -2095 3920 -2020
rect 3720 -2135 3800 -2095
rect 3840 -2135 3920 -2095
rect 3720 -2220 3920 -2135
rect 4070 -2095 4270 -2020
rect 4070 -2135 4150 -2095
rect 4190 -2135 4270 -2095
rect 4070 -2220 4270 -2135
rect 4420 -2095 4620 -2020
rect 4420 -2135 4500 -2095
rect 4540 -2135 4620 -2095
rect 4420 -2220 4620 -2135
rect 4770 -2095 4970 -2020
rect 4770 -2135 4850 -2095
rect 4890 -2135 4970 -2095
rect 4770 -2220 4970 -2135
<< mimcapcontact >>
rect -3200 3815 -3160 3855
rect -2850 3815 -2810 3855
rect -2500 3815 -2460 3855
rect -2150 3815 -2110 3855
rect -1800 3815 -1760 3855
rect -1450 3815 -1410 3855
rect -1100 3815 -1060 3855
rect -750 3815 -710 3855
rect -400 3815 -360 3855
rect -50 3815 -10 3855
rect 300 3815 340 3855
rect 650 3815 690 3855
rect 1000 3815 1040 3855
rect 1350 3815 1390 3855
rect 1700 3815 1740 3855
rect 2050 3815 2090 3855
rect 2400 3815 2440 3855
rect 2750 3815 2790 3855
rect 3100 3815 3140 3855
rect 3450 3815 3490 3855
rect 3800 3815 3840 3855
rect 4150 3815 4190 3855
rect 4500 3815 4540 3855
rect 4850 3815 4890 3855
rect -3200 3465 -3160 3505
rect -2850 3465 -2810 3505
rect -2500 3465 -2460 3505
rect -2150 3465 -2110 3505
rect -1800 3465 -1760 3505
rect -1450 3465 -1410 3505
rect -1100 3465 -1060 3505
rect -750 3465 -710 3505
rect -400 3465 -360 3505
rect -50 3465 -10 3505
rect 300 3465 340 3505
rect 650 3465 690 3505
rect 1000 3465 1040 3505
rect 1350 3465 1390 3505
rect 1700 3465 1740 3505
rect 2050 3465 2090 3505
rect 2400 3465 2440 3505
rect 2750 3465 2790 3505
rect 3100 3465 3140 3505
rect 3450 3465 3490 3505
rect 3800 3465 3840 3505
rect 4150 3465 4190 3505
rect 4500 3465 4540 3505
rect 4850 3465 4890 3505
rect -3200 3115 -3160 3155
rect -2850 3115 -2810 3155
rect -2500 3115 -2460 3155
rect -2150 3115 -2110 3155
rect -1800 3115 -1760 3155
rect -1450 3115 -1410 3155
rect -1100 3115 -1060 3155
rect -750 3115 -710 3155
rect -400 3115 -360 3155
rect -50 3105 -10 3145
rect 300 3105 340 3145
rect 650 3105 690 3145
rect 1000 3105 1040 3145
rect 1350 3105 1390 3145
rect 1700 3105 1740 3145
rect 2050 3115 2090 3155
rect 2400 3115 2440 3155
rect 2750 3115 2790 3155
rect 3100 3115 3140 3155
rect 3450 3115 3490 3155
rect 3800 3115 3840 3155
rect 4150 3115 4190 3155
rect 4500 3115 4540 3155
rect 4850 3115 4890 3155
rect -3200 2765 -3160 2805
rect -2850 2765 -2810 2805
rect -2500 2765 -2460 2805
rect -2150 2765 -2110 2805
rect -1800 2765 -1760 2805
rect -1450 2765 -1410 2805
rect -1100 2765 -1060 2805
rect -750 2765 -710 2805
rect 2400 2765 2440 2805
rect 2750 2765 2790 2805
rect 3100 2765 3140 2805
rect 3450 2765 3490 2805
rect 3800 2765 3840 2805
rect 4150 2765 4190 2805
rect 4500 2765 4540 2805
rect 4850 2765 4890 2805
rect -3200 2415 -3160 2455
rect -2850 2415 -2810 2455
rect -2500 2415 -2460 2455
rect -2150 2415 -2110 2455
rect -1800 2415 -1760 2455
rect -1450 2415 -1410 2455
rect -1100 2415 -1060 2455
rect -750 2415 -710 2455
rect 2400 2415 2440 2455
rect 2750 2415 2790 2455
rect 3100 2415 3140 2455
rect 3450 2415 3490 2455
rect 3800 2415 3840 2455
rect 4150 2415 4190 2455
rect 4500 2415 4540 2455
rect 4850 2415 4890 2455
rect -3200 2065 -3160 2105
rect -2850 2065 -2810 2105
rect -2500 2065 -2460 2105
rect -2150 2065 -2110 2105
rect -1800 2065 -1760 2105
rect 3450 2065 3490 2105
rect 3800 2065 3840 2105
rect 4150 2065 4190 2105
rect 4500 2065 4540 2105
rect 4850 2065 4890 2105
rect -3200 1715 -3160 1755
rect -2850 1715 -2810 1755
rect -2500 1715 -2460 1755
rect -2150 1715 -2110 1755
rect -1800 1715 -1760 1755
rect 3450 1715 3490 1755
rect 3800 1715 3840 1755
rect 4150 1715 4190 1755
rect 4500 1715 4540 1755
rect 4850 1715 4890 1755
rect -3200 1365 -3160 1405
rect -2850 1365 -2810 1405
rect -2500 1365 -2460 1405
rect -2150 1365 -2110 1405
rect -1800 1365 -1760 1405
rect 3450 1365 3490 1405
rect 3800 1365 3840 1405
rect 4150 1365 4190 1405
rect 4500 1365 4540 1405
rect 4850 1365 4890 1405
rect -3200 1015 -3160 1055
rect -2850 1015 -2810 1055
rect -2500 1015 -2460 1055
rect -2150 1015 -2110 1055
rect -1800 1015 -1760 1055
rect 3450 1015 3490 1055
rect 3800 1015 3840 1055
rect 4150 1015 4190 1055
rect 4500 1015 4540 1055
rect 4850 1015 4890 1055
rect -3200 665 -3160 705
rect -2850 665 -2810 705
rect -2500 665 -2460 705
rect -2150 665 -2110 705
rect -1800 665 -1760 705
rect 3450 665 3490 705
rect 3800 665 3840 705
rect 4150 665 4190 705
rect 4500 665 4540 705
rect 4850 665 4890 705
rect -3200 315 -3160 355
rect -2850 315 -2810 355
rect -2500 315 -2460 355
rect -2150 315 -2110 355
rect -1800 315 -1760 355
rect 3450 315 3490 355
rect 3800 315 3840 355
rect 4150 315 4190 355
rect 4500 315 4540 355
rect 4850 315 4890 355
rect -3200 -35 -3160 5
rect -2850 -35 -2810 5
rect -2500 -35 -2460 5
rect -2150 -35 -2110 5
rect -1800 -35 -1760 5
rect 3450 -35 3490 5
rect 3800 -35 3840 5
rect 4150 -35 4190 5
rect 4500 -35 4540 5
rect 4850 -35 4890 5
rect -3200 -385 -3160 -345
rect -2850 -385 -2810 -345
rect -2500 -385 -2460 -345
rect -2150 -385 -2110 -345
rect -1800 -385 -1760 -345
rect 3450 -385 3490 -345
rect 3800 -385 3840 -345
rect 4150 -385 4190 -345
rect 4500 -385 4540 -345
rect 4850 -385 4890 -345
rect -3200 -735 -3160 -695
rect -2850 -735 -2810 -695
rect -2500 -735 -2460 -695
rect -2150 -735 -2110 -695
rect -1800 -735 -1760 -695
rect 3450 -735 3490 -695
rect 3800 -735 3840 -695
rect 4150 -735 4190 -695
rect 4500 -735 4540 -695
rect 4850 -735 4890 -695
rect -3200 -1085 -3160 -1045
rect -2850 -1085 -2810 -1045
rect -2500 -1085 -2460 -1045
rect -2150 -1085 -2110 -1045
rect -1800 -1085 -1760 -1045
rect 3450 -1085 3490 -1045
rect 3800 -1085 3840 -1045
rect 4150 -1085 4190 -1045
rect 4500 -1085 4540 -1045
rect 4850 -1085 4890 -1045
rect -3200 -1435 -3160 -1395
rect -2850 -1435 -2810 -1395
rect -2500 -1435 -2460 -1395
rect -2150 -1435 -2110 -1395
rect -1800 -1435 -1760 -1395
rect -1450 -1435 -1410 -1395
rect -1100 -1435 -1060 -1395
rect -750 -1435 -710 -1395
rect -400 -1435 -360 -1395
rect -50 -1435 -10 -1395
rect 300 -1435 340 -1395
rect 650 -1435 690 -1395
rect 1000 -1435 1040 -1395
rect 1350 -1435 1390 -1395
rect 1700 -1435 1740 -1395
rect 2050 -1435 2090 -1395
rect 2400 -1435 2440 -1395
rect 2750 -1435 2790 -1395
rect 3100 -1435 3140 -1395
rect 3450 -1435 3490 -1395
rect 3800 -1435 3840 -1395
rect 4150 -1435 4190 -1395
rect 4500 -1435 4540 -1395
rect 4850 -1435 4890 -1395
rect -3200 -1785 -3160 -1745
rect -2850 -1785 -2810 -1745
rect -2500 -1785 -2460 -1745
rect -2150 -1785 -2110 -1745
rect -1800 -1785 -1760 -1745
rect -1450 -1785 -1410 -1745
rect -1100 -1785 -1060 -1745
rect -750 -1785 -710 -1745
rect -400 -1785 -360 -1745
rect -50 -1785 -10 -1745
rect 300 -1785 340 -1745
rect 650 -1785 690 -1745
rect 1000 -1785 1040 -1745
rect 1350 -1785 1390 -1745
rect 1700 -1785 1740 -1745
rect 2050 -1785 2090 -1745
rect 2400 -1785 2440 -1745
rect 2750 -1785 2790 -1745
rect 3100 -1785 3140 -1745
rect 3450 -1785 3490 -1745
rect 3800 -1785 3840 -1745
rect 4150 -1785 4190 -1745
rect 4500 -1785 4540 -1745
rect 4850 -1785 4890 -1745
rect -3200 -2135 -3160 -2095
rect -2850 -2135 -2810 -2095
rect -2500 -2135 -2460 -2095
rect -2150 -2135 -2110 -2095
rect -1800 -2135 -1760 -2095
rect -1450 -2135 -1410 -2095
rect -1100 -2135 -1060 -2095
rect -750 -2135 -710 -2095
rect -400 -2135 -360 -2095
rect -50 -2135 -10 -2095
rect 300 -2135 340 -2095
rect 650 -2135 690 -2095
rect 1000 -2135 1040 -2095
rect 1350 -2135 1390 -2095
rect 1700 -2135 1740 -2095
rect 2050 -2135 2090 -2095
rect 2400 -2135 2440 -2095
rect 2750 -2135 2790 -2095
rect 3100 -2135 3140 -2095
rect 3450 -2135 3490 -2095
rect 3800 -2135 3840 -2095
rect 4150 -2135 4190 -2095
rect 4500 -2135 4540 -2095
rect 4850 -2135 4890 -2095
<< metal4 >>
rect -3850 4280 5140 4285
rect -3850 4240 825 4280
rect 865 4240 5140 4280
rect -3850 4235 5140 4240
rect -3205 3855 -2455 3860
rect -3205 3815 -3200 3855
rect -3160 3815 -2850 3855
rect -2810 3815 -2500 3855
rect -2460 3815 -2455 3855
rect -3205 3810 -2455 3815
rect -2505 3510 -2455 3810
rect -2155 3855 -2105 3860
rect -2155 3815 -2150 3855
rect -2110 3815 -2105 3855
rect -2155 3510 -2105 3815
rect -1805 3855 -1755 3860
rect -1805 3815 -1800 3855
rect -1760 3815 -1755 3855
rect -1805 3510 -1755 3815
rect -1455 3855 -1405 3860
rect -1455 3815 -1450 3855
rect -1410 3815 -1405 3855
rect -1455 3510 -1405 3815
rect -1105 3855 -1055 3860
rect -1105 3815 -1100 3855
rect -1060 3815 -1055 3855
rect -1105 3510 -1055 3815
rect -755 3855 -705 3860
rect -755 3815 -750 3855
rect -710 3815 -705 3855
rect -755 3510 -705 3815
rect -405 3855 -355 3860
rect -405 3815 -400 3855
rect -360 3815 -355 3855
rect -405 3510 -355 3815
rect -55 3855 -5 3860
rect -55 3815 -50 3855
rect -10 3815 -5 3855
rect -55 3510 -5 3815
rect 295 3855 345 3860
rect 295 3815 300 3855
rect 340 3815 345 3855
rect 295 3510 345 3815
rect 645 3855 695 3860
rect 645 3815 650 3855
rect 690 3815 695 3855
rect 645 3510 695 3815
rect -3205 3505 695 3510
rect -3205 3465 -3200 3505
rect -3160 3465 -2850 3505
rect -2810 3465 -2500 3505
rect -2460 3465 -2150 3505
rect -2110 3465 -1800 3505
rect -1760 3465 -1450 3505
rect -1410 3465 -1100 3505
rect -1060 3465 -750 3505
rect -710 3465 -400 3505
rect -360 3465 -50 3505
rect -10 3465 300 3505
rect 340 3465 650 3505
rect 690 3465 695 3505
rect -3205 3460 695 3465
rect -2505 3160 -2455 3460
rect -3205 3155 -2105 3160
rect -3205 3115 -3200 3155
rect -3160 3115 -2850 3155
rect -2810 3115 -2500 3155
rect -2460 3115 -2150 3155
rect -2110 3115 -2105 3155
rect -3205 3110 -2105 3115
rect -1805 3155 -1755 3460
rect -1805 3115 -1800 3155
rect -1760 3115 -1755 3155
rect -2505 2810 -2455 3110
rect -3205 2805 -2105 2810
rect -3205 2765 -3200 2805
rect -3160 2765 -2850 2805
rect -2810 2765 -2500 2805
rect -2460 2765 -2150 2805
rect -2110 2765 -2105 2805
rect -3205 2760 -2105 2765
rect -1805 2805 -1755 3115
rect -1805 2765 -1800 2805
rect -1760 2765 -1755 2805
rect -1805 2760 -1755 2765
rect -1455 3155 -1405 3460
rect -1455 3115 -1450 3155
rect -1410 3115 -1405 3155
rect -1455 2805 -1405 3115
rect -1455 2765 -1450 2805
rect -1410 2765 -1405 2805
rect -2505 2460 -2455 2760
rect -3205 2455 -1755 2460
rect -3205 2415 -3200 2455
rect -3160 2415 -2850 2455
rect -2810 2415 -2500 2455
rect -2460 2415 -2150 2455
rect -2110 2415 -1800 2455
rect -1760 2415 -1755 2455
rect -3205 2410 -1755 2415
rect -1455 2455 -1405 2765
rect -1455 2415 -1450 2455
rect -1410 2415 -1405 2455
rect -1455 2410 -1405 2415
rect -1105 3155 -1055 3460
rect -1105 3115 -1100 3155
rect -1060 3115 -1055 3155
rect -1105 2805 -1055 3115
rect -1105 2765 -1100 2805
rect -1060 2765 -1055 2805
rect -1105 2455 -1055 2765
rect -1105 2415 -1100 2455
rect -1060 2415 -1055 2455
rect -1105 2410 -1055 2415
rect -755 3155 -705 3460
rect -755 3115 -750 3155
rect -710 3115 -705 3155
rect -755 2805 -705 3115
rect -405 3155 -355 3460
rect -405 3115 -400 3155
rect -360 3115 -355 3155
rect -405 3110 -355 3115
rect -55 3145 -5 3460
rect -55 3105 -50 3145
rect -10 3105 -5 3145
rect -55 3100 -5 3105
rect 295 3145 345 3460
rect 295 3105 300 3145
rect 340 3105 345 3145
rect 295 3100 345 3105
rect 645 3145 695 3460
rect 645 3105 650 3145
rect 690 3105 695 3145
rect 645 3100 695 3105
rect 995 3855 1045 3860
rect 995 3815 1000 3855
rect 1040 3815 1045 3855
rect 995 3510 1045 3815
rect 1345 3855 1395 3860
rect 1345 3815 1350 3855
rect 1390 3815 1395 3855
rect 1345 3510 1395 3815
rect 1695 3855 1745 3860
rect 1695 3815 1700 3855
rect 1740 3815 1745 3855
rect 1695 3510 1745 3815
rect 2045 3855 2095 3860
rect 2045 3815 2050 3855
rect 2090 3815 2095 3855
rect 2045 3510 2095 3815
rect 2395 3855 2445 3860
rect 2395 3815 2400 3855
rect 2440 3815 2445 3855
rect 2395 3510 2445 3815
rect 2745 3855 2795 3860
rect 2745 3815 2750 3855
rect 2790 3815 2795 3855
rect 2745 3510 2795 3815
rect 3095 3855 3145 3860
rect 3095 3815 3100 3855
rect 3140 3815 3145 3855
rect 3095 3510 3145 3815
rect 3445 3855 3495 3860
rect 3445 3815 3450 3855
rect 3490 3815 3495 3855
rect 3445 3510 3495 3815
rect 3795 3855 3845 3860
rect 3795 3815 3800 3855
rect 3840 3815 3845 3855
rect 3795 3510 3845 3815
rect 4145 3855 4895 3860
rect 4145 3815 4150 3855
rect 4190 3815 4500 3855
rect 4540 3815 4850 3855
rect 4890 3815 4895 3855
rect 4145 3810 4895 3815
rect 4145 3510 4195 3810
rect 995 3505 4895 3510
rect 995 3465 1000 3505
rect 1040 3465 1350 3505
rect 1390 3465 1700 3505
rect 1740 3465 2050 3505
rect 2090 3465 2400 3505
rect 2440 3465 2750 3505
rect 2790 3465 3100 3505
rect 3140 3465 3450 3505
rect 3490 3465 3800 3505
rect 3840 3465 4150 3505
rect 4190 3465 4500 3505
rect 4540 3465 4850 3505
rect 4890 3465 4895 3505
rect 995 3460 4895 3465
rect 995 3145 1045 3460
rect 995 3105 1000 3145
rect 1040 3105 1045 3145
rect 995 3100 1045 3105
rect 1345 3145 1395 3460
rect 1345 3105 1350 3145
rect 1390 3105 1395 3145
rect 1345 3100 1395 3105
rect 1695 3145 1745 3460
rect 1695 3105 1700 3145
rect 1740 3105 1745 3145
rect 2045 3155 2095 3460
rect 2045 3115 2050 3155
rect 2090 3115 2095 3155
rect 2045 3110 2095 3115
rect 2395 3155 2445 3460
rect 2395 3115 2400 3155
rect 2440 3115 2445 3155
rect 1695 3100 1745 3105
rect -755 2765 -750 2805
rect -710 2765 -705 2805
rect -755 2455 -705 2765
rect -755 2415 -750 2455
rect -710 2415 -705 2455
rect -755 2410 -705 2415
rect 2395 2805 2445 3115
rect 2395 2765 2400 2805
rect 2440 2765 2445 2805
rect 2395 2455 2445 2765
rect 2395 2415 2400 2455
rect 2440 2415 2445 2455
rect 2395 2410 2445 2415
rect 2745 3155 2795 3460
rect 2745 3115 2750 3155
rect 2790 3115 2795 3155
rect 2745 2805 2795 3115
rect 2745 2765 2750 2805
rect 2790 2765 2795 2805
rect 2745 2455 2795 2765
rect 2745 2415 2750 2455
rect 2790 2415 2795 2455
rect 2745 2410 2795 2415
rect 3095 3155 3145 3460
rect 3095 3115 3100 3155
rect 3140 3115 3145 3155
rect 3095 2805 3145 3115
rect 3095 2765 3100 2805
rect 3140 2765 3145 2805
rect 3095 2455 3145 2765
rect 3445 3155 3495 3460
rect 4145 3160 4195 3460
rect 3445 3115 3450 3155
rect 3490 3115 3495 3155
rect 3445 2805 3495 3115
rect 3795 3155 4895 3160
rect 3795 3115 3800 3155
rect 3840 3115 4150 3155
rect 4190 3115 4500 3155
rect 4540 3115 4850 3155
rect 4890 3115 4895 3155
rect 3795 3110 4895 3115
rect 4145 2810 4195 3110
rect 3445 2765 3450 2805
rect 3490 2765 3495 2805
rect 3445 2760 3495 2765
rect 3795 2805 4895 2810
rect 3795 2765 3800 2805
rect 3840 2765 4150 2805
rect 4190 2765 4500 2805
rect 4540 2765 4850 2805
rect 4890 2765 4895 2805
rect 3795 2760 4895 2765
rect 4145 2460 4195 2760
rect 3095 2415 3100 2455
rect 3140 2415 3145 2455
rect 3095 2410 3145 2415
rect 3445 2455 4895 2460
rect 3445 2415 3450 2455
rect 3490 2415 3800 2455
rect 3840 2415 4150 2455
rect 4190 2415 4500 2455
rect 4540 2415 4850 2455
rect 4890 2415 4895 2455
rect 3445 2410 4895 2415
rect -2505 2110 -2455 2410
rect 4145 2110 4195 2410
rect -3205 2105 -1755 2110
rect -3205 2065 -3200 2105
rect -3160 2065 -2850 2105
rect -2810 2065 -2500 2105
rect -2460 2065 -2150 2105
rect -2110 2065 -1800 2105
rect -1760 2065 -1755 2105
rect -3205 2060 -1755 2065
rect 3445 2105 4895 2110
rect 3445 2065 3450 2105
rect 3490 2065 3800 2105
rect 3840 2065 4150 2105
rect 4190 2065 4500 2105
rect 4540 2065 4850 2105
rect 4890 2065 4895 2105
rect 3445 2060 4895 2065
rect -2505 1760 -2455 2060
rect 4145 1760 4195 2060
rect -3205 1755 -1755 1760
rect -3205 1715 -3200 1755
rect -3160 1715 -2850 1755
rect -2810 1715 -2500 1755
rect -2460 1715 -2150 1755
rect -2110 1715 -1800 1755
rect -1760 1715 -1755 1755
rect -3205 1710 -1755 1715
rect 3445 1755 4895 1760
rect 3445 1715 3450 1755
rect 3490 1715 3800 1755
rect 3840 1715 4150 1755
rect 4190 1715 4500 1755
rect 4540 1715 4850 1755
rect 4890 1715 4895 1755
rect 3445 1710 4895 1715
rect -2505 1410 -2455 1710
rect 4145 1410 4195 1710
rect -3205 1405 -1755 1410
rect -3205 1365 -3200 1405
rect -3160 1365 -2850 1405
rect -2810 1365 -2500 1405
rect -2460 1365 -2150 1405
rect -2110 1365 -1800 1405
rect -1760 1365 -1755 1405
rect -3205 1360 -1755 1365
rect 3445 1405 4895 1410
rect 3445 1365 3450 1405
rect 3490 1365 3800 1405
rect 3840 1365 4150 1405
rect 4190 1365 4500 1405
rect 4540 1365 4850 1405
rect 4890 1365 4895 1405
rect 3445 1360 4895 1365
rect -2505 1060 -2455 1360
rect 4145 1060 4195 1360
rect -3205 1055 -1755 1060
rect -3205 1015 -3200 1055
rect -3160 1015 -2850 1055
rect -2810 1015 -2500 1055
rect -2460 1015 -2150 1055
rect -2110 1015 -1800 1055
rect -1760 1015 -1755 1055
rect -3205 1010 -1755 1015
rect 3445 1055 4895 1060
rect 3445 1015 3450 1055
rect 3490 1015 3800 1055
rect 3840 1015 4150 1055
rect 4190 1015 4500 1055
rect 4540 1015 4850 1055
rect 4890 1015 4895 1055
rect 3445 1010 4895 1015
rect -2505 710 -2455 1010
rect 4145 710 4195 1010
rect -3205 705 -1755 710
rect -3205 665 -3200 705
rect -3160 665 -2850 705
rect -2810 665 -2500 705
rect -2460 665 -2150 705
rect -2110 665 -1800 705
rect -1760 665 -1755 705
rect -3205 660 -1755 665
rect 3445 705 4895 710
rect 3445 665 3450 705
rect 3490 665 3800 705
rect 3840 665 4150 705
rect 4190 665 4500 705
rect 4540 665 4850 705
rect 4890 665 4895 705
rect 3445 660 4895 665
rect -2505 360 -2455 660
rect 4145 360 4195 660
rect -3205 355 -1495 360
rect -3205 315 -3200 355
rect -3160 315 -2850 355
rect -2810 315 -2500 355
rect -2460 315 -2150 355
rect -2110 315 -1800 355
rect -1760 315 -1540 355
rect -1500 315 -1495 355
rect -3205 310 -1495 315
rect 3185 355 4895 360
rect 3185 315 3190 355
rect 3230 315 3450 355
rect 3490 315 3800 355
rect 3840 315 4150 355
rect 4190 315 4500 355
rect 4540 315 4850 355
rect 4890 315 4895 355
rect 3185 310 4895 315
rect -2505 10 -2455 310
rect 4145 10 4195 310
rect -3205 5 -1755 10
rect -3205 -35 -3200 5
rect -3160 -35 -2850 5
rect -2810 -35 -2500 5
rect -2460 -35 -2150 5
rect -2110 -35 -1800 5
rect -1760 -35 -1755 5
rect -3205 -40 -1755 -35
rect 3445 5 4895 10
rect 3445 -35 3450 5
rect 3490 -35 3800 5
rect 3840 -35 4150 5
rect 4190 -35 4500 5
rect 4540 -35 4850 5
rect 4890 -35 4895 5
rect 3445 -40 4895 -35
rect -2505 -340 -2455 -40
rect 4145 -340 4195 -40
rect -3205 -345 -1755 -340
rect -3205 -385 -3200 -345
rect -3160 -385 -2850 -345
rect -2810 -385 -2500 -345
rect -2460 -385 -2150 -345
rect -2110 -385 -1800 -345
rect -1760 -385 -1755 -345
rect -3205 -390 -1755 -385
rect 3445 -345 4895 -340
rect 3445 -385 3450 -345
rect 3490 -385 3800 -345
rect 3840 -385 4150 -345
rect 4190 -385 4500 -345
rect 4540 -385 4850 -345
rect 4890 -385 4895 -345
rect 3445 -390 4895 -385
rect -2505 -690 -2455 -390
rect 4145 -690 4195 -390
rect -3205 -695 -1755 -690
rect -3205 -735 -3200 -695
rect -3160 -735 -2850 -695
rect -2810 -735 -2500 -695
rect -2460 -735 -2150 -695
rect -2110 -735 -1800 -695
rect -1760 -735 -1755 -695
rect -3205 -740 -1755 -735
rect 3445 -695 4895 -690
rect 3445 -735 3450 -695
rect 3490 -735 3800 -695
rect 3840 -735 4150 -695
rect 4190 -735 4500 -695
rect 4540 -735 4850 -695
rect 4890 -735 4895 -695
rect 3445 -740 4895 -735
rect -2505 -1040 -2455 -740
rect 4145 -1040 4195 -740
rect -3205 -1045 -1755 -1040
rect -3205 -1085 -3200 -1045
rect -3160 -1085 -2850 -1045
rect -2810 -1085 -2500 -1045
rect -2460 -1085 -2150 -1045
rect -2110 -1085 -1800 -1045
rect -1760 -1085 -1755 -1045
rect -3205 -1090 -1755 -1085
rect 3445 -1045 4895 -1040
rect 3445 -1085 3450 -1045
rect 3490 -1085 3800 -1045
rect 3840 -1085 4150 -1045
rect 4190 -1085 4500 -1045
rect 4540 -1085 4850 -1045
rect 4890 -1085 4895 -1045
rect 3445 -1090 4895 -1085
rect -2505 -1390 -2455 -1090
rect 4145 -1390 4195 -1090
rect -3205 -1395 -1755 -1390
rect -3205 -1435 -3200 -1395
rect -3160 -1435 -2850 -1395
rect -2810 -1435 -2500 -1395
rect -2460 -1435 -2150 -1395
rect -2110 -1435 -1800 -1395
rect -1760 -1435 -1755 -1395
rect -3205 -1440 -1755 -1435
rect -1455 -1395 -1405 -1390
rect -1455 -1435 -1450 -1395
rect -1410 -1435 -1405 -1395
rect -2505 -1740 -2455 -1440
rect -1455 -1740 -1405 -1435
rect -1105 -1395 -1055 -1390
rect -1105 -1435 -1100 -1395
rect -1060 -1435 -1055 -1395
rect -1105 -1740 -1055 -1435
rect -755 -1395 -705 -1390
rect -755 -1435 -750 -1395
rect -710 -1435 -705 -1395
rect -755 -1740 -705 -1435
rect -405 -1395 -355 -1390
rect -405 -1435 -400 -1395
rect -360 -1435 -355 -1395
rect -405 -1740 -355 -1435
rect -55 -1395 -5 -1390
rect -55 -1435 -50 -1395
rect -10 -1435 -5 -1395
rect -55 -1740 -5 -1435
rect 295 -1395 345 -1390
rect 295 -1435 300 -1395
rect 340 -1435 345 -1395
rect 295 -1740 345 -1435
rect 645 -1395 695 -1390
rect 645 -1435 650 -1395
rect 690 -1435 695 -1395
rect 645 -1740 695 -1435
rect -3205 -1745 695 -1740
rect -3205 -1785 -3200 -1745
rect -3160 -1785 -2850 -1745
rect -2810 -1785 -2500 -1745
rect -2460 -1785 -2150 -1745
rect -2110 -1785 -1800 -1745
rect -1760 -1785 -1450 -1745
rect -1410 -1785 -1100 -1745
rect -1060 -1785 -750 -1745
rect -710 -1785 -400 -1745
rect -360 -1785 -50 -1745
rect -10 -1785 300 -1745
rect 340 -1785 650 -1745
rect 690 -1785 695 -1745
rect -3205 -1790 695 -1785
rect -2505 -2090 -2455 -1790
rect -3205 -2095 -2455 -2090
rect -3205 -2135 -3200 -2095
rect -3160 -2135 -2850 -2095
rect -2810 -2135 -2500 -2095
rect -2460 -2135 -2455 -2095
rect -3205 -2140 -2455 -2135
rect -2155 -2095 -2105 -1790
rect -2155 -2135 -2150 -2095
rect -2110 -2135 -2105 -2095
rect -2155 -2140 -2105 -2135
rect -1805 -2095 -1755 -1790
rect -1805 -2135 -1800 -2095
rect -1760 -2135 -1755 -2095
rect -1805 -2140 -1755 -2135
rect -1455 -2095 -1405 -1790
rect -1455 -2135 -1450 -2095
rect -1410 -2135 -1405 -2095
rect -1455 -2140 -1405 -2135
rect -1105 -2095 -1055 -1790
rect -1105 -2135 -1100 -2095
rect -1060 -2135 -1055 -2095
rect -1105 -2140 -1055 -2135
rect -755 -2095 -705 -1790
rect -755 -2135 -750 -2095
rect -710 -2135 -705 -2095
rect -755 -2140 -705 -2135
rect -405 -2095 -355 -1790
rect -405 -2135 -400 -2095
rect -360 -2135 -355 -2095
rect -405 -2140 -355 -2135
rect -55 -2095 -5 -1790
rect -55 -2135 -50 -2095
rect -10 -2135 -5 -2095
rect -55 -2140 -5 -2135
rect 295 -2095 345 -1790
rect 295 -2135 300 -2095
rect 340 -2135 345 -2095
rect 295 -2140 345 -2135
rect 645 -2095 695 -1790
rect 645 -2135 650 -2095
rect 690 -2135 695 -2095
rect 645 -2140 695 -2135
rect 995 -1395 1045 -1390
rect 995 -1435 1000 -1395
rect 1040 -1435 1045 -1395
rect 995 -1740 1045 -1435
rect 1345 -1395 1395 -1390
rect 1345 -1435 1350 -1395
rect 1390 -1435 1395 -1395
rect 1345 -1740 1395 -1435
rect 1695 -1395 1745 -1390
rect 1695 -1435 1700 -1395
rect 1740 -1435 1745 -1395
rect 1695 -1740 1745 -1435
rect 2045 -1395 2095 -1390
rect 2045 -1435 2050 -1395
rect 2090 -1435 2095 -1395
rect 2045 -1740 2095 -1435
rect 2395 -1395 2445 -1390
rect 2395 -1435 2400 -1395
rect 2440 -1435 2445 -1395
rect 2395 -1740 2445 -1435
rect 2745 -1395 2795 -1390
rect 2745 -1435 2750 -1395
rect 2790 -1435 2795 -1395
rect 2745 -1740 2795 -1435
rect 3095 -1395 3145 -1390
rect 3095 -1435 3100 -1395
rect 3140 -1435 3145 -1395
rect 3095 -1740 3145 -1435
rect 3445 -1395 4895 -1390
rect 3445 -1435 3450 -1395
rect 3490 -1435 3800 -1395
rect 3840 -1435 4150 -1395
rect 4190 -1435 4500 -1395
rect 4540 -1435 4850 -1395
rect 4890 -1435 4895 -1395
rect 3445 -1440 4895 -1435
rect 4145 -1740 4195 -1440
rect 995 -1745 4895 -1740
rect 995 -1785 1000 -1745
rect 1040 -1785 1350 -1745
rect 1390 -1785 1700 -1745
rect 1740 -1785 2050 -1745
rect 2090 -1785 2400 -1745
rect 2440 -1785 2750 -1745
rect 2790 -1785 3100 -1745
rect 3140 -1785 3450 -1745
rect 3490 -1785 3800 -1745
rect 3840 -1785 4150 -1745
rect 4190 -1785 4500 -1745
rect 4540 -1785 4850 -1745
rect 4890 -1785 4895 -1745
rect 995 -1790 4895 -1785
rect 995 -2095 1045 -1790
rect 995 -2135 1000 -2095
rect 1040 -2135 1045 -2095
rect 995 -2140 1045 -2135
rect 1345 -2095 1395 -1790
rect 1345 -2135 1350 -2095
rect 1390 -2135 1395 -2095
rect 1345 -2140 1395 -2135
rect 1695 -2095 1745 -1790
rect 1695 -2135 1700 -2095
rect 1740 -2135 1745 -2095
rect 1695 -2140 1745 -2135
rect 2045 -2095 2095 -1790
rect 2045 -2135 2050 -2095
rect 2090 -2135 2095 -2095
rect 2045 -2140 2095 -2135
rect 2395 -2095 2445 -1790
rect 2395 -2135 2400 -2095
rect 2440 -2135 2445 -2095
rect 2395 -2140 2445 -2135
rect 2745 -2095 2795 -1790
rect 2745 -2135 2750 -2095
rect 2790 -2135 2795 -2095
rect 2745 -2140 2795 -2135
rect 3095 -2095 3145 -1790
rect 3095 -2135 3100 -2095
rect 3140 -2135 3145 -2095
rect 3095 -2140 3145 -2135
rect 3445 -2095 3495 -1790
rect 3445 -2135 3450 -2095
rect 3490 -2135 3495 -2095
rect 3445 -2140 3495 -2135
rect 3795 -2095 3845 -1790
rect 3795 -2135 3800 -2095
rect 3840 -2135 3845 -2095
rect 3795 -2140 3845 -2135
rect 4145 -2090 4195 -1790
rect 4145 -2095 4895 -2090
rect 4145 -2135 4150 -2095
rect 4190 -2135 4500 -2095
rect 4540 -2135 4850 -2095
rect 4890 -2135 4895 -2095
rect 4145 -2140 4895 -2135
rect -3850 -2420 5140 -2415
rect -3850 -2460 825 -2420
rect 865 -2460 5140 -2420
rect -3850 -2465 5140 -2460
<< labels >>
flabel metal1 3210 -335 3210 -335 5 FreeSans 240 0 0 -80 VOUT-
port 9 s
flabel metal1 2860 400 2860 400 1 FreeSans 240 0 0 80 V_CMFB_S1
port 2 n
flabel metal1 2815 290 2815 290 1 FreeSans 240 0 0 80 V_CMFB_S2
port 7 n
flabel metal3 3100 1595 3100 1595 7 FreeSans 240 0 -80 0 cap_res_X
flabel metal1 1960 305 1960 305 5 FreeSans 240 0 0 -80 X
flabel metal1 1890 2135 1890 2135 3 FreeSans 240 0 80 0 VD3
flabel metal2 845 655 845 655 1 FreeSans 240 0 0 80 Vb1
port 6 n
flabel metal1 -1520 -335 -1520 -335 5 FreeSans 240 0 0 -80 VOUT+
port 10 s
flabel metal1 -1170 400 -1170 400 1 FreeSans 240 0 0 80 V_CMFB_S3
port 3 n
flabel metal1 -1125 290 -1125 290 1 FreeSans 240 0 0 80 V_CMFB_S4
port 8 n
flabel metal3 -1410 1610 -1410 1610 3 FreeSans 240 0 80 0 cap_res_Y
flabel metal1 -200 2135 -200 2135 7 FreeSans 240 0 -80 0 VD4
flabel metal1 1170 -280 1170 -280 3 FreeSans 240 0 80 0 V_source
flabel metal2 1550 -245 1550 -245 1 FreeSans 240 0 0 80 V_b_2nd_stage
flabel metal4 -3850 4260 -3850 4260 7 FreeSans 240 0 -80 0 VDDA
port 1 w
flabel metal4 -3850 -2440 -3850 -2440 7 FreeSans 240 0 -80 0 GNDA
port 16 w
flabel metal1 2415 1610 2415 1610 3 FreeSans 240 0 80 0 Vb3
port 4 e
flabel metal1 320 1655 320 1655 7 FreeSans 240 0 -80 0 Vb2
port 5 w
flabel metal2 1310 2775 1310 2775 1 FreeSans 240 0 0 80 Vb2_Vb3
flabel metal2 400 2775 400 2775 1 FreeSans 240 0 0 80 Vb2_2
flabel metal1 1175 1300 1175 1300 3 FreeSans 240 0 80 0 V_err_p
flabel metal1 605 1295 605 1295 3 FreeSans 240 0 80 0 V_err_mir_p
flabel metal2 -90 1120 -90 1120 7 FreeSans 240 0 -80 0 V_err_amp_ref
port 12 w
flabel metal1 890 1315 890 1315 7 FreeSans 240 0 -80 0 V_err_gate
port 13 w
flabel metal2 805 1250 805 1250 1 FreeSans 240 0 0 80 V_tot
flabel metal1 1530 1060 1530 1060 3 FreeSans 240 0 80 0 err_amp_mir
flabel metal1 1180 995 1180 995 5 FreeSans 240 0 0 -80 err_amp_out
flabel metal1 -270 305 -270 305 5 FreeSans 240 0 0 -80 Y
flabel metal1 865 -310 865 -310 3 FreeSans 240 0 80 0 V_p_mir
flabel metal2 1715 165 1715 165 3 FreeSans 240 0 80 0 VIN-
flabel metal2 -25 165 -25 165 7 FreeSans 240 0 -80 0 VIN+
flabel metal1 905 245 905 245 7 FreeSans 240 0 -80 0 V_tail_gate
flabel metal1 1375 295 1375 295 3 FreeSans 240 0 80 0 VD1
flabel metal1 315 300 315 300 7 FreeSans 240 0 -80 0 VD2
<< end >>
