* PEX produced on Wed Jul 16 10:17:22 AM CEST 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from bgr_9.ext - technology: sky130A

.subckt bgr_9 VDDA ERR_AMP_REF V_CMFB_S3 VB1_CUR_BIAS TAIL_CUR_MIR_BIAS V_CMFB_S1
+ ERR_AMP_CUR_BIAS VB3_CUR_BIAS V_CMFB_S4 V_CMFB_S2 VB2_CUR_BIAS GNDA
X0 1st_Vout_2.t11 cap_res2.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X1 TAIL_CUR_MIR_BIAS.t3 PFET_GATE_10uA.t10 VDDA.t114 VDDA.t113 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X2 GNDA.t79 NFET_GATE_10uA.t5 V_CMFB_S2.t1 GNDA.t78 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X3 VB1_CUR_BIAS.t0 PFET_GATE_10uA.t11 VDDA.t112 VDDA.t111 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X4 V_mir2.t14 V_mir2.t13 VDDA.t193 VDDA.t192 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X5 VB2_CUR_BIAS.t5 NFET_GATE_10uA.t6 GNDA.t77 GNDA.t76 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X6 a_38570_n6504.t1 a_38690_n7778.t1 GNDA.t28 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X7 GNDA.t112 GNDA.t110 V_CMFB_S2.t0 GNDA.t111 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X8 1st_Vout_1.t11 cap_res1.t20 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X9 GNDA.t75 NFET_GATE_10uA.t7 V_CMFB_S4.t2 GNDA.t74 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X10 V_p_1.t8 Vin+.t6 1st_Vout_1.t1 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X11 VB2_CUR_BIAS.t4 NFET_GATE_10uA.t8 GNDA.t73 GNDA.t72 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X12 V_p_2.t6 ERR_AMP_REF.t7 V_mir2.t16 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X13 1st_Vout_1.t12 cap_res1.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X14 GNDA.t6 START_UP_NFET1.t0 START_UP_NFET1.t1 GNDA.t5 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=10
X15 VDDA.t170 VDDA.t168 V_CMFB_S1.t5 VDDA.t169 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X16 V_TOP.t2 START_UP.t6 Vin-.t4 VDDA.t57 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X17 V_CMFB_S3.t5 VDDA.t165 VDDA.t167 VDDA.t166 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X18 GNDA.t71 NFET_GATE_10uA.t9 VB3_CUR_BIAS.t4 GNDA.t70 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X19 VB3_CUR_BIAS.t3 NFET_GATE_10uA.t10 GNDA.t69 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X20 NFET_GATE_10uA.t0 GNDA.t107 GNDA.t109 GNDA.t108 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X21 1st_Vout_1.t13 cap_res1.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X22 GNDA.t67 NFET_GATE_10uA.t3 NFET_GATE_10uA.t4 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X23 1st_Vout_2.t10 V_mir2.t17 VDDA.t188 VDDA.t187 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X24 V_p_1.t1 Vin-.t8 V_mir1.t16 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X25 V_p_2.t10 VDDA.t212 GNDA.t39 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X26 1st_Vout_2.t12 cap_res2.t19 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X27 V_CUR_REF_REG.t0 a_32320_n7778.t0 GNDA.t10 sky130_fd_pr__res_xhigh_po_0p35 l=4
X28 VB2_CUR_BIAS.t7 GNDA.t104 GNDA.t106 GNDA.t105 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X29 1st_Vout_2.t13 cap_res2.t18 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X30 V_CUR_REF_REG.t1 PFET_GATE_10uA.t12 VDDA.t110 VDDA.t109 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X31 1st_Vout_2.t14 cap_res2.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X32 VDDA.t80 V_TOP.t14 ERR_AMP_REF.t3 VDDA.t79 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X33 1st_Vout_2.t15 cap_res2.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X34 VDDA.t108 PFET_GATE_10uA.t13 V_CMFB_S1.t3 VDDA.t107 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X35 1st_Vout_2.t16 cap_res2.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X36 VB2_CUR_BIAS.t3 NFET_GATE_10uA.t11 GNDA.t65 GNDA.t64 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X37 1st_Vout_1.t14 cap_res1.t17 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X38 1st_Vout_2.t17 cap_res2.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X39 1st_Vout_2.t18 cap_res2.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X40 1st_Vout_1.t15 cap_res1.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X41 VDDA.t34 V_mir1.t10 V_mir1.t11 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X42 Vin+.t2 V_TOP.t15 VDDA.t40 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X43 1st_Vout_1.t16 cap_res1.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X44 V_TOP.t16 VDDA.t75 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X45 V_mir1.t15 Vin-.t9 V_p_1.t0 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X46 1st_Vout_1.t17 cap_res1.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X47 1st_Vout_1.t18 cap_res1.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X48 NFET_GATE_10uA.t2 VDDA.t162 VDDA.t164 VDDA.t163 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X49 VDDA.t205 V_mir2.t11 V_mir2.t12 VDDA.t204 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X50 V_TOP.t17 VDDA.t15 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X51 ERR_AMP_REF.t5 VDDA.t159 VDDA.t161 VDDA.t160 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=1.2 ps=6.8 w=3 l=0.5
X52 V_mir1.t14 Vin-.t10 V_p_1.t3 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X53 1st_Vout_1.t10 V_mir1.t17 VDDA.t210 VDDA.t209 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X54 V_TOP.t18 VDDA.t78 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X55 1st_Vout_2.t19 cap_res2.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X56 V_CMFB_S3.t3 PFET_GATE_10uA.t14 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X57 VDDA.t67 V_TOP.t19 Vin+.t3 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X58 V_TOP.t20 VDDA.t51 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 Vin+.t1 GNDA.t9 sky130_fd_pr__res_xhigh_po_0p35 l=2.3
X60 PFET_GATE_10uA.t8 1st_Vout_2.t20 VDDA.t182 VDDA.t181 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X61 1st_Vout_1.t7 Vin+.t7 V_p_1.t7 GNDA.t24 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X62 VDDA.t7 V_mir2.t18 1st_Vout_2.t3 VDDA.t6 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X63 GNDA.t103 GNDA.t101 VB3_CUR_BIAS.t5 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X64 VDDA.t180 1st_Vout_2.t21 PFET_GATE_10uA.t6 VDDA.t179 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X65 V_p_1.t6 Vin+.t8 1st_Vout_1.t5 GNDA.t16 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X66 V_CMFB_S3.t2 PFET_GATE_10uA.t15 VDDA.t104 VDDA.t103 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X67 VDDA.t158 VDDA.t156 V_TOP.t6 VDDA.t157 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X68 V_CMFB_S2.t3 NFET_GATE_10uA.t12 GNDA.t63 GNDA.t62 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X69 V_CMFB_S2.t2 NFET_GATE_10uA.t13 GNDA.t61 GNDA.t60 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X70 V_CMFB_S1.t2 PFET_GATE_10uA.t16 VDDA.t102 VDDA.t101 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X71 Vin+.t4 a_38040_n7928.t1 GNDA.t12 sky130_fd_pr__res_xhigh_po_0p35 l=6
X72 VDDA.t100 PFET_GATE_10uA.t17 TAIL_CUR_MIR_BIAS.t2 VDDA.t99 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X73 1st_Vout_1.t8 V_mir1.t18 VDDA.t184 VDDA.t183 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X74 V_mir1.t9 V_mir1.t8 VDDA.t197 VDDA.t196 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X75 V_TOP.t21 VDDA.t22 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X76 GNDA.t37 VDDA.t213 PFET_GATE_10uA.t1 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1 ps=5.8 w=2.5 l=5
X77 VDDA.t26 1st_Vout_1.t19 V_TOP.t13 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X78 PFET_GATE_10uA.t4 1st_Vout_2.t22 VDDA.t178 VDDA.t177 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X79 V_p_2.t5 ERR_AMP_REF.t8 V_mir2.t1 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.2 ps=1.8 w=0.5 l=0.2
X80 V_TOP.t7 VDDA.t214 GNDA.t36 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=1 pd=5.8 as=1.01 ps=6.15 w=2.5 l=5
X81 V_TOP.t22 VDDA.t41 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X82 VB3_CUR_BIAS.t2 NFET_GATE_10uA.t14 GNDA.t59 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X83 GNDA.t57 NFET_GATE_10uA.t15 ERR_AMP_CUR_BIAS.t1 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X84 VDDA.t36 V_mir1.t19 1st_Vout_1.t4 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X85 V_p_1.t5 Vin+.t9 1st_Vout_1.t6 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X86 1st_Vout_2.t23 cap_res2.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X87 1st_Vout_2.t24 cap_res2.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X88 V_CMFB_S1.t4 VDDA.t153 VDDA.t155 VDDA.t154 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X89 VDDA.t9 V_mir2.t19 1st_Vout_2.t4 VDDA.t8 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X90 1st_Vout_2.t25 cap_res2.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X91 VDDA.t176 1st_Vout_2.t26 PFET_GATE_10uA.t9 VDDA.t175 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X92 V_p_2.t7 V_CUR_REF_REG.t3 1st_Vout_2.t7 GNDA.t26 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X93 VDDA.t98 PFET_GATE_10uA.t18 TAIL_CUR_MIR_BIAS.t1 VDDA.t97 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X94 1st_Vout_1.t20 cap_res1.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X95 VDDA.t152 VDDA.t149 VDDA.t151 VDDA.t150 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.15
X96 V_TOP.t5 VDDA.t146 VDDA.t148 VDDA.t147 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X97 1st_Vout_2.t27 cap_res2.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X98 VDDA.t145 VDDA.t143 VB1_CUR_BIAS.t1 VDDA.t144 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X99 1st_Vout_1.t21 cap_res1.t11 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X100 V_TOP.t23 VDDA.t30 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X101 V_CMFB_S4.t1 NFET_GATE_10uA.t16 GNDA.t55 GNDA.t54 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X102 V_mir2.t10 V_mir2.t9 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X103 1st_Vout_1.t22 cap_res1.t10 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X104 GNDA.t53 NFET_GATE_10uA.t17 V_CMFB_S4.t0 GNDA.t52 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X105 1st_Vout_2.t5 V_mir2.t20 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X106 1st_Vout_1.t23 cap_res1.t9 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X107 GNDA.t85 GNDA.t98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X108 V_TOP.t24 VDDA.t27 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X109 1st_Vout_2.t28 cap_res2.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X110 Vin-.t0 a_32970_n7928.t0 GNDA.t4 sky130_fd_pr__res_xhigh_po_0p35 l=6
X111 GNDA.t85 GNDA.t99 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X112 VDDA.t142 VDDA.t140 V_TOP.t4 VDDA.t141 sky130_fd_pr__pfet_01v8 ad=0.45 pd=2.9 as=0.2 ps=1.4 w=1 l=0.15
X113 VDDA.t208 V_TOP.t25 Vin-.t6 VDDA.t207 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X114 V_TOP.t26 VDDA.t16 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X115 VDDA.t139 VDDA.t136 VDDA.t138 VDDA.t137 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0 ps=0 w=2 l=0.15
X116 a_32440_n6570.t1 a_32320_n7778.t1 GNDA.t30 sky130_fd_pr__res_xhigh_po_0p35 l=4
X117 GNDA.t85 GNDA.t100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X118 ERR_AMP_REF.t6 V_TOP.t27 VDDA.t195 VDDA.t194 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X119 VDDA.t5 V_mir1.t20 1st_Vout_1.t0 VDDA.t4 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X120 1st_Vout_2.t9 V_CUR_REF_REG.t4 V_p_2.t9 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X121 VDDA.t84 V_mir1.t6 V_mir1.t7 VDDA.t83 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X122 Vin+.t5 V_TOP.t28 VDDA.t201 VDDA.t200 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X123 V_mir1.t13 Vin-.t11 V_p_1.t10 GNDA.t35 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X124 V_TOP.t29 VDDA.t206 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X125 a_38570_n6504.t0 GNDA.t29 GNDA.t28 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X126 a_33090_n6320.t0 GNDA.t8 GNDA.t7 sky130_fd_pr__res_xhigh_po_0p35 l=6
X127 VDDA.t135 VDDA.t133 V_CUR_REF_REG.t2 VDDA.t134 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X128 V_mir1.t5 V_mir1.t4 VDDA.t43 VDDA.t42 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X129 VDDA.t132 VDDA.t130 PFET_GATE_10uA.t2 VDDA.t131 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.2
X130 GNDA.t34 VDDA.t215 V_p_1.t9 GNDA.t33 sky130_fd_pr__nfet_01v8 ad=1.01 pd=6.15 as=1 ps=5.8 w=2.5 l=5
X131 V_CMFB_S1.t1 PFET_GATE_10uA.t19 VDDA.t96 VDDA.t95 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X132 Vin-.t5 START_UP.t7 V_TOP.t1 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X133 V_TOP.t12 1st_Vout_1.t24 VDDA.t199 VDDA.t198 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X134 V_mir2.t15 ERR_AMP_REF.t9 V_p_2.t4 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X135 Vin-.t2 V_TOP.t30 VDDA.t45 VDDA.t44 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X136 a_37920_n6320.t1 GNDA.t82 GNDA.t12 sky130_fd_pr__res_xhigh_po_0p35 l=6
X137 V_mir2.t8 V_mir2.t7 VDDA.t190 VDDA.t189 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X138 PFET_GATE_10uA.t0 cap_res2.t0 GNDA.t22 sky130_fd_pr__res_high_po_0p35 l=2.05
X139 VDDA.t50 V_TOP.t31 START_UP.t0 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X140 1st_Vout_2.t6 V_mir2.t21 VDDA.t54 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X141 V_TOP.t32 VDDA.t191 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X142 VDDA.t174 1st_Vout_2.t29 PFET_GATE_10uA.t5 VDDA.t173 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X143 V_TOP.t0 cap_res1.t0 GNDA.t3 sky130_fd_pr__res_high_po_0p35 l=2.05
X144 V_TOP.t33 VDDA.t14 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X145 VDDA.t3 V_TOP.t34 ERR_AMP_REF.t0 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X146 VDDA.t47 V_mir2.t5 V_mir2.t6 VDDA.t46 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X147 VDDA.t94 PFET_GATE_10uA.t20 NFET_GATE_10uA.t1 VDDA.t93 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X148 V_TOP.t35 VDDA.t13 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X149 1st_Vout_2.t30 cap_res2.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X150 GNDA.t51 NFET_GATE_10uA.t18 VB2_CUR_BIAS.t2 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X151 V_TOP.t36 VDDA.t21 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X152 VDDA.t61 V_TOP.t37 START_UP.t2 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X153 GNDA.t97 GNDA.t95 VB2_CUR_BIAS.t6 GNDA.t96 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X154 VDDA.t129 VDDA.t127 V_CMFB_S3.t4 VDDA.t128 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X155 START_UP_NFET1.t1 START_UP.t4 START_UP.t5 GNDA.t18 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=10
X156 1st_Vout_1.t25 cap_res1.t8 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X157 PFET_GATE_10uA.t3 VDDA.t124 VDDA.t126 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.2
X158 1st_Vout_2.t31 cap_res2.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X159 V_p_1.t2 Vin-.t12 V_mir1.t12 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X160 V_p_2.t1 V_CUR_REF_REG.t5 1st_Vout_2.t2 GNDA.t1 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X161 START_UP.t1 V_TOP.t38 VDDA.t56 VDDA.t55 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X162 1st_Vout_1.t26 cap_res1.t7 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X163 V_TOP.t39 VDDA.t74 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X164 VB3_CUR_BIAS.t1 NFET_GATE_10uA.t19 GNDA.t49 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X165 1st_Vout_1.t27 cap_res1.t6 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X166 GNDA.t47 NFET_GATE_10uA.t20 VB3_CUR_BIAS.t0 GNDA.t46 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X167 ERR_AMP_CUR_BIAS.t0 NFET_GATE_10uA.t21 GNDA.t45 GNDA.t44 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X168 ERR_AMP_REF.t2 V_TOP.t40 VDDA.t77 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X169 V_TOP.t11 1st_Vout_1.t28 VDDA.t186 VDDA.t185 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X170 V_p_2.t3 ERR_AMP_REF.t10 V_mir2.t0 GNDA.t14 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X171 1st_Vout_1.t29 cap_res1.t5 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X172 1st_Vout_1.t3 V_mir1.t21 VDDA.t32 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X173 ERR_AMP_REF.t1 a_38690_n7778.t0 GNDA.t28 sky130_fd_pr__res_xhigh_po_0p35 l=4.33
X174 START_UP.t3 V_TOP.t41 VDDA.t65 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X175 VDDA.t203 V_mir1.t2 V_mir1.t3 VDDA.t202 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X176 GNDA.t43 NFET_GATE_10uA.t22 VB2_CUR_BIAS.t1 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X177 GNDA.t85 GNDA.t93 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X178 VDDA.t92 PFET_GATE_10uA.t21 V_CMFB_S3.t1 VDDA.t91 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X179 GNDA.t85 GNDA.t94 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X180 VDDA.t11 1st_Vout_1.t30 V_TOP.t10 VDDA.t10 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X181 V_TOP.t3 VDDA.t121 VDDA.t123 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X182 VDDA.t71 V_mir2.t3 V_mir2.t4 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X183 GNDA.t41 NFET_GATE_10uA.t23 VB2_CUR_BIAS.t0 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X184 V_CMFB_S4.t3 GNDA.t90 GNDA.t92 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X185 VDDA.t73 V_TOP.t42 Vin-.t3 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X186 1st_Vout_1.t31 cap_res1.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X187 VDDA.t1 V_mir2.t22 1st_Vout_2.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X188 a_33090_n6320.t1 a_32970_n7928.t1 GNDA.t23 sky130_fd_pr__res_xhigh_po_0p35 l=6
X189 GNDA.t85 GNDA.t89 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X190 VDDA.t120 VDDA.t118 VDDA.t120 VDDA.t119 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0 ps=0 w=2 l=0.15
X191 VDDA.t18 V_TOP.t43 Vin+.t0 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X192 PFET_GATE_10uA.t7 1st_Vout_2.t32 VDDA.t172 VDDA.t171 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X193 1st_Vout_2.t33 cap_res2.t4 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X194 V_TOP.t44 VDDA.t24 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X195 VDDA.t90 PFET_GATE_10uA.t22 V_CMFB_S3.t0 VDDA.t89 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X196 1st_Vout_2.t34 cap_res2.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X197 1st_Vout_1.t9 Vin+.t10 V_p_1.t4 GNDA.t80 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X198 V_mir2.t2 ERR_AMP_REF.t11 V_p_2.t2 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X199 VDDA.t88 PFET_GATE_10uA.t23 V_CMFB_S1.t0 VDDA.t87 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.15
X200 V_TOP.t9 1st_Vout_1.t32 VDDA.t59 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X201 1st_Vout_2.t35 cap_res2.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X202 Vin-.t1 V_TOP.t45 VDDA.t38 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.6 pd=3.4 as=0.6 ps=3.4 w=3 l=0.5
X203 1st_Vout_1.t33 cap_res1.t3 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X204 TAIL_CUR_MIR_BIAS.t0 PFET_GATE_10uA.t24 VDDA.t86 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.4 ps=2.4 w=2 l=0.15
X205 GNDA.t85 GNDA.t86 Vin-.t7 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X206 1st_Vout_2.t8 V_CUR_REF_REG.t6 V_p_2.t8 GNDA.t31 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.8 as=0.1 ps=0.9 w=0.5 l=0.2
X207 1st_Vout_1.t34 cap_res1.t2 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X208 1st_Vout_1.t35 cap_res1.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X209 a_37920_n6320.t0 a_38040_n7928.t0 GNDA.t12 sky130_fd_pr__res_xhigh_po_0p35 l=6
X210 GNDA.t88 GNDA.t87 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X211 VDDA.t63 1st_Vout_1.t36 V_TOP.t8 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X212 V_TOP.t46 VDDA.t12 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X213 1st_Vout_2.t1 V_CUR_REF_REG.t7 V_p_2.t0 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.9 as=0.1 ps=0.9 w=0.5 l=0.2
X214 VDDA.t117 VDDA.t115 ERR_AMP_REF.t4 VDDA.t116 sky130_fd_pr__pfet_01v8 ad=1.2 pd=6.8 as=0.6 ps=3.4 w=3 l=0.5
X215 VDDA.t29 V_mir1.t22 1st_Vout_1.t2 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
X216 V_TOP.t47 VDDA.t23 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X217 GNDA.t85 GNDA.t84 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__pnp_05v5_W3p40L3p40
**devattr s=462400,2720
X218 V_TOP.t48 VDDA.t211 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X219 1st_Vout_2.t36 cap_res2.t1 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X220 a_32440_n6570.t0 GNDA.t21 GNDA.t20 sky130_fd_pr__res_xhigh_po_0p35 l=4
X221 V_TOP.t49 VDDA.t48 sky130_fd_pr__cap_mim_m3_1 l=2 w=2
X222 V_mir1.t1 V_mir1.t0 VDDA.t82 VDDA.t81 sky130_fd_pr__pfet_01v8 ad=0.2 pd=1.4 as=0.2 ps=1.4 w=1 l=0.2
R0 1st_Vout_2 1st_Vout_2.t29 354.854
R1 1st_Vout_2.n0 1st_Vout_2.t22 346.8
R2 1st_Vout_2 1st_Vout_2.n11 344.95
R3 1st_Vout_2.n0 1st_Vout_2.n4 344.95
R4 1st_Vout_2.n2 1st_Vout_2.n6 340.45
R5 1st_Vout_2.n8 1st_Vout_2.t8 275.909
R6 1st_Vout_2.n8 1st_Vout_2.n7 227.909
R7 1st_Vout_2.n2 1st_Vout_2.n9 222.034
R8 1st_Vout_2.n5 1st_Vout_2.t20 184.097
R9 1st_Vout_2.n5 1st_Vout_2.t26 184.097
R10 1st_Vout_2.n10 1st_Vout_2.t32 184.097
R11 1st_Vout_2.n10 1st_Vout_2.t21 184.097
R12 1st_Vout_2.n0 1st_Vout_2.n5 166.05
R13 1st_Vout_2 1st_Vout_2.n10 166.05
R14 1st_Vout_2.n0 1st_Vout_2.n3 52.9634
R15 1st_Vout_2.n9 1st_Vout_2.t7 48.0005
R16 1st_Vout_2.n9 1st_Vout_2.t1 48.0005
R17 1st_Vout_2.n7 1st_Vout_2.t2 48.0005
R18 1st_Vout_2.n7 1st_Vout_2.t9 48.0005
R19 1st_Vout_2.n6 1st_Vout_2.t4 39.4005
R20 1st_Vout_2.n6 1st_Vout_2.t5 39.4005
R21 1st_Vout_2.n11 1st_Vout_2.t3 39.4005
R22 1st_Vout_2.n11 1st_Vout_2.t10 39.4005
R23 1st_Vout_2.n4 1st_Vout_2.t0 39.4005
R24 1st_Vout_2.n4 1st_Vout_2.t6 39.4005
R25 1st_Vout_2 1st_Vout_2.n0 5.6255
R26 1st_Vout_2 1st_Vout_2.n2 5.28175
R27 1st_Vout_2.n1 1st_Vout_2.t27 4.8295
R28 1st_Vout_2.n1 1st_Vout_2.t11 4.8295
R29 1st_Vout_2.n1 1st_Vout_2.t18 4.8295
R30 1st_Vout_2.n1 1st_Vout_2.t31 4.8295
R31 1st_Vout_2.n1 1st_Vout_2.t35 4.8295
R32 1st_Vout_2.n1 1st_Vout_2.t24 4.8295
R33 1st_Vout_2.n3 1st_Vout_2.t16 4.8295
R34 1st_Vout_2.n3 1st_Vout_2.t30 4.8295
R35 1st_Vout_2.n3 1st_Vout_2.t28 4.8295
R36 1st_Vout_2.n2 1st_Vout_2.n8 4.5005
R37 1st_Vout_2.n1 1st_Vout_2.t25 4.5005
R38 1st_Vout_2.n1 1st_Vout_2.t23 4.5005
R39 1st_Vout_2.n1 1st_Vout_2.t17 4.5005
R40 1st_Vout_2.n1 1st_Vout_2.t15 4.5005
R41 1st_Vout_2.n1 1st_Vout_2.t34 4.5005
R42 1st_Vout_2.n1 1st_Vout_2.t33 4.5005
R43 1st_Vout_2.n3 1st_Vout_2.t13 4.5005
R44 1st_Vout_2.n3 1st_Vout_2.t12 4.5005
R45 1st_Vout_2.n3 1st_Vout_2.t19 4.5005
R46 1st_Vout_2.n3 1st_Vout_2.t36 4.5005
R47 1st_Vout_2.n3 1st_Vout_2.t14 4.5005
R48 1st_Vout_2.n3 1st_Vout_2.n1 3.1025
R49 cap_res2 cap_res2.t0 121.05
R50 cap_res2 cap_res2.t12 0.194375
R51 cap_res2.t1 cap_res2.t17 0.1603
R52 cap_res2.t19 cap_res2.t6 0.1603
R53 cap_res2.t4 cap_res2.t10 0.1603
R54 cap_res2.t16 cap_res2.t5 0.1603
R55 cap_res2.t11 cap_res2.t20 0.1603
R56 cap_res2.n1 cap_res2.t9 0.159278
R57 cap_res2.n2 cap_res2.t14 0.159278
R58 cap_res2.n3 cap_res2.t3 0.159278
R59 cap_res2.n4 cap_res2.t18 0.159278
R60 cap_res2.n4 cap_res2.t1 0.1368
R61 cap_res2.n4 cap_res2.t7 0.1368
R62 cap_res2.n3 cap_res2.t19 0.1368
R63 cap_res2.n3 cap_res2.t15 0.1368
R64 cap_res2.n2 cap_res2.t4 0.1368
R65 cap_res2.n2 cap_res2.t2 0.1368
R66 cap_res2.n1 cap_res2.t16 0.1368
R67 cap_res2.n1 cap_res2.t13 0.1368
R68 cap_res2.n0 cap_res2.t11 0.1368
R69 cap_res2.n0 cap_res2.t8 0.1368
R70 cap_res2.t9 cap_res2.n0 0.00152174
R71 cap_res2.t14 cap_res2.n1 0.00152174
R72 cap_res2.t3 cap_res2.n2 0.00152174
R73 cap_res2.t18 cap_res2.n3 0.00152174
R74 cap_res2.t12 cap_res2.n4 0.00152174
R75 PFET_GATE_10uA.n3 PFET_GATE_10uA.t11 565.114
R76 PFET_GATE_10uA.n19 PFET_GATE_10uA.t10 530.201
R77 PFET_GATE_10uA.n21 PFET_GATE_10uA.t17 409.7
R78 PFET_GATE_10uA.n16 PFET_GATE_10uA.t23 369.534
R79 PFET_GATE_10uA.n15 PFET_GATE_10uA.t19 369.534
R80 PFET_GATE_10uA.n1 PFET_GATE_10uA.t22 369.534
R81 PFET_GATE_10uA.n0 PFET_GATE_10uA.t14 369.534
R82 PFET_GATE_10uA.n19 PFET_GATE_10uA.t18 353.467
R83 PFET_GATE_10uA.n20 PFET_GATE_10uA.t24 353.467
R84 PFET_GATE_10uA.n6 PFET_GATE_10uA.n4 346.825
R85 PFET_GATE_10uA.n8 PFET_GATE_10uA.n7 344.7
R86 PFET_GATE_10uA.n6 PFET_GATE_10uA.n5 344.7
R87 PFET_GATE_10uA.n11 PFET_GATE_10uA.n10 340.2
R88 PFET_GATE_10uA.n14 PFET_GATE_10uA.t20 325.351
R89 PFET_GATE_10uA.n18 PFET_GATE_10uA.n14 202.364
R90 PFET_GATE_10uA.n16 PFET_GATE_10uA.t16 192.8
R91 PFET_GATE_10uA.n15 PFET_GATE_10uA.t13 192.8
R92 PFET_GATE_10uA.n14 PFET_GATE_10uA.t12 192.8
R93 PFET_GATE_10uA.n1 PFET_GATE_10uA.t15 192.8
R94 PFET_GATE_10uA.n0 PFET_GATE_10uA.t21 192.8
R95 PFET_GATE_10uA.n20 PFET_GATE_10uA.n19 176.733
R96 PFET_GATE_10uA.n13 PFET_GATE_10uA.n2 168.166
R97 PFET_GATE_10uA PFET_GATE_10uA.n21 166.071
R98 PFET_GATE_10uA.n18 PFET_GATE_10uA.n17 166.071
R99 PFET_GATE_10uA.n3 PFET_GATE_10uA.t0 137.386
R100 PFET_GATE_10uA.n9 PFET_GATE_10uA.t1 116.584
R101 PFET_GATE_10uA.n21 PFET_GATE_10uA.n20 56.2338
R102 PFET_GATE_10uA.n17 PFET_GATE_10uA.n16 56.2338
R103 PFET_GATE_10uA.n17 PFET_GATE_10uA.n15 56.2338
R104 PFET_GATE_10uA.n2 PFET_GATE_10uA.n1 56.2338
R105 PFET_GATE_10uA.n2 PFET_GATE_10uA.n0 56.2338
R106 PFET_GATE_10uA.n10 PFET_GATE_10uA.t5 39.4005
R107 PFET_GATE_10uA.n10 PFET_GATE_10uA.t3 39.4005
R108 PFET_GATE_10uA.n7 PFET_GATE_10uA.t6 39.4005
R109 PFET_GATE_10uA.n7 PFET_GATE_10uA.t7 39.4005
R110 PFET_GATE_10uA.n5 PFET_GATE_10uA.t9 39.4005
R111 PFET_GATE_10uA.n5 PFET_GATE_10uA.t8 39.4005
R112 PFET_GATE_10uA.n4 PFET_GATE_10uA.t2 39.4005
R113 PFET_GATE_10uA.n4 PFET_GATE_10uA.t4 39.4005
R114 PFET_GATE_10uA.n13 PFET_GATE_10uA.n12 27.5005
R115 PFET_GATE_10uA.n12 PFET_GATE_10uA.n11 9.53175
R116 PFET_GATE_10uA PFET_GATE_10uA.n18 5.2505
R117 PFET_GATE_10uA.n11 PFET_GATE_10uA.n9 4.5005
R118 PFET_GATE_10uA PFET_GATE_10uA.n13 2.34425
R119 PFET_GATE_10uA.n8 PFET_GATE_10uA.n6 2.1255
R120 PFET_GATE_10uA.n9 PFET_GATE_10uA.n8 2.1255
R121 PFET_GATE_10uA.n12 PFET_GATE_10uA.n3 1.78175
R122 VDDA.n102 VDDA.t141 683.365
R123 VDDA.n94 VDDA.t131 660
R124 VDDA.t125 VDDA.n93 660
R125 VDDA.n88 VDDA.t157 660
R126 VDDA.t147 VDDA.n87 660
R127 VDDA.n36 VDDA.t128 643.037
R128 VDDA.t166 VDDA.n35 643.037
R129 VDDA.n24 VDDA.t169 643.037
R130 VDDA.t154 VDDA.n23 643.037
R131 VDDA.n18 VDDA.t134 643.037
R132 VDDA.t163 VDDA.n17 643.037
R133 VDDA.t122 VDDA.n101 643.037
R134 VDDA.n126 VDDA.t149 611.909
R135 VDDA.n28 VDDA.t136 601.867
R136 VDDA.n31 VDDA.t118 601.867
R137 VDDA.n123 VDDA.t143 579.775
R138 VDDA.n100 VDDA.t121 413.084
R139 VDDA.n103 VDDA.t140 413.084
R140 VDDA.n34 VDDA.t165 409.067
R141 VDDA.n37 VDDA.t127 409.067
R142 VDDA.n22 VDDA.t153 409.067
R143 VDDA.n16 VDDA.t162 409.067
R144 VDDA.n19 VDDA.t133 409.067
R145 VDDA.t131 VDDA.t177 407.144
R146 VDDA.t177 VDDA.t204 407.144
R147 VDDA.t204 VDDA.t192 407.144
R148 VDDA.t192 VDDA.t0 407.144
R149 VDDA.t0 VDDA.t53 407.144
R150 VDDA.t53 VDDA.t175 407.144
R151 VDDA.t175 VDDA.t181 407.144
R152 VDDA.t181 VDDA.t70 407.144
R153 VDDA.t70 VDDA.t189 407.144
R154 VDDA.t189 VDDA.t8 407.144
R155 VDDA.t8 VDDA.t19 407.144
R156 VDDA.t19 VDDA.t179 407.144
R157 VDDA.t179 VDDA.t171 407.144
R158 VDDA.t171 VDDA.t46 407.144
R159 VDDA.t46 VDDA.t68 407.144
R160 VDDA.t68 VDDA.t6 407.144
R161 VDDA.t6 VDDA.t187 407.144
R162 VDDA.t187 VDDA.t173 407.144
R163 VDDA.t173 VDDA.t125 407.144
R164 VDDA.t157 VDDA.t58 407.144
R165 VDDA.t58 VDDA.t28 407.144
R166 VDDA.t28 VDDA.t31 407.144
R167 VDDA.t31 VDDA.t83 407.144
R168 VDDA.t83 VDDA.t196 407.144
R169 VDDA.t196 VDDA.t62 407.144
R170 VDDA.t62 VDDA.t185 407.144
R171 VDDA.t185 VDDA.t4 407.144
R172 VDDA.t4 VDDA.t183 407.144
R173 VDDA.t183 VDDA.t33 407.144
R174 VDDA.t33 VDDA.t81 407.144
R175 VDDA.t81 VDDA.t10 407.144
R176 VDDA.t10 VDDA.t198 407.144
R177 VDDA.t198 VDDA.t35 407.144
R178 VDDA.t35 VDDA.t209 407.144
R179 VDDA.t209 VDDA.t202 407.144
R180 VDDA.t202 VDDA.t42 407.144
R181 VDDA.t42 VDDA.t25 407.144
R182 VDDA.t25 VDDA.t147 407.144
R183 VDDA.n25 VDDA.t168 390.322
R184 VDDA.t128 VDDA.t105 373.214
R185 VDDA.t105 VDDA.t91 373.214
R186 VDDA.t91 VDDA.t103 373.214
R187 VDDA.t103 VDDA.t89 373.214
R188 VDDA.t89 VDDA.t166 373.214
R189 VDDA.t169 VDDA.t95 373.214
R190 VDDA.t95 VDDA.t107 373.214
R191 VDDA.t107 VDDA.t101 373.214
R192 VDDA.t101 VDDA.t87 373.214
R193 VDDA.t87 VDDA.t154 373.214
R194 VDDA.t134 VDDA.t109 373.214
R195 VDDA.t109 VDDA.t93 373.214
R196 VDDA.t93 VDDA.t163 373.214
R197 VDDA.t141 VDDA.t57 373.214
R198 VDDA.t57 VDDA.t52 373.214
R199 VDDA.t52 VDDA.t122 373.214
R200 VDDA.n122 VDDA.t115 360.868
R201 VDDA.n105 VDDA.t159 360.868
R202 VDDA.n89 VDDA.t156 358.858
R203 VDDA.n51 VDDA.n50 347.104
R204 VDDA.n53 VDDA.n52 347.104
R205 VDDA.n55 VDDA.n54 347.104
R206 VDDA.n57 VDDA.n56 347.104
R207 VDDA.n59 VDDA.n58 347.104
R208 VDDA.n61 VDDA.n60 347.104
R209 VDDA.n63 VDDA.n62 347.104
R210 VDDA.n65 VDDA.n64 347.104
R211 VDDA.n67 VDDA.n66 347.104
R212 VDDA.n69 VDDA.n68 347.104
R213 VDDA.n71 VDDA.n70 347.104
R214 VDDA.n73 VDDA.n72 347.104
R215 VDDA.n75 VDDA.n74 347.104
R216 VDDA.n77 VDDA.n76 347.104
R217 VDDA.n79 VDDA.n78 347.104
R218 VDDA.n81 VDDA.n80 347.104
R219 VDDA.n83 VDDA.n82 347.104
R220 VDDA.n85 VDDA.n84 347.104
R221 VDDA.n11 VDDA.n10 345.127
R222 VDDA.n13 VDDA.n12 345.127
R223 VDDA.n15 VDDA.n14 345.127
R224 VDDA.n1 VDDA.n0 344.7
R225 VDDA.n3 VDDA.n2 344.7
R226 VDDA.n30 VDDA.t119 341.188
R227 VDDA.t137 VDDA.n29 341.188
R228 VDDA.t144 VDDA.n124 341.188
R229 VDDA.n125 VDDA.t150 341.188
R230 VDDA.n24 VDDA.t170 332.267
R231 VDDA.n23 VDDA.t155 332.267
R232 VDDA.n18 VDDA.t135 332.267
R233 VDDA.n17 VDDA.t164 332.267
R234 VDDA.n36 VDDA.t129 332.084
R235 VDDA.n35 VDDA.t167 332.084
R236 VDDA.n102 VDDA.t142 331.901
R237 VDDA.n101 VDDA.t123 331.901
R238 VDDA.n94 VDDA.t132 331.901
R239 VDDA.n93 VDDA.t126 331.901
R240 VDDA.n88 VDDA.t158 331.901
R241 VDDA.n87 VDDA.t148 331.901
R242 VDDA.t116 VDDA.n98 280.798
R243 VDDA.n99 VDDA.t160 280.798
R244 VDDA.t194 VDDA.t116 240.845
R245 VDDA.t49 VDDA.t194 240.845
R246 VDDA.t55 VDDA.t49 240.845
R247 VDDA.t72 VDDA.t55 240.845
R248 VDDA.t37 VDDA.t72 240.845
R249 VDDA.t66 VDDA.t37 240.845
R250 VDDA.t200 VDDA.t66 240.845
R251 VDDA.t2 VDDA.t200 240.845
R252 VDDA.t76 VDDA.t2 240.845
R253 VDDA.t17 VDDA.t76 240.845
R254 VDDA.t39 VDDA.t17 240.845
R255 VDDA.t207 VDDA.t39 240.845
R256 VDDA.t44 VDDA.t207 240.845
R257 VDDA.t60 VDDA.t44 240.845
R258 VDDA.t64 VDDA.t60 240.845
R259 VDDA.t79 VDDA.t64 240.845
R260 VDDA.t160 VDDA.t79 240.845
R261 VDDA.t119 VDDA.t99 217.708
R262 VDDA.t99 VDDA.t85 217.708
R263 VDDA.t85 VDDA.t97 217.708
R264 VDDA.t97 VDDA.t113 217.708
R265 VDDA.t113 VDDA.t137 217.708
R266 VDDA.t111 VDDA.t144 217.708
R267 VDDA.t150 VDDA.t111 217.708
R268 VDDA.n5 VDDA.n4 190.534
R269 VDDA.n7 VDDA.n6 190.534
R270 VDDA.n9 VDDA.n8 190.534
R271 VDDA.n129 VDDA.n128 186.034
R272 VDDA.n92 VDDA.t124 179.43
R273 VDDA.n86 VDDA.t146 179.43
R274 VDDA.n95 VDDA.t130 179.358
R275 VDDA.n46 VDDA.t215 169.55
R276 VDDA.n48 VDDA.t212 165.8
R277 VDDA.n47 VDDA.t213 165.8
R278 VDDA.n46 VDDA.t214 165.8
R279 VDDA.n107 VDDA.n106 147.792
R280 VDDA.n109 VDDA.n108 147.792
R281 VDDA.n111 VDDA.n110 147.792
R282 VDDA.n113 VDDA.n112 147.792
R283 VDDA.n115 VDDA.n114 147.792
R284 VDDA.n117 VDDA.n116 147.792
R285 VDDA.n119 VDDA.n118 147.792
R286 VDDA.n121 VDDA.n120 147.792
R287 VDDA.n30 VDDA.t120 136.701
R288 VDDA.n29 VDDA.t139 136.701
R289 VDDA.n124 VDDA.t145 136.701
R290 VDDA.n125 VDDA.t152 136.701
R291 VDDA.n107 VDDA.n105 99.2005
R292 VDDA.n122 VDDA.n121 99.2005
R293 VDDA.n109 VDDA.n107 96.0005
R294 VDDA.n111 VDDA.n109 96.0005
R295 VDDA.n113 VDDA.n111 96.0005
R296 VDDA.n115 VDDA.n113 96.0005
R297 VDDA.n117 VDDA.n115 96.0005
R298 VDDA.n119 VDDA.n117 96.0005
R299 VDDA.n121 VDDA.n119 96.0005
R300 VDDA.n98 VDDA.t117 86.2588
R301 VDDA.n99 VDDA.t161 86.2588
R302 VDDA.n0 VDDA.t106 39.4005
R303 VDDA.n0 VDDA.t92 39.4005
R304 VDDA.n2 VDDA.t104 39.4005
R305 VDDA.n2 VDDA.t90 39.4005
R306 VDDA.n10 VDDA.t96 39.4005
R307 VDDA.n10 VDDA.t108 39.4005
R308 VDDA.n12 VDDA.t102 39.4005
R309 VDDA.n12 VDDA.t88 39.4005
R310 VDDA.n14 VDDA.t110 39.4005
R311 VDDA.n14 VDDA.t94 39.4005
R312 VDDA.n50 VDDA.t178 39.4005
R313 VDDA.n50 VDDA.t205 39.4005
R314 VDDA.n52 VDDA.t193 39.4005
R315 VDDA.n52 VDDA.t1 39.4005
R316 VDDA.n54 VDDA.t54 39.4005
R317 VDDA.n54 VDDA.t176 39.4005
R318 VDDA.n56 VDDA.t182 39.4005
R319 VDDA.n56 VDDA.t71 39.4005
R320 VDDA.n58 VDDA.t190 39.4005
R321 VDDA.n58 VDDA.t9 39.4005
R322 VDDA.n60 VDDA.t20 39.4005
R323 VDDA.n60 VDDA.t180 39.4005
R324 VDDA.n62 VDDA.t172 39.4005
R325 VDDA.n62 VDDA.t47 39.4005
R326 VDDA.n64 VDDA.t69 39.4005
R327 VDDA.n64 VDDA.t7 39.4005
R328 VDDA.n66 VDDA.t188 39.4005
R329 VDDA.n66 VDDA.t174 39.4005
R330 VDDA.n68 VDDA.t59 39.4005
R331 VDDA.n68 VDDA.t29 39.4005
R332 VDDA.n70 VDDA.t32 39.4005
R333 VDDA.n70 VDDA.t84 39.4005
R334 VDDA.n72 VDDA.t197 39.4005
R335 VDDA.n72 VDDA.t63 39.4005
R336 VDDA.n74 VDDA.t186 39.4005
R337 VDDA.n74 VDDA.t5 39.4005
R338 VDDA.n76 VDDA.t184 39.4005
R339 VDDA.n76 VDDA.t34 39.4005
R340 VDDA.n78 VDDA.t82 39.4005
R341 VDDA.n78 VDDA.t11 39.4005
R342 VDDA.n80 VDDA.t199 39.4005
R343 VDDA.n80 VDDA.t36 39.4005
R344 VDDA.n82 VDDA.t210 39.4005
R345 VDDA.n82 VDDA.t203 39.4005
R346 VDDA.n84 VDDA.t43 39.4005
R347 VDDA.n84 VDDA.t26 39.4005
R348 VDDA.n31 VDDA.n30 36.5719
R349 VDDA.n29 VDDA.n28 36.5719
R350 VDDA.n126 VDDA.n125 36.5719
R351 VDDA.n124 VDDA.n123 36.5719
R352 VDDA.n122 VDDA.n98 35.0481
R353 VDDA.n105 VDDA.n99 35.0481
R354 VDDA.n45 VDDA.n39 33.7847
R355 VDDA.n37 VDDA.n36 27.2462
R356 VDDA.n35 VDDA.n34 27.2462
R357 VDDA.n25 VDDA.n24 27.2462
R358 VDDA.n23 VDDA.n22 27.2462
R359 VDDA.n19 VDDA.n18 27.2462
R360 VDDA.n17 VDDA.n16 27.2462
R361 VDDA.n86 VDDA.n85 26.5117
R362 VDDA.n96 VDDA.n95 25.8913
R363 VDDA.n92 VDDA.n91 25.8867
R364 VDDA.n101 VDDA.n100 25.2957
R365 VDDA.n89 VDDA.n88 25.2957
R366 VDDA.n45 VDDA.t206 19.9244
R367 VDDA.t120 VDDA.n5 19.7005
R368 VDDA.n5 VDDA.t100 19.7005
R369 VDDA.n6 VDDA.t86 19.7005
R370 VDDA.n6 VDDA.t98 19.7005
R371 VDDA.n8 VDDA.t114 19.7005
R372 VDDA.n8 VDDA.t138 19.7005
R373 VDDA.n128 VDDA.t112 19.7005
R374 VDDA.n128 VDDA.t151 19.7005
R375 VDDA.n130 VDDA.n122 16.3005
R376 VDDA.n105 VDDA.n104 15.6443
R377 VDDA.n104 VDDA.n100 15.488
R378 VDDA.n103 VDDA.n102 14.9338
R379 VDDA.n127 VDDA.n123 14.363
R380 VDDA.n16 VDDA.n15 14.2693
R381 VDDA.n104 VDDA.n103 14.238
R382 VDDA.n127 VDDA.n126 14.0818
R383 VDDA.n90 VDDA.n89 14.0713
R384 VDDA.n34 VDDA.n33 13.8005
R385 VDDA.n28 VDDA.n27 13.8005
R386 VDDA.n22 VDDA.n21 13.8005
R387 VDDA.n20 VDDA.n19 13.8005
R388 VDDA.n26 VDDA.n25 13.8005
R389 VDDA.n32 VDDA.n31 13.8005
R390 VDDA.n38 VDDA.n37 13.8005
R391 VDDA.n106 VDDA.t65 13.1338
R392 VDDA.n106 VDDA.t80 13.1338
R393 VDDA.n108 VDDA.t45 13.1338
R394 VDDA.n108 VDDA.t61 13.1338
R395 VDDA.n110 VDDA.t40 13.1338
R396 VDDA.n110 VDDA.t208 13.1338
R397 VDDA.n112 VDDA.t77 13.1338
R398 VDDA.n112 VDDA.t18 13.1338
R399 VDDA.n114 VDDA.t201 13.1338
R400 VDDA.n114 VDDA.t3 13.1338
R401 VDDA.n116 VDDA.t38 13.1338
R402 VDDA.n116 VDDA.t67 13.1338
R403 VDDA.n118 VDDA.t56 13.1338
R404 VDDA.n118 VDDA.t73 13.1338
R405 VDDA.n120 VDDA.t195 13.1338
R406 VDDA.n120 VDDA.t50 13.1338
R407 VDDA.n93 VDDA.n92 12.6486
R408 VDDA.n87 VDDA.n86 12.6486
R409 VDDA.n95 VDDA.n94 12.6436
R410 VDDA.n39 VDDA.n38 11.4105
R411 VDDA.n49 VDDA.n48 11.348
R412 VDDA.n131 VDDA.n130 9.7855
R413 VDDA.n97 VDDA.n96 8.973
R414 VDDA.n130 VDDA.n129 4.7505
R415 VDDA.n49 VDDA.n45 4.5595
R416 VDDA.n129 VDDA.n127 4.5005
R417 VDDA.n47 VDDA.n46 4.3755
R418 VDDA.n48 VDDA.n47 3.7505
R419 VDDA.n27 VDDA.n26 2.78175
R420 VDDA.n33 VDDA.n32 2.78175
R421 VDDA.n21 VDDA.n20 2.063
R422 VDDA.n91 VDDA.n90 1.8755
R423 VDDA.n97 VDDA.n49 0.840625
R424 VDDA.n131 VDDA.n97 0.74075
R425 VDDA.n20 VDDA.n15 0.65675
R426 VDDA.n85 VDDA.n83 0.6255
R427 VDDA.n83 VDDA.n81 0.6255
R428 VDDA.n81 VDDA.n79 0.6255
R429 VDDA.n79 VDDA.n77 0.6255
R430 VDDA.n77 VDDA.n75 0.6255
R431 VDDA.n75 VDDA.n73 0.6255
R432 VDDA.n73 VDDA.n71 0.6255
R433 VDDA.n71 VDDA.n69 0.6255
R434 VDDA.n90 VDDA.n69 0.6255
R435 VDDA.n91 VDDA.n67 0.6255
R436 VDDA.n67 VDDA.n65 0.6255
R437 VDDA.n65 VDDA.n63 0.6255
R438 VDDA.n63 VDDA.n61 0.6255
R439 VDDA.n61 VDDA.n59 0.6255
R440 VDDA.n59 VDDA.n57 0.6255
R441 VDDA.n57 VDDA.n55 0.6255
R442 VDDA.n55 VDDA.n53 0.6255
R443 VDDA.n53 VDDA.n51 0.6255
R444 VDDA.n96 VDDA.n51 0.6255
R445 VDDA.n21 VDDA.n13 0.563
R446 VDDA.n13 VDDA.n11 0.563
R447 VDDA.n26 VDDA.n11 0.563
R448 VDDA.n9 VDDA.n7 0.563
R449 VDDA.n7 VDDA.n4 0.563
R450 VDDA.n33 VDDA.n3 0.563
R451 VDDA.n3 VDDA.n1 0.563
R452 VDDA.n38 VDDA.n1 0.563
R453 VDDA VDDA.n131 0.41175
R454 VDDA.n27 VDDA.n9 0.28175
R455 VDDA.n32 VDDA.n4 0.28175
R456 VDDA.t74 VDDA.t30 0.1603
R457 VDDA.t15 VDDA.t75 0.1603
R458 VDDA.t211 VDDA.t12 0.1603
R459 VDDA.t51 VDDA.t78 0.1603
R460 VDDA.t16 VDDA.t27 0.1603
R461 VDDA.n41 VDDA.t23 0.159278
R462 VDDA.n42 VDDA.t13 0.159278
R463 VDDA.n43 VDDA.t22 0.159278
R464 VDDA.n44 VDDA.t191 0.159278
R465 VDDA.n44 VDDA.t74 0.1368
R466 VDDA.n44 VDDA.t24 0.1368
R467 VDDA.n43 VDDA.t15 0.1368
R468 VDDA.n43 VDDA.t14 0.1368
R469 VDDA.n42 VDDA.t211 0.1368
R470 VDDA.n42 VDDA.t41 0.1368
R471 VDDA.n41 VDDA.t51 0.1368
R472 VDDA.n41 VDDA.t21 0.1368
R473 VDDA.n40 VDDA.t16 0.1368
R474 VDDA.n40 VDDA.t48 0.1368
R475 VDDA VDDA.n39 0.135625
R476 VDDA.t23 VDDA.n40 0.00152174
R477 VDDA.t13 VDDA.n41 0.00152174
R478 VDDA.t22 VDDA.n42 0.00152174
R479 VDDA.t191 VDDA.n43 0.00152174
R480 VDDA.t206 VDDA.n44 0.00152174
R481 TAIL_CUR_MIR_BIAS.n2 TAIL_CUR_MIR_BIAS.n0 264.63
R482 TAIL_CUR_MIR_BIAS.n2 TAIL_CUR_MIR_BIAS.n1 117.001
R483 TAIL_CUR_MIR_BIAS TAIL_CUR_MIR_BIAS.n2 73.188
R484 TAIL_CUR_MIR_BIAS.n1 TAIL_CUR_MIR_BIAS.t1 19.7005
R485 TAIL_CUR_MIR_BIAS.n1 TAIL_CUR_MIR_BIAS.t3 19.7005
R486 TAIL_CUR_MIR_BIAS.n0 TAIL_CUR_MIR_BIAS.t2 19.7005
R487 TAIL_CUR_MIR_BIAS.n0 TAIL_CUR_MIR_BIAS.t0 19.7005
R488 NFET_GATE_10uA.n19 NFET_GATE_10uA.n0 396.791
R489 NFET_GATE_10uA.n19 NFET_GATE_10uA.t3 384.967
R490 NFET_GATE_10uA.n10 NFET_GATE_10uA.t22 369.534
R491 NFET_GATE_10uA.n9 NFET_GATE_10uA.t13 369.534
R492 NFET_GATE_10uA.n7 NFET_GATE_10uA.t17 369.534
R493 NFET_GATE_10uA.n4 NFET_GATE_10uA.t8 369.534
R494 NFET_GATE_10uA.n1 NFET_GATE_10uA.t19 369.534
R495 NFET_GATE_10uA.t3 NFET_GATE_10uA.n18 369.534
R496 NFET_GATE_10uA.n10 NFET_GATE_10uA.t12 192.8
R497 NFET_GATE_10uA.n11 NFET_GATE_10uA.t5 192.8
R498 NFET_GATE_10uA.n12 NFET_GATE_10uA.t6 192.8
R499 NFET_GATE_10uA.n9 NFET_GATE_10uA.t18 192.8
R500 NFET_GATE_10uA.n7 NFET_GATE_10uA.t11 192.8
R501 NFET_GATE_10uA.n6 NFET_GATE_10uA.t23 192.8
R502 NFET_GATE_10uA.n5 NFET_GATE_10uA.t16 192.8
R503 NFET_GATE_10uA.n4 NFET_GATE_10uA.t7 192.8
R504 NFET_GATE_10uA.n3 NFET_GATE_10uA.t20 192.8
R505 NFET_GATE_10uA.n2 NFET_GATE_10uA.t14 192.8
R506 NFET_GATE_10uA.n1 NFET_GATE_10uA.t9 192.8
R507 NFET_GATE_10uA.n18 NFET_GATE_10uA.t21 192.8
R508 NFET_GATE_10uA.n17 NFET_GATE_10uA.t15 192.8
R509 NFET_GATE_10uA.n16 NFET_GATE_10uA.t10 192.8
R510 NFET_GATE_10uA.n12 NFET_GATE_10uA.n11 176.733
R511 NFET_GATE_10uA.n11 NFET_GATE_10uA.n10 176.733
R512 NFET_GATE_10uA.n5 NFET_GATE_10uA.n4 176.733
R513 NFET_GATE_10uA.n6 NFET_GATE_10uA.n5 176.733
R514 NFET_GATE_10uA.n2 NFET_GATE_10uA.n1 176.733
R515 NFET_GATE_10uA.n3 NFET_GATE_10uA.n2 176.733
R516 NFET_GATE_10uA.n17 NFET_GATE_10uA.n16 176.733
R517 NFET_GATE_10uA.n18 NFET_GATE_10uA.n17 176.733
R518 NFET_GATE_10uA.n14 NFET_GATE_10uA.n13 169.852
R519 NFET_GATE_10uA.n14 NFET_GATE_10uA.n8 169.852
R520 NFET_GATE_10uA.n15 NFET_GATE_10uA.n14 166.133
R521 NFET_GATE_10uA.n20 NFET_GATE_10uA.n19 132.5
R522 NFET_GATE_10uA.n13 NFET_GATE_10uA.n12 56.2338
R523 NFET_GATE_10uA.n13 NFET_GATE_10uA.n9 56.2338
R524 NFET_GATE_10uA.n8 NFET_GATE_10uA.n7 56.2338
R525 NFET_GATE_10uA.n8 NFET_GATE_10uA.n6 56.2338
R526 NFET_GATE_10uA.n15 NFET_GATE_10uA.n3 56.2338
R527 NFET_GATE_10uA.n16 NFET_GATE_10uA.n15 56.2338
R528 NFET_GATE_10uA.n0 NFET_GATE_10uA.t1 39.4005
R529 NFET_GATE_10uA.n0 NFET_GATE_10uA.t2 39.4005
R530 NFET_GATE_10uA.n20 NFET_GATE_10uA.t4 24.0005
R531 NFET_GATE_10uA.t0 NFET_GATE_10uA.n20 24.0005
R532 V_CMFB_S2.n2 V_CMFB_S2.n0 150.451
R533 V_CMFB_S2.n2 V_CMFB_S2.n1 140.201
R534 V_CMFB_S2 V_CMFB_S2.n2 37.563
R535 V_CMFB_S2.n1 V_CMFB_S2.t1 24.0005
R536 V_CMFB_S2.n1 V_CMFB_S2.t3 24.0005
R537 V_CMFB_S2.n0 V_CMFB_S2.t0 24.0005
R538 V_CMFB_S2.n0 V_CMFB_S2.t2 24.0005
R539 GNDA.n2019 GNDA.n2018 11953.3
R540 GNDA.n2019 GNDA.n16 11949.5
R541 GNDA.n208 GNDA.n207 11663.5
R542 GNDA.n206 GNDA.n18 11348.7
R543 GNDA.n210 GNDA.n205 11202.2
R544 GNDA.n209 GNDA.n16 10235.4
R545 GNDA.n206 GNDA.n205 10120
R546 GNDA.n207 GNDA.n17 5394.83
R547 GNDA.n209 GNDA.n208 5305.86
R548 GNDA.n2017 GNDA.n18 4721.86
R549 GNDA.n2018 GNDA.n2017 4497.78
R550 GNDA.n211 GNDA.n210 4387.43
R551 GNDA.n207 GNDA.n206 4120.63
R552 GNDA.n208 GNDA.n205 4120.63
R553 GNDA.n2018 GNDA.n17 4106.67
R554 GNDA.n2021 GNDA.n2019 3974.19
R555 GNDA.n211 GNDA.n16 3962.24
R556 GNDA.n210 GNDA.n209 2913.51
R557 GNDA.n18 GNDA.n17 2443.04
R558 GNDA.n2017 GNDA.n2016 2374.29
R559 GNDA.n1507 GNDA.n211 2243.1
R560 GNDA.n1373 GNDA.n1217 1367.21
R561 GNDA.n2016 GNDA.t33 1311.87
R562 GNDA.n1809 GNDA.n1806 1185.07
R563 GNDA.n1809 GNDA.n1808 1185.07
R564 GNDA.n1507 GNDA.n1506 1104.89
R565 GNDA.n221 GNDA.n217 669.307
R566 GNDA.n945 GNDA.n22 585
R567 GNDA.n969 GNDA.n818 585
R568 GNDA.n967 GNDA.n966 585
R569 GNDA.n965 GNDA.n820 585
R570 GNDA.n964 GNDA.n963 585
R571 GNDA.n961 GNDA.n821 585
R572 GNDA.n959 GNDA.n958 585
R573 GNDA.n957 GNDA.n822 585
R574 GNDA.n956 GNDA.n955 585
R575 GNDA.n953 GNDA.n823 585
R576 GNDA.n951 GNDA.n950 585
R577 GNDA.n949 GNDA.n824 585
R578 GNDA.n1994 GNDA.n1993 585
R579 GNDA.n1995 GNDA.n29 585
R580 GNDA.n1997 GNDA.n1996 585
R581 GNDA.n1999 GNDA.n27 585
R582 GNDA.n2001 GNDA.n2000 585
R583 GNDA.n2002 GNDA.n26 585
R584 GNDA.n2004 GNDA.n2003 585
R585 GNDA.n2006 GNDA.n24 585
R586 GNDA.n2008 GNDA.n2007 585
R587 GNDA.n2009 GNDA.n23 585
R588 GNDA.n2011 GNDA.n2010 585
R589 GNDA.n1352 GNDA.n1351 585
R590 GNDA.n1351 GNDA.n1350 585
R591 GNDA.n1352 GNDA.n1228 585
R592 GNDA.n1228 GNDA.n1227 585
R593 GNDA.n1354 GNDA.n1353 585
R594 GNDA.n1355 GNDA.n1354 585
R595 GNDA.n1226 GNDA.n1225 585
R596 GNDA.n1356 GNDA.n1226 585
R597 GNDA.n1360 GNDA.n1359 585
R598 GNDA.n1359 GNDA.n1358 585
R599 GNDA.n1361 GNDA.n1224 585
R600 GNDA.n1357 GNDA.n1224 585
R601 GNDA.n1363 GNDA.n1362 585
R602 GNDA.n1363 GNDA.n1211 585
R603 GNDA.n1364 GNDA.n1223 585
R604 GNDA.n1364 GNDA.n1212 585
R605 GNDA.n1367 GNDA.n1366 585
R606 GNDA.n1366 GNDA.n1365 585
R607 GNDA.n1368 GNDA.n1222 585
R608 GNDA.n1222 GNDA.n1221 585
R609 GNDA.n1370 GNDA.n1369 585
R610 GNDA.n1371 GNDA.n1370 585
R611 GNDA.n1220 GNDA.n1219 585
R612 GNDA.n1372 GNDA.n1220 585
R613 GNDA.n1375 GNDA.n1374 585
R614 GNDA.n1374 GNDA.n1373 585
R615 GNDA.n539 GNDA.n538 585
R616 GNDA.n538 GNDA.n51 585
R617 GNDA.n539 GNDA.n537 585
R618 GNDA.n537 GNDA.n536 585
R619 GNDA.n477 GNDA.n476 585
R620 GNDA.n535 GNDA.n477 585
R621 GNDA.n533 GNDA.n532 585
R622 GNDA.n534 GNDA.n533 585
R623 GNDA.n531 GNDA.n479 585
R624 GNDA.n479 GNDA.n478 585
R625 GNDA.n530 GNDA.n529 585
R626 GNDA.n529 GNDA.n528 585
R627 GNDA.n527 GNDA.n480 585
R628 GNDA.n527 GNDA.n58 585
R629 GNDA.n526 GNDA.n525 585
R630 GNDA.n526 GNDA.n59 585
R631 GNDA.n524 GNDA.n481 585
R632 GNDA.n484 GNDA.n481 585
R633 GNDA.n523 GNDA.n522 585
R634 GNDA.n522 GNDA.n521 585
R635 GNDA.n483 GNDA.n482 585
R636 GNDA.n520 GNDA.n483 585
R637 GNDA.n518 GNDA.n517 585
R638 GNDA.n519 GNDA.n518 585
R639 GNDA.n516 GNDA.n486 585
R640 GNDA.n486 GNDA.n485 585
R641 GNDA.n204 GNDA.n202 585
R642 GNDA.n1559 GNDA.n204 585
R643 GNDA.n1557 GNDA.n1556 585
R644 GNDA.n1558 GNDA.n1557 585
R645 GNDA.n1555 GNDA.n1509 585
R646 GNDA.n1509 GNDA.n1508 585
R647 GNDA.n1554 GNDA.n1553 585
R648 GNDA.n1553 GNDA.n1552 585
R649 GNDA.n1551 GNDA.n1510 585
R650 GNDA.n1551 GNDA.n65 585
R651 GNDA.n1550 GNDA.n1549 585
R652 GNDA.n1550 GNDA.n66 585
R653 GNDA.n1548 GNDA.n1511 585
R654 GNDA.n1514 GNDA.n1511 585
R655 GNDA.n1547 GNDA.n1546 585
R656 GNDA.n1546 GNDA.n1545 585
R657 GNDA.n1513 GNDA.n1512 585
R658 GNDA.n1544 GNDA.n1513 585
R659 GNDA.n1542 GNDA.n1541 585
R660 GNDA.n1543 GNDA.n1542 585
R661 GNDA.n1540 GNDA.n1515 585
R662 GNDA.n1515 GNDA.n52 585
R663 GNDA.n172 GNDA.n20 585
R664 GNDA.n1830 GNDA.n20 585
R665 GNDA.n1833 GNDA.n1832 585
R666 GNDA.n1832 GNDA.n1831 585
R667 GNDA.n175 GNDA.n174 585
R668 GNDA.n1829 GNDA.n175 585
R669 GNDA.n1827 GNDA.n1826 585
R670 GNDA.n1828 GNDA.n1827 585
R671 GNDA.n1821 GNDA.n176 585
R672 GNDA.n1813 GNDA.n176 585
R673 GNDA.n1816 GNDA.n1815 585
R674 GNDA.n1815 GNDA.n1814 585
R675 GNDA.n178 GNDA.n177 585
R676 GNDA.n193 GNDA.n178 585
R677 GNDA.n191 GNDA.n190 585
R678 GNDA.n192 GNDA.n191 585
R679 GNDA.n185 GNDA.n183 585
R680 GNDA.n183 GNDA.n182 585
R681 GNDA.n179 GNDA.n151 585
R682 GNDA.n181 GNDA.n179 585
R683 GNDA.n1889 GNDA.n149 585
R684 GNDA.n180 GNDA.n149 585
R685 GNDA.n1892 GNDA.n1891 585
R686 GNDA.n1893 GNDA.n1892 585
R687 GNDA.n2015 GNDA.n2014 585
R688 GNDA.n1691 GNDA.n1690 585
R689 GNDA.n1712 GNDA.n1711 585
R690 GNDA.n1706 GNDA.n196 585
R691 GNDA.n1901 GNDA.n1900 585
R692 GNDA.n1895 GNDA.n1894 585
R693 GNDA.n139 GNDA.n19 585
R694 GNDA.n1506 GNDA.n1505 585
R695 GNDA.n631 GNDA.n630 585
R696 GNDA.n628 GNDA.n627 585
R697 GNDA.n626 GNDA.n625 585
R698 GNDA.n600 GNDA.n450 585
R699 GNDA.n606 GNDA.n605 585
R700 GNDA.n608 GNDA.n599 585
R701 GNDA.n610 GNDA.n609 585
R702 GNDA.n596 GNDA.n595 585
R703 GNDA.n616 GNDA.n615 585
R704 GNDA.n619 GNDA.n618 585
R705 GNDA.n594 GNDA.n473 585
R706 GNDA.n592 GNDA.n591 585
R707 GNDA.n755 GNDA.n754 585
R708 GNDA.n752 GNDA.n751 585
R709 GNDA.n637 GNDA.n636 585
R710 GNDA.n745 GNDA.n744 585
R711 GNDA.n742 GNDA.n741 585
R712 GNDA.n731 GNDA.n730 585
R713 GNDA.n733 GNDA.n732 585
R714 GNDA.n728 GNDA.n644 585
R715 GNDA.n727 GNDA.n726 585
R716 GNDA.n717 GNDA.n646 585
R717 GNDA.n719 GNDA.n718 585
R718 GNDA.n715 GNDA.n714 585
R719 GNDA.n944 GNDA.n825 585
R720 GNDA.n942 GNDA.n941 585
R721 GNDA.n861 GNDA.n826 585
R722 GNDA.n859 GNDA.n858 585
R723 GNDA.n871 GNDA.n870 585
R724 GNDA.n873 GNDA.n856 585
R725 GNDA.n875 GNDA.n874 585
R726 GNDA.n852 GNDA.n851 585
R727 GNDA.n882 GNDA.n881 585
R728 GNDA.n885 GNDA.n884 585
R729 GNDA.n850 GNDA.n846 585
R730 GNDA.n848 GNDA.n756 585
R731 GNDA.n1517 GNDA.n1516 585
R732 GNDA.n1519 GNDA.n1518 585
R733 GNDA.n1521 GNDA.n1520 585
R734 GNDA.n1523 GNDA.n1522 585
R735 GNDA.n1525 GNDA.n1524 585
R736 GNDA.n1527 GNDA.n1526 585
R737 GNDA.n1529 GNDA.n1528 585
R738 GNDA.n1531 GNDA.n1530 585
R739 GNDA.n1533 GNDA.n1532 585
R740 GNDA.n1535 GNDA.n1534 585
R741 GNDA.n1537 GNDA.n1536 585
R742 GNDA.n1539 GNDA.n1538 585
R743 GNDA.n1942 GNDA.n1941 585
R744 GNDA.n1944 GNDA.n1943 585
R745 GNDA.n1946 GNDA.n1945 585
R746 GNDA.n1948 GNDA.n1947 585
R747 GNDA.n1950 GNDA.n1949 585
R748 GNDA.n1952 GNDA.n1951 585
R749 GNDA.n1954 GNDA.n1953 585
R750 GNDA.n1956 GNDA.n1955 585
R751 GNDA.n1958 GNDA.n1957 585
R752 GNDA.n1960 GNDA.n1959 585
R753 GNDA.n1962 GNDA.n1961 585
R754 GNDA.n1964 GNDA.n1963 585
R755 GNDA.n1992 GNDA.n30 585
R756 GNDA.n101 GNDA.n32 585
R757 GNDA.n103 GNDA.n102 585
R758 GNDA.n105 GNDA.n104 585
R759 GNDA.n107 GNDA.n106 585
R760 GNDA.n109 GNDA.n108 585
R761 GNDA.n111 GNDA.n110 585
R762 GNDA.n113 GNDA.n112 585
R763 GNDA.n115 GNDA.n114 585
R764 GNDA.n117 GNDA.n116 585
R765 GNDA.n119 GNDA.n118 585
R766 GNDA.n121 GNDA.n120 585
R767 GNDA.n1286 GNDA.n1059 585
R768 GNDA.n1289 GNDA.n1288 585
R769 GNDA.n1285 GNDA.n1255 585
R770 GNDA.n1283 GNDA.n1282 585
R771 GNDA.n1277 GNDA.n1256 585
R772 GNDA.n1272 GNDA.n1271 585
R773 GNDA.n1269 GNDA.n1257 585
R774 GNDA.n1267 GNDA.n1266 585
R775 GNDA.n1261 GNDA.n1259 585
R776 GNDA.n1232 GNDA.n1230 585
R777 GNDA.n1346 GNDA.n1345 585
R778 GNDA.n1348 GNDA.n1229 585
R779 GNDA.n495 GNDA.n431 585
R780 GNDA.n497 GNDA.n493 585
R781 GNDA.n499 GNDA.n498 585
R782 GNDA.n500 GNDA.n492 585
R783 GNDA.n502 GNDA.n501 585
R784 GNDA.n504 GNDA.n490 585
R785 GNDA.n506 GNDA.n505 585
R786 GNDA.n507 GNDA.n489 585
R787 GNDA.n509 GNDA.n508 585
R788 GNDA.n511 GNDA.n488 585
R789 GNDA.n512 GNDA.n487 585
R790 GNDA.n515 GNDA.n514 585
R791 GNDA.n808 GNDA.n807 585
R792 GNDA.n805 GNDA.n781 585
R793 GNDA.n804 GNDA.n803 585
R794 GNDA.n802 GNDA.n801 585
R795 GNDA.n800 GNDA.n783 585
R796 GNDA.n798 GNDA.n797 585
R797 GNDA.n796 GNDA.n784 585
R798 GNDA.n795 GNDA.n794 585
R799 GNDA.n792 GNDA.n785 585
R800 GNDA.n790 GNDA.n789 585
R801 GNDA.n788 GNDA.n787 585
R802 GNDA.n434 GNDA.n430 585
R803 GNDA.n971 GNDA.n970 585
R804 GNDA.n972 GNDA.n817 585
R805 GNDA.n974 GNDA.n973 585
R806 GNDA.n976 GNDA.n815 585
R807 GNDA.n978 GNDA.n977 585
R808 GNDA.n979 GNDA.n814 585
R809 GNDA.n981 GNDA.n980 585
R810 GNDA.n983 GNDA.n812 585
R811 GNDA.n985 GNDA.n984 585
R812 GNDA.n986 GNDA.n811 585
R813 GNDA.n988 GNDA.n987 585
R814 GNDA.n990 GNDA.n810 585
R815 GNDA.n1399 GNDA.n1398 585
R816 GNDA.n1398 GNDA.n1397 585
R817 GNDA.n1196 GNDA.n1195 585
R818 GNDA.n1396 GNDA.n1196 585
R819 GNDA.n1394 GNDA.n1393 585
R820 GNDA.n1395 GNDA.n1394 585
R821 GNDA.n1392 GNDA.n1198 585
R822 GNDA.n1198 GNDA.n1197 585
R823 GNDA.n1391 GNDA.n1390 585
R824 GNDA.n1390 GNDA.n1389 585
R825 GNDA.n1200 GNDA.n1199 585
R826 GNDA.n1388 GNDA.n1200 585
R827 GNDA.n1386 GNDA.n1385 585
R828 GNDA.n1387 GNDA.n1386 585
R829 GNDA.n1384 GNDA.n1214 585
R830 GNDA.n1214 GNDA.n1213 585
R831 GNDA.n1383 GNDA.n1382 585
R832 GNDA.n1382 GNDA.n1381 585
R833 GNDA.n1216 GNDA.n1215 585
R834 GNDA.n1380 GNDA.n1216 585
R835 GNDA.n1378 GNDA.n1377 585
R836 GNDA.n1379 GNDA.n1378 585
R837 GNDA.n1376 GNDA.n1218 585
R838 GNDA.n1218 GNDA.n1217 585
R839 GNDA.n406 GNDA.n405 585
R840 GNDA.n405 GNDA.n54 585
R841 GNDA.n407 GNDA.n252 585
R842 GNDA.n252 GNDA.n251 585
R843 GNDA.n409 GNDA.n408 585
R844 GNDA.n410 GNDA.n409 585
R845 GNDA.n250 GNDA.n249 585
R846 GNDA.n411 GNDA.n250 585
R847 GNDA.n414 GNDA.n413 585
R848 GNDA.n413 GNDA.n412 585
R849 GNDA.n415 GNDA.n248 585
R850 GNDA.n248 GNDA.n57 585
R851 GNDA.n417 GNDA.n416 585
R852 GNDA.n417 GNDA.n56 585
R853 GNDA.n418 GNDA.n247 585
R854 GNDA.n419 GNDA.n418 585
R855 GNDA.n422 GNDA.n421 585
R856 GNDA.n421 GNDA.n420 585
R857 GNDA.n423 GNDA.n246 585
R858 GNDA.n246 GNDA.n245 585
R859 GNDA.n425 GNDA.n424 585
R860 GNDA.n426 GNDA.n425 585
R861 GNDA.n230 GNDA.n227 585
R862 GNDA.n427 GNDA.n230 585
R863 GNDA.n404 GNDA.n253 585
R864 GNDA.n404 GNDA.n22 585
R865 GNDA.n403 GNDA.n254 585
R866 GNDA.n401 GNDA.n400 585
R867 GNDA.n399 GNDA.n255 585
R868 GNDA.n398 GNDA.n397 585
R869 GNDA.n395 GNDA.n256 585
R870 GNDA.n393 GNDA.n392 585
R871 GNDA.n391 GNDA.n257 585
R872 GNDA.n390 GNDA.n389 585
R873 GNDA.n387 GNDA.n258 585
R874 GNDA.n385 GNDA.n384 585
R875 GNDA.n380 GNDA.n260 585
R876 GNDA.n378 GNDA.n377 585
R877 GNDA.n297 GNDA.n261 585
R878 GNDA.n295 GNDA.n294 585
R879 GNDA.n307 GNDA.n306 585
R880 GNDA.n309 GNDA.n292 585
R881 GNDA.n311 GNDA.n310 585
R882 GNDA.n288 GNDA.n287 585
R883 GNDA.n318 GNDA.n317 585
R884 GNDA.n321 GNDA.n320 585
R885 GNDA.n286 GNDA.n281 585
R886 GNDA.n284 GNDA.n283 585
R887 GNDA.n383 GNDA.n382 585
R888 GNDA.n383 GNDA.n259 585
R889 GNDA.n1084 GNDA.n242 585
R890 GNDA.n1119 GNDA.n1118 585
R891 GNDA.n1116 GNDA.n1086 585
R892 GNDA.n1114 GNDA.n1113 585
R893 GNDA.n1108 GNDA.n1087 585
R894 GNDA.n1103 GNDA.n1102 585
R895 GNDA.n1100 GNDA.n1088 585
R896 GNDA.n1098 GNDA.n1097 585
R897 GNDA.n1092 GNDA.n1090 585
R898 GNDA.n1062 GNDA.n1061 585
R899 GNDA.n1176 GNDA.n1175 585
R900 GNDA.n1179 GNDA.n1178 585
R901 GNDA.n1445 GNDA.n243 585
R902 GNDA.n1445 GNDA.n1444 585
R903 GNDA.n1482 GNDA.n229 585
R904 GNDA.n1471 GNDA.n228 585
R905 GNDA.n1472 GNDA.n231 585
R906 GNDA.n1475 GNDA.n1474 585
R907 GNDA.n1469 GNDA.n233 585
R908 GNDA.n1467 GNDA.n1466 585
R909 GNDA.n235 GNDA.n234 585
R910 GNDA.n1460 GNDA.n1459 585
R911 GNDA.n1457 GNDA.n237 585
R912 GNDA.n1455 GNDA.n1454 585
R913 GNDA.n239 GNDA.n238 585
R914 GNDA.n1448 GNDA.n1447 585
R915 GNDA.n428 GNDA.n243 585
R916 GNDA.n1444 GNDA.n428 585
R917 GNDA.n1449 GNDA.n1448 585
R918 GNDA.n1451 GNDA.n239 585
R919 GNDA.n1454 GNDA.n1453 585
R920 GNDA.n237 GNDA.n236 585
R921 GNDA.n1461 GNDA.n1460 585
R922 GNDA.n1463 GNDA.n235 585
R923 GNDA.n1466 GNDA.n1465 585
R924 GNDA.n233 GNDA.n232 585
R925 GNDA.n1476 GNDA.n1475 585
R926 GNDA.n1478 GNDA.n231 585
R927 GNDA.n1479 GNDA.n228 585
R928 GNDA.n1482 GNDA.n1481 585
R929 GNDA.n1016 GNDA.n633 585
R930 GNDA.n1019 GNDA.n633 585
R931 GNDA.n993 GNDA.n780 585
R932 GNDA.n994 GNDA.n778 585
R933 GNDA.n995 GNDA.n777 585
R934 GNDA.n775 GNDA.n773 585
R935 GNDA.n1001 GNDA.n772 585
R936 GNDA.n1002 GNDA.n770 585
R937 GNDA.n1003 GNDA.n769 585
R938 GNDA.n767 GNDA.n765 585
R939 GNDA.n1008 GNDA.n764 585
R940 GNDA.n1009 GNDA.n762 585
R941 GNDA.n761 GNDA.n758 585
R942 GNDA.n1014 GNDA.n757 585
R943 GNDA.n1017 GNDA.n1016 585
R944 GNDA.n1019 GNDA.n1017 585
R945 GNDA.n1014 GNDA.n1013 585
R946 GNDA.n1011 GNDA.n758 585
R947 GNDA.n1010 GNDA.n1009 585
R948 GNDA.n1008 GNDA.n1007 585
R949 GNDA.n1006 GNDA.n765 585
R950 GNDA.n1004 GNDA.n1003 585
R951 GNDA.n1002 GNDA.n766 585
R952 GNDA.n1001 GNDA.n1000 585
R953 GNDA.n998 GNDA.n773 585
R954 GNDA.n996 GNDA.n995 585
R955 GNDA.n994 GNDA.n774 585
R956 GNDA.n993 GNDA.n992 585
R957 GNDA.n1903 GNDA.n134 585
R958 GNDA.n1903 GNDA.n1902 585
R959 GNDA.n1940 GNDA.n1939 585
R960 GNDA.n1928 GNDA.n100 585
R961 GNDA.n1929 GNDA.n122 585
R962 GNDA.n1932 GNDA.n1931 585
R963 GNDA.n1927 GNDA.n124 585
R964 GNDA.n1925 GNDA.n1924 585
R965 GNDA.n126 GNDA.n125 585
R966 GNDA.n1918 GNDA.n1917 585
R967 GNDA.n1915 GNDA.n128 585
R968 GNDA.n1913 GNDA.n1912 585
R969 GNDA.n130 GNDA.n129 585
R970 GNDA.n1906 GNDA.n1905 585
R971 GNDA.n147 GNDA.n134 585
R972 GNDA.n148 GNDA.n147 585
R973 GNDA.n1907 GNDA.n1906 585
R974 GNDA.n1909 GNDA.n130 585
R975 GNDA.n1912 GNDA.n1911 585
R976 GNDA.n128 GNDA.n127 585
R977 GNDA.n1919 GNDA.n1918 585
R978 GNDA.n1921 GNDA.n126 585
R979 GNDA.n1924 GNDA.n1923 585
R980 GNDA.n124 GNDA.n123 585
R981 GNDA.n1933 GNDA.n1932 585
R982 GNDA.n1935 GNDA.n122 585
R983 GNDA.n1936 GNDA.n100 585
R984 GNDA.n1939 GNDA.n1938 585
R985 GNDA.n1737 GNDA.n133 585
R986 GNDA.n135 GNDA.n133 585
R987 GNDA.n9 GNDA.n6 585
R988 GNDA.n1807 GNDA.n6 585
R989 GNDA.n2037 GNDA.n2036 585
R990 GNDA.n2038 GNDA.n2037 585
R991 GNDA.n7 GNDA.n5 585
R992 GNDA.n2039 GNDA.n5 585
R993 GNDA.n2042 GNDA.n2041 585
R994 GNDA.n2041 GNDA.n2040 585
R995 GNDA.n11 GNDA.n4 585
R996 GNDA.n2020 GNDA.n4 585
R997 GNDA.n2024 GNDA.n2023 585
R998 GNDA.n2023 GNDA.n2022 585
R999 GNDA.n15 GNDA.n14 585
R1000 GNDA.n1795 GNDA.n15 585
R1001 GNDA.n1798 GNDA.n1797 585
R1002 GNDA.n1797 GNDA.n1796 585
R1003 GNDA.n1723 GNDA.n1720 585
R1004 GNDA.n1794 GNDA.n1720 585
R1005 GNDA.n1804 GNDA.n1803 585
R1006 GNDA.n1805 GNDA.n1804 585
R1007 GNDA.n1721 GNDA.n1719 585
R1008 GNDA.n1719 GNDA.n1718 585
R1009 GNDA.n1585 GNDA.n197 585
R1010 GNDA.n1626 GNDA.n197 585
R1011 GNDA.n1629 GNDA.n1628 585
R1012 GNDA.n1628 GNDA.n1627 585
R1013 GNDA.n1588 GNDA.n1587 585
R1014 GNDA.n1625 GNDA.n1588 585
R1015 GNDA.n1623 GNDA.n1622 585
R1016 GNDA.n1624 GNDA.n1623 585
R1017 GNDA.n1617 GNDA.n1589 585
R1018 GNDA.n1609 GNDA.n1589 585
R1019 GNDA.n1612 GNDA.n1611 585
R1020 GNDA.n1611 GNDA.n1610 585
R1021 GNDA.n1591 GNDA.n1590 585
R1022 GNDA.n1606 GNDA.n1591 585
R1023 GNDA.n1604 GNDA.n1603 585
R1024 GNDA.n1605 GNDA.n1604 585
R1025 GNDA.n1598 GNDA.n1596 585
R1026 GNDA.n1596 GNDA.n1595 585
R1027 GNDA.n1592 GNDA.n1564 585
R1028 GNDA.n1594 GNDA.n1592 585
R1029 GNDA.n1685 GNDA.n201 585
R1030 GNDA.n1593 GNDA.n201 585
R1031 GNDA.n1688 GNDA.n1687 585
R1032 GNDA.n1689 GNDA.n1688 585
R1033 GNDA.n1562 GNDA.n203 585
R1034 GNDA.n203 GNDA.n199 585
R1035 GNDA.n1562 GNDA.n1561 585
R1036 GNDA.n1561 GNDA.n1560 585
R1037 GNDA.n1715 GNDA.n1714 585
R1038 GNDA.n1714 GNDA.n1713 585
R1039 GNDA.n1966 GNDA.n96 585
R1040 GNDA.n1967 GNDA.n94 585
R1041 GNDA.n1970 GNDA.n93 585
R1042 GNDA.n1971 GNDA.n91 585
R1043 GNDA.n1974 GNDA.n90 585
R1044 GNDA.n1975 GNDA.n88 585
R1045 GNDA.n1978 GNDA.n87 585
R1046 GNDA.n1979 GNDA.n85 585
R1047 GNDA.n1982 GNDA.n84 585
R1048 GNDA.n1984 GNDA.n82 585
R1049 GNDA.n1985 GNDA.n81 585
R1050 GNDA.n1986 GNDA.n79 585
R1051 GNDA.n1716 GNDA.n1715 585
R1052 GNDA.n1717 GNDA.n1716 585
R1053 GNDA.n1987 GNDA.n1986 585
R1054 GNDA.n1985 GNDA.n76 585
R1055 GNDA.n1984 GNDA.n1983 585
R1056 GNDA.n1982 GNDA.n1981 585
R1057 GNDA.n1980 GNDA.n1979 585
R1058 GNDA.n1978 GNDA.n1977 585
R1059 GNDA.n1976 GNDA.n1975 585
R1060 GNDA.n1974 GNDA.n1973 585
R1061 GNDA.n1972 GNDA.n1971 585
R1062 GNDA.n1970 GNDA.n1969 585
R1063 GNDA.n1968 GNDA.n1967 585
R1064 GNDA.n1966 GNDA.n1965 585
R1065 GNDA.n1020 GNDA.n632 585
R1066 GNDA.n1020 GNDA.n1019 585
R1067 GNDA.n1057 GNDA.n433 585
R1068 GNDA.n1046 GNDA.n432 585
R1069 GNDA.n1047 GNDA.n435 585
R1070 GNDA.n1050 GNDA.n1049 585
R1071 GNDA.n1044 GNDA.n437 585
R1072 GNDA.n1042 GNDA.n1041 585
R1073 GNDA.n439 GNDA.n438 585
R1074 GNDA.n1035 GNDA.n1034 585
R1075 GNDA.n1032 GNDA.n441 585
R1076 GNDA.n1030 GNDA.n1029 585
R1077 GNDA.n443 GNDA.n442 585
R1078 GNDA.n1023 GNDA.n1022 585
R1079 GNDA.n1018 GNDA.n632 585
R1080 GNDA.n1019 GNDA.n1018 585
R1081 GNDA.n1024 GNDA.n1023 585
R1082 GNDA.n1026 GNDA.n443 585
R1083 GNDA.n1029 GNDA.n1028 585
R1084 GNDA.n441 GNDA.n440 585
R1085 GNDA.n1036 GNDA.n1035 585
R1086 GNDA.n1038 GNDA.n439 585
R1087 GNDA.n1041 GNDA.n1040 585
R1088 GNDA.n437 GNDA.n436 585
R1089 GNDA.n1051 GNDA.n1050 585
R1090 GNDA.n1053 GNDA.n435 585
R1091 GNDA.n1054 GNDA.n432 585
R1092 GNDA.n1057 GNDA.n1056 585
R1093 GNDA.n1442 GNDA.n244 585
R1094 GNDA.n1444 GNDA.n244 585
R1095 GNDA.n1419 GNDA.n1194 585
R1096 GNDA.n1420 GNDA.n1193 585
R1097 GNDA.n1421 GNDA.n1192 585
R1098 GNDA.n1207 GNDA.n1190 585
R1099 GNDA.n1427 GNDA.n1189 585
R1100 GNDA.n1428 GNDA.n1188 585
R1101 GNDA.n1429 GNDA.n1187 585
R1102 GNDA.n1204 GNDA.n1185 585
R1103 GNDA.n1434 GNDA.n1184 585
R1104 GNDA.n1435 GNDA.n1183 585
R1105 GNDA.n1201 GNDA.n1181 585
R1106 GNDA.n1440 GNDA.n1180 585
R1107 GNDA.n1443 GNDA.n1442 585
R1108 GNDA.n1444 GNDA.n1443 585
R1109 GNDA.n1440 GNDA.n1439 585
R1110 GNDA.n1437 GNDA.n1181 585
R1111 GNDA.n1436 GNDA.n1435 585
R1112 GNDA.n1434 GNDA.n1433 585
R1113 GNDA.n1432 GNDA.n1185 585
R1114 GNDA.n1430 GNDA.n1429 585
R1115 GNDA.n1428 GNDA.n1186 585
R1116 GNDA.n1427 GNDA.n1426 585
R1117 GNDA.n1424 GNDA.n1190 585
R1118 GNDA.n1422 GNDA.n1421 585
R1119 GNDA.n1420 GNDA.n1191 585
R1120 GNDA.n1419 GNDA.n1418 585
R1121 GNDA.n1484 GNDA.n226 585
R1122 GNDA.n226 GNDA.n225 585
R1123 GNDA.n1486 GNDA.n1485 585
R1124 GNDA.n1487 GNDA.n1486 585
R1125 GNDA.n224 GNDA.n223 585
R1126 GNDA.n1488 GNDA.n224 585
R1127 GNDA.n1491 GNDA.n1490 585
R1128 GNDA.n1490 GNDA.n1489 585
R1129 GNDA.n1492 GNDA.n220 585
R1130 GNDA.n220 GNDA.n218 585
R1131 GNDA.n1494 GNDA.n1493 585
R1132 GNDA.n1495 GNDA.n1494 585
R1133 GNDA.n1406 GNDA.n219 585
R1134 GNDA.n219 GNDA.n216 585
R1135 GNDA.n1409 GNDA.n1408 585
R1136 GNDA.n1408 GNDA.n1407 585
R1137 GNDA.n1410 GNDA.n1404 585
R1138 GNDA.n1404 GNDA.n1403 585
R1139 GNDA.n1412 GNDA.n1411 585
R1140 GNDA.n1413 GNDA.n1412 585
R1141 GNDA.n1405 GNDA.n1401 585
R1142 GNDA.n1414 GNDA.n1401 585
R1143 GNDA.n1416 GNDA.n1402 585
R1144 GNDA.n1416 GNDA.n1415 585
R1145 GNDA.n213 GNDA.n212 585
R1146 GNDA.n1497 GNDA.n1496 585
R1147 GNDA.n1496 GNDA.t85 585
R1148 GNDA.n1692 GNDA.t95 409.067
R1149 GNDA.n1710 GNDA.t90 409.067
R1150 GNDA.n1707 GNDA.t101 409.067
R1151 GNDA.n1899 GNDA.t107 409.067
R1152 GNDA.n1896 GNDA.t110 409.067
R1153 GNDA.n140 GNDA.t104 409.067
R1154 GNDA.n136 GNDA.n67 370.214
R1155 GNDA.n70 GNDA.n69 370.214
R1156 GNDA.n136 GNDA.n68 365.957
R1157 GNDA.n1989 GNDA.n70 365.957
R1158 GNDA.t85 GNDA.n214 172.876
R1159 GNDA.t85 GNDA.n68 327.661
R1160 GNDA.t85 GNDA.n1989 327.661
R1161 GNDA.t85 GNDA.n61 172.876
R1162 GNDA.t85 GNDA.n63 172.876
R1163 GNDA.t85 GNDA.n55 172.876
R1164 GNDA.t85 GNDA.n1210 172.615
R1165 GNDA.t85 GNDA.n67 323.404
R1166 GNDA.t85 GNDA.n69 323.404
R1167 GNDA.t85 GNDA.n60 172.615
R1168 GNDA.t85 GNDA.n62 172.615
R1169 GNDA.t85 GNDA.n215 172.615
R1170 GNDA.t85 GNDA.n52 274.089
R1171 GNDA.n381 GNDA.n22 263.904
R1172 GNDA.n948 GNDA.n947 263.904
R1173 GNDA.n2013 GNDA.n21 263.904
R1174 GNDA.n1418 GNDA.n1416 257.466
R1175 GNDA.n1965 GNDA.n1964 257.466
R1176 GNDA.n1056 GNDA.n434 257.466
R1177 GNDA.n1938 GNDA.n121 257.466
R1178 GNDA.n992 GNDA.n990 257.466
R1179 GNDA.n1538 GNDA.n1515 257.466
R1180 GNDA.n514 GNDA.n486 257.466
R1181 GNDA.n1374 GNDA.n1218 257.466
R1182 GNDA.n1481 GNDA.n230 257.466
R1183 GNDA.n968 GNDA.n22 254.34
R1184 GNDA.n962 GNDA.n22 254.34
R1185 GNDA.n960 GNDA.n22 254.34
R1186 GNDA.n954 GNDA.n22 254.34
R1187 GNDA.n952 GNDA.n22 254.34
R1188 GNDA.n946 GNDA.n22 254.34
R1189 GNDA.n31 GNDA.n22 254.34
R1190 GNDA.n1998 GNDA.n22 254.34
R1191 GNDA.n28 GNDA.n22 254.34
R1192 GNDA.n2005 GNDA.n22 254.34
R1193 GNDA.n25 GNDA.n22 254.34
R1194 GNDA.n2012 GNDA.n22 254.34
R1195 GNDA.n446 GNDA.n50 254.34
R1196 GNDA.n449 GNDA.n50 254.34
R1197 GNDA.n607 GNDA.n50 254.34
R1198 GNDA.n598 GNDA.n50 254.34
R1199 GNDA.n617 GNDA.n50 254.34
R1200 GNDA.n593 GNDA.n50 254.34
R1201 GNDA.n753 GNDA.n50 254.34
R1202 GNDA.n743 GNDA.n50 254.34
R1203 GNDA.n641 GNDA.n50 254.34
R1204 GNDA.n729 GNDA.n50 254.34
R1205 GNDA.n645 GNDA.n50 254.34
R1206 GNDA.n716 GNDA.n50 254.34
R1207 GNDA.n943 GNDA.n50 254.34
R1208 GNDA.n857 GNDA.n50 254.34
R1209 GNDA.n872 GNDA.n50 254.34
R1210 GNDA.n855 GNDA.n50 254.34
R1211 GNDA.n883 GNDA.n50 254.34
R1212 GNDA.n849 GNDA.n50 254.34
R1213 GNDA.n1990 GNDA.n49 254.34
R1214 GNDA.n1990 GNDA.n48 254.34
R1215 GNDA.n1990 GNDA.n47 254.34
R1216 GNDA.n1990 GNDA.n46 254.34
R1217 GNDA.n1990 GNDA.n45 254.34
R1218 GNDA.n1990 GNDA.n44 254.34
R1219 GNDA.n1990 GNDA.n43 254.34
R1220 GNDA.n1990 GNDA.n42 254.34
R1221 GNDA.n1990 GNDA.n41 254.34
R1222 GNDA.n1990 GNDA.n40 254.34
R1223 GNDA.n1990 GNDA.n39 254.34
R1224 GNDA.n1990 GNDA.n38 254.34
R1225 GNDA.n1991 GNDA.n1990 254.34
R1226 GNDA.n1990 GNDA.n37 254.34
R1227 GNDA.n1990 GNDA.n36 254.34
R1228 GNDA.n1990 GNDA.n35 254.34
R1229 GNDA.n1990 GNDA.n34 254.34
R1230 GNDA.n1990 GNDA.n33 254.34
R1231 GNDA.n1287 GNDA.n53 254.34
R1232 GNDA.n1284 GNDA.n53 254.34
R1233 GNDA.n1270 GNDA.n53 254.34
R1234 GNDA.n1268 GNDA.n53 254.34
R1235 GNDA.n1258 GNDA.n53 254.34
R1236 GNDA.n1347 GNDA.n53 254.34
R1237 GNDA.n496 GNDA.n64 254.34
R1238 GNDA.n494 GNDA.n64 254.34
R1239 GNDA.n503 GNDA.n64 254.34
R1240 GNDA.n491 GNDA.n64 254.34
R1241 GNDA.n510 GNDA.n64 254.34
R1242 GNDA.n513 GNDA.n64 254.34
R1243 GNDA.n806 GNDA.n64 254.34
R1244 GNDA.n782 GNDA.n64 254.34
R1245 GNDA.n799 GNDA.n64 254.34
R1246 GNDA.n793 GNDA.n64 254.34
R1247 GNDA.n791 GNDA.n64 254.34
R1248 GNDA.n786 GNDA.n64 254.34
R1249 GNDA.n819 GNDA.n64 254.34
R1250 GNDA.n975 GNDA.n64 254.34
R1251 GNDA.n816 GNDA.n64 254.34
R1252 GNDA.n982 GNDA.n64 254.34
R1253 GNDA.n813 GNDA.n64 254.34
R1254 GNDA.n989 GNDA.n64 254.34
R1255 GNDA.n402 GNDA.n22 254.34
R1256 GNDA.n396 GNDA.n22 254.34
R1257 GNDA.n394 GNDA.n22 254.34
R1258 GNDA.n388 GNDA.n22 254.34
R1259 GNDA.n386 GNDA.n22 254.34
R1260 GNDA.n379 GNDA.n53 254.34
R1261 GNDA.n293 GNDA.n53 254.34
R1262 GNDA.n308 GNDA.n53 254.34
R1263 GNDA.n291 GNDA.n53 254.34
R1264 GNDA.n319 GNDA.n53 254.34
R1265 GNDA.n285 GNDA.n53 254.34
R1266 GNDA.n1117 GNDA.n53 254.34
R1267 GNDA.n1115 GNDA.n53 254.34
R1268 GNDA.n1101 GNDA.n53 254.34
R1269 GNDA.n1099 GNDA.n53 254.34
R1270 GNDA.n1089 GNDA.n53 254.34
R1271 GNDA.n1177 GNDA.n53 254.34
R1272 GNDA.n1470 GNDA.n215 254.34
R1273 GNDA.n1473 GNDA.n215 254.34
R1274 GNDA.n1468 GNDA.n215 254.34
R1275 GNDA.n1458 GNDA.n215 254.34
R1276 GNDA.n1456 GNDA.n215 254.34
R1277 GNDA.n1446 GNDA.n215 254.34
R1278 GNDA.n1450 GNDA.n55 254.34
R1279 GNDA.n1452 GNDA.n55 254.34
R1280 GNDA.n1462 GNDA.n55 254.34
R1281 GNDA.n1464 GNDA.n55 254.34
R1282 GNDA.n1477 GNDA.n55 254.34
R1283 GNDA.n1480 GNDA.n55 254.34
R1284 GNDA.n779 GNDA.n60 254.34
R1285 GNDA.n776 GNDA.n60 254.34
R1286 GNDA.n771 GNDA.n60 254.34
R1287 GNDA.n768 GNDA.n60 254.34
R1288 GNDA.n763 GNDA.n60 254.34
R1289 GNDA.n760 GNDA.n60 254.34
R1290 GNDA.n1012 GNDA.n61 254.34
R1291 GNDA.n759 GNDA.n61 254.34
R1292 GNDA.n1005 GNDA.n61 254.34
R1293 GNDA.n999 GNDA.n61 254.34
R1294 GNDA.n997 GNDA.n61 254.34
R1295 GNDA.n991 GNDA.n61 254.34
R1296 GNDA.n99 GNDA.n67 254.34
R1297 GNDA.n1930 GNDA.n67 254.34
R1298 GNDA.n1926 GNDA.n67 254.34
R1299 GNDA.n1916 GNDA.n67 254.34
R1300 GNDA.n1914 GNDA.n67 254.34
R1301 GNDA.n1904 GNDA.n67 254.34
R1302 GNDA.n1908 GNDA.n68 254.34
R1303 GNDA.n1910 GNDA.n68 254.34
R1304 GNDA.n1920 GNDA.n68 254.34
R1305 GNDA.n1922 GNDA.n68 254.34
R1306 GNDA.n1934 GNDA.n68 254.34
R1307 GNDA.n1937 GNDA.n68 254.34
R1308 GNDA.n95 GNDA.n69 254.34
R1309 GNDA.n92 GNDA.n69 254.34
R1310 GNDA.n89 GNDA.n69 254.34
R1311 GNDA.n86 GNDA.n69 254.34
R1312 GNDA.n83 GNDA.n69 254.34
R1313 GNDA.n80 GNDA.n69 254.34
R1314 GNDA.n1989 GNDA.n1988 254.34
R1315 GNDA.n1989 GNDA.n75 254.34
R1316 GNDA.n1989 GNDA.n74 254.34
R1317 GNDA.n1989 GNDA.n73 254.34
R1318 GNDA.n1989 GNDA.n72 254.34
R1319 GNDA.n1989 GNDA.n71 254.34
R1320 GNDA.n1045 GNDA.n62 254.34
R1321 GNDA.n1048 GNDA.n62 254.34
R1322 GNDA.n1043 GNDA.n62 254.34
R1323 GNDA.n1033 GNDA.n62 254.34
R1324 GNDA.n1031 GNDA.n62 254.34
R1325 GNDA.n1021 GNDA.n62 254.34
R1326 GNDA.n1025 GNDA.n63 254.34
R1327 GNDA.n1027 GNDA.n63 254.34
R1328 GNDA.n1037 GNDA.n63 254.34
R1329 GNDA.n1039 GNDA.n63 254.34
R1330 GNDA.n1052 GNDA.n63 254.34
R1331 GNDA.n1055 GNDA.n63 254.34
R1332 GNDA.n1210 GNDA.n1209 254.34
R1333 GNDA.n1210 GNDA.n1208 254.34
R1334 GNDA.n1210 GNDA.n1206 254.34
R1335 GNDA.n1210 GNDA.n1205 254.34
R1336 GNDA.n1210 GNDA.n1203 254.34
R1337 GNDA.n1210 GNDA.n1202 254.34
R1338 GNDA.n1438 GNDA.n214 254.34
R1339 GNDA.n1182 GNDA.n214 254.34
R1340 GNDA.n1431 GNDA.n214 254.34
R1341 GNDA.n1425 GNDA.n214 254.34
R1342 GNDA.n1423 GNDA.n214 254.34
R1343 GNDA.n1417 GNDA.n214 254.34
R1344 GNDA.n229 GNDA.n226 251.614
R1345 GNDA.n1941 GNDA.n1940 251.614
R1346 GNDA.n807 GNDA.n780 251.614
R1347 GNDA.n1993 GNDA.n1992 251.614
R1348 GNDA.n970 GNDA.n969 251.614
R1349 GNDA.n1516 GNDA.n96 251.614
R1350 GNDA.n495 GNDA.n433 251.614
R1351 GNDA.n1398 GNDA.n1194 251.614
R1352 GNDA.n405 GNDA.n404 251.614
R1353 GNDA.t85 GNDA.n217 250.349
R1354 GNDA.n485 GNDA.t12 248.139
R1355 GNDA.t10 GNDA.t3 224.626
R1356 GNDA.n1632 GNDA.n1631 221.667
R1357 GNDA.n1122 GNDA.n1121 221.667
R1358 GNDA.n749 GNDA.n638 221.667
R1359 GNDA.n1836 GNDA.n1835 221.667
R1360 GNDA.n938 GNDA.n829 221.667
R1361 GNDA.n461 GNDA.n452 221.667
R1362 GNDA.n1292 GNDA.n1291 221.667
R1363 GNDA.n374 GNDA.n264 221.667
R1364 GNDA.n2034 GNDA.n10 221.667
R1365 GNDA.t4 GNDA.t20 219.279
R1366 GNDA.n22 GNDA.t7 215
R1367 GNDA.n1506 GNDA.t38 205.945
R1368 GNDA.n1496 GNDA.n213 197
R1369 GNDA.n1178 GNDA.n429 195.049
R1370 GNDA.n1719 GNDA.n77 195.049
R1371 GNDA.n715 GNDA.n444 195.049
R1372 GNDA.n1892 GNDA.n131 195.049
R1373 GNDA.n848 GNDA.n634 195.049
R1374 GNDA.n1688 GNDA.n200 195.049
R1375 GNDA.n592 GNDA.n475 195.049
R1376 GNDA.n1349 GNDA.n1348 195.049
R1377 GNDA.n284 GNDA.n240 195.049
R1378 GNDA.n1608 GNDA.n1607 195
R1379 GNDA.n1812 GNDA.n1811 195
R1380 GNDA.n1445 GNDA.n242 187.249
R1381 GNDA.n1903 GNDA.n133 187.249
R1382 GNDA.n754 GNDA.n633 187.249
R1383 GNDA.n2014 GNDA.n20 187.249
R1384 GNDA.n945 GNDA.n944 187.249
R1385 GNDA.n1714 GNDA.n197 187.249
R1386 GNDA.n1020 GNDA.n631 187.249
R1387 GNDA.n1286 GNDA.n244 187.249
R1388 GNDA.n382 GNDA.n380 187.249
R1389 GNDA.n1649 GNDA.n1648 185
R1390 GNDA.n1647 GNDA.n1646 185
R1391 GNDA.n1645 GNDA.n1644 185
R1392 GNDA.n1643 GNDA.n1642 185
R1393 GNDA.n1641 GNDA.n1640 185
R1394 GNDA.n1639 GNDA.n1638 185
R1395 GNDA.n1637 GNDA.n1636 185
R1396 GNDA.n1635 GNDA.n1634 185
R1397 GNDA.n1633 GNDA.n1632 185
R1398 GNDA.n1651 GNDA.n1650 185
R1399 GNDA.n1652 GNDA.n1574 185
R1400 GNDA.t100 GNDA.n1574 185
R1401 GNDA.n1654 GNDA.n1653 185
R1402 GNDA.n1656 GNDA.n1655 185
R1403 GNDA.n1658 GNDA.n1657 185
R1404 GNDA.n1660 GNDA.n1659 185
R1405 GNDA.n1662 GNDA.n1661 185
R1406 GNDA.n1664 GNDA.n1663 185
R1407 GNDA.n1666 GNDA.n1665 185
R1408 GNDA.n1565 GNDA.n1563 185
R1409 GNDA.n1681 GNDA.n1680 185
R1410 GNDA.n1679 GNDA.n1584 185
R1411 GNDA.n1678 GNDA.n1677 185
R1412 GNDA.n1676 GNDA.n1675 185
R1413 GNDA.n1674 GNDA.n1673 185
R1414 GNDA.n1672 GNDA.n1671 185
R1415 GNDA.n1670 GNDA.n1669 185
R1416 GNDA.n1668 GNDA.n1667 185
R1417 GNDA.n1139 GNDA.n1138 185
R1418 GNDA.n1137 GNDA.n1136 185
R1419 GNDA.n1135 GNDA.n1134 185
R1420 GNDA.n1133 GNDA.n1132 185
R1421 GNDA.n1131 GNDA.n1130 185
R1422 GNDA.n1129 GNDA.n1128 185
R1423 GNDA.n1127 GNDA.n1126 185
R1424 GNDA.n1125 GNDA.n1124 185
R1425 GNDA.n1123 GNDA.n1122 185
R1426 GNDA.n1141 GNDA.n1140 185
R1427 GNDA.n1142 GNDA.n1072 185
R1428 GNDA.t87 GNDA.n1072 185
R1429 GNDA.n1144 GNDA.n1143 185
R1430 GNDA.n1146 GNDA.n1145 185
R1431 GNDA.n1148 GNDA.n1147 185
R1432 GNDA.n1150 GNDA.n1149 185
R1433 GNDA.n1152 GNDA.n1151 185
R1434 GNDA.n1154 GNDA.n1153 185
R1435 GNDA.n1156 GNDA.n1155 185
R1436 GNDA.n1083 GNDA.n1063 185
R1437 GNDA.n1171 GNDA.n1170 185
R1438 GNDA.n1169 GNDA.n1082 185
R1439 GNDA.n1168 GNDA.n1167 185
R1440 GNDA.n1166 GNDA.n1165 185
R1441 GNDA.n1164 GNDA.n1163 185
R1442 GNDA.n1162 GNDA.n1161 185
R1443 GNDA.n1160 GNDA.n1159 185
R1444 GNDA.n1158 GNDA.n1157 185
R1445 GNDA.n676 GNDA.n656 185
R1446 GNDA.n675 GNDA.n674 185
R1447 GNDA.n673 GNDA.n672 185
R1448 GNDA.n671 GNDA.n658 185
R1449 GNDA.n669 GNDA.n668 185
R1450 GNDA.n667 GNDA.n659 185
R1451 GNDA.n666 GNDA.n665 185
R1452 GNDA.n663 GNDA.n661 185
R1453 GNDA.n660 GNDA.n638 185
R1454 GNDA.n679 GNDA.n678 185
R1455 GNDA.n680 GNDA.n655 185
R1456 GNDA.n655 GNDA.t86 185
R1457 GNDA.n682 GNDA.n681 185
R1458 GNDA.n684 GNDA.n654 185
R1459 GNDA.n687 GNDA.n686 185
R1460 GNDA.n688 GNDA.n653 185
R1461 GNDA.n690 GNDA.n689 185
R1462 GNDA.n692 GNDA.n652 185
R1463 GNDA.n695 GNDA.n694 185
R1464 GNDA.n712 GNDA.n647 185
R1465 GNDA.n711 GNDA.n710 185
R1466 GNDA.n708 GNDA.n648 185
R1467 GNDA.n706 GNDA.n705 185
R1468 GNDA.n704 GNDA.n649 185
R1469 GNDA.n703 GNDA.n702 185
R1470 GNDA.n700 GNDA.n650 185
R1471 GNDA.n698 GNDA.n697 185
R1472 GNDA.n696 GNDA.n651 185
R1473 GNDA.n750 GNDA.n749 185
R1474 GNDA.n747 GNDA.n746 185
R1475 GNDA.n640 GNDA.n639 185
R1476 GNDA.n740 GNDA.n739 185
R1477 GNDA.n737 GNDA.n642 185
R1478 GNDA.n735 GNDA.n734 185
R1479 GNDA.n725 GNDA.n643 185
R1480 GNDA.n724 GNDA.n723 185
R1481 GNDA.n721 GNDA.n720 185
R1482 GNDA.n721 GNDA.t86 185
R1483 GNDA.n1853 GNDA.n1852 185
R1484 GNDA.n1851 GNDA.n1850 185
R1485 GNDA.n1849 GNDA.n1848 185
R1486 GNDA.n1847 GNDA.n1846 185
R1487 GNDA.n1845 GNDA.n1844 185
R1488 GNDA.n1843 GNDA.n1842 185
R1489 GNDA.n1841 GNDA.n1840 185
R1490 GNDA.n1839 GNDA.n1838 185
R1491 GNDA.n1837 GNDA.n1836 185
R1492 GNDA.n1855 GNDA.n1854 185
R1493 GNDA.n1856 GNDA.n161 185
R1494 GNDA.t89 GNDA.n161 185
R1495 GNDA.n1858 GNDA.n1857 185
R1496 GNDA.n1860 GNDA.n1859 185
R1497 GNDA.n1862 GNDA.n1861 185
R1498 GNDA.n1864 GNDA.n1863 185
R1499 GNDA.n1866 GNDA.n1865 185
R1500 GNDA.n1868 GNDA.n1867 185
R1501 GNDA.n1870 GNDA.n1869 185
R1502 GNDA.n152 GNDA.n150 185
R1503 GNDA.n1885 GNDA.n1884 185
R1504 GNDA.n1883 GNDA.n171 185
R1505 GNDA.n1882 GNDA.n1881 185
R1506 GNDA.n1880 GNDA.n1879 185
R1507 GNDA.n1878 GNDA.n1877 185
R1508 GNDA.n1876 GNDA.n1875 185
R1509 GNDA.n1874 GNDA.n1873 185
R1510 GNDA.n1872 GNDA.n1871 185
R1511 GNDA.n1835 GNDA.n1834 185
R1512 GNDA.n1825 GNDA.n1824 185
R1513 GNDA.n1823 GNDA.n1822 185
R1514 GNDA.n1820 GNDA.n1819 185
R1515 GNDA.n1818 GNDA.n1817 185
R1516 GNDA.n189 GNDA.n188 185
R1517 GNDA.n187 GNDA.n186 185
R1518 GNDA.n184 GNDA.n153 185
R1519 GNDA.n1888 GNDA.n1887 185
R1520 GNDA.n1887 GNDA.t89 185
R1521 GNDA.n924 GNDA.n834 185
R1522 GNDA.n926 GNDA.n925 185
R1523 GNDA.n928 GNDA.n832 185
R1524 GNDA.n930 GNDA.n929 185
R1525 GNDA.n931 GNDA.n831 185
R1526 GNDA.n933 GNDA.n932 185
R1527 GNDA.n935 GNDA.n830 185
R1528 GNDA.n936 GNDA.n828 185
R1529 GNDA.n939 GNDA.n938 185
R1530 GNDA.n923 GNDA.n922 185
R1531 GNDA.n920 GNDA.n835 185
R1532 GNDA.n920 GNDA.t93 185
R1533 GNDA.n919 GNDA.n836 185
R1534 GNDA.n917 GNDA.n916 185
R1535 GNDA.n915 GNDA.n837 185
R1536 GNDA.n914 GNDA.n913 185
R1537 GNDA.n911 GNDA.n838 185
R1538 GNDA.n909 GNDA.n908 185
R1539 GNDA.n907 GNDA.n839 185
R1540 GNDA.n890 GNDA.n889 185
R1541 GNDA.n891 GNDA.n843 185
R1542 GNDA.n893 GNDA.n892 185
R1543 GNDA.n895 GNDA.n842 185
R1544 GNDA.n898 GNDA.n897 185
R1545 GNDA.n899 GNDA.n841 185
R1546 GNDA.n901 GNDA.n900 185
R1547 GNDA.n903 GNDA.n840 185
R1548 GNDA.n906 GNDA.n905 185
R1549 GNDA.n829 GNDA.n827 185
R1550 GNDA.n863 GNDA.n862 185
R1551 GNDA.n869 GNDA.n868 185
R1552 GNDA.n866 GNDA.n865 185
R1553 GNDA.n864 GNDA.n854 185
R1554 GNDA.n877 GNDA.n876 185
R1555 GNDA.n880 GNDA.n879 185
R1556 GNDA.n847 GNDA.n845 185
R1557 GNDA.n887 GNDA.n886 185
R1558 GNDA.n887 GNDA.t93 185
R1559 GNDA.n555 GNDA.n554 185
R1560 GNDA.n553 GNDA.n552 185
R1561 GNDA.n551 GNDA.n550 185
R1562 GNDA.n549 GNDA.n548 185
R1563 GNDA.n547 GNDA.n546 185
R1564 GNDA.n545 GNDA.n544 185
R1565 GNDA.n543 GNDA.n542 185
R1566 GNDA.n541 GNDA.n540 185
R1567 GNDA.n461 GNDA.n447 185
R1568 GNDA.n557 GNDA.n556 185
R1569 GNDA.n558 GNDA.n459 185
R1570 GNDA.t98 GNDA.n459 185
R1571 GNDA.n560 GNDA.n559 185
R1572 GNDA.n562 GNDA.n561 185
R1573 GNDA.n564 GNDA.n563 185
R1574 GNDA.n566 GNDA.n565 185
R1575 GNDA.n568 GNDA.n567 185
R1576 GNDA.n570 GNDA.n569 185
R1577 GNDA.n572 GNDA.n571 185
R1578 GNDA.n589 GNDA.n471 185
R1579 GNDA.n588 GNDA.n587 185
R1580 GNDA.n586 GNDA.n585 185
R1581 GNDA.n584 GNDA.n583 185
R1582 GNDA.n582 GNDA.n581 185
R1583 GNDA.n580 GNDA.n579 185
R1584 GNDA.n578 GNDA.n577 185
R1585 GNDA.n576 GNDA.n575 185
R1586 GNDA.n574 GNDA.n573 185
R1587 GNDA.n452 GNDA.n448 185
R1588 GNDA.n624 GNDA.n623 185
R1589 GNDA.n604 GNDA.n451 185
R1590 GNDA.n603 GNDA.n602 185
R1591 GNDA.n601 GNDA.n597 185
R1592 GNDA.n612 GNDA.n611 185
R1593 GNDA.n614 GNDA.n613 185
R1594 GNDA.n474 GNDA.n472 185
R1595 GNDA.n621 GNDA.n620 185
R1596 GNDA.t98 GNDA.n621 185
R1597 GNDA.n1309 GNDA.n1308 185
R1598 GNDA.n1307 GNDA.n1306 185
R1599 GNDA.n1305 GNDA.n1304 185
R1600 GNDA.n1303 GNDA.n1302 185
R1601 GNDA.n1301 GNDA.n1300 185
R1602 GNDA.n1299 GNDA.n1298 185
R1603 GNDA.n1297 GNDA.n1296 185
R1604 GNDA.n1295 GNDA.n1294 185
R1605 GNDA.n1293 GNDA.n1292 185
R1606 GNDA.n1311 GNDA.n1310 185
R1607 GNDA.n1312 GNDA.n1242 185
R1608 GNDA.t99 GNDA.n1242 185
R1609 GNDA.n1314 GNDA.n1313 185
R1610 GNDA.n1316 GNDA.n1315 185
R1611 GNDA.n1318 GNDA.n1317 185
R1612 GNDA.n1320 GNDA.n1319 185
R1613 GNDA.n1322 GNDA.n1321 185
R1614 GNDA.n1324 GNDA.n1323 185
R1615 GNDA.n1326 GNDA.n1325 185
R1616 GNDA.n1253 GNDA.n1233 185
R1617 GNDA.n1341 GNDA.n1340 185
R1618 GNDA.n1339 GNDA.n1252 185
R1619 GNDA.n1338 GNDA.n1337 185
R1620 GNDA.n1336 GNDA.n1335 185
R1621 GNDA.n1334 GNDA.n1333 185
R1622 GNDA.n1332 GNDA.n1331 185
R1623 GNDA.n1330 GNDA.n1329 185
R1624 GNDA.n1328 GNDA.n1327 185
R1625 GNDA.n1291 GNDA.n1290 185
R1626 GNDA.n1281 GNDA.n1280 185
R1627 GNDA.n1279 GNDA.n1278 185
R1628 GNDA.n1276 GNDA.n1275 185
R1629 GNDA.n1274 GNDA.n1273 185
R1630 GNDA.n1265 GNDA.n1264 185
R1631 GNDA.n1263 GNDA.n1262 185
R1632 GNDA.n1260 GNDA.n1234 185
R1633 GNDA.n1344 GNDA.n1343 185
R1634 GNDA.n1343 GNDA.t99 185
R1635 GNDA.n360 GNDA.n269 185
R1636 GNDA.n362 GNDA.n361 185
R1637 GNDA.n364 GNDA.n267 185
R1638 GNDA.n366 GNDA.n365 185
R1639 GNDA.n367 GNDA.n266 185
R1640 GNDA.n369 GNDA.n368 185
R1641 GNDA.n371 GNDA.n265 185
R1642 GNDA.n372 GNDA.n263 185
R1643 GNDA.n375 GNDA.n374 185
R1644 GNDA.n359 GNDA.n358 185
R1645 GNDA.n356 GNDA.n270 185
R1646 GNDA.n356 GNDA.t94 185
R1647 GNDA.n355 GNDA.n271 185
R1648 GNDA.n353 GNDA.n352 185
R1649 GNDA.n351 GNDA.n272 185
R1650 GNDA.n350 GNDA.n349 185
R1651 GNDA.n347 GNDA.n273 185
R1652 GNDA.n345 GNDA.n344 185
R1653 GNDA.n343 GNDA.n274 185
R1654 GNDA.n326 GNDA.n325 185
R1655 GNDA.n327 GNDA.n278 185
R1656 GNDA.n329 GNDA.n328 185
R1657 GNDA.n331 GNDA.n277 185
R1658 GNDA.n334 GNDA.n333 185
R1659 GNDA.n335 GNDA.n276 185
R1660 GNDA.n337 GNDA.n336 185
R1661 GNDA.n339 GNDA.n275 185
R1662 GNDA.n342 GNDA.n341 185
R1663 GNDA.n264 GNDA.n262 185
R1664 GNDA.n299 GNDA.n298 185
R1665 GNDA.n305 GNDA.n304 185
R1666 GNDA.n302 GNDA.n301 185
R1667 GNDA.n300 GNDA.n290 185
R1668 GNDA.n313 GNDA.n312 185
R1669 GNDA.n316 GNDA.n315 185
R1670 GNDA.n282 GNDA.n280 185
R1671 GNDA.n323 GNDA.n322 185
R1672 GNDA.n323 GNDA.t94 185
R1673 GNDA.n1121 GNDA.n1120 185
R1674 GNDA.n1112 GNDA.n1111 185
R1675 GNDA.n1110 GNDA.n1109 185
R1676 GNDA.n1107 GNDA.n1106 185
R1677 GNDA.n1105 GNDA.n1104 185
R1678 GNDA.n1096 GNDA.n1095 185
R1679 GNDA.n1094 GNDA.n1093 185
R1680 GNDA.n1091 GNDA.n1064 185
R1681 GNDA.n1174 GNDA.n1173 185
R1682 GNDA.n1173 GNDA.t87 185
R1683 GNDA.n1755 GNDA.n1733 185
R1684 GNDA.n1754 GNDA.n1753 185
R1685 GNDA.n1752 GNDA.n1751 185
R1686 GNDA.n1750 GNDA.n1735 185
R1687 GNDA.n1748 GNDA.n1747 185
R1688 GNDA.n1746 GNDA.n1736 185
R1689 GNDA.n1745 GNDA.n1744 185
R1690 GNDA.n1742 GNDA.n1740 185
R1691 GNDA.n1739 GNDA.n10 185
R1692 GNDA.n1758 GNDA.n1757 185
R1693 GNDA.n1759 GNDA.n1732 185
R1694 GNDA.n1732 GNDA.t84 185
R1695 GNDA.n1761 GNDA.n1760 185
R1696 GNDA.n1763 GNDA.n1731 185
R1697 GNDA.n1766 GNDA.n1765 185
R1698 GNDA.n1767 GNDA.n1730 185
R1699 GNDA.n1769 GNDA.n1768 185
R1700 GNDA.n1771 GNDA.n1729 185
R1701 GNDA.n1774 GNDA.n1773 185
R1702 GNDA.n1791 GNDA.n1790 185
R1703 GNDA.n1789 GNDA.n1788 185
R1704 GNDA.n1787 GNDA.n1725 185
R1705 GNDA.n1785 GNDA.n1784 185
R1706 GNDA.n1783 GNDA.n1726 185
R1707 GNDA.n1782 GNDA.n1781 185
R1708 GNDA.n1779 GNDA.n1727 185
R1709 GNDA.n1777 GNDA.n1776 185
R1710 GNDA.n1775 GNDA.n1728 185
R1711 GNDA.n2035 GNDA.n2034 185
R1712 GNDA.n2032 GNDA.n8 185
R1713 GNDA.n2031 GNDA.n3 185
R1714 GNDA.n2029 GNDA.n2 185
R1715 GNDA.n2028 GNDA.n12 185
R1716 GNDA.n2026 GNDA.n2025 185
R1717 GNDA.n1793 GNDA.n13 185
R1718 GNDA.n1800 GNDA.n1799 185
R1719 GNDA.n1802 GNDA.n1801 185
R1720 GNDA.n1801 GNDA.t84 185
R1721 GNDA.n1631 GNDA.n1630 185
R1722 GNDA.n1621 GNDA.n1620 185
R1723 GNDA.n1619 GNDA.n1618 185
R1724 GNDA.n1616 GNDA.n1615 185
R1725 GNDA.n1614 GNDA.n1613 185
R1726 GNDA.n1602 GNDA.n1601 185
R1727 GNDA.n1600 GNDA.n1599 185
R1728 GNDA.n1597 GNDA.n1566 185
R1729 GNDA.n1684 GNDA.n1683 185
R1730 GNDA.n1683 GNDA.t100 185
R1731 GNDA.n1415 GNDA.t85 183.948
R1732 GNDA.t85 GNDA.n427 183.948
R1733 GNDA.t85 GNDA.n51 180.023
R1734 GNDA.n1397 GNDA.t85 180.013
R1735 GNDA.t85 GNDA.n225 180.013
R1736 GNDA.n1455 GNDA.n238 175.546
R1737 GNDA.n1459 GNDA.n1457 175.546
R1738 GNDA.n1467 GNDA.n234 175.546
R1739 GNDA.n1474 GNDA.n1469 175.546
R1740 GNDA.n1472 GNDA.n1471 175.546
R1741 GNDA.n1416 GNDA.n1401 175.546
R1742 GNDA.n1412 GNDA.n1401 175.546
R1743 GNDA.n1412 GNDA.n1404 175.546
R1744 GNDA.n1408 GNDA.n1404 175.546
R1745 GNDA.n1408 GNDA.n219 175.546
R1746 GNDA.n1494 GNDA.n219 175.546
R1747 GNDA.n1494 GNDA.n220 175.546
R1748 GNDA.n1490 GNDA.n220 175.546
R1749 GNDA.n1490 GNDA.n224 175.546
R1750 GNDA.n1486 GNDA.n224 175.546
R1751 GNDA.n1486 GNDA.n226 175.546
R1752 GNDA.n1437 GNDA.n1436 175.546
R1753 GNDA.n1433 GNDA.n1432 175.546
R1754 GNDA.n1430 GNDA.n1186 175.546
R1755 GNDA.n1426 GNDA.n1424 175.546
R1756 GNDA.n1422 GNDA.n1191 175.546
R1757 GNDA.n1176 GNDA.n1061 175.546
R1758 GNDA.n1098 GNDA.n1090 175.546
R1759 GNDA.n1102 GNDA.n1100 175.546
R1760 GNDA.n1114 GNDA.n1087 175.546
R1761 GNDA.n1118 GNDA.n1116 175.546
R1762 GNDA.n1983 GNDA.n76 175.546
R1763 GNDA.n1981 GNDA.n1980 175.546
R1764 GNDA.n1977 GNDA.n1976 175.546
R1765 GNDA.n1973 GNDA.n1972 175.546
R1766 GNDA.n1969 GNDA.n1968 175.546
R1767 GNDA.n1804 GNDA.n1719 175.546
R1768 GNDA.n1804 GNDA.n1720 175.546
R1769 GNDA.n1797 GNDA.n1720 175.546
R1770 GNDA.n1797 GNDA.n15 175.546
R1771 GNDA.n2023 GNDA.n15 175.546
R1772 GNDA.n2023 GNDA.n4 175.546
R1773 GNDA.n2041 GNDA.n4 175.546
R1774 GNDA.n2041 GNDA.n5 175.546
R1775 GNDA.n2037 GNDA.n5 175.546
R1776 GNDA.n2037 GNDA.n6 175.546
R1777 GNDA.n133 GNDA.n6 175.546
R1778 GNDA.n1913 GNDA.n129 175.546
R1779 GNDA.n1917 GNDA.n1915 175.546
R1780 GNDA.n1925 GNDA.n125 175.546
R1781 GNDA.n1931 GNDA.n1927 175.546
R1782 GNDA.n1929 GNDA.n1928 175.546
R1783 GNDA.n1961 GNDA.n1960 175.546
R1784 GNDA.n1957 GNDA.n1956 175.546
R1785 GNDA.n1953 GNDA.n1952 175.546
R1786 GNDA.n1949 GNDA.n1948 175.546
R1787 GNDA.n1945 GNDA.n1944 175.546
R1788 GNDA.n762 GNDA.n761 175.546
R1789 GNDA.n767 GNDA.n764 175.546
R1790 GNDA.n770 GNDA.n769 175.546
R1791 GNDA.n775 GNDA.n772 175.546
R1792 GNDA.n778 GNDA.n777 175.546
R1793 GNDA.n790 GNDA.n787 175.546
R1794 GNDA.n794 GNDA.n792 175.546
R1795 GNDA.n798 GNDA.n784 175.546
R1796 GNDA.n801 GNDA.n800 175.546
R1797 GNDA.n805 GNDA.n804 175.546
R1798 GNDA.n1028 GNDA.n1026 175.546
R1799 GNDA.n1036 GNDA.n440 175.546
R1800 GNDA.n1040 GNDA.n1038 175.546
R1801 GNDA.n1051 GNDA.n436 175.546
R1802 GNDA.n1054 GNDA.n1053 175.546
R1803 GNDA.n718 GNDA.n717 175.546
R1804 GNDA.n728 GNDA.n727 175.546
R1805 GNDA.n732 GNDA.n731 175.546
R1806 GNDA.n744 GNDA.n742 175.546
R1807 GNDA.n752 GNDA.n636 175.546
R1808 GNDA.n1892 GNDA.n149 175.546
R1809 GNDA.n179 GNDA.n149 175.546
R1810 GNDA.n183 GNDA.n179 175.546
R1811 GNDA.n191 GNDA.n183 175.546
R1812 GNDA.n191 GNDA.n178 175.546
R1813 GNDA.n1815 GNDA.n178 175.546
R1814 GNDA.n1815 GNDA.n176 175.546
R1815 GNDA.n1827 GNDA.n176 175.546
R1816 GNDA.n1827 GNDA.n175 175.546
R1817 GNDA.n1832 GNDA.n175 175.546
R1818 GNDA.n1832 GNDA.n20 175.546
R1819 GNDA.n1911 GNDA.n1909 175.546
R1820 GNDA.n1919 GNDA.n127 175.546
R1821 GNDA.n1923 GNDA.n1921 175.546
R1822 GNDA.n1933 GNDA.n123 175.546
R1823 GNDA.n1936 GNDA.n1935 175.546
R1824 GNDA.n118 GNDA.n117 175.546
R1825 GNDA.n114 GNDA.n113 175.546
R1826 GNDA.n110 GNDA.n109 175.546
R1827 GNDA.n106 GNDA.n105 175.546
R1828 GNDA.n102 GNDA.n32 175.546
R1829 GNDA.n2011 GNDA.n23 175.546
R1830 GNDA.n2007 GNDA.n2006 175.546
R1831 GNDA.n2004 GNDA.n26 175.546
R1832 GNDA.n2000 GNDA.n1999 175.546
R1833 GNDA.n1997 GNDA.n29 175.546
R1834 GNDA.n951 GNDA.n824 175.546
R1835 GNDA.n955 GNDA.n953 175.546
R1836 GNDA.n959 GNDA.n822 175.546
R1837 GNDA.n963 GNDA.n961 175.546
R1838 GNDA.n967 GNDA.n820 175.546
R1839 GNDA.n988 GNDA.n811 175.546
R1840 GNDA.n984 GNDA.n983 175.546
R1841 GNDA.n981 GNDA.n814 175.546
R1842 GNDA.n977 GNDA.n976 175.546
R1843 GNDA.n974 GNDA.n817 175.546
R1844 GNDA.n1011 GNDA.n1010 175.546
R1845 GNDA.n1007 GNDA.n1006 175.546
R1846 GNDA.n1004 GNDA.n766 175.546
R1847 GNDA.n1000 GNDA.n998 175.546
R1848 GNDA.n996 GNDA.n774 175.546
R1849 GNDA.n884 GNDA.n850 175.546
R1850 GNDA.n882 GNDA.n851 175.546
R1851 GNDA.n874 GNDA.n873 175.546
R1852 GNDA.n871 GNDA.n858 175.546
R1853 GNDA.n942 GNDA.n826 175.546
R1854 GNDA.n1688 GNDA.n201 175.546
R1855 GNDA.n1592 GNDA.n201 175.546
R1856 GNDA.n1596 GNDA.n1592 175.546
R1857 GNDA.n1604 GNDA.n1596 175.546
R1858 GNDA.n1604 GNDA.n1591 175.546
R1859 GNDA.n1611 GNDA.n1591 175.546
R1860 GNDA.n1611 GNDA.n1589 175.546
R1861 GNDA.n1623 GNDA.n1589 175.546
R1862 GNDA.n1623 GNDA.n1588 175.546
R1863 GNDA.n1628 GNDA.n1588 175.546
R1864 GNDA.n1628 GNDA.n197 175.546
R1865 GNDA.n82 GNDA.n81 175.546
R1866 GNDA.n85 GNDA.n84 175.546
R1867 GNDA.n88 GNDA.n87 175.546
R1868 GNDA.n91 GNDA.n90 175.546
R1869 GNDA.n94 GNDA.n93 175.546
R1870 GNDA.n1536 GNDA.n1535 175.546
R1871 GNDA.n1532 GNDA.n1531 175.546
R1872 GNDA.n1528 GNDA.n1527 175.546
R1873 GNDA.n1524 GNDA.n1523 175.546
R1874 GNDA.n1520 GNDA.n1519 175.546
R1875 GNDA.n1561 GNDA.n204 175.546
R1876 GNDA.n1557 GNDA.n204 175.546
R1877 GNDA.n1557 GNDA.n1509 175.546
R1878 GNDA.n1553 GNDA.n1509 175.546
R1879 GNDA.n1553 GNDA.n1551 175.546
R1880 GNDA.n1551 GNDA.n1550 175.546
R1881 GNDA.n1550 GNDA.n1511 175.546
R1882 GNDA.n1546 GNDA.n1511 175.546
R1883 GNDA.n1546 GNDA.n1513 175.546
R1884 GNDA.n1542 GNDA.n1513 175.546
R1885 GNDA.n1542 GNDA.n1515 175.546
R1886 GNDA.n1030 GNDA.n442 175.546
R1887 GNDA.n1034 GNDA.n1032 175.546
R1888 GNDA.n1042 GNDA.n438 175.546
R1889 GNDA.n1049 GNDA.n1044 175.546
R1890 GNDA.n1047 GNDA.n1046 175.546
R1891 GNDA.n512 GNDA.n511 175.546
R1892 GNDA.n509 GNDA.n489 175.546
R1893 GNDA.n505 GNDA.n504 175.546
R1894 GNDA.n502 GNDA.n492 175.546
R1895 GNDA.n498 GNDA.n497 175.546
R1896 GNDA.n537 GNDA.n477 175.546
R1897 GNDA.n533 GNDA.n477 175.546
R1898 GNDA.n533 GNDA.n479 175.546
R1899 GNDA.n529 GNDA.n479 175.546
R1900 GNDA.n529 GNDA.n527 175.546
R1901 GNDA.n527 GNDA.n526 175.546
R1902 GNDA.n526 GNDA.n481 175.546
R1903 GNDA.n522 GNDA.n481 175.546
R1904 GNDA.n522 GNDA.n483 175.546
R1905 GNDA.n518 GNDA.n483 175.546
R1906 GNDA.n518 GNDA.n486 175.546
R1907 GNDA.n618 GNDA.n594 175.546
R1908 GNDA.n616 GNDA.n595 175.546
R1909 GNDA.n609 GNDA.n608 175.546
R1910 GNDA.n606 GNDA.n600 175.546
R1911 GNDA.n627 GNDA.n626 175.546
R1912 GNDA.n1201 GNDA.n1183 175.546
R1913 GNDA.n1204 GNDA.n1184 175.546
R1914 GNDA.n1188 GNDA.n1187 175.546
R1915 GNDA.n1207 GNDA.n1189 175.546
R1916 GNDA.n1193 GNDA.n1192 175.546
R1917 GNDA.n1378 GNDA.n1218 175.546
R1918 GNDA.n1378 GNDA.n1216 175.546
R1919 GNDA.n1382 GNDA.n1216 175.546
R1920 GNDA.n1382 GNDA.n1214 175.546
R1921 GNDA.n1386 GNDA.n1214 175.546
R1922 GNDA.n1386 GNDA.n1200 175.546
R1923 GNDA.n1390 GNDA.n1200 175.546
R1924 GNDA.n1390 GNDA.n1198 175.546
R1925 GNDA.n1394 GNDA.n1198 175.546
R1926 GNDA.n1394 GNDA.n1196 175.546
R1927 GNDA.n1398 GNDA.n1196 175.546
R1928 GNDA.n1354 GNDA.n1228 175.546
R1929 GNDA.n1354 GNDA.n1226 175.546
R1930 GNDA.n1359 GNDA.n1226 175.546
R1931 GNDA.n1359 GNDA.n1224 175.546
R1932 GNDA.n1363 GNDA.n1224 175.546
R1933 GNDA.n1364 GNDA.n1363 175.546
R1934 GNDA.n1366 GNDA.n1364 175.546
R1935 GNDA.n1366 GNDA.n1222 175.546
R1936 GNDA.n1370 GNDA.n1222 175.546
R1937 GNDA.n1370 GNDA.n1220 175.546
R1938 GNDA.n1374 GNDA.n1220 175.546
R1939 GNDA.n1346 GNDA.n1230 175.546
R1940 GNDA.n1267 GNDA.n1259 175.546
R1941 GNDA.n1271 GNDA.n1269 175.546
R1942 GNDA.n1283 GNDA.n1256 175.546
R1943 GNDA.n1288 GNDA.n1285 175.546
R1944 GNDA.n1453 GNDA.n1451 175.546
R1945 GNDA.n1461 GNDA.n236 175.546
R1946 GNDA.n1465 GNDA.n1463 175.546
R1947 GNDA.n1476 GNDA.n232 175.546
R1948 GNDA.n1479 GNDA.n1478 175.546
R1949 GNDA.n320 GNDA.n286 175.546
R1950 GNDA.n318 GNDA.n287 175.546
R1951 GNDA.n310 GNDA.n309 175.546
R1952 GNDA.n307 GNDA.n294 175.546
R1953 GNDA.n378 GNDA.n261 175.546
R1954 GNDA.n385 GNDA.n259 175.546
R1955 GNDA.n389 GNDA.n387 175.546
R1956 GNDA.n393 GNDA.n257 175.546
R1957 GNDA.n397 GNDA.n395 175.546
R1958 GNDA.n401 GNDA.n255 175.546
R1959 GNDA.n404 GNDA.n403 175.546
R1960 GNDA.n425 GNDA.n230 175.546
R1961 GNDA.n425 GNDA.n246 175.546
R1962 GNDA.n421 GNDA.n246 175.546
R1963 GNDA.n421 GNDA.n418 175.546
R1964 GNDA.n418 GNDA.n417 175.546
R1965 GNDA.n417 GNDA.n248 175.546
R1966 GNDA.n413 GNDA.n248 175.546
R1967 GNDA.n413 GNDA.n250 175.546
R1968 GNDA.n409 GNDA.n250 175.546
R1969 GNDA.n409 GNDA.n252 175.546
R1970 GNDA.n405 GNDA.n252 175.546
R1971 GNDA.n1683 GNDA.n1565 163.333
R1972 GNDA.n1173 GNDA.n1063 163.333
R1973 GNDA.n721 GNDA.n647 163.333
R1974 GNDA.n1887 GNDA.n152 163.333
R1975 GNDA.n889 GNDA.n887 163.333
R1976 GNDA.n621 GNDA.n471 163.333
R1977 GNDA.n1343 GNDA.n1233 163.333
R1978 GNDA.n325 GNDA.n323 163.333
R1979 GNDA.n1801 GNDA.n1791 163.333
R1980 GNDA.n1683 GNDA.n1566 150
R1981 GNDA.n1601 GNDA.n1600 150
R1982 GNDA.n1615 GNDA.n1614 150
R1983 GNDA.n1620 GNDA.n1619 150
R1984 GNDA.n1681 GNDA.n1584 150
R1985 GNDA.n1677 GNDA.n1676 150
R1986 GNDA.n1673 GNDA.n1672 150
R1987 GNDA.n1669 GNDA.n1668 150
R1988 GNDA.n1665 GNDA.n1664 150
R1989 GNDA.n1661 GNDA.n1660 150
R1990 GNDA.n1657 GNDA.n1656 150
R1991 GNDA.n1653 GNDA.n1574 150
R1992 GNDA.n1650 GNDA.n1574 150
R1993 GNDA.n1636 GNDA.n1635 150
R1994 GNDA.n1640 GNDA.n1639 150
R1995 GNDA.n1644 GNDA.n1643 150
R1996 GNDA.n1648 GNDA.n1647 150
R1997 GNDA.n1173 GNDA.n1064 150
R1998 GNDA.n1095 GNDA.n1094 150
R1999 GNDA.n1106 GNDA.n1105 150
R2000 GNDA.n1111 GNDA.n1110 150
R2001 GNDA.n1171 GNDA.n1082 150
R2002 GNDA.n1167 GNDA.n1166 150
R2003 GNDA.n1163 GNDA.n1162 150
R2004 GNDA.n1159 GNDA.n1158 150
R2005 GNDA.n1155 GNDA.n1154 150
R2006 GNDA.n1151 GNDA.n1150 150
R2007 GNDA.n1147 GNDA.n1146 150
R2008 GNDA.n1143 GNDA.n1072 150
R2009 GNDA.n1140 GNDA.n1072 150
R2010 GNDA.n1126 GNDA.n1125 150
R2011 GNDA.n1130 GNDA.n1129 150
R2012 GNDA.n1134 GNDA.n1133 150
R2013 GNDA.n1138 GNDA.n1137 150
R2014 GNDA.n723 GNDA.n721 150
R2015 GNDA.n735 GNDA.n643 150
R2016 GNDA.n739 GNDA.n737 150
R2017 GNDA.n747 GNDA.n639 150
R2018 GNDA.n710 GNDA.n708 150
R2019 GNDA.n706 GNDA.n649 150
R2020 GNDA.n702 GNDA.n700 150
R2021 GNDA.n698 GNDA.n651 150
R2022 GNDA.n694 GNDA.n692 150
R2023 GNDA.n690 GNDA.n653 150
R2024 GNDA.n686 GNDA.n684 150
R2025 GNDA.n682 GNDA.n655 150
R2026 GNDA.n678 GNDA.n655 150
R2027 GNDA.n665 GNDA.n663 150
R2028 GNDA.n669 GNDA.n659 150
R2029 GNDA.n672 GNDA.n671 150
R2030 GNDA.n676 GNDA.n675 150
R2031 GNDA.n1887 GNDA.n153 150
R2032 GNDA.n188 GNDA.n187 150
R2033 GNDA.n1819 GNDA.n1818 150
R2034 GNDA.n1824 GNDA.n1823 150
R2035 GNDA.n1885 GNDA.n171 150
R2036 GNDA.n1881 GNDA.n1880 150
R2037 GNDA.n1877 GNDA.n1876 150
R2038 GNDA.n1873 GNDA.n1872 150
R2039 GNDA.n1869 GNDA.n1868 150
R2040 GNDA.n1865 GNDA.n1864 150
R2041 GNDA.n1861 GNDA.n1860 150
R2042 GNDA.n1857 GNDA.n161 150
R2043 GNDA.n1854 GNDA.n161 150
R2044 GNDA.n1840 GNDA.n1839 150
R2045 GNDA.n1844 GNDA.n1843 150
R2046 GNDA.n1848 GNDA.n1847 150
R2047 GNDA.n1852 GNDA.n1851 150
R2048 GNDA.n887 GNDA.n845 150
R2049 GNDA.n879 GNDA.n877 150
R2050 GNDA.n866 GNDA.n864 150
R2051 GNDA.n868 GNDA.n863 150
R2052 GNDA.n893 GNDA.n843 150
R2053 GNDA.n897 GNDA.n895 150
R2054 GNDA.n901 GNDA.n841 150
R2055 GNDA.n905 GNDA.n903 150
R2056 GNDA.n909 GNDA.n839 150
R2057 GNDA.n913 GNDA.n911 150
R2058 GNDA.n917 GNDA.n837 150
R2059 GNDA.n920 GNDA.n919 150
R2060 GNDA.n922 GNDA.n920 150
R2061 GNDA.n936 GNDA.n935 150
R2062 GNDA.n933 GNDA.n831 150
R2063 GNDA.n929 GNDA.n928 150
R2064 GNDA.n926 GNDA.n834 150
R2065 GNDA.n621 GNDA.n472 150
R2066 GNDA.n613 GNDA.n612 150
R2067 GNDA.n602 GNDA.n601 150
R2068 GNDA.n623 GNDA.n451 150
R2069 GNDA.n587 GNDA.n586 150
R2070 GNDA.n583 GNDA.n582 150
R2071 GNDA.n579 GNDA.n578 150
R2072 GNDA.n575 GNDA.n574 150
R2073 GNDA.n571 GNDA.n570 150
R2074 GNDA.n567 GNDA.n566 150
R2075 GNDA.n563 GNDA.n562 150
R2076 GNDA.n559 GNDA.n459 150
R2077 GNDA.n556 GNDA.n459 150
R2078 GNDA.n542 GNDA.n541 150
R2079 GNDA.n546 GNDA.n545 150
R2080 GNDA.n550 GNDA.n549 150
R2081 GNDA.n554 GNDA.n553 150
R2082 GNDA.n1343 GNDA.n1234 150
R2083 GNDA.n1264 GNDA.n1263 150
R2084 GNDA.n1275 GNDA.n1274 150
R2085 GNDA.n1280 GNDA.n1279 150
R2086 GNDA.n1341 GNDA.n1252 150
R2087 GNDA.n1337 GNDA.n1336 150
R2088 GNDA.n1333 GNDA.n1332 150
R2089 GNDA.n1329 GNDA.n1328 150
R2090 GNDA.n1325 GNDA.n1324 150
R2091 GNDA.n1321 GNDA.n1320 150
R2092 GNDA.n1317 GNDA.n1316 150
R2093 GNDA.n1313 GNDA.n1242 150
R2094 GNDA.n1310 GNDA.n1242 150
R2095 GNDA.n1296 GNDA.n1295 150
R2096 GNDA.n1300 GNDA.n1299 150
R2097 GNDA.n1304 GNDA.n1303 150
R2098 GNDA.n1308 GNDA.n1307 150
R2099 GNDA.n323 GNDA.n280 150
R2100 GNDA.n315 GNDA.n313 150
R2101 GNDA.n302 GNDA.n300 150
R2102 GNDA.n304 GNDA.n299 150
R2103 GNDA.n329 GNDA.n278 150
R2104 GNDA.n333 GNDA.n331 150
R2105 GNDA.n337 GNDA.n276 150
R2106 GNDA.n341 GNDA.n339 150
R2107 GNDA.n345 GNDA.n274 150
R2108 GNDA.n349 GNDA.n347 150
R2109 GNDA.n353 GNDA.n272 150
R2110 GNDA.n356 GNDA.n355 150
R2111 GNDA.n358 GNDA.n356 150
R2112 GNDA.n372 GNDA.n371 150
R2113 GNDA.n369 GNDA.n266 150
R2114 GNDA.n365 GNDA.n364 150
R2115 GNDA.n362 GNDA.n269 150
R2116 GNDA.n1801 GNDA.n1800 150
R2117 GNDA.n2026 GNDA.n13 150
R2118 GNDA.n2029 GNDA.n2028 150
R2119 GNDA.n2032 GNDA.n2031 150
R2120 GNDA.n1788 GNDA.n1787 150
R2121 GNDA.n1785 GNDA.n1726 150
R2122 GNDA.n1781 GNDA.n1779 150
R2123 GNDA.n1777 GNDA.n1728 150
R2124 GNDA.n1773 GNDA.n1771 150
R2125 GNDA.n1769 GNDA.n1730 150
R2126 GNDA.n1765 GNDA.n1763 150
R2127 GNDA.n1761 GNDA.n1732 150
R2128 GNDA.n1757 GNDA.n1732 150
R2129 GNDA.n1744 GNDA.n1742 150
R2130 GNDA.n1748 GNDA.n1736 150
R2131 GNDA.n1751 GNDA.n1750 150
R2132 GNDA.n1755 GNDA.n1754 150
R2133 GNDA.n1560 GNDA.n1559 145.964
R2134 GNDA.n1559 GNDA.n1558 145.964
R2135 GNDA.n1558 GNDA.n1508 145.964
R2136 GNDA.n1552 GNDA.n1508 145.964
R2137 GNDA.n1552 GNDA.n65 145.964
R2138 GNDA.n1514 GNDA.n66 145.964
R2139 GNDA.n1545 GNDA.n1514 145.964
R2140 GNDA.n1545 GNDA.n1544 145.964
R2141 GNDA.n1544 GNDA.n1543 145.964
R2142 GNDA.n1543 GNDA.n52 145.964
R2143 GNDA.n536 GNDA.n51 145.964
R2144 GNDA.n536 GNDA.n535 145.964
R2145 GNDA.n535 GNDA.n534 145.964
R2146 GNDA.n534 GNDA.n478 145.964
R2147 GNDA.n528 GNDA.n478 145.964
R2148 GNDA.n528 GNDA.n58 145.964
R2149 GNDA.n484 GNDA.n59 145.964
R2150 GNDA.n521 GNDA.n484 145.964
R2151 GNDA.n521 GNDA.n520 145.964
R2152 GNDA.n520 GNDA.n519 145.964
R2153 GNDA.n519 GNDA.n485 145.964
R2154 GNDA.n1350 GNDA.t22 145.964
R2155 GNDA.n1350 GNDA.n1227 145.964
R2156 GNDA.n1355 GNDA.n1227 145.964
R2157 GNDA.n1356 GNDA.n1355 145.964
R2158 GNDA.n1358 GNDA.n1356 145.964
R2159 GNDA.n1358 GNDA.n1357 145.964
R2160 GNDA.n1357 GNDA.n1211 145.964
R2161 GNDA.n1365 GNDA.n1212 145.964
R2162 GNDA.n1365 GNDA.n1221 145.964
R2163 GNDA.n1371 GNDA.n1221 145.964
R2164 GNDA.n1372 GNDA.n1371 145.964
R2165 GNDA.n1373 GNDA.n1372 145.964
R2166 GNDA.n1695 GNDA.n1694 144.701
R2167 GNDA.n1697 GNDA.n1696 144.701
R2168 GNDA.n1699 GNDA.n1698 144.701
R2169 GNDA.n1705 GNDA.n1704 144.701
R2170 GNDA.n1703 GNDA.n1702 144.701
R2171 GNDA.n1701 GNDA.n1700 144.701
R2172 GNDA.n138 GNDA.n137 144.701
R2173 GNDA.n146 GNDA.n145 144.701
R2174 GNDA.n144 GNDA.n143 144.701
R2175 GNDA.n142 GNDA.n141 144.701
R2176 GNDA.n2013 GNDA.n2012 133.517
R2177 GNDA.n947 GNDA.n946 133.517
R2178 GNDA.n1447 GNDA.n1445 126.782
R2179 GNDA.n1905 GNDA.n1903 126.782
R2180 GNDA.n757 GNDA.n633 126.782
R2181 GNDA.n1714 GNDA.n79 126.782
R2182 GNDA.n1022 GNDA.n1020 126.782
R2183 GNDA.n1180 GNDA.n244 126.782
R2184 GNDA.n1439 GNDA.n429 124.832
R2185 GNDA.n1987 GNDA.n77 124.832
R2186 GNDA.n1024 GNDA.n444 124.832
R2187 GNDA.n1907 GNDA.n131 124.832
R2188 GNDA.n1013 GNDA.n634 124.832
R2189 GNDA.n1561 GNDA.n200 124.832
R2190 GNDA.n537 GNDA.n475 124.832
R2191 GNDA.n1349 GNDA.n1228 124.832
R2192 GNDA.n1449 GNDA.n240 124.832
R2193 GNDA.n1505 GNDA.t6 122.189
R2194 GNDA.n1691 GNDA.t97 116.501
R2195 GNDA.n1711 GNDA.t92 116.501
R2196 GNDA.n1706 GNDA.t103 116.501
R2197 GNDA.n1900 GNDA.t109 116.501
R2198 GNDA.n1895 GNDA.t112 116.501
R2199 GNDA.n139 GNDA.t106 116.501
R2200 GNDA.n1501 GNDA.t8 116.073
R2201 GNDA.n1499 GNDA.t29 115.105
R2202 GNDA.n1498 GNDA.t82 114.635
R2203 GNDA.n1501 GNDA.t21 114.635
R2204 GNDA.n1 GNDA.n50 14.555
R2205 GNDA.n0 GNDA.n53 14.555
R2206 GNDA.t102 GNDA.n1717 101.942
R2207 GNDA.t85 GNDA.n66 98.9316
R2208 GNDA.t85 GNDA.n59 98.9316
R2209 GNDA.t85 GNDA.n1212 98.9316
R2210 GNDA.n1902 GNDA.n135 98.8538
R2211 GNDA.n1690 GNDA.n199 96.7943
R2212 GNDA.n2015 GNDA.n19 95.7646
R2213 GNDA.n1627 GNDA.n1626 92.6754
R2214 GNDA.n1893 GNDA.t111 90.616
R2215 GNDA.n1379 GNDA.n1217 88.5317
R2216 GNDA.n1380 GNDA.n1379 88.5317
R2217 GNDA.n1381 GNDA.n1380 88.5317
R2218 GNDA.n1381 GNDA.n1213 88.5317
R2219 GNDA.n1387 GNDA.n1213 88.5317
R2220 GNDA.n1389 GNDA.n1388 88.5317
R2221 GNDA.n1389 GNDA.n1197 88.5317
R2222 GNDA.n1395 GNDA.n1197 88.5317
R2223 GNDA.n1396 GNDA.n1395 88.5317
R2224 GNDA.n1397 GNDA.n1396 88.5317
R2225 GNDA.n1415 GNDA.n1414 88.5317
R2226 GNDA.n1414 GNDA.n1413 88.5317
R2227 GNDA.n1413 GNDA.n1403 88.5317
R2228 GNDA.n1407 GNDA.n1403 88.5317
R2229 GNDA.n1407 GNDA.n216 88.5317
R2230 GNDA.n1495 GNDA.n218 88.5317
R2231 GNDA.n1489 GNDA.n218 88.5317
R2232 GNDA.n1489 GNDA.n1488 88.5317
R2233 GNDA.n1488 GNDA.n1487 88.5317
R2234 GNDA.n1487 GNDA.n225 88.5317
R2235 GNDA.n427 GNDA.n426 88.5317
R2236 GNDA.n426 GNDA.n245 88.5317
R2237 GNDA.n420 GNDA.n245 88.5317
R2238 GNDA.n420 GNDA.n419 88.5317
R2239 GNDA.n419 GNDA.n56 88.5317
R2240 GNDA.n412 GNDA.n57 88.5317
R2241 GNDA.n412 GNDA.n411 88.5317
R2242 GNDA.n411 GNDA.n410 88.5317
R2243 GNDA.n410 GNDA.n251 88.5317
R2244 GNDA.n251 GNDA.n54 88.5317
R2245 GNDA.n2040 GNDA.t68 84.4377
R2246 GNDA.n217 GNDA.n213 84.306
R2247 GNDA.t1 GNDA.t5 82.3782
R2248 GNDA.t18 GNDA.t24 82.3782
R2249 GNDA.n1795 GNDA.t46 80.3188
R2250 GNDA.n1446 GNDA.n238 76.3222
R2251 GNDA.n1457 GNDA.n1456 76.3222
R2252 GNDA.n1458 GNDA.n234 76.3222
R2253 GNDA.n1469 GNDA.n1468 76.3222
R2254 GNDA.n1473 GNDA.n1472 76.3222
R2255 GNDA.n1470 GNDA.n229 76.3222
R2256 GNDA.n1439 GNDA.n1438 76.3222
R2257 GNDA.n1436 GNDA.n1182 76.3222
R2258 GNDA.n1432 GNDA.n1431 76.3222
R2259 GNDA.n1425 GNDA.n1186 76.3222
R2260 GNDA.n1424 GNDA.n1423 76.3222
R2261 GNDA.n1417 GNDA.n1191 76.3222
R2262 GNDA.n1177 GNDA.n1176 76.3222
R2263 GNDA.n1090 GNDA.n1089 76.3222
R2264 GNDA.n1100 GNDA.n1099 76.3222
R2265 GNDA.n1101 GNDA.n1087 76.3222
R2266 GNDA.n1116 GNDA.n1115 76.3222
R2267 GNDA.n1117 GNDA.n242 76.3222
R2268 GNDA.n1988 GNDA.n1987 76.3222
R2269 GNDA.n1983 GNDA.n75 76.3222
R2270 GNDA.n1980 GNDA.n74 76.3222
R2271 GNDA.n1976 GNDA.n73 76.3222
R2272 GNDA.n1972 GNDA.n72 76.3222
R2273 GNDA.n1968 GNDA.n71 76.3222
R2274 GNDA.n1904 GNDA.n129 76.3222
R2275 GNDA.n1915 GNDA.n1914 76.3222
R2276 GNDA.n1916 GNDA.n125 76.3222
R2277 GNDA.n1927 GNDA.n1926 76.3222
R2278 GNDA.n1930 GNDA.n1929 76.3222
R2279 GNDA.n1940 GNDA.n99 76.3222
R2280 GNDA.n1961 GNDA.n38 76.3222
R2281 GNDA.n1957 GNDA.n39 76.3222
R2282 GNDA.n1953 GNDA.n40 76.3222
R2283 GNDA.n1949 GNDA.n41 76.3222
R2284 GNDA.n1945 GNDA.n42 76.3222
R2285 GNDA.n1941 GNDA.n43 76.3222
R2286 GNDA.n761 GNDA.n760 76.3222
R2287 GNDA.n764 GNDA.n763 76.3222
R2288 GNDA.n769 GNDA.n768 76.3222
R2289 GNDA.n772 GNDA.n771 76.3222
R2290 GNDA.n777 GNDA.n776 76.3222
R2291 GNDA.n780 GNDA.n779 76.3222
R2292 GNDA.n787 GNDA.n786 76.3222
R2293 GNDA.n792 GNDA.n791 76.3222
R2294 GNDA.n793 GNDA.n784 76.3222
R2295 GNDA.n800 GNDA.n799 76.3222
R2296 GNDA.n804 GNDA.n782 76.3222
R2297 GNDA.n807 GNDA.n806 76.3222
R2298 GNDA.n1025 GNDA.n1024 76.3222
R2299 GNDA.n1028 GNDA.n1027 76.3222
R2300 GNDA.n1037 GNDA.n1036 76.3222
R2301 GNDA.n1040 GNDA.n1039 76.3222
R2302 GNDA.n1052 GNDA.n1051 76.3222
R2303 GNDA.n1055 GNDA.n1054 76.3222
R2304 GNDA.n718 GNDA.n716 76.3222
R2305 GNDA.n727 GNDA.n645 76.3222
R2306 GNDA.n732 GNDA.n729 76.3222
R2307 GNDA.n742 GNDA.n641 76.3222
R2308 GNDA.n743 GNDA.n636 76.3222
R2309 GNDA.n754 GNDA.n753 76.3222
R2310 GNDA.n1908 GNDA.n1907 76.3222
R2311 GNDA.n1911 GNDA.n1910 76.3222
R2312 GNDA.n1920 GNDA.n1919 76.3222
R2313 GNDA.n1923 GNDA.n1922 76.3222
R2314 GNDA.n1934 GNDA.n1933 76.3222
R2315 GNDA.n1937 GNDA.n1936 76.3222
R2316 GNDA.n118 GNDA.n33 76.3222
R2317 GNDA.n114 GNDA.n34 76.3222
R2318 GNDA.n110 GNDA.n35 76.3222
R2319 GNDA.n106 GNDA.n36 76.3222
R2320 GNDA.n102 GNDA.n37 76.3222
R2321 GNDA.n1992 GNDA.n1991 76.3222
R2322 GNDA.n2012 GNDA.n2011 76.3222
R2323 GNDA.n2007 GNDA.n25 76.3222
R2324 GNDA.n2005 GNDA.n2004 76.3222
R2325 GNDA.n2000 GNDA.n28 76.3222
R2326 GNDA.n1998 GNDA.n1997 76.3222
R2327 GNDA.n1993 GNDA.n31 76.3222
R2328 GNDA.n946 GNDA.n824 76.3222
R2329 GNDA.n953 GNDA.n952 76.3222
R2330 GNDA.n954 GNDA.n822 76.3222
R2331 GNDA.n961 GNDA.n960 76.3222
R2332 GNDA.n962 GNDA.n820 76.3222
R2333 GNDA.n969 GNDA.n968 76.3222
R2334 GNDA.n989 GNDA.n988 76.3222
R2335 GNDA.n984 GNDA.n813 76.3222
R2336 GNDA.n982 GNDA.n981 76.3222
R2337 GNDA.n977 GNDA.n816 76.3222
R2338 GNDA.n975 GNDA.n974 76.3222
R2339 GNDA.n970 GNDA.n819 76.3222
R2340 GNDA.n1013 GNDA.n1012 76.3222
R2341 GNDA.n1010 GNDA.n759 76.3222
R2342 GNDA.n1006 GNDA.n1005 76.3222
R2343 GNDA.n999 GNDA.n766 76.3222
R2344 GNDA.n998 GNDA.n997 76.3222
R2345 GNDA.n991 GNDA.n774 76.3222
R2346 GNDA.n850 GNDA.n849 76.3222
R2347 GNDA.n883 GNDA.n882 76.3222
R2348 GNDA.n874 GNDA.n855 76.3222
R2349 GNDA.n872 GNDA.n871 76.3222
R2350 GNDA.n857 GNDA.n826 76.3222
R2351 GNDA.n944 GNDA.n943 76.3222
R2352 GNDA.n968 GNDA.n967 76.3222
R2353 GNDA.n963 GNDA.n962 76.3222
R2354 GNDA.n960 GNDA.n959 76.3222
R2355 GNDA.n955 GNDA.n954 76.3222
R2356 GNDA.n952 GNDA.n951 76.3222
R2357 GNDA.n31 GNDA.n29 76.3222
R2358 GNDA.n1999 GNDA.n1998 76.3222
R2359 GNDA.n28 GNDA.n26 76.3222
R2360 GNDA.n2006 GNDA.n2005 76.3222
R2361 GNDA.n25 GNDA.n23 76.3222
R2362 GNDA.n81 GNDA.n80 76.3222
R2363 GNDA.n84 GNDA.n83 76.3222
R2364 GNDA.n87 GNDA.n86 76.3222
R2365 GNDA.n90 GNDA.n89 76.3222
R2366 GNDA.n93 GNDA.n92 76.3222
R2367 GNDA.n96 GNDA.n95 76.3222
R2368 GNDA.n1536 GNDA.n44 76.3222
R2369 GNDA.n1532 GNDA.n45 76.3222
R2370 GNDA.n1528 GNDA.n46 76.3222
R2371 GNDA.n1524 GNDA.n47 76.3222
R2372 GNDA.n1520 GNDA.n48 76.3222
R2373 GNDA.n1516 GNDA.n49 76.3222
R2374 GNDA.n1021 GNDA.n442 76.3222
R2375 GNDA.n1032 GNDA.n1031 76.3222
R2376 GNDA.n1033 GNDA.n438 76.3222
R2377 GNDA.n1044 GNDA.n1043 76.3222
R2378 GNDA.n1048 GNDA.n1047 76.3222
R2379 GNDA.n1045 GNDA.n433 76.3222
R2380 GNDA.n513 GNDA.n512 76.3222
R2381 GNDA.n510 GNDA.n509 76.3222
R2382 GNDA.n505 GNDA.n491 76.3222
R2383 GNDA.n503 GNDA.n502 76.3222
R2384 GNDA.n498 GNDA.n494 76.3222
R2385 GNDA.n496 GNDA.n495 76.3222
R2386 GNDA.n594 GNDA.n593 76.3222
R2387 GNDA.n617 GNDA.n616 76.3222
R2388 GNDA.n609 GNDA.n598 76.3222
R2389 GNDA.n607 GNDA.n606 76.3222
R2390 GNDA.n626 GNDA.n449 76.3222
R2391 GNDA.n631 GNDA.n446 76.3222
R2392 GNDA.n1202 GNDA.n1201 76.3222
R2393 GNDA.n1203 GNDA.n1184 76.3222
R2394 GNDA.n1205 GNDA.n1187 76.3222
R2395 GNDA.n1206 GNDA.n1189 76.3222
R2396 GNDA.n1208 GNDA.n1192 76.3222
R2397 GNDA.n1209 GNDA.n1194 76.3222
R2398 GNDA.n1347 GNDA.n1346 76.3222
R2399 GNDA.n1259 GNDA.n1258 76.3222
R2400 GNDA.n1269 GNDA.n1268 76.3222
R2401 GNDA.n1270 GNDA.n1256 76.3222
R2402 GNDA.n1285 GNDA.n1284 76.3222
R2403 GNDA.n1287 GNDA.n1286 76.3222
R2404 GNDA.n627 GNDA.n446 76.3222
R2405 GNDA.n600 GNDA.n449 76.3222
R2406 GNDA.n608 GNDA.n607 76.3222
R2407 GNDA.n598 GNDA.n595 76.3222
R2408 GNDA.n618 GNDA.n617 76.3222
R2409 GNDA.n593 GNDA.n592 76.3222
R2410 GNDA.n753 GNDA.n752 76.3222
R2411 GNDA.n744 GNDA.n743 76.3222
R2412 GNDA.n731 GNDA.n641 76.3222
R2413 GNDA.n729 GNDA.n728 76.3222
R2414 GNDA.n717 GNDA.n645 76.3222
R2415 GNDA.n716 GNDA.n715 76.3222
R2416 GNDA.n943 GNDA.n942 76.3222
R2417 GNDA.n858 GNDA.n857 76.3222
R2418 GNDA.n873 GNDA.n872 76.3222
R2419 GNDA.n855 GNDA.n851 76.3222
R2420 GNDA.n884 GNDA.n883 76.3222
R2421 GNDA.n849 GNDA.n848 76.3222
R2422 GNDA.n1519 GNDA.n49 76.3222
R2423 GNDA.n1523 GNDA.n48 76.3222
R2424 GNDA.n1527 GNDA.n47 76.3222
R2425 GNDA.n1531 GNDA.n46 76.3222
R2426 GNDA.n1535 GNDA.n45 76.3222
R2427 GNDA.n1538 GNDA.n44 76.3222
R2428 GNDA.n1944 GNDA.n43 76.3222
R2429 GNDA.n1948 GNDA.n42 76.3222
R2430 GNDA.n1952 GNDA.n41 76.3222
R2431 GNDA.n1956 GNDA.n40 76.3222
R2432 GNDA.n1960 GNDA.n39 76.3222
R2433 GNDA.n1964 GNDA.n38 76.3222
R2434 GNDA.n1991 GNDA.n32 76.3222
R2435 GNDA.n105 GNDA.n37 76.3222
R2436 GNDA.n109 GNDA.n36 76.3222
R2437 GNDA.n113 GNDA.n35 76.3222
R2438 GNDA.n117 GNDA.n34 76.3222
R2439 GNDA.n121 GNDA.n33 76.3222
R2440 GNDA.n1288 GNDA.n1287 76.3222
R2441 GNDA.n1284 GNDA.n1283 76.3222
R2442 GNDA.n1271 GNDA.n1270 76.3222
R2443 GNDA.n1268 GNDA.n1267 76.3222
R2444 GNDA.n1258 GNDA.n1230 76.3222
R2445 GNDA.n1348 GNDA.n1347 76.3222
R2446 GNDA.n497 GNDA.n496 76.3222
R2447 GNDA.n494 GNDA.n492 76.3222
R2448 GNDA.n504 GNDA.n503 76.3222
R2449 GNDA.n491 GNDA.n489 76.3222
R2450 GNDA.n511 GNDA.n510 76.3222
R2451 GNDA.n514 GNDA.n513 76.3222
R2452 GNDA.n806 GNDA.n805 76.3222
R2453 GNDA.n801 GNDA.n782 76.3222
R2454 GNDA.n799 GNDA.n798 76.3222
R2455 GNDA.n794 GNDA.n793 76.3222
R2456 GNDA.n791 GNDA.n790 76.3222
R2457 GNDA.n786 GNDA.n434 76.3222
R2458 GNDA.n819 GNDA.n817 76.3222
R2459 GNDA.n976 GNDA.n975 76.3222
R2460 GNDA.n816 GNDA.n814 76.3222
R2461 GNDA.n983 GNDA.n982 76.3222
R2462 GNDA.n813 GNDA.n811 76.3222
R2463 GNDA.n990 GNDA.n989 76.3222
R2464 GNDA.n1450 GNDA.n1449 76.3222
R2465 GNDA.n1453 GNDA.n1452 76.3222
R2466 GNDA.n1462 GNDA.n1461 76.3222
R2467 GNDA.n1465 GNDA.n1464 76.3222
R2468 GNDA.n1477 GNDA.n1476 76.3222
R2469 GNDA.n1480 GNDA.n1479 76.3222
R2470 GNDA.n286 GNDA.n285 76.3222
R2471 GNDA.n319 GNDA.n318 76.3222
R2472 GNDA.n310 GNDA.n291 76.3222
R2473 GNDA.n308 GNDA.n307 76.3222
R2474 GNDA.n293 GNDA.n261 76.3222
R2475 GNDA.n380 GNDA.n379 76.3222
R2476 GNDA.n386 GNDA.n385 76.3222
R2477 GNDA.n389 GNDA.n388 76.3222
R2478 GNDA.n394 GNDA.n393 76.3222
R2479 GNDA.n397 GNDA.n396 76.3222
R2480 GNDA.n402 GNDA.n401 76.3222
R2481 GNDA.n403 GNDA.n402 76.3222
R2482 GNDA.n396 GNDA.n255 76.3222
R2483 GNDA.n395 GNDA.n394 76.3222
R2484 GNDA.n388 GNDA.n257 76.3222
R2485 GNDA.n387 GNDA.n386 76.3222
R2486 GNDA.n379 GNDA.n378 76.3222
R2487 GNDA.n294 GNDA.n293 76.3222
R2488 GNDA.n309 GNDA.n308 76.3222
R2489 GNDA.n291 GNDA.n287 76.3222
R2490 GNDA.n320 GNDA.n319 76.3222
R2491 GNDA.n285 GNDA.n284 76.3222
R2492 GNDA.n1118 GNDA.n1117 76.3222
R2493 GNDA.n1115 GNDA.n1114 76.3222
R2494 GNDA.n1102 GNDA.n1101 76.3222
R2495 GNDA.n1099 GNDA.n1098 76.3222
R2496 GNDA.n1089 GNDA.n1061 76.3222
R2497 GNDA.n1178 GNDA.n1177 76.3222
R2498 GNDA.n1471 GNDA.n1470 76.3222
R2499 GNDA.n1474 GNDA.n1473 76.3222
R2500 GNDA.n1468 GNDA.n1467 76.3222
R2501 GNDA.n1459 GNDA.n1458 76.3222
R2502 GNDA.n1456 GNDA.n1455 76.3222
R2503 GNDA.n1447 GNDA.n1446 76.3222
R2504 GNDA.n1451 GNDA.n1450 76.3222
R2505 GNDA.n1452 GNDA.n236 76.3222
R2506 GNDA.n1463 GNDA.n1462 76.3222
R2507 GNDA.n1464 GNDA.n232 76.3222
R2508 GNDA.n1478 GNDA.n1477 76.3222
R2509 GNDA.n1481 GNDA.n1480 76.3222
R2510 GNDA.n779 GNDA.n778 76.3222
R2511 GNDA.n776 GNDA.n775 76.3222
R2512 GNDA.n771 GNDA.n770 76.3222
R2513 GNDA.n768 GNDA.n767 76.3222
R2514 GNDA.n763 GNDA.n762 76.3222
R2515 GNDA.n760 GNDA.n757 76.3222
R2516 GNDA.n1012 GNDA.n1011 76.3222
R2517 GNDA.n1007 GNDA.n759 76.3222
R2518 GNDA.n1005 GNDA.n1004 76.3222
R2519 GNDA.n1000 GNDA.n999 76.3222
R2520 GNDA.n997 GNDA.n996 76.3222
R2521 GNDA.n992 GNDA.n991 76.3222
R2522 GNDA.n1928 GNDA.n99 76.3222
R2523 GNDA.n1931 GNDA.n1930 76.3222
R2524 GNDA.n1926 GNDA.n1925 76.3222
R2525 GNDA.n1917 GNDA.n1916 76.3222
R2526 GNDA.n1914 GNDA.n1913 76.3222
R2527 GNDA.n1905 GNDA.n1904 76.3222
R2528 GNDA.n1909 GNDA.n1908 76.3222
R2529 GNDA.n1910 GNDA.n127 76.3222
R2530 GNDA.n1921 GNDA.n1920 76.3222
R2531 GNDA.n1922 GNDA.n123 76.3222
R2532 GNDA.n1935 GNDA.n1934 76.3222
R2533 GNDA.n1938 GNDA.n1937 76.3222
R2534 GNDA.n95 GNDA.n94 76.3222
R2535 GNDA.n92 GNDA.n91 76.3222
R2536 GNDA.n89 GNDA.n88 76.3222
R2537 GNDA.n86 GNDA.n85 76.3222
R2538 GNDA.n83 GNDA.n82 76.3222
R2539 GNDA.n80 GNDA.n79 76.3222
R2540 GNDA.n1988 GNDA.n76 76.3222
R2541 GNDA.n1981 GNDA.n75 76.3222
R2542 GNDA.n1977 GNDA.n74 76.3222
R2543 GNDA.n1973 GNDA.n73 76.3222
R2544 GNDA.n1969 GNDA.n72 76.3222
R2545 GNDA.n1965 GNDA.n71 76.3222
R2546 GNDA.n1046 GNDA.n1045 76.3222
R2547 GNDA.n1049 GNDA.n1048 76.3222
R2548 GNDA.n1043 GNDA.n1042 76.3222
R2549 GNDA.n1034 GNDA.n1033 76.3222
R2550 GNDA.n1031 GNDA.n1030 76.3222
R2551 GNDA.n1022 GNDA.n1021 76.3222
R2552 GNDA.n1026 GNDA.n1025 76.3222
R2553 GNDA.n1027 GNDA.n440 76.3222
R2554 GNDA.n1038 GNDA.n1037 76.3222
R2555 GNDA.n1039 GNDA.n436 76.3222
R2556 GNDA.n1053 GNDA.n1052 76.3222
R2557 GNDA.n1056 GNDA.n1055 76.3222
R2558 GNDA.n1209 GNDA.n1193 76.3222
R2559 GNDA.n1208 GNDA.n1207 76.3222
R2560 GNDA.n1206 GNDA.n1188 76.3222
R2561 GNDA.n1205 GNDA.n1204 76.3222
R2562 GNDA.n1203 GNDA.n1183 76.3222
R2563 GNDA.n1202 GNDA.n1180 76.3222
R2564 GNDA.n1438 GNDA.n1437 76.3222
R2565 GNDA.n1433 GNDA.n1182 76.3222
R2566 GNDA.n1431 GNDA.n1430 76.3222
R2567 GNDA.n1426 GNDA.n1425 76.3222
R2568 GNDA.n1423 GNDA.n1422 76.3222
R2569 GNDA.n1418 GNDA.n1417 76.3222
R2570 GNDA.n1650 GNDA.n1575 76.062
R2571 GNDA.n1648 GNDA.n1575 76.062
R2572 GNDA.n1140 GNDA.n1073 76.062
R2573 GNDA.n1138 GNDA.n1073 76.062
R2574 GNDA.n678 GNDA.n677 76.062
R2575 GNDA.n677 GNDA.n676 76.062
R2576 GNDA.n1854 GNDA.n162 76.062
R2577 GNDA.n1852 GNDA.n162 76.062
R2578 GNDA.n922 GNDA.n921 76.062
R2579 GNDA.n921 GNDA.n834 76.062
R2580 GNDA.n556 GNDA.n460 76.062
R2581 GNDA.n554 GNDA.n460 76.062
R2582 GNDA.n1310 GNDA.n1243 76.062
R2583 GNDA.n1308 GNDA.n1243 76.062
R2584 GNDA.n358 GNDA.n357 76.062
R2585 GNDA.n357 GNDA.n269 76.062
R2586 GNDA.n1757 GNDA.n1756 76.062
R2587 GNDA.n1756 GNDA.n1755 76.062
R2588 GNDA.n1668 GNDA.n1580 74.5978
R2589 GNDA.n1665 GNDA.n1580 74.5978
R2590 GNDA.n1158 GNDA.n1078 74.5978
R2591 GNDA.n1155 GNDA.n1078 74.5978
R2592 GNDA.n693 GNDA.n651 74.5978
R2593 GNDA.n694 GNDA.n693 74.5978
R2594 GNDA.n1872 GNDA.n167 74.5978
R2595 GNDA.n1869 GNDA.n167 74.5978
R2596 GNDA.n905 GNDA.n904 74.5978
R2597 GNDA.n904 GNDA.n839 74.5978
R2598 GNDA.n574 GNDA.n466 74.5978
R2599 GNDA.n571 GNDA.n466 74.5978
R2600 GNDA.n1328 GNDA.n1248 74.5978
R2601 GNDA.n1325 GNDA.n1248 74.5978
R2602 GNDA.n341 GNDA.n340 74.5978
R2603 GNDA.n340 GNDA.n274 74.5978
R2604 GNDA.n1772 GNDA.n1728 74.5978
R2605 GNDA.n1773 GNDA.n1772 74.5978
R2606 GNDA.n1794 GNDA.t48 74.1404
R2607 GNDA.n2038 GNDA.t66 70.0216
R2608 GNDA.t100 GNDA.n1579 65.8183
R2609 GNDA.t100 GNDA.n1578 65.8183
R2610 GNDA.t100 GNDA.n1577 65.8183
R2611 GNDA.t100 GNDA.n1576 65.8183
R2612 GNDA.t100 GNDA.n1572 65.8183
R2613 GNDA.t100 GNDA.n1570 65.8183
R2614 GNDA.t100 GNDA.n1568 65.8183
R2615 GNDA.t100 GNDA.n1682 65.8183
R2616 GNDA.t100 GNDA.n1583 65.8183
R2617 GNDA.t100 GNDA.n1582 65.8183
R2618 GNDA.t100 GNDA.n1581 65.8183
R2619 GNDA.t87 GNDA.n1077 65.8183
R2620 GNDA.t87 GNDA.n1076 65.8183
R2621 GNDA.t87 GNDA.n1075 65.8183
R2622 GNDA.t87 GNDA.n1074 65.8183
R2623 GNDA.t87 GNDA.n1070 65.8183
R2624 GNDA.t87 GNDA.n1068 65.8183
R2625 GNDA.t87 GNDA.n1066 65.8183
R2626 GNDA.t87 GNDA.n1172 65.8183
R2627 GNDA.t87 GNDA.n1081 65.8183
R2628 GNDA.t87 GNDA.n1080 65.8183
R2629 GNDA.t87 GNDA.n1079 65.8183
R2630 GNDA.n657 GNDA.t86 65.8183
R2631 GNDA.n670 GNDA.t86 65.8183
R2632 GNDA.n664 GNDA.t86 65.8183
R2633 GNDA.n662 GNDA.t86 65.8183
R2634 GNDA.n683 GNDA.t86 65.8183
R2635 GNDA.n685 GNDA.t86 65.8183
R2636 GNDA.n691 GNDA.t86 65.8183
R2637 GNDA.n709 GNDA.t86 65.8183
R2638 GNDA.n707 GNDA.t86 65.8183
R2639 GNDA.n701 GNDA.t86 65.8183
R2640 GNDA.n699 GNDA.t86 65.8183
R2641 GNDA.n748 GNDA.t86 65.8183
R2642 GNDA.n738 GNDA.t86 65.8183
R2643 GNDA.n736 GNDA.t86 65.8183
R2644 GNDA.n722 GNDA.t86 65.8183
R2645 GNDA.t89 GNDA.n166 65.8183
R2646 GNDA.t89 GNDA.n165 65.8183
R2647 GNDA.t89 GNDA.n164 65.8183
R2648 GNDA.t89 GNDA.n163 65.8183
R2649 GNDA.t89 GNDA.n159 65.8183
R2650 GNDA.t89 GNDA.n157 65.8183
R2651 GNDA.t89 GNDA.n155 65.8183
R2652 GNDA.t89 GNDA.n1886 65.8183
R2653 GNDA.t89 GNDA.n170 65.8183
R2654 GNDA.t89 GNDA.n169 65.8183
R2655 GNDA.t89 GNDA.n168 65.8183
R2656 GNDA.t89 GNDA.n160 65.8183
R2657 GNDA.t89 GNDA.n158 65.8183
R2658 GNDA.t89 GNDA.n156 65.8183
R2659 GNDA.t89 GNDA.n154 65.8183
R2660 GNDA.n927 GNDA.t93 65.8183
R2661 GNDA.n833 GNDA.t93 65.8183
R2662 GNDA.n934 GNDA.t93 65.8183
R2663 GNDA.n937 GNDA.t93 65.8183
R2664 GNDA.n918 GNDA.t93 65.8183
R2665 GNDA.n912 GNDA.t93 65.8183
R2666 GNDA.n910 GNDA.t93 65.8183
R2667 GNDA.n888 GNDA.t93 65.8183
R2668 GNDA.n894 GNDA.t93 65.8183
R2669 GNDA.n896 GNDA.t93 65.8183
R2670 GNDA.n902 GNDA.t93 65.8183
R2671 GNDA.n860 GNDA.t93 65.8183
R2672 GNDA.n867 GNDA.t93 65.8183
R2673 GNDA.n853 GNDA.t93 65.8183
R2674 GNDA.n878 GNDA.t93 65.8183
R2675 GNDA.t98 GNDA.n465 65.8183
R2676 GNDA.t98 GNDA.n464 65.8183
R2677 GNDA.t98 GNDA.n463 65.8183
R2678 GNDA.t98 GNDA.n462 65.8183
R2679 GNDA.t98 GNDA.n458 65.8183
R2680 GNDA.t98 GNDA.n456 65.8183
R2681 GNDA.t98 GNDA.n454 65.8183
R2682 GNDA.t98 GNDA.n470 65.8183
R2683 GNDA.t98 GNDA.n469 65.8183
R2684 GNDA.t98 GNDA.n468 65.8183
R2685 GNDA.t98 GNDA.n467 65.8183
R2686 GNDA.n622 GNDA.t98 65.8183
R2687 GNDA.t98 GNDA.n457 65.8183
R2688 GNDA.t98 GNDA.n455 65.8183
R2689 GNDA.t98 GNDA.n453 65.8183
R2690 GNDA.t99 GNDA.n1247 65.8183
R2691 GNDA.t99 GNDA.n1246 65.8183
R2692 GNDA.t99 GNDA.n1245 65.8183
R2693 GNDA.t99 GNDA.n1244 65.8183
R2694 GNDA.t99 GNDA.n1240 65.8183
R2695 GNDA.t99 GNDA.n1238 65.8183
R2696 GNDA.t99 GNDA.n1236 65.8183
R2697 GNDA.t99 GNDA.n1342 65.8183
R2698 GNDA.t99 GNDA.n1251 65.8183
R2699 GNDA.t99 GNDA.n1250 65.8183
R2700 GNDA.t99 GNDA.n1249 65.8183
R2701 GNDA.t99 GNDA.n1241 65.8183
R2702 GNDA.t99 GNDA.n1239 65.8183
R2703 GNDA.t99 GNDA.n1237 65.8183
R2704 GNDA.t99 GNDA.n1235 65.8183
R2705 GNDA.n363 GNDA.t94 65.8183
R2706 GNDA.n268 GNDA.t94 65.8183
R2707 GNDA.n370 GNDA.t94 65.8183
R2708 GNDA.n373 GNDA.t94 65.8183
R2709 GNDA.n354 GNDA.t94 65.8183
R2710 GNDA.n348 GNDA.t94 65.8183
R2711 GNDA.n346 GNDA.t94 65.8183
R2712 GNDA.n324 GNDA.t94 65.8183
R2713 GNDA.n330 GNDA.t94 65.8183
R2714 GNDA.n332 GNDA.t94 65.8183
R2715 GNDA.n338 GNDA.t94 65.8183
R2716 GNDA.n296 GNDA.t94 65.8183
R2717 GNDA.n303 GNDA.t94 65.8183
R2718 GNDA.n289 GNDA.t94 65.8183
R2719 GNDA.n314 GNDA.t94 65.8183
R2720 GNDA.t87 GNDA.n1071 65.8183
R2721 GNDA.t87 GNDA.n1069 65.8183
R2722 GNDA.t87 GNDA.n1067 65.8183
R2723 GNDA.t87 GNDA.n1065 65.8183
R2724 GNDA.n1734 GNDA.t84 65.8183
R2725 GNDA.n1749 GNDA.t84 65.8183
R2726 GNDA.n1743 GNDA.t84 65.8183
R2727 GNDA.n1741 GNDA.t84 65.8183
R2728 GNDA.n1762 GNDA.t84 65.8183
R2729 GNDA.n1764 GNDA.t84 65.8183
R2730 GNDA.n1770 GNDA.t84 65.8183
R2731 GNDA.n1724 GNDA.t84 65.8183
R2732 GNDA.n1786 GNDA.t84 65.8183
R2733 GNDA.n1780 GNDA.t84 65.8183
R2734 GNDA.n1778 GNDA.t84 65.8183
R2735 GNDA.n2033 GNDA.t84 65.8183
R2736 GNDA.n2030 GNDA.t84 65.8183
R2737 GNDA.n2027 GNDA.t84 65.8183
R2738 GNDA.n1792 GNDA.t84 65.8183
R2739 GNDA.t100 GNDA.n1573 65.8183
R2740 GNDA.t100 GNDA.n1571 65.8183
R2741 GNDA.t100 GNDA.n1569 65.8183
R2742 GNDA.t100 GNDA.n1567 65.8183
R2743 GNDA.t7 GNDA.t23 64.1794
R2744 GNDA.t23 GNDA.t4 64.1794
R2745 GNDA.t20 GNDA.t30 64.1794
R2746 GNDA.t40 GNDA.n1609 63.8432
R2747 GNDA.t56 GNDA.n2039 63.8432
R2748 GNDA.n1829 GNDA.t42 63.8432
R2749 GNDA.n1560 GNDA.n1507 61.6297
R2750 GNDA.n1 GNDA.t85 32.9056
R2751 GNDA.n0 GNDA.t85 32.9056
R2752 GNDA.t72 GNDA.n1594 59.7243
R2753 GNDA.n1796 GNDA.t58 59.7243
R2754 GNDA.t76 GNDA.n192 59.7243
R2755 GNDA.n182 GNDA.t13 58.6946
R2756 GNDA.t80 GNDA.n1813 58.6946
R2757 GNDA.t16 GNDA.n1830 58.6946
R2758 GNDA.n2016 GNDA.t30 58.2964
R2759 GNDA.n382 GNDA.n381 57.1945
R2760 GNDA.n381 GNDA.n259 57.1945
R2761 GNDA.n947 GNDA.n945 57.1945
R2762 GNDA.n2014 GNDA.n2013 57.1945
R2763 GNDA.t81 GNDA.t74 56.6352
R2764 GNDA.n1808 GNDA.t108 56.6352
R2765 GNDA.t62 GNDA.t19 56.6352
R2766 GNDA.n1894 GNDA.n148 55.6055
R2767 GNDA.t100 GNDA.n1580 55.2026
R2768 GNDA.t87 GNDA.n1078 55.2026
R2769 GNDA.n693 GNDA.t86 55.2026
R2770 GNDA.t89 GNDA.n167 55.2026
R2771 GNDA.n904 GNDA.t93 55.2026
R2772 GNDA.t98 GNDA.n466 55.2026
R2773 GNDA.t99 GNDA.n1248 55.2026
R2774 GNDA.n340 GNDA.t94 55.2026
R2775 GNDA.n1772 GNDA.t84 55.2026
R2776 GNDA.n1689 GNDA.t31 54.5757
R2777 GNDA.t26 GNDA.n1605 54.5757
R2778 GNDA.t27 GNDA.n1624 54.5757
R2779 GNDA.n1713 GNDA.n1712 54.5757
R2780 GNDA.n1806 GNDA.n1718 54.5757
R2781 GNDA.t100 GNDA.n1575 54.4705
R2782 GNDA.t87 GNDA.n1073 54.4705
R2783 GNDA.n677 GNDA.t86 54.4705
R2784 GNDA.t89 GNDA.n162 54.4705
R2785 GNDA.n921 GNDA.t93 54.4705
R2786 GNDA.t98 GNDA.n460 54.4705
R2787 GNDA.t99 GNDA.n1243 54.4705
R2788 GNDA.n357 GNDA.t94 54.4705
R2789 GNDA.n1756 GNDA.t84 54.4705
R2790 GNDA.n1796 GNDA.t70 53.546
R2791 GNDA.n1567 GNDA.n1566 53.3664
R2792 GNDA.n1601 GNDA.n1569 53.3664
R2793 GNDA.n1615 GNDA.n1571 53.3664
R2794 GNDA.n1620 GNDA.n1573 53.3664
R2795 GNDA.n1682 GNDA.n1565 53.3664
R2796 GNDA.n1584 GNDA.n1583 53.3664
R2797 GNDA.n1676 GNDA.n1582 53.3664
R2798 GNDA.n1672 GNDA.n1581 53.3664
R2799 GNDA.n1664 GNDA.n1568 53.3664
R2800 GNDA.n1660 GNDA.n1570 53.3664
R2801 GNDA.n1656 GNDA.n1572 53.3664
R2802 GNDA.n1635 GNDA.n1576 53.3664
R2803 GNDA.n1639 GNDA.n1577 53.3664
R2804 GNDA.n1643 GNDA.n1578 53.3664
R2805 GNDA.n1647 GNDA.n1579 53.3664
R2806 GNDA.n1644 GNDA.n1579 53.3664
R2807 GNDA.n1640 GNDA.n1578 53.3664
R2808 GNDA.n1636 GNDA.n1577 53.3664
R2809 GNDA.n1632 GNDA.n1576 53.3664
R2810 GNDA.n1653 GNDA.n1572 53.3664
R2811 GNDA.n1657 GNDA.n1570 53.3664
R2812 GNDA.n1661 GNDA.n1568 53.3664
R2813 GNDA.n1682 GNDA.n1681 53.3664
R2814 GNDA.n1677 GNDA.n1583 53.3664
R2815 GNDA.n1673 GNDA.n1582 53.3664
R2816 GNDA.n1669 GNDA.n1581 53.3664
R2817 GNDA.n1065 GNDA.n1064 53.3664
R2818 GNDA.n1095 GNDA.n1067 53.3664
R2819 GNDA.n1106 GNDA.n1069 53.3664
R2820 GNDA.n1111 GNDA.n1071 53.3664
R2821 GNDA.n1172 GNDA.n1063 53.3664
R2822 GNDA.n1082 GNDA.n1081 53.3664
R2823 GNDA.n1166 GNDA.n1080 53.3664
R2824 GNDA.n1162 GNDA.n1079 53.3664
R2825 GNDA.n1154 GNDA.n1066 53.3664
R2826 GNDA.n1150 GNDA.n1068 53.3664
R2827 GNDA.n1146 GNDA.n1070 53.3664
R2828 GNDA.n1125 GNDA.n1074 53.3664
R2829 GNDA.n1129 GNDA.n1075 53.3664
R2830 GNDA.n1133 GNDA.n1076 53.3664
R2831 GNDA.n1137 GNDA.n1077 53.3664
R2832 GNDA.n1134 GNDA.n1077 53.3664
R2833 GNDA.n1130 GNDA.n1076 53.3664
R2834 GNDA.n1126 GNDA.n1075 53.3664
R2835 GNDA.n1122 GNDA.n1074 53.3664
R2836 GNDA.n1143 GNDA.n1070 53.3664
R2837 GNDA.n1147 GNDA.n1068 53.3664
R2838 GNDA.n1151 GNDA.n1066 53.3664
R2839 GNDA.n1172 GNDA.n1171 53.3664
R2840 GNDA.n1167 GNDA.n1081 53.3664
R2841 GNDA.n1163 GNDA.n1080 53.3664
R2842 GNDA.n1159 GNDA.n1079 53.3664
R2843 GNDA.n723 GNDA.n722 53.3664
R2844 GNDA.n736 GNDA.n735 53.3664
R2845 GNDA.n739 GNDA.n738 53.3664
R2846 GNDA.n748 GNDA.n747 53.3664
R2847 GNDA.n709 GNDA.n647 53.3664
R2848 GNDA.n708 GNDA.n707 53.3664
R2849 GNDA.n701 GNDA.n649 53.3664
R2850 GNDA.n700 GNDA.n699 53.3664
R2851 GNDA.n692 GNDA.n691 53.3664
R2852 GNDA.n685 GNDA.n653 53.3664
R2853 GNDA.n684 GNDA.n683 53.3664
R2854 GNDA.n663 GNDA.n662 53.3664
R2855 GNDA.n664 GNDA.n659 53.3664
R2856 GNDA.n671 GNDA.n670 53.3664
R2857 GNDA.n675 GNDA.n657 53.3664
R2858 GNDA.n672 GNDA.n657 53.3664
R2859 GNDA.n670 GNDA.n669 53.3664
R2860 GNDA.n665 GNDA.n664 53.3664
R2861 GNDA.n662 GNDA.n638 53.3664
R2862 GNDA.n683 GNDA.n682 53.3664
R2863 GNDA.n686 GNDA.n685 53.3664
R2864 GNDA.n691 GNDA.n690 53.3664
R2865 GNDA.n710 GNDA.n709 53.3664
R2866 GNDA.n707 GNDA.n706 53.3664
R2867 GNDA.n702 GNDA.n701 53.3664
R2868 GNDA.n699 GNDA.n698 53.3664
R2869 GNDA.n749 GNDA.n748 53.3664
R2870 GNDA.n738 GNDA.n639 53.3664
R2871 GNDA.n737 GNDA.n736 53.3664
R2872 GNDA.n722 GNDA.n643 53.3664
R2873 GNDA.n154 GNDA.n153 53.3664
R2874 GNDA.n188 GNDA.n156 53.3664
R2875 GNDA.n1819 GNDA.n158 53.3664
R2876 GNDA.n1824 GNDA.n160 53.3664
R2877 GNDA.n1886 GNDA.n152 53.3664
R2878 GNDA.n171 GNDA.n170 53.3664
R2879 GNDA.n1880 GNDA.n169 53.3664
R2880 GNDA.n1876 GNDA.n168 53.3664
R2881 GNDA.n1868 GNDA.n155 53.3664
R2882 GNDA.n1864 GNDA.n157 53.3664
R2883 GNDA.n1860 GNDA.n159 53.3664
R2884 GNDA.n1839 GNDA.n163 53.3664
R2885 GNDA.n1843 GNDA.n164 53.3664
R2886 GNDA.n1847 GNDA.n165 53.3664
R2887 GNDA.n1851 GNDA.n166 53.3664
R2888 GNDA.n1848 GNDA.n166 53.3664
R2889 GNDA.n1844 GNDA.n165 53.3664
R2890 GNDA.n1840 GNDA.n164 53.3664
R2891 GNDA.n1836 GNDA.n163 53.3664
R2892 GNDA.n1857 GNDA.n159 53.3664
R2893 GNDA.n1861 GNDA.n157 53.3664
R2894 GNDA.n1865 GNDA.n155 53.3664
R2895 GNDA.n1886 GNDA.n1885 53.3664
R2896 GNDA.n1881 GNDA.n170 53.3664
R2897 GNDA.n1877 GNDA.n169 53.3664
R2898 GNDA.n1873 GNDA.n168 53.3664
R2899 GNDA.n1835 GNDA.n160 53.3664
R2900 GNDA.n1823 GNDA.n158 53.3664
R2901 GNDA.n1818 GNDA.n156 53.3664
R2902 GNDA.n187 GNDA.n154 53.3664
R2903 GNDA.n878 GNDA.n845 53.3664
R2904 GNDA.n877 GNDA.n853 53.3664
R2905 GNDA.n867 GNDA.n866 53.3664
R2906 GNDA.n863 GNDA.n860 53.3664
R2907 GNDA.n889 GNDA.n888 53.3664
R2908 GNDA.n894 GNDA.n893 53.3664
R2909 GNDA.n897 GNDA.n896 53.3664
R2910 GNDA.n902 GNDA.n901 53.3664
R2911 GNDA.n910 GNDA.n909 53.3664
R2912 GNDA.n913 GNDA.n912 53.3664
R2913 GNDA.n918 GNDA.n917 53.3664
R2914 GNDA.n937 GNDA.n936 53.3664
R2915 GNDA.n934 GNDA.n933 53.3664
R2916 GNDA.n929 GNDA.n833 53.3664
R2917 GNDA.n927 GNDA.n926 53.3664
R2918 GNDA.n928 GNDA.n927 53.3664
R2919 GNDA.n833 GNDA.n831 53.3664
R2920 GNDA.n935 GNDA.n934 53.3664
R2921 GNDA.n938 GNDA.n937 53.3664
R2922 GNDA.n919 GNDA.n918 53.3664
R2923 GNDA.n912 GNDA.n837 53.3664
R2924 GNDA.n911 GNDA.n910 53.3664
R2925 GNDA.n888 GNDA.n843 53.3664
R2926 GNDA.n895 GNDA.n894 53.3664
R2927 GNDA.n896 GNDA.n841 53.3664
R2928 GNDA.n903 GNDA.n902 53.3664
R2929 GNDA.n860 GNDA.n829 53.3664
R2930 GNDA.n868 GNDA.n867 53.3664
R2931 GNDA.n864 GNDA.n853 53.3664
R2932 GNDA.n879 GNDA.n878 53.3664
R2933 GNDA.n472 GNDA.n453 53.3664
R2934 GNDA.n612 GNDA.n455 53.3664
R2935 GNDA.n602 GNDA.n457 53.3664
R2936 GNDA.n623 GNDA.n622 53.3664
R2937 GNDA.n471 GNDA.n470 53.3664
R2938 GNDA.n586 GNDA.n469 53.3664
R2939 GNDA.n582 GNDA.n468 53.3664
R2940 GNDA.n578 GNDA.n467 53.3664
R2941 GNDA.n570 GNDA.n454 53.3664
R2942 GNDA.n566 GNDA.n456 53.3664
R2943 GNDA.n562 GNDA.n458 53.3664
R2944 GNDA.n541 GNDA.n462 53.3664
R2945 GNDA.n545 GNDA.n463 53.3664
R2946 GNDA.n549 GNDA.n464 53.3664
R2947 GNDA.n553 GNDA.n465 53.3664
R2948 GNDA.n550 GNDA.n465 53.3664
R2949 GNDA.n546 GNDA.n464 53.3664
R2950 GNDA.n542 GNDA.n463 53.3664
R2951 GNDA.n462 GNDA.n461 53.3664
R2952 GNDA.n559 GNDA.n458 53.3664
R2953 GNDA.n563 GNDA.n456 53.3664
R2954 GNDA.n567 GNDA.n454 53.3664
R2955 GNDA.n587 GNDA.n470 53.3664
R2956 GNDA.n583 GNDA.n469 53.3664
R2957 GNDA.n579 GNDA.n468 53.3664
R2958 GNDA.n575 GNDA.n467 53.3664
R2959 GNDA.n622 GNDA.n452 53.3664
R2960 GNDA.n457 GNDA.n451 53.3664
R2961 GNDA.n601 GNDA.n455 53.3664
R2962 GNDA.n613 GNDA.n453 53.3664
R2963 GNDA.n1235 GNDA.n1234 53.3664
R2964 GNDA.n1264 GNDA.n1237 53.3664
R2965 GNDA.n1275 GNDA.n1239 53.3664
R2966 GNDA.n1280 GNDA.n1241 53.3664
R2967 GNDA.n1342 GNDA.n1233 53.3664
R2968 GNDA.n1252 GNDA.n1251 53.3664
R2969 GNDA.n1336 GNDA.n1250 53.3664
R2970 GNDA.n1332 GNDA.n1249 53.3664
R2971 GNDA.n1324 GNDA.n1236 53.3664
R2972 GNDA.n1320 GNDA.n1238 53.3664
R2973 GNDA.n1316 GNDA.n1240 53.3664
R2974 GNDA.n1295 GNDA.n1244 53.3664
R2975 GNDA.n1299 GNDA.n1245 53.3664
R2976 GNDA.n1303 GNDA.n1246 53.3664
R2977 GNDA.n1307 GNDA.n1247 53.3664
R2978 GNDA.n1304 GNDA.n1247 53.3664
R2979 GNDA.n1300 GNDA.n1246 53.3664
R2980 GNDA.n1296 GNDA.n1245 53.3664
R2981 GNDA.n1292 GNDA.n1244 53.3664
R2982 GNDA.n1313 GNDA.n1240 53.3664
R2983 GNDA.n1317 GNDA.n1238 53.3664
R2984 GNDA.n1321 GNDA.n1236 53.3664
R2985 GNDA.n1342 GNDA.n1341 53.3664
R2986 GNDA.n1337 GNDA.n1251 53.3664
R2987 GNDA.n1333 GNDA.n1250 53.3664
R2988 GNDA.n1329 GNDA.n1249 53.3664
R2989 GNDA.n1291 GNDA.n1241 53.3664
R2990 GNDA.n1279 GNDA.n1239 53.3664
R2991 GNDA.n1274 GNDA.n1237 53.3664
R2992 GNDA.n1263 GNDA.n1235 53.3664
R2993 GNDA.n314 GNDA.n280 53.3664
R2994 GNDA.n313 GNDA.n289 53.3664
R2995 GNDA.n303 GNDA.n302 53.3664
R2996 GNDA.n299 GNDA.n296 53.3664
R2997 GNDA.n325 GNDA.n324 53.3664
R2998 GNDA.n330 GNDA.n329 53.3664
R2999 GNDA.n333 GNDA.n332 53.3664
R3000 GNDA.n338 GNDA.n337 53.3664
R3001 GNDA.n346 GNDA.n345 53.3664
R3002 GNDA.n349 GNDA.n348 53.3664
R3003 GNDA.n354 GNDA.n353 53.3664
R3004 GNDA.n373 GNDA.n372 53.3664
R3005 GNDA.n370 GNDA.n369 53.3664
R3006 GNDA.n365 GNDA.n268 53.3664
R3007 GNDA.n363 GNDA.n362 53.3664
R3008 GNDA.n364 GNDA.n363 53.3664
R3009 GNDA.n268 GNDA.n266 53.3664
R3010 GNDA.n371 GNDA.n370 53.3664
R3011 GNDA.n374 GNDA.n373 53.3664
R3012 GNDA.n355 GNDA.n354 53.3664
R3013 GNDA.n348 GNDA.n272 53.3664
R3014 GNDA.n347 GNDA.n346 53.3664
R3015 GNDA.n324 GNDA.n278 53.3664
R3016 GNDA.n331 GNDA.n330 53.3664
R3017 GNDA.n332 GNDA.n276 53.3664
R3018 GNDA.n339 GNDA.n338 53.3664
R3019 GNDA.n296 GNDA.n264 53.3664
R3020 GNDA.n304 GNDA.n303 53.3664
R3021 GNDA.n300 GNDA.n289 53.3664
R3022 GNDA.n315 GNDA.n314 53.3664
R3023 GNDA.n1121 GNDA.n1071 53.3664
R3024 GNDA.n1110 GNDA.n1069 53.3664
R3025 GNDA.n1105 GNDA.n1067 53.3664
R3026 GNDA.n1094 GNDA.n1065 53.3664
R3027 GNDA.n1800 GNDA.n1792 53.3664
R3028 GNDA.n2027 GNDA.n2026 53.3664
R3029 GNDA.n2030 GNDA.n2029 53.3664
R3030 GNDA.n2033 GNDA.n2032 53.3664
R3031 GNDA.n1791 GNDA.n1724 53.3664
R3032 GNDA.n1787 GNDA.n1786 53.3664
R3033 GNDA.n1780 GNDA.n1726 53.3664
R3034 GNDA.n1779 GNDA.n1778 53.3664
R3035 GNDA.n1771 GNDA.n1770 53.3664
R3036 GNDA.n1764 GNDA.n1730 53.3664
R3037 GNDA.n1763 GNDA.n1762 53.3664
R3038 GNDA.n1742 GNDA.n1741 53.3664
R3039 GNDA.n1743 GNDA.n1736 53.3664
R3040 GNDA.n1750 GNDA.n1749 53.3664
R3041 GNDA.n1754 GNDA.n1734 53.3664
R3042 GNDA.n1751 GNDA.n1734 53.3664
R3043 GNDA.n1749 GNDA.n1748 53.3664
R3044 GNDA.n1744 GNDA.n1743 53.3664
R3045 GNDA.n1741 GNDA.n10 53.3664
R3046 GNDA.n1762 GNDA.n1761 53.3664
R3047 GNDA.n1765 GNDA.n1764 53.3664
R3048 GNDA.n1770 GNDA.n1769 53.3664
R3049 GNDA.n1788 GNDA.n1724 53.3664
R3050 GNDA.n1786 GNDA.n1785 53.3664
R3051 GNDA.n1781 GNDA.n1780 53.3664
R3052 GNDA.n1778 GNDA.n1777 53.3664
R3053 GNDA.n2034 GNDA.n2033 53.3664
R3054 GNDA.n2031 GNDA.n2030 53.3664
R3055 GNDA.n2028 GNDA.n2027 53.3664
R3056 GNDA.n1792 GNDA.n13 53.3664
R3057 GNDA.n1631 GNDA.n1573 53.3664
R3058 GNDA.n1619 GNDA.n1571 53.3664
R3059 GNDA.n1614 GNDA.n1569 53.3664
R3060 GNDA.n1600 GNDA.n1567 53.3664
R3061 GNDA.n196 GNDA.n70 51.4866
R3062 GNDA.n1901 GNDA.n136 51.4866
R3063 GNDA.n1811 GNDA.n1810 51.0266
R3064 GNDA.n2039 GNDA.t44 49.4271
R3065 GNDA.n1713 GNDA.t15 48.3974
R3066 GNDA.n1990 GNDA.t85 47.6748
R3067 GNDA.t85 GNDA.n64 47.6748
R3068 GNDA.n148 GNDA.t35 47.3677
R3069 GNDA.t85 GNDA.n65 47.0333
R3070 GNDA.t85 GNDA.n58 47.0333
R3071 GNDA.t85 GNDA.n1211 47.0333
R3072 GNDA.n1607 GNDA.n195 46.9641
R3073 GNDA.t14 GNDA.t96 46.338
R3074 GNDA.t105 GNDA.t25 46.338
R3075 GNDA.n1388 GNDA.t85 46.2335
R3076 GNDA.t85 GNDA.n1495 46.2335
R3077 GNDA.t85 GNDA.n57 46.2335
R3078 GNDA.n1624 GNDA.t64 43.2488
R3079 GNDA.t44 GNDA.n2038 43.2488
R3080 GNDA.n1831 GNDA.t105 43.2488
R3081 GNDA.t85 GNDA.n1387 42.2987
R3082 GNDA.t85 GNDA.n216 42.2987
R3083 GNDA.t85 GNDA.n56 42.2987
R3084 GNDA.t9 GNDA.n2020 42.2191
R3085 GNDA.t15 GNDA.n70 41.1894
R3086 GNDA.t35 GNDA.n136 41.1894
R3087 GNDA.t85 GNDA.n22 40.6472
R3088 GNDA.n1607 GNDA.t37 40.4338
R3089 GNDA.n1607 GNDA.t39 40.4338
R3090 GNDA.t96 GNDA.n1593 39.1299
R3091 GNDA.t70 GNDA.n1794 39.1299
R3092 GNDA.n2022 GNDA.n2021 39.1299
R3093 GNDA.n182 GNDA.t50 39.1299
R3094 GNDA.n194 GNDA.t36 38.6076
R3095 GNDA.n194 GNDA.t34 38.6076
R3096 GNDA.n1593 GNDA.t31 38.1002
R3097 GNDA.n1606 GNDA.t26 38.1002
R3098 GNDA.n1806 GNDA.n1805 38.1002
R3099 GNDA.n1902 GNDA.n1901 38.1002
R3100 GNDA.n1717 GNDA.n196 37.0705
R3101 GNDA.t85 GNDA.t54 36.0408
R3102 GNDA.t78 GNDA.t85 36.0408
R3103 GNDA.n1808 GNDA.n1807 33.9813
R3104 GNDA.n1814 GNDA.t80 33.9813
R3105 GNDA.n1831 GNDA.t16 33.9813
R3106 GNDA.n1595 GNDA.t72 32.9516
R3107 GNDA.t58 GNDA.n1795 32.9516
R3108 GNDA.n193 GNDA.t76 32.9516
R3109 GNDA.t22 GNDA.t28 32.4369
R3110 GNDA.n1505 GNDA.n1504 32.3063
R3111 GNDA.n1610 GNDA.t40 28.8327
R3112 GNDA.n2040 GNDA.t56 28.8327
R3113 GNDA.t42 GNDA.n1828 28.8327
R3114 GNDA.t17 GNDA.n1893 27.803
R3115 GNDA.n192 GNDA.t11 27.803
R3116 GNDA.n1828 GNDA.t19 27.803
R3117 GNDA.n1651 GNDA.n1649 27.5561
R3118 GNDA.n1141 GNDA.n1139 27.5561
R3119 GNDA.n679 GNDA.n656 27.5561
R3120 GNDA.n1855 GNDA.n1853 27.5561
R3121 GNDA.n924 GNDA.n923 27.5561
R3122 GNDA.n557 GNDA.n555 27.5561
R3123 GNDA.n1311 GNDA.n1309 27.5561
R3124 GNDA.n360 GNDA.n359 27.5561
R3125 GNDA.n1758 GNDA.n1733 27.5561
R3126 GNDA.n1019 GNDA.n1 8.60107
R3127 GNDA.n1444 GNDA.n0 8.60107
R3128 GNDA.n1667 GNDA.n1666 26.6672
R3129 GNDA.n1157 GNDA.n1156 26.6672
R3130 GNDA.n696 GNDA.n695 26.6672
R3131 GNDA.n1871 GNDA.n1870 26.6672
R3132 GNDA.n907 GNDA.n906 26.6672
R3133 GNDA.n573 GNDA.n572 26.6672
R3134 GNDA.n1327 GNDA.n1326 26.6672
R3135 GNDA.n343 GNDA.n342 26.6672
R3136 GNDA.n1775 GNDA.n1774 26.6672
R3137 GNDA.t85 GNDA.t12 25.9496
R3138 GNDA.t83 GNDA.t64 25.7435
R3139 GNDA.t50 GNDA.t11 25.7435
R3140 GNDA.n1694 GNDA.t73 24.0005
R3141 GNDA.n1694 GNDA.t75 24.0005
R3142 GNDA.n1696 GNDA.t55 24.0005
R3143 GNDA.n1696 GNDA.t41 24.0005
R3144 GNDA.n1698 GNDA.t65 24.0005
R3145 GNDA.n1698 GNDA.t53 24.0005
R3146 GNDA.n1704 GNDA.t49 24.0005
R3147 GNDA.n1704 GNDA.t71 24.0005
R3148 GNDA.n1702 GNDA.t59 24.0005
R3149 GNDA.n1702 GNDA.t47 24.0005
R3150 GNDA.n1700 GNDA.t69 24.0005
R3151 GNDA.n1700 GNDA.t57 24.0005
R3152 GNDA.n137 GNDA.t45 24.0005
R3153 GNDA.n137 GNDA.t67 24.0005
R3154 GNDA.n145 GNDA.t61 24.0005
R3155 GNDA.n145 GNDA.t51 24.0005
R3156 GNDA.n143 GNDA.t77 24.0005
R3157 GNDA.n143 GNDA.t79 24.0005
R3158 GNDA.n141 GNDA.t63 24.0005
R3159 GNDA.n141 GNDA.t43 24.0005
R3160 GNDA.n1595 GNDA.t81 23.6841
R3161 GNDA.n1609 GNDA.t83 23.6841
R3162 GNDA.n1626 GNDA.t32 23.6841
R3163 GNDA.n1711 GNDA.n1710 23.1624
R3164 GNDA.n1707 GNDA.n1706 23.1624
R3165 GNDA.n1900 GNDA.n1899 23.1624
R3166 GNDA.n1896 GNDA.n1895 23.1624
R3167 GNDA.n140 GNDA.n139 23.1624
R3168 GNDA.n1692 GNDA.n1691 23.1624
R3169 GNDA.n1625 GNDA.t52 22.6544
R3170 GNDA.n1807 GNDA.t66 22.6544
R3171 GNDA.n1498 GNDA.n1497 21.0192
R3172 GNDA.n1608 GNDA.t85 20.5949
R3173 GNDA.t0 GNDA.n1608 20.5949
R3174 GNDA.n1712 GNDA.t32 20.5949
R3175 GNDA.n1894 GNDA.t17 20.5949
R3176 GNDA.n1812 GNDA.t2 20.5949
R3177 GNDA.t85 GNDA.n1812 20.5949
R3178 GNDA.t85 GNDA.n54 19.6741
R3179 GNDA.n222 GNDA.n221 18.5605
R3180 GNDA.n1805 GNDA.t48 18.5355
R3181 GNDA.t60 GNDA.n181 18.5355
R3182 GNDA GNDA.n1502 18.1546
R3183 GNDA.n1540 GNDA.n1539 17.455
R3184 GNDA.n516 GNDA.n515 17.455
R3185 GNDA.n1376 GNDA.n1375 17.455
R3186 GNDA.n1994 GNDA.n30 17.0672
R3187 GNDA.n971 GNDA.n818 17.0672
R3188 GNDA.n406 GNDA.n253 17.0672
R3189 GNDA.n809 GNDA.n243 16.7235
R3190 GNDA.n1016 GNDA.n98 16.7235
R3191 GNDA.n632 GNDA.n97 16.7235
R3192 GNDA.n1442 GNDA.n1058 16.7235
R3193 GNDA.n1634 GNDA.n1633 16.0005
R3194 GNDA.n1637 GNDA.n1634 16.0005
R3195 GNDA.n1638 GNDA.n1637 16.0005
R3196 GNDA.n1641 GNDA.n1638 16.0005
R3197 GNDA.n1642 GNDA.n1641 16.0005
R3198 GNDA.n1645 GNDA.n1642 16.0005
R3199 GNDA.n1646 GNDA.n1645 16.0005
R3200 GNDA.n1649 GNDA.n1646 16.0005
R3201 GNDA.n1666 GNDA.n1663 16.0005
R3202 GNDA.n1663 GNDA.n1662 16.0005
R3203 GNDA.n1662 GNDA.n1659 16.0005
R3204 GNDA.n1659 GNDA.n1658 16.0005
R3205 GNDA.n1658 GNDA.n1655 16.0005
R3206 GNDA.n1655 GNDA.n1654 16.0005
R3207 GNDA.n1654 GNDA.n1652 16.0005
R3208 GNDA.n1652 GNDA.n1651 16.0005
R3209 GNDA.n1680 GNDA.n1563 16.0005
R3210 GNDA.n1680 GNDA.n1679 16.0005
R3211 GNDA.n1679 GNDA.n1678 16.0005
R3212 GNDA.n1678 GNDA.n1675 16.0005
R3213 GNDA.n1675 GNDA.n1674 16.0005
R3214 GNDA.n1674 GNDA.n1671 16.0005
R3215 GNDA.n1671 GNDA.n1670 16.0005
R3216 GNDA.n1670 GNDA.n1667 16.0005
R3217 GNDA.n1124 GNDA.n1123 16.0005
R3218 GNDA.n1127 GNDA.n1124 16.0005
R3219 GNDA.n1128 GNDA.n1127 16.0005
R3220 GNDA.n1131 GNDA.n1128 16.0005
R3221 GNDA.n1132 GNDA.n1131 16.0005
R3222 GNDA.n1135 GNDA.n1132 16.0005
R3223 GNDA.n1136 GNDA.n1135 16.0005
R3224 GNDA.n1139 GNDA.n1136 16.0005
R3225 GNDA.n1156 GNDA.n1153 16.0005
R3226 GNDA.n1153 GNDA.n1152 16.0005
R3227 GNDA.n1152 GNDA.n1149 16.0005
R3228 GNDA.n1149 GNDA.n1148 16.0005
R3229 GNDA.n1148 GNDA.n1145 16.0005
R3230 GNDA.n1145 GNDA.n1144 16.0005
R3231 GNDA.n1144 GNDA.n1142 16.0005
R3232 GNDA.n1142 GNDA.n1141 16.0005
R3233 GNDA.n1170 GNDA.n1083 16.0005
R3234 GNDA.n1170 GNDA.n1169 16.0005
R3235 GNDA.n1169 GNDA.n1168 16.0005
R3236 GNDA.n1168 GNDA.n1165 16.0005
R3237 GNDA.n1165 GNDA.n1164 16.0005
R3238 GNDA.n1164 GNDA.n1161 16.0005
R3239 GNDA.n1161 GNDA.n1160 16.0005
R3240 GNDA.n1160 GNDA.n1157 16.0005
R3241 GNDA.n661 GNDA.n660 16.0005
R3242 GNDA.n666 GNDA.n661 16.0005
R3243 GNDA.n667 GNDA.n666 16.0005
R3244 GNDA.n668 GNDA.n667 16.0005
R3245 GNDA.n668 GNDA.n658 16.0005
R3246 GNDA.n673 GNDA.n658 16.0005
R3247 GNDA.n674 GNDA.n673 16.0005
R3248 GNDA.n674 GNDA.n656 16.0005
R3249 GNDA.n695 GNDA.n652 16.0005
R3250 GNDA.n689 GNDA.n652 16.0005
R3251 GNDA.n689 GNDA.n688 16.0005
R3252 GNDA.n688 GNDA.n687 16.0005
R3253 GNDA.n687 GNDA.n654 16.0005
R3254 GNDA.n681 GNDA.n654 16.0005
R3255 GNDA.n681 GNDA.n680 16.0005
R3256 GNDA.n680 GNDA.n679 16.0005
R3257 GNDA.n712 GNDA.n711 16.0005
R3258 GNDA.n711 GNDA.n648 16.0005
R3259 GNDA.n705 GNDA.n648 16.0005
R3260 GNDA.n705 GNDA.n704 16.0005
R3261 GNDA.n704 GNDA.n703 16.0005
R3262 GNDA.n703 GNDA.n650 16.0005
R3263 GNDA.n697 GNDA.n650 16.0005
R3264 GNDA.n697 GNDA.n696 16.0005
R3265 GNDA.n1838 GNDA.n1837 16.0005
R3266 GNDA.n1841 GNDA.n1838 16.0005
R3267 GNDA.n1842 GNDA.n1841 16.0005
R3268 GNDA.n1845 GNDA.n1842 16.0005
R3269 GNDA.n1846 GNDA.n1845 16.0005
R3270 GNDA.n1849 GNDA.n1846 16.0005
R3271 GNDA.n1850 GNDA.n1849 16.0005
R3272 GNDA.n1853 GNDA.n1850 16.0005
R3273 GNDA.n1870 GNDA.n1867 16.0005
R3274 GNDA.n1867 GNDA.n1866 16.0005
R3275 GNDA.n1866 GNDA.n1863 16.0005
R3276 GNDA.n1863 GNDA.n1862 16.0005
R3277 GNDA.n1862 GNDA.n1859 16.0005
R3278 GNDA.n1859 GNDA.n1858 16.0005
R3279 GNDA.n1858 GNDA.n1856 16.0005
R3280 GNDA.n1856 GNDA.n1855 16.0005
R3281 GNDA.n1884 GNDA.n150 16.0005
R3282 GNDA.n1884 GNDA.n1883 16.0005
R3283 GNDA.n1883 GNDA.n1882 16.0005
R3284 GNDA.n1882 GNDA.n1879 16.0005
R3285 GNDA.n1879 GNDA.n1878 16.0005
R3286 GNDA.n1878 GNDA.n1875 16.0005
R3287 GNDA.n1875 GNDA.n1874 16.0005
R3288 GNDA.n1874 GNDA.n1871 16.0005
R3289 GNDA.n939 GNDA.n828 16.0005
R3290 GNDA.n830 GNDA.n828 16.0005
R3291 GNDA.n932 GNDA.n830 16.0005
R3292 GNDA.n932 GNDA.n931 16.0005
R3293 GNDA.n931 GNDA.n930 16.0005
R3294 GNDA.n930 GNDA.n832 16.0005
R3295 GNDA.n925 GNDA.n832 16.0005
R3296 GNDA.n925 GNDA.n924 16.0005
R3297 GNDA.n908 GNDA.n907 16.0005
R3298 GNDA.n908 GNDA.n838 16.0005
R3299 GNDA.n914 GNDA.n838 16.0005
R3300 GNDA.n915 GNDA.n914 16.0005
R3301 GNDA.n916 GNDA.n915 16.0005
R3302 GNDA.n916 GNDA.n836 16.0005
R3303 GNDA.n836 GNDA.n835 16.0005
R3304 GNDA.n923 GNDA.n835 16.0005
R3305 GNDA.n891 GNDA.n890 16.0005
R3306 GNDA.n892 GNDA.n891 16.0005
R3307 GNDA.n892 GNDA.n842 16.0005
R3308 GNDA.n898 GNDA.n842 16.0005
R3309 GNDA.n899 GNDA.n898 16.0005
R3310 GNDA.n900 GNDA.n899 16.0005
R3311 GNDA.n900 GNDA.n840 16.0005
R3312 GNDA.n906 GNDA.n840 16.0005
R3313 GNDA.n540 GNDA.n447 16.0005
R3314 GNDA.n543 GNDA.n540 16.0005
R3315 GNDA.n544 GNDA.n543 16.0005
R3316 GNDA.n547 GNDA.n544 16.0005
R3317 GNDA.n548 GNDA.n547 16.0005
R3318 GNDA.n551 GNDA.n548 16.0005
R3319 GNDA.n552 GNDA.n551 16.0005
R3320 GNDA.n555 GNDA.n552 16.0005
R3321 GNDA.n572 GNDA.n569 16.0005
R3322 GNDA.n569 GNDA.n568 16.0005
R3323 GNDA.n568 GNDA.n565 16.0005
R3324 GNDA.n565 GNDA.n564 16.0005
R3325 GNDA.n564 GNDA.n561 16.0005
R3326 GNDA.n561 GNDA.n560 16.0005
R3327 GNDA.n560 GNDA.n558 16.0005
R3328 GNDA.n558 GNDA.n557 16.0005
R3329 GNDA.n589 GNDA.n588 16.0005
R3330 GNDA.n588 GNDA.n585 16.0005
R3331 GNDA.n585 GNDA.n584 16.0005
R3332 GNDA.n584 GNDA.n581 16.0005
R3333 GNDA.n581 GNDA.n580 16.0005
R3334 GNDA.n580 GNDA.n577 16.0005
R3335 GNDA.n577 GNDA.n576 16.0005
R3336 GNDA.n576 GNDA.n573 16.0005
R3337 GNDA.n1294 GNDA.n1293 16.0005
R3338 GNDA.n1297 GNDA.n1294 16.0005
R3339 GNDA.n1298 GNDA.n1297 16.0005
R3340 GNDA.n1301 GNDA.n1298 16.0005
R3341 GNDA.n1302 GNDA.n1301 16.0005
R3342 GNDA.n1305 GNDA.n1302 16.0005
R3343 GNDA.n1306 GNDA.n1305 16.0005
R3344 GNDA.n1309 GNDA.n1306 16.0005
R3345 GNDA.n1326 GNDA.n1323 16.0005
R3346 GNDA.n1323 GNDA.n1322 16.0005
R3347 GNDA.n1322 GNDA.n1319 16.0005
R3348 GNDA.n1319 GNDA.n1318 16.0005
R3349 GNDA.n1318 GNDA.n1315 16.0005
R3350 GNDA.n1315 GNDA.n1314 16.0005
R3351 GNDA.n1314 GNDA.n1312 16.0005
R3352 GNDA.n1312 GNDA.n1311 16.0005
R3353 GNDA.n1340 GNDA.n1253 16.0005
R3354 GNDA.n1340 GNDA.n1339 16.0005
R3355 GNDA.n1339 GNDA.n1338 16.0005
R3356 GNDA.n1338 GNDA.n1335 16.0005
R3357 GNDA.n1335 GNDA.n1334 16.0005
R3358 GNDA.n1334 GNDA.n1331 16.0005
R3359 GNDA.n1331 GNDA.n1330 16.0005
R3360 GNDA.n1330 GNDA.n1327 16.0005
R3361 GNDA.n375 GNDA.n263 16.0005
R3362 GNDA.n265 GNDA.n263 16.0005
R3363 GNDA.n368 GNDA.n265 16.0005
R3364 GNDA.n368 GNDA.n367 16.0005
R3365 GNDA.n367 GNDA.n366 16.0005
R3366 GNDA.n366 GNDA.n267 16.0005
R3367 GNDA.n361 GNDA.n267 16.0005
R3368 GNDA.n361 GNDA.n360 16.0005
R3369 GNDA.n344 GNDA.n343 16.0005
R3370 GNDA.n344 GNDA.n273 16.0005
R3371 GNDA.n350 GNDA.n273 16.0005
R3372 GNDA.n351 GNDA.n350 16.0005
R3373 GNDA.n352 GNDA.n351 16.0005
R3374 GNDA.n352 GNDA.n271 16.0005
R3375 GNDA.n271 GNDA.n270 16.0005
R3376 GNDA.n359 GNDA.n270 16.0005
R3377 GNDA.n327 GNDA.n326 16.0005
R3378 GNDA.n328 GNDA.n327 16.0005
R3379 GNDA.n328 GNDA.n277 16.0005
R3380 GNDA.n334 GNDA.n277 16.0005
R3381 GNDA.n335 GNDA.n334 16.0005
R3382 GNDA.n336 GNDA.n335 16.0005
R3383 GNDA.n336 GNDA.n275 16.0005
R3384 GNDA.n342 GNDA.n275 16.0005
R3385 GNDA.n1740 GNDA.n1739 16.0005
R3386 GNDA.n1745 GNDA.n1740 16.0005
R3387 GNDA.n1746 GNDA.n1745 16.0005
R3388 GNDA.n1747 GNDA.n1746 16.0005
R3389 GNDA.n1747 GNDA.n1735 16.0005
R3390 GNDA.n1752 GNDA.n1735 16.0005
R3391 GNDA.n1753 GNDA.n1752 16.0005
R3392 GNDA.n1753 GNDA.n1733 16.0005
R3393 GNDA.n1774 GNDA.n1729 16.0005
R3394 GNDA.n1768 GNDA.n1729 16.0005
R3395 GNDA.n1768 GNDA.n1767 16.0005
R3396 GNDA.n1767 GNDA.n1766 16.0005
R3397 GNDA.n1766 GNDA.n1731 16.0005
R3398 GNDA.n1760 GNDA.n1731 16.0005
R3399 GNDA.n1760 GNDA.n1759 16.0005
R3400 GNDA.n1759 GNDA.n1758 16.0005
R3401 GNDA.n1790 GNDA.n1789 16.0005
R3402 GNDA.n1789 GNDA.n1725 16.0005
R3403 GNDA.n1784 GNDA.n1725 16.0005
R3404 GNDA.n1784 GNDA.n1783 16.0005
R3405 GNDA.n1783 GNDA.n1782 16.0005
R3406 GNDA.n1782 GNDA.n1727 16.0005
R3407 GNDA.n1776 GNDA.n1727 16.0005
R3408 GNDA.n1776 GNDA.n1775 16.0005
R3409 GNDA.n221 GNDA.n212 16.0005
R3410 GNDA.n1497 GNDA.n212 16.0005
R3411 GNDA.n1502 GNDA.n1500 15.4932
R3412 GNDA.t52 GNDA.t27 15.4463
R3413 GNDA.t13 GNDA.t60 15.4463
R3414 GNDA.n142 GNDA.n140 14.363
R3415 GNDA.n1710 GNDA.n1709 13.8005
R3416 GNDA.n1708 GNDA.n1707 13.8005
R3417 GNDA.n1899 GNDA.n1898 13.8005
R3418 GNDA.n1897 GNDA.n1896 13.8005
R3419 GNDA.n1693 GNDA.n1692 13.8005
R3420 GNDA.n1503 GNDA.n195 12.7542
R3421 GNDA.n1605 GNDA.t74 12.3572
R3422 GNDA.n2022 GNDA.t46 12.3572
R3423 GNDA.n1814 GNDA.t78 12.3572
R3424 GNDA.n1810 GNDA.n1809 12.2193
R3425 GNDA.n788 GNDA.n430 11.6369
R3426 GNDA.n789 GNDA.n788 11.6369
R3427 GNDA.n789 GNDA.n785 11.6369
R3428 GNDA.n795 GNDA.n785 11.6369
R3429 GNDA.n796 GNDA.n795 11.6369
R3430 GNDA.n797 GNDA.n796 11.6369
R3431 GNDA.n797 GNDA.n783 11.6369
R3432 GNDA.n802 GNDA.n783 11.6369
R3433 GNDA.n803 GNDA.n802 11.6369
R3434 GNDA.n803 GNDA.n781 11.6369
R3435 GNDA.n808 GNDA.n781 11.6369
R3436 GNDA.n1963 GNDA.n1962 11.6369
R3437 GNDA.n1962 GNDA.n1959 11.6369
R3438 GNDA.n1959 GNDA.n1958 11.6369
R3439 GNDA.n1958 GNDA.n1955 11.6369
R3440 GNDA.n1955 GNDA.n1954 11.6369
R3441 GNDA.n1954 GNDA.n1951 11.6369
R3442 GNDA.n1951 GNDA.n1950 11.6369
R3443 GNDA.n1950 GNDA.n1947 11.6369
R3444 GNDA.n1947 GNDA.n1946 11.6369
R3445 GNDA.n1946 GNDA.n1943 11.6369
R3446 GNDA.n1943 GNDA.n1942 11.6369
R3447 GNDA.n120 GNDA.n119 11.6369
R3448 GNDA.n119 GNDA.n116 11.6369
R3449 GNDA.n116 GNDA.n115 11.6369
R3450 GNDA.n115 GNDA.n112 11.6369
R3451 GNDA.n112 GNDA.n111 11.6369
R3452 GNDA.n111 GNDA.n108 11.6369
R3453 GNDA.n108 GNDA.n107 11.6369
R3454 GNDA.n107 GNDA.n104 11.6369
R3455 GNDA.n104 GNDA.n103 11.6369
R3456 GNDA.n103 GNDA.n101 11.6369
R3457 GNDA.n101 GNDA.n30 11.6369
R3458 GNDA.n2010 GNDA.n2009 11.6369
R3459 GNDA.n2009 GNDA.n2008 11.6369
R3460 GNDA.n2008 GNDA.n24 11.6369
R3461 GNDA.n2003 GNDA.n24 11.6369
R3462 GNDA.n2003 GNDA.n2002 11.6369
R3463 GNDA.n2002 GNDA.n2001 11.6369
R3464 GNDA.n2001 GNDA.n27 11.6369
R3465 GNDA.n1996 GNDA.n27 11.6369
R3466 GNDA.n1996 GNDA.n1995 11.6369
R3467 GNDA.n1995 GNDA.n1994 11.6369
R3468 GNDA.n987 GNDA.n810 11.6369
R3469 GNDA.n987 GNDA.n986 11.6369
R3470 GNDA.n986 GNDA.n985 11.6369
R3471 GNDA.n985 GNDA.n812 11.6369
R3472 GNDA.n980 GNDA.n812 11.6369
R3473 GNDA.n980 GNDA.n979 11.6369
R3474 GNDA.n979 GNDA.n978 11.6369
R3475 GNDA.n978 GNDA.n815 11.6369
R3476 GNDA.n973 GNDA.n815 11.6369
R3477 GNDA.n973 GNDA.n972 11.6369
R3478 GNDA.n972 GNDA.n971 11.6369
R3479 GNDA.n950 GNDA.n949 11.6369
R3480 GNDA.n950 GNDA.n823 11.6369
R3481 GNDA.n956 GNDA.n823 11.6369
R3482 GNDA.n957 GNDA.n956 11.6369
R3483 GNDA.n958 GNDA.n957 11.6369
R3484 GNDA.n958 GNDA.n821 11.6369
R3485 GNDA.n964 GNDA.n821 11.6369
R3486 GNDA.n965 GNDA.n964 11.6369
R3487 GNDA.n966 GNDA.n965 11.6369
R3488 GNDA.n966 GNDA.n818 11.6369
R3489 GNDA.n1539 GNDA.n1537 11.6369
R3490 GNDA.n1537 GNDA.n1534 11.6369
R3491 GNDA.n1534 GNDA.n1533 11.6369
R3492 GNDA.n1533 GNDA.n1530 11.6369
R3493 GNDA.n1530 GNDA.n1529 11.6369
R3494 GNDA.n1529 GNDA.n1526 11.6369
R3495 GNDA.n1526 GNDA.n1525 11.6369
R3496 GNDA.n1525 GNDA.n1522 11.6369
R3497 GNDA.n1522 GNDA.n1521 11.6369
R3498 GNDA.n1521 GNDA.n1518 11.6369
R3499 GNDA.n1518 GNDA.n1517 11.6369
R3500 GNDA.n1556 GNDA.n202 11.6369
R3501 GNDA.n1556 GNDA.n1555 11.6369
R3502 GNDA.n1555 GNDA.n1554 11.6369
R3503 GNDA.n1554 GNDA.n1510 11.6369
R3504 GNDA.n1549 GNDA.n1510 11.6369
R3505 GNDA.n1549 GNDA.n1548 11.6369
R3506 GNDA.n1548 GNDA.n1547 11.6369
R3507 GNDA.n1547 GNDA.n1512 11.6369
R3508 GNDA.n1541 GNDA.n1512 11.6369
R3509 GNDA.n1541 GNDA.n1540 11.6369
R3510 GNDA.n515 GNDA.n487 11.6369
R3511 GNDA.n488 GNDA.n487 11.6369
R3512 GNDA.n508 GNDA.n488 11.6369
R3513 GNDA.n508 GNDA.n507 11.6369
R3514 GNDA.n507 GNDA.n506 11.6369
R3515 GNDA.n506 GNDA.n490 11.6369
R3516 GNDA.n501 GNDA.n490 11.6369
R3517 GNDA.n501 GNDA.n500 11.6369
R3518 GNDA.n500 GNDA.n499 11.6369
R3519 GNDA.n499 GNDA.n493 11.6369
R3520 GNDA.n493 GNDA.n431 11.6369
R3521 GNDA.n532 GNDA.n476 11.6369
R3522 GNDA.n532 GNDA.n531 11.6369
R3523 GNDA.n531 GNDA.n530 11.6369
R3524 GNDA.n530 GNDA.n480 11.6369
R3525 GNDA.n525 GNDA.n480 11.6369
R3526 GNDA.n525 GNDA.n524 11.6369
R3527 GNDA.n524 GNDA.n523 11.6369
R3528 GNDA.n523 GNDA.n482 11.6369
R3529 GNDA.n517 GNDA.n482 11.6369
R3530 GNDA.n517 GNDA.n516 11.6369
R3531 GNDA.n1377 GNDA.n1376 11.6369
R3532 GNDA.n1377 GNDA.n1215 11.6369
R3533 GNDA.n1383 GNDA.n1215 11.6369
R3534 GNDA.n1384 GNDA.n1383 11.6369
R3535 GNDA.n1385 GNDA.n1384 11.6369
R3536 GNDA.n1385 GNDA.n1199 11.6369
R3537 GNDA.n1391 GNDA.n1199 11.6369
R3538 GNDA.n1392 GNDA.n1391 11.6369
R3539 GNDA.n1393 GNDA.n1392 11.6369
R3540 GNDA.n1393 GNDA.n1195 11.6369
R3541 GNDA.n1399 GNDA.n1195 11.6369
R3542 GNDA.n1353 GNDA.n1225 11.6369
R3543 GNDA.n1360 GNDA.n1225 11.6369
R3544 GNDA.n1361 GNDA.n1360 11.6369
R3545 GNDA.n1362 GNDA.n1361 11.6369
R3546 GNDA.n1362 GNDA.n1223 11.6369
R3547 GNDA.n1367 GNDA.n1223 11.6369
R3548 GNDA.n1368 GNDA.n1367 11.6369
R3549 GNDA.n1369 GNDA.n1368 11.6369
R3550 GNDA.n1369 GNDA.n1219 11.6369
R3551 GNDA.n1375 GNDA.n1219 11.6369
R3552 GNDA.n424 GNDA.n227 11.6369
R3553 GNDA.n424 GNDA.n423 11.6369
R3554 GNDA.n423 GNDA.n422 11.6369
R3555 GNDA.n422 GNDA.n247 11.6369
R3556 GNDA.n416 GNDA.n247 11.6369
R3557 GNDA.n416 GNDA.n415 11.6369
R3558 GNDA.n415 GNDA.n414 11.6369
R3559 GNDA.n414 GNDA.n249 11.6369
R3560 GNDA.n408 GNDA.n249 11.6369
R3561 GNDA.n408 GNDA.n407 11.6369
R3562 GNDA.n407 GNDA.n406 11.6369
R3563 GNDA.n384 GNDA.n258 11.6369
R3564 GNDA.n390 GNDA.n258 11.6369
R3565 GNDA.n391 GNDA.n390 11.6369
R3566 GNDA.n392 GNDA.n391 11.6369
R3567 GNDA.n392 GNDA.n256 11.6369
R3568 GNDA.n398 GNDA.n256 11.6369
R3569 GNDA.n399 GNDA.n398 11.6369
R3570 GNDA.n400 GNDA.n399 11.6369
R3571 GNDA.n400 GNDA.n254 11.6369
R3572 GNDA.n254 GNDA.n253 11.6369
R3573 GNDA.n1405 GNDA.n1402 11.6369
R3574 GNDA.n1411 GNDA.n1405 11.6369
R3575 GNDA.n1411 GNDA.n1410 11.6369
R3576 GNDA.n1410 GNDA.n1409 11.6369
R3577 GNDA.n1409 GNDA.n1406 11.6369
R3578 GNDA.n1493 GNDA.n1492 11.6369
R3579 GNDA.n1492 GNDA.n1491 11.6369
R3580 GNDA.n1491 GNDA.n223 11.6369
R3581 GNDA.n1485 GNDA.n223 11.6369
R3582 GNDA.n1485 GNDA.n1484 11.6369
R3583 GNDA.n1693 GNDA.n198 11.3792
R3584 GNDA.t54 GNDA.n1606 8.23827
R3585 GNDA.n2020 GNDA.t68 8.23827
R3586 GNDA.n1813 GNDA.t62 8.23827
R3587 GNDA.n1500 GNDA.n1499 7.56675
R3588 GNDA.n1502 GNDA.n1501 7.56675
R3589 GNDA.n1690 GNDA.n1689 7.20855
R3590 GNDA.n1594 GNDA.t14 7.20855
R3591 GNDA.n1610 GNDA.t0 7.20855
R3592 GNDA.n181 GNDA.t18 7.20855
R3593 GNDA.t33 GNDA.n2015 7.20855
R3594 GNDA.n1058 GNDA.n430 6.72373
R3595 GNDA.n1963 GNDA.n97 6.72373
R3596 GNDA.n120 GNDA.n98 6.72373
R3597 GNDA.n810 GNDA.n809 6.72373
R3598 GNDA.n1483 GNDA.n227 6.72373
R3599 GNDA.n1402 GNDA.n1400 6.72373
R3600 GNDA.n809 GNDA.n808 6.20656
R3601 GNDA.n1942 GNDA.n98 6.20656
R3602 GNDA.n1517 GNDA.n97 6.20656
R3603 GNDA.n1058 GNDA.n431 6.20656
R3604 GNDA.n1400 GNDA.n1399 6.20656
R3605 GNDA.n1484 GNDA.n1483 6.20656
R3606 GNDA.t38 GNDA.n199 6.17883
R3607 GNDA.t85 GNDA.t9 6.17883
R3608 GNDA.n1493 GNDA.n222 6.07727
R3609 GNDA.n2016 GNDA.t10 5.88357
R3610 GNDA.n1406 GNDA.n222 5.5601
R3611 GNDA.n1686 GNDA.n1563 5.51161
R3612 GNDA.n1083 GNDA.n1060 5.51161
R3613 GNDA.n713 GNDA.n712 5.51161
R3614 GNDA.n1890 GNDA.n150 5.51161
R3615 GNDA.n890 GNDA.n844 5.51161
R3616 GNDA.n590 GNDA.n589 5.51161
R3617 GNDA.n1253 GNDA.n1231 5.51161
R3618 GNDA.n326 GNDA.n279 5.51161
R3619 GNDA.n1790 GNDA.n1722 5.51161
R3620 GNDA.n591 GNDA.n539 5.1717
R3621 GNDA.n1352 GNDA.n1229 5.1717
R3622 GNDA.n1687 GNDA.n1562 5.1717
R3623 GNDA.t91 GNDA.t1 5.14911
R3624 GNDA.n2021 GNDA.t85 5.14911
R3625 GNDA.n172 GNDA.n21 4.9157
R3626 GNDA.n948 GNDA.n825 4.9157
R3627 GNDA.n383 GNDA.n260 4.9157
R3628 GNDA.n1448 GNDA.n239 4.26717
R3629 GNDA.n1454 GNDA.n239 4.26717
R3630 GNDA.n1454 GNDA.n237 4.26717
R3631 GNDA.n1460 GNDA.n237 4.26717
R3632 GNDA.n1460 GNDA.n235 4.26717
R3633 GNDA.n1466 GNDA.n235 4.26717
R3634 GNDA.n1466 GNDA.n233 4.26717
R3635 GNDA.n1475 GNDA.n233 4.26717
R3636 GNDA.n1475 GNDA.n231 4.26717
R3637 GNDA.n231 GNDA.n228 4.26717
R3638 GNDA.n1482 GNDA.n228 4.26717
R3639 GNDA.n1014 GNDA.n758 4.26717
R3640 GNDA.n1009 GNDA.n758 4.26717
R3641 GNDA.n1009 GNDA.n1008 4.26717
R3642 GNDA.n1008 GNDA.n765 4.26717
R3643 GNDA.n1003 GNDA.n765 4.26717
R3644 GNDA.n1003 GNDA.n1002 4.26717
R3645 GNDA.n1002 GNDA.n1001 4.26717
R3646 GNDA.n1001 GNDA.n773 4.26717
R3647 GNDA.n995 GNDA.n773 4.26717
R3648 GNDA.n995 GNDA.n994 4.26717
R3649 GNDA.n994 GNDA.n993 4.26717
R3650 GNDA.n1906 GNDA.n130 4.26717
R3651 GNDA.n1912 GNDA.n130 4.26717
R3652 GNDA.n1912 GNDA.n128 4.26717
R3653 GNDA.n1918 GNDA.n128 4.26717
R3654 GNDA.n1918 GNDA.n126 4.26717
R3655 GNDA.n1924 GNDA.n126 4.26717
R3656 GNDA.n1924 GNDA.n124 4.26717
R3657 GNDA.n1932 GNDA.n124 4.26717
R3658 GNDA.n1932 GNDA.n122 4.26717
R3659 GNDA.n122 GNDA.n100 4.26717
R3660 GNDA.n1939 GNDA.n100 4.26717
R3661 GNDA.n1986 GNDA.n1985 4.26717
R3662 GNDA.n1985 GNDA.n1984 4.26717
R3663 GNDA.n1984 GNDA.n1982 4.26717
R3664 GNDA.n1982 GNDA.n1979 4.26717
R3665 GNDA.n1979 GNDA.n1978 4.26717
R3666 GNDA.n1978 GNDA.n1975 4.26717
R3667 GNDA.n1975 GNDA.n1974 4.26717
R3668 GNDA.n1974 GNDA.n1971 4.26717
R3669 GNDA.n1971 GNDA.n1970 4.26717
R3670 GNDA.n1970 GNDA.n1967 4.26717
R3671 GNDA.n1967 GNDA.n1966 4.26717
R3672 GNDA.n1023 GNDA.n443 4.26717
R3673 GNDA.n1029 GNDA.n443 4.26717
R3674 GNDA.n1029 GNDA.n441 4.26717
R3675 GNDA.n1035 GNDA.n441 4.26717
R3676 GNDA.n1035 GNDA.n439 4.26717
R3677 GNDA.n1041 GNDA.n439 4.26717
R3678 GNDA.n1041 GNDA.n437 4.26717
R3679 GNDA.n1050 GNDA.n437 4.26717
R3680 GNDA.n1050 GNDA.n435 4.26717
R3681 GNDA.n435 GNDA.n432 4.26717
R3682 GNDA.n1057 GNDA.n432 4.26717
R3683 GNDA.n1440 GNDA.n1181 4.26717
R3684 GNDA.n1435 GNDA.n1181 4.26717
R3685 GNDA.n1435 GNDA.n1434 4.26717
R3686 GNDA.n1434 GNDA.n1185 4.26717
R3687 GNDA.n1429 GNDA.n1185 4.26717
R3688 GNDA.n1429 GNDA.n1428 4.26717
R3689 GNDA.n1428 GNDA.n1427 4.26717
R3690 GNDA.n1427 GNDA.n1190 4.26717
R3691 GNDA.n1421 GNDA.n1190 4.26717
R3692 GNDA.n1421 GNDA.n1420 4.26717
R3693 GNDA.n1420 GNDA.n1419 4.26717
R3694 GNDA.n1810 GNDA.n195 4.063
R3695 GNDA.n1483 GNDA.n1482 3.98272
R3696 GNDA.n993 GNDA.n809 3.98272
R3697 GNDA.n1939 GNDA.n98 3.98272
R3698 GNDA.n1966 GNDA.n97 3.98272
R3699 GNDA.n1058 GNDA.n1057 3.98272
R3700 GNDA.n1419 GNDA.n1400 3.98272
R3701 GNDA.n720 GNDA.n646 3.7893
R3702 GNDA.n726 GNDA.n724 3.7893
R3703 GNDA.n725 GNDA.n644 3.7893
R3704 GNDA.n734 GNDA.n733 3.7893
R3705 GNDA.n730 GNDA.n642 3.7893
R3706 GNDA.n745 GNDA.n640 3.7893
R3707 GNDA.n746 GNDA.n637 3.7893
R3708 GNDA.n751 GNDA.n750 3.7893
R3709 GNDA.n1888 GNDA.n151 3.7893
R3710 GNDA.n185 GNDA.n184 3.7893
R3711 GNDA.n190 GNDA.n186 3.7893
R3712 GNDA.n189 GNDA.n177 3.7893
R3713 GNDA.n1817 GNDA.n1816 3.7893
R3714 GNDA.n1826 GNDA.n1822 3.7893
R3715 GNDA.n1825 GNDA.n174 3.7893
R3716 GNDA.n1834 GNDA.n1833 3.7893
R3717 GNDA.n886 GNDA.n885 3.7893
R3718 GNDA.n881 GNDA.n847 3.7893
R3719 GNDA.n880 GNDA.n852 3.7893
R3720 GNDA.n876 GNDA.n875 3.7893
R3721 GNDA.n856 GNDA.n854 3.7893
R3722 GNDA.n869 GNDA.n859 3.7893
R3723 GNDA.n862 GNDA.n861 3.7893
R3724 GNDA.n941 GNDA.n827 3.7893
R3725 GNDA.n620 GNDA.n619 3.7893
R3726 GNDA.n615 GNDA.n474 3.7893
R3727 GNDA.n614 GNDA.n596 3.7893
R3728 GNDA.n611 GNDA.n610 3.7893
R3729 GNDA.n599 GNDA.n597 3.7893
R3730 GNDA.n604 GNDA.n450 3.7893
R3731 GNDA.n625 GNDA.n624 3.7893
R3732 GNDA.n628 GNDA.n448 3.7893
R3733 GNDA.n1344 GNDA.n1232 3.7893
R3734 GNDA.n1261 GNDA.n1260 3.7893
R3735 GNDA.n1266 GNDA.n1262 3.7893
R3736 GNDA.n1265 GNDA.n1257 3.7893
R3737 GNDA.n1273 GNDA.n1272 3.7893
R3738 GNDA.n1282 GNDA.n1278 3.7893
R3739 GNDA.n1281 GNDA.n1255 3.7893
R3740 GNDA.n1290 GNDA.n1289 3.7893
R3741 GNDA.n322 GNDA.n321 3.7893
R3742 GNDA.n317 GNDA.n282 3.7893
R3743 GNDA.n316 GNDA.n288 3.7893
R3744 GNDA.n312 GNDA.n311 3.7893
R3745 GNDA.n292 GNDA.n290 3.7893
R3746 GNDA.n305 GNDA.n295 3.7893
R3747 GNDA.n298 GNDA.n297 3.7893
R3748 GNDA.n377 GNDA.n262 3.7893
R3749 GNDA.n1174 GNDA.n1062 3.7893
R3750 GNDA.n1092 GNDA.n1091 3.7893
R3751 GNDA.n1097 GNDA.n1093 3.7893
R3752 GNDA.n1096 GNDA.n1088 3.7893
R3753 GNDA.n1104 GNDA.n1103 3.7893
R3754 GNDA.n1113 GNDA.n1109 3.7893
R3755 GNDA.n1112 GNDA.n1086 3.7893
R3756 GNDA.n1120 GNDA.n1119 3.7893
R3757 GNDA.n1802 GNDA.n1723 3.7893
R3758 GNDA.n1799 GNDA.n1798 3.7893
R3759 GNDA.n1793 GNDA.n14 3.7893
R3760 GNDA.n2025 GNDA.n2024 3.7893
R3761 GNDA.n12 GNDA.n11 3.7893
R3762 GNDA.n7 GNDA.n3 3.7893
R3763 GNDA.n2036 GNDA.n8 3.7893
R3764 GNDA.n2035 GNDA.n9 3.7893
R3765 GNDA.n1684 GNDA.n1564 3.7893
R3766 GNDA.n1598 GNDA.n1597 3.7893
R3767 GNDA.n1603 GNDA.n1599 3.7893
R3768 GNDA.n1602 GNDA.n1590 3.7893
R3769 GNDA.n1613 GNDA.n1612 3.7893
R3770 GNDA.n1622 GNDA.n1618 3.7893
R3771 GNDA.n1621 GNDA.n1587 3.7893
R3772 GNDA.n1630 GNDA.n1629 3.7893
R3773 GNDA.n1500 GNDA.n198 3.51962
R3774 GNDA.t5 GNDA.n1625 3.08966
R3775 GNDA.t24 GNDA.n180 3.08966
R3776 GNDA.t2 GNDA.n193 3.08966
R3777 GNDA.t25 GNDA.n1829 3.08966
R3778 GNDA.n1830 GNDA.n19 3.08966
R3779 GNDA.n741 GNDA 2.9189
R3780 GNDA.n1821 GNDA 2.9189
R3781 GNDA.n870 GNDA 2.9189
R3782 GNDA.n605 GNDA 2.9189
R3783 GNDA.n1277 GNDA 2.9189
R3784 GNDA.n306 GNDA 2.9189
R3785 GNDA.n1108 GNDA 2.9189
R3786 GNDA GNDA.n2042 2.9189
R3787 GNDA.n1617 GNDA 2.9189
R3788 GNDA.n714 GNDA.n445 2.6629
R3789 GNDA.n755 GNDA.n635 2.6629
R3790 GNDA.n1891 GNDA.n132 2.6629
R3791 GNDA.n173 GNDA.n172 2.6629
R3792 GNDA.n1015 GNDA.n756 2.6629
R3793 GNDA.n940 GNDA.n825 2.6629
R3794 GNDA.n630 GNDA.n629 2.6629
R3795 GNDA.n1254 GNDA.n1059 2.6629
R3796 GNDA.n283 GNDA.n241 2.6629
R3797 GNDA.n376 GNDA.n260 2.6629
R3798 GNDA.n1441 GNDA.n1179 2.6629
R3799 GNDA.n1085 GNDA.n1084 2.6629
R3800 GNDA.n1721 GNDA.n78 2.6629
R3801 GNDA.n1738 GNDA.n1737 2.6629
R3802 GNDA.n1586 GNDA.n1585 2.6629
R3803 GNDA.n714 GNDA.n713 2.4581
R3804 GNDA.n1015 GNDA.n755 2.4581
R3805 GNDA.n1891 GNDA.n1890 2.4581
R3806 GNDA.n844 GNDA.n756 2.4581
R3807 GNDA.n591 GNDA.n590 2.4581
R3808 GNDA.n630 GNDA.n445 2.4581
R3809 GNDA.n1231 GNDA.n1229 2.4581
R3810 GNDA.n1441 GNDA.n1059 2.4581
R3811 GNDA.n283 GNDA.n279 2.4581
R3812 GNDA.n1179 GNDA.n1060 2.4581
R3813 GNDA.n1084 GNDA.n241 2.4581
R3814 GNDA.n1722 GNDA.n1721 2.4581
R3815 GNDA.n1737 GNDA.n132 2.4581
R3816 GNDA.n1687 GNDA.n1686 2.4581
R3817 GNDA.n1585 GNDA.n78 2.4581
R3818 GNDA.n1448 GNDA.n241 2.18124
R3819 GNDA.n1015 GNDA.n1014 2.18124
R3820 GNDA.n1906 GNDA.n132 2.18124
R3821 GNDA.n1986 GNDA.n78 2.18124
R3822 GNDA.n1023 GNDA.n445 2.18124
R3823 GNDA.n1441 GNDA.n1440 2.18124
R3824 GNDA.n719 GNDA.n713 2.1509
R3825 GNDA.n1890 GNDA.n1889 2.1509
R3826 GNDA.n846 GNDA.n844 2.1509
R3827 GNDA.n590 GNDA.n473 2.1509
R3828 GNDA.n1345 GNDA.n1231 2.1509
R3829 GNDA.n281 GNDA.n279 2.1509
R3830 GNDA.n1175 GNDA.n1060 2.1509
R3831 GNDA.n1803 GNDA.n1722 2.1509
R3832 GNDA.n1686 GNDA.n1685 2.1509
R3833 GNDA.n1633 GNDA.n1586 2.13383
R3834 GNDA.n1123 GNDA.n1085 2.13383
R3835 GNDA.n660 GNDA.n635 2.13383
R3836 GNDA.n1837 GNDA.n173 2.13383
R3837 GNDA.n940 GNDA.n939 2.13383
R3838 GNDA.n629 GNDA.n447 2.13383
R3839 GNDA.n1293 GNDA.n1254 2.13383
R3840 GNDA.n376 GNDA.n375 2.13383
R3841 GNDA.n1739 GNDA.n1738 2.13383
R3842 GNDA.n1503 GNDA 2.09787
R3843 GNDA.n243 GNDA.n241 2.08643
R3844 GNDA.n1016 GNDA.n1015 2.08643
R3845 GNDA.n134 GNDA.n132 2.08643
R3846 GNDA.n1715 GNDA.n78 2.08643
R3847 GNDA.n632 GNDA.n445 2.08643
R3848 GNDA.n1442 GNDA.n1441 2.08643
R3849 GNDA.n1627 GNDA.t91 2.05994
R3850 GNDA.n1718 GNDA.t102 2.05994
R3851 GNDA.t108 GNDA.n135 2.05994
R3852 GNDA.n180 GNDA.t111 2.05994
R3853 GNDA.n1443 GNDA.n429 1.951
R3854 GNDA.n1716 GNDA.n77 1.951
R3855 GNDA.n1018 GNDA.n444 1.951
R3856 GNDA.n147 GNDA.n131 1.951
R3857 GNDA.n1017 GNDA.n634 1.951
R3858 GNDA.n203 GNDA.n200 1.951
R3859 GNDA.n538 GNDA.n475 1.951
R3860 GNDA.n1351 GNDA.n1349 1.951
R3861 GNDA.n428 GNDA.n240 1.951
R3862 GNDA.n751 GNDA.n635 1.9461
R3863 GNDA.n1833 GNDA.n173 1.9461
R3864 GNDA.n941 GNDA.n940 1.9461
R3865 GNDA.n629 GNDA.n628 1.9461
R3866 GNDA.n1289 GNDA.n1254 1.9461
R3867 GNDA.n377 GNDA.n376 1.9461
R3868 GNDA.n1119 GNDA.n1085 1.9461
R3869 GNDA.n1738 GNDA.n9 1.9461
R3870 GNDA.n1629 GNDA.n1586 1.9461
R3871 GNDA.n1499 GNDA.n1498 1.90675
R3872 GNDA.t85 GNDA.t28 1.62232
R3873 GNDA.n2010 GNDA.n21 1.52512
R3874 GNDA.n949 GNDA.n948 1.52512
R3875 GNDA.n384 GNDA.n383 1.52512
R3876 GNDA.n1562 GNDA.n202 1.42272
R3877 GNDA.n539 GNDA.n476 1.42272
R3878 GNDA.n1353 GNDA.n1352 1.42272
R3879 GNDA.n1898 GNDA.n1897 0.96925
R3880 GNDA.n1709 GNDA.n1708 0.96925
R3881 GNDA.n1811 GNDA.n194 0.914368
R3882 GNDA GNDA.n740 0.8709
R3883 GNDA GNDA.n1820 0.8709
R3884 GNDA.n865 GNDA 0.8709
R3885 GNDA GNDA.n603 0.8709
R3886 GNDA GNDA.n1276 0.8709
R3887 GNDA.n301 GNDA 0.8709
R3888 GNDA GNDA.n1107 0.8709
R3889 GNDA GNDA.n2 0.8709
R3890 GNDA GNDA.n1616 0.8709
R3891 GNDA.n720 GNDA.n719 0.8197
R3892 GNDA.n724 GNDA.n646 0.8197
R3893 GNDA.n726 GNDA.n725 0.8197
R3894 GNDA.n734 GNDA.n644 0.8197
R3895 GNDA.n733 GNDA.n642 0.8197
R3896 GNDA.n741 GNDA.n640 0.8197
R3897 GNDA.n746 GNDA.n745 0.8197
R3898 GNDA.n750 GNDA.n637 0.8197
R3899 GNDA.n1889 GNDA.n1888 0.8197
R3900 GNDA.n184 GNDA.n151 0.8197
R3901 GNDA.n186 GNDA.n185 0.8197
R3902 GNDA.n190 GNDA.n189 0.8197
R3903 GNDA.n1817 GNDA.n177 0.8197
R3904 GNDA.n1822 GNDA.n1821 0.8197
R3905 GNDA.n1826 GNDA.n1825 0.8197
R3906 GNDA.n1834 GNDA.n174 0.8197
R3907 GNDA.n886 GNDA.n846 0.8197
R3908 GNDA.n885 GNDA.n847 0.8197
R3909 GNDA.n881 GNDA.n880 0.8197
R3910 GNDA.n876 GNDA.n852 0.8197
R3911 GNDA.n875 GNDA.n854 0.8197
R3912 GNDA.n870 GNDA.n869 0.8197
R3913 GNDA.n862 GNDA.n859 0.8197
R3914 GNDA.n861 GNDA.n827 0.8197
R3915 GNDA.n620 GNDA.n473 0.8197
R3916 GNDA.n619 GNDA.n474 0.8197
R3917 GNDA.n615 GNDA.n614 0.8197
R3918 GNDA.n611 GNDA.n596 0.8197
R3919 GNDA.n610 GNDA.n597 0.8197
R3920 GNDA.n605 GNDA.n604 0.8197
R3921 GNDA.n624 GNDA.n450 0.8197
R3922 GNDA.n625 GNDA.n448 0.8197
R3923 GNDA.n1345 GNDA.n1344 0.8197
R3924 GNDA.n1260 GNDA.n1232 0.8197
R3925 GNDA.n1262 GNDA.n1261 0.8197
R3926 GNDA.n1266 GNDA.n1265 0.8197
R3927 GNDA.n1273 GNDA.n1257 0.8197
R3928 GNDA.n1278 GNDA.n1277 0.8197
R3929 GNDA.n1282 GNDA.n1281 0.8197
R3930 GNDA.n1290 GNDA.n1255 0.8197
R3931 GNDA.n322 GNDA.n281 0.8197
R3932 GNDA.n321 GNDA.n282 0.8197
R3933 GNDA.n317 GNDA.n316 0.8197
R3934 GNDA.n312 GNDA.n288 0.8197
R3935 GNDA.n311 GNDA.n290 0.8197
R3936 GNDA.n306 GNDA.n305 0.8197
R3937 GNDA.n298 GNDA.n295 0.8197
R3938 GNDA.n297 GNDA.n262 0.8197
R3939 GNDA.n1175 GNDA.n1174 0.8197
R3940 GNDA.n1091 GNDA.n1062 0.8197
R3941 GNDA.n1093 GNDA.n1092 0.8197
R3942 GNDA.n1097 GNDA.n1096 0.8197
R3943 GNDA.n1104 GNDA.n1088 0.8197
R3944 GNDA.n1109 GNDA.n1108 0.8197
R3945 GNDA.n1113 GNDA.n1112 0.8197
R3946 GNDA.n1120 GNDA.n1086 0.8197
R3947 GNDA.n1803 GNDA.n1802 0.8197
R3948 GNDA.n1799 GNDA.n1723 0.8197
R3949 GNDA.n1798 GNDA.n1793 0.8197
R3950 GNDA.n2025 GNDA.n14 0.8197
R3951 GNDA.n2024 GNDA.n12 0.8197
R3952 GNDA.n2042 GNDA.n3 0.8197
R3953 GNDA.n8 GNDA.n7 0.8197
R3954 GNDA.n2036 GNDA.n2035 0.8197
R3955 GNDA.n1685 GNDA.n1684 0.8197
R3956 GNDA.n1597 GNDA.n1564 0.8197
R3957 GNDA.n1599 GNDA.n1598 0.8197
R3958 GNDA.n1603 GNDA.n1602 0.8197
R3959 GNDA.n1613 GNDA.n1590 0.8197
R3960 GNDA.n1618 GNDA.n1617 0.8197
R3961 GNDA.n1622 GNDA.n1621 0.8197
R3962 GNDA.n1630 GNDA.n1587 0.8197
R3963 GNDA.n144 GNDA.n142 0.563
R3964 GNDA.n146 GNDA.n144 0.563
R3965 GNDA.n1897 GNDA.n146 0.563
R3966 GNDA.n1898 GNDA.n138 0.563
R3967 GNDA.n1701 GNDA.n138 0.563
R3968 GNDA.n1703 GNDA.n1701 0.563
R3969 GNDA.n1705 GNDA.n1703 0.563
R3970 GNDA.n1708 GNDA.n1705 0.563
R3971 GNDA.n1709 GNDA.n1699 0.563
R3972 GNDA.n1699 GNDA.n1697 0.563
R3973 GNDA.n1697 GNDA.n1695 0.563
R3974 GNDA.n1695 GNDA.n1693 0.563
R3975 GNDA.n730 GNDA 0.5125
R3976 GNDA.n1816 GNDA 0.5125
R3977 GNDA GNDA.n856 0.5125
R3978 GNDA GNDA.n599 0.5125
R3979 GNDA.n1272 GNDA 0.5125
R3980 GNDA GNDA.n292 0.5125
R3981 GNDA.n1103 GNDA 0.5125
R3982 GNDA.n11 GNDA 0.5125
R3983 GNDA.n1612 GNDA 0.5125
R3984 GNDA.n740 GNDA 0.3077
R3985 GNDA.n1820 GNDA 0.3077
R3986 GNDA.n865 GNDA 0.3077
R3987 GNDA.n603 GNDA 0.3077
R3988 GNDA.n1276 GNDA 0.3077
R3989 GNDA.n301 GNDA 0.3077
R3990 GNDA.n1107 GNDA 0.3077
R3991 GNDA GNDA.n2 0.3077
R3992 GNDA.n1616 GNDA 0.3077
R3993 GNDA.n1504 GNDA.n1503 0.276625
R3994 GNDA.n1504 GNDA.n198 0.22375
R3995 VB1_CUR_BIAS VB1_CUR_BIAS.n0 202.94
R3996 VB1_CUR_BIAS.n0 VB1_CUR_BIAS.t1 19.7005
R3997 VB1_CUR_BIAS.n0 VB1_CUR_BIAS.t0 19.7005
R3998 V_mir2.n9 V_mir2.n5 330.901
R3999 V_mir2.n4 V_mir2.n0 330.901
R4000 V_mir2.n20 V_mir2.n19 330.901
R4001 V_mir2.n16 V_mir2.t21 310.488
R4002 V_mir2.n6 V_mir2.t20 310.488
R4003 V_mir2.n1 V_mir2.t17 310.488
R4004 V_mir2.n12 V_mir2.t1 278.312
R4005 V_mir2.n12 V_mir2.n11 228.939
R4006 V_mir2.n13 V_mir2.n10 224.439
R4007 V_mir2.n18 V_mir2.t11 184.097
R4008 V_mir2.n8 V_mir2.t3 184.097
R4009 V_mir2.n3 V_mir2.t5 184.097
R4010 V_mir2.n17 V_mir2.n16 167.094
R4011 V_mir2.n7 V_mir2.n6 167.094
R4012 V_mir2.n2 V_mir2.n1 167.094
R4013 V_mir2.n9 V_mir2.n8 152
R4014 V_mir2.n4 V_mir2.n3 152
R4015 V_mir2.n19 V_mir2.n18 152
R4016 V_mir2.n16 V_mir2.t22 120.501
R4017 V_mir2.n17 V_mir2.t13 120.501
R4018 V_mir2.n6 V_mir2.t19 120.501
R4019 V_mir2.n7 V_mir2.t7 120.501
R4020 V_mir2.n1 V_mir2.t18 120.501
R4021 V_mir2.n2 V_mir2.t9 120.501
R4022 V_mir2.n11 V_mir2.t16 48.0005
R4023 V_mir2.n11 V_mir2.t2 48.0005
R4024 V_mir2.n10 V_mir2.t0 48.0005
R4025 V_mir2.n10 V_mir2.t15 48.0005
R4026 V_mir2.n18 V_mir2.n17 40.7027
R4027 V_mir2.n8 V_mir2.n7 40.7027
R4028 V_mir2.n3 V_mir2.n2 40.7027
R4029 V_mir2.n5 V_mir2.t4 39.4005
R4030 V_mir2.n5 V_mir2.t8 39.4005
R4031 V_mir2.n0 V_mir2.t6 39.4005
R4032 V_mir2.n0 V_mir2.t10 39.4005
R4033 V_mir2.n20 V_mir2.t12 39.4005
R4034 V_mir2.t14 V_mir2.n20 39.4005
R4035 V_mir2.n15 V_mir2.n4 15.8005
R4036 V_mir2.n19 V_mir2.n15 15.8005
R4037 V_mir2.n14 V_mir2.n9 9.3005
R4038 V_mir2.n13 V_mir2.n12 5.8755
R4039 V_mir2.n15 V_mir2.n14 4.5005
R4040 V_mir2.n14 V_mir2.n13 0.78175
R4041 VB2_CUR_BIAS.n2 VB2_CUR_BIAS.n0 146.482
R4042 VB2_CUR_BIAS.n6 VB2_CUR_BIAS.n5 145.232
R4043 VB2_CUR_BIAS.n4 VB2_CUR_BIAS.n3 145.232
R4044 VB2_CUR_BIAS.n2 VB2_CUR_BIAS.n1 145.232
R4045 VB2_CUR_BIAS VB2_CUR_BIAS.n6 29.688
R4046 VB2_CUR_BIAS.n5 VB2_CUR_BIAS.t1 24.0005
R4047 VB2_CUR_BIAS.n5 VB2_CUR_BIAS.t7 24.0005
R4048 VB2_CUR_BIAS.n3 VB2_CUR_BIAS.t2 24.0005
R4049 VB2_CUR_BIAS.n3 VB2_CUR_BIAS.t5 24.0005
R4050 VB2_CUR_BIAS.n1 VB2_CUR_BIAS.t0 24.0005
R4051 VB2_CUR_BIAS.n1 VB2_CUR_BIAS.t3 24.0005
R4052 VB2_CUR_BIAS.n0 VB2_CUR_BIAS.t6 24.0005
R4053 VB2_CUR_BIAS.n0 VB2_CUR_BIAS.t4 24.0005
R4054 VB2_CUR_BIAS.n4 VB2_CUR_BIAS.n2 7.563
R4055 VB2_CUR_BIAS.n6 VB2_CUR_BIAS.n4 1.2505
R4056 a_38570_n6504.t0 a_38570_n6504.t1 178.133
R4057 a_38690_n7778.t0 a_38690_n7778.t1 178.133
R4058 1st_Vout_1.n1 1st_Vout_1.t32 355.293
R4059 1st_Vout_1.n0 1st_Vout_1.t19 346.8
R4060 1st_Vout_1.n0 1st_Vout_1.n10 344.95
R4061 1st_Vout_1.n1 1st_Vout_1.n8 344.95
R4062 1st_Vout_1.n12 1st_Vout_1.n3 340.45
R4063 1st_Vout_1.n6 1st_Vout_1.t5 275.909
R4064 1st_Vout_1.n6 1st_Vout_1.n5 227.909
R4065 1st_Vout_1.n3 1st_Vout_1.n7 222.034
R4066 1st_Vout_1.n11 1st_Vout_1.t24 184.097
R4067 1st_Vout_1.n11 1st_Vout_1.t30 184.097
R4068 1st_Vout_1.n9 1st_Vout_1.t28 184.097
R4069 1st_Vout_1.n9 1st_Vout_1.t36 184.097
R4070 1st_Vout_1.n0 1st_Vout_1.n11 166.05
R4071 1st_Vout_1.n1 1st_Vout_1.n9 166.05
R4072 1st_Vout_1.n0 1st_Vout_1.n4 54.2759
R4073 1st_Vout_1.n7 1st_Vout_1.t1 48.0005
R4074 1st_Vout_1.n7 1st_Vout_1.t9 48.0005
R4075 1st_Vout_1.n5 1st_Vout_1.t6 48.0005
R4076 1st_Vout_1.n5 1st_Vout_1.t7 48.0005
R4077 1st_Vout_1.n10 1st_Vout_1.t4 39.4005
R4078 1st_Vout_1.n10 1st_Vout_1.t10 39.4005
R4079 1st_Vout_1.n8 1st_Vout_1.t2 39.4005
R4080 1st_Vout_1.n8 1st_Vout_1.t3 39.4005
R4081 1st_Vout_1.t0 1st_Vout_1.n12 39.4005
R4082 1st_Vout_1.n12 1st_Vout_1.t8 39.4005
R4083 1st_Vout_1.n3 1st_Vout_1.n1 5.28175
R4084 1st_Vout_1.n1 1st_Vout_1.n0 5.188
R4085 1st_Vout_1.n2 1st_Vout_1.t23 4.8295
R4086 1st_Vout_1.n2 1st_Vout_1.t11 4.8295
R4087 1st_Vout_1.n2 1st_Vout_1.t18 4.8295
R4088 1st_Vout_1.n2 1st_Vout_1.t27 4.8295
R4089 1st_Vout_1.n2 1st_Vout_1.t34 4.8295
R4090 1st_Vout_1.n2 1st_Vout_1.t20 4.8295
R4091 1st_Vout_1.n4 1st_Vout_1.t15 4.8295
R4092 1st_Vout_1.n4 1st_Vout_1.t25 4.8295
R4093 1st_Vout_1.n4 1st_Vout_1.t31 4.8295
R4094 1st_Vout_1.n2 1st_Vout_1.t21 4.5005
R4095 1st_Vout_1.n2 1st_Vout_1.t12 4.5005
R4096 1st_Vout_1.n2 1st_Vout_1.t16 4.5005
R4097 1st_Vout_1.n2 1st_Vout_1.t29 4.5005
R4098 1st_Vout_1.n2 1st_Vout_1.t33 4.5005
R4099 1st_Vout_1.n2 1st_Vout_1.t22 4.5005
R4100 1st_Vout_1.n4 1st_Vout_1.t14 4.5005
R4101 1st_Vout_1.n4 1st_Vout_1.t26 4.5005
R4102 1st_Vout_1.n4 1st_Vout_1.t17 4.5005
R4103 1st_Vout_1.n4 1st_Vout_1.t35 4.5005
R4104 1st_Vout_1.n4 1st_Vout_1.t13 4.5005
R4105 1st_Vout_1.n3 1st_Vout_1.n6 4.5005
R4106 1st_Vout_1.n4 1st_Vout_1.n2 3.1025
R4107 cap_res1.t0 cap_res1.t18 121.245
R4108 cap_res1.t1 cap_res1.t14 0.1603
R4109 cap_res1.t17 cap_res1.t16 0.1603
R4110 cap_res1.t3 cap_res1.t2 0.1603
R4111 cap_res1.t15 cap_res1.t13 0.1603
R4112 cap_res1.t11 cap_res1.t9 0.1603
R4113 cap_res1.n1 cap_res1.t19 0.159278
R4114 cap_res1.n2 cap_res1.t5 0.159278
R4115 cap_res1.n3 cap_res1.t10 0.159278
R4116 cap_res1.n4 cap_res1.t7 0.159278
R4117 cap_res1.n4 cap_res1.t4 0.1368
R4118 cap_res1.n4 cap_res1.t1 0.1368
R4119 cap_res1.n3 cap_res1.t8 0.1368
R4120 cap_res1.n3 cap_res1.t17 0.1368
R4121 cap_res1.n2 cap_res1.t12 0.1368
R4122 cap_res1.n2 cap_res1.t3 0.1368
R4123 cap_res1.n1 cap_res1.t6 0.1368
R4124 cap_res1.n1 cap_res1.t15 0.1368
R4125 cap_res1.n0 cap_res1.t20 0.1368
R4126 cap_res1.n0 cap_res1.t11 0.1368
R4127 cap_res1.t19 cap_res1.n0 0.00152174
R4128 cap_res1.t5 cap_res1.n1 0.00152174
R4129 cap_res1.t10 cap_res1.n2 0.00152174
R4130 cap_res1.t7 cap_res1.n3 0.00152174
R4131 cap_res1.t18 cap_res1.n4 0.00152174
R4132 V_CMFB_S4.n2 V_CMFB_S4.n0 150.451
R4133 V_CMFB_S4.n2 V_CMFB_S4.n1 140.201
R4134 V_CMFB_S4 V_CMFB_S4.n2 37.563
R4135 V_CMFB_S4.n1 V_CMFB_S4.t2 24.0005
R4136 V_CMFB_S4.n1 V_CMFB_S4.t1 24.0005
R4137 V_CMFB_S4.n0 V_CMFB_S4.t0 24.0005
R4138 V_CMFB_S4.n0 V_CMFB_S4.t3 24.0005
R4139 Vin+.n3 Vin+.n2 526.183
R4140 Vin+.n1 Vin+.n0 514.134
R4141 Vin+.n0 Vin+.t9 303.259
R4142 Vin+.n5 Vin+.n3 227.169
R4143 Vin+.n0 Vin+.t7 174.726
R4144 Vin+.n1 Vin+.t6 174.726
R4145 Vin+.n2 Vin+.t10 174.726
R4146 Vin+.n7 Vin+.n6 167.993
R4147 Vin+.n5 Vin+.n4 167.993
R4148 Vin+.t1 Vin+.n8 158.989
R4149 Vin+.n2 Vin+.n1 128.534
R4150 Vin+.n8 Vin+.t4 119.067
R4151 Vin+.n3 Vin+.t8 96.4005
R4152 Vin+.n8 Vin+.n7 35.0317
R4153 Vin+.n6 Vin+.t3 13.1338
R4154 Vin+.n6 Vin+.t5 13.1338
R4155 Vin+.n4 Vin+.t0 13.1338
R4156 Vin+.n4 Vin+.t2 13.1338
R4157 Vin+.n7 Vin+.n5 2.1255
R4158 V_p_1.n5 V_p_1.n3 263.933
R4159 V_p_1.n2 V_p_1.n0 263.933
R4160 V_p_1.n5 V_p_1.n4 206.333
R4161 V_p_1.n2 V_p_1.n1 206.333
R4162 V_p_1.n7 V_p_1.n6 206.333
R4163 V_p_1.n6 V_p_1.t9 134.474
R4164 V_p_1.n6 V_p_1.n2 57.6005
R4165 V_p_1.n6 V_p_1.n5 57.6005
R4166 V_p_1.n3 V_p_1.t10 48.0005
R4167 V_p_1.n3 V_p_1.t5 48.0005
R4168 V_p_1.n4 V_p_1.t7 48.0005
R4169 V_p_1.n4 V_p_1.t1 48.0005
R4170 V_p_1.n0 V_p_1.t3 48.0005
R4171 V_p_1.n0 V_p_1.t6 48.0005
R4172 V_p_1.n1 V_p_1.t4 48.0005
R4173 V_p_1.n1 V_p_1.t2 48.0005
R4174 V_p_1.n7 V_p_1.t0 48.0005
R4175 V_p_1.t8 V_p_1.n7 48.0005
R4176 ERR_AMP_REF.n0 ERR_AMP_REF.t8 688.859
R4177 ERR_AMP_REF.n2 ERR_AMP_REF.n1 514.134
R4178 ERR_AMP_REF.n4 ERR_AMP_REF.n3 214.056
R4179 ERR_AMP_REF.n0 ERR_AMP_REF.t11 174.726
R4180 ERR_AMP_REF.n1 ERR_AMP_REF.t7 174.726
R4181 ERR_AMP_REF.n2 ERR_AMP_REF.t9 174.726
R4182 ERR_AMP_REF.n3 ERR_AMP_REF.t10 174.726
R4183 ERR_AMP_REF.n7 ERR_AMP_REF.n5 173.149
R4184 ERR_AMP_REF.n9 ERR_AMP_REF.n8 168.774
R4185 ERR_AMP_REF.n7 ERR_AMP_REF.n6 168.774
R4186 ERR_AMP_REF.n1 ERR_AMP_REF.n0 128.534
R4187 ERR_AMP_REF.n3 ERR_AMP_REF.n2 128.534
R4188 ERR_AMP_REF.n4 ERR_AMP_REF.t1 125.736
R4189 ERR_AMP_REF.n8 ERR_AMP_REF.t4 13.1338
R4190 ERR_AMP_REF.n8 ERR_AMP_REF.t6 13.1338
R4191 ERR_AMP_REF.n6 ERR_AMP_REF.t0 13.1338
R4192 ERR_AMP_REF.n6 ERR_AMP_REF.t2 13.1338
R4193 ERR_AMP_REF.n5 ERR_AMP_REF.t3 13.1338
R4194 ERR_AMP_REF.n5 ERR_AMP_REF.t5 13.1338
R4195 ERR_AMP_REF.n10 ERR_AMP_REF.n9 10.0317
R4196 ERR_AMP_REF ERR_AMP_REF.n10 8.09425
R4197 ERR_AMP_REF.n9 ERR_AMP_REF.n7 4.3755
R4198 ERR_AMP_REF.n10 ERR_AMP_REF.n4 3.03175
R4199 V_p_2.n5 V_p_2.n3 263.933
R4200 V_p_2.n2 V_p_2.n0 263.933
R4201 V_p_2.n5 V_p_2.n4 206.333
R4202 V_p_2.n2 V_p_2.n1 206.333
R4203 V_p_2.n7 V_p_2.n6 206.333
R4204 V_p_2 V_p_2.t10 120.677
R4205 V_p_2.n7 V_p_2.n2 57.6005
R4206 V_p_2.n7 V_p_2.n5 57.6005
R4207 V_p_2.n3 V_p_2.t8 48.0005
R4208 V_p_2.n3 V_p_2.t3 48.0005
R4209 V_p_2.n4 V_p_2.t4 48.0005
R4210 V_p_2.n4 V_p_2.t7 48.0005
R4211 V_p_2.n0 V_p_2.t9 48.0005
R4212 V_p_2.n0 V_p_2.t5 48.0005
R4213 V_p_2.n1 V_p_2.t2 48.0005
R4214 V_p_2.n1 V_p_2.t1 48.0005
R4215 V_p_2.n6 V_p_2.t0 48.0005
R4216 V_p_2.n6 V_p_2.t6 48.0005
R4217 V_p_2 V_p_2.n7 13.7338
R4218 START_UP_NFET1.t1 START_UP_NFET1.t0 183.816
R4219 V_CMFB_S1.n2 V_CMFB_S1.n0 344.837
R4220 V_CMFB_S1.n2 V_CMFB_S1.n1 344.274
R4221 V_CMFB_S1.n4 V_CMFB_S1.n3 292.5
R4222 V_CMFB_S1.n4 V_CMFB_S1.n2 52.3363
R4223 V_CMFB_S1 V_CMFB_S1.n4 52.1563
R4224 V_CMFB_S1.n3 V_CMFB_S1.t5 39.4005
R4225 V_CMFB_S1.n3 V_CMFB_S1.t1 39.4005
R4226 V_CMFB_S1.n1 V_CMFB_S1.t3 39.4005
R4227 V_CMFB_S1.n1 V_CMFB_S1.t2 39.4005
R4228 V_CMFB_S1.n0 V_CMFB_S1.t0 39.4005
R4229 V_CMFB_S1.n0 V_CMFB_S1.t4 39.4005
R4230 START_UP.n1 START_UP.t7 238.322
R4231 START_UP.n1 START_UP.t6 238.322
R4232 START_UP.n5 START_UP.n4 175.118
R4233 START_UP.n4 START_UP.n3 168.493
R4234 START_UP.n2 START_UP.n1 166.925
R4235 START_UP.n0 START_UP.t5 116.501
R4236 START_UP.n0 START_UP.t4 82.7833
R4237 START_UP.n2 START_UP.n0 49.3505
R4238 START_UP.n3 START_UP.t2 13.1338
R4239 START_UP.n3 START_UP.t3 13.1338
R4240 START_UP.t0 START_UP.n5 13.1338
R4241 START_UP.n5 START_UP.t1 13.1338
R4242 START_UP.n4 START_UP.n2 4.21925
R4243 Vin-.n7 Vin-.t11 688.859
R4244 Vin-.n9 Vin-.n8 514.134
R4245 Vin-.n6 Vin-.n5 356.95
R4246 Vin-.n11 Vin-.n10 213.4
R4247 Vin-.n7 Vin-.t8 174.726
R4248 Vin-.n8 Vin-.t9 174.726
R4249 Vin-.n9 Vin-.t12 174.726
R4250 Vin-.n10 Vin-.t10 174.726
R4251 Vin-.n4 Vin-.n2 172.585
R4252 Vin-.n4 Vin-.n3 168.21
R4253 Vin-.n8 Vin-.n7 128.534
R4254 Vin-.n10 Vin-.n9 128.534
R4255 Vin-.n12 Vin-.t0 119.099
R4256 Vin-.n1 Vin-.n0 83.5719
R4257 Vin-.n17 Vin-.n1 73.682
R4258 Vin-.n5 Vin-.t4 39.4005
R4259 Vin-.n5 Vin-.t5 39.4005
R4260 Vin-.n14 Vin-.t7 36.6632
R4261 Vin-.n13 Vin-.n12 28.813
R4262 Vin-.t7 Vin-.n1 25.7843
R4263 Vin-.n12 Vin-.n11 16.188
R4264 Vin-.n3 Vin-.t6 13.1338
R4265 Vin-.n3 Vin-.t2 13.1338
R4266 Vin-.n2 Vin-.t3 13.1338
R4267 Vin-.n2 Vin-.t1 13.1338
R4268 Vin-.n11 Vin-.n6 11.2193
R4269 Vin-.n6 Vin-.n4 3.8755
R4270 Vin-.n15 Vin-.n14 1.80777
R4271 Vin-.n16 Vin-.n15 1.5505
R4272 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter Vin-.n17 1.07742
R4273 Vin-.n14 Vin-.n13 1.04793
R4274 Vin-.n17 Vin-.n16 0.763532
R4275 Vin-.n15 Vin-.n0 0.590702
R4276 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter Vin-.n0 0.498483
R4277 Vin-.n16 Vin-.n13 0.0106786
R4278 V_TOP.n0 V_TOP.t14 369.534
R4279 V_TOP.n22 V_TOP.n20 345.389
R4280 V_TOP.n19 V_TOP.n18 344.7
R4281 V_TOP.n22 V_TOP.n21 344.7
R4282 V_TOP.n27 V_TOP.n26 344.7
R4283 V_TOP.n29 V_TOP.n28 344.7
R4284 V_TOP.n24 V_TOP.n23 340.2
R4285 V_TOP.n1 V_TOP.n0 224.934
R4286 V_TOP.n2 V_TOP.n1 224.934
R4287 V_TOP.n3 V_TOP.n2 224.934
R4288 V_TOP.n4 V_TOP.n3 224.934
R4289 V_TOP.n5 V_TOP.n4 224.934
R4290 V_TOP.n39 V_TOP.n38 224.934
R4291 V_TOP.n38 V_TOP.n37 224.934
R4292 V_TOP.n37 V_TOP.n36 224.934
R4293 V_TOP.n36 V_TOP.n35 224.934
R4294 V_TOP.n35 V_TOP.n34 224.934
R4295 V_TOP.n34 V_TOP.n33 224.934
R4296 V_TOP.n33 V_TOP.n32 224.934
R4297 V_TOP V_TOP.t27 214.222
R4298 V_TOP.n31 V_TOP.n30 163.175
R4299 V_TOP.n0 V_TOP.t41 144.601
R4300 V_TOP.n1 V_TOP.t37 144.601
R4301 V_TOP.n2 V_TOP.t30 144.601
R4302 V_TOP.n3 V_TOP.t25 144.601
R4303 V_TOP.n4 V_TOP.t15 144.601
R4304 V_TOP.n5 V_TOP.t43 144.601
R4305 V_TOP.n39 V_TOP.t31 144.601
R4306 V_TOP.n38 V_TOP.t38 144.601
R4307 V_TOP.n37 V_TOP.t42 144.601
R4308 V_TOP.n36 V_TOP.t45 144.601
R4309 V_TOP.n35 V_TOP.t19 144.601
R4310 V_TOP.n34 V_TOP.t28 144.601
R4311 V_TOP.n33 V_TOP.t34 144.601
R4312 V_TOP.n32 V_TOP.t40 144.601
R4313 V_TOP.n30 V_TOP.t7 111.397
R4314 V_TOP.n17 V_TOP.t0 108.424
R4315 V_TOP.n31 V_TOP.n5 69.6227
R4316 V_TOP V_TOP.n39 69.6227
R4317 V_TOP.n32 V_TOP.n31 69.6227
R4318 V_TOP.n18 V_TOP.t13 39.4005
R4319 V_TOP.n18 V_TOP.t5 39.4005
R4320 V_TOP.n23 V_TOP.t10 39.4005
R4321 V_TOP.n23 V_TOP.t12 39.4005
R4322 V_TOP.n21 V_TOP.t4 39.4005
R4323 V_TOP.n21 V_TOP.t2 39.4005
R4324 V_TOP.n20 V_TOP.t1 39.4005
R4325 V_TOP.n20 V_TOP.t3 39.4005
R4326 V_TOP.n26 V_TOP.t8 39.4005
R4327 V_TOP.n26 V_TOP.t11 39.4005
R4328 V_TOP.n28 V_TOP.t6 39.4005
R4329 V_TOP.n28 V_TOP.t9 39.4005
R4330 V_TOP.n17 V_TOP.n16 37.1479
R4331 V_TOP.n19 V_TOP.n17 27.8371
R4332 V_TOP.n24 V_TOP.n22 8.313
R4333 V_TOP.n30 V_TOP.n29 5.188
R4334 V_TOP.n7 V_TOP.t49 4.8295
R4335 V_TOP.n6 V_TOP.t24 4.8295
R4336 V_TOP.n9 V_TOP.t36 4.8295
R4337 V_TOP.n8 V_TOP.t18 4.8295
R4338 V_TOP.n11 V_TOP.t22 4.8295
R4339 V_TOP.n10 V_TOP.t46 4.8295
R4340 V_TOP.n13 V_TOP.t33 4.8295
R4341 V_TOP.n12 V_TOP.t16 4.8295
R4342 V_TOP.n14 V_TOP.t44 4.8295
R4343 V_TOP.n7 V_TOP.t47 4.5005
R4344 V_TOP.n6 V_TOP.t26 4.5005
R4345 V_TOP.n9 V_TOP.t35 4.5005
R4346 V_TOP.n8 V_TOP.t20 4.5005
R4347 V_TOP.n11 V_TOP.t21 4.5005
R4348 V_TOP.n10 V_TOP.t48 4.5005
R4349 V_TOP.n13 V_TOP.t32 4.5005
R4350 V_TOP.n12 V_TOP.t17 4.5005
R4351 V_TOP.n14 V_TOP.t29 4.5005
R4352 V_TOP.n15 V_TOP.t39 4.5005
R4353 V_TOP.n16 V_TOP.t23 4.5005
R4354 V_TOP.n25 V_TOP.n24 4.5005
R4355 V_TOP.n29 V_TOP.n27 2.1255
R4356 V_TOP.n27 V_TOP.n25 2.1255
R4357 V_TOP.n25 V_TOP.n19 2.1255
R4358 V_TOP.n7 V_TOP.n6 0.3295
R4359 V_TOP.n9 V_TOP.n8 0.3295
R4360 V_TOP.n11 V_TOP.n10 0.3295
R4361 V_TOP.n13 V_TOP.n12 0.3295
R4362 V_TOP.n15 V_TOP.n14 0.3295
R4363 V_TOP.n16 V_TOP.n15 0.3295
R4364 V_TOP.n9 V_TOP.n7 0.2825
R4365 V_TOP.n11 V_TOP.n9 0.2825
R4366 V_TOP.n13 V_TOP.n11 0.2825
R4367 V_TOP.n14 V_TOP.n13 0.2825
R4368 V_CMFB_S3.n2 V_CMFB_S3.n0 345.264
R4369 V_CMFB_S3.n2 V_CMFB_S3.n1 344.7
R4370 V_CMFB_S3.n4 V_CMFB_S3.n3 292.5
R4371 V_CMFB_S3.n4 V_CMFB_S3.n2 52.763
R4372 V_CMFB_S3 V_CMFB_S3.n4 51.7297
R4373 V_CMFB_S3.n3 V_CMFB_S3.t0 39.4005
R4374 V_CMFB_S3.n3 V_CMFB_S3.t5 39.4005
R4375 V_CMFB_S3.n1 V_CMFB_S3.t1 39.4005
R4376 V_CMFB_S3.n1 V_CMFB_S3.t2 39.4005
R4377 V_CMFB_S3.n0 V_CMFB_S3.t4 39.4005
R4378 V_CMFB_S3.n0 V_CMFB_S3.t3 39.4005
R4379 VB3_CUR_BIAS.n2 VB3_CUR_BIAS.n1 145.262
R4380 VB3_CUR_BIAS.n2 VB3_CUR_BIAS.n0 145.262
R4381 VB3_CUR_BIAS.n4 VB3_CUR_BIAS.n3 140.201
R4382 VB3_CUR_BIAS VB3_CUR_BIAS.n4 41.063
R4383 VB3_CUR_BIAS.n3 VB3_CUR_BIAS.t4 24.0005
R4384 VB3_CUR_BIAS.n3 VB3_CUR_BIAS.t2 24.0005
R4385 VB3_CUR_BIAS.n1 VB3_CUR_BIAS.t0 24.0005
R4386 VB3_CUR_BIAS.n1 VB3_CUR_BIAS.t3 24.0005
R4387 VB3_CUR_BIAS.n0 VB3_CUR_BIAS.t5 24.0005
R4388 VB3_CUR_BIAS.n0 VB3_CUR_BIAS.t1 24.0005
R4389 VB3_CUR_BIAS.n4 VB3_CUR_BIAS.n2 4.5005
R4390 V_mir1.n9 V_mir1.n5 330.901
R4391 V_mir1.n4 V_mir1.n0 330.901
R4392 V_mir1.n20 V_mir1.n19 330.901
R4393 V_mir1.n16 V_mir1.t20 310.488
R4394 V_mir1.n6 V_mir1.t19 310.488
R4395 V_mir1.n1 V_mir1.t22 310.488
R4396 V_mir1.n13 V_mir1.t13 278.312
R4397 V_mir1.n13 V_mir1.n12 228.939
R4398 V_mir1.n14 V_mir1.n11 224.439
R4399 V_mir1.n18 V_mir1.t0 184.097
R4400 V_mir1.n8 V_mir1.t4 184.097
R4401 V_mir1.n3 V_mir1.t8 184.097
R4402 V_mir1.n17 V_mir1.n16 167.094
R4403 V_mir1.n7 V_mir1.n6 167.094
R4404 V_mir1.n2 V_mir1.n1 167.094
R4405 V_mir1.n9 V_mir1.n8 152
R4406 V_mir1.n4 V_mir1.n3 152
R4407 V_mir1.n19 V_mir1.n18 152
R4408 V_mir1.n16 V_mir1.t18 120.501
R4409 V_mir1.n17 V_mir1.t10 120.501
R4410 V_mir1.n6 V_mir1.t17 120.501
R4411 V_mir1.n7 V_mir1.t2 120.501
R4412 V_mir1.n1 V_mir1.t21 120.501
R4413 V_mir1.n2 V_mir1.t6 120.501
R4414 V_mir1.n12 V_mir1.t16 48.0005
R4415 V_mir1.n12 V_mir1.t15 48.0005
R4416 V_mir1.n11 V_mir1.t12 48.0005
R4417 V_mir1.n11 V_mir1.t14 48.0005
R4418 V_mir1.n18 V_mir1.n17 40.7027
R4419 V_mir1.n8 V_mir1.n7 40.7027
R4420 V_mir1.n3 V_mir1.n2 40.7027
R4421 V_mir1.n5 V_mir1.t3 39.4005
R4422 V_mir1.n5 V_mir1.t5 39.4005
R4423 V_mir1.n0 V_mir1.t7 39.4005
R4424 V_mir1.n0 V_mir1.t9 39.4005
R4425 V_mir1.t11 V_mir1.n20 39.4005
R4426 V_mir1.n20 V_mir1.t1 39.4005
R4427 V_mir1.n10 V_mir1.n9 15.8005
R4428 V_mir1.n10 V_mir1.n4 15.8005
R4429 V_mir1.n19 V_mir1.n15 9.3005
R4430 V_mir1.n14 V_mir1.n13 5.8755
R4431 V_mir1.n15 V_mir1.n10 4.5005
R4432 V_mir1.n15 V_mir1.n14 0.78175
R4433 V_CUR_REF_REG.n4 V_CUR_REF_REG.n3 526.183
R4434 V_CUR_REF_REG.n2 V_CUR_REF_REG.n1 514.134
R4435 V_CUR_REF_REG.n5 V_CUR_REF_REG.n0 378.053
R4436 V_CUR_REF_REG.n1 V_CUR_REF_REG.t4 303.259
R4437 V_CUR_REF_REG.n5 V_CUR_REF_REG.n4 210.169
R4438 V_CUR_REF_REG.n1 V_CUR_REF_REG.t5 174.726
R4439 V_CUR_REF_REG.n2 V_CUR_REF_REG.t7 174.726
R4440 V_CUR_REF_REG.n3 V_CUR_REF_REG.t3 174.726
R4441 V_CUR_REF_REG.t0 V_CUR_REF_REG.n5 153.474
R4442 V_CUR_REF_REG.n3 V_CUR_REF_REG.n2 128.534
R4443 V_CUR_REF_REG.n4 V_CUR_REF_REG.t6 96.4005
R4444 V_CUR_REF_REG.n0 V_CUR_REF_REG.t2 39.4005
R4445 V_CUR_REF_REG.n0 V_CUR_REF_REG.t1 39.4005
R4446 a_32320_n7778.t0 a_32320_n7778.t1 178.133
R4447 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t0 195.608
R4448 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 83.5719
R4449 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 83.5719
R4450 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 83.5719
R4451 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 83.5719
R4452 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 83.5719
R4453 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 83.5719
R4454 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 83.5719
R4455 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 83.5719
R4456 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 83.5719
R4457 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 83.5719
R4458 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 83.5719
R4459 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 83.5719
R4460 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 83.5719
R4461 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 83.5719
R4462 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 83.5719
R4463 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 83.5719
R4464 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 83.5719
R4465 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 83.5719
R4466 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 83.5719
R4467 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 83.5719
R4468 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 73.682
R4469 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 73.682
R4470 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 73.3165
R4471 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 73.3165
R4472 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 73.3165
R4473 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 73.3165
R4474 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 73.3165
R4475 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 73.3165
R4476 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 73.19
R4477 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 73.19
R4478 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 73.19
R4479 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 73.19
R4480 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 73.19
R4481 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 73.19
R4482 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 36.6632
R4483 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 36.6632
R4484 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n53 26.074
R4485 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n89 26.074
R4486 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n74 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 26.074
R4487 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n104 26.074
R4488 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n9 26.074
R4489 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n4 26.074
R4490 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n57 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 25.7843
R4491 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n91 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 25.7843
R4492 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n28 25.7843
R4493 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t7 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n33 25.7843
R4494 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n108 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 25.7843
R4495 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n13 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 25.7843
R4496 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n125 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 25.7843
R4497 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t6 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n49 25.7843
R4498 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4499 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4500 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4501 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 9.3005
R4502 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4503 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4504 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4505 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 9.3005
R4506 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4507 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4508 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4509 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 9.3005
R4510 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4511 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4512 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4513 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 9.3005
R4514 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4515 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4516 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4517 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R4518 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 9.3005
R4519 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 9.3005
R4520 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 9.3005
R4521 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 9.3005
R4522 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 9.3005
R4523 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 9.3005
R4524 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4525 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4526 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4527 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 9.3005
R4528 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R4529 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4530 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4531 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4532 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 9.3005
R4533 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 9.3005
R4534 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4535 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4536 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4537 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 9.3005
R4538 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4539 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4540 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4541 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 9.3005
R4542 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4543 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4544 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4545 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 9.3005
R4546 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 9.3005
R4547 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 9.3005
R4548 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 9.3005
R4549 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 9.3005
R4550 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 9.3005
R4551 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 9.3005
R4552 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 4.64654
R4553 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 4.64654
R4554 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 4.64654
R4555 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 4.64654
R4556 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 4.64654
R4557 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 4.64654
R4558 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 4.64654
R4559 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 4.64654
R4560 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 4.64654
R4561 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 2.36206
R4562 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 2.36206
R4563 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 2.36206
R4564 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 2.36206
R4565 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 2.19742
R4566 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 2.19742
R4567 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 2.19742
R4568 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 2.19742
R4569 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.80777
R4570 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 1.80777
R4571 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 1.5505
R4572 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 1.5505
R4573 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 1.5505
R4574 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 1.5505
R4575 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 1.5505
R4576 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 1.5505
R4577 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 1.5505
R4578 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 1.5505
R4579 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 1.5505
R4580 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 1.5505
R4581 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 1.5505
R4582 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 1.5505
R4583 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 1.5505
R4584 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 1.5505
R4585 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 1.5505
R4586 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 1.5505
R4587 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 1.5505
R4588 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 1.5505
R4589 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 1.19225
R4590 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n26 1.19225
R4591 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n72 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 1.19225
R4592 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 1.19225
R4593 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n120 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 1.19225
R4594 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n133 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 1.19225
R4595 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 1.07742
R4596 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 1.07742
R4597 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 1.07024
R4598 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 1.07024
R4599 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 1.07024
R4600 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 1.07024
R4601 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 1.07024
R4602 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 1.07024
R4603 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n50 1.04793
R4604 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n34 1.04793
R4605 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 1.0237
R4606 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n82 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 1.0237
R4607 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n69 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 1.0237
R4608 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 1.0237
R4609 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n124 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 1.0237
R4610 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n1 1.0237
R4611 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n36 0.959578
R4612 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n86 0.959578
R4613 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n31 0.959578
R4614 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n17 0.959578
R4615 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n119 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 0.959578
R4616 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n132 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 0.959578
R4617 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n52 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 0.885803
R4618 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n88 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 0.885803
R4619 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n75 0.885803
R4620 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n103 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.885803
R4621 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n118 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 0.885803
R4622 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n131 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 0.885803
R4623 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n59 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n58 0.812055
R4624 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n110 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n109 0.812055
R4625 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n54 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n39 0.77514
R4626 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n87 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n25 0.77514
R4627 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n76 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n29 0.77514
R4628 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n105 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n21 0.77514
R4629 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n117 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n10 0.77514
R4630 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n130 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n5 0.77514
R4631 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n11 0.763532
R4632 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n24 0.763532
R4633 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n38 0.756696
R4634 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n81 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R4635 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n68 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R4636 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n20 0.756696
R4637 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n123 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.756696
R4638 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n137 0.756696
R4639 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n62 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n40 0.647417
R4640 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n113 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n22 0.647417
R4641 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n37 0.590702
R4642 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n93 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 0.590702
R4643 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n79 0.590702
R4644 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n66 0.590702
R4645 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n18 0.590702
R4646 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n15 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 0.590702
R4647 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n127 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 0.590702
R4648 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n48 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.590702
R4649 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n56 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4650 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n92 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4651 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n80 0.498483
R4652 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n67 0.498483
R4653 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n107 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4654 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n14 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4655 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n126 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.498483
R4656 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n0 0.498483
R4657 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t8 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n55 0.290206
R4658 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t4 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n90 0.290206
R4659 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n73 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t2 0.290206
R4660 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t5 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n106 0.290206
R4661 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t3 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n12 0.290206
R4662 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.t1 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n7 0.290206
R4663 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 0.154071
R4664 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 0.154071
R4665 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 0.154071
R4666 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 0.154071
R4667 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 0.137464
R4668 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 0.137464
R4669 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 0.134964
R4670 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 0.134964
R4671 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0183571
R4672 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n136 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n135 0.0183571
R4673 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n134 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R4674 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n3 0.0183571
R4675 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n129 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 0.0183571
R4676 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n128 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R4677 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n122 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n6 0.0183571
R4678 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n121 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 0.0183571
R4679 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n8 0.0183571
R4680 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.0183571
R4681 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n70 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n32 0.0183571
R4682 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n71 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.0183571
R4683 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n30 0.0183571
R4684 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n77 0.0183571
R4685 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n78 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 0.0183571
R4686 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n83 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n27 0.0183571
R4687 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n84 0.0183571
R4688 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n85 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.0183571
R4689 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n51 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n2 0.0106786
R4690 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n16 0.0106786
R4691 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n65 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n64 0.0106786
R4692 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n94 0.0106786
R4693 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 0.0106786
R4694 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n114 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R4695 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 0.00992001
R4696 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 0.00992001
R4697 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 0.00992001
R4698 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n96 0.00992001
R4699 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n19 0.00992001
R4700 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n99 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n98 0.00992001
R4701 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n102 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n100 0.00992001
R4702 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n101 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n97 0.00992001
R4703 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n112 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n111 0.00992001
R4704 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n61 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 0.00992001
R4705 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 0.00992001
R4706 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 0.00992001
R4707 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n63 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.00992001
R4708 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n60 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.00992001
R4709 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n43 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n42 0.00992001
R4710 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n46 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n41 0.00992001
R4711 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n47 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n35 0.00992001
R4712 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n116 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n115 0.00817857
R4713 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n95 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n23 0.00817857
R4714 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n45 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter.n44 0.00817857
R4715 a_38040_n7928.t0 a_38040_n7928.t1 178.133
R4716 ERR_AMP_CUR_BIAS ERR_AMP_CUR_BIAS.n0 180.794
R4717 ERR_AMP_CUR_BIAS.n0 ERR_AMP_CUR_BIAS.t1 24.0005
R4718 ERR_AMP_CUR_BIAS.n0 ERR_AMP_CUR_BIAS.t0 24.0005
R4719 a_32970_n7928.t0 a_32970_n7928.t1 178.133
R4720 a_32440_n6570.t0 a_32440_n6570.t1 178.133
R4721 a_33090_n6320.t0 a_33090_n6320.t1 178.133
R4722 a_37920_n6320.t0 a_37920_n6320.t1 178.133
C0 VB1_CUR_BIAS PFET_GATE_10uA 0.151852f
C1 V_TOP 1st_Vout_2 0.073737f
C2 VDDA VB2_CUR_BIAS 0.011895f
C3 cap_res2 1st_Vout_2 7.78879f
C4 V_CMFB_S1 TAIL_CUR_MIR_BIAS 0.021516f
C5 VB2_CUR_BIAS V_CMFB_S2 1.66154f
C6 PFET_GATE_10uA ERR_AMP_CUR_BIAS 0.011616f
C7 1st_Vout_2 ERR_AMP_REF 0.670874f
C8 V_p_2 1st_Vout_2 0.311653f
C9 1st_Vout_2 VDDA 1.53362f
C10 VB3_CUR_BIAS PFET_GATE_10uA 1.13474f
C11 V_CMFB_S3 TAIL_CUR_MIR_BIAS 0.015021f
C12 VB2_CUR_BIAS ERR_AMP_CUR_BIAS 1.86293f
C13 cap_res2 V_TOP 0.01893f
C14 ERR_AMP_REF V_CMFB_S4 0.03827f
C15 VDDA V_CMFB_S1 0.785042f
C16 VB2_CUR_BIAS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.011598f
C17 V_CMFB_S4 VDDA 0.232993f
C18 V_TOP ERR_AMP_REF 0.583702f
C19 VB3_CUR_BIAS VB2_CUR_BIAS 0.383231f
C20 V_TOP VDDA 13.526401f
C21 VDDA TAIL_CUR_MIR_BIAS 0.831217f
C22 V_CMFB_S3 VDDA 0.783868f
C23 cap_res2 VDDA 1.06733f
C24 V_CMFB_S3 VB1_CUR_BIAS 0.017903f
C25 V_TOP V_CMFB_S2 0.503779f
C26 V_p_2 ERR_AMP_REF 0.124262f
C27 1st_Vout_2 VB3_CUR_BIAS 0.042806f
C28 ERR_AMP_REF VDDA 1.53646f
C29 V_p_2 VDDA 0.566952f
C30 ERR_AMP_REF VB1_CUR_BIAS 0.200016f
C31 V_TOP ERR_AMP_CUR_BIAS 0.08195f
C32 VB3_CUR_BIAS V_CMFB_S4 0.818388f
C33 VB1_CUR_BIAS VDDA 0.566908f
C34 V_TOP sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.055802f
C35 VDDA V_CMFB_S2 0.03011f
C36 1st_Vout_2 PFET_GATE_10uA 1.5028f
C37 VDDA ERR_AMP_CUR_BIAS 0.056576f
C38 ERR_AMP_REF VB3_CUR_BIAS 0.414647f
C39 V_CMFB_S1 PFET_GATE_10uA 0.216843f
C40 VDDA sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter 0.046803f
C41 V_CMFB_S4 PFET_GATE_10uA 0.137571f
C42 VB3_CUR_BIAS VDDA 0.183515f
C43 V_CMFB_S2 ERR_AMP_CUR_BIAS 0.063017f
C44 V_TOP PFET_GATE_10uA 0.212258f
C45 TAIL_CUR_MIR_BIAS PFET_GATE_10uA 0.237552f
C46 V_CMFB_S3 PFET_GATE_10uA 0.356974f
C47 V_CMFB_S4 VB2_CUR_BIAS 0.559002f
C48 V_TOP VB2_CUR_BIAS 0.936691f
C49 ERR_AMP_REF PFET_GATE_10uA 1.67029f
C50 VB3_CUR_BIAS ERR_AMP_CUR_BIAS 0.096717f
C51 V_p_2 PFET_GATE_10uA 0.010026f
C52 VDDA PFET_GATE_10uA 8.289901f
C53 1st_Vout_2 V_CMFB_S4 1.40961f
C54 V_CMFB_S4 GNDA 3.39236f
C55 VB3_CUR_BIAS GNDA 2.31377f
C56 ERR_AMP_CUR_BIAS GNDA 4.2973f
C57 V_CMFB_S2 GNDA 2.64392f
C58 VB2_CUR_BIAS GNDA 2.86051f
C59 VB1_CUR_BIAS GNDA 0.664246f
C60 ERR_AMP_REF GNDA 3.916142f
C61 V_CMFB_S3 GNDA 0.551428f
C62 TAIL_CUR_MIR_BIAS GNDA 0.40902f
C63 V_CMFB_S1 GNDA 0.588375f
C64 VDDA GNDA 74.79788f
C65 cap_res2 GNDA 6.69715f
C66 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_25.Emitter GNDA 17.900902f
C67 V_p_2 GNDA 0.764548f
C68 1st_Vout_2 GNDA 8.084408f
C69 V_TOP GNDA 9.886665f
C70 PFET_GATE_10uA GNDA 6.606697f
C71 ERR_AMP_CUR_BIAS.t1 GNDA 0.029966f
C72 ERR_AMP_CUR_BIAS.t0 GNDA 0.029966f
C73 ERR_AMP_CUR_BIAS.n0 GNDA 0.446705f
C74 V_mir1.t1 GNDA 0.019293f
C75 V_mir1.t7 GNDA 0.019293f
C76 V_mir1.t9 GNDA 0.019293f
C77 V_mir1.n0 GNDA 0.044322f
C78 V_mir1.t6 GNDA 0.023151f
C79 V_mir1.t21 GNDA 0.023151f
C80 V_mir1.t22 GNDA 0.037369f
C81 V_mir1.n1 GNDA 0.041731f
C82 V_mir1.n2 GNDA 0.028507f
C83 V_mir1.t8 GNDA 0.02939f
C84 V_mir1.n3 GNDA 0.044354f
C85 V_mir1.n4 GNDA 0.109787f
C86 V_mir1.t3 GNDA 0.019293f
C87 V_mir1.t5 GNDA 0.019293f
C88 V_mir1.n5 GNDA 0.044322f
C89 V_mir1.t2 GNDA 0.023151f
C90 V_mir1.t17 GNDA 0.023151f
C91 V_mir1.t19 GNDA 0.037369f
C92 V_mir1.n6 GNDA 0.041731f
C93 V_mir1.n7 GNDA 0.028507f
C94 V_mir1.t4 GNDA 0.02939f
C95 V_mir1.n8 GNDA 0.044354f
C96 V_mir1.n9 GNDA 0.110886f
C97 V_mir1.n10 GNDA 0.381359f
C98 V_mir1.n11 GNDA 0.025223f
C99 V_mir1.t13 GNDA 0.041163f
C100 V_mir1.n12 GNDA 0.027381f
C101 V_mir1.n13 GNDA 0.451535f
C102 V_mir1.n14 GNDA 0.146338f
C103 V_mir1.n15 GNDA 0.051125f
C104 V_mir1.t10 GNDA 0.023151f
C105 V_mir1.t18 GNDA 0.023151f
C106 V_mir1.t20 GNDA 0.037369f
C107 V_mir1.n16 GNDA 0.041731f
C108 V_mir1.n17 GNDA 0.028507f
C109 V_mir1.t0 GNDA 0.02939f
C110 V_mir1.n18 GNDA 0.044354f
C111 V_mir1.n19 GNDA 0.084938f
C112 V_mir1.n20 GNDA 0.044322f
C113 V_mir1.t11 GNDA 0.019293f
C114 V_TOP.t27 GNDA 0.112091f
C115 V_TOP.t31 GNDA 0.097271f
C116 V_TOP.t38 GNDA 0.097271f
C117 V_TOP.t42 GNDA 0.097271f
C118 V_TOP.t45 GNDA 0.097271f
C119 V_TOP.t19 GNDA 0.097271f
C120 V_TOP.t28 GNDA 0.097271f
C121 V_TOP.t34 GNDA 0.097271f
C122 V_TOP.t40 GNDA 0.097271f
C123 V_TOP.t43 GNDA 0.097271f
C124 V_TOP.t15 GNDA 0.097271f
C125 V_TOP.t25 GNDA 0.097271f
C126 V_TOP.t30 GNDA 0.097271f
C127 V_TOP.t37 GNDA 0.097271f
C128 V_TOP.t41 GNDA 0.097271f
C129 V_TOP.t14 GNDA 0.127158f
C130 V_TOP.n0 GNDA 0.071091f
C131 V_TOP.n1 GNDA 0.051878f
C132 V_TOP.n2 GNDA 0.051878f
C133 V_TOP.n3 GNDA 0.051878f
C134 V_TOP.n4 GNDA 0.051878f
C135 V_TOP.n5 GNDA 0.048377f
C136 V_TOP.t7 GNDA 0.126138f
C137 V_TOP.t49 GNDA 0.37687f
C138 V_TOP.t47 GNDA 0.370558f
C139 V_TOP.t24 GNDA 0.37687f
C140 V_TOP.t26 GNDA 0.370558f
C141 V_TOP.n6 GNDA 0.248447f
C142 V_TOP.n7 GNDA 0.317927f
C143 V_TOP.t36 GNDA 0.37687f
C144 V_TOP.t35 GNDA 0.370558f
C145 V_TOP.t18 GNDA 0.37687f
C146 V_TOP.t20 GNDA 0.370558f
C147 V_TOP.n8 GNDA 0.248447f
C148 V_TOP.n9 GNDA 0.387406f
C149 V_TOP.t22 GNDA 0.37687f
C150 V_TOP.t21 GNDA 0.370558f
C151 V_TOP.t46 GNDA 0.37687f
C152 V_TOP.t48 GNDA 0.370558f
C153 V_TOP.n10 GNDA 0.248447f
C154 V_TOP.n11 GNDA 0.387406f
C155 V_TOP.t33 GNDA 0.37687f
C156 V_TOP.t32 GNDA 0.370558f
C157 V_TOP.t16 GNDA 0.37687f
C158 V_TOP.t17 GNDA 0.370558f
C159 V_TOP.n12 GNDA 0.248447f
C160 V_TOP.n13 GNDA 0.387406f
C161 V_TOP.t44 GNDA 0.37687f
C162 V_TOP.t29 GNDA 0.370558f
C163 V_TOP.n14 GNDA 0.317927f
C164 V_TOP.t39 GNDA 0.370558f
C165 V_TOP.n15 GNDA 0.162119f
C166 V_TOP.t23 GNDA 0.370558f
C167 V_TOP.n16 GNDA 0.554811f
C168 V_TOP.t0 GNDA 0.104243f
C169 V_TOP.n17 GNDA 0.73814f
C170 V_TOP.n18 GNDA 0.023109f
C171 V_TOP.n19 GNDA 0.422529f
C172 V_TOP.n20 GNDA 0.023262f
C173 V_TOP.n21 GNDA 0.023109f
C174 V_TOP.n22 GNDA 0.213681f
C175 V_TOP.n23 GNDA 0.022398f
C176 V_TOP.n24 GNDA 0.129796f
C177 V_TOP.n25 GNDA 0.074112f
C178 V_TOP.n26 GNDA 0.023109f
C179 V_TOP.n27 GNDA 0.127893f
C180 V_TOP.n28 GNDA 0.023109f
C181 V_TOP.n29 GNDA 0.126677f
C182 V_TOP.n30 GNDA 0.277504f
C183 V_TOP.n31 GNDA 0.019602f
C184 V_TOP.n32 GNDA 0.048377f
C185 V_TOP.n33 GNDA 0.051878f
C186 V_TOP.n34 GNDA 0.051878f
C187 V_TOP.n35 GNDA 0.051878f
C188 V_TOP.n36 GNDA 0.051878f
C189 V_TOP.n37 GNDA 0.051878f
C190 V_TOP.n38 GNDA 0.051878f
C191 V_TOP.n39 GNDA 0.048377f
C192 Vin-.n0 GNDA 0.046896f
C193 Vin-.n1 GNDA 0.320511f
C194 Vin-.t3 GNDA 0.027487f
C195 Vin-.t1 GNDA 0.027487f
C196 Vin-.n2 GNDA 0.099751f
C197 Vin-.t6 GNDA 0.027487f
C198 Vin-.t2 GNDA 0.027487f
C199 Vin-.n3 GNDA 0.09553f
C200 Vin-.n4 GNDA 0.383788f
C201 Vin-.n5 GNDA 0.028037f
C202 Vin-.n6 GNDA 0.371517f
C203 Vin-.t11 GNDA 0.022665f
C204 Vin-.n7 GNDA 0.026583f
C205 Vin-.n8 GNDA 0.021761f
C206 Vin-.n9 GNDA 0.021761f
C207 Vin-.n10 GNDA 0.037011f
C208 Vin-.n11 GNDA 0.505034f
C209 Vin-.t0 GNDA 0.120899f
C210 Vin-.n12 GNDA 0.678321f
C211 Vin-.n13 GNDA 1.35751f
C212 Vin-.t7 GNDA 0.333763f
C213 Vin-.n14 GNDA 0.298273f
C214 Vin-.n15 GNDA 0.124261f
C215 Vin-.n16 GNDA 0.587205f
C216 Vin-.n17 GNDA 0.373496f
C217 sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_23.Emitter GNDA 0.083247f
C218 START_UP.t1 GNDA 0.027731f
C219 START_UP.t4 GNDA 1.11411f
C220 START_UP.t5 GNDA 0.031262f
C221 START_UP.n0 GNDA 0.808511f
C222 START_UP.t6 GNDA 0.010421f
C223 START_UP.t7 GNDA 0.010421f
C224 START_UP.n1 GNDA 0.029418f
C225 START_UP.n2 GNDA 0.512458f
C226 START_UP.t2 GNDA 0.027731f
C227 START_UP.t3 GNDA 0.027731f
C228 START_UP.n3 GNDA 0.096735f
C229 START_UP.n4 GNDA 0.471093f
C230 START_UP.n5 GNDA 0.104651f
C231 START_UP.t0 GNDA 0.027731f
C232 ERR_AMP_REF.t1 GNDA 0.146345f
C233 ERR_AMP_REF.t8 GNDA 0.022576f
C234 ERR_AMP_REF.n0 GNDA 0.026478f
C235 ERR_AMP_REF.n1 GNDA 0.021675f
C236 ERR_AMP_REF.n2 GNDA 0.021675f
C237 ERR_AMP_REF.n3 GNDA 0.037766f
C238 ERR_AMP_REF.n4 GNDA 0.765165f
C239 ERR_AMP_REF.t3 GNDA 0.027379f
C240 ERR_AMP_REF.t5 GNDA 0.027379f
C241 ERR_AMP_REF.n5 GNDA 0.100461f
C242 ERR_AMP_REF.t0 GNDA 0.027379f
C243 ERR_AMP_REF.t2 GNDA 0.027379f
C244 ERR_AMP_REF.n6 GNDA 0.095873f
C245 ERR_AMP_REF.n7 GNDA 0.420606f
C246 ERR_AMP_REF.t4 GNDA 0.027379f
C247 ERR_AMP_REF.t6 GNDA 0.027379f
C248 ERR_AMP_REF.n8 GNDA 0.095873f
C249 ERR_AMP_REF.n9 GNDA 0.302474f
C250 ERR_AMP_REF.n10 GNDA 0.22496f
C251 Vin+.t8 GNDA 0.010641f
C252 Vin+.t9 GNDA 0.025236f
C253 Vin+.t7 GNDA 0.016404f
C254 Vin+.n0 GNDA 0.054125f
C255 Vin+.t6 GNDA 0.016404f
C256 Vin+.n1 GNDA 0.042119f
C257 Vin+.t10 GNDA 0.016404f
C258 Vin+.n2 GNDA 0.042687f
C259 Vin+.n3 GNDA 0.130116f
C260 Vin+.t0 GNDA 0.053203f
C261 Vin+.t2 GNDA 0.053203f
C262 Vin+.n4 GNDA 0.183813f
C263 Vin+.n5 GNDA 1.26385f
C264 Vin+.t3 GNDA 0.053203f
C265 Vin+.t5 GNDA 0.053203f
C266 Vin+.n6 GNDA 0.183813f
C267 Vin+.n7 GNDA 1.0517f
C268 Vin+.t4 GNDA 0.233821f
C269 Vin+.n8 GNDA 1.743f
C270 Vin+.t1 GNDA 0.173052f
C271 cap_res1.t14 GNDA 0.349634f
C272 cap_res1.t1 GNDA 0.350901f
C273 cap_res1.t4 GNDA 0.332137f
C274 cap_res1.t16 GNDA 0.349634f
C275 cap_res1.t17 GNDA 0.350901f
C276 cap_res1.t8 GNDA 0.332137f
C277 cap_res1.t2 GNDA 0.349634f
C278 cap_res1.t3 GNDA 0.350901f
C279 cap_res1.t12 GNDA 0.332137f
C280 cap_res1.t13 GNDA 0.349634f
C281 cap_res1.t15 GNDA 0.350901f
C282 cap_res1.t6 GNDA 0.332137f
C283 cap_res1.t9 GNDA 0.349634f
C284 cap_res1.t11 GNDA 0.350901f
C285 cap_res1.t20 GNDA 0.332137f
C286 cap_res1.n0 GNDA 0.23436f
C287 cap_res1.t19 GNDA 0.186633f
C288 cap_res1.n1 GNDA 0.254286f
C289 cap_res1.t5 GNDA 0.186633f
C290 cap_res1.n2 GNDA 0.254286f
C291 cap_res1.t10 GNDA 0.186633f
C292 cap_res1.n3 GNDA 0.254286f
C293 cap_res1.t7 GNDA 0.186633f
C294 cap_res1.n4 GNDA 0.254286f
C295 cap_res1.t18 GNDA 0.355331f
C296 cap_res1.t0 GNDA 0.083274f
C297 1st_Vout_1.n0 GNDA 0.902606f
C298 1st_Vout_1.n1 GNDA 0.290245f
C299 1st_Vout_1.n2 GNDA 1.74831f
C300 1st_Vout_1.n3 GNDA 0.12751f
C301 1st_Vout_1.n4 GNDA 1.79885f
C302 1st_Vout_1.n5 GNDA 0.012728f
C303 1st_Vout_1.t5 GNDA 0.018559f
C304 1st_Vout_1.n6 GNDA 0.192525f
C305 1st_Vout_1.n7 GNDA 0.011517f
C306 1st_Vout_1.t32 GNDA 0.021148f
C307 1st_Vout_1.n8 GNDA 0.022249f
C308 1st_Vout_1.t36 GNDA 0.013423f
C309 1st_Vout_1.t28 GNDA 0.013423f
C310 1st_Vout_1.n9 GNDA 0.029862f
C311 1st_Vout_1.t17 GNDA 0.35246f
C312 1st_Vout_1.t23 GNDA 0.358463f
C313 1st_Vout_1.t21 GNDA 0.35246f
C314 1st_Vout_1.t12 GNDA 0.35246f
C315 1st_Vout_1.t11 GNDA 0.358463f
C316 1st_Vout_1.t18 GNDA 0.358463f
C317 1st_Vout_1.t16 GNDA 0.35246f
C318 1st_Vout_1.t29 GNDA 0.35246f
C319 1st_Vout_1.t27 GNDA 0.358463f
C320 1st_Vout_1.t34 GNDA 0.358463f
C321 1st_Vout_1.t33 GNDA 0.35246f
C322 1st_Vout_1.t22 GNDA 0.35246f
C323 1st_Vout_1.t20 GNDA 0.358463f
C324 1st_Vout_1.t15 GNDA 0.358463f
C325 1st_Vout_1.t14 GNDA 0.35246f
C326 1st_Vout_1.t26 GNDA 0.35246f
C327 1st_Vout_1.t25 GNDA 0.358463f
C328 1st_Vout_1.t31 GNDA 0.358463f
C329 1st_Vout_1.t13 GNDA 0.35246f
C330 1st_Vout_1.t35 GNDA 0.35246f
C331 1st_Vout_1.t19 GNDA 0.023025f
C332 1st_Vout_1.n10 GNDA 0.022249f
C333 1st_Vout_1.t30 GNDA 0.013423f
C334 1st_Vout_1.t24 GNDA 0.013423f
C335 1st_Vout_1.n11 GNDA 0.029862f
C336 1st_Vout_1.n12 GNDA 0.021343f
C337 V_mir2.t12 GNDA 0.019293f
C338 V_mir2.t6 GNDA 0.019293f
C339 V_mir2.t10 GNDA 0.019293f
C340 V_mir2.n0 GNDA 0.044322f
C341 V_mir2.t5 GNDA 0.02939f
C342 V_mir2.t9 GNDA 0.023151f
C343 V_mir2.t18 GNDA 0.023151f
C344 V_mir2.t17 GNDA 0.037369f
C345 V_mir2.n1 GNDA 0.041731f
C346 V_mir2.n2 GNDA 0.028507f
C347 V_mir2.n3 GNDA 0.044354f
C348 V_mir2.n4 GNDA 0.109787f
C349 V_mir2.t4 GNDA 0.019293f
C350 V_mir2.t8 GNDA 0.019293f
C351 V_mir2.n5 GNDA 0.044322f
C352 V_mir2.t3 GNDA 0.02939f
C353 V_mir2.t7 GNDA 0.023151f
C354 V_mir2.t19 GNDA 0.023151f
C355 V_mir2.t20 GNDA 0.037369f
C356 V_mir2.n6 GNDA 0.041731f
C357 V_mir2.n7 GNDA 0.028507f
C358 V_mir2.n8 GNDA 0.044354f
C359 V_mir2.n9 GNDA 0.084938f
C360 V_mir2.n10 GNDA 0.025223f
C361 V_mir2.t1 GNDA 0.041163f
C362 V_mir2.n11 GNDA 0.027381f
C363 V_mir2.n12 GNDA 0.451535f
C364 V_mir2.n13 GNDA 0.146338f
C365 V_mir2.n14 GNDA 0.051125f
C366 V_mir2.n15 GNDA 0.381359f
C367 V_mir2.t11 GNDA 0.02939f
C368 V_mir2.t13 GNDA 0.023151f
C369 V_mir2.t22 GNDA 0.023151f
C370 V_mir2.t21 GNDA 0.037369f
C371 V_mir2.n16 GNDA 0.041731f
C372 V_mir2.n17 GNDA 0.028507f
C373 V_mir2.n18 GNDA 0.044354f
C374 V_mir2.n19 GNDA 0.110886f
C375 V_mir2.n20 GNDA 0.044322f
C376 V_mir2.t14 GNDA 0.019293f
C377 NFET_GATE_10uA.t4 GNDA 0.01675f
C378 NFET_GATE_10uA.t1 GNDA 0.01675f
C379 NFET_GATE_10uA.t2 GNDA 0.01675f
C380 NFET_GATE_10uA.n0 GNDA 0.183066f
C381 NFET_GATE_10uA.t21 GNDA 0.016332f
C382 NFET_GATE_10uA.t15 GNDA 0.016332f
C383 NFET_GATE_10uA.t10 GNDA 0.016332f
C384 NFET_GATE_10uA.t20 GNDA 0.016332f
C385 NFET_GATE_10uA.t14 GNDA 0.016332f
C386 NFET_GATE_10uA.t9 GNDA 0.016332f
C387 NFET_GATE_10uA.t19 GNDA 0.024143f
C388 NFET_GATE_10uA.n1 GNDA 0.029878f
C389 NFET_GATE_10uA.n2 GNDA 0.021357f
C390 NFET_GATE_10uA.n3 GNDA 0.018081f
C391 NFET_GATE_10uA.t23 GNDA 0.016332f
C392 NFET_GATE_10uA.t16 GNDA 0.016332f
C393 NFET_GATE_10uA.t7 GNDA 0.016332f
C394 NFET_GATE_10uA.t8 GNDA 0.024143f
C395 NFET_GATE_10uA.n4 GNDA 0.029878f
C396 NFET_GATE_10uA.n5 GNDA 0.021357f
C397 NFET_GATE_10uA.n6 GNDA 0.018081f
C398 NFET_GATE_10uA.t11 GNDA 0.016332f
C399 NFET_GATE_10uA.t17 GNDA 0.024143f
C400 NFET_GATE_10uA.n7 GNDA 0.026602f
C401 NFET_GATE_10uA.n8 GNDA 0.029239f
C402 NFET_GATE_10uA.t18 GNDA 0.016332f
C403 NFET_GATE_10uA.t13 GNDA 0.024143f
C404 NFET_GATE_10uA.n9 GNDA 0.026602f
C405 NFET_GATE_10uA.t6 GNDA 0.016332f
C406 NFET_GATE_10uA.t5 GNDA 0.016332f
C407 NFET_GATE_10uA.t12 GNDA 0.016332f
C408 NFET_GATE_10uA.t22 GNDA 0.024143f
C409 NFET_GATE_10uA.n10 GNDA 0.029878f
C410 NFET_GATE_10uA.n11 GNDA 0.021357f
C411 NFET_GATE_10uA.n12 GNDA 0.018081f
C412 NFET_GATE_10uA.n13 GNDA 0.029239f
C413 NFET_GATE_10uA.n14 GNDA 0.67829f
C414 NFET_GATE_10uA.n15 GNDA 0.024928f
C415 NFET_GATE_10uA.n16 GNDA 0.018081f
C416 NFET_GATE_10uA.n17 GNDA 0.021357f
C417 NFET_GATE_10uA.n18 GNDA 0.029878f
C418 NFET_GATE_10uA.t3 GNDA 0.038251f
C419 NFET_GATE_10uA.n19 GNDA 1.72301f
C420 NFET_GATE_10uA.n20 GNDA 0.047154f
C421 NFET_GATE_10uA.t0 GNDA 0.01675f
C422 VDDA.n1 GNDA 0.035114f
C423 VDDA.t129 GNDA 0.014539f
C424 VDDA.n3 GNDA 0.035114f
C425 VDDA.n4 GNDA 0.038803f
C426 VDDA.n5 GNDA 0.024404f
C427 VDDA.t120 GNDA 0.03643f
C428 VDDA.t136 GNDA 0.012055f
C429 VDDA.n6 GNDA 0.024404f
C430 VDDA.n7 GNDA 0.040597f
C431 VDDA.n8 GNDA 0.024404f
C432 VDDA.n9 GNDA 0.038803f
C433 VDDA.n11 GNDA 0.03511f
C434 VDDA.t170 GNDA 0.014546f
C435 VDDA.n13 GNDA 0.03511f
C436 VDDA.n15 GNDA 0.047561f
C437 VDDA.t135 GNDA 0.014546f
C438 VDDA.n16 GNDA 0.016575f
C439 VDDA.t164 GNDA 0.014546f
C440 VDDA.n17 GNDA 0.04151f
C441 VDDA.t163 GNDA 0.043746f
C442 VDDA.t93 GNDA 0.030706f
C443 VDDA.t109 GNDA 0.030706f
C444 VDDA.t134 GNDA 0.043746f
C445 VDDA.n18 GNDA 0.04151f
C446 VDDA.n19 GNDA 0.016152f
C447 VDDA.n20 GNDA 0.026432f
C448 VDDA.n21 GNDA 0.025834f
C449 VDDA.n22 GNDA 0.016152f
C450 VDDA.t155 GNDA 0.014546f
C451 VDDA.n23 GNDA 0.04151f
C452 VDDA.t154 GNDA 0.043746f
C453 VDDA.t87 GNDA 0.030706f
C454 VDDA.t101 GNDA 0.030706f
C455 VDDA.t107 GNDA 0.030706f
C456 VDDA.t95 GNDA 0.030706f
C457 VDDA.t169 GNDA 0.043746f
C458 VDDA.n24 GNDA 0.04151f
C459 VDDA.n25 GNDA 0.016401f
C460 VDDA.n26 GNDA 0.03042f
C461 VDDA.n27 GNDA 0.028625f
C462 VDDA.n28 GNDA 0.023301f
C463 VDDA.t139 GNDA 0.028454f
C464 VDDA.n29 GNDA 0.077857f
C465 VDDA.t137 GNDA 0.07047f
C466 VDDA.t113 GNDA 0.052639f
C467 VDDA.t97 GNDA 0.052639f
C468 VDDA.t85 GNDA 0.052639f
C469 VDDA.t99 GNDA 0.052639f
C470 VDDA.t119 GNDA 0.07047f
C471 VDDA.n30 GNDA 0.077857f
C472 VDDA.t118 GNDA 0.012055f
C473 VDDA.n31 GNDA 0.023301f
C474 VDDA.n32 GNDA 0.028625f
C475 VDDA.n33 GNDA 0.03042f
C476 VDDA.n34 GNDA 0.016152f
C477 VDDA.t167 GNDA 0.014539f
C478 VDDA.n35 GNDA 0.041518f
C479 VDDA.t166 GNDA 0.043746f
C480 VDDA.t89 GNDA 0.030706f
C481 VDDA.t103 GNDA 0.030706f
C482 VDDA.t91 GNDA 0.030706f
C483 VDDA.t105 GNDA 0.030706f
C484 VDDA.t128 GNDA 0.043746f
C485 VDDA.n36 GNDA 0.041518f
C486 VDDA.n37 GNDA 0.016152f
C487 VDDA.n38 GNDA 0.080642f
C488 VDDA.n39 GNDA 1.73385f
C489 VDDA.t24 GNDA 0.211762f
C490 VDDA.t30 GNDA 0.222918f
C491 VDDA.t74 GNDA 0.223726f
C492 VDDA.t14 GNDA 0.211762f
C493 VDDA.t75 GNDA 0.222918f
C494 VDDA.t15 GNDA 0.223726f
C495 VDDA.t41 GNDA 0.211762f
C496 VDDA.t12 GNDA 0.222918f
C497 VDDA.t211 GNDA 0.223726f
C498 VDDA.t21 GNDA 0.211762f
C499 VDDA.t78 GNDA 0.222918f
C500 VDDA.t51 GNDA 0.223726f
C501 VDDA.t48 GNDA 0.211762f
C502 VDDA.t27 GNDA 0.222918f
C503 VDDA.t16 GNDA 0.223726f
C504 VDDA.n40 GNDA 0.149422f
C505 VDDA.t23 GNDA 0.118993f
C506 VDDA.n41 GNDA 0.162126f
C507 VDDA.t13 GNDA 0.118993f
C508 VDDA.n42 GNDA 0.162126f
C509 VDDA.t22 GNDA 0.118993f
C510 VDDA.n43 GNDA 0.162126f
C511 VDDA.t191 GNDA 0.118993f
C512 VDDA.n44 GNDA 0.162126f
C513 VDDA.t206 GNDA 0.208455f
C514 VDDA.n45 GNDA 2.14591f
C515 VDDA.t215 GNDA 0.505599f
C516 VDDA.t214 GNDA 0.504696f
C517 VDDA.n46 GNDA 0.107884f
C518 VDDA.t213 GNDA 0.504762f
C519 VDDA.n47 GNDA 0.068683f
C520 VDDA.t212 GNDA 0.504762f
C521 VDDA.n48 GNDA 0.108311f
C522 VDDA.n49 GNDA 0.40581f
C523 VDDA.n50 GNDA 0.010047f
C524 VDDA.n51 GNDA 0.040598f
C525 VDDA.t132 GNDA 0.014531f
C526 VDDA.t126 GNDA 0.014531f
C527 VDDA.n52 GNDA 0.010047f
C528 VDDA.n53 GNDA 0.040598f
C529 VDDA.n54 GNDA 0.010047f
C530 VDDA.n55 GNDA 0.040598f
C531 VDDA.n56 GNDA 0.010047f
C532 VDDA.n57 GNDA 0.040598f
C533 VDDA.n58 GNDA 0.010047f
C534 VDDA.n59 GNDA 0.040598f
C535 VDDA.n60 GNDA 0.010047f
C536 VDDA.n61 GNDA 0.040598f
C537 VDDA.n62 GNDA 0.010047f
C538 VDDA.n63 GNDA 0.040598f
C539 VDDA.n64 GNDA 0.010047f
C540 VDDA.n65 GNDA 0.040598f
C541 VDDA.n66 GNDA 0.010047f
C542 VDDA.n67 GNDA 0.040598f
C543 VDDA.n68 GNDA 0.010047f
C544 VDDA.n69 GNDA 0.040598f
C545 VDDA.t158 GNDA 0.014531f
C546 VDDA.t148 GNDA 0.014531f
C547 VDDA.n70 GNDA 0.010047f
C548 VDDA.n71 GNDA 0.040598f
C549 VDDA.n72 GNDA 0.010047f
C550 VDDA.n73 GNDA 0.040598f
C551 VDDA.n74 GNDA 0.010047f
C552 VDDA.n75 GNDA 0.040598f
C553 VDDA.n76 GNDA 0.010047f
C554 VDDA.n77 GNDA 0.040598f
C555 VDDA.n78 GNDA 0.010047f
C556 VDDA.n79 GNDA 0.040598f
C557 VDDA.n80 GNDA 0.010047f
C558 VDDA.n81 GNDA 0.040598f
C559 VDDA.n82 GNDA 0.010047f
C560 VDDA.n83 GNDA 0.040598f
C561 VDDA.n84 GNDA 0.010047f
C562 VDDA.n85 GNDA 0.066091f
C563 VDDA.t146 GNDA 0.014962f
C564 VDDA.n87 GNDA 0.053494f
C565 VDDA.t147 GNDA 0.04579f
C566 VDDA.t25 GNDA 0.033498f
C567 VDDA.t42 GNDA 0.033498f
C568 VDDA.t202 GNDA 0.033498f
C569 VDDA.t209 GNDA 0.033498f
C570 VDDA.t35 GNDA 0.033498f
C571 VDDA.t198 GNDA 0.033498f
C572 VDDA.t10 GNDA 0.033498f
C573 VDDA.t81 GNDA 0.033498f
C574 VDDA.t33 GNDA 0.033498f
C575 VDDA.t183 GNDA 0.033498f
C576 VDDA.t4 GNDA 0.033498f
C577 VDDA.t185 GNDA 0.033498f
C578 VDDA.t62 GNDA 0.033498f
C579 VDDA.t196 GNDA 0.033498f
C580 VDDA.t83 GNDA 0.033498f
C581 VDDA.t31 GNDA 0.033498f
C582 VDDA.t28 GNDA 0.033498f
C583 VDDA.t58 GNDA 0.033498f
C584 VDDA.t157 GNDA 0.046573f
C585 VDDA.n88 GNDA 0.044543f
C586 VDDA.n89 GNDA 0.016582f
C587 VDDA.n90 GNDA 0.029705f
C588 VDDA.n91 GNDA 0.037274f
C589 VDDA.t124 GNDA 0.014962f
C590 VDDA.n93 GNDA 0.053494f
C591 VDDA.t125 GNDA 0.04579f
C592 VDDA.t173 GNDA 0.033498f
C593 VDDA.t187 GNDA 0.033498f
C594 VDDA.t6 GNDA 0.033498f
C595 VDDA.t68 GNDA 0.033498f
C596 VDDA.t46 GNDA 0.033498f
C597 VDDA.t171 GNDA 0.033498f
C598 VDDA.t179 GNDA 0.033498f
C599 VDDA.t19 GNDA 0.033498f
C600 VDDA.t8 GNDA 0.033498f
C601 VDDA.t189 GNDA 0.033498f
C602 VDDA.t70 GNDA 0.033498f
C603 VDDA.t181 GNDA 0.033498f
C604 VDDA.t175 GNDA 0.033498f
C605 VDDA.t53 GNDA 0.033498f
C606 VDDA.t0 GNDA 0.033498f
C607 VDDA.t192 GNDA 0.033498f
C608 VDDA.t204 GNDA 0.033498f
C609 VDDA.t177 GNDA 0.033498f
C610 VDDA.t131 GNDA 0.04579f
C611 VDDA.n94 GNDA 0.0536f
C612 VDDA.t130 GNDA 0.014956f
C613 VDDA.n96 GNDA 0.076414f
C614 VDDA.n97 GNDA 0.132736f
C615 VDDA.t117 GNDA 0.042389f
C616 VDDA.n98 GNDA 0.120669f
C617 VDDA.t115 GNDA 0.057046f
C618 VDDA.t161 GNDA 0.042389f
C619 VDDA.t116 GNDA 0.137557f
C620 VDDA.t194 GNDA 0.12741f
C621 VDDA.t49 GNDA 0.12741f
C622 VDDA.t55 GNDA 0.12741f
C623 VDDA.t72 GNDA 0.12741f
C624 VDDA.t37 GNDA 0.12741f
C625 VDDA.t66 GNDA 0.12741f
C626 VDDA.t200 GNDA 0.12741f
C627 VDDA.t2 GNDA 0.12741f
C628 VDDA.t76 GNDA 0.12741f
C629 VDDA.t17 GNDA 0.12741f
C630 VDDA.t39 GNDA 0.12741f
C631 VDDA.t207 GNDA 0.12741f
C632 VDDA.t44 GNDA 0.12741f
C633 VDDA.t60 GNDA 0.12741f
C634 VDDA.t64 GNDA 0.12741f
C635 VDDA.t79 GNDA 0.12741f
C636 VDDA.t160 GNDA 0.137557f
C637 VDDA.n99 GNDA 0.120669f
C638 VDDA.n100 GNDA 0.019858f
C639 VDDA.t123 GNDA 0.014531f
C640 VDDA.n101 GNDA 0.041786f
C641 VDDA.t122 GNDA 0.043746f
C642 VDDA.t52 GNDA 0.030706f
C643 VDDA.t57 GNDA 0.030706f
C644 VDDA.t141 GNDA 0.045332f
C645 VDDA.t142 GNDA 0.016288f
C646 VDDA.n102 GNDA 0.047845f
C647 VDDA.n103 GNDA 0.016634f
C648 VDDA.n104 GNDA 0.077576f
C649 VDDA.t159 GNDA 0.057046f
C650 VDDA.n105 GNDA 0.045873f
C651 VDDA.t65 GNDA 0.011963f
C652 VDDA.t80 GNDA 0.011963f
C653 VDDA.n106 GNDA 0.037979f
C654 VDDA.n107 GNDA 0.037667f
C655 VDDA.t45 GNDA 0.011963f
C656 VDDA.t61 GNDA 0.011963f
C657 VDDA.n108 GNDA 0.037979f
C658 VDDA.n109 GNDA 0.03739f
C659 VDDA.t40 GNDA 0.011963f
C660 VDDA.t208 GNDA 0.011963f
C661 VDDA.n110 GNDA 0.037979f
C662 VDDA.n111 GNDA 0.03739f
C663 VDDA.t77 GNDA 0.011963f
C664 VDDA.t18 GNDA 0.011963f
C665 VDDA.n112 GNDA 0.037979f
C666 VDDA.n113 GNDA 0.03739f
C667 VDDA.t201 GNDA 0.011963f
C668 VDDA.t3 GNDA 0.011963f
C669 VDDA.n114 GNDA 0.037979f
C670 VDDA.n115 GNDA 0.03739f
C671 VDDA.t38 GNDA 0.011963f
C672 VDDA.t67 GNDA 0.011963f
C673 VDDA.n116 GNDA 0.037979f
C674 VDDA.n117 GNDA 0.03739f
C675 VDDA.t56 GNDA 0.011963f
C676 VDDA.t73 GNDA 0.011963f
C677 VDDA.n118 GNDA 0.037979f
C678 VDDA.n119 GNDA 0.03739f
C679 VDDA.t195 GNDA 0.011963f
C680 VDDA.t50 GNDA 0.011963f
C681 VDDA.n120 GNDA 0.037979f
C682 VDDA.n121 GNDA 0.037667f
C683 VDDA.n122 GNDA 0.047284f
C684 VDDA.t143 GNDA 0.011471f
C685 VDDA.n123 GNDA 0.022519f
C686 VDDA.t152 GNDA 0.028454f
C687 VDDA.t145 GNDA 0.028454f
C688 VDDA.n124 GNDA 0.077857f
C689 VDDA.t144 GNDA 0.07047f
C690 VDDA.t111 GNDA 0.052639f
C691 VDDA.t150 GNDA 0.07047f
C692 VDDA.n125 GNDA 0.077857f
C693 VDDA.t149 GNDA 0.011742f
C694 VDDA.n126 GNDA 0.022552f
C695 VDDA.n127 GNDA 0.034557f
C696 VDDA.n128 GNDA 0.023711f
C697 VDDA.n129 GNDA 0.036924f
C698 VDDA.n130 GNDA 0.099782f
C699 VDDA.n131 GNDA 0.108299f
C700 PFET_GATE_10uA.t21 GNDA 0.020941f
C701 PFET_GATE_10uA.t14 GNDA 0.030957f
C702 PFET_GATE_10uA.n0 GNDA 0.034111f
C703 PFET_GATE_10uA.t15 GNDA 0.020941f
C704 PFET_GATE_10uA.t22 GNDA 0.030957f
C705 PFET_GATE_10uA.n1 GNDA 0.034111f
C706 PFET_GATE_10uA.n2 GNDA 0.034221f
C707 PFET_GATE_10uA.t0 GNDA 0.472888f
C708 PFET_GATE_10uA.t11 GNDA 0.055245f
C709 PFET_GATE_10uA.n3 GNDA 1.93329f
C710 PFET_GATE_10uA.t2 GNDA 0.021478f
C711 PFET_GATE_10uA.t4 GNDA 0.021478f
C712 PFET_GATE_10uA.n4 GNDA 0.054974f
C713 PFET_GATE_10uA.t9 GNDA 0.021478f
C714 PFET_GATE_10uA.t8 GNDA 0.021478f
C715 PFET_GATE_10uA.n5 GNDA 0.053578f
C716 PFET_GATE_10uA.n6 GNDA 0.522912f
C717 PFET_GATE_10uA.t6 GNDA 0.021478f
C718 PFET_GATE_10uA.t7 GNDA 0.021478f
C719 PFET_GATE_10uA.n7 GNDA 0.053578f
C720 PFET_GATE_10uA.n8 GNDA 0.29652f
C721 PFET_GATE_10uA.t1 GNDA 0.31282f
C722 PFET_GATE_10uA.n9 GNDA 0.606455f
C723 PFET_GATE_10uA.t5 GNDA 0.021478f
C724 PFET_GATE_10uA.t3 GNDA 0.021478f
C725 PFET_GATE_10uA.n10 GNDA 0.051929f
C726 PFET_GATE_10uA.n11 GNDA 0.276412f
C727 PFET_GATE_10uA.n12 GNDA 0.777893f
C728 PFET_GATE_10uA.n13 GNDA 0.762338f
C729 PFET_GATE_10uA.t12 GNDA 0.020941f
C730 PFET_GATE_10uA.t20 GNDA 0.031004f
C731 PFET_GATE_10uA.n14 GNDA 0.06665f
C732 PFET_GATE_10uA.t13 GNDA 0.020941f
C733 PFET_GATE_10uA.t19 GNDA 0.030957f
C734 PFET_GATE_10uA.n15 GNDA 0.034111f
C735 PFET_GATE_10uA.t16 GNDA 0.020941f
C736 PFET_GATE_10uA.t23 GNDA 0.030957f
C737 PFET_GATE_10uA.n16 GNDA 0.034111f
C738 PFET_GATE_10uA.n17 GNDA 0.031825f
C739 PFET_GATE_10uA.n18 GNDA 0.658801f
C740 PFET_GATE_10uA.t17 GNDA 0.048508f
C741 PFET_GATE_10uA.t24 GNDA 0.045105f
C742 PFET_GATE_10uA.t18 GNDA 0.045105f
C743 PFET_GATE_10uA.t10 GNDA 0.05477f
C744 PFET_GATE_10uA.n19 GNDA 0.05477f
C745 PFET_GATE_10uA.n20 GNDA 0.03124f
C746 PFET_GATE_10uA.n21 GNDA 0.053217f
C747 cap_res2.t7 GNDA 0.340877f
C748 cap_res2.t17 GNDA 0.358835f
C749 cap_res2.t1 GNDA 0.360135f
C750 cap_res2.t15 GNDA 0.340877f
C751 cap_res2.t6 GNDA 0.358835f
C752 cap_res2.t19 GNDA 0.360135f
C753 cap_res2.t2 GNDA 0.340877f
C754 cap_res2.t10 GNDA 0.358835f
C755 cap_res2.t4 GNDA 0.360135f
C756 cap_res2.t13 GNDA 0.340877f
C757 cap_res2.t5 GNDA 0.358835f
C758 cap_res2.t16 GNDA 0.360135f
C759 cap_res2.t8 GNDA 0.340877f
C760 cap_res2.t20 GNDA 0.358835f
C761 cap_res2.t11 GNDA 0.360135f
C762 cap_res2.n0 GNDA 0.240527f
C763 cap_res2.t9 GNDA 0.191544f
C764 cap_res2.n1 GNDA 0.260978f
C765 cap_res2.t14 GNDA 0.191544f
C766 cap_res2.n2 GNDA 0.260978f
C767 cap_res2.t3 GNDA 0.191544f
C768 cap_res2.n3 GNDA 0.260978f
C769 cap_res2.t18 GNDA 0.191544f
C770 cap_res2.n4 GNDA 0.260978f
C771 cap_res2.t12 GNDA 0.179549f
C772 cap_res2.t0 GNDA 0.085169f
C773 1st_Vout_2.n0 GNDA 0.722974f
C774 1st_Vout_2.n1 GNDA 1.43086f
C775 1st_Vout_2.n2 GNDA 0.104357f
C776 1st_Vout_2.n3 GNDA 1.45767f
C777 1st_Vout_2.t27 GNDA 0.293375f
C778 1st_Vout_2.t25 GNDA 0.288462f
C779 1st_Vout_2.t11 GNDA 0.293375f
C780 1st_Vout_2.t23 GNDA 0.288462f
C781 1st_Vout_2.t18 GNDA 0.293375f
C782 1st_Vout_2.t17 GNDA 0.288462f
C783 1st_Vout_2.t31 GNDA 0.293375f
C784 1st_Vout_2.t15 GNDA 0.288462f
C785 1st_Vout_2.t35 GNDA 0.293375f
C786 1st_Vout_2.t34 GNDA 0.288462f
C787 1st_Vout_2.t24 GNDA 0.293375f
C788 1st_Vout_2.t33 GNDA 0.288462f
C789 1st_Vout_2.t16 GNDA 0.293375f
C790 1st_Vout_2.t13 GNDA 0.288462f
C791 1st_Vout_2.t30 GNDA 0.293375f
C792 1st_Vout_2.t12 GNDA 0.288462f
C793 1st_Vout_2.t28 GNDA 0.293375f
C794 1st_Vout_2.t19 GNDA 0.288462f
C795 1st_Vout_2.t36 GNDA 0.288462f
C796 1st_Vout_2.t14 GNDA 0.288462f
C797 1st_Vout_2.t22 GNDA 0.018845f
C798 1st_Vout_2.n4 GNDA 0.018209f
C799 1st_Vout_2.t26 GNDA 0.010986f
C800 1st_Vout_2.t20 GNDA 0.010986f
C801 1st_Vout_2.n5 GNDA 0.024439f
C802 1st_Vout_2.n6 GNDA 0.017468f
C803 1st_Vout_2.t8 GNDA 0.015189f
C804 1st_Vout_2.n7 GNDA 0.010417f
C805 1st_Vout_2.n8 GNDA 0.157567f
C806 1st_Vout_2.t21 GNDA 0.010986f
C807 1st_Vout_2.t32 GNDA 0.010986f
C808 1st_Vout_2.n10 GNDA 0.024439f
C809 1st_Vout_2.n11 GNDA 0.018209f
C810 1st_Vout_2.t29 GNDA 0.017243f
.ends

