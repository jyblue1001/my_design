* PEX produced on Sat Feb  1 12:21:39 PM CET 2025 using /foss/tools/osic-multitool/iic-pex.sh with m=3 and s=1
* NGSPICE file created from vco2_2.ext - technology: sky130A

.subckt vco2_2
X0 a_82_186.t1 a_38_n62.t2 V_OSC.t1 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.22
X1 a_636_n552.t2 V_CONT GNDA.t13 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X2 a_1190_n552.t1 V_OSC.t2 a_592_n62.t1 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.22
X3 a_82_186.t0 GNDA.t14 VDDA.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.15
X4 GNDA.t12 V_CONT a_n746_764.t2 GNDA.t11 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X5 VDDA.t6 a_n746_764.t0 a_n746_764.t1 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X6 a_82_n552.t1 a_38_n62.t3 V_OSC.t0 GNDA.t7 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.22
X7 a_1190_n552.t0 VDDA.t17 GNDA.t5 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.15
X8 a_1190_n552.t2 V_CONT GNDA.t10 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X9 a_636_186.t1 a_592_n62.t2 a_38_n62.t0 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.22
X10 a_82_n552.t0 VDDA.t18 GNDA.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.15
X11 a_82_n552.t2 V_CONT GNDA.t9 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X12 a_636_186.t0 a_n746_764.t3 VDDA.t14 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X13 a_636_n552.t1 a_592_n62.t3 a_38_n62.t1 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.22
X14 a_82_186.t2 a_n746_764.t4 VDDA.t16 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X15 a_1190_186.t0 V_OSC.t3 a_592_n62.t0 VDDA.t12 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.22
X16 a_1190_186.t1 a_n746_764.t5 VDDA.t4 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=1.5
X17 a_636_186.t2 GNDA.t15 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.15
X18 a_1190_186.t2 GNDA.t16 VDDA.t2 VDDA.t1 sky130_fd_pr__pfet_01v8 ad=0.43 pd=2.72 as=0.43 ps=2.72 w=0.86 l=0.15
X19 a_636_n552.t0 VDDA.t19 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.215 pd=1.86 as=0.215 ps=1.86 w=0.43 l=0.15
R0 a_38_n62.n1 a_38_n62.n0 770.567
R1 a_38_n62.t0 a_38_n62.n1 374.728
R2 a_38_n62.n1 a_38_n62.t1 271.567
R3 a_38_n62.n0 a_38_n62.t2 135.837
R4 a_38_n62.n0 a_38_n62.t3 84.3505
R5 V_OSC.n1 V_OSC.n0 2387.29
R6 V_OSC.t1 V_OSC.n1 374.728
R7 V_OSC.n1 V_OSC.t0 271.567
R8 V_OSC.n0 V_OSC.t3 135.837
R9 V_OSC.n0 V_OSC.t2 84.3505
R10 a_82_186.n0 a_82_186.t1 398.087
R11 a_82_186.t0 a_82_186.n0 349.767
R12 a_82_186.n0 a_82_186.t2 212.364
R13 VDDA.n1 VDDA.t17 1007.38
R14 VDDA.n2 VDDA.t18 618.567
R15 VDDA.t15 VDDA.t5 488.219
R16 VDDA.t9 VDDA.t3 480.288
R17 VDDA.n3 VDDA.n2 357.406
R18 VDDA VDDA.t2 354.445
R19 VDDA VDDA.t8 354.418
R20 VDDA.n3 VDDA.t10 349.767
R21 VDDA.n0 VDDA.t7 341.048
R22 VDDA.n2 VDDA.n1 308.481
R23 VDDA.n3 VDDA.n0 185
R24 VDDA VDDA.t6 143.486
R25 VDDA VDDA.t16 143.486
R26 VDDA VDDA.t14 143.486
R27 VDDA VDDA.t4 143.486
R28 VDDA.n0 VDDA.t13 139.239
R29 VDDA.n1 VDDA.t19 117.287
R30 VDDA.t12 VDDA.t1 6.16933
R31 VDDA.t0 VDDA.t9 6.16933
R32 VDDA.t7 VDDA.t11 6.16933
R33 VDDA VDDA.n3 2.50857
R34 VDDA.t3 VDDA.t12 1.76302
R35 VDDA.t13 VDDA.t0 1.76302
R36 VDDA.t11 VDDA.t15 1.76302
R37 GNDA.t7 GNDA.t11 2665.66
R38 GNDA.t6 GNDA.t2 2599.14
R39 GNDA.n1 GNDA.t0 1848.38
R40 GNDA.n4 GNDA.n1 1170
R41 GNDA.n2 GNDA.t14 1076.47
R42 GNDA.n1 GNDA.t8 750.756
R43 GNDA.n3 GNDA.n2 504.493
R44 GNDA.n3 GNDA.t16 491.64
R45 GNDA.n4 GNDA.n3 352.723
R46 GNDA GNDA.t3 264.067
R47 GNDA GNDA.t1 264.067
R48 GNDA.n0 GNDA.t5 258.902
R49 GNDA.n2 GNDA.t15 186.374
R50 GNDA GNDA.t9 127.15
R51 GNDA GNDA.t13 127.15
R52 GNDA GNDA.t10 127.15
R53 GNDA GNDA.t12 127.15
R54 GNDA.t8 GNDA.t4 33.2618
R55 GNDA.t0 GNDA.t6 33.2618
R56 GNDA.t2 GNDA.t7 33.2618
R57 GNDA.n0 GNDA.n4 4.13491
R58 GNDA.n0 GNDA 3.12085
R59 a_636_n552.n0 a_636_n552.t1 289.967
R60 a_636_n552.n0 a_636_n552.t0 254.768
R61 a_636_n552.t2 a_636_n552.n0 161.701
R62 a_592_n62.n1 a_592_n62.n0 776.994
R63 a_592_n62.t0 a_592_n62.n1 374.728
R64 a_592_n62.n1 a_592_n62.t1 271.567
R65 a_592_n62.n0 a_592_n62.t2 135.837
R66 a_592_n62.n0 a_592_n62.t3 84.3505
R67 a_1190_n552.n0 a_1190_n552.t1 289.967
R68 a_1190_n552.n0 a_1190_n552.t0 254.768
R69 a_1190_n552.t2 a_1190_n552.n0 161.701
R70 a_n746_764.t2 a_n746_764.n2 466.82
R71 a_n746_764.n2 a_n746_764.t0 225.869
R72 a_n746_764.n2 a_n746_764.t1 225.786
R73 a_n746_764.t0 a_n746_764.n1 188.501
R74 a_n746_764.n0 a_n746_764.t5 188.501
R75 a_n746_764.n1 a_n746_764.n0 107.442
R76 a_n746_764.n1 a_n746_764.t4 81.0592
R77 a_n746_764.n0 a_n746_764.t3 81.0592
R78 a_82_n552.n0 a_82_n552.t1 289.967
R79 a_82_n552.n0 a_82_n552.t0 254.768
R80 a_82_n552.t2 a_82_n552.n0 161.701
R81 a_636_186.n0 a_636_186.t1 398.087
R82 a_636_186.t2 a_636_186.n0 349.767
R83 a_636_186.n0 a_636_186.t0 212.364
R84 a_1190_186.n0 a_1190_186.t0 398.087
R85 a_1190_186.t2 a_1190_186.n0 349.767
R86 a_1190_186.n0 a_1190_186.t1 212.364
C0 VDDA V_CONT 0.063762f
C1 V_CONT GNDA 1.51311f
C2 VDDA GNDA 10.900789f
C3 a_n746_764.t1 GNDA 0.153998f
C4 a_n746_764.t5 GNDA 0.465957f
C5 a_n746_764.t3 GNDA 0.365904f
C6 a_n746_764.n0 GNDA 0.27731f
C7 a_n746_764.t4 GNDA 0.365904f
C8 a_n746_764.n1 GNDA 0.276948f
C9 a_n746_764.t0 GNDA 0.518928f
C10 a_n746_764.n2 GNDA 0.237652f
C11 a_n746_764.t2 GNDA 0.137401f
C12 VDDA.t4 GNDA 0.022852f
C13 VDDA.t1 GNDA 0.195936f
C14 VDDA.t3 GNDA 0.191046f
C15 VDDA.t9 GNDA 0.192792f
C16 VDDA.t13 GNDA 0.055882f
C17 VDDA.t5 GNDA 0.444959f
C18 VDDA.t15 GNDA 0.194189f
C19 VDDA.t7 GNDA 0.137609f
C20 VDDA.n0 GNDA 0.184775f
C21 VDDA.n2 GNDA 0.015998f
C22 VDDA.n3 GNDA 0.023552f
C23 VDDA.t14 GNDA 0.022852f
C24 VDDA.t16 GNDA 0.022852f
C25 VDDA.t6 GNDA 0.022852f
.ends

