* NGSPICE file created from nor2.ext - technology: sky130A

**.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

**.subckt nor2
Xsky130_fd_sc_hd__nor2_1_1 sky130_fd_sc_hd__nor2_1_1/A sky130_fd_sc_hd__nor2_1_1/B
+ sky130_fd_sc_hd__nor2_1_1/VGND VSUBS sky130_fd_sc_hd__nor2_1_1/VPB sky130_fd_sc_hd__nor2_1_1/VPWR
+ sky130_fd_sc_hd__nor2_1_1/Y sky130_fd_sc_hd__nor2_1
Xsky130_fd_sc_hd__nor2_1_0 sky130_fd_sc_hd__nor2_1_0/A sky130_fd_sc_hd__nor2_1_1/Y
+ sky130_fd_sc_hd__nor2_1_1/VGND VSUBS sky130_fd_sc_hd__nor2_1_1/VPB sky130_fd_sc_hd__nor2_1_1/VPWR
+ sky130_fd_sc_hd__nor2_1_1/B sky130_fd_sc_hd__nor2_1
.ends

