* PEX produced on Mon Feb 17 06:40:18 PM CET 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from pfd_cp_lf_magic.ext - technology: sky130A

.subckt pfd_cp_lf_magic V_OUT VDDA GNDA F_REF F_VCO I_IN
X0 a_6400_6270.t2 a_6400_6270.t1 GNDA.t92 GNDA.t91 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X1 VDDA.t75 opamp_cell_4_0.n_left.t6 opamp_cell_4_0.n_right.t4 VDDA.t74 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X2 VDDA.t83 opamp_cell_4_0.n_right.t5 pfd_8_0.opamp_out.t9 VDDA.t82 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X3 GNDA.t31 a_6380_5710.t4 a_6380_5710.t5 GNDA.t30 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X4 a_6500_6300.t8 a_6500_6300.t6 a_6500_6300.t7 GNDA.t29 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X5 pfd_8_0.DOWN_b.t1 VDDA.t129 pfd_8_0.DOWN_PFD_b.t3 GNDA.t39 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X6 a_870_1400.t1 pfd_8_0.QA_b.t3 VDDA.t124 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X7 a_6500_6300.t12 a_6400_6270.t9 GNDA.t90 GNDA.t89 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X8 a_6150_5090.t8 opamp_cell_4_0.p_bias.t9 VDDA.t63 VDDA.t62 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X9 pfd_8_0.DOWN.t1 pfd_8_0.DOWN_b.t2 VDDA.t8 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X10 V_OUT.t4 pfd_8_0.UP_input.t3 VDDA.t48 VDDA.t47 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X11 opamp_cell_4_0.p_bias.t7 opamp_cell_4_0.p_bias.t6 VDDA.t55 VDDA.t54 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X12 a_6150_5090.t11 V_OUT.t8 a_6380_5710.t1 VDDA.t53 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X13 VDDA.t117 VDDA.t114 VDDA.t116 VDDA.t115 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X14 a_2350_1400.t0 pfd_8_0.before_Reset.t3 GNDA.t74 GNDA.t73 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X15 pfd_8_0.DOWN.t0 pfd_8_0.DOWN_b.t3 GNDA.t49 GNDA.t48 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X16 GNDA.t134 GNDA.t131 GNDA.t133 GNDA.t132 sky130_fd_pr__nfet_01v8 ad=0.625 pd=3.5 as=0 ps=0 w=1.25 l=0.5
X17 a_n30_1400.t1 F_REF.t0 VDDA.t30 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X18 pfd_8_0.opamp_out.t3 a_6670_5090.t5 GNDA.t28 GNDA.t27 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X19 GNDA.t5 pfd_8_0.QA.t3 pfd_8_0.QA_b.t1 GNDA.t4 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X20 GNDA.t88 a_6400_6270.t10 a_6500_6300.t11 GNDA.t87 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X21 pfd_8_0.DOWN_input.t0 pfd_8_0.DOWN_b.t4 I_IN.t0 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X22 pfd_8_0.opamp_out.t8 opamp_cell_4_0.n_right.t6 VDDA.t81 VDDA.t80 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X23 a_1910_2020.t0 pfd_8_0.QB.t3 GNDA.t1 GNDA.t0 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X24 a_6500_6300.t5 a_6500_6300.t4 a_6500_6300.t5 GNDA.t141 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X25 pfd_8_0.UP.t1 pfd_8_0.UP_PFD_b.t2 VDDA.t20 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X26 pfd_8_0.UP_input.t1 pfd_8_0.UP.t2 pfd_8_0.opamp_out.t4 GNDA.t55 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X27 pfd_8_0.QA.t2 pfd_8_0.QA_b.t4 GNDA.t143 GNDA.t142 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X28 pfd_8_0.opamp_out.t10 a_9540_3974.t1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X29 pfd_8_0.DOWN_input.t2 pfd_8_0.DOWN.t3 I_IN.t1 GNDA.t58 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X30 a_1390_1400.t1 pfd_8_0.E.t3 pfd_8_0.E_b.t1 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X31 a_870_640.t0 pfd_8_0.QB_b.t3 VDDA.t127 VDDA.t123 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X32 VDDA.t113 VDDA.t111 VDDA.t113 VDDA.t112 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X33 VDDA.t29 a_2530_190.t2 a_2200_190.t1 VDDA.t28 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X34 GNDA.t130 GNDA.t127 GNDA.t129 GNDA.t128 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X35 pfd_8_0.DOWN_input.t1 pfd_8_0.DOWN_b.t5 GNDA.t147 GNDA.t146 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X36 GNDA.t149 a_2530_190.t3 a_2200_190.t0 GNDA.t148 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X37 pfd_8_0.F.t1 pfd_8_0.QB_b.t4 GNDA.t153 GNDA.t152 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X38 pfd_8_0.UP_b.t0 pfd_8_0.UP.t3 GNDA.t54 GNDA.t53 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X39 GNDA.t9 pfd_8_0.E_b.t3 pfd_8_0.E.t0 GNDA.t8 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X40 a_1390_640.t0 pfd_8_0.F.t3 pfd_8_0.F_b.t1 VDDA.t31 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X41 VDDA.t110 VDDA.t107 VDDA.t109 VDDA.t108 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X42 a_2350_1400.t1 pfd_8_0.before_Reset.t4 VDDA.t119 VDDA.t118 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X43 pfd_8_0.F_b.t2 pfd_8_0.F.t4 GNDA.t76 GNDA.t75 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X44 VDDA.t128 pfd_8_0.F.t5 a_490_640.t0 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X45 pfd_8_0.QA_b.t2 pfd_8_0.QA.t4 a_n30_1400.t0 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X46 GNDA.t126 GNDA.t124 GNDA.t126 GNDA.t125 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X47 opamp_cell_4_0.n_right.t2 opamp_cell_4_0.VIN+.t6 a_6500_6300.t1 GNDA.t42 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X48 VDDA.t106 VDDA.t104 VDDA.t106 VDDA.t105 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X49 GNDA.t136 pfd_8_0.F.t6 pfd_8_0.QB.t0 GNDA.t135 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X50 pfd_8_0.before_Reset.t0 pfd_8_0.QB.t4 VDDA.t6 VDDA.t5 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.805 ps=5 w=2 l=0.15
X51 GNDA.t123 GNDA.t121 GNDA.t123 GNDA.t122 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0 ps=0 w=1.25 l=0.5
X52 a_6150_5090.t4 a_6150_5090.t3 a_6150_5090.t4 VDDA.t35 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X53 opamp_cell_4_0.n_right.t3 opamp_cell_4_0.n_left.t7 VDDA.t73 VDDA.t72 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X54 pfd_8_0.UP_input.t2 pfd_8_0.UP_b.t3 pfd_8_0.opamp_out.t5 VDDA.t66 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X55 a_490_1400.t0 pfd_8_0.QA_b.t5 pfd_8_0.QA.t1 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X56 a_6380_5710.t3 a_6380_5710.t2 GNDA.t41 GNDA.t40 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X57 GNDA.t44 pfd_8_0.Reset.t2 pfd_8_0.E_b.t0 GNDA.t43 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X58 opamp_cell_4_0.p_bias.t5 opamp_cell_4_0.p_bias.t4 VDDA.t57 VDDA.t56 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X59 opamp_cell_4_0.VIN+.t3 pfd_8_0.opamp_out.t11 VDDA.t50 VDDA.t49 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X60 a_2530_190.t0 a_2350_1400.t2 GNDA.t57 GNDA.t56 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X61 a_6150_5090.t7 opamp_cell_4_0.p_bias.t10 VDDA.t4 VDDA.t3 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X62 VDDA.t103 VDDA.t101 VDDA.t103 VDDA.t102 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X63 a_6380_5710.t0 V_OUT.t9 a_6150_5090.t10 VDDA.t52 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X64 GNDA.t86 a_6400_6270.t5 a_6400_6270.t6 GNDA.t85 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X65 GNDA.t156 V_OUT.t7 sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X66 pfd_8_0.E.t1 pfd_8_0.E_b.t4 a_870_1400.t0 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X67 a_6500_6300.t3 V_OUT.t10 opamp_cell_4_0.n_left.t1 GNDA.t68 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X68 pfd_8_0.UP_b.t1 pfd_8_0.UP.t4 VDDA.t120 VDDA.t7 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X69 GNDA.t84 a_6400_6270.t7 a_6400_6270.t8 GNDA.t83 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X70 VDDA.t100 VDDA.t98 VDDA.t99 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=1.25 pd=6 as=0 ps=0 w=2.5 l=0.5
X71 VDDA.t14 a_1870_190.t2 pfd_8_0.Reset.t1 VDDA.t13 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X72 VDDA.t40 pfd_8_0.opamp_out.t12 opamp_cell_4_0.VIN+.t2 VDDA.t39 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X73 VDDA.t71 opamp_cell_4_0.n_left.t2 opamp_cell_4_0.n_left.t3 VDDA.t70 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X74 VDDA.t46 pfd_8_0.UP_input.t4 V_OUT.t3 VDDA.t45 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X75 GNDA.t82 a_6400_6270.t11 a_6500_6300.t10 GNDA.t81 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X76 VDDA.t59 opamp_cell_4_0.p_bias.t11 a_6150_5090.t6 VDDA.t58 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X77 V_OUT.t6 pfd_8_0.DOWN_input.t3 GNDA.t64 GNDA.t63 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X78 GNDA.t120 GNDA.t117 GNDA.t119 GNDA.t118 sky130_fd_pr__nfet_01v8 ad=0.25 pd=2 as=0 ps=0 w=0.5 l=0.15
X79 GNDA.t11 a_1870_190.t3 pfd_8_0.Reset.t0 GNDA.t10 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X80 pfd_8_0.opamp_out.t1 a_6670_5090.t6 GNDA.t16 GNDA.t15 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X81 opamp_cell_4_0.n_right.t0 a_9540_3974.t0 GNDA.t12 sky130_fd_pr__res_xhigh_po_0p35 l=1.14
X82 GNDA.t116 GNDA.t114 GNDA.t116 GNDA.t115 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X83 a_6150_5090.t2 a_6150_5090.t0 a_6150_5090.t1 VDDA.t36 sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0 ps=0 w=1 l=0.15
X84 a_6500_6300.t9 a_6400_6270.t12 GNDA.t80 GNDA.t79 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X85 opamp_cell_4_0.VIN+.t1 pfd_8_0.opamp_out.t13 VDDA.t1 VDDA.t0 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X86 pfd_8_0.before_Reset.t1 pfd_8_0.QA.t5 a_1910_2020.t1 GNDA.t38 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X87 pfd_8_0.opamp_out.t7 opamp_cell_4_0.n_right.t7 VDDA.t79 VDDA.t78 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X88 V_OUT.t0 loop_filter_2_0.R1_C1.t0 GNDA.t47 sky130_fd_pr__res_xhigh_po_0p35 l=7.52
X89 GNDA.t113 GNDA.t111 GNDA.t113 GNDA.t112 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X90 pfd_8_0.UP_PFD_b.t0 pfd_8_0.QA.t6 GNDA.t138 GNDA.t137 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X91 opamp_cell_4_0.p_bias.t8 a_6400_6270.t0 GNDA.t52 sky130_fd_pr__res_xhigh_po_5p73 l=1
X92 a_6400_6270.t4 a_6400_6270.t3 GNDA.t78 GNDA.t77 sky130_fd_pr__nfet_01v8 ad=0.3125 pd=1.75 as=0.3125 ps=1.75 w=1.25 l=0.5
X93 opamp_cell_4_0.n_left.t0 V_OUT.t11 a_6500_6300.t2 GNDA.t65 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X94 GNDA.t110 GNDA.t108 GNDA.t110 GNDA.t109 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0 ps=0 w=0.5 l=0.15
X95 GNDA.t46 pfd_8_0.E.t4 pfd_8_0.QA.t0 GNDA.t45 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X96 pfd_8_0.F.t2 pfd_8_0.F_b.t3 a_870_640.t1 VDDA.t25 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X97 VDDA.t24 pfd_8_0.Reset.t3 a_1390_1400.t0 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X98 GNDA.t107 GNDA.t105 GNDA.t107 GNDA.t106 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0 ps=0 w=2 l=0.6
X99 GNDA.t104 GNDA.t101 GNDA.t103 GNDA.t102 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X100 pfd_8_0.UP_input.t5 pfd_8_0.UP_b.t2 sky130_fd_pr__cap_mim_m3_1 l=6.3 w=7
X101 a_2530_190.t1 a_2350_1400.t3 VDDA.t10 VDDA.t9 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X102 VDDA.t97 VDDA.t95 VDDA.t97 VDDA.t96 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0 ps=0 w=1 l=0.15
X103 a_9540_6900.t0 a_6670_5090.t0 GNDA.t24 sky130_fd_pr__res_xhigh_po_0p35 l=0.86
X104 opamp_cell_4_0.n_left.t5 opamp_cell_4_0.n_left.t4 VDDA.t69 VDDA.t68 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X105 GNDA.t100 GNDA.t97 GNDA.t99 GNDA.t98 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X106 GNDA.t23 pfd_8_0.F_b.t4 pfd_8_0.F.t0 GNDA.t22 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X107 GNDA.t62 pfd_8_0.DOWN_input.t4 V_OUT.t5 GNDA.t61 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X108 pfd_8_0.QB_b.t0 pfd_8_0.QB.t5 a_n30_640.t1 VDDA.t2 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X109 VDDA.t34 pfd_8_0.opamp_out.t14 opamp_cell_4_0.VIN+.t0 VDDA.t33 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X110 VDDA.t94 VDDA.t91 VDDA.t93 VDDA.t92 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X111 pfd_8_0.opamp_out.t15 a_9540_6900.t1 sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X112 VDDA.t121 pfd_8_0.Reset.t4 a_1390_640.t1 VDDA.t23 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X113 GNDA.t18 I_IN.t6 opamp_cell_4_0.VIN+.t5 GNDA.t17 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X114 pfd_8_0.UP_input.t0 pfd_8_0.UP.t5 VDDA.t27 VDDA.t26 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X115 GNDA.t140 a_6380_5710.t6 a_6670_5090.t4 GNDA.t139 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X116 GNDA.t70 pfd_8_0.QB.t6 pfd_8_0.QB_b.t1 GNDA.t69 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X117 GNDA.t20 I_IN.t4 I_IN.t5 GNDA.t19 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X118 GNDA.t35 pfd_8_0.Reset.t5 pfd_8_0.F_b.t0 GNDA.t34 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.2 ps=1.4 w=1 l=0.15
X119 GNDA.t14 a_6670_5090.t7 pfd_8_0.opamp_out.t0 GNDA.t13 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X120 a_6150_5090.t12 opamp_cell_4_0.VIN+.t7 a_6670_5090.t2 VDDA.t67 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X121 VDDA.t90 VDDA.t87 VDDA.t89 VDDA.t88 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X122 pfd_8_0.E.t2 pfd_8_0.QA_b.t6 GNDA.t33 GNDA.t32 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X123 VDDA.t77 opamp_cell_4_0.n_right.t8 pfd_8_0.opamp_out.t6 VDDA.t76 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X124 VDDA.t86 VDDA.t84 VDDA.t86 VDDA.t85 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0 ps=0 w=2.5 l=0.5
X125 VDDA.t22 pfd_8_0.QA.t7 pfd_8_0.before_Reset.t2 VDDA.t21 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X126 opamp_cell_4_0.VIN+.t4 I_IN.t7 GNDA.t7 GNDA.t6 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X127 a_n30_640.t0 F_VCO.t0 VDDA.t16 VDDA.t15 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X128 pfd_8_0.UP_PFD_b.t1 pfd_8_0.QA.t8 VDDA.t18 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X129 VDDA.t126 pfd_8_0.E.t5 a_490_1400.t1 VDDA.t125 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.4 ps=2.4 w=2 l=0.15
X130 I_IN.t3 I_IN.t2 GNDA.t67 GNDA.t66 sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X131 VDDA.t12 a_2200_190.t2 a_1870_190.t1 VDDA.t11 sky130_fd_pr__pfet_01v8 ad=0.8 pd=4.8 as=0.8 ps=4.8 w=2 l=0.15
X132 V_OUT.t2 pfd_8_0.UP_input.t6 VDDA.t44 VDDA.t43 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X133 pfd_8_0.QA_b.t0 F_REF.t1 GNDA.t3 GNDA.t2 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X134 a_6670_5090.t3 a_6380_5710.t7 GNDA.t145 GNDA.t144 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X135 pfd_8_0.QB_b.t2 F_VCO.t1 GNDA.t51 GNDA.t50 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X136 a_490_640.t1 pfd_8_0.QB_b.t5 pfd_8_0.QB.t1 VDDA.t122 sky130_fd_pr__pfet_01v8 ad=0.4 pd=2.4 as=0.8 ps=4.8 w=2 l=0.15
X137 GNDA.t157 loop_filter_2_0.R1_C1.t1 sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X138 GNDA.t37 a_2200_190.t3 a_1870_190.t0 GNDA.t36 sky130_fd_pr__nfet_01v8 ad=0.4 pd=2.8 as=0.4 ps=2.8 w=1 l=0.15
X139 VDDA.t61 opamp_cell_4_0.p_bias.t2 opamp_cell_4_0.p_bias.t3 VDDA.t60 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X140 pfd_8_0.DOWN_input.t5 pfd_8_0.DOWN.t2 sky130_fd_pr__cap_mim_m3_1 l=2.6 w=3.8
X141 pfd_8_0.QB.t2 pfd_8_0.QB_b.t6 GNDA.t155 GNDA.t154 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X142 pfd_8_0.DOWN_PFD_b.t1 pfd_8_0.QB.t7 VDDA.t51 VDDA.t17 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
X143 a_6670_5090.t1 opamp_cell_4_0.VIN+.t8 a_6150_5090.t9 VDDA.t32 sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X144 pfd_8_0.UP.t0 pfd_8_0.UP_PFD_b.t3 GNDA.t72 GNDA.t71 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X145 VDDA.t38 opamp_cell_4_0.p_bias.t0 opamp_cell_4_0.p_bias.t1 VDDA.t37 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X146 a_6500_6300.t0 opamp_cell_4_0.VIN+.t9 opamp_cell_4_0.n_right.t1 GNDA.t21 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X147 GNDA.t26 a_6670_5090.t8 pfd_8_0.opamp_out.t2 GNDA.t25 sky130_fd_pr__nfet_01v8 ad=0.125 pd=1 as=0.125 ps=1 w=0.5 l=0.15
X148 pfd_8_0.DOWN_PFD_b.t0 pfd_8_0.QB.t8 GNDA.t60 GNDA.t59 sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X149 VDDA.t42 pfd_8_0.UP_input.t7 V_OUT.t1 VDDA.t41 sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.5 ps=2.5 w=2 l=0.6
X150 pfd_8_0.E_b.t2 pfd_8_0.E.t6 GNDA.t151 GNDA.t150 sky130_fd_pr__nfet_01v8 ad=0.2 pd=1.4 as=0.4 ps=2.8 w=1 l=0.15
X151 VDDA.t65 opamp_cell_4_0.p_bias.t12 a_6150_5090.t5 VDDA.t64 sky130_fd_pr__pfet_01v8 ad=0.625 pd=3 as=0.625 ps=3 w=2.5 l=0.5
X152 GNDA.t96 GNDA.t93 GNDA.t95 GNDA.t94 sky130_fd_pr__nfet_01v8 ad=1 pd=5 as=0 ps=0 w=2 l=0.6
X153 pfd_8_0.DOWN_b.t0 GNDA.t158 pfd_8_0.DOWN_PFD_b.t2 VDDA.t19 sky130_fd_pr__pfet_01v8 ad=1 pd=5 as=1 ps=5 w=2 l=0.15
R0 a_6400_6270.n4 a_6400_6270.t12 317.317
R1 a_6400_6270.n2 a_6400_6270.t11 317.317
R2 a_6400_6270.n5 a_6400_6270.n4 257.067
R3 a_6400_6270.n3 a_6400_6270.n2 257.067
R4 a_6400_6270.n10 a_6400_6270.n9 257.067
R5 a_6400_6270.t0 a_6400_6270.n12 194.478
R6 a_6400_6270.n8 a_6400_6270.n7 152
R7 a_6400_6270.n12 a_6400_6270.n11 152
R8 a_6400_6270.n1 a_6400_6270.n0 120.981
R9 a_6400_6270.n7 a_6400_6270.n6 117.781
R10 a_6400_6270.n7 a_6400_6270.n1 108.8
R11 a_6400_6270.n8 a_6400_6270.n5 85.6894
R12 a_6400_6270.n11 a_6400_6270.n3 85.6894
R13 a_6400_6270.n11 a_6400_6270.n10 85.6894
R14 a_6400_6270.n9 a_6400_6270.n8 85.6894
R15 a_6400_6270.n4 a_6400_6270.t10 60.2505
R16 a_6400_6270.n5 a_6400_6270.t3 60.2505
R17 a_6400_6270.n2 a_6400_6270.t9 60.2505
R18 a_6400_6270.n3 a_6400_6270.t7 60.2505
R19 a_6400_6270.n10 a_6400_6270.t1 60.2505
R20 a_6400_6270.n9 a_6400_6270.t5 60.2505
R21 a_6400_6270.n6 a_6400_6270.t6 24.0005
R22 a_6400_6270.n6 a_6400_6270.t4 24.0005
R23 a_6400_6270.n0 a_6400_6270.t8 24.0005
R24 a_6400_6270.n0 a_6400_6270.t2 24.0005
R25 a_6400_6270.n12 a_6400_6270.n1 3.2005
R26 GNDA.n246 GNDA.n77 35793.3
R27 GNDA.n396 GNDA.n395 18430.6
R28 GNDA.t55 GNDA.n311 1397.16
R29 GNDA.n261 GNDA.n260 1186
R30 GNDA.n58 GNDA.n50 1186
R31 GNDA.n256 GNDA.n255 1186
R32 GNDA.n251 GNDA.n250 1186
R33 GNDA.n246 GNDA.n245 1170
R34 GNDA.t12 GNDA.t47 1026.12
R35 GNDA.n173 GNDA.n172 669.307
R36 GNDA.n175 GNDA.n94 669.307
R37 GNDA.n168 GNDA.n167 669.307
R38 GNDA.n165 GNDA.n98 669.307
R39 GNDA.n119 GNDA.n118 669.307
R40 GNDA.n123 GNDA.n122 669.307
R41 GNDA.n360 GNDA.n359 585.003
R42 GNDA.n398 GNDA.n397 585.003
R43 GNDA.n395 GNDA.n394 585.001
R44 GNDA.n362 GNDA.n361 585.001
R45 GNDA.n357 GNDA.n356 585.001
R46 GNDA.n313 GNDA.n312 585.001
R47 GNDA.n315 GNDA.n314 585.001
R48 GNDA.n206 GNDA.n205 585.001
R49 GNDA.n208 GNDA.n207 585.001
R50 GNDA.n214 GNDA.n23 585.001
R51 GNDA.n403 GNDA.n402 585.001
R52 GNDA.n401 GNDA.n19 585.001
R53 GNDA.n400 GNDA.n16 585.001
R54 GNDA.n399 GNDA.n13 585.001
R55 GNDA.n396 GNDA.n2 585.001
R56 GNDA.n319 GNDA.n318 585.001
R57 GNDA.n317 GNDA.n47 585.001
R58 GNDA.n316 GNDA.n44 585.001
R59 GNDA.n259 GNDA.n258 585.001
R60 GNDA.n311 GNDA.n310 585.001
R61 GNDA.n120 GNDA.n117 585
R62 GNDA.n121 GNDA.n114 585
R63 GNDA.n102 GNDA.n99 585
R64 GNDA.n105 GNDA.n104 585
R65 GNDA.n97 GNDA.n96 585
R66 GNDA.n177 GNDA.n176 585
R67 GNDA.n203 GNDA.n202 585
R68 GNDA.n204 GNDA.n203 585
R69 GNDA.n201 GNDA.n86 585
R70 GNDA.n199 GNDA.n198 585
R71 GNDA.n197 GNDA.n85 585
R72 GNDA.n204 GNDA.n85 585
R73 GNDA.n212 GNDA.t158 566.966
R74 GNDA.n247 GNDA.t12 491.574
R75 GNDA.t146 GNDA.n204 450.389
R76 GNDA.n170 GNDA.t105 336.329
R77 GNDA.n170 GNDA.t97 336.329
R78 GNDA.n100 GNDA.t111 336.329
R79 GNDA.n100 GNDA.t101 336.329
R80 GNDA.n259 GNDA.t141 333.075
R81 GNDA.n196 GNDA.t93 320.7
R82 GNDA.n124 GNDA.t114 320.7
R83 GNDA.n248 GNDA.t108 304.634
R84 GNDA.n262 GNDA.t127 304.634
R85 GNDA.n59 GNDA.t117 304.634
R86 GNDA.n254 GNDA.t124 304.634
R87 GNDA.t150 GNDA.t8 296.906
R88 GNDA.t142 GNDA.t4 296.906
R89 GNDA.n257 GNDA.t121 292.584
R90 GNDA.n309 GNDA.t131 292.584
R91 GNDA.t91 GNDA.n256 290.373
R92 GNDA.t109 GNDA.n251 281.832
R93 GNDA.n260 GNDA.t128 281.832
R94 GNDA.t29 GNDA.t91 264.752
R95 GNDA.t132 GNDA.n50 256.212
R96 GNDA.n119 GNDA.n77 250.349
R97 GNDA.n122 GNDA.n77 250.349
R98 GNDA.n169 GNDA.n168 250.349
R99 GNDA.n169 GNDA.n98 250.349
R100 GNDA.n174 GNDA.n173 250.349
R101 GNDA.n175 GNDA.n174 250.349
R102 GNDA.n204 GNDA.n84 250.349
R103 GNDA.n250 GNDA.t110 245
R104 GNDA.n261 GNDA.t130 245
R105 GNDA.n58 GNDA.t120 245
R106 GNDA.n255 GNDA.t126 245
R107 GNDA.t85 GNDA.t125 230.59
R108 GNDA.t13 GNDA.t109 222.05
R109 GNDA.t15 GNDA.t13 222.05
R110 GNDA.t25 GNDA.t15 222.05
R111 GNDA.t27 GNDA.t25 222.05
R112 GNDA.t128 GNDA.t27 222.05
R113 GNDA.n260 GNDA.n259 222.05
R114 GNDA.t42 GNDA.t68 222.05
R115 GNDA.t139 GNDA.t144 222.05
R116 GNDA.t40 GNDA.t118 222.05
R117 GNDA.t122 GNDA.t21 213.51
R118 GNDA.t87 GNDA.t30 213.51
R119 GNDA.t53 GNDA.t55 210.007
R120 GNDA.n316 GNDA.t56 206.387
R121 GNDA.n264 GNDA.n74 204.201
R122 GNDA.n61 GNDA.n56 204.201
R123 GNDA.n60 GNDA.n57 204.201
R124 GNDA.n253 GNDA.n252 204.201
R125 GNDA.n263 GNDA.n76 204.201
R126 GNDA.n249 GNDA.n75 204.201
R127 GNDA.n3 GNDA.t70 198.058
R128 GNDA.n444 GNDA.t155 198.058
R129 GNDA.n432 GNDA.t23 198.058
R130 GNDA.n11 GNDA.t76 198.058
R131 GNDA.n388 GNDA.t5 198.058
R132 GNDA.n26 GNDA.t143 198.058
R133 GNDA.n374 GNDA.t9 198.058
R134 GNDA.n369 GNDA.t151 198.058
R135 GNDA.n176 GNDA.n97 197
R136 GNDA.n104 GNDA.n99 197
R137 GNDA.n121 GNDA.n120 197
R138 GNDA.n203 GNDA.n86 197
R139 GNDA.n198 GNDA.n85 197
R140 GNDA.t89 GNDA.t65 196.429
R141 GNDA.n172 GNDA.n171 185
R142 GNDA.n171 GNDA.n94 185
R143 GNDA.n167 GNDA.n166 185
R144 GNDA.n166 GNDA.n165 185
R145 GNDA.n118 GNDA.n115 185
R146 GNDA.n123 GNDA.n115 185
R147 GNDA.n202 GNDA.n87 185
R148 GNDA.n197 GNDA.n87 185
R149 GNDA.n318 GNDA.t71 170.179
R150 GNDA.n317 GNDA.t137 170.179
R151 GNDA.n172 GNDA.n170 166.63
R152 GNDA.n167 GNDA.n100 166.63
R153 GNDA.n251 GNDA.n247 153.727
R154 GNDA.t65 GNDA.t83 145.186
R155 GNDA.n315 GNDA.t73 141.212
R156 GNDA.n313 GNDA.t38 141.212
R157 GNDA.t75 GNDA.t22 137.921
R158 GNDA.t154 GNDA.t69 137.921
R159 GNDA.n258 GNDA.t123 134.501
R160 GNDA.n310 GNDA.t134 134.501
R161 GNDA.t39 GNDA.t59 131.194
R162 GNDA.n7 GNDA.t136 130.713
R163 GNDA.n394 GNDA.t3 130.001
R164 GNDA.n362 GNDA.t44 130.001
R165 GNDA.n356 GNDA.t1 130.001
R166 GNDA.n312 GNDA.t74 130.001
R167 GNDA.n314 GNDA.t57 130.001
R168 GNDA.n2 GNDA.t51 130.001
R169 GNDA.n13 GNDA.t35 130.001
R170 GNDA.n16 GNDA.t11 130.001
R171 GNDA.n19 GNDA.t37 130.001
R172 GNDA.n403 GNDA.t149 130.001
R173 GNDA.n358 GNDA.t33 130.001
R174 GNDA.n28 GNDA.t46 130.001
R175 GNDA.n8 GNDA.t153 130.001
R176 GNDA.t21 GNDA.t81 128.107
R177 GNDA.t30 GNDA.t79 128.107
R178 GNDA.n44 GNDA.t138 122.501
R179 GNDA.n47 GNDA.t72 122.501
R180 GNDA.n319 GNDA.t54 122.501
R181 GNDA.n214 GNDA.t60 122.501
R182 GNDA.n208 GNDA.t49 122.501
R183 GNDA.n205 GNDA.t147 122.501
R184 GNDA.n318 GNDA.t53 112.246
R185 GNDA.t71 GNDA.n317 112.246
R186 GNDA.t137 GNDA.n316 112.246
R187 GNDA.t125 GNDA.t77 111.025
R188 GNDA.t77 GNDA.t139 111.025
R189 GNDA.n361 GNDA.n357 101.382
R190 GNDA.n269 GNDA.n72 97.8707
R191 GNDA.n276 GNDA.n69 97.8707
R192 GNDA.n283 GNDA.n66 97.8707
R193 GNDA.n290 GNDA.n63 97.8707
R194 GNDA.n298 GNDA.n54 97.8707
R195 GNDA.t56 GNDA.n315 97.7622
R196 GNDA.t73 GNDA.n313 97.7622
R197 GNDA.n357 GNDA.t0 97.7622
R198 GNDA.n361 GNDA.t43 97.7622
R199 GNDA.t32 GNDA.n360 97.7622
R200 GNDA.n360 GNDA.t45 97.7622
R201 GNDA.n395 GNDA.t2 97.7622
R202 GNDA.t48 GNDA.t58 97.554
R203 GNDA.t81 GNDA.t42 93.9446
R204 GNDA.n133 GNDA.n110 92.2612
R205 GNDA.n126 GNDA.n113 92.2612
R206 GNDA.n159 GNDA.n139 92.2612
R207 GNDA.n153 GNDA.n142 92.2612
R208 GNDA.n181 GNDA.n180 92.2612
R209 GNDA.n188 GNDA.n187 92.2612
R210 GNDA.n171 GNDA.n95 91.3721
R211 GNDA.n179 GNDA.n93 91.3721
R212 GNDA.n179 GNDA.n178 91.3721
R213 GNDA.n166 GNDA.n103 91.3721
R214 GNDA.n138 GNDA.n101 91.3721
R215 GNDA.n138 GNDA.n106 91.3721
R216 GNDA.n116 GNDA.n115 90.7567
R217 GNDA.n200 GNDA.n87 90.7567
R218 GNDA.t10 GNDA.n399 89.1442
R219 GNDA.n402 GNDA.n23 87.4623
R220 GNDA.n311 GNDA.n50 85.4042
R221 GNDA.n120 GNDA.n119 84.306
R222 GNDA.n122 GNDA.n121 84.306
R223 GNDA.n168 GNDA.n99 84.306
R224 GNDA.n104 GNDA.n98 84.306
R225 GNDA.n173 GNDA.n97 84.306
R226 GNDA.n176 GNDA.n175 84.306
R227 GNDA.n86 GNDA.n84 84.306
R228 GNDA.n198 GNDA.n84 84.306
R229 GNDA.n253 GNDA.n61 83.2005
R230 GNDA.n61 GNDA.n60 83.2005
R231 GNDA.n78 GNDA.t156 79.6829
R232 GNDA.t38 GNDA.t0 79.6582
R233 GNDA.t43 GNDA.t150 79.6582
R234 GNDA.t8 GNDA.t32 79.6582
R235 GNDA.t45 GNDA.t142 79.6582
R236 GNDA.t4 GNDA.t2 79.6582
R237 GNDA.t83 GNDA.t29 76.8638
R238 GNDA.n78 GNDA.t157 76.4829
R239 GNDA.t58 GNDA.n206 75.6886
R240 GNDA.n207 GNDA.t39 75.6886
R241 GNDA.t61 GNDA.t115 70.6574
R242 GNDA.t63 GNDA.t61 70.6574
R243 GNDA.t102 GNDA.t63 70.6574
R244 GNDA.t17 GNDA.t112 70.6574
R245 GNDA.t6 GNDA.t17 70.6574
R246 GNDA.t98 GNDA.t6 70.6574
R247 GNDA.t106 GNDA.t19 70.6574
R248 GNDA.t19 GNDA.t66 70.6574
R249 GNDA.t66 GNDA.t94 70.6574
R250 GNDA.t115 GNDA.n77 67.4458
R251 GNDA.n169 GNDA.t102 67.4458
R252 GNDA.t112 GNDA.n169 67.4458
R253 GNDA.n174 GNDA.t98 67.4458
R254 GNDA.n174 GNDA.t106 67.4458
R255 GNDA.n204 GNDA.t94 67.4458
R256 GNDA.n264 GNDA.n75 66.5605
R257 GNDA.n264 GNDA.n263 66.5605
R258 GNDA.n265 GNDA.n264 65.9634
R259 GNDA.t148 GNDA.n401 65.5968
R260 GNDA.t36 GNDA.n400 65.5968
R261 GNDA.n394 GNDA.n393 60.29
R262 GNDA.n363 GNDA.n362 60.29
R263 GNDA.n356 GNDA.n355 60.29
R264 GNDA.n312 GNDA.n38 60.29
R265 GNDA.n314 GNDA.n40 60.29
R266 GNDA.n404 GNDA.n403 60.29
R267 GNDA.n411 GNDA.n19 60.29
R268 GNDA.n417 GNDA.n16 60.29
R269 GNDA.n424 GNDA.n13 60.29
R270 GNDA.n452 GNDA.n2 60.29
R271 GNDA.n74 GNDA.t16 60.0005
R272 GNDA.n74 GNDA.t26 60.0005
R273 GNDA.n56 GNDA.t145 60.0005
R274 GNDA.n56 GNDA.t31 60.0005
R275 GNDA.n57 GNDA.t41 60.0005
R276 GNDA.n57 GNDA.t119 60.0005
R277 GNDA.n252 GNDA.t126 60.0005
R278 GNDA.n252 GNDA.t140 60.0005
R279 GNDA.n76 GNDA.t28 60.0005
R280 GNDA.n76 GNDA.t129 60.0005
R281 GNDA.t110 GNDA.n249 60.0005
R282 GNDA.n249 GNDA.t14 60.0005
R283 GNDA.n333 GNDA.n44 59.5478
R284 GNDA.n326 GNDA.n47 59.5478
R285 GNDA.n320 GNDA.n319 59.5478
R286 GNDA.t47 GNDA.n246 59.2402
R287 GNDA.n233 GNDA.n208 58.9809
R288 GNDA.n221 GNDA.n214 58.9809
R289 GNDA.n205 GNDA.n80 58.9809
R290 GNDA.n206 GNDA.t146 55.5051
R291 GNDA.n207 GNDA.t48 55.5051
R292 GNDA.t59 GNDA.n23 55.5051
R293 GNDA.n380 GNDA.n28 54.4005
R294 GNDA.n358 GNDA.n29 54.4005
R295 GNDA.n437 GNDA.n8 54.4005
R296 GNDA.n439 GNDA.n7 54.4005
R297 GNDA.t52 GNDA.t40 52.9508
R298 GNDA.n256 GNDA.t85 51.2427
R299 GNDA.n247 GNDA.t24 46.9276
R300 GNDA.n402 GNDA.t148 45.4133
R301 GNDA.n401 GNDA.t36 45.4133
R302 GNDA.n400 GNDA.t10 45.4133
R303 GNDA.n399 GNDA.t34 45.4133
R304 GNDA.t152 GNDA.n398 45.4133
R305 GNDA.n398 GNDA.t135 45.4133
R306 GNDA.t50 GNDA.n396 45.4133
R307 GNDA GNDA.n244 41.8937
R308 GNDA.n294 GNDA.n61 41.6005
R309 GNDA.n194 GNDA.n192 41.3005
R310 GNDA.t79 GNDA.t52 40.9943
R311 GNDA.n266 GNDA.n265 39.4985
R312 GNDA.t34 GNDA.t75 37.0036
R313 GNDA.t22 GNDA.t152 37.0036
R314 GNDA.t135 GNDA.t154 37.0036
R315 GNDA.t69 GNDA.t50 37.0036
R316 GNDA.n393 GNDA.n0 33.0991
R317 GNDA.n453 GNDA.n452 33.0991
R318 GNDA.n134 GNDA.n133 32.0005
R319 GNDA.n134 GNDA.n107 32.0005
R320 GNDA.n128 GNDA.n127 32.0005
R321 GNDA.n128 GNDA.n111 32.0005
R322 GNDA.n132 GNDA.n111 32.0005
R323 GNDA.n160 GNDA.n108 32.0005
R324 GNDA.n158 GNDA.n140 32.0005
R325 GNDA.n154 GNDA.n140 32.0005
R326 GNDA.n154 GNDA.n153 32.0005
R327 GNDA.n152 GNDA.n143 32.0005
R328 GNDA.n148 GNDA.n143 32.0005
R329 GNDA.n147 GNDA.n146 32.0005
R330 GNDA.n146 GNDA.n92 32.0005
R331 GNDA.n185 GNDA.n90 32.0005
R332 GNDA.n186 GNDA.n185 32.0005
R333 GNDA.n195 GNDA.n88 32.0005
R334 GNDA.n266 GNDA.n71 32.0005
R335 GNDA.n271 GNDA.n71 32.0005
R336 GNDA.n272 GNDA.n271 32.0005
R337 GNDA.n273 GNDA.n272 32.0005
R338 GNDA.n273 GNDA.n68 32.0005
R339 GNDA.n278 GNDA.n68 32.0005
R340 GNDA.n279 GNDA.n278 32.0005
R341 GNDA.n280 GNDA.n279 32.0005
R342 GNDA.n280 GNDA.n65 32.0005
R343 GNDA.n285 GNDA.n65 32.0005
R344 GNDA.n286 GNDA.n285 32.0005
R345 GNDA.n287 GNDA.n286 32.0005
R346 GNDA.n287 GNDA.n62 32.0005
R347 GNDA.n292 GNDA.n62 32.0005
R348 GNDA.n293 GNDA.n292 32.0005
R349 GNDA.n295 GNDA.n53 32.0005
R350 GNDA.n300 GNDA.n53 32.0005
R351 GNDA.n301 GNDA.n300 32.0005
R352 GNDA.n306 GNDA.n301 32.0005
R353 GNDA.n306 GNDA.n305 32.0005
R354 GNDA.n305 GNDA.n304 32.0005
R355 GNDA.n320 GNDA.n48 32.0005
R356 GNDA.n324 GNDA.n48 32.0005
R357 GNDA.n325 GNDA.n324 32.0005
R358 GNDA.n327 GNDA.n45 32.0005
R359 GNDA.n331 GNDA.n45 32.0005
R360 GNDA.n332 GNDA.n331 32.0005
R361 GNDA.n334 GNDA.n42 32.0005
R362 GNDA.n338 GNDA.n42 32.0005
R363 GNDA.n339 GNDA.n338 32.0005
R364 GNDA.n340 GNDA.n339 32.0005
R365 GNDA.n344 GNDA.n343 32.0005
R366 GNDA.n345 GNDA.n344 32.0005
R367 GNDA.n349 GNDA.n348 32.0005
R368 GNDA.n350 GNDA.n349 32.0005
R369 GNDA.n350 GNDA.n36 32.0005
R370 GNDA.n354 GNDA.n35 32.0005
R371 GNDA.n364 GNDA.n35 32.0005
R372 GNDA.n368 GNDA.n33 32.0005
R373 GNDA.n369 GNDA.n368 32.0005
R374 GNDA.n370 GNDA.n369 32.0005
R375 GNDA.n370 GNDA.n31 32.0005
R376 GNDA.n374 GNDA.n31 32.0005
R377 GNDA.n375 GNDA.n374 32.0005
R378 GNDA.n376 GNDA.n375 32.0005
R379 GNDA.n382 GNDA.n381 32.0005
R380 GNDA.n382 GNDA.n26 32.0005
R381 GNDA.n386 GNDA.n26 32.0005
R382 GNDA.n387 GNDA.n386 32.0005
R383 GNDA.n388 GNDA.n387 32.0005
R384 GNDA.n388 GNDA.n24 32.0005
R385 GNDA.n392 GNDA.n24 32.0005
R386 GNDA.n241 GNDA.n240 32.0005
R387 GNDA.n240 GNDA.n239 32.0005
R388 GNDA.n239 GNDA.n82 32.0005
R389 GNDA.n235 GNDA.n82 32.0005
R390 GNDA.n235 GNDA.n234 32.0005
R391 GNDA.n234 GNDA.n233 32.0005
R392 GNDA.n233 GNDA.n209 32.0005
R393 GNDA.n229 GNDA.n209 32.0005
R394 GNDA.n229 GNDA.n228 32.0005
R395 GNDA.n228 GNDA.n227 32.0005
R396 GNDA.n227 GNDA.n211 32.0005
R397 GNDA.n223 GNDA.n211 32.0005
R398 GNDA.n223 GNDA.n222 32.0005
R399 GNDA.n220 GNDA.n215 32.0005
R400 GNDA.n216 GNDA.n215 32.0005
R401 GNDA.n216 GNDA.n22 32.0005
R402 GNDA.n405 GNDA.n22 32.0005
R403 GNDA.n409 GNDA.n20 32.0005
R404 GNDA.n410 GNDA.n409 32.0005
R405 GNDA.n412 GNDA.n17 32.0005
R406 GNDA.n416 GNDA.n17 32.0005
R407 GNDA.n419 GNDA.n418 32.0005
R408 GNDA.n419 GNDA.n14 32.0005
R409 GNDA.n423 GNDA.n14 32.0005
R410 GNDA.n426 GNDA.n425 32.0005
R411 GNDA.n426 GNDA.n11 32.0005
R412 GNDA.n430 GNDA.n11 32.0005
R413 GNDA.n431 GNDA.n430 32.0005
R414 GNDA.n432 GNDA.n431 32.0005
R415 GNDA.n432 GNDA.n9 32.0005
R416 GNDA.n436 GNDA.n9 32.0005
R417 GNDA.n440 GNDA.n5 32.0005
R418 GNDA.n444 GNDA.n5 32.0005
R419 GNDA.n445 GNDA.n444 32.0005
R420 GNDA.n446 GNDA.n445 32.0005
R421 GNDA.n446 GNDA.n3 32.0005
R422 GNDA.n450 GNDA.n3 32.0005
R423 GNDA.n451 GNDA.n450 32.0005
R424 GNDA.n147 GNDA.n94 29.0291
R425 GNDA.n165 GNDA.n164 29.0291
R426 GNDA.n326 GNDA.n325 28.8005
R427 GNDA.n343 GNDA.n40 28.8005
R428 GNDA.n262 GNDA.n261 27.2005
R429 GNDA.n250 GNDA.n248 27.2005
R430 GNDA.t68 GNDA.t89 25.6216
R431 GNDA.t118 GNDA.t132 25.6216
R432 GNDA.n164 GNDA.n108 25.6005
R433 GNDA.n181 GNDA.n90 25.6005
R434 GNDA.n188 GNDA.n186 25.6005
R435 GNDA.n59 GNDA.n58 25.6005
R436 GNDA.n255 GNDA.n254 25.6005
R437 GNDA.n295 GNDA.n294 25.6005
R438 GNDA.n304 GNDA 25.6005
R439 GNDA.n333 GNDA.n332 25.6005
R440 GNDA.n355 GNDA.n36 25.6005
R441 GNDA.n364 GNDA.n363 25.6005
R442 GNDA.n379 GNDA.n29 25.6005
R443 GNDA.n380 GNDA.n379 25.6005
R444 GNDA.n241 GNDA.n80 25.6005
R445 GNDA.n222 GNDA.n221 25.6005
R446 GNDA.n404 GNDA.n20 25.6005
R447 GNDA.n417 GNDA.n416 25.6005
R448 GNDA.n424 GNDA.n423 25.6005
R449 GNDA.n438 GNDA.n437 25.6005
R450 GNDA.n258 GNDA.n257 24.8279
R451 GNDA.n310 GNDA.n309 24.8279
R452 GNDA.t123 GNDA.n72 24.0005
R453 GNDA.n72 GNDA.t82 24.0005
R454 GNDA.n69 GNDA.t90 24.0005
R455 GNDA.n69 GNDA.t84 24.0005
R456 GNDA.n66 GNDA.t92 24.0005
R457 GNDA.n66 GNDA.t86 24.0005
R458 GNDA.n63 GNDA.t78 24.0005
R459 GNDA.n63 GNDA.t88 24.0005
R460 GNDA.n54 GNDA.t80 24.0005
R461 GNDA.n54 GNDA.t133 24.0005
R462 GNDA.n439 GNDA.n438 22.4005
R463 GNDA.n125 GNDA.n124 20.9665
R464 GNDA.n160 GNDA.n159 19.2005
R465 GNDA.n159 GNDA.n158 19.2005
R466 GNDA.n348 GNDA.n38 19.2005
R467 GNDA.n411 GNDA.n410 16.0005
R468 GNDA.n412 GNDA.n411 16.0005
R469 GNDA.n302 GNDA 15.7005
R470 GNDA.n124 GNDA.n123 15.6449
R471 GNDA.n197 GNDA.n196 15.6449
R472 GNDA.n110 GNDA.t64 15.0005
R473 GNDA.n110 GNDA.t103 15.0005
R474 GNDA.t116 GNDA.n113 15.0005
R475 GNDA.n113 GNDA.t62 15.0005
R476 GNDA.n139 GNDA.t113 15.0005
R477 GNDA.n139 GNDA.t18 15.0005
R478 GNDA.n142 GNDA.t7 15.0005
R479 GNDA.n142 GNDA.t99 15.0005
R480 GNDA.n180 GNDA.t107 15.0005
R481 GNDA.n180 GNDA.t20 15.0005
R482 GNDA.n187 GNDA.t67 15.0005
R483 GNDA.n187 GNDA.t95 15.0005
R484 GNDA.t107 GNDA.n179 15.0005
R485 GNDA.n171 GNDA.t100 15.0005
R486 GNDA.t113 GNDA.n138 15.0005
R487 GNDA.n166 GNDA.t104 15.0005
R488 GNDA.n115 GNDA.t116 15.0005
R489 GNDA.n87 GNDA.t96 15.0005
R490 GNDA.n196 GNDA.n195 14.4005
R491 GNDA.n263 GNDA.n262 14.0805
R492 GNDA.n248 GNDA.n75 14.0805
R493 GNDA.n243 GNDA.n80 13.9181
R494 GNDA.n302 GNDA.n49 13.506
R495 GNDA.n321 GNDA.n49 12.8163
R496 GNDA.n164 GNDA.n107 12.8005
R497 GNDA.n127 GNDA.n126 12.8005
R498 GNDA.n181 GNDA.n92 12.8005
R499 GNDA.n188 GNDA.n88 12.8005
R500 GNDA.n60 GNDA.n59 12.8005
R501 GNDA.n254 GNDA.n253 12.8005
R502 GNDA.n345 GNDA.n38 12.8005
R503 GNDA GNDA.n0 12.7806
R504 GNDA GNDA.n453 11.8829
R505 GNDA.n192 GNDA.n79 11.8187
R506 GNDA.n244 GNDA.n243 11.7212
R507 GNDA.n440 GNDA.n439 9.6005
R508 GNDA.n257 GNDA.n73 9.58175
R509 GNDA.n309 GNDA.n308 9.58175
R510 GNDA.n267 GNDA.n266 9.3005
R511 GNDA.n268 GNDA.n71 9.3005
R512 GNDA.n271 GNDA.n270 9.3005
R513 GNDA.n272 GNDA.n70 9.3005
R514 GNDA.n274 GNDA.n273 9.3005
R515 GNDA.n275 GNDA.n68 9.3005
R516 GNDA.n278 GNDA.n277 9.3005
R517 GNDA.n279 GNDA.n67 9.3005
R518 GNDA.n281 GNDA.n280 9.3005
R519 GNDA.n282 GNDA.n65 9.3005
R520 GNDA.n285 GNDA.n284 9.3005
R521 GNDA.n286 GNDA.n64 9.3005
R522 GNDA.n288 GNDA.n287 9.3005
R523 GNDA.n289 GNDA.n62 9.3005
R524 GNDA.n292 GNDA.n291 9.3005
R525 GNDA.n293 GNDA.n55 9.3005
R526 GNDA.n296 GNDA.n295 9.3005
R527 GNDA.n297 GNDA.n53 9.3005
R528 GNDA.n300 GNDA.n299 9.3005
R529 GNDA.n301 GNDA.n51 9.3005
R530 GNDA.n307 GNDA.n306 9.3005
R531 GNDA.n305 GNDA.n52 9.3005
R532 GNDA.n304 GNDA.n303 9.3005
R533 GNDA.n322 GNDA.n48 9.3005
R534 GNDA.n324 GNDA.n323 9.3005
R535 GNDA.n325 GNDA.n46 9.3005
R536 GNDA.n328 GNDA.n327 9.3005
R537 GNDA.n329 GNDA.n45 9.3005
R538 GNDA.n331 GNDA.n330 9.3005
R539 GNDA.n332 GNDA.n43 9.3005
R540 GNDA.n335 GNDA.n334 9.3005
R541 GNDA.n336 GNDA.n42 9.3005
R542 GNDA.n338 GNDA.n337 9.3005
R543 GNDA.n339 GNDA.n41 9.3005
R544 GNDA.n341 GNDA.n340 9.3005
R545 GNDA.n343 GNDA.n342 9.3005
R546 GNDA.n344 GNDA.n39 9.3005
R547 GNDA.n346 GNDA.n345 9.3005
R548 GNDA.n348 GNDA.n347 9.3005
R549 GNDA.n349 GNDA.n37 9.3005
R550 GNDA.n351 GNDA.n350 9.3005
R551 GNDA.n352 GNDA.n36 9.3005
R552 GNDA.n354 GNDA.n353 9.3005
R553 GNDA.n35 GNDA.n34 9.3005
R554 GNDA.n365 GNDA.n364 9.3005
R555 GNDA.n366 GNDA.n33 9.3005
R556 GNDA.n368 GNDA.n367 9.3005
R557 GNDA.n369 GNDA.n32 9.3005
R558 GNDA.n371 GNDA.n370 9.3005
R559 GNDA.n372 GNDA.n31 9.3005
R560 GNDA.n374 GNDA.n373 9.3005
R561 GNDA.n375 GNDA.n30 9.3005
R562 GNDA.n377 GNDA.n376 9.3005
R563 GNDA.n379 GNDA.n378 9.3005
R564 GNDA.n381 GNDA.n27 9.3005
R565 GNDA.n383 GNDA.n382 9.3005
R566 GNDA.n384 GNDA.n26 9.3005
R567 GNDA.n386 GNDA.n385 9.3005
R568 GNDA.n387 GNDA.n25 9.3005
R569 GNDA.n389 GNDA.n388 9.3005
R570 GNDA.n390 GNDA.n24 9.3005
R571 GNDA.n392 GNDA.n391 9.3005
R572 GNDA.n194 GNDA.n193 9.3005
R573 GNDA.n195 GNDA.n191 9.3005
R574 GNDA.n190 GNDA.n88 9.3005
R575 GNDA.n189 GNDA.n188 9.3005
R576 GNDA.n186 GNDA.n89 9.3005
R577 GNDA.n185 GNDA.n184 9.3005
R578 GNDA.n183 GNDA.n90 9.3005
R579 GNDA.n182 GNDA.n181 9.3005
R580 GNDA.n92 GNDA.n91 9.3005
R581 GNDA.n146 GNDA.n145 9.3005
R582 GNDA.n147 GNDA.n144 9.3005
R583 GNDA.n127 GNDA.n112 9.3005
R584 GNDA.n129 GNDA.n128 9.3005
R585 GNDA.n130 GNDA.n111 9.3005
R586 GNDA.n132 GNDA.n131 9.3005
R587 GNDA.n133 GNDA.n109 9.3005
R588 GNDA.n135 GNDA.n134 9.3005
R589 GNDA.n136 GNDA.n107 9.3005
R590 GNDA.n164 GNDA.n163 9.3005
R591 GNDA.n162 GNDA.n108 9.3005
R592 GNDA.n161 GNDA.n160 9.3005
R593 GNDA.n159 GNDA.n137 9.3005
R594 GNDA.n158 GNDA.n157 9.3005
R595 GNDA.n156 GNDA.n140 9.3005
R596 GNDA.n155 GNDA.n154 9.3005
R597 GNDA.n153 GNDA.n141 9.3005
R598 GNDA.n152 GNDA.n151 9.3005
R599 GNDA.n150 GNDA.n143 9.3005
R600 GNDA.n149 GNDA.n148 9.3005
R601 GNDA.n242 GNDA.n241 9.3005
R602 GNDA.n240 GNDA.n81 9.3005
R603 GNDA.n239 GNDA.n238 9.3005
R604 GNDA.n237 GNDA.n82 9.3005
R605 GNDA.n236 GNDA.n235 9.3005
R606 GNDA.n234 GNDA.n83 9.3005
R607 GNDA.n233 GNDA.n232 9.3005
R608 GNDA.n231 GNDA.n209 9.3005
R609 GNDA.n230 GNDA.n229 9.3005
R610 GNDA.n228 GNDA.n210 9.3005
R611 GNDA.n227 GNDA.n226 9.3005
R612 GNDA.n225 GNDA.n211 9.3005
R613 GNDA.n224 GNDA.n223 9.3005
R614 GNDA.n222 GNDA.n213 9.3005
R615 GNDA.n220 GNDA.n219 9.3005
R616 GNDA.n218 GNDA.n215 9.3005
R617 GNDA.n217 GNDA.n216 9.3005
R618 GNDA.n22 GNDA.n21 9.3005
R619 GNDA.n406 GNDA.n405 9.3005
R620 GNDA.n407 GNDA.n20 9.3005
R621 GNDA.n409 GNDA.n408 9.3005
R622 GNDA.n410 GNDA.n18 9.3005
R623 GNDA.n413 GNDA.n412 9.3005
R624 GNDA.n414 GNDA.n17 9.3005
R625 GNDA.n416 GNDA.n415 9.3005
R626 GNDA.n418 GNDA.n15 9.3005
R627 GNDA.n420 GNDA.n419 9.3005
R628 GNDA.n421 GNDA.n14 9.3005
R629 GNDA.n423 GNDA.n422 9.3005
R630 GNDA.n425 GNDA.n12 9.3005
R631 GNDA.n427 GNDA.n426 9.3005
R632 GNDA.n428 GNDA.n11 9.3005
R633 GNDA.n430 GNDA.n429 9.3005
R634 GNDA.n431 GNDA.n10 9.3005
R635 GNDA.n433 GNDA.n432 9.3005
R636 GNDA.n434 GNDA.n9 9.3005
R637 GNDA.n436 GNDA.n435 9.3005
R638 GNDA.n438 GNDA.n6 9.3005
R639 GNDA.n441 GNDA.n440 9.3005
R640 GNDA.n442 GNDA.n5 9.3005
R641 GNDA.n444 GNDA.n443 9.3005
R642 GNDA.n445 GNDA.n4 9.3005
R643 GNDA.n447 GNDA.n446 9.3005
R644 GNDA.n448 GNDA.n3 9.3005
R645 GNDA.n450 GNDA.n449 9.3005
R646 GNDA.n451 GNDA.n1 9.3005
R647 GNDA.n245 GNDA.n78 8.9605
R648 GNDA.t141 GNDA.t122 8.54087
R649 GNDA.t144 GNDA.t87 8.54087
R650 GNDA.n321 GNDA.n320 7.49888
R651 GNDA.n118 GNDA.n117 7.11161
R652 GNDA.n123 GNDA.n114 7.11161
R653 GNDA.n202 GNDA.n201 7.11161
R654 GNDA.n199 GNDA.n197 7.11161
R655 GNDA.n126 GNDA.n125 6.69883
R656 GNDA.n133 GNDA.n132 6.4005
R657 GNDA.n153 GNDA.n152 6.4005
R658 GNDA.n148 GNDA.n147 6.4005
R659 GNDA.n245 GNDA 6.4005
R660 GNDA.n294 GNDA.n293 6.4005
R661 GNDA.n334 GNDA.n333 6.4005
R662 GNDA.n355 GNDA.n354 6.4005
R663 GNDA.n363 GNDA.n33 6.4005
R664 GNDA.n376 GNDA.n29 6.4005
R665 GNDA.n381 GNDA.n380 6.4005
R666 GNDA.n393 GNDA.n392 6.4005
R667 GNDA.n221 GNDA.n220 6.4005
R668 GNDA.n405 GNDA.n404 6.4005
R669 GNDA.n418 GNDA.n417 6.4005
R670 GNDA.n425 GNDA.n424 6.4005
R671 GNDA.n437 GNDA.n436 6.4005
R672 GNDA.n452 GNDA.n451 6.4005
R673 GNDA.n195 GNDA.n194 6.4005
R674 GNDA.n359 GNDA.n358 5.68939
R675 GNDA.n359 GNDA.n28 5.68939
R676 GNDA.n397 GNDA.n8 5.68939
R677 GNDA.n397 GNDA.n7 4.97828
R678 GNDA.n117 GNDA.n116 3.48951
R679 GNDA.n116 GNDA.n114 3.48951
R680 GNDA.n201 GNDA.n200 3.48951
R681 GNDA.n200 GNDA.n199 3.48951
R682 GNDA.n327 GNDA.n326 3.2005
R683 GNDA.n340 GNDA.n40 3.2005
R684 GNDA.n96 GNDA.n93 2.25882
R685 GNDA.n96 GNDA.n95 2.25882
R686 GNDA.n178 GNDA.n94 2.25882
R687 GNDA.n177 GNDA.n95 2.25882
R688 GNDA.n172 GNDA.n93 2.25882
R689 GNDA.n178 GNDA.n177 2.25882
R690 GNDA.n102 GNDA.n101 2.25882
R691 GNDA.n103 GNDA.n102 2.25882
R692 GNDA.n165 GNDA.n106 2.25882
R693 GNDA.n105 GNDA.n103 2.25882
R694 GNDA.n167 GNDA.n101 2.25882
R695 GNDA.n106 GNDA.n105 2.25882
R696 GNDA.n79 GNDA.n49 1.0063
R697 GNDA.n125 GNDA.n112 0.703977
R698 GNDA.n322 GNDA.n321 0.193977
R699 GNDA.n391 GNDA.n0 0.193881
R700 GNDA.n453 GNDA.n1 0.193881
R701 GNDA.n243 GNDA.n242 0.193695
R702 GNDA.n303 GNDA.n302 0.188
R703 GNDA.n268 GNDA.n267 0.15675
R704 GNDA.n270 GNDA.n70 0.15675
R705 GNDA.n274 GNDA.n70 0.15675
R706 GNDA.n275 GNDA.n274 0.15675
R707 GNDA.n277 GNDA.n67 0.15675
R708 GNDA.n281 GNDA.n67 0.15675
R709 GNDA.n282 GNDA.n281 0.15675
R710 GNDA.n284 GNDA.n64 0.15675
R711 GNDA.n288 GNDA.n64 0.15675
R712 GNDA.n289 GNDA.n288 0.15675
R713 GNDA.n291 GNDA.n55 0.15675
R714 GNDA.n296 GNDA.n55 0.15675
R715 GNDA.n297 GNDA.n296 0.15675
R716 GNDA.n299 GNDA.n51 0.15675
R717 GNDA.n307 GNDA.n52 0.15675
R718 GNDA.n303 GNDA.n52 0.15675
R719 GNDA.n323 GNDA.n322 0.15675
R720 GNDA.n323 GNDA.n46 0.15675
R721 GNDA.n328 GNDA.n46 0.15675
R722 GNDA.n329 GNDA.n328 0.15675
R723 GNDA.n330 GNDA.n329 0.15675
R724 GNDA.n330 GNDA.n43 0.15675
R725 GNDA.n335 GNDA.n43 0.15675
R726 GNDA.n336 GNDA.n335 0.15675
R727 GNDA.n337 GNDA.n336 0.15675
R728 GNDA.n337 GNDA.n41 0.15675
R729 GNDA.n341 GNDA.n41 0.15675
R730 GNDA.n342 GNDA.n341 0.15675
R731 GNDA.n342 GNDA.n39 0.15675
R732 GNDA.n346 GNDA.n39 0.15675
R733 GNDA.n347 GNDA.n346 0.15675
R734 GNDA.n347 GNDA.n37 0.15675
R735 GNDA.n351 GNDA.n37 0.15675
R736 GNDA.n352 GNDA.n351 0.15675
R737 GNDA.n353 GNDA.n352 0.15675
R738 GNDA.n353 GNDA.n34 0.15675
R739 GNDA.n365 GNDA.n34 0.15675
R740 GNDA.n366 GNDA.n365 0.15675
R741 GNDA.n367 GNDA.n366 0.15675
R742 GNDA.n367 GNDA.n32 0.15675
R743 GNDA.n371 GNDA.n32 0.15675
R744 GNDA.n372 GNDA.n371 0.15675
R745 GNDA.n373 GNDA.n372 0.15675
R746 GNDA.n373 GNDA.n30 0.15675
R747 GNDA.n377 GNDA.n30 0.15675
R748 GNDA.n378 GNDA.n377 0.15675
R749 GNDA.n378 GNDA.n27 0.15675
R750 GNDA.n383 GNDA.n27 0.15675
R751 GNDA.n384 GNDA.n383 0.15675
R752 GNDA.n385 GNDA.n384 0.15675
R753 GNDA.n385 GNDA.n25 0.15675
R754 GNDA.n389 GNDA.n25 0.15675
R755 GNDA.n390 GNDA.n389 0.15675
R756 GNDA.n391 GNDA.n390 0.15675
R757 GNDA.n129 GNDA.n112 0.15675
R758 GNDA.n130 GNDA.n129 0.15675
R759 GNDA.n131 GNDA.n130 0.15675
R760 GNDA.n131 GNDA.n109 0.15675
R761 GNDA.n135 GNDA.n109 0.15675
R762 GNDA.n136 GNDA.n135 0.15675
R763 GNDA.n163 GNDA.n136 0.15675
R764 GNDA.n163 GNDA.n162 0.15675
R765 GNDA.n162 GNDA.n161 0.15675
R766 GNDA.n161 GNDA.n137 0.15675
R767 GNDA.n157 GNDA.n137 0.15675
R768 GNDA.n157 GNDA.n156 0.15675
R769 GNDA.n156 GNDA.n155 0.15675
R770 GNDA.n155 GNDA.n141 0.15675
R771 GNDA.n151 GNDA.n141 0.15675
R772 GNDA.n151 GNDA.n150 0.15675
R773 GNDA.n150 GNDA.n149 0.15675
R774 GNDA.n149 GNDA.n144 0.15675
R775 GNDA.n145 GNDA.n144 0.15675
R776 GNDA.n145 GNDA.n91 0.15675
R777 GNDA.n182 GNDA.n91 0.15675
R778 GNDA.n183 GNDA.n182 0.15675
R779 GNDA.n184 GNDA.n183 0.15675
R780 GNDA.n184 GNDA.n89 0.15675
R781 GNDA.n189 GNDA.n89 0.15675
R782 GNDA.n190 GNDA.n189 0.15675
R783 GNDA.n191 GNDA.n190 0.15675
R784 GNDA.n193 GNDA.n191 0.15675
R785 GNDA.n242 GNDA.n81 0.15675
R786 GNDA.n238 GNDA.n81 0.15675
R787 GNDA.n238 GNDA.n237 0.15675
R788 GNDA.n237 GNDA.n236 0.15675
R789 GNDA.n236 GNDA.n83 0.15675
R790 GNDA.n232 GNDA.n83 0.15675
R791 GNDA.n232 GNDA.n231 0.15675
R792 GNDA.n231 GNDA.n230 0.15675
R793 GNDA.n230 GNDA.n210 0.15675
R794 GNDA.n226 GNDA.n225 0.15675
R795 GNDA.n225 GNDA.n224 0.15675
R796 GNDA.n224 GNDA.n213 0.15675
R797 GNDA.n219 GNDA.n213 0.15675
R798 GNDA.n219 GNDA.n218 0.15675
R799 GNDA.n218 GNDA.n217 0.15675
R800 GNDA.n217 GNDA.n21 0.15675
R801 GNDA.n406 GNDA.n21 0.15675
R802 GNDA.n407 GNDA.n406 0.15675
R803 GNDA.n408 GNDA.n407 0.15675
R804 GNDA.n408 GNDA.n18 0.15675
R805 GNDA.n413 GNDA.n18 0.15675
R806 GNDA.n414 GNDA.n413 0.15675
R807 GNDA.n415 GNDA.n414 0.15675
R808 GNDA.n415 GNDA.n15 0.15675
R809 GNDA.n420 GNDA.n15 0.15675
R810 GNDA.n421 GNDA.n420 0.15675
R811 GNDA.n422 GNDA.n421 0.15675
R812 GNDA.n422 GNDA.n12 0.15675
R813 GNDA.n427 GNDA.n12 0.15675
R814 GNDA.n428 GNDA.n427 0.15675
R815 GNDA.n429 GNDA.n428 0.15675
R816 GNDA.n429 GNDA.n10 0.15675
R817 GNDA.n433 GNDA.n10 0.15675
R818 GNDA.n434 GNDA.n433 0.15675
R819 GNDA.n435 GNDA.n434 0.15675
R820 GNDA.n435 GNDA.n6 0.15675
R821 GNDA.n441 GNDA.n6 0.15675
R822 GNDA.n442 GNDA.n441 0.15675
R823 GNDA.n443 GNDA.n442 0.15675
R824 GNDA.n443 GNDA.n4 0.15675
R825 GNDA.n447 GNDA.n4 0.15675
R826 GNDA.n448 GNDA.n447 0.15675
R827 GNDA.n449 GNDA.n448 0.15675
R828 GNDA.n449 GNDA.n1 0.15675
R829 GNDA.n265 GNDA.n73 0.131895
R830 GNDA.n193 GNDA 0.1255
R831 GNDA.n212 GNDA.n210 0.109875
R832 GNDA.n244 GNDA.n79 0.0945
R833 GNDA.n269 GNDA.n268 0.09425
R834 GNDA.n276 GNDA.n275 0.09425
R835 GNDA.n283 GNDA.n282 0.09425
R836 GNDA.n290 GNDA.n289 0.09425
R837 GNDA.n298 GNDA.n297 0.09425
R838 GNDA.n308 GNDA.n51 0.09425
R839 GNDA.n267 GNDA.n73 0.063
R840 GNDA.n270 GNDA.n269 0.063
R841 GNDA.n277 GNDA.n276 0.063
R842 GNDA.n284 GNDA.n283 0.063
R843 GNDA.n291 GNDA.n290 0.063
R844 GNDA.n299 GNDA.n298 0.063
R845 GNDA.n308 GNDA.n307 0.063
R846 GNDA GNDA.n192 0.063
R847 GNDA.n226 GNDA.n212 0.047375
R848 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t6 401.668
R849 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.n4 325.248
R850 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n0 313
R851 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.t4 252.248
R852 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.n1 208.868
R853 opamp_cell_4_0.n_left.n2 opamp_cell_4_0.n_left.t2 192.8
R854 opamp_cell_4_0.n_left.n1 opamp_cell_4_0.n_left.t7 192.8
R855 opamp_cell_4_0.n_left.n4 opamp_cell_4_0.n_left.n3 152
R856 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t1 60.0005
R857 opamp_cell_4_0.n_left.n0 opamp_cell_4_0.n_left.t0 60.0005
R858 opamp_cell_4_0.n_left.n3 opamp_cell_4_0.n_left.n2 59.4472
R859 opamp_cell_4_0.n_left.t3 opamp_cell_4_0.n_left.n5 49.2505
R860 opamp_cell_4_0.n_left.n5 opamp_cell_4_0.n_left.t5 49.2505
R861 opamp_cell_4_0.n_right.t0 opamp_cell_4_0.n_right.n6 1010.36
R862 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.n2 416.101
R863 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n1 354.048
R864 opamp_cell_4_0.n_right.n3 opamp_cell_4_0.n_right.t6 289.2
R865 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.t5 289.2
R866 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.t7 289.2
R867 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.t8 289.2
R868 opamp_cell_4_0.n_right.n2 opamp_cell_4_0.n_right.n0 284.2
R869 opamp_cell_4_0.n_right.n6 opamp_cell_4_0.n_right.n5 208.868
R870 opamp_cell_4_0.n_right.n5 opamp_cell_4_0.n_right.n4 208.868
R871 opamp_cell_4_0.n_right.n4 opamp_cell_4_0.n_right.n3 208.868
R872 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t1 60.0005
R873 opamp_cell_4_0.n_right.n0 opamp_cell_4_0.n_right.t2 60.0005
R874 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t4 49.2505
R875 opamp_cell_4_0.n_right.n1 opamp_cell_4_0.n_right.t3 49.2505
R876 VDDA.n164 VDDA.n130 3803.21
R877 VDDA.n261 VDDA.t26 2266.27
R878 VDDA.n441 VDDA.n433 831.25
R879 VDDA.n436 VDDA.n435 831.25
R880 VDDA.n452 VDDA.n444 831.25
R881 VDDA.n447 VDDA.n446 831.25
R882 VDDA.n151 VDDA.n150 585
R883 VDDA.n263 VDDA.n60 585
R884 VDDA.n256 VDDA.n60 585
R885 VDDA.n200 VDDA.n199 585
R886 VDDA.n199 VDDA.n198 585
R887 VDDA.n362 VDDA.n357 585
R888 VDDA.n357 VDDA.n48 585
R889 VDDA.n291 VDDA.n55 585
R890 VDDA.n286 VDDA.n55 585
R891 VDDA.n348 VDDA.n343 585
R892 VDDA.n343 VDDA.n45 585
R893 VDDA.n328 VDDA.n42 585
R894 VDDA.n328 VDDA.n327 585
R895 VDDA.n339 VDDA.n334 585
R896 VDDA.n334 VDDA.n41 585
R897 VDDA.n434 VDDA.n433 585
R898 VDDA.n438 VDDA.n436 585
R899 VDDA.n445 VDDA.n444 585
R900 VDDA.n449 VDDA.n447 585
R901 VDDA.n366 VDDA.n50 585
R902 VDDA.n351 VDDA.n50 585
R903 VDDA.n253 VDDA.n246 585
R904 VDDA.n169 VDDA.n168 585
R905 VDDA.n169 VDDA.n125 585
R906 VDDA.n440 VDDA.t127 465.079
R907 VDDA.t127 VDDA.n439 465.079
R908 VDDA.n451 VDDA.t124 465.079
R909 VDDA.t124 VDDA.n450 465.079
R910 VDDA.n313 VDDA.t10 464.281
R911 VDDA.t10 VDDA.n312 464.281
R912 VDDA.n29 VDDA.t119 464.281
R913 VDDA.t119 VDDA.n26 464.281
R914 VDDA.n474 VDDA.t6 464.281
R915 VDDA.t6 VDDA.n18 464.281
R916 VDDA.t121 VDDA.n457 464.281
R917 VDDA.n458 VDDA.t121 464.281
R918 VDDA.n468 VDDA.t24 464.281
R919 VDDA.t24 VDDA.n467 464.281
R920 VDDA.t16 VDDA.n417 464.281
R921 VDDA.n418 VDDA.t16 464.281
R922 VDDA.n428 VDDA.t30 464.281
R923 VDDA.t30 VDDA.n427 464.281
R924 VDDA.n408 VDDA.t14 464.281
R925 VDDA.t14 VDDA.n407 464.281
R926 VDDA.t12 VDDA.n301 464.281
R927 VDDA.n302 VDDA.t12 464.281
R928 VDDA.t29 VDDA.n317 464.281
R929 VDDA.n318 VDDA.t29 464.281
R930 VDDA.n371 VDDA.t129 415.336
R931 VDDA.n157 VDDA.t95 384.967
R932 VDDA.n161 VDDA.t107 384.967
R933 VDDA.n205 VDDA.t114 384.967
R934 VDDA.n133 VDDA.t111 384.967
R935 VDDA.n150 VDDA.t84 374.878
R936 VDDA.n245 VDDA.t98 352.834
R937 VDDA.t97 VDDA.n130 341.991
R938 VDDA.n134 VDDA.t113 341.752
R939 VDDA.n162 VDDA.t110 341.752
R940 VDDA.n204 VDDA.t117 341.752
R941 VDDA.n197 VDDA.t104 336.329
R942 VDDA.n197 VDDA.t87 336.329
R943 VDDA.n126 VDDA.t101 320.7
R944 VDDA.n264 VDDA.t91 320.7
R945 VDDA.n158 VDDA.n156 315.647
R946 VDDA.n207 VDDA.n81 315.647
R947 VDDA.n132 VDDA.n82 315.647
R948 VDDA.n206 VDDA.n83 315.647
R949 VDDA.n159 VDDA.n138 315.647
R950 VDDA.n160 VDDA.n137 315.647
R951 VDDA.n23 VDDA.t22 315.25
R952 VDDA.t31 VDDA.t25 314.113
R953 VDDA.t122 VDDA.t2 314.113
R954 VDDA.n199 VDDA.n89 291.363
R955 VDDA.n195 VDDA.n87 291.363
R956 VDDA.n196 VDDA.n195 291.363
R957 VDDA.n151 VDDA.n140 290.733
R958 VDDA.n151 VDDA.n141 290.733
R959 VDDA.n257 VDDA.n60 290.733
R960 VDDA.n360 VDDA.n357 290.733
R961 VDDA.n289 VDDA.n55 290.733
R962 VDDA.n346 VDDA.n343 290.733
R963 VDDA.n329 VDDA.n328 290.733
R964 VDDA.n337 VDDA.n334 290.733
R965 VDDA.n352 VDDA.n50 290.733
R966 VDDA.n251 VDDA.n246 290.733
R967 VDDA.n247 VDDA.n246 290.733
R968 VDDA.n169 VDDA.n124 290.733
R969 VDDA.n429 VDDA.n428 243.698
R970 VDDA.n469 VDDA.n468 243.698
R971 VDDA.n475 VDDA.n474 243.698
R972 VDDA.n29 VDDA.n28 243.698
R973 VDDA.n314 VDDA.n313 243.698
R974 VDDA.n407 VDDA.n21 243.698
R975 VDDA.n302 VDDA.n299 243.698
R976 VDDA.n318 VDDA.n297 243.698
R977 VDDA.n458 VDDA.n455 243.698
R978 VDDA.n418 VDDA.n415 243.698
R979 VDDA.n414 VDDA.n1 238.367
R980 VDDA.n453 VDDA.n452 238.367
R981 VDDA.n446 VDDA.n413 238.367
R982 VDDA.n412 VDDA.n13 238.367
R983 VDDA.n478 VDDA.n477 238.367
R984 VDDA.n34 VDDA.n33 238.367
R985 VDDA.n298 VDDA.n38 238.367
R986 VDDA.n422 VDDA.n2 238.367
R987 VDDA.n442 VDDA.n441 238.367
R988 VDDA.n462 VDDA.n14 238.367
R989 VDDA.n410 VDDA.n409 238.367
R990 VDDA.n306 VDDA.n25 238.367
R991 VDDA.n322 VDDA.n37 238.367
R992 VDDA.n435 VDDA.n431 238.367
R993 VDDA.n143 VDDA.n141 233.841
R994 VDDA.n247 VDDA.n63 233.841
R995 VDDA.n254 VDDA.n253 230.308
R996 VDDA.n150 VDDA.n149 230.308
R997 VDDA.n263 VDDA.n262 230.308
R998 VDDA.n260 VDDA.n256 230.308
R999 VDDA.n201 VDDA.n200 230.308
R1000 VDDA.n198 VDDA.n84 230.308
R1001 VDDA.n340 VDDA.n339 230.308
R1002 VDDA.n296 VDDA.n41 230.308
R1003 VDDA.n349 VDDA.n348 230.308
R1004 VDDA.n295 VDDA.n45 230.308
R1005 VDDA.n363 VDDA.n362 230.308
R1006 VDDA.n294 VDDA.n48 230.308
R1007 VDDA.n292 VDDA.n291 230.308
R1008 VDDA.n286 VDDA.n53 230.308
R1009 VDDA.n332 VDDA.n42 230.308
R1010 VDDA.n366 VDDA.n365 230.308
R1011 VDDA.n355 VDDA.n351 230.308
R1012 VDDA.n327 VDDA.n324 230.308
R1013 VDDA.t7 VDDA.t66 222.178
R1014 VDDA.n341 VDDA.n323 199.195
R1015 VDDA.n98 VDDA.n97 196.502
R1016 VDDA.n95 VDDA.n94 196.502
R1017 VDDA.n194 VDDA.n193 196.502
R1018 VDDA.n185 VDDA.n117 196.502
R1019 VDDA.n178 VDDA.n120 196.502
R1020 VDDA.n171 VDDA.n170 196.502
R1021 VDDA.n163 VDDA.n162 185.001
R1022 VDDA.n135 VDDA.n134 185.001
R1023 VDDA.n204 VDDA.n203 185.001
R1024 VDDA.n52 VDDA.n51 185
R1025 VDDA.n354 VDDA.n353 185
R1026 VDDA.n331 VDDA.n330 185
R1027 VDDA.n326 VDDA.n325 185
R1028 VDDA.n321 VDDA.n320 185
R1029 VDDA.n319 VDDA.n316 185
R1030 VDDA.n305 VDDA.n304 185
R1031 VDDA.n303 VDDA.n300 185
R1032 VDDA.n404 VDDA.n22 185
R1033 VDDA.n406 VDDA.n405 185
R1034 VDDA.n461 VDDA.n460 185
R1035 VDDA.n459 VDDA.n456 185
R1036 VDDA.n434 VDDA.n432 185
R1037 VDDA.n438 VDDA.n437 185
R1038 VDDA.n421 VDDA.n420 185
R1039 VDDA.n419 VDDA.n416 185
R1040 VDDA.n290 VDDA.n54 185
R1041 VDDA.n288 VDDA.n287 185
R1042 VDDA.n361 VDDA.n356 185
R1043 VDDA.n359 VDDA.n358 185
R1044 VDDA.n347 VDDA.n342 185
R1045 VDDA.n345 VDDA.n344 185
R1046 VDDA.n338 VDDA.n333 185
R1047 VDDA.n336 VDDA.n335 185
R1048 VDDA.n309 VDDA.n308 185
R1049 VDDA.n311 VDDA.n310 185
R1050 VDDA.n30 VDDA.n27 185
R1051 VDDA.n32 VDDA.n31 185
R1052 VDDA.n473 VDDA.n471 185
R1053 VDDA.n472 VDDA.n19 185
R1054 VDDA.n464 VDDA.n463 185
R1055 VDDA.n466 VDDA.n465 185
R1056 VDDA.n445 VDDA.n443 185
R1057 VDDA.n449 VDDA.n448 185
R1058 VDDA.n424 VDDA.n423 185
R1059 VDDA.n426 VDDA.n425 185
R1060 VDDA.n88 VDDA.n85 185
R1061 VDDA.n91 VDDA.n90 185
R1062 VDDA.n62 VDDA.n61 185
R1063 VDDA.n259 VDDA.n258 185
R1064 VDDA.n148 VDDA.n142 185
R1065 VDDA.n147 VDDA.n146 185
R1066 VDDA.n147 VDDA.n136 185
R1067 VDDA.n145 VDDA.n144 185
R1068 VDDA.n252 VDDA.n65 185
R1069 VDDA.n250 VDDA.n64 185
R1070 VDDA.n255 VDDA.n64 185
R1071 VDDA.n249 VDDA.n248 185
R1072 VDDA.n168 VDDA.n127 185
R1073 VDDA.n164 VDDA.n127 185
R1074 VDDA.n167 VDDA.n166 185
R1075 VDDA.n129 VDDA.n128 185
R1076 VDDA.n131 VDDA.n125 185
R1077 VDDA.n164 VDDA.n131 185
R1078 VDDA.t66 VDDA.n293 172.38
R1079 VDDA.n364 VDDA.t19 172.38
R1080 VDDA.n350 VDDA.t17 172.38
R1081 VDDA.n198 VDDA.n197 166.63
R1082 VDDA.n425 VDDA.n423 150
R1083 VDDA.n448 VDDA.n443 150
R1084 VDDA.n465 VDDA.n463 150
R1085 VDDA.n471 VDDA.n19 150
R1086 VDDA.n32 VDDA.n27 150
R1087 VDDA.n310 VDDA.n308 150
R1088 VDDA.n421 VDDA.n416 150
R1089 VDDA.n437 VDDA.n432 150
R1090 VDDA.n461 VDDA.n456 150
R1091 VDDA.n405 VDDA.n22 150
R1092 VDDA.n305 VDDA.n300 150
R1093 VDDA.n321 VDDA.n316 150
R1094 VDDA.n315 VDDA.n307 137.904
R1095 VDDA.n411 VDDA.n20 137.904
R1096 VDDA.n293 VDDA.t26 126.412
R1097 VDDA.n364 VDDA.t7 126.412
R1098 VDDA.t19 VDDA.n350 126.412
R1099 VDDA.t17 VDDA.n341 126.412
R1100 VDDA.t128 VDDA.n433 123.126
R1101 VDDA.n436 VDDA.t128 123.126
R1102 VDDA.t126 VDDA.n444 123.126
R1103 VDDA.n447 VDDA.t126 123.126
R1104 VDDA.n65 VDDA.n64 120.001
R1105 VDDA.n248 VDDA.n64 120.001
R1106 VDDA.n148 VDDA.n147 120.001
R1107 VDDA.n147 VDDA.n144 120.001
R1108 VDDA.n259 VDDA.n62 120.001
R1109 VDDA.n90 VDDA.n85 120.001
R1110 VDDA.n335 VDDA.n333 120.001
R1111 VDDA.n344 VDDA.n342 120.001
R1112 VDDA.n358 VDDA.n356 120.001
R1113 VDDA.n287 VDDA.n54 120.001
R1114 VDDA.n331 VDDA.n325 120.001
R1115 VDDA.n354 VDDA.n52 120.001
R1116 VDDA.n166 VDDA.n127 120.001
R1117 VDDA.n131 VDDA.n129 120.001
R1118 VDDA.n233 VDDA.n69 119.737
R1119 VDDA.n226 VDDA.n72 119.737
R1120 VDDA.n219 VDDA.n75 119.737
R1121 VDDA.n212 VDDA.n78 119.737
R1122 VDDA.n154 VDDA.n152 119.737
R1123 VDDA.n476 VDDA.n470 107.258
R1124 VDDA.n470 VDDA.t23 103.427
R1125 VDDA.t123 VDDA.n454 103.427
R1126 VDDA.n454 VDDA.t125 103.427
R1127 VDDA.t15 VDDA.n430 103.427
R1128 VDDA.n476 VDDA.t13 95.7666
R1129 VDDA.t9 VDDA.t28 91.936
R1130 VDDA.t118 VDDA.t11 91.936
R1131 VDDA.t5 VDDA.t21 84.2747
R1132 VDDA.t23 VDDA.t31 84.2747
R1133 VDDA.t25 VDDA.t123 84.2747
R1134 VDDA.t125 VDDA.t122 84.2747
R1135 VDDA.t2 VDDA.t15 84.2747
R1136 VDDA.n207 VDDA.n82 83.2005
R1137 VDDA.n207 VDDA.n206 83.2005
R1138 VDDA.n159 VDDA.n158 83.2005
R1139 VDDA.n160 VDDA.n159 83.2005
R1140 VDDA.n365 VDDA.n364 69.8479
R1141 VDDA.n364 VDDA.n355 69.8479
R1142 VDDA.n341 VDDA.n332 69.8479
R1143 VDDA.n341 VDDA.n324 69.8479
R1144 VDDA.n293 VDDA.n292 69.8479
R1145 VDDA.n293 VDDA.n53 69.8479
R1146 VDDA.n364 VDDA.n363 69.8479
R1147 VDDA.n364 VDDA.n294 69.8479
R1148 VDDA.n350 VDDA.n349 69.8479
R1149 VDDA.n350 VDDA.n295 69.8479
R1150 VDDA.n341 VDDA.n340 69.8479
R1151 VDDA.n341 VDDA.n296 69.8479
R1152 VDDA.n202 VDDA.n201 69.8479
R1153 VDDA.n202 VDDA.n84 69.8479
R1154 VDDA.n262 VDDA.n261 69.8479
R1155 VDDA.n261 VDDA.n260 69.8479
R1156 VDDA.n149 VDDA.n136 69.8479
R1157 VDDA.n143 VDDA.n136 69.8479
R1158 VDDA.n255 VDDA.n254 69.8479
R1159 VDDA.n255 VDDA.n63 69.8479
R1160 VDDA.n165 VDDA.n164 69.8479
R1161 VDDA.n159 VDDA.n155 69.3203
R1162 VDDA.n323 VDDA.n322 65.8183
R1163 VDDA.n323 VDDA.n297 65.8183
R1164 VDDA.n307 VDDA.n306 65.8183
R1165 VDDA.n307 VDDA.n299 65.8183
R1166 VDDA.n411 VDDA.n410 65.8183
R1167 VDDA.n411 VDDA.n21 65.8183
R1168 VDDA.n470 VDDA.n462 65.8183
R1169 VDDA.n470 VDDA.n455 65.8183
R1170 VDDA.n454 VDDA.n442 65.8183
R1171 VDDA.n454 VDDA.n431 65.8183
R1172 VDDA.n430 VDDA.n422 65.8183
R1173 VDDA.n430 VDDA.n415 65.8183
R1174 VDDA.n315 VDDA.n314 65.8183
R1175 VDDA.n315 VDDA.n298 65.8183
R1176 VDDA.n28 VDDA.n20 65.8183
R1177 VDDA.n33 VDDA.n20 65.8183
R1178 VDDA.n476 VDDA.n475 65.8183
R1179 VDDA.n477 VDDA.n476 65.8183
R1180 VDDA.n470 VDDA.n469 65.8183
R1181 VDDA.n470 VDDA.n412 65.8183
R1182 VDDA.n454 VDDA.n453 65.8183
R1183 VDDA.n454 VDDA.n413 65.8183
R1184 VDDA.n430 VDDA.n429 65.8183
R1185 VDDA.n430 VDDA.n414 65.8183
R1186 VDDA.n389 VDDA.n38 58.0576
R1187 VDDA.n396 VDDA.n34 58.0576
R1188 VDDA.n479 VDDA.n478 58.0576
R1189 VDDA.n485 VDDA.n14 58.0576
R1190 VDDA.n485 VDDA.n13 58.0576
R1191 VDDA.n513 VDDA.n2 58.0576
R1192 VDDA.n513 VDDA.n1 58.0576
R1193 VDDA.n409 VDDA.n403 58.0576
R1194 VDDA.n397 VDDA.n25 58.0576
R1195 VDDA.n390 VDDA.n37 58.0576
R1196 VDDA.n367 VDDA.n48 57.2449
R1197 VDDA.n286 VDDA.n285 57.2449
R1198 VDDA.n374 VDDA.n45 57.2449
R1199 VDDA.n381 VDDA.n42 57.2449
R1200 VDDA.n381 VDDA.n41 57.2449
R1201 VDDA.n367 VDDA.n366 57.2449
R1202 VDDA.n498 VDDA.n8 54.4005
R1203 VDDA.n498 VDDA.n7 54.4005
R1204 VDDA.n500 VDDA.n7 54.4005
R1205 VDDA.n500 VDDA.n8 54.4005
R1206 VDDA.n416 VDDA.n415 53.3664
R1207 VDDA.n437 VDDA.n431 53.3664
R1208 VDDA.n456 VDDA.n455 53.3664
R1209 VDDA.n322 VDDA.n321 53.3664
R1210 VDDA.n316 VDDA.n297 53.3664
R1211 VDDA.n306 VDDA.n305 53.3664
R1212 VDDA.n300 VDDA.n299 53.3664
R1213 VDDA.n410 VDDA.n22 53.3664
R1214 VDDA.n405 VDDA.n21 53.3664
R1215 VDDA.n462 VDDA.n461 53.3664
R1216 VDDA.n442 VDDA.n432 53.3664
R1217 VDDA.n422 VDDA.n421 53.3664
R1218 VDDA.n314 VDDA.n308 53.3664
R1219 VDDA.n310 VDDA.n298 53.3664
R1220 VDDA.n28 VDDA.n27 53.3664
R1221 VDDA.n33 VDDA.n32 53.3664
R1222 VDDA.n475 VDDA.n471 53.3664
R1223 VDDA.n477 VDDA.n19 53.3664
R1224 VDDA.n469 VDDA.n463 53.3664
R1225 VDDA.n465 VDDA.n412 53.3664
R1226 VDDA.n453 VDDA.n443 53.3664
R1227 VDDA.n448 VDDA.n413 53.3664
R1228 VDDA.n429 VDDA.n423 53.3664
R1229 VDDA.n425 VDDA.n414 53.3664
R1230 VDDA.n156 VDDA.t97 49.2505
R1231 VDDA.n156 VDDA.t77 49.2505
R1232 VDDA.n81 VDDA.t73 49.2505
R1233 VDDA.n81 VDDA.t71 49.2505
R1234 VDDA.t113 VDDA.n132 49.2505
R1235 VDDA.n132 VDDA.t75 49.2505
R1236 VDDA.n83 VDDA.t69 49.2505
R1237 VDDA.n83 VDDA.t116 49.2505
R1238 VDDA.n138 VDDA.t79 49.2505
R1239 VDDA.n138 VDDA.t83 49.2505
R1240 VDDA.n137 VDDA.t81 49.2505
R1241 VDDA.n137 VDDA.t109 49.2505
R1242 VDDA.n248 VDDA.n63 45.3071
R1243 VDDA.n144 VDDA.n143 45.3071
R1244 VDDA.n325 VDDA.n324 45.3071
R1245 VDDA.n355 VDDA.n354 45.3071
R1246 VDDA.n365 VDDA.n52 45.3071
R1247 VDDA.n332 VDDA.n331 45.3071
R1248 VDDA.n292 VDDA.n54 45.3071
R1249 VDDA.n287 VDDA.n53 45.3071
R1250 VDDA.n363 VDDA.n356 45.3071
R1251 VDDA.n358 VDDA.n294 45.3071
R1252 VDDA.n349 VDDA.n342 45.3071
R1253 VDDA.n344 VDDA.n295 45.3071
R1254 VDDA.n340 VDDA.n333 45.3071
R1255 VDDA.n335 VDDA.n296 45.3071
R1256 VDDA.n201 VDDA.n85 45.3071
R1257 VDDA.n90 VDDA.n84 45.3071
R1258 VDDA.n262 VDDA.n62 45.3071
R1259 VDDA.n260 VDDA.n259 45.3071
R1260 VDDA.n149 VDDA.n148 45.3071
R1261 VDDA.n254 VDDA.n65 45.3071
R1262 VDDA.n166 VDDA.n165 45.3071
R1263 VDDA.n165 VDDA.n129 45.3071
R1264 VDDA.n208 VDDA.n207 41.6005
R1265 VDDA.n155 VDDA.n139 39.4988
R1266 VDDA.n271 VDDA.n270 38.1005
R1267 VDDA.t108 VDDA.n163 38.0466
R1268 VDDA.n514 VDDA.n513 34.9005
R1269 VDDA.t60 VDDA.t49 32.2821
R1270 VDDA.n200 VDDA.n86 32.2291
R1271 VDDA.n266 VDDA.n57 32.0005
R1272 VDDA.n270 VDDA.n57 32.0005
R1273 VDDA.n104 VDDA.n103 32.0005
R1274 VDDA.n103 VDDA.n102 32.0005
R1275 VDDA.n110 VDDA.n92 32.0005
R1276 VDDA.n110 VDDA.n109 32.0005
R1277 VDDA.n109 VDDA.n108 32.0005
R1278 VDDA.n192 VDDA.n114 32.0005
R1279 VDDA.n187 VDDA.n186 32.0005
R1280 VDDA.n180 VDDA.n179 32.0005
R1281 VDDA.n180 VDDA.n118 32.0005
R1282 VDDA.n184 VDDA.n118 32.0005
R1283 VDDA.n173 VDDA.n172 32.0005
R1284 VDDA.n173 VDDA.n121 32.0005
R1285 VDDA.n177 VDDA.n121 32.0005
R1286 VDDA.n284 VDDA.n274 32.0005
R1287 VDDA.n280 VDDA.n274 32.0005
R1288 VDDA.n280 VDDA.n279 32.0005
R1289 VDDA.n279 VDDA.n278 32.0005
R1290 VDDA.n278 VDDA.n49 32.0005
R1291 VDDA.n367 VDDA.n49 32.0005
R1292 VDDA.n368 VDDA.n367 32.0005
R1293 VDDA.n368 VDDA.n46 32.0005
R1294 VDDA.n373 VDDA.n46 32.0005
R1295 VDDA.n376 VDDA.n375 32.0005
R1296 VDDA.n376 VDDA.n43 32.0005
R1297 VDDA.n380 VDDA.n43 32.0005
R1298 VDDA.n383 VDDA.n382 32.0005
R1299 VDDA.n383 VDDA.n39 32.0005
R1300 VDDA.n387 VDDA.n39 32.0005
R1301 VDDA.n388 VDDA.n387 32.0005
R1302 VDDA.n391 VDDA.n35 32.0005
R1303 VDDA.n395 VDDA.n35 32.0005
R1304 VDDA.n399 VDDA.n398 32.0005
R1305 VDDA.n480 VDDA.n17 32.0005
R1306 VDDA.n484 VDDA.n15 32.0005
R1307 VDDA.n487 VDDA.n486 32.0005
R1308 VDDA.n487 VDDA.n11 32.0005
R1309 VDDA.n491 VDDA.n11 32.0005
R1310 VDDA.n492 VDDA.n491 32.0005
R1311 VDDA.n493 VDDA.n492 32.0005
R1312 VDDA.n493 VDDA.n9 32.0005
R1313 VDDA.n497 VDDA.n9 32.0005
R1314 VDDA.n501 VDDA.n5 32.0005
R1315 VDDA.n505 VDDA.n5 32.0005
R1316 VDDA.n506 VDDA.n505 32.0005
R1317 VDDA.n507 VDDA.n506 32.0005
R1318 VDDA.n507 VDDA.n3 32.0005
R1319 VDDA.n511 VDDA.n3 32.0005
R1320 VDDA.n512 VDDA.n511 32.0005
R1321 VDDA.n139 VDDA.n80 32.0005
R1322 VDDA.n209 VDDA.n80 32.0005
R1323 VDDA.n214 VDDA.n77 32.0005
R1324 VDDA.n215 VDDA.n214 32.0005
R1325 VDDA.n216 VDDA.n215 32.0005
R1326 VDDA.n216 VDDA.n74 32.0005
R1327 VDDA.n221 VDDA.n74 32.0005
R1328 VDDA.n222 VDDA.n221 32.0005
R1329 VDDA.n223 VDDA.n222 32.0005
R1330 VDDA.n223 VDDA.n71 32.0005
R1331 VDDA.n228 VDDA.n71 32.0005
R1332 VDDA.n229 VDDA.n228 32.0005
R1333 VDDA.n230 VDDA.n229 32.0005
R1334 VDDA.n230 VDDA.n68 32.0005
R1335 VDDA.n235 VDDA.n68 32.0005
R1336 VDDA.n236 VDDA.n235 32.0005
R1337 VDDA.n242 VDDA.n236 32.0005
R1338 VDDA.n242 VDDA.n241 32.0005
R1339 VDDA.n241 VDDA.n240 32.0005
R1340 VDDA.n240 VDDA.n237 32.0005
R1341 VDDA.n162 VDDA.n161 30.754
R1342 VDDA.n205 VDDA.n204 30.754
R1343 VDDA.n134 VDDA.n133 30.186
R1344 VDDA.t96 VDDA.t76 29.9762
R1345 VDDA.t78 VDDA.t82 29.9762
R1346 VDDA.t53 VDDA.t52 29.9762
R1347 VDDA.n157 VDDA.n130 29.9467
R1348 VDDA.t80 VDDA.t43 28.8233
R1349 VDDA.n265 VDDA.n59 28.8005
R1350 VDDA.n104 VDDA.n95 28.8005
R1351 VDDA.n193 VDDA.n192 28.8005
R1352 VDDA.n374 VDDA.n373 28.8005
R1353 VDDA.t33 VDDA.t56 27.6704
R1354 VDDA.t58 VDDA.t32 26.5175
R1355 VDDA.n285 VDDA.n284 25.6005
R1356 VDDA.n381 VDDA.n380 25.6005
R1357 VDDA.n391 VDDA.n390 25.6005
R1358 VDDA.n403 VDDA.n402 25.6005
R1359 VDDA.n479 VDDA.n15 25.6005
R1360 VDDA.n485 VDDA.n484 25.6005
R1361 VDDA.n499 VDDA.n498 25.6005
R1362 VDDA.n500 VDDA.n499 25.6005
R1363 VDDA.n209 VDDA.n208 25.6005
R1364 VDDA.n237 VDDA 25.6005
R1365 VDDA.t41 VDDA.n135 25.3646
R1366 VDDA.n97 VDDA.t1 24.6255
R1367 VDDA.n97 VDDA.t93 24.6255
R1368 VDDA.n94 VDDA.t50 24.6255
R1369 VDDA.n94 VDDA.t40 24.6255
R1370 VDDA.t106 VDDA.n194 24.6255
R1371 VDDA.n194 VDDA.t34 24.6255
R1372 VDDA.n117 VDDA.t48 24.6255
R1373 VDDA.n117 VDDA.t89 24.6255
R1374 VDDA.n120 VDDA.t44 24.6255
R1375 VDDA.n120 VDDA.t42 24.6255
R1376 VDDA.n170 VDDA.t103 24.6255
R1377 VDDA.n170 VDDA.t46 24.6255
R1378 VDDA.t103 VDDA.n169 24.6255
R1379 VDDA.n60 VDDA.t94 24.6255
R1380 VDDA.n195 VDDA.t106 24.6255
R1381 VDDA.n199 VDDA.t90 24.6255
R1382 VDDA.n50 VDDA.t8 24.6255
R1383 VDDA.n357 VDDA.t120 24.6255
R1384 VDDA.n55 VDDA.t27 24.6255
R1385 VDDA.n343 VDDA.t20 24.6255
R1386 VDDA.n328 VDDA.t51 24.6255
R1387 VDDA.n334 VDDA.t18 24.6255
R1388 VDDA.n126 VDDA.n123 24.361
R1389 VDDA.t35 VDDA.t39 24.2117
R1390 VDDA.t92 VDDA.t36 24.2117
R1391 VDDA.n102 VDDA.n98 22.4005
R1392 VDDA.n186 VDDA.n185 22.4005
R1393 VDDA.n187 VDDA.n86 22.4005
R1394 VDDA.n253 VDDA.n245 22.0449
R1395 VDDA.t45 VDDA.t80 21.9058
R1396 VDDA.t88 VDDA.t72 21.9058
R1397 VDDA.t37 VDDA.t70 21.9058
R1398 VDDA.n255 VDDA.t36 21.9058
R1399 VDDA.n202 VDDA.t3 20.7529
R1400 VDDA.t86 VDDA.n151 19.7005
R1401 VDDA.n246 VDDA.t100 19.7005
R1402 VDDA.n69 VDDA.t63 19.7005
R1403 VDDA.n69 VDDA.t99 19.7005
R1404 VDDA.n72 VDDA.t55 19.7005
R1405 VDDA.n72 VDDA.t59 19.7005
R1406 VDDA.n75 VDDA.t57 19.7005
R1407 VDDA.n75 VDDA.t61 19.7005
R1408 VDDA.n78 VDDA.t4 19.7005
R1409 VDDA.n78 VDDA.t38 19.7005
R1410 VDDA.n152 VDDA.t86 19.7005
R1411 VDDA.n152 VDDA.t65 19.7005
R1412 VDDA.t112 VDDA.t64 19.6
R1413 VDDA.n399 VDDA.n23 19.2005
R1414 VDDA.n265 VDDA.n264 17.6005
R1415 VDDA.t76 VDDA.t102 17.2942
R1416 VDDA.n203 VDDA.t60 16.1413
R1417 VDDA.n98 VDDA.n59 16.0005
R1418 VDDA.n114 VDDA.n86 16.0005
R1419 VDDA.n185 VDDA.n184 16.0005
R1420 VDDA.n172 VDDA.n171 16.0005
R1421 VDDA.n398 VDDA.n397 16.0005
R1422 VDDA.n161 VDDA.n160 16.0005
R1423 VDDA.n206 VDDA.n205 16.0005
R1424 VDDA.n133 VDDA.n82 16.0005
R1425 VDDA.n158 VDDA.n157 16.0005
R1426 VDDA VDDA.n56 15.7005
R1427 VDDA.n264 VDDA.n263 15.6449
R1428 VDDA.n168 VDDA.n126 15.6449
R1429 VDDA.t105 VDDA.t68 14.9884
R1430 VDDA.t115 VDDA.t105 14.9884
R1431 VDDA.t32 VDDA.t0 14.9884
R1432 VDDA.n285 VDDA.n273 13.8989
R1433 VDDA.t85 VDDA.t47 13.8355
R1434 VDDA.t49 VDDA.t54 13.8355
R1435 VDDA.n272 VDDA.n56 13.0501
R1436 VDDA.n396 VDDA.n395 12.8005
R1437 VDDA.n402 VDDA.n23 12.8005
R1438 VDDA.t102 VDDA.t78 12.6825
R1439 VDDA.t47 VDDA.t112 12.6825
R1440 VDDA.t54 VDDA.t35 12.6825
R1441 VDDA.n273 VDDA.n272 12.4261
R1442 VDDA.n272 VDDA.n271 11.7059
R1443 VDDA.n135 VDDA.t85 11.5296
R1444 VDDA.n323 VDDA.t9 11.4924
R1445 VDDA.t28 VDDA.n315 11.4924
R1446 VDDA.n307 VDDA.t118 11.4924
R1447 VDDA.t11 VDDA.n20 11.4924
R1448 VDDA.t21 VDDA.n411 11.4924
R1449 VDDA.t64 VDDA.t74 10.3767
R1450 VDDA.t62 VDDA.t53 10.3767
R1451 VDDA.n245 VDDA.n244 9.613
R1452 VDDA.n266 VDDA.n265 9.6005
R1453 VDDA.n193 VDDA.n92 9.6005
R1454 VDDA.n108 VDDA.n95 9.6005
R1455 VDDA.n238 VDDA.n237 9.3005
R1456 VDDA.n240 VDDA.n239 9.3005
R1457 VDDA.n241 VDDA.n67 9.3005
R1458 VDDA.n243 VDDA.n242 9.3005
R1459 VDDA.n236 VDDA.n66 9.3005
R1460 VDDA.n235 VDDA.n234 9.3005
R1461 VDDA.n232 VDDA.n68 9.3005
R1462 VDDA.n231 VDDA.n230 9.3005
R1463 VDDA.n229 VDDA.n70 9.3005
R1464 VDDA.n228 VDDA.n227 9.3005
R1465 VDDA.n225 VDDA.n71 9.3005
R1466 VDDA.n224 VDDA.n223 9.3005
R1467 VDDA.n222 VDDA.n73 9.3005
R1468 VDDA.n221 VDDA.n220 9.3005
R1469 VDDA.n218 VDDA.n74 9.3005
R1470 VDDA.n217 VDDA.n216 9.3005
R1471 VDDA.n215 VDDA.n76 9.3005
R1472 VDDA.n214 VDDA.n213 9.3005
R1473 VDDA.n211 VDDA.n77 9.3005
R1474 VDDA.n153 VDDA.n139 9.3005
R1475 VDDA.n80 VDDA.n79 9.3005
R1476 VDDA.n210 VDDA.n209 9.3005
R1477 VDDA.n172 VDDA.n122 9.3005
R1478 VDDA.n174 VDDA.n173 9.3005
R1479 VDDA.n175 VDDA.n121 9.3005
R1480 VDDA.n177 VDDA.n176 9.3005
R1481 VDDA.n179 VDDA.n119 9.3005
R1482 VDDA.n181 VDDA.n180 9.3005
R1483 VDDA.n182 VDDA.n118 9.3005
R1484 VDDA.n184 VDDA.n183 9.3005
R1485 VDDA.n185 VDDA.n116 9.3005
R1486 VDDA.n186 VDDA.n115 9.3005
R1487 VDDA.n188 VDDA.n187 9.3005
R1488 VDDA.n189 VDDA.n86 9.3005
R1489 VDDA.n190 VDDA.n114 9.3005
R1490 VDDA.n192 VDDA.n191 9.3005
R1491 VDDA.n193 VDDA.n113 9.3005
R1492 VDDA.n112 VDDA.n92 9.3005
R1493 VDDA.n111 VDDA.n110 9.3005
R1494 VDDA.n109 VDDA.n93 9.3005
R1495 VDDA.n108 VDDA.n107 9.3005
R1496 VDDA.n106 VDDA.n95 9.3005
R1497 VDDA.n105 VDDA.n104 9.3005
R1498 VDDA.n103 VDDA.n96 9.3005
R1499 VDDA.n102 VDDA.n101 9.3005
R1500 VDDA.n100 VDDA.n98 9.3005
R1501 VDDA.n99 VDDA.n59 9.3005
R1502 VDDA.n265 VDDA.n58 9.3005
R1503 VDDA.n267 VDDA.n266 9.3005
R1504 VDDA.n268 VDDA.n57 9.3005
R1505 VDDA.n270 VDDA.n269 9.3005
R1506 VDDA.n284 VDDA.n283 9.3005
R1507 VDDA.n282 VDDA.n274 9.3005
R1508 VDDA.n281 VDDA.n280 9.3005
R1509 VDDA.n279 VDDA.n275 9.3005
R1510 VDDA.n278 VDDA.n277 9.3005
R1511 VDDA.n276 VDDA.n49 9.3005
R1512 VDDA.n367 VDDA.n47 9.3005
R1513 VDDA.n369 VDDA.n368 9.3005
R1514 VDDA.n370 VDDA.n46 9.3005
R1515 VDDA.n373 VDDA.n372 9.3005
R1516 VDDA.n375 VDDA.n44 9.3005
R1517 VDDA.n377 VDDA.n376 9.3005
R1518 VDDA.n378 VDDA.n43 9.3005
R1519 VDDA.n380 VDDA.n379 9.3005
R1520 VDDA.n382 VDDA.n40 9.3005
R1521 VDDA.n384 VDDA.n383 9.3005
R1522 VDDA.n385 VDDA.n39 9.3005
R1523 VDDA.n387 VDDA.n386 9.3005
R1524 VDDA.n388 VDDA.n36 9.3005
R1525 VDDA.n392 VDDA.n391 9.3005
R1526 VDDA.n393 VDDA.n35 9.3005
R1527 VDDA.n395 VDDA.n394 9.3005
R1528 VDDA.n398 VDDA.n24 9.3005
R1529 VDDA.n400 VDDA.n399 9.3005
R1530 VDDA.n402 VDDA.n401 9.3005
R1531 VDDA.n17 VDDA.n16 9.3005
R1532 VDDA.n481 VDDA.n480 9.3005
R1533 VDDA.n482 VDDA.n15 9.3005
R1534 VDDA.n484 VDDA.n483 9.3005
R1535 VDDA.n486 VDDA.n12 9.3005
R1536 VDDA.n488 VDDA.n487 9.3005
R1537 VDDA.n489 VDDA.n11 9.3005
R1538 VDDA.n491 VDDA.n490 9.3005
R1539 VDDA.n492 VDDA.n10 9.3005
R1540 VDDA.n494 VDDA.n493 9.3005
R1541 VDDA.n495 VDDA.n9 9.3005
R1542 VDDA.n497 VDDA.n496 9.3005
R1543 VDDA.n499 VDDA.n6 9.3005
R1544 VDDA.n502 VDDA.n501 9.3005
R1545 VDDA.n503 VDDA.n5 9.3005
R1546 VDDA.n505 VDDA.n504 9.3005
R1547 VDDA.n506 VDDA.n4 9.3005
R1548 VDDA.n508 VDDA.n507 9.3005
R1549 VDDA.n509 VDDA.n3 9.3005
R1550 VDDA.n511 VDDA.n510 9.3005
R1551 VDDA.n512 VDDA.n0 9.3005
R1552 VDDA.n136 VDDA.t41 9.2238
R1553 VDDA.n311 VDDA.n309 9.14336
R1554 VDDA.n31 VDDA.n30 9.14336
R1555 VDDA.n473 VDDA.n472 9.14336
R1556 VDDA.n460 VDDA.n459 9.14336
R1557 VDDA.n466 VDDA.n464 9.14336
R1558 VDDA.n420 VDDA.n419 9.14336
R1559 VDDA.n426 VDDA.n424 9.14336
R1560 VDDA.n406 VDDA.n404 9.14336
R1561 VDDA.n304 VDDA.n303 9.14336
R1562 VDDA.n320 VDDA.n319 9.14336
R1563 VDDA.t82 VDDA.t45 8.07089
R1564 VDDA.t74 VDDA.t88 8.07089
R1565 VDDA.t68 VDDA.t37 8.07089
R1566 VDDA.t56 VDDA.t115 8.07089
R1567 VDDA.t13 VDDA.t5 7.66179
R1568 VDDA.n150 VDDA.n142 7.11161
R1569 VDDA.n146 VDDA.n145 7.11161
R1570 VDDA.n263 VDDA.n61 7.11161
R1571 VDDA.n258 VDDA.n256 7.11161
R1572 VDDA.n362 VDDA.n361 7.11161
R1573 VDDA.n359 VDDA.n48 7.11161
R1574 VDDA.n291 VDDA.n290 7.11161
R1575 VDDA.n288 VDDA.n286 7.11161
R1576 VDDA.n348 VDDA.n347 7.11161
R1577 VDDA.n345 VDDA.n45 7.11161
R1578 VDDA.n330 VDDA.n42 7.11161
R1579 VDDA.n327 VDDA.n326 7.11161
R1580 VDDA.n339 VDDA.n338 7.11161
R1581 VDDA.n336 VDDA.n41 7.11161
R1582 VDDA.n366 VDDA.n51 7.11161
R1583 VDDA.n353 VDDA.n351 7.11161
R1584 VDDA.n253 VDDA.n252 7.11161
R1585 VDDA.n250 VDDA.n249 7.11161
R1586 VDDA.n168 VDDA.n167 7.11161
R1587 VDDA.n128 VDDA.n125 7.11161
R1588 VDDA.n171 VDDA.n123 6.54033
R1589 VDDA.n382 VDDA.n381 6.4005
R1590 VDDA.n403 VDDA.n17 6.4005
R1591 VDDA.n480 VDDA.n479 6.4005
R1592 VDDA.n486 VDDA.n485 6.4005
R1593 VDDA.n498 VDDA.n497 6.4005
R1594 VDDA.n501 VDDA.n500 6.4005
R1595 VDDA.n513 VDDA.n512 6.4005
R1596 VDDA.n208 VDDA.n77 6.4005
R1597 VDDA.n438 VDDA.n434 5.81868
R1598 VDDA.n449 VDDA.n445 5.81868
R1599 VDDA.t72 VDDA.t3 5.76506
R1600 VDDA.t39 VDDA.t67 5.76506
R1601 VDDA.t52 VDDA.t92 5.76506
R1602 VDDA.n312 VDDA.n38 5.33286
R1603 VDDA.n34 VDDA.n26 5.33286
R1604 VDDA.n478 VDDA.n18 5.33286
R1605 VDDA.n457 VDDA.n14 5.33286
R1606 VDDA.n467 VDDA.n13 5.33286
R1607 VDDA.n417 VDDA.n2 5.33286
R1608 VDDA.n427 VDDA.n1 5.33286
R1609 VDDA.n409 VDDA.n408 5.33286
R1610 VDDA.n301 VDDA.n25 5.33286
R1611 VDDA.n317 VDDA.n37 5.33286
R1612 VDDA.t0 VDDA.t62 4.61215
R1613 VDDA.n313 VDDA.n309 3.75335
R1614 VDDA.n312 VDDA.n311 3.75335
R1615 VDDA.n30 VDDA.n29 3.75335
R1616 VDDA.n31 VDDA.n26 3.75335
R1617 VDDA.n474 VDDA.n473 3.75335
R1618 VDDA.n472 VDDA.n18 3.75335
R1619 VDDA.n460 VDDA.n457 3.75335
R1620 VDDA.n459 VDDA.n458 3.75335
R1621 VDDA.n468 VDDA.n464 3.75335
R1622 VDDA.n467 VDDA.n466 3.75335
R1623 VDDA.n420 VDDA.n417 3.75335
R1624 VDDA.n419 VDDA.n418 3.75335
R1625 VDDA.n428 VDDA.n424 3.75335
R1626 VDDA.n427 VDDA.n426 3.75335
R1627 VDDA.n408 VDDA.n404 3.75335
R1628 VDDA.n407 VDDA.n406 3.75335
R1629 VDDA.n304 VDDA.n301 3.75335
R1630 VDDA.n303 VDDA.n302 3.75335
R1631 VDDA.n320 VDDA.n317 3.75335
R1632 VDDA.n319 VDDA.n318 3.75335
R1633 VDDA.n142 VDDA.n140 3.53508
R1634 VDDA.n145 VDDA.n141 3.53508
R1635 VDDA.n146 VDDA.n140 3.53508
R1636 VDDA.n257 VDDA.n61 3.53508
R1637 VDDA.n258 VDDA.n257 3.53508
R1638 VDDA.n361 VDDA.n360 3.53508
R1639 VDDA.n360 VDDA.n359 3.53508
R1640 VDDA.n290 VDDA.n289 3.53508
R1641 VDDA.n289 VDDA.n288 3.53508
R1642 VDDA.n347 VDDA.n346 3.53508
R1643 VDDA.n346 VDDA.n345 3.53508
R1644 VDDA.n330 VDDA.n329 3.53508
R1645 VDDA.n329 VDDA.n326 3.53508
R1646 VDDA.n338 VDDA.n337 3.53508
R1647 VDDA.n337 VDDA.n336 3.53508
R1648 VDDA.n352 VDDA.n51 3.53508
R1649 VDDA.n353 VDDA.n352 3.53508
R1650 VDDA.n252 VDDA.n251 3.53508
R1651 VDDA.n249 VDDA.n247 3.53508
R1652 VDDA.n251 VDDA.n250 3.53508
R1653 VDDA.n167 VDDA.n124 3.53508
R1654 VDDA.n128 VDDA.n124 3.53508
R1655 VDDA.t70 VDDA.n202 3.45924
R1656 VDDA.t67 VDDA.t58 3.45924
R1657 VDDA.n441 VDDA.n440 3.40194
R1658 VDDA.n439 VDDA.n435 3.40194
R1659 VDDA.n452 VDDA.n451 3.40194
R1660 VDDA.n450 VDDA.n446 3.40194
R1661 VDDA.n179 VDDA.n178 3.2005
R1662 VDDA.n178 VDDA.n177 3.2005
R1663 VDDA.n375 VDDA.n374 3.2005
R1664 VDDA.n389 VDDA.n388 3.2005
R1665 VDDA.n390 VDDA.n389 3.2005
R1666 VDDA.n397 VDDA.n396 3.2005
R1667 VDDA.n440 VDDA.n434 2.39444
R1668 VDDA.n439 VDDA.n438 2.39444
R1669 VDDA.n451 VDDA.n445 2.39444
R1670 VDDA.n450 VDDA.n449 2.39444
R1671 VDDA.n441 VDDA.n8 2.32777
R1672 VDDA.n446 VDDA.n7 2.32777
R1673 VDDA.n163 VDDA.n136 2.30633
R1674 VDDA.n203 VDDA.t33 2.30633
R1675 VDDA.n261 VDDA.n255 2.30633
R1676 VDDA.n88 VDDA.n87 2.27782
R1677 VDDA.n89 VDDA.n88 2.27782
R1678 VDDA.n198 VDDA.n196 2.27782
R1679 VDDA.n91 VDDA.n89 2.27782
R1680 VDDA.n200 VDDA.n87 2.27782
R1681 VDDA.n196 VDDA.n91 2.27782
R1682 VDDA.n164 VDDA.t96 1.15341
R1683 VDDA.t43 VDDA.t108 1.15341
R1684 VDDA.n123 VDDA.n122 0.703395
R1685 VDDA.n283 VDDA.n273 0.193974
R1686 VDDA.n238 VDDA.n56 0.188
R1687 VDDA.n153 VDDA.n79 0.15675
R1688 VDDA.n210 VDDA.n79 0.15675
R1689 VDDA.n211 VDDA.n210 0.15675
R1690 VDDA.n213 VDDA.n76 0.15675
R1691 VDDA.n217 VDDA.n76 0.15675
R1692 VDDA.n218 VDDA.n217 0.15675
R1693 VDDA.n220 VDDA.n73 0.15675
R1694 VDDA.n224 VDDA.n73 0.15675
R1695 VDDA.n225 VDDA.n224 0.15675
R1696 VDDA.n227 VDDA.n70 0.15675
R1697 VDDA.n231 VDDA.n70 0.15675
R1698 VDDA.n232 VDDA.n231 0.15675
R1699 VDDA.n234 VDDA.n66 0.15675
R1700 VDDA.n243 VDDA.n67 0.15675
R1701 VDDA.n239 VDDA.n67 0.15675
R1702 VDDA.n239 VDDA.n238 0.15675
R1703 VDDA.n174 VDDA.n122 0.15675
R1704 VDDA.n175 VDDA.n174 0.15675
R1705 VDDA.n176 VDDA.n175 0.15675
R1706 VDDA.n176 VDDA.n119 0.15675
R1707 VDDA.n181 VDDA.n119 0.15675
R1708 VDDA.n182 VDDA.n181 0.15675
R1709 VDDA.n183 VDDA.n182 0.15675
R1710 VDDA.n183 VDDA.n116 0.15675
R1711 VDDA.n116 VDDA.n115 0.15675
R1712 VDDA.n188 VDDA.n115 0.15675
R1713 VDDA.n189 VDDA.n188 0.15675
R1714 VDDA.n190 VDDA.n189 0.15675
R1715 VDDA.n191 VDDA.n190 0.15675
R1716 VDDA.n191 VDDA.n113 0.15675
R1717 VDDA.n113 VDDA.n112 0.15675
R1718 VDDA.n112 VDDA.n111 0.15675
R1719 VDDA.n111 VDDA.n93 0.15675
R1720 VDDA.n107 VDDA.n93 0.15675
R1721 VDDA.n107 VDDA.n106 0.15675
R1722 VDDA.n106 VDDA.n105 0.15675
R1723 VDDA.n105 VDDA.n96 0.15675
R1724 VDDA.n101 VDDA.n96 0.15675
R1725 VDDA.n101 VDDA.n100 0.15675
R1726 VDDA.n100 VDDA.n99 0.15675
R1727 VDDA.n99 VDDA.n58 0.15675
R1728 VDDA.n267 VDDA.n58 0.15675
R1729 VDDA.n268 VDDA.n267 0.15675
R1730 VDDA.n269 VDDA.n268 0.15675
R1731 VDDA.n283 VDDA.n282 0.15675
R1732 VDDA.n282 VDDA.n281 0.15675
R1733 VDDA.n281 VDDA.n275 0.15675
R1734 VDDA.n277 VDDA.n275 0.15675
R1735 VDDA.n277 VDDA.n276 0.15675
R1736 VDDA.n276 VDDA.n47 0.15675
R1737 VDDA.n369 VDDA.n47 0.15675
R1738 VDDA.n370 VDDA.n369 0.15675
R1739 VDDA.n372 VDDA.n44 0.15675
R1740 VDDA.n377 VDDA.n44 0.15675
R1741 VDDA.n378 VDDA.n377 0.15675
R1742 VDDA.n379 VDDA.n378 0.15675
R1743 VDDA.n379 VDDA.n40 0.15675
R1744 VDDA.n384 VDDA.n40 0.15675
R1745 VDDA.n385 VDDA.n384 0.15675
R1746 VDDA.n386 VDDA.n385 0.15675
R1747 VDDA.n386 VDDA.n36 0.15675
R1748 VDDA.n392 VDDA.n36 0.15675
R1749 VDDA.n393 VDDA.n392 0.15675
R1750 VDDA.n394 VDDA.n393 0.15675
R1751 VDDA.n394 VDDA.n24 0.15675
R1752 VDDA.n400 VDDA.n24 0.15675
R1753 VDDA.n401 VDDA.n400 0.15675
R1754 VDDA.n401 VDDA.n16 0.15675
R1755 VDDA.n481 VDDA.n16 0.15675
R1756 VDDA.n482 VDDA.n481 0.15675
R1757 VDDA.n483 VDDA.n482 0.15675
R1758 VDDA.n483 VDDA.n12 0.15675
R1759 VDDA.n488 VDDA.n12 0.15675
R1760 VDDA.n489 VDDA.n488 0.15675
R1761 VDDA.n490 VDDA.n489 0.15675
R1762 VDDA.n490 VDDA.n10 0.15675
R1763 VDDA.n494 VDDA.n10 0.15675
R1764 VDDA.n495 VDDA.n494 0.15675
R1765 VDDA.n496 VDDA.n495 0.15675
R1766 VDDA.n496 VDDA.n6 0.15675
R1767 VDDA.n502 VDDA.n6 0.15675
R1768 VDDA.n503 VDDA.n502 0.15675
R1769 VDDA.n504 VDDA.n503 0.15675
R1770 VDDA.n504 VDDA.n4 0.15675
R1771 VDDA.n508 VDDA.n4 0.15675
R1772 VDDA.n509 VDDA.n508 0.15675
R1773 VDDA.n510 VDDA.n509 0.15675
R1774 VDDA.n510 VDDA.n0 0.15675
R1775 VDDA.n514 VDDA.n0 0.15675
R1776 VDDA VDDA.n514 0.1255
R1777 VDDA.n269 VDDA 0.122375
R1778 VDDA.n155 VDDA.n154 0.100307
R1779 VDDA.n154 VDDA.n153 0.09425
R1780 VDDA.n213 VDDA.n212 0.09425
R1781 VDDA.n220 VDDA.n219 0.09425
R1782 VDDA.n227 VDDA.n226 0.09425
R1783 VDDA.n234 VDDA.n233 0.09425
R1784 VDDA.n244 VDDA.n243 0.09425
R1785 VDDA.n371 VDDA.n370 0.078625
R1786 VDDA.n372 VDDA.n371 0.078625
R1787 VDDA.n212 VDDA.n211 0.063
R1788 VDDA.n219 VDDA.n218 0.063
R1789 VDDA.n226 VDDA.n225 0.063
R1790 VDDA.n233 VDDA.n232 0.063
R1791 VDDA.n244 VDDA.n66 0.063
R1792 VDDA.n271 VDDA 0.0505
R1793 opamp_cell_4_0.VOUT pfd_8_0.opamp_out.n6 3993.6
R1794 pfd_8_0.opamp_out.n6 pfd_8_0.opamp_out.n4 823.75
R1795 pfd_8_0.opamp_out.n6 pfd_8_0.opamp_out.n5 753.326
R1796 pfd_8_0.opamp_out.n13 pfd_8_0.opamp_out.n12 424.447
R1797 pfd_8_0.opamp_out.n13 pfd_8_0.opamp_out.n11 354.048
R1798 pfd_8_0.opamp_out.n9 pfd_8_0.opamp_out.n8 313
R1799 pfd_8_0.opamp_out.t14 pfd_8_0.opamp_out.n0 297.233
R1800 pfd_8_0.opamp_out.n1 pfd_8_0.opamp_out.t14 297.233
R1801 pfd_8_0.opamp_out.n2 pfd_8_0.opamp_out.t13 297.233
R1802 pfd_8_0.opamp_out.n5 pfd_8_0.opamp_out.t5 281.596
R1803 pfd_8_0.opamp_out.n9 pfd_8_0.opamp_out.n7 242.601
R1804 pfd_8_0.opamp_out.n10 pfd_8_0.opamp_out.n9 220.8
R1805 pfd_8_0.opamp_out.n14 pfd_8_0.opamp_out.n13 220.8
R1806 pfd_8_0.opamp_out.n2 pfd_8_0.opamp_out.n1 216.9
R1807 pfd_8_0.opamp_out.n3 pfd_8_0.opamp_out.n0 216.9
R1808 charge_pump_cell_6_0.opamp_out pfd_8_0.opamp_out.n3 176.733
R1809 pfd_8_0.opamp_out.n5 pfd_8_0.opamp_out.t4 118.666
R1810 pfd_8_0.opamp_out.n1 pfd_8_0.opamp_out.t11 80.3338
R1811 pfd_8_0.opamp_out.t11 pfd_8_0.opamp_out.n0 80.3338
R1812 pfd_8_0.opamp_out.t12 pfd_8_0.opamp_out.n2 80.3338
R1813 pfd_8_0.opamp_out.n3 pfd_8_0.opamp_out.t12 80.3338
R1814 pfd_8_0.opamp_out.n4 pfd_8_0.opamp_out.t13 80.3338
R1815 pfd_8_0.opamp_out.n10 pfd_8_0.opamp_out.t15 70.0829
R1816 pfd_8_0.opamp_out.n15 pfd_8_0.opamp_out.n14 64.0005
R1817 pfd_8_0.opamp_out.n14 pfd_8_0.opamp_out.t10 63.6829
R1818 pfd_8_0.opamp_out.n15 pfd_8_0.opamp_out.n10 60.8005
R1819 pfd_8_0.opamp_out.n7 pfd_8_0.opamp_out.t0 60.0005
R1820 pfd_8_0.opamp_out.n7 pfd_8_0.opamp_out.t1 60.0005
R1821 pfd_8_0.opamp_out.n8 pfd_8_0.opamp_out.t2 60.0005
R1822 pfd_8_0.opamp_out.n8 pfd_8_0.opamp_out.t3 60.0005
R1823 pfd_8_0.opamp_out.n11 pfd_8_0.opamp_out.t6 49.2505
R1824 pfd_8_0.opamp_out.n11 pfd_8_0.opamp_out.t7 49.2505
R1825 pfd_8_0.opamp_out.n12 pfd_8_0.opamp_out.t9 49.2505
R1826 pfd_8_0.opamp_out.n12 pfd_8_0.opamp_out.t8 49.2505
R1827 pfd_8_0.opamp_out.n4 charge_pump_cell_6_0.opamp_out 16.0672
R1828 opamp_cell_4_0.VOUT pfd_8_0.opamp_out.n15 6.4005
R1829 a_6380_5710.n4 a_6380_5710.n0 427.647
R1830 a_6380_5710.n1 a_6380_5710.t6 321.334
R1831 a_6380_5710.n5 a_6380_5710.n4 210.601
R1832 a_6380_5710.n2 a_6380_5710.n1 208.868
R1833 a_6380_5710.n3 a_6380_5710.t2 174.056
R1834 a_6380_5710.n4 a_6380_5710.n3 152
R1835 a_6380_5710.n1 a_6380_5710.t7 112.468
R1836 a_6380_5710.n2 a_6380_5710.t4 112.468
R1837 a_6380_5710.n3 a_6380_5710.n2 61.5894
R1838 a_6380_5710.n5 a_6380_5710.t5 60.0005
R1839 a_6380_5710.t3 a_6380_5710.n5 60.0005
R1840 a_6380_5710.n0 a_6380_5710.t1 49.2505
R1841 a_6380_5710.n0 a_6380_5710.t0 49.2505
R1842 a_6500_6300.n7 a_6500_6300.n5 482.582
R1843 a_6500_6300.n10 a_6500_6300.t6 304.634
R1844 a_6500_6300.n3 a_6500_6300.t4 304.634
R1845 a_6500_6300.t8 a_6500_6300.n10 277.914
R1846 a_6500_6300.n3 a_6500_6300.t5 276.289
R1847 a_6500_6300.n8 a_6500_6300.n1 204.201
R1848 a_6500_6300.n4 a_6500_6300.n2 204.201
R1849 a_6500_6300.n9 a_6500_6300.n0 204.201
R1850 a_6500_6300.n7 a_6500_6300.n6 120.981
R1851 a_6500_6300.n8 a_6500_6300.n4 74.6672
R1852 a_6500_6300.n9 a_6500_6300.n8 74.6672
R1853 a_6500_6300.n1 a_6500_6300.t1 60.0005
R1854 a_6500_6300.n1 a_6500_6300.t3 60.0005
R1855 a_6500_6300.t5 a_6500_6300.n2 60.0005
R1856 a_6500_6300.n2 a_6500_6300.t0 60.0005
R1857 a_6500_6300.n0 a_6500_6300.t2 60.0005
R1858 a_6500_6300.n0 a_6500_6300.t7 60.0005
R1859 a_6500_6300.n8 a_6500_6300.n7 37.763
R1860 a_6500_6300.n5 a_6500_6300.t11 24.0005
R1861 a_6500_6300.n5 a_6500_6300.t9 24.0005
R1862 a_6500_6300.n6 a_6500_6300.t10 24.0005
R1863 a_6500_6300.n6 a_6500_6300.t12 24.0005
R1864 a_6500_6300.n4 a_6500_6300.n3 16.0005
R1865 a_6500_6300.n10 a_6500_6300.n9 16.0005
R1866 pfd_8_0.DOWN_PFD_b.t1 pfd_8_0.DOWN_PFD_b.n1 203.528
R1867 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t2 203.528
R1868 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.t0 183.935
R1869 pfd_8_0.DOWN_PFD_b.n0 pfd_8_0.DOWN_PFD_b.t3 183.935
R1870 pfd_8_0.DOWN_PFD_b.n1 pfd_8_0.DOWN_PFD_b.n0 83.2005
R1871 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t5 1028.27
R1872 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.n1 569.734
R1873 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.n0 465.933
R1874 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t3 401.668
R1875 pfd_8_0.DOWN_b.n0 pfd_8_0.DOWN_b.t4 385.601
R1876 pfd_8_0.DOWN_b.n1 pfd_8_0.DOWN_b.t2 385.601
R1877 pfd_8_0.DOWN_b.t0 pfd_8_0.DOWN_b.n2 211.847
R1878 pfd_8_0.DOWN_b.n2 pfd_8_0.DOWN_b.t1 173.055
R1879 pfd_8_0.QA_b.t4 pfd_8_0.QA_b.t6 1188.93
R1880 pfd_8_0.QA_b pfd_8_0.QA_b.n2 837.38
R1881 pfd_8_0.QA_b.t6 pfd_8_0.QA_b.t3 835.467
R1882 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t5 562.333
R1883 pfd_8_0.QA_b pfd_8_0.QA_b.n0 482
R1884 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.n1 247.917
R1885 pfd_8_0.QA_b.n0 pfd_8_0.QA_b.t4 224.934
R1886 pfd_8_0.QA_b.n2 pfd_8_0.QA_b.t2 221.411
R1887 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t1 24.0005
R1888 pfd_8_0.QA_b.n1 pfd_8_0.QA_b.t0 24.0005
R1889 a_870_1400.t0 a_870_1400.t1 39.4005
R1890 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.t8 918.318
R1891 opamp_cell_4_0.p_bias opamp_cell_4_0.p_bias.n11 540.801
R1892 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t9 377.567
R1893 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t12 377.567
R1894 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.n8 257.067
R1895 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.n6 257.067
R1896 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.n3 257.067
R1897 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n0 154.321
R1898 opamp_cell_4_0.p_bias.n2 opamp_cell_4_0.p_bias.n1 154.321
R1899 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n2 152
R1900 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n10 152
R1901 opamp_cell_4_0.p_bias.n8 opamp_cell_4_0.p_bias.t11 120.501
R1902 opamp_cell_4_0.p_bias.n9 opamp_cell_4_0.p_bias.t6 120.501
R1903 opamp_cell_4_0.p_bias.n7 opamp_cell_4_0.p_bias.t2 120.501
R1904 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.t4 120.501
R1905 opamp_cell_4_0.p_bias.n3 opamp_cell_4_0.p_bias.t10 120.501
R1906 opamp_cell_4_0.p_bias.n4 opamp_cell_4_0.p_bias.t0 120.501
R1907 opamp_cell_4_0.p_bias.n11 opamp_cell_4_0.p_bias.n2 115.201
R1908 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n9 85.6894
R1909 opamp_cell_4_0.p_bias.n10 opamp_cell_4_0.p_bias.n7 85.6894
R1910 opamp_cell_4_0.p_bias.n6 opamp_cell_4_0.p_bias.n5 85.6894
R1911 opamp_cell_4_0.p_bias.n5 opamp_cell_4_0.p_bias.n4 85.6894
R1912 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t3 19.7005
R1913 opamp_cell_4_0.p_bias.n0 opamp_cell_4_0.p_bias.t7 19.7005
R1914 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t1 19.7005
R1915 opamp_cell_4_0.p_bias.n1 opamp_cell_4_0.p_bias.t5 19.7005
R1916 a_6150_5090.n8 a_6150_5090.n6 522.322
R1917 a_6150_5090.n3 a_6150_5090.t0 384.967
R1918 a_6150_5090.n0 a_6150_5090.t3 384.967
R1919 a_6150_5090.n3 a_6150_5090.t2 379.166
R1920 a_6150_5090.t4 a_6150_5090.n0 376.56
R1921 a_6150_5090.n5 a_6150_5090.n1 315.647
R1922 a_6150_5090.n4 a_6150_5090.n2 315.647
R1923 a_6150_5090.n11 a_6150_5090.n10 314.502
R1924 a_6150_5090.n8 a_6150_5090.n7 160.721
R1925 a_6150_5090.n5 a_6150_5090.n4 83.2005
R1926 a_6150_5090.n1 a_6150_5090.t9 49.2505
R1927 a_6150_5090.n1 a_6150_5090.t11 49.2505
R1928 a_6150_5090.n2 a_6150_5090.t10 49.2505
R1929 a_6150_5090.n2 a_6150_5090.t1 49.2505
R1930 a_6150_5090.t4 a_6150_5090.n11 49.2505
R1931 a_6150_5090.n11 a_6150_5090.t12 49.2505
R1932 a_6150_5090.n10 a_6150_5090.n9 42.6672
R1933 a_6150_5090.n9 a_6150_5090.n8 37.763
R1934 a_6150_5090.n9 a_6150_5090.n5 23.4672
R1935 a_6150_5090.n6 a_6150_5090.t5 19.7005
R1936 a_6150_5090.n6 a_6150_5090.t7 19.7005
R1937 a_6150_5090.n7 a_6150_5090.t6 19.7005
R1938 a_6150_5090.n7 a_6150_5090.t8 19.7005
R1939 a_6150_5090.n4 a_6150_5090.n3 16.0005
R1940 a_6150_5090.n10 a_6150_5090.n0 16.0005
R1941 pfd_8_0.DOWN.t3 pfd_8_0.DOWN.n0 605.311
R1942 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN.t3 398.807
R1943 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t1 240.327
R1944 pfd_8_0.DOWN.n0 pfd_8_0.DOWN.t0 148.736
R1945 charge_pump_cell_6_0.DOWN pfd_8_0.DOWN.t2 12.0821
R1946 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.t5 326.658
R1947 pfd_8_0.UP_input.n4 pfd_8_0.UP_input.t4 297.233
R1948 pfd_8_0.UP_input.t3 pfd_8_0.UP_input.n5 297.233
R1949 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.n1 257.067
R1950 pfd_8_0.UP_input.n0 pfd_8_0.UP_input.t2 241.928
R1951 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.n1 226.942
R1952 pfd_8_0.UP_input.n3 pfd_8_0.UP_input.n2 226.942
R1953 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.n6 225.417
R1954 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.n4 216.9
R1955 pfd_8_0.UP_input.t0 pfd_8_0.UP_input.n7 209.928
R1956 pfd_8_0.UP_input.n0 pfd_8_0.UP_input.t1 145.536
R1957 pfd_8_0.UP_input.n7 pfd_8_0.UP_input.n0 144
R1958 pfd_8_0.UP_input.n2 pfd_8_0.UP_input.t4 92.3838
R1959 pfd_8_0.UP_input.n6 pfd_8_0.UP_input.t3 92.3838
R1960 pfd_8_0.UP_input.n4 pfd_8_0.UP_input.t6 80.3338
R1961 pfd_8_0.UP_input.t6 pfd_8_0.UP_input.n3 80.3338
R1962 pfd_8_0.UP_input.n5 pfd_8_0.UP_input.t7 80.3338
R1963 pfd_8_0.UP_input.t7 pfd_8_0.UP_input.n1 80.3338
R1964 V_OUT.n2 V_OUT.n1 2008.33
R1965 V_OUT.n10 V_OUT 1614.79
R1966 V_OUT V_OUT.n2 618.567
R1967 V_OUT.n0 V_OUT.t8 401.668
R1968 V_OUT.n2 V_OUT.n0 369.534
R1969 V_OUT.n1 V_OUT.t10 321.334
R1970 V_OUT.n5 V_OUT.n4 242.903
R1971 V_OUT.n0 V_OUT.t9 192.8
R1972 V_OUT.n5 V_OUT.n3 172.502
R1973 V_OUT.n9 V_OUT.t0 164.118
R1974 V_OUT.n10 V_OUT.n7 113.178
R1975 V_OUT.n1 V_OUT.t11 112.468
R1976 V_OUT.n7 V_OUT.n6 106.662
R1977 V_OUT.n3 V_OUT.t3 24.6255
R1978 V_OUT.n3 V_OUT.t2 24.6255
R1979 V_OUT.n4 V_OUT.t1 24.6255
R1980 V_OUT.n4 V_OUT.t4 24.6255
R1981 V_OUT.n7 V_OUT.n5 19.2005
R1982 V_OUT.n6 V_OUT.t5 15.0005
R1983 V_OUT.n6 V_OUT.t6 15.0005
R1984 V_OUT.n9 V_OUT.t7 8.246
R1985 V_OUT.n10 V_OUT.n9 1.4505
R1986 V_OUT V_OUT.n10 0.063
R1987 V_OUT.n10 V_OUT.n8 0.063
R1988 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.n0 481.334
R1989 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t4 465.933
R1990 pfd_8_0.before_Reset.n0 pfd_8_0.before_Reset.t3 321.334
R1991 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.n1 226.889
R1992 pfd_8_0.before_Reset.n1 pfd_8_0.before_Reset.t1 172.458
R1993 pfd_8_0.before_Reset.n2 pfd_8_0.before_Reset.t2 19.7005
R1994 pfd_8_0.before_Reset.t0 pfd_8_0.before_Reset.n2 19.7005
R1995 a_2350_1400.t1 a_2350_1400.n2 500.086
R1996 a_2350_1400.n1 a_2350_1400.n0 473.334
R1997 a_2350_1400.n0 a_2350_1400.t3 465.933
R1998 a_2350_1400.t1 a_2350_1400.n2 461.389
R1999 a_2350_1400.n0 a_2350_1400.t2 321.334
R2000 a_2350_1400.n1 a_2350_1400.t0 177.577
R2001 a_2350_1400.n2 a_2350_1400.n1 48.3899
R2002 F_REF.n0 F_REF.t0 514.134
R2003 F_REF.n0 F_REF.t1 273.134
R2004 F_REF F_REF.n0 216.9
R2005 a_n30_1400.t0 a_n30_1400.t1 39.4005
R2006 a_6670_5090.t0 a_6670_5090.n6 1112.76
R2007 a_6670_5090.n3 a_6670_5090.n2 416.863
R2008 a_6670_5090.n2 a_6670_5090.n1 366.848
R2009 a_6670_5090.n2 a_6670_5090.n0 271.401
R2010 a_6670_5090.n3 a_6670_5090.t5 208.868
R2011 a_6670_5090.n6 a_6670_5090.t7 208.868
R2012 a_6670_5090.n5 a_6670_5090.t6 208.868
R2013 a_6670_5090.n4 a_6670_5090.t8 208.868
R2014 a_6670_5090.n6 a_6670_5090.n5 208.868
R2015 a_6670_5090.n5 a_6670_5090.n4 208.868
R2016 a_6670_5090.n4 a_6670_5090.n3 193.804
R2017 a_6670_5090.n0 a_6670_5090.t4 60.0005
R2018 a_6670_5090.n0 a_6670_5090.t3 60.0005
R2019 a_6670_5090.n1 a_6670_5090.t2 49.2505
R2020 a_6670_5090.n1 a_6670_5090.t1 49.2505
R2021 pfd_8_0.QA.t5 pfd_8_0.QA.t7 835.467
R2022 pfd_8_0.QA.n2 pfd_8_0.QA.t4 517.347
R2023 pfd_8_0.QA.n0 pfd_8_0.QA.t8 465.933
R2024 pfd_8_0.QA.n1 pfd_8_0.QA.n0 454.031
R2025 pfd_8_0.QA.n1 pfd_8_0.QA.t5 394.267
R2026 pfd_8_0.QA.n0 pfd_8_0.QA.t6 321.334
R2027 pfd_8_0.QA.n4 pfd_8_0.QA.n3 244.715
R2028 pfd_8_0.QA.n2 pfd_8_0.QA.t3 228.148
R2029 pfd_8_0.QA.n4 pfd_8_0.QA.t1 221.411
R2030 pfd_8_0.QA.n5 pfd_8_0.QA.n2 216
R2031 pfd_8_0.QA.n5 pfd_8_0.QA.n4 201.573
R2032 pfd_8_0.QA pfd_8_0.QA.n5 60.8005
R2033 pfd_8_0.QA pfd_8_0.QA.n1 56.1505
R2034 pfd_8_0.QA.n3 pfd_8_0.QA.t0 24.0005
R2035 pfd_8_0.QA.n3 pfd_8_0.QA.t2 24.0005
R2036 I_IN.n2 I_IN.n1 1269.42
R2037 I_IN I_IN.n5 589.356
R2038 I_IN.n2 I_IN.t2 275.325
R2039 I_IN.n4 I_IN.n3 248.4
R2040 I_IN.n5 I_IN.t1 238.892
R2041 I_IN I_IN.n4 214.4
R2042 I_IN.n5 I_IN.t0 161.371
R2043 I_IN.n1 I_IN.t6 151.792
R2044 I_IN.n3 I_IN.t4 140.583
R2045 I_IN.n3 I_IN.t2 140.583
R2046 I_IN.n4 I_IN.n0 98.6614
R2047 I_IN.t4 I_IN.n2 80.3338
R2048 I_IN.n1 I_IN.t7 44.2902
R2049 I_IN.n0 I_IN.t5 15.0005
R2050 I_IN.n0 I_IN.t3 15.0005
R2051 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n1 539.794
R2052 pfd_8_0.DOWN_input.t3 pfd_8_0.DOWN_input.t4 377.567
R2053 pfd_8_0.DOWN_input.n0 pfd_8_0.DOWN_input.t5 326.658
R2054 pfd_8_0.DOWN_input.n2 pfd_8_0.DOWN_input.t0 229.127
R2055 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.n0 196.817
R2056 pfd_8_0.DOWN_input.n2 pfd_8_0.DOWN_input.t2 158.335
R2057 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.t1 158.335
R2058 pfd_8_0.DOWN_input.n3 pfd_8_0.DOWN_input.n2 124.8
R2059 pfd_8_0.DOWN_input.t4 pfd_8_0.DOWN_input.n0 92.3838
R2060 pfd_8_0.DOWN_input.n1 pfd_8_0.DOWN_input.t3 92.3838
R2061 pfd_8_0.DOWN_input pfd_8_0.DOWN_input.n3 6.4005
R2062 pfd_8_0.QB.t4 pfd_8_0.QB.t3 835.467
R2063 pfd_8_0.QB.n1 pfd_8_0.QB.t4 564.496
R2064 pfd_8_0.QB.n2 pfd_8_0.QB.t5 517.347
R2065 pfd_8_0.QB.n0 pfd_8_0.QB.t7 514.134
R2066 pfd_8_0.QB.n1 pfd_8_0.QB.n0 455.219
R2067 pfd_8_0.QB.n5 pfd_8_0.QB.n2 363.2
R2068 pfd_8_0.QB.n0 pfd_8_0.QB.t8 273.134
R2069 pfd_8_0.QB.n4 pfd_8_0.QB.n3 244.716
R2070 pfd_8_0.QB.n2 pfd_8_0.QB.t6 228.148
R2071 pfd_8_0.QB.n4 pfd_8_0.QB.t1 221.411
R2072 pfd_8_0.QB.n5 pfd_8_0.QB.n4 54.3734
R2073 pfd_8_0.QB pfd_8_0.QB.n1 26.7568
R2074 pfd_8_0.QB.n3 pfd_8_0.QB.t0 24.0005
R2075 pfd_8_0.QB.n3 pfd_8_0.QB.t2 24.0005
R2076 pfd_8_0.QB pfd_8_0.QB.n5 6.4005
R2077 a_1910_2020.t0 a_1910_2020.t1 48.0005
R2078 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t2 441.834
R2079 pfd_8_0.UP_PFD_b.n0 pfd_8_0.UP_PFD_b.t3 313.3
R2080 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.n0 235.201
R2081 pfd_8_0.UP_PFD_b.t1 pfd_8_0.UP_PFD_b.n1 219.528
R2082 pfd_8_0.UP_PFD_b.n1 pfd_8_0.UP_PFD_b.t0 167.935
R2083 pfd_8_0.UP.n0 pfd_8_0.UP.t5 1205
R2084 pfd_8_0.UP.n2 pfd_8_0.UP.t4 522.168
R2085 pfd_8_0.UP.n1 pfd_8_0.UP.n0 441.834
R2086 pfd_8_0.UP.n3 pfd_8_0.UP.n2 235.201
R2087 pfd_8_0.UP.t1 pfd_8_0.UP.n3 229.127
R2088 pfd_8_0.UP.n1 pfd_8_0.UP.t3 217.905
R2089 pfd_8_0.UP.n0 pfd_8_0.UP.t2 208.868
R2090 pfd_8_0.UP.n3 pfd_8_0.UP.t0 158.335
R2091 pfd_8_0.UP.n2 pfd_8_0.UP.n1 15.063
R2092 a_9540_3974.t0 a_9540_3974.t1 323.964
R2093 pfd_8_0.E.n4 pfd_8_0.E.n0 1319.38
R2094 pfd_8_0.E.n0 pfd_8_0.E.t3 562.333
R2095 pfd_8_0.E.n2 pfd_8_0.E.t5 388.813
R2096 pfd_8_0.E.n2 pfd_8_0.E.t4 356.68
R2097 pfd_8_0.E.n3 pfd_8_0.E.n2 232
R2098 pfd_8_0.E.n0 pfd_8_0.E.t6 224.934
R2099 pfd_8_0.E.t1 pfd_8_0.E.n4 221.411
R2100 pfd_8_0.E.n3 pfd_8_0.E.n1 157.278
R2101 pfd_8_0.E.n4 pfd_8_0.E.n3 90.64
R2102 pfd_8_0.E.n1 pfd_8_0.E.t0 24.0005
R2103 pfd_8_0.E.n1 pfd_8_0.E.t2 24.0005
R2104 pfd_8_0.E_b.n0 pfd_8_0.E_b.t4 517.347
R2105 pfd_8_0.E_b.n2 pfd_8_0.E_b.n0 417.574
R2106 pfd_8_0.E_b.n2 pfd_8_0.E_b.n1 244.716
R2107 pfd_8_0.E_b.n0 pfd_8_0.E_b.t3 228.148
R2108 pfd_8_0.E_b.t1 pfd_8_0.E_b.n2 221.411
R2109 pfd_8_0.E_b.n1 pfd_8_0.E_b.t0 24.0005
R2110 pfd_8_0.E_b.n1 pfd_8_0.E_b.t2 24.0005
R2111 a_1390_1400.t0 a_1390_1400.t1 39.4005
R2112 pfd_8_0.QB_b.t6 pfd_8_0.QB_b.t4 1188.93
R2113 pfd_8_0.QB_b pfd_8_0.QB_b.n2 899.734
R2114 pfd_8_0.QB_b.t4 pfd_8_0.QB_b.t3 835.467
R2115 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t5 562.333
R2116 pfd_8_0.QB_b pfd_8_0.QB_b.n1 419.647
R2117 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.n0 247.917
R2118 pfd_8_0.QB_b.n2 pfd_8_0.QB_b.t6 224.934
R2119 pfd_8_0.QB_b.n1 pfd_8_0.QB_b.t0 221.411
R2120 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t1 24.0005
R2121 pfd_8_0.QB_b.n0 pfd_8_0.QB_b.t2 24.0005
R2122 a_870_640.t0 a_870_640.t1 39.4005
R2123 a_2530_190.t1 a_2530_190.n2 500.086
R2124 a_2530_190.n0 a_2530_190.t2 465.933
R2125 a_2530_190.t1 a_2530_190.n2 461.389
R2126 a_2530_190.n1 a_2530_190.n0 392.623
R2127 a_2530_190.n0 a_2530_190.t3 321.334
R2128 a_2530_190.n1 a_2530_190.t0 177.577
R2129 a_2530_190.n2 a_2530_190.n1 48.3899
R2130 a_2200_190.t1 a_2200_190.n2 500.086
R2131 a_2200_190.n1 a_2200_190.n0 473.334
R2132 a_2200_190.n0 a_2200_190.t2 465.933
R2133 a_2200_190.t1 a_2200_190.n2 461.389
R2134 a_2200_190.n0 a_2200_190.t3 321.334
R2135 a_2200_190.n1 a_2200_190.t0 177.577
R2136 a_2200_190.n2 a_2200_190.n1 48.3898
R2137 pfd_8_0.F.n4 pfd_8_0.F.n0 1319.38
R2138 pfd_8_0.F.n0 pfd_8_0.F.t3 562.333
R2139 pfd_8_0.F.n2 pfd_8_0.F.t5 388.813
R2140 pfd_8_0.F.n2 pfd_8_0.F.t6 356.68
R2141 pfd_8_0.F.n3 pfd_8_0.F.n2 232
R2142 pfd_8_0.F.n0 pfd_8_0.F.t4 224.934
R2143 pfd_8_0.F.t2 pfd_8_0.F.n4 221.411
R2144 pfd_8_0.F.n3 pfd_8_0.F.n1 157.278
R2145 pfd_8_0.F.n4 pfd_8_0.F.n3 90.64
R2146 pfd_8_0.F.n1 pfd_8_0.F.t0 24.0005
R2147 pfd_8_0.F.n1 pfd_8_0.F.t1 24.0005
R2148 charge_pump_cell_6_0.UP_b pfd_8_0.UP_b.n1 485.846
R2149 pfd_8_0.UP_b.n1 pfd_8_0.UP_b.n0 409.067
R2150 pfd_8_0.UP_b.n1 pfd_8_0.UP_b.t3 369.534
R2151 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t1 209.928
R2152 pfd_8_0.UP_b.n0 pfd_8_0.UP_b.t0 177.536
R2153 charge_pump_cell_6_0.UP_b pfd_8_0.UP_b.t2 12.0774
R2154 pfd_8_0.F_b.n0 pfd_8_0.F_b.t3 517.347
R2155 pfd_8_0.F_b.n2 pfd_8_0.F_b.n0 417.574
R2156 pfd_8_0.F_b.n2 pfd_8_0.F_b.n1 244.716
R2157 pfd_8_0.F_b.n0 pfd_8_0.F_b.t4 228.148
R2158 pfd_8_0.F_b.t1 pfd_8_0.F_b.n2 221.411
R2159 pfd_8_0.F_b.n1 pfd_8_0.F_b.t0 24.0005
R2160 pfd_8_0.F_b.n1 pfd_8_0.F_b.t2 24.0005
R2161 a_1390_640.t0 a_1390_640.t1 39.4005
R2162 a_490_640.t0 a_490_640.t1 39.4005
R2163 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n7 933.13
R2164 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t8 377.567
R2165 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t9 297.233
R2166 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n1 243.44
R2167 opamp_cell_4_0.VIN+.n2 opamp_cell_4_0.VIN+.n0 224.496
R2168 opamp_cell_4_0.VIN+.n0 opamp_cell_4_0.VIN+.t7 216.9
R2169 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.n4 196.262
R2170 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n3 172.502
R2171 opamp_cell_4_0.VIN+.n6 opamp_cell_4_0.VIN+.n5 172.5
R2172 opamp_cell_4_0.VIN+.n1 opamp_cell_4_0.VIN+.t6 136.567
R2173 opamp_cell_4_0.VIN+.n7 opamp_cell_4_0.VIN+.n6 70.4005
R2174 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t2 24.6255
R2175 opamp_cell_4_0.VIN+.n3 opamp_cell_4_0.VIN+.t1 24.6255
R2176 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.t0 24.6255
R2177 opamp_cell_4_0.VIN+.n5 opamp_cell_4_0.VIN+.t3 24.6255
R2178 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t5 15.0005
R2179 opamp_cell_4_0.VIN+.n4 opamp_cell_4_0.VIN+.t4 15.0005
R2180 opamp_cell_4_0.VIN+ opamp_cell_4_0.VIN+.n2 3.438
R2181 a_490_1400.t0 a_490_1400.t1 39.4005
R2182 pfd_8_0.Reset.n1 pfd_8_0.Reset.t3 562.333
R2183 pfd_8_0.Reset.n2 pfd_8_0.Reset.n1 480.45
R2184 pfd_8_0.Reset.n0 pfd_8_0.Reset.t4 417.733
R2185 pfd_8_0.Reset.n0 pfd_8_0.Reset.t5 369.534
R2186 pfd_8_0.Reset.n3 pfd_8_0.Reset.n2 328.733
R2187 pfd_8_0.Reset.t1 pfd_8_0.Reset.n3 288.37
R2188 pfd_8_0.Reset.n1 pfd_8_0.Reset.t2 224.934
R2189 pfd_8_0.Reset.n3 pfd_8_0.Reset.t0 177.577
R2190 pfd_8_0.Reset.n2 pfd_8_0.Reset.n0 176.733
R2191 a_1870_190.t1 a_1870_190.n2 500.086
R2192 a_1870_190.n1 a_1870_190.n0 473.334
R2193 a_1870_190.n0 a_1870_190.t2 465.933
R2194 a_1870_190.t1 a_1870_190.n2 461.389
R2195 a_1870_190.n0 a_1870_190.t3 321.334
R2196 a_1870_190.n1 a_1870_190.t0 177.577
R2197 a_1870_190.n2 a_1870_190.n1 48.3898
R2198 loop_filter_2_0.R1_C1.t0 loop_filter_2_0.R1_C1.t1 167.429
R2199 a_9540_6900.t0 a_9540_6900.t1 245.883
R2200 a_n30_640.t0 a_n30_640.t1 39.4005
R2201 F_VCO.n0 F_VCO.t0 514.134
R2202 F_VCO.n0 F_VCO.t1 273.134
R2203 F_VCO F_VCO.n0 216.9
C0 pfd_8_0.DOWN_input I_IN 0.581394f
C1 F_REF pfd_8_0.QA_b 0.027208f
C2 VDDA opamp_cell_4_0.p_bias 3.3163f
C3 pfd_8_0.DOWN_input opamp_cell_4_0.VIN+ 0.132099f
C4 opamp_cell_4_0.VIN+ V_OUT 1.18544f
C5 opamp_cell_4_0.VIN+ I_IN 0.544835f
C6 VDDA pfd_8_0.QA_b 0.52066f
C7 opamp_cell_4_0.p_bias V_OUT 0.049138f
C8 pfd_8_0.QB_b F_VCO 0.027208f
C9 F_REF pfd_8_0.QA 0.056f
C10 F_VCO pfd_8_0.QB 0.056153f
C11 pfd_8_0.QA pfd_8_0.QB 0.074487f
C12 opamp_cell_4_0.VIN+ opamp_cell_4_0.p_bias 0.498662f
C13 VDDA F_VCO 0.098386f
C14 VDDA pfd_8_0.QA 0.550605f
C15 pfd_8_0.QB_b pfd_8_0.QB 0.388258f
C16 VDDA F_REF 0.098433f
C17 VDDA pfd_8_0.QB_b 0.511838f
C18 VDDA pfd_8_0.QB 2.74984f
C19 VDDA pfd_8_0.DOWN_input 0.168412f
C20 VDDA V_OUT 1.44907f
C21 pfd_8_0.QA_b pfd_8_0.QA 0.422694f
C22 VDDA I_IN 0.452819f
C23 VDDA opamp_cell_4_0.VIN+ 1.06587f
C24 pfd_8_0.DOWN_input V_OUT 0.406052f
C25 I_IN GNDA 3.05246f
C26 F_VCO GNDA 0.277756f
C27 F_REF GNDA 0.277756f
C28 V_OUT GNDA 26.45354f
C29 VDDA GNDA 65.93004f
C30 pfd_8_0.DOWN_input GNDA 3.21297f
C31 pfd_8_0.QB_b GNDA 1.06334f
C32 pfd_8_0.QB GNDA 1.3083f
C33 pfd_8_0.QA GNDA 3.10074f
C34 pfd_8_0.QA_b GNDA 1.05138f
C35 opamp_cell_4_0.VIN+ GNDA 2.71146f
C36 opamp_cell_4_0.p_bias GNDA 3.153184f
C37 loop_filter_2_0.R1_C1.t1 GNDA 2.39887f
C38 pfd_8_0.QB.t7 GNDA 0.066708f
C39 pfd_8_0.QB.t8 GNDA 0.031333f
C40 pfd_8_0.QB.n0 GNDA 0.096363f
C41 pfd_8_0.QB.t3 GNDA 0.066708f
C42 pfd_8_0.QB.t4 GNDA 0.100569f
C43 pfd_8_0.QB.n1 GNDA 1.20598f
C44 pfd_8_0.QB.t5 GNDA 0.067367f
C45 pfd_8_0.QB.t6 GNDA 0.029539f
C46 pfd_8_0.QB.n2 GNDA 0.170164f
C47 pfd_8_0.QB.t1 GNDA 0.14186f
C48 pfd_8_0.QB.t0 GNDA 0.026953f
C49 pfd_8_0.QB.t2 GNDA 0.026953f
C50 pfd_8_0.QB.n3 GNDA 0.143916f
C51 pfd_8_0.QB.n4 GNDA 0.255686f
C52 pfd_8_0.QB.n5 GNDA 0.218372f
C53 V_OUT.t7 GNDA 2.24688f
C54 V_OUT.n9 GNDA 0.049845f
C55 V_OUT.n10 GNDA 0.069037f
C56 pfd_8_0.UP_input.t1 GNDA 0.019943f
C57 pfd_8_0.UP_input.t2 GNDA 0.048355f
C58 pfd_8_0.UP_input.n0 GNDA 0.059297f
C59 pfd_8_0.UP_input.n1 GNDA 0.022544f
C60 pfd_8_0.UP_input.t7 GNDA 0.024945f
C61 pfd_8_0.UP_input.t4 GNDA 0.042895f
C62 pfd_8_0.UP_input.t5 GNDA 1.97861f
C63 pfd_8_0.UP_input.n2 GNDA 0.043722f
C64 pfd_8_0.UP_input.n3 GNDA 0.022544f
C65 pfd_8_0.UP_input.t6 GNDA 0.024945f
C66 pfd_8_0.UP_input.n4 GNDA 0.030069f
C67 pfd_8_0.UP_input.n5 GNDA 0.030069f
C68 pfd_8_0.UP_input.t3 GNDA 0.042895f
C69 pfd_8_0.UP_input.n6 GNDA 0.039471f
C70 pfd_8_0.UP_input.n7 GNDA 0.22578f
C71 pfd_8_0.UP_input.t0 GNDA 0.043912f
C72 a_6150_5090.t3 GNDA 0.030769f
C73 a_6150_5090.n0 GNDA 0.124795f
C74 a_6150_5090.t12 GNDA 0.020325f
C75 a_6150_5090.t9 GNDA 0.020325f
C76 a_6150_5090.t11 GNDA 0.020325f
C77 a_6150_5090.n1 GNDA 0.044943f
C78 a_6150_5090.t10 GNDA 0.020325f
C79 a_6150_5090.t1 GNDA 0.020325f
C80 a_6150_5090.n2 GNDA 0.044943f
C81 a_6150_5090.t2 GNDA 0.077457f
C82 a_6150_5090.t0 GNDA 0.030769f
C83 a_6150_5090.n3 GNDA 0.097952f
C84 a_6150_5090.n4 GNDA 0.087903f
C85 a_6150_5090.n5 GNDA 0.089425f
C86 a_6150_5090.t5 GNDA 0.050813f
C87 a_6150_5090.t7 GNDA 0.050813f
C88 a_6150_5090.n6 GNDA 0.295522f
C89 a_6150_5090.t6 GNDA 0.050813f
C90 a_6150_5090.t8 GNDA 0.050813f
C91 a_6150_5090.n7 GNDA 0.144587f
C92 a_6150_5090.n8 GNDA 0.360746f
C93 a_6150_5090.n9 GNDA 0.13437f
C94 a_6150_5090.n10 GNDA 0.085474f
C95 a_6150_5090.n11 GNDA 0.045257f
C96 a_6150_5090.t4 GNDA 0.100208f
C97 opamp_cell_4_0.p_bias.t8 GNDA 1.892f
C98 opamp_cell_4_0.p_bias.t3 GNDA 0.022409f
C99 opamp_cell_4_0.p_bias.t7 GNDA 0.022409f
C100 opamp_cell_4_0.p_bias.n0 GNDA 0.061525f
C101 opamp_cell_4_0.p_bias.t1 GNDA 0.022409f
C102 opamp_cell_4_0.p_bias.t5 GNDA 0.022409f
C103 opamp_cell_4_0.p_bias.n1 GNDA 0.061525f
C104 opamp_cell_4_0.p_bias.n2 GNDA 0.07795f
C105 opamp_cell_4_0.p_bias.t2 GNDA 0.061849f
C106 opamp_cell_4_0.p_bias.t4 GNDA 0.061849f
C107 opamp_cell_4_0.p_bias.t0 GNDA 0.061849f
C108 opamp_cell_4_0.p_bias.t10 GNDA 0.061849f
C109 opamp_cell_4_0.p_bias.t12 GNDA 0.085041f
C110 opamp_cell_4_0.p_bias.n3 GNDA 0.047622f
C111 opamp_cell_4_0.p_bias.n4 GNDA 0.033793f
C112 opamp_cell_4_0.p_bias.n5 GNDA 0.014521f
C113 opamp_cell_4_0.p_bias.n6 GNDA 0.033793f
C114 opamp_cell_4_0.p_bias.n7 GNDA 0.033793f
C115 opamp_cell_4_0.p_bias.t6 GNDA 0.061849f
C116 opamp_cell_4_0.p_bias.t11 GNDA 0.061849f
C117 opamp_cell_4_0.p_bias.t9 GNDA 0.085041f
C118 opamp_cell_4_0.p_bias.n8 GNDA 0.047622f
C119 opamp_cell_4_0.p_bias.n9 GNDA 0.033793f
C120 opamp_cell_4_0.p_bias.n10 GNDA 0.014521f
C121 opamp_cell_4_0.p_bias.n11 GNDA 0.137263f
C122 pfd_8_0.opamp_out.t13 GNDA 0.016624f
C123 pfd_8_0.opamp_out.n0 GNDA 0.012184f
C124 pfd_8_0.opamp_out.t14 GNDA 0.02314f
C125 pfd_8_0.opamp_out.t11 GNDA 0.010108f
C126 pfd_8_0.opamp_out.n1 GNDA 0.012184f
C127 pfd_8_0.opamp_out.n2 GNDA 0.012184f
C128 pfd_8_0.opamp_out.t12 GNDA 0.010108f
C129 pfd_8_0.opamp_out.n4 GNDA 0.01577f
C130 pfd_8_0.opamp_out.t5 GNDA 0.021617f
C131 pfd_8_0.opamp_out.n5 GNDA 0.039426f
C132 pfd_8_0.opamp_out.n6 GNDA 0.150316f
C133 pfd_8_0.opamp_out.t15 GNDA 1.72189f
C134 pfd_8_0.opamp_out.n9 GNDA 0.017323f
C135 pfd_8_0.opamp_out.n10 GNDA 0.014909f
C136 pfd_8_0.opamp_out.t10 GNDA 1.72116f
C137 pfd_8_0.opamp_out.n13 GNDA 0.023291f
C138 pfd_8_0.opamp_out.n14 GNDA 0.015404f
C139 opamp_cell_4_0.VOUT GNDA 0.10585f
C140 VDDA.n1 GNDA 0.010245f
C141 VDDA.n2 GNDA 0.010245f
C142 VDDA.n13 GNDA 0.010245f
C143 VDDA.n14 GNDA 0.010245f
C144 VDDA.n20 GNDA 0.062647f
C145 VDDA.t22 GNDA 0.015729f
C146 VDDA.n23 GNDA 0.017227f
C147 VDDA.n25 GNDA 0.010245f
C148 VDDA.t119 GNDA 0.010929f
C149 VDDA.n29 GNDA 0.010093f
C150 VDDA.n34 GNDA 0.010245f
C151 VDDA.n37 GNDA 0.010245f
C152 VDDA.n38 GNDA 0.010245f
C153 VDDA.n41 GNDA 0.010995f
C154 VDDA.n42 GNDA 0.010995f
C155 VDDA.n45 GNDA 0.010995f
C156 VDDA.n48 GNDA 0.010995f
C157 VDDA.n50 GNDA 0.015545f
C158 VDDA.t26 GNDA 0.339085f
C159 VDDA.n55 GNDA 0.015545f
C160 VDDA.n56 GNDA 0.035604f
C161 VDDA.n60 GNDA 0.015545f
C162 VDDA.t36 GNDA 0.213486f
C163 VDDA.t98 GNDA 0.025667f
C164 VDDA.n69 GNDA 0.013565f
C165 VDDA.n72 GNDA 0.013565f
C166 VDDA.n75 GNDA 0.013565f
C167 VDDA.n78 GNDA 0.013565f
C168 VDDA.n82 GNDA 0.011205f
C169 VDDA.t3 GNDA 0.122755f
C170 VDDA.n88 GNDA 0.014509f
C171 VDDA.n91 GNDA 0.014509f
C172 VDDA.n94 GNDA 0.014982f
C173 VDDA.n95 GNDA 0.021082f
C174 VDDA.n97 GNDA 0.014982f
C175 VDDA.n98 GNDA 0.021082f
C176 VDDA.n117 GNDA 0.014982f
C177 VDDA.n120 GNDA 0.014982f
C178 VDDA.n122 GNDA 0.013328f
C179 VDDA.t101 GNDA 0.025829f
C180 VDDA.n126 GNDA 0.010158f
C181 VDDA.n130 GNDA 0.068227f
C182 VDDA.t72 GNDA 0.128092f
C183 VDDA.t88 GNDA 0.138766f
C184 VDDA.t74 GNDA 0.085395f
C185 VDDA.t64 GNDA 0.138766f
C186 VDDA.t112 GNDA 0.149441f
C187 VDDA.t47 GNDA 0.122755f
C188 VDDA.t85 GNDA 0.117418f
C189 VDDA.t113 GNDA 0.011882f
C190 VDDA.n134 GNDA 0.023158f
C191 VDDA.n135 GNDA 0.176059f
C192 VDDA.t41 GNDA 0.160115f
C193 VDDA.n136 GNDA 0.053372f
C194 VDDA.t84 GNDA 0.026192f
C195 VDDA.n150 GNDA 0.018302f
C196 VDDA.n151 GNDA 0.019431f
C197 VDDA.t86 GNDA 0.012954f
C198 VDDA.n152 GNDA 0.013565f
C199 VDDA.n154 GNDA 0.046819f
C200 VDDA.n155 GNDA 0.046596f
C201 VDDA.t97 GNDA 0.011911f
C202 VDDA.n158 GNDA 0.011205f
C203 VDDA.n159 GNDA 0.016038f
C204 VDDA.n160 GNDA 0.011205f
C205 VDDA.n162 GNDA 0.019491f
C206 VDDA.n163 GNDA 0.192062f
C207 VDDA.t108 GNDA 0.181463f
C208 VDDA.t43 GNDA 0.138766f
C209 VDDA.t80 GNDA 0.234835f
C210 VDDA.t45 GNDA 0.138766f
C211 VDDA.t82 GNDA 0.176126f
C212 VDDA.t78 GNDA 0.197475f
C213 VDDA.t102 GNDA 0.138766f
C214 VDDA.t76 GNDA 0.218824f
C215 VDDA.t96 GNDA 0.144103f
C216 VDDA.n164 GNDA 0.289573f
C217 VDDA.n169 GNDA 0.015545f
C218 VDDA.t103 GNDA 0.010363f
C219 VDDA.n170 GNDA 0.014982f
C220 VDDA.n171 GNDA 0.02135f
C221 VDDA.n178 GNDA 0.020046f
C222 VDDA.n185 GNDA 0.021082f
C223 VDDA.n193 GNDA 0.021082f
C224 VDDA.n194 GNDA 0.014982f
C225 VDDA.t106 GNDA 0.010363f
C226 VDDA.n195 GNDA 0.015545f
C227 VDDA.t87 GNDA 0.024372f
C228 VDDA.t104 GNDA 0.024372f
C229 VDDA.n197 GNDA 0.01098f
C230 VDDA.n198 GNDA 0.018711f
C231 VDDA.n199 GNDA 0.015545f
C232 VDDA.n200 GNDA 0.017627f
C233 VDDA.n202 GNDA 0.11208f
C234 VDDA.t70 GNDA 0.117418f
C235 VDDA.t37 GNDA 0.138766f
C236 VDDA.t68 GNDA 0.106743f
C237 VDDA.t105 GNDA 0.138766f
C238 VDDA.t115 GNDA 0.106743f
C239 VDDA.t56 GNDA 0.165452f
C240 VDDA.t33 GNDA 0.138766f
C241 VDDA.t92 GNDA 0.138766f
C242 VDDA.t52 GNDA 0.165452f
C243 VDDA.t53 GNDA 0.186801f
C244 VDDA.t62 GNDA 0.069383f
C245 VDDA.t0 GNDA 0.090732f
C246 VDDA.t32 GNDA 0.192138f
C247 VDDA.t58 GNDA 0.138766f
C248 VDDA.t67 GNDA 0.042697f
C249 VDDA.t39 GNDA 0.138766f
C250 VDDA.t35 GNDA 0.170789f
C251 VDDA.t54 GNDA 0.122755f
C252 VDDA.t49 GNDA 0.213486f
C253 VDDA.t60 GNDA 0.224161f
C254 VDDA.n203 GNDA 0.090656f
C255 VDDA.n204 GNDA 0.019491f
C256 VDDA.n206 GNDA 0.011205f
C257 VDDA.n207 GNDA 0.01448f
C258 VDDA.n212 GNDA 0.045403f
C259 VDDA.n219 GNDA 0.045403f
C260 VDDA.n226 GNDA 0.045403f
C261 VDDA.n233 GNDA 0.045403f
C262 VDDA.n246 GNDA 0.019431f
C263 VDDA.n255 GNDA 0.11208f
C264 VDDA.n261 GNDA 0.532116f
C265 VDDA.n263 GNDA 0.010431f
C266 VDDA.t91 GNDA 0.025829f
C267 VDDA.n271 GNDA 0.025615f
C268 VDDA.n272 GNDA 0.256051f
C269 VDDA.n273 GNDA 0.044213f
C270 VDDA.n286 GNDA 0.010995f
C271 VDDA.n293 GNDA 0.125294f
C272 VDDA.t66 GNDA 0.165452f
C273 VDDA.t7 GNDA 0.146176f
C274 VDDA.t11 GNDA 0.043371f
C275 VDDA.t118 GNDA 0.043371f
C276 VDDA.t12 GNDA 0.010929f
C277 VDDA.n302 GNDA 0.010093f
C278 VDDA.n307 GNDA 0.062647f
C279 VDDA.t10 GNDA 0.010929f
C280 VDDA.n313 GNDA 0.010093f
C281 VDDA.n315 GNDA 0.062647f
C282 VDDA.t28 GNDA 0.043371f
C283 VDDA.t9 GNDA 0.043371f
C284 VDDA.t29 GNDA 0.010929f
C285 VDDA.n318 GNDA 0.010093f
C286 VDDA.n323 GNDA 0.088348f
C287 VDDA.n328 GNDA 0.015545f
C288 VDDA.n334 GNDA 0.015545f
C289 VDDA.n341 GNDA 0.136538f
C290 VDDA.t17 GNDA 0.125294f
C291 VDDA.n343 GNDA 0.015545f
C292 VDDA.n350 GNDA 0.125294f
C293 VDDA.t19 GNDA 0.125294f
C294 VDDA.n357 GNDA 0.015545f
C295 VDDA.n364 GNDA 0.125294f
C296 VDDA.n366 GNDA 0.010995f
C297 VDDA.n371 GNDA 0.039908f
C298 VDDA.n407 GNDA 0.010093f
C299 VDDA.t14 GNDA 0.010929f
C300 VDDA.n409 GNDA 0.010245f
C301 VDDA.n411 GNDA 0.062647f
C302 VDDA.t21 GNDA 0.040158f
C303 VDDA.t5 GNDA 0.038552f
C304 VDDA.t13 GNDA 0.043371f
C305 VDDA.t16 GNDA 0.010929f
C306 VDDA.n418 GNDA 0.010093f
C307 VDDA.t30 GNDA 0.010929f
C308 VDDA.n428 GNDA 0.010093f
C309 VDDA.n430 GNDA 0.094773f
C310 VDDA.t15 GNDA 0.07871f
C311 VDDA.t2 GNDA 0.167058f
C312 VDDA.t122 GNDA 0.167058f
C313 VDDA.t125 GNDA 0.07871f
C314 VDDA.n434 GNDA 0.0114f
C315 VDDA.n435 GNDA 0.013644f
C316 VDDA.n438 GNDA 0.0114f
C317 VDDA.t127 GNDA 0.010935f
C318 VDDA.n441 GNDA 0.011364f
C319 VDDA.n445 GNDA 0.0114f
C320 VDDA.n446 GNDA 0.011364f
C321 VDDA.n449 GNDA 0.0114f
C322 VDDA.t124 GNDA 0.010935f
C323 VDDA.n452 GNDA 0.013644f
C324 VDDA.n454 GNDA 0.086742f
C325 VDDA.t123 GNDA 0.07871f
C326 VDDA.t25 GNDA 0.167058f
C327 VDDA.t31 GNDA 0.167058f
C328 VDDA.t23 GNDA 0.07871f
C329 VDDA.t121 GNDA 0.010929f
C330 VDDA.n458 GNDA 0.010093f
C331 VDDA.t24 GNDA 0.010929f
C332 VDDA.n468 GNDA 0.010093f
C333 VDDA.n470 GNDA 0.088348f
C334 VDDA.t6 GNDA 0.010875f
C335 VDDA.n474 GNDA 0.010093f
C336 VDDA.n476 GNDA 0.085135f
C337 VDDA.n478 GNDA 0.010051f
.ends

