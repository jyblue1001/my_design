magic
tech sky130A
timestamp 1746550971
<< nwell >>
rect 2450 1960 4655 2820
<< pwell >>
rect 2710 1560 3750 1660
<< nmos >>
rect 2750 1560 2810 1660
rect 2850 1560 2910 1660
rect 2950 1560 3010 1660
rect 3050 1560 3110 1660
rect 3150 1560 3210 1660
rect 3250 1560 3310 1660
rect 3350 1560 3410 1660
rect 3450 1560 3510 1660
rect 3550 1560 3610 1660
rect 3650 1560 3710 1660
rect 2770 985 3170 1385
rect 3290 985 3690 1385
rect 2720 755 3720 855
<< pmos >>
rect 2550 2400 2610 2800
rect 2650 2400 2710 2800
rect 2750 2400 2810 2800
rect 2850 2400 2910 2800
rect 2950 2400 3010 2800
rect 3050 2400 3110 2800
rect 3150 2400 3210 2800
rect 3250 2400 3310 2800
rect 3350 2400 3410 2800
rect 3450 2400 3510 2800
rect 3550 2400 3610 2800
rect 3650 2400 3710 2800
rect 3750 2400 3810 2800
rect 3850 2400 3910 2800
rect 2550 1980 2610 2180
rect 2650 1980 2710 2180
rect 2750 1980 2810 2180
rect 2850 1980 2910 2180
rect 2950 1980 3010 2180
rect 3050 1980 3110 2180
rect 3150 1980 3210 2180
rect 3250 1980 3310 2180
rect 3350 1980 3410 2180
rect 3450 1980 3510 2180
rect 3550 1980 3610 2180
rect 3650 1980 3710 2180
rect 3750 1980 3810 2180
rect 3850 1980 3910 2180
rect 4415 1980 4430 2180
rect 4540 1980 4555 2180
<< ndiff >>
rect 2710 1645 2750 1660
rect 2710 1625 2720 1645
rect 2740 1625 2750 1645
rect 2710 1595 2750 1625
rect 2710 1575 2720 1595
rect 2740 1575 2750 1595
rect 2710 1560 2750 1575
rect 2810 1645 2850 1660
rect 2810 1625 2820 1645
rect 2840 1625 2850 1645
rect 2810 1595 2850 1625
rect 2810 1575 2820 1595
rect 2840 1575 2850 1595
rect 2810 1560 2850 1575
rect 2910 1645 2950 1660
rect 2910 1625 2920 1645
rect 2940 1625 2950 1645
rect 2910 1595 2950 1625
rect 2910 1575 2920 1595
rect 2940 1575 2950 1595
rect 2910 1560 2950 1575
rect 3010 1645 3050 1660
rect 3010 1625 3020 1645
rect 3040 1625 3050 1645
rect 3010 1595 3050 1625
rect 3010 1575 3020 1595
rect 3040 1575 3050 1595
rect 3010 1560 3050 1575
rect 3110 1645 3150 1660
rect 3110 1625 3120 1645
rect 3140 1625 3150 1645
rect 3110 1595 3150 1625
rect 3110 1575 3120 1595
rect 3140 1575 3150 1595
rect 3110 1560 3150 1575
rect 3210 1645 3250 1660
rect 3210 1625 3220 1645
rect 3240 1625 3250 1645
rect 3210 1595 3250 1625
rect 3210 1575 3220 1595
rect 3240 1575 3250 1595
rect 3210 1560 3250 1575
rect 3310 1645 3350 1660
rect 3310 1625 3320 1645
rect 3340 1625 3350 1645
rect 3310 1595 3350 1625
rect 3310 1575 3320 1595
rect 3340 1575 3350 1595
rect 3310 1560 3350 1575
rect 3410 1645 3450 1660
rect 3410 1625 3420 1645
rect 3440 1625 3450 1645
rect 3410 1595 3450 1625
rect 3410 1575 3420 1595
rect 3440 1575 3450 1595
rect 3410 1560 3450 1575
rect 3510 1645 3550 1660
rect 3510 1625 3520 1645
rect 3540 1625 3550 1645
rect 3510 1595 3550 1625
rect 3510 1575 3520 1595
rect 3540 1575 3550 1595
rect 3510 1560 3550 1575
rect 3610 1645 3650 1660
rect 3610 1625 3620 1645
rect 3640 1625 3650 1645
rect 3610 1595 3650 1625
rect 3610 1575 3620 1595
rect 3640 1575 3650 1595
rect 3610 1560 3650 1575
rect 3710 1645 3750 1660
rect 3710 1625 3720 1645
rect 3740 1625 3750 1645
rect 3710 1595 3750 1625
rect 3710 1575 3720 1595
rect 3740 1575 3750 1595
rect 3710 1560 3750 1575
rect 2730 1370 2770 1385
rect 2730 1350 2740 1370
rect 2760 1350 2770 1370
rect 2730 1320 2770 1350
rect 2730 1300 2740 1320
rect 2760 1300 2770 1320
rect 2730 1270 2770 1300
rect 2730 1250 2740 1270
rect 2760 1250 2770 1270
rect 2730 1220 2770 1250
rect 2730 1200 2740 1220
rect 2760 1200 2770 1220
rect 2730 1170 2770 1200
rect 2730 1150 2740 1170
rect 2760 1150 2770 1170
rect 2730 1120 2770 1150
rect 2730 1100 2740 1120
rect 2760 1100 2770 1120
rect 2730 1070 2770 1100
rect 2730 1050 2740 1070
rect 2760 1050 2770 1070
rect 2730 1020 2770 1050
rect 2730 1000 2740 1020
rect 2760 1000 2770 1020
rect 2730 985 2770 1000
rect 3170 1370 3210 1385
rect 3250 1370 3290 1385
rect 3170 1350 3180 1370
rect 3200 1350 3210 1370
rect 3250 1350 3260 1370
rect 3280 1350 3290 1370
rect 3170 1320 3210 1350
rect 3250 1320 3290 1350
rect 3170 1300 3180 1320
rect 3200 1300 3210 1320
rect 3250 1300 3260 1320
rect 3280 1300 3290 1320
rect 3170 1270 3210 1300
rect 3250 1270 3290 1300
rect 3170 1250 3180 1270
rect 3200 1250 3210 1270
rect 3250 1250 3260 1270
rect 3280 1250 3290 1270
rect 3170 1220 3210 1250
rect 3250 1220 3290 1250
rect 3170 1200 3180 1220
rect 3200 1200 3210 1220
rect 3250 1200 3260 1220
rect 3280 1200 3290 1220
rect 3170 1170 3210 1200
rect 3250 1170 3290 1200
rect 3170 1150 3180 1170
rect 3200 1150 3210 1170
rect 3250 1150 3260 1170
rect 3280 1150 3290 1170
rect 3170 1120 3210 1150
rect 3250 1120 3290 1150
rect 3170 1100 3180 1120
rect 3200 1100 3210 1120
rect 3250 1100 3260 1120
rect 3280 1100 3290 1120
rect 3170 1070 3210 1100
rect 3250 1070 3290 1100
rect 3170 1050 3180 1070
rect 3200 1050 3210 1070
rect 3250 1050 3260 1070
rect 3280 1050 3290 1070
rect 3170 1020 3210 1050
rect 3250 1020 3290 1050
rect 3170 1000 3180 1020
rect 3200 1000 3210 1020
rect 3250 1000 3260 1020
rect 3280 1000 3290 1020
rect 3170 985 3210 1000
rect 3250 985 3290 1000
rect 3690 1370 3730 1385
rect 3690 1350 3700 1370
rect 3720 1350 3730 1370
rect 3690 1320 3730 1350
rect 3690 1300 3700 1320
rect 3720 1300 3730 1320
rect 3690 1270 3730 1300
rect 3690 1250 3700 1270
rect 3720 1250 3730 1270
rect 3690 1220 3730 1250
rect 3690 1200 3700 1220
rect 3720 1200 3730 1220
rect 3690 1170 3730 1200
rect 3690 1150 3700 1170
rect 3720 1150 3730 1170
rect 3690 1120 3730 1150
rect 3690 1100 3700 1120
rect 3720 1100 3730 1120
rect 3690 1070 3730 1100
rect 3690 1050 3700 1070
rect 3720 1050 3730 1070
rect 3690 1020 3730 1050
rect 3690 1000 3700 1020
rect 3720 1000 3730 1020
rect 3690 985 3730 1000
rect 2680 840 2720 855
rect 2680 820 2690 840
rect 2710 820 2720 840
rect 2680 790 2720 820
rect 2680 770 2690 790
rect 2710 770 2720 790
rect 2680 755 2720 770
rect 3720 840 3760 855
rect 3720 820 3730 840
rect 3750 820 3760 840
rect 3720 790 3760 820
rect 3720 770 3730 790
rect 3750 770 3760 790
rect 3720 755 3760 770
<< pdiff >>
rect 2510 2785 2550 2800
rect 2510 2765 2520 2785
rect 2540 2765 2550 2785
rect 2510 2735 2550 2765
rect 2510 2715 2520 2735
rect 2540 2715 2550 2735
rect 2510 2685 2550 2715
rect 2510 2665 2520 2685
rect 2540 2665 2550 2685
rect 2510 2635 2550 2665
rect 2510 2615 2520 2635
rect 2540 2615 2550 2635
rect 2510 2585 2550 2615
rect 2510 2565 2520 2585
rect 2540 2565 2550 2585
rect 2510 2535 2550 2565
rect 2510 2515 2520 2535
rect 2540 2515 2550 2535
rect 2510 2485 2550 2515
rect 2510 2465 2520 2485
rect 2540 2465 2550 2485
rect 2510 2435 2550 2465
rect 2510 2415 2520 2435
rect 2540 2415 2550 2435
rect 2510 2400 2550 2415
rect 2610 2785 2650 2800
rect 2610 2765 2620 2785
rect 2640 2765 2650 2785
rect 2610 2735 2650 2765
rect 2610 2715 2620 2735
rect 2640 2715 2650 2735
rect 2610 2685 2650 2715
rect 2610 2665 2620 2685
rect 2640 2665 2650 2685
rect 2610 2635 2650 2665
rect 2610 2615 2620 2635
rect 2640 2615 2650 2635
rect 2610 2585 2650 2615
rect 2610 2565 2620 2585
rect 2640 2565 2650 2585
rect 2610 2535 2650 2565
rect 2610 2515 2620 2535
rect 2640 2515 2650 2535
rect 2610 2485 2650 2515
rect 2610 2465 2620 2485
rect 2640 2465 2650 2485
rect 2610 2435 2650 2465
rect 2610 2415 2620 2435
rect 2640 2415 2650 2435
rect 2610 2400 2650 2415
rect 2710 2785 2750 2800
rect 2710 2765 2720 2785
rect 2740 2765 2750 2785
rect 2710 2735 2750 2765
rect 2710 2715 2720 2735
rect 2740 2715 2750 2735
rect 2710 2685 2750 2715
rect 2710 2665 2720 2685
rect 2740 2665 2750 2685
rect 2710 2635 2750 2665
rect 2710 2615 2720 2635
rect 2740 2615 2750 2635
rect 2710 2585 2750 2615
rect 2710 2565 2720 2585
rect 2740 2565 2750 2585
rect 2710 2535 2750 2565
rect 2710 2515 2720 2535
rect 2740 2515 2750 2535
rect 2710 2485 2750 2515
rect 2710 2465 2720 2485
rect 2740 2465 2750 2485
rect 2710 2435 2750 2465
rect 2710 2415 2720 2435
rect 2740 2415 2750 2435
rect 2710 2400 2750 2415
rect 2810 2785 2850 2800
rect 2810 2765 2820 2785
rect 2840 2765 2850 2785
rect 2810 2735 2850 2765
rect 2810 2715 2820 2735
rect 2840 2715 2850 2735
rect 2810 2685 2850 2715
rect 2810 2665 2820 2685
rect 2840 2665 2850 2685
rect 2810 2635 2850 2665
rect 2810 2615 2820 2635
rect 2840 2615 2850 2635
rect 2810 2585 2850 2615
rect 2810 2565 2820 2585
rect 2840 2565 2850 2585
rect 2810 2535 2850 2565
rect 2810 2515 2820 2535
rect 2840 2515 2850 2535
rect 2810 2485 2850 2515
rect 2810 2465 2820 2485
rect 2840 2465 2850 2485
rect 2810 2435 2850 2465
rect 2810 2415 2820 2435
rect 2840 2415 2850 2435
rect 2810 2400 2850 2415
rect 2910 2785 2950 2800
rect 2910 2765 2920 2785
rect 2940 2765 2950 2785
rect 2910 2735 2950 2765
rect 2910 2715 2920 2735
rect 2940 2715 2950 2735
rect 2910 2685 2950 2715
rect 2910 2665 2920 2685
rect 2940 2665 2950 2685
rect 2910 2635 2950 2665
rect 2910 2615 2920 2635
rect 2940 2615 2950 2635
rect 2910 2585 2950 2615
rect 2910 2565 2920 2585
rect 2940 2565 2950 2585
rect 2910 2535 2950 2565
rect 2910 2515 2920 2535
rect 2940 2515 2950 2535
rect 2910 2485 2950 2515
rect 2910 2465 2920 2485
rect 2940 2465 2950 2485
rect 2910 2435 2950 2465
rect 2910 2415 2920 2435
rect 2940 2415 2950 2435
rect 2910 2400 2950 2415
rect 3010 2785 3050 2800
rect 3010 2765 3020 2785
rect 3040 2765 3050 2785
rect 3010 2735 3050 2765
rect 3010 2715 3020 2735
rect 3040 2715 3050 2735
rect 3010 2685 3050 2715
rect 3010 2665 3020 2685
rect 3040 2665 3050 2685
rect 3010 2635 3050 2665
rect 3010 2615 3020 2635
rect 3040 2615 3050 2635
rect 3010 2585 3050 2615
rect 3010 2565 3020 2585
rect 3040 2565 3050 2585
rect 3010 2535 3050 2565
rect 3010 2515 3020 2535
rect 3040 2515 3050 2535
rect 3010 2485 3050 2515
rect 3010 2465 3020 2485
rect 3040 2465 3050 2485
rect 3010 2435 3050 2465
rect 3010 2415 3020 2435
rect 3040 2415 3050 2435
rect 3010 2400 3050 2415
rect 3110 2785 3150 2800
rect 3110 2765 3120 2785
rect 3140 2765 3150 2785
rect 3110 2735 3150 2765
rect 3110 2715 3120 2735
rect 3140 2715 3150 2735
rect 3110 2685 3150 2715
rect 3110 2665 3120 2685
rect 3140 2665 3150 2685
rect 3110 2635 3150 2665
rect 3110 2615 3120 2635
rect 3140 2615 3150 2635
rect 3110 2585 3150 2615
rect 3110 2565 3120 2585
rect 3140 2565 3150 2585
rect 3110 2535 3150 2565
rect 3110 2515 3120 2535
rect 3140 2515 3150 2535
rect 3110 2485 3150 2515
rect 3110 2465 3120 2485
rect 3140 2465 3150 2485
rect 3110 2435 3150 2465
rect 3110 2415 3120 2435
rect 3140 2415 3150 2435
rect 3110 2400 3150 2415
rect 3210 2785 3250 2800
rect 3210 2765 3220 2785
rect 3240 2765 3250 2785
rect 3210 2735 3250 2765
rect 3210 2715 3220 2735
rect 3240 2715 3250 2735
rect 3210 2685 3250 2715
rect 3210 2665 3220 2685
rect 3240 2665 3250 2685
rect 3210 2635 3250 2665
rect 3210 2615 3220 2635
rect 3240 2615 3250 2635
rect 3210 2585 3250 2615
rect 3210 2565 3220 2585
rect 3240 2565 3250 2585
rect 3210 2535 3250 2565
rect 3210 2515 3220 2535
rect 3240 2515 3250 2535
rect 3210 2485 3250 2515
rect 3210 2465 3220 2485
rect 3240 2465 3250 2485
rect 3210 2435 3250 2465
rect 3210 2415 3220 2435
rect 3240 2415 3250 2435
rect 3210 2400 3250 2415
rect 3310 2785 3350 2800
rect 3310 2765 3320 2785
rect 3340 2765 3350 2785
rect 3310 2735 3350 2765
rect 3310 2715 3320 2735
rect 3340 2715 3350 2735
rect 3310 2685 3350 2715
rect 3310 2665 3320 2685
rect 3340 2665 3350 2685
rect 3310 2635 3350 2665
rect 3310 2615 3320 2635
rect 3340 2615 3350 2635
rect 3310 2585 3350 2615
rect 3310 2565 3320 2585
rect 3340 2565 3350 2585
rect 3310 2535 3350 2565
rect 3310 2515 3320 2535
rect 3340 2515 3350 2535
rect 3310 2485 3350 2515
rect 3310 2465 3320 2485
rect 3340 2465 3350 2485
rect 3310 2435 3350 2465
rect 3310 2415 3320 2435
rect 3340 2415 3350 2435
rect 3310 2400 3350 2415
rect 3410 2785 3450 2800
rect 3410 2765 3420 2785
rect 3440 2765 3450 2785
rect 3410 2735 3450 2765
rect 3410 2715 3420 2735
rect 3440 2715 3450 2735
rect 3410 2685 3450 2715
rect 3410 2665 3420 2685
rect 3440 2665 3450 2685
rect 3410 2635 3450 2665
rect 3410 2615 3420 2635
rect 3440 2615 3450 2635
rect 3410 2585 3450 2615
rect 3410 2565 3420 2585
rect 3440 2565 3450 2585
rect 3410 2535 3450 2565
rect 3410 2515 3420 2535
rect 3440 2515 3450 2535
rect 3410 2485 3450 2515
rect 3410 2465 3420 2485
rect 3440 2465 3450 2485
rect 3410 2435 3450 2465
rect 3410 2415 3420 2435
rect 3440 2415 3450 2435
rect 3410 2400 3450 2415
rect 3510 2785 3550 2800
rect 3510 2765 3520 2785
rect 3540 2765 3550 2785
rect 3510 2735 3550 2765
rect 3510 2715 3520 2735
rect 3540 2715 3550 2735
rect 3510 2685 3550 2715
rect 3510 2665 3520 2685
rect 3540 2665 3550 2685
rect 3510 2635 3550 2665
rect 3510 2615 3520 2635
rect 3540 2615 3550 2635
rect 3510 2585 3550 2615
rect 3510 2565 3520 2585
rect 3540 2565 3550 2585
rect 3510 2535 3550 2565
rect 3510 2515 3520 2535
rect 3540 2515 3550 2535
rect 3510 2485 3550 2515
rect 3510 2465 3520 2485
rect 3540 2465 3550 2485
rect 3510 2435 3550 2465
rect 3510 2415 3520 2435
rect 3540 2415 3550 2435
rect 3510 2400 3550 2415
rect 3610 2785 3650 2800
rect 3610 2765 3620 2785
rect 3640 2765 3650 2785
rect 3610 2735 3650 2765
rect 3610 2715 3620 2735
rect 3640 2715 3650 2735
rect 3610 2685 3650 2715
rect 3610 2665 3620 2685
rect 3640 2665 3650 2685
rect 3610 2635 3650 2665
rect 3610 2615 3620 2635
rect 3640 2615 3650 2635
rect 3610 2585 3650 2615
rect 3610 2565 3620 2585
rect 3640 2565 3650 2585
rect 3610 2535 3650 2565
rect 3610 2515 3620 2535
rect 3640 2515 3650 2535
rect 3610 2485 3650 2515
rect 3610 2465 3620 2485
rect 3640 2465 3650 2485
rect 3610 2435 3650 2465
rect 3610 2415 3620 2435
rect 3640 2415 3650 2435
rect 3610 2400 3650 2415
rect 3710 2785 3750 2800
rect 3710 2765 3720 2785
rect 3740 2765 3750 2785
rect 3710 2735 3750 2765
rect 3710 2715 3720 2735
rect 3740 2715 3750 2735
rect 3710 2685 3750 2715
rect 3710 2665 3720 2685
rect 3740 2665 3750 2685
rect 3710 2635 3750 2665
rect 3710 2615 3720 2635
rect 3740 2615 3750 2635
rect 3710 2585 3750 2615
rect 3710 2565 3720 2585
rect 3740 2565 3750 2585
rect 3710 2535 3750 2565
rect 3710 2515 3720 2535
rect 3740 2515 3750 2535
rect 3710 2485 3750 2515
rect 3710 2465 3720 2485
rect 3740 2465 3750 2485
rect 3710 2435 3750 2465
rect 3710 2415 3720 2435
rect 3740 2415 3750 2435
rect 3710 2400 3750 2415
rect 3810 2785 3850 2800
rect 3810 2765 3820 2785
rect 3840 2765 3850 2785
rect 3810 2735 3850 2765
rect 3810 2715 3820 2735
rect 3840 2715 3850 2735
rect 3810 2685 3850 2715
rect 3810 2665 3820 2685
rect 3840 2665 3850 2685
rect 3810 2635 3850 2665
rect 3810 2615 3820 2635
rect 3840 2615 3850 2635
rect 3810 2585 3850 2615
rect 3810 2565 3820 2585
rect 3840 2565 3850 2585
rect 3810 2535 3850 2565
rect 3810 2515 3820 2535
rect 3840 2515 3850 2535
rect 3810 2485 3850 2515
rect 3810 2465 3820 2485
rect 3840 2465 3850 2485
rect 3810 2435 3850 2465
rect 3810 2415 3820 2435
rect 3840 2415 3850 2435
rect 3810 2400 3850 2415
rect 3910 2785 3950 2800
rect 3910 2765 3920 2785
rect 3940 2765 3950 2785
rect 3910 2735 3950 2765
rect 3910 2715 3920 2735
rect 3940 2715 3950 2735
rect 3910 2685 3950 2715
rect 3910 2665 3920 2685
rect 3940 2665 3950 2685
rect 3910 2635 3950 2665
rect 3910 2615 3920 2635
rect 3940 2615 3950 2635
rect 3910 2585 3950 2615
rect 3910 2565 3920 2585
rect 3940 2565 3950 2585
rect 3910 2535 3950 2565
rect 3910 2515 3920 2535
rect 3940 2515 3950 2535
rect 3910 2485 3950 2515
rect 3910 2465 3920 2485
rect 3940 2465 3950 2485
rect 3910 2435 3950 2465
rect 3910 2415 3920 2435
rect 3940 2415 3950 2435
rect 3910 2400 3950 2415
rect 2510 2165 2550 2180
rect 2510 2145 2520 2165
rect 2540 2145 2550 2165
rect 2510 2115 2550 2145
rect 2510 2095 2520 2115
rect 2540 2095 2550 2115
rect 2510 2065 2550 2095
rect 2510 2045 2520 2065
rect 2540 2045 2550 2065
rect 2510 2015 2550 2045
rect 2510 1995 2520 2015
rect 2540 1995 2550 2015
rect 2510 1980 2550 1995
rect 2610 2165 2650 2180
rect 2610 2145 2620 2165
rect 2640 2145 2650 2165
rect 2610 2115 2650 2145
rect 2610 2095 2620 2115
rect 2640 2095 2650 2115
rect 2610 2065 2650 2095
rect 2610 2045 2620 2065
rect 2640 2045 2650 2065
rect 2610 2015 2650 2045
rect 2610 1995 2620 2015
rect 2640 1995 2650 2015
rect 2610 1980 2650 1995
rect 2710 2165 2750 2180
rect 2710 2145 2720 2165
rect 2740 2145 2750 2165
rect 2710 2115 2750 2145
rect 2710 2095 2720 2115
rect 2740 2095 2750 2115
rect 2710 2065 2750 2095
rect 2710 2045 2720 2065
rect 2740 2045 2750 2065
rect 2710 2015 2750 2045
rect 2710 1995 2720 2015
rect 2740 1995 2750 2015
rect 2710 1980 2750 1995
rect 2810 2165 2850 2180
rect 2810 2145 2820 2165
rect 2840 2145 2850 2165
rect 2810 2115 2850 2145
rect 2810 2095 2820 2115
rect 2840 2095 2850 2115
rect 2810 2065 2850 2095
rect 2810 2045 2820 2065
rect 2840 2045 2850 2065
rect 2810 2015 2850 2045
rect 2810 1995 2820 2015
rect 2840 1995 2850 2015
rect 2810 1980 2850 1995
rect 2910 2165 2950 2180
rect 2910 2145 2920 2165
rect 2940 2145 2950 2165
rect 2910 2115 2950 2145
rect 2910 2095 2920 2115
rect 2940 2095 2950 2115
rect 2910 2065 2950 2095
rect 2910 2045 2920 2065
rect 2940 2045 2950 2065
rect 2910 2015 2950 2045
rect 2910 1995 2920 2015
rect 2940 1995 2950 2015
rect 2910 1980 2950 1995
rect 3010 2165 3050 2180
rect 3010 2145 3020 2165
rect 3040 2145 3050 2165
rect 3010 2115 3050 2145
rect 3010 2095 3020 2115
rect 3040 2095 3050 2115
rect 3010 2065 3050 2095
rect 3010 2045 3020 2065
rect 3040 2045 3050 2065
rect 3010 2015 3050 2045
rect 3010 1995 3020 2015
rect 3040 1995 3050 2015
rect 3010 1980 3050 1995
rect 3110 2165 3150 2180
rect 3110 2145 3120 2165
rect 3140 2145 3150 2165
rect 3110 2115 3150 2145
rect 3110 2095 3120 2115
rect 3140 2095 3150 2115
rect 3110 2065 3150 2095
rect 3110 2045 3120 2065
rect 3140 2045 3150 2065
rect 3110 2015 3150 2045
rect 3110 1995 3120 2015
rect 3140 1995 3150 2015
rect 3110 1980 3150 1995
rect 3210 2165 3250 2180
rect 3210 2145 3220 2165
rect 3240 2145 3250 2165
rect 3210 2115 3250 2145
rect 3210 2095 3220 2115
rect 3240 2095 3250 2115
rect 3210 2065 3250 2095
rect 3210 2045 3220 2065
rect 3240 2045 3250 2065
rect 3210 2015 3250 2045
rect 3210 1995 3220 2015
rect 3240 1995 3250 2015
rect 3210 1980 3250 1995
rect 3310 2165 3350 2180
rect 3310 2145 3320 2165
rect 3340 2145 3350 2165
rect 3310 2115 3350 2145
rect 3310 2095 3320 2115
rect 3340 2095 3350 2115
rect 3310 2065 3350 2095
rect 3310 2045 3320 2065
rect 3340 2045 3350 2065
rect 3310 2015 3350 2045
rect 3310 1995 3320 2015
rect 3340 1995 3350 2015
rect 3310 1980 3350 1995
rect 3410 2165 3450 2180
rect 3410 2145 3420 2165
rect 3440 2145 3450 2165
rect 3410 2115 3450 2145
rect 3410 2095 3420 2115
rect 3440 2095 3450 2115
rect 3410 2065 3450 2095
rect 3410 2045 3420 2065
rect 3440 2045 3450 2065
rect 3410 2015 3450 2045
rect 3410 1995 3420 2015
rect 3440 1995 3450 2015
rect 3410 1980 3450 1995
rect 3510 2165 3550 2180
rect 3510 2145 3520 2165
rect 3540 2145 3550 2165
rect 3510 2115 3550 2145
rect 3510 2095 3520 2115
rect 3540 2095 3550 2115
rect 3510 2065 3550 2095
rect 3510 2045 3520 2065
rect 3540 2045 3550 2065
rect 3510 2015 3550 2045
rect 3510 1995 3520 2015
rect 3540 1995 3550 2015
rect 3510 1980 3550 1995
rect 3610 2165 3650 2180
rect 3610 2145 3620 2165
rect 3640 2145 3650 2165
rect 3610 2115 3650 2145
rect 3610 2095 3620 2115
rect 3640 2095 3650 2115
rect 3610 2065 3650 2095
rect 3610 2045 3620 2065
rect 3640 2045 3650 2065
rect 3610 2015 3650 2045
rect 3610 1995 3620 2015
rect 3640 1995 3650 2015
rect 3610 1980 3650 1995
rect 3710 2165 3750 2180
rect 3710 2145 3720 2165
rect 3740 2145 3750 2165
rect 3710 2115 3750 2145
rect 3710 2095 3720 2115
rect 3740 2095 3750 2115
rect 3710 2065 3750 2095
rect 3710 2045 3720 2065
rect 3740 2045 3750 2065
rect 3710 2015 3750 2045
rect 3710 1995 3720 2015
rect 3740 1995 3750 2015
rect 3710 1980 3750 1995
rect 3810 2165 3850 2180
rect 3810 2145 3820 2165
rect 3840 2145 3850 2165
rect 3810 2115 3850 2145
rect 3810 2095 3820 2115
rect 3840 2095 3850 2115
rect 3810 2065 3850 2095
rect 3810 2045 3820 2065
rect 3840 2045 3850 2065
rect 3810 2015 3850 2045
rect 3810 1995 3820 2015
rect 3840 1995 3850 2015
rect 3810 1980 3850 1995
rect 3910 2165 3950 2180
rect 3910 2145 3920 2165
rect 3940 2145 3950 2165
rect 3910 2115 3950 2145
rect 3910 2095 3920 2115
rect 3940 2095 3950 2115
rect 3910 2065 3950 2095
rect 3910 2045 3920 2065
rect 3940 2045 3950 2065
rect 3910 2015 3950 2045
rect 3910 1995 3920 2015
rect 3940 1995 3950 2015
rect 3910 1980 3950 1995
rect 4375 2165 4415 2180
rect 4375 2145 4385 2165
rect 4405 2145 4415 2165
rect 4375 2115 4415 2145
rect 4375 2095 4385 2115
rect 4405 2095 4415 2115
rect 4375 2065 4415 2095
rect 4375 2045 4385 2065
rect 4405 2045 4415 2065
rect 4375 2015 4415 2045
rect 4375 1995 4385 2015
rect 4405 1995 4415 2015
rect 4375 1980 4415 1995
rect 4430 2165 4470 2180
rect 4430 2145 4440 2165
rect 4460 2145 4470 2165
rect 4430 2115 4470 2145
rect 4430 2095 4440 2115
rect 4460 2095 4470 2115
rect 4430 2065 4470 2095
rect 4430 2045 4440 2065
rect 4460 2045 4470 2065
rect 4430 2015 4470 2045
rect 4430 1995 4440 2015
rect 4460 1995 4470 2015
rect 4430 1980 4470 1995
rect 4500 2165 4540 2180
rect 4500 2145 4510 2165
rect 4530 2145 4540 2165
rect 4500 2115 4540 2145
rect 4500 2095 4510 2115
rect 4530 2095 4540 2115
rect 4500 2065 4540 2095
rect 4500 2045 4510 2065
rect 4530 2045 4540 2065
rect 4500 2015 4540 2045
rect 4500 1995 4510 2015
rect 4530 1995 4540 2015
rect 4500 1980 4540 1995
rect 4555 2165 4595 2180
rect 4555 2145 4565 2165
rect 4585 2145 4595 2165
rect 4555 2115 4595 2145
rect 4555 2095 4565 2115
rect 4585 2095 4595 2115
rect 4555 2065 4595 2095
rect 4555 2045 4565 2065
rect 4585 2045 4595 2065
rect 4555 2015 4595 2045
rect 4555 1995 4565 2015
rect 4585 1995 4595 2015
rect 4555 1980 4595 1995
<< ndiffc >>
rect 2720 1625 2740 1645
rect 2720 1575 2740 1595
rect 2820 1625 2840 1645
rect 2820 1575 2840 1595
rect 2920 1625 2940 1645
rect 2920 1575 2940 1595
rect 3020 1625 3040 1645
rect 3020 1575 3040 1595
rect 3120 1625 3140 1645
rect 3120 1575 3140 1595
rect 3220 1625 3240 1645
rect 3220 1575 3240 1595
rect 3320 1625 3340 1645
rect 3320 1575 3340 1595
rect 3420 1625 3440 1645
rect 3420 1575 3440 1595
rect 3520 1625 3540 1645
rect 3520 1575 3540 1595
rect 3620 1625 3640 1645
rect 3620 1575 3640 1595
rect 3720 1625 3740 1645
rect 3720 1575 3740 1595
rect 2740 1350 2760 1370
rect 2740 1300 2760 1320
rect 2740 1250 2760 1270
rect 2740 1200 2760 1220
rect 2740 1150 2760 1170
rect 2740 1100 2760 1120
rect 2740 1050 2760 1070
rect 2740 1000 2760 1020
rect 3180 1350 3200 1370
rect 3260 1350 3280 1370
rect 3180 1300 3200 1320
rect 3260 1300 3280 1320
rect 3180 1250 3200 1270
rect 3260 1250 3280 1270
rect 3180 1200 3200 1220
rect 3260 1200 3280 1220
rect 3180 1150 3200 1170
rect 3260 1150 3280 1170
rect 3180 1100 3200 1120
rect 3260 1100 3280 1120
rect 3180 1050 3200 1070
rect 3260 1050 3280 1070
rect 3180 1000 3200 1020
rect 3260 1000 3280 1020
rect 3700 1350 3720 1370
rect 3700 1300 3720 1320
rect 3700 1250 3720 1270
rect 3700 1200 3720 1220
rect 3700 1150 3720 1170
rect 3700 1100 3720 1120
rect 3700 1050 3720 1070
rect 3700 1000 3720 1020
rect 2690 820 2710 840
rect 2690 770 2710 790
rect 3730 820 3750 840
rect 3730 770 3750 790
<< pdiffc >>
rect 2520 2765 2540 2785
rect 2520 2715 2540 2735
rect 2520 2665 2540 2685
rect 2520 2615 2540 2635
rect 2520 2565 2540 2585
rect 2520 2515 2540 2535
rect 2520 2465 2540 2485
rect 2520 2415 2540 2435
rect 2620 2765 2640 2785
rect 2620 2715 2640 2735
rect 2620 2665 2640 2685
rect 2620 2615 2640 2635
rect 2620 2565 2640 2585
rect 2620 2515 2640 2535
rect 2620 2465 2640 2485
rect 2620 2415 2640 2435
rect 2720 2765 2740 2785
rect 2720 2715 2740 2735
rect 2720 2665 2740 2685
rect 2720 2615 2740 2635
rect 2720 2565 2740 2585
rect 2720 2515 2740 2535
rect 2720 2465 2740 2485
rect 2720 2415 2740 2435
rect 2820 2765 2840 2785
rect 2820 2715 2840 2735
rect 2820 2665 2840 2685
rect 2820 2615 2840 2635
rect 2820 2565 2840 2585
rect 2820 2515 2840 2535
rect 2820 2465 2840 2485
rect 2820 2415 2840 2435
rect 2920 2765 2940 2785
rect 2920 2715 2940 2735
rect 2920 2665 2940 2685
rect 2920 2615 2940 2635
rect 2920 2565 2940 2585
rect 2920 2515 2940 2535
rect 2920 2465 2940 2485
rect 2920 2415 2940 2435
rect 3020 2765 3040 2785
rect 3020 2715 3040 2735
rect 3020 2665 3040 2685
rect 3020 2615 3040 2635
rect 3020 2565 3040 2585
rect 3020 2515 3040 2535
rect 3020 2465 3040 2485
rect 3020 2415 3040 2435
rect 3120 2765 3140 2785
rect 3120 2715 3140 2735
rect 3120 2665 3140 2685
rect 3120 2615 3140 2635
rect 3120 2565 3140 2585
rect 3120 2515 3140 2535
rect 3120 2465 3140 2485
rect 3120 2415 3140 2435
rect 3220 2765 3240 2785
rect 3220 2715 3240 2735
rect 3220 2665 3240 2685
rect 3220 2615 3240 2635
rect 3220 2565 3240 2585
rect 3220 2515 3240 2535
rect 3220 2465 3240 2485
rect 3220 2415 3240 2435
rect 3320 2765 3340 2785
rect 3320 2715 3340 2735
rect 3320 2665 3340 2685
rect 3320 2615 3340 2635
rect 3320 2565 3340 2585
rect 3320 2515 3340 2535
rect 3320 2465 3340 2485
rect 3320 2415 3340 2435
rect 3420 2765 3440 2785
rect 3420 2715 3440 2735
rect 3420 2665 3440 2685
rect 3420 2615 3440 2635
rect 3420 2565 3440 2585
rect 3420 2515 3440 2535
rect 3420 2465 3440 2485
rect 3420 2415 3440 2435
rect 3520 2765 3540 2785
rect 3520 2715 3540 2735
rect 3520 2665 3540 2685
rect 3520 2615 3540 2635
rect 3520 2565 3540 2585
rect 3520 2515 3540 2535
rect 3520 2465 3540 2485
rect 3520 2415 3540 2435
rect 3620 2765 3640 2785
rect 3620 2715 3640 2735
rect 3620 2665 3640 2685
rect 3620 2615 3640 2635
rect 3620 2565 3640 2585
rect 3620 2515 3640 2535
rect 3620 2465 3640 2485
rect 3620 2415 3640 2435
rect 3720 2765 3740 2785
rect 3720 2715 3740 2735
rect 3720 2665 3740 2685
rect 3720 2615 3740 2635
rect 3720 2565 3740 2585
rect 3720 2515 3740 2535
rect 3720 2465 3740 2485
rect 3720 2415 3740 2435
rect 3820 2765 3840 2785
rect 3820 2715 3840 2735
rect 3820 2665 3840 2685
rect 3820 2615 3840 2635
rect 3820 2565 3840 2585
rect 3820 2515 3840 2535
rect 3820 2465 3840 2485
rect 3820 2415 3840 2435
rect 3920 2765 3940 2785
rect 3920 2715 3940 2735
rect 3920 2665 3940 2685
rect 3920 2615 3940 2635
rect 3920 2565 3940 2585
rect 3920 2515 3940 2535
rect 3920 2465 3940 2485
rect 3920 2415 3940 2435
rect 2520 2145 2540 2165
rect 2520 2095 2540 2115
rect 2520 2045 2540 2065
rect 2520 1995 2540 2015
rect 2620 2145 2640 2165
rect 2620 2095 2640 2115
rect 2620 2045 2640 2065
rect 2620 1995 2640 2015
rect 2720 2145 2740 2165
rect 2720 2095 2740 2115
rect 2720 2045 2740 2065
rect 2720 1995 2740 2015
rect 2820 2145 2840 2165
rect 2820 2095 2840 2115
rect 2820 2045 2840 2065
rect 2820 1995 2840 2015
rect 2920 2145 2940 2165
rect 2920 2095 2940 2115
rect 2920 2045 2940 2065
rect 2920 1995 2940 2015
rect 3020 2145 3040 2165
rect 3020 2095 3040 2115
rect 3020 2045 3040 2065
rect 3020 1995 3040 2015
rect 3120 2145 3140 2165
rect 3120 2095 3140 2115
rect 3120 2045 3140 2065
rect 3120 1995 3140 2015
rect 3220 2145 3240 2165
rect 3220 2095 3240 2115
rect 3220 2045 3240 2065
rect 3220 1995 3240 2015
rect 3320 2145 3340 2165
rect 3320 2095 3340 2115
rect 3320 2045 3340 2065
rect 3320 1995 3340 2015
rect 3420 2145 3440 2165
rect 3420 2095 3440 2115
rect 3420 2045 3440 2065
rect 3420 1995 3440 2015
rect 3520 2145 3540 2165
rect 3520 2095 3540 2115
rect 3520 2045 3540 2065
rect 3520 1995 3540 2015
rect 3620 2145 3640 2165
rect 3620 2095 3640 2115
rect 3620 2045 3640 2065
rect 3620 1995 3640 2015
rect 3720 2145 3740 2165
rect 3720 2095 3740 2115
rect 3720 2045 3740 2065
rect 3720 1995 3740 2015
rect 3820 2145 3840 2165
rect 3820 2095 3840 2115
rect 3820 2045 3840 2065
rect 3820 1995 3840 2015
rect 3920 2145 3940 2165
rect 3920 2095 3940 2115
rect 3920 2045 3940 2065
rect 3920 1995 3940 2015
rect 4385 2145 4405 2165
rect 4385 2095 4405 2115
rect 4385 2045 4405 2065
rect 4385 1995 4405 2015
rect 4440 2145 4460 2165
rect 4440 2095 4460 2115
rect 4440 2045 4460 2065
rect 4440 1995 4460 2015
rect 4510 2145 4530 2165
rect 4510 2095 4530 2115
rect 4510 2045 4530 2065
rect 4510 1995 4530 2015
rect 4565 2145 4585 2165
rect 4565 2095 4585 2115
rect 4565 2045 4585 2065
rect 4565 1995 4585 2015
<< psubdiff >>
rect 3210 1370 3250 1385
rect 3210 1350 3220 1370
rect 3240 1350 3250 1370
rect 3210 1320 3250 1350
rect 3210 1300 3220 1320
rect 3240 1300 3250 1320
rect 3210 1270 3250 1300
rect 3210 1250 3220 1270
rect 3240 1250 3250 1270
rect 3210 1220 3250 1250
rect 3210 1200 3220 1220
rect 3240 1200 3250 1220
rect 3210 1170 3250 1200
rect 3210 1150 3220 1170
rect 3240 1150 3250 1170
rect 3210 1120 3250 1150
rect 3210 1100 3220 1120
rect 3240 1100 3250 1120
rect 3210 1070 3250 1100
rect 3210 1050 3220 1070
rect 3240 1050 3250 1070
rect 3210 1020 3250 1050
rect 3210 1000 3220 1020
rect 3240 1000 3250 1020
rect 3210 985 3250 1000
rect 645 820 695 835
rect 645 800 660 820
rect 680 800 695 820
rect 645 770 695 800
rect 645 750 660 770
rect 680 750 695 770
rect 3760 840 3800 855
rect 3760 820 3770 840
rect 3790 820 3800 840
rect 3760 790 3800 820
rect 3760 770 3770 790
rect 3790 770 3800 790
rect 3760 755 3800 770
rect 645 720 695 750
rect 645 700 660 720
rect 680 700 695 720
rect 645 685 695 700
<< nsubdiff >>
rect 2470 2785 2510 2800
rect 2470 2765 2480 2785
rect 2500 2765 2510 2785
rect 2470 2735 2510 2765
rect 2470 2715 2480 2735
rect 2500 2715 2510 2735
rect 2470 2685 2510 2715
rect 2470 2665 2480 2685
rect 2500 2665 2510 2685
rect 2470 2635 2510 2665
rect 2470 2615 2480 2635
rect 2500 2615 2510 2635
rect 2470 2585 2510 2615
rect 2470 2565 2480 2585
rect 2500 2565 2510 2585
rect 2470 2535 2510 2565
rect 2470 2515 2480 2535
rect 2500 2515 2510 2535
rect 2470 2485 2510 2515
rect 2470 2465 2480 2485
rect 2500 2465 2510 2485
rect 2470 2435 2510 2465
rect 2470 2415 2480 2435
rect 2500 2415 2510 2435
rect 2470 2400 2510 2415
rect 3950 2785 3990 2800
rect 3950 2765 3960 2785
rect 3980 2765 3990 2785
rect 3950 2735 3990 2765
rect 3950 2715 3960 2735
rect 3980 2715 3990 2735
rect 3950 2685 3990 2715
rect 3950 2665 3960 2685
rect 3980 2665 3990 2685
rect 3950 2635 3990 2665
rect 3950 2615 3960 2635
rect 3980 2615 3990 2635
rect 3950 2585 3990 2615
rect 3950 2565 3960 2585
rect 3980 2565 3990 2585
rect 3950 2535 3990 2565
rect 3950 2515 3960 2535
rect 3980 2515 3990 2535
rect 3950 2485 3990 2515
rect 3950 2465 3960 2485
rect 3980 2465 3990 2485
rect 3950 2435 3990 2465
rect 3950 2415 3960 2435
rect 3980 2415 3990 2435
rect 3950 2400 3990 2415
rect 2470 2165 2510 2180
rect 2470 2145 2480 2165
rect 2500 2145 2510 2165
rect 2470 2115 2510 2145
rect 2470 2095 2480 2115
rect 2500 2095 2510 2115
rect 2470 2065 2510 2095
rect 2470 2045 2480 2065
rect 2500 2045 2510 2065
rect 2470 2015 2510 2045
rect 2470 1995 2480 2015
rect 2500 1995 2510 2015
rect 2470 1980 2510 1995
rect 3950 2165 3990 2180
rect 3950 2145 3960 2165
rect 3980 2145 3990 2165
rect 3950 2115 3990 2145
rect 3950 2095 3960 2115
rect 3980 2095 3990 2115
rect 3950 2065 3990 2095
rect 3950 2045 3960 2065
rect 3980 2045 3990 2065
rect 3950 2015 3990 2045
rect 3950 1995 3960 2015
rect 3980 1995 3990 2015
rect 3950 1980 3990 1995
<< psubdiffcont >>
rect 3220 1350 3240 1370
rect 3220 1300 3240 1320
rect 3220 1250 3240 1270
rect 3220 1200 3240 1220
rect 3220 1150 3240 1170
rect 3220 1100 3240 1120
rect 3220 1050 3240 1070
rect 3220 1000 3240 1020
rect 660 800 680 820
rect 660 750 680 770
rect 3770 820 3790 840
rect 3770 770 3790 790
rect 660 700 680 720
<< nsubdiffcont >>
rect 2480 2765 2500 2785
rect 2480 2715 2500 2735
rect 2480 2665 2500 2685
rect 2480 2615 2500 2635
rect 2480 2565 2500 2585
rect 2480 2515 2500 2535
rect 2480 2465 2500 2485
rect 2480 2415 2500 2435
rect 3960 2765 3980 2785
rect 3960 2715 3980 2735
rect 3960 2665 3980 2685
rect 3960 2615 3980 2635
rect 3960 2565 3980 2585
rect 3960 2515 3980 2535
rect 3960 2465 3980 2485
rect 3960 2415 3980 2435
rect 2480 2145 2500 2165
rect 2480 2095 2500 2115
rect 2480 2045 2500 2065
rect 2480 1995 2500 2015
rect 3960 2145 3980 2165
rect 3960 2095 3980 2115
rect 3960 2045 3980 2065
rect 3960 1995 3980 2015
<< poly >>
rect 2560 2845 2600 2855
rect 2560 2825 2570 2845
rect 2590 2825 2600 2845
rect 2560 2815 2600 2825
rect 3860 2845 3900 2855
rect 3860 2825 3870 2845
rect 3890 2825 3900 2845
rect 3860 2815 3900 2825
rect 2550 2800 2610 2815
rect 2650 2800 2710 2815
rect 2750 2800 2810 2815
rect 2850 2800 2910 2815
rect 2950 2800 3010 2815
rect 3050 2800 3110 2815
rect 3150 2800 3210 2815
rect 3250 2800 3310 2815
rect 3350 2800 3410 2815
rect 3450 2800 3510 2815
rect 3550 2800 3610 2815
rect 3650 2800 3710 2815
rect 3750 2800 3810 2815
rect 3850 2800 3910 2815
rect 2550 2385 2610 2400
rect 2650 2390 2710 2400
rect 2750 2390 2810 2400
rect 2850 2390 2910 2400
rect 2950 2390 3010 2400
rect 3050 2390 3110 2400
rect 3150 2390 3210 2400
rect 3250 2390 3310 2400
rect 3350 2390 3410 2400
rect 3450 2390 3510 2400
rect 3550 2390 3610 2400
rect 3650 2390 3710 2400
rect 3750 2390 3810 2400
rect 2650 2375 3810 2390
rect 3850 2385 3910 2400
rect 3760 2355 3770 2375
rect 3790 2355 3800 2375
rect 3760 2345 3800 2355
rect 4515 2265 4555 2275
rect 4515 2245 4525 2265
rect 4545 2245 4555 2265
rect 4515 2235 4555 2245
rect 2560 2225 2600 2235
rect 2560 2205 2570 2225
rect 2590 2205 2600 2225
rect 2560 2195 2600 2205
rect 3860 2225 3900 2235
rect 3860 2205 3870 2225
rect 3890 2205 3900 2225
rect 3860 2195 3900 2205
rect 2550 2180 2610 2195
rect 2650 2180 2710 2195
rect 2750 2180 2810 2195
rect 2850 2180 2910 2195
rect 2950 2180 3010 2195
rect 3050 2180 3110 2195
rect 3150 2180 3210 2195
rect 3250 2180 3310 2195
rect 3350 2180 3410 2195
rect 3450 2180 3510 2195
rect 3550 2180 3610 2195
rect 3650 2180 3710 2195
rect 3750 2180 3810 2195
rect 3850 2180 3910 2195
rect 4415 2180 4430 2195
rect 4540 2180 4555 2235
rect 2550 1965 2610 1980
rect 2650 1965 2710 1980
rect 2750 1970 2810 1980
rect 2850 1970 2910 1980
rect 2950 1970 3010 1980
rect 3050 1970 3110 1980
rect 2670 1915 2690 1965
rect 2750 1955 3110 1970
rect 3150 1970 3210 1980
rect 3250 1970 3310 1980
rect 3150 1955 3310 1970
rect 3350 1970 3410 1980
rect 3450 1970 3510 1980
rect 3550 1970 3610 1980
rect 3650 1970 3710 1980
rect 3350 1955 3710 1970
rect 3750 1965 3810 1980
rect 3850 1965 3910 1980
rect 2810 1950 2850 1955
rect 2810 1930 2820 1950
rect 2840 1930 2850 1950
rect 2810 1920 2850 1930
rect 3170 1915 3190 1955
rect 3270 1915 3290 1955
rect 3610 1950 3650 1955
rect 3610 1930 3620 1950
rect 3640 1930 3650 1950
rect 3610 1920 3650 1930
rect 3770 1915 3790 1965
rect 4415 1940 4430 1980
rect 4540 1965 4555 1980
rect 4485 1940 4525 1950
rect 4415 1920 4495 1940
rect 4515 1920 4525 1940
rect 2660 1905 2700 1915
rect 2660 1885 2670 1905
rect 2690 1885 2700 1905
rect 2660 1875 2700 1885
rect 3160 1905 3200 1915
rect 3160 1885 3170 1905
rect 3190 1885 3200 1905
rect 3160 1875 3200 1885
rect 3260 1905 3300 1915
rect 3260 1885 3270 1905
rect 3290 1885 3300 1905
rect 3260 1875 3300 1885
rect 3760 1905 3800 1915
rect 4485 1910 4525 1920
rect 3760 1885 3770 1905
rect 3790 1885 3800 1905
rect 3760 1875 3800 1885
rect 2860 1700 2900 1710
rect 2860 1680 2870 1700
rect 2890 1680 2900 1700
rect 3160 1700 3200 1710
rect 3160 1685 3170 1700
rect 2860 1675 2900 1680
rect 3150 1680 3170 1685
rect 3190 1685 3200 1700
rect 3260 1700 3300 1710
rect 3260 1685 3270 1700
rect 3190 1680 3270 1685
rect 3290 1685 3300 1700
rect 3560 1700 3600 1710
rect 3290 1680 3310 1685
rect 2750 1660 2810 1675
rect 2850 1660 2910 1675
rect 2950 1660 3010 1675
rect 3050 1660 3110 1675
rect 3150 1670 3310 1680
rect 3560 1680 3570 1700
rect 3590 1680 3600 1700
rect 3560 1675 3600 1680
rect 3150 1660 3210 1670
rect 3250 1660 3310 1670
rect 3350 1660 3410 1675
rect 3450 1660 3510 1675
rect 3550 1660 3610 1675
rect 3650 1660 3710 1675
rect 2750 1545 2810 1560
rect 2850 1545 2910 1560
rect 2950 1550 3010 1560
rect 3050 1550 3110 1560
rect 2760 1540 2800 1545
rect 2760 1520 2770 1540
rect 2790 1520 2800 1540
rect 2950 1535 3110 1550
rect 3150 1545 3210 1560
rect 3250 1545 3310 1560
rect 3350 1550 3410 1560
rect 3450 1550 3510 1560
rect 3350 1535 3510 1550
rect 3550 1545 3610 1560
rect 3650 1545 3710 1560
rect 3660 1540 3700 1545
rect 2760 1510 2800 1520
rect 3010 1515 3020 1535
rect 3040 1515 3050 1535
rect 3010 1505 3050 1515
rect 3410 1515 3420 1535
rect 3440 1515 3450 1535
rect 3410 1505 3450 1515
rect 3660 1520 3670 1540
rect 3690 1520 3700 1540
rect 3660 1510 3700 1520
rect 2770 1430 3170 1440
rect 2770 1410 2780 1430
rect 2800 1410 2820 1430
rect 2840 1410 2860 1430
rect 2880 1410 2900 1430
rect 2920 1410 2940 1430
rect 2960 1410 2980 1430
rect 3000 1410 3020 1430
rect 3040 1410 3060 1430
rect 3080 1410 3100 1430
rect 3120 1410 3140 1430
rect 3160 1410 3170 1430
rect 2770 1385 3170 1410
rect 3290 1430 3690 1440
rect 3290 1410 3300 1430
rect 3320 1410 3340 1430
rect 3360 1410 3380 1430
rect 3400 1410 3420 1430
rect 3440 1410 3460 1430
rect 3480 1410 3500 1430
rect 3520 1410 3540 1430
rect 3560 1410 3580 1430
rect 3600 1410 3620 1430
rect 3640 1410 3660 1430
rect 3680 1410 3690 1430
rect 3290 1385 3690 1410
rect 2770 970 3170 985
rect 3290 970 3690 985
rect 2720 900 2760 910
rect 2720 880 2730 900
rect 2750 880 2760 900
rect 2720 870 2760 880
rect 2800 900 2840 910
rect 2800 880 2810 900
rect 2830 880 2840 900
rect 2800 870 2840 880
rect 2880 900 2920 910
rect 2880 880 2890 900
rect 2910 880 2920 900
rect 2880 870 2920 880
rect 2960 900 3000 910
rect 2960 880 2970 900
rect 2990 880 3000 900
rect 2960 870 3000 880
rect 3040 900 3080 910
rect 3040 880 3050 900
rect 3070 880 3080 900
rect 3040 870 3080 880
rect 3120 900 3160 910
rect 3120 880 3130 900
rect 3150 880 3160 900
rect 3120 870 3160 880
rect 3200 900 3240 910
rect 3200 880 3210 900
rect 3230 880 3240 900
rect 3200 870 3240 880
rect 3280 900 3320 910
rect 3280 880 3290 900
rect 3310 880 3320 900
rect 3280 870 3320 880
rect 3360 900 3400 910
rect 3360 880 3370 900
rect 3390 880 3400 900
rect 3360 870 3400 880
rect 3440 900 3480 910
rect 3440 880 3450 900
rect 3470 880 3480 900
rect 3440 870 3480 880
rect 3520 900 3560 910
rect 3520 880 3530 900
rect 3550 880 3560 900
rect 3520 870 3560 880
rect 3600 900 3640 910
rect 3600 880 3610 900
rect 3630 880 3640 900
rect 3600 870 3640 880
rect 3680 900 3720 910
rect 3680 880 3690 900
rect 3710 880 3720 900
rect 3680 870 3720 880
rect 2720 855 3720 870
rect 2720 740 3720 755
<< polycont >>
rect 2570 2825 2590 2845
rect 3870 2825 3890 2845
rect 3770 2355 3790 2375
rect 4525 2245 4545 2265
rect 2570 2205 2590 2225
rect 3870 2205 3890 2225
rect 2820 1930 2840 1950
rect 3620 1930 3640 1950
rect 4495 1920 4515 1940
rect 2670 1885 2690 1905
rect 3170 1885 3190 1905
rect 3270 1885 3290 1905
rect 3770 1885 3790 1905
rect 2870 1680 2890 1700
rect 3170 1680 3190 1700
rect 3270 1680 3290 1700
rect 3570 1680 3590 1700
rect 2770 1520 2790 1540
rect 3020 1515 3040 1535
rect 3420 1515 3440 1535
rect 3670 1520 3690 1540
rect 2780 1410 2800 1430
rect 2820 1410 2840 1430
rect 2860 1410 2880 1430
rect 2900 1410 2920 1430
rect 2940 1410 2960 1430
rect 2980 1410 3000 1430
rect 3020 1410 3040 1430
rect 3060 1410 3080 1430
rect 3100 1410 3120 1430
rect 3140 1410 3160 1430
rect 3300 1410 3320 1430
rect 3340 1410 3360 1430
rect 3380 1410 3400 1430
rect 3420 1410 3440 1430
rect 3460 1410 3480 1430
rect 3500 1410 3520 1430
rect 3540 1410 3560 1430
rect 3580 1410 3600 1430
rect 3620 1410 3640 1430
rect 3660 1410 3680 1430
rect 2730 880 2750 900
rect 2810 880 2830 900
rect 2890 880 2910 900
rect 2970 880 2990 900
rect 3050 880 3070 900
rect 3130 880 3150 900
rect 3210 880 3230 900
rect 3290 880 3310 900
rect 3370 880 3390 900
rect 3450 880 3470 900
rect 3530 880 3550 900
rect 3610 880 3630 900
rect 3690 880 3710 900
<< xpolycontact >>
rect 1005 2560 1225 2595
rect 1895 2560 2115 2595
rect 1005 2500 1225 2535
rect 1895 2500 2115 2535
rect 1005 2440 1225 2475
rect 1895 2440 2115 2475
rect 1005 2380 1225 2415
rect 1895 2380 2115 2415
rect 1005 2320 1225 2355
rect 1895 2320 2115 2355
rect 1005 1975 1225 2010
rect 1895 1975 2115 2010
rect 1005 1915 1225 1950
rect 1895 1915 2115 1950
rect 1005 1855 1225 1890
rect 1895 1855 2115 1890
rect 1005 1795 1225 1830
rect 1895 1795 2115 1830
rect 1005 1735 1225 1770
rect 1895 1735 2115 1770
rect 1005 1505 1225 1540
rect 1575 1505 1795 1540
rect 1005 1445 1225 1480
rect 1895 1445 2115 1480
rect 1005 1385 1225 1420
rect 1895 1385 2115 1420
rect 1005 1325 1225 1360
rect 1895 1325 2115 1360
rect 1005 1265 1225 1300
rect 1895 1265 2115 1300
rect 1005 1205 1225 1240
rect 1895 1205 2115 1240
<< xpolyres >>
rect 1225 2560 1895 2595
rect 1225 2500 1895 2535
rect 1225 2440 1895 2475
rect 1225 2380 1895 2415
rect 1225 2320 1895 2355
rect 1225 1975 1895 2010
rect 1225 1915 1895 1950
rect 1225 1855 1895 1890
rect 1225 1795 1895 1830
rect 1225 1735 1895 1770
rect 1225 1505 1575 1540
rect 1225 1445 1895 1480
rect 1225 1385 1895 1420
rect 1225 1325 1895 1360
rect 1225 1265 1895 1300
rect 1225 1205 1895 1240
<< locali >>
rect 2510 2845 2610 2855
rect 2510 2825 2520 2845
rect 2540 2825 2570 2845
rect 2590 2825 2610 2845
rect 2510 2815 2610 2825
rect 2710 2845 2750 2855
rect 2710 2825 2720 2845
rect 2740 2825 2750 2845
rect 2710 2815 2750 2825
rect 2910 2845 2950 2855
rect 2910 2825 2920 2845
rect 2940 2825 2950 2845
rect 2910 2815 2950 2825
rect 3110 2845 3150 2855
rect 3110 2825 3120 2845
rect 3140 2825 3150 2845
rect 3110 2815 3150 2825
rect 3210 2845 3250 2855
rect 3210 2825 3220 2845
rect 3240 2825 3250 2845
rect 3210 2815 3250 2825
rect 3310 2845 3350 2855
rect 3310 2825 3320 2845
rect 3340 2825 3350 2845
rect 3310 2815 3350 2825
rect 3510 2845 3550 2855
rect 3510 2825 3520 2845
rect 3540 2825 3550 2845
rect 3510 2815 3550 2825
rect 3710 2845 3750 2855
rect 3710 2825 3720 2845
rect 3740 2825 3750 2845
rect 3710 2815 3750 2825
rect 3850 2845 3950 2855
rect 3850 2825 3870 2845
rect 3890 2825 3920 2845
rect 3940 2825 3950 2845
rect 3850 2815 3950 2825
rect 2520 2795 2540 2815
rect 2720 2795 2740 2815
rect 2920 2795 2940 2815
rect 3120 2795 3140 2815
rect 3220 2795 3240 2815
rect 3320 2795 3340 2815
rect 3520 2795 3540 2815
rect 3720 2795 3740 2815
rect 3920 2795 3940 2815
rect 2475 2785 2545 2795
rect 2475 2765 2480 2785
rect 2500 2765 2520 2785
rect 2540 2765 2545 2785
rect 2475 2735 2545 2765
rect 2475 2715 2480 2735
rect 2500 2715 2520 2735
rect 2540 2715 2545 2735
rect 2475 2685 2545 2715
rect 2475 2665 2480 2685
rect 2500 2665 2520 2685
rect 2540 2665 2545 2685
rect 2475 2635 2545 2665
rect 2475 2615 2480 2635
rect 2500 2615 2520 2635
rect 2540 2615 2545 2635
rect 945 2585 1005 2595
rect 945 2565 955 2585
rect 975 2565 1005 2585
rect 945 2560 1005 2565
rect 945 2555 985 2560
rect 1895 2535 2115 2560
rect 2475 2585 2545 2615
rect 2475 2565 2480 2585
rect 2500 2565 2520 2585
rect 2540 2565 2545 2585
rect 2475 2535 2545 2565
rect 2475 2515 2480 2535
rect 2500 2515 2520 2535
rect 2540 2515 2545 2535
rect 1005 2475 1225 2500
rect 2475 2485 2545 2515
rect 1895 2415 2115 2440
rect 2475 2465 2480 2485
rect 2500 2465 2520 2485
rect 2540 2465 2545 2485
rect 2475 2435 2545 2465
rect 2475 2415 2480 2435
rect 2500 2415 2520 2435
rect 2540 2415 2545 2435
rect 2475 2405 2545 2415
rect 2615 2785 2645 2795
rect 2615 2765 2620 2785
rect 2640 2765 2645 2785
rect 2615 2735 2645 2765
rect 2615 2715 2620 2735
rect 2640 2715 2645 2735
rect 2615 2685 2645 2715
rect 2615 2665 2620 2685
rect 2640 2665 2645 2685
rect 2615 2635 2645 2665
rect 2615 2615 2620 2635
rect 2640 2615 2645 2635
rect 2615 2585 2645 2615
rect 2615 2565 2620 2585
rect 2640 2565 2645 2585
rect 2615 2535 2645 2565
rect 2615 2515 2620 2535
rect 2640 2515 2645 2535
rect 2615 2485 2645 2515
rect 2615 2465 2620 2485
rect 2640 2465 2645 2485
rect 2615 2435 2645 2465
rect 2615 2415 2620 2435
rect 2640 2415 2645 2435
rect 2615 2405 2645 2415
rect 2715 2785 2745 2795
rect 2715 2765 2720 2785
rect 2740 2765 2745 2785
rect 2715 2735 2745 2765
rect 2715 2715 2720 2735
rect 2740 2715 2745 2735
rect 2715 2685 2745 2715
rect 2715 2665 2720 2685
rect 2740 2665 2745 2685
rect 2715 2635 2745 2665
rect 2715 2615 2720 2635
rect 2740 2615 2745 2635
rect 2715 2585 2745 2615
rect 2715 2565 2720 2585
rect 2740 2565 2745 2585
rect 2715 2535 2745 2565
rect 2715 2515 2720 2535
rect 2740 2515 2745 2535
rect 2715 2485 2745 2515
rect 2715 2465 2720 2485
rect 2740 2465 2745 2485
rect 2715 2435 2745 2465
rect 2715 2415 2720 2435
rect 2740 2415 2745 2435
rect 2715 2405 2745 2415
rect 2815 2785 2845 2795
rect 2815 2765 2820 2785
rect 2840 2765 2845 2785
rect 2815 2735 2845 2765
rect 2815 2715 2820 2735
rect 2840 2715 2845 2735
rect 2815 2685 2845 2715
rect 2815 2665 2820 2685
rect 2840 2665 2845 2685
rect 2815 2635 2845 2665
rect 2815 2615 2820 2635
rect 2840 2615 2845 2635
rect 2815 2585 2845 2615
rect 2815 2565 2820 2585
rect 2840 2565 2845 2585
rect 2815 2535 2845 2565
rect 2815 2515 2820 2535
rect 2840 2515 2845 2535
rect 2815 2485 2845 2515
rect 2815 2465 2820 2485
rect 2840 2465 2845 2485
rect 2815 2435 2845 2465
rect 2815 2415 2820 2435
rect 2840 2415 2845 2435
rect 2815 2405 2845 2415
rect 2915 2785 2945 2795
rect 2915 2765 2920 2785
rect 2940 2765 2945 2785
rect 2915 2735 2945 2765
rect 2915 2715 2920 2735
rect 2940 2715 2945 2735
rect 2915 2685 2945 2715
rect 2915 2665 2920 2685
rect 2940 2665 2945 2685
rect 2915 2635 2945 2665
rect 2915 2615 2920 2635
rect 2940 2615 2945 2635
rect 2915 2585 2945 2615
rect 2915 2565 2920 2585
rect 2940 2565 2945 2585
rect 2915 2535 2945 2565
rect 2915 2515 2920 2535
rect 2940 2515 2945 2535
rect 2915 2485 2945 2515
rect 2915 2465 2920 2485
rect 2940 2465 2945 2485
rect 2915 2435 2945 2465
rect 2915 2415 2920 2435
rect 2940 2415 2945 2435
rect 2915 2405 2945 2415
rect 3015 2785 3045 2795
rect 3015 2765 3020 2785
rect 3040 2765 3045 2785
rect 3015 2735 3045 2765
rect 3015 2715 3020 2735
rect 3040 2715 3045 2735
rect 3015 2685 3045 2715
rect 3015 2665 3020 2685
rect 3040 2665 3045 2685
rect 3015 2635 3045 2665
rect 3015 2615 3020 2635
rect 3040 2615 3045 2635
rect 3015 2585 3045 2615
rect 3015 2565 3020 2585
rect 3040 2565 3045 2585
rect 3015 2535 3045 2565
rect 3015 2515 3020 2535
rect 3040 2515 3045 2535
rect 3015 2485 3045 2515
rect 3015 2465 3020 2485
rect 3040 2465 3045 2485
rect 3015 2435 3045 2465
rect 3015 2415 3020 2435
rect 3040 2415 3045 2435
rect 3015 2405 3045 2415
rect 3115 2785 3145 2795
rect 3115 2765 3120 2785
rect 3140 2765 3145 2785
rect 3115 2735 3145 2765
rect 3115 2715 3120 2735
rect 3140 2715 3145 2735
rect 3115 2685 3145 2715
rect 3115 2665 3120 2685
rect 3140 2665 3145 2685
rect 3115 2635 3145 2665
rect 3115 2615 3120 2635
rect 3140 2615 3145 2635
rect 3115 2585 3145 2615
rect 3115 2565 3120 2585
rect 3140 2565 3145 2585
rect 3115 2535 3145 2565
rect 3115 2515 3120 2535
rect 3140 2515 3145 2535
rect 3115 2485 3145 2515
rect 3115 2465 3120 2485
rect 3140 2465 3145 2485
rect 3115 2435 3145 2465
rect 3115 2415 3120 2435
rect 3140 2415 3145 2435
rect 3115 2405 3145 2415
rect 3215 2785 3245 2795
rect 3215 2765 3220 2785
rect 3240 2765 3245 2785
rect 3215 2735 3245 2765
rect 3215 2715 3220 2735
rect 3240 2715 3245 2735
rect 3215 2685 3245 2715
rect 3215 2665 3220 2685
rect 3240 2665 3245 2685
rect 3215 2635 3245 2665
rect 3215 2615 3220 2635
rect 3240 2615 3245 2635
rect 3215 2585 3245 2615
rect 3215 2565 3220 2585
rect 3240 2565 3245 2585
rect 3215 2535 3245 2565
rect 3215 2515 3220 2535
rect 3240 2515 3245 2535
rect 3215 2485 3245 2515
rect 3215 2465 3220 2485
rect 3240 2465 3245 2485
rect 3215 2435 3245 2465
rect 3215 2415 3220 2435
rect 3240 2415 3245 2435
rect 3215 2405 3245 2415
rect 3315 2785 3345 2795
rect 3315 2765 3320 2785
rect 3340 2765 3345 2785
rect 3315 2735 3345 2765
rect 3315 2715 3320 2735
rect 3340 2715 3345 2735
rect 3315 2685 3345 2715
rect 3315 2665 3320 2685
rect 3340 2665 3345 2685
rect 3315 2635 3345 2665
rect 3315 2615 3320 2635
rect 3340 2615 3345 2635
rect 3315 2585 3345 2615
rect 3315 2565 3320 2585
rect 3340 2565 3345 2585
rect 3315 2535 3345 2565
rect 3315 2515 3320 2535
rect 3340 2515 3345 2535
rect 3315 2485 3345 2515
rect 3315 2465 3320 2485
rect 3340 2465 3345 2485
rect 3315 2435 3345 2465
rect 3315 2415 3320 2435
rect 3340 2415 3345 2435
rect 3315 2405 3345 2415
rect 3415 2785 3445 2795
rect 3415 2765 3420 2785
rect 3440 2765 3445 2785
rect 3415 2735 3445 2765
rect 3415 2715 3420 2735
rect 3440 2715 3445 2735
rect 3415 2685 3445 2715
rect 3415 2665 3420 2685
rect 3440 2665 3445 2685
rect 3415 2635 3445 2665
rect 3415 2615 3420 2635
rect 3440 2615 3445 2635
rect 3415 2585 3445 2615
rect 3415 2565 3420 2585
rect 3440 2565 3445 2585
rect 3415 2535 3445 2565
rect 3415 2515 3420 2535
rect 3440 2515 3445 2535
rect 3415 2485 3445 2515
rect 3415 2465 3420 2485
rect 3440 2465 3445 2485
rect 3415 2435 3445 2465
rect 3415 2415 3420 2435
rect 3440 2415 3445 2435
rect 3415 2405 3445 2415
rect 3515 2785 3545 2795
rect 3515 2765 3520 2785
rect 3540 2765 3545 2785
rect 3515 2735 3545 2765
rect 3515 2715 3520 2735
rect 3540 2715 3545 2735
rect 3515 2685 3545 2715
rect 3515 2665 3520 2685
rect 3540 2665 3545 2685
rect 3515 2635 3545 2665
rect 3515 2615 3520 2635
rect 3540 2615 3545 2635
rect 3515 2585 3545 2615
rect 3515 2565 3520 2585
rect 3540 2565 3545 2585
rect 3515 2535 3545 2565
rect 3515 2515 3520 2535
rect 3540 2515 3545 2535
rect 3515 2485 3545 2515
rect 3515 2465 3520 2485
rect 3540 2465 3545 2485
rect 3515 2435 3545 2465
rect 3515 2415 3520 2435
rect 3540 2415 3545 2435
rect 3515 2405 3545 2415
rect 3615 2785 3645 2795
rect 3615 2765 3620 2785
rect 3640 2765 3645 2785
rect 3615 2735 3645 2765
rect 3615 2715 3620 2735
rect 3640 2715 3645 2735
rect 3615 2685 3645 2715
rect 3615 2665 3620 2685
rect 3640 2665 3645 2685
rect 3615 2635 3645 2665
rect 3615 2615 3620 2635
rect 3640 2615 3645 2635
rect 3615 2585 3645 2615
rect 3615 2565 3620 2585
rect 3640 2565 3645 2585
rect 3615 2535 3645 2565
rect 3615 2515 3620 2535
rect 3640 2515 3645 2535
rect 3615 2485 3645 2515
rect 3615 2465 3620 2485
rect 3640 2465 3645 2485
rect 3615 2435 3645 2465
rect 3615 2415 3620 2435
rect 3640 2415 3645 2435
rect 3615 2405 3645 2415
rect 3715 2785 3745 2795
rect 3715 2765 3720 2785
rect 3740 2765 3745 2785
rect 3715 2735 3745 2765
rect 3715 2715 3720 2735
rect 3740 2715 3745 2735
rect 3715 2685 3745 2715
rect 3715 2665 3720 2685
rect 3740 2665 3745 2685
rect 3715 2635 3745 2665
rect 3715 2615 3720 2635
rect 3740 2615 3745 2635
rect 3715 2585 3745 2615
rect 3715 2565 3720 2585
rect 3740 2565 3745 2585
rect 3715 2535 3745 2565
rect 3715 2515 3720 2535
rect 3740 2515 3745 2535
rect 3715 2485 3745 2515
rect 3715 2465 3720 2485
rect 3740 2465 3745 2485
rect 3715 2435 3745 2465
rect 3715 2415 3720 2435
rect 3740 2415 3745 2435
rect 3715 2405 3745 2415
rect 3815 2785 3845 2795
rect 3815 2765 3820 2785
rect 3840 2765 3845 2785
rect 3815 2735 3845 2765
rect 3815 2715 3820 2735
rect 3840 2715 3845 2735
rect 3815 2685 3845 2715
rect 3815 2665 3820 2685
rect 3840 2665 3845 2685
rect 3815 2635 3845 2665
rect 3815 2615 3820 2635
rect 3840 2615 3845 2635
rect 3815 2585 3845 2615
rect 3815 2565 3820 2585
rect 3840 2565 3845 2585
rect 3815 2535 3845 2565
rect 3815 2515 3820 2535
rect 3840 2515 3845 2535
rect 3815 2485 3845 2515
rect 3815 2465 3820 2485
rect 3840 2465 3845 2485
rect 3815 2435 3845 2465
rect 3815 2415 3820 2435
rect 3840 2415 3845 2435
rect 3815 2405 3845 2415
rect 3915 2785 3985 2795
rect 3915 2765 3920 2785
rect 3940 2765 3960 2785
rect 3980 2765 3985 2785
rect 3915 2735 3985 2765
rect 3915 2715 3920 2735
rect 3940 2715 3960 2735
rect 3980 2715 3985 2735
rect 3915 2685 3985 2715
rect 3915 2665 3920 2685
rect 3940 2665 3960 2685
rect 3980 2665 3985 2685
rect 3915 2635 3985 2665
rect 3915 2615 3920 2635
rect 3940 2615 3960 2635
rect 3980 2615 3985 2635
rect 3915 2585 3985 2615
rect 3915 2565 3920 2585
rect 3940 2565 3960 2585
rect 3980 2565 3985 2585
rect 3915 2535 3985 2565
rect 3915 2515 3920 2535
rect 3940 2515 3960 2535
rect 3980 2515 3985 2535
rect 3915 2485 3985 2515
rect 3915 2465 3920 2485
rect 3940 2465 3960 2485
rect 3980 2465 3985 2485
rect 3915 2435 3985 2465
rect 3915 2415 3920 2435
rect 3940 2415 3960 2435
rect 3980 2415 3985 2435
rect 3915 2405 3985 2415
rect 1005 2355 1225 2380
rect 1895 2290 2115 2320
rect 2620 2295 2640 2405
rect 2820 2340 2840 2405
rect 3020 2385 3040 2405
rect 3010 2375 3050 2385
rect 3010 2355 3020 2375
rect 3040 2355 3050 2375
rect 3010 2345 3050 2355
rect 2820 2330 2860 2340
rect 2820 2310 2830 2330
rect 2850 2310 2860 2330
rect 2820 2300 2860 2310
rect 3220 2295 3240 2405
rect 3420 2385 3440 2405
rect 3410 2375 3450 2385
rect 3410 2355 3420 2375
rect 3440 2355 3450 2375
rect 3410 2345 3450 2355
rect 3620 2340 3640 2405
rect 3760 2375 3800 2385
rect 3760 2355 3770 2375
rect 3790 2355 3800 2375
rect 3760 2345 3800 2355
rect 3600 2330 3640 2340
rect 3600 2310 3610 2330
rect 3630 2310 3640 2330
rect 3600 2300 3640 2310
rect 3820 2295 3840 2405
rect 1895 2270 1905 2290
rect 1925 2270 1950 2290
rect 1970 2270 1995 2290
rect 2015 2270 2040 2290
rect 2060 2270 2085 2290
rect 2105 2270 2115 2290
rect 1895 2260 2115 2270
rect 2610 2285 2650 2295
rect 2610 2265 2620 2285
rect 2640 2265 2650 2285
rect 2610 2255 2650 2265
rect 3210 2285 3250 2295
rect 3210 2265 3220 2285
rect 3240 2265 3250 2285
rect 3210 2255 3250 2265
rect 3810 2285 3850 2295
rect 3810 2265 3820 2285
rect 3840 2265 3850 2285
rect 3810 2255 3850 2265
rect 4375 2275 4415 2285
rect 4375 2255 4385 2275
rect 4405 2265 4555 2275
rect 4405 2255 4525 2265
rect 4375 2245 4415 2255
rect 4515 2245 4525 2255
rect 4545 2245 4555 2265
rect 2510 2225 2610 2235
rect 2510 2205 2520 2225
rect 2540 2205 2570 2225
rect 2590 2205 2610 2225
rect 2510 2195 2610 2205
rect 2710 2225 2750 2235
rect 2710 2205 2720 2225
rect 2740 2205 2750 2225
rect 2710 2195 2750 2205
rect 2910 2225 2950 2235
rect 2910 2205 2920 2225
rect 2940 2205 2950 2225
rect 2910 2195 2950 2205
rect 3110 2225 3150 2235
rect 3110 2205 3120 2225
rect 3140 2205 3150 2225
rect 3110 2195 3150 2205
rect 3310 2225 3350 2235
rect 3310 2205 3320 2225
rect 3340 2205 3350 2225
rect 3310 2195 3350 2205
rect 3510 2225 3550 2235
rect 3510 2205 3520 2225
rect 3540 2205 3550 2225
rect 3510 2195 3550 2205
rect 3710 2225 3750 2235
rect 3710 2205 3720 2225
rect 3740 2205 3750 2225
rect 3710 2195 3750 2205
rect 3860 2225 3950 2235
rect 3860 2205 3870 2225
rect 3890 2205 3920 2225
rect 3940 2205 3950 2225
rect 3860 2195 3950 2205
rect 2520 2175 2540 2195
rect 2720 2175 2740 2195
rect 2920 2175 2940 2195
rect 3120 2175 3140 2195
rect 3320 2175 3340 2195
rect 3520 2175 3540 2195
rect 3720 2175 3740 2195
rect 3920 2175 3940 2195
rect 4385 2175 4405 2245
rect 4515 2235 4555 2245
rect 4585 2225 4625 2235
rect 4585 2205 4595 2225
rect 4615 2205 4625 2225
rect 4585 2195 4625 2205
rect 4595 2175 4615 2195
rect 2475 2165 2545 2175
rect 2475 2145 2480 2165
rect 2500 2145 2520 2165
rect 2540 2145 2545 2165
rect 2475 2115 2545 2145
rect 2475 2095 2480 2115
rect 2500 2095 2520 2115
rect 2540 2095 2545 2115
rect 2475 2065 2545 2095
rect 2475 2045 2480 2065
rect 2500 2045 2520 2065
rect 2540 2045 2545 2065
rect 2475 2015 2545 2045
rect 945 2000 1005 2010
rect 945 1980 955 2000
rect 975 1980 1005 2000
rect 945 1975 1005 1980
rect 2475 1995 2480 2015
rect 2500 1995 2520 2015
rect 2540 1995 2545 2015
rect 2475 1985 2545 1995
rect 2615 2165 2645 2175
rect 2615 2145 2620 2165
rect 2640 2145 2645 2165
rect 2615 2115 2645 2145
rect 2615 2095 2620 2115
rect 2640 2095 2645 2115
rect 2615 2065 2645 2095
rect 2615 2045 2620 2065
rect 2640 2045 2645 2065
rect 2615 2015 2645 2045
rect 2615 1995 2620 2015
rect 2640 1995 2645 2015
rect 2615 1985 2645 1995
rect 2715 2165 2745 2175
rect 2715 2145 2720 2165
rect 2740 2145 2745 2165
rect 2715 2115 2745 2145
rect 2715 2095 2720 2115
rect 2740 2095 2745 2115
rect 2715 2065 2745 2095
rect 2715 2045 2720 2065
rect 2740 2045 2745 2065
rect 2715 2015 2745 2045
rect 2715 1995 2720 2015
rect 2740 1995 2745 2015
rect 2715 1985 2745 1995
rect 2815 2165 2845 2175
rect 2815 2145 2820 2165
rect 2840 2145 2845 2165
rect 2815 2115 2845 2145
rect 2815 2095 2820 2115
rect 2840 2095 2845 2115
rect 2815 2065 2845 2095
rect 2815 2045 2820 2065
rect 2840 2045 2845 2065
rect 2815 2015 2845 2045
rect 2815 1995 2820 2015
rect 2840 1995 2845 2015
rect 2815 1985 2845 1995
rect 2915 2165 2945 2175
rect 2915 2145 2920 2165
rect 2940 2145 2945 2165
rect 2915 2115 2945 2145
rect 2915 2095 2920 2115
rect 2940 2095 2945 2115
rect 2915 2065 2945 2095
rect 2915 2045 2920 2065
rect 2940 2045 2945 2065
rect 2915 2015 2945 2045
rect 2915 1995 2920 2015
rect 2940 1995 2945 2015
rect 2915 1985 2945 1995
rect 3015 2165 3045 2175
rect 3015 2145 3020 2165
rect 3040 2145 3045 2165
rect 3015 2115 3045 2145
rect 3015 2095 3020 2115
rect 3040 2095 3045 2115
rect 3015 2065 3045 2095
rect 3015 2045 3020 2065
rect 3040 2045 3045 2065
rect 3015 2015 3045 2045
rect 3015 1995 3020 2015
rect 3040 1995 3045 2015
rect 3015 1985 3045 1995
rect 3115 2165 3145 2175
rect 3115 2145 3120 2165
rect 3140 2145 3145 2165
rect 3115 2115 3145 2145
rect 3115 2095 3120 2115
rect 3140 2095 3145 2115
rect 3115 2065 3145 2095
rect 3115 2045 3120 2065
rect 3140 2045 3145 2065
rect 3115 2015 3145 2045
rect 3115 1995 3120 2015
rect 3140 1995 3145 2015
rect 3115 1985 3145 1995
rect 3215 2165 3245 2175
rect 3215 2145 3220 2165
rect 3240 2145 3245 2165
rect 3215 2115 3245 2145
rect 3215 2095 3220 2115
rect 3240 2095 3245 2115
rect 3215 2065 3245 2095
rect 3215 2045 3220 2065
rect 3240 2045 3245 2065
rect 3215 2015 3245 2045
rect 3215 1995 3220 2015
rect 3240 1995 3245 2015
rect 3215 1985 3245 1995
rect 3315 2165 3345 2175
rect 3315 2145 3320 2165
rect 3340 2145 3345 2165
rect 3315 2115 3345 2145
rect 3315 2095 3320 2115
rect 3340 2095 3345 2115
rect 3315 2065 3345 2095
rect 3315 2045 3320 2065
rect 3340 2045 3345 2065
rect 3315 2015 3345 2045
rect 3315 1995 3320 2015
rect 3340 1995 3345 2015
rect 3315 1985 3345 1995
rect 3415 2165 3445 2175
rect 3415 2145 3420 2165
rect 3440 2145 3445 2165
rect 3415 2115 3445 2145
rect 3415 2095 3420 2115
rect 3440 2095 3445 2115
rect 3415 2065 3445 2095
rect 3415 2045 3420 2065
rect 3440 2045 3445 2065
rect 3415 2015 3445 2045
rect 3415 1995 3420 2015
rect 3440 1995 3445 2015
rect 3415 1985 3445 1995
rect 3515 2165 3545 2175
rect 3515 2145 3520 2165
rect 3540 2145 3545 2165
rect 3515 2115 3545 2145
rect 3515 2095 3520 2115
rect 3540 2095 3545 2115
rect 3515 2065 3545 2095
rect 3515 2045 3520 2065
rect 3540 2045 3545 2065
rect 3515 2015 3545 2045
rect 3515 1995 3520 2015
rect 3540 1995 3545 2015
rect 3515 1985 3545 1995
rect 3615 2165 3645 2175
rect 3615 2145 3620 2165
rect 3640 2145 3645 2165
rect 3615 2115 3645 2145
rect 3615 2095 3620 2115
rect 3640 2095 3645 2115
rect 3615 2065 3645 2095
rect 3615 2045 3620 2065
rect 3640 2045 3645 2065
rect 3615 2015 3645 2045
rect 3615 1995 3620 2015
rect 3640 1995 3645 2015
rect 3615 1985 3645 1995
rect 3715 2165 3745 2175
rect 3715 2145 3720 2165
rect 3740 2145 3745 2165
rect 3715 2115 3745 2145
rect 3715 2095 3720 2115
rect 3740 2095 3745 2115
rect 3715 2065 3745 2095
rect 3715 2045 3720 2065
rect 3740 2045 3745 2065
rect 3715 2015 3745 2045
rect 3715 1995 3720 2015
rect 3740 1995 3745 2015
rect 3715 1985 3745 1995
rect 3815 2165 3845 2175
rect 3815 2145 3820 2165
rect 3840 2145 3845 2165
rect 3815 2115 3845 2145
rect 3815 2095 3820 2115
rect 3840 2095 3845 2115
rect 3815 2065 3845 2095
rect 3815 2045 3820 2065
rect 3840 2045 3845 2065
rect 3815 2015 3845 2045
rect 3815 1995 3820 2015
rect 3840 1995 3845 2015
rect 3815 1985 3845 1995
rect 3915 2165 3985 2175
rect 3915 2145 3920 2165
rect 3940 2145 3960 2165
rect 3980 2145 3985 2165
rect 3915 2115 3985 2145
rect 3915 2095 3920 2115
rect 3940 2095 3960 2115
rect 3980 2095 3985 2115
rect 3915 2065 3985 2095
rect 3915 2045 3920 2065
rect 3940 2045 3960 2065
rect 3980 2045 3985 2065
rect 3915 2015 3985 2045
rect 3915 1995 3920 2015
rect 3940 1995 3960 2015
rect 3980 1995 3985 2015
rect 3915 1985 3985 1995
rect 4380 2165 4410 2175
rect 4380 2145 4385 2165
rect 4405 2145 4410 2165
rect 4380 2115 4410 2145
rect 4380 2095 4385 2115
rect 4405 2095 4410 2115
rect 4380 2065 4410 2095
rect 4380 2045 4385 2065
rect 4405 2045 4410 2065
rect 4380 2015 4410 2045
rect 4380 1995 4385 2015
rect 4405 1995 4410 2015
rect 4380 1985 4410 1995
rect 4435 2165 4465 2175
rect 4435 2145 4440 2165
rect 4460 2145 4465 2165
rect 4435 2115 4465 2145
rect 4435 2095 4440 2115
rect 4460 2095 4465 2115
rect 4435 2065 4465 2095
rect 4435 2045 4440 2065
rect 4460 2045 4465 2065
rect 4435 2015 4465 2045
rect 4435 1995 4440 2015
rect 4460 1995 4465 2015
rect 4435 1985 4465 1995
rect 4505 2165 4535 2175
rect 4505 2145 4510 2165
rect 4530 2145 4535 2165
rect 4505 2115 4535 2145
rect 4505 2095 4510 2115
rect 4530 2095 4535 2115
rect 4505 2065 4535 2095
rect 4505 2045 4510 2065
rect 4530 2045 4535 2065
rect 4505 2015 4535 2045
rect 4505 1995 4510 2015
rect 4530 1995 4535 2015
rect 4505 1985 4535 1995
rect 4560 2165 4615 2175
rect 4560 2145 4565 2165
rect 4585 2145 4615 2165
rect 4560 2115 4595 2145
rect 4560 2095 4565 2115
rect 4585 2095 4595 2115
rect 4560 2065 4595 2095
rect 4560 2045 4565 2065
rect 4585 2045 4595 2065
rect 4560 2015 4595 2045
rect 4560 1995 4565 2015
rect 4585 1995 4595 2015
rect 4560 1985 4595 1995
rect 945 1970 985 1975
rect 1895 1950 2115 1975
rect 1005 1890 1225 1915
rect 2620 1860 2640 1985
rect 2820 1960 2840 1985
rect 2810 1950 2850 1960
rect 2810 1930 2820 1950
rect 2840 1930 2850 1950
rect 2810 1920 2850 1930
rect 3020 1915 3040 1985
rect 2660 1905 2700 1915
rect 2660 1885 2670 1905
rect 2690 1885 2700 1905
rect 2660 1875 2700 1885
rect 3010 1905 3050 1915
rect 3010 1885 3020 1905
rect 3040 1885 3050 1905
rect 3010 1875 3050 1885
rect 3160 1905 3200 1915
rect 3160 1885 3170 1905
rect 3190 1885 3200 1905
rect 3160 1875 3200 1885
rect 3220 1860 3240 1985
rect 3420 1915 3440 1985
rect 3620 1960 3640 1985
rect 3610 1950 3650 1960
rect 3610 1930 3620 1950
rect 3640 1930 3650 1950
rect 3610 1920 3650 1930
rect 3260 1905 3300 1915
rect 3260 1885 3270 1905
rect 3290 1885 3300 1905
rect 3260 1875 3300 1885
rect 3410 1905 3450 1915
rect 3410 1885 3420 1905
rect 3440 1885 3450 1905
rect 3410 1875 3450 1885
rect 3760 1905 3800 1915
rect 3760 1885 3770 1905
rect 3790 1885 3800 1905
rect 3760 1875 3800 1885
rect 3820 1860 3840 1985
rect 1895 1830 2115 1855
rect 2610 1850 2650 1860
rect 2610 1830 2620 1850
rect 2640 1830 2650 1850
rect 2610 1820 2650 1830
rect 3210 1850 3250 1860
rect 3210 1830 3220 1850
rect 3240 1830 3250 1850
rect 3210 1820 3250 1830
rect 3810 1850 3850 1860
rect 3810 1830 3820 1850
rect 3840 1830 3850 1850
rect 3810 1820 3850 1830
rect 1005 1770 1225 1795
rect 2810 1790 2850 1800
rect 2810 1770 2820 1790
rect 2840 1770 2850 1790
rect 2810 1760 2850 1770
rect 3210 1790 3250 1800
rect 3210 1770 3220 1790
rect 3240 1770 3250 1790
rect 3210 1760 3250 1770
rect 3610 1790 3650 1800
rect 3610 1770 3620 1790
rect 3640 1770 3650 1790
rect 3610 1760 3650 1770
rect 1895 1705 2115 1735
rect 1895 1685 1905 1705
rect 1925 1685 1950 1705
rect 1970 1685 1995 1705
rect 2015 1685 2040 1705
rect 2060 1685 2085 1705
rect 2105 1685 2115 1705
rect 1895 1675 2115 1685
rect 2820 1655 2840 1760
rect 3010 1745 3050 1755
rect 3010 1725 3020 1745
rect 3040 1725 3050 1745
rect 3010 1715 3050 1725
rect 2860 1700 2900 1710
rect 2860 1680 2870 1700
rect 2890 1680 2900 1700
rect 2860 1670 2900 1680
rect 3020 1655 3040 1715
rect 3160 1700 3200 1710
rect 3160 1680 3170 1700
rect 3190 1680 3200 1700
rect 3160 1670 3200 1680
rect 3220 1655 3240 1760
rect 3410 1745 3450 1755
rect 3410 1725 3420 1745
rect 3440 1725 3450 1745
rect 3410 1715 3450 1725
rect 3260 1700 3300 1710
rect 3260 1680 3270 1700
rect 3290 1680 3300 1700
rect 3260 1670 3300 1680
rect 3420 1655 3440 1715
rect 3560 1700 3600 1710
rect 3560 1680 3570 1700
rect 3590 1680 3600 1700
rect 3560 1670 3600 1680
rect 3620 1655 3640 1760
rect 4440 1710 4460 1985
rect 4505 1950 4525 1985
rect 4485 1940 4525 1950
rect 4485 1920 4495 1940
rect 4515 1920 4525 1940
rect 4485 1910 4525 1920
rect 4430 1700 4470 1710
rect 4430 1680 4440 1700
rect 4460 1680 4470 1700
rect 4430 1670 4470 1680
rect 2715 1645 2745 1655
rect 2715 1630 2720 1645
rect 2675 1625 2720 1630
rect 2740 1625 2745 1645
rect 2675 1620 2745 1625
rect 2675 1600 2685 1620
rect 2705 1600 2745 1620
rect 2675 1595 2745 1600
rect 2675 1590 2720 1595
rect 2715 1575 2720 1590
rect 2740 1575 2745 1595
rect 2715 1565 2745 1575
rect 2815 1645 2845 1655
rect 2815 1625 2820 1645
rect 2840 1625 2845 1645
rect 2815 1595 2845 1625
rect 2815 1575 2820 1595
rect 2840 1575 2845 1595
rect 2815 1565 2845 1575
rect 2915 1645 2945 1655
rect 2915 1625 2920 1645
rect 2940 1625 2945 1645
rect 2915 1595 2945 1625
rect 2915 1575 2920 1595
rect 2940 1575 2945 1595
rect 2915 1565 2945 1575
rect 3015 1645 3045 1655
rect 3015 1625 3020 1645
rect 3040 1625 3045 1645
rect 3015 1595 3045 1625
rect 3015 1575 3020 1595
rect 3040 1575 3045 1595
rect 3015 1565 3045 1575
rect 3115 1645 3145 1655
rect 3115 1625 3120 1645
rect 3140 1625 3145 1645
rect 3115 1595 3145 1625
rect 3115 1575 3120 1595
rect 3140 1575 3145 1595
rect 3115 1565 3145 1575
rect 3215 1645 3245 1655
rect 3215 1625 3220 1645
rect 3240 1625 3245 1645
rect 3215 1595 3245 1625
rect 3215 1575 3220 1595
rect 3240 1575 3245 1595
rect 3215 1565 3245 1575
rect 3315 1645 3345 1655
rect 3315 1625 3320 1645
rect 3340 1625 3345 1645
rect 3315 1595 3345 1625
rect 3315 1575 3320 1595
rect 3340 1575 3345 1595
rect 3315 1565 3345 1575
rect 3415 1645 3445 1655
rect 3415 1625 3420 1645
rect 3440 1625 3445 1645
rect 3415 1595 3445 1625
rect 3415 1575 3420 1595
rect 3440 1575 3445 1595
rect 3415 1565 3445 1575
rect 3515 1645 3545 1655
rect 3515 1625 3520 1645
rect 3540 1625 3545 1645
rect 3515 1595 3545 1625
rect 3515 1575 3520 1595
rect 3540 1575 3545 1595
rect 3515 1565 3545 1575
rect 3615 1645 3645 1655
rect 3615 1625 3620 1645
rect 3640 1625 3645 1645
rect 3615 1595 3645 1625
rect 3615 1575 3620 1595
rect 3640 1575 3645 1595
rect 3615 1565 3645 1575
rect 3715 1645 3745 1655
rect 3715 1625 3720 1645
rect 3740 1625 3745 1645
rect 3715 1595 3745 1625
rect 3715 1575 3720 1595
rect 3740 1575 3745 1595
rect 3715 1565 3745 1575
rect 2720 1540 2740 1565
rect 2760 1540 2800 1550
rect 945 1530 1005 1540
rect 945 1510 955 1530
rect 975 1510 1005 1530
rect 945 1505 1005 1510
rect 1795 1530 2115 1540
rect 1795 1510 1905 1530
rect 1925 1510 1950 1530
rect 1970 1510 1995 1530
rect 2015 1510 2040 1530
rect 2060 1510 2085 1530
rect 2105 1510 2115 1530
rect 2720 1520 2770 1540
rect 2790 1520 2800 1540
rect 2760 1510 2800 1520
rect 1795 1505 2115 1510
rect 945 1500 985 1505
rect 1895 1480 2115 1505
rect 2920 1500 2940 1565
rect 3010 1535 3050 1545
rect 3010 1515 3020 1535
rect 3040 1515 3050 1535
rect 3010 1505 3050 1515
rect 3120 1500 3140 1565
rect 3320 1500 3340 1565
rect 3410 1535 3450 1545
rect 3410 1515 3420 1535
rect 3440 1515 3450 1535
rect 3410 1505 3450 1515
rect 3520 1500 3540 1565
rect 3660 1540 3700 1550
rect 3720 1540 3740 1565
rect 3660 1520 3670 1540
rect 3690 1520 3740 1540
rect 3660 1510 3700 1520
rect 2910 1490 2950 1500
rect 2910 1470 2920 1490
rect 2940 1470 2950 1490
rect 2910 1460 2950 1470
rect 3110 1490 3150 1500
rect 3110 1470 3120 1490
rect 3140 1470 3150 1490
rect 3110 1460 3150 1470
rect 3310 1490 3350 1500
rect 3310 1470 3320 1490
rect 3340 1470 3350 1490
rect 3310 1460 3350 1470
rect 3510 1490 3550 1500
rect 3510 1470 3520 1490
rect 3540 1470 3550 1490
rect 3510 1460 3550 1470
rect 1005 1420 1225 1445
rect 2920 1440 2940 1460
rect 3120 1440 3140 1460
rect 2735 1430 3170 1440
rect 1895 1360 2115 1385
rect 2735 1410 2780 1430
rect 2800 1410 2820 1430
rect 2840 1410 2860 1430
rect 2880 1410 2900 1430
rect 2920 1410 2940 1430
rect 2960 1410 2980 1430
rect 3000 1410 3020 1430
rect 3040 1410 3060 1430
rect 3080 1410 3100 1430
rect 3120 1410 3140 1430
rect 3160 1410 3170 1430
rect 2735 1400 3170 1410
rect 3290 1430 3730 1440
rect 3290 1410 3300 1430
rect 3320 1410 3340 1430
rect 3360 1410 3380 1430
rect 3400 1410 3420 1430
rect 3440 1410 3460 1430
rect 3480 1410 3500 1430
rect 3520 1410 3540 1430
rect 3560 1410 3580 1430
rect 3600 1410 3620 1430
rect 3640 1410 3660 1430
rect 3680 1410 3700 1430
rect 3720 1410 3730 1430
rect 3290 1400 3730 1410
rect 2735 1370 2765 1400
rect 2735 1350 2740 1370
rect 2760 1350 2765 1370
rect 1005 1300 1225 1325
rect 2735 1320 2765 1350
rect 2735 1300 2740 1320
rect 2760 1300 2765 1320
rect 945 1240 985 1245
rect 1895 1240 2115 1265
rect 945 1235 1005 1240
rect 945 1215 955 1235
rect 975 1215 1005 1235
rect 945 1205 1005 1215
rect 2735 1270 2765 1300
rect 2735 1250 2740 1270
rect 2760 1250 2765 1270
rect 2735 1220 2765 1250
rect 2735 1200 2740 1220
rect 2760 1200 2765 1220
rect 2735 1170 2765 1200
rect 2735 1150 2740 1170
rect 2760 1150 2765 1170
rect 2735 1120 2765 1150
rect 2735 1100 2740 1120
rect 2760 1100 2765 1120
rect 2735 1070 2765 1100
rect 2735 1050 2740 1070
rect 2760 1050 2765 1070
rect 2735 1020 2765 1050
rect 2735 1000 2740 1020
rect 2760 1000 2765 1020
rect 2735 990 2765 1000
rect 3175 1370 3285 1380
rect 3175 1350 3180 1370
rect 3200 1350 3220 1370
rect 3240 1350 3260 1370
rect 3280 1350 3285 1370
rect 3175 1320 3285 1350
rect 3175 1300 3180 1320
rect 3200 1300 3220 1320
rect 3240 1300 3260 1320
rect 3280 1300 3285 1320
rect 3175 1270 3285 1300
rect 3175 1250 3180 1270
rect 3200 1250 3220 1270
rect 3240 1250 3260 1270
rect 3280 1250 3285 1270
rect 3175 1220 3285 1250
rect 3175 1200 3180 1220
rect 3200 1200 3220 1220
rect 3240 1200 3260 1220
rect 3280 1200 3285 1220
rect 3175 1170 3285 1200
rect 3175 1150 3180 1170
rect 3200 1150 3220 1170
rect 3240 1150 3260 1170
rect 3280 1150 3285 1170
rect 3175 1120 3285 1150
rect 3175 1100 3180 1120
rect 3200 1100 3220 1120
rect 3240 1100 3260 1120
rect 3280 1100 3285 1120
rect 3175 1070 3285 1100
rect 3175 1050 3180 1070
rect 3200 1050 3220 1070
rect 3240 1050 3260 1070
rect 3280 1050 3285 1070
rect 3175 1020 3285 1050
rect 3175 1000 3180 1020
rect 3200 1000 3220 1020
rect 3240 1000 3260 1020
rect 3280 1000 3285 1020
rect 3175 990 3285 1000
rect 3695 1370 3725 1400
rect 3695 1350 3700 1370
rect 3720 1350 3725 1370
rect 3695 1320 3725 1350
rect 3695 1300 3700 1320
rect 3720 1300 3725 1320
rect 3695 1270 3725 1300
rect 3695 1250 3700 1270
rect 3720 1250 3725 1270
rect 3695 1220 3725 1250
rect 3695 1200 3700 1220
rect 3720 1200 3725 1220
rect 3695 1170 3725 1200
rect 3695 1150 3700 1170
rect 3720 1150 3725 1170
rect 3695 1120 3725 1150
rect 3695 1100 3700 1120
rect 3720 1100 3725 1120
rect 3695 1070 3725 1100
rect 3695 1050 3700 1070
rect 3720 1050 3725 1070
rect 3695 1020 3725 1050
rect 3695 1000 3700 1020
rect 3720 1000 3725 1020
rect 3695 990 3725 1000
rect 3180 970 3200 990
rect 3220 970 3240 990
rect 3260 970 3280 990
rect 3170 960 3290 970
rect 3170 940 3180 960
rect 3200 940 3220 960
rect 3240 940 3260 960
rect 3280 940 3290 960
rect 3170 930 3290 940
rect 2690 900 3760 910
rect 2690 880 2730 900
rect 2750 880 2810 900
rect 2830 880 2890 900
rect 2910 880 2970 900
rect 2990 880 3050 900
rect 3070 880 3130 900
rect 3150 880 3210 900
rect 3230 880 3290 900
rect 3310 880 3370 900
rect 3390 880 3450 900
rect 3470 880 3530 900
rect 3550 880 3610 900
rect 3630 880 3690 900
rect 3710 880 3730 900
rect 3750 880 3760 900
rect 2690 870 3760 880
rect 2690 850 2710 870
rect 2685 840 2715 850
rect 650 820 690 830
rect 650 800 660 820
rect 680 800 690 820
rect 650 770 690 800
rect 650 750 660 770
rect 680 750 690 770
rect 2685 820 2690 840
rect 2710 820 2715 840
rect 2685 790 2715 820
rect 2685 770 2690 790
rect 2710 770 2715 790
rect 2685 760 2715 770
rect 3725 840 3795 850
rect 3725 820 3730 840
rect 3750 820 3770 840
rect 3790 825 3795 840
rect 3790 820 3835 825
rect 3725 815 3835 820
rect 3725 795 3805 815
rect 3825 795 3835 815
rect 3725 790 3835 795
rect 3725 770 3730 790
rect 3750 770 3770 790
rect 3790 785 3835 790
rect 3790 770 3795 785
rect 3725 760 3795 770
rect 650 720 690 750
rect 650 700 660 720
rect 680 700 690 720
rect 650 660 690 700
rect 5 535 4740 660
rect 650 10 690 535
rect 1330 10 1370 535
rect 2010 10 2050 535
rect 2690 10 2730 535
rect 3370 10 3410 535
rect 4050 10 4090 535
<< viali >>
rect 2520 2825 2540 2845
rect 2720 2825 2740 2845
rect 2920 2825 2940 2845
rect 3120 2825 3140 2845
rect 3220 2825 3240 2845
rect 3320 2825 3340 2845
rect 3520 2825 3540 2845
rect 3720 2825 3740 2845
rect 3920 2825 3940 2845
rect 955 2565 975 2585
rect 3020 2355 3040 2375
rect 2830 2310 2850 2330
rect 3420 2355 3440 2375
rect 3770 2355 3790 2375
rect 3610 2310 3630 2330
rect 1905 2270 1925 2290
rect 1950 2270 1970 2290
rect 1995 2270 2015 2290
rect 2040 2270 2060 2290
rect 2085 2270 2105 2290
rect 2620 2265 2640 2285
rect 3220 2265 3240 2285
rect 3820 2265 3840 2285
rect 4385 2255 4405 2275
rect 2520 2205 2540 2225
rect 2720 2205 2740 2225
rect 2920 2205 2940 2225
rect 3120 2205 3140 2225
rect 3320 2205 3340 2225
rect 3520 2205 3540 2225
rect 3720 2205 3740 2225
rect 3920 2205 3940 2225
rect 4595 2205 4615 2225
rect 955 1980 975 2000
rect 2820 1930 2840 1950
rect 2670 1885 2690 1905
rect 3020 1885 3040 1905
rect 3170 1885 3190 1905
rect 3620 1930 3640 1950
rect 3270 1885 3290 1905
rect 3420 1885 3440 1905
rect 3770 1885 3790 1905
rect 2620 1830 2640 1850
rect 3220 1830 3240 1850
rect 3820 1830 3840 1850
rect 2820 1770 2840 1790
rect 3220 1770 3240 1790
rect 3620 1770 3640 1790
rect 1905 1685 1925 1705
rect 1950 1685 1970 1705
rect 1995 1685 2015 1705
rect 2040 1685 2060 1705
rect 2085 1685 2105 1705
rect 3020 1725 3040 1745
rect 2870 1680 2890 1700
rect 3170 1680 3190 1700
rect 3420 1725 3440 1745
rect 3270 1680 3290 1700
rect 3570 1680 3590 1700
rect 4495 1920 4515 1940
rect 4440 1680 4460 1700
rect 2685 1600 2705 1620
rect 955 1510 975 1530
rect 1905 1510 1925 1530
rect 1950 1510 1970 1530
rect 1995 1510 2015 1530
rect 2040 1510 2060 1530
rect 2085 1510 2105 1530
rect 3020 1515 3040 1535
rect 3420 1515 3440 1535
rect 3670 1520 3690 1540
rect 2920 1470 2940 1490
rect 3120 1470 3140 1490
rect 3320 1470 3340 1490
rect 3520 1470 3540 1490
rect 3700 1410 3720 1430
rect 955 1215 975 1235
rect 3180 940 3200 960
rect 3220 940 3240 960
rect 3260 940 3280 960
rect 3730 880 3750 900
rect 660 800 680 820
rect 3805 795 3825 815
<< metal1 >>
rect 3220 2855 3240 3165
rect 2510 2850 2550 2855
rect 2510 2820 2515 2850
rect 2545 2820 2550 2850
rect 2510 2815 2550 2820
rect 2710 2850 2750 2855
rect 2710 2820 2715 2850
rect 2745 2820 2750 2850
rect 2710 2815 2750 2820
rect 2910 2850 2950 2855
rect 2910 2820 2915 2850
rect 2945 2820 2950 2850
rect 2910 2815 2950 2820
rect 3110 2850 3150 2855
rect 3110 2820 3115 2850
rect 3145 2820 3150 2850
rect 3110 2815 3150 2820
rect 3210 2845 3250 2855
rect 3210 2825 3220 2845
rect 3240 2825 3250 2845
rect 3210 2815 3250 2825
rect 3310 2850 3350 2855
rect 3310 2820 3315 2850
rect 3345 2820 3350 2850
rect 3310 2815 3350 2820
rect 3510 2850 3550 2855
rect 3510 2820 3515 2850
rect 3545 2820 3550 2850
rect 3510 2815 3550 2820
rect 3710 2850 3750 2855
rect 3710 2820 3715 2850
rect 3745 2820 3750 2850
rect 3710 2815 3750 2820
rect 3910 2850 3950 2855
rect 3910 2820 3915 2850
rect 3945 2820 3950 2850
rect 3910 2815 3950 2820
rect 945 2590 985 2595
rect 945 2560 950 2590
rect 980 2560 985 2590
rect 945 2555 985 2560
rect 2150 2380 2190 2385
rect 2150 2350 2155 2380
rect 2185 2350 2190 2380
rect 2150 2345 2190 2350
rect 3010 2380 3050 2385
rect 3010 2350 3015 2380
rect 3045 2350 3050 2380
rect 3010 2345 3050 2350
rect 3410 2380 3450 2385
rect 3410 2350 3415 2380
rect 3445 2350 3450 2380
rect 3410 2345 3450 2350
rect 3760 2380 3800 2385
rect 3760 2350 3765 2380
rect 3795 2350 3800 2380
rect 3760 2345 3800 2350
rect 4375 2380 4415 2385
rect 4375 2350 4380 2380
rect 4410 2350 4415 2380
rect 4375 2345 4415 2350
rect 1895 2295 2115 2300
rect 1895 2265 1900 2295
rect 2110 2265 2115 2295
rect 1895 2260 2115 2265
rect 945 2005 985 2010
rect 945 1975 950 2005
rect 980 1975 985 2005
rect 945 1970 985 1975
rect 465 1710 505 1715
rect 465 1680 470 1710
rect 500 1680 505 1710
rect 465 725 505 1680
rect 1895 1710 2115 1715
rect 2160 1710 2180 2345
rect 2295 2335 2335 2340
rect 2295 2305 2300 2335
rect 2330 2305 2335 2335
rect 2295 2300 2335 2305
rect 2820 2335 2860 2340
rect 2820 2305 2825 2335
rect 2855 2305 2860 2335
rect 2820 2300 2860 2305
rect 3600 2335 3640 2340
rect 3600 2305 3605 2335
rect 3635 2305 3640 2335
rect 3600 2300 3640 2305
rect 1895 1680 1900 1710
rect 2110 1680 2115 1710
rect 1895 1675 2115 1680
rect 2150 1705 2190 1710
rect 2150 1675 2155 1705
rect 2185 1675 2190 1705
rect 2150 1670 2190 1675
rect 2305 1545 2325 2300
rect 2610 2290 2650 2295
rect 2610 2260 2615 2290
rect 2645 2260 2650 2290
rect 2610 2255 2650 2260
rect 3210 2290 3250 2295
rect 3210 2260 3215 2290
rect 3245 2260 3250 2290
rect 3210 2255 3250 2260
rect 3810 2290 3850 2295
rect 3810 2260 3815 2290
rect 3845 2260 3850 2290
rect 4385 2285 4405 2345
rect 3810 2255 3850 2260
rect 4375 2275 4415 2285
rect 4375 2255 4385 2275
rect 4405 2255 4415 2275
rect 4375 2245 4415 2255
rect 2510 2230 2550 2235
rect 2510 2200 2515 2230
rect 2545 2200 2550 2230
rect 2510 2195 2550 2200
rect 2710 2230 2750 2235
rect 2710 2200 2715 2230
rect 2745 2200 2750 2230
rect 2710 2195 2750 2200
rect 2910 2230 2950 2235
rect 2910 2200 2915 2230
rect 2945 2200 2950 2230
rect 2910 2195 2950 2200
rect 3110 2230 3150 2235
rect 3110 2200 3115 2230
rect 3145 2200 3150 2230
rect 3110 2195 3150 2200
rect 3310 2230 3350 2235
rect 3310 2200 3315 2230
rect 3345 2200 3350 2230
rect 3310 2195 3350 2200
rect 3510 2230 3550 2235
rect 3510 2200 3515 2230
rect 3545 2200 3550 2230
rect 3510 2195 3550 2200
rect 3710 2230 3750 2235
rect 3710 2200 3715 2230
rect 3745 2200 3750 2230
rect 3710 2195 3750 2200
rect 3910 2230 3950 2235
rect 3910 2200 3915 2230
rect 3945 2200 3950 2230
rect 3910 2195 3950 2200
rect 4585 2230 4625 2235
rect 4585 2200 4590 2230
rect 4620 2200 4625 2230
rect 4585 2195 4625 2200
rect 2810 1955 2850 1960
rect 2810 1925 2815 1955
rect 2845 1925 2850 1955
rect 2810 1920 2850 1925
rect 3610 1955 3650 1960
rect 3610 1925 3615 1955
rect 3645 1925 3650 1955
rect 3610 1920 3650 1925
rect 4485 1940 4525 1950
rect 4485 1920 4495 1940
rect 4515 1920 4525 1940
rect 2660 1910 2700 1915
rect 2660 1880 2665 1910
rect 2695 1880 2700 1910
rect 2660 1875 2700 1880
rect 2610 1855 2650 1860
rect 2610 1825 2615 1855
rect 2645 1825 2650 1855
rect 2610 1820 2650 1825
rect 2820 1800 2840 1920
rect 3010 1910 3050 1915
rect 3010 1880 3015 1910
rect 3045 1880 3050 1910
rect 3010 1875 3050 1880
rect 3160 1910 3200 1915
rect 3160 1880 3165 1910
rect 3195 1880 3200 1910
rect 3160 1875 3200 1880
rect 3260 1910 3300 1915
rect 3260 1880 3265 1910
rect 3295 1880 3300 1910
rect 3260 1875 3300 1880
rect 3410 1910 3450 1915
rect 3410 1880 3415 1910
rect 3445 1880 3450 1910
rect 3410 1875 3450 1880
rect 3760 1910 3800 1915
rect 4485 1910 4525 1920
rect 3760 1880 3765 1910
rect 3795 1880 3800 1910
rect 3760 1875 3800 1880
rect 3210 1855 3250 1860
rect 3210 1825 3215 1855
rect 3245 1825 3250 1855
rect 3210 1820 3250 1825
rect 2810 1795 2850 1800
rect 2810 1765 2815 1795
rect 2845 1765 2850 1795
rect 2810 1760 2850 1765
rect 3210 1795 3250 1800
rect 3210 1765 3215 1795
rect 3245 1765 3250 1795
rect 3210 1760 3250 1765
rect 3420 1755 3440 1875
rect 3810 1855 3850 1860
rect 3810 1825 3815 1855
rect 3845 1825 3850 1855
rect 3810 1820 3850 1825
rect 3610 1795 3650 1800
rect 3610 1765 3615 1795
rect 3645 1765 3650 1795
rect 3610 1760 3650 1765
rect 3010 1750 3050 1755
rect 3010 1720 3015 1750
rect 3045 1720 3050 1750
rect 3010 1715 3050 1720
rect 3410 1750 3450 1755
rect 3410 1720 3415 1750
rect 3445 1720 3450 1750
rect 3410 1715 3450 1720
rect 2860 1705 2900 1710
rect 2860 1675 2865 1705
rect 2895 1675 2900 1705
rect 2860 1670 2900 1675
rect 3160 1705 3200 1710
rect 3160 1675 3165 1705
rect 3195 1675 3200 1705
rect 3160 1670 3200 1675
rect 3260 1705 3300 1710
rect 3260 1675 3265 1705
rect 3295 1675 3300 1705
rect 3260 1670 3300 1675
rect 3560 1705 3600 1710
rect 3560 1675 3565 1705
rect 3595 1675 3600 1705
rect 3560 1670 3600 1675
rect 2675 1625 2715 1630
rect 2675 1595 2680 1625
rect 2710 1595 2715 1625
rect 2675 1590 2715 1595
rect 3660 1545 3700 1550
rect 2295 1540 2335 1545
rect 835 1535 875 1540
rect 835 1505 840 1535
rect 870 1505 875 1535
rect 650 825 690 830
rect 650 795 655 825
rect 685 795 690 825
rect 650 790 690 795
rect 155 160 505 725
rect 835 725 875 1505
rect 945 1535 985 1540
rect 945 1505 950 1535
rect 980 1505 985 1535
rect 945 1500 985 1505
rect 1895 1535 2115 1540
rect 1895 1505 1900 1535
rect 2110 1505 2115 1535
rect 2295 1510 2300 1540
rect 2330 1510 2335 1540
rect 2295 1505 2335 1510
rect 3010 1540 3050 1545
rect 3010 1510 3015 1540
rect 3045 1510 3050 1540
rect 3010 1505 3050 1510
rect 3410 1540 3450 1545
rect 3410 1510 3415 1540
rect 3445 1510 3450 1540
rect 3660 1515 3665 1545
rect 3695 1515 3700 1545
rect 3660 1510 3700 1515
rect 3410 1505 3450 1510
rect 1895 1500 2115 1505
rect 2910 1495 2950 1500
rect 2910 1465 2915 1495
rect 2945 1465 2950 1495
rect 2910 1460 2950 1465
rect 3110 1495 3150 1500
rect 3110 1465 3115 1495
rect 3145 1465 3150 1495
rect 3110 1460 3150 1465
rect 3310 1495 3350 1500
rect 3310 1465 3315 1495
rect 3345 1465 3350 1495
rect 3310 1460 3350 1465
rect 3510 1495 3550 1500
rect 3510 1465 3515 1495
rect 3545 1465 3550 1495
rect 3510 1460 3550 1465
rect 3820 1440 3840 1820
rect 4430 1705 4470 1710
rect 4430 1675 4435 1705
rect 4465 1675 4470 1705
rect 4430 1670 4470 1675
rect 3690 1435 3730 1440
rect 3690 1405 3695 1435
rect 3725 1405 3730 1435
rect 3690 1400 3730 1405
rect 3810 1435 3850 1440
rect 3810 1405 3815 1435
rect 3845 1405 3850 1435
rect 3810 1400 3850 1405
rect 945 1240 985 1245
rect 945 1210 950 1240
rect 980 1210 985 1240
rect 945 1205 985 1210
rect 3170 965 3290 970
rect 3170 935 3175 965
rect 3205 935 3215 965
rect 3245 935 3255 965
rect 3285 935 3290 965
rect 3170 930 3290 935
rect 4505 910 4525 1910
rect 3720 905 3760 910
rect 3720 875 3725 905
rect 3755 875 3760 905
rect 3720 870 3760 875
rect 4495 905 4535 910
rect 4495 875 4500 905
rect 4530 875 4535 905
rect 4495 870 4535 875
rect 3795 820 3835 825
rect 3795 790 3800 820
rect 3830 790 3835 820
rect 3795 785 3835 790
rect 835 690 4585 725
rect 835 160 1185 690
rect 1515 160 1865 690
rect 2195 160 2545 690
rect 2875 160 3225 690
rect 3555 160 3905 690
rect 4235 160 4585 690
<< via1 >>
rect 2515 2845 2545 2850
rect 2515 2825 2520 2845
rect 2520 2825 2540 2845
rect 2540 2825 2545 2845
rect 2515 2820 2545 2825
rect 2715 2845 2745 2850
rect 2715 2825 2720 2845
rect 2720 2825 2740 2845
rect 2740 2825 2745 2845
rect 2715 2820 2745 2825
rect 2915 2845 2945 2850
rect 2915 2825 2920 2845
rect 2920 2825 2940 2845
rect 2940 2825 2945 2845
rect 2915 2820 2945 2825
rect 3115 2845 3145 2850
rect 3115 2825 3120 2845
rect 3120 2825 3140 2845
rect 3140 2825 3145 2845
rect 3115 2820 3145 2825
rect 3315 2845 3345 2850
rect 3315 2825 3320 2845
rect 3320 2825 3340 2845
rect 3340 2825 3345 2845
rect 3315 2820 3345 2825
rect 3515 2845 3545 2850
rect 3515 2825 3520 2845
rect 3520 2825 3540 2845
rect 3540 2825 3545 2845
rect 3515 2820 3545 2825
rect 3715 2845 3745 2850
rect 3715 2825 3720 2845
rect 3720 2825 3740 2845
rect 3740 2825 3745 2845
rect 3715 2820 3745 2825
rect 3915 2845 3945 2850
rect 3915 2825 3920 2845
rect 3920 2825 3940 2845
rect 3940 2825 3945 2845
rect 3915 2820 3945 2825
rect 950 2585 980 2590
rect 950 2565 955 2585
rect 955 2565 975 2585
rect 975 2565 980 2585
rect 950 2560 980 2565
rect 2155 2350 2185 2380
rect 3015 2375 3045 2380
rect 3015 2355 3020 2375
rect 3020 2355 3040 2375
rect 3040 2355 3045 2375
rect 3015 2350 3045 2355
rect 3415 2375 3445 2380
rect 3415 2355 3420 2375
rect 3420 2355 3440 2375
rect 3440 2355 3445 2375
rect 3415 2350 3445 2355
rect 3765 2375 3795 2380
rect 3765 2355 3770 2375
rect 3770 2355 3790 2375
rect 3790 2355 3795 2375
rect 3765 2350 3795 2355
rect 4380 2350 4410 2380
rect 1900 2290 2110 2295
rect 1900 2270 1905 2290
rect 1905 2270 1925 2290
rect 1925 2270 1950 2290
rect 1950 2270 1970 2290
rect 1970 2270 1995 2290
rect 1995 2270 2015 2290
rect 2015 2270 2040 2290
rect 2040 2270 2060 2290
rect 2060 2270 2085 2290
rect 2085 2270 2105 2290
rect 2105 2270 2110 2290
rect 1900 2265 2110 2270
rect 950 2000 980 2005
rect 950 1980 955 2000
rect 955 1980 975 2000
rect 975 1980 980 2000
rect 950 1975 980 1980
rect 470 1680 500 1710
rect 2300 2305 2330 2335
rect 2825 2330 2855 2335
rect 2825 2310 2830 2330
rect 2830 2310 2850 2330
rect 2850 2310 2855 2330
rect 2825 2305 2855 2310
rect 3605 2330 3635 2335
rect 3605 2310 3610 2330
rect 3610 2310 3630 2330
rect 3630 2310 3635 2330
rect 3605 2305 3635 2310
rect 1900 1705 2110 1710
rect 1900 1685 1905 1705
rect 1905 1685 1925 1705
rect 1925 1685 1950 1705
rect 1950 1685 1970 1705
rect 1970 1685 1995 1705
rect 1995 1685 2015 1705
rect 2015 1685 2040 1705
rect 2040 1685 2060 1705
rect 2060 1685 2085 1705
rect 2085 1685 2105 1705
rect 2105 1685 2110 1705
rect 1900 1680 2110 1685
rect 2155 1675 2185 1705
rect 2615 2285 2645 2290
rect 2615 2265 2620 2285
rect 2620 2265 2640 2285
rect 2640 2265 2645 2285
rect 2615 2260 2645 2265
rect 3215 2285 3245 2290
rect 3215 2265 3220 2285
rect 3220 2265 3240 2285
rect 3240 2265 3245 2285
rect 3215 2260 3245 2265
rect 3815 2285 3845 2290
rect 3815 2265 3820 2285
rect 3820 2265 3840 2285
rect 3840 2265 3845 2285
rect 3815 2260 3845 2265
rect 2515 2225 2545 2230
rect 2515 2205 2520 2225
rect 2520 2205 2540 2225
rect 2540 2205 2545 2225
rect 2515 2200 2545 2205
rect 2715 2225 2745 2230
rect 2715 2205 2720 2225
rect 2720 2205 2740 2225
rect 2740 2205 2745 2225
rect 2715 2200 2745 2205
rect 2915 2225 2945 2230
rect 2915 2205 2920 2225
rect 2920 2205 2940 2225
rect 2940 2205 2945 2225
rect 2915 2200 2945 2205
rect 3115 2225 3145 2230
rect 3115 2205 3120 2225
rect 3120 2205 3140 2225
rect 3140 2205 3145 2225
rect 3115 2200 3145 2205
rect 3315 2225 3345 2230
rect 3315 2205 3320 2225
rect 3320 2205 3340 2225
rect 3340 2205 3345 2225
rect 3315 2200 3345 2205
rect 3515 2225 3545 2230
rect 3515 2205 3520 2225
rect 3520 2205 3540 2225
rect 3540 2205 3545 2225
rect 3515 2200 3545 2205
rect 3715 2225 3745 2230
rect 3715 2205 3720 2225
rect 3720 2205 3740 2225
rect 3740 2205 3745 2225
rect 3715 2200 3745 2205
rect 3915 2225 3945 2230
rect 3915 2205 3920 2225
rect 3920 2205 3940 2225
rect 3940 2205 3945 2225
rect 3915 2200 3945 2205
rect 4590 2225 4620 2230
rect 4590 2205 4595 2225
rect 4595 2205 4615 2225
rect 4615 2205 4620 2225
rect 4590 2200 4620 2205
rect 2815 1950 2845 1955
rect 2815 1930 2820 1950
rect 2820 1930 2840 1950
rect 2840 1930 2845 1950
rect 2815 1925 2845 1930
rect 3615 1950 3645 1955
rect 3615 1930 3620 1950
rect 3620 1930 3640 1950
rect 3640 1930 3645 1950
rect 3615 1925 3645 1930
rect 2665 1905 2695 1910
rect 2665 1885 2670 1905
rect 2670 1885 2690 1905
rect 2690 1885 2695 1905
rect 2665 1880 2695 1885
rect 2615 1850 2645 1855
rect 2615 1830 2620 1850
rect 2620 1830 2640 1850
rect 2640 1830 2645 1850
rect 2615 1825 2645 1830
rect 3015 1905 3045 1910
rect 3015 1885 3020 1905
rect 3020 1885 3040 1905
rect 3040 1885 3045 1905
rect 3015 1880 3045 1885
rect 3165 1905 3195 1910
rect 3165 1885 3170 1905
rect 3170 1885 3190 1905
rect 3190 1885 3195 1905
rect 3165 1880 3195 1885
rect 3265 1905 3295 1910
rect 3265 1885 3270 1905
rect 3270 1885 3290 1905
rect 3290 1885 3295 1905
rect 3265 1880 3295 1885
rect 3415 1905 3445 1910
rect 3415 1885 3420 1905
rect 3420 1885 3440 1905
rect 3440 1885 3445 1905
rect 3415 1880 3445 1885
rect 3765 1905 3795 1910
rect 3765 1885 3770 1905
rect 3770 1885 3790 1905
rect 3790 1885 3795 1905
rect 3765 1880 3795 1885
rect 3215 1850 3245 1855
rect 3215 1830 3220 1850
rect 3220 1830 3240 1850
rect 3240 1830 3245 1850
rect 3215 1825 3245 1830
rect 2815 1790 2845 1795
rect 2815 1770 2820 1790
rect 2820 1770 2840 1790
rect 2840 1770 2845 1790
rect 2815 1765 2845 1770
rect 3215 1790 3245 1795
rect 3215 1770 3220 1790
rect 3220 1770 3240 1790
rect 3240 1770 3245 1790
rect 3215 1765 3245 1770
rect 3815 1850 3845 1855
rect 3815 1830 3820 1850
rect 3820 1830 3840 1850
rect 3840 1830 3845 1850
rect 3815 1825 3845 1830
rect 3615 1790 3645 1795
rect 3615 1770 3620 1790
rect 3620 1770 3640 1790
rect 3640 1770 3645 1790
rect 3615 1765 3645 1770
rect 3015 1745 3045 1750
rect 3015 1725 3020 1745
rect 3020 1725 3040 1745
rect 3040 1725 3045 1745
rect 3015 1720 3045 1725
rect 3415 1745 3445 1750
rect 3415 1725 3420 1745
rect 3420 1725 3440 1745
rect 3440 1725 3445 1745
rect 3415 1720 3445 1725
rect 2865 1700 2895 1705
rect 2865 1680 2870 1700
rect 2870 1680 2890 1700
rect 2890 1680 2895 1700
rect 2865 1675 2895 1680
rect 3165 1700 3195 1705
rect 3165 1680 3170 1700
rect 3170 1680 3190 1700
rect 3190 1680 3195 1700
rect 3165 1675 3195 1680
rect 3265 1700 3295 1705
rect 3265 1680 3270 1700
rect 3270 1680 3290 1700
rect 3290 1680 3295 1700
rect 3265 1675 3295 1680
rect 3565 1700 3595 1705
rect 3565 1680 3570 1700
rect 3570 1680 3590 1700
rect 3590 1680 3595 1700
rect 3565 1675 3595 1680
rect 2680 1620 2710 1625
rect 2680 1600 2685 1620
rect 2685 1600 2705 1620
rect 2705 1600 2710 1620
rect 2680 1595 2710 1600
rect 840 1505 870 1535
rect 655 820 685 825
rect 655 800 660 820
rect 660 800 680 820
rect 680 800 685 820
rect 655 795 685 800
rect 950 1530 980 1535
rect 950 1510 955 1530
rect 955 1510 975 1530
rect 975 1510 980 1530
rect 950 1505 980 1510
rect 1900 1530 2110 1535
rect 1900 1510 1905 1530
rect 1905 1510 1925 1530
rect 1925 1510 1950 1530
rect 1950 1510 1970 1530
rect 1970 1510 1995 1530
rect 1995 1510 2015 1530
rect 2015 1510 2040 1530
rect 2040 1510 2060 1530
rect 2060 1510 2085 1530
rect 2085 1510 2105 1530
rect 2105 1510 2110 1530
rect 1900 1505 2110 1510
rect 2300 1510 2330 1540
rect 3015 1535 3045 1540
rect 3015 1515 3020 1535
rect 3020 1515 3040 1535
rect 3040 1515 3045 1535
rect 3015 1510 3045 1515
rect 3415 1535 3445 1540
rect 3415 1515 3420 1535
rect 3420 1515 3440 1535
rect 3440 1515 3445 1535
rect 3415 1510 3445 1515
rect 3665 1540 3695 1545
rect 3665 1520 3670 1540
rect 3670 1520 3690 1540
rect 3690 1520 3695 1540
rect 3665 1515 3695 1520
rect 2915 1490 2945 1495
rect 2915 1470 2920 1490
rect 2920 1470 2940 1490
rect 2940 1470 2945 1490
rect 2915 1465 2945 1470
rect 3115 1490 3145 1495
rect 3115 1470 3120 1490
rect 3120 1470 3140 1490
rect 3140 1470 3145 1490
rect 3115 1465 3145 1470
rect 3315 1490 3345 1495
rect 3315 1470 3320 1490
rect 3320 1470 3340 1490
rect 3340 1470 3345 1490
rect 3315 1465 3345 1470
rect 3515 1490 3545 1495
rect 3515 1470 3520 1490
rect 3520 1470 3540 1490
rect 3540 1470 3545 1490
rect 3515 1465 3545 1470
rect 4435 1700 4465 1705
rect 4435 1680 4440 1700
rect 4440 1680 4460 1700
rect 4460 1680 4465 1700
rect 4435 1675 4465 1680
rect 3695 1430 3725 1435
rect 3695 1410 3700 1430
rect 3700 1410 3720 1430
rect 3720 1410 3725 1430
rect 3695 1405 3725 1410
rect 3815 1405 3845 1435
rect 950 1235 980 1240
rect 950 1215 955 1235
rect 955 1215 975 1235
rect 975 1215 980 1235
rect 950 1210 980 1215
rect 3175 960 3205 965
rect 3175 940 3180 960
rect 3180 940 3200 960
rect 3200 940 3205 960
rect 3175 935 3205 940
rect 3215 960 3245 965
rect 3215 940 3220 960
rect 3220 940 3240 960
rect 3240 940 3245 960
rect 3215 935 3245 940
rect 3255 960 3285 965
rect 3255 940 3260 960
rect 3260 940 3280 960
rect 3280 940 3285 960
rect 3255 935 3285 940
rect 3725 900 3755 905
rect 3725 880 3730 900
rect 3730 880 3750 900
rect 3750 880 3755 900
rect 3725 875 3755 880
rect 4500 875 4530 905
rect 3800 815 3830 820
rect 3800 795 3805 815
rect 3805 795 3825 815
rect 3825 795 3830 815
rect 3800 790 3830 795
<< metal2 >>
rect -130 2975 -90 2980
rect -130 2945 -125 2975
rect -95 2945 -90 2975
rect -130 2940 -90 2945
rect 4830 2975 4870 2980
rect 4830 2945 4835 2975
rect 4865 2945 4870 2975
rect 4830 2940 4870 2945
rect -130 2850 -90 2855
rect -130 2820 -125 2850
rect -95 2845 -90 2850
rect 2510 2850 2550 2855
rect 2510 2845 2515 2850
rect -95 2825 2515 2845
rect -95 2820 -90 2825
rect -130 2815 -90 2820
rect 2510 2820 2515 2825
rect 2545 2845 2550 2850
rect 2710 2850 2750 2855
rect 2710 2845 2715 2850
rect 2545 2825 2715 2845
rect 2545 2820 2550 2825
rect 2510 2815 2550 2820
rect 2710 2820 2715 2825
rect 2745 2845 2750 2850
rect 2910 2850 2950 2855
rect 2910 2845 2915 2850
rect 2745 2825 2915 2845
rect 2745 2820 2750 2825
rect 2710 2815 2750 2820
rect 2910 2820 2915 2825
rect 2945 2845 2950 2850
rect 3110 2850 3150 2855
rect 3110 2845 3115 2850
rect 2945 2825 3115 2845
rect 2945 2820 2950 2825
rect 2910 2815 2950 2820
rect 3110 2820 3115 2825
rect 3145 2845 3150 2850
rect 3310 2850 3350 2855
rect 3310 2845 3315 2850
rect 3145 2825 3210 2845
rect 3250 2825 3315 2845
rect 3145 2820 3150 2825
rect 3110 2815 3150 2820
rect 3310 2820 3315 2825
rect 3345 2845 3350 2850
rect 3510 2850 3550 2855
rect 3510 2845 3515 2850
rect 3345 2825 3515 2845
rect 3345 2820 3350 2825
rect 3310 2815 3350 2820
rect 3510 2820 3515 2825
rect 3545 2845 3550 2850
rect 3710 2850 3750 2855
rect 3710 2845 3715 2850
rect 3545 2825 3715 2845
rect 3545 2820 3550 2825
rect 3510 2815 3550 2820
rect 3710 2820 3715 2825
rect 3745 2845 3750 2850
rect 3910 2850 3950 2855
rect 3910 2845 3915 2850
rect 3745 2825 3915 2845
rect 3745 2820 3750 2825
rect 3710 2815 3750 2820
rect 3910 2820 3915 2825
rect 3945 2845 3950 2850
rect 4830 2850 4870 2855
rect 4830 2845 4835 2850
rect 3945 2825 4835 2845
rect 3945 2820 3950 2825
rect 3910 2815 3950 2820
rect 4830 2820 4835 2825
rect 4865 2820 4870 2850
rect 4830 2815 4870 2820
rect -55 2590 985 2595
rect -55 2560 -50 2590
rect -20 2560 950 2590
rect 980 2560 985 2590
rect -55 2555 985 2560
rect 2150 2380 2190 2385
rect 2150 2350 2155 2380
rect 2185 2375 2190 2380
rect 3010 2380 3050 2385
rect 3010 2375 3015 2380
rect 2185 2355 3015 2375
rect 2185 2350 2190 2355
rect 2150 2345 2190 2350
rect 3010 2350 3015 2355
rect 3045 2375 3050 2380
rect 3410 2380 3450 2385
rect 3410 2375 3415 2380
rect 3045 2355 3415 2375
rect 3045 2350 3050 2355
rect 3010 2345 3050 2350
rect 3410 2350 3415 2355
rect 3445 2350 3450 2380
rect 3410 2345 3450 2350
rect 3760 2380 3800 2385
rect 3760 2350 3765 2380
rect 3795 2375 3800 2380
rect 4375 2380 4415 2385
rect 4375 2375 4380 2380
rect 3795 2355 4380 2375
rect 3795 2350 3800 2355
rect 3760 2345 3800 2350
rect 4375 2350 4380 2355
rect 4410 2350 4415 2380
rect 4375 2345 4415 2350
rect 2295 2335 2335 2340
rect 2295 2305 2300 2335
rect 2330 2330 2335 2335
rect 2820 2335 2860 2340
rect 2820 2330 2825 2335
rect 2330 2310 2825 2330
rect 2330 2305 2335 2310
rect 2295 2300 2335 2305
rect 2820 2305 2825 2310
rect 2855 2330 2860 2335
rect 3600 2335 3640 2340
rect 3600 2330 3605 2335
rect 2855 2310 3605 2330
rect 2855 2305 2860 2310
rect 2820 2300 2860 2305
rect 3600 2305 3605 2310
rect 3635 2305 3640 2335
rect 3600 2300 3640 2305
rect 1895 2295 2115 2300
rect 1895 2265 1900 2295
rect 2110 2285 2115 2295
rect 2610 2290 2650 2295
rect 2610 2285 2615 2290
rect 2110 2265 2615 2285
rect 1895 2260 2115 2265
rect 2610 2260 2615 2265
rect 2645 2285 2650 2290
rect 3210 2290 3250 2295
rect 3210 2285 3215 2290
rect 2645 2265 3215 2285
rect 2645 2260 2650 2265
rect 2610 2255 2650 2260
rect 3210 2260 3215 2265
rect 3245 2285 3250 2290
rect 3810 2290 3850 2295
rect 3810 2285 3815 2290
rect 3245 2265 3815 2285
rect 3245 2260 3250 2265
rect 3210 2255 3250 2260
rect 3810 2260 3815 2265
rect 3845 2260 3850 2290
rect 3810 2255 3850 2260
rect -130 2230 -90 2235
rect -130 2200 -125 2230
rect -95 2225 -90 2230
rect 2510 2230 2550 2235
rect 2510 2225 2515 2230
rect -95 2205 2515 2225
rect -95 2200 -90 2205
rect -130 2195 -90 2200
rect 2510 2200 2515 2205
rect 2545 2225 2550 2230
rect 2710 2230 2750 2235
rect 2710 2225 2715 2230
rect 2545 2205 2715 2225
rect 2545 2200 2550 2205
rect 2510 2195 2550 2200
rect 2710 2200 2715 2205
rect 2745 2225 2750 2230
rect 2910 2230 2950 2235
rect 2910 2225 2915 2230
rect 2745 2205 2915 2225
rect 2745 2200 2750 2205
rect 2710 2195 2750 2200
rect 2910 2200 2915 2205
rect 2945 2225 2950 2230
rect 3110 2230 3150 2235
rect 3110 2225 3115 2230
rect 2945 2205 3115 2225
rect 2945 2200 2950 2205
rect 2910 2195 2950 2200
rect 3110 2200 3115 2205
rect 3145 2225 3150 2230
rect 3310 2230 3350 2235
rect 3310 2225 3315 2230
rect 3145 2205 3315 2225
rect 3145 2200 3150 2205
rect 3110 2195 3150 2200
rect 3310 2200 3315 2205
rect 3345 2225 3350 2230
rect 3510 2230 3550 2235
rect 3510 2225 3515 2230
rect 3345 2205 3515 2225
rect 3345 2200 3350 2205
rect 3310 2195 3350 2200
rect 3510 2200 3515 2205
rect 3545 2225 3550 2230
rect 3710 2230 3750 2235
rect 3710 2225 3715 2230
rect 3545 2205 3715 2225
rect 3545 2200 3550 2205
rect 3510 2195 3550 2200
rect 3710 2200 3715 2205
rect 3745 2225 3750 2230
rect 3910 2230 3950 2235
rect 3910 2225 3915 2230
rect 3745 2205 3915 2225
rect 3745 2200 3750 2205
rect 3710 2195 3750 2200
rect 3910 2200 3915 2205
rect 3945 2200 3950 2230
rect 3910 2195 3950 2200
rect 4585 2230 4625 2235
rect 4585 2200 4590 2230
rect 4620 2225 4625 2230
rect 4830 2230 4870 2235
rect 4830 2225 4835 2230
rect 4620 2205 4835 2225
rect 4620 2200 4625 2205
rect 4585 2195 4625 2200
rect 4830 2200 4835 2205
rect 4865 2200 4870 2230
rect 4830 2195 4870 2200
rect -55 2005 985 2010
rect -55 1975 -50 2005
rect -20 1975 950 2005
rect 980 1975 985 2005
rect -55 1970 985 1975
rect 2810 1955 2850 1960
rect 2810 1925 2815 1955
rect 2845 1950 2850 1955
rect 3610 1955 3650 1960
rect 3610 1950 3615 1955
rect 2845 1930 3615 1950
rect 2845 1925 2850 1930
rect 2810 1920 2850 1925
rect 3610 1925 3615 1930
rect 3645 1925 3650 1955
rect 3610 1920 3650 1925
rect 2660 1910 2700 1915
rect 2660 1880 2665 1910
rect 2695 1905 2700 1910
rect 3010 1910 3050 1915
rect 3010 1905 3015 1910
rect 2695 1885 3015 1905
rect 2695 1880 2700 1885
rect 2660 1875 2700 1880
rect 3010 1880 3015 1885
rect 3045 1905 3050 1910
rect 3160 1910 3200 1915
rect 3160 1905 3165 1910
rect 3045 1885 3165 1905
rect 3045 1880 3050 1885
rect 3010 1875 3050 1880
rect 3160 1880 3165 1885
rect 3195 1905 3200 1910
rect 3260 1910 3300 1915
rect 3260 1905 3265 1910
rect 3195 1885 3265 1905
rect 3195 1880 3200 1885
rect 3160 1875 3200 1880
rect 3260 1880 3265 1885
rect 3295 1905 3300 1910
rect 3410 1910 3450 1915
rect 3410 1905 3415 1910
rect 3295 1885 3415 1905
rect 3295 1880 3300 1885
rect 3260 1875 3300 1880
rect 3410 1880 3415 1885
rect 3445 1905 3450 1910
rect 3760 1910 3800 1915
rect 3760 1905 3765 1910
rect 3445 1885 3765 1905
rect 3445 1880 3450 1885
rect 3410 1875 3450 1880
rect 3760 1880 3765 1885
rect 3795 1880 3800 1910
rect 3760 1875 3800 1880
rect 2610 1855 2650 1860
rect 2610 1825 2615 1855
rect 2645 1850 2650 1855
rect 3210 1855 3250 1860
rect 3210 1850 3215 1855
rect 2645 1830 3215 1850
rect 2645 1825 2650 1830
rect 2610 1820 2650 1825
rect 3210 1825 3215 1830
rect 3245 1850 3250 1855
rect 3810 1855 3850 1860
rect 3810 1850 3815 1855
rect 3245 1830 3815 1850
rect 3245 1825 3250 1830
rect 3210 1820 3250 1825
rect 3810 1825 3815 1830
rect 3845 1825 3850 1855
rect 3810 1820 3850 1825
rect 2810 1795 2850 1800
rect 2810 1765 2815 1795
rect 2845 1790 2850 1795
rect 3210 1795 3250 1800
rect 3210 1790 3215 1795
rect 2845 1770 3215 1790
rect 2845 1765 2850 1770
rect 2810 1760 2850 1765
rect 3210 1765 3215 1770
rect 3245 1790 3250 1795
rect 3610 1795 3650 1800
rect 3610 1790 3615 1795
rect 3245 1770 3615 1790
rect 3245 1765 3250 1770
rect 3210 1760 3250 1765
rect 3610 1765 3615 1770
rect 3645 1765 3650 1795
rect 3610 1760 3650 1765
rect 3010 1750 3050 1755
rect 3010 1720 3015 1750
rect 3045 1745 3050 1750
rect 3410 1750 3450 1755
rect 3410 1745 3415 1750
rect 3045 1725 3415 1745
rect 3045 1720 3050 1725
rect 3010 1715 3050 1720
rect 3410 1720 3415 1725
rect 3445 1720 3450 1750
rect 3410 1715 3450 1720
rect 465 1710 2115 1715
rect 465 1680 470 1710
rect 500 1680 1900 1710
rect 2110 1700 2115 1710
rect 2150 1705 2190 1710
rect 2150 1700 2155 1705
rect 2110 1680 2155 1700
rect 465 1675 2115 1680
rect 2150 1675 2155 1680
rect 2185 1700 2190 1705
rect 2860 1705 2900 1710
rect 2860 1700 2865 1705
rect 2185 1680 2865 1700
rect 2185 1675 2190 1680
rect 2150 1670 2190 1675
rect 2860 1675 2865 1680
rect 2895 1700 2900 1705
rect 3160 1705 3200 1710
rect 3160 1700 3165 1705
rect 2895 1680 3165 1700
rect 2895 1675 2900 1680
rect 2860 1670 2900 1675
rect 3160 1675 3165 1680
rect 3195 1700 3200 1705
rect 3260 1705 3300 1710
rect 3260 1700 3265 1705
rect 3195 1680 3265 1700
rect 3195 1675 3200 1680
rect 3160 1670 3200 1675
rect 3260 1675 3265 1680
rect 3295 1700 3300 1705
rect 3560 1705 3600 1710
rect 3560 1700 3565 1705
rect 3295 1680 3565 1700
rect 3295 1675 3300 1680
rect 3260 1670 3300 1675
rect 3560 1675 3565 1680
rect 3595 1700 3600 1705
rect 4430 1705 4470 1710
rect 4430 1700 4435 1705
rect 3595 1680 4435 1700
rect 3595 1675 3600 1680
rect 3560 1670 3600 1675
rect 4430 1675 4435 1680
rect 4465 1675 4470 1705
rect 4430 1670 4470 1675
rect -55 1625 -15 1630
rect -55 1595 -50 1625
rect -20 1620 -15 1625
rect 2675 1625 2715 1630
rect 2675 1620 2680 1625
rect -20 1600 2680 1620
rect -20 1595 -15 1600
rect -55 1590 -15 1595
rect 2675 1595 2680 1600
rect 2710 1595 2715 1625
rect 2675 1590 2715 1595
rect 3660 1545 3700 1550
rect 2295 1540 2335 1545
rect 835 1535 985 1540
rect 835 1505 840 1535
rect 870 1505 950 1535
rect 980 1505 985 1535
rect 835 1500 985 1505
rect 1895 1535 2115 1540
rect 2295 1535 2300 1540
rect 1895 1505 1900 1535
rect 2110 1515 2300 1535
rect 2110 1505 2115 1515
rect 2295 1510 2300 1515
rect 2330 1535 2335 1540
rect 3010 1540 3050 1545
rect 3010 1535 3015 1540
rect 2330 1515 3015 1535
rect 2330 1510 2335 1515
rect 2295 1505 2335 1510
rect 3010 1510 3015 1515
rect 3045 1535 3050 1540
rect 3410 1540 3450 1545
rect 3410 1535 3415 1540
rect 3045 1515 3415 1535
rect 3045 1510 3050 1515
rect 3010 1505 3050 1510
rect 3410 1510 3415 1515
rect 3445 1510 3450 1540
rect 3660 1515 3665 1545
rect 3695 1540 3700 1545
rect 4755 1545 4795 1550
rect 4755 1540 4760 1545
rect 3695 1520 4760 1540
rect 3695 1515 3700 1520
rect 3660 1510 3700 1515
rect 4755 1515 4760 1520
rect 4790 1515 4795 1545
rect 4755 1510 4795 1515
rect 3410 1505 3450 1510
rect 1895 1500 2115 1505
rect 2910 1495 2950 1500
rect 2910 1465 2915 1495
rect 2945 1490 2950 1495
rect 3110 1495 3150 1500
rect 3110 1490 3115 1495
rect 2945 1470 3115 1490
rect 2945 1465 2950 1470
rect 2910 1460 2950 1465
rect 3110 1465 3115 1470
rect 3145 1490 3150 1495
rect 3310 1495 3350 1500
rect 3310 1490 3315 1495
rect 3145 1470 3315 1490
rect 3145 1465 3150 1470
rect 3110 1460 3150 1465
rect 3310 1465 3315 1470
rect 3345 1490 3350 1495
rect 3510 1495 3550 1500
rect 3510 1490 3515 1495
rect 3345 1470 3515 1490
rect 3345 1465 3350 1470
rect 3310 1460 3350 1465
rect 3510 1465 3515 1470
rect 3545 1465 3550 1495
rect 3510 1460 3550 1465
rect 3690 1435 3730 1440
rect 3690 1405 3695 1435
rect 3725 1430 3730 1435
rect 3810 1435 3850 1440
rect 3810 1430 3815 1435
rect 3725 1410 3815 1430
rect 3725 1405 3730 1410
rect 3690 1400 3730 1405
rect 3810 1405 3815 1410
rect 3845 1405 3850 1435
rect 3810 1400 3850 1405
rect -55 1240 985 1245
rect -55 1210 -50 1240
rect -20 1210 950 1240
rect 980 1210 985 1240
rect -55 1205 985 1210
rect -55 965 -15 970
rect -55 935 -50 965
rect -20 960 -15 965
rect 3170 965 3290 970
rect 3170 960 3175 965
rect -20 940 3175 960
rect -20 935 -15 940
rect -55 930 -15 935
rect 3170 935 3175 940
rect 3205 935 3215 965
rect 3245 935 3255 965
rect 3285 960 3290 965
rect 4755 965 4795 970
rect 4755 960 4760 965
rect 3285 940 4760 960
rect 3285 935 3290 940
rect 3170 930 3290 935
rect 4755 935 4760 940
rect 4790 935 4795 965
rect 4755 930 4795 935
rect 3720 905 3760 910
rect 3720 875 3725 905
rect 3755 900 3760 905
rect 4495 905 4535 910
rect 4495 900 4500 905
rect 3755 880 4500 900
rect 3755 875 3760 880
rect 3720 870 3760 875
rect 4495 875 4500 880
rect 4530 875 4535 905
rect 4495 870 4535 875
rect -55 825 -15 830
rect -55 795 -50 825
rect -20 820 -15 825
rect 650 825 690 830
rect 650 820 655 825
rect -20 800 655 820
rect -20 795 -15 800
rect -55 790 -15 795
rect 650 795 655 800
rect 685 795 690 825
rect 650 790 690 795
rect 3795 820 3835 825
rect 3795 790 3800 820
rect 3830 815 3835 820
rect 4755 820 4795 825
rect 4755 815 4760 820
rect 3830 795 4760 815
rect 3830 790 3835 795
rect 3795 785 3835 790
rect 4755 790 4760 795
rect 4790 790 4795 820
rect 4755 785 4795 790
rect -130 -90 -90 -85
rect -130 -120 -125 -90
rect -95 -120 -90 -90
rect -130 -125 -90 -120
<< via2 >>
rect -125 2945 -95 2975
rect 4835 2945 4865 2975
rect -125 2820 -95 2850
rect 4835 2820 4865 2850
rect -50 2560 -20 2590
rect -125 2200 -95 2230
rect 4835 2200 4865 2230
rect -50 1975 -20 2005
rect -50 1595 -20 1625
rect 4760 1515 4790 1545
rect -50 1210 -20 1240
rect -50 935 -20 965
rect 4760 935 4790 965
rect -50 795 -20 825
rect 4760 790 4790 820
rect -125 -120 -95 -90
<< metal3 >>
rect -135 2980 -85 2985
rect -135 2940 -130 2980
rect -90 2940 -85 2980
rect -135 2935 -85 2940
rect 4825 2980 4875 2985
rect 4825 2940 4830 2980
rect 4870 2940 4875 2980
rect 4825 2935 4875 2940
rect -130 2850 -90 2935
rect -60 2905 -10 2910
rect -60 2865 -55 2905
rect -15 2865 -10 2905
rect -60 2860 -10 2865
rect 4750 2905 4800 2910
rect 4750 2865 4755 2905
rect 4795 2865 4800 2905
rect 4750 2860 4800 2865
rect -130 2820 -125 2850
rect -95 2820 -90 2850
rect -130 2230 -90 2820
rect -130 2200 -125 2230
rect -95 2200 -90 2230
rect -130 -80 -90 2200
rect -55 2590 -15 2860
rect -55 2560 -50 2590
rect -20 2560 -15 2590
rect -55 2005 -15 2560
rect -55 1975 -50 2005
rect -20 1975 -15 2005
rect -55 1625 -15 1975
rect -55 1595 -50 1625
rect -20 1595 -15 1625
rect -55 1240 -15 1595
rect -55 1210 -50 1240
rect -20 1210 -15 1240
rect -55 965 -15 1210
rect -55 935 -50 965
rect -20 935 -15 965
rect -55 825 -15 935
rect -55 795 -50 825
rect -20 795 -15 825
rect -55 -5 -15 795
rect 4755 1545 4795 2860
rect 4755 1515 4760 1545
rect 4790 1515 4795 1545
rect 4755 965 4795 1515
rect 4755 935 4760 965
rect 4790 935 4795 965
rect 4755 820 4795 935
rect 4755 790 4760 820
rect 4790 790 4795 820
rect 4755 -5 4795 790
rect 4830 2850 4870 2935
rect 4830 2820 4835 2850
rect 4865 2820 4870 2850
rect 4830 2230 4870 2820
rect 4830 2200 4835 2230
rect 4865 2200 4870 2230
rect -60 -10 -10 -5
rect -60 -50 -55 -10
rect -15 -50 -10 -10
rect -60 -55 -10 -50
rect 4750 -10 4800 -5
rect 4750 -50 4755 -10
rect 4795 -50 4800 -10
rect 4750 -55 4800 -50
rect 4830 -80 4870 2200
rect -135 -85 -85 -80
rect -135 -125 -130 -85
rect -90 -125 -85 -85
rect -135 -130 -85 -125
rect 4825 -85 4875 -80
rect 4825 -125 4830 -85
rect 4870 -125 4875 -85
rect 4825 -130 4875 -125
<< via3 >>
rect -130 2975 -90 2980
rect -130 2945 -125 2975
rect -125 2945 -95 2975
rect -95 2945 -90 2975
rect -130 2940 -90 2945
rect 4830 2975 4870 2980
rect 4830 2945 4835 2975
rect 4835 2945 4865 2975
rect 4865 2945 4870 2975
rect 4830 2940 4870 2945
rect -55 2865 -15 2905
rect 4755 2865 4795 2905
rect -55 -50 -15 -10
rect 4755 -50 4795 -10
rect -130 -90 -90 -85
rect -130 -120 -125 -90
rect -125 -120 -95 -90
rect -95 -120 -90 -90
rect -130 -125 -90 -120
rect 4830 -125 4870 -85
<< metal4 >>
rect -135 2980 -85 2985
rect 4825 2980 4875 2985
rect -135 2940 -130 2980
rect -90 2940 4830 2980
rect 4870 2940 4875 2980
rect -135 2935 -85 2940
rect 4825 2935 4875 2940
rect -60 2905 -10 2910
rect 4750 2905 4800 2910
rect -60 2865 -55 2905
rect -15 2865 4755 2905
rect 4795 2865 4800 2905
rect -60 2860 -10 2865
rect 4750 2860 4800 2865
rect -60 -10 -10 -5
rect 4750 -10 4800 -5
rect -60 -50 -55 -10
rect -15 -50 4755 -10
rect 4795 -50 4800 -10
rect -60 -55 -10 -50
rect 4750 -55 4800 -50
rect -135 -85 -85 -80
rect 4825 -85 4875 -80
rect -135 -125 -130 -85
rect -90 -125 4830 -85
rect 4870 -125 4875 -85
rect -135 -130 -85 -125
rect 4825 -130 4875 -125
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1723858470
transform 1 0 675 0 1 0
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1723858470
transform 1 0 -5 0 1 0
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
timestamp 1723858470
transform 1 0 1355 0 1 0
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1723858470
transform 1 0 2035 0 1 0
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1723858470
transform 1 0 2715 0 1 0
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5
timestamp 1723858470
transform 1 0 3395 0 1 0
box 0 0 670 670
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6
timestamp 1723858470
transform 1 0 4075 0 1 0
box 0 0 670 670
<< labels >>
flabel metal3 4870 1400 4870 1400 3 FreeSans 800 0 80 0 VDDA
port 1 e
flabel metal3 4795 1175 4795 1175 3 FreeSans 800 0 80 0 GNDA
port 6 e
flabel metal1 4525 1615 4525 1615 3 FreeSans 400 0 80 0 start_up
flabel metal2 2285 1515 2285 1515 5 FreeSans 400 0 0 -80 Vin+
flabel metal1 875 1040 875 1040 3 FreeSans 400 0 80 0 Vbe2
flabel metal1 3230 3165 3230 3165 1 FreeSans 800 0 0 400 V_out
port 5 n
flabel locali 2920 1450 2920 1450 7 FreeSans 400 0 -80 0 V_p
flabel metal2 2285 1680 2285 1680 5 FreeSans 400 0 0 -80 Vin-
flabel metal1 4415 2365 4415 2365 3 FreeSans 400 0 80 0 V_TOP
<< end >>
