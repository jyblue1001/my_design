* PEX produced on Mon Feb 17 04:12:37 PM CET 2025 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from loop_filter_2.ext - technology: sky130A

.subckt loop_filter_magic V_OUT GNDA
X0 GNDA.t1 V_OUT.t1 sky130_fd_pr__cap_mim_m3_1 l=60 w=13.8
X1 GNDA.t2 R1_C1.t1 sky130_fd_pr__cap_mim_m3_1 l=60 w=69.8
X2 V_OUT.t0 R1_C1.t0 GNDA.t0 sky130_fd_pr__res_xhigh_po_0p35 l=7.52
R0 GNDA GNDA.t0 3597.15
R1 GNDA GNDA.t1 84.2543
R2 GNDA GNDA.t2 81.0543
R3 V_OUT V_OUT.t0 162.983
R4 V_OUT.n1 V_OUT.t1 8.3085
R5 V_OUT V_OUT.n1 1.07193
R6 V_OUT.n1 V_OUT.n0 0.7505
R7 R1_C1.t0 R1_C1.t1 167.429
C0 V_OUT GNDA 19.821081f
C1 R1_C1.t1 GNDA 2.39887f
C2 V_OUT.t1 GNDA 2.34592f
C3 V_OUT.n1 GNDA 0.011043f
.ends

