magic
tech sky130A
timestamp 1738049277
<< nwell >>
rect 945 100 2035 655
<< nmos >>
rect 1045 -125 1060 -75
rect 1110 -125 1125 -75
rect 1175 -125 1190 -75
rect 1240 -125 1255 -75
rect 1405 -125 1420 -75
rect 1470 -125 1485 -75
rect 1535 -125 1550 -75
rect 1600 -125 1615 -75
rect 1755 -125 1770 -75
rect 1820 -125 1835 -75
rect 1885 -125 1900 -75
rect 1950 -125 1965 -75
rect 1615 -520 1665 -270
rect 1715 -520 1765 -270
rect 1815 -520 1865 -270
rect 1915 -520 1965 -270
<< pmos >>
rect 1095 330 1145 580
rect 1195 330 1245 580
rect 1295 330 1345 580
rect 1395 330 1445 580
rect 1495 330 1545 580
rect 1595 330 1645 580
rect 1695 330 1745 580
rect 1795 330 1845 580
rect 1045 125 1060 225
rect 1110 125 1125 225
rect 1175 125 1190 225
rect 1240 125 1255 225
rect 1405 125 1420 225
rect 1470 125 1485 225
rect 1535 125 1550 225
rect 1600 125 1615 225
rect 1755 125 1770 225
rect 1820 125 1835 225
rect 1885 125 1900 225
rect 1950 125 1965 225
<< ndiff >>
rect 995 -90 1045 -75
rect 995 -110 1010 -90
rect 1030 -110 1045 -90
rect 995 -125 1045 -110
rect 1060 -90 1110 -75
rect 1060 -110 1075 -90
rect 1095 -110 1110 -90
rect 1060 -125 1110 -110
rect 1125 -90 1175 -75
rect 1125 -110 1140 -90
rect 1160 -110 1175 -90
rect 1125 -125 1175 -110
rect 1190 -90 1240 -75
rect 1190 -110 1205 -90
rect 1225 -110 1240 -90
rect 1190 -125 1240 -110
rect 1255 -90 1305 -75
rect 1255 -110 1270 -90
rect 1290 -110 1305 -90
rect 1255 -125 1305 -110
rect 1355 -90 1405 -75
rect 1355 -110 1370 -90
rect 1390 -110 1405 -90
rect 1355 -125 1405 -110
rect 1420 -90 1470 -75
rect 1420 -110 1435 -90
rect 1455 -110 1470 -90
rect 1420 -125 1470 -110
rect 1485 -90 1535 -75
rect 1485 -110 1500 -90
rect 1520 -110 1535 -90
rect 1485 -125 1535 -110
rect 1550 -90 1600 -75
rect 1550 -110 1565 -90
rect 1585 -110 1600 -90
rect 1550 -125 1600 -110
rect 1615 -90 1665 -75
rect 1615 -110 1630 -90
rect 1650 -110 1665 -90
rect 1615 -125 1665 -110
rect 1705 -90 1755 -75
rect 1705 -110 1720 -90
rect 1740 -110 1755 -90
rect 1705 -125 1755 -110
rect 1770 -90 1820 -75
rect 1770 -110 1785 -90
rect 1805 -110 1820 -90
rect 1770 -125 1820 -110
rect 1835 -90 1885 -75
rect 1835 -110 1850 -90
rect 1870 -110 1885 -90
rect 1835 -125 1885 -110
rect 1900 -90 1950 -75
rect 1900 -110 1915 -90
rect 1935 -110 1950 -90
rect 1900 -125 1950 -110
rect 1965 -90 2015 -75
rect 1965 -110 1980 -90
rect 2000 -110 2015 -90
rect 1965 -125 2015 -110
rect 1565 -285 1615 -270
rect 1565 -505 1580 -285
rect 1600 -505 1615 -285
rect 1565 -520 1615 -505
rect 1665 -285 1715 -270
rect 1665 -505 1680 -285
rect 1700 -505 1715 -285
rect 1665 -520 1715 -505
rect 1765 -285 1815 -270
rect 1765 -505 1780 -285
rect 1800 -505 1815 -285
rect 1765 -520 1815 -505
rect 1865 -285 1915 -270
rect 1865 -505 1880 -285
rect 1900 -505 1915 -285
rect 1865 -520 1915 -505
rect 1965 -285 2015 -270
rect 1965 -505 1980 -285
rect 2000 -505 2015 -285
rect 1965 -520 2015 -505
<< pdiff >>
rect 1045 565 1095 580
rect 1045 345 1060 565
rect 1080 345 1095 565
rect 1045 330 1095 345
rect 1145 565 1195 580
rect 1145 345 1160 565
rect 1180 345 1195 565
rect 1145 330 1195 345
rect 1245 565 1295 580
rect 1245 345 1260 565
rect 1280 345 1295 565
rect 1245 330 1295 345
rect 1345 565 1395 580
rect 1345 345 1360 565
rect 1380 345 1395 565
rect 1345 330 1395 345
rect 1445 565 1495 580
rect 1445 345 1460 565
rect 1480 345 1495 565
rect 1445 330 1495 345
rect 1545 565 1595 580
rect 1545 345 1560 565
rect 1580 345 1595 565
rect 1545 330 1595 345
rect 1645 565 1695 580
rect 1645 345 1660 565
rect 1680 345 1695 565
rect 1645 330 1695 345
rect 1745 565 1795 580
rect 1745 345 1760 565
rect 1780 345 1795 565
rect 1745 330 1795 345
rect 1845 565 1895 580
rect 1845 345 1860 565
rect 1880 345 1895 565
rect 1845 330 1895 345
rect 995 210 1045 225
rect 995 140 1010 210
rect 1030 140 1045 210
rect 995 125 1045 140
rect 1060 210 1110 225
rect 1060 140 1075 210
rect 1095 140 1110 210
rect 1060 125 1110 140
rect 1125 210 1175 225
rect 1125 140 1140 210
rect 1160 140 1175 210
rect 1125 125 1175 140
rect 1190 210 1240 225
rect 1190 140 1205 210
rect 1225 140 1240 210
rect 1190 125 1240 140
rect 1255 210 1305 225
rect 1255 140 1270 210
rect 1290 140 1305 210
rect 1255 125 1305 140
rect 1355 210 1405 225
rect 1355 140 1370 210
rect 1390 140 1405 210
rect 1355 125 1405 140
rect 1420 210 1470 225
rect 1420 140 1435 210
rect 1455 140 1470 210
rect 1420 125 1470 140
rect 1485 210 1535 225
rect 1485 140 1500 210
rect 1520 140 1535 210
rect 1485 125 1535 140
rect 1550 210 1600 225
rect 1550 140 1565 210
rect 1585 140 1600 210
rect 1550 125 1600 140
rect 1615 210 1665 225
rect 1615 140 1630 210
rect 1650 140 1665 210
rect 1615 125 1665 140
rect 1705 210 1755 225
rect 1705 140 1720 210
rect 1740 140 1755 210
rect 1705 125 1755 140
rect 1770 210 1820 225
rect 1770 140 1785 210
rect 1805 140 1820 210
rect 1770 125 1820 140
rect 1835 210 1885 225
rect 1835 140 1850 210
rect 1870 140 1885 210
rect 1835 125 1885 140
rect 1900 210 1950 225
rect 1900 140 1915 210
rect 1935 140 1950 210
rect 1900 125 1950 140
rect 1965 210 2015 225
rect 1965 140 1980 210
rect 2000 140 2015 210
rect 1965 125 2015 140
<< ndiffc >>
rect 1010 -110 1030 -90
rect 1075 -110 1095 -90
rect 1140 -110 1160 -90
rect 1205 -110 1225 -90
rect 1270 -110 1290 -90
rect 1370 -110 1390 -90
rect 1435 -110 1455 -90
rect 1500 -110 1520 -90
rect 1565 -110 1585 -90
rect 1630 -110 1650 -90
rect 1720 -110 1740 -90
rect 1785 -110 1805 -90
rect 1850 -110 1870 -90
rect 1915 -110 1935 -90
rect 1980 -110 2000 -90
rect 1580 -505 1600 -285
rect 1680 -505 1700 -285
rect 1780 -505 1800 -285
rect 1880 -505 1900 -285
rect 1980 -505 2000 -285
<< pdiffc >>
rect 1060 345 1080 565
rect 1160 345 1180 565
rect 1260 345 1280 565
rect 1360 345 1380 565
rect 1460 345 1480 565
rect 1560 345 1580 565
rect 1660 345 1680 565
rect 1760 345 1780 565
rect 1860 345 1880 565
rect 1010 140 1030 210
rect 1075 140 1095 210
rect 1140 140 1160 210
rect 1205 140 1225 210
rect 1270 140 1290 210
rect 1370 140 1390 210
rect 1435 140 1455 210
rect 1500 140 1520 210
rect 1565 140 1585 210
rect 1630 140 1650 210
rect 1720 140 1740 210
rect 1785 140 1805 210
rect 1850 140 1870 210
rect 1915 140 1935 210
rect 1980 140 2000 210
<< poly >>
rect 1245 630 1295 645
rect 1245 610 1260 630
rect 1280 610 1295 630
rect 1245 605 1295 610
rect 1645 630 1695 645
rect 1645 610 1660 630
rect 1680 610 1695 630
rect 1645 605 1695 610
rect 1095 590 1845 605
rect 1095 580 1145 590
rect 1195 580 1245 590
rect 1295 580 1345 590
rect 1395 580 1445 590
rect 1495 580 1545 590
rect 1595 580 1645 590
rect 1695 580 1745 590
rect 1795 580 1845 590
rect 1095 315 1145 330
rect 1195 315 1245 330
rect 1295 315 1345 330
rect 1395 315 1445 330
rect 1495 315 1545 330
rect 1595 315 1645 330
rect 1695 315 1745 330
rect 1795 315 1845 330
rect 755 280 1155 290
rect 755 275 935 280
rect 925 260 935 275
rect 955 275 1155 280
rect 955 260 965 275
rect 925 250 965 260
rect 1140 250 1155 275
rect 1045 225 1060 240
rect 1110 235 1190 250
rect 1110 225 1125 235
rect 1175 225 1190 235
rect 1240 225 1255 240
rect 1405 225 1420 240
rect 1470 225 1485 240
rect 1535 225 1550 240
rect 1600 225 1615 240
rect 1755 225 1770 240
rect 1820 225 1835 240
rect 1885 225 1900 240
rect 1950 225 1965 240
rect 1045 85 1060 125
rect 1110 110 1125 125
rect 1175 110 1190 125
rect 1240 85 1255 125
rect 1405 115 1420 125
rect 1470 115 1485 125
rect 1535 115 1550 125
rect 1600 115 1615 125
rect 1405 100 1615 115
rect 1755 110 1770 125
rect 1820 110 1835 125
rect 1885 110 1900 125
rect 1950 110 1965 125
rect 1925 100 1965 110
rect 825 70 1255 85
rect 1490 80 1500 100
rect 1520 80 1530 100
rect 1490 70 1530 80
rect 1925 80 1935 100
rect 1955 80 1965 100
rect 1925 70 1965 80
rect 825 -205 840 70
rect 1270 35 1965 45
rect 1270 15 1280 35
rect 1300 30 1965 35
rect 1300 15 1310 30
rect 1270 5 1310 15
rect 925 -5 965 5
rect 925 -25 935 -5
rect 955 -20 965 -5
rect 1410 -5 1450 5
rect 1410 -20 1420 -5
rect 955 -25 1420 -20
rect 1440 -20 1450 -5
rect 1440 -25 1615 -20
rect 925 -35 1615 -25
rect 1045 -75 1060 -60
rect 1110 -75 1125 -60
rect 1175 -75 1190 -60
rect 1240 -75 1255 -60
rect 1405 -75 1420 -35
rect 1470 -75 1485 -60
rect 1535 -75 1550 -60
rect 1600 -75 1615 -35
rect 1950 -50 1965 30
rect 1755 -65 1965 -50
rect 1755 -75 1770 -65
rect 1820 -75 1835 -65
rect 1885 -75 1900 -65
rect 1950 -75 1965 -65
rect 1045 -135 1060 -125
rect 1110 -135 1125 -125
rect 1175 -135 1190 -125
rect 1240 -135 1255 -125
rect 1045 -150 1255 -135
rect 1405 -140 1420 -125
rect 1470 -135 1485 -125
rect 1535 -135 1550 -125
rect 1470 -150 1550 -135
rect 1600 -140 1615 -125
rect 1755 -140 1770 -125
rect 1820 -140 1835 -125
rect 1885 -140 1900 -125
rect 1950 -140 1965 -125
rect 1130 -170 1140 -150
rect 1160 -170 1170 -150
rect 1130 -180 1170 -170
rect 1470 -205 1485 -150
rect 760 -220 1485 -205
rect 1615 -270 1665 -255
rect 1715 -270 1765 -255
rect 1815 -270 1865 -255
rect 1915 -270 1965 -255
rect 1615 -530 1665 -520
rect 1715 -530 1765 -520
rect 1815 -530 1865 -520
rect 1915 -530 1965 -520
rect 1615 -545 1965 -530
rect 1615 -550 1780 -545
rect 1770 -565 1780 -550
rect 1800 -550 1965 -545
rect 1800 -565 1810 -550
rect 1770 -575 1810 -565
<< polycont >>
rect 1260 610 1280 630
rect 1660 610 1680 630
rect 935 260 955 280
rect 1500 80 1520 100
rect 1935 80 1955 100
rect 1280 15 1300 35
rect 935 -25 955 -5
rect 1420 -25 1440 -5
rect 1140 -170 1160 -150
rect 1780 -565 1800 -545
<< xpolycontact >>
rect 2070 645 2105 865
rect 2070 310 2105 530
rect 1020 -555 1240 -270
rect 1290 -555 1510 -270
rect 2070 -500 2105 -280
rect 2070 -805 2105 -585
<< xpolyres >>
rect 2070 530 2105 645
rect 1240 -555 1290 -270
rect 2070 -585 2105 -500
<< locali >>
rect 2125 920 2165 930
rect 2085 900 2135 920
rect 2155 900 2165 920
rect 2085 865 2105 900
rect 2125 890 2165 900
rect 1245 630 1295 645
rect 1245 620 1260 630
rect 865 610 1260 620
rect 1280 620 1295 630
rect 1645 630 1695 645
rect 1645 620 1660 630
rect 1280 610 1660 620
rect 1680 610 1695 630
rect 865 595 1695 610
rect 865 -270 885 595
rect 1260 575 1280 595
rect 1660 575 1680 595
rect 1050 565 1090 575
rect 1050 345 1060 565
rect 1080 345 1090 565
rect 1050 335 1090 345
rect 1150 565 1190 575
rect 1150 345 1160 565
rect 1180 345 1190 565
rect 1150 335 1190 345
rect 1250 565 1290 575
rect 1250 345 1260 565
rect 1280 345 1290 565
rect 1250 335 1290 345
rect 1350 565 1390 575
rect 1350 345 1360 565
rect 1380 345 1390 565
rect 1350 335 1390 345
rect 1450 565 1490 575
rect 1450 345 1460 565
rect 1480 345 1490 565
rect 1450 335 1490 345
rect 1550 565 1590 575
rect 1550 345 1560 565
rect 1580 345 1590 565
rect 1550 335 1590 345
rect 1650 565 1690 575
rect 1650 345 1660 565
rect 1680 345 1690 565
rect 1650 335 1690 345
rect 1750 565 1790 575
rect 1750 345 1760 565
rect 1780 345 1790 565
rect 1750 335 1790 345
rect 1850 565 1890 575
rect 1850 345 1860 565
rect 1880 345 1890 565
rect 1850 335 1890 345
rect 1060 315 1080 335
rect 1460 315 1480 335
rect 1860 315 1880 335
rect 1060 295 1880 315
rect 925 280 965 290
rect 925 260 935 280
rect 955 260 965 280
rect 925 250 965 260
rect 945 5 965 250
rect 1075 220 1095 295
rect 1205 220 1225 295
rect 2085 260 2105 310
rect 1720 240 2105 260
rect 1720 220 1740 240
rect 1850 220 1870 240
rect 1980 220 2000 240
rect 1000 210 1040 220
rect 1000 140 1010 210
rect 1030 140 1040 210
rect 1000 130 1040 140
rect 1065 210 1105 220
rect 1065 140 1075 210
rect 1095 140 1105 210
rect 1065 130 1105 140
rect 1130 210 1170 220
rect 1130 140 1140 210
rect 1160 140 1170 210
rect 1130 130 1170 140
rect 1195 210 1235 220
rect 1195 140 1205 210
rect 1225 140 1235 210
rect 1195 130 1235 140
rect 1260 210 1300 220
rect 1260 140 1270 210
rect 1290 140 1300 210
rect 1260 130 1300 140
rect 1360 210 1400 220
rect 1360 140 1370 210
rect 1390 140 1400 210
rect 1360 130 1400 140
rect 1425 210 1465 220
rect 1425 140 1435 210
rect 1455 140 1465 210
rect 1425 130 1465 140
rect 1490 210 1530 220
rect 1490 140 1500 210
rect 1520 140 1530 210
rect 1490 130 1530 140
rect 1555 210 1595 220
rect 1555 140 1565 210
rect 1585 140 1595 210
rect 1555 130 1595 140
rect 1620 210 1660 220
rect 1620 140 1630 210
rect 1650 140 1660 210
rect 1620 130 1660 140
rect 1710 210 1750 220
rect 1710 140 1720 210
rect 1740 140 1750 210
rect 1710 130 1750 140
rect 1775 210 1815 220
rect 1775 140 1785 210
rect 1805 140 1815 210
rect 1775 130 1815 140
rect 1840 210 1880 220
rect 1840 140 1850 210
rect 1870 140 1880 210
rect 1840 130 1880 140
rect 1905 210 1945 220
rect 1905 140 1915 210
rect 1935 140 1945 210
rect 1905 130 1945 140
rect 1970 210 2010 220
rect 1970 140 1980 210
rect 2000 140 2010 210
rect 1970 130 2010 140
rect 2125 155 2165 165
rect 2125 135 2135 155
rect 2155 135 2165 155
rect 925 -5 965 5
rect 925 -25 935 -5
rect 955 -25 965 -5
rect 925 -35 965 -25
rect 1010 -80 1030 130
rect 1140 -80 1160 130
rect 1270 45 1290 130
rect 1270 35 1310 45
rect 1270 15 1280 35
rect 1300 15 1310 35
rect 1270 5 1310 15
rect 1270 -80 1290 5
rect 1370 -80 1390 130
rect 1500 110 1520 130
rect 1630 110 1650 130
rect 2125 125 2165 135
rect 1490 100 1530 110
rect 1490 80 1500 100
rect 1520 80 1530 100
rect 1490 70 1530 80
rect 1630 100 1965 110
rect 1630 90 1935 100
rect 1410 -5 1450 5
rect 1410 -25 1420 -5
rect 1440 -25 1450 -5
rect 1410 -35 1450 -25
rect 1500 -80 1520 70
rect 1630 -80 1650 90
rect 1925 80 1935 90
rect 1955 80 1965 100
rect 1925 70 1965 80
rect 2125 35 2145 125
rect 2125 15 3055 35
rect 2125 -80 2145 15
rect 1000 -90 1040 -80
rect 1000 -110 1010 -90
rect 1030 -110 1040 -90
rect 1000 -120 1040 -110
rect 1065 -90 1105 -80
rect 1065 -110 1075 -90
rect 1095 -110 1105 -90
rect 1065 -120 1105 -110
rect 1130 -90 1170 -80
rect 1130 -110 1140 -90
rect 1160 -110 1170 -90
rect 1130 -120 1170 -110
rect 1195 -90 1235 -80
rect 1195 -110 1205 -90
rect 1225 -110 1235 -90
rect 1195 -120 1235 -110
rect 1260 -90 1300 -80
rect 1260 -110 1270 -90
rect 1290 -110 1300 -90
rect 1260 -120 1300 -110
rect 1360 -90 1400 -80
rect 1360 -110 1370 -90
rect 1390 -110 1400 -90
rect 1360 -120 1400 -110
rect 1425 -90 1465 -80
rect 1425 -110 1435 -90
rect 1455 -110 1465 -90
rect 1425 -120 1465 -110
rect 1490 -90 1530 -80
rect 1490 -110 1500 -90
rect 1520 -110 1530 -90
rect 1490 -120 1530 -110
rect 1555 -90 1595 -80
rect 1555 -110 1565 -90
rect 1585 -110 1595 -90
rect 1555 -120 1595 -110
rect 1620 -90 1660 -80
rect 1620 -110 1630 -90
rect 1650 -110 1660 -90
rect 1620 -120 1660 -110
rect 1710 -90 1750 -80
rect 1710 -110 1720 -90
rect 1740 -110 1750 -90
rect 1710 -120 1750 -110
rect 1775 -90 1815 -80
rect 1775 -110 1785 -90
rect 1805 -110 1815 -90
rect 1775 -120 1815 -110
rect 1840 -90 1880 -80
rect 1840 -110 1850 -90
rect 1870 -110 1880 -90
rect 1840 -120 1880 -110
rect 1905 -90 1945 -80
rect 1905 -110 1915 -90
rect 1935 -110 1945 -90
rect 1905 -120 1945 -110
rect 1970 -90 2010 -80
rect 1970 -110 1980 -90
rect 2000 -110 2010 -90
rect 1970 -120 2010 -110
rect 2125 -90 2165 -80
rect 2125 -110 2135 -90
rect 2155 -110 2165 -90
rect 2125 -120 2165 -110
rect 1140 -140 1160 -120
rect 1435 -140 1455 -120
rect 1565 -140 1585 -120
rect 1720 -140 1740 -120
rect 1850 -140 1870 -120
rect 1980 -140 2000 -120
rect 1130 -150 1170 -140
rect 1130 -170 1140 -150
rect 1160 -170 1170 -150
rect 1435 -160 1700 -140
rect 1720 -160 2105 -140
rect 1130 -180 1170 -170
rect 1680 -235 1700 -160
rect 1580 -255 2000 -235
rect 865 -290 1020 -270
rect 1580 -275 1600 -255
rect 1980 -275 2000 -255
rect 1570 -285 1610 -275
rect 1570 -505 1580 -285
rect 1600 -505 1610 -285
rect 1570 -515 1610 -505
rect 1670 -285 1710 -275
rect 1670 -505 1680 -285
rect 1700 -505 1710 -285
rect 1670 -515 1710 -505
rect 1770 -285 1810 -275
rect 1770 -505 1780 -285
rect 1800 -505 1810 -285
rect 1770 -515 1810 -505
rect 1870 -285 1910 -275
rect 1870 -505 1880 -285
rect 1900 -505 1910 -285
rect 1870 -515 1910 -505
rect 1970 -285 2010 -275
rect 2085 -280 2105 -160
rect 1970 -505 1980 -285
rect 2000 -505 2010 -285
rect 1970 -515 2010 -505
rect 1780 -535 1800 -515
rect 1510 -545 1810 -535
rect 1510 -555 1780 -545
rect 1770 -565 1780 -555
rect 1800 -565 1810 -545
rect 1770 -575 1810 -565
rect 2085 -855 2105 -805
rect 2125 -855 2165 -845
rect 2085 -875 2135 -855
rect 2155 -875 2165 -855
rect 2125 -885 2165 -875
<< viali >>
rect 2135 900 2155 920
rect 1160 345 1180 565
rect 1360 345 1380 565
rect 1560 345 1580 565
rect 1760 345 1780 565
rect 1435 140 1455 210
rect 1565 140 1585 210
rect 1785 140 1805 210
rect 1915 140 1935 210
rect 2135 135 2155 155
rect 1075 -110 1095 -90
rect 1205 -110 1225 -90
rect 1785 -110 1805 -90
rect 1915 -110 1935 -90
rect 2135 -110 2155 -90
rect 1680 -505 1700 -285
rect 1880 -505 1900 -285
rect 2135 -875 2155 -855
<< metal1 >>
rect 2125 920 2165 930
rect 2125 900 2135 920
rect 2155 900 2165 920
rect 2125 890 2165 900
rect 915 565 2055 655
rect 915 345 1160 565
rect 1180 345 1360 565
rect 1380 345 1560 565
rect 1580 345 1760 565
rect 1780 345 2055 565
rect 915 210 2055 345
rect 915 140 1435 210
rect 1455 140 1565 210
rect 1585 140 1785 210
rect 1805 140 1915 210
rect 1935 140 2055 210
rect 915 100 2055 140
rect 2125 155 2165 165
rect 2125 135 2135 155
rect 2155 135 2165 155
rect 2125 125 2165 135
rect 1490 70 1530 100
rect 915 -90 2055 -35
rect 915 -110 1075 -90
rect 1095 -110 1205 -90
rect 1225 -110 1785 -90
rect 1805 -110 1915 -90
rect 1935 -110 2055 -90
rect 915 -285 2055 -110
rect 2125 -90 2165 -80
rect 2125 -110 2135 -90
rect 2155 -110 2165 -90
rect 2125 -120 2165 -110
rect 915 -505 1680 -285
rect 1700 -505 1880 -285
rect 1900 -505 2055 -285
rect 915 -575 2055 -505
rect 2125 -855 2165 -845
rect 2125 -875 2135 -855
rect 2155 -875 2165 -855
rect 2125 -885 2165 -875
<< metal3 >>
rect 2125 890 3010 935
rect 2180 105 3010 890
rect 2180 -845 3010 -60
rect 2125 -890 3010 -845
<< mimcap >>
rect 2195 165 2995 920
rect 2195 130 2205 165
rect 2240 130 2995 165
rect 2195 120 2995 130
rect 2195 -85 2995 -75
rect 2195 -120 2205 -85
rect 2240 -120 2995 -85
rect 2195 -875 2995 -120
<< mimcapcontact >>
rect 2205 130 2240 165
rect 2205 -120 2240 -85
<< metal4 >>
rect 2125 165 2245 170
rect 2125 130 2205 165
rect 2240 130 2245 165
rect 2125 125 2245 130
rect 2125 -85 2245 -80
rect 2125 -120 2205 -85
rect 2240 -120 2245 -85
rect 2125 -125 2245 -120
<< labels >>
flabel poly 760 -210 760 -210 7 FreeSans 400 0 0 0 VIN-
flabel poly 755 280 755 280 7 FreeSans 400 0 0 0 VIN+
flabel locali 3055 20 3055 20 3 FreeSans 400 0 0 0 VOUT
flabel metal1 915 -405 915 -405 7 FreeSans 400 0 0 0 GNDA
flabel metal1 915 465 915 465 7 FreeSans 400 0 0 0 VDDA
<< end >>
